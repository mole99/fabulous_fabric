module top(
    input  wire        clk,
    input  wire [47:0] io_in,
    output wire [47:0] io_out,
    output wire [47:0] io_oeb
);

    wire [31:0] sram_do, sram0_do, sram2_do, sram2_do, sram3_do, sram4_do, sram5_do, sram6_do, sram7_do;

    EF_SRAM_1024x32_wrapper0 sram0 (
        .AD     (io_in[9:0]),
        .BEN    (32'hFFFFFFFF),
        .DI     ({4'd0, io_in[31:0]}),
        .EN     (1'b1),
        .R_WB   (1'b1),
        .DO     (sram0_do)
    );
    
    EF_SRAM_1024x32_wrapper1 sram1 (
        .AD     (io_in[9:0]),
        .BEN    (32'hFFFFFFFF),
        .DI     ({4'd0, io_in[31:0]}),
        .EN     (1'b1),
        .R_WB   (1'b1),
        .DO     (sram1_do)
    );
    
    EF_SRAM_1024x32_wrapper2 sram2 (
        .AD     (io_in[9:0]),
        .BEN    (32'hFFFFFFFF),
        .DI     ({4'd0, io_in[31:0]}),
        .EN     (1'b1),
        .R_WB   (1'b1),
        .DO     (sram2_do)
    );
    
    EF_SRAM_1024x32_wrapper3 sram3 (
        .AD     (io_in[9:0]),
        .BEN    (32'hFFFFFFFF),
        .DI     ({4'd0, io_in[31:0]}),
        .EN     (1'b1),
        .R_WB   (1'b1),
        .DO     (sram3_do)
    );
    
    EF_SRAM_1024x32_wrapper4 sram4 (
        .AD     (io_in[9:0]),
        .BEN    (32'hFFFFFFFF),
        .DI     ({4'd0, io_in[31:0]}),
        .EN     (1'b1),
        .R_WB   (1'b1),
        .DO     (sram4_do)
    );
    
    EF_SRAM_1024x32_wrapper5 sram5 (
        .AD     (io_in[9:0]),
        .BEN    (32'hFFFFFFFF),
        .DI     ({4'd0, io_in[31:0]}),
        .EN     (1'b1),
        .R_WB   (1'b1),
        .DO     (sram5_do)
    );
    
    EF_SRAM_1024x32_wrapper6 sram6 (
        .AD     (io_in[9:0]),
        .BEN    (32'hFFFFFFFF),
        .DI     ({4'd0, io_in[31:0]}),
        .EN     (1'b1),
        .R_WB   (1'b1),
        .DO     (sram6_do)
    );
    
    EF_SRAM_1024x32_wrapper7 sram7 (
        .AD     (io_in[9:0]),
        .BEN    (32'hFFFFFFFF),
        .DI     ({4'd0, io_in[31:0]}),
        .EN     (1'b1),
        .R_WB   (1'b1),
        .DO     (sram7_do)
    );
    
    always_comb begin
        case (io_in[12:10])
            3'd0:  sram_do = sram0_do;
            3'd1:  sram_do = sram1_do;
            3'd2:  sram_do = sram2_do;
            3'd3:  sram_do = sram3_do;
            3'd4:  sram_do = sram4_do;
            3'd5:  sram_do = sram5_do;
            3'd6:  sram_do = sram6_do;
            3'd7:  sram_do = sram7_do;
            default: sram_do = 'x;
        endcase
    end
    
    assign io_out = {16'd0, sram_do};

endmodule

module EF_SRAM_1024x32_wrapper0 (
    input  [ 9:0] AD,
    input  [31:0] BEN,
    input  [31:0] DI,
    input         EN,
    input         R_WB,
    output [31:0] DO
);
    (* keep, BEL="X11Y2.A" *) EF_SRAM_1024x32 i_EF_SRAM_1024x32 (
        .AD0    (AD[0]),
        .AD1    (AD[1]),
        .AD2    (AD[2]),
        .AD3    (AD[3]),
        .AD4    (AD[4]),
        .AD5    (AD[5]),
        .AD6    (AD[6]),
        .AD7    (AD[7]),
        .AD8    (AD[8]),
        .AD9    (AD[9]),
        
        .BEN0   (BEN[0]),
        .BEN1   (BEN[1]),
        .BEN2   (BEN[2]),
        .BEN3   (BEN[3]),
        .BEN4   (BEN[4]),
        .BEN5   (BEN[5]),
        .BEN6   (BEN[6]),
        .BEN7   (BEN[7]),
        .BEN8   (BEN[8]),
        .BEN9   (BEN[9]),
        .BEN10   (BEN[10]),
        .BEN11   (BEN[11]),
        .BEN12   (BEN[12]),
        .BEN13   (BEN[13]),
        .BEN14   (BEN[14]),
        .BEN15   (BEN[15]),
        .BEN16   (BEN[16]),
        .BEN17   (BEN[17]),
        .BEN18   (BEN[18]),
        .BEN19   (BEN[19]),
        .BEN20   (BEN[20]),
        .BEN21   (BEN[21]),
        .BEN22   (BEN[22]),
        .BEN23   (BEN[23]),
        .BEN24   (BEN[24]),
        .BEN25   (BEN[25]),
        .BEN26   (BEN[26]),
        .BEN27   (BEN[27]),
        .BEN28   (BEN[28]),
        .BEN29   (BEN[29]),
        .BEN30   (BEN[30]),
        .BEN31   (BEN[31]),
        
        .DI0    (DI[0]),
        .DI1    (DI[1]),
        .DI2    (DI[2]),
        .DI3    (DI[3]),
        .DI4    (DI[4]),
        .DI5    (DI[5]),
        .DI6    (DI[6]),
        .DI7    (DI[7]),
        .DI8    (DI[8]),
        .DI9    (DI[9]),
        .DI10    (DI[10]),
        .DI11    (DI[11]),
        .DI12    (DI[12]),
        .DI13    (DI[13]),
        .DI14    (DI[14]),
        .DI15    (DI[15]),
        .DI16    (DI[16]),
        .DI17    (DI[17]),
        .DI18    (DI[18]),
        .DI19    (DI[19]),
        .DI20    (DI[20]),
        .DI21    (DI[21]),
        .DI22    (DI[22]),
        .DI23    (DI[23]),
        .DI24    (DI[24]),
        .DI25    (DI[25]),
        .DI26    (DI[26]),
        .DI27    (DI[27]),
        .DI28    (DI[28]),
        .DI29    (DI[29]),
        .DI30    (DI[30]),
        .DI31    (DI[31]),
        
        .EN     (EN),

        .R_WB   (R_WB),
        
        .DO0    (DO[0]),
        .DO1    (DO[1]),
        .DO2    (DO[2]),
        .DO3    (DO[3]),
        .DO4    (DO[4]),
        .DO5    (DO[5]),
        .DO6    (DO[6]),
        .DO7    (DO[7]),
        .DO8    (DO[8]),
        .DO9    (DO[9]),
        .DO10    (DO[10]),
        .DO11    (DO[11]),
        .DO12    (DO[12]),
        .DO13    (DO[13]),
        .DO14    (DO[14]),
        .DO15    (DO[15]),
        .DO16    (DO[16]),
        .DO17    (DO[17]),
        .DO18    (DO[18]),
        .DO19    (DO[19]),
        .DO20    (DO[20]),
        .DO21    (DO[21]),
        .DO22    (DO[22]),
        .DO23    (DO[23]),
        .DO24    (DO[24]),
        .DO25    (DO[25]),
        .DO26    (DO[26]),
        .DO27    (DO[27]),
        .DO28    (DO[28]),
        .DO29    (DO[29]),
        .DO30    (DO[30]),
        .DO31    (DO[31])
    );

endmodule

module EF_SRAM_1024x32_wrapper1 (
    input  [ 9:0] AD,
    input  [31:0] BEN,
    input  [31:0] DI,
    input         EN,
    input         R_WB,
    output [31:0] DO
);
    (* keep, BEL="X11Y4.A" *) EF_SRAM_1024x32 i_EF_SRAM_1024x32 (
        .AD0    (AD[0]),
        .AD1    (AD[1]),
        .AD2    (AD[2]),
        .AD3    (AD[3]),
        .AD4    (AD[4]),
        .AD5    (AD[5]),
        .AD6    (AD[6]),
        .AD7    (AD[7]),
        .AD8    (AD[8]),
        .AD9    (AD[9]),
        
        .BEN0   (BEN[0]),
        .BEN1   (BEN[1]),
        .BEN2   (BEN[2]),
        .BEN3   (BEN[3]),
        .BEN4   (BEN[4]),
        .BEN5   (BEN[5]),
        .BEN6   (BEN[6]),
        .BEN7   (BEN[7]),
        .BEN8   (BEN[8]),
        .BEN9   (BEN[9]),
        .BEN10   (BEN[10]),
        .BEN11   (BEN[11]),
        .BEN12   (BEN[12]),
        .BEN13   (BEN[13]),
        .BEN14   (BEN[14]),
        .BEN15   (BEN[15]),
        .BEN16   (BEN[16]),
        .BEN17   (BEN[17]),
        .BEN18   (BEN[18]),
        .BEN19   (BEN[19]),
        .BEN20   (BEN[20]),
        .BEN21   (BEN[21]),
        .BEN22   (BEN[22]),
        .BEN23   (BEN[23]),
        .BEN24   (BEN[24]),
        .BEN25   (BEN[25]),
        .BEN26   (BEN[26]),
        .BEN27   (BEN[27]),
        .BEN28   (BEN[28]),
        .BEN29   (BEN[29]),
        .BEN30   (BEN[30]),
        .BEN31   (BEN[31]),
        
        .DI0    (DI[0]),
        .DI1    (DI[1]),
        .DI2    (DI[2]),
        .DI3    (DI[3]),
        .DI4    (DI[4]),
        .DI5    (DI[5]),
        .DI6    (DI[6]),
        .DI7    (DI[7]),
        .DI8    (DI[8]),
        .DI9    (DI[9]),
        .DI10    (DI[10]),
        .DI11    (DI[11]),
        .DI12    (DI[12]),
        .DI13    (DI[13]),
        .DI14    (DI[14]),
        .DI15    (DI[15]),
        .DI16    (DI[16]),
        .DI17    (DI[17]),
        .DI18    (DI[18]),
        .DI19    (DI[19]),
        .DI20    (DI[20]),
        .DI21    (DI[21]),
        .DI22    (DI[22]),
        .DI23    (DI[23]),
        .DI24    (DI[24]),
        .DI25    (DI[25]),
        .DI26    (DI[26]),
        .DI27    (DI[27]),
        .DI28    (DI[28]),
        .DI29    (DI[29]),
        .DI30    (DI[30]),
        .DI31    (DI[31]),
        
        .EN     (EN),

        .R_WB   (R_WB),
        
        .DO0    (DO[0]),
        .DO1    (DO[1]),
        .DO2    (DO[2]),
        .DO3    (DO[3]),
        .DO4    (DO[4]),
        .DO5    (DO[5]),
        .DO6    (DO[6]),
        .DO7    (DO[7]),
        .DO8    (DO[8]),
        .DO9    (DO[9]),
        .DO10    (DO[10]),
        .DO11    (DO[11]),
        .DO12    (DO[12]),
        .DO13    (DO[13]),
        .DO14    (DO[14]),
        .DO15    (DO[15]),
        .DO16    (DO[16]),
        .DO17    (DO[17]),
        .DO18    (DO[18]),
        .DO19    (DO[19]),
        .DO20    (DO[20]),
        .DO21    (DO[21]),
        .DO22    (DO[22]),
        .DO23    (DO[23]),
        .DO24    (DO[24]),
        .DO25    (DO[25]),
        .DO26    (DO[26]),
        .DO27    (DO[27]),
        .DO28    (DO[28]),
        .DO29    (DO[29]),
        .DO30    (DO[30]),
        .DO31    (DO[31])
    );

endmodule

module EF_SRAM_1024x32_wrapper2 (
    input  [ 9:0] AD,
    input  [31:0] BEN,
    input  [31:0] DI,
    input         EN,
    input         R_WB,
    output [31:0] DO
);
    (* keep, BEL="X11Y6.A" *) EF_SRAM_1024x32 i_EF_SRAM_1024x32 (
        .AD0    (AD[0]),
        .AD1    (AD[1]),
        .AD2    (AD[2]),
        .AD3    (AD[3]),
        .AD4    (AD[4]),
        .AD5    (AD[5]),
        .AD6    (AD[6]),
        .AD7    (AD[7]),
        .AD8    (AD[8]),
        .AD9    (AD[9]),
        
        .BEN0   (BEN[0]),
        .BEN1   (BEN[1]),
        .BEN2   (BEN[2]),
        .BEN3   (BEN[3]),
        .BEN4   (BEN[4]),
        .BEN5   (BEN[5]),
        .BEN6   (BEN[6]),
        .BEN7   (BEN[7]),
        .BEN8   (BEN[8]),
        .BEN9   (BEN[9]),
        .BEN10   (BEN[10]),
        .BEN11   (BEN[11]),
        .BEN12   (BEN[12]),
        .BEN13   (BEN[13]),
        .BEN14   (BEN[14]),
        .BEN15   (BEN[15]),
        .BEN16   (BEN[16]),
        .BEN17   (BEN[17]),
        .BEN18   (BEN[18]),
        .BEN19   (BEN[19]),
        .BEN20   (BEN[20]),
        .BEN21   (BEN[21]),
        .BEN22   (BEN[22]),
        .BEN23   (BEN[23]),
        .BEN24   (BEN[24]),
        .BEN25   (BEN[25]),
        .BEN26   (BEN[26]),
        .BEN27   (BEN[27]),
        .BEN28   (BEN[28]),
        .BEN29   (BEN[29]),
        .BEN30   (BEN[30]),
        .BEN31   (BEN[31]),
        
        .DI0    (DI[0]),
        .DI1    (DI[1]),
        .DI2    (DI[2]),
        .DI3    (DI[3]),
        .DI4    (DI[4]),
        .DI5    (DI[5]),
        .DI6    (DI[6]),
        .DI7    (DI[7]),
        .DI8    (DI[8]),
        .DI9    (DI[9]),
        .DI10    (DI[10]),
        .DI11    (DI[11]),
        .DI12    (DI[12]),
        .DI13    (DI[13]),
        .DI14    (DI[14]),
        .DI15    (DI[15]),
        .DI16    (DI[16]),
        .DI17    (DI[17]),
        .DI18    (DI[18]),
        .DI19    (DI[19]),
        .DI20    (DI[20]),
        .DI21    (DI[21]),
        .DI22    (DI[22]),
        .DI23    (DI[23]),
        .DI24    (DI[24]),
        .DI25    (DI[25]),
        .DI26    (DI[26]),
        .DI27    (DI[27]),
        .DI28    (DI[28]),
        .DI29    (DI[29]),
        .DI30    (DI[30]),
        .DI31    (DI[31]),
        
        .EN     (EN),

        .R_WB   (R_WB),
        
        .DO0    (DO[0]),
        .DO1    (DO[1]),
        .DO2    (DO[2]),
        .DO3    (DO[3]),
        .DO4    (DO[4]),
        .DO5    (DO[5]),
        .DO6    (DO[6]),
        .DO7    (DO[7]),
        .DO8    (DO[8]),
        .DO9    (DO[9]),
        .DO10    (DO[10]),
        .DO11    (DO[11]),
        .DO12    (DO[12]),
        .DO13    (DO[13]),
        .DO14    (DO[14]),
        .DO15    (DO[15]),
        .DO16    (DO[16]),
        .DO17    (DO[17]),
        .DO18    (DO[18]),
        .DO19    (DO[19]),
        .DO20    (DO[20]),
        .DO21    (DO[21]),
        .DO22    (DO[22]),
        .DO23    (DO[23]),
        .DO24    (DO[24]),
        .DO25    (DO[25]),
        .DO26    (DO[26]),
        .DO27    (DO[27]),
        .DO28    (DO[28]),
        .DO29    (DO[29]),
        .DO30    (DO[30]),
        .DO31    (DO[31])
    );

endmodule

module EF_SRAM_1024x32_wrapper3 (
    input  [ 9:0] AD,
    input  [31:0] BEN,
    input  [31:0] DI,
    input         EN,
    input         R_WB,
    output [31:0] DO
);
    (* keep, BEL="X11Y8.A" *) EF_SRAM_1024x32 i_EF_SRAM_1024x32 (
        .AD0    (AD[0]),
        .AD1    (AD[1]),
        .AD2    (AD[2]),
        .AD3    (AD[3]),
        .AD4    (AD[4]),
        .AD5    (AD[5]),
        .AD6    (AD[6]),
        .AD7    (AD[7]),
        .AD8    (AD[8]),
        .AD9    (AD[9]),
        
        .BEN0   (BEN[0]),
        .BEN1   (BEN[1]),
        .BEN2   (BEN[2]),
        .BEN3   (BEN[3]),
        .BEN4   (BEN[4]),
        .BEN5   (BEN[5]),
        .BEN6   (BEN[6]),
        .BEN7   (BEN[7]),
        .BEN8   (BEN[8]),
        .BEN9   (BEN[9]),
        .BEN10   (BEN[10]),
        .BEN11   (BEN[11]),
        .BEN12   (BEN[12]),
        .BEN13   (BEN[13]),
        .BEN14   (BEN[14]),
        .BEN15   (BEN[15]),
        .BEN16   (BEN[16]),
        .BEN17   (BEN[17]),
        .BEN18   (BEN[18]),
        .BEN19   (BEN[19]),
        .BEN20   (BEN[20]),
        .BEN21   (BEN[21]),
        .BEN22   (BEN[22]),
        .BEN23   (BEN[23]),
        .BEN24   (BEN[24]),
        .BEN25   (BEN[25]),
        .BEN26   (BEN[26]),
        .BEN27   (BEN[27]),
        .BEN28   (BEN[28]),
        .BEN29   (BEN[29]),
        .BEN30   (BEN[30]),
        .BEN31   (BEN[31]),
        
        .DI0    (DI[0]),
        .DI1    (DI[1]),
        .DI2    (DI[2]),
        .DI3    (DI[3]),
        .DI4    (DI[4]),
        .DI5    (DI[5]),
        .DI6    (DI[6]),
        .DI7    (DI[7]),
        .DI8    (DI[8]),
        .DI9    (DI[9]),
        .DI10    (DI[10]),
        .DI11    (DI[11]),
        .DI12    (DI[12]),
        .DI13    (DI[13]),
        .DI14    (DI[14]),
        .DI15    (DI[15]),
        .DI16    (DI[16]),
        .DI17    (DI[17]),
        .DI18    (DI[18]),
        .DI19    (DI[19]),
        .DI20    (DI[20]),
        .DI21    (DI[21]),
        .DI22    (DI[22]),
        .DI23    (DI[23]),
        .DI24    (DI[24]),
        .DI25    (DI[25]),
        .DI26    (DI[26]),
        .DI27    (DI[27]),
        .DI28    (DI[28]),
        .DI29    (DI[29]),
        .DI30    (DI[30]),
        .DI31    (DI[31]),
        
        .EN     (EN),

        .R_WB   (R_WB),
        
        .DO0    (DO[0]),
        .DO1    (DO[1]),
        .DO2    (DO[2]),
        .DO3    (DO[3]),
        .DO4    (DO[4]),
        .DO5    (DO[5]),
        .DO6    (DO[6]),
        .DO7    (DO[7]),
        .DO8    (DO[8]),
        .DO9    (DO[9]),
        .DO10    (DO[10]),
        .DO11    (DO[11]),
        .DO12    (DO[12]),
        .DO13    (DO[13]),
        .DO14    (DO[14]),
        .DO15    (DO[15]),
        .DO16    (DO[16]),
        .DO17    (DO[17]),
        .DO18    (DO[18]),
        .DO19    (DO[19]),
        .DO20    (DO[20]),
        .DO21    (DO[21]),
        .DO22    (DO[22]),
        .DO23    (DO[23]),
        .DO24    (DO[24]),
        .DO25    (DO[25]),
        .DO26    (DO[26]),
        .DO27    (DO[27]),
        .DO28    (DO[28]),
        .DO29    (DO[29]),
        .DO30    (DO[30]),
        .DO31    (DO[31])
    );

endmodule

module EF_SRAM_1024x32_wrapper4 (
    input  [ 9:0] AD,
    input  [31:0] BEN,
    input  [31:0] DI,
    input         EN,
    input         R_WB,
    output [31:0] DO
);
    (* keep, BEL="X11Y10.A" *) EF_SRAM_1024x32 i_EF_SRAM_1024x32 (
        .AD0    (AD[0]),
        .AD1    (AD[1]),
        .AD2    (AD[2]),
        .AD3    (AD[3]),
        .AD4    (AD[4]),
        .AD5    (AD[5]),
        .AD6    (AD[6]),
        .AD7    (AD[7]),
        .AD8    (AD[8]),
        .AD9    (AD[9]),
        
        .BEN0   (BEN[0]),
        .BEN1   (BEN[1]),
        .BEN2   (BEN[2]),
        .BEN3   (BEN[3]),
        .BEN4   (BEN[4]),
        .BEN5   (BEN[5]),
        .BEN6   (BEN[6]),
        .BEN7   (BEN[7]),
        .BEN8   (BEN[8]),
        .BEN9   (BEN[9]),
        .BEN10   (BEN[10]),
        .BEN11   (BEN[11]),
        .BEN12   (BEN[12]),
        .BEN13   (BEN[13]),
        .BEN14   (BEN[14]),
        .BEN15   (BEN[15]),
        .BEN16   (BEN[16]),
        .BEN17   (BEN[17]),
        .BEN18   (BEN[18]),
        .BEN19   (BEN[19]),
        .BEN20   (BEN[20]),
        .BEN21   (BEN[21]),
        .BEN22   (BEN[22]),
        .BEN23   (BEN[23]),
        .BEN24   (BEN[24]),
        .BEN25   (BEN[25]),
        .BEN26   (BEN[26]),
        .BEN27   (BEN[27]),
        .BEN28   (BEN[28]),
        .BEN29   (BEN[29]),
        .BEN30   (BEN[30]),
        .BEN31   (BEN[31]),
        
        .DI0    (DI[0]),
        .DI1    (DI[1]),
        .DI2    (DI[2]),
        .DI3    (DI[3]),
        .DI4    (DI[4]),
        .DI5    (DI[5]),
        .DI6    (DI[6]),
        .DI7    (DI[7]),
        .DI8    (DI[8]),
        .DI9    (DI[9]),
        .DI10    (DI[10]),
        .DI11    (DI[11]),
        .DI12    (DI[12]),
        .DI13    (DI[13]),
        .DI14    (DI[14]),
        .DI15    (DI[15]),
        .DI16    (DI[16]),
        .DI17    (DI[17]),
        .DI18    (DI[18]),
        .DI19    (DI[19]),
        .DI20    (DI[20]),
        .DI21    (DI[21]),
        .DI22    (DI[22]),
        .DI23    (DI[23]),
        .DI24    (DI[24]),
        .DI25    (DI[25]),
        .DI26    (DI[26]),
        .DI27    (DI[27]),
        .DI28    (DI[28]),
        .DI29    (DI[29]),
        .DI30    (DI[30]),
        .DI31    (DI[31]),
        
        .EN     (EN),

        .R_WB   (R_WB),
        
        .DO0    (DO[0]),
        .DO1    (DO[1]),
        .DO2    (DO[2]),
        .DO3    (DO[3]),
        .DO4    (DO[4]),
        .DO5    (DO[5]),
        .DO6    (DO[6]),
        .DO7    (DO[7]),
        .DO8    (DO[8]),
        .DO9    (DO[9]),
        .DO10    (DO[10]),
        .DO11    (DO[11]),
        .DO12    (DO[12]),
        .DO13    (DO[13]),
        .DO14    (DO[14]),
        .DO15    (DO[15]),
        .DO16    (DO[16]),
        .DO17    (DO[17]),
        .DO18    (DO[18]),
        .DO19    (DO[19]),
        .DO20    (DO[20]),
        .DO21    (DO[21]),
        .DO22    (DO[22]),
        .DO23    (DO[23]),
        .DO24    (DO[24]),
        .DO25    (DO[25]),
        .DO26    (DO[26]),
        .DO27    (DO[27]),
        .DO28    (DO[28]),
        .DO29    (DO[29]),
        .DO30    (DO[30]),
        .DO31    (DO[31])
    );

endmodule

module EF_SRAM_1024x32_wrapper5 (
    input  [ 9:0] AD,
    input  [31:0] BEN,
    input  [31:0] DI,
    input         EN,
    input         R_WB,
    output [31:0] DO
);
    (* keep, BEL="X11Y12.A" *) EF_SRAM_1024x32 i_EF_SRAM_1024x32 (
        .AD0    (AD[0]),
        .AD1    (AD[1]),
        .AD2    (AD[2]),
        .AD3    (AD[3]),
        .AD4    (AD[4]),
        .AD5    (AD[5]),
        .AD6    (AD[6]),
        .AD7    (AD[7]),
        .AD8    (AD[8]),
        .AD9    (AD[9]),
        
        .BEN0   (BEN[0]),
        .BEN1   (BEN[1]),
        .BEN2   (BEN[2]),
        .BEN3   (BEN[3]),
        .BEN4   (BEN[4]),
        .BEN5   (BEN[5]),
        .BEN6   (BEN[6]),
        .BEN7   (BEN[7]),
        .BEN8   (BEN[8]),
        .BEN9   (BEN[9]),
        .BEN10   (BEN[10]),
        .BEN11   (BEN[11]),
        .BEN12   (BEN[12]),
        .BEN13   (BEN[13]),
        .BEN14   (BEN[14]),
        .BEN15   (BEN[15]),
        .BEN16   (BEN[16]),
        .BEN17   (BEN[17]),
        .BEN18   (BEN[18]),
        .BEN19   (BEN[19]),
        .BEN20   (BEN[20]),
        .BEN21   (BEN[21]),
        .BEN22   (BEN[22]),
        .BEN23   (BEN[23]),
        .BEN24   (BEN[24]),
        .BEN25   (BEN[25]),
        .BEN26   (BEN[26]),
        .BEN27   (BEN[27]),
        .BEN28   (BEN[28]),
        .BEN29   (BEN[29]),
        .BEN30   (BEN[30]),
        .BEN31   (BEN[31]),
        
        .DI0    (DI[0]),
        .DI1    (DI[1]),
        .DI2    (DI[2]),
        .DI3    (DI[3]),
        .DI4    (DI[4]),
        .DI5    (DI[5]),
        .DI6    (DI[6]),
        .DI7    (DI[7]),
        .DI8    (DI[8]),
        .DI9    (DI[9]),
        .DI10    (DI[10]),
        .DI11    (DI[11]),
        .DI12    (DI[12]),
        .DI13    (DI[13]),
        .DI14    (DI[14]),
        .DI15    (DI[15]),
        .DI16    (DI[16]),
        .DI17    (DI[17]),
        .DI18    (DI[18]),
        .DI19    (DI[19]),
        .DI20    (DI[20]),
        .DI21    (DI[21]),
        .DI22    (DI[22]),
        .DI23    (DI[23]),
        .DI24    (DI[24]),
        .DI25    (DI[25]),
        .DI26    (DI[26]),
        .DI27    (DI[27]),
        .DI28    (DI[28]),
        .DI29    (DI[29]),
        .DI30    (DI[30]),
        .DI31    (DI[31]),
        
        .EN     (EN),

        .R_WB   (R_WB),
        
        .DO0    (DO[0]),
        .DO1    (DO[1]),
        .DO2    (DO[2]),
        .DO3    (DO[3]),
        .DO4    (DO[4]),
        .DO5    (DO[5]),
        .DO6    (DO[6]),
        .DO7    (DO[7]),
        .DO8    (DO[8]),
        .DO9    (DO[9]),
        .DO10    (DO[10]),
        .DO11    (DO[11]),
        .DO12    (DO[12]),
        .DO13    (DO[13]),
        .DO14    (DO[14]),
        .DO15    (DO[15]),
        .DO16    (DO[16]),
        .DO17    (DO[17]),
        .DO18    (DO[18]),
        .DO19    (DO[19]),
        .DO20    (DO[20]),
        .DO21    (DO[21]),
        .DO22    (DO[22]),
        .DO23    (DO[23]),
        .DO24    (DO[24]),
        .DO25    (DO[25]),
        .DO26    (DO[26]),
        .DO27    (DO[27]),
        .DO28    (DO[28]),
        .DO29    (DO[29]),
        .DO30    (DO[30]),
        .DO31    (DO[31])
    );

endmodule

module EF_SRAM_1024x32_wrapper6 (
    input  [ 9:0] AD,
    input  [31:0] BEN,
    input  [31:0] DI,
    input         EN,
    input         R_WB,
    output [31:0] DO
);
    (* keep, BEL="X11Y14.A" *) EF_SRAM_1024x32 i_EF_SRAM_1024x32 (
        .AD0    (AD[0]),
        .AD1    (AD[1]),
        .AD2    (AD[2]),
        .AD3    (AD[3]),
        .AD4    (AD[4]),
        .AD5    (AD[5]),
        .AD6    (AD[6]),
        .AD7    (AD[7]),
        .AD8    (AD[8]),
        .AD9    (AD[9]),
        
        .BEN0   (BEN[0]),
        .BEN1   (BEN[1]),
        .BEN2   (BEN[2]),
        .BEN3   (BEN[3]),
        .BEN4   (BEN[4]),
        .BEN5   (BEN[5]),
        .BEN6   (BEN[6]),
        .BEN7   (BEN[7]),
        .BEN8   (BEN[8]),
        .BEN9   (BEN[9]),
        .BEN10   (BEN[10]),
        .BEN11   (BEN[11]),
        .BEN12   (BEN[12]),
        .BEN13   (BEN[13]),
        .BEN14   (BEN[14]),
        .BEN15   (BEN[15]),
        .BEN16   (BEN[16]),
        .BEN17   (BEN[17]),
        .BEN18   (BEN[18]),
        .BEN19   (BEN[19]),
        .BEN20   (BEN[20]),
        .BEN21   (BEN[21]),
        .BEN22   (BEN[22]),
        .BEN23   (BEN[23]),
        .BEN24   (BEN[24]),
        .BEN25   (BEN[25]),
        .BEN26   (BEN[26]),
        .BEN27   (BEN[27]),
        .BEN28   (BEN[28]),
        .BEN29   (BEN[29]),
        .BEN30   (BEN[30]),
        .BEN31   (BEN[31]),
        
        .DI0    (DI[0]),
        .DI1    (DI[1]),
        .DI2    (DI[2]),
        .DI3    (DI[3]),
        .DI4    (DI[4]),
        .DI5    (DI[5]),
        .DI6    (DI[6]),
        .DI7    (DI[7]),
        .DI8    (DI[8]),
        .DI9    (DI[9]),
        .DI10    (DI[10]),
        .DI11    (DI[11]),
        .DI12    (DI[12]),
        .DI13    (DI[13]),
        .DI14    (DI[14]),
        .DI15    (DI[15]),
        .DI16    (DI[16]),
        .DI17    (DI[17]),
        .DI18    (DI[18]),
        .DI19    (DI[19]),
        .DI20    (DI[20]),
        .DI21    (DI[21]),
        .DI22    (DI[22]),
        .DI23    (DI[23]),
        .DI24    (DI[24]),
        .DI25    (DI[25]),
        .DI26    (DI[26]),
        .DI27    (DI[27]),
        .DI28    (DI[28]),
        .DI29    (DI[29]),
        .DI30    (DI[30]),
        .DI31    (DI[31]),
        
        .EN     (EN),

        .R_WB   (R_WB),
        
        .DO0    (DO[0]),
        .DO1    (DO[1]),
        .DO2    (DO[2]),
        .DO3    (DO[3]),
        .DO4    (DO[4]),
        .DO5    (DO[5]),
        .DO6    (DO[6]),
        .DO7    (DO[7]),
        .DO8    (DO[8]),
        .DO9    (DO[9]),
        .DO10    (DO[10]),
        .DO11    (DO[11]),
        .DO12    (DO[12]),
        .DO13    (DO[13]),
        .DO14    (DO[14]),
        .DO15    (DO[15]),
        .DO16    (DO[16]),
        .DO17    (DO[17]),
        .DO18    (DO[18]),
        .DO19    (DO[19]),
        .DO20    (DO[20]),
        .DO21    (DO[21]),
        .DO22    (DO[22]),
        .DO23    (DO[23]),
        .DO24    (DO[24]),
        .DO25    (DO[25]),
        .DO26    (DO[26]),
        .DO27    (DO[27]),
        .DO28    (DO[28]),
        .DO29    (DO[29]),
        .DO30    (DO[30]),
        .DO31    (DO[31])
    );

endmodule

module EF_SRAM_1024x32_wrapper7 (
    input  [ 9:0] AD,
    input  [31:0] BEN,
    input  [31:0] DI,
    input         EN,
    input         R_WB,
    output [31:0] DO
);
    (* keep, BEL="X11Y16.A" *) EF_SRAM_1024x32 i_EF_SRAM_1024x32 (
        .AD0    (AD[0]),
        .AD1    (AD[1]),
        .AD2    (AD[2]),
        .AD3    (AD[3]),
        .AD4    (AD[4]),
        .AD5    (AD[5]),
        .AD6    (AD[6]),
        .AD7    (AD[7]),
        .AD8    (AD[8]),
        .AD9    (AD[9]),
        
        .BEN0   (BEN[0]),
        .BEN1   (BEN[1]),
        .BEN2   (BEN[2]),
        .BEN3   (BEN[3]),
        .BEN4   (BEN[4]),
        .BEN5   (BEN[5]),
        .BEN6   (BEN[6]),
        .BEN7   (BEN[7]),
        .BEN8   (BEN[8]),
        .BEN9   (BEN[9]),
        .BEN10   (BEN[10]),
        .BEN11   (BEN[11]),
        .BEN12   (BEN[12]),
        .BEN13   (BEN[13]),
        .BEN14   (BEN[14]),
        .BEN15   (BEN[15]),
        .BEN16   (BEN[16]),
        .BEN17   (BEN[17]),
        .BEN18   (BEN[18]),
        .BEN19   (BEN[19]),
        .BEN20   (BEN[20]),
        .BEN21   (BEN[21]),
        .BEN22   (BEN[22]),
        .BEN23   (BEN[23]),
        .BEN24   (BEN[24]),
        .BEN25   (BEN[25]),
        .BEN26   (BEN[26]),
        .BEN27   (BEN[27]),
        .BEN28   (BEN[28]),
        .BEN29   (BEN[29]),
        .BEN30   (BEN[30]),
        .BEN31   (BEN[31]),
        
        .DI0    (DI[0]),
        .DI1    (DI[1]),
        .DI2    (DI[2]),
        .DI3    (DI[3]),
        .DI4    (DI[4]),
        .DI5    (DI[5]),
        .DI6    (DI[6]),
        .DI7    (DI[7]),
        .DI8    (DI[8]),
        .DI9    (DI[9]),
        .DI10    (DI[10]),
        .DI11    (DI[11]),
        .DI12    (DI[12]),
        .DI13    (DI[13]),
        .DI14    (DI[14]),
        .DI15    (DI[15]),
        .DI16    (DI[16]),
        .DI17    (DI[17]),
        .DI18    (DI[18]),
        .DI19    (DI[19]),
        .DI20    (DI[20]),
        .DI21    (DI[21]),
        .DI22    (DI[22]),
        .DI23    (DI[23]),
        .DI24    (DI[24]),
        .DI25    (DI[25]),
        .DI26    (DI[26]),
        .DI27    (DI[27]),
        .DI28    (DI[28]),
        .DI29    (DI[29]),
        .DI30    (DI[30]),
        .DI31    (DI[31]),
        
        .EN     (EN),

        .R_WB   (R_WB),
        
        .DO0    (DO[0]),
        .DO1    (DO[1]),
        .DO2    (DO[2]),
        .DO3    (DO[3]),
        .DO4    (DO[4]),
        .DO5    (DO[5]),
        .DO6    (DO[6]),
        .DO7    (DO[7]),
        .DO8    (DO[8]),
        .DO9    (DO[9]),
        .DO10    (DO[10]),
        .DO11    (DO[11]),
        .DO12    (DO[12]),
        .DO13    (DO[13]),
        .DO14    (DO[14]),
        .DO15    (DO[15]),
        .DO16    (DO[16]),
        .DO17    (DO[17]),
        .DO18    (DO[18]),
        .DO19    (DO[19]),
        .DO20    (DO[20]),
        .DO21    (DO[21]),
        .DO22    (DO[22]),
        .DO23    (DO[23]),
        .DO24    (DO[24]),
        .DO25    (DO[25]),
        .DO26    (DO[26]),
        .DO27    (DO[27]),
        .DO28    (DO[28]),
        .DO29    (DO[29]),
        .DO30    (DO[30]),
        .DO31    (DO[31])
    );

endmodule
