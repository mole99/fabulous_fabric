VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO eFPGA
  CLASS BLOCK ;
  FOREIGN eFPGA ;
  ORIGIN 0.000 0.000 ;
  SIZE 2263.200 BY 3511.680 ;
  PIN FrameData[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 3453.880 0.480 3454.280 ;
    END
  END FrameData[0]
  PIN FrameData[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2822.200 0.860 2822.600 ;
    END
  END FrameData[100]
  PIN FrameData[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2827.240 0.860 2827.640 ;
    END
  END FrameData[101]
  PIN FrameData[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2832.280 0.930 2832.680 ;
    END
  END FrameData[102]
  PIN FrameData[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2837.320 0.860 2837.720 ;
    END
  END FrameData[103]
  PIN FrameData[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2842.360 0.930 2842.760 ;
    END
  END FrameData[104]
  PIN FrameData[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2847.400 0.930 2847.800 ;
    END
  END FrameData[105]
  PIN FrameData[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2852.440 0.930 2852.840 ;
    END
  END FrameData[106]
  PIN FrameData[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2857.480 0.930 2857.880 ;
    END
  END FrameData[107]
  PIN FrameData[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2862.520 0.930 2862.920 ;
    END
  END FrameData[108]
  PIN FrameData[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2867.560 0.860 2867.960 ;
    END
  END FrameData[109]
  PIN FrameData[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 3470.680 0.480 3471.080 ;
    END
  END FrameData[10]
  PIN FrameData[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2872.600 0.860 2873.000 ;
    END
  END FrameData[110]
  PIN FrameData[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2877.640 0.930 2878.040 ;
    END
  END FrameData[111]
  PIN FrameData[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2882.680 0.860 2883.080 ;
    END
  END FrameData[112]
  PIN FrameData[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2887.720 0.860 2888.120 ;
    END
  END FrameData[113]
  PIN FrameData[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2892.760 0.930 2893.160 ;
    END
  END FrameData[114]
  PIN FrameData[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2897.800 0.860 2898.200 ;
    END
  END FrameData[115]
  PIN FrameData[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2902.840 0.860 2903.240 ;
    END
  END FrameData[116]
  PIN FrameData[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2907.880 0.930 2908.280 ;
    END
  END FrameData[117]
  PIN FrameData[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2912.920 0.860 2913.320 ;
    END
  END FrameData[118]
  PIN FrameData[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2917.960 0.860 2918.360 ;
    END
  END FrameData[119]
  PIN FrameData[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 3472.360 0.480 3472.760 ;
    END
  END FrameData[11]
  PIN FrameData[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2923.000 0.930 2923.400 ;
    END
  END FrameData[120]
  PIN FrameData[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2928.040 0.860 2928.440 ;
    END
  END FrameData[121]
  PIN FrameData[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2933.080 0.860 2933.480 ;
    END
  END FrameData[122]
  PIN FrameData[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2938.120 0.930 2938.520 ;
    END
  END FrameData[123]
  PIN FrameData[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2943.160 0.860 2943.560 ;
    END
  END FrameData[124]
  PIN FrameData[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2948.200 0.860 2948.600 ;
    END
  END FrameData[125]
  PIN FrameData[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2953.240 0.930 2953.640 ;
    END
  END FrameData[126]
  PIN FrameData[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2958.280 0.930 2958.680 ;
    END
  END FrameData[127]
  PIN FrameData[128]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2560.120 0.930 2560.520 ;
    END
  END FrameData[128]
  PIN FrameData[129]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2565.160 0.860 2565.560 ;
    END
  END FrameData[129]
  PIN FrameData[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 3474.040 0.480 3474.440 ;
    END
  END FrameData[12]
  PIN FrameData[130]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2570.200 0.860 2570.600 ;
    END
  END FrameData[130]
  PIN FrameData[131]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2575.240 0.860 2575.640 ;
    END
  END FrameData[131]
  PIN FrameData[132]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2580.280 0.860 2580.680 ;
    END
  END FrameData[132]
  PIN FrameData[133]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2585.320 0.860 2585.720 ;
    END
  END FrameData[133]
  PIN FrameData[134]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2590.360 0.930 2590.760 ;
    END
  END FrameData[134]
  PIN FrameData[135]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2595.400 0.860 2595.800 ;
    END
  END FrameData[135]
  PIN FrameData[136]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2600.440 0.930 2600.840 ;
    END
  END FrameData[136]
  PIN FrameData[137]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2605.480 0.930 2605.880 ;
    END
  END FrameData[137]
  PIN FrameData[138]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2610.520 0.930 2610.920 ;
    END
  END FrameData[138]
  PIN FrameData[139]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2615.560 0.930 2615.960 ;
    END
  END FrameData[139]
  PIN FrameData[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 3475.720 0.480 3476.120 ;
    END
  END FrameData[13]
  PIN FrameData[140]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2620.600 0.930 2621.000 ;
    END
  END FrameData[140]
  PIN FrameData[141]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2625.640 0.860 2626.040 ;
    END
  END FrameData[141]
  PIN FrameData[142]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2630.680 0.860 2631.080 ;
    END
  END FrameData[142]
  PIN FrameData[143]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2635.720 0.930 2636.120 ;
    END
  END FrameData[143]
  PIN FrameData[144]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2640.760 0.860 2641.160 ;
    END
  END FrameData[144]
  PIN FrameData[145]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2645.800 0.860 2646.200 ;
    END
  END FrameData[145]
  PIN FrameData[146]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2650.840 0.930 2651.240 ;
    END
  END FrameData[146]
  PIN FrameData[147]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2655.880 0.860 2656.280 ;
    END
  END FrameData[147]
  PIN FrameData[148]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2660.920 0.860 2661.320 ;
    END
  END FrameData[148]
  PIN FrameData[149]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2665.960 0.930 2666.360 ;
    END
  END FrameData[149]
  PIN FrameData[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 3477.400 0.480 3477.800 ;
    END
  END FrameData[14]
  PIN FrameData[150]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2671.000 0.860 2671.400 ;
    END
  END FrameData[150]
  PIN FrameData[151]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2676.040 0.860 2676.440 ;
    END
  END FrameData[151]
  PIN FrameData[152]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2681.080 0.930 2681.480 ;
    END
  END FrameData[152]
  PIN FrameData[153]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2686.120 0.860 2686.520 ;
    END
  END FrameData[153]
  PIN FrameData[154]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2691.160 0.860 2691.560 ;
    END
  END FrameData[154]
  PIN FrameData[155]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2696.200 0.930 2696.600 ;
    END
  END FrameData[155]
  PIN FrameData[156]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2701.240 0.860 2701.640 ;
    END
  END FrameData[156]
  PIN FrameData[157]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2706.280 0.860 2706.680 ;
    END
  END FrameData[157]
  PIN FrameData[158]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2711.320 0.930 2711.720 ;
    END
  END FrameData[158]
  PIN FrameData[159]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2716.360 0.930 2716.760 ;
    END
  END FrameData[159]
  PIN FrameData[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 3479.080 0.480 3479.480 ;
    END
  END FrameData[15]
  PIN FrameData[160]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2318.200 0.930 2318.600 ;
    END
  END FrameData[160]
  PIN FrameData[161]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2323.240 0.860 2323.640 ;
    END
  END FrameData[161]
  PIN FrameData[162]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2328.280 0.860 2328.680 ;
    END
  END FrameData[162]
  PIN FrameData[163]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2333.320 0.860 2333.720 ;
    END
  END FrameData[163]
  PIN FrameData[164]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2338.360 0.860 2338.760 ;
    END
  END FrameData[164]
  PIN FrameData[165]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2343.400 0.860 2343.800 ;
    END
  END FrameData[165]
  PIN FrameData[166]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2348.440 0.930 2348.840 ;
    END
  END FrameData[166]
  PIN FrameData[167]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2353.480 0.860 2353.880 ;
    END
  END FrameData[167]
  PIN FrameData[168]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2358.520 0.930 2358.920 ;
    END
  END FrameData[168]
  PIN FrameData[169]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2363.560 0.930 2363.960 ;
    END
  END FrameData[169]
  PIN FrameData[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 3480.760 0.480 3481.160 ;
    END
  END FrameData[16]
  PIN FrameData[170]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2368.600 0.930 2369.000 ;
    END
  END FrameData[170]
  PIN FrameData[171]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2373.640 0.930 2374.040 ;
    END
  END FrameData[171]
  PIN FrameData[172]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2378.680 0.930 2379.080 ;
    END
  END FrameData[172]
  PIN FrameData[173]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2383.720 0.860 2384.120 ;
    END
  END FrameData[173]
  PIN FrameData[174]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2388.760 0.860 2389.160 ;
    END
  END FrameData[174]
  PIN FrameData[175]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2393.800 0.930 2394.200 ;
    END
  END FrameData[175]
  PIN FrameData[176]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2398.840 0.860 2399.240 ;
    END
  END FrameData[176]
  PIN FrameData[177]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2403.880 0.860 2404.280 ;
    END
  END FrameData[177]
  PIN FrameData[178]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2408.920 0.930 2409.320 ;
    END
  END FrameData[178]
  PIN FrameData[179]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2413.960 0.860 2414.360 ;
    END
  END FrameData[179]
  PIN FrameData[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 3482.440 0.480 3482.840 ;
    END
  END FrameData[17]
  PIN FrameData[180]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2419.000 0.860 2419.400 ;
    END
  END FrameData[180]
  PIN FrameData[181]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2424.040 0.930 2424.440 ;
    END
  END FrameData[181]
  PIN FrameData[182]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2429.080 0.860 2429.480 ;
    END
  END FrameData[182]
  PIN FrameData[183]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2434.120 0.860 2434.520 ;
    END
  END FrameData[183]
  PIN FrameData[184]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2439.160 0.930 2439.560 ;
    END
  END FrameData[184]
  PIN FrameData[185]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2444.200 0.860 2444.600 ;
    END
  END FrameData[185]
  PIN FrameData[186]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2449.240 0.860 2449.640 ;
    END
  END FrameData[186]
  PIN FrameData[187]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2454.280 0.930 2454.680 ;
    END
  END FrameData[187]
  PIN FrameData[188]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2459.320 0.860 2459.720 ;
    END
  END FrameData[188]
  PIN FrameData[189]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2464.360 0.860 2464.760 ;
    END
  END FrameData[189]
  PIN FrameData[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 3484.120 0.480 3484.520 ;
    END
  END FrameData[18]
  PIN FrameData[190]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2469.400 0.930 2469.800 ;
    END
  END FrameData[190]
  PIN FrameData[191]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2474.440 0.930 2474.840 ;
    END
  END FrameData[191]
  PIN FrameData[192]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2076.280 0.930 2076.680 ;
    END
  END FrameData[192]
  PIN FrameData[193]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2081.320 0.860 2081.720 ;
    END
  END FrameData[193]
  PIN FrameData[194]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2086.360 0.860 2086.760 ;
    END
  END FrameData[194]
  PIN FrameData[195]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2091.400 0.860 2091.800 ;
    END
  END FrameData[195]
  PIN FrameData[196]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2096.440 0.860 2096.840 ;
    END
  END FrameData[196]
  PIN FrameData[197]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2101.480 0.860 2101.880 ;
    END
  END FrameData[197]
  PIN FrameData[198]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2106.520 0.930 2106.920 ;
    END
  END FrameData[198]
  PIN FrameData[199]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2111.560 0.860 2111.960 ;
    END
  END FrameData[199]
  PIN FrameData[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 3485.800 0.480 3486.200 ;
    END
  END FrameData[19]
  PIN FrameData[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 3455.560 0.480 3455.960 ;
    END
  END FrameData[1]
  PIN FrameData[200]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2116.600 0.930 2117.000 ;
    END
  END FrameData[200]
  PIN FrameData[201]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2121.640 0.930 2122.040 ;
    END
  END FrameData[201]
  PIN FrameData[202]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2126.680 0.930 2127.080 ;
    END
  END FrameData[202]
  PIN FrameData[203]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2131.720 0.930 2132.120 ;
    END
  END FrameData[203]
  PIN FrameData[204]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2136.760 0.930 2137.160 ;
    END
  END FrameData[204]
  PIN FrameData[205]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2141.800 0.860 2142.200 ;
    END
  END FrameData[205]
  PIN FrameData[206]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2146.840 0.860 2147.240 ;
    END
  END FrameData[206]
  PIN FrameData[207]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2151.880 0.930 2152.280 ;
    END
  END FrameData[207]
  PIN FrameData[208]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2156.920 0.860 2157.320 ;
    END
  END FrameData[208]
  PIN FrameData[209]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2161.960 0.860 2162.360 ;
    END
  END FrameData[209]
  PIN FrameData[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 3487.480 0.480 3487.880 ;
    END
  END FrameData[20]
  PIN FrameData[210]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2167.000 0.930 2167.400 ;
    END
  END FrameData[210]
  PIN FrameData[211]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2172.040 0.860 2172.440 ;
    END
  END FrameData[211]
  PIN FrameData[212]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2177.080 0.860 2177.480 ;
    END
  END FrameData[212]
  PIN FrameData[213]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2182.120 0.930 2182.520 ;
    END
  END FrameData[213]
  PIN FrameData[214]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2187.160 0.860 2187.560 ;
    END
  END FrameData[214]
  PIN FrameData[215]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2192.200 0.860 2192.600 ;
    END
  END FrameData[215]
  PIN FrameData[216]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2197.240 0.930 2197.640 ;
    END
  END FrameData[216]
  PIN FrameData[217]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2202.280 0.860 2202.680 ;
    END
  END FrameData[217]
  PIN FrameData[218]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2207.320 0.860 2207.720 ;
    END
  END FrameData[218]
  PIN FrameData[219]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2212.360 0.930 2212.760 ;
    END
  END FrameData[219]
  PIN FrameData[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 3489.160 0.480 3489.560 ;
    END
  END FrameData[21]
  PIN FrameData[220]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2217.400 0.860 2217.800 ;
    END
  END FrameData[220]
  PIN FrameData[221]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2222.440 0.860 2222.840 ;
    END
  END FrameData[221]
  PIN FrameData[222]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2227.480 0.930 2227.880 ;
    END
  END FrameData[222]
  PIN FrameData[223]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2232.520 0.930 2232.920 ;
    END
  END FrameData[223]
  PIN FrameData[224]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1834.360 0.930 1834.760 ;
    END
  END FrameData[224]
  PIN FrameData[225]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1839.400 0.860 1839.800 ;
    END
  END FrameData[225]
  PIN FrameData[226]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1844.440 0.860 1844.840 ;
    END
  END FrameData[226]
  PIN FrameData[227]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1849.480 0.860 1849.880 ;
    END
  END FrameData[227]
  PIN FrameData[228]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1854.520 0.860 1854.920 ;
    END
  END FrameData[228]
  PIN FrameData[229]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1859.560 0.860 1859.960 ;
    END
  END FrameData[229]
  PIN FrameData[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 3490.840 0.480 3491.240 ;
    END
  END FrameData[22]
  PIN FrameData[230]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1864.600 0.930 1865.000 ;
    END
  END FrameData[230]
  PIN FrameData[231]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1869.640 0.860 1870.040 ;
    END
  END FrameData[231]
  PIN FrameData[232]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1874.680 0.930 1875.080 ;
    END
  END FrameData[232]
  PIN FrameData[233]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1879.720 0.930 1880.120 ;
    END
  END FrameData[233]
  PIN FrameData[234]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1884.760 0.930 1885.160 ;
    END
  END FrameData[234]
  PIN FrameData[235]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1889.800 0.930 1890.200 ;
    END
  END FrameData[235]
  PIN FrameData[236]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1894.840 0.930 1895.240 ;
    END
  END FrameData[236]
  PIN FrameData[237]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1899.880 0.860 1900.280 ;
    END
  END FrameData[237]
  PIN FrameData[238]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1904.920 0.860 1905.320 ;
    END
  END FrameData[238]
  PIN FrameData[239]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1909.960 0.930 1910.360 ;
    END
  END FrameData[239]
  PIN FrameData[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 3492.520 0.480 3492.920 ;
    END
  END FrameData[23]
  PIN FrameData[240]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1915.000 0.860 1915.400 ;
    END
  END FrameData[240]
  PIN FrameData[241]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1920.040 0.860 1920.440 ;
    END
  END FrameData[241]
  PIN FrameData[242]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1925.080 0.930 1925.480 ;
    END
  END FrameData[242]
  PIN FrameData[243]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1930.120 0.860 1930.520 ;
    END
  END FrameData[243]
  PIN FrameData[244]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1935.160 0.860 1935.560 ;
    END
  END FrameData[244]
  PIN FrameData[245]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1940.200 0.930 1940.600 ;
    END
  END FrameData[245]
  PIN FrameData[246]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1945.240 0.860 1945.640 ;
    END
  END FrameData[246]
  PIN FrameData[247]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1950.280 0.860 1950.680 ;
    END
  END FrameData[247]
  PIN FrameData[248]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1955.320 0.930 1955.720 ;
    END
  END FrameData[248]
  PIN FrameData[249]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1960.360 0.860 1960.760 ;
    END
  END FrameData[249]
  PIN FrameData[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 3494.200 0.480 3494.600 ;
    END
  END FrameData[24]
  PIN FrameData[250]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1965.400 0.860 1965.800 ;
    END
  END FrameData[250]
  PIN FrameData[251]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1970.440 0.930 1970.840 ;
    END
  END FrameData[251]
  PIN FrameData[252]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1975.480 0.860 1975.880 ;
    END
  END FrameData[252]
  PIN FrameData[253]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1980.520 0.860 1980.920 ;
    END
  END FrameData[253]
  PIN FrameData[254]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1985.560 0.930 1985.960 ;
    END
  END FrameData[254]
  PIN FrameData[255]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1990.600 0.930 1991.000 ;
    END
  END FrameData[255]
  PIN FrameData[256]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1592.440 0.930 1592.840 ;
    END
  END FrameData[256]
  PIN FrameData[257]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1597.480 0.860 1597.880 ;
    END
  END FrameData[257]
  PIN FrameData[258]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1602.520 0.860 1602.920 ;
    END
  END FrameData[258]
  PIN FrameData[259]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1607.560 0.860 1607.960 ;
    END
  END FrameData[259]
  PIN FrameData[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 3495.880 0.480 3496.280 ;
    END
  END FrameData[25]
  PIN FrameData[260]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1612.600 0.860 1613.000 ;
    END
  END FrameData[260]
  PIN FrameData[261]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1617.640 0.860 1618.040 ;
    END
  END FrameData[261]
  PIN FrameData[262]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1622.680 0.930 1623.080 ;
    END
  END FrameData[262]
  PIN FrameData[263]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1627.720 0.860 1628.120 ;
    END
  END FrameData[263]
  PIN FrameData[264]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1632.760 0.930 1633.160 ;
    END
  END FrameData[264]
  PIN FrameData[265]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1637.800 0.930 1638.200 ;
    END
  END FrameData[265]
  PIN FrameData[266]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1642.840 0.930 1643.240 ;
    END
  END FrameData[266]
  PIN FrameData[267]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1647.880 0.930 1648.280 ;
    END
  END FrameData[267]
  PIN FrameData[268]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1652.920 0.930 1653.320 ;
    END
  END FrameData[268]
  PIN FrameData[269]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1657.960 0.860 1658.360 ;
    END
  END FrameData[269]
  PIN FrameData[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 3497.560 0.480 3497.960 ;
    END
  END FrameData[26]
  PIN FrameData[270]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1663.000 0.860 1663.400 ;
    END
  END FrameData[270]
  PIN FrameData[271]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1668.040 0.930 1668.440 ;
    END
  END FrameData[271]
  PIN FrameData[272]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1673.080 0.860 1673.480 ;
    END
  END FrameData[272]
  PIN FrameData[273]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1678.120 0.860 1678.520 ;
    END
  END FrameData[273]
  PIN FrameData[274]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1683.160 0.930 1683.560 ;
    END
  END FrameData[274]
  PIN FrameData[275]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1688.200 0.860 1688.600 ;
    END
  END FrameData[275]
  PIN FrameData[276]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1693.240 0.860 1693.640 ;
    END
  END FrameData[276]
  PIN FrameData[277]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1698.280 0.930 1698.680 ;
    END
  END FrameData[277]
  PIN FrameData[278]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1703.320 0.860 1703.720 ;
    END
  END FrameData[278]
  PIN FrameData[279]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1708.360 0.860 1708.760 ;
    END
  END FrameData[279]
  PIN FrameData[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 3499.240 0.480 3499.640 ;
    END
  END FrameData[27]
  PIN FrameData[280]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1713.400 0.930 1713.800 ;
    END
  END FrameData[280]
  PIN FrameData[281]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1718.440 0.860 1718.840 ;
    END
  END FrameData[281]
  PIN FrameData[282]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1723.480 0.860 1723.880 ;
    END
  END FrameData[282]
  PIN FrameData[283]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1728.520 0.930 1728.920 ;
    END
  END FrameData[283]
  PIN FrameData[284]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1733.560 0.860 1733.960 ;
    END
  END FrameData[284]
  PIN FrameData[285]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1738.600 0.860 1739.000 ;
    END
  END FrameData[285]
  PIN FrameData[286]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1743.640 0.930 1744.040 ;
    END
  END FrameData[286]
  PIN FrameData[287]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1748.680 0.930 1749.080 ;
    END
  END FrameData[287]
  PIN FrameData[288]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1350.520 0.930 1350.920 ;
    END
  END FrameData[288]
  PIN FrameData[289]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1355.560 0.860 1355.960 ;
    END
  END FrameData[289]
  PIN FrameData[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 3500.920 0.480 3501.320 ;
    END
  END FrameData[28]
  PIN FrameData[290]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1360.600 0.860 1361.000 ;
    END
  END FrameData[290]
  PIN FrameData[291]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1365.640 0.860 1366.040 ;
    END
  END FrameData[291]
  PIN FrameData[292]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1370.680 0.860 1371.080 ;
    END
  END FrameData[292]
  PIN FrameData[293]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1375.720 0.860 1376.120 ;
    END
  END FrameData[293]
  PIN FrameData[294]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1380.760 0.930 1381.160 ;
    END
  END FrameData[294]
  PIN FrameData[295]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1385.800 0.860 1386.200 ;
    END
  END FrameData[295]
  PIN FrameData[296]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1390.840 0.930 1391.240 ;
    END
  END FrameData[296]
  PIN FrameData[297]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1395.880 0.930 1396.280 ;
    END
  END FrameData[297]
  PIN FrameData[298]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1400.920 0.930 1401.320 ;
    END
  END FrameData[298]
  PIN FrameData[299]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1405.960 0.930 1406.360 ;
    END
  END FrameData[299]
  PIN FrameData[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 3502.600 0.480 3503.000 ;
    END
  END FrameData[29]
  PIN FrameData[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 3457.240 0.480 3457.640 ;
    END
  END FrameData[2]
  PIN FrameData[300]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1411.000 0.930 1411.400 ;
    END
  END FrameData[300]
  PIN FrameData[301]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1416.040 0.860 1416.440 ;
    END
  END FrameData[301]
  PIN FrameData[302]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1421.080 0.860 1421.480 ;
    END
  END FrameData[302]
  PIN FrameData[303]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1426.120 0.930 1426.520 ;
    END
  END FrameData[303]
  PIN FrameData[304]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1431.160 0.860 1431.560 ;
    END
  END FrameData[304]
  PIN FrameData[305]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1436.200 0.860 1436.600 ;
    END
  END FrameData[305]
  PIN FrameData[306]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1441.240 0.930 1441.640 ;
    END
  END FrameData[306]
  PIN FrameData[307]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1446.280 0.860 1446.680 ;
    END
  END FrameData[307]
  PIN FrameData[308]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1451.320 0.860 1451.720 ;
    END
  END FrameData[308]
  PIN FrameData[309]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1456.360 0.930 1456.760 ;
    END
  END FrameData[309]
  PIN FrameData[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 3504.280 0.480 3504.680 ;
    END
  END FrameData[30]
  PIN FrameData[310]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1461.400 0.860 1461.800 ;
    END
  END FrameData[310]
  PIN FrameData[311]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1466.440 0.860 1466.840 ;
    END
  END FrameData[311]
  PIN FrameData[312]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1471.480 0.930 1471.880 ;
    END
  END FrameData[312]
  PIN FrameData[313]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1476.520 0.860 1476.920 ;
    END
  END FrameData[313]
  PIN FrameData[314]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1481.560 0.860 1481.960 ;
    END
  END FrameData[314]
  PIN FrameData[315]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1486.600 0.930 1487.000 ;
    END
  END FrameData[315]
  PIN FrameData[316]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1491.640 0.860 1492.040 ;
    END
  END FrameData[316]
  PIN FrameData[317]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1496.680 0.860 1497.080 ;
    END
  END FrameData[317]
  PIN FrameData[318]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1501.720 0.930 1502.120 ;
    END
  END FrameData[318]
  PIN FrameData[319]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1506.760 0.930 1507.160 ;
    END
  END FrameData[319]
  PIN FrameData[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 3505.960 0.480 3506.360 ;
    END
  END FrameData[31]
  PIN FrameData[320]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1108.600 0.930 1109.000 ;
    END
  END FrameData[320]
  PIN FrameData[321]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1113.640 0.860 1114.040 ;
    END
  END FrameData[321]
  PIN FrameData[322]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1118.680 0.860 1119.080 ;
    END
  END FrameData[322]
  PIN FrameData[323]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1123.720 0.860 1124.120 ;
    END
  END FrameData[323]
  PIN FrameData[324]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1128.760 0.860 1129.160 ;
    END
  END FrameData[324]
  PIN FrameData[325]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1133.800 0.860 1134.200 ;
    END
  END FrameData[325]
  PIN FrameData[326]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1138.840 0.930 1139.240 ;
    END
  END FrameData[326]
  PIN FrameData[327]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1143.880 0.860 1144.280 ;
    END
  END FrameData[327]
  PIN FrameData[328]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1148.920 0.930 1149.320 ;
    END
  END FrameData[328]
  PIN FrameData[329]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1153.960 0.930 1154.360 ;
    END
  END FrameData[329]
  PIN FrameData[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 3285.880 0.930 3286.280 ;
    END
  END FrameData[32]
  PIN FrameData[330]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1159.000 0.930 1159.400 ;
    END
  END FrameData[330]
  PIN FrameData[331]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1164.040 0.930 1164.440 ;
    END
  END FrameData[331]
  PIN FrameData[332]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1169.080 0.930 1169.480 ;
    END
  END FrameData[332]
  PIN FrameData[333]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1174.120 0.860 1174.520 ;
    END
  END FrameData[333]
  PIN FrameData[334]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1179.160 0.860 1179.560 ;
    END
  END FrameData[334]
  PIN FrameData[335]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1184.200 0.930 1184.600 ;
    END
  END FrameData[335]
  PIN FrameData[336]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1189.240 0.860 1189.640 ;
    END
  END FrameData[336]
  PIN FrameData[337]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1194.280 0.860 1194.680 ;
    END
  END FrameData[337]
  PIN FrameData[338]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1199.320 0.930 1199.720 ;
    END
  END FrameData[338]
  PIN FrameData[339]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1204.360 0.860 1204.760 ;
    END
  END FrameData[339]
  PIN FrameData[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 3290.920 0.860 3291.320 ;
    END
  END FrameData[33]
  PIN FrameData[340]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1209.400 0.860 1209.800 ;
    END
  END FrameData[340]
  PIN FrameData[341]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1214.440 0.930 1214.840 ;
    END
  END FrameData[341]
  PIN FrameData[342]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1219.480 0.860 1219.880 ;
    END
  END FrameData[342]
  PIN FrameData[343]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1224.520 0.860 1224.920 ;
    END
  END FrameData[343]
  PIN FrameData[344]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1229.560 0.930 1229.960 ;
    END
  END FrameData[344]
  PIN FrameData[345]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1234.600 0.860 1235.000 ;
    END
  END FrameData[345]
  PIN FrameData[346]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1239.640 0.860 1240.040 ;
    END
  END FrameData[346]
  PIN FrameData[347]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1244.680 0.930 1245.080 ;
    END
  END FrameData[347]
  PIN FrameData[348]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1249.720 0.860 1250.120 ;
    END
  END FrameData[348]
  PIN FrameData[349]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1254.760 0.860 1255.160 ;
    END
  END FrameData[349]
  PIN FrameData[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 3295.960 0.860 3296.360 ;
    END
  END FrameData[34]
  PIN FrameData[350]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1259.800 0.930 1260.200 ;
    END
  END FrameData[350]
  PIN FrameData[351]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1264.840 0.930 1265.240 ;
    END
  END FrameData[351]
  PIN FrameData[352]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 866.680 0.930 867.080 ;
    END
  END FrameData[352]
  PIN FrameData[353]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 871.720 0.860 872.120 ;
    END
  END FrameData[353]
  PIN FrameData[354]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 876.760 0.860 877.160 ;
    END
  END FrameData[354]
  PIN FrameData[355]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 881.800 0.860 882.200 ;
    END
  END FrameData[355]
  PIN FrameData[356]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 886.840 0.860 887.240 ;
    END
  END FrameData[356]
  PIN FrameData[357]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 891.880 0.860 892.280 ;
    END
  END FrameData[357]
  PIN FrameData[358]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 896.920 0.930 897.320 ;
    END
  END FrameData[358]
  PIN FrameData[359]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 901.960 0.860 902.360 ;
    END
  END FrameData[359]
  PIN FrameData[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 3301.000 0.860 3301.400 ;
    END
  END FrameData[35]
  PIN FrameData[360]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 907.000 0.930 907.400 ;
    END
  END FrameData[360]
  PIN FrameData[361]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 912.040 0.930 912.440 ;
    END
  END FrameData[361]
  PIN FrameData[362]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 917.080 0.930 917.480 ;
    END
  END FrameData[362]
  PIN FrameData[363]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 922.120 0.930 922.520 ;
    END
  END FrameData[363]
  PIN FrameData[364]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 927.160 0.930 927.560 ;
    END
  END FrameData[364]
  PIN FrameData[365]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 932.200 0.860 932.600 ;
    END
  END FrameData[365]
  PIN FrameData[366]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 937.240 0.860 937.640 ;
    END
  END FrameData[366]
  PIN FrameData[367]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 942.280 0.930 942.680 ;
    END
  END FrameData[367]
  PIN FrameData[368]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 947.320 0.860 947.720 ;
    END
  END FrameData[368]
  PIN FrameData[369]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 952.360 0.860 952.760 ;
    END
  END FrameData[369]
  PIN FrameData[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 3306.040 0.860 3306.440 ;
    END
  END FrameData[36]
  PIN FrameData[370]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 957.400 0.930 957.800 ;
    END
  END FrameData[370]
  PIN FrameData[371]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 962.440 0.860 962.840 ;
    END
  END FrameData[371]
  PIN FrameData[372]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 967.480 0.860 967.880 ;
    END
  END FrameData[372]
  PIN FrameData[373]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 972.520 0.930 972.920 ;
    END
  END FrameData[373]
  PIN FrameData[374]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 977.560 0.860 977.960 ;
    END
  END FrameData[374]
  PIN FrameData[375]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 982.600 0.860 983.000 ;
    END
  END FrameData[375]
  PIN FrameData[376]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 987.640 0.930 988.040 ;
    END
  END FrameData[376]
  PIN FrameData[377]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 992.680 0.860 993.080 ;
    END
  END FrameData[377]
  PIN FrameData[378]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 997.720 0.860 998.120 ;
    END
  END FrameData[378]
  PIN FrameData[379]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1002.760 0.930 1003.160 ;
    END
  END FrameData[379]
  PIN FrameData[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 3311.080 0.860 3311.480 ;
    END
  END FrameData[37]
  PIN FrameData[380]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1007.800 0.860 1008.200 ;
    END
  END FrameData[380]
  PIN FrameData[381]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1012.840 0.860 1013.240 ;
    END
  END FrameData[381]
  PIN FrameData[382]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1017.880 0.930 1018.280 ;
    END
  END FrameData[382]
  PIN FrameData[383]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1022.920 0.930 1023.320 ;
    END
  END FrameData[383]
  PIN FrameData[384]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 624.760 0.930 625.160 ;
    END
  END FrameData[384]
  PIN FrameData[385]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 629.800 0.860 630.200 ;
    END
  END FrameData[385]
  PIN FrameData[386]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 634.840 0.860 635.240 ;
    END
  END FrameData[386]
  PIN FrameData[387]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 639.880 0.860 640.280 ;
    END
  END FrameData[387]
  PIN FrameData[388]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 644.920 0.860 645.320 ;
    END
  END FrameData[388]
  PIN FrameData[389]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 649.960 0.860 650.360 ;
    END
  END FrameData[389]
  PIN FrameData[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 3316.120 0.930 3316.520 ;
    END
  END FrameData[38]
  PIN FrameData[390]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 655.000 0.930 655.400 ;
    END
  END FrameData[390]
  PIN FrameData[391]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 660.040 0.860 660.440 ;
    END
  END FrameData[391]
  PIN FrameData[392]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 665.080 0.930 665.480 ;
    END
  END FrameData[392]
  PIN FrameData[393]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 670.120 0.930 670.520 ;
    END
  END FrameData[393]
  PIN FrameData[394]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 675.160 0.930 675.560 ;
    END
  END FrameData[394]
  PIN FrameData[395]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 680.200 0.930 680.600 ;
    END
  END FrameData[395]
  PIN FrameData[396]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 685.240 0.930 685.640 ;
    END
  END FrameData[396]
  PIN FrameData[397]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 690.280 0.860 690.680 ;
    END
  END FrameData[397]
  PIN FrameData[398]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 695.320 0.860 695.720 ;
    END
  END FrameData[398]
  PIN FrameData[399]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 700.360 0.930 700.760 ;
    END
  END FrameData[399]
  PIN FrameData[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 3321.160 0.860 3321.560 ;
    END
  END FrameData[39]
  PIN FrameData[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 3458.920 0.480 3459.320 ;
    END
  END FrameData[3]
  PIN FrameData[400]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 705.400 0.860 705.800 ;
    END
  END FrameData[400]
  PIN FrameData[401]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 710.440 0.860 710.840 ;
    END
  END FrameData[401]
  PIN FrameData[402]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 715.480 0.930 715.880 ;
    END
  END FrameData[402]
  PIN FrameData[403]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 720.520 0.860 720.920 ;
    END
  END FrameData[403]
  PIN FrameData[404]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 725.560 0.860 725.960 ;
    END
  END FrameData[404]
  PIN FrameData[405]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 730.600 0.930 731.000 ;
    END
  END FrameData[405]
  PIN FrameData[406]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 735.640 0.860 736.040 ;
    END
  END FrameData[406]
  PIN FrameData[407]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 740.680 0.860 741.080 ;
    END
  END FrameData[407]
  PIN FrameData[408]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 745.720 0.930 746.120 ;
    END
  END FrameData[408]
  PIN FrameData[409]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 750.760 0.860 751.160 ;
    END
  END FrameData[409]
  PIN FrameData[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 3326.200 0.930 3326.600 ;
    END
  END FrameData[40]
  PIN FrameData[410]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 755.800 0.860 756.200 ;
    END
  END FrameData[410]
  PIN FrameData[411]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 760.840 0.930 761.240 ;
    END
  END FrameData[411]
  PIN FrameData[412]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 765.880 0.860 766.280 ;
    END
  END FrameData[412]
  PIN FrameData[413]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 770.920 0.860 771.320 ;
    END
  END FrameData[413]
  PIN FrameData[414]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 775.960 0.930 776.360 ;
    END
  END FrameData[414]
  PIN FrameData[415]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 781.000 0.930 781.400 ;
    END
  END FrameData[415]
  PIN FrameData[416]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 382.840 0.930 383.240 ;
    END
  END FrameData[416]
  PIN FrameData[417]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 387.880 0.860 388.280 ;
    END
  END FrameData[417]
  PIN FrameData[418]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 392.920 0.860 393.320 ;
    END
  END FrameData[418]
  PIN FrameData[419]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 397.960 0.860 398.360 ;
    END
  END FrameData[419]
  PIN FrameData[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 3331.240 0.930 3331.640 ;
    END
  END FrameData[41]
  PIN FrameData[420]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 403.000 0.860 403.400 ;
    END
  END FrameData[420]
  PIN FrameData[421]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 408.040 0.860 408.440 ;
    END
  END FrameData[421]
  PIN FrameData[422]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 413.080 0.930 413.480 ;
    END
  END FrameData[422]
  PIN FrameData[423]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 418.120 0.860 418.520 ;
    END
  END FrameData[423]
  PIN FrameData[424]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 423.160 0.930 423.560 ;
    END
  END FrameData[424]
  PIN FrameData[425]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 428.200 0.930 428.600 ;
    END
  END FrameData[425]
  PIN FrameData[426]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 433.240 0.930 433.640 ;
    END
  END FrameData[426]
  PIN FrameData[427]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 438.280 0.930 438.680 ;
    END
  END FrameData[427]
  PIN FrameData[428]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 443.320 0.930 443.720 ;
    END
  END FrameData[428]
  PIN FrameData[429]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 448.360 0.860 448.760 ;
    END
  END FrameData[429]
  PIN FrameData[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 3336.280 0.930 3336.680 ;
    END
  END FrameData[42]
  PIN FrameData[430]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 453.400 0.860 453.800 ;
    END
  END FrameData[430]
  PIN FrameData[431]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 458.440 0.930 458.840 ;
    END
  END FrameData[431]
  PIN FrameData[432]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 463.480 0.860 463.880 ;
    END
  END FrameData[432]
  PIN FrameData[433]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 468.520 0.860 468.920 ;
    END
  END FrameData[433]
  PIN FrameData[434]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 473.560 0.930 473.960 ;
    END
  END FrameData[434]
  PIN FrameData[435]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 478.600 0.860 479.000 ;
    END
  END FrameData[435]
  PIN FrameData[436]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 483.640 0.860 484.040 ;
    END
  END FrameData[436]
  PIN FrameData[437]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 488.680 0.930 489.080 ;
    END
  END FrameData[437]
  PIN FrameData[438]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 493.720 0.860 494.120 ;
    END
  END FrameData[438]
  PIN FrameData[439]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 498.760 0.860 499.160 ;
    END
  END FrameData[439]
  PIN FrameData[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 3341.320 0.930 3341.720 ;
    END
  END FrameData[43]
  PIN FrameData[440]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 503.800 0.930 504.200 ;
    END
  END FrameData[440]
  PIN FrameData[441]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 508.840 0.860 509.240 ;
    END
  END FrameData[441]
  PIN FrameData[442]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 513.880 0.860 514.280 ;
    END
  END FrameData[442]
  PIN FrameData[443]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 518.920 0.930 519.320 ;
    END
  END FrameData[443]
  PIN FrameData[444]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 523.960 0.860 524.360 ;
    END
  END FrameData[444]
  PIN FrameData[445]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 529.000 0.860 529.400 ;
    END
  END FrameData[445]
  PIN FrameData[446]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 534.040 0.930 534.440 ;
    END
  END FrameData[446]
  PIN FrameData[447]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 539.080 0.930 539.480 ;
    END
  END FrameData[447]
  PIN FrameData[448]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 140.920 0.930 141.320 ;
    END
  END FrameData[448]
  PIN FrameData[449]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 145.960 0.860 146.360 ;
    END
  END FrameData[449]
  PIN FrameData[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 3346.360 0.930 3346.760 ;
    END
  END FrameData[44]
  PIN FrameData[450]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 151.000 0.860 151.400 ;
    END
  END FrameData[450]
  PIN FrameData[451]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 156.040 0.860 156.440 ;
    END
  END FrameData[451]
  PIN FrameData[452]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 161.080 0.860 161.480 ;
    END
  END FrameData[452]
  PIN FrameData[453]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 166.120 0.860 166.520 ;
    END
  END FrameData[453]
  PIN FrameData[454]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 171.160 0.930 171.560 ;
    END
  END FrameData[454]
  PIN FrameData[455]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 176.200 0.860 176.600 ;
    END
  END FrameData[455]
  PIN FrameData[456]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 181.240 0.930 181.640 ;
    END
  END FrameData[456]
  PIN FrameData[457]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 186.280 0.930 186.680 ;
    END
  END FrameData[457]
  PIN FrameData[458]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 191.320 0.930 191.720 ;
    END
  END FrameData[458]
  PIN FrameData[459]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 196.360 0.930 196.760 ;
    END
  END FrameData[459]
  PIN FrameData[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 3351.400 0.860 3351.800 ;
    END
  END FrameData[45]
  PIN FrameData[460]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 201.400 0.930 201.800 ;
    END
  END FrameData[460]
  PIN FrameData[461]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 206.440 0.860 206.840 ;
    END
  END FrameData[461]
  PIN FrameData[462]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 211.480 0.860 211.880 ;
    END
  END FrameData[462]
  PIN FrameData[463]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 216.520 0.930 216.920 ;
    END
  END FrameData[463]
  PIN FrameData[464]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 221.560 0.860 221.960 ;
    END
  END FrameData[464]
  PIN FrameData[465]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 226.600 0.860 227.000 ;
    END
  END FrameData[465]
  PIN FrameData[466]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 231.640 0.930 232.040 ;
    END
  END FrameData[466]
  PIN FrameData[467]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 236.680 0.860 237.080 ;
    END
  END FrameData[467]
  PIN FrameData[468]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 241.720 0.860 242.120 ;
    END
  END FrameData[468]
  PIN FrameData[469]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 246.760 0.930 247.160 ;
    END
  END FrameData[469]
  PIN FrameData[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 3356.440 0.860 3356.840 ;
    END
  END FrameData[46]
  PIN FrameData[470]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 251.800 0.860 252.200 ;
    END
  END FrameData[470]
  PIN FrameData[471]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 256.840 0.860 257.240 ;
    END
  END FrameData[471]
  PIN FrameData[472]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 261.880 0.930 262.280 ;
    END
  END FrameData[472]
  PIN FrameData[473]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 266.920 0.860 267.320 ;
    END
  END FrameData[473]
  PIN FrameData[474]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 271.960 0.860 272.360 ;
    END
  END FrameData[474]
  PIN FrameData[475]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 277.000 0.930 277.400 ;
    END
  END FrameData[475]
  PIN FrameData[476]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 282.040 0.860 282.440 ;
    END
  END FrameData[476]
  PIN FrameData[477]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 287.080 0.860 287.480 ;
    END
  END FrameData[477]
  PIN FrameData[478]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 292.120 0.930 292.520 ;
    END
  END FrameData[478]
  PIN FrameData[479]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 297.160 0.930 297.560 ;
    END
  END FrameData[479]
  PIN FrameData[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 3361.480 0.930 3361.880 ;
    END
  END FrameData[47]
  PIN FrameData[480]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 6.940 0.480 7.340 ;
    END
  END FrameData[480]
  PIN FrameData[481]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 8.620 0.480 9.020 ;
    END
  END FrameData[481]
  PIN FrameData[482]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 10.300 0.480 10.700 ;
    END
  END FrameData[482]
  PIN FrameData[483]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 11.980 0.480 12.380 ;
    END
  END FrameData[483]
  PIN FrameData[484]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 13.660 0.480 14.060 ;
    END
  END FrameData[484]
  PIN FrameData[485]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 15.340 0.480 15.740 ;
    END
  END FrameData[485]
  PIN FrameData[486]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 17.020 0.480 17.420 ;
    END
  END FrameData[486]
  PIN FrameData[487]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 18.700 0.480 19.100 ;
    END
  END FrameData[487]
  PIN FrameData[488]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 20.380 0.480 20.780 ;
    END
  END FrameData[488]
  PIN FrameData[489]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 22.060 0.480 22.460 ;
    END
  END FrameData[489]
  PIN FrameData[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 3366.520 0.860 3366.920 ;
    END
  END FrameData[48]
  PIN FrameData[490]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 23.740 0.480 24.140 ;
    END
  END FrameData[490]
  PIN FrameData[491]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 25.420 0.480 25.820 ;
    END
  END FrameData[491]
  PIN FrameData[492]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 27.100 0.480 27.500 ;
    END
  END FrameData[492]
  PIN FrameData[493]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 28.780 0.480 29.180 ;
    END
  END FrameData[493]
  PIN FrameData[494]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 30.460 0.480 30.860 ;
    END
  END FrameData[494]
  PIN FrameData[495]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 32.140 0.480 32.540 ;
    END
  END FrameData[495]
  PIN FrameData[496]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.397500 ;
    ANTENNADIFFAREA 4.030800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 33.820 0.480 34.220 ;
    END
  END FrameData[496]
  PIN FrameData[497]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 35.500 0.480 35.900 ;
    END
  END FrameData[497]
  PIN FrameData[498]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 37.180 0.480 37.580 ;
    END
  END FrameData[498]
  PIN FrameData[499]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 38.860 0.480 39.260 ;
    END
  END FrameData[499]
  PIN FrameData[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 3371.560 0.860 3371.960 ;
    END
  END FrameData[49]
  PIN FrameData[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 3460.600 0.480 3461.000 ;
    END
  END FrameData[4]
  PIN FrameData[500]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 40.540 0.480 40.940 ;
    END
  END FrameData[500]
  PIN FrameData[501]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.397500 ;
    ANTENNADIFFAREA 4.030800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 42.220 0.480 42.620 ;
    END
  END FrameData[501]
  PIN FrameData[502]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 43.900 0.480 44.300 ;
    END
  END FrameData[502]
  PIN FrameData[503]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 45.580 0.480 45.980 ;
    END
  END FrameData[503]
  PIN FrameData[504]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 6.264700 ;
    ANTENNADIFFAREA 20.153999 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 47.260 0.480 47.660 ;
    END
  END FrameData[504]
  PIN FrameData[505]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 6.264700 ;
    ANTENNADIFFAREA 20.153999 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 48.940 0.480 49.340 ;
    END
  END FrameData[505]
  PIN FrameData[506]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 6.264700 ;
    ANTENNADIFFAREA 20.153999 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 50.620 0.480 51.020 ;
    END
  END FrameData[506]
  PIN FrameData[507]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 5.656300 ;
    ANTENNADIFFAREA 18.138599 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 52.300 0.480 52.700 ;
    END
  END FrameData[507]
  PIN FrameData[508]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 53.980 0.480 54.380 ;
    END
  END FrameData[508]
  PIN FrameData[509]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.397500 ;
    ANTENNADIFFAREA 4.030800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 55.660 0.480 56.060 ;
    END
  END FrameData[509]
  PIN FrameData[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 3376.600 0.930 3377.000 ;
    END
  END FrameData[50]
  PIN FrameData[510]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 57.340 0.480 57.740 ;
    END
  END FrameData[510]
  PIN FrameData[511]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 59.020 0.480 59.420 ;
    END
  END FrameData[511]
  PIN FrameData[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 3381.640 0.860 3382.040 ;
    END
  END FrameData[51]
  PIN FrameData[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 3386.680 0.860 3387.080 ;
    END
  END FrameData[52]
  PIN FrameData[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 3391.720 0.930 3392.120 ;
    END
  END FrameData[53]
  PIN FrameData[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 3396.760 0.860 3397.160 ;
    END
  END FrameData[54]
  PIN FrameData[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 3401.800 0.860 3402.200 ;
    END
  END FrameData[55]
  PIN FrameData[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 3406.840 0.930 3407.240 ;
    END
  END FrameData[56]
  PIN FrameData[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 3411.880 0.860 3412.280 ;
    END
  END FrameData[57]
  PIN FrameData[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 3416.920 0.860 3417.320 ;
    END
  END FrameData[58]
  PIN FrameData[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 3421.960 0.930 3422.360 ;
    END
  END FrameData[59]
  PIN FrameData[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 3462.280 0.480 3462.680 ;
    END
  END FrameData[5]
  PIN FrameData[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 3427.000 0.860 3427.400 ;
    END
  END FrameData[60]
  PIN FrameData[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 3432.040 0.860 3432.440 ;
    END
  END FrameData[61]
  PIN FrameData[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 3437.080 0.930 3437.480 ;
    END
  END FrameData[62]
  PIN FrameData[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 3442.120 0.930 3442.520 ;
    END
  END FrameData[63]
  PIN FrameData[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 3043.960 0.930 3044.360 ;
    END
  END FrameData[64]
  PIN FrameData[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 3049.000 0.860 3049.400 ;
    END
  END FrameData[65]
  PIN FrameData[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 3054.040 0.860 3054.440 ;
    END
  END FrameData[66]
  PIN FrameData[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 3059.080 0.860 3059.480 ;
    END
  END FrameData[67]
  PIN FrameData[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 3064.120 0.860 3064.520 ;
    END
  END FrameData[68]
  PIN FrameData[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 3069.160 0.860 3069.560 ;
    END
  END FrameData[69]
  PIN FrameData[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 3463.960 0.480 3464.360 ;
    END
  END FrameData[6]
  PIN FrameData[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 3074.200 0.930 3074.600 ;
    END
  END FrameData[70]
  PIN FrameData[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 3079.240 0.860 3079.640 ;
    END
  END FrameData[71]
  PIN FrameData[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 3084.280 0.930 3084.680 ;
    END
  END FrameData[72]
  PIN FrameData[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 3089.320 0.930 3089.720 ;
    END
  END FrameData[73]
  PIN FrameData[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 3094.360 0.930 3094.760 ;
    END
  END FrameData[74]
  PIN FrameData[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 3099.400 0.930 3099.800 ;
    END
  END FrameData[75]
  PIN FrameData[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 3104.440 0.930 3104.840 ;
    END
  END FrameData[76]
  PIN FrameData[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 3109.480 0.860 3109.880 ;
    END
  END FrameData[77]
  PIN FrameData[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 3114.520 0.860 3114.920 ;
    END
  END FrameData[78]
  PIN FrameData[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 3119.560 0.930 3119.960 ;
    END
  END FrameData[79]
  PIN FrameData[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 3465.640 0.480 3466.040 ;
    END
  END FrameData[7]
  PIN FrameData[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 3124.600 0.860 3125.000 ;
    END
  END FrameData[80]
  PIN FrameData[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 3129.640 0.860 3130.040 ;
    END
  END FrameData[81]
  PIN FrameData[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 3134.680 0.930 3135.080 ;
    END
  END FrameData[82]
  PIN FrameData[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 3139.720 0.860 3140.120 ;
    END
  END FrameData[83]
  PIN FrameData[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 3144.760 0.860 3145.160 ;
    END
  END FrameData[84]
  PIN FrameData[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 3149.800 0.930 3150.200 ;
    END
  END FrameData[85]
  PIN FrameData[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 3154.840 0.860 3155.240 ;
    END
  END FrameData[86]
  PIN FrameData[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 3159.880 0.860 3160.280 ;
    END
  END FrameData[87]
  PIN FrameData[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 3164.920 0.930 3165.320 ;
    END
  END FrameData[88]
  PIN FrameData[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 3169.960 0.860 3170.360 ;
    END
  END FrameData[89]
  PIN FrameData[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 3467.320 0.480 3467.720 ;
    END
  END FrameData[8]
  PIN FrameData[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 3175.000 0.860 3175.400 ;
    END
  END FrameData[90]
  PIN FrameData[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 3180.040 0.930 3180.440 ;
    END
  END FrameData[91]
  PIN FrameData[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 3185.080 0.860 3185.480 ;
    END
  END FrameData[92]
  PIN FrameData[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 3190.120 0.860 3190.520 ;
    END
  END FrameData[93]
  PIN FrameData[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 3195.160 0.930 3195.560 ;
    END
  END FrameData[94]
  PIN FrameData[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 3200.200 0.930 3200.600 ;
    END
  END FrameData[95]
  PIN FrameData[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2802.040 0.930 2802.440 ;
    END
  END FrameData[96]
  PIN FrameData[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2807.080 0.860 2807.480 ;
    END
  END FrameData[97]
  PIN FrameData[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2812.120 0.860 2812.520 ;
    END
  END FrameData[98]
  PIN FrameData[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2817.160 0.860 2817.560 ;
    END
  END FrameData[99]
  PIN FrameData[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 3469.000 0.480 3469.400 ;
    END
  END FrameData[9]
  PIN FrameStrobe[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 8.440 0.000 8.840 0.400 ;
    END
  END FrameStrobe[0]
  PIN FrameStrobe[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1173.400 0.000 1173.800 0.480 ;
    END
  END FrameStrobe[100]
  PIN FrameStrobe[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1177.240 0.000 1177.640 0.480 ;
    END
  END FrameStrobe[101]
  PIN FrameStrobe[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1181.080 0.000 1181.480 0.480 ;
    END
  END FrameStrobe[102]
  PIN FrameStrobe[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1184.920 0.000 1185.320 0.480 ;
    END
  END FrameStrobe[103]
  PIN FrameStrobe[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1188.760 0.000 1189.160 0.480 ;
    END
  END FrameStrobe[104]
  PIN FrameStrobe[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1192.600 0.000 1193.000 0.480 ;
    END
  END FrameStrobe[105]
  PIN FrameStrobe[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1196.440 0.000 1196.840 0.480 ;
    END
  END FrameStrobe[106]
  PIN FrameStrobe[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1200.280 0.000 1200.680 0.480 ;
    END
  END FrameStrobe[107]
  PIN FrameStrobe[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1204.120 0.000 1204.520 0.480 ;
    END
  END FrameStrobe[108]
  PIN FrameStrobe[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1207.960 0.000 1208.360 0.480 ;
    END
  END FrameStrobe[109]
  PIN FrameStrobe[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 37.240 0.000 37.640 0.400 ;
    END
  END FrameStrobe[10]
  PIN FrameStrobe[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1211.800 0.000 1212.200 0.480 ;
    END
  END FrameStrobe[110]
  PIN FrameStrobe[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1215.640 0.000 1216.040 0.480 ;
    END
  END FrameStrobe[111]
  PIN FrameStrobe[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1219.480 0.000 1219.880 0.480 ;
    END
  END FrameStrobe[112]
  PIN FrameStrobe[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1223.320 0.000 1223.720 0.480 ;
    END
  END FrameStrobe[113]
  PIN FrameStrobe[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1227.160 0.000 1227.560 0.480 ;
    END
  END FrameStrobe[114]
  PIN FrameStrobe[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1231.000 0.000 1231.400 0.480 ;
    END
  END FrameStrobe[115]
  PIN FrameStrobe[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1234.840 0.000 1235.240 0.480 ;
    END
  END FrameStrobe[116]
  PIN FrameStrobe[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1238.680 0.000 1239.080 0.480 ;
    END
  END FrameStrobe[117]
  PIN FrameStrobe[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1242.520 0.000 1242.920 0.480 ;
    END
  END FrameStrobe[118]
  PIN FrameStrobe[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1246.360 0.000 1246.760 0.480 ;
    END
  END FrameStrobe[119]
  PIN FrameStrobe[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 40.120 0.000 40.520 0.400 ;
    END
  END FrameStrobe[11]
  PIN FrameStrobe[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1405.240 0.000 1405.640 0.480 ;
    END
  END FrameStrobe[120]
  PIN FrameStrobe[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1409.080 0.000 1409.480 0.480 ;
    END
  END FrameStrobe[121]
  PIN FrameStrobe[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1412.920 0.000 1413.320 0.480 ;
    END
  END FrameStrobe[122]
  PIN FrameStrobe[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1416.760 0.000 1417.160 0.480 ;
    END
  END FrameStrobe[123]
  PIN FrameStrobe[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1420.600 0.000 1421.000 0.480 ;
    END
  END FrameStrobe[124]
  PIN FrameStrobe[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1424.440 0.000 1424.840 0.480 ;
    END
  END FrameStrobe[125]
  PIN FrameStrobe[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1428.280 0.000 1428.680 0.480 ;
    END
  END FrameStrobe[126]
  PIN FrameStrobe[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1432.120 0.000 1432.520 0.480 ;
    END
  END FrameStrobe[127]
  PIN FrameStrobe[128]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1435.960 0.000 1436.360 0.480 ;
    END
  END FrameStrobe[128]
  PIN FrameStrobe[129]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1439.800 0.000 1440.200 0.480 ;
    END
  END FrameStrobe[129]
  PIN FrameStrobe[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 43.000 0.000 43.400 0.400 ;
    END
  END FrameStrobe[12]
  PIN FrameStrobe[130]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1443.640 0.000 1444.040 0.480 ;
    END
  END FrameStrobe[130]
  PIN FrameStrobe[131]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1447.480 0.000 1447.880 0.480 ;
    END
  END FrameStrobe[131]
  PIN FrameStrobe[132]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1451.320 0.000 1451.720 0.480 ;
    END
  END FrameStrobe[132]
  PIN FrameStrobe[133]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1455.160 0.000 1455.560 0.480 ;
    END
  END FrameStrobe[133]
  PIN FrameStrobe[134]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1459.000 0.000 1459.400 0.480 ;
    END
  END FrameStrobe[134]
  PIN FrameStrobe[135]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1462.840 0.000 1463.240 0.480 ;
    END
  END FrameStrobe[135]
  PIN FrameStrobe[136]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1466.680 0.000 1467.080 0.480 ;
    END
  END FrameStrobe[136]
  PIN FrameStrobe[137]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1470.520 0.000 1470.920 0.480 ;
    END
  END FrameStrobe[137]
  PIN FrameStrobe[138]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1474.360 0.000 1474.760 0.480 ;
    END
  END FrameStrobe[138]
  PIN FrameStrobe[139]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1478.200 0.000 1478.600 0.480 ;
    END
  END FrameStrobe[139]
  PIN FrameStrobe[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 45.880 0.000 46.280 0.400 ;
    END
  END FrameStrobe[13]
  PIN FrameStrobe[140]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1514.200 0.000 1514.600 0.480 ;
    END
  END FrameStrobe[140]
  PIN FrameStrobe[141]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1522.840 0.000 1523.240 0.480 ;
    END
  END FrameStrobe[141]
  PIN FrameStrobe[142]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1531.480 0.000 1531.880 0.480 ;
    END
  END FrameStrobe[142]
  PIN FrameStrobe[143]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1540.120 0.000 1540.520 0.480 ;
    END
  END FrameStrobe[143]
  PIN FrameStrobe[144]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1548.760 0.000 1549.160 0.480 ;
    END
  END FrameStrobe[144]
  PIN FrameStrobe[145]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1557.400 0.000 1557.800 0.480 ;
    END
  END FrameStrobe[145]
  PIN FrameStrobe[146]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1566.040 0.000 1566.440 0.480 ;
    END
  END FrameStrobe[146]
  PIN FrameStrobe[147]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1574.680 0.000 1575.080 0.480 ;
    END
  END FrameStrobe[147]
  PIN FrameStrobe[148]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1583.320 0.000 1583.720 0.480 ;
    END
  END FrameStrobe[148]
  PIN FrameStrobe[149]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1591.960 0.000 1592.360 0.480 ;
    END
  END FrameStrobe[149]
  PIN FrameStrobe[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 48.760 0.000 49.160 0.400 ;
    END
  END FrameStrobe[14]
  PIN FrameStrobe[150]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1600.600 0.000 1601.000 0.480 ;
    END
  END FrameStrobe[150]
  PIN FrameStrobe[151]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1609.240 0.000 1609.640 0.480 ;
    END
  END FrameStrobe[151]
  PIN FrameStrobe[152]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1617.880 0.000 1618.280 0.480 ;
    END
  END FrameStrobe[152]
  PIN FrameStrobe[153]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1626.520 0.000 1626.920 0.480 ;
    END
  END FrameStrobe[153]
  PIN FrameStrobe[154]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1635.160 0.000 1635.560 0.480 ;
    END
  END FrameStrobe[154]
  PIN FrameStrobe[155]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1643.800 0.000 1644.200 0.480 ;
    END
  END FrameStrobe[155]
  PIN FrameStrobe[156]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1652.440 0.000 1652.840 0.480 ;
    END
  END FrameStrobe[156]
  PIN FrameStrobe[157]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1661.080 0.000 1661.480 0.480 ;
    END
  END FrameStrobe[157]
  PIN FrameStrobe[158]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1669.720 0.000 1670.120 0.480 ;
    END
  END FrameStrobe[158]
  PIN FrameStrobe[159]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1678.360 0.000 1678.760 0.480 ;
    END
  END FrameStrobe[159]
  PIN FrameStrobe[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 51.640 0.000 52.040 0.400 ;
    END
  END FrameStrobe[15]
  PIN FrameStrobe[160]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1833.400 0.000 1833.800 0.480 ;
    END
  END FrameStrobe[160]
  PIN FrameStrobe[161]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1837.240 0.000 1837.640 0.480 ;
    END
  END FrameStrobe[161]
  PIN FrameStrobe[162]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1841.080 0.000 1841.480 0.480 ;
    END
  END FrameStrobe[162]
  PIN FrameStrobe[163]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1844.920 0.000 1845.320 0.480 ;
    END
  END FrameStrobe[163]
  PIN FrameStrobe[164]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1848.760 0.000 1849.160 0.480 ;
    END
  END FrameStrobe[164]
  PIN FrameStrobe[165]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1852.600 0.000 1853.000 0.480 ;
    END
  END FrameStrobe[165]
  PIN FrameStrobe[166]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1856.440 0.000 1856.840 0.480 ;
    END
  END FrameStrobe[166]
  PIN FrameStrobe[167]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1860.280 0.000 1860.680 0.480 ;
    END
  END FrameStrobe[167]
  PIN FrameStrobe[168]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1864.120 0.000 1864.520 0.480 ;
    END
  END FrameStrobe[168]
  PIN FrameStrobe[169]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1867.960 0.000 1868.360 0.480 ;
    END
  END FrameStrobe[169]
  PIN FrameStrobe[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 54.520 0.000 54.920 0.400 ;
    END
  END FrameStrobe[16]
  PIN FrameStrobe[170]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1871.800 0.000 1872.200 0.480 ;
    END
  END FrameStrobe[170]
  PIN FrameStrobe[171]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1875.640 0.000 1876.040 0.480 ;
    END
  END FrameStrobe[171]
  PIN FrameStrobe[172]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1879.480 0.000 1879.880 0.480 ;
    END
  END FrameStrobe[172]
  PIN FrameStrobe[173]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1883.320 0.000 1883.720 0.480 ;
    END
  END FrameStrobe[173]
  PIN FrameStrobe[174]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1887.160 0.000 1887.560 0.480 ;
    END
  END FrameStrobe[174]
  PIN FrameStrobe[175]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1891.000 0.000 1891.400 0.480 ;
    END
  END FrameStrobe[175]
  PIN FrameStrobe[176]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1894.840 0.000 1895.240 0.480 ;
    END
  END FrameStrobe[176]
  PIN FrameStrobe[177]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1898.680 0.000 1899.080 0.480 ;
    END
  END FrameStrobe[177]
  PIN FrameStrobe[178]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1902.520 0.000 1902.920 0.480 ;
    END
  END FrameStrobe[178]
  PIN FrameStrobe[179]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1906.360 0.000 1906.760 0.480 ;
    END
  END FrameStrobe[179]
  PIN FrameStrobe[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 57.400 0.000 57.800 0.400 ;
    END
  END FrameStrobe[17]
  PIN FrameStrobe[180]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 2065.240 0.000 2065.640 0.480 ;
    END
  END FrameStrobe[180]
  PIN FrameStrobe[181]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 2069.080 0.000 2069.480 0.480 ;
    END
  END FrameStrobe[181]
  PIN FrameStrobe[182]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 2072.920 0.000 2073.320 0.480 ;
    END
  END FrameStrobe[182]
  PIN FrameStrobe[183]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 2076.760 0.000 2077.160 0.480 ;
    END
  END FrameStrobe[183]
  PIN FrameStrobe[184]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 2080.600 0.000 2081.000 0.480 ;
    END
  END FrameStrobe[184]
  PIN FrameStrobe[185]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 2084.440 0.000 2084.840 0.480 ;
    END
  END FrameStrobe[185]
  PIN FrameStrobe[186]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 2088.280 0.000 2088.680 0.480 ;
    END
  END FrameStrobe[186]
  PIN FrameStrobe[187]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 2092.120 0.000 2092.520 0.480 ;
    END
  END FrameStrobe[187]
  PIN FrameStrobe[188]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 2095.960 0.000 2096.360 0.480 ;
    END
  END FrameStrobe[188]
  PIN FrameStrobe[189]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 2099.800 0.000 2100.200 0.480 ;
    END
  END FrameStrobe[189]
  PIN FrameStrobe[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 60.280 0.000 60.680 0.400 ;
    END
  END FrameStrobe[18]
  PIN FrameStrobe[190]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 2103.640 0.000 2104.040 0.480 ;
    END
  END FrameStrobe[190]
  PIN FrameStrobe[191]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 2107.480 0.000 2107.880 0.480 ;
    END
  END FrameStrobe[191]
  PIN FrameStrobe[192]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 2111.320 0.000 2111.720 0.480 ;
    END
  END FrameStrobe[192]
  PIN FrameStrobe[193]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 2115.160 0.000 2115.560 0.480 ;
    END
  END FrameStrobe[193]
  PIN FrameStrobe[194]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 2119.000 0.000 2119.400 0.480 ;
    END
  END FrameStrobe[194]
  PIN FrameStrobe[195]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 2122.840 0.000 2123.240 0.480 ;
    END
  END FrameStrobe[195]
  PIN FrameStrobe[196]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 2126.680 0.000 2127.080 0.480 ;
    END
  END FrameStrobe[196]
  PIN FrameStrobe[197]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 2130.520 0.000 2130.920 0.480 ;
    END
  END FrameStrobe[197]
  PIN FrameStrobe[198]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 2134.360 0.000 2134.760 0.480 ;
    END
  END FrameStrobe[198]
  PIN FrameStrobe[199]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 2138.200 0.000 2138.600 0.480 ;
    END
  END FrameStrobe[199]
  PIN FrameStrobe[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 63.160 0.000 63.560 0.400 ;
    END
  END FrameStrobe[19]
  PIN FrameStrobe[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 11.320 0.000 11.720 0.400 ;
    END
  END FrameStrobe[1]
  PIN FrameStrobe[200]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 2164.600 0.000 2165.000 0.400 ;
    END
  END FrameStrobe[200]
  PIN FrameStrobe[201]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 2169.400 0.000 2169.800 0.400 ;
    END
  END FrameStrobe[201]
  PIN FrameStrobe[202]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 2174.200 0.000 2174.600 0.400 ;
    END
  END FrameStrobe[202]
  PIN FrameStrobe[203]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 2179.000 0.000 2179.400 0.400 ;
    END
  END FrameStrobe[203]
  PIN FrameStrobe[204]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 2183.800 0.000 2184.200 0.400 ;
    END
  END FrameStrobe[204]
  PIN FrameStrobe[205]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 2188.600 0.000 2189.000 0.400 ;
    END
  END FrameStrobe[205]
  PIN FrameStrobe[206]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 2193.400 0.000 2193.800 0.400 ;
    END
  END FrameStrobe[206]
  PIN FrameStrobe[207]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 2198.200 0.000 2198.600 0.400 ;
    END
  END FrameStrobe[207]
  PIN FrameStrobe[208]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 2203.000 0.000 2203.400 0.400 ;
    END
  END FrameStrobe[208]
  PIN FrameStrobe[209]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 2207.800 0.000 2208.200 0.400 ;
    END
  END FrameStrobe[209]
  PIN FrameStrobe[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 89.560 0.000 89.960 0.480 ;
    END
  END FrameStrobe[20]
  PIN FrameStrobe[210]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 2212.600 0.000 2213.000 0.400 ;
    END
  END FrameStrobe[210]
  PIN FrameStrobe[211]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 2217.400 0.000 2217.800 0.400 ;
    END
  END FrameStrobe[211]
  PIN FrameStrobe[212]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 2222.200 0.000 2222.600 0.400 ;
    END
  END FrameStrobe[212]
  PIN FrameStrobe[213]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 2227.000 0.000 2227.400 0.400 ;
    END
  END FrameStrobe[213]
  PIN FrameStrobe[214]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 2231.800 0.000 2232.200 0.400 ;
    END
  END FrameStrobe[214]
  PIN FrameStrobe[215]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 2236.600 0.000 2237.000 0.400 ;
    END
  END FrameStrobe[215]
  PIN FrameStrobe[216]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 2241.400 0.000 2241.800 0.400 ;
    END
  END FrameStrobe[216]
  PIN FrameStrobe[217]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 2246.200 0.000 2246.600 0.400 ;
    END
  END FrameStrobe[217]
  PIN FrameStrobe[218]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 2251.000 0.000 2251.400 0.400 ;
    END
  END FrameStrobe[218]
  PIN FrameStrobe[219]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 2255.800 0.000 2256.200 0.400 ;
    END
  END FrameStrobe[219]
  PIN FrameStrobe[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 100.120 0.000 100.520 0.480 ;
    END
  END FrameStrobe[21]
  PIN FrameStrobe[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 110.680 0.000 111.080 0.480 ;
    END
  END FrameStrobe[22]
  PIN FrameStrobe[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 121.240 0.000 121.640 0.480 ;
    END
  END FrameStrobe[23]
  PIN FrameStrobe[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 131.800 0.000 132.200 0.480 ;
    END
  END FrameStrobe[24]
  PIN FrameStrobe[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 142.360 0.000 142.760 0.480 ;
    END
  END FrameStrobe[25]
  PIN FrameStrobe[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 152.920 0.000 153.320 0.480 ;
    END
  END FrameStrobe[26]
  PIN FrameStrobe[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 163.480 0.000 163.880 0.480 ;
    END
  END FrameStrobe[27]
  PIN FrameStrobe[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 174.040 0.000 174.440 0.480 ;
    END
  END FrameStrobe[28]
  PIN FrameStrobe[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 184.600 0.000 185.000 0.480 ;
    END
  END FrameStrobe[29]
  PIN FrameStrobe[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 14.200 0.000 14.600 0.400 ;
    END
  END FrameStrobe[2]
  PIN FrameStrobe[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 195.160 0.000 195.560 0.480 ;
    END
  END FrameStrobe[30]
  PIN FrameStrobe[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 205.720 0.000 206.120 0.480 ;
    END
  END FrameStrobe[31]
  PIN FrameStrobe[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 216.280 0.000 216.680 0.480 ;
    END
  END FrameStrobe[32]
  PIN FrameStrobe[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 226.840 0.000 227.240 0.480 ;
    END
  END FrameStrobe[33]
  PIN FrameStrobe[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 237.400 0.000 237.800 0.480 ;
    END
  END FrameStrobe[34]
  PIN FrameStrobe[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 247.960 0.000 248.360 0.480 ;
    END
  END FrameStrobe[35]
  PIN FrameStrobe[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 258.520 0.000 258.920 0.480 ;
    END
  END FrameStrobe[36]
  PIN FrameStrobe[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 269.080 0.000 269.480 0.480 ;
    END
  END FrameStrobe[37]
  PIN FrameStrobe[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 279.640 0.000 280.040 0.480 ;
    END
  END FrameStrobe[38]
  PIN FrameStrobe[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 290.200 0.000 290.600 0.480 ;
    END
  END FrameStrobe[39]
  PIN FrameStrobe[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 17.080 0.000 17.480 0.400 ;
    END
  END FrameStrobe[3]
  PIN FrameStrobe[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 374.200 0.000 374.600 0.480 ;
    END
  END FrameStrobe[40]
  PIN FrameStrobe[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 381.880 0.000 382.280 0.480 ;
    END
  END FrameStrobe[41]
  PIN FrameStrobe[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 389.560 0.000 389.960 0.480 ;
    END
  END FrameStrobe[42]
  PIN FrameStrobe[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 397.240 0.000 397.640 0.480 ;
    END
  END FrameStrobe[43]
  PIN FrameStrobe[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 404.920 0.000 405.320 0.480 ;
    END
  END FrameStrobe[44]
  PIN FrameStrobe[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 412.600 0.000 413.000 0.480 ;
    END
  END FrameStrobe[45]
  PIN FrameStrobe[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 420.280 0.000 420.680 0.480 ;
    END
  END FrameStrobe[46]
  PIN FrameStrobe[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 427.960 0.000 428.360 0.480 ;
    END
  END FrameStrobe[47]
  PIN FrameStrobe[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 435.640 0.000 436.040 0.480 ;
    END
  END FrameStrobe[48]
  PIN FrameStrobe[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 443.320 0.000 443.720 0.480 ;
    END
  END FrameStrobe[49]
  PIN FrameStrobe[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 19.960 0.000 20.360 0.400 ;
    END
  END FrameStrobe[4]
  PIN FrameStrobe[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 451.000 0.000 451.400 0.480 ;
    END
  END FrameStrobe[50]
  PIN FrameStrobe[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 458.680 0.000 459.080 0.480 ;
    END
  END FrameStrobe[51]
  PIN FrameStrobe[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 466.360 0.000 466.760 0.480 ;
    END
  END FrameStrobe[52]
  PIN FrameStrobe[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 474.040 0.000 474.440 0.480 ;
    END
  END FrameStrobe[53]
  PIN FrameStrobe[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 481.720 0.000 482.120 0.480 ;
    END
  END FrameStrobe[54]
  PIN FrameStrobe[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 489.400 0.000 489.800 0.480 ;
    END
  END FrameStrobe[55]
  PIN FrameStrobe[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 497.080 0.000 497.480 0.480 ;
    END
  END FrameStrobe[56]
  PIN FrameStrobe[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 504.760 0.000 505.160 0.480 ;
    END
  END FrameStrobe[57]
  PIN FrameStrobe[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 512.440 0.000 512.840 0.480 ;
    END
  END FrameStrobe[58]
  PIN FrameStrobe[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 520.120 0.000 520.520 0.480 ;
    END
  END FrameStrobe[59]
  PIN FrameStrobe[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 22.840 0.000 23.240 0.400 ;
    END
  END FrameStrobe[5]
  PIN FrameStrobe[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.361400 ;
    PORT
      LAYER Metal3 ;
        RECT 591.640 0.000 592.040 0.480 ;
    END
  END FrameStrobe[60]
  PIN FrameStrobe[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 600.280 0.000 600.680 0.480 ;
    END
  END FrameStrobe[61]
  PIN FrameStrobe[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 608.920 0.000 609.320 0.480 ;
    END
  END FrameStrobe[62]
  PIN FrameStrobe[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 617.560 0.000 617.960 0.480 ;
    END
  END FrameStrobe[63]
  PIN FrameStrobe[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 626.200 0.000 626.600 0.480 ;
    END
  END FrameStrobe[64]
  PIN FrameStrobe[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 634.840 0.000 635.240 0.480 ;
    END
  END FrameStrobe[65]
  PIN FrameStrobe[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 643.480 0.000 643.880 0.480 ;
    END
  END FrameStrobe[66]
  PIN FrameStrobe[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 652.120 0.000 652.520 0.480 ;
    END
  END FrameStrobe[67]
  PIN FrameStrobe[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 660.760 0.000 661.160 0.480 ;
    END
  END FrameStrobe[68]
  PIN FrameStrobe[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 669.400 0.000 669.800 0.480 ;
    END
  END FrameStrobe[69]
  PIN FrameStrobe[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 25.720 0.000 26.120 0.400 ;
    END
  END FrameStrobe[6]
  PIN FrameStrobe[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 678.040 0.000 678.440 0.480 ;
    END
  END FrameStrobe[70]
  PIN FrameStrobe[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 686.680 0.000 687.080 0.480 ;
    END
  END FrameStrobe[71]
  PIN FrameStrobe[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 695.320 0.000 695.720 0.480 ;
    END
  END FrameStrobe[72]
  PIN FrameStrobe[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 703.960 0.000 704.360 0.480 ;
    END
  END FrameStrobe[73]
  PIN FrameStrobe[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 712.600 0.000 713.000 0.480 ;
    END
  END FrameStrobe[74]
  PIN FrameStrobe[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 721.240 0.000 721.640 0.480 ;
    END
  END FrameStrobe[75]
  PIN FrameStrobe[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 729.880 0.000 730.280 0.480 ;
    END
  END FrameStrobe[76]
  PIN FrameStrobe[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 738.520 0.000 738.920 0.480 ;
    END
  END FrameStrobe[77]
  PIN FrameStrobe[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 747.160 0.000 747.560 0.480 ;
    END
  END FrameStrobe[78]
  PIN FrameStrobe[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 755.800 0.000 756.200 0.480 ;
    END
  END FrameStrobe[79]
  PIN FrameStrobe[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 28.600 0.000 29.000 0.400 ;
    END
  END FrameStrobe[7]
  PIN FrameStrobe[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 785.080 0.000 785.480 0.480 ;
    END
  END FrameStrobe[80]
  PIN FrameStrobe[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 797.560 0.000 797.960 0.480 ;
    END
  END FrameStrobe[81]
  PIN FrameStrobe[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 810.040 0.000 810.440 0.480 ;
    END
  END FrameStrobe[82]
  PIN FrameStrobe[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 822.520 0.000 822.920 0.480 ;
    END
  END FrameStrobe[83]
  PIN FrameStrobe[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 835.000 0.000 835.400 0.480 ;
    END
  END FrameStrobe[84]
  PIN FrameStrobe[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 847.480 0.000 847.880 0.480 ;
    END
  END FrameStrobe[85]
  PIN FrameStrobe[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 859.960 0.000 860.360 0.480 ;
    END
  END FrameStrobe[86]
  PIN FrameStrobe[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 872.440 0.000 872.840 0.480 ;
    END
  END FrameStrobe[87]
  PIN FrameStrobe[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 884.920 0.000 885.320 0.480 ;
    END
  END FrameStrobe[88]
  PIN FrameStrobe[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 897.400 0.000 897.800 0.480 ;
    END
  END FrameStrobe[89]
  PIN FrameStrobe[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 31.480 0.000 31.880 0.400 ;
    END
  END FrameStrobe[8]
  PIN FrameStrobe[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 909.880 0.000 910.280 0.480 ;
    END
  END FrameStrobe[90]
  PIN FrameStrobe[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 922.360 0.000 922.760 0.480 ;
    END
  END FrameStrobe[91]
  PIN FrameStrobe[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 934.840 0.000 935.240 0.480 ;
    END
  END FrameStrobe[92]
  PIN FrameStrobe[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 947.320 0.000 947.720 0.480 ;
    END
  END FrameStrobe[93]
  PIN FrameStrobe[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 959.800 0.000 960.200 0.480 ;
    END
  END FrameStrobe[94]
  PIN FrameStrobe[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 972.280 0.000 972.680 0.480 ;
    END
  END FrameStrobe[95]
  PIN FrameStrobe[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 984.760 0.000 985.160 0.480 ;
    END
  END FrameStrobe[96]
  PIN FrameStrobe[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 997.240 0.000 997.640 0.480 ;
    END
  END FrameStrobe[97]
  PIN FrameStrobe[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1009.720 0.000 1010.120 0.480 ;
    END
  END FrameStrobe[98]
  PIN FrameStrobe[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1022.200 0.000 1022.600 0.480 ;
    END
  END FrameStrobe[99]
  PIN FrameStrobe[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 34.360 0.000 34.760 0.400 ;
    END
  END FrameStrobe[9]
  PIN Tile_X0Y10_A_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1043.080 0.930 1043.480 ;
    END
  END Tile_X0Y10_A_I_top
  PIN Tile_X0Y10_A_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1038.040 0.860 1038.440 ;
    END
  END Tile_X0Y10_A_O_top
  PIN Tile_X0Y10_A_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1048.120 0.860 1048.520 ;
    END
  END Tile_X0Y10_A_T_top
  PIN Tile_X0Y10_A_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1068.280 0.930 1068.680 ;
    END
  END Tile_X0Y10_A_config_C_bit0
  PIN Tile_X0Y10_A_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1073.320 0.930 1073.720 ;
    END
  END Tile_X0Y10_A_config_C_bit1
  PIN Tile_X0Y10_A_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1078.360 0.860 1078.760 ;
    END
  END Tile_X0Y10_A_config_C_bit2
  PIN Tile_X0Y10_A_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1083.400 0.930 1083.800 ;
    END
  END Tile_X0Y10_A_config_C_bit3
  PIN Tile_X0Y10_B_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1058.200 0.930 1058.600 ;
    END
  END Tile_X0Y10_B_I_top
  PIN Tile_X0Y10_B_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1053.160 0.930 1053.560 ;
    END
  END Tile_X0Y10_B_O_top
  PIN Tile_X0Y10_B_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1063.240 0.930 1063.640 ;
    END
  END Tile_X0Y10_B_T_top
  PIN Tile_X0Y10_B_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1088.440 0.930 1088.840 ;
    END
  END Tile_X0Y10_B_config_C_bit0
  PIN Tile_X0Y10_B_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1093.480 0.930 1093.880 ;
    END
  END Tile_X0Y10_B_config_C_bit1
  PIN Tile_X0Y10_B_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1098.520 0.860 1098.920 ;
    END
  END Tile_X0Y10_B_config_C_bit2
  PIN Tile_X0Y10_B_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1103.560 0.930 1103.960 ;
    END
  END Tile_X0Y10_B_config_C_bit3
  PIN Tile_X0Y11_A_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 801.160 0.930 801.560 ;
    END
  END Tile_X0Y11_A_I_top
  PIN Tile_X0Y11_A_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 796.120 0.860 796.520 ;
    END
  END Tile_X0Y11_A_O_top
  PIN Tile_X0Y11_A_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 806.200 0.860 806.600 ;
    END
  END Tile_X0Y11_A_T_top
  PIN Tile_X0Y11_A_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 826.360 0.930 826.760 ;
    END
  END Tile_X0Y11_A_config_C_bit0
  PIN Tile_X0Y11_A_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 831.400 0.930 831.800 ;
    END
  END Tile_X0Y11_A_config_C_bit1
  PIN Tile_X0Y11_A_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 836.440 0.860 836.840 ;
    END
  END Tile_X0Y11_A_config_C_bit2
  PIN Tile_X0Y11_A_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 841.480 0.930 841.880 ;
    END
  END Tile_X0Y11_A_config_C_bit3
  PIN Tile_X0Y11_B_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 816.280 0.930 816.680 ;
    END
  END Tile_X0Y11_B_I_top
  PIN Tile_X0Y11_B_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 811.240 0.930 811.640 ;
    END
  END Tile_X0Y11_B_O_top
  PIN Tile_X0Y11_B_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 821.320 0.930 821.720 ;
    END
  END Tile_X0Y11_B_T_top
  PIN Tile_X0Y11_B_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 846.520 0.930 846.920 ;
    END
  END Tile_X0Y11_B_config_C_bit0
  PIN Tile_X0Y11_B_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 851.560 0.930 851.960 ;
    END
  END Tile_X0Y11_B_config_C_bit1
  PIN Tile_X0Y11_B_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 856.600 0.860 857.000 ;
    END
  END Tile_X0Y11_B_config_C_bit2
  PIN Tile_X0Y11_B_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 861.640 0.930 862.040 ;
    END
  END Tile_X0Y11_B_config_C_bit3
  PIN Tile_X0Y12_A_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 559.240 0.930 559.640 ;
    END
  END Tile_X0Y12_A_I_top
  PIN Tile_X0Y12_A_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 554.200 0.860 554.600 ;
    END
  END Tile_X0Y12_A_O_top
  PIN Tile_X0Y12_A_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 564.280 0.860 564.680 ;
    END
  END Tile_X0Y12_A_T_top
  PIN Tile_X0Y12_A_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 584.440 0.930 584.840 ;
    END
  END Tile_X0Y12_A_config_C_bit0
  PIN Tile_X0Y12_A_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 589.480 0.930 589.880 ;
    END
  END Tile_X0Y12_A_config_C_bit1
  PIN Tile_X0Y12_A_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 594.520 0.860 594.920 ;
    END
  END Tile_X0Y12_A_config_C_bit2
  PIN Tile_X0Y12_A_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 599.560 0.930 599.960 ;
    END
  END Tile_X0Y12_A_config_C_bit3
  PIN Tile_X0Y12_B_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 574.360 0.930 574.760 ;
    END
  END Tile_X0Y12_B_I_top
  PIN Tile_X0Y12_B_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 569.320 0.930 569.720 ;
    END
  END Tile_X0Y12_B_O_top
  PIN Tile_X0Y12_B_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 579.400 0.930 579.800 ;
    END
  END Tile_X0Y12_B_T_top
  PIN Tile_X0Y12_B_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 604.600 0.930 605.000 ;
    END
  END Tile_X0Y12_B_config_C_bit0
  PIN Tile_X0Y12_B_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 609.640 0.930 610.040 ;
    END
  END Tile_X0Y12_B_config_C_bit1
  PIN Tile_X0Y12_B_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 614.680 0.860 615.080 ;
    END
  END Tile_X0Y12_B_config_C_bit2
  PIN Tile_X0Y12_B_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 619.720 0.930 620.120 ;
    END
  END Tile_X0Y12_B_config_C_bit3
  PIN Tile_X0Y13_A_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 317.320 0.930 317.720 ;
    END
  END Tile_X0Y13_A_I_top
  PIN Tile_X0Y13_A_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 312.280 0.860 312.680 ;
    END
  END Tile_X0Y13_A_O_top
  PIN Tile_X0Y13_A_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 322.360 0.860 322.760 ;
    END
  END Tile_X0Y13_A_T_top
  PIN Tile_X0Y13_A_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 342.520 0.930 342.920 ;
    END
  END Tile_X0Y13_A_config_C_bit0
  PIN Tile_X0Y13_A_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 347.560 0.930 347.960 ;
    END
  END Tile_X0Y13_A_config_C_bit1
  PIN Tile_X0Y13_A_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 352.600 0.860 353.000 ;
    END
  END Tile_X0Y13_A_config_C_bit2
  PIN Tile_X0Y13_A_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 357.640 0.930 358.040 ;
    END
  END Tile_X0Y13_A_config_C_bit3
  PIN Tile_X0Y13_B_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 332.440 0.930 332.840 ;
    END
  END Tile_X0Y13_B_I_top
  PIN Tile_X0Y13_B_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 327.400 0.930 327.800 ;
    END
  END Tile_X0Y13_B_O_top
  PIN Tile_X0Y13_B_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 337.480 0.930 337.880 ;
    END
  END Tile_X0Y13_B_T_top
  PIN Tile_X0Y13_B_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 362.680 0.930 363.080 ;
    END
  END Tile_X0Y13_B_config_C_bit0
  PIN Tile_X0Y13_B_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 367.720 0.930 368.120 ;
    END
  END Tile_X0Y13_B_config_C_bit1
  PIN Tile_X0Y13_B_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 372.760 0.860 373.160 ;
    END
  END Tile_X0Y13_B_config_C_bit2
  PIN Tile_X0Y13_B_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 377.800 0.930 378.200 ;
    END
  END Tile_X0Y13_B_config_C_bit3
  PIN Tile_X0Y14_A_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 75.400 0.930 75.800 ;
    END
  END Tile_X0Y14_A_I_top
  PIN Tile_X0Y14_A_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 66.160 0.480 66.560 ;
    END
  END Tile_X0Y14_A_O_top
  PIN Tile_X0Y14_A_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 80.440 0.860 80.840 ;
    END
  END Tile_X0Y14_A_T_top
  PIN Tile_X0Y14_A_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 100.600 0.930 101.000 ;
    END
  END Tile_X0Y14_A_config_C_bit0
  PIN Tile_X0Y14_A_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 105.640 0.930 106.040 ;
    END
  END Tile_X0Y14_A_config_C_bit1
  PIN Tile_X0Y14_A_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 110.680 0.860 111.080 ;
    END
  END Tile_X0Y14_A_config_C_bit2
  PIN Tile_X0Y14_A_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 115.720 0.930 116.120 ;
    END
  END Tile_X0Y14_A_config_C_bit3
  PIN Tile_X0Y14_B_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 90.520 0.930 90.920 ;
    END
  END Tile_X0Y14_B_I_top
  PIN Tile_X0Y14_B_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 85.480 0.930 85.880 ;
    END
  END Tile_X0Y14_B_O_top
  PIN Tile_X0Y14_B_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 95.560 0.930 95.960 ;
    END
  END Tile_X0Y14_B_T_top
  PIN Tile_X0Y14_B_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 120.760 0.930 121.160 ;
    END
  END Tile_X0Y14_B_config_C_bit0
  PIN Tile_X0Y14_B_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 125.800 0.930 126.200 ;
    END
  END Tile_X0Y14_B_config_C_bit1
  PIN Tile_X0Y14_B_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 130.840 0.860 131.240 ;
    END
  END Tile_X0Y14_B_config_C_bit2
  PIN Tile_X0Y14_B_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 135.880 0.930 136.280 ;
    END
  END Tile_X0Y14_B_config_C_bit3
  PIN Tile_X0Y1_A_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 3220.360 0.930 3220.760 ;
    END
  END Tile_X0Y1_A_I_top
  PIN Tile_X0Y1_A_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 3215.320 0.860 3215.720 ;
    END
  END Tile_X0Y1_A_O_top
  PIN Tile_X0Y1_A_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 3225.400 0.860 3225.800 ;
    END
  END Tile_X0Y1_A_T_top
  PIN Tile_X0Y1_A_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 3245.560 0.930 3245.960 ;
    END
  END Tile_X0Y1_A_config_C_bit0
  PIN Tile_X0Y1_A_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 3250.600 0.930 3251.000 ;
    END
  END Tile_X0Y1_A_config_C_bit1
  PIN Tile_X0Y1_A_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 3255.640 0.860 3256.040 ;
    END
  END Tile_X0Y1_A_config_C_bit2
  PIN Tile_X0Y1_A_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 3260.680 0.930 3261.080 ;
    END
  END Tile_X0Y1_A_config_C_bit3
  PIN Tile_X0Y1_B_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 3235.480 0.930 3235.880 ;
    END
  END Tile_X0Y1_B_I_top
  PIN Tile_X0Y1_B_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 3230.440 0.930 3230.840 ;
    END
  END Tile_X0Y1_B_O_top
  PIN Tile_X0Y1_B_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 3240.520 0.930 3240.920 ;
    END
  END Tile_X0Y1_B_T_top
  PIN Tile_X0Y1_B_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 3265.720 0.930 3266.120 ;
    END
  END Tile_X0Y1_B_config_C_bit0
  PIN Tile_X0Y1_B_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 3270.760 0.930 3271.160 ;
    END
  END Tile_X0Y1_B_config_C_bit1
  PIN Tile_X0Y1_B_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 3275.800 0.860 3276.200 ;
    END
  END Tile_X0Y1_B_config_C_bit2
  PIN Tile_X0Y1_B_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 3280.840 0.930 3281.240 ;
    END
  END Tile_X0Y1_B_config_C_bit3
  PIN Tile_X0Y2_A_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2978.440 0.930 2978.840 ;
    END
  END Tile_X0Y2_A_I_top
  PIN Tile_X0Y2_A_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2973.400 0.860 2973.800 ;
    END
  END Tile_X0Y2_A_O_top
  PIN Tile_X0Y2_A_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2983.480 0.860 2983.880 ;
    END
  END Tile_X0Y2_A_T_top
  PIN Tile_X0Y2_A_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 3003.640 0.930 3004.040 ;
    END
  END Tile_X0Y2_A_config_C_bit0
  PIN Tile_X0Y2_A_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 3008.680 0.930 3009.080 ;
    END
  END Tile_X0Y2_A_config_C_bit1
  PIN Tile_X0Y2_A_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 3013.720 0.860 3014.120 ;
    END
  END Tile_X0Y2_A_config_C_bit2
  PIN Tile_X0Y2_A_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 3018.760 0.930 3019.160 ;
    END
  END Tile_X0Y2_A_config_C_bit3
  PIN Tile_X0Y2_B_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2993.560 0.930 2993.960 ;
    END
  END Tile_X0Y2_B_I_top
  PIN Tile_X0Y2_B_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2988.520 0.930 2988.920 ;
    END
  END Tile_X0Y2_B_O_top
  PIN Tile_X0Y2_B_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2998.600 0.930 2999.000 ;
    END
  END Tile_X0Y2_B_T_top
  PIN Tile_X0Y2_B_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 3023.800 0.930 3024.200 ;
    END
  END Tile_X0Y2_B_config_C_bit0
  PIN Tile_X0Y2_B_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 3028.840 0.930 3029.240 ;
    END
  END Tile_X0Y2_B_config_C_bit1
  PIN Tile_X0Y2_B_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 3033.880 0.860 3034.280 ;
    END
  END Tile_X0Y2_B_config_C_bit2
  PIN Tile_X0Y2_B_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 3038.920 0.930 3039.320 ;
    END
  END Tile_X0Y2_B_config_C_bit3
  PIN Tile_X0Y3_A_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2736.520 0.930 2736.920 ;
    END
  END Tile_X0Y3_A_I_top
  PIN Tile_X0Y3_A_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2731.480 0.860 2731.880 ;
    END
  END Tile_X0Y3_A_O_top
  PIN Tile_X0Y3_A_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2741.560 0.860 2741.960 ;
    END
  END Tile_X0Y3_A_T_top
  PIN Tile_X0Y3_A_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2761.720 0.930 2762.120 ;
    END
  END Tile_X0Y3_A_config_C_bit0
  PIN Tile_X0Y3_A_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2766.760 0.930 2767.160 ;
    END
  END Tile_X0Y3_A_config_C_bit1
  PIN Tile_X0Y3_A_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2771.800 0.860 2772.200 ;
    END
  END Tile_X0Y3_A_config_C_bit2
  PIN Tile_X0Y3_A_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2776.840 0.930 2777.240 ;
    END
  END Tile_X0Y3_A_config_C_bit3
  PIN Tile_X0Y3_B_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2751.640 0.930 2752.040 ;
    END
  END Tile_X0Y3_B_I_top
  PIN Tile_X0Y3_B_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2746.600 0.930 2747.000 ;
    END
  END Tile_X0Y3_B_O_top
  PIN Tile_X0Y3_B_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2756.680 0.930 2757.080 ;
    END
  END Tile_X0Y3_B_T_top
  PIN Tile_X0Y3_B_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2781.880 0.930 2782.280 ;
    END
  END Tile_X0Y3_B_config_C_bit0
  PIN Tile_X0Y3_B_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2786.920 0.930 2787.320 ;
    END
  END Tile_X0Y3_B_config_C_bit1
  PIN Tile_X0Y3_B_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2791.960 0.860 2792.360 ;
    END
  END Tile_X0Y3_B_config_C_bit2
  PIN Tile_X0Y3_B_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2797.000 0.930 2797.400 ;
    END
  END Tile_X0Y3_B_config_C_bit3
  PIN Tile_X0Y4_A_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2494.600 0.930 2495.000 ;
    END
  END Tile_X0Y4_A_I_top
  PIN Tile_X0Y4_A_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2489.560 0.860 2489.960 ;
    END
  END Tile_X0Y4_A_O_top
  PIN Tile_X0Y4_A_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2499.640 0.860 2500.040 ;
    END
  END Tile_X0Y4_A_T_top
  PIN Tile_X0Y4_A_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2519.800 0.930 2520.200 ;
    END
  END Tile_X0Y4_A_config_C_bit0
  PIN Tile_X0Y4_A_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2524.840 0.930 2525.240 ;
    END
  END Tile_X0Y4_A_config_C_bit1
  PIN Tile_X0Y4_A_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2529.880 0.860 2530.280 ;
    END
  END Tile_X0Y4_A_config_C_bit2
  PIN Tile_X0Y4_A_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2534.920 0.930 2535.320 ;
    END
  END Tile_X0Y4_A_config_C_bit3
  PIN Tile_X0Y4_B_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2509.720 0.930 2510.120 ;
    END
  END Tile_X0Y4_B_I_top
  PIN Tile_X0Y4_B_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2504.680 0.930 2505.080 ;
    END
  END Tile_X0Y4_B_O_top
  PIN Tile_X0Y4_B_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2514.760 0.930 2515.160 ;
    END
  END Tile_X0Y4_B_T_top
  PIN Tile_X0Y4_B_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2539.960 0.930 2540.360 ;
    END
  END Tile_X0Y4_B_config_C_bit0
  PIN Tile_X0Y4_B_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2545.000 0.930 2545.400 ;
    END
  END Tile_X0Y4_B_config_C_bit1
  PIN Tile_X0Y4_B_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2550.040 0.860 2550.440 ;
    END
  END Tile_X0Y4_B_config_C_bit2
  PIN Tile_X0Y4_B_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2555.080 0.930 2555.480 ;
    END
  END Tile_X0Y4_B_config_C_bit3
  PIN Tile_X0Y5_A_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2252.680 0.930 2253.080 ;
    END
  END Tile_X0Y5_A_I_top
  PIN Tile_X0Y5_A_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2247.640 0.860 2248.040 ;
    END
  END Tile_X0Y5_A_O_top
  PIN Tile_X0Y5_A_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2257.720 0.860 2258.120 ;
    END
  END Tile_X0Y5_A_T_top
  PIN Tile_X0Y5_A_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2277.880 0.930 2278.280 ;
    END
  END Tile_X0Y5_A_config_C_bit0
  PIN Tile_X0Y5_A_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2282.920 0.930 2283.320 ;
    END
  END Tile_X0Y5_A_config_C_bit1
  PIN Tile_X0Y5_A_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2287.960 0.860 2288.360 ;
    END
  END Tile_X0Y5_A_config_C_bit2
  PIN Tile_X0Y5_A_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2293.000 0.930 2293.400 ;
    END
  END Tile_X0Y5_A_config_C_bit3
  PIN Tile_X0Y5_B_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2267.800 0.930 2268.200 ;
    END
  END Tile_X0Y5_B_I_top
  PIN Tile_X0Y5_B_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2262.760 0.930 2263.160 ;
    END
  END Tile_X0Y5_B_O_top
  PIN Tile_X0Y5_B_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2272.840 0.930 2273.240 ;
    END
  END Tile_X0Y5_B_T_top
  PIN Tile_X0Y5_B_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2298.040 0.930 2298.440 ;
    END
  END Tile_X0Y5_B_config_C_bit0
  PIN Tile_X0Y5_B_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2303.080 0.930 2303.480 ;
    END
  END Tile_X0Y5_B_config_C_bit1
  PIN Tile_X0Y5_B_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2308.120 0.860 2308.520 ;
    END
  END Tile_X0Y5_B_config_C_bit2
  PIN Tile_X0Y5_B_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2313.160 0.930 2313.560 ;
    END
  END Tile_X0Y5_B_config_C_bit3
  PIN Tile_X0Y6_A_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2010.760 0.930 2011.160 ;
    END
  END Tile_X0Y6_A_I_top
  PIN Tile_X0Y6_A_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2005.720 0.860 2006.120 ;
    END
  END Tile_X0Y6_A_O_top
  PIN Tile_X0Y6_A_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2015.800 0.860 2016.200 ;
    END
  END Tile_X0Y6_A_T_top
  PIN Tile_X0Y6_A_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2035.960 0.930 2036.360 ;
    END
  END Tile_X0Y6_A_config_C_bit0
  PIN Tile_X0Y6_A_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2041.000 0.930 2041.400 ;
    END
  END Tile_X0Y6_A_config_C_bit1
  PIN Tile_X0Y6_A_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2046.040 0.860 2046.440 ;
    END
  END Tile_X0Y6_A_config_C_bit2
  PIN Tile_X0Y6_A_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2051.080 0.930 2051.480 ;
    END
  END Tile_X0Y6_A_config_C_bit3
  PIN Tile_X0Y6_B_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2025.880 0.930 2026.280 ;
    END
  END Tile_X0Y6_B_I_top
  PIN Tile_X0Y6_B_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2020.840 0.930 2021.240 ;
    END
  END Tile_X0Y6_B_O_top
  PIN Tile_X0Y6_B_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2030.920 0.930 2031.320 ;
    END
  END Tile_X0Y6_B_T_top
  PIN Tile_X0Y6_B_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2056.120 0.930 2056.520 ;
    END
  END Tile_X0Y6_B_config_C_bit0
  PIN Tile_X0Y6_B_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2061.160 0.930 2061.560 ;
    END
  END Tile_X0Y6_B_config_C_bit1
  PIN Tile_X0Y6_B_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2066.200 0.860 2066.600 ;
    END
  END Tile_X0Y6_B_config_C_bit2
  PIN Tile_X0Y6_B_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2071.240 0.930 2071.640 ;
    END
  END Tile_X0Y6_B_config_C_bit3
  PIN Tile_X0Y7_A_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1768.840 0.930 1769.240 ;
    END
  END Tile_X0Y7_A_I_top
  PIN Tile_X0Y7_A_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1763.800 0.860 1764.200 ;
    END
  END Tile_X0Y7_A_O_top
  PIN Tile_X0Y7_A_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1773.880 0.860 1774.280 ;
    END
  END Tile_X0Y7_A_T_top
  PIN Tile_X0Y7_A_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1794.040 0.930 1794.440 ;
    END
  END Tile_X0Y7_A_config_C_bit0
  PIN Tile_X0Y7_A_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1799.080 0.930 1799.480 ;
    END
  END Tile_X0Y7_A_config_C_bit1
  PIN Tile_X0Y7_A_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1804.120 0.860 1804.520 ;
    END
  END Tile_X0Y7_A_config_C_bit2
  PIN Tile_X0Y7_A_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1809.160 0.930 1809.560 ;
    END
  END Tile_X0Y7_A_config_C_bit3
  PIN Tile_X0Y7_B_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1783.960 0.930 1784.360 ;
    END
  END Tile_X0Y7_B_I_top
  PIN Tile_X0Y7_B_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1778.920 0.930 1779.320 ;
    END
  END Tile_X0Y7_B_O_top
  PIN Tile_X0Y7_B_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1789.000 0.930 1789.400 ;
    END
  END Tile_X0Y7_B_T_top
  PIN Tile_X0Y7_B_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1814.200 0.930 1814.600 ;
    END
  END Tile_X0Y7_B_config_C_bit0
  PIN Tile_X0Y7_B_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1819.240 0.930 1819.640 ;
    END
  END Tile_X0Y7_B_config_C_bit1
  PIN Tile_X0Y7_B_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1824.280 0.860 1824.680 ;
    END
  END Tile_X0Y7_B_config_C_bit2
  PIN Tile_X0Y7_B_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1829.320 0.930 1829.720 ;
    END
  END Tile_X0Y7_B_config_C_bit3
  PIN Tile_X0Y8_A_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1526.920 0.930 1527.320 ;
    END
  END Tile_X0Y8_A_I_top
  PIN Tile_X0Y8_A_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1521.880 0.860 1522.280 ;
    END
  END Tile_X0Y8_A_O_top
  PIN Tile_X0Y8_A_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1531.960 0.860 1532.360 ;
    END
  END Tile_X0Y8_A_T_top
  PIN Tile_X0Y8_A_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1552.120 0.930 1552.520 ;
    END
  END Tile_X0Y8_A_config_C_bit0
  PIN Tile_X0Y8_A_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1557.160 0.930 1557.560 ;
    END
  END Tile_X0Y8_A_config_C_bit1
  PIN Tile_X0Y8_A_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1562.200 0.860 1562.600 ;
    END
  END Tile_X0Y8_A_config_C_bit2
  PIN Tile_X0Y8_A_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1567.240 0.930 1567.640 ;
    END
  END Tile_X0Y8_A_config_C_bit3
  PIN Tile_X0Y8_B_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1542.040 0.930 1542.440 ;
    END
  END Tile_X0Y8_B_I_top
  PIN Tile_X0Y8_B_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1537.000 0.930 1537.400 ;
    END
  END Tile_X0Y8_B_O_top
  PIN Tile_X0Y8_B_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1547.080 0.930 1547.480 ;
    END
  END Tile_X0Y8_B_T_top
  PIN Tile_X0Y8_B_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1572.280 0.930 1572.680 ;
    END
  END Tile_X0Y8_B_config_C_bit0
  PIN Tile_X0Y8_B_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1577.320 0.930 1577.720 ;
    END
  END Tile_X0Y8_B_config_C_bit1
  PIN Tile_X0Y8_B_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1582.360 0.860 1582.760 ;
    END
  END Tile_X0Y8_B_config_C_bit2
  PIN Tile_X0Y8_B_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1587.400 0.930 1587.800 ;
    END
  END Tile_X0Y8_B_config_C_bit3
  PIN Tile_X0Y9_A_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1285.000 0.930 1285.400 ;
    END
  END Tile_X0Y9_A_I_top
  PIN Tile_X0Y9_A_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1279.960 0.860 1280.360 ;
    END
  END Tile_X0Y9_A_O_top
  PIN Tile_X0Y9_A_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1290.040 0.860 1290.440 ;
    END
  END Tile_X0Y9_A_T_top
  PIN Tile_X0Y9_A_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1310.200 0.930 1310.600 ;
    END
  END Tile_X0Y9_A_config_C_bit0
  PIN Tile_X0Y9_A_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1315.240 0.930 1315.640 ;
    END
  END Tile_X0Y9_A_config_C_bit1
  PIN Tile_X0Y9_A_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1320.280 0.860 1320.680 ;
    END
  END Tile_X0Y9_A_config_C_bit2
  PIN Tile_X0Y9_A_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1325.320 0.930 1325.720 ;
    END
  END Tile_X0Y9_A_config_C_bit3
  PIN Tile_X0Y9_B_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1300.120 0.930 1300.520 ;
    END
  END Tile_X0Y9_B_I_top
  PIN Tile_X0Y9_B_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1295.080 0.930 1295.480 ;
    END
  END Tile_X0Y9_B_O_top
  PIN Tile_X0Y9_B_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1305.160 0.930 1305.560 ;
    END
  END Tile_X0Y9_B_T_top
  PIN Tile_X0Y9_B_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1330.360 0.930 1330.760 ;
    END
  END Tile_X0Y9_B_config_C_bit0
  PIN Tile_X0Y9_B_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1335.400 0.930 1335.800 ;
    END
  END Tile_X0Y9_B_config_C_bit1
  PIN Tile_X0Y9_B_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1340.440 0.860 1340.840 ;
    END
  END Tile_X0Y9_B_config_C_bit2
  PIN Tile_X0Y9_B_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1345.480 0.930 1345.880 ;
    END
  END Tile_X0Y9_B_config_C_bit3
  PIN Tile_X10Y10_ADDR_SRAM0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1133.800 2263.200 1134.200 ;
    END
  END Tile_X10Y10_ADDR_SRAM0
  PIN Tile_X10Y10_ADDR_SRAM1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.340 1136.320 2263.200 1136.720 ;
    END
  END Tile_X10Y10_ADDR_SRAM1
  PIN Tile_X10Y10_ADDR_SRAM2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1138.840 2263.200 1139.240 ;
    END
  END Tile_X10Y10_ADDR_SRAM2
  PIN Tile_X10Y10_ADDR_SRAM3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1141.360 2263.200 1141.760 ;
    END
  END Tile_X10Y10_ADDR_SRAM3
  PIN Tile_X10Y10_ADDR_SRAM4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1143.880 2263.200 1144.280 ;
    END
  END Tile_X10Y10_ADDR_SRAM4
  PIN Tile_X10Y10_ADDR_SRAM5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1146.400 2263.200 1146.800 ;
    END
  END Tile_X10Y10_ADDR_SRAM5
  PIN Tile_X10Y10_ADDR_SRAM6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1148.920 2263.200 1149.320 ;
    END
  END Tile_X10Y10_ADDR_SRAM6
  PIN Tile_X10Y10_ADDR_SRAM7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1151.440 2263.200 1151.840 ;
    END
  END Tile_X10Y10_ADDR_SRAM7
  PIN Tile_X10Y10_ADDR_SRAM8
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1153.960 2263.200 1154.360 ;
    END
  END Tile_X10Y10_ADDR_SRAM8
  PIN Tile_X10Y10_ADDR_SRAM9
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1156.480 2263.200 1156.880 ;
    END
  END Tile_X10Y10_ADDR_SRAM9
  PIN Tile_X10Y10_BM_SRAM0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1159.000 2263.200 1159.400 ;
    END
  END Tile_X10Y10_BM_SRAM0
  PIN Tile_X10Y10_BM_SRAM1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1161.520 2263.200 1161.920 ;
    END
  END Tile_X10Y10_BM_SRAM1
  PIN Tile_X10Y10_BM_SRAM10
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1184.200 2263.200 1184.600 ;
    END
  END Tile_X10Y10_BM_SRAM10
  PIN Tile_X10Y10_BM_SRAM11
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1186.720 2263.200 1187.120 ;
    END
  END Tile_X10Y10_BM_SRAM11
  PIN Tile_X10Y10_BM_SRAM12
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1189.240 2263.200 1189.640 ;
    END
  END Tile_X10Y10_BM_SRAM12
  PIN Tile_X10Y10_BM_SRAM13
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1191.760 2263.200 1192.160 ;
    END
  END Tile_X10Y10_BM_SRAM13
  PIN Tile_X10Y10_BM_SRAM14
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1194.280 2263.200 1194.680 ;
    END
  END Tile_X10Y10_BM_SRAM14
  PIN Tile_X10Y10_BM_SRAM15
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1196.800 2263.200 1197.200 ;
    END
  END Tile_X10Y10_BM_SRAM15
  PIN Tile_X10Y10_BM_SRAM16
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1199.320 2263.200 1199.720 ;
    END
  END Tile_X10Y10_BM_SRAM16
  PIN Tile_X10Y10_BM_SRAM17
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1201.840 2263.200 1202.240 ;
    END
  END Tile_X10Y10_BM_SRAM17
  PIN Tile_X10Y10_BM_SRAM18
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1204.360 2263.200 1204.760 ;
    END
  END Tile_X10Y10_BM_SRAM18
  PIN Tile_X10Y10_BM_SRAM19
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1206.880 2263.200 1207.280 ;
    END
  END Tile_X10Y10_BM_SRAM19
  PIN Tile_X10Y10_BM_SRAM2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1164.040 2263.200 1164.440 ;
    END
  END Tile_X10Y10_BM_SRAM2
  PIN Tile_X10Y10_BM_SRAM20
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1209.400 2263.200 1209.800 ;
    END
  END Tile_X10Y10_BM_SRAM20
  PIN Tile_X10Y10_BM_SRAM21
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1211.920 2263.200 1212.320 ;
    END
  END Tile_X10Y10_BM_SRAM21
  PIN Tile_X10Y10_BM_SRAM22
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1214.440 2263.200 1214.840 ;
    END
  END Tile_X10Y10_BM_SRAM22
  PIN Tile_X10Y10_BM_SRAM23
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1216.960 2263.200 1217.360 ;
    END
  END Tile_X10Y10_BM_SRAM23
  PIN Tile_X10Y10_BM_SRAM24
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1219.480 2263.200 1219.880 ;
    END
  END Tile_X10Y10_BM_SRAM24
  PIN Tile_X10Y10_BM_SRAM25
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1222.000 2263.200 1222.400 ;
    END
  END Tile_X10Y10_BM_SRAM25
  PIN Tile_X10Y10_BM_SRAM26
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1224.520 2263.200 1224.920 ;
    END
  END Tile_X10Y10_BM_SRAM26
  PIN Tile_X10Y10_BM_SRAM27
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1227.040 2263.200 1227.440 ;
    END
  END Tile_X10Y10_BM_SRAM27
  PIN Tile_X10Y10_BM_SRAM28
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1229.560 2263.200 1229.960 ;
    END
  END Tile_X10Y10_BM_SRAM28
  PIN Tile_X10Y10_BM_SRAM29
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1232.080 2263.200 1232.480 ;
    END
  END Tile_X10Y10_BM_SRAM29
  PIN Tile_X10Y10_BM_SRAM3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1166.560 2263.200 1166.960 ;
    END
  END Tile_X10Y10_BM_SRAM3
  PIN Tile_X10Y10_BM_SRAM30
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1234.600 2263.200 1235.000 ;
    END
  END Tile_X10Y10_BM_SRAM30
  PIN Tile_X10Y10_BM_SRAM31
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1237.120 2263.200 1237.520 ;
    END
  END Tile_X10Y10_BM_SRAM31
  PIN Tile_X10Y10_BM_SRAM4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1169.080 2263.200 1169.480 ;
    END
  END Tile_X10Y10_BM_SRAM4
  PIN Tile_X10Y10_BM_SRAM5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1171.600 2263.200 1172.000 ;
    END
  END Tile_X10Y10_BM_SRAM5
  PIN Tile_X10Y10_BM_SRAM6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1174.120 2263.200 1174.520 ;
    END
  END Tile_X10Y10_BM_SRAM6
  PIN Tile_X10Y10_BM_SRAM7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1176.640 2263.200 1177.040 ;
    END
  END Tile_X10Y10_BM_SRAM7
  PIN Tile_X10Y10_BM_SRAM8
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1179.160 2263.200 1179.560 ;
    END
  END Tile_X10Y10_BM_SRAM8
  PIN Tile_X10Y10_BM_SRAM9
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1181.680 2263.200 1182.080 ;
    END
  END Tile_X10Y10_BM_SRAM9
  PIN Tile_X10Y10_CLK_SRAM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1239.640 2263.200 1240.040 ;
    END
  END Tile_X10Y10_CLK_SRAM
  PIN Tile_X10Y10_CONFIGURED_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1050.640 2263.200 1051.040 ;
    END
  END Tile_X10Y10_CONFIGURED_top
  PIN Tile_X10Y10_DIN_SRAM0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1242.160 2263.200 1242.560 ;
    END
  END Tile_X10Y10_DIN_SRAM0
  PIN Tile_X10Y10_DIN_SRAM1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1244.680 2263.200 1245.080 ;
    END
  END Tile_X10Y10_DIN_SRAM1
  PIN Tile_X10Y10_DIN_SRAM10
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1267.360 2263.200 1267.760 ;
    END
  END Tile_X10Y10_DIN_SRAM10
  PIN Tile_X10Y10_DIN_SRAM11
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1269.880 2263.200 1270.280 ;
    END
  END Tile_X10Y10_DIN_SRAM11
  PIN Tile_X10Y10_DIN_SRAM12
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1272.400 2263.200 1272.800 ;
    END
  END Tile_X10Y10_DIN_SRAM12
  PIN Tile_X10Y10_DIN_SRAM13
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1274.920 2263.200 1275.320 ;
    END
  END Tile_X10Y10_DIN_SRAM13
  PIN Tile_X10Y10_DIN_SRAM14
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1277.440 2263.200 1277.840 ;
    END
  END Tile_X10Y10_DIN_SRAM14
  PIN Tile_X10Y10_DIN_SRAM15
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1279.960 2263.200 1280.360 ;
    END
  END Tile_X10Y10_DIN_SRAM15
  PIN Tile_X10Y10_DIN_SRAM16
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1282.480 2263.200 1282.880 ;
    END
  END Tile_X10Y10_DIN_SRAM16
  PIN Tile_X10Y10_DIN_SRAM17
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1285.000 2263.200 1285.400 ;
    END
  END Tile_X10Y10_DIN_SRAM17
  PIN Tile_X10Y10_DIN_SRAM18
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1287.520 2263.200 1287.920 ;
    END
  END Tile_X10Y10_DIN_SRAM18
  PIN Tile_X10Y10_DIN_SRAM19
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1290.040 2263.200 1290.440 ;
    END
  END Tile_X10Y10_DIN_SRAM19
  PIN Tile_X10Y10_DIN_SRAM2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1247.200 2263.200 1247.600 ;
    END
  END Tile_X10Y10_DIN_SRAM2
  PIN Tile_X10Y10_DIN_SRAM20
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1292.560 2263.200 1292.960 ;
    END
  END Tile_X10Y10_DIN_SRAM20
  PIN Tile_X10Y10_DIN_SRAM21
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1295.080 2263.200 1295.480 ;
    END
  END Tile_X10Y10_DIN_SRAM21
  PIN Tile_X10Y10_DIN_SRAM22
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1297.600 2263.200 1298.000 ;
    END
  END Tile_X10Y10_DIN_SRAM22
  PIN Tile_X10Y10_DIN_SRAM23
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1300.120 2263.200 1300.520 ;
    END
  END Tile_X10Y10_DIN_SRAM23
  PIN Tile_X10Y10_DIN_SRAM24
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1302.640 2263.200 1303.040 ;
    END
  END Tile_X10Y10_DIN_SRAM24
  PIN Tile_X10Y10_DIN_SRAM25
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1305.160 2263.200 1305.560 ;
    END
  END Tile_X10Y10_DIN_SRAM25
  PIN Tile_X10Y10_DIN_SRAM26
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1307.680 2263.200 1308.080 ;
    END
  END Tile_X10Y10_DIN_SRAM26
  PIN Tile_X10Y10_DIN_SRAM27
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1310.200 2263.200 1310.600 ;
    END
  END Tile_X10Y10_DIN_SRAM27
  PIN Tile_X10Y10_DIN_SRAM28
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1312.720 2263.200 1313.120 ;
    END
  END Tile_X10Y10_DIN_SRAM28
  PIN Tile_X10Y10_DIN_SRAM29
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1315.240 2263.200 1315.640 ;
    END
  END Tile_X10Y10_DIN_SRAM29
  PIN Tile_X10Y10_DIN_SRAM3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1249.720 2263.200 1250.120 ;
    END
  END Tile_X10Y10_DIN_SRAM3
  PIN Tile_X10Y10_DIN_SRAM30
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1317.760 2263.200 1318.160 ;
    END
  END Tile_X10Y10_DIN_SRAM30
  PIN Tile_X10Y10_DIN_SRAM31
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1320.280 2263.200 1320.680 ;
    END
  END Tile_X10Y10_DIN_SRAM31
  PIN Tile_X10Y10_DIN_SRAM4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1252.240 2263.200 1252.640 ;
    END
  END Tile_X10Y10_DIN_SRAM4
  PIN Tile_X10Y10_DIN_SRAM5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1254.760 2263.200 1255.160 ;
    END
  END Tile_X10Y10_DIN_SRAM5
  PIN Tile_X10Y10_DIN_SRAM6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1257.280 2263.200 1257.680 ;
    END
  END Tile_X10Y10_DIN_SRAM6
  PIN Tile_X10Y10_DIN_SRAM7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1259.800 2263.200 1260.200 ;
    END
  END Tile_X10Y10_DIN_SRAM7
  PIN Tile_X10Y10_DIN_SRAM8
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1262.320 2263.200 1262.720 ;
    END
  END Tile_X10Y10_DIN_SRAM8
  PIN Tile_X10Y10_DIN_SRAM9
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1264.840 2263.200 1265.240 ;
    END
  END Tile_X10Y10_DIN_SRAM9
  PIN Tile_X10Y10_DOUT_SRAM0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1053.160 2263.200 1053.560 ;
    END
  END Tile_X10Y10_DOUT_SRAM0
  PIN Tile_X10Y10_DOUT_SRAM1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1055.680 2263.200 1056.080 ;
    END
  END Tile_X10Y10_DOUT_SRAM1
  PIN Tile_X10Y10_DOUT_SRAM10
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1078.360 2263.200 1078.760 ;
    END
  END Tile_X10Y10_DOUT_SRAM10
  PIN Tile_X10Y10_DOUT_SRAM11
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1080.880 2263.200 1081.280 ;
    END
  END Tile_X10Y10_DOUT_SRAM11
  PIN Tile_X10Y10_DOUT_SRAM12
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1083.400 2263.200 1083.800 ;
    END
  END Tile_X10Y10_DOUT_SRAM12
  PIN Tile_X10Y10_DOUT_SRAM13
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1085.920 2263.200 1086.320 ;
    END
  END Tile_X10Y10_DOUT_SRAM13
  PIN Tile_X10Y10_DOUT_SRAM14
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1088.440 2263.200 1088.840 ;
    END
  END Tile_X10Y10_DOUT_SRAM14
  PIN Tile_X10Y10_DOUT_SRAM15
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1090.960 2263.200 1091.360 ;
    END
  END Tile_X10Y10_DOUT_SRAM15
  PIN Tile_X10Y10_DOUT_SRAM16
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1093.480 2263.200 1093.880 ;
    END
  END Tile_X10Y10_DOUT_SRAM16
  PIN Tile_X10Y10_DOUT_SRAM17
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1096.000 2263.200 1096.400 ;
    END
  END Tile_X10Y10_DOUT_SRAM17
  PIN Tile_X10Y10_DOUT_SRAM18
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1098.520 2263.200 1098.920 ;
    END
  END Tile_X10Y10_DOUT_SRAM18
  PIN Tile_X10Y10_DOUT_SRAM19
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1101.040 2263.200 1101.440 ;
    END
  END Tile_X10Y10_DOUT_SRAM19
  PIN Tile_X10Y10_DOUT_SRAM2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1058.200 2263.200 1058.600 ;
    END
  END Tile_X10Y10_DOUT_SRAM2
  PIN Tile_X10Y10_DOUT_SRAM20
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1103.560 2263.200 1103.960 ;
    END
  END Tile_X10Y10_DOUT_SRAM20
  PIN Tile_X10Y10_DOUT_SRAM21
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1106.080 2263.200 1106.480 ;
    END
  END Tile_X10Y10_DOUT_SRAM21
  PIN Tile_X10Y10_DOUT_SRAM22
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1108.600 2263.200 1109.000 ;
    END
  END Tile_X10Y10_DOUT_SRAM22
  PIN Tile_X10Y10_DOUT_SRAM23
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1111.120 2263.200 1111.520 ;
    END
  END Tile_X10Y10_DOUT_SRAM23
  PIN Tile_X10Y10_DOUT_SRAM24
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1113.640 2263.200 1114.040 ;
    END
  END Tile_X10Y10_DOUT_SRAM24
  PIN Tile_X10Y10_DOUT_SRAM25
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1116.160 2263.200 1116.560 ;
    END
  END Tile_X10Y10_DOUT_SRAM25
  PIN Tile_X10Y10_DOUT_SRAM26
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1118.680 2263.200 1119.080 ;
    END
  END Tile_X10Y10_DOUT_SRAM26
  PIN Tile_X10Y10_DOUT_SRAM27
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1121.200 2263.200 1121.600 ;
    END
  END Tile_X10Y10_DOUT_SRAM27
  PIN Tile_X10Y10_DOUT_SRAM28
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1123.720 2263.200 1124.120 ;
    END
  END Tile_X10Y10_DOUT_SRAM28
  PIN Tile_X10Y10_DOUT_SRAM29
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1126.240 2263.200 1126.640 ;
    END
  END Tile_X10Y10_DOUT_SRAM29
  PIN Tile_X10Y10_DOUT_SRAM3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1060.720 2263.200 1061.120 ;
    END
  END Tile_X10Y10_DOUT_SRAM3
  PIN Tile_X10Y10_DOUT_SRAM30
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1128.760 2263.200 1129.160 ;
    END
  END Tile_X10Y10_DOUT_SRAM30
  PIN Tile_X10Y10_DOUT_SRAM31
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1131.280 2263.200 1131.680 ;
    END
  END Tile_X10Y10_DOUT_SRAM31
  PIN Tile_X10Y10_DOUT_SRAM4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1063.240 2263.200 1063.640 ;
    END
  END Tile_X10Y10_DOUT_SRAM4
  PIN Tile_X10Y10_DOUT_SRAM5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1065.760 2263.200 1066.160 ;
    END
  END Tile_X10Y10_DOUT_SRAM5
  PIN Tile_X10Y10_DOUT_SRAM6
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1068.280 2263.200 1068.680 ;
    END
  END Tile_X10Y10_DOUT_SRAM6
  PIN Tile_X10Y10_DOUT_SRAM7
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1070.800 2263.200 1071.200 ;
    END
  END Tile_X10Y10_DOUT_SRAM7
  PIN Tile_X10Y10_DOUT_SRAM8
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1073.320 2263.200 1073.720 ;
    END
  END Tile_X10Y10_DOUT_SRAM8
  PIN Tile_X10Y10_DOUT_SRAM9
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1075.840 2263.200 1076.240 ;
    END
  END Tile_X10Y10_DOUT_SRAM9
  PIN Tile_X10Y10_MEN_SRAM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1322.800 2263.200 1323.200 ;
    END
  END Tile_X10Y10_MEN_SRAM
  PIN Tile_X10Y10_REN_SRAM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1325.320 2263.200 1325.720 ;
    END
  END Tile_X10Y10_REN_SRAM
  PIN Tile_X10Y10_TIE_HIGH_SRAM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.392700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1327.840 2263.200 1328.240 ;
    END
  END Tile_X10Y10_TIE_HIGH_SRAM
  PIN Tile_X10Y10_TIE_LOW_SRAM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1330.360 2263.200 1330.760 ;
    END
  END Tile_X10Y10_TIE_LOW_SRAM
  PIN Tile_X10Y10_WEN_SRAM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1332.880 2263.200 1333.280 ;
    END
  END Tile_X10Y10_WEN_SRAM
  PIN Tile_X10Y12_ADDR_SRAM0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 649.960 2263.200 650.360 ;
    END
  END Tile_X10Y12_ADDR_SRAM0
  PIN Tile_X10Y12_ADDR_SRAM1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.340 652.480 2263.200 652.880 ;
    END
  END Tile_X10Y12_ADDR_SRAM1
  PIN Tile_X10Y12_ADDR_SRAM2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 655.000 2263.200 655.400 ;
    END
  END Tile_X10Y12_ADDR_SRAM2
  PIN Tile_X10Y12_ADDR_SRAM3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 657.520 2263.200 657.920 ;
    END
  END Tile_X10Y12_ADDR_SRAM3
  PIN Tile_X10Y12_ADDR_SRAM4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 660.040 2263.200 660.440 ;
    END
  END Tile_X10Y12_ADDR_SRAM4
  PIN Tile_X10Y12_ADDR_SRAM5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 662.560 2263.200 662.960 ;
    END
  END Tile_X10Y12_ADDR_SRAM5
  PIN Tile_X10Y12_ADDR_SRAM6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 665.080 2263.200 665.480 ;
    END
  END Tile_X10Y12_ADDR_SRAM6
  PIN Tile_X10Y12_ADDR_SRAM7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 667.600 2263.200 668.000 ;
    END
  END Tile_X10Y12_ADDR_SRAM7
  PIN Tile_X10Y12_ADDR_SRAM8
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 670.120 2263.200 670.520 ;
    END
  END Tile_X10Y12_ADDR_SRAM8
  PIN Tile_X10Y12_ADDR_SRAM9
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 672.640 2263.200 673.040 ;
    END
  END Tile_X10Y12_ADDR_SRAM9
  PIN Tile_X10Y12_BM_SRAM0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 675.160 2263.200 675.560 ;
    END
  END Tile_X10Y12_BM_SRAM0
  PIN Tile_X10Y12_BM_SRAM1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 677.680 2263.200 678.080 ;
    END
  END Tile_X10Y12_BM_SRAM1
  PIN Tile_X10Y12_BM_SRAM10
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 700.360 2263.200 700.760 ;
    END
  END Tile_X10Y12_BM_SRAM10
  PIN Tile_X10Y12_BM_SRAM11
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 702.880 2263.200 703.280 ;
    END
  END Tile_X10Y12_BM_SRAM11
  PIN Tile_X10Y12_BM_SRAM12
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 705.400 2263.200 705.800 ;
    END
  END Tile_X10Y12_BM_SRAM12
  PIN Tile_X10Y12_BM_SRAM13
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 707.920 2263.200 708.320 ;
    END
  END Tile_X10Y12_BM_SRAM13
  PIN Tile_X10Y12_BM_SRAM14
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 710.440 2263.200 710.840 ;
    END
  END Tile_X10Y12_BM_SRAM14
  PIN Tile_X10Y12_BM_SRAM15
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 712.960 2263.200 713.360 ;
    END
  END Tile_X10Y12_BM_SRAM15
  PIN Tile_X10Y12_BM_SRAM16
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 715.480 2263.200 715.880 ;
    END
  END Tile_X10Y12_BM_SRAM16
  PIN Tile_X10Y12_BM_SRAM17
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 718.000 2263.200 718.400 ;
    END
  END Tile_X10Y12_BM_SRAM17
  PIN Tile_X10Y12_BM_SRAM18
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 720.520 2263.200 720.920 ;
    END
  END Tile_X10Y12_BM_SRAM18
  PIN Tile_X10Y12_BM_SRAM19
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 723.040 2263.200 723.440 ;
    END
  END Tile_X10Y12_BM_SRAM19
  PIN Tile_X10Y12_BM_SRAM2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 680.200 2263.200 680.600 ;
    END
  END Tile_X10Y12_BM_SRAM2
  PIN Tile_X10Y12_BM_SRAM20
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 725.560 2263.200 725.960 ;
    END
  END Tile_X10Y12_BM_SRAM20
  PIN Tile_X10Y12_BM_SRAM21
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 728.080 2263.200 728.480 ;
    END
  END Tile_X10Y12_BM_SRAM21
  PIN Tile_X10Y12_BM_SRAM22
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 730.600 2263.200 731.000 ;
    END
  END Tile_X10Y12_BM_SRAM22
  PIN Tile_X10Y12_BM_SRAM23
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 733.120 2263.200 733.520 ;
    END
  END Tile_X10Y12_BM_SRAM23
  PIN Tile_X10Y12_BM_SRAM24
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 735.640 2263.200 736.040 ;
    END
  END Tile_X10Y12_BM_SRAM24
  PIN Tile_X10Y12_BM_SRAM25
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 738.160 2263.200 738.560 ;
    END
  END Tile_X10Y12_BM_SRAM25
  PIN Tile_X10Y12_BM_SRAM26
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 740.680 2263.200 741.080 ;
    END
  END Tile_X10Y12_BM_SRAM26
  PIN Tile_X10Y12_BM_SRAM27
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 743.200 2263.200 743.600 ;
    END
  END Tile_X10Y12_BM_SRAM27
  PIN Tile_X10Y12_BM_SRAM28
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 745.720 2263.200 746.120 ;
    END
  END Tile_X10Y12_BM_SRAM28
  PIN Tile_X10Y12_BM_SRAM29
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 748.240 2263.200 748.640 ;
    END
  END Tile_X10Y12_BM_SRAM29
  PIN Tile_X10Y12_BM_SRAM3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 682.720 2263.200 683.120 ;
    END
  END Tile_X10Y12_BM_SRAM3
  PIN Tile_X10Y12_BM_SRAM30
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 750.760 2263.200 751.160 ;
    END
  END Tile_X10Y12_BM_SRAM30
  PIN Tile_X10Y12_BM_SRAM31
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 753.280 2263.200 753.680 ;
    END
  END Tile_X10Y12_BM_SRAM31
  PIN Tile_X10Y12_BM_SRAM4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 685.240 2263.200 685.640 ;
    END
  END Tile_X10Y12_BM_SRAM4
  PIN Tile_X10Y12_BM_SRAM5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 687.760 2263.200 688.160 ;
    END
  END Tile_X10Y12_BM_SRAM5
  PIN Tile_X10Y12_BM_SRAM6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 690.280 2263.200 690.680 ;
    END
  END Tile_X10Y12_BM_SRAM6
  PIN Tile_X10Y12_BM_SRAM7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 692.800 2263.200 693.200 ;
    END
  END Tile_X10Y12_BM_SRAM7
  PIN Tile_X10Y12_BM_SRAM8
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 695.320 2263.200 695.720 ;
    END
  END Tile_X10Y12_BM_SRAM8
  PIN Tile_X10Y12_BM_SRAM9
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 697.840 2263.200 698.240 ;
    END
  END Tile_X10Y12_BM_SRAM9
  PIN Tile_X10Y12_CLK_SRAM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 755.800 2263.200 756.200 ;
    END
  END Tile_X10Y12_CLK_SRAM
  PIN Tile_X10Y12_CONFIGURED_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 566.800 2263.200 567.200 ;
    END
  END Tile_X10Y12_CONFIGURED_top
  PIN Tile_X10Y12_DIN_SRAM0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 758.320 2263.200 758.720 ;
    END
  END Tile_X10Y12_DIN_SRAM0
  PIN Tile_X10Y12_DIN_SRAM1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 760.840 2263.200 761.240 ;
    END
  END Tile_X10Y12_DIN_SRAM1
  PIN Tile_X10Y12_DIN_SRAM10
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 783.520 2263.200 783.920 ;
    END
  END Tile_X10Y12_DIN_SRAM10
  PIN Tile_X10Y12_DIN_SRAM11
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 786.040 2263.200 786.440 ;
    END
  END Tile_X10Y12_DIN_SRAM11
  PIN Tile_X10Y12_DIN_SRAM12
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 788.560 2263.200 788.960 ;
    END
  END Tile_X10Y12_DIN_SRAM12
  PIN Tile_X10Y12_DIN_SRAM13
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 791.080 2263.200 791.480 ;
    END
  END Tile_X10Y12_DIN_SRAM13
  PIN Tile_X10Y12_DIN_SRAM14
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 793.600 2263.200 794.000 ;
    END
  END Tile_X10Y12_DIN_SRAM14
  PIN Tile_X10Y12_DIN_SRAM15
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 796.120 2263.200 796.520 ;
    END
  END Tile_X10Y12_DIN_SRAM15
  PIN Tile_X10Y12_DIN_SRAM16
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 798.640 2263.200 799.040 ;
    END
  END Tile_X10Y12_DIN_SRAM16
  PIN Tile_X10Y12_DIN_SRAM17
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 801.160 2263.200 801.560 ;
    END
  END Tile_X10Y12_DIN_SRAM17
  PIN Tile_X10Y12_DIN_SRAM18
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 803.680 2263.200 804.080 ;
    END
  END Tile_X10Y12_DIN_SRAM18
  PIN Tile_X10Y12_DIN_SRAM19
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 806.200 2263.200 806.600 ;
    END
  END Tile_X10Y12_DIN_SRAM19
  PIN Tile_X10Y12_DIN_SRAM2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 763.360 2263.200 763.760 ;
    END
  END Tile_X10Y12_DIN_SRAM2
  PIN Tile_X10Y12_DIN_SRAM20
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 808.720 2263.200 809.120 ;
    END
  END Tile_X10Y12_DIN_SRAM20
  PIN Tile_X10Y12_DIN_SRAM21
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 811.240 2263.200 811.640 ;
    END
  END Tile_X10Y12_DIN_SRAM21
  PIN Tile_X10Y12_DIN_SRAM22
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 813.760 2263.200 814.160 ;
    END
  END Tile_X10Y12_DIN_SRAM22
  PIN Tile_X10Y12_DIN_SRAM23
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 816.280 2263.200 816.680 ;
    END
  END Tile_X10Y12_DIN_SRAM23
  PIN Tile_X10Y12_DIN_SRAM24
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 818.800 2263.200 819.200 ;
    END
  END Tile_X10Y12_DIN_SRAM24
  PIN Tile_X10Y12_DIN_SRAM25
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 821.320 2263.200 821.720 ;
    END
  END Tile_X10Y12_DIN_SRAM25
  PIN Tile_X10Y12_DIN_SRAM26
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 823.840 2263.200 824.240 ;
    END
  END Tile_X10Y12_DIN_SRAM26
  PIN Tile_X10Y12_DIN_SRAM27
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 826.360 2263.200 826.760 ;
    END
  END Tile_X10Y12_DIN_SRAM27
  PIN Tile_X10Y12_DIN_SRAM28
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 828.880 2263.200 829.280 ;
    END
  END Tile_X10Y12_DIN_SRAM28
  PIN Tile_X10Y12_DIN_SRAM29
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 831.400 2263.200 831.800 ;
    END
  END Tile_X10Y12_DIN_SRAM29
  PIN Tile_X10Y12_DIN_SRAM3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 765.880 2263.200 766.280 ;
    END
  END Tile_X10Y12_DIN_SRAM3
  PIN Tile_X10Y12_DIN_SRAM30
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 833.920 2263.200 834.320 ;
    END
  END Tile_X10Y12_DIN_SRAM30
  PIN Tile_X10Y12_DIN_SRAM31
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 836.440 2263.200 836.840 ;
    END
  END Tile_X10Y12_DIN_SRAM31
  PIN Tile_X10Y12_DIN_SRAM4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 768.400 2263.200 768.800 ;
    END
  END Tile_X10Y12_DIN_SRAM4
  PIN Tile_X10Y12_DIN_SRAM5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 770.920 2263.200 771.320 ;
    END
  END Tile_X10Y12_DIN_SRAM5
  PIN Tile_X10Y12_DIN_SRAM6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 773.440 2263.200 773.840 ;
    END
  END Tile_X10Y12_DIN_SRAM6
  PIN Tile_X10Y12_DIN_SRAM7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 775.960 2263.200 776.360 ;
    END
  END Tile_X10Y12_DIN_SRAM7
  PIN Tile_X10Y12_DIN_SRAM8
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 778.480 2263.200 778.880 ;
    END
  END Tile_X10Y12_DIN_SRAM8
  PIN Tile_X10Y12_DIN_SRAM9
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 781.000 2263.200 781.400 ;
    END
  END Tile_X10Y12_DIN_SRAM9
  PIN Tile_X10Y12_DOUT_SRAM0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 569.320 2263.200 569.720 ;
    END
  END Tile_X10Y12_DOUT_SRAM0
  PIN Tile_X10Y12_DOUT_SRAM1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 571.840 2263.200 572.240 ;
    END
  END Tile_X10Y12_DOUT_SRAM1
  PIN Tile_X10Y12_DOUT_SRAM10
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 594.520 2263.200 594.920 ;
    END
  END Tile_X10Y12_DOUT_SRAM10
  PIN Tile_X10Y12_DOUT_SRAM11
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 597.040 2263.200 597.440 ;
    END
  END Tile_X10Y12_DOUT_SRAM11
  PIN Tile_X10Y12_DOUT_SRAM12
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 599.560 2263.200 599.960 ;
    END
  END Tile_X10Y12_DOUT_SRAM12
  PIN Tile_X10Y12_DOUT_SRAM13
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 602.080 2263.200 602.480 ;
    END
  END Tile_X10Y12_DOUT_SRAM13
  PIN Tile_X10Y12_DOUT_SRAM14
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 604.600 2263.200 605.000 ;
    END
  END Tile_X10Y12_DOUT_SRAM14
  PIN Tile_X10Y12_DOUT_SRAM15
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 607.120 2263.200 607.520 ;
    END
  END Tile_X10Y12_DOUT_SRAM15
  PIN Tile_X10Y12_DOUT_SRAM16
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 609.640 2263.200 610.040 ;
    END
  END Tile_X10Y12_DOUT_SRAM16
  PIN Tile_X10Y12_DOUT_SRAM17
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 612.160 2263.200 612.560 ;
    END
  END Tile_X10Y12_DOUT_SRAM17
  PIN Tile_X10Y12_DOUT_SRAM18
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 614.680 2263.200 615.080 ;
    END
  END Tile_X10Y12_DOUT_SRAM18
  PIN Tile_X10Y12_DOUT_SRAM19
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 617.200 2263.200 617.600 ;
    END
  END Tile_X10Y12_DOUT_SRAM19
  PIN Tile_X10Y12_DOUT_SRAM2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 574.360 2263.200 574.760 ;
    END
  END Tile_X10Y12_DOUT_SRAM2
  PIN Tile_X10Y12_DOUT_SRAM20
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 619.720 2263.200 620.120 ;
    END
  END Tile_X10Y12_DOUT_SRAM20
  PIN Tile_X10Y12_DOUT_SRAM21
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 622.240 2263.200 622.640 ;
    END
  END Tile_X10Y12_DOUT_SRAM21
  PIN Tile_X10Y12_DOUT_SRAM22
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 624.760 2263.200 625.160 ;
    END
  END Tile_X10Y12_DOUT_SRAM22
  PIN Tile_X10Y12_DOUT_SRAM23
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 627.280 2263.200 627.680 ;
    END
  END Tile_X10Y12_DOUT_SRAM23
  PIN Tile_X10Y12_DOUT_SRAM24
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 629.800 2263.200 630.200 ;
    END
  END Tile_X10Y12_DOUT_SRAM24
  PIN Tile_X10Y12_DOUT_SRAM25
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 632.320 2263.200 632.720 ;
    END
  END Tile_X10Y12_DOUT_SRAM25
  PIN Tile_X10Y12_DOUT_SRAM26
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 634.840 2263.200 635.240 ;
    END
  END Tile_X10Y12_DOUT_SRAM26
  PIN Tile_X10Y12_DOUT_SRAM27
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 637.360 2263.200 637.760 ;
    END
  END Tile_X10Y12_DOUT_SRAM27
  PIN Tile_X10Y12_DOUT_SRAM28
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 639.880 2263.200 640.280 ;
    END
  END Tile_X10Y12_DOUT_SRAM28
  PIN Tile_X10Y12_DOUT_SRAM29
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 642.400 2263.200 642.800 ;
    END
  END Tile_X10Y12_DOUT_SRAM29
  PIN Tile_X10Y12_DOUT_SRAM3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 576.880 2263.200 577.280 ;
    END
  END Tile_X10Y12_DOUT_SRAM3
  PIN Tile_X10Y12_DOUT_SRAM30
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 644.920 2263.200 645.320 ;
    END
  END Tile_X10Y12_DOUT_SRAM30
  PIN Tile_X10Y12_DOUT_SRAM31
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 647.440 2263.200 647.840 ;
    END
  END Tile_X10Y12_DOUT_SRAM31
  PIN Tile_X10Y12_DOUT_SRAM4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 579.400 2263.200 579.800 ;
    END
  END Tile_X10Y12_DOUT_SRAM4
  PIN Tile_X10Y12_DOUT_SRAM5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 581.920 2263.200 582.320 ;
    END
  END Tile_X10Y12_DOUT_SRAM5
  PIN Tile_X10Y12_DOUT_SRAM6
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 584.440 2263.200 584.840 ;
    END
  END Tile_X10Y12_DOUT_SRAM6
  PIN Tile_X10Y12_DOUT_SRAM7
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 586.960 2263.200 587.360 ;
    END
  END Tile_X10Y12_DOUT_SRAM7
  PIN Tile_X10Y12_DOUT_SRAM8
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 589.480 2263.200 589.880 ;
    END
  END Tile_X10Y12_DOUT_SRAM8
  PIN Tile_X10Y12_DOUT_SRAM9
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 592.000 2263.200 592.400 ;
    END
  END Tile_X10Y12_DOUT_SRAM9
  PIN Tile_X10Y12_MEN_SRAM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 838.960 2263.200 839.360 ;
    END
  END Tile_X10Y12_MEN_SRAM
  PIN Tile_X10Y12_REN_SRAM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 841.480 2263.200 841.880 ;
    END
  END Tile_X10Y12_REN_SRAM
  PIN Tile_X10Y12_TIE_HIGH_SRAM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.392700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 844.000 2263.200 844.400 ;
    END
  END Tile_X10Y12_TIE_HIGH_SRAM
  PIN Tile_X10Y12_TIE_LOW_SRAM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 846.520 2263.200 846.920 ;
    END
  END Tile_X10Y12_TIE_LOW_SRAM
  PIN Tile_X10Y12_WEN_SRAM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 849.040 2263.200 849.440 ;
    END
  END Tile_X10Y12_WEN_SRAM
  PIN Tile_X10Y14_ADDR_SRAM0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 166.120 2263.200 166.520 ;
    END
  END Tile_X10Y14_ADDR_SRAM0
  PIN Tile_X10Y14_ADDR_SRAM1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.340 168.640 2263.200 169.040 ;
    END
  END Tile_X10Y14_ADDR_SRAM1
  PIN Tile_X10Y14_ADDR_SRAM2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 171.160 2263.200 171.560 ;
    END
  END Tile_X10Y14_ADDR_SRAM2
  PIN Tile_X10Y14_ADDR_SRAM3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 173.680 2263.200 174.080 ;
    END
  END Tile_X10Y14_ADDR_SRAM3
  PIN Tile_X10Y14_ADDR_SRAM4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 176.200 2263.200 176.600 ;
    END
  END Tile_X10Y14_ADDR_SRAM4
  PIN Tile_X10Y14_ADDR_SRAM5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 178.720 2263.200 179.120 ;
    END
  END Tile_X10Y14_ADDR_SRAM5
  PIN Tile_X10Y14_ADDR_SRAM6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 181.240 2263.200 181.640 ;
    END
  END Tile_X10Y14_ADDR_SRAM6
  PIN Tile_X10Y14_ADDR_SRAM7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 183.760 2263.200 184.160 ;
    END
  END Tile_X10Y14_ADDR_SRAM7
  PIN Tile_X10Y14_ADDR_SRAM8
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 186.280 2263.200 186.680 ;
    END
  END Tile_X10Y14_ADDR_SRAM8
  PIN Tile_X10Y14_ADDR_SRAM9
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 188.800 2263.200 189.200 ;
    END
  END Tile_X10Y14_ADDR_SRAM9
  PIN Tile_X10Y14_BM_SRAM0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 191.320 2263.200 191.720 ;
    END
  END Tile_X10Y14_BM_SRAM0
  PIN Tile_X10Y14_BM_SRAM1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 193.840 2263.200 194.240 ;
    END
  END Tile_X10Y14_BM_SRAM1
  PIN Tile_X10Y14_BM_SRAM10
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 216.520 2263.200 216.920 ;
    END
  END Tile_X10Y14_BM_SRAM10
  PIN Tile_X10Y14_BM_SRAM11
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 219.040 2263.200 219.440 ;
    END
  END Tile_X10Y14_BM_SRAM11
  PIN Tile_X10Y14_BM_SRAM12
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 221.560 2263.200 221.960 ;
    END
  END Tile_X10Y14_BM_SRAM12
  PIN Tile_X10Y14_BM_SRAM13
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 224.080 2263.200 224.480 ;
    END
  END Tile_X10Y14_BM_SRAM13
  PIN Tile_X10Y14_BM_SRAM14
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 226.600 2263.200 227.000 ;
    END
  END Tile_X10Y14_BM_SRAM14
  PIN Tile_X10Y14_BM_SRAM15
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 229.120 2263.200 229.520 ;
    END
  END Tile_X10Y14_BM_SRAM15
  PIN Tile_X10Y14_BM_SRAM16
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 231.640 2263.200 232.040 ;
    END
  END Tile_X10Y14_BM_SRAM16
  PIN Tile_X10Y14_BM_SRAM17
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 234.160 2263.200 234.560 ;
    END
  END Tile_X10Y14_BM_SRAM17
  PIN Tile_X10Y14_BM_SRAM18
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 236.680 2263.200 237.080 ;
    END
  END Tile_X10Y14_BM_SRAM18
  PIN Tile_X10Y14_BM_SRAM19
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 239.200 2263.200 239.600 ;
    END
  END Tile_X10Y14_BM_SRAM19
  PIN Tile_X10Y14_BM_SRAM2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 196.360 2263.200 196.760 ;
    END
  END Tile_X10Y14_BM_SRAM2
  PIN Tile_X10Y14_BM_SRAM20
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 241.720 2263.200 242.120 ;
    END
  END Tile_X10Y14_BM_SRAM20
  PIN Tile_X10Y14_BM_SRAM21
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 244.240 2263.200 244.640 ;
    END
  END Tile_X10Y14_BM_SRAM21
  PIN Tile_X10Y14_BM_SRAM22
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 246.760 2263.200 247.160 ;
    END
  END Tile_X10Y14_BM_SRAM22
  PIN Tile_X10Y14_BM_SRAM23
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 249.280 2263.200 249.680 ;
    END
  END Tile_X10Y14_BM_SRAM23
  PIN Tile_X10Y14_BM_SRAM24
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 251.800 2263.200 252.200 ;
    END
  END Tile_X10Y14_BM_SRAM24
  PIN Tile_X10Y14_BM_SRAM25
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 254.320 2263.200 254.720 ;
    END
  END Tile_X10Y14_BM_SRAM25
  PIN Tile_X10Y14_BM_SRAM26
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 256.840 2263.200 257.240 ;
    END
  END Tile_X10Y14_BM_SRAM26
  PIN Tile_X10Y14_BM_SRAM27
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 259.360 2263.200 259.760 ;
    END
  END Tile_X10Y14_BM_SRAM27
  PIN Tile_X10Y14_BM_SRAM28
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 261.880 2263.200 262.280 ;
    END
  END Tile_X10Y14_BM_SRAM28
  PIN Tile_X10Y14_BM_SRAM29
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 264.400 2263.200 264.800 ;
    END
  END Tile_X10Y14_BM_SRAM29
  PIN Tile_X10Y14_BM_SRAM3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 198.880 2263.200 199.280 ;
    END
  END Tile_X10Y14_BM_SRAM3
  PIN Tile_X10Y14_BM_SRAM30
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 266.920 2263.200 267.320 ;
    END
  END Tile_X10Y14_BM_SRAM30
  PIN Tile_X10Y14_BM_SRAM31
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 269.440 2263.200 269.840 ;
    END
  END Tile_X10Y14_BM_SRAM31
  PIN Tile_X10Y14_BM_SRAM4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 201.400 2263.200 201.800 ;
    END
  END Tile_X10Y14_BM_SRAM4
  PIN Tile_X10Y14_BM_SRAM5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 203.920 2263.200 204.320 ;
    END
  END Tile_X10Y14_BM_SRAM5
  PIN Tile_X10Y14_BM_SRAM6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 206.440 2263.200 206.840 ;
    END
  END Tile_X10Y14_BM_SRAM6
  PIN Tile_X10Y14_BM_SRAM7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 208.960 2263.200 209.360 ;
    END
  END Tile_X10Y14_BM_SRAM7
  PIN Tile_X10Y14_BM_SRAM8
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 211.480 2263.200 211.880 ;
    END
  END Tile_X10Y14_BM_SRAM8
  PIN Tile_X10Y14_BM_SRAM9
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 214.000 2263.200 214.400 ;
    END
  END Tile_X10Y14_BM_SRAM9
  PIN Tile_X10Y14_CLK_SRAM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 271.960 2263.200 272.360 ;
    END
  END Tile_X10Y14_CLK_SRAM
  PIN Tile_X10Y14_CONFIGURED_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 82.960 2263.200 83.360 ;
    END
  END Tile_X10Y14_CONFIGURED_top
  PIN Tile_X10Y14_DIN_SRAM0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 274.480 2263.200 274.880 ;
    END
  END Tile_X10Y14_DIN_SRAM0
  PIN Tile_X10Y14_DIN_SRAM1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 277.000 2263.200 277.400 ;
    END
  END Tile_X10Y14_DIN_SRAM1
  PIN Tile_X10Y14_DIN_SRAM10
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 299.680 2263.200 300.080 ;
    END
  END Tile_X10Y14_DIN_SRAM10
  PIN Tile_X10Y14_DIN_SRAM11
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 302.200 2263.200 302.600 ;
    END
  END Tile_X10Y14_DIN_SRAM11
  PIN Tile_X10Y14_DIN_SRAM12
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 304.720 2263.200 305.120 ;
    END
  END Tile_X10Y14_DIN_SRAM12
  PIN Tile_X10Y14_DIN_SRAM13
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 307.240 2263.200 307.640 ;
    END
  END Tile_X10Y14_DIN_SRAM13
  PIN Tile_X10Y14_DIN_SRAM14
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 309.760 2263.200 310.160 ;
    END
  END Tile_X10Y14_DIN_SRAM14
  PIN Tile_X10Y14_DIN_SRAM15
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 312.280 2263.200 312.680 ;
    END
  END Tile_X10Y14_DIN_SRAM15
  PIN Tile_X10Y14_DIN_SRAM16
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 314.800 2263.200 315.200 ;
    END
  END Tile_X10Y14_DIN_SRAM16
  PIN Tile_X10Y14_DIN_SRAM17
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 317.320 2263.200 317.720 ;
    END
  END Tile_X10Y14_DIN_SRAM17
  PIN Tile_X10Y14_DIN_SRAM18
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 319.840 2263.200 320.240 ;
    END
  END Tile_X10Y14_DIN_SRAM18
  PIN Tile_X10Y14_DIN_SRAM19
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 322.360 2263.200 322.760 ;
    END
  END Tile_X10Y14_DIN_SRAM19
  PIN Tile_X10Y14_DIN_SRAM2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 279.520 2263.200 279.920 ;
    END
  END Tile_X10Y14_DIN_SRAM2
  PIN Tile_X10Y14_DIN_SRAM20
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 324.880 2263.200 325.280 ;
    END
  END Tile_X10Y14_DIN_SRAM20
  PIN Tile_X10Y14_DIN_SRAM21
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 327.400 2263.200 327.800 ;
    END
  END Tile_X10Y14_DIN_SRAM21
  PIN Tile_X10Y14_DIN_SRAM22
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 329.920 2263.200 330.320 ;
    END
  END Tile_X10Y14_DIN_SRAM22
  PIN Tile_X10Y14_DIN_SRAM23
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 332.440 2263.200 332.840 ;
    END
  END Tile_X10Y14_DIN_SRAM23
  PIN Tile_X10Y14_DIN_SRAM24
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 334.960 2263.200 335.360 ;
    END
  END Tile_X10Y14_DIN_SRAM24
  PIN Tile_X10Y14_DIN_SRAM25
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 337.480 2263.200 337.880 ;
    END
  END Tile_X10Y14_DIN_SRAM25
  PIN Tile_X10Y14_DIN_SRAM26
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 340.000 2263.200 340.400 ;
    END
  END Tile_X10Y14_DIN_SRAM26
  PIN Tile_X10Y14_DIN_SRAM27
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 342.520 2263.200 342.920 ;
    END
  END Tile_X10Y14_DIN_SRAM27
  PIN Tile_X10Y14_DIN_SRAM28
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 345.040 2263.200 345.440 ;
    END
  END Tile_X10Y14_DIN_SRAM28
  PIN Tile_X10Y14_DIN_SRAM29
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 347.560 2263.200 347.960 ;
    END
  END Tile_X10Y14_DIN_SRAM29
  PIN Tile_X10Y14_DIN_SRAM3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 282.040 2263.200 282.440 ;
    END
  END Tile_X10Y14_DIN_SRAM3
  PIN Tile_X10Y14_DIN_SRAM30
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 350.080 2263.200 350.480 ;
    END
  END Tile_X10Y14_DIN_SRAM30
  PIN Tile_X10Y14_DIN_SRAM31
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 352.600 2263.200 353.000 ;
    END
  END Tile_X10Y14_DIN_SRAM31
  PIN Tile_X10Y14_DIN_SRAM4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 284.560 2263.200 284.960 ;
    END
  END Tile_X10Y14_DIN_SRAM4
  PIN Tile_X10Y14_DIN_SRAM5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 287.080 2263.200 287.480 ;
    END
  END Tile_X10Y14_DIN_SRAM5
  PIN Tile_X10Y14_DIN_SRAM6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 289.600 2263.200 290.000 ;
    END
  END Tile_X10Y14_DIN_SRAM6
  PIN Tile_X10Y14_DIN_SRAM7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 292.120 2263.200 292.520 ;
    END
  END Tile_X10Y14_DIN_SRAM7
  PIN Tile_X10Y14_DIN_SRAM8
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 294.640 2263.200 295.040 ;
    END
  END Tile_X10Y14_DIN_SRAM8
  PIN Tile_X10Y14_DIN_SRAM9
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 297.160 2263.200 297.560 ;
    END
  END Tile_X10Y14_DIN_SRAM9
  PIN Tile_X10Y14_DOUT_SRAM0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 85.480 2263.200 85.880 ;
    END
  END Tile_X10Y14_DOUT_SRAM0
  PIN Tile_X10Y14_DOUT_SRAM1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 88.000 2263.200 88.400 ;
    END
  END Tile_X10Y14_DOUT_SRAM1
  PIN Tile_X10Y14_DOUT_SRAM10
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 110.680 2263.200 111.080 ;
    END
  END Tile_X10Y14_DOUT_SRAM10
  PIN Tile_X10Y14_DOUT_SRAM11
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 113.200 2263.200 113.600 ;
    END
  END Tile_X10Y14_DOUT_SRAM11
  PIN Tile_X10Y14_DOUT_SRAM12
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 115.720 2263.200 116.120 ;
    END
  END Tile_X10Y14_DOUT_SRAM12
  PIN Tile_X10Y14_DOUT_SRAM13
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 118.240 2263.200 118.640 ;
    END
  END Tile_X10Y14_DOUT_SRAM13
  PIN Tile_X10Y14_DOUT_SRAM14
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 120.760 2263.200 121.160 ;
    END
  END Tile_X10Y14_DOUT_SRAM14
  PIN Tile_X10Y14_DOUT_SRAM15
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 123.280 2263.200 123.680 ;
    END
  END Tile_X10Y14_DOUT_SRAM15
  PIN Tile_X10Y14_DOUT_SRAM16
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 125.800 2263.200 126.200 ;
    END
  END Tile_X10Y14_DOUT_SRAM16
  PIN Tile_X10Y14_DOUT_SRAM17
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 128.320 2263.200 128.720 ;
    END
  END Tile_X10Y14_DOUT_SRAM17
  PIN Tile_X10Y14_DOUT_SRAM18
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 130.840 2263.200 131.240 ;
    END
  END Tile_X10Y14_DOUT_SRAM18
  PIN Tile_X10Y14_DOUT_SRAM19
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 133.360 2263.200 133.760 ;
    END
  END Tile_X10Y14_DOUT_SRAM19
  PIN Tile_X10Y14_DOUT_SRAM2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 90.520 2263.200 90.920 ;
    END
  END Tile_X10Y14_DOUT_SRAM2
  PIN Tile_X10Y14_DOUT_SRAM20
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 135.880 2263.200 136.280 ;
    END
  END Tile_X10Y14_DOUT_SRAM20
  PIN Tile_X10Y14_DOUT_SRAM21
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 138.400 2263.200 138.800 ;
    END
  END Tile_X10Y14_DOUT_SRAM21
  PIN Tile_X10Y14_DOUT_SRAM22
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 140.920 2263.200 141.320 ;
    END
  END Tile_X10Y14_DOUT_SRAM22
  PIN Tile_X10Y14_DOUT_SRAM23
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 143.440 2263.200 143.840 ;
    END
  END Tile_X10Y14_DOUT_SRAM23
  PIN Tile_X10Y14_DOUT_SRAM24
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 145.960 2263.200 146.360 ;
    END
  END Tile_X10Y14_DOUT_SRAM24
  PIN Tile_X10Y14_DOUT_SRAM25
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 148.480 2263.200 148.880 ;
    END
  END Tile_X10Y14_DOUT_SRAM25
  PIN Tile_X10Y14_DOUT_SRAM26
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 151.000 2263.200 151.400 ;
    END
  END Tile_X10Y14_DOUT_SRAM26
  PIN Tile_X10Y14_DOUT_SRAM27
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 153.520 2263.200 153.920 ;
    END
  END Tile_X10Y14_DOUT_SRAM27
  PIN Tile_X10Y14_DOUT_SRAM28
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 156.040 2263.200 156.440 ;
    END
  END Tile_X10Y14_DOUT_SRAM28
  PIN Tile_X10Y14_DOUT_SRAM29
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 158.560 2263.200 158.960 ;
    END
  END Tile_X10Y14_DOUT_SRAM29
  PIN Tile_X10Y14_DOUT_SRAM3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 93.040 2263.200 93.440 ;
    END
  END Tile_X10Y14_DOUT_SRAM3
  PIN Tile_X10Y14_DOUT_SRAM30
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 161.080 2263.200 161.480 ;
    END
  END Tile_X10Y14_DOUT_SRAM30
  PIN Tile_X10Y14_DOUT_SRAM31
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 163.600 2263.200 164.000 ;
    END
  END Tile_X10Y14_DOUT_SRAM31
  PIN Tile_X10Y14_DOUT_SRAM4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 95.560 2263.200 95.960 ;
    END
  END Tile_X10Y14_DOUT_SRAM4
  PIN Tile_X10Y14_DOUT_SRAM5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 98.080 2263.200 98.480 ;
    END
  END Tile_X10Y14_DOUT_SRAM5
  PIN Tile_X10Y14_DOUT_SRAM6
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 100.600 2263.200 101.000 ;
    END
  END Tile_X10Y14_DOUT_SRAM6
  PIN Tile_X10Y14_DOUT_SRAM7
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 103.120 2263.200 103.520 ;
    END
  END Tile_X10Y14_DOUT_SRAM7
  PIN Tile_X10Y14_DOUT_SRAM8
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 105.640 2263.200 106.040 ;
    END
  END Tile_X10Y14_DOUT_SRAM8
  PIN Tile_X10Y14_DOUT_SRAM9
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 108.160 2263.200 108.560 ;
    END
  END Tile_X10Y14_DOUT_SRAM9
  PIN Tile_X10Y14_MEN_SRAM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 355.120 2263.200 355.520 ;
    END
  END Tile_X10Y14_MEN_SRAM
  PIN Tile_X10Y14_REN_SRAM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 357.640 2263.200 358.040 ;
    END
  END Tile_X10Y14_REN_SRAM
  PIN Tile_X10Y14_TIE_HIGH_SRAM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.392700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 360.160 2263.200 360.560 ;
    END
  END Tile_X10Y14_TIE_HIGH_SRAM
  PIN Tile_X10Y14_TIE_LOW_SRAM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 362.680 2263.200 363.080 ;
    END
  END Tile_X10Y14_TIE_LOW_SRAM
  PIN Tile_X10Y14_WEN_SRAM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 365.200 2263.200 365.600 ;
    END
  END Tile_X10Y14_WEN_SRAM
  PIN Tile_X10Y2_ADDR_SRAM0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 3069.160 2263.200 3069.560 ;
    END
  END Tile_X10Y2_ADDR_SRAM0
  PIN Tile_X10Y2_ADDR_SRAM1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.340 3071.680 2263.200 3072.080 ;
    END
  END Tile_X10Y2_ADDR_SRAM1
  PIN Tile_X10Y2_ADDR_SRAM2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 3074.200 2263.200 3074.600 ;
    END
  END Tile_X10Y2_ADDR_SRAM2
  PIN Tile_X10Y2_ADDR_SRAM3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 3076.720 2263.200 3077.120 ;
    END
  END Tile_X10Y2_ADDR_SRAM3
  PIN Tile_X10Y2_ADDR_SRAM4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 3079.240 2263.200 3079.640 ;
    END
  END Tile_X10Y2_ADDR_SRAM4
  PIN Tile_X10Y2_ADDR_SRAM5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 3081.760 2263.200 3082.160 ;
    END
  END Tile_X10Y2_ADDR_SRAM5
  PIN Tile_X10Y2_ADDR_SRAM6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 3084.280 2263.200 3084.680 ;
    END
  END Tile_X10Y2_ADDR_SRAM6
  PIN Tile_X10Y2_ADDR_SRAM7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 3086.800 2263.200 3087.200 ;
    END
  END Tile_X10Y2_ADDR_SRAM7
  PIN Tile_X10Y2_ADDR_SRAM8
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 3089.320 2263.200 3089.720 ;
    END
  END Tile_X10Y2_ADDR_SRAM8
  PIN Tile_X10Y2_ADDR_SRAM9
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 3091.840 2263.200 3092.240 ;
    END
  END Tile_X10Y2_ADDR_SRAM9
  PIN Tile_X10Y2_BM_SRAM0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 3094.360 2263.200 3094.760 ;
    END
  END Tile_X10Y2_BM_SRAM0
  PIN Tile_X10Y2_BM_SRAM1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 3096.880 2263.200 3097.280 ;
    END
  END Tile_X10Y2_BM_SRAM1
  PIN Tile_X10Y2_BM_SRAM10
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 3119.560 2263.200 3119.960 ;
    END
  END Tile_X10Y2_BM_SRAM10
  PIN Tile_X10Y2_BM_SRAM11
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 3122.080 2263.200 3122.480 ;
    END
  END Tile_X10Y2_BM_SRAM11
  PIN Tile_X10Y2_BM_SRAM12
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 3124.600 2263.200 3125.000 ;
    END
  END Tile_X10Y2_BM_SRAM12
  PIN Tile_X10Y2_BM_SRAM13
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 3127.120 2263.200 3127.520 ;
    END
  END Tile_X10Y2_BM_SRAM13
  PIN Tile_X10Y2_BM_SRAM14
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 3129.640 2263.200 3130.040 ;
    END
  END Tile_X10Y2_BM_SRAM14
  PIN Tile_X10Y2_BM_SRAM15
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 3132.160 2263.200 3132.560 ;
    END
  END Tile_X10Y2_BM_SRAM15
  PIN Tile_X10Y2_BM_SRAM16
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 3134.680 2263.200 3135.080 ;
    END
  END Tile_X10Y2_BM_SRAM16
  PIN Tile_X10Y2_BM_SRAM17
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 3137.200 2263.200 3137.600 ;
    END
  END Tile_X10Y2_BM_SRAM17
  PIN Tile_X10Y2_BM_SRAM18
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 3139.720 2263.200 3140.120 ;
    END
  END Tile_X10Y2_BM_SRAM18
  PIN Tile_X10Y2_BM_SRAM19
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 3142.240 2263.200 3142.640 ;
    END
  END Tile_X10Y2_BM_SRAM19
  PIN Tile_X10Y2_BM_SRAM2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 3099.400 2263.200 3099.800 ;
    END
  END Tile_X10Y2_BM_SRAM2
  PIN Tile_X10Y2_BM_SRAM20
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 3144.760 2263.200 3145.160 ;
    END
  END Tile_X10Y2_BM_SRAM20
  PIN Tile_X10Y2_BM_SRAM21
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 3147.280 2263.200 3147.680 ;
    END
  END Tile_X10Y2_BM_SRAM21
  PIN Tile_X10Y2_BM_SRAM22
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 3149.800 2263.200 3150.200 ;
    END
  END Tile_X10Y2_BM_SRAM22
  PIN Tile_X10Y2_BM_SRAM23
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 3152.320 2263.200 3152.720 ;
    END
  END Tile_X10Y2_BM_SRAM23
  PIN Tile_X10Y2_BM_SRAM24
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 3154.840 2263.200 3155.240 ;
    END
  END Tile_X10Y2_BM_SRAM24
  PIN Tile_X10Y2_BM_SRAM25
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 3157.360 2263.200 3157.760 ;
    END
  END Tile_X10Y2_BM_SRAM25
  PIN Tile_X10Y2_BM_SRAM26
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 3159.880 2263.200 3160.280 ;
    END
  END Tile_X10Y2_BM_SRAM26
  PIN Tile_X10Y2_BM_SRAM27
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 3162.400 2263.200 3162.800 ;
    END
  END Tile_X10Y2_BM_SRAM27
  PIN Tile_X10Y2_BM_SRAM28
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 3164.920 2263.200 3165.320 ;
    END
  END Tile_X10Y2_BM_SRAM28
  PIN Tile_X10Y2_BM_SRAM29
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 3167.440 2263.200 3167.840 ;
    END
  END Tile_X10Y2_BM_SRAM29
  PIN Tile_X10Y2_BM_SRAM3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 3101.920 2263.200 3102.320 ;
    END
  END Tile_X10Y2_BM_SRAM3
  PIN Tile_X10Y2_BM_SRAM30
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 3169.960 2263.200 3170.360 ;
    END
  END Tile_X10Y2_BM_SRAM30
  PIN Tile_X10Y2_BM_SRAM31
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 3172.480 2263.200 3172.880 ;
    END
  END Tile_X10Y2_BM_SRAM31
  PIN Tile_X10Y2_BM_SRAM4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 3104.440 2263.200 3104.840 ;
    END
  END Tile_X10Y2_BM_SRAM4
  PIN Tile_X10Y2_BM_SRAM5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 3106.960 2263.200 3107.360 ;
    END
  END Tile_X10Y2_BM_SRAM5
  PIN Tile_X10Y2_BM_SRAM6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 3109.480 2263.200 3109.880 ;
    END
  END Tile_X10Y2_BM_SRAM6
  PIN Tile_X10Y2_BM_SRAM7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 3112.000 2263.200 3112.400 ;
    END
  END Tile_X10Y2_BM_SRAM7
  PIN Tile_X10Y2_BM_SRAM8
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 3114.520 2263.200 3114.920 ;
    END
  END Tile_X10Y2_BM_SRAM8
  PIN Tile_X10Y2_BM_SRAM9
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 3117.040 2263.200 3117.440 ;
    END
  END Tile_X10Y2_BM_SRAM9
  PIN Tile_X10Y2_CLK_SRAM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 3175.000 2263.200 3175.400 ;
    END
  END Tile_X10Y2_CLK_SRAM
  PIN Tile_X10Y2_CONFIGURED_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2986.000 2263.200 2986.400 ;
    END
  END Tile_X10Y2_CONFIGURED_top
  PIN Tile_X10Y2_DIN_SRAM0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 3177.520 2263.200 3177.920 ;
    END
  END Tile_X10Y2_DIN_SRAM0
  PIN Tile_X10Y2_DIN_SRAM1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 3180.040 2263.200 3180.440 ;
    END
  END Tile_X10Y2_DIN_SRAM1
  PIN Tile_X10Y2_DIN_SRAM10
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 3202.720 2263.200 3203.120 ;
    END
  END Tile_X10Y2_DIN_SRAM10
  PIN Tile_X10Y2_DIN_SRAM11
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 3205.240 2263.200 3205.640 ;
    END
  END Tile_X10Y2_DIN_SRAM11
  PIN Tile_X10Y2_DIN_SRAM12
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 3207.760 2263.200 3208.160 ;
    END
  END Tile_X10Y2_DIN_SRAM12
  PIN Tile_X10Y2_DIN_SRAM13
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 3210.280 2263.200 3210.680 ;
    END
  END Tile_X10Y2_DIN_SRAM13
  PIN Tile_X10Y2_DIN_SRAM14
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 3212.800 2263.200 3213.200 ;
    END
  END Tile_X10Y2_DIN_SRAM14
  PIN Tile_X10Y2_DIN_SRAM15
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 3215.320 2263.200 3215.720 ;
    END
  END Tile_X10Y2_DIN_SRAM15
  PIN Tile_X10Y2_DIN_SRAM16
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 3217.840 2263.200 3218.240 ;
    END
  END Tile_X10Y2_DIN_SRAM16
  PIN Tile_X10Y2_DIN_SRAM17
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 3220.360 2263.200 3220.760 ;
    END
  END Tile_X10Y2_DIN_SRAM17
  PIN Tile_X10Y2_DIN_SRAM18
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 3222.880 2263.200 3223.280 ;
    END
  END Tile_X10Y2_DIN_SRAM18
  PIN Tile_X10Y2_DIN_SRAM19
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 3225.400 2263.200 3225.800 ;
    END
  END Tile_X10Y2_DIN_SRAM19
  PIN Tile_X10Y2_DIN_SRAM2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 3182.560 2263.200 3182.960 ;
    END
  END Tile_X10Y2_DIN_SRAM2
  PIN Tile_X10Y2_DIN_SRAM20
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 3227.920 2263.200 3228.320 ;
    END
  END Tile_X10Y2_DIN_SRAM20
  PIN Tile_X10Y2_DIN_SRAM21
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 3230.440 2263.200 3230.840 ;
    END
  END Tile_X10Y2_DIN_SRAM21
  PIN Tile_X10Y2_DIN_SRAM22
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 3232.960 2263.200 3233.360 ;
    END
  END Tile_X10Y2_DIN_SRAM22
  PIN Tile_X10Y2_DIN_SRAM23
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 3235.480 2263.200 3235.880 ;
    END
  END Tile_X10Y2_DIN_SRAM23
  PIN Tile_X10Y2_DIN_SRAM24
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 3238.000 2263.200 3238.400 ;
    END
  END Tile_X10Y2_DIN_SRAM24
  PIN Tile_X10Y2_DIN_SRAM25
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 3240.520 2263.200 3240.920 ;
    END
  END Tile_X10Y2_DIN_SRAM25
  PIN Tile_X10Y2_DIN_SRAM26
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 3243.040 2263.200 3243.440 ;
    END
  END Tile_X10Y2_DIN_SRAM26
  PIN Tile_X10Y2_DIN_SRAM27
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 3245.560 2263.200 3245.960 ;
    END
  END Tile_X10Y2_DIN_SRAM27
  PIN Tile_X10Y2_DIN_SRAM28
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 3248.080 2263.200 3248.480 ;
    END
  END Tile_X10Y2_DIN_SRAM28
  PIN Tile_X10Y2_DIN_SRAM29
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 3250.600 2263.200 3251.000 ;
    END
  END Tile_X10Y2_DIN_SRAM29
  PIN Tile_X10Y2_DIN_SRAM3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 3185.080 2263.200 3185.480 ;
    END
  END Tile_X10Y2_DIN_SRAM3
  PIN Tile_X10Y2_DIN_SRAM30
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 3253.120 2263.200 3253.520 ;
    END
  END Tile_X10Y2_DIN_SRAM30
  PIN Tile_X10Y2_DIN_SRAM31
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 3255.640 2263.200 3256.040 ;
    END
  END Tile_X10Y2_DIN_SRAM31
  PIN Tile_X10Y2_DIN_SRAM4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 3187.600 2263.200 3188.000 ;
    END
  END Tile_X10Y2_DIN_SRAM4
  PIN Tile_X10Y2_DIN_SRAM5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 3190.120 2263.200 3190.520 ;
    END
  END Tile_X10Y2_DIN_SRAM5
  PIN Tile_X10Y2_DIN_SRAM6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 3192.640 2263.200 3193.040 ;
    END
  END Tile_X10Y2_DIN_SRAM6
  PIN Tile_X10Y2_DIN_SRAM7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 3195.160 2263.200 3195.560 ;
    END
  END Tile_X10Y2_DIN_SRAM7
  PIN Tile_X10Y2_DIN_SRAM8
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 3197.680 2263.200 3198.080 ;
    END
  END Tile_X10Y2_DIN_SRAM8
  PIN Tile_X10Y2_DIN_SRAM9
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 3200.200 2263.200 3200.600 ;
    END
  END Tile_X10Y2_DIN_SRAM9
  PIN Tile_X10Y2_DOUT_SRAM0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2988.520 2263.200 2988.920 ;
    END
  END Tile_X10Y2_DOUT_SRAM0
  PIN Tile_X10Y2_DOUT_SRAM1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2991.040 2263.200 2991.440 ;
    END
  END Tile_X10Y2_DOUT_SRAM1
  PIN Tile_X10Y2_DOUT_SRAM10
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 3013.720 2263.200 3014.120 ;
    END
  END Tile_X10Y2_DOUT_SRAM10
  PIN Tile_X10Y2_DOUT_SRAM11
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 3016.240 2263.200 3016.640 ;
    END
  END Tile_X10Y2_DOUT_SRAM11
  PIN Tile_X10Y2_DOUT_SRAM12
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 3018.760 2263.200 3019.160 ;
    END
  END Tile_X10Y2_DOUT_SRAM12
  PIN Tile_X10Y2_DOUT_SRAM13
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 3021.280 2263.200 3021.680 ;
    END
  END Tile_X10Y2_DOUT_SRAM13
  PIN Tile_X10Y2_DOUT_SRAM14
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 3023.800 2263.200 3024.200 ;
    END
  END Tile_X10Y2_DOUT_SRAM14
  PIN Tile_X10Y2_DOUT_SRAM15
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 3026.320 2263.200 3026.720 ;
    END
  END Tile_X10Y2_DOUT_SRAM15
  PIN Tile_X10Y2_DOUT_SRAM16
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 3028.840 2263.200 3029.240 ;
    END
  END Tile_X10Y2_DOUT_SRAM16
  PIN Tile_X10Y2_DOUT_SRAM17
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 3031.360 2263.200 3031.760 ;
    END
  END Tile_X10Y2_DOUT_SRAM17
  PIN Tile_X10Y2_DOUT_SRAM18
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 3033.880 2263.200 3034.280 ;
    END
  END Tile_X10Y2_DOUT_SRAM18
  PIN Tile_X10Y2_DOUT_SRAM19
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 3036.400 2263.200 3036.800 ;
    END
  END Tile_X10Y2_DOUT_SRAM19
  PIN Tile_X10Y2_DOUT_SRAM2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2993.560 2263.200 2993.960 ;
    END
  END Tile_X10Y2_DOUT_SRAM2
  PIN Tile_X10Y2_DOUT_SRAM20
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 3038.920 2263.200 3039.320 ;
    END
  END Tile_X10Y2_DOUT_SRAM20
  PIN Tile_X10Y2_DOUT_SRAM21
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 3041.440 2263.200 3041.840 ;
    END
  END Tile_X10Y2_DOUT_SRAM21
  PIN Tile_X10Y2_DOUT_SRAM22
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 3043.960 2263.200 3044.360 ;
    END
  END Tile_X10Y2_DOUT_SRAM22
  PIN Tile_X10Y2_DOUT_SRAM23
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 3046.480 2263.200 3046.880 ;
    END
  END Tile_X10Y2_DOUT_SRAM23
  PIN Tile_X10Y2_DOUT_SRAM24
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 3049.000 2263.200 3049.400 ;
    END
  END Tile_X10Y2_DOUT_SRAM24
  PIN Tile_X10Y2_DOUT_SRAM25
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 3051.520 2263.200 3051.920 ;
    END
  END Tile_X10Y2_DOUT_SRAM25
  PIN Tile_X10Y2_DOUT_SRAM26
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 3054.040 2263.200 3054.440 ;
    END
  END Tile_X10Y2_DOUT_SRAM26
  PIN Tile_X10Y2_DOUT_SRAM27
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 3056.560 2263.200 3056.960 ;
    END
  END Tile_X10Y2_DOUT_SRAM27
  PIN Tile_X10Y2_DOUT_SRAM28
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 3059.080 2263.200 3059.480 ;
    END
  END Tile_X10Y2_DOUT_SRAM28
  PIN Tile_X10Y2_DOUT_SRAM29
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 3061.600 2263.200 3062.000 ;
    END
  END Tile_X10Y2_DOUT_SRAM29
  PIN Tile_X10Y2_DOUT_SRAM3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2996.080 2263.200 2996.480 ;
    END
  END Tile_X10Y2_DOUT_SRAM3
  PIN Tile_X10Y2_DOUT_SRAM30
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 3064.120 2263.200 3064.520 ;
    END
  END Tile_X10Y2_DOUT_SRAM30
  PIN Tile_X10Y2_DOUT_SRAM31
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 3066.640 2263.200 3067.040 ;
    END
  END Tile_X10Y2_DOUT_SRAM31
  PIN Tile_X10Y2_DOUT_SRAM4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2998.600 2263.200 2999.000 ;
    END
  END Tile_X10Y2_DOUT_SRAM4
  PIN Tile_X10Y2_DOUT_SRAM5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 3001.120 2263.200 3001.520 ;
    END
  END Tile_X10Y2_DOUT_SRAM5
  PIN Tile_X10Y2_DOUT_SRAM6
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 3003.640 2263.200 3004.040 ;
    END
  END Tile_X10Y2_DOUT_SRAM6
  PIN Tile_X10Y2_DOUT_SRAM7
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 3006.160 2263.200 3006.560 ;
    END
  END Tile_X10Y2_DOUT_SRAM7
  PIN Tile_X10Y2_DOUT_SRAM8
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 3008.680 2263.200 3009.080 ;
    END
  END Tile_X10Y2_DOUT_SRAM8
  PIN Tile_X10Y2_DOUT_SRAM9
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 3011.200 2263.200 3011.600 ;
    END
  END Tile_X10Y2_DOUT_SRAM9
  PIN Tile_X10Y2_MEN_SRAM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 3258.160 2263.200 3258.560 ;
    END
  END Tile_X10Y2_MEN_SRAM
  PIN Tile_X10Y2_REN_SRAM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 3260.680 2263.200 3261.080 ;
    END
  END Tile_X10Y2_REN_SRAM
  PIN Tile_X10Y2_TIE_HIGH_SRAM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.392700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 3263.200 2263.200 3263.600 ;
    END
  END Tile_X10Y2_TIE_HIGH_SRAM
  PIN Tile_X10Y2_TIE_LOW_SRAM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 3265.720 2263.200 3266.120 ;
    END
  END Tile_X10Y2_TIE_LOW_SRAM
  PIN Tile_X10Y2_WEN_SRAM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 3268.240 2263.200 3268.640 ;
    END
  END Tile_X10Y2_WEN_SRAM
  PIN Tile_X10Y4_ADDR_SRAM0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2585.320 2263.200 2585.720 ;
    END
  END Tile_X10Y4_ADDR_SRAM0
  PIN Tile_X10Y4_ADDR_SRAM1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.340 2587.840 2263.200 2588.240 ;
    END
  END Tile_X10Y4_ADDR_SRAM1
  PIN Tile_X10Y4_ADDR_SRAM2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2590.360 2263.200 2590.760 ;
    END
  END Tile_X10Y4_ADDR_SRAM2
  PIN Tile_X10Y4_ADDR_SRAM3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2592.880 2263.200 2593.280 ;
    END
  END Tile_X10Y4_ADDR_SRAM3
  PIN Tile_X10Y4_ADDR_SRAM4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2595.400 2263.200 2595.800 ;
    END
  END Tile_X10Y4_ADDR_SRAM4
  PIN Tile_X10Y4_ADDR_SRAM5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2597.920 2263.200 2598.320 ;
    END
  END Tile_X10Y4_ADDR_SRAM5
  PIN Tile_X10Y4_ADDR_SRAM6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2600.440 2263.200 2600.840 ;
    END
  END Tile_X10Y4_ADDR_SRAM6
  PIN Tile_X10Y4_ADDR_SRAM7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2602.960 2263.200 2603.360 ;
    END
  END Tile_X10Y4_ADDR_SRAM7
  PIN Tile_X10Y4_ADDR_SRAM8
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2605.480 2263.200 2605.880 ;
    END
  END Tile_X10Y4_ADDR_SRAM8
  PIN Tile_X10Y4_ADDR_SRAM9
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2608.000 2263.200 2608.400 ;
    END
  END Tile_X10Y4_ADDR_SRAM9
  PIN Tile_X10Y4_BM_SRAM0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2610.520 2263.200 2610.920 ;
    END
  END Tile_X10Y4_BM_SRAM0
  PIN Tile_X10Y4_BM_SRAM1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2613.040 2263.200 2613.440 ;
    END
  END Tile_X10Y4_BM_SRAM1
  PIN Tile_X10Y4_BM_SRAM10
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2635.720 2263.200 2636.120 ;
    END
  END Tile_X10Y4_BM_SRAM10
  PIN Tile_X10Y4_BM_SRAM11
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2638.240 2263.200 2638.640 ;
    END
  END Tile_X10Y4_BM_SRAM11
  PIN Tile_X10Y4_BM_SRAM12
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2640.760 2263.200 2641.160 ;
    END
  END Tile_X10Y4_BM_SRAM12
  PIN Tile_X10Y4_BM_SRAM13
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2643.280 2263.200 2643.680 ;
    END
  END Tile_X10Y4_BM_SRAM13
  PIN Tile_X10Y4_BM_SRAM14
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2645.800 2263.200 2646.200 ;
    END
  END Tile_X10Y4_BM_SRAM14
  PIN Tile_X10Y4_BM_SRAM15
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2648.320 2263.200 2648.720 ;
    END
  END Tile_X10Y4_BM_SRAM15
  PIN Tile_X10Y4_BM_SRAM16
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2650.840 2263.200 2651.240 ;
    END
  END Tile_X10Y4_BM_SRAM16
  PIN Tile_X10Y4_BM_SRAM17
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2653.360 2263.200 2653.760 ;
    END
  END Tile_X10Y4_BM_SRAM17
  PIN Tile_X10Y4_BM_SRAM18
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2655.880 2263.200 2656.280 ;
    END
  END Tile_X10Y4_BM_SRAM18
  PIN Tile_X10Y4_BM_SRAM19
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2658.400 2263.200 2658.800 ;
    END
  END Tile_X10Y4_BM_SRAM19
  PIN Tile_X10Y4_BM_SRAM2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2615.560 2263.200 2615.960 ;
    END
  END Tile_X10Y4_BM_SRAM2
  PIN Tile_X10Y4_BM_SRAM20
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2660.920 2263.200 2661.320 ;
    END
  END Tile_X10Y4_BM_SRAM20
  PIN Tile_X10Y4_BM_SRAM21
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2663.440 2263.200 2663.840 ;
    END
  END Tile_X10Y4_BM_SRAM21
  PIN Tile_X10Y4_BM_SRAM22
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2665.960 2263.200 2666.360 ;
    END
  END Tile_X10Y4_BM_SRAM22
  PIN Tile_X10Y4_BM_SRAM23
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2668.480 2263.200 2668.880 ;
    END
  END Tile_X10Y4_BM_SRAM23
  PIN Tile_X10Y4_BM_SRAM24
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2671.000 2263.200 2671.400 ;
    END
  END Tile_X10Y4_BM_SRAM24
  PIN Tile_X10Y4_BM_SRAM25
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2673.520 2263.200 2673.920 ;
    END
  END Tile_X10Y4_BM_SRAM25
  PIN Tile_X10Y4_BM_SRAM26
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2676.040 2263.200 2676.440 ;
    END
  END Tile_X10Y4_BM_SRAM26
  PIN Tile_X10Y4_BM_SRAM27
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2678.560 2263.200 2678.960 ;
    END
  END Tile_X10Y4_BM_SRAM27
  PIN Tile_X10Y4_BM_SRAM28
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2681.080 2263.200 2681.480 ;
    END
  END Tile_X10Y4_BM_SRAM28
  PIN Tile_X10Y4_BM_SRAM29
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2683.600 2263.200 2684.000 ;
    END
  END Tile_X10Y4_BM_SRAM29
  PIN Tile_X10Y4_BM_SRAM3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2618.080 2263.200 2618.480 ;
    END
  END Tile_X10Y4_BM_SRAM3
  PIN Tile_X10Y4_BM_SRAM30
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2686.120 2263.200 2686.520 ;
    END
  END Tile_X10Y4_BM_SRAM30
  PIN Tile_X10Y4_BM_SRAM31
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2688.640 2263.200 2689.040 ;
    END
  END Tile_X10Y4_BM_SRAM31
  PIN Tile_X10Y4_BM_SRAM4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2620.600 2263.200 2621.000 ;
    END
  END Tile_X10Y4_BM_SRAM4
  PIN Tile_X10Y4_BM_SRAM5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2623.120 2263.200 2623.520 ;
    END
  END Tile_X10Y4_BM_SRAM5
  PIN Tile_X10Y4_BM_SRAM6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2625.640 2263.200 2626.040 ;
    END
  END Tile_X10Y4_BM_SRAM6
  PIN Tile_X10Y4_BM_SRAM7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2628.160 2263.200 2628.560 ;
    END
  END Tile_X10Y4_BM_SRAM7
  PIN Tile_X10Y4_BM_SRAM8
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2630.680 2263.200 2631.080 ;
    END
  END Tile_X10Y4_BM_SRAM8
  PIN Tile_X10Y4_BM_SRAM9
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2633.200 2263.200 2633.600 ;
    END
  END Tile_X10Y4_BM_SRAM9
  PIN Tile_X10Y4_CLK_SRAM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2691.160 2263.200 2691.560 ;
    END
  END Tile_X10Y4_CLK_SRAM
  PIN Tile_X10Y4_CONFIGURED_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2502.160 2263.200 2502.560 ;
    END
  END Tile_X10Y4_CONFIGURED_top
  PIN Tile_X10Y4_DIN_SRAM0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2693.680 2263.200 2694.080 ;
    END
  END Tile_X10Y4_DIN_SRAM0
  PIN Tile_X10Y4_DIN_SRAM1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2696.200 2263.200 2696.600 ;
    END
  END Tile_X10Y4_DIN_SRAM1
  PIN Tile_X10Y4_DIN_SRAM10
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2718.880 2263.200 2719.280 ;
    END
  END Tile_X10Y4_DIN_SRAM10
  PIN Tile_X10Y4_DIN_SRAM11
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2721.400 2263.200 2721.800 ;
    END
  END Tile_X10Y4_DIN_SRAM11
  PIN Tile_X10Y4_DIN_SRAM12
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2723.920 2263.200 2724.320 ;
    END
  END Tile_X10Y4_DIN_SRAM12
  PIN Tile_X10Y4_DIN_SRAM13
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2726.440 2263.200 2726.840 ;
    END
  END Tile_X10Y4_DIN_SRAM13
  PIN Tile_X10Y4_DIN_SRAM14
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2728.960 2263.200 2729.360 ;
    END
  END Tile_X10Y4_DIN_SRAM14
  PIN Tile_X10Y4_DIN_SRAM15
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2731.480 2263.200 2731.880 ;
    END
  END Tile_X10Y4_DIN_SRAM15
  PIN Tile_X10Y4_DIN_SRAM16
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2734.000 2263.200 2734.400 ;
    END
  END Tile_X10Y4_DIN_SRAM16
  PIN Tile_X10Y4_DIN_SRAM17
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2736.520 2263.200 2736.920 ;
    END
  END Tile_X10Y4_DIN_SRAM17
  PIN Tile_X10Y4_DIN_SRAM18
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2739.040 2263.200 2739.440 ;
    END
  END Tile_X10Y4_DIN_SRAM18
  PIN Tile_X10Y4_DIN_SRAM19
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2741.560 2263.200 2741.960 ;
    END
  END Tile_X10Y4_DIN_SRAM19
  PIN Tile_X10Y4_DIN_SRAM2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2698.720 2263.200 2699.120 ;
    END
  END Tile_X10Y4_DIN_SRAM2
  PIN Tile_X10Y4_DIN_SRAM20
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2744.080 2263.200 2744.480 ;
    END
  END Tile_X10Y4_DIN_SRAM20
  PIN Tile_X10Y4_DIN_SRAM21
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2746.600 2263.200 2747.000 ;
    END
  END Tile_X10Y4_DIN_SRAM21
  PIN Tile_X10Y4_DIN_SRAM22
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2749.120 2263.200 2749.520 ;
    END
  END Tile_X10Y4_DIN_SRAM22
  PIN Tile_X10Y4_DIN_SRAM23
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2751.640 2263.200 2752.040 ;
    END
  END Tile_X10Y4_DIN_SRAM23
  PIN Tile_X10Y4_DIN_SRAM24
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2754.160 2263.200 2754.560 ;
    END
  END Tile_X10Y4_DIN_SRAM24
  PIN Tile_X10Y4_DIN_SRAM25
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2756.680 2263.200 2757.080 ;
    END
  END Tile_X10Y4_DIN_SRAM25
  PIN Tile_X10Y4_DIN_SRAM26
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2759.200 2263.200 2759.600 ;
    END
  END Tile_X10Y4_DIN_SRAM26
  PIN Tile_X10Y4_DIN_SRAM27
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2761.720 2263.200 2762.120 ;
    END
  END Tile_X10Y4_DIN_SRAM27
  PIN Tile_X10Y4_DIN_SRAM28
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2764.240 2263.200 2764.640 ;
    END
  END Tile_X10Y4_DIN_SRAM28
  PIN Tile_X10Y4_DIN_SRAM29
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2766.760 2263.200 2767.160 ;
    END
  END Tile_X10Y4_DIN_SRAM29
  PIN Tile_X10Y4_DIN_SRAM3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2701.240 2263.200 2701.640 ;
    END
  END Tile_X10Y4_DIN_SRAM3
  PIN Tile_X10Y4_DIN_SRAM30
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2769.280 2263.200 2769.680 ;
    END
  END Tile_X10Y4_DIN_SRAM30
  PIN Tile_X10Y4_DIN_SRAM31
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2771.800 2263.200 2772.200 ;
    END
  END Tile_X10Y4_DIN_SRAM31
  PIN Tile_X10Y4_DIN_SRAM4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2703.760 2263.200 2704.160 ;
    END
  END Tile_X10Y4_DIN_SRAM4
  PIN Tile_X10Y4_DIN_SRAM5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2706.280 2263.200 2706.680 ;
    END
  END Tile_X10Y4_DIN_SRAM5
  PIN Tile_X10Y4_DIN_SRAM6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2708.800 2263.200 2709.200 ;
    END
  END Tile_X10Y4_DIN_SRAM6
  PIN Tile_X10Y4_DIN_SRAM7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2711.320 2263.200 2711.720 ;
    END
  END Tile_X10Y4_DIN_SRAM7
  PIN Tile_X10Y4_DIN_SRAM8
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2713.840 2263.200 2714.240 ;
    END
  END Tile_X10Y4_DIN_SRAM8
  PIN Tile_X10Y4_DIN_SRAM9
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2716.360 2263.200 2716.760 ;
    END
  END Tile_X10Y4_DIN_SRAM9
  PIN Tile_X10Y4_DOUT_SRAM0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2504.680 2263.200 2505.080 ;
    END
  END Tile_X10Y4_DOUT_SRAM0
  PIN Tile_X10Y4_DOUT_SRAM1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2507.200 2263.200 2507.600 ;
    END
  END Tile_X10Y4_DOUT_SRAM1
  PIN Tile_X10Y4_DOUT_SRAM10
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2529.880 2263.200 2530.280 ;
    END
  END Tile_X10Y4_DOUT_SRAM10
  PIN Tile_X10Y4_DOUT_SRAM11
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2532.400 2263.200 2532.800 ;
    END
  END Tile_X10Y4_DOUT_SRAM11
  PIN Tile_X10Y4_DOUT_SRAM12
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2534.920 2263.200 2535.320 ;
    END
  END Tile_X10Y4_DOUT_SRAM12
  PIN Tile_X10Y4_DOUT_SRAM13
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2537.440 2263.200 2537.840 ;
    END
  END Tile_X10Y4_DOUT_SRAM13
  PIN Tile_X10Y4_DOUT_SRAM14
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2539.960 2263.200 2540.360 ;
    END
  END Tile_X10Y4_DOUT_SRAM14
  PIN Tile_X10Y4_DOUT_SRAM15
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2542.480 2263.200 2542.880 ;
    END
  END Tile_X10Y4_DOUT_SRAM15
  PIN Tile_X10Y4_DOUT_SRAM16
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2545.000 2263.200 2545.400 ;
    END
  END Tile_X10Y4_DOUT_SRAM16
  PIN Tile_X10Y4_DOUT_SRAM17
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2547.520 2263.200 2547.920 ;
    END
  END Tile_X10Y4_DOUT_SRAM17
  PIN Tile_X10Y4_DOUT_SRAM18
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2550.040 2263.200 2550.440 ;
    END
  END Tile_X10Y4_DOUT_SRAM18
  PIN Tile_X10Y4_DOUT_SRAM19
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2552.560 2263.200 2552.960 ;
    END
  END Tile_X10Y4_DOUT_SRAM19
  PIN Tile_X10Y4_DOUT_SRAM2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2509.720 2263.200 2510.120 ;
    END
  END Tile_X10Y4_DOUT_SRAM2
  PIN Tile_X10Y4_DOUT_SRAM20
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2555.080 2263.200 2555.480 ;
    END
  END Tile_X10Y4_DOUT_SRAM20
  PIN Tile_X10Y4_DOUT_SRAM21
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2557.600 2263.200 2558.000 ;
    END
  END Tile_X10Y4_DOUT_SRAM21
  PIN Tile_X10Y4_DOUT_SRAM22
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2560.120 2263.200 2560.520 ;
    END
  END Tile_X10Y4_DOUT_SRAM22
  PIN Tile_X10Y4_DOUT_SRAM23
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2562.640 2263.200 2563.040 ;
    END
  END Tile_X10Y4_DOUT_SRAM23
  PIN Tile_X10Y4_DOUT_SRAM24
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2565.160 2263.200 2565.560 ;
    END
  END Tile_X10Y4_DOUT_SRAM24
  PIN Tile_X10Y4_DOUT_SRAM25
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2567.680 2263.200 2568.080 ;
    END
  END Tile_X10Y4_DOUT_SRAM25
  PIN Tile_X10Y4_DOUT_SRAM26
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2570.200 2263.200 2570.600 ;
    END
  END Tile_X10Y4_DOUT_SRAM26
  PIN Tile_X10Y4_DOUT_SRAM27
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2572.720 2263.200 2573.120 ;
    END
  END Tile_X10Y4_DOUT_SRAM27
  PIN Tile_X10Y4_DOUT_SRAM28
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2575.240 2263.200 2575.640 ;
    END
  END Tile_X10Y4_DOUT_SRAM28
  PIN Tile_X10Y4_DOUT_SRAM29
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2577.760 2263.200 2578.160 ;
    END
  END Tile_X10Y4_DOUT_SRAM29
  PIN Tile_X10Y4_DOUT_SRAM3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2512.240 2263.200 2512.640 ;
    END
  END Tile_X10Y4_DOUT_SRAM3
  PIN Tile_X10Y4_DOUT_SRAM30
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2580.280 2263.200 2580.680 ;
    END
  END Tile_X10Y4_DOUT_SRAM30
  PIN Tile_X10Y4_DOUT_SRAM31
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2582.800 2263.200 2583.200 ;
    END
  END Tile_X10Y4_DOUT_SRAM31
  PIN Tile_X10Y4_DOUT_SRAM4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2514.760 2263.200 2515.160 ;
    END
  END Tile_X10Y4_DOUT_SRAM4
  PIN Tile_X10Y4_DOUT_SRAM5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2517.280 2263.200 2517.680 ;
    END
  END Tile_X10Y4_DOUT_SRAM5
  PIN Tile_X10Y4_DOUT_SRAM6
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2519.800 2263.200 2520.200 ;
    END
  END Tile_X10Y4_DOUT_SRAM6
  PIN Tile_X10Y4_DOUT_SRAM7
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2522.320 2263.200 2522.720 ;
    END
  END Tile_X10Y4_DOUT_SRAM7
  PIN Tile_X10Y4_DOUT_SRAM8
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2524.840 2263.200 2525.240 ;
    END
  END Tile_X10Y4_DOUT_SRAM8
  PIN Tile_X10Y4_DOUT_SRAM9
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2527.360 2263.200 2527.760 ;
    END
  END Tile_X10Y4_DOUT_SRAM9
  PIN Tile_X10Y4_MEN_SRAM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2774.320 2263.200 2774.720 ;
    END
  END Tile_X10Y4_MEN_SRAM
  PIN Tile_X10Y4_REN_SRAM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2776.840 2263.200 2777.240 ;
    END
  END Tile_X10Y4_REN_SRAM
  PIN Tile_X10Y4_TIE_HIGH_SRAM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.392700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2779.360 2263.200 2779.760 ;
    END
  END Tile_X10Y4_TIE_HIGH_SRAM
  PIN Tile_X10Y4_TIE_LOW_SRAM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2781.880 2263.200 2782.280 ;
    END
  END Tile_X10Y4_TIE_LOW_SRAM
  PIN Tile_X10Y4_WEN_SRAM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2784.400 2263.200 2784.800 ;
    END
  END Tile_X10Y4_WEN_SRAM
  PIN Tile_X10Y6_ADDR_SRAM0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2101.480 2263.200 2101.880 ;
    END
  END Tile_X10Y6_ADDR_SRAM0
  PIN Tile_X10Y6_ADDR_SRAM1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.340 2104.000 2263.200 2104.400 ;
    END
  END Tile_X10Y6_ADDR_SRAM1
  PIN Tile_X10Y6_ADDR_SRAM2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2106.520 2263.200 2106.920 ;
    END
  END Tile_X10Y6_ADDR_SRAM2
  PIN Tile_X10Y6_ADDR_SRAM3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2109.040 2263.200 2109.440 ;
    END
  END Tile_X10Y6_ADDR_SRAM3
  PIN Tile_X10Y6_ADDR_SRAM4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2111.560 2263.200 2111.960 ;
    END
  END Tile_X10Y6_ADDR_SRAM4
  PIN Tile_X10Y6_ADDR_SRAM5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2114.080 2263.200 2114.480 ;
    END
  END Tile_X10Y6_ADDR_SRAM5
  PIN Tile_X10Y6_ADDR_SRAM6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2116.600 2263.200 2117.000 ;
    END
  END Tile_X10Y6_ADDR_SRAM6
  PIN Tile_X10Y6_ADDR_SRAM7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2119.120 2263.200 2119.520 ;
    END
  END Tile_X10Y6_ADDR_SRAM7
  PIN Tile_X10Y6_ADDR_SRAM8
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2121.640 2263.200 2122.040 ;
    END
  END Tile_X10Y6_ADDR_SRAM8
  PIN Tile_X10Y6_ADDR_SRAM9
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2124.160 2263.200 2124.560 ;
    END
  END Tile_X10Y6_ADDR_SRAM9
  PIN Tile_X10Y6_BM_SRAM0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2126.680 2263.200 2127.080 ;
    END
  END Tile_X10Y6_BM_SRAM0
  PIN Tile_X10Y6_BM_SRAM1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2129.200 2263.200 2129.600 ;
    END
  END Tile_X10Y6_BM_SRAM1
  PIN Tile_X10Y6_BM_SRAM10
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2151.880 2263.200 2152.280 ;
    END
  END Tile_X10Y6_BM_SRAM10
  PIN Tile_X10Y6_BM_SRAM11
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2154.400 2263.200 2154.800 ;
    END
  END Tile_X10Y6_BM_SRAM11
  PIN Tile_X10Y6_BM_SRAM12
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2156.920 2263.200 2157.320 ;
    END
  END Tile_X10Y6_BM_SRAM12
  PIN Tile_X10Y6_BM_SRAM13
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2159.440 2263.200 2159.840 ;
    END
  END Tile_X10Y6_BM_SRAM13
  PIN Tile_X10Y6_BM_SRAM14
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2161.960 2263.200 2162.360 ;
    END
  END Tile_X10Y6_BM_SRAM14
  PIN Tile_X10Y6_BM_SRAM15
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2164.480 2263.200 2164.880 ;
    END
  END Tile_X10Y6_BM_SRAM15
  PIN Tile_X10Y6_BM_SRAM16
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2167.000 2263.200 2167.400 ;
    END
  END Tile_X10Y6_BM_SRAM16
  PIN Tile_X10Y6_BM_SRAM17
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2169.520 2263.200 2169.920 ;
    END
  END Tile_X10Y6_BM_SRAM17
  PIN Tile_X10Y6_BM_SRAM18
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2172.040 2263.200 2172.440 ;
    END
  END Tile_X10Y6_BM_SRAM18
  PIN Tile_X10Y6_BM_SRAM19
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2174.560 2263.200 2174.960 ;
    END
  END Tile_X10Y6_BM_SRAM19
  PIN Tile_X10Y6_BM_SRAM2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2131.720 2263.200 2132.120 ;
    END
  END Tile_X10Y6_BM_SRAM2
  PIN Tile_X10Y6_BM_SRAM20
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2177.080 2263.200 2177.480 ;
    END
  END Tile_X10Y6_BM_SRAM20
  PIN Tile_X10Y6_BM_SRAM21
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2179.600 2263.200 2180.000 ;
    END
  END Tile_X10Y6_BM_SRAM21
  PIN Tile_X10Y6_BM_SRAM22
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2182.120 2263.200 2182.520 ;
    END
  END Tile_X10Y6_BM_SRAM22
  PIN Tile_X10Y6_BM_SRAM23
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2184.640 2263.200 2185.040 ;
    END
  END Tile_X10Y6_BM_SRAM23
  PIN Tile_X10Y6_BM_SRAM24
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2187.160 2263.200 2187.560 ;
    END
  END Tile_X10Y6_BM_SRAM24
  PIN Tile_X10Y6_BM_SRAM25
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2189.680 2263.200 2190.080 ;
    END
  END Tile_X10Y6_BM_SRAM25
  PIN Tile_X10Y6_BM_SRAM26
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2192.200 2263.200 2192.600 ;
    END
  END Tile_X10Y6_BM_SRAM26
  PIN Tile_X10Y6_BM_SRAM27
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2194.720 2263.200 2195.120 ;
    END
  END Tile_X10Y6_BM_SRAM27
  PIN Tile_X10Y6_BM_SRAM28
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2197.240 2263.200 2197.640 ;
    END
  END Tile_X10Y6_BM_SRAM28
  PIN Tile_X10Y6_BM_SRAM29
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2199.760 2263.200 2200.160 ;
    END
  END Tile_X10Y6_BM_SRAM29
  PIN Tile_X10Y6_BM_SRAM3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2134.240 2263.200 2134.640 ;
    END
  END Tile_X10Y6_BM_SRAM3
  PIN Tile_X10Y6_BM_SRAM30
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2202.280 2263.200 2202.680 ;
    END
  END Tile_X10Y6_BM_SRAM30
  PIN Tile_X10Y6_BM_SRAM31
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2204.800 2263.200 2205.200 ;
    END
  END Tile_X10Y6_BM_SRAM31
  PIN Tile_X10Y6_BM_SRAM4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2136.760 2263.200 2137.160 ;
    END
  END Tile_X10Y6_BM_SRAM4
  PIN Tile_X10Y6_BM_SRAM5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2139.280 2263.200 2139.680 ;
    END
  END Tile_X10Y6_BM_SRAM5
  PIN Tile_X10Y6_BM_SRAM6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2141.800 2263.200 2142.200 ;
    END
  END Tile_X10Y6_BM_SRAM6
  PIN Tile_X10Y6_BM_SRAM7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2144.320 2263.200 2144.720 ;
    END
  END Tile_X10Y6_BM_SRAM7
  PIN Tile_X10Y6_BM_SRAM8
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2146.840 2263.200 2147.240 ;
    END
  END Tile_X10Y6_BM_SRAM8
  PIN Tile_X10Y6_BM_SRAM9
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2149.360 2263.200 2149.760 ;
    END
  END Tile_X10Y6_BM_SRAM9
  PIN Tile_X10Y6_CLK_SRAM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2207.320 2263.200 2207.720 ;
    END
  END Tile_X10Y6_CLK_SRAM
  PIN Tile_X10Y6_CONFIGURED_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2018.320 2263.200 2018.720 ;
    END
  END Tile_X10Y6_CONFIGURED_top
  PIN Tile_X10Y6_DIN_SRAM0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2209.840 2263.200 2210.240 ;
    END
  END Tile_X10Y6_DIN_SRAM0
  PIN Tile_X10Y6_DIN_SRAM1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2212.360 2263.200 2212.760 ;
    END
  END Tile_X10Y6_DIN_SRAM1
  PIN Tile_X10Y6_DIN_SRAM10
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2235.040 2263.200 2235.440 ;
    END
  END Tile_X10Y6_DIN_SRAM10
  PIN Tile_X10Y6_DIN_SRAM11
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2237.560 2263.200 2237.960 ;
    END
  END Tile_X10Y6_DIN_SRAM11
  PIN Tile_X10Y6_DIN_SRAM12
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2240.080 2263.200 2240.480 ;
    END
  END Tile_X10Y6_DIN_SRAM12
  PIN Tile_X10Y6_DIN_SRAM13
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2242.600 2263.200 2243.000 ;
    END
  END Tile_X10Y6_DIN_SRAM13
  PIN Tile_X10Y6_DIN_SRAM14
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2245.120 2263.200 2245.520 ;
    END
  END Tile_X10Y6_DIN_SRAM14
  PIN Tile_X10Y6_DIN_SRAM15
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2247.640 2263.200 2248.040 ;
    END
  END Tile_X10Y6_DIN_SRAM15
  PIN Tile_X10Y6_DIN_SRAM16
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2250.160 2263.200 2250.560 ;
    END
  END Tile_X10Y6_DIN_SRAM16
  PIN Tile_X10Y6_DIN_SRAM17
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2252.680 2263.200 2253.080 ;
    END
  END Tile_X10Y6_DIN_SRAM17
  PIN Tile_X10Y6_DIN_SRAM18
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2255.200 2263.200 2255.600 ;
    END
  END Tile_X10Y6_DIN_SRAM18
  PIN Tile_X10Y6_DIN_SRAM19
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2257.720 2263.200 2258.120 ;
    END
  END Tile_X10Y6_DIN_SRAM19
  PIN Tile_X10Y6_DIN_SRAM2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2214.880 2263.200 2215.280 ;
    END
  END Tile_X10Y6_DIN_SRAM2
  PIN Tile_X10Y6_DIN_SRAM20
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2260.240 2263.200 2260.640 ;
    END
  END Tile_X10Y6_DIN_SRAM20
  PIN Tile_X10Y6_DIN_SRAM21
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2262.760 2263.200 2263.160 ;
    END
  END Tile_X10Y6_DIN_SRAM21
  PIN Tile_X10Y6_DIN_SRAM22
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2265.280 2263.200 2265.680 ;
    END
  END Tile_X10Y6_DIN_SRAM22
  PIN Tile_X10Y6_DIN_SRAM23
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2267.800 2263.200 2268.200 ;
    END
  END Tile_X10Y6_DIN_SRAM23
  PIN Tile_X10Y6_DIN_SRAM24
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2270.320 2263.200 2270.720 ;
    END
  END Tile_X10Y6_DIN_SRAM24
  PIN Tile_X10Y6_DIN_SRAM25
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2272.840 2263.200 2273.240 ;
    END
  END Tile_X10Y6_DIN_SRAM25
  PIN Tile_X10Y6_DIN_SRAM26
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2275.360 2263.200 2275.760 ;
    END
  END Tile_X10Y6_DIN_SRAM26
  PIN Tile_X10Y6_DIN_SRAM27
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2277.880 2263.200 2278.280 ;
    END
  END Tile_X10Y6_DIN_SRAM27
  PIN Tile_X10Y6_DIN_SRAM28
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2280.400 2263.200 2280.800 ;
    END
  END Tile_X10Y6_DIN_SRAM28
  PIN Tile_X10Y6_DIN_SRAM29
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2282.920 2263.200 2283.320 ;
    END
  END Tile_X10Y6_DIN_SRAM29
  PIN Tile_X10Y6_DIN_SRAM3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2217.400 2263.200 2217.800 ;
    END
  END Tile_X10Y6_DIN_SRAM3
  PIN Tile_X10Y6_DIN_SRAM30
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2285.440 2263.200 2285.840 ;
    END
  END Tile_X10Y6_DIN_SRAM30
  PIN Tile_X10Y6_DIN_SRAM31
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2287.960 2263.200 2288.360 ;
    END
  END Tile_X10Y6_DIN_SRAM31
  PIN Tile_X10Y6_DIN_SRAM4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2219.920 2263.200 2220.320 ;
    END
  END Tile_X10Y6_DIN_SRAM4
  PIN Tile_X10Y6_DIN_SRAM5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2222.440 2263.200 2222.840 ;
    END
  END Tile_X10Y6_DIN_SRAM5
  PIN Tile_X10Y6_DIN_SRAM6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2224.960 2263.200 2225.360 ;
    END
  END Tile_X10Y6_DIN_SRAM6
  PIN Tile_X10Y6_DIN_SRAM7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2227.480 2263.200 2227.880 ;
    END
  END Tile_X10Y6_DIN_SRAM7
  PIN Tile_X10Y6_DIN_SRAM8
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2230.000 2263.200 2230.400 ;
    END
  END Tile_X10Y6_DIN_SRAM8
  PIN Tile_X10Y6_DIN_SRAM9
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2232.520 2263.200 2232.920 ;
    END
  END Tile_X10Y6_DIN_SRAM9
  PIN Tile_X10Y6_DOUT_SRAM0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2020.840 2263.200 2021.240 ;
    END
  END Tile_X10Y6_DOUT_SRAM0
  PIN Tile_X10Y6_DOUT_SRAM1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2023.360 2263.200 2023.760 ;
    END
  END Tile_X10Y6_DOUT_SRAM1
  PIN Tile_X10Y6_DOUT_SRAM10
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2046.040 2263.200 2046.440 ;
    END
  END Tile_X10Y6_DOUT_SRAM10
  PIN Tile_X10Y6_DOUT_SRAM11
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2048.560 2263.200 2048.960 ;
    END
  END Tile_X10Y6_DOUT_SRAM11
  PIN Tile_X10Y6_DOUT_SRAM12
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2051.080 2263.200 2051.480 ;
    END
  END Tile_X10Y6_DOUT_SRAM12
  PIN Tile_X10Y6_DOUT_SRAM13
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2053.600 2263.200 2054.000 ;
    END
  END Tile_X10Y6_DOUT_SRAM13
  PIN Tile_X10Y6_DOUT_SRAM14
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2056.120 2263.200 2056.520 ;
    END
  END Tile_X10Y6_DOUT_SRAM14
  PIN Tile_X10Y6_DOUT_SRAM15
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2058.640 2263.200 2059.040 ;
    END
  END Tile_X10Y6_DOUT_SRAM15
  PIN Tile_X10Y6_DOUT_SRAM16
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2061.160 2263.200 2061.560 ;
    END
  END Tile_X10Y6_DOUT_SRAM16
  PIN Tile_X10Y6_DOUT_SRAM17
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2063.680 2263.200 2064.080 ;
    END
  END Tile_X10Y6_DOUT_SRAM17
  PIN Tile_X10Y6_DOUT_SRAM18
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2066.200 2263.200 2066.600 ;
    END
  END Tile_X10Y6_DOUT_SRAM18
  PIN Tile_X10Y6_DOUT_SRAM19
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2068.720 2263.200 2069.120 ;
    END
  END Tile_X10Y6_DOUT_SRAM19
  PIN Tile_X10Y6_DOUT_SRAM2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2025.880 2263.200 2026.280 ;
    END
  END Tile_X10Y6_DOUT_SRAM2
  PIN Tile_X10Y6_DOUT_SRAM20
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2071.240 2263.200 2071.640 ;
    END
  END Tile_X10Y6_DOUT_SRAM20
  PIN Tile_X10Y6_DOUT_SRAM21
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2073.760 2263.200 2074.160 ;
    END
  END Tile_X10Y6_DOUT_SRAM21
  PIN Tile_X10Y6_DOUT_SRAM22
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2076.280 2263.200 2076.680 ;
    END
  END Tile_X10Y6_DOUT_SRAM22
  PIN Tile_X10Y6_DOUT_SRAM23
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2078.800 2263.200 2079.200 ;
    END
  END Tile_X10Y6_DOUT_SRAM23
  PIN Tile_X10Y6_DOUT_SRAM24
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2081.320 2263.200 2081.720 ;
    END
  END Tile_X10Y6_DOUT_SRAM24
  PIN Tile_X10Y6_DOUT_SRAM25
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2083.840 2263.200 2084.240 ;
    END
  END Tile_X10Y6_DOUT_SRAM25
  PIN Tile_X10Y6_DOUT_SRAM26
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2086.360 2263.200 2086.760 ;
    END
  END Tile_X10Y6_DOUT_SRAM26
  PIN Tile_X10Y6_DOUT_SRAM27
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2088.880 2263.200 2089.280 ;
    END
  END Tile_X10Y6_DOUT_SRAM27
  PIN Tile_X10Y6_DOUT_SRAM28
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2091.400 2263.200 2091.800 ;
    END
  END Tile_X10Y6_DOUT_SRAM28
  PIN Tile_X10Y6_DOUT_SRAM29
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2093.920 2263.200 2094.320 ;
    END
  END Tile_X10Y6_DOUT_SRAM29
  PIN Tile_X10Y6_DOUT_SRAM3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2028.400 2263.200 2028.800 ;
    END
  END Tile_X10Y6_DOUT_SRAM3
  PIN Tile_X10Y6_DOUT_SRAM30
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2096.440 2263.200 2096.840 ;
    END
  END Tile_X10Y6_DOUT_SRAM30
  PIN Tile_X10Y6_DOUT_SRAM31
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2098.960 2263.200 2099.360 ;
    END
  END Tile_X10Y6_DOUT_SRAM31
  PIN Tile_X10Y6_DOUT_SRAM4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2030.920 2263.200 2031.320 ;
    END
  END Tile_X10Y6_DOUT_SRAM4
  PIN Tile_X10Y6_DOUT_SRAM5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2033.440 2263.200 2033.840 ;
    END
  END Tile_X10Y6_DOUT_SRAM5
  PIN Tile_X10Y6_DOUT_SRAM6
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2035.960 2263.200 2036.360 ;
    END
  END Tile_X10Y6_DOUT_SRAM6
  PIN Tile_X10Y6_DOUT_SRAM7
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2038.480 2263.200 2038.880 ;
    END
  END Tile_X10Y6_DOUT_SRAM7
  PIN Tile_X10Y6_DOUT_SRAM8
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2041.000 2263.200 2041.400 ;
    END
  END Tile_X10Y6_DOUT_SRAM8
  PIN Tile_X10Y6_DOUT_SRAM9
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2043.520 2263.200 2043.920 ;
    END
  END Tile_X10Y6_DOUT_SRAM9
  PIN Tile_X10Y6_MEN_SRAM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2290.480 2263.200 2290.880 ;
    END
  END Tile_X10Y6_MEN_SRAM
  PIN Tile_X10Y6_REN_SRAM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2293.000 2263.200 2293.400 ;
    END
  END Tile_X10Y6_REN_SRAM
  PIN Tile_X10Y6_TIE_HIGH_SRAM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.392700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2295.520 2263.200 2295.920 ;
    END
  END Tile_X10Y6_TIE_HIGH_SRAM
  PIN Tile_X10Y6_TIE_LOW_SRAM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2298.040 2263.200 2298.440 ;
    END
  END Tile_X10Y6_TIE_LOW_SRAM
  PIN Tile_X10Y6_WEN_SRAM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 2300.560 2263.200 2300.960 ;
    END
  END Tile_X10Y6_WEN_SRAM
  PIN Tile_X10Y8_ADDR_SRAM0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1617.640 2263.200 1618.040 ;
    END
  END Tile_X10Y8_ADDR_SRAM0
  PIN Tile_X10Y8_ADDR_SRAM1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.340 1620.160 2263.200 1620.560 ;
    END
  END Tile_X10Y8_ADDR_SRAM1
  PIN Tile_X10Y8_ADDR_SRAM2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1622.680 2263.200 1623.080 ;
    END
  END Tile_X10Y8_ADDR_SRAM2
  PIN Tile_X10Y8_ADDR_SRAM3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1625.200 2263.200 1625.600 ;
    END
  END Tile_X10Y8_ADDR_SRAM3
  PIN Tile_X10Y8_ADDR_SRAM4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1627.720 2263.200 1628.120 ;
    END
  END Tile_X10Y8_ADDR_SRAM4
  PIN Tile_X10Y8_ADDR_SRAM5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1630.240 2263.200 1630.640 ;
    END
  END Tile_X10Y8_ADDR_SRAM5
  PIN Tile_X10Y8_ADDR_SRAM6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1632.760 2263.200 1633.160 ;
    END
  END Tile_X10Y8_ADDR_SRAM6
  PIN Tile_X10Y8_ADDR_SRAM7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1635.280 2263.200 1635.680 ;
    END
  END Tile_X10Y8_ADDR_SRAM7
  PIN Tile_X10Y8_ADDR_SRAM8
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1637.800 2263.200 1638.200 ;
    END
  END Tile_X10Y8_ADDR_SRAM8
  PIN Tile_X10Y8_ADDR_SRAM9
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1640.320 2263.200 1640.720 ;
    END
  END Tile_X10Y8_ADDR_SRAM9
  PIN Tile_X10Y8_BM_SRAM0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1642.840 2263.200 1643.240 ;
    END
  END Tile_X10Y8_BM_SRAM0
  PIN Tile_X10Y8_BM_SRAM1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1645.360 2263.200 1645.760 ;
    END
  END Tile_X10Y8_BM_SRAM1
  PIN Tile_X10Y8_BM_SRAM10
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1668.040 2263.200 1668.440 ;
    END
  END Tile_X10Y8_BM_SRAM10
  PIN Tile_X10Y8_BM_SRAM11
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1670.560 2263.200 1670.960 ;
    END
  END Tile_X10Y8_BM_SRAM11
  PIN Tile_X10Y8_BM_SRAM12
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1673.080 2263.200 1673.480 ;
    END
  END Tile_X10Y8_BM_SRAM12
  PIN Tile_X10Y8_BM_SRAM13
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1675.600 2263.200 1676.000 ;
    END
  END Tile_X10Y8_BM_SRAM13
  PIN Tile_X10Y8_BM_SRAM14
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1678.120 2263.200 1678.520 ;
    END
  END Tile_X10Y8_BM_SRAM14
  PIN Tile_X10Y8_BM_SRAM15
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1680.640 2263.200 1681.040 ;
    END
  END Tile_X10Y8_BM_SRAM15
  PIN Tile_X10Y8_BM_SRAM16
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1683.160 2263.200 1683.560 ;
    END
  END Tile_X10Y8_BM_SRAM16
  PIN Tile_X10Y8_BM_SRAM17
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1685.680 2263.200 1686.080 ;
    END
  END Tile_X10Y8_BM_SRAM17
  PIN Tile_X10Y8_BM_SRAM18
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1688.200 2263.200 1688.600 ;
    END
  END Tile_X10Y8_BM_SRAM18
  PIN Tile_X10Y8_BM_SRAM19
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1690.720 2263.200 1691.120 ;
    END
  END Tile_X10Y8_BM_SRAM19
  PIN Tile_X10Y8_BM_SRAM2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1647.880 2263.200 1648.280 ;
    END
  END Tile_X10Y8_BM_SRAM2
  PIN Tile_X10Y8_BM_SRAM20
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1693.240 2263.200 1693.640 ;
    END
  END Tile_X10Y8_BM_SRAM20
  PIN Tile_X10Y8_BM_SRAM21
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1695.760 2263.200 1696.160 ;
    END
  END Tile_X10Y8_BM_SRAM21
  PIN Tile_X10Y8_BM_SRAM22
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1698.280 2263.200 1698.680 ;
    END
  END Tile_X10Y8_BM_SRAM22
  PIN Tile_X10Y8_BM_SRAM23
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1700.800 2263.200 1701.200 ;
    END
  END Tile_X10Y8_BM_SRAM23
  PIN Tile_X10Y8_BM_SRAM24
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1703.320 2263.200 1703.720 ;
    END
  END Tile_X10Y8_BM_SRAM24
  PIN Tile_X10Y8_BM_SRAM25
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1705.840 2263.200 1706.240 ;
    END
  END Tile_X10Y8_BM_SRAM25
  PIN Tile_X10Y8_BM_SRAM26
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1708.360 2263.200 1708.760 ;
    END
  END Tile_X10Y8_BM_SRAM26
  PIN Tile_X10Y8_BM_SRAM27
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1710.880 2263.200 1711.280 ;
    END
  END Tile_X10Y8_BM_SRAM27
  PIN Tile_X10Y8_BM_SRAM28
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1713.400 2263.200 1713.800 ;
    END
  END Tile_X10Y8_BM_SRAM28
  PIN Tile_X10Y8_BM_SRAM29
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1715.920 2263.200 1716.320 ;
    END
  END Tile_X10Y8_BM_SRAM29
  PIN Tile_X10Y8_BM_SRAM3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1650.400 2263.200 1650.800 ;
    END
  END Tile_X10Y8_BM_SRAM3
  PIN Tile_X10Y8_BM_SRAM30
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1718.440 2263.200 1718.840 ;
    END
  END Tile_X10Y8_BM_SRAM30
  PIN Tile_X10Y8_BM_SRAM31
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1720.960 2263.200 1721.360 ;
    END
  END Tile_X10Y8_BM_SRAM31
  PIN Tile_X10Y8_BM_SRAM4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1652.920 2263.200 1653.320 ;
    END
  END Tile_X10Y8_BM_SRAM4
  PIN Tile_X10Y8_BM_SRAM5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1655.440 2263.200 1655.840 ;
    END
  END Tile_X10Y8_BM_SRAM5
  PIN Tile_X10Y8_BM_SRAM6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1657.960 2263.200 1658.360 ;
    END
  END Tile_X10Y8_BM_SRAM6
  PIN Tile_X10Y8_BM_SRAM7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1660.480 2263.200 1660.880 ;
    END
  END Tile_X10Y8_BM_SRAM7
  PIN Tile_X10Y8_BM_SRAM8
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1663.000 2263.200 1663.400 ;
    END
  END Tile_X10Y8_BM_SRAM8
  PIN Tile_X10Y8_BM_SRAM9
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1665.520 2263.200 1665.920 ;
    END
  END Tile_X10Y8_BM_SRAM9
  PIN Tile_X10Y8_CLK_SRAM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1723.480 2263.200 1723.880 ;
    END
  END Tile_X10Y8_CLK_SRAM
  PIN Tile_X10Y8_CONFIGURED_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1534.480 2263.200 1534.880 ;
    END
  END Tile_X10Y8_CONFIGURED_top
  PIN Tile_X10Y8_DIN_SRAM0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1726.000 2263.200 1726.400 ;
    END
  END Tile_X10Y8_DIN_SRAM0
  PIN Tile_X10Y8_DIN_SRAM1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1728.520 2263.200 1728.920 ;
    END
  END Tile_X10Y8_DIN_SRAM1
  PIN Tile_X10Y8_DIN_SRAM10
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1751.200 2263.200 1751.600 ;
    END
  END Tile_X10Y8_DIN_SRAM10
  PIN Tile_X10Y8_DIN_SRAM11
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1753.720 2263.200 1754.120 ;
    END
  END Tile_X10Y8_DIN_SRAM11
  PIN Tile_X10Y8_DIN_SRAM12
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1756.240 2263.200 1756.640 ;
    END
  END Tile_X10Y8_DIN_SRAM12
  PIN Tile_X10Y8_DIN_SRAM13
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1758.760 2263.200 1759.160 ;
    END
  END Tile_X10Y8_DIN_SRAM13
  PIN Tile_X10Y8_DIN_SRAM14
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1761.280 2263.200 1761.680 ;
    END
  END Tile_X10Y8_DIN_SRAM14
  PIN Tile_X10Y8_DIN_SRAM15
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1763.800 2263.200 1764.200 ;
    END
  END Tile_X10Y8_DIN_SRAM15
  PIN Tile_X10Y8_DIN_SRAM16
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1766.320 2263.200 1766.720 ;
    END
  END Tile_X10Y8_DIN_SRAM16
  PIN Tile_X10Y8_DIN_SRAM17
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1768.840 2263.200 1769.240 ;
    END
  END Tile_X10Y8_DIN_SRAM17
  PIN Tile_X10Y8_DIN_SRAM18
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1771.360 2263.200 1771.760 ;
    END
  END Tile_X10Y8_DIN_SRAM18
  PIN Tile_X10Y8_DIN_SRAM19
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1773.880 2263.200 1774.280 ;
    END
  END Tile_X10Y8_DIN_SRAM19
  PIN Tile_X10Y8_DIN_SRAM2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1731.040 2263.200 1731.440 ;
    END
  END Tile_X10Y8_DIN_SRAM2
  PIN Tile_X10Y8_DIN_SRAM20
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1776.400 2263.200 1776.800 ;
    END
  END Tile_X10Y8_DIN_SRAM20
  PIN Tile_X10Y8_DIN_SRAM21
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1778.920 2263.200 1779.320 ;
    END
  END Tile_X10Y8_DIN_SRAM21
  PIN Tile_X10Y8_DIN_SRAM22
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1781.440 2263.200 1781.840 ;
    END
  END Tile_X10Y8_DIN_SRAM22
  PIN Tile_X10Y8_DIN_SRAM23
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1783.960 2263.200 1784.360 ;
    END
  END Tile_X10Y8_DIN_SRAM23
  PIN Tile_X10Y8_DIN_SRAM24
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1786.480 2263.200 1786.880 ;
    END
  END Tile_X10Y8_DIN_SRAM24
  PIN Tile_X10Y8_DIN_SRAM25
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1789.000 2263.200 1789.400 ;
    END
  END Tile_X10Y8_DIN_SRAM25
  PIN Tile_X10Y8_DIN_SRAM26
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1791.520 2263.200 1791.920 ;
    END
  END Tile_X10Y8_DIN_SRAM26
  PIN Tile_X10Y8_DIN_SRAM27
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1794.040 2263.200 1794.440 ;
    END
  END Tile_X10Y8_DIN_SRAM27
  PIN Tile_X10Y8_DIN_SRAM28
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1796.560 2263.200 1796.960 ;
    END
  END Tile_X10Y8_DIN_SRAM28
  PIN Tile_X10Y8_DIN_SRAM29
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1799.080 2263.200 1799.480 ;
    END
  END Tile_X10Y8_DIN_SRAM29
  PIN Tile_X10Y8_DIN_SRAM3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1733.560 2263.200 1733.960 ;
    END
  END Tile_X10Y8_DIN_SRAM3
  PIN Tile_X10Y8_DIN_SRAM30
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1801.600 2263.200 1802.000 ;
    END
  END Tile_X10Y8_DIN_SRAM30
  PIN Tile_X10Y8_DIN_SRAM31
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1804.120 2263.200 1804.520 ;
    END
  END Tile_X10Y8_DIN_SRAM31
  PIN Tile_X10Y8_DIN_SRAM4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1736.080 2263.200 1736.480 ;
    END
  END Tile_X10Y8_DIN_SRAM4
  PIN Tile_X10Y8_DIN_SRAM5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1738.600 2263.200 1739.000 ;
    END
  END Tile_X10Y8_DIN_SRAM5
  PIN Tile_X10Y8_DIN_SRAM6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1741.120 2263.200 1741.520 ;
    END
  END Tile_X10Y8_DIN_SRAM6
  PIN Tile_X10Y8_DIN_SRAM7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1743.640 2263.200 1744.040 ;
    END
  END Tile_X10Y8_DIN_SRAM7
  PIN Tile_X10Y8_DIN_SRAM8
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1746.160 2263.200 1746.560 ;
    END
  END Tile_X10Y8_DIN_SRAM8
  PIN Tile_X10Y8_DIN_SRAM9
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1748.680 2263.200 1749.080 ;
    END
  END Tile_X10Y8_DIN_SRAM9
  PIN Tile_X10Y8_DOUT_SRAM0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1537.000 2263.200 1537.400 ;
    END
  END Tile_X10Y8_DOUT_SRAM0
  PIN Tile_X10Y8_DOUT_SRAM1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1539.520 2263.200 1539.920 ;
    END
  END Tile_X10Y8_DOUT_SRAM1
  PIN Tile_X10Y8_DOUT_SRAM10
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1562.200 2263.200 1562.600 ;
    END
  END Tile_X10Y8_DOUT_SRAM10
  PIN Tile_X10Y8_DOUT_SRAM11
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1564.720 2263.200 1565.120 ;
    END
  END Tile_X10Y8_DOUT_SRAM11
  PIN Tile_X10Y8_DOUT_SRAM12
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1567.240 2263.200 1567.640 ;
    END
  END Tile_X10Y8_DOUT_SRAM12
  PIN Tile_X10Y8_DOUT_SRAM13
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1569.760 2263.200 1570.160 ;
    END
  END Tile_X10Y8_DOUT_SRAM13
  PIN Tile_X10Y8_DOUT_SRAM14
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1572.280 2263.200 1572.680 ;
    END
  END Tile_X10Y8_DOUT_SRAM14
  PIN Tile_X10Y8_DOUT_SRAM15
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1574.800 2263.200 1575.200 ;
    END
  END Tile_X10Y8_DOUT_SRAM15
  PIN Tile_X10Y8_DOUT_SRAM16
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1577.320 2263.200 1577.720 ;
    END
  END Tile_X10Y8_DOUT_SRAM16
  PIN Tile_X10Y8_DOUT_SRAM17
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1579.840 2263.200 1580.240 ;
    END
  END Tile_X10Y8_DOUT_SRAM17
  PIN Tile_X10Y8_DOUT_SRAM18
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1582.360 2263.200 1582.760 ;
    END
  END Tile_X10Y8_DOUT_SRAM18
  PIN Tile_X10Y8_DOUT_SRAM19
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1584.880 2263.200 1585.280 ;
    END
  END Tile_X10Y8_DOUT_SRAM19
  PIN Tile_X10Y8_DOUT_SRAM2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1542.040 2263.200 1542.440 ;
    END
  END Tile_X10Y8_DOUT_SRAM2
  PIN Tile_X10Y8_DOUT_SRAM20
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1587.400 2263.200 1587.800 ;
    END
  END Tile_X10Y8_DOUT_SRAM20
  PIN Tile_X10Y8_DOUT_SRAM21
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1589.920 2263.200 1590.320 ;
    END
  END Tile_X10Y8_DOUT_SRAM21
  PIN Tile_X10Y8_DOUT_SRAM22
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1592.440 2263.200 1592.840 ;
    END
  END Tile_X10Y8_DOUT_SRAM22
  PIN Tile_X10Y8_DOUT_SRAM23
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1594.960 2263.200 1595.360 ;
    END
  END Tile_X10Y8_DOUT_SRAM23
  PIN Tile_X10Y8_DOUT_SRAM24
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1597.480 2263.200 1597.880 ;
    END
  END Tile_X10Y8_DOUT_SRAM24
  PIN Tile_X10Y8_DOUT_SRAM25
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1600.000 2263.200 1600.400 ;
    END
  END Tile_X10Y8_DOUT_SRAM25
  PIN Tile_X10Y8_DOUT_SRAM26
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1602.520 2263.200 1602.920 ;
    END
  END Tile_X10Y8_DOUT_SRAM26
  PIN Tile_X10Y8_DOUT_SRAM27
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1605.040 2263.200 1605.440 ;
    END
  END Tile_X10Y8_DOUT_SRAM27
  PIN Tile_X10Y8_DOUT_SRAM28
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1607.560 2263.200 1607.960 ;
    END
  END Tile_X10Y8_DOUT_SRAM28
  PIN Tile_X10Y8_DOUT_SRAM29
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1610.080 2263.200 1610.480 ;
    END
  END Tile_X10Y8_DOUT_SRAM29
  PIN Tile_X10Y8_DOUT_SRAM3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1544.560 2263.200 1544.960 ;
    END
  END Tile_X10Y8_DOUT_SRAM3
  PIN Tile_X10Y8_DOUT_SRAM30
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1612.600 2263.200 1613.000 ;
    END
  END Tile_X10Y8_DOUT_SRAM30
  PIN Tile_X10Y8_DOUT_SRAM31
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1615.120 2263.200 1615.520 ;
    END
  END Tile_X10Y8_DOUT_SRAM31
  PIN Tile_X10Y8_DOUT_SRAM4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1547.080 2263.200 1547.480 ;
    END
  END Tile_X10Y8_DOUT_SRAM4
  PIN Tile_X10Y8_DOUT_SRAM5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1549.600 2263.200 1550.000 ;
    END
  END Tile_X10Y8_DOUT_SRAM5
  PIN Tile_X10Y8_DOUT_SRAM6
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1552.120 2263.200 1552.520 ;
    END
  END Tile_X10Y8_DOUT_SRAM6
  PIN Tile_X10Y8_DOUT_SRAM7
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1554.640 2263.200 1555.040 ;
    END
  END Tile_X10Y8_DOUT_SRAM7
  PIN Tile_X10Y8_DOUT_SRAM8
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1557.160 2263.200 1557.560 ;
    END
  END Tile_X10Y8_DOUT_SRAM8
  PIN Tile_X10Y8_DOUT_SRAM9
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1559.680 2263.200 1560.080 ;
    END
  END Tile_X10Y8_DOUT_SRAM9
  PIN Tile_X10Y8_MEN_SRAM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1806.640 2263.200 1807.040 ;
    END
  END Tile_X10Y8_MEN_SRAM
  PIN Tile_X10Y8_REN_SRAM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1809.160 2263.200 1809.560 ;
    END
  END Tile_X10Y8_REN_SRAM
  PIN Tile_X10Y8_TIE_HIGH_SRAM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.392700 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1811.680 2263.200 1812.080 ;
    END
  END Tile_X10Y8_TIE_HIGH_SRAM
  PIN Tile_X10Y8_TIE_LOW_SRAM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1814.200 2263.200 1814.600 ;
    END
  END Tile_X10Y8_TIE_LOW_SRAM
  PIN Tile_X10Y8_WEN_SRAM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 2262.270 1816.720 2263.200 1817.120 ;
    END
  END Tile_X10Y8_WEN_SRAM
  PIN Tile_X1Y0_A_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 92.440 3510.800 92.840 3511.680 ;
    END
  END Tile_X1Y0_A_I_top
  PIN Tile_X1Y0_A_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 86.680 3510.800 87.080 3511.680 ;
    END
  END Tile_X1Y0_A_O_top
  PIN Tile_X1Y0_A_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 98.200 3510.800 98.600 3511.680 ;
    END
  END Tile_X1Y0_A_T_top
  PIN Tile_X1Y0_A_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 121.240 3510.800 121.640 3511.680 ;
    END
  END Tile_X1Y0_A_config_C_bit0
  PIN Tile_X1Y0_A_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 127.000 3510.800 127.400 3511.680 ;
    END
  END Tile_X1Y0_A_config_C_bit1
  PIN Tile_X1Y0_A_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 132.760 3510.800 133.160 3511.680 ;
    END
  END Tile_X1Y0_A_config_C_bit2
  PIN Tile_X1Y0_A_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 138.520 3510.800 138.920 3511.680 ;
    END
  END Tile_X1Y0_A_config_C_bit3
  PIN Tile_X1Y0_B_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 109.720 3510.800 110.120 3511.680 ;
    END
  END Tile_X1Y0_B_I_top
  PIN Tile_X1Y0_B_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 103.960 3510.800 104.360 3511.680 ;
    END
  END Tile_X1Y0_B_O_top
  PIN Tile_X1Y0_B_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 115.480 3510.800 115.880 3511.680 ;
    END
  END Tile_X1Y0_B_T_top
  PIN Tile_X1Y0_B_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 144.280 3510.800 144.680 3511.680 ;
    END
  END Tile_X1Y0_B_config_C_bit0
  PIN Tile_X1Y0_B_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 150.040 3510.800 150.440 3511.680 ;
    END
  END Tile_X1Y0_B_config_C_bit1
  PIN Tile_X1Y0_B_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 155.800 3510.800 156.200 3511.680 ;
    END
  END Tile_X1Y0_B_config_C_bit2
  PIN Tile_X1Y0_B_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 161.560 3510.800 161.960 3511.680 ;
    END
  END Tile_X1Y0_B_config_C_bit3
  PIN Tile_X2Y0_A_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 324.280 3510.800 324.680 3511.680 ;
    END
  END Tile_X2Y0_A_I_top
  PIN Tile_X2Y0_A_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 318.520 3510.800 318.920 3511.680 ;
    END
  END Tile_X2Y0_A_O_top
  PIN Tile_X2Y0_A_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 330.040 3510.800 330.440 3511.680 ;
    END
  END Tile_X2Y0_A_T_top
  PIN Tile_X2Y0_A_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 353.080 3510.800 353.480 3511.680 ;
    END
  END Tile_X2Y0_A_config_C_bit0
  PIN Tile_X2Y0_A_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 358.840 3510.800 359.240 3511.680 ;
    END
  END Tile_X2Y0_A_config_C_bit1
  PIN Tile_X2Y0_A_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 364.600 3510.800 365.000 3511.680 ;
    END
  END Tile_X2Y0_A_config_C_bit2
  PIN Tile_X2Y0_A_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 370.360 3510.800 370.760 3511.680 ;
    END
  END Tile_X2Y0_A_config_C_bit3
  PIN Tile_X2Y0_B_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 341.560 3510.800 341.960 3511.680 ;
    END
  END Tile_X2Y0_B_I_top
  PIN Tile_X2Y0_B_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 335.800 3510.800 336.200 3511.680 ;
    END
  END Tile_X2Y0_B_O_top
  PIN Tile_X2Y0_B_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 347.320 3510.800 347.720 3511.680 ;
    END
  END Tile_X2Y0_B_T_top
  PIN Tile_X2Y0_B_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 376.120 3510.800 376.520 3511.680 ;
    END
  END Tile_X2Y0_B_config_C_bit0
  PIN Tile_X2Y0_B_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 381.880 3510.800 382.280 3511.680 ;
    END
  END Tile_X2Y0_B_config_C_bit1
  PIN Tile_X2Y0_B_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 387.640 3510.800 388.040 3511.680 ;
    END
  END Tile_X2Y0_B_config_C_bit2
  PIN Tile_X2Y0_B_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 393.400 3510.800 393.800 3511.680 ;
    END
  END Tile_X2Y0_B_config_C_bit3
  PIN Tile_X2Y15_BOOT_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 328.120 0.000 328.520 0.480 ;
    END
  END Tile_X2Y15_BOOT_top
  PIN Tile_X2Y15_CONFIGURED_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 312.760 0.000 313.160 0.480 ;
    END
  END Tile_X2Y15_CONFIGURED_top
  PIN Tile_X2Y15_RESET_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 320.440 0.000 320.840 0.480 ;
    END
  END Tile_X2Y15_RESET_top
  PIN Tile_X2Y15_SLOT_top0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 335.800 0.000 336.200 0.480 ;
    END
  END Tile_X2Y15_SLOT_top0
  PIN Tile_X2Y15_SLOT_top1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 343.480 0.000 343.880 0.480 ;
    END
  END Tile_X2Y15_SLOT_top1
  PIN Tile_X2Y15_SLOT_top2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 351.160 0.000 351.560 0.480 ;
    END
  END Tile_X2Y15_SLOT_top2
  PIN Tile_X2Y15_SLOT_top3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 358.840 0.000 359.240 0.480 ;
    END
  END Tile_X2Y15_SLOT_top3
  PIN Tile_X3Y15_CONFIGURED_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 539.800 0.000 540.200 0.480 ;
    END
  END Tile_X3Y15_CONFIGURED_top
  PIN Tile_X3Y15_IRQ_top0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 548.440 0.000 548.840 0.480 ;
    END
  END Tile_X3Y15_IRQ_top0
  PIN Tile_X3Y15_IRQ_top1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 557.080 0.000 557.480 0.480 ;
    END
  END Tile_X3Y15_IRQ_top1
  PIN Tile_X3Y15_IRQ_top2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 565.720 0.000 566.120 0.480 ;
    END
  END Tile_X3Y15_IRQ_top2
  PIN Tile_X3Y15_IRQ_top3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 574.360 0.000 574.760 0.480 ;
    END
  END Tile_X3Y15_IRQ_top3
  PIN Tile_X5Y15_I_top0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 1108.120 0.000 1108.520 0.480 ;
    END
  END Tile_X5Y15_I_top0
  PIN Tile_X5Y15_I_top1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 1111.960 0.000 1112.360 0.480 ;
    END
  END Tile_X5Y15_I_top1
  PIN Tile_X5Y15_I_top10
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.520 0.000 1146.920 0.480 ;
    END
  END Tile_X5Y15_I_top10
  PIN Tile_X5Y15_I_top11
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 1150.360 0.000 1150.760 0.480 ;
    END
  END Tile_X5Y15_I_top11
  PIN Tile_X5Y15_I_top12
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 1154.200 0.000 1154.600 0.480 ;
    END
  END Tile_X5Y15_I_top12
  PIN Tile_X5Y15_I_top13
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 1158.040 0.000 1158.440 0.480 ;
    END
  END Tile_X5Y15_I_top13
  PIN Tile_X5Y15_I_top14
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 1161.880 0.000 1162.280 0.480 ;
    END
  END Tile_X5Y15_I_top14
  PIN Tile_X5Y15_I_top15
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 1165.720 0.000 1166.120 0.480 ;
    END
  END Tile_X5Y15_I_top15
  PIN Tile_X5Y15_I_top2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 1115.800 0.000 1116.200 0.480 ;
    END
  END Tile_X5Y15_I_top2
  PIN Tile_X5Y15_I_top3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 1119.640 0.000 1120.040 0.480 ;
    END
  END Tile_X5Y15_I_top3
  PIN Tile_X5Y15_I_top4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 1123.480 0.000 1123.880 0.480 ;
    END
  END Tile_X5Y15_I_top4
  PIN Tile_X5Y15_I_top5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 1127.320 0.000 1127.720 0.480 ;
    END
  END Tile_X5Y15_I_top5
  PIN Tile_X5Y15_I_top6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 1131.160 0.000 1131.560 0.480 ;
    END
  END Tile_X5Y15_I_top6
  PIN Tile_X5Y15_I_top7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 1135.000 0.000 1135.400 0.480 ;
    END
  END Tile_X5Y15_I_top7
  PIN Tile_X5Y15_I_top8
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 1138.840 0.000 1139.240 0.480 ;
    END
  END Tile_X5Y15_I_top8
  PIN Tile_X5Y15_I_top9
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 1142.680 0.000 1143.080 0.480 ;
    END
  END Tile_X5Y15_I_top9
  PIN Tile_X5Y15_O_top0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1046.680 0.000 1047.080 0.480 ;
    END
  END Tile_X5Y15_O_top0
  PIN Tile_X5Y15_O_top1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1050.520 0.000 1050.920 0.480 ;
    END
  END Tile_X5Y15_O_top1
  PIN Tile_X5Y15_O_top10
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1085.080 0.000 1085.480 0.480 ;
    END
  END Tile_X5Y15_O_top10
  PIN Tile_X5Y15_O_top11
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1088.920 0.000 1089.320 0.480 ;
    END
  END Tile_X5Y15_O_top11
  PIN Tile_X5Y15_O_top12
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1092.760 0.000 1093.160 0.480 ;
    END
  END Tile_X5Y15_O_top12
  PIN Tile_X5Y15_O_top13
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1096.600 0.000 1097.000 0.480 ;
    END
  END Tile_X5Y15_O_top13
  PIN Tile_X5Y15_O_top14
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1100.440 0.000 1100.840 0.480 ;
    END
  END Tile_X5Y15_O_top14
  PIN Tile_X5Y15_O_top15
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1104.280 0.000 1104.680 0.480 ;
    END
  END Tile_X5Y15_O_top15
  PIN Tile_X5Y15_O_top2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1054.360 0.000 1054.760 0.480 ;
    END
  END Tile_X5Y15_O_top2
  PIN Tile_X5Y15_O_top3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1058.200 0.000 1058.600 0.480 ;
    END
  END Tile_X5Y15_O_top3
  PIN Tile_X5Y15_O_top4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1062.040 0.000 1062.440 0.480 ;
    END
  END Tile_X5Y15_O_top4
  PIN Tile_X5Y15_O_top5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1065.880 0.000 1066.280 0.480 ;
    END
  END Tile_X5Y15_O_top5
  PIN Tile_X5Y15_O_top6
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1069.720 0.000 1070.120 0.480 ;
    END
  END Tile_X5Y15_O_top6
  PIN Tile_X5Y15_O_top7
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1073.560 0.000 1073.960 0.480 ;
    END
  END Tile_X5Y15_O_top7
  PIN Tile_X5Y15_O_top8
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1077.400 0.000 1077.800 0.480 ;
    END
  END Tile_X5Y15_O_top8
  PIN Tile_X5Y15_O_top9
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1081.240 0.000 1081.640 0.480 ;
    END
  END Tile_X5Y15_O_top9
  PIN Tile_X6Y15_I_top0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 1339.960 0.000 1340.360 0.480 ;
    END
  END Tile_X6Y15_I_top0
  PIN Tile_X6Y15_I_top1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 1343.800 0.000 1344.200 0.480 ;
    END
  END Tile_X6Y15_I_top1
  PIN Tile_X6Y15_I_top10
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 1378.360 0.000 1378.760 0.480 ;
    END
  END Tile_X6Y15_I_top10
  PIN Tile_X6Y15_I_top11
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 1382.200 0.000 1382.600 0.480 ;
    END
  END Tile_X6Y15_I_top11
  PIN Tile_X6Y15_I_top12
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 1386.040 0.000 1386.440 0.480 ;
    END
  END Tile_X6Y15_I_top12
  PIN Tile_X6Y15_I_top13
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 1389.880 0.000 1390.280 0.480 ;
    END
  END Tile_X6Y15_I_top13
  PIN Tile_X6Y15_I_top14
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 1393.720 0.000 1394.120 0.480 ;
    END
  END Tile_X6Y15_I_top14
  PIN Tile_X6Y15_I_top15
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 1397.560 0.000 1397.960 0.480 ;
    END
  END Tile_X6Y15_I_top15
  PIN Tile_X6Y15_I_top2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 1347.640 0.000 1348.040 0.480 ;
    END
  END Tile_X6Y15_I_top2
  PIN Tile_X6Y15_I_top3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 1351.480 0.000 1351.880 0.480 ;
    END
  END Tile_X6Y15_I_top3
  PIN Tile_X6Y15_I_top4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 1355.320 0.000 1355.720 0.480 ;
    END
  END Tile_X6Y15_I_top4
  PIN Tile_X6Y15_I_top5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 1359.160 0.000 1359.560 0.480 ;
    END
  END Tile_X6Y15_I_top5
  PIN Tile_X6Y15_I_top6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 1363.000 0.000 1363.400 0.480 ;
    END
  END Tile_X6Y15_I_top6
  PIN Tile_X6Y15_I_top7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 1366.840 0.000 1367.240 0.480 ;
    END
  END Tile_X6Y15_I_top7
  PIN Tile_X6Y15_I_top8
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 1370.680 0.000 1371.080 0.480 ;
    END
  END Tile_X6Y15_I_top8
  PIN Tile_X6Y15_I_top9
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 1374.520 0.000 1374.920 0.480 ;
    END
  END Tile_X6Y15_I_top9
  PIN Tile_X6Y15_O_top0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1278.520 0.000 1278.920 0.480 ;
    END
  END Tile_X6Y15_O_top0
  PIN Tile_X6Y15_O_top1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1282.360 0.000 1282.760 0.480 ;
    END
  END Tile_X6Y15_O_top1
  PIN Tile_X6Y15_O_top10
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1316.920 0.000 1317.320 0.480 ;
    END
  END Tile_X6Y15_O_top10
  PIN Tile_X6Y15_O_top11
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1320.760 0.000 1321.160 0.480 ;
    END
  END Tile_X6Y15_O_top11
  PIN Tile_X6Y15_O_top12
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1324.600 0.000 1325.000 0.480 ;
    END
  END Tile_X6Y15_O_top12
  PIN Tile_X6Y15_O_top13
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1328.440 0.000 1328.840 0.480 ;
    END
  END Tile_X6Y15_O_top13
  PIN Tile_X6Y15_O_top14
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1332.280 0.000 1332.680 0.480 ;
    END
  END Tile_X6Y15_O_top14
  PIN Tile_X6Y15_O_top15
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1336.120 0.000 1336.520 0.480 ;
    END
  END Tile_X6Y15_O_top15
  PIN Tile_X6Y15_O_top2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1286.200 0.000 1286.600 0.480 ;
    END
  END Tile_X6Y15_O_top2
  PIN Tile_X6Y15_O_top3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1290.040 0.000 1290.440 0.480 ;
    END
  END Tile_X6Y15_O_top3
  PIN Tile_X6Y15_O_top4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1293.880 0.000 1294.280 0.480 ;
    END
  END Tile_X6Y15_O_top4
  PIN Tile_X6Y15_O_top5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1297.720 0.000 1298.120 0.480 ;
    END
  END Tile_X6Y15_O_top5
  PIN Tile_X6Y15_O_top6
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1301.560 0.000 1301.960 0.480 ;
    END
  END Tile_X6Y15_O_top6
  PIN Tile_X6Y15_O_top7
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1305.400 0.000 1305.800 0.480 ;
    END
  END Tile_X6Y15_O_top7
  PIN Tile_X6Y15_O_top8
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1309.240 0.000 1309.640 0.480 ;
    END
  END Tile_X6Y15_O_top8
  PIN Tile_X6Y15_O_top9
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1313.080 0.000 1313.480 0.480 ;
    END
  END Tile_X6Y15_O_top9
  PIN Tile_X8Y15_I_top0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 1768.120 0.000 1768.520 0.480 ;
    END
  END Tile_X8Y15_I_top0
  PIN Tile_X8Y15_I_top1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 1771.960 0.000 1772.360 0.480 ;
    END
  END Tile_X8Y15_I_top1
  PIN Tile_X8Y15_I_top10
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 1806.520 0.000 1806.920 0.480 ;
    END
  END Tile_X8Y15_I_top10
  PIN Tile_X8Y15_I_top11
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 1810.360 0.000 1810.760 0.480 ;
    END
  END Tile_X8Y15_I_top11
  PIN Tile_X8Y15_I_top12
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 1814.200 0.000 1814.600 0.480 ;
    END
  END Tile_X8Y15_I_top12
  PIN Tile_X8Y15_I_top13
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 1818.040 0.000 1818.440 0.480 ;
    END
  END Tile_X8Y15_I_top13
  PIN Tile_X8Y15_I_top14
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 1821.880 0.000 1822.280 0.480 ;
    END
  END Tile_X8Y15_I_top14
  PIN Tile_X8Y15_I_top15
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 1825.720 0.000 1826.120 0.480 ;
    END
  END Tile_X8Y15_I_top15
  PIN Tile_X8Y15_I_top2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 1775.800 0.000 1776.200 0.480 ;
    END
  END Tile_X8Y15_I_top2
  PIN Tile_X8Y15_I_top3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 1779.640 0.000 1780.040 0.480 ;
    END
  END Tile_X8Y15_I_top3
  PIN Tile_X8Y15_I_top4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 1783.480 0.000 1783.880 0.480 ;
    END
  END Tile_X8Y15_I_top4
  PIN Tile_X8Y15_I_top5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 1787.320 0.000 1787.720 0.480 ;
    END
  END Tile_X8Y15_I_top5
  PIN Tile_X8Y15_I_top6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 1791.160 0.000 1791.560 0.480 ;
    END
  END Tile_X8Y15_I_top6
  PIN Tile_X8Y15_I_top7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 1795.000 0.000 1795.400 0.480 ;
    END
  END Tile_X8Y15_I_top7
  PIN Tile_X8Y15_I_top8
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 1798.840 0.000 1799.240 0.480 ;
    END
  END Tile_X8Y15_I_top8
  PIN Tile_X8Y15_I_top9
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 1802.680 0.000 1803.080 0.480 ;
    END
  END Tile_X8Y15_I_top9
  PIN Tile_X8Y15_O_top0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1706.680 0.000 1707.080 0.480 ;
    END
  END Tile_X8Y15_O_top0
  PIN Tile_X8Y15_O_top1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1710.520 0.000 1710.920 0.480 ;
    END
  END Tile_X8Y15_O_top1
  PIN Tile_X8Y15_O_top10
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1745.080 0.000 1745.480 0.480 ;
    END
  END Tile_X8Y15_O_top10
  PIN Tile_X8Y15_O_top11
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1748.920 0.000 1749.320 0.480 ;
    END
  END Tile_X8Y15_O_top11
  PIN Tile_X8Y15_O_top12
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1752.760 0.000 1753.160 0.480 ;
    END
  END Tile_X8Y15_O_top12
  PIN Tile_X8Y15_O_top13
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1756.600 0.000 1757.000 0.480 ;
    END
  END Tile_X8Y15_O_top13
  PIN Tile_X8Y15_O_top14
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1760.440 0.000 1760.840 0.480 ;
    END
  END Tile_X8Y15_O_top14
  PIN Tile_X8Y15_O_top15
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1764.280 0.000 1764.680 0.480 ;
    END
  END Tile_X8Y15_O_top15
  PIN Tile_X8Y15_O_top2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1714.360 0.000 1714.760 0.480 ;
    END
  END Tile_X8Y15_O_top2
  PIN Tile_X8Y15_O_top3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1718.200 0.000 1718.600 0.480 ;
    END
  END Tile_X8Y15_O_top3
  PIN Tile_X8Y15_O_top4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1722.040 0.000 1722.440 0.480 ;
    END
  END Tile_X8Y15_O_top4
  PIN Tile_X8Y15_O_top5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1725.880 0.000 1726.280 0.480 ;
    END
  END Tile_X8Y15_O_top5
  PIN Tile_X8Y15_O_top6
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1729.720 0.000 1730.120 0.480 ;
    END
  END Tile_X8Y15_O_top6
  PIN Tile_X8Y15_O_top7
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1733.560 0.000 1733.960 0.480 ;
    END
  END Tile_X8Y15_O_top7
  PIN Tile_X8Y15_O_top8
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1737.400 0.000 1737.800 0.480 ;
    END
  END Tile_X8Y15_O_top8
  PIN Tile_X8Y15_O_top9
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1741.240 0.000 1741.640 0.480 ;
    END
  END Tile_X8Y15_O_top9
  PIN Tile_X9Y15_I_top0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 1999.960 0.000 2000.360 0.480 ;
    END
  END Tile_X9Y15_I_top0
  PIN Tile_X9Y15_I_top1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 2003.800 0.000 2004.200 0.480 ;
    END
  END Tile_X9Y15_I_top1
  PIN Tile_X9Y15_I_top10
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 2038.360 0.000 2038.760 0.480 ;
    END
  END Tile_X9Y15_I_top10
  PIN Tile_X9Y15_I_top11
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 2042.200 0.000 2042.600 0.480 ;
    END
  END Tile_X9Y15_I_top11
  PIN Tile_X9Y15_I_top12
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 2046.040 0.000 2046.440 0.480 ;
    END
  END Tile_X9Y15_I_top12
  PIN Tile_X9Y15_I_top13
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 2049.880 0.000 2050.280 0.480 ;
    END
  END Tile_X9Y15_I_top13
  PIN Tile_X9Y15_I_top14
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 2053.720 0.000 2054.120 0.480 ;
    END
  END Tile_X9Y15_I_top14
  PIN Tile_X9Y15_I_top15
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 2057.560 0.000 2057.960 0.480 ;
    END
  END Tile_X9Y15_I_top15
  PIN Tile_X9Y15_I_top2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 2007.640 0.000 2008.040 0.480 ;
    END
  END Tile_X9Y15_I_top2
  PIN Tile_X9Y15_I_top3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 2011.480 0.000 2011.880 0.480 ;
    END
  END Tile_X9Y15_I_top3
  PIN Tile_X9Y15_I_top4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 2015.320 0.000 2015.720 0.480 ;
    END
  END Tile_X9Y15_I_top4
  PIN Tile_X9Y15_I_top5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 2019.160 0.000 2019.560 0.480 ;
    END
  END Tile_X9Y15_I_top5
  PIN Tile_X9Y15_I_top6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 2023.000 0.000 2023.400 0.480 ;
    END
  END Tile_X9Y15_I_top6
  PIN Tile_X9Y15_I_top7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 2026.840 0.000 2027.240 0.480 ;
    END
  END Tile_X9Y15_I_top7
  PIN Tile_X9Y15_I_top8
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 2030.680 0.000 2031.080 0.480 ;
    END
  END Tile_X9Y15_I_top8
  PIN Tile_X9Y15_I_top9
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 2034.520 0.000 2034.920 0.480 ;
    END
  END Tile_X9Y15_I_top9
  PIN Tile_X9Y15_O_top0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1938.520 0.000 1938.920 0.480 ;
    END
  END Tile_X9Y15_O_top0
  PIN Tile_X9Y15_O_top1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1942.360 0.000 1942.760 0.480 ;
    END
  END Tile_X9Y15_O_top1
  PIN Tile_X9Y15_O_top10
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1976.920 0.000 1977.320 0.480 ;
    END
  END Tile_X9Y15_O_top10
  PIN Tile_X9Y15_O_top11
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1980.760 0.000 1981.160 0.480 ;
    END
  END Tile_X9Y15_O_top11
  PIN Tile_X9Y15_O_top12
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1984.600 0.000 1985.000 0.480 ;
    END
  END Tile_X9Y15_O_top12
  PIN Tile_X9Y15_O_top13
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1988.440 0.000 1988.840 0.480 ;
    END
  END Tile_X9Y15_O_top13
  PIN Tile_X9Y15_O_top14
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1992.280 0.000 1992.680 0.480 ;
    END
  END Tile_X9Y15_O_top14
  PIN Tile_X9Y15_O_top15
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1996.120 0.000 1996.520 0.480 ;
    END
  END Tile_X9Y15_O_top15
  PIN Tile_X9Y15_O_top2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1946.200 0.000 1946.600 0.480 ;
    END
  END Tile_X9Y15_O_top2
  PIN Tile_X9Y15_O_top3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1950.040 0.000 1950.440 0.480 ;
    END
  END Tile_X9Y15_O_top3
  PIN Tile_X9Y15_O_top4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1953.880 0.000 1954.280 0.480 ;
    END
  END Tile_X9Y15_O_top4
  PIN Tile_X9Y15_O_top5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1957.720 0.000 1958.120 0.480 ;
    END
  END Tile_X9Y15_O_top5
  PIN Tile_X9Y15_O_top6
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1961.560 0.000 1961.960 0.480 ;
    END
  END Tile_X9Y15_O_top6
  PIN Tile_X9Y15_O_top7
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1965.400 0.000 1965.800 0.480 ;
    END
  END Tile_X9Y15_O_top7
  PIN Tile_X9Y15_O_top8
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1969.240 0.000 1969.640 0.480 ;
    END
  END Tile_X9Y15_O_top8
  PIN Tile_X9Y15_O_top9
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 1973.080 0.000 1973.480 0.480 ;
    END
  END Tile_X9Y15_O_top9
  PIN UserCLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.440100 ;
    PORT
      LAYER Metal3 ;
        RECT 5.560 0.000 5.960 0.400 ;
    END
  END UserCLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal5 ;
        RECT 24.940 4.200 27.140 3511.200 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 93.580 4.200 95.780 3511.200 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 169.180 4.200 171.380 3511.200 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 244.780 4.200 246.980 3511.200 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 325.420 4.200 327.620 3511.200 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 401.020 4.200 403.220 3511.200 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 476.620 4.200 478.820 3511.200 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 557.260 4.200 559.460 3511.200 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 632.860 4.200 635.060 3511.200 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 708.460 4.200 710.660 3511.200 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 789.100 4.200 791.300 3511.200 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 864.700 4.200 866.900 3511.200 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 940.300 4.200 942.500 3511.200 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1015.900 4.200 1018.100 3511.200 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1055.500 4.200 1057.700 3511.200 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1131.100 4.200 1133.300 3511.200 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1206.700 4.200 1208.900 3511.200 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1287.340 4.200 1289.540 3511.200 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1362.940 4.200 1365.140 3511.200 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1438.540 4.200 1440.740 3511.200 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1519.180 4.200 1521.380 3511.200 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1594.780 4.200 1596.980 3511.200 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1670.380 4.200 1672.580 3511.200 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1715.500 4.200 1717.700 3511.200 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1791.100 4.200 1793.300 3511.200 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1866.700 4.200 1868.900 3511.200 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1947.340 4.200 1949.540 3511.200 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2022.940 4.200 2025.140 3511.200 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2098.540 4.200 2100.740 3511.200 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2179.180 4.200 2181.380 3511.200 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal5 ;
        RECT 18.740 4.200 20.940 3511.200 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 87.380 4.200 89.580 3511.200 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 162.980 4.200 165.180 3511.200 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 238.580 4.200 240.780 3511.200 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 319.220 4.200 321.420 3511.200 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 394.820 4.200 397.020 3511.200 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 470.420 4.200 472.620 3511.200 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 551.060 4.200 553.260 3511.200 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 626.660 4.200 628.860 3511.200 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 702.260 4.200 704.460 3511.200 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 782.900 4.200 785.100 3511.200 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 858.500 4.200 860.700 3511.200 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 934.100 4.200 936.300 3511.200 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1009.700 4.200 1011.900 3511.200 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1049.300 4.200 1051.500 3511.200 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1124.900 4.200 1127.100 3511.200 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1200.500 4.200 1202.700 3511.200 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1281.140 4.200 1283.340 3511.200 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1356.740 4.200 1358.940 3511.200 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1432.340 4.200 1434.540 3511.200 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1512.980 4.200 1515.180 3511.200 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1588.580 4.200 1590.780 3511.200 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1664.180 4.200 1666.380 3511.200 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1709.300 4.200 1711.500 3511.200 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1784.900 4.200 1787.100 3511.200 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1860.500 4.200 1862.700 3511.200 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1941.140 4.200 1943.340 3511.200 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2016.740 4.200 2018.940 3511.200 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2092.340 4.200 2094.540 3511.200 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2172.980 4.200 2175.180 3511.200 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2248.580 4.200 2250.780 3511.200 ;
    END
  END VPWR
  OBS
      LAYER GatPoly ;
        RECT 6.240 11.610 2256.960 3503.370 ;
      LAYER Metal1 ;
        RECT 6.240 11.540 2256.980 3503.440 ;
      LAYER Metal2 ;
        RECT 0.140 3506.570 2262.720 3508.780 ;
        RECT 0.690 3505.750 2262.720 3506.570 ;
        RECT 0.140 3504.890 2262.720 3505.750 ;
        RECT 0.690 3504.070 2262.720 3504.890 ;
        RECT 0.140 3503.210 2262.720 3504.070 ;
        RECT 0.690 3502.390 2262.720 3503.210 ;
        RECT 0.140 3501.530 2262.720 3502.390 ;
        RECT 0.690 3500.710 2262.720 3501.530 ;
        RECT 0.140 3499.850 2262.720 3500.710 ;
        RECT 0.690 3499.030 2262.720 3499.850 ;
        RECT 0.140 3498.170 2262.720 3499.030 ;
        RECT 0.690 3497.350 2262.720 3498.170 ;
        RECT 0.140 3496.490 2262.720 3497.350 ;
        RECT 0.690 3495.670 2262.720 3496.490 ;
        RECT 0.140 3494.810 2262.720 3495.670 ;
        RECT 0.690 3493.990 2262.720 3494.810 ;
        RECT 0.140 3493.130 2262.720 3493.990 ;
        RECT 0.690 3492.310 2262.720 3493.130 ;
        RECT 0.140 3491.450 2262.720 3492.310 ;
        RECT 0.690 3490.630 2262.720 3491.450 ;
        RECT 0.140 3489.770 2262.720 3490.630 ;
        RECT 0.690 3488.950 2262.720 3489.770 ;
        RECT 0.140 3488.090 2262.720 3488.950 ;
        RECT 0.690 3487.270 2262.720 3488.090 ;
        RECT 0.140 3486.410 2262.720 3487.270 ;
        RECT 0.690 3485.590 2262.720 3486.410 ;
        RECT 0.140 3484.730 2262.720 3485.590 ;
        RECT 0.690 3483.910 2262.720 3484.730 ;
        RECT 0.140 3483.050 2262.720 3483.910 ;
        RECT 0.690 3482.230 2262.720 3483.050 ;
        RECT 0.140 3481.370 2262.720 3482.230 ;
        RECT 0.690 3480.550 2262.720 3481.370 ;
        RECT 0.140 3479.690 2262.720 3480.550 ;
        RECT 0.690 3478.870 2262.720 3479.690 ;
        RECT 0.140 3478.010 2262.720 3478.870 ;
        RECT 0.690 3477.190 2262.720 3478.010 ;
        RECT 0.140 3476.330 2262.720 3477.190 ;
        RECT 0.690 3475.510 2262.720 3476.330 ;
        RECT 0.140 3474.650 2262.720 3475.510 ;
        RECT 0.690 3473.830 2262.720 3474.650 ;
        RECT 0.140 3472.970 2262.720 3473.830 ;
        RECT 0.690 3472.150 2262.720 3472.970 ;
        RECT 0.140 3471.290 2262.720 3472.150 ;
        RECT 0.690 3470.470 2262.720 3471.290 ;
        RECT 0.140 3469.610 2262.720 3470.470 ;
        RECT 0.690 3468.790 2262.720 3469.610 ;
        RECT 0.140 3467.930 2262.720 3468.790 ;
        RECT 0.690 3467.110 2262.720 3467.930 ;
        RECT 0.140 3466.250 2262.720 3467.110 ;
        RECT 0.690 3465.430 2262.720 3466.250 ;
        RECT 0.140 3464.570 2262.720 3465.430 ;
        RECT 0.690 3463.750 2262.720 3464.570 ;
        RECT 0.140 3462.890 2262.720 3463.750 ;
        RECT 0.690 3462.070 2262.720 3462.890 ;
        RECT 0.140 3461.210 2262.720 3462.070 ;
        RECT 0.690 3460.390 2262.720 3461.210 ;
        RECT 0.140 3459.530 2262.720 3460.390 ;
        RECT 0.690 3458.710 2262.720 3459.530 ;
        RECT 0.140 3457.850 2262.720 3458.710 ;
        RECT 0.690 3457.030 2262.720 3457.850 ;
        RECT 0.140 3456.170 2262.720 3457.030 ;
        RECT 0.690 3455.350 2262.720 3456.170 ;
        RECT 0.140 3454.490 2262.720 3455.350 ;
        RECT 0.690 3453.670 2262.720 3454.490 ;
        RECT 0.140 3442.730 2262.720 3453.670 ;
        RECT 1.140 3441.910 2262.720 3442.730 ;
        RECT 0.140 3437.690 2262.720 3441.910 ;
        RECT 1.140 3436.870 2262.720 3437.690 ;
        RECT 0.140 3432.650 2262.720 3436.870 ;
        RECT 1.070 3431.830 2262.720 3432.650 ;
        RECT 0.140 3427.610 2262.720 3431.830 ;
        RECT 1.070 3426.790 2262.720 3427.610 ;
        RECT 0.140 3422.570 2262.720 3426.790 ;
        RECT 1.140 3421.750 2262.720 3422.570 ;
        RECT 0.140 3417.530 2262.720 3421.750 ;
        RECT 1.070 3416.710 2262.720 3417.530 ;
        RECT 0.140 3412.490 2262.720 3416.710 ;
        RECT 1.070 3411.670 2262.720 3412.490 ;
        RECT 0.140 3407.450 2262.720 3411.670 ;
        RECT 1.140 3406.630 2262.720 3407.450 ;
        RECT 0.140 3402.410 2262.720 3406.630 ;
        RECT 1.070 3401.590 2262.720 3402.410 ;
        RECT 0.140 3397.370 2262.720 3401.590 ;
        RECT 1.070 3396.550 2262.720 3397.370 ;
        RECT 0.140 3392.330 2262.720 3396.550 ;
        RECT 1.140 3391.510 2262.720 3392.330 ;
        RECT 0.140 3387.290 2262.720 3391.510 ;
        RECT 1.070 3386.470 2262.720 3387.290 ;
        RECT 0.140 3382.250 2262.720 3386.470 ;
        RECT 1.070 3381.430 2262.720 3382.250 ;
        RECT 0.140 3377.210 2262.720 3381.430 ;
        RECT 1.140 3376.390 2262.720 3377.210 ;
        RECT 0.140 3372.170 2262.720 3376.390 ;
        RECT 1.070 3371.350 2262.720 3372.170 ;
        RECT 0.140 3367.130 2262.720 3371.350 ;
        RECT 1.070 3366.310 2262.720 3367.130 ;
        RECT 0.140 3362.090 2262.720 3366.310 ;
        RECT 1.140 3361.270 2262.720 3362.090 ;
        RECT 0.140 3357.050 2262.720 3361.270 ;
        RECT 1.070 3356.230 2262.720 3357.050 ;
        RECT 0.140 3352.010 2262.720 3356.230 ;
        RECT 1.070 3351.190 2262.720 3352.010 ;
        RECT 0.140 3346.970 2262.720 3351.190 ;
        RECT 1.140 3346.150 2262.720 3346.970 ;
        RECT 0.140 3341.930 2262.720 3346.150 ;
        RECT 1.140 3341.110 2262.720 3341.930 ;
        RECT 0.140 3336.890 2262.720 3341.110 ;
        RECT 1.140 3336.070 2262.720 3336.890 ;
        RECT 0.140 3331.850 2262.720 3336.070 ;
        RECT 1.140 3331.030 2262.720 3331.850 ;
        RECT 0.140 3326.810 2262.720 3331.030 ;
        RECT 1.140 3325.990 2262.720 3326.810 ;
        RECT 0.140 3321.770 2262.720 3325.990 ;
        RECT 1.070 3320.950 2262.720 3321.770 ;
        RECT 0.140 3316.730 2262.720 3320.950 ;
        RECT 1.140 3315.910 2262.720 3316.730 ;
        RECT 0.140 3311.690 2262.720 3315.910 ;
        RECT 1.070 3310.870 2262.720 3311.690 ;
        RECT 0.140 3306.650 2262.720 3310.870 ;
        RECT 1.070 3305.830 2262.720 3306.650 ;
        RECT 0.140 3301.610 2262.720 3305.830 ;
        RECT 1.070 3300.790 2262.720 3301.610 ;
        RECT 0.140 3296.570 2262.720 3300.790 ;
        RECT 1.070 3295.750 2262.720 3296.570 ;
        RECT 0.140 3291.530 2262.720 3295.750 ;
        RECT 1.070 3290.710 2262.720 3291.530 ;
        RECT 0.140 3286.490 2262.720 3290.710 ;
        RECT 1.140 3285.670 2262.720 3286.490 ;
        RECT 0.140 3281.450 2262.720 3285.670 ;
        RECT 1.140 3280.630 2262.720 3281.450 ;
        RECT 0.140 3276.410 2262.720 3280.630 ;
        RECT 1.070 3275.590 2262.720 3276.410 ;
        RECT 0.140 3271.370 2262.720 3275.590 ;
        RECT 1.140 3270.550 2262.720 3271.370 ;
        RECT 0.140 3268.850 2262.720 3270.550 ;
        RECT 0.140 3268.030 2262.060 3268.850 ;
        RECT 0.140 3266.330 2262.720 3268.030 ;
        RECT 1.140 3265.510 2262.060 3266.330 ;
        RECT 0.140 3263.810 2262.720 3265.510 ;
        RECT 0.140 3262.990 2262.060 3263.810 ;
        RECT 0.140 3261.290 2262.720 3262.990 ;
        RECT 1.140 3260.470 2262.060 3261.290 ;
        RECT 0.140 3258.770 2262.720 3260.470 ;
        RECT 0.140 3257.950 2262.060 3258.770 ;
        RECT 0.140 3256.250 2262.720 3257.950 ;
        RECT 1.070 3255.430 2262.060 3256.250 ;
        RECT 0.140 3253.730 2262.720 3255.430 ;
        RECT 0.140 3252.910 2262.060 3253.730 ;
        RECT 0.140 3251.210 2262.720 3252.910 ;
        RECT 1.140 3250.390 2262.060 3251.210 ;
        RECT 0.140 3248.690 2262.720 3250.390 ;
        RECT 0.140 3247.870 2262.060 3248.690 ;
        RECT 0.140 3246.170 2262.720 3247.870 ;
        RECT 1.140 3245.350 2262.060 3246.170 ;
        RECT 0.140 3243.650 2262.720 3245.350 ;
        RECT 0.140 3242.830 2262.060 3243.650 ;
        RECT 0.140 3241.130 2262.720 3242.830 ;
        RECT 1.140 3240.310 2262.060 3241.130 ;
        RECT 0.140 3238.610 2262.720 3240.310 ;
        RECT 0.140 3237.790 2262.060 3238.610 ;
        RECT 0.140 3236.090 2262.720 3237.790 ;
        RECT 1.140 3235.270 2262.060 3236.090 ;
        RECT 0.140 3233.570 2262.720 3235.270 ;
        RECT 0.140 3232.750 2262.060 3233.570 ;
        RECT 0.140 3231.050 2262.720 3232.750 ;
        RECT 1.140 3230.230 2262.060 3231.050 ;
        RECT 0.140 3228.530 2262.720 3230.230 ;
        RECT 0.140 3227.710 2262.060 3228.530 ;
        RECT 0.140 3226.010 2262.720 3227.710 ;
        RECT 1.070 3225.190 2262.060 3226.010 ;
        RECT 0.140 3223.490 2262.720 3225.190 ;
        RECT 0.140 3222.670 2262.060 3223.490 ;
        RECT 0.140 3220.970 2262.720 3222.670 ;
        RECT 1.140 3220.150 2262.060 3220.970 ;
        RECT 0.140 3218.450 2262.720 3220.150 ;
        RECT 0.140 3217.630 2262.060 3218.450 ;
        RECT 0.140 3215.930 2262.720 3217.630 ;
        RECT 1.070 3215.110 2262.060 3215.930 ;
        RECT 0.140 3213.410 2262.720 3215.110 ;
        RECT 0.140 3212.590 2262.060 3213.410 ;
        RECT 0.140 3210.890 2262.720 3212.590 ;
        RECT 0.140 3210.070 2262.060 3210.890 ;
        RECT 0.140 3208.370 2262.720 3210.070 ;
        RECT 0.140 3207.550 2262.060 3208.370 ;
        RECT 0.140 3205.850 2262.720 3207.550 ;
        RECT 0.140 3205.030 2262.060 3205.850 ;
        RECT 0.140 3203.330 2262.720 3205.030 ;
        RECT 0.140 3202.510 2262.060 3203.330 ;
        RECT 0.140 3200.810 2262.720 3202.510 ;
        RECT 1.140 3199.990 2262.060 3200.810 ;
        RECT 0.140 3198.290 2262.720 3199.990 ;
        RECT 0.140 3197.470 2262.060 3198.290 ;
        RECT 0.140 3195.770 2262.720 3197.470 ;
        RECT 1.140 3194.950 2262.060 3195.770 ;
        RECT 0.140 3193.250 2262.720 3194.950 ;
        RECT 0.140 3192.430 2262.060 3193.250 ;
        RECT 0.140 3190.730 2262.720 3192.430 ;
        RECT 1.070 3189.910 2262.060 3190.730 ;
        RECT 0.140 3188.210 2262.720 3189.910 ;
        RECT 0.140 3187.390 2262.060 3188.210 ;
        RECT 0.140 3185.690 2262.720 3187.390 ;
        RECT 1.070 3184.870 2262.060 3185.690 ;
        RECT 0.140 3183.170 2262.720 3184.870 ;
        RECT 0.140 3182.350 2262.060 3183.170 ;
        RECT 0.140 3180.650 2262.720 3182.350 ;
        RECT 1.140 3179.830 2262.060 3180.650 ;
        RECT 0.140 3178.130 2262.720 3179.830 ;
        RECT 0.140 3177.310 2262.060 3178.130 ;
        RECT 0.140 3175.610 2262.720 3177.310 ;
        RECT 1.070 3174.790 2262.060 3175.610 ;
        RECT 0.140 3173.090 2262.720 3174.790 ;
        RECT 0.140 3172.270 2262.060 3173.090 ;
        RECT 0.140 3170.570 2262.720 3172.270 ;
        RECT 1.070 3169.750 2262.060 3170.570 ;
        RECT 0.140 3168.050 2262.720 3169.750 ;
        RECT 0.140 3167.230 2262.060 3168.050 ;
        RECT 0.140 3165.530 2262.720 3167.230 ;
        RECT 1.140 3164.710 2262.060 3165.530 ;
        RECT 0.140 3163.010 2262.720 3164.710 ;
        RECT 0.140 3162.190 2262.060 3163.010 ;
        RECT 0.140 3160.490 2262.720 3162.190 ;
        RECT 1.070 3159.670 2262.060 3160.490 ;
        RECT 0.140 3157.970 2262.720 3159.670 ;
        RECT 0.140 3157.150 2262.060 3157.970 ;
        RECT 0.140 3155.450 2262.720 3157.150 ;
        RECT 1.070 3154.630 2262.060 3155.450 ;
        RECT 0.140 3152.930 2262.720 3154.630 ;
        RECT 0.140 3152.110 2262.060 3152.930 ;
        RECT 0.140 3150.410 2262.720 3152.110 ;
        RECT 1.140 3149.590 2262.060 3150.410 ;
        RECT 0.140 3147.890 2262.720 3149.590 ;
        RECT 0.140 3147.070 2262.060 3147.890 ;
        RECT 0.140 3145.370 2262.720 3147.070 ;
        RECT 1.070 3144.550 2262.060 3145.370 ;
        RECT 0.140 3142.850 2262.720 3144.550 ;
        RECT 0.140 3142.030 2262.060 3142.850 ;
        RECT 0.140 3140.330 2262.720 3142.030 ;
        RECT 1.070 3139.510 2262.060 3140.330 ;
        RECT 0.140 3137.810 2262.720 3139.510 ;
        RECT 0.140 3136.990 2262.060 3137.810 ;
        RECT 0.140 3135.290 2262.720 3136.990 ;
        RECT 1.140 3134.470 2262.060 3135.290 ;
        RECT 0.140 3132.770 2262.720 3134.470 ;
        RECT 0.140 3131.950 2262.060 3132.770 ;
        RECT 0.140 3130.250 2262.720 3131.950 ;
        RECT 1.070 3129.430 2262.060 3130.250 ;
        RECT 0.140 3127.730 2262.720 3129.430 ;
        RECT 0.140 3126.910 2262.060 3127.730 ;
        RECT 0.140 3125.210 2262.720 3126.910 ;
        RECT 1.070 3124.390 2262.060 3125.210 ;
        RECT 0.140 3122.690 2262.720 3124.390 ;
        RECT 0.140 3121.870 2262.060 3122.690 ;
        RECT 0.140 3120.170 2262.720 3121.870 ;
        RECT 1.140 3119.350 2262.060 3120.170 ;
        RECT 0.140 3117.650 2262.720 3119.350 ;
        RECT 0.140 3116.830 2262.060 3117.650 ;
        RECT 0.140 3115.130 2262.720 3116.830 ;
        RECT 1.070 3114.310 2262.060 3115.130 ;
        RECT 0.140 3112.610 2262.720 3114.310 ;
        RECT 0.140 3111.790 2262.060 3112.610 ;
        RECT 0.140 3110.090 2262.720 3111.790 ;
        RECT 1.070 3109.270 2262.060 3110.090 ;
        RECT 0.140 3107.570 2262.720 3109.270 ;
        RECT 0.140 3106.750 2262.060 3107.570 ;
        RECT 0.140 3105.050 2262.720 3106.750 ;
        RECT 1.140 3104.230 2262.060 3105.050 ;
        RECT 0.140 3102.530 2262.720 3104.230 ;
        RECT 0.140 3101.710 2262.060 3102.530 ;
        RECT 0.140 3100.010 2262.720 3101.710 ;
        RECT 1.140 3099.190 2262.060 3100.010 ;
        RECT 0.140 3097.490 2262.720 3099.190 ;
        RECT 0.140 3096.670 2262.060 3097.490 ;
        RECT 0.140 3094.970 2262.720 3096.670 ;
        RECT 1.140 3094.150 2262.060 3094.970 ;
        RECT 0.140 3092.450 2262.720 3094.150 ;
        RECT 0.140 3091.630 2262.060 3092.450 ;
        RECT 0.140 3089.930 2262.720 3091.630 ;
        RECT 1.140 3089.110 2262.060 3089.930 ;
        RECT 0.140 3087.410 2262.720 3089.110 ;
        RECT 0.140 3086.590 2262.060 3087.410 ;
        RECT 0.140 3084.890 2262.720 3086.590 ;
        RECT 1.140 3084.070 2262.060 3084.890 ;
        RECT 0.140 3082.370 2262.720 3084.070 ;
        RECT 0.140 3081.550 2262.060 3082.370 ;
        RECT 0.140 3079.850 2262.720 3081.550 ;
        RECT 1.070 3079.030 2262.060 3079.850 ;
        RECT 0.140 3077.330 2262.720 3079.030 ;
        RECT 0.140 3076.510 2262.060 3077.330 ;
        RECT 0.140 3074.810 2262.720 3076.510 ;
        RECT 1.140 3073.990 2262.060 3074.810 ;
        RECT 0.140 3072.290 2262.720 3073.990 ;
        RECT 0.140 3071.470 2262.130 3072.290 ;
        RECT 0.140 3069.770 2262.720 3071.470 ;
        RECT 1.070 3068.950 2262.060 3069.770 ;
        RECT 0.140 3067.250 2262.720 3068.950 ;
        RECT 0.140 3066.430 2262.060 3067.250 ;
        RECT 0.140 3064.730 2262.720 3066.430 ;
        RECT 1.070 3063.910 2262.060 3064.730 ;
        RECT 0.140 3062.210 2262.720 3063.910 ;
        RECT 0.140 3061.390 2262.060 3062.210 ;
        RECT 0.140 3059.690 2262.720 3061.390 ;
        RECT 1.070 3058.870 2262.060 3059.690 ;
        RECT 0.140 3057.170 2262.720 3058.870 ;
        RECT 0.140 3056.350 2262.060 3057.170 ;
        RECT 0.140 3054.650 2262.720 3056.350 ;
        RECT 1.070 3053.830 2262.060 3054.650 ;
        RECT 0.140 3052.130 2262.720 3053.830 ;
        RECT 0.140 3051.310 2262.060 3052.130 ;
        RECT 0.140 3049.610 2262.720 3051.310 ;
        RECT 1.070 3048.790 2262.060 3049.610 ;
        RECT 0.140 3047.090 2262.720 3048.790 ;
        RECT 0.140 3046.270 2262.060 3047.090 ;
        RECT 0.140 3044.570 2262.720 3046.270 ;
        RECT 1.140 3043.750 2262.060 3044.570 ;
        RECT 0.140 3042.050 2262.720 3043.750 ;
        RECT 0.140 3041.230 2262.060 3042.050 ;
        RECT 0.140 3039.530 2262.720 3041.230 ;
        RECT 1.140 3038.710 2262.060 3039.530 ;
        RECT 0.140 3037.010 2262.720 3038.710 ;
        RECT 0.140 3036.190 2262.060 3037.010 ;
        RECT 0.140 3034.490 2262.720 3036.190 ;
        RECT 1.070 3033.670 2262.060 3034.490 ;
        RECT 0.140 3031.970 2262.720 3033.670 ;
        RECT 0.140 3031.150 2262.060 3031.970 ;
        RECT 0.140 3029.450 2262.720 3031.150 ;
        RECT 1.140 3028.630 2262.060 3029.450 ;
        RECT 0.140 3026.930 2262.720 3028.630 ;
        RECT 0.140 3026.110 2262.060 3026.930 ;
        RECT 0.140 3024.410 2262.720 3026.110 ;
        RECT 1.140 3023.590 2262.060 3024.410 ;
        RECT 0.140 3021.890 2262.720 3023.590 ;
        RECT 0.140 3021.070 2262.060 3021.890 ;
        RECT 0.140 3019.370 2262.720 3021.070 ;
        RECT 1.140 3018.550 2262.060 3019.370 ;
        RECT 0.140 3016.850 2262.720 3018.550 ;
        RECT 0.140 3016.030 2262.060 3016.850 ;
        RECT 0.140 3014.330 2262.720 3016.030 ;
        RECT 1.070 3013.510 2262.060 3014.330 ;
        RECT 0.140 3011.810 2262.720 3013.510 ;
        RECT 0.140 3010.990 2262.060 3011.810 ;
        RECT 0.140 3009.290 2262.720 3010.990 ;
        RECT 1.140 3008.470 2262.060 3009.290 ;
        RECT 0.140 3006.770 2262.720 3008.470 ;
        RECT 0.140 3005.950 2262.060 3006.770 ;
        RECT 0.140 3004.250 2262.720 3005.950 ;
        RECT 1.140 3003.430 2262.060 3004.250 ;
        RECT 0.140 3001.730 2262.720 3003.430 ;
        RECT 0.140 3000.910 2262.060 3001.730 ;
        RECT 0.140 2999.210 2262.720 3000.910 ;
        RECT 1.140 2998.390 2262.060 2999.210 ;
        RECT 0.140 2996.690 2262.720 2998.390 ;
        RECT 0.140 2995.870 2262.060 2996.690 ;
        RECT 0.140 2994.170 2262.720 2995.870 ;
        RECT 1.140 2993.350 2262.060 2994.170 ;
        RECT 0.140 2991.650 2262.720 2993.350 ;
        RECT 0.140 2990.830 2262.060 2991.650 ;
        RECT 0.140 2989.130 2262.720 2990.830 ;
        RECT 1.140 2988.310 2262.060 2989.130 ;
        RECT 0.140 2986.610 2262.720 2988.310 ;
        RECT 0.140 2985.790 2262.060 2986.610 ;
        RECT 0.140 2984.090 2262.720 2985.790 ;
        RECT 1.070 2983.270 2262.720 2984.090 ;
        RECT 0.140 2979.050 2262.720 2983.270 ;
        RECT 1.140 2978.230 2262.720 2979.050 ;
        RECT 0.140 2974.010 2262.720 2978.230 ;
        RECT 1.070 2973.190 2262.720 2974.010 ;
        RECT 0.140 2958.890 2262.720 2973.190 ;
        RECT 1.140 2958.070 2262.720 2958.890 ;
        RECT 0.140 2953.850 2262.720 2958.070 ;
        RECT 1.140 2953.030 2262.720 2953.850 ;
        RECT 0.140 2948.810 2262.720 2953.030 ;
        RECT 1.070 2947.990 2262.720 2948.810 ;
        RECT 0.140 2943.770 2262.720 2947.990 ;
        RECT 1.070 2942.950 2262.720 2943.770 ;
        RECT 0.140 2938.730 2262.720 2942.950 ;
        RECT 1.140 2937.910 2262.720 2938.730 ;
        RECT 0.140 2933.690 2262.720 2937.910 ;
        RECT 1.070 2932.870 2262.720 2933.690 ;
        RECT 0.140 2928.650 2262.720 2932.870 ;
        RECT 1.070 2927.830 2262.720 2928.650 ;
        RECT 0.140 2923.610 2262.720 2927.830 ;
        RECT 1.140 2922.790 2262.720 2923.610 ;
        RECT 0.140 2918.570 2262.720 2922.790 ;
        RECT 1.070 2917.750 2262.720 2918.570 ;
        RECT 0.140 2913.530 2262.720 2917.750 ;
        RECT 1.070 2912.710 2262.720 2913.530 ;
        RECT 0.140 2908.490 2262.720 2912.710 ;
        RECT 1.140 2907.670 2262.720 2908.490 ;
        RECT 0.140 2903.450 2262.720 2907.670 ;
        RECT 1.070 2902.630 2262.720 2903.450 ;
        RECT 0.140 2898.410 2262.720 2902.630 ;
        RECT 1.070 2897.590 2262.720 2898.410 ;
        RECT 0.140 2893.370 2262.720 2897.590 ;
        RECT 1.140 2892.550 2262.720 2893.370 ;
        RECT 0.140 2888.330 2262.720 2892.550 ;
        RECT 1.070 2887.510 2262.720 2888.330 ;
        RECT 0.140 2883.290 2262.720 2887.510 ;
        RECT 1.070 2882.470 2262.720 2883.290 ;
        RECT 0.140 2878.250 2262.720 2882.470 ;
        RECT 1.140 2877.430 2262.720 2878.250 ;
        RECT 0.140 2873.210 2262.720 2877.430 ;
        RECT 1.070 2872.390 2262.720 2873.210 ;
        RECT 0.140 2868.170 2262.720 2872.390 ;
        RECT 1.070 2867.350 2262.720 2868.170 ;
        RECT 0.140 2863.130 2262.720 2867.350 ;
        RECT 1.140 2862.310 2262.720 2863.130 ;
        RECT 0.140 2858.090 2262.720 2862.310 ;
        RECT 1.140 2857.270 2262.720 2858.090 ;
        RECT 0.140 2853.050 2262.720 2857.270 ;
        RECT 1.140 2852.230 2262.720 2853.050 ;
        RECT 0.140 2848.010 2262.720 2852.230 ;
        RECT 1.140 2847.190 2262.720 2848.010 ;
        RECT 0.140 2842.970 2262.720 2847.190 ;
        RECT 1.140 2842.150 2262.720 2842.970 ;
        RECT 0.140 2837.930 2262.720 2842.150 ;
        RECT 1.070 2837.110 2262.720 2837.930 ;
        RECT 0.140 2832.890 2262.720 2837.110 ;
        RECT 1.140 2832.070 2262.720 2832.890 ;
        RECT 0.140 2827.850 2262.720 2832.070 ;
        RECT 1.070 2827.030 2262.720 2827.850 ;
        RECT 0.140 2822.810 2262.720 2827.030 ;
        RECT 1.070 2821.990 2262.720 2822.810 ;
        RECT 0.140 2817.770 2262.720 2821.990 ;
        RECT 1.070 2816.950 2262.720 2817.770 ;
        RECT 0.140 2812.730 2262.720 2816.950 ;
        RECT 1.070 2811.910 2262.720 2812.730 ;
        RECT 0.140 2807.690 2262.720 2811.910 ;
        RECT 1.070 2806.870 2262.720 2807.690 ;
        RECT 0.140 2802.650 2262.720 2806.870 ;
        RECT 1.140 2801.830 2262.720 2802.650 ;
        RECT 0.140 2797.610 2262.720 2801.830 ;
        RECT 1.140 2796.790 2262.720 2797.610 ;
        RECT 0.140 2792.570 2262.720 2796.790 ;
        RECT 1.070 2791.750 2262.720 2792.570 ;
        RECT 0.140 2787.530 2262.720 2791.750 ;
        RECT 1.140 2786.710 2262.720 2787.530 ;
        RECT 0.140 2785.010 2262.720 2786.710 ;
        RECT 0.140 2784.190 2262.060 2785.010 ;
        RECT 0.140 2782.490 2262.720 2784.190 ;
        RECT 1.140 2781.670 2262.060 2782.490 ;
        RECT 0.140 2779.970 2262.720 2781.670 ;
        RECT 0.140 2779.150 2262.060 2779.970 ;
        RECT 0.140 2777.450 2262.720 2779.150 ;
        RECT 1.140 2776.630 2262.060 2777.450 ;
        RECT 0.140 2774.930 2262.720 2776.630 ;
        RECT 0.140 2774.110 2262.060 2774.930 ;
        RECT 0.140 2772.410 2262.720 2774.110 ;
        RECT 1.070 2771.590 2262.060 2772.410 ;
        RECT 0.140 2769.890 2262.720 2771.590 ;
        RECT 0.140 2769.070 2262.060 2769.890 ;
        RECT 0.140 2767.370 2262.720 2769.070 ;
        RECT 1.140 2766.550 2262.060 2767.370 ;
        RECT 0.140 2764.850 2262.720 2766.550 ;
        RECT 0.140 2764.030 2262.060 2764.850 ;
        RECT 0.140 2762.330 2262.720 2764.030 ;
        RECT 1.140 2761.510 2262.060 2762.330 ;
        RECT 0.140 2759.810 2262.720 2761.510 ;
        RECT 0.140 2758.990 2262.060 2759.810 ;
        RECT 0.140 2757.290 2262.720 2758.990 ;
        RECT 1.140 2756.470 2262.060 2757.290 ;
        RECT 0.140 2754.770 2262.720 2756.470 ;
        RECT 0.140 2753.950 2262.060 2754.770 ;
        RECT 0.140 2752.250 2262.720 2753.950 ;
        RECT 1.140 2751.430 2262.060 2752.250 ;
        RECT 0.140 2749.730 2262.720 2751.430 ;
        RECT 0.140 2748.910 2262.060 2749.730 ;
        RECT 0.140 2747.210 2262.720 2748.910 ;
        RECT 1.140 2746.390 2262.060 2747.210 ;
        RECT 0.140 2744.690 2262.720 2746.390 ;
        RECT 0.140 2743.870 2262.060 2744.690 ;
        RECT 0.140 2742.170 2262.720 2743.870 ;
        RECT 1.070 2741.350 2262.060 2742.170 ;
        RECT 0.140 2739.650 2262.720 2741.350 ;
        RECT 0.140 2738.830 2262.060 2739.650 ;
        RECT 0.140 2737.130 2262.720 2738.830 ;
        RECT 1.140 2736.310 2262.060 2737.130 ;
        RECT 0.140 2734.610 2262.720 2736.310 ;
        RECT 0.140 2733.790 2262.060 2734.610 ;
        RECT 0.140 2732.090 2262.720 2733.790 ;
        RECT 1.070 2731.270 2262.060 2732.090 ;
        RECT 0.140 2729.570 2262.720 2731.270 ;
        RECT 0.140 2728.750 2262.060 2729.570 ;
        RECT 0.140 2727.050 2262.720 2728.750 ;
        RECT 0.140 2726.230 2262.060 2727.050 ;
        RECT 0.140 2724.530 2262.720 2726.230 ;
        RECT 0.140 2723.710 2262.060 2724.530 ;
        RECT 0.140 2722.010 2262.720 2723.710 ;
        RECT 0.140 2721.190 2262.060 2722.010 ;
        RECT 0.140 2719.490 2262.720 2721.190 ;
        RECT 0.140 2718.670 2262.060 2719.490 ;
        RECT 0.140 2716.970 2262.720 2718.670 ;
        RECT 1.140 2716.150 2262.060 2716.970 ;
        RECT 0.140 2714.450 2262.720 2716.150 ;
        RECT 0.140 2713.630 2262.060 2714.450 ;
        RECT 0.140 2711.930 2262.720 2713.630 ;
        RECT 1.140 2711.110 2262.060 2711.930 ;
        RECT 0.140 2709.410 2262.720 2711.110 ;
        RECT 0.140 2708.590 2262.060 2709.410 ;
        RECT 0.140 2706.890 2262.720 2708.590 ;
        RECT 1.070 2706.070 2262.060 2706.890 ;
        RECT 0.140 2704.370 2262.720 2706.070 ;
        RECT 0.140 2703.550 2262.060 2704.370 ;
        RECT 0.140 2701.850 2262.720 2703.550 ;
        RECT 1.070 2701.030 2262.060 2701.850 ;
        RECT 0.140 2699.330 2262.720 2701.030 ;
        RECT 0.140 2698.510 2262.060 2699.330 ;
        RECT 0.140 2696.810 2262.720 2698.510 ;
        RECT 1.140 2695.990 2262.060 2696.810 ;
        RECT 0.140 2694.290 2262.720 2695.990 ;
        RECT 0.140 2693.470 2262.060 2694.290 ;
        RECT 0.140 2691.770 2262.720 2693.470 ;
        RECT 1.070 2690.950 2262.060 2691.770 ;
        RECT 0.140 2689.250 2262.720 2690.950 ;
        RECT 0.140 2688.430 2262.060 2689.250 ;
        RECT 0.140 2686.730 2262.720 2688.430 ;
        RECT 1.070 2685.910 2262.060 2686.730 ;
        RECT 0.140 2684.210 2262.720 2685.910 ;
        RECT 0.140 2683.390 2262.060 2684.210 ;
        RECT 0.140 2681.690 2262.720 2683.390 ;
        RECT 1.140 2680.870 2262.060 2681.690 ;
        RECT 0.140 2679.170 2262.720 2680.870 ;
        RECT 0.140 2678.350 2262.060 2679.170 ;
        RECT 0.140 2676.650 2262.720 2678.350 ;
        RECT 1.070 2675.830 2262.060 2676.650 ;
        RECT 0.140 2674.130 2262.720 2675.830 ;
        RECT 0.140 2673.310 2262.060 2674.130 ;
        RECT 0.140 2671.610 2262.720 2673.310 ;
        RECT 1.070 2670.790 2262.060 2671.610 ;
        RECT 0.140 2669.090 2262.720 2670.790 ;
        RECT 0.140 2668.270 2262.060 2669.090 ;
        RECT 0.140 2666.570 2262.720 2668.270 ;
        RECT 1.140 2665.750 2262.060 2666.570 ;
        RECT 0.140 2664.050 2262.720 2665.750 ;
        RECT 0.140 2663.230 2262.060 2664.050 ;
        RECT 0.140 2661.530 2262.720 2663.230 ;
        RECT 1.070 2660.710 2262.060 2661.530 ;
        RECT 0.140 2659.010 2262.720 2660.710 ;
        RECT 0.140 2658.190 2262.060 2659.010 ;
        RECT 0.140 2656.490 2262.720 2658.190 ;
        RECT 1.070 2655.670 2262.060 2656.490 ;
        RECT 0.140 2653.970 2262.720 2655.670 ;
        RECT 0.140 2653.150 2262.060 2653.970 ;
        RECT 0.140 2651.450 2262.720 2653.150 ;
        RECT 1.140 2650.630 2262.060 2651.450 ;
        RECT 0.140 2648.930 2262.720 2650.630 ;
        RECT 0.140 2648.110 2262.060 2648.930 ;
        RECT 0.140 2646.410 2262.720 2648.110 ;
        RECT 1.070 2645.590 2262.060 2646.410 ;
        RECT 0.140 2643.890 2262.720 2645.590 ;
        RECT 0.140 2643.070 2262.060 2643.890 ;
        RECT 0.140 2641.370 2262.720 2643.070 ;
        RECT 1.070 2640.550 2262.060 2641.370 ;
        RECT 0.140 2638.850 2262.720 2640.550 ;
        RECT 0.140 2638.030 2262.060 2638.850 ;
        RECT 0.140 2636.330 2262.720 2638.030 ;
        RECT 1.140 2635.510 2262.060 2636.330 ;
        RECT 0.140 2633.810 2262.720 2635.510 ;
        RECT 0.140 2632.990 2262.060 2633.810 ;
        RECT 0.140 2631.290 2262.720 2632.990 ;
        RECT 1.070 2630.470 2262.060 2631.290 ;
        RECT 0.140 2628.770 2262.720 2630.470 ;
        RECT 0.140 2627.950 2262.060 2628.770 ;
        RECT 0.140 2626.250 2262.720 2627.950 ;
        RECT 1.070 2625.430 2262.060 2626.250 ;
        RECT 0.140 2623.730 2262.720 2625.430 ;
        RECT 0.140 2622.910 2262.060 2623.730 ;
        RECT 0.140 2621.210 2262.720 2622.910 ;
        RECT 1.140 2620.390 2262.060 2621.210 ;
        RECT 0.140 2618.690 2262.720 2620.390 ;
        RECT 0.140 2617.870 2262.060 2618.690 ;
        RECT 0.140 2616.170 2262.720 2617.870 ;
        RECT 1.140 2615.350 2262.060 2616.170 ;
        RECT 0.140 2613.650 2262.720 2615.350 ;
        RECT 0.140 2612.830 2262.060 2613.650 ;
        RECT 0.140 2611.130 2262.720 2612.830 ;
        RECT 1.140 2610.310 2262.060 2611.130 ;
        RECT 0.140 2608.610 2262.720 2610.310 ;
        RECT 0.140 2607.790 2262.060 2608.610 ;
        RECT 0.140 2606.090 2262.720 2607.790 ;
        RECT 1.140 2605.270 2262.060 2606.090 ;
        RECT 0.140 2603.570 2262.720 2605.270 ;
        RECT 0.140 2602.750 2262.060 2603.570 ;
        RECT 0.140 2601.050 2262.720 2602.750 ;
        RECT 1.140 2600.230 2262.060 2601.050 ;
        RECT 0.140 2598.530 2262.720 2600.230 ;
        RECT 0.140 2597.710 2262.060 2598.530 ;
        RECT 0.140 2596.010 2262.720 2597.710 ;
        RECT 1.070 2595.190 2262.060 2596.010 ;
        RECT 0.140 2593.490 2262.720 2595.190 ;
        RECT 0.140 2592.670 2262.060 2593.490 ;
        RECT 0.140 2590.970 2262.720 2592.670 ;
        RECT 1.140 2590.150 2262.060 2590.970 ;
        RECT 0.140 2588.450 2262.720 2590.150 ;
        RECT 0.140 2587.630 2262.130 2588.450 ;
        RECT 0.140 2585.930 2262.720 2587.630 ;
        RECT 1.070 2585.110 2262.060 2585.930 ;
        RECT 0.140 2583.410 2262.720 2585.110 ;
        RECT 0.140 2582.590 2262.060 2583.410 ;
        RECT 0.140 2580.890 2262.720 2582.590 ;
        RECT 1.070 2580.070 2262.060 2580.890 ;
        RECT 0.140 2578.370 2262.720 2580.070 ;
        RECT 0.140 2577.550 2262.060 2578.370 ;
        RECT 0.140 2575.850 2262.720 2577.550 ;
        RECT 1.070 2575.030 2262.060 2575.850 ;
        RECT 0.140 2573.330 2262.720 2575.030 ;
        RECT 0.140 2572.510 2262.060 2573.330 ;
        RECT 0.140 2570.810 2262.720 2572.510 ;
        RECT 1.070 2569.990 2262.060 2570.810 ;
        RECT 0.140 2568.290 2262.720 2569.990 ;
        RECT 0.140 2567.470 2262.060 2568.290 ;
        RECT 0.140 2565.770 2262.720 2567.470 ;
        RECT 1.070 2564.950 2262.060 2565.770 ;
        RECT 0.140 2563.250 2262.720 2564.950 ;
        RECT 0.140 2562.430 2262.060 2563.250 ;
        RECT 0.140 2560.730 2262.720 2562.430 ;
        RECT 1.140 2559.910 2262.060 2560.730 ;
        RECT 0.140 2558.210 2262.720 2559.910 ;
        RECT 0.140 2557.390 2262.060 2558.210 ;
        RECT 0.140 2555.690 2262.720 2557.390 ;
        RECT 1.140 2554.870 2262.060 2555.690 ;
        RECT 0.140 2553.170 2262.720 2554.870 ;
        RECT 0.140 2552.350 2262.060 2553.170 ;
        RECT 0.140 2550.650 2262.720 2552.350 ;
        RECT 1.070 2549.830 2262.060 2550.650 ;
        RECT 0.140 2548.130 2262.720 2549.830 ;
        RECT 0.140 2547.310 2262.060 2548.130 ;
        RECT 0.140 2545.610 2262.720 2547.310 ;
        RECT 1.140 2544.790 2262.060 2545.610 ;
        RECT 0.140 2543.090 2262.720 2544.790 ;
        RECT 0.140 2542.270 2262.060 2543.090 ;
        RECT 0.140 2540.570 2262.720 2542.270 ;
        RECT 1.140 2539.750 2262.060 2540.570 ;
        RECT 0.140 2538.050 2262.720 2539.750 ;
        RECT 0.140 2537.230 2262.060 2538.050 ;
        RECT 0.140 2535.530 2262.720 2537.230 ;
        RECT 1.140 2534.710 2262.060 2535.530 ;
        RECT 0.140 2533.010 2262.720 2534.710 ;
        RECT 0.140 2532.190 2262.060 2533.010 ;
        RECT 0.140 2530.490 2262.720 2532.190 ;
        RECT 1.070 2529.670 2262.060 2530.490 ;
        RECT 0.140 2527.970 2262.720 2529.670 ;
        RECT 0.140 2527.150 2262.060 2527.970 ;
        RECT 0.140 2525.450 2262.720 2527.150 ;
        RECT 1.140 2524.630 2262.060 2525.450 ;
        RECT 0.140 2522.930 2262.720 2524.630 ;
        RECT 0.140 2522.110 2262.060 2522.930 ;
        RECT 0.140 2520.410 2262.720 2522.110 ;
        RECT 1.140 2519.590 2262.060 2520.410 ;
        RECT 0.140 2517.890 2262.720 2519.590 ;
        RECT 0.140 2517.070 2262.060 2517.890 ;
        RECT 0.140 2515.370 2262.720 2517.070 ;
        RECT 1.140 2514.550 2262.060 2515.370 ;
        RECT 0.140 2512.850 2262.720 2514.550 ;
        RECT 0.140 2512.030 2262.060 2512.850 ;
        RECT 0.140 2510.330 2262.720 2512.030 ;
        RECT 1.140 2509.510 2262.060 2510.330 ;
        RECT 0.140 2507.810 2262.720 2509.510 ;
        RECT 0.140 2506.990 2262.060 2507.810 ;
        RECT 0.140 2505.290 2262.720 2506.990 ;
        RECT 1.140 2504.470 2262.060 2505.290 ;
        RECT 0.140 2502.770 2262.720 2504.470 ;
        RECT 0.140 2501.950 2262.060 2502.770 ;
        RECT 0.140 2500.250 2262.720 2501.950 ;
        RECT 1.070 2499.430 2262.720 2500.250 ;
        RECT 0.140 2495.210 2262.720 2499.430 ;
        RECT 1.140 2494.390 2262.720 2495.210 ;
        RECT 0.140 2490.170 2262.720 2494.390 ;
        RECT 1.070 2489.350 2262.720 2490.170 ;
        RECT 0.140 2475.050 2262.720 2489.350 ;
        RECT 1.140 2474.230 2262.720 2475.050 ;
        RECT 0.140 2470.010 2262.720 2474.230 ;
        RECT 1.140 2469.190 2262.720 2470.010 ;
        RECT 0.140 2464.970 2262.720 2469.190 ;
        RECT 1.070 2464.150 2262.720 2464.970 ;
        RECT 0.140 2459.930 2262.720 2464.150 ;
        RECT 1.070 2459.110 2262.720 2459.930 ;
        RECT 0.140 2454.890 2262.720 2459.110 ;
        RECT 1.140 2454.070 2262.720 2454.890 ;
        RECT 0.140 2449.850 2262.720 2454.070 ;
        RECT 1.070 2449.030 2262.720 2449.850 ;
        RECT 0.140 2444.810 2262.720 2449.030 ;
        RECT 1.070 2443.990 2262.720 2444.810 ;
        RECT 0.140 2439.770 2262.720 2443.990 ;
        RECT 1.140 2438.950 2262.720 2439.770 ;
        RECT 0.140 2434.730 2262.720 2438.950 ;
        RECT 1.070 2433.910 2262.720 2434.730 ;
        RECT 0.140 2429.690 2262.720 2433.910 ;
        RECT 1.070 2428.870 2262.720 2429.690 ;
        RECT 0.140 2424.650 2262.720 2428.870 ;
        RECT 1.140 2423.830 2262.720 2424.650 ;
        RECT 0.140 2419.610 2262.720 2423.830 ;
        RECT 1.070 2418.790 2262.720 2419.610 ;
        RECT 0.140 2414.570 2262.720 2418.790 ;
        RECT 1.070 2413.750 2262.720 2414.570 ;
        RECT 0.140 2409.530 2262.720 2413.750 ;
        RECT 1.140 2408.710 2262.720 2409.530 ;
        RECT 0.140 2404.490 2262.720 2408.710 ;
        RECT 1.070 2403.670 2262.720 2404.490 ;
        RECT 0.140 2399.450 2262.720 2403.670 ;
        RECT 1.070 2398.630 2262.720 2399.450 ;
        RECT 0.140 2394.410 2262.720 2398.630 ;
        RECT 1.140 2393.590 2262.720 2394.410 ;
        RECT 0.140 2389.370 2262.720 2393.590 ;
        RECT 1.070 2388.550 2262.720 2389.370 ;
        RECT 0.140 2384.330 2262.720 2388.550 ;
        RECT 1.070 2383.510 2262.720 2384.330 ;
        RECT 0.140 2379.290 2262.720 2383.510 ;
        RECT 1.140 2378.470 2262.720 2379.290 ;
        RECT 0.140 2374.250 2262.720 2378.470 ;
        RECT 1.140 2373.430 2262.720 2374.250 ;
        RECT 0.140 2369.210 2262.720 2373.430 ;
        RECT 1.140 2368.390 2262.720 2369.210 ;
        RECT 0.140 2364.170 2262.720 2368.390 ;
        RECT 1.140 2363.350 2262.720 2364.170 ;
        RECT 0.140 2359.130 2262.720 2363.350 ;
        RECT 1.140 2358.310 2262.720 2359.130 ;
        RECT 0.140 2354.090 2262.720 2358.310 ;
        RECT 1.070 2353.270 2262.720 2354.090 ;
        RECT 0.140 2349.050 2262.720 2353.270 ;
        RECT 1.140 2348.230 2262.720 2349.050 ;
        RECT 0.140 2344.010 2262.720 2348.230 ;
        RECT 1.070 2343.190 2262.720 2344.010 ;
        RECT 0.140 2338.970 2262.720 2343.190 ;
        RECT 1.070 2338.150 2262.720 2338.970 ;
        RECT 0.140 2333.930 2262.720 2338.150 ;
        RECT 1.070 2333.110 2262.720 2333.930 ;
        RECT 0.140 2328.890 2262.720 2333.110 ;
        RECT 1.070 2328.070 2262.720 2328.890 ;
        RECT 0.140 2323.850 2262.720 2328.070 ;
        RECT 1.070 2323.030 2262.720 2323.850 ;
        RECT 0.140 2318.810 2262.720 2323.030 ;
        RECT 1.140 2317.990 2262.720 2318.810 ;
        RECT 0.140 2313.770 2262.720 2317.990 ;
        RECT 1.140 2312.950 2262.720 2313.770 ;
        RECT 0.140 2308.730 2262.720 2312.950 ;
        RECT 1.070 2307.910 2262.720 2308.730 ;
        RECT 0.140 2303.690 2262.720 2307.910 ;
        RECT 1.140 2302.870 2262.720 2303.690 ;
        RECT 0.140 2301.170 2262.720 2302.870 ;
        RECT 0.140 2300.350 2262.060 2301.170 ;
        RECT 0.140 2298.650 2262.720 2300.350 ;
        RECT 1.140 2297.830 2262.060 2298.650 ;
        RECT 0.140 2296.130 2262.720 2297.830 ;
        RECT 0.140 2295.310 2262.060 2296.130 ;
        RECT 0.140 2293.610 2262.720 2295.310 ;
        RECT 1.140 2292.790 2262.060 2293.610 ;
        RECT 0.140 2291.090 2262.720 2292.790 ;
        RECT 0.140 2290.270 2262.060 2291.090 ;
        RECT 0.140 2288.570 2262.720 2290.270 ;
        RECT 1.070 2287.750 2262.060 2288.570 ;
        RECT 0.140 2286.050 2262.720 2287.750 ;
        RECT 0.140 2285.230 2262.060 2286.050 ;
        RECT 0.140 2283.530 2262.720 2285.230 ;
        RECT 1.140 2282.710 2262.060 2283.530 ;
        RECT 0.140 2281.010 2262.720 2282.710 ;
        RECT 0.140 2280.190 2262.060 2281.010 ;
        RECT 0.140 2278.490 2262.720 2280.190 ;
        RECT 1.140 2277.670 2262.060 2278.490 ;
        RECT 0.140 2275.970 2262.720 2277.670 ;
        RECT 0.140 2275.150 2262.060 2275.970 ;
        RECT 0.140 2273.450 2262.720 2275.150 ;
        RECT 1.140 2272.630 2262.060 2273.450 ;
        RECT 0.140 2270.930 2262.720 2272.630 ;
        RECT 0.140 2270.110 2262.060 2270.930 ;
        RECT 0.140 2268.410 2262.720 2270.110 ;
        RECT 1.140 2267.590 2262.060 2268.410 ;
        RECT 0.140 2265.890 2262.720 2267.590 ;
        RECT 0.140 2265.070 2262.060 2265.890 ;
        RECT 0.140 2263.370 2262.720 2265.070 ;
        RECT 1.140 2262.550 2262.060 2263.370 ;
        RECT 0.140 2260.850 2262.720 2262.550 ;
        RECT 0.140 2260.030 2262.060 2260.850 ;
        RECT 0.140 2258.330 2262.720 2260.030 ;
        RECT 1.070 2257.510 2262.060 2258.330 ;
        RECT 0.140 2255.810 2262.720 2257.510 ;
        RECT 0.140 2254.990 2262.060 2255.810 ;
        RECT 0.140 2253.290 2262.720 2254.990 ;
        RECT 1.140 2252.470 2262.060 2253.290 ;
        RECT 0.140 2250.770 2262.720 2252.470 ;
        RECT 0.140 2249.950 2262.060 2250.770 ;
        RECT 0.140 2248.250 2262.720 2249.950 ;
        RECT 1.070 2247.430 2262.060 2248.250 ;
        RECT 0.140 2245.730 2262.720 2247.430 ;
        RECT 0.140 2244.910 2262.060 2245.730 ;
        RECT 0.140 2243.210 2262.720 2244.910 ;
        RECT 0.140 2242.390 2262.060 2243.210 ;
        RECT 0.140 2240.690 2262.720 2242.390 ;
        RECT 0.140 2239.870 2262.060 2240.690 ;
        RECT 0.140 2238.170 2262.720 2239.870 ;
        RECT 0.140 2237.350 2262.060 2238.170 ;
        RECT 0.140 2235.650 2262.720 2237.350 ;
        RECT 0.140 2234.830 2262.060 2235.650 ;
        RECT 0.140 2233.130 2262.720 2234.830 ;
        RECT 1.140 2232.310 2262.060 2233.130 ;
        RECT 0.140 2230.610 2262.720 2232.310 ;
        RECT 0.140 2229.790 2262.060 2230.610 ;
        RECT 0.140 2228.090 2262.720 2229.790 ;
        RECT 1.140 2227.270 2262.060 2228.090 ;
        RECT 0.140 2225.570 2262.720 2227.270 ;
        RECT 0.140 2224.750 2262.060 2225.570 ;
        RECT 0.140 2223.050 2262.720 2224.750 ;
        RECT 1.070 2222.230 2262.060 2223.050 ;
        RECT 0.140 2220.530 2262.720 2222.230 ;
        RECT 0.140 2219.710 2262.060 2220.530 ;
        RECT 0.140 2218.010 2262.720 2219.710 ;
        RECT 1.070 2217.190 2262.060 2218.010 ;
        RECT 0.140 2215.490 2262.720 2217.190 ;
        RECT 0.140 2214.670 2262.060 2215.490 ;
        RECT 0.140 2212.970 2262.720 2214.670 ;
        RECT 1.140 2212.150 2262.060 2212.970 ;
        RECT 0.140 2210.450 2262.720 2212.150 ;
        RECT 0.140 2209.630 2262.060 2210.450 ;
        RECT 0.140 2207.930 2262.720 2209.630 ;
        RECT 1.070 2207.110 2262.060 2207.930 ;
        RECT 0.140 2205.410 2262.720 2207.110 ;
        RECT 0.140 2204.590 2262.060 2205.410 ;
        RECT 0.140 2202.890 2262.720 2204.590 ;
        RECT 1.070 2202.070 2262.060 2202.890 ;
        RECT 0.140 2200.370 2262.720 2202.070 ;
        RECT 0.140 2199.550 2262.060 2200.370 ;
        RECT 0.140 2197.850 2262.720 2199.550 ;
        RECT 1.140 2197.030 2262.060 2197.850 ;
        RECT 0.140 2195.330 2262.720 2197.030 ;
        RECT 0.140 2194.510 2262.060 2195.330 ;
        RECT 0.140 2192.810 2262.720 2194.510 ;
        RECT 1.070 2191.990 2262.060 2192.810 ;
        RECT 0.140 2190.290 2262.720 2191.990 ;
        RECT 0.140 2189.470 2262.060 2190.290 ;
        RECT 0.140 2187.770 2262.720 2189.470 ;
        RECT 1.070 2186.950 2262.060 2187.770 ;
        RECT 0.140 2185.250 2262.720 2186.950 ;
        RECT 0.140 2184.430 2262.060 2185.250 ;
        RECT 0.140 2182.730 2262.720 2184.430 ;
        RECT 1.140 2181.910 2262.060 2182.730 ;
        RECT 0.140 2180.210 2262.720 2181.910 ;
        RECT 0.140 2179.390 2262.060 2180.210 ;
        RECT 0.140 2177.690 2262.720 2179.390 ;
        RECT 1.070 2176.870 2262.060 2177.690 ;
        RECT 0.140 2175.170 2262.720 2176.870 ;
        RECT 0.140 2174.350 2262.060 2175.170 ;
        RECT 0.140 2172.650 2262.720 2174.350 ;
        RECT 1.070 2171.830 2262.060 2172.650 ;
        RECT 0.140 2170.130 2262.720 2171.830 ;
        RECT 0.140 2169.310 2262.060 2170.130 ;
        RECT 0.140 2167.610 2262.720 2169.310 ;
        RECT 1.140 2166.790 2262.060 2167.610 ;
        RECT 0.140 2165.090 2262.720 2166.790 ;
        RECT 0.140 2164.270 2262.060 2165.090 ;
        RECT 0.140 2162.570 2262.720 2164.270 ;
        RECT 1.070 2161.750 2262.060 2162.570 ;
        RECT 0.140 2160.050 2262.720 2161.750 ;
        RECT 0.140 2159.230 2262.060 2160.050 ;
        RECT 0.140 2157.530 2262.720 2159.230 ;
        RECT 1.070 2156.710 2262.060 2157.530 ;
        RECT 0.140 2155.010 2262.720 2156.710 ;
        RECT 0.140 2154.190 2262.060 2155.010 ;
        RECT 0.140 2152.490 2262.720 2154.190 ;
        RECT 1.140 2151.670 2262.060 2152.490 ;
        RECT 0.140 2149.970 2262.720 2151.670 ;
        RECT 0.140 2149.150 2262.060 2149.970 ;
        RECT 0.140 2147.450 2262.720 2149.150 ;
        RECT 1.070 2146.630 2262.060 2147.450 ;
        RECT 0.140 2144.930 2262.720 2146.630 ;
        RECT 0.140 2144.110 2262.060 2144.930 ;
        RECT 0.140 2142.410 2262.720 2144.110 ;
        RECT 1.070 2141.590 2262.060 2142.410 ;
        RECT 0.140 2139.890 2262.720 2141.590 ;
        RECT 0.140 2139.070 2262.060 2139.890 ;
        RECT 0.140 2137.370 2262.720 2139.070 ;
        RECT 1.140 2136.550 2262.060 2137.370 ;
        RECT 0.140 2134.850 2262.720 2136.550 ;
        RECT 0.140 2134.030 2262.060 2134.850 ;
        RECT 0.140 2132.330 2262.720 2134.030 ;
        RECT 1.140 2131.510 2262.060 2132.330 ;
        RECT 0.140 2129.810 2262.720 2131.510 ;
        RECT 0.140 2128.990 2262.060 2129.810 ;
        RECT 0.140 2127.290 2262.720 2128.990 ;
        RECT 1.140 2126.470 2262.060 2127.290 ;
        RECT 0.140 2124.770 2262.720 2126.470 ;
        RECT 0.140 2123.950 2262.060 2124.770 ;
        RECT 0.140 2122.250 2262.720 2123.950 ;
        RECT 1.140 2121.430 2262.060 2122.250 ;
        RECT 0.140 2119.730 2262.720 2121.430 ;
        RECT 0.140 2118.910 2262.060 2119.730 ;
        RECT 0.140 2117.210 2262.720 2118.910 ;
        RECT 1.140 2116.390 2262.060 2117.210 ;
        RECT 0.140 2114.690 2262.720 2116.390 ;
        RECT 0.140 2113.870 2262.060 2114.690 ;
        RECT 0.140 2112.170 2262.720 2113.870 ;
        RECT 1.070 2111.350 2262.060 2112.170 ;
        RECT 0.140 2109.650 2262.720 2111.350 ;
        RECT 0.140 2108.830 2262.060 2109.650 ;
        RECT 0.140 2107.130 2262.720 2108.830 ;
        RECT 1.140 2106.310 2262.060 2107.130 ;
        RECT 0.140 2104.610 2262.720 2106.310 ;
        RECT 0.140 2103.790 2262.130 2104.610 ;
        RECT 0.140 2102.090 2262.720 2103.790 ;
        RECT 1.070 2101.270 2262.060 2102.090 ;
        RECT 0.140 2099.570 2262.720 2101.270 ;
        RECT 0.140 2098.750 2262.060 2099.570 ;
        RECT 0.140 2097.050 2262.720 2098.750 ;
        RECT 1.070 2096.230 2262.060 2097.050 ;
        RECT 0.140 2094.530 2262.720 2096.230 ;
        RECT 0.140 2093.710 2262.060 2094.530 ;
        RECT 0.140 2092.010 2262.720 2093.710 ;
        RECT 1.070 2091.190 2262.060 2092.010 ;
        RECT 0.140 2089.490 2262.720 2091.190 ;
        RECT 0.140 2088.670 2262.060 2089.490 ;
        RECT 0.140 2086.970 2262.720 2088.670 ;
        RECT 1.070 2086.150 2262.060 2086.970 ;
        RECT 0.140 2084.450 2262.720 2086.150 ;
        RECT 0.140 2083.630 2262.060 2084.450 ;
        RECT 0.140 2081.930 2262.720 2083.630 ;
        RECT 1.070 2081.110 2262.060 2081.930 ;
        RECT 0.140 2079.410 2262.720 2081.110 ;
        RECT 0.140 2078.590 2262.060 2079.410 ;
        RECT 0.140 2076.890 2262.720 2078.590 ;
        RECT 1.140 2076.070 2262.060 2076.890 ;
        RECT 0.140 2074.370 2262.720 2076.070 ;
        RECT 0.140 2073.550 2262.060 2074.370 ;
        RECT 0.140 2071.850 2262.720 2073.550 ;
        RECT 1.140 2071.030 2262.060 2071.850 ;
        RECT 0.140 2069.330 2262.720 2071.030 ;
        RECT 0.140 2068.510 2262.060 2069.330 ;
        RECT 0.140 2066.810 2262.720 2068.510 ;
        RECT 1.070 2065.990 2262.060 2066.810 ;
        RECT 0.140 2064.290 2262.720 2065.990 ;
        RECT 0.140 2063.470 2262.060 2064.290 ;
        RECT 0.140 2061.770 2262.720 2063.470 ;
        RECT 1.140 2060.950 2262.060 2061.770 ;
        RECT 0.140 2059.250 2262.720 2060.950 ;
        RECT 0.140 2058.430 2262.060 2059.250 ;
        RECT 0.140 2056.730 2262.720 2058.430 ;
        RECT 1.140 2055.910 2262.060 2056.730 ;
        RECT 0.140 2054.210 2262.720 2055.910 ;
        RECT 0.140 2053.390 2262.060 2054.210 ;
        RECT 0.140 2051.690 2262.720 2053.390 ;
        RECT 1.140 2050.870 2262.060 2051.690 ;
        RECT 0.140 2049.170 2262.720 2050.870 ;
        RECT 0.140 2048.350 2262.060 2049.170 ;
        RECT 0.140 2046.650 2262.720 2048.350 ;
        RECT 1.070 2045.830 2262.060 2046.650 ;
        RECT 0.140 2044.130 2262.720 2045.830 ;
        RECT 0.140 2043.310 2262.060 2044.130 ;
        RECT 0.140 2041.610 2262.720 2043.310 ;
        RECT 1.140 2040.790 2262.060 2041.610 ;
        RECT 0.140 2039.090 2262.720 2040.790 ;
        RECT 0.140 2038.270 2262.060 2039.090 ;
        RECT 0.140 2036.570 2262.720 2038.270 ;
        RECT 1.140 2035.750 2262.060 2036.570 ;
        RECT 0.140 2034.050 2262.720 2035.750 ;
        RECT 0.140 2033.230 2262.060 2034.050 ;
        RECT 0.140 2031.530 2262.720 2033.230 ;
        RECT 1.140 2030.710 2262.060 2031.530 ;
        RECT 0.140 2029.010 2262.720 2030.710 ;
        RECT 0.140 2028.190 2262.060 2029.010 ;
        RECT 0.140 2026.490 2262.720 2028.190 ;
        RECT 1.140 2025.670 2262.060 2026.490 ;
        RECT 0.140 2023.970 2262.720 2025.670 ;
        RECT 0.140 2023.150 2262.060 2023.970 ;
        RECT 0.140 2021.450 2262.720 2023.150 ;
        RECT 1.140 2020.630 2262.060 2021.450 ;
        RECT 0.140 2018.930 2262.720 2020.630 ;
        RECT 0.140 2018.110 2262.060 2018.930 ;
        RECT 0.140 2016.410 2262.720 2018.110 ;
        RECT 1.070 2015.590 2262.720 2016.410 ;
        RECT 0.140 2011.370 2262.720 2015.590 ;
        RECT 1.140 2010.550 2262.720 2011.370 ;
        RECT 0.140 2006.330 2262.720 2010.550 ;
        RECT 1.070 2005.510 2262.720 2006.330 ;
        RECT 0.140 1991.210 2262.720 2005.510 ;
        RECT 1.140 1990.390 2262.720 1991.210 ;
        RECT 0.140 1986.170 2262.720 1990.390 ;
        RECT 1.140 1985.350 2262.720 1986.170 ;
        RECT 0.140 1981.130 2262.720 1985.350 ;
        RECT 1.070 1980.310 2262.720 1981.130 ;
        RECT 0.140 1976.090 2262.720 1980.310 ;
        RECT 1.070 1975.270 2262.720 1976.090 ;
        RECT 0.140 1971.050 2262.720 1975.270 ;
        RECT 1.140 1970.230 2262.720 1971.050 ;
        RECT 0.140 1966.010 2262.720 1970.230 ;
        RECT 1.070 1965.190 2262.720 1966.010 ;
        RECT 0.140 1960.970 2262.720 1965.190 ;
        RECT 1.070 1960.150 2262.720 1960.970 ;
        RECT 0.140 1955.930 2262.720 1960.150 ;
        RECT 1.140 1955.110 2262.720 1955.930 ;
        RECT 0.140 1950.890 2262.720 1955.110 ;
        RECT 1.070 1950.070 2262.720 1950.890 ;
        RECT 0.140 1945.850 2262.720 1950.070 ;
        RECT 1.070 1945.030 2262.720 1945.850 ;
        RECT 0.140 1940.810 2262.720 1945.030 ;
        RECT 1.140 1939.990 2262.720 1940.810 ;
        RECT 0.140 1935.770 2262.720 1939.990 ;
        RECT 1.070 1934.950 2262.720 1935.770 ;
        RECT 0.140 1930.730 2262.720 1934.950 ;
        RECT 1.070 1929.910 2262.720 1930.730 ;
        RECT 0.140 1925.690 2262.720 1929.910 ;
        RECT 1.140 1924.870 2262.720 1925.690 ;
        RECT 0.140 1920.650 2262.720 1924.870 ;
        RECT 1.070 1919.830 2262.720 1920.650 ;
        RECT 0.140 1915.610 2262.720 1919.830 ;
        RECT 1.070 1914.790 2262.720 1915.610 ;
        RECT 0.140 1910.570 2262.720 1914.790 ;
        RECT 1.140 1909.750 2262.720 1910.570 ;
        RECT 0.140 1905.530 2262.720 1909.750 ;
        RECT 1.070 1904.710 2262.720 1905.530 ;
        RECT 0.140 1900.490 2262.720 1904.710 ;
        RECT 1.070 1899.670 2262.720 1900.490 ;
        RECT 0.140 1895.450 2262.720 1899.670 ;
        RECT 1.140 1894.630 2262.720 1895.450 ;
        RECT 0.140 1890.410 2262.720 1894.630 ;
        RECT 1.140 1889.590 2262.720 1890.410 ;
        RECT 0.140 1885.370 2262.720 1889.590 ;
        RECT 1.140 1884.550 2262.720 1885.370 ;
        RECT 0.140 1880.330 2262.720 1884.550 ;
        RECT 1.140 1879.510 2262.720 1880.330 ;
        RECT 0.140 1875.290 2262.720 1879.510 ;
        RECT 1.140 1874.470 2262.720 1875.290 ;
        RECT 0.140 1870.250 2262.720 1874.470 ;
        RECT 1.070 1869.430 2262.720 1870.250 ;
        RECT 0.140 1865.210 2262.720 1869.430 ;
        RECT 1.140 1864.390 2262.720 1865.210 ;
        RECT 0.140 1860.170 2262.720 1864.390 ;
        RECT 1.070 1859.350 2262.720 1860.170 ;
        RECT 0.140 1855.130 2262.720 1859.350 ;
        RECT 1.070 1854.310 2262.720 1855.130 ;
        RECT 0.140 1850.090 2262.720 1854.310 ;
        RECT 1.070 1849.270 2262.720 1850.090 ;
        RECT 0.140 1845.050 2262.720 1849.270 ;
        RECT 1.070 1844.230 2262.720 1845.050 ;
        RECT 0.140 1840.010 2262.720 1844.230 ;
        RECT 1.070 1839.190 2262.720 1840.010 ;
        RECT 0.140 1834.970 2262.720 1839.190 ;
        RECT 1.140 1834.150 2262.720 1834.970 ;
        RECT 0.140 1829.930 2262.720 1834.150 ;
        RECT 1.140 1829.110 2262.720 1829.930 ;
        RECT 0.140 1824.890 2262.720 1829.110 ;
        RECT 1.070 1824.070 2262.720 1824.890 ;
        RECT 0.140 1819.850 2262.720 1824.070 ;
        RECT 1.140 1819.030 2262.720 1819.850 ;
        RECT 0.140 1817.330 2262.720 1819.030 ;
        RECT 0.140 1816.510 2262.060 1817.330 ;
        RECT 0.140 1814.810 2262.720 1816.510 ;
        RECT 1.140 1813.990 2262.060 1814.810 ;
        RECT 0.140 1812.290 2262.720 1813.990 ;
        RECT 0.140 1811.470 2262.060 1812.290 ;
        RECT 0.140 1809.770 2262.720 1811.470 ;
        RECT 1.140 1808.950 2262.060 1809.770 ;
        RECT 0.140 1807.250 2262.720 1808.950 ;
        RECT 0.140 1806.430 2262.060 1807.250 ;
        RECT 0.140 1804.730 2262.720 1806.430 ;
        RECT 1.070 1803.910 2262.060 1804.730 ;
        RECT 0.140 1802.210 2262.720 1803.910 ;
        RECT 0.140 1801.390 2262.060 1802.210 ;
        RECT 0.140 1799.690 2262.720 1801.390 ;
        RECT 1.140 1798.870 2262.060 1799.690 ;
        RECT 0.140 1797.170 2262.720 1798.870 ;
        RECT 0.140 1796.350 2262.060 1797.170 ;
        RECT 0.140 1794.650 2262.720 1796.350 ;
        RECT 1.140 1793.830 2262.060 1794.650 ;
        RECT 0.140 1792.130 2262.720 1793.830 ;
        RECT 0.140 1791.310 2262.060 1792.130 ;
        RECT 0.140 1789.610 2262.720 1791.310 ;
        RECT 1.140 1788.790 2262.060 1789.610 ;
        RECT 0.140 1787.090 2262.720 1788.790 ;
        RECT 0.140 1786.270 2262.060 1787.090 ;
        RECT 0.140 1784.570 2262.720 1786.270 ;
        RECT 1.140 1783.750 2262.060 1784.570 ;
        RECT 0.140 1782.050 2262.720 1783.750 ;
        RECT 0.140 1781.230 2262.060 1782.050 ;
        RECT 0.140 1779.530 2262.720 1781.230 ;
        RECT 1.140 1778.710 2262.060 1779.530 ;
        RECT 0.140 1777.010 2262.720 1778.710 ;
        RECT 0.140 1776.190 2262.060 1777.010 ;
        RECT 0.140 1774.490 2262.720 1776.190 ;
        RECT 1.070 1773.670 2262.060 1774.490 ;
        RECT 0.140 1771.970 2262.720 1773.670 ;
        RECT 0.140 1771.150 2262.060 1771.970 ;
        RECT 0.140 1769.450 2262.720 1771.150 ;
        RECT 1.140 1768.630 2262.060 1769.450 ;
        RECT 0.140 1766.930 2262.720 1768.630 ;
        RECT 0.140 1766.110 2262.060 1766.930 ;
        RECT 0.140 1764.410 2262.720 1766.110 ;
        RECT 1.070 1763.590 2262.060 1764.410 ;
        RECT 0.140 1761.890 2262.720 1763.590 ;
        RECT 0.140 1761.070 2262.060 1761.890 ;
        RECT 0.140 1759.370 2262.720 1761.070 ;
        RECT 0.140 1758.550 2262.060 1759.370 ;
        RECT 0.140 1756.850 2262.720 1758.550 ;
        RECT 0.140 1756.030 2262.060 1756.850 ;
        RECT 0.140 1754.330 2262.720 1756.030 ;
        RECT 0.140 1753.510 2262.060 1754.330 ;
        RECT 0.140 1751.810 2262.720 1753.510 ;
        RECT 0.140 1750.990 2262.060 1751.810 ;
        RECT 0.140 1749.290 2262.720 1750.990 ;
        RECT 1.140 1748.470 2262.060 1749.290 ;
        RECT 0.140 1746.770 2262.720 1748.470 ;
        RECT 0.140 1745.950 2262.060 1746.770 ;
        RECT 0.140 1744.250 2262.720 1745.950 ;
        RECT 1.140 1743.430 2262.060 1744.250 ;
        RECT 0.140 1741.730 2262.720 1743.430 ;
        RECT 0.140 1740.910 2262.060 1741.730 ;
        RECT 0.140 1739.210 2262.720 1740.910 ;
        RECT 1.070 1738.390 2262.060 1739.210 ;
        RECT 0.140 1736.690 2262.720 1738.390 ;
        RECT 0.140 1735.870 2262.060 1736.690 ;
        RECT 0.140 1734.170 2262.720 1735.870 ;
        RECT 1.070 1733.350 2262.060 1734.170 ;
        RECT 0.140 1731.650 2262.720 1733.350 ;
        RECT 0.140 1730.830 2262.060 1731.650 ;
        RECT 0.140 1729.130 2262.720 1730.830 ;
        RECT 1.140 1728.310 2262.060 1729.130 ;
        RECT 0.140 1726.610 2262.720 1728.310 ;
        RECT 0.140 1725.790 2262.060 1726.610 ;
        RECT 0.140 1724.090 2262.720 1725.790 ;
        RECT 1.070 1723.270 2262.060 1724.090 ;
        RECT 0.140 1721.570 2262.720 1723.270 ;
        RECT 0.140 1720.750 2262.060 1721.570 ;
        RECT 0.140 1719.050 2262.720 1720.750 ;
        RECT 1.070 1718.230 2262.060 1719.050 ;
        RECT 0.140 1716.530 2262.720 1718.230 ;
        RECT 0.140 1715.710 2262.060 1716.530 ;
        RECT 0.140 1714.010 2262.720 1715.710 ;
        RECT 1.140 1713.190 2262.060 1714.010 ;
        RECT 0.140 1711.490 2262.720 1713.190 ;
        RECT 0.140 1710.670 2262.060 1711.490 ;
        RECT 0.140 1708.970 2262.720 1710.670 ;
        RECT 1.070 1708.150 2262.060 1708.970 ;
        RECT 0.140 1706.450 2262.720 1708.150 ;
        RECT 0.140 1705.630 2262.060 1706.450 ;
        RECT 0.140 1703.930 2262.720 1705.630 ;
        RECT 1.070 1703.110 2262.060 1703.930 ;
        RECT 0.140 1701.410 2262.720 1703.110 ;
        RECT 0.140 1700.590 2262.060 1701.410 ;
        RECT 0.140 1698.890 2262.720 1700.590 ;
        RECT 1.140 1698.070 2262.060 1698.890 ;
        RECT 0.140 1696.370 2262.720 1698.070 ;
        RECT 0.140 1695.550 2262.060 1696.370 ;
        RECT 0.140 1693.850 2262.720 1695.550 ;
        RECT 1.070 1693.030 2262.060 1693.850 ;
        RECT 0.140 1691.330 2262.720 1693.030 ;
        RECT 0.140 1690.510 2262.060 1691.330 ;
        RECT 0.140 1688.810 2262.720 1690.510 ;
        RECT 1.070 1687.990 2262.060 1688.810 ;
        RECT 0.140 1686.290 2262.720 1687.990 ;
        RECT 0.140 1685.470 2262.060 1686.290 ;
        RECT 0.140 1683.770 2262.720 1685.470 ;
        RECT 1.140 1682.950 2262.060 1683.770 ;
        RECT 0.140 1681.250 2262.720 1682.950 ;
        RECT 0.140 1680.430 2262.060 1681.250 ;
        RECT 0.140 1678.730 2262.720 1680.430 ;
        RECT 1.070 1677.910 2262.060 1678.730 ;
        RECT 0.140 1676.210 2262.720 1677.910 ;
        RECT 0.140 1675.390 2262.060 1676.210 ;
        RECT 0.140 1673.690 2262.720 1675.390 ;
        RECT 1.070 1672.870 2262.060 1673.690 ;
        RECT 0.140 1671.170 2262.720 1672.870 ;
        RECT 0.140 1670.350 2262.060 1671.170 ;
        RECT 0.140 1668.650 2262.720 1670.350 ;
        RECT 1.140 1667.830 2262.060 1668.650 ;
        RECT 0.140 1666.130 2262.720 1667.830 ;
        RECT 0.140 1665.310 2262.060 1666.130 ;
        RECT 0.140 1663.610 2262.720 1665.310 ;
        RECT 1.070 1662.790 2262.060 1663.610 ;
        RECT 0.140 1661.090 2262.720 1662.790 ;
        RECT 0.140 1660.270 2262.060 1661.090 ;
        RECT 0.140 1658.570 2262.720 1660.270 ;
        RECT 1.070 1657.750 2262.060 1658.570 ;
        RECT 0.140 1656.050 2262.720 1657.750 ;
        RECT 0.140 1655.230 2262.060 1656.050 ;
        RECT 0.140 1653.530 2262.720 1655.230 ;
        RECT 1.140 1652.710 2262.060 1653.530 ;
        RECT 0.140 1651.010 2262.720 1652.710 ;
        RECT 0.140 1650.190 2262.060 1651.010 ;
        RECT 0.140 1648.490 2262.720 1650.190 ;
        RECT 1.140 1647.670 2262.060 1648.490 ;
        RECT 0.140 1645.970 2262.720 1647.670 ;
        RECT 0.140 1645.150 2262.060 1645.970 ;
        RECT 0.140 1643.450 2262.720 1645.150 ;
        RECT 1.140 1642.630 2262.060 1643.450 ;
        RECT 0.140 1640.930 2262.720 1642.630 ;
        RECT 0.140 1640.110 2262.060 1640.930 ;
        RECT 0.140 1638.410 2262.720 1640.110 ;
        RECT 1.140 1637.590 2262.060 1638.410 ;
        RECT 0.140 1635.890 2262.720 1637.590 ;
        RECT 0.140 1635.070 2262.060 1635.890 ;
        RECT 0.140 1633.370 2262.720 1635.070 ;
        RECT 1.140 1632.550 2262.060 1633.370 ;
        RECT 0.140 1630.850 2262.720 1632.550 ;
        RECT 0.140 1630.030 2262.060 1630.850 ;
        RECT 0.140 1628.330 2262.720 1630.030 ;
        RECT 1.070 1627.510 2262.060 1628.330 ;
        RECT 0.140 1625.810 2262.720 1627.510 ;
        RECT 0.140 1624.990 2262.060 1625.810 ;
        RECT 0.140 1623.290 2262.720 1624.990 ;
        RECT 1.140 1622.470 2262.060 1623.290 ;
        RECT 0.140 1620.770 2262.720 1622.470 ;
        RECT 0.140 1619.950 2262.130 1620.770 ;
        RECT 0.140 1618.250 2262.720 1619.950 ;
        RECT 1.070 1617.430 2262.060 1618.250 ;
        RECT 0.140 1615.730 2262.720 1617.430 ;
        RECT 0.140 1614.910 2262.060 1615.730 ;
        RECT 0.140 1613.210 2262.720 1614.910 ;
        RECT 1.070 1612.390 2262.060 1613.210 ;
        RECT 0.140 1610.690 2262.720 1612.390 ;
        RECT 0.140 1609.870 2262.060 1610.690 ;
        RECT 0.140 1608.170 2262.720 1609.870 ;
        RECT 1.070 1607.350 2262.060 1608.170 ;
        RECT 0.140 1605.650 2262.720 1607.350 ;
        RECT 0.140 1604.830 2262.060 1605.650 ;
        RECT 0.140 1603.130 2262.720 1604.830 ;
        RECT 1.070 1602.310 2262.060 1603.130 ;
        RECT 0.140 1600.610 2262.720 1602.310 ;
        RECT 0.140 1599.790 2262.060 1600.610 ;
        RECT 0.140 1598.090 2262.720 1599.790 ;
        RECT 1.070 1597.270 2262.060 1598.090 ;
        RECT 0.140 1595.570 2262.720 1597.270 ;
        RECT 0.140 1594.750 2262.060 1595.570 ;
        RECT 0.140 1593.050 2262.720 1594.750 ;
        RECT 1.140 1592.230 2262.060 1593.050 ;
        RECT 0.140 1590.530 2262.720 1592.230 ;
        RECT 0.140 1589.710 2262.060 1590.530 ;
        RECT 0.140 1588.010 2262.720 1589.710 ;
        RECT 1.140 1587.190 2262.060 1588.010 ;
        RECT 0.140 1585.490 2262.720 1587.190 ;
        RECT 0.140 1584.670 2262.060 1585.490 ;
        RECT 0.140 1582.970 2262.720 1584.670 ;
        RECT 1.070 1582.150 2262.060 1582.970 ;
        RECT 0.140 1580.450 2262.720 1582.150 ;
        RECT 0.140 1579.630 2262.060 1580.450 ;
        RECT 0.140 1577.930 2262.720 1579.630 ;
        RECT 1.140 1577.110 2262.060 1577.930 ;
        RECT 0.140 1575.410 2262.720 1577.110 ;
        RECT 0.140 1574.590 2262.060 1575.410 ;
        RECT 0.140 1572.890 2262.720 1574.590 ;
        RECT 1.140 1572.070 2262.060 1572.890 ;
        RECT 0.140 1570.370 2262.720 1572.070 ;
        RECT 0.140 1569.550 2262.060 1570.370 ;
        RECT 0.140 1567.850 2262.720 1569.550 ;
        RECT 1.140 1567.030 2262.060 1567.850 ;
        RECT 0.140 1565.330 2262.720 1567.030 ;
        RECT 0.140 1564.510 2262.060 1565.330 ;
        RECT 0.140 1562.810 2262.720 1564.510 ;
        RECT 1.070 1561.990 2262.060 1562.810 ;
        RECT 0.140 1560.290 2262.720 1561.990 ;
        RECT 0.140 1559.470 2262.060 1560.290 ;
        RECT 0.140 1557.770 2262.720 1559.470 ;
        RECT 1.140 1556.950 2262.060 1557.770 ;
        RECT 0.140 1555.250 2262.720 1556.950 ;
        RECT 0.140 1554.430 2262.060 1555.250 ;
        RECT 0.140 1552.730 2262.720 1554.430 ;
        RECT 1.140 1551.910 2262.060 1552.730 ;
        RECT 0.140 1550.210 2262.720 1551.910 ;
        RECT 0.140 1549.390 2262.060 1550.210 ;
        RECT 0.140 1547.690 2262.720 1549.390 ;
        RECT 1.140 1546.870 2262.060 1547.690 ;
        RECT 0.140 1545.170 2262.720 1546.870 ;
        RECT 0.140 1544.350 2262.060 1545.170 ;
        RECT 0.140 1542.650 2262.720 1544.350 ;
        RECT 1.140 1541.830 2262.060 1542.650 ;
        RECT 0.140 1540.130 2262.720 1541.830 ;
        RECT 0.140 1539.310 2262.060 1540.130 ;
        RECT 0.140 1537.610 2262.720 1539.310 ;
        RECT 1.140 1536.790 2262.060 1537.610 ;
        RECT 0.140 1535.090 2262.720 1536.790 ;
        RECT 0.140 1534.270 2262.060 1535.090 ;
        RECT 0.140 1532.570 2262.720 1534.270 ;
        RECT 1.070 1531.750 2262.720 1532.570 ;
        RECT 0.140 1527.530 2262.720 1531.750 ;
        RECT 1.140 1526.710 2262.720 1527.530 ;
        RECT 0.140 1522.490 2262.720 1526.710 ;
        RECT 1.070 1521.670 2262.720 1522.490 ;
        RECT 0.140 1507.370 2262.720 1521.670 ;
        RECT 1.140 1506.550 2262.720 1507.370 ;
        RECT 0.140 1502.330 2262.720 1506.550 ;
        RECT 1.140 1501.510 2262.720 1502.330 ;
        RECT 0.140 1497.290 2262.720 1501.510 ;
        RECT 1.070 1496.470 2262.720 1497.290 ;
        RECT 0.140 1492.250 2262.720 1496.470 ;
        RECT 1.070 1491.430 2262.720 1492.250 ;
        RECT 0.140 1487.210 2262.720 1491.430 ;
        RECT 1.140 1486.390 2262.720 1487.210 ;
        RECT 0.140 1482.170 2262.720 1486.390 ;
        RECT 1.070 1481.350 2262.720 1482.170 ;
        RECT 0.140 1477.130 2262.720 1481.350 ;
        RECT 1.070 1476.310 2262.720 1477.130 ;
        RECT 0.140 1472.090 2262.720 1476.310 ;
        RECT 1.140 1471.270 2262.720 1472.090 ;
        RECT 0.140 1467.050 2262.720 1471.270 ;
        RECT 1.070 1466.230 2262.720 1467.050 ;
        RECT 0.140 1462.010 2262.720 1466.230 ;
        RECT 1.070 1461.190 2262.720 1462.010 ;
        RECT 0.140 1456.970 2262.720 1461.190 ;
        RECT 1.140 1456.150 2262.720 1456.970 ;
        RECT 0.140 1451.930 2262.720 1456.150 ;
        RECT 1.070 1451.110 2262.720 1451.930 ;
        RECT 0.140 1446.890 2262.720 1451.110 ;
        RECT 1.070 1446.070 2262.720 1446.890 ;
        RECT 0.140 1441.850 2262.720 1446.070 ;
        RECT 1.140 1441.030 2262.720 1441.850 ;
        RECT 0.140 1436.810 2262.720 1441.030 ;
        RECT 1.070 1435.990 2262.720 1436.810 ;
        RECT 0.140 1431.770 2262.720 1435.990 ;
        RECT 1.070 1430.950 2262.720 1431.770 ;
        RECT 0.140 1426.730 2262.720 1430.950 ;
        RECT 1.140 1425.910 2262.720 1426.730 ;
        RECT 0.140 1421.690 2262.720 1425.910 ;
        RECT 1.070 1420.870 2262.720 1421.690 ;
        RECT 0.140 1416.650 2262.720 1420.870 ;
        RECT 1.070 1415.830 2262.720 1416.650 ;
        RECT 0.140 1411.610 2262.720 1415.830 ;
        RECT 1.140 1410.790 2262.720 1411.610 ;
        RECT 0.140 1406.570 2262.720 1410.790 ;
        RECT 1.140 1405.750 2262.720 1406.570 ;
        RECT 0.140 1401.530 2262.720 1405.750 ;
        RECT 1.140 1400.710 2262.720 1401.530 ;
        RECT 0.140 1396.490 2262.720 1400.710 ;
        RECT 1.140 1395.670 2262.720 1396.490 ;
        RECT 0.140 1391.450 2262.720 1395.670 ;
        RECT 1.140 1390.630 2262.720 1391.450 ;
        RECT 0.140 1386.410 2262.720 1390.630 ;
        RECT 1.070 1385.590 2262.720 1386.410 ;
        RECT 0.140 1381.370 2262.720 1385.590 ;
        RECT 1.140 1380.550 2262.720 1381.370 ;
        RECT 0.140 1376.330 2262.720 1380.550 ;
        RECT 1.070 1375.510 2262.720 1376.330 ;
        RECT 0.140 1371.290 2262.720 1375.510 ;
        RECT 1.070 1370.470 2262.720 1371.290 ;
        RECT 0.140 1366.250 2262.720 1370.470 ;
        RECT 1.070 1365.430 2262.720 1366.250 ;
        RECT 0.140 1361.210 2262.720 1365.430 ;
        RECT 1.070 1360.390 2262.720 1361.210 ;
        RECT 0.140 1356.170 2262.720 1360.390 ;
        RECT 1.070 1355.350 2262.720 1356.170 ;
        RECT 0.140 1351.130 2262.720 1355.350 ;
        RECT 1.140 1350.310 2262.720 1351.130 ;
        RECT 0.140 1346.090 2262.720 1350.310 ;
        RECT 1.140 1345.270 2262.720 1346.090 ;
        RECT 0.140 1341.050 2262.720 1345.270 ;
        RECT 1.070 1340.230 2262.720 1341.050 ;
        RECT 0.140 1336.010 2262.720 1340.230 ;
        RECT 1.140 1335.190 2262.720 1336.010 ;
        RECT 0.140 1333.490 2262.720 1335.190 ;
        RECT 0.140 1332.670 2262.060 1333.490 ;
        RECT 0.140 1330.970 2262.720 1332.670 ;
        RECT 1.140 1330.150 2262.060 1330.970 ;
        RECT 0.140 1328.450 2262.720 1330.150 ;
        RECT 0.140 1327.630 2262.060 1328.450 ;
        RECT 0.140 1325.930 2262.720 1327.630 ;
        RECT 1.140 1325.110 2262.060 1325.930 ;
        RECT 0.140 1323.410 2262.720 1325.110 ;
        RECT 0.140 1322.590 2262.060 1323.410 ;
        RECT 0.140 1320.890 2262.720 1322.590 ;
        RECT 1.070 1320.070 2262.060 1320.890 ;
        RECT 0.140 1318.370 2262.720 1320.070 ;
        RECT 0.140 1317.550 2262.060 1318.370 ;
        RECT 0.140 1315.850 2262.720 1317.550 ;
        RECT 1.140 1315.030 2262.060 1315.850 ;
        RECT 0.140 1313.330 2262.720 1315.030 ;
        RECT 0.140 1312.510 2262.060 1313.330 ;
        RECT 0.140 1310.810 2262.720 1312.510 ;
        RECT 1.140 1309.990 2262.060 1310.810 ;
        RECT 0.140 1308.290 2262.720 1309.990 ;
        RECT 0.140 1307.470 2262.060 1308.290 ;
        RECT 0.140 1305.770 2262.720 1307.470 ;
        RECT 1.140 1304.950 2262.060 1305.770 ;
        RECT 0.140 1303.250 2262.720 1304.950 ;
        RECT 0.140 1302.430 2262.060 1303.250 ;
        RECT 0.140 1300.730 2262.720 1302.430 ;
        RECT 1.140 1299.910 2262.060 1300.730 ;
        RECT 0.140 1298.210 2262.720 1299.910 ;
        RECT 0.140 1297.390 2262.060 1298.210 ;
        RECT 0.140 1295.690 2262.720 1297.390 ;
        RECT 1.140 1294.870 2262.060 1295.690 ;
        RECT 0.140 1293.170 2262.720 1294.870 ;
        RECT 0.140 1292.350 2262.060 1293.170 ;
        RECT 0.140 1290.650 2262.720 1292.350 ;
        RECT 1.070 1289.830 2262.060 1290.650 ;
        RECT 0.140 1288.130 2262.720 1289.830 ;
        RECT 0.140 1287.310 2262.060 1288.130 ;
        RECT 0.140 1285.610 2262.720 1287.310 ;
        RECT 1.140 1284.790 2262.060 1285.610 ;
        RECT 0.140 1283.090 2262.720 1284.790 ;
        RECT 0.140 1282.270 2262.060 1283.090 ;
        RECT 0.140 1280.570 2262.720 1282.270 ;
        RECT 1.070 1279.750 2262.060 1280.570 ;
        RECT 0.140 1278.050 2262.720 1279.750 ;
        RECT 0.140 1277.230 2262.060 1278.050 ;
        RECT 0.140 1275.530 2262.720 1277.230 ;
        RECT 0.140 1274.710 2262.060 1275.530 ;
        RECT 0.140 1273.010 2262.720 1274.710 ;
        RECT 0.140 1272.190 2262.060 1273.010 ;
        RECT 0.140 1270.490 2262.720 1272.190 ;
        RECT 0.140 1269.670 2262.060 1270.490 ;
        RECT 0.140 1267.970 2262.720 1269.670 ;
        RECT 0.140 1267.150 2262.060 1267.970 ;
        RECT 0.140 1265.450 2262.720 1267.150 ;
        RECT 1.140 1264.630 2262.060 1265.450 ;
        RECT 0.140 1262.930 2262.720 1264.630 ;
        RECT 0.140 1262.110 2262.060 1262.930 ;
        RECT 0.140 1260.410 2262.720 1262.110 ;
        RECT 1.140 1259.590 2262.060 1260.410 ;
        RECT 0.140 1257.890 2262.720 1259.590 ;
        RECT 0.140 1257.070 2262.060 1257.890 ;
        RECT 0.140 1255.370 2262.720 1257.070 ;
        RECT 1.070 1254.550 2262.060 1255.370 ;
        RECT 0.140 1252.850 2262.720 1254.550 ;
        RECT 0.140 1252.030 2262.060 1252.850 ;
        RECT 0.140 1250.330 2262.720 1252.030 ;
        RECT 1.070 1249.510 2262.060 1250.330 ;
        RECT 0.140 1247.810 2262.720 1249.510 ;
        RECT 0.140 1246.990 2262.060 1247.810 ;
        RECT 0.140 1245.290 2262.720 1246.990 ;
        RECT 1.140 1244.470 2262.060 1245.290 ;
        RECT 0.140 1242.770 2262.720 1244.470 ;
        RECT 0.140 1241.950 2262.060 1242.770 ;
        RECT 0.140 1240.250 2262.720 1241.950 ;
        RECT 1.070 1239.430 2262.060 1240.250 ;
        RECT 0.140 1237.730 2262.720 1239.430 ;
        RECT 0.140 1236.910 2262.060 1237.730 ;
        RECT 0.140 1235.210 2262.720 1236.910 ;
        RECT 1.070 1234.390 2262.060 1235.210 ;
        RECT 0.140 1232.690 2262.720 1234.390 ;
        RECT 0.140 1231.870 2262.060 1232.690 ;
        RECT 0.140 1230.170 2262.720 1231.870 ;
        RECT 1.140 1229.350 2262.060 1230.170 ;
        RECT 0.140 1227.650 2262.720 1229.350 ;
        RECT 0.140 1226.830 2262.060 1227.650 ;
        RECT 0.140 1225.130 2262.720 1226.830 ;
        RECT 1.070 1224.310 2262.060 1225.130 ;
        RECT 0.140 1222.610 2262.720 1224.310 ;
        RECT 0.140 1221.790 2262.060 1222.610 ;
        RECT 0.140 1220.090 2262.720 1221.790 ;
        RECT 1.070 1219.270 2262.060 1220.090 ;
        RECT 0.140 1217.570 2262.720 1219.270 ;
        RECT 0.140 1216.750 2262.060 1217.570 ;
        RECT 0.140 1215.050 2262.720 1216.750 ;
        RECT 1.140 1214.230 2262.060 1215.050 ;
        RECT 0.140 1212.530 2262.720 1214.230 ;
        RECT 0.140 1211.710 2262.060 1212.530 ;
        RECT 0.140 1210.010 2262.720 1211.710 ;
        RECT 1.070 1209.190 2262.060 1210.010 ;
        RECT 0.140 1207.490 2262.720 1209.190 ;
        RECT 0.140 1206.670 2262.060 1207.490 ;
        RECT 0.140 1204.970 2262.720 1206.670 ;
        RECT 1.070 1204.150 2262.060 1204.970 ;
        RECT 0.140 1202.450 2262.720 1204.150 ;
        RECT 0.140 1201.630 2262.060 1202.450 ;
        RECT 0.140 1199.930 2262.720 1201.630 ;
        RECT 1.140 1199.110 2262.060 1199.930 ;
        RECT 0.140 1197.410 2262.720 1199.110 ;
        RECT 0.140 1196.590 2262.060 1197.410 ;
        RECT 0.140 1194.890 2262.720 1196.590 ;
        RECT 1.070 1194.070 2262.060 1194.890 ;
        RECT 0.140 1192.370 2262.720 1194.070 ;
        RECT 0.140 1191.550 2262.060 1192.370 ;
        RECT 0.140 1189.850 2262.720 1191.550 ;
        RECT 1.070 1189.030 2262.060 1189.850 ;
        RECT 0.140 1187.330 2262.720 1189.030 ;
        RECT 0.140 1186.510 2262.060 1187.330 ;
        RECT 0.140 1184.810 2262.720 1186.510 ;
        RECT 1.140 1183.990 2262.060 1184.810 ;
        RECT 0.140 1182.290 2262.720 1183.990 ;
        RECT 0.140 1181.470 2262.060 1182.290 ;
        RECT 0.140 1179.770 2262.720 1181.470 ;
        RECT 1.070 1178.950 2262.060 1179.770 ;
        RECT 0.140 1177.250 2262.720 1178.950 ;
        RECT 0.140 1176.430 2262.060 1177.250 ;
        RECT 0.140 1174.730 2262.720 1176.430 ;
        RECT 1.070 1173.910 2262.060 1174.730 ;
        RECT 0.140 1172.210 2262.720 1173.910 ;
        RECT 0.140 1171.390 2262.060 1172.210 ;
        RECT 0.140 1169.690 2262.720 1171.390 ;
        RECT 1.140 1168.870 2262.060 1169.690 ;
        RECT 0.140 1167.170 2262.720 1168.870 ;
        RECT 0.140 1166.350 2262.060 1167.170 ;
        RECT 0.140 1164.650 2262.720 1166.350 ;
        RECT 1.140 1163.830 2262.060 1164.650 ;
        RECT 0.140 1162.130 2262.720 1163.830 ;
        RECT 0.140 1161.310 2262.060 1162.130 ;
        RECT 0.140 1159.610 2262.720 1161.310 ;
        RECT 1.140 1158.790 2262.060 1159.610 ;
        RECT 0.140 1157.090 2262.720 1158.790 ;
        RECT 0.140 1156.270 2262.060 1157.090 ;
        RECT 0.140 1154.570 2262.720 1156.270 ;
        RECT 1.140 1153.750 2262.060 1154.570 ;
        RECT 0.140 1152.050 2262.720 1153.750 ;
        RECT 0.140 1151.230 2262.060 1152.050 ;
        RECT 0.140 1149.530 2262.720 1151.230 ;
        RECT 1.140 1148.710 2262.060 1149.530 ;
        RECT 0.140 1147.010 2262.720 1148.710 ;
        RECT 0.140 1146.190 2262.060 1147.010 ;
        RECT 0.140 1144.490 2262.720 1146.190 ;
        RECT 1.070 1143.670 2262.060 1144.490 ;
        RECT 0.140 1141.970 2262.720 1143.670 ;
        RECT 0.140 1141.150 2262.060 1141.970 ;
        RECT 0.140 1139.450 2262.720 1141.150 ;
        RECT 1.140 1138.630 2262.060 1139.450 ;
        RECT 0.140 1136.930 2262.720 1138.630 ;
        RECT 0.140 1136.110 2262.130 1136.930 ;
        RECT 0.140 1134.410 2262.720 1136.110 ;
        RECT 1.070 1133.590 2262.060 1134.410 ;
        RECT 0.140 1131.890 2262.720 1133.590 ;
        RECT 0.140 1131.070 2262.060 1131.890 ;
        RECT 0.140 1129.370 2262.720 1131.070 ;
        RECT 1.070 1128.550 2262.060 1129.370 ;
        RECT 0.140 1126.850 2262.720 1128.550 ;
        RECT 0.140 1126.030 2262.060 1126.850 ;
        RECT 0.140 1124.330 2262.720 1126.030 ;
        RECT 1.070 1123.510 2262.060 1124.330 ;
        RECT 0.140 1121.810 2262.720 1123.510 ;
        RECT 0.140 1120.990 2262.060 1121.810 ;
        RECT 0.140 1119.290 2262.720 1120.990 ;
        RECT 1.070 1118.470 2262.060 1119.290 ;
        RECT 0.140 1116.770 2262.720 1118.470 ;
        RECT 0.140 1115.950 2262.060 1116.770 ;
        RECT 0.140 1114.250 2262.720 1115.950 ;
        RECT 1.070 1113.430 2262.060 1114.250 ;
        RECT 0.140 1111.730 2262.720 1113.430 ;
        RECT 0.140 1110.910 2262.060 1111.730 ;
        RECT 0.140 1109.210 2262.720 1110.910 ;
        RECT 1.140 1108.390 2262.060 1109.210 ;
        RECT 0.140 1106.690 2262.720 1108.390 ;
        RECT 0.140 1105.870 2262.060 1106.690 ;
        RECT 0.140 1104.170 2262.720 1105.870 ;
        RECT 1.140 1103.350 2262.060 1104.170 ;
        RECT 0.140 1101.650 2262.720 1103.350 ;
        RECT 0.140 1100.830 2262.060 1101.650 ;
        RECT 0.140 1099.130 2262.720 1100.830 ;
        RECT 1.070 1098.310 2262.060 1099.130 ;
        RECT 0.140 1096.610 2262.720 1098.310 ;
        RECT 0.140 1095.790 2262.060 1096.610 ;
        RECT 0.140 1094.090 2262.720 1095.790 ;
        RECT 1.140 1093.270 2262.060 1094.090 ;
        RECT 0.140 1091.570 2262.720 1093.270 ;
        RECT 0.140 1090.750 2262.060 1091.570 ;
        RECT 0.140 1089.050 2262.720 1090.750 ;
        RECT 1.140 1088.230 2262.060 1089.050 ;
        RECT 0.140 1086.530 2262.720 1088.230 ;
        RECT 0.140 1085.710 2262.060 1086.530 ;
        RECT 0.140 1084.010 2262.720 1085.710 ;
        RECT 1.140 1083.190 2262.060 1084.010 ;
        RECT 0.140 1081.490 2262.720 1083.190 ;
        RECT 0.140 1080.670 2262.060 1081.490 ;
        RECT 0.140 1078.970 2262.720 1080.670 ;
        RECT 1.070 1078.150 2262.060 1078.970 ;
        RECT 0.140 1076.450 2262.720 1078.150 ;
        RECT 0.140 1075.630 2262.060 1076.450 ;
        RECT 0.140 1073.930 2262.720 1075.630 ;
        RECT 1.140 1073.110 2262.060 1073.930 ;
        RECT 0.140 1071.410 2262.720 1073.110 ;
        RECT 0.140 1070.590 2262.060 1071.410 ;
        RECT 0.140 1068.890 2262.720 1070.590 ;
        RECT 1.140 1068.070 2262.060 1068.890 ;
        RECT 0.140 1066.370 2262.720 1068.070 ;
        RECT 0.140 1065.550 2262.060 1066.370 ;
        RECT 0.140 1063.850 2262.720 1065.550 ;
        RECT 1.140 1063.030 2262.060 1063.850 ;
        RECT 0.140 1061.330 2262.720 1063.030 ;
        RECT 0.140 1060.510 2262.060 1061.330 ;
        RECT 0.140 1058.810 2262.720 1060.510 ;
        RECT 1.140 1057.990 2262.060 1058.810 ;
        RECT 0.140 1056.290 2262.720 1057.990 ;
        RECT 0.140 1055.470 2262.060 1056.290 ;
        RECT 0.140 1053.770 2262.720 1055.470 ;
        RECT 1.140 1052.950 2262.060 1053.770 ;
        RECT 0.140 1051.250 2262.720 1052.950 ;
        RECT 0.140 1050.430 2262.060 1051.250 ;
        RECT 0.140 1048.730 2262.720 1050.430 ;
        RECT 1.070 1047.910 2262.720 1048.730 ;
        RECT 0.140 1043.690 2262.720 1047.910 ;
        RECT 1.140 1042.870 2262.720 1043.690 ;
        RECT 0.140 1038.650 2262.720 1042.870 ;
        RECT 1.070 1037.830 2262.720 1038.650 ;
        RECT 0.140 1023.530 2262.720 1037.830 ;
        RECT 1.140 1022.710 2262.720 1023.530 ;
        RECT 0.140 1018.490 2262.720 1022.710 ;
        RECT 1.140 1017.670 2262.720 1018.490 ;
        RECT 0.140 1013.450 2262.720 1017.670 ;
        RECT 1.070 1012.630 2262.720 1013.450 ;
        RECT 0.140 1008.410 2262.720 1012.630 ;
        RECT 1.070 1007.590 2262.720 1008.410 ;
        RECT 0.140 1003.370 2262.720 1007.590 ;
        RECT 1.140 1002.550 2262.720 1003.370 ;
        RECT 0.140 998.330 2262.720 1002.550 ;
        RECT 1.070 997.510 2262.720 998.330 ;
        RECT 0.140 993.290 2262.720 997.510 ;
        RECT 1.070 992.470 2262.720 993.290 ;
        RECT 0.140 988.250 2262.720 992.470 ;
        RECT 1.140 987.430 2262.720 988.250 ;
        RECT 0.140 983.210 2262.720 987.430 ;
        RECT 1.070 982.390 2262.720 983.210 ;
        RECT 0.140 978.170 2262.720 982.390 ;
        RECT 1.070 977.350 2262.720 978.170 ;
        RECT 0.140 973.130 2262.720 977.350 ;
        RECT 1.140 972.310 2262.720 973.130 ;
        RECT 0.140 968.090 2262.720 972.310 ;
        RECT 1.070 967.270 2262.720 968.090 ;
        RECT 0.140 963.050 2262.720 967.270 ;
        RECT 1.070 962.230 2262.720 963.050 ;
        RECT 0.140 958.010 2262.720 962.230 ;
        RECT 1.140 957.190 2262.720 958.010 ;
        RECT 0.140 952.970 2262.720 957.190 ;
        RECT 1.070 952.150 2262.720 952.970 ;
        RECT 0.140 947.930 2262.720 952.150 ;
        RECT 1.070 947.110 2262.720 947.930 ;
        RECT 0.140 942.890 2262.720 947.110 ;
        RECT 1.140 942.070 2262.720 942.890 ;
        RECT 0.140 937.850 2262.720 942.070 ;
        RECT 1.070 937.030 2262.720 937.850 ;
        RECT 0.140 932.810 2262.720 937.030 ;
        RECT 1.070 931.990 2262.720 932.810 ;
        RECT 0.140 927.770 2262.720 931.990 ;
        RECT 1.140 926.950 2262.720 927.770 ;
        RECT 0.140 922.730 2262.720 926.950 ;
        RECT 1.140 921.910 2262.720 922.730 ;
        RECT 0.140 917.690 2262.720 921.910 ;
        RECT 1.140 916.870 2262.720 917.690 ;
        RECT 0.140 912.650 2262.720 916.870 ;
        RECT 1.140 911.830 2262.720 912.650 ;
        RECT 0.140 907.610 2262.720 911.830 ;
        RECT 1.140 906.790 2262.720 907.610 ;
        RECT 0.140 902.570 2262.720 906.790 ;
        RECT 1.070 901.750 2262.720 902.570 ;
        RECT 0.140 897.530 2262.720 901.750 ;
        RECT 1.140 896.710 2262.720 897.530 ;
        RECT 0.140 892.490 2262.720 896.710 ;
        RECT 1.070 891.670 2262.720 892.490 ;
        RECT 0.140 887.450 2262.720 891.670 ;
        RECT 1.070 886.630 2262.720 887.450 ;
        RECT 0.140 882.410 2262.720 886.630 ;
        RECT 1.070 881.590 2262.720 882.410 ;
        RECT 0.140 877.370 2262.720 881.590 ;
        RECT 1.070 876.550 2262.720 877.370 ;
        RECT 0.140 872.330 2262.720 876.550 ;
        RECT 1.070 871.510 2262.720 872.330 ;
        RECT 0.140 867.290 2262.720 871.510 ;
        RECT 1.140 866.470 2262.720 867.290 ;
        RECT 0.140 862.250 2262.720 866.470 ;
        RECT 1.140 861.430 2262.720 862.250 ;
        RECT 0.140 857.210 2262.720 861.430 ;
        RECT 1.070 856.390 2262.720 857.210 ;
        RECT 0.140 852.170 2262.720 856.390 ;
        RECT 1.140 851.350 2262.720 852.170 ;
        RECT 0.140 849.650 2262.720 851.350 ;
        RECT 0.140 848.830 2262.060 849.650 ;
        RECT 0.140 847.130 2262.720 848.830 ;
        RECT 1.140 846.310 2262.060 847.130 ;
        RECT 0.140 844.610 2262.720 846.310 ;
        RECT 0.140 843.790 2262.060 844.610 ;
        RECT 0.140 842.090 2262.720 843.790 ;
        RECT 1.140 841.270 2262.060 842.090 ;
        RECT 0.140 839.570 2262.720 841.270 ;
        RECT 0.140 838.750 2262.060 839.570 ;
        RECT 0.140 837.050 2262.720 838.750 ;
        RECT 1.070 836.230 2262.060 837.050 ;
        RECT 0.140 834.530 2262.720 836.230 ;
        RECT 0.140 833.710 2262.060 834.530 ;
        RECT 0.140 832.010 2262.720 833.710 ;
        RECT 1.140 831.190 2262.060 832.010 ;
        RECT 0.140 829.490 2262.720 831.190 ;
        RECT 0.140 828.670 2262.060 829.490 ;
        RECT 0.140 826.970 2262.720 828.670 ;
        RECT 1.140 826.150 2262.060 826.970 ;
        RECT 0.140 824.450 2262.720 826.150 ;
        RECT 0.140 823.630 2262.060 824.450 ;
        RECT 0.140 821.930 2262.720 823.630 ;
        RECT 1.140 821.110 2262.060 821.930 ;
        RECT 0.140 819.410 2262.720 821.110 ;
        RECT 0.140 818.590 2262.060 819.410 ;
        RECT 0.140 816.890 2262.720 818.590 ;
        RECT 1.140 816.070 2262.060 816.890 ;
        RECT 0.140 814.370 2262.720 816.070 ;
        RECT 0.140 813.550 2262.060 814.370 ;
        RECT 0.140 811.850 2262.720 813.550 ;
        RECT 1.140 811.030 2262.060 811.850 ;
        RECT 0.140 809.330 2262.720 811.030 ;
        RECT 0.140 808.510 2262.060 809.330 ;
        RECT 0.140 806.810 2262.720 808.510 ;
        RECT 1.070 805.990 2262.060 806.810 ;
        RECT 0.140 804.290 2262.720 805.990 ;
        RECT 0.140 803.470 2262.060 804.290 ;
        RECT 0.140 801.770 2262.720 803.470 ;
        RECT 1.140 800.950 2262.060 801.770 ;
        RECT 0.140 799.250 2262.720 800.950 ;
        RECT 0.140 798.430 2262.060 799.250 ;
        RECT 0.140 796.730 2262.720 798.430 ;
        RECT 1.070 795.910 2262.060 796.730 ;
        RECT 0.140 794.210 2262.720 795.910 ;
        RECT 0.140 793.390 2262.060 794.210 ;
        RECT 0.140 791.690 2262.720 793.390 ;
        RECT 0.140 790.870 2262.060 791.690 ;
        RECT 0.140 789.170 2262.720 790.870 ;
        RECT 0.140 788.350 2262.060 789.170 ;
        RECT 0.140 786.650 2262.720 788.350 ;
        RECT 0.140 785.830 2262.060 786.650 ;
        RECT 0.140 784.130 2262.720 785.830 ;
        RECT 0.140 783.310 2262.060 784.130 ;
        RECT 0.140 781.610 2262.720 783.310 ;
        RECT 1.140 780.790 2262.060 781.610 ;
        RECT 0.140 779.090 2262.720 780.790 ;
        RECT 0.140 778.270 2262.060 779.090 ;
        RECT 0.140 776.570 2262.720 778.270 ;
        RECT 1.140 775.750 2262.060 776.570 ;
        RECT 0.140 774.050 2262.720 775.750 ;
        RECT 0.140 773.230 2262.060 774.050 ;
        RECT 0.140 771.530 2262.720 773.230 ;
        RECT 1.070 770.710 2262.060 771.530 ;
        RECT 0.140 769.010 2262.720 770.710 ;
        RECT 0.140 768.190 2262.060 769.010 ;
        RECT 0.140 766.490 2262.720 768.190 ;
        RECT 1.070 765.670 2262.060 766.490 ;
        RECT 0.140 763.970 2262.720 765.670 ;
        RECT 0.140 763.150 2262.060 763.970 ;
        RECT 0.140 761.450 2262.720 763.150 ;
        RECT 1.140 760.630 2262.060 761.450 ;
        RECT 0.140 758.930 2262.720 760.630 ;
        RECT 0.140 758.110 2262.060 758.930 ;
        RECT 0.140 756.410 2262.720 758.110 ;
        RECT 1.070 755.590 2262.060 756.410 ;
        RECT 0.140 753.890 2262.720 755.590 ;
        RECT 0.140 753.070 2262.060 753.890 ;
        RECT 0.140 751.370 2262.720 753.070 ;
        RECT 1.070 750.550 2262.060 751.370 ;
        RECT 0.140 748.850 2262.720 750.550 ;
        RECT 0.140 748.030 2262.060 748.850 ;
        RECT 0.140 746.330 2262.720 748.030 ;
        RECT 1.140 745.510 2262.060 746.330 ;
        RECT 0.140 743.810 2262.720 745.510 ;
        RECT 0.140 742.990 2262.060 743.810 ;
        RECT 0.140 741.290 2262.720 742.990 ;
        RECT 1.070 740.470 2262.060 741.290 ;
        RECT 0.140 738.770 2262.720 740.470 ;
        RECT 0.140 737.950 2262.060 738.770 ;
        RECT 0.140 736.250 2262.720 737.950 ;
        RECT 1.070 735.430 2262.060 736.250 ;
        RECT 0.140 733.730 2262.720 735.430 ;
        RECT 0.140 732.910 2262.060 733.730 ;
        RECT 0.140 731.210 2262.720 732.910 ;
        RECT 1.140 730.390 2262.060 731.210 ;
        RECT 0.140 728.690 2262.720 730.390 ;
        RECT 0.140 727.870 2262.060 728.690 ;
        RECT 0.140 726.170 2262.720 727.870 ;
        RECT 1.070 725.350 2262.060 726.170 ;
        RECT 0.140 723.650 2262.720 725.350 ;
        RECT 0.140 722.830 2262.060 723.650 ;
        RECT 0.140 721.130 2262.720 722.830 ;
        RECT 1.070 720.310 2262.060 721.130 ;
        RECT 0.140 718.610 2262.720 720.310 ;
        RECT 0.140 717.790 2262.060 718.610 ;
        RECT 0.140 716.090 2262.720 717.790 ;
        RECT 1.140 715.270 2262.060 716.090 ;
        RECT 0.140 713.570 2262.720 715.270 ;
        RECT 0.140 712.750 2262.060 713.570 ;
        RECT 0.140 711.050 2262.720 712.750 ;
        RECT 1.070 710.230 2262.060 711.050 ;
        RECT 0.140 708.530 2262.720 710.230 ;
        RECT 0.140 707.710 2262.060 708.530 ;
        RECT 0.140 706.010 2262.720 707.710 ;
        RECT 1.070 705.190 2262.060 706.010 ;
        RECT 0.140 703.490 2262.720 705.190 ;
        RECT 0.140 702.670 2262.060 703.490 ;
        RECT 0.140 700.970 2262.720 702.670 ;
        RECT 1.140 700.150 2262.060 700.970 ;
        RECT 0.140 698.450 2262.720 700.150 ;
        RECT 0.140 697.630 2262.060 698.450 ;
        RECT 0.140 695.930 2262.720 697.630 ;
        RECT 1.070 695.110 2262.060 695.930 ;
        RECT 0.140 693.410 2262.720 695.110 ;
        RECT 0.140 692.590 2262.060 693.410 ;
        RECT 0.140 690.890 2262.720 692.590 ;
        RECT 1.070 690.070 2262.060 690.890 ;
        RECT 0.140 688.370 2262.720 690.070 ;
        RECT 0.140 687.550 2262.060 688.370 ;
        RECT 0.140 685.850 2262.720 687.550 ;
        RECT 1.140 685.030 2262.060 685.850 ;
        RECT 0.140 683.330 2262.720 685.030 ;
        RECT 0.140 682.510 2262.060 683.330 ;
        RECT 0.140 680.810 2262.720 682.510 ;
        RECT 1.140 679.990 2262.060 680.810 ;
        RECT 0.140 678.290 2262.720 679.990 ;
        RECT 0.140 677.470 2262.060 678.290 ;
        RECT 0.140 675.770 2262.720 677.470 ;
        RECT 1.140 674.950 2262.060 675.770 ;
        RECT 0.140 673.250 2262.720 674.950 ;
        RECT 0.140 672.430 2262.060 673.250 ;
        RECT 0.140 670.730 2262.720 672.430 ;
        RECT 1.140 669.910 2262.060 670.730 ;
        RECT 0.140 668.210 2262.720 669.910 ;
        RECT 0.140 667.390 2262.060 668.210 ;
        RECT 0.140 665.690 2262.720 667.390 ;
        RECT 1.140 664.870 2262.060 665.690 ;
        RECT 0.140 663.170 2262.720 664.870 ;
        RECT 0.140 662.350 2262.060 663.170 ;
        RECT 0.140 660.650 2262.720 662.350 ;
        RECT 1.070 659.830 2262.060 660.650 ;
        RECT 0.140 658.130 2262.720 659.830 ;
        RECT 0.140 657.310 2262.060 658.130 ;
        RECT 0.140 655.610 2262.720 657.310 ;
        RECT 1.140 654.790 2262.060 655.610 ;
        RECT 0.140 653.090 2262.720 654.790 ;
        RECT 0.140 652.270 2262.130 653.090 ;
        RECT 0.140 650.570 2262.720 652.270 ;
        RECT 1.070 649.750 2262.060 650.570 ;
        RECT 0.140 648.050 2262.720 649.750 ;
        RECT 0.140 647.230 2262.060 648.050 ;
        RECT 0.140 645.530 2262.720 647.230 ;
        RECT 1.070 644.710 2262.060 645.530 ;
        RECT 0.140 643.010 2262.720 644.710 ;
        RECT 0.140 642.190 2262.060 643.010 ;
        RECT 0.140 640.490 2262.720 642.190 ;
        RECT 1.070 639.670 2262.060 640.490 ;
        RECT 0.140 637.970 2262.720 639.670 ;
        RECT 0.140 637.150 2262.060 637.970 ;
        RECT 0.140 635.450 2262.720 637.150 ;
        RECT 1.070 634.630 2262.060 635.450 ;
        RECT 0.140 632.930 2262.720 634.630 ;
        RECT 0.140 632.110 2262.060 632.930 ;
        RECT 0.140 630.410 2262.720 632.110 ;
        RECT 1.070 629.590 2262.060 630.410 ;
        RECT 0.140 627.890 2262.720 629.590 ;
        RECT 0.140 627.070 2262.060 627.890 ;
        RECT 0.140 625.370 2262.720 627.070 ;
        RECT 1.140 624.550 2262.060 625.370 ;
        RECT 0.140 622.850 2262.720 624.550 ;
        RECT 0.140 622.030 2262.060 622.850 ;
        RECT 0.140 620.330 2262.720 622.030 ;
        RECT 1.140 619.510 2262.060 620.330 ;
        RECT 0.140 617.810 2262.720 619.510 ;
        RECT 0.140 616.990 2262.060 617.810 ;
        RECT 0.140 615.290 2262.720 616.990 ;
        RECT 1.070 614.470 2262.060 615.290 ;
        RECT 0.140 612.770 2262.720 614.470 ;
        RECT 0.140 611.950 2262.060 612.770 ;
        RECT 0.140 610.250 2262.720 611.950 ;
        RECT 1.140 609.430 2262.060 610.250 ;
        RECT 0.140 607.730 2262.720 609.430 ;
        RECT 0.140 606.910 2262.060 607.730 ;
        RECT 0.140 605.210 2262.720 606.910 ;
        RECT 1.140 604.390 2262.060 605.210 ;
        RECT 0.140 602.690 2262.720 604.390 ;
        RECT 0.140 601.870 2262.060 602.690 ;
        RECT 0.140 600.170 2262.720 601.870 ;
        RECT 1.140 599.350 2262.060 600.170 ;
        RECT 0.140 597.650 2262.720 599.350 ;
        RECT 0.140 596.830 2262.060 597.650 ;
        RECT 0.140 595.130 2262.720 596.830 ;
        RECT 1.070 594.310 2262.060 595.130 ;
        RECT 0.140 592.610 2262.720 594.310 ;
        RECT 0.140 591.790 2262.060 592.610 ;
        RECT 0.140 590.090 2262.720 591.790 ;
        RECT 1.140 589.270 2262.060 590.090 ;
        RECT 0.140 587.570 2262.720 589.270 ;
        RECT 0.140 586.750 2262.060 587.570 ;
        RECT 0.140 585.050 2262.720 586.750 ;
        RECT 1.140 584.230 2262.060 585.050 ;
        RECT 0.140 582.530 2262.720 584.230 ;
        RECT 0.140 581.710 2262.060 582.530 ;
        RECT 0.140 580.010 2262.720 581.710 ;
        RECT 1.140 579.190 2262.060 580.010 ;
        RECT 0.140 577.490 2262.720 579.190 ;
        RECT 0.140 576.670 2262.060 577.490 ;
        RECT 0.140 574.970 2262.720 576.670 ;
        RECT 1.140 574.150 2262.060 574.970 ;
        RECT 0.140 572.450 2262.720 574.150 ;
        RECT 0.140 571.630 2262.060 572.450 ;
        RECT 0.140 569.930 2262.720 571.630 ;
        RECT 1.140 569.110 2262.060 569.930 ;
        RECT 0.140 567.410 2262.720 569.110 ;
        RECT 0.140 566.590 2262.060 567.410 ;
        RECT 0.140 564.890 2262.720 566.590 ;
        RECT 1.070 564.070 2262.720 564.890 ;
        RECT 0.140 559.850 2262.720 564.070 ;
        RECT 1.140 559.030 2262.720 559.850 ;
        RECT 0.140 554.810 2262.720 559.030 ;
        RECT 1.070 553.990 2262.720 554.810 ;
        RECT 0.140 539.690 2262.720 553.990 ;
        RECT 1.140 538.870 2262.720 539.690 ;
        RECT 0.140 534.650 2262.720 538.870 ;
        RECT 1.140 533.830 2262.720 534.650 ;
        RECT 0.140 529.610 2262.720 533.830 ;
        RECT 1.070 528.790 2262.720 529.610 ;
        RECT 0.140 524.570 2262.720 528.790 ;
        RECT 1.070 523.750 2262.720 524.570 ;
        RECT 0.140 519.530 2262.720 523.750 ;
        RECT 1.140 518.710 2262.720 519.530 ;
        RECT 0.140 514.490 2262.720 518.710 ;
        RECT 1.070 513.670 2262.720 514.490 ;
        RECT 0.140 509.450 2262.720 513.670 ;
        RECT 1.070 508.630 2262.720 509.450 ;
        RECT 0.140 504.410 2262.720 508.630 ;
        RECT 1.140 503.590 2262.720 504.410 ;
        RECT 0.140 499.370 2262.720 503.590 ;
        RECT 1.070 498.550 2262.720 499.370 ;
        RECT 0.140 494.330 2262.720 498.550 ;
        RECT 1.070 493.510 2262.720 494.330 ;
        RECT 0.140 489.290 2262.720 493.510 ;
        RECT 1.140 488.470 2262.720 489.290 ;
        RECT 0.140 484.250 2262.720 488.470 ;
        RECT 1.070 483.430 2262.720 484.250 ;
        RECT 0.140 479.210 2262.720 483.430 ;
        RECT 1.070 478.390 2262.720 479.210 ;
        RECT 0.140 474.170 2262.720 478.390 ;
        RECT 1.140 473.350 2262.720 474.170 ;
        RECT 0.140 469.130 2262.720 473.350 ;
        RECT 1.070 468.310 2262.720 469.130 ;
        RECT 0.140 464.090 2262.720 468.310 ;
        RECT 1.070 463.270 2262.720 464.090 ;
        RECT 0.140 459.050 2262.720 463.270 ;
        RECT 1.140 458.230 2262.720 459.050 ;
        RECT 0.140 454.010 2262.720 458.230 ;
        RECT 1.070 453.190 2262.720 454.010 ;
        RECT 0.140 448.970 2262.720 453.190 ;
        RECT 1.070 448.150 2262.720 448.970 ;
        RECT 0.140 443.930 2262.720 448.150 ;
        RECT 1.140 443.110 2262.720 443.930 ;
        RECT 0.140 438.890 2262.720 443.110 ;
        RECT 1.140 438.070 2262.720 438.890 ;
        RECT 0.140 433.850 2262.720 438.070 ;
        RECT 1.140 433.030 2262.720 433.850 ;
        RECT 0.140 428.810 2262.720 433.030 ;
        RECT 1.140 427.990 2262.720 428.810 ;
        RECT 0.140 423.770 2262.720 427.990 ;
        RECT 1.140 422.950 2262.720 423.770 ;
        RECT 0.140 418.730 2262.720 422.950 ;
        RECT 1.070 417.910 2262.720 418.730 ;
        RECT 0.140 413.690 2262.720 417.910 ;
        RECT 1.140 412.870 2262.720 413.690 ;
        RECT 0.140 408.650 2262.720 412.870 ;
        RECT 1.070 407.830 2262.720 408.650 ;
        RECT 0.140 403.610 2262.720 407.830 ;
        RECT 1.070 402.790 2262.720 403.610 ;
        RECT 0.140 398.570 2262.720 402.790 ;
        RECT 1.070 397.750 2262.720 398.570 ;
        RECT 0.140 393.530 2262.720 397.750 ;
        RECT 1.070 392.710 2262.720 393.530 ;
        RECT 0.140 388.490 2262.720 392.710 ;
        RECT 1.070 387.670 2262.720 388.490 ;
        RECT 0.140 383.450 2262.720 387.670 ;
        RECT 1.140 382.630 2262.720 383.450 ;
        RECT 0.140 378.410 2262.720 382.630 ;
        RECT 1.140 377.590 2262.720 378.410 ;
        RECT 0.140 373.370 2262.720 377.590 ;
        RECT 1.070 372.550 2262.720 373.370 ;
        RECT 0.140 368.330 2262.720 372.550 ;
        RECT 1.140 367.510 2262.720 368.330 ;
        RECT 0.140 365.810 2262.720 367.510 ;
        RECT 0.140 364.990 2262.060 365.810 ;
        RECT 0.140 363.290 2262.720 364.990 ;
        RECT 1.140 362.470 2262.060 363.290 ;
        RECT 0.140 360.770 2262.720 362.470 ;
        RECT 0.140 359.950 2262.060 360.770 ;
        RECT 0.140 358.250 2262.720 359.950 ;
        RECT 1.140 357.430 2262.060 358.250 ;
        RECT 0.140 355.730 2262.720 357.430 ;
        RECT 0.140 354.910 2262.060 355.730 ;
        RECT 0.140 353.210 2262.720 354.910 ;
        RECT 1.070 352.390 2262.060 353.210 ;
        RECT 0.140 350.690 2262.720 352.390 ;
        RECT 0.140 349.870 2262.060 350.690 ;
        RECT 0.140 348.170 2262.720 349.870 ;
        RECT 1.140 347.350 2262.060 348.170 ;
        RECT 0.140 345.650 2262.720 347.350 ;
        RECT 0.140 344.830 2262.060 345.650 ;
        RECT 0.140 343.130 2262.720 344.830 ;
        RECT 1.140 342.310 2262.060 343.130 ;
        RECT 0.140 340.610 2262.720 342.310 ;
        RECT 0.140 339.790 2262.060 340.610 ;
        RECT 0.140 338.090 2262.720 339.790 ;
        RECT 1.140 337.270 2262.060 338.090 ;
        RECT 0.140 335.570 2262.720 337.270 ;
        RECT 0.140 334.750 2262.060 335.570 ;
        RECT 0.140 333.050 2262.720 334.750 ;
        RECT 1.140 332.230 2262.060 333.050 ;
        RECT 0.140 330.530 2262.720 332.230 ;
        RECT 0.140 329.710 2262.060 330.530 ;
        RECT 0.140 328.010 2262.720 329.710 ;
        RECT 1.140 327.190 2262.060 328.010 ;
        RECT 0.140 325.490 2262.720 327.190 ;
        RECT 0.140 324.670 2262.060 325.490 ;
        RECT 0.140 322.970 2262.720 324.670 ;
        RECT 1.070 322.150 2262.060 322.970 ;
        RECT 0.140 320.450 2262.720 322.150 ;
        RECT 0.140 319.630 2262.060 320.450 ;
        RECT 0.140 317.930 2262.720 319.630 ;
        RECT 1.140 317.110 2262.060 317.930 ;
        RECT 0.140 315.410 2262.720 317.110 ;
        RECT 0.140 314.590 2262.060 315.410 ;
        RECT 0.140 312.890 2262.720 314.590 ;
        RECT 1.070 312.070 2262.060 312.890 ;
        RECT 0.140 310.370 2262.720 312.070 ;
        RECT 0.140 309.550 2262.060 310.370 ;
        RECT 0.140 307.850 2262.720 309.550 ;
        RECT 0.140 307.030 2262.060 307.850 ;
        RECT 0.140 305.330 2262.720 307.030 ;
        RECT 0.140 304.510 2262.060 305.330 ;
        RECT 0.140 302.810 2262.720 304.510 ;
        RECT 0.140 301.990 2262.060 302.810 ;
        RECT 0.140 300.290 2262.720 301.990 ;
        RECT 0.140 299.470 2262.060 300.290 ;
        RECT 0.140 297.770 2262.720 299.470 ;
        RECT 1.140 296.950 2262.060 297.770 ;
        RECT 0.140 295.250 2262.720 296.950 ;
        RECT 0.140 294.430 2262.060 295.250 ;
        RECT 0.140 292.730 2262.720 294.430 ;
        RECT 1.140 291.910 2262.060 292.730 ;
        RECT 0.140 290.210 2262.720 291.910 ;
        RECT 0.140 289.390 2262.060 290.210 ;
        RECT 0.140 287.690 2262.720 289.390 ;
        RECT 1.070 286.870 2262.060 287.690 ;
        RECT 0.140 285.170 2262.720 286.870 ;
        RECT 0.140 284.350 2262.060 285.170 ;
        RECT 0.140 282.650 2262.720 284.350 ;
        RECT 1.070 281.830 2262.060 282.650 ;
        RECT 0.140 280.130 2262.720 281.830 ;
        RECT 0.140 279.310 2262.060 280.130 ;
        RECT 0.140 277.610 2262.720 279.310 ;
        RECT 1.140 276.790 2262.060 277.610 ;
        RECT 0.140 275.090 2262.720 276.790 ;
        RECT 0.140 274.270 2262.060 275.090 ;
        RECT 0.140 272.570 2262.720 274.270 ;
        RECT 1.070 271.750 2262.060 272.570 ;
        RECT 0.140 270.050 2262.720 271.750 ;
        RECT 0.140 269.230 2262.060 270.050 ;
        RECT 0.140 267.530 2262.720 269.230 ;
        RECT 1.070 266.710 2262.060 267.530 ;
        RECT 0.140 265.010 2262.720 266.710 ;
        RECT 0.140 264.190 2262.060 265.010 ;
        RECT 0.140 262.490 2262.720 264.190 ;
        RECT 1.140 261.670 2262.060 262.490 ;
        RECT 0.140 259.970 2262.720 261.670 ;
        RECT 0.140 259.150 2262.060 259.970 ;
        RECT 0.140 257.450 2262.720 259.150 ;
        RECT 1.070 256.630 2262.060 257.450 ;
        RECT 0.140 254.930 2262.720 256.630 ;
        RECT 0.140 254.110 2262.060 254.930 ;
        RECT 0.140 252.410 2262.720 254.110 ;
        RECT 1.070 251.590 2262.060 252.410 ;
        RECT 0.140 249.890 2262.720 251.590 ;
        RECT 0.140 249.070 2262.060 249.890 ;
        RECT 0.140 247.370 2262.720 249.070 ;
        RECT 1.140 246.550 2262.060 247.370 ;
        RECT 0.140 244.850 2262.720 246.550 ;
        RECT 0.140 244.030 2262.060 244.850 ;
        RECT 0.140 242.330 2262.720 244.030 ;
        RECT 1.070 241.510 2262.060 242.330 ;
        RECT 0.140 239.810 2262.720 241.510 ;
        RECT 0.140 238.990 2262.060 239.810 ;
        RECT 0.140 237.290 2262.720 238.990 ;
        RECT 1.070 236.470 2262.060 237.290 ;
        RECT 0.140 234.770 2262.720 236.470 ;
        RECT 0.140 233.950 2262.060 234.770 ;
        RECT 0.140 232.250 2262.720 233.950 ;
        RECT 1.140 231.430 2262.060 232.250 ;
        RECT 0.140 229.730 2262.720 231.430 ;
        RECT 0.140 228.910 2262.060 229.730 ;
        RECT 0.140 227.210 2262.720 228.910 ;
        RECT 1.070 226.390 2262.060 227.210 ;
        RECT 0.140 224.690 2262.720 226.390 ;
        RECT 0.140 223.870 2262.060 224.690 ;
        RECT 0.140 222.170 2262.720 223.870 ;
        RECT 1.070 221.350 2262.060 222.170 ;
        RECT 0.140 219.650 2262.720 221.350 ;
        RECT 0.140 218.830 2262.060 219.650 ;
        RECT 0.140 217.130 2262.720 218.830 ;
        RECT 1.140 216.310 2262.060 217.130 ;
        RECT 0.140 214.610 2262.720 216.310 ;
        RECT 0.140 213.790 2262.060 214.610 ;
        RECT 0.140 212.090 2262.720 213.790 ;
        RECT 1.070 211.270 2262.060 212.090 ;
        RECT 0.140 209.570 2262.720 211.270 ;
        RECT 0.140 208.750 2262.060 209.570 ;
        RECT 0.140 207.050 2262.720 208.750 ;
        RECT 1.070 206.230 2262.060 207.050 ;
        RECT 0.140 204.530 2262.720 206.230 ;
        RECT 0.140 203.710 2262.060 204.530 ;
        RECT 0.140 202.010 2262.720 203.710 ;
        RECT 1.140 201.190 2262.060 202.010 ;
        RECT 0.140 199.490 2262.720 201.190 ;
        RECT 0.140 198.670 2262.060 199.490 ;
        RECT 0.140 196.970 2262.720 198.670 ;
        RECT 1.140 196.150 2262.060 196.970 ;
        RECT 0.140 194.450 2262.720 196.150 ;
        RECT 0.140 193.630 2262.060 194.450 ;
        RECT 0.140 191.930 2262.720 193.630 ;
        RECT 1.140 191.110 2262.060 191.930 ;
        RECT 0.140 189.410 2262.720 191.110 ;
        RECT 0.140 188.590 2262.060 189.410 ;
        RECT 0.140 186.890 2262.720 188.590 ;
        RECT 1.140 186.070 2262.060 186.890 ;
        RECT 0.140 184.370 2262.720 186.070 ;
        RECT 0.140 183.550 2262.060 184.370 ;
        RECT 0.140 181.850 2262.720 183.550 ;
        RECT 1.140 181.030 2262.060 181.850 ;
        RECT 0.140 179.330 2262.720 181.030 ;
        RECT 0.140 178.510 2262.060 179.330 ;
        RECT 0.140 176.810 2262.720 178.510 ;
        RECT 1.070 175.990 2262.060 176.810 ;
        RECT 0.140 174.290 2262.720 175.990 ;
        RECT 0.140 173.470 2262.060 174.290 ;
        RECT 0.140 171.770 2262.720 173.470 ;
        RECT 1.140 170.950 2262.060 171.770 ;
        RECT 0.140 169.250 2262.720 170.950 ;
        RECT 0.140 168.430 2262.130 169.250 ;
        RECT 0.140 166.730 2262.720 168.430 ;
        RECT 1.070 165.910 2262.060 166.730 ;
        RECT 0.140 164.210 2262.720 165.910 ;
        RECT 0.140 163.390 2262.060 164.210 ;
        RECT 0.140 161.690 2262.720 163.390 ;
        RECT 1.070 160.870 2262.060 161.690 ;
        RECT 0.140 159.170 2262.720 160.870 ;
        RECT 0.140 158.350 2262.060 159.170 ;
        RECT 0.140 156.650 2262.720 158.350 ;
        RECT 1.070 155.830 2262.060 156.650 ;
        RECT 0.140 154.130 2262.720 155.830 ;
        RECT 0.140 153.310 2262.060 154.130 ;
        RECT 0.140 151.610 2262.720 153.310 ;
        RECT 1.070 150.790 2262.060 151.610 ;
        RECT 0.140 149.090 2262.720 150.790 ;
        RECT 0.140 148.270 2262.060 149.090 ;
        RECT 0.140 146.570 2262.720 148.270 ;
        RECT 1.070 145.750 2262.060 146.570 ;
        RECT 0.140 144.050 2262.720 145.750 ;
        RECT 0.140 143.230 2262.060 144.050 ;
        RECT 0.140 141.530 2262.720 143.230 ;
        RECT 1.140 140.710 2262.060 141.530 ;
        RECT 0.140 139.010 2262.720 140.710 ;
        RECT 0.140 138.190 2262.060 139.010 ;
        RECT 0.140 136.490 2262.720 138.190 ;
        RECT 1.140 135.670 2262.060 136.490 ;
        RECT 0.140 133.970 2262.720 135.670 ;
        RECT 0.140 133.150 2262.060 133.970 ;
        RECT 0.140 131.450 2262.720 133.150 ;
        RECT 1.070 130.630 2262.060 131.450 ;
        RECT 0.140 128.930 2262.720 130.630 ;
        RECT 0.140 128.110 2262.060 128.930 ;
        RECT 0.140 126.410 2262.720 128.110 ;
        RECT 1.140 125.590 2262.060 126.410 ;
        RECT 0.140 123.890 2262.720 125.590 ;
        RECT 0.140 123.070 2262.060 123.890 ;
        RECT 0.140 121.370 2262.720 123.070 ;
        RECT 1.140 120.550 2262.060 121.370 ;
        RECT 0.140 118.850 2262.720 120.550 ;
        RECT 0.140 118.030 2262.060 118.850 ;
        RECT 0.140 116.330 2262.720 118.030 ;
        RECT 1.140 115.510 2262.060 116.330 ;
        RECT 0.140 113.810 2262.720 115.510 ;
        RECT 0.140 112.990 2262.060 113.810 ;
        RECT 0.140 111.290 2262.720 112.990 ;
        RECT 1.070 110.470 2262.060 111.290 ;
        RECT 0.140 108.770 2262.720 110.470 ;
        RECT 0.140 107.950 2262.060 108.770 ;
        RECT 0.140 106.250 2262.720 107.950 ;
        RECT 1.140 105.430 2262.060 106.250 ;
        RECT 0.140 103.730 2262.720 105.430 ;
        RECT 0.140 102.910 2262.060 103.730 ;
        RECT 0.140 101.210 2262.720 102.910 ;
        RECT 1.140 100.390 2262.060 101.210 ;
        RECT 0.140 98.690 2262.720 100.390 ;
        RECT 0.140 97.870 2262.060 98.690 ;
        RECT 0.140 96.170 2262.720 97.870 ;
        RECT 1.140 95.350 2262.060 96.170 ;
        RECT 0.140 93.650 2262.720 95.350 ;
        RECT 0.140 92.830 2262.060 93.650 ;
        RECT 0.140 91.130 2262.720 92.830 ;
        RECT 1.140 90.310 2262.060 91.130 ;
        RECT 0.140 88.610 2262.720 90.310 ;
        RECT 0.140 87.790 2262.060 88.610 ;
        RECT 0.140 86.090 2262.720 87.790 ;
        RECT 1.140 85.270 2262.060 86.090 ;
        RECT 0.140 83.570 2262.720 85.270 ;
        RECT 0.140 82.750 2262.060 83.570 ;
        RECT 0.140 81.050 2262.720 82.750 ;
        RECT 1.070 80.230 2262.720 81.050 ;
        RECT 0.140 76.010 2262.720 80.230 ;
        RECT 1.140 75.190 2262.720 76.010 ;
        RECT 0.140 66.770 2262.720 75.190 ;
        RECT 0.690 65.950 2262.720 66.770 ;
        RECT 0.140 59.630 2262.720 65.950 ;
        RECT 0.690 58.810 2262.720 59.630 ;
        RECT 0.140 57.950 2262.720 58.810 ;
        RECT 0.690 57.130 2262.720 57.950 ;
        RECT 0.140 56.270 2262.720 57.130 ;
        RECT 0.690 55.450 2262.720 56.270 ;
        RECT 0.140 54.590 2262.720 55.450 ;
        RECT 0.690 53.770 2262.720 54.590 ;
        RECT 0.140 52.910 2262.720 53.770 ;
        RECT 0.690 52.090 2262.720 52.910 ;
        RECT 0.140 51.230 2262.720 52.090 ;
        RECT 0.690 50.410 2262.720 51.230 ;
        RECT 0.140 49.550 2262.720 50.410 ;
        RECT 0.690 48.730 2262.720 49.550 ;
        RECT 0.140 47.870 2262.720 48.730 ;
        RECT 0.690 47.050 2262.720 47.870 ;
        RECT 0.140 46.190 2262.720 47.050 ;
        RECT 0.690 45.370 2262.720 46.190 ;
        RECT 0.140 44.510 2262.720 45.370 ;
        RECT 0.690 43.690 2262.720 44.510 ;
        RECT 0.140 42.830 2262.720 43.690 ;
        RECT 0.690 42.010 2262.720 42.830 ;
        RECT 0.140 41.150 2262.720 42.010 ;
        RECT 0.690 40.330 2262.720 41.150 ;
        RECT 0.140 39.470 2262.720 40.330 ;
        RECT 0.690 38.650 2262.720 39.470 ;
        RECT 0.140 37.790 2262.720 38.650 ;
        RECT 0.690 36.970 2262.720 37.790 ;
        RECT 0.140 36.110 2262.720 36.970 ;
        RECT 0.690 35.290 2262.720 36.110 ;
        RECT 0.140 34.430 2262.720 35.290 ;
        RECT 0.690 33.610 2262.720 34.430 ;
        RECT 0.140 32.750 2262.720 33.610 ;
        RECT 0.690 31.930 2262.720 32.750 ;
        RECT 0.140 31.070 2262.720 31.930 ;
        RECT 0.690 30.250 2262.720 31.070 ;
        RECT 0.140 29.390 2262.720 30.250 ;
        RECT 0.690 28.570 2262.720 29.390 ;
        RECT 0.140 27.710 2262.720 28.570 ;
        RECT 0.690 26.890 2262.720 27.710 ;
        RECT 0.140 26.030 2262.720 26.890 ;
        RECT 0.690 25.210 2262.720 26.030 ;
        RECT 0.140 24.350 2262.720 25.210 ;
        RECT 0.690 23.530 2262.720 24.350 ;
        RECT 0.140 22.670 2262.720 23.530 ;
        RECT 0.690 21.850 2262.720 22.670 ;
        RECT 0.140 20.990 2262.720 21.850 ;
        RECT 0.690 20.170 2262.720 20.990 ;
        RECT 0.140 19.310 2262.720 20.170 ;
        RECT 0.690 18.490 2262.720 19.310 ;
        RECT 0.140 17.630 2262.720 18.490 ;
        RECT 0.690 16.810 2262.720 17.630 ;
        RECT 0.140 15.950 2262.720 16.810 ;
        RECT 0.690 15.130 2262.720 15.950 ;
        RECT 0.140 14.270 2262.720 15.130 ;
        RECT 0.690 13.450 2262.720 14.270 ;
        RECT 0.140 12.590 2262.720 13.450 ;
        RECT 0.690 11.770 2262.720 12.590 ;
        RECT 0.140 10.910 2262.720 11.770 ;
        RECT 0.690 10.090 2262.720 10.910 ;
        RECT 0.140 9.230 2262.720 10.090 ;
        RECT 0.690 8.410 2262.720 9.230 ;
        RECT 0.140 7.550 2262.720 8.410 ;
        RECT 0.690 6.730 2262.720 7.550 ;
        RECT 0.140 4.520 2262.720 6.730 ;
      LAYER Metal3 ;
        RECT 0.860 3510.590 86.470 3511.200 ;
        RECT 87.290 3510.590 92.230 3511.200 ;
        RECT 93.050 3510.590 97.990 3511.200 ;
        RECT 98.810 3510.590 103.750 3511.200 ;
        RECT 104.570 3510.590 109.510 3511.200 ;
        RECT 110.330 3510.590 115.270 3511.200 ;
        RECT 116.090 3510.590 121.030 3511.200 ;
        RECT 121.850 3510.590 126.790 3511.200 ;
        RECT 127.610 3510.590 132.550 3511.200 ;
        RECT 133.370 3510.590 138.310 3511.200 ;
        RECT 139.130 3510.590 144.070 3511.200 ;
        RECT 144.890 3510.590 149.830 3511.200 ;
        RECT 150.650 3510.590 155.590 3511.200 ;
        RECT 156.410 3510.590 161.350 3511.200 ;
        RECT 162.170 3510.590 318.310 3511.200 ;
        RECT 319.130 3510.590 324.070 3511.200 ;
        RECT 324.890 3510.590 329.830 3511.200 ;
        RECT 330.650 3510.590 335.590 3511.200 ;
        RECT 336.410 3510.590 341.350 3511.200 ;
        RECT 342.170 3510.590 347.110 3511.200 ;
        RECT 347.930 3510.590 352.870 3511.200 ;
        RECT 353.690 3510.590 358.630 3511.200 ;
        RECT 359.450 3510.590 364.390 3511.200 ;
        RECT 365.210 3510.590 370.150 3511.200 ;
        RECT 370.970 3510.590 375.910 3511.200 ;
        RECT 376.730 3510.590 381.670 3511.200 ;
        RECT 382.490 3510.590 387.430 3511.200 ;
        RECT 388.250 3510.590 393.190 3511.200 ;
        RECT 394.010 3510.590 2262.340 3511.200 ;
        RECT 0.860 0.690 2262.340 3510.590 ;
        RECT 0.860 0.610 89.350 0.690 ;
        RECT 0.860 0.275 5.350 0.610 ;
        RECT 6.170 0.275 8.230 0.610 ;
        RECT 9.050 0.275 11.110 0.610 ;
        RECT 11.930 0.275 13.990 0.610 ;
        RECT 14.810 0.275 16.870 0.610 ;
        RECT 17.690 0.275 19.750 0.610 ;
        RECT 20.570 0.275 22.630 0.610 ;
        RECT 23.450 0.275 25.510 0.610 ;
        RECT 26.330 0.275 28.390 0.610 ;
        RECT 29.210 0.275 31.270 0.610 ;
        RECT 32.090 0.275 34.150 0.610 ;
        RECT 34.970 0.275 37.030 0.610 ;
        RECT 37.850 0.275 39.910 0.610 ;
        RECT 40.730 0.275 42.790 0.610 ;
        RECT 43.610 0.275 45.670 0.610 ;
        RECT 46.490 0.275 48.550 0.610 ;
        RECT 49.370 0.275 51.430 0.610 ;
        RECT 52.250 0.275 54.310 0.610 ;
        RECT 55.130 0.275 57.190 0.610 ;
        RECT 58.010 0.275 60.070 0.610 ;
        RECT 60.890 0.275 62.950 0.610 ;
        RECT 63.770 0.275 89.350 0.610 ;
        RECT 90.170 0.275 99.910 0.690 ;
        RECT 100.730 0.275 110.470 0.690 ;
        RECT 111.290 0.275 121.030 0.690 ;
        RECT 121.850 0.275 131.590 0.690 ;
        RECT 132.410 0.275 142.150 0.690 ;
        RECT 142.970 0.275 152.710 0.690 ;
        RECT 153.530 0.275 163.270 0.690 ;
        RECT 164.090 0.275 173.830 0.690 ;
        RECT 174.650 0.275 184.390 0.690 ;
        RECT 185.210 0.275 194.950 0.690 ;
        RECT 195.770 0.275 205.510 0.690 ;
        RECT 206.330 0.275 216.070 0.690 ;
        RECT 216.890 0.275 226.630 0.690 ;
        RECT 227.450 0.275 237.190 0.690 ;
        RECT 238.010 0.275 247.750 0.690 ;
        RECT 248.570 0.275 258.310 0.690 ;
        RECT 259.130 0.275 268.870 0.690 ;
        RECT 269.690 0.275 279.430 0.690 ;
        RECT 280.250 0.275 289.990 0.690 ;
        RECT 290.810 0.275 312.550 0.690 ;
        RECT 313.370 0.275 320.230 0.690 ;
        RECT 321.050 0.275 327.910 0.690 ;
        RECT 328.730 0.275 335.590 0.690 ;
        RECT 336.410 0.275 343.270 0.690 ;
        RECT 344.090 0.275 350.950 0.690 ;
        RECT 351.770 0.275 358.630 0.690 ;
        RECT 359.450 0.275 373.990 0.690 ;
        RECT 374.810 0.275 381.670 0.690 ;
        RECT 382.490 0.275 389.350 0.690 ;
        RECT 390.170 0.275 397.030 0.690 ;
        RECT 397.850 0.275 404.710 0.690 ;
        RECT 405.530 0.275 412.390 0.690 ;
        RECT 413.210 0.275 420.070 0.690 ;
        RECT 420.890 0.275 427.750 0.690 ;
        RECT 428.570 0.275 435.430 0.690 ;
        RECT 436.250 0.275 443.110 0.690 ;
        RECT 443.930 0.275 450.790 0.690 ;
        RECT 451.610 0.275 458.470 0.690 ;
        RECT 459.290 0.275 466.150 0.690 ;
        RECT 466.970 0.275 473.830 0.690 ;
        RECT 474.650 0.275 481.510 0.690 ;
        RECT 482.330 0.275 489.190 0.690 ;
        RECT 490.010 0.275 496.870 0.690 ;
        RECT 497.690 0.275 504.550 0.690 ;
        RECT 505.370 0.275 512.230 0.690 ;
        RECT 513.050 0.275 519.910 0.690 ;
        RECT 520.730 0.275 539.590 0.690 ;
        RECT 540.410 0.275 548.230 0.690 ;
        RECT 549.050 0.275 556.870 0.690 ;
        RECT 557.690 0.275 565.510 0.690 ;
        RECT 566.330 0.275 574.150 0.690 ;
        RECT 574.970 0.275 591.430 0.690 ;
        RECT 592.250 0.275 600.070 0.690 ;
        RECT 600.890 0.275 608.710 0.690 ;
        RECT 609.530 0.275 617.350 0.690 ;
        RECT 618.170 0.275 625.990 0.690 ;
        RECT 626.810 0.275 634.630 0.690 ;
        RECT 635.450 0.275 643.270 0.690 ;
        RECT 644.090 0.275 651.910 0.690 ;
        RECT 652.730 0.275 660.550 0.690 ;
        RECT 661.370 0.275 669.190 0.690 ;
        RECT 670.010 0.275 677.830 0.690 ;
        RECT 678.650 0.275 686.470 0.690 ;
        RECT 687.290 0.275 695.110 0.690 ;
        RECT 695.930 0.275 703.750 0.690 ;
        RECT 704.570 0.275 712.390 0.690 ;
        RECT 713.210 0.275 721.030 0.690 ;
        RECT 721.850 0.275 729.670 0.690 ;
        RECT 730.490 0.275 738.310 0.690 ;
        RECT 739.130 0.275 746.950 0.690 ;
        RECT 747.770 0.275 755.590 0.690 ;
        RECT 756.410 0.275 784.870 0.690 ;
        RECT 785.690 0.275 797.350 0.690 ;
        RECT 798.170 0.275 809.830 0.690 ;
        RECT 810.650 0.275 822.310 0.690 ;
        RECT 823.130 0.275 834.790 0.690 ;
        RECT 835.610 0.275 847.270 0.690 ;
        RECT 848.090 0.275 859.750 0.690 ;
        RECT 860.570 0.275 872.230 0.690 ;
        RECT 873.050 0.275 884.710 0.690 ;
        RECT 885.530 0.275 897.190 0.690 ;
        RECT 898.010 0.275 909.670 0.690 ;
        RECT 910.490 0.275 922.150 0.690 ;
        RECT 922.970 0.275 934.630 0.690 ;
        RECT 935.450 0.275 947.110 0.690 ;
        RECT 947.930 0.275 959.590 0.690 ;
        RECT 960.410 0.275 972.070 0.690 ;
        RECT 972.890 0.275 984.550 0.690 ;
        RECT 985.370 0.275 997.030 0.690 ;
        RECT 997.850 0.275 1009.510 0.690 ;
        RECT 1010.330 0.275 1021.990 0.690 ;
        RECT 1022.810 0.275 1046.470 0.690 ;
        RECT 1047.290 0.275 1050.310 0.690 ;
        RECT 1051.130 0.275 1054.150 0.690 ;
        RECT 1054.970 0.275 1057.990 0.690 ;
        RECT 1058.810 0.275 1061.830 0.690 ;
        RECT 1062.650 0.275 1065.670 0.690 ;
        RECT 1066.490 0.275 1069.510 0.690 ;
        RECT 1070.330 0.275 1073.350 0.690 ;
        RECT 1074.170 0.275 1077.190 0.690 ;
        RECT 1078.010 0.275 1081.030 0.690 ;
        RECT 1081.850 0.275 1084.870 0.690 ;
        RECT 1085.690 0.275 1088.710 0.690 ;
        RECT 1089.530 0.275 1092.550 0.690 ;
        RECT 1093.370 0.275 1096.390 0.690 ;
        RECT 1097.210 0.275 1100.230 0.690 ;
        RECT 1101.050 0.275 1104.070 0.690 ;
        RECT 1104.890 0.275 1107.910 0.690 ;
        RECT 1108.730 0.275 1111.750 0.690 ;
        RECT 1112.570 0.275 1115.590 0.690 ;
        RECT 1116.410 0.275 1119.430 0.690 ;
        RECT 1120.250 0.275 1123.270 0.690 ;
        RECT 1124.090 0.275 1127.110 0.690 ;
        RECT 1127.930 0.275 1130.950 0.690 ;
        RECT 1131.770 0.275 1134.790 0.690 ;
        RECT 1135.610 0.275 1138.630 0.690 ;
        RECT 1139.450 0.275 1142.470 0.690 ;
        RECT 1143.290 0.275 1146.310 0.690 ;
        RECT 1147.130 0.275 1150.150 0.690 ;
        RECT 1150.970 0.275 1153.990 0.690 ;
        RECT 1154.810 0.275 1157.830 0.690 ;
        RECT 1158.650 0.275 1161.670 0.690 ;
        RECT 1162.490 0.275 1165.510 0.690 ;
        RECT 1166.330 0.275 1173.190 0.690 ;
        RECT 1174.010 0.275 1177.030 0.690 ;
        RECT 1177.850 0.275 1180.870 0.690 ;
        RECT 1181.690 0.275 1184.710 0.690 ;
        RECT 1185.530 0.275 1188.550 0.690 ;
        RECT 1189.370 0.275 1192.390 0.690 ;
        RECT 1193.210 0.275 1196.230 0.690 ;
        RECT 1197.050 0.275 1200.070 0.690 ;
        RECT 1200.890 0.275 1203.910 0.690 ;
        RECT 1204.730 0.275 1207.750 0.690 ;
        RECT 1208.570 0.275 1211.590 0.690 ;
        RECT 1212.410 0.275 1215.430 0.690 ;
        RECT 1216.250 0.275 1219.270 0.690 ;
        RECT 1220.090 0.275 1223.110 0.690 ;
        RECT 1223.930 0.275 1226.950 0.690 ;
        RECT 1227.770 0.275 1230.790 0.690 ;
        RECT 1231.610 0.275 1234.630 0.690 ;
        RECT 1235.450 0.275 1238.470 0.690 ;
        RECT 1239.290 0.275 1242.310 0.690 ;
        RECT 1243.130 0.275 1246.150 0.690 ;
        RECT 1246.970 0.275 1278.310 0.690 ;
        RECT 1279.130 0.275 1282.150 0.690 ;
        RECT 1282.970 0.275 1285.990 0.690 ;
        RECT 1286.810 0.275 1289.830 0.690 ;
        RECT 1290.650 0.275 1293.670 0.690 ;
        RECT 1294.490 0.275 1297.510 0.690 ;
        RECT 1298.330 0.275 1301.350 0.690 ;
        RECT 1302.170 0.275 1305.190 0.690 ;
        RECT 1306.010 0.275 1309.030 0.690 ;
        RECT 1309.850 0.275 1312.870 0.690 ;
        RECT 1313.690 0.275 1316.710 0.690 ;
        RECT 1317.530 0.275 1320.550 0.690 ;
        RECT 1321.370 0.275 1324.390 0.690 ;
        RECT 1325.210 0.275 1328.230 0.690 ;
        RECT 1329.050 0.275 1332.070 0.690 ;
        RECT 1332.890 0.275 1335.910 0.690 ;
        RECT 1336.730 0.275 1339.750 0.690 ;
        RECT 1340.570 0.275 1343.590 0.690 ;
        RECT 1344.410 0.275 1347.430 0.690 ;
        RECT 1348.250 0.275 1351.270 0.690 ;
        RECT 1352.090 0.275 1355.110 0.690 ;
        RECT 1355.930 0.275 1358.950 0.690 ;
        RECT 1359.770 0.275 1362.790 0.690 ;
        RECT 1363.610 0.275 1366.630 0.690 ;
        RECT 1367.450 0.275 1370.470 0.690 ;
        RECT 1371.290 0.275 1374.310 0.690 ;
        RECT 1375.130 0.275 1378.150 0.690 ;
        RECT 1378.970 0.275 1381.990 0.690 ;
        RECT 1382.810 0.275 1385.830 0.690 ;
        RECT 1386.650 0.275 1389.670 0.690 ;
        RECT 1390.490 0.275 1393.510 0.690 ;
        RECT 1394.330 0.275 1397.350 0.690 ;
        RECT 1398.170 0.275 1405.030 0.690 ;
        RECT 1405.850 0.275 1408.870 0.690 ;
        RECT 1409.690 0.275 1412.710 0.690 ;
        RECT 1413.530 0.275 1416.550 0.690 ;
        RECT 1417.370 0.275 1420.390 0.690 ;
        RECT 1421.210 0.275 1424.230 0.690 ;
        RECT 1425.050 0.275 1428.070 0.690 ;
        RECT 1428.890 0.275 1431.910 0.690 ;
        RECT 1432.730 0.275 1435.750 0.690 ;
        RECT 1436.570 0.275 1439.590 0.690 ;
        RECT 1440.410 0.275 1443.430 0.690 ;
        RECT 1444.250 0.275 1447.270 0.690 ;
        RECT 1448.090 0.275 1451.110 0.690 ;
        RECT 1451.930 0.275 1454.950 0.690 ;
        RECT 1455.770 0.275 1458.790 0.690 ;
        RECT 1459.610 0.275 1462.630 0.690 ;
        RECT 1463.450 0.275 1466.470 0.690 ;
        RECT 1467.290 0.275 1470.310 0.690 ;
        RECT 1471.130 0.275 1474.150 0.690 ;
        RECT 1474.970 0.275 1477.990 0.690 ;
        RECT 1478.810 0.275 1513.990 0.690 ;
        RECT 1514.810 0.275 1522.630 0.690 ;
        RECT 1523.450 0.275 1531.270 0.690 ;
        RECT 1532.090 0.275 1539.910 0.690 ;
        RECT 1540.730 0.275 1548.550 0.690 ;
        RECT 1549.370 0.275 1557.190 0.690 ;
        RECT 1558.010 0.275 1565.830 0.690 ;
        RECT 1566.650 0.275 1574.470 0.690 ;
        RECT 1575.290 0.275 1583.110 0.690 ;
        RECT 1583.930 0.275 1591.750 0.690 ;
        RECT 1592.570 0.275 1600.390 0.690 ;
        RECT 1601.210 0.275 1609.030 0.690 ;
        RECT 1609.850 0.275 1617.670 0.690 ;
        RECT 1618.490 0.275 1626.310 0.690 ;
        RECT 1627.130 0.275 1634.950 0.690 ;
        RECT 1635.770 0.275 1643.590 0.690 ;
        RECT 1644.410 0.275 1652.230 0.690 ;
        RECT 1653.050 0.275 1660.870 0.690 ;
        RECT 1661.690 0.275 1669.510 0.690 ;
        RECT 1670.330 0.275 1678.150 0.690 ;
        RECT 1678.970 0.275 1706.470 0.690 ;
        RECT 1707.290 0.275 1710.310 0.690 ;
        RECT 1711.130 0.275 1714.150 0.690 ;
        RECT 1714.970 0.275 1717.990 0.690 ;
        RECT 1718.810 0.275 1721.830 0.690 ;
        RECT 1722.650 0.275 1725.670 0.690 ;
        RECT 1726.490 0.275 1729.510 0.690 ;
        RECT 1730.330 0.275 1733.350 0.690 ;
        RECT 1734.170 0.275 1737.190 0.690 ;
        RECT 1738.010 0.275 1741.030 0.690 ;
        RECT 1741.850 0.275 1744.870 0.690 ;
        RECT 1745.690 0.275 1748.710 0.690 ;
        RECT 1749.530 0.275 1752.550 0.690 ;
        RECT 1753.370 0.275 1756.390 0.690 ;
        RECT 1757.210 0.275 1760.230 0.690 ;
        RECT 1761.050 0.275 1764.070 0.690 ;
        RECT 1764.890 0.275 1767.910 0.690 ;
        RECT 1768.730 0.275 1771.750 0.690 ;
        RECT 1772.570 0.275 1775.590 0.690 ;
        RECT 1776.410 0.275 1779.430 0.690 ;
        RECT 1780.250 0.275 1783.270 0.690 ;
        RECT 1784.090 0.275 1787.110 0.690 ;
        RECT 1787.930 0.275 1790.950 0.690 ;
        RECT 1791.770 0.275 1794.790 0.690 ;
        RECT 1795.610 0.275 1798.630 0.690 ;
        RECT 1799.450 0.275 1802.470 0.690 ;
        RECT 1803.290 0.275 1806.310 0.690 ;
        RECT 1807.130 0.275 1810.150 0.690 ;
        RECT 1810.970 0.275 1813.990 0.690 ;
        RECT 1814.810 0.275 1817.830 0.690 ;
        RECT 1818.650 0.275 1821.670 0.690 ;
        RECT 1822.490 0.275 1825.510 0.690 ;
        RECT 1826.330 0.275 1833.190 0.690 ;
        RECT 1834.010 0.275 1837.030 0.690 ;
        RECT 1837.850 0.275 1840.870 0.690 ;
        RECT 1841.690 0.275 1844.710 0.690 ;
        RECT 1845.530 0.275 1848.550 0.690 ;
        RECT 1849.370 0.275 1852.390 0.690 ;
        RECT 1853.210 0.275 1856.230 0.690 ;
        RECT 1857.050 0.275 1860.070 0.690 ;
        RECT 1860.890 0.275 1863.910 0.690 ;
        RECT 1864.730 0.275 1867.750 0.690 ;
        RECT 1868.570 0.275 1871.590 0.690 ;
        RECT 1872.410 0.275 1875.430 0.690 ;
        RECT 1876.250 0.275 1879.270 0.690 ;
        RECT 1880.090 0.275 1883.110 0.690 ;
        RECT 1883.930 0.275 1886.950 0.690 ;
        RECT 1887.770 0.275 1890.790 0.690 ;
        RECT 1891.610 0.275 1894.630 0.690 ;
        RECT 1895.450 0.275 1898.470 0.690 ;
        RECT 1899.290 0.275 1902.310 0.690 ;
        RECT 1903.130 0.275 1906.150 0.690 ;
        RECT 1906.970 0.275 1938.310 0.690 ;
        RECT 1939.130 0.275 1942.150 0.690 ;
        RECT 1942.970 0.275 1945.990 0.690 ;
        RECT 1946.810 0.275 1949.830 0.690 ;
        RECT 1950.650 0.275 1953.670 0.690 ;
        RECT 1954.490 0.275 1957.510 0.690 ;
        RECT 1958.330 0.275 1961.350 0.690 ;
        RECT 1962.170 0.275 1965.190 0.690 ;
        RECT 1966.010 0.275 1969.030 0.690 ;
        RECT 1969.850 0.275 1972.870 0.690 ;
        RECT 1973.690 0.275 1976.710 0.690 ;
        RECT 1977.530 0.275 1980.550 0.690 ;
        RECT 1981.370 0.275 1984.390 0.690 ;
        RECT 1985.210 0.275 1988.230 0.690 ;
        RECT 1989.050 0.275 1992.070 0.690 ;
        RECT 1992.890 0.275 1995.910 0.690 ;
        RECT 1996.730 0.275 1999.750 0.690 ;
        RECT 2000.570 0.275 2003.590 0.690 ;
        RECT 2004.410 0.275 2007.430 0.690 ;
        RECT 2008.250 0.275 2011.270 0.690 ;
        RECT 2012.090 0.275 2015.110 0.690 ;
        RECT 2015.930 0.275 2018.950 0.690 ;
        RECT 2019.770 0.275 2022.790 0.690 ;
        RECT 2023.610 0.275 2026.630 0.690 ;
        RECT 2027.450 0.275 2030.470 0.690 ;
        RECT 2031.290 0.275 2034.310 0.690 ;
        RECT 2035.130 0.275 2038.150 0.690 ;
        RECT 2038.970 0.275 2041.990 0.690 ;
        RECT 2042.810 0.275 2045.830 0.690 ;
        RECT 2046.650 0.275 2049.670 0.690 ;
        RECT 2050.490 0.275 2053.510 0.690 ;
        RECT 2054.330 0.275 2057.350 0.690 ;
        RECT 2058.170 0.275 2065.030 0.690 ;
        RECT 2065.850 0.275 2068.870 0.690 ;
        RECT 2069.690 0.275 2072.710 0.690 ;
        RECT 2073.530 0.275 2076.550 0.690 ;
        RECT 2077.370 0.275 2080.390 0.690 ;
        RECT 2081.210 0.275 2084.230 0.690 ;
        RECT 2085.050 0.275 2088.070 0.690 ;
        RECT 2088.890 0.275 2091.910 0.690 ;
        RECT 2092.730 0.275 2095.750 0.690 ;
        RECT 2096.570 0.275 2099.590 0.690 ;
        RECT 2100.410 0.275 2103.430 0.690 ;
        RECT 2104.250 0.275 2107.270 0.690 ;
        RECT 2108.090 0.275 2111.110 0.690 ;
        RECT 2111.930 0.275 2114.950 0.690 ;
        RECT 2115.770 0.275 2118.790 0.690 ;
        RECT 2119.610 0.275 2122.630 0.690 ;
        RECT 2123.450 0.275 2126.470 0.690 ;
        RECT 2127.290 0.275 2130.310 0.690 ;
        RECT 2131.130 0.275 2134.150 0.690 ;
        RECT 2134.970 0.275 2137.990 0.690 ;
        RECT 2138.810 0.610 2262.340 0.690 ;
        RECT 2138.810 0.275 2164.390 0.610 ;
        RECT 2165.210 0.275 2169.190 0.610 ;
        RECT 2170.010 0.275 2173.990 0.610 ;
        RECT 2174.810 0.275 2178.790 0.610 ;
        RECT 2179.610 0.275 2183.590 0.610 ;
        RECT 2184.410 0.275 2188.390 0.610 ;
        RECT 2189.210 0.275 2193.190 0.610 ;
        RECT 2194.010 0.275 2197.990 0.610 ;
        RECT 2198.810 0.275 2202.790 0.610 ;
        RECT 2203.610 0.275 2207.590 0.610 ;
        RECT 2208.410 0.275 2212.390 0.610 ;
        RECT 2213.210 0.275 2217.190 0.610 ;
        RECT 2218.010 0.275 2221.990 0.610 ;
        RECT 2222.810 0.275 2226.790 0.610 ;
        RECT 2227.610 0.275 2231.590 0.610 ;
        RECT 2232.410 0.275 2236.390 0.610 ;
        RECT 2237.210 0.275 2241.190 0.610 ;
        RECT 2242.010 0.275 2245.990 0.610 ;
        RECT 2246.810 0.275 2250.790 0.610 ;
        RECT 2251.610 0.275 2255.590 0.610 ;
        RECT 2256.410 0.275 2262.340 0.610 ;
      LAYER Metal4 ;
        RECT 5.615 0.320 2262.385 3505.000 ;
      LAYER Metal5 ;
        RECT 7.580 4.200 18.530 3511.200 ;
        RECT 21.150 4.200 24.730 3511.200 ;
        RECT 27.350 4.200 87.170 3511.200 ;
        RECT 89.790 4.200 93.370 3511.200 ;
        RECT 95.990 4.200 162.770 3511.200 ;
        RECT 165.390 4.200 168.970 3511.200 ;
        RECT 171.590 4.200 238.370 3511.200 ;
        RECT 240.990 4.200 244.570 3511.200 ;
        RECT 247.190 4.200 319.010 3511.200 ;
        RECT 321.630 4.200 325.210 3511.200 ;
        RECT 327.830 4.200 394.610 3511.200 ;
        RECT 397.230 4.200 400.810 3511.200 ;
        RECT 403.430 4.200 470.210 3511.200 ;
        RECT 472.830 4.200 476.410 3511.200 ;
        RECT 479.030 4.200 550.850 3511.200 ;
        RECT 553.470 4.200 557.050 3511.200 ;
        RECT 559.670 4.200 626.450 3511.200 ;
        RECT 629.070 4.200 632.650 3511.200 ;
        RECT 635.270 4.200 702.050 3511.200 ;
        RECT 704.670 4.200 708.250 3511.200 ;
        RECT 710.870 4.200 782.690 3511.200 ;
        RECT 785.310 4.200 788.890 3511.200 ;
        RECT 791.510 4.200 858.290 3511.200 ;
        RECT 860.910 4.200 864.490 3511.200 ;
        RECT 867.110 4.200 933.890 3511.200 ;
        RECT 936.510 4.200 940.090 3511.200 ;
        RECT 942.710 4.200 1009.490 3511.200 ;
        RECT 1012.110 4.200 1015.690 3511.200 ;
        RECT 1018.310 4.200 1049.090 3511.200 ;
        RECT 1051.710 4.200 1055.290 3511.200 ;
        RECT 1057.910 4.200 1124.690 3511.200 ;
        RECT 1127.310 4.200 1130.890 3511.200 ;
        RECT 1133.510 4.200 1200.290 3511.200 ;
        RECT 1202.910 4.200 1206.490 3511.200 ;
        RECT 1209.110 4.200 1280.930 3511.200 ;
        RECT 1283.550 4.200 1287.130 3511.200 ;
        RECT 1289.750 4.200 1356.530 3511.200 ;
        RECT 1359.150 4.200 1362.730 3511.200 ;
        RECT 1365.350 4.200 1432.130 3511.200 ;
        RECT 1434.750 4.200 1438.330 3511.200 ;
        RECT 1440.950 4.200 1512.770 3511.200 ;
        RECT 1515.390 4.200 1518.970 3511.200 ;
        RECT 1521.590 4.200 1588.370 3511.200 ;
        RECT 1590.990 4.200 1594.570 3511.200 ;
        RECT 1597.190 4.200 1663.970 3511.200 ;
        RECT 1666.590 4.200 1670.170 3511.200 ;
        RECT 1672.790 4.200 1709.090 3511.200 ;
        RECT 1711.710 4.200 1715.290 3511.200 ;
        RECT 1717.910 4.200 1784.690 3511.200 ;
        RECT 1787.310 4.200 1790.890 3511.200 ;
        RECT 1793.510 4.200 1860.290 3511.200 ;
        RECT 1862.910 4.200 1866.490 3511.200 ;
        RECT 1869.110 4.200 1940.930 3511.200 ;
        RECT 1943.550 4.200 1947.130 3511.200 ;
        RECT 1949.750 4.200 2016.530 3511.200 ;
        RECT 2019.150 4.200 2022.730 3511.200 ;
        RECT 2025.350 4.200 2092.130 3511.200 ;
        RECT 2094.750 4.200 2098.330 3511.200 ;
        RECT 2100.950 4.200 2172.770 3511.200 ;
        RECT 2175.390 4.200 2178.970 3511.200 ;
        RECT 2181.590 4.200 2248.370 3511.200 ;
        RECT 2250.990 4.200 2262.340 3511.200 ;
  END
END eFPGA
END LIBRARY

