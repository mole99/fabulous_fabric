`default_nettype none

module fabric_wrapper #(
    	parameter FrameBitsPerRow = 32,
	parameter MaxFramesPerCol = 20,
	
	parameter NumColumns = 11,
	parameter NumRows = 16,
	
    parameter FABRIC_NUM_IO_WEST = 28,
    parameter FABRIC_NUM_IO_NORTH = 4
)(
    input clk_i,
    
    // Configuration
    input  logic [(FrameBitsPerRow*NumRows)-1:0]    FrameData_i,
    input  logic [(MaxFramesPerCol*NumColumns)-1:0] FrameStrobe_i,
    
    // Fabric is configured
    input                                configured_i,
    
    // I/Os West
    input  [FABRIC_NUM_IO_WEST-1:0]      fabric_io_west_in_i,
    output [FABRIC_NUM_IO_WEST-1:0]      fabric_io_west_out_o,
    output [FABRIC_NUM_IO_WEST-1:0]      fabric_io_west_oe_o,

    // I/O West config
    output [FABRIC_NUM_IO_WEST-1:0]      fabric_io_west_config_bit0_o,
    output [FABRIC_NUM_IO_WEST-1:0]      fabric_io_west_config_bit1_o,
    output [FABRIC_NUM_IO_WEST-1:0]      fabric_io_west_config_bit2_o,
    output [FABRIC_NUM_IO_WEST-1:0]      fabric_io_west_config_bit3_o,

    // I/Os North
    input  [FABRIC_NUM_IO_NORTH-1:0]      fabric_io_north_in_i,
    output [FABRIC_NUM_IO_NORTH-1:0]      fabric_io_north_out_o,
    output [FABRIC_NUM_IO_NORTH-1:0]      fabric_io_north_oe_o,

    // I/O North config
    output [FABRIC_NUM_IO_NORTH-1:0]      fabric_io_north_config_bit0_o,
    output [FABRIC_NUM_IO_NORTH-1:0]      fabric_io_north_config_bit1_o,
    output [FABRIC_NUM_IO_NORTH-1:0]      fabric_io_north_config_bit2_o,
    output [FABRIC_NUM_IO_NORTH-1:0]      fabric_io_north_config_bit3_o,

    // WARMBOOT
    output        fabric_warmboot_boot_o,
    output  [3:0] fabric_warmboot_slot_o,
    input         fabric_warmboot_reset_i,

    // CPU_IRQ
    output  [3:0] fabric_irq_o,

    // CPU_IF - Selector
    input  logic            fabric_xif_or_periph_i,
    
    // Custom instruction interface
    input  logic [31:0]     fabric_rs1_i,
    input  logic [31:0]     fabric_rs2_i,
    output logic [31:0]     fabric_result_o,
    
    // Bus interface
    output logic            fabric_gnt_o,
    input  logic            fabric_req_i,
    output logic            fabric_rvalid_o,
    input  logic            fabric_we_i,
    input  logic [ 3:0]     fabric_be_i,
    input  logic [23:0]     fabric_addr_i,
    input  logic [31:0]     fabric_wdata_i,
    output logic [31:0]     fabric_rdata_o
);
    // SRAM 0
    logic [31:0] fabric_sram0_dout_i;
    logic [9 :0] fabric_sram0_addr_o;
    logic [31:0] fabric_sram0_bm_o;
    logic [31:0] fabric_sram0_din_o;
    logic        fabric_sram0_wen_o;
    logic        fabric_sram0_men_o;
    logic        fabric_sram0_ren_o;
    logic        fabric_sram0_clk_o;
    logic        fabric_sram0_tie_high_o;
    logic        fabric_sram0_tie_low_o;

    // SRAM 1
    logic [31:0] fabric_sram1_dout_i;
    logic [9 :0] fabric_sram1_addr_o;
    logic [31:0] fabric_sram1_bm_o;
    logic [31:0] fabric_sram1_din_o;
    logic        fabric_sram1_wen_o;
    logic        fabric_sram1_men_o;
    logic        fabric_sram1_ren_o;
    logic        fabric_sram1_clk_o;
    logic        fabric_sram1_tie_high_o;
    logic        fabric_sram1_tie_low_o;

    // SRAM 2
    logic [31:0] fabric_sram2_dout_i;
    logic [9 :0] fabric_sram2_addr_o;
    logic [31:0] fabric_sram2_bm_o;
    logic [31:0] fabric_sram2_din_o;
    logic        fabric_sram2_wen_o;
    logic        fabric_sram2_men_o;
    logic        fabric_sram2_ren_o;
    logic        fabric_sram2_clk_o;
    logic        fabric_sram2_tie_high_o;
    logic        fabric_sram2_tie_low_o;

    // SRAM 3
    logic [31:0] fabric_sram3_dout_i;
    logic [9 :0] fabric_sram3_addr_o;
    logic [31:0] fabric_sram3_bm_o;
    logic [31:0] fabric_sram3_din_o;
    logic        fabric_sram3_wen_o;
    logic        fabric_sram3_men_o;
    logic        fabric_sram3_ren_o;
    logic        fabric_sram3_clk_o;
    logic        fabric_sram3_tie_high_o;
    logic        fabric_sram3_tie_low_o;

    // SRAM 4
    logic [31:0] fabric_sram4_dout_i;
    logic [9 :0] fabric_sram4_addr_o;
    logic [31:0] fabric_sram4_bm_o;
    logic [31:0] fabric_sram4_din_o;
    logic        fabric_sram4_wen_o;
    logic        fabric_sram4_men_o;
    logic        fabric_sram4_ren_o;
    logic        fabric_sram4_clk_o;
    logic        fabric_sram4_tie_high_o;
    logic        fabric_sram4_tie_low_o;

    // SRAM 5
    logic [31:0] fabric_sram5_dout_i;
    logic [9 :0] fabric_sram5_addr_o;
    logic [31:0] fabric_sram5_bm_o;
    logic [31:0] fabric_sram5_din_o;
    logic        fabric_sram5_wen_o;
    logic        fabric_sram5_men_o;
    logic        fabric_sram5_ren_o;
    logic        fabric_sram5_clk_o;
    logic        fabric_sram5_tie_high_o;
    logic        fabric_sram5_tie_low_o;

    // SRAM 6
    logic [31:0] fabric_sram6_dout_i;
    logic [9 :0] fabric_sram6_addr_o;
    logic [31:0] fabric_sram6_bm_o;
    logic [31:0] fabric_sram6_din_o;
    logic        fabric_sram6_wen_o;
    logic        fabric_sram6_men_o;
    logic        fabric_sram6_ren_o;
    logic        fabric_sram6_clk_o;
    logic        fabric_sram6_tie_high_o;
    logic        fabric_sram6_tie_low_o;

    // CPU_IF
    logic [63:0] fabric_cpu_i;
    logic [63:0] fabric_cpu_o;
    
    logic fabric_req_d;
    always_ff @(posedge clk_i) begin
        fabric_req_d <= fabric_req_i;
    end
    
    // CPU_IF muxing
    always_comb begin
        // Custom instruction interface selected
        if (fabric_xif_or_periph_i == 1'b0) begin
            // XIF connected to CPU_IF
            fabric_cpu_i    = {fabric_rs2_i, fabric_rs1_i};
            fabric_result_o = fabric_cpu_o[31:0];

            // Default values for peripheral
            fabric_gnt_o    = fabric_req_i;
            fabric_rvalid_o = fabric_req_d;
            fabric_rdata_o  = 32'hDEADBEEF;

        // Bus interface selected
        end else begin
            // Periperhal connected to CPU_IF
            fabric_cpu_i = {2'b0, fabric_req_i, fabric_we_i, fabric_be_i, fabric_addr_i, fabric_wdata_i};

            fabric_gnt_o    = fabric_cpu_o[33];
            fabric_rvalid_o = fabric_cpu_o[32];
            fabric_rdata_o  = fabric_cpu_o[31:0];

            // Default value for XIF
            fabric_result_o = 32'hDEADBEEF;
        end
    end
    
    eFPGA
    //#(
    //    .MaxFramesPerCol(MaxFramesPerCol),
    //    .FrameBitsPerRow(FrameBitsPerRow)
    //)
    eFPGA
    (
        .FrameData      (FrameData_i),
        .FrameStrobe    (FrameStrobe_i),
        .UserCLK        (clk_i),

        // West I/Os
        .Tile_X0Y1_A_O_top(fabric_io_west_in_i[27]),
        .Tile_X0Y1_A_I_top(fabric_io_west_out_o[27]),
        .Tile_X0Y1_A_T_top(fabric_io_west_oe_o[27]),

        .Tile_X0Y1_B_O_top(fabric_io_west_in_i[26]),
        .Tile_X0Y1_B_I_top(fabric_io_west_out_o[26]),
        .Tile_X0Y1_B_T_top(fabric_io_west_oe_o[26]),

        .Tile_X0Y1_A_config_C_bit0(fabric_io_west_config_bit0_o[27]),
        .Tile_X0Y1_A_config_C_bit1(fabric_io_west_config_bit1_o[27]),
        .Tile_X0Y1_A_config_C_bit2(fabric_io_west_config_bit2_o[27]),
        .Tile_X0Y1_A_config_C_bit3(fabric_io_west_config_bit3_o[27]),

        .Tile_X0Y1_B_config_C_bit0(fabric_io_west_config_bit0_o[26]),
        .Tile_X0Y1_B_config_C_bit1(fabric_io_west_config_bit1_o[26]),
        .Tile_X0Y1_B_config_C_bit2(fabric_io_west_config_bit2_o[26]),
        .Tile_X0Y1_B_config_C_bit3(fabric_io_west_config_bit3_o[26]),

        .Tile_X0Y2_A_O_top(fabric_io_west_in_i[25]),
        .Tile_X0Y2_A_I_top(fabric_io_west_out_o[25]),
        .Tile_X0Y2_A_T_top(fabric_io_west_oe_o[25]),

        .Tile_X0Y2_B_O_top(fabric_io_west_in_i[24]),
        .Tile_X0Y2_B_I_top(fabric_io_west_out_o[24]),
        .Tile_X0Y2_B_T_top(fabric_io_west_oe_o[24]),

        .Tile_X0Y2_A_config_C_bit0(fabric_io_west_config_bit0_o[25]),
        .Tile_X0Y2_A_config_C_bit1(fabric_io_west_config_bit1_o[25]),
        .Tile_X0Y2_A_config_C_bit2(fabric_io_west_config_bit2_o[25]),
        .Tile_X0Y2_A_config_C_bit3(fabric_io_west_config_bit3_o[25]),

        .Tile_X0Y2_B_config_C_bit0(fabric_io_west_config_bit0_o[24]),
        .Tile_X0Y2_B_config_C_bit1(fabric_io_west_config_bit1_o[24]),
        .Tile_X0Y2_B_config_C_bit2(fabric_io_west_config_bit2_o[24]),
        .Tile_X0Y2_B_config_C_bit3(fabric_io_west_config_bit3_o[24]),

        .Tile_X0Y3_A_O_top(fabric_io_west_in_i[23]),
        .Tile_X0Y3_A_I_top(fabric_io_west_out_o[23]),
        .Tile_X0Y3_A_T_top(fabric_io_west_oe_o[23]),

        .Tile_X0Y3_B_O_top(fabric_io_west_in_i[22]),
        .Tile_X0Y3_B_I_top(fabric_io_west_out_o[22]),
        .Tile_X0Y3_B_T_top(fabric_io_west_oe_o[22]),

        .Tile_X0Y3_A_config_C_bit0(fabric_io_west_config_bit0_o[23]),
        .Tile_X0Y3_A_config_C_bit1(fabric_io_west_config_bit1_o[23]),
        .Tile_X0Y3_A_config_C_bit2(fabric_io_west_config_bit2_o[23]),
        .Tile_X0Y3_A_config_C_bit3(fabric_io_west_config_bit3_o[23]),

        .Tile_X0Y3_B_config_C_bit0(fabric_io_west_config_bit0_o[22]),
        .Tile_X0Y3_B_config_C_bit1(fabric_io_west_config_bit1_o[22]),
        .Tile_X0Y3_B_config_C_bit2(fabric_io_west_config_bit2_o[22]),
        .Tile_X0Y3_B_config_C_bit3(fabric_io_west_config_bit3_o[22]),

        .Tile_X0Y4_A_O_top(fabric_io_west_in_i[21]),
        .Tile_X0Y4_A_I_top(fabric_io_west_out_o[21]),
        .Tile_X0Y4_A_T_top(fabric_io_west_oe_o[21]),

        .Tile_X0Y4_B_O_top(fabric_io_west_in_i[20]),
        .Tile_X0Y4_B_I_top(fabric_io_west_out_o[20]),
        .Tile_X0Y4_B_T_top(fabric_io_west_oe_o[20]),

        .Tile_X0Y4_A_config_C_bit0(fabric_io_west_config_bit0_o[21]),
        .Tile_X0Y4_A_config_C_bit1(fabric_io_west_config_bit1_o[21]),
        .Tile_X0Y4_A_config_C_bit2(fabric_io_west_config_bit2_o[21]),
        .Tile_X0Y4_A_config_C_bit3(fabric_io_west_config_bit3_o[21]),

        .Tile_X0Y4_B_config_C_bit0(fabric_io_west_config_bit0_o[20]),
        .Tile_X0Y4_B_config_C_bit1(fabric_io_west_config_bit1_o[20]),
        .Tile_X0Y4_B_config_C_bit2(fabric_io_west_config_bit2_o[20]),
        .Tile_X0Y4_B_config_C_bit3(fabric_io_west_config_bit3_o[20]),

        .Tile_X0Y5_A_O_top(fabric_io_west_in_i[19]),
        .Tile_X0Y5_A_I_top(fabric_io_west_out_o[19]),
        .Tile_X0Y5_A_T_top(fabric_io_west_oe_o[19]),

        .Tile_X0Y5_B_O_top(fabric_io_west_in_i[18]),
        .Tile_X0Y5_B_I_top(fabric_io_west_out_o[18]),
        .Tile_X0Y5_B_T_top(fabric_io_west_oe_o[18]),

        .Tile_X0Y5_A_config_C_bit0(fabric_io_west_config_bit0_o[19]),
        .Tile_X0Y5_A_config_C_bit1(fabric_io_west_config_bit1_o[19]),
        .Tile_X0Y5_A_config_C_bit2(fabric_io_west_config_bit2_o[19]),
        .Tile_X0Y5_A_config_C_bit3(fabric_io_west_config_bit3_o[19]),

        .Tile_X0Y5_B_config_C_bit0(fabric_io_west_config_bit0_o[18]),
        .Tile_X0Y5_B_config_C_bit1(fabric_io_west_config_bit1_o[18]),
        .Tile_X0Y5_B_config_C_bit2(fabric_io_west_config_bit2_o[18]),
        .Tile_X0Y5_B_config_C_bit3(fabric_io_west_config_bit3_o[18]),

        .Tile_X0Y6_A_O_top(fabric_io_west_in_i[17]),
        .Tile_X0Y6_A_I_top(fabric_io_west_out_o[17]),
        .Tile_X0Y6_A_T_top(fabric_io_west_oe_o[17]),

        .Tile_X0Y6_B_O_top(fabric_io_west_in_i[16]),
        .Tile_X0Y6_B_I_top(fabric_io_west_out_o[16]),
        .Tile_X0Y6_B_T_top(fabric_io_west_oe_o[16]),

        .Tile_X0Y6_A_config_C_bit0(fabric_io_west_config_bit0_o[17]),
        .Tile_X0Y6_A_config_C_bit1(fabric_io_west_config_bit1_o[17]),
        .Tile_X0Y6_A_config_C_bit2(fabric_io_west_config_bit2_o[17]),
        .Tile_X0Y6_A_config_C_bit3(fabric_io_west_config_bit3_o[17]),

        .Tile_X0Y6_B_config_C_bit0(fabric_io_west_config_bit0_o[16]),
        .Tile_X0Y6_B_config_C_bit1(fabric_io_west_config_bit1_o[16]),
        .Tile_X0Y6_B_config_C_bit2(fabric_io_west_config_bit2_o[16]),
        .Tile_X0Y6_B_config_C_bit3(fabric_io_west_config_bit3_o[16]),

        .Tile_X0Y7_A_O_top(fabric_io_west_in_i[15]),
        .Tile_X0Y7_A_I_top(fabric_io_west_out_o[15]),
        .Tile_X0Y7_A_T_top(fabric_io_west_oe_o[15]),

        .Tile_X0Y7_B_O_top(fabric_io_west_in_i[14]),
        .Tile_X0Y7_B_I_top(fabric_io_west_out_o[14]),
        .Tile_X0Y7_B_T_top(fabric_io_west_oe_o[14]),

        .Tile_X0Y7_A_config_C_bit0(fabric_io_west_config_bit0_o[15]),
        .Tile_X0Y7_A_config_C_bit1(fabric_io_west_config_bit1_o[15]),
        .Tile_X0Y7_A_config_C_bit2(fabric_io_west_config_bit2_o[15]),
        .Tile_X0Y7_A_config_C_bit3(fabric_io_west_config_bit3_o[15]),

        .Tile_X0Y7_B_config_C_bit0(fabric_io_west_config_bit0_o[14]),
        .Tile_X0Y7_B_config_C_bit1(fabric_io_west_config_bit1_o[14]),
        .Tile_X0Y7_B_config_C_bit2(fabric_io_west_config_bit2_o[14]),
        .Tile_X0Y7_B_config_C_bit3(fabric_io_west_config_bit3_o[14]),

        .Tile_X0Y8_A_O_top(fabric_io_west_in_i[13]),
        .Tile_X0Y8_A_I_top(fabric_io_west_out_o[13]),
        .Tile_X0Y8_A_T_top(fabric_io_west_oe_o[13]),

        .Tile_X0Y8_B_O_top(fabric_io_west_in_i[12]),
        .Tile_X0Y8_B_I_top(fabric_io_west_out_o[12]),
        .Tile_X0Y8_B_T_top(fabric_io_west_oe_o[12]),

        .Tile_X0Y8_A_config_C_bit0(fabric_io_west_config_bit0_o[13]),
        .Tile_X0Y8_A_config_C_bit1(fabric_io_west_config_bit1_o[13]),
        .Tile_X0Y8_A_config_C_bit2(fabric_io_west_config_bit2_o[13]),
        .Tile_X0Y8_A_config_C_bit3(fabric_io_west_config_bit3_o[13]),

        .Tile_X0Y8_B_config_C_bit0(fabric_io_west_config_bit0_o[12]),
        .Tile_X0Y8_B_config_C_bit1(fabric_io_west_config_bit1_o[12]),
        .Tile_X0Y8_B_config_C_bit2(fabric_io_west_config_bit2_o[12]),
        .Tile_X0Y8_B_config_C_bit3(fabric_io_west_config_bit3_o[12]),

        .Tile_X0Y9_A_O_top(fabric_io_west_in_i[11]),
        .Tile_X0Y9_A_I_top(fabric_io_west_out_o[11]),
        .Tile_X0Y9_A_T_top(fabric_io_west_oe_o[11]),

        .Tile_X0Y9_B_O_top(fabric_io_west_in_i[10]),
        .Tile_X0Y9_B_I_top(fabric_io_west_out_o[10]),
        .Tile_X0Y9_B_T_top(fabric_io_west_oe_o[10]),

        .Tile_X0Y9_A_config_C_bit0(fabric_io_west_config_bit0_o[11]),
        .Tile_X0Y9_A_config_C_bit1(fabric_io_west_config_bit1_o[11]),
        .Tile_X0Y9_A_config_C_bit2(fabric_io_west_config_bit2_o[11]),
        .Tile_X0Y9_A_config_C_bit3(fabric_io_west_config_bit3_o[11]),

        .Tile_X0Y9_B_config_C_bit0(fabric_io_west_config_bit0_o[10]),
        .Tile_X0Y9_B_config_C_bit1(fabric_io_west_config_bit1_o[10]),
        .Tile_X0Y9_B_config_C_bit2(fabric_io_west_config_bit2_o[10]),
        .Tile_X0Y9_B_config_C_bit3(fabric_io_west_config_bit3_o[10]),

        .Tile_X0Y10_A_O_top(fabric_io_west_in_i[9]),
        .Tile_X0Y10_A_I_top(fabric_io_west_out_o[9]),
        .Tile_X0Y10_A_T_top(fabric_io_west_oe_o[9]),

        .Tile_X0Y10_B_O_top(fabric_io_west_in_i[8]),
        .Tile_X0Y10_B_I_top(fabric_io_west_out_o[8]),
        .Tile_X0Y10_B_T_top(fabric_io_west_oe_o[8]),

        .Tile_X0Y10_A_config_C_bit0(fabric_io_west_config_bit0_o[9]),
        .Tile_X0Y10_A_config_C_bit1(fabric_io_west_config_bit1_o[9]),
        .Tile_X0Y10_A_config_C_bit2(fabric_io_west_config_bit2_o[9]),
        .Tile_X0Y10_A_config_C_bit3(fabric_io_west_config_bit3_o[9]),

        .Tile_X0Y10_B_config_C_bit0(fabric_io_west_config_bit0_o[8]),
        .Tile_X0Y10_B_config_C_bit1(fabric_io_west_config_bit1_o[8]),
        .Tile_X0Y10_B_config_C_bit2(fabric_io_west_config_bit2_o[8]),
        .Tile_X0Y10_B_config_C_bit3(fabric_io_west_config_bit3_o[8]),

        .Tile_X0Y11_A_O_top(fabric_io_west_in_i[7]),
        .Tile_X0Y11_A_I_top(fabric_io_west_out_o[7]),
        .Tile_X0Y11_A_T_top(fabric_io_west_oe_o[7]),

        .Tile_X0Y11_B_O_top(fabric_io_west_in_i[6]),
        .Tile_X0Y11_B_I_top(fabric_io_west_out_o[6]),
        .Tile_X0Y11_B_T_top(fabric_io_west_oe_o[6]),

        .Tile_X0Y11_A_config_C_bit0(fabric_io_west_config_bit0_o[7]),
        .Tile_X0Y11_A_config_C_bit1(fabric_io_west_config_bit1_o[7]),
        .Tile_X0Y11_A_config_C_bit2(fabric_io_west_config_bit2_o[7]),
        .Tile_X0Y11_A_config_C_bit3(fabric_io_west_config_bit3_o[7]),

        .Tile_X0Y11_B_config_C_bit0(fabric_io_west_config_bit0_o[6]),
        .Tile_X0Y11_B_config_C_bit1(fabric_io_west_config_bit1_o[6]),
        .Tile_X0Y11_B_config_C_bit2(fabric_io_west_config_bit2_o[6]),
        .Tile_X0Y11_B_config_C_bit3(fabric_io_west_config_bit3_o[6]),

        .Tile_X0Y12_A_O_top(fabric_io_west_in_i[5]),
        .Tile_X0Y12_A_I_top(fabric_io_west_out_o[5]),
        .Tile_X0Y12_A_T_top(fabric_io_west_oe_o[5]),

        .Tile_X0Y12_B_O_top(fabric_io_west_in_i[4]),
        .Tile_X0Y12_B_I_top(fabric_io_west_out_o[4]),
        .Tile_X0Y12_B_T_top(fabric_io_west_oe_o[4]),

        .Tile_X0Y12_A_config_C_bit0(fabric_io_west_config_bit0_o[5]),
        .Tile_X0Y12_A_config_C_bit1(fabric_io_west_config_bit1_o[5]),
        .Tile_X0Y12_A_config_C_bit2(fabric_io_west_config_bit2_o[5]),
        .Tile_X0Y12_A_config_C_bit3(fabric_io_west_config_bit3_o[5]),

        .Tile_X0Y12_B_config_C_bit0(fabric_io_west_config_bit0_o[4]),
        .Tile_X0Y12_B_config_C_bit1(fabric_io_west_config_bit1_o[4]),
        .Tile_X0Y12_B_config_C_bit2(fabric_io_west_config_bit2_o[4]),
        .Tile_X0Y12_B_config_C_bit3(fabric_io_west_config_bit3_o[4]),

        .Tile_X0Y13_A_O_top(fabric_io_west_in_i[3]),
        .Tile_X0Y13_A_I_top(fabric_io_west_out_o[3]),
        .Tile_X0Y13_A_T_top(fabric_io_west_oe_o[3]),

        .Tile_X0Y13_B_O_top(fabric_io_west_in_i[2]),
        .Tile_X0Y13_B_I_top(fabric_io_west_out_o[2]),
        .Tile_X0Y13_B_T_top(fabric_io_west_oe_o[2]),

        .Tile_X0Y13_A_config_C_bit0(fabric_io_west_config_bit0_o[3]),
        .Tile_X0Y13_A_config_C_bit1(fabric_io_west_config_bit1_o[3]),
        .Tile_X0Y13_A_config_C_bit2(fabric_io_west_config_bit2_o[3]),
        .Tile_X0Y13_A_config_C_bit3(fabric_io_west_config_bit3_o[3]),

        .Tile_X0Y13_B_config_C_bit0(fabric_io_west_config_bit0_o[2]),
        .Tile_X0Y13_B_config_C_bit1(fabric_io_west_config_bit1_o[2]),
        .Tile_X0Y13_B_config_C_bit2(fabric_io_west_config_bit2_o[2]),
        .Tile_X0Y13_B_config_C_bit3(fabric_io_west_config_bit3_o[2]),

        .Tile_X0Y14_A_O_top(fabric_io_west_in_i[1]),
        .Tile_X0Y14_A_I_top(fabric_io_west_out_o[1]),
        .Tile_X0Y14_A_T_top(fabric_io_west_oe_o[1]),

        .Tile_X0Y14_B_O_top(fabric_io_west_in_i[0]),
        .Tile_X0Y14_B_I_top(fabric_io_west_out_o[0]),
        .Tile_X0Y14_B_T_top(fabric_io_west_oe_o[0]),

        .Tile_X0Y14_A_config_C_bit0(fabric_io_west_config_bit0_o[1]),
        .Tile_X0Y14_A_config_C_bit1(fabric_io_west_config_bit1_o[1]),
        .Tile_X0Y14_A_config_C_bit2(fabric_io_west_config_bit2_o[1]),
        .Tile_X0Y14_A_config_C_bit3(fabric_io_west_config_bit3_o[1]),

        .Tile_X0Y14_B_config_C_bit0(fabric_io_west_config_bit0_o[0]),
        .Tile_X0Y14_B_config_C_bit1(fabric_io_west_config_bit1_o[0]),
        .Tile_X0Y14_B_config_C_bit2(fabric_io_west_config_bit2_o[0]),
        .Tile_X0Y14_B_config_C_bit3(fabric_io_west_config_bit3_o[0]),

        // North I/Os
        .Tile_X1Y0_A_O_top(fabric_io_north_in_i[1]),
        .Tile_X1Y0_A_I_top(fabric_io_north_out_o[1]),
        .Tile_X1Y0_A_T_top(fabric_io_north_oe_o[1]),

        .Tile_X1Y0_B_O_top(fabric_io_north_in_i[0]),
        .Tile_X1Y0_B_I_top(fabric_io_north_out_o[0]),
        .Tile_X1Y0_B_T_top(fabric_io_north_oe_o[0]),

        .Tile_X1Y0_A_config_C_bit0(fabric_io_north_config_bit0_o[1]),
        .Tile_X1Y0_A_config_C_bit1(fabric_io_north_config_bit1_o[1]),
        .Tile_X1Y0_A_config_C_bit2(fabric_io_north_config_bit2_o[1]),
        .Tile_X1Y0_A_config_C_bit3(fabric_io_north_config_bit3_o[1]),

        .Tile_X1Y0_B_config_C_bit0(fabric_io_north_config_bit0_o[0]),
        .Tile_X1Y0_B_config_C_bit1(fabric_io_north_config_bit1_o[0]),
        .Tile_X1Y0_B_config_C_bit2(fabric_io_north_config_bit2_o[0]),
        .Tile_X1Y0_B_config_C_bit3(fabric_io_north_config_bit3_o[0]),

        .Tile_X2Y0_A_O_top(fabric_io_north_in_i[3]),
        .Tile_X2Y0_A_I_top(fabric_io_north_out_o[3]),
        .Tile_X2Y0_A_T_top(fabric_io_north_oe_o[3]),

        .Tile_X2Y0_B_O_top(fabric_io_north_in_i[2]),
        .Tile_X2Y0_B_I_top(fabric_io_north_out_o[2]),
        .Tile_X2Y0_B_T_top(fabric_io_north_oe_o[2]),

        .Tile_X2Y0_A_config_C_bit0(fabric_io_north_config_bit0_o[3]),
        .Tile_X2Y0_A_config_C_bit1(fabric_io_north_config_bit1_o[3]),
        .Tile_X2Y0_A_config_C_bit2(fabric_io_north_config_bit2_o[3]),
        .Tile_X2Y0_A_config_C_bit3(fabric_io_north_config_bit3_o[3]),

        .Tile_X2Y0_B_config_C_bit0(fabric_io_north_config_bit0_o[2]),
        .Tile_X2Y0_B_config_C_bit1(fabric_io_north_config_bit1_o[2]),
        .Tile_X2Y0_B_config_C_bit2(fabric_io_north_config_bit2_o[2]),
        .Tile_X2Y0_B_config_C_bit3(fabric_io_north_config_bit3_o[2]),

        // WARMBOOT
        .Tile_X2Y15_RESET_top(fabric_warmboot_reset_i),
        .Tile_X2Y15_BOOT_top(fabric_warmboot_boot_o),
        .Tile_X2Y15_SLOT_top0(fabric_warmboot_slot_o[0]),
        .Tile_X2Y15_SLOT_top1(fabric_warmboot_slot_o[1]),
        .Tile_X2Y15_SLOT_top2(fabric_warmboot_slot_o[2]),
        .Tile_X2Y15_SLOT_top3(fabric_warmboot_slot_o[3]),
        .Tile_X2Y15_CONFIGURED_top(configured_i),

        // IRQ
        .Tile_X3Y15_IRQ_top0(fabric_irq_o[0]),
        .Tile_X3Y15_IRQ_top1(fabric_irq_o[1]),
        .Tile_X3Y15_IRQ_top2(fabric_irq_o[2]),
        .Tile_X3Y15_IRQ_top3(fabric_irq_o[3]),
        .Tile_X3Y15_CONFIGURED_top(configured_i),

        // CPU_IF 0
        .Tile_X5Y15_I_top0(fabric_cpu_o[0]),
        .Tile_X5Y15_I_top1(fabric_cpu_o[1]),
        .Tile_X5Y15_I_top2(fabric_cpu_o[2]),
        .Tile_X5Y15_I_top3(fabric_cpu_o[3]),
        .Tile_X5Y15_I_top4(fabric_cpu_o[4]),
        .Tile_X5Y15_I_top5(fabric_cpu_o[5]),
        .Tile_X5Y15_I_top6(fabric_cpu_o[6]),
        .Tile_X5Y15_I_top7(fabric_cpu_o[7]),
        .Tile_X5Y15_I_top8(fabric_cpu_o[8]),
        .Tile_X5Y15_I_top9(fabric_cpu_o[9]),
        .Tile_X5Y15_I_top10(fabric_cpu_o[10]),
        .Tile_X5Y15_I_top11(fabric_cpu_o[11]),
        .Tile_X5Y15_I_top12(fabric_cpu_o[12]),
        .Tile_X5Y15_I_top13(fabric_cpu_o[13]),
        .Tile_X5Y15_I_top14(fabric_cpu_o[14]),
        .Tile_X5Y15_I_top15(fabric_cpu_o[15]),
        .Tile_X5Y15_O_top0(fabric_cpu_i[0]),
        .Tile_X5Y15_O_top1(fabric_cpu_i[1]),
        .Tile_X5Y15_O_top2(fabric_cpu_i[2]),
        .Tile_X5Y15_O_top3(fabric_cpu_i[3]),
        .Tile_X5Y15_O_top4(fabric_cpu_i[4]),
        .Tile_X5Y15_O_top5(fabric_cpu_i[5]),
        .Tile_X5Y15_O_top6(fabric_cpu_i[6]),
        .Tile_X5Y15_O_top7(fabric_cpu_i[7]),
        .Tile_X5Y15_O_top8(fabric_cpu_i[8]),
        .Tile_X5Y15_O_top9(fabric_cpu_i[9]),
        .Tile_X5Y15_O_top10(fabric_cpu_i[10]),
        .Tile_X5Y15_O_top11(fabric_cpu_i[11]),
        .Tile_X5Y15_O_top12(fabric_cpu_i[12]),
        .Tile_X5Y15_O_top13(fabric_cpu_i[13]),
        .Tile_X5Y15_O_top14(fabric_cpu_i[14]),
        .Tile_X5Y15_O_top15(fabric_cpu_i[15]),

        // CPU_IF 1
        .Tile_X6Y15_I_top0(fabric_cpu_o[16]),
        .Tile_X6Y15_I_top1(fabric_cpu_o[17]),
        .Tile_X6Y15_I_top2(fabric_cpu_o[18]),
        .Tile_X6Y15_I_top3(fabric_cpu_o[19]),
        .Tile_X6Y15_I_top4(fabric_cpu_o[20]),
        .Tile_X6Y15_I_top5(fabric_cpu_o[21]),
        .Tile_X6Y15_I_top6(fabric_cpu_o[22]),
        .Tile_X6Y15_I_top7(fabric_cpu_o[23]),
        .Tile_X6Y15_I_top8(fabric_cpu_o[24]),
        .Tile_X6Y15_I_top9(fabric_cpu_o[25]),
        .Tile_X6Y15_I_top10(fabric_cpu_o[26]),
        .Tile_X6Y15_I_top11(fabric_cpu_o[27]),
        .Tile_X6Y15_I_top12(fabric_cpu_o[28]),
        .Tile_X6Y15_I_top13(fabric_cpu_o[29]),
        .Tile_X6Y15_I_top14(fabric_cpu_o[30]),
        .Tile_X6Y15_I_top15(fabric_cpu_o[31]),
        .Tile_X6Y15_O_top0(fabric_cpu_i[16]),
        .Tile_X6Y15_O_top1(fabric_cpu_i[17]),
        .Tile_X6Y15_O_top2(fabric_cpu_i[18]),
        .Tile_X6Y15_O_top3(fabric_cpu_i[19]),
        .Tile_X6Y15_O_top4(fabric_cpu_i[20]),
        .Tile_X6Y15_O_top5(fabric_cpu_i[21]),
        .Tile_X6Y15_O_top6(fabric_cpu_i[22]),
        .Tile_X6Y15_O_top7(fabric_cpu_i[23]),
        .Tile_X6Y15_O_top8(fabric_cpu_i[24]),
        .Tile_X6Y15_O_top9(fabric_cpu_i[25]),
        .Tile_X6Y15_O_top10(fabric_cpu_i[26]),
        .Tile_X6Y15_O_top11(fabric_cpu_i[27]),
        .Tile_X6Y15_O_top12(fabric_cpu_i[28]),
        .Tile_X6Y15_O_top13(fabric_cpu_i[29]),
        .Tile_X6Y15_O_top14(fabric_cpu_i[30]),
        .Tile_X6Y15_O_top15(fabric_cpu_i[31]),

        // CPU_IF 2
        .Tile_X8Y15_I_top0(fabric_cpu_o[32]),
        .Tile_X8Y15_I_top1(fabric_cpu_o[33]),
        .Tile_X8Y15_I_top2(fabric_cpu_o[34]),
        .Tile_X8Y15_I_top3(fabric_cpu_o[35]),
        .Tile_X8Y15_I_top4(fabric_cpu_o[36]),
        .Tile_X8Y15_I_top5(fabric_cpu_o[37]),
        .Tile_X8Y15_I_top6(fabric_cpu_o[38]),
        .Tile_X8Y15_I_top7(fabric_cpu_o[39]),
        .Tile_X8Y15_I_top8(fabric_cpu_o[40]),
        .Tile_X8Y15_I_top9(fabric_cpu_o[41]),
        .Tile_X8Y15_I_top10(fabric_cpu_o[42]),
        .Tile_X8Y15_I_top11(fabric_cpu_o[43]),
        .Tile_X8Y15_I_top12(fabric_cpu_o[44]),
        .Tile_X8Y15_I_top13(fabric_cpu_o[45]),
        .Tile_X8Y15_I_top14(fabric_cpu_o[46]),
        .Tile_X8Y15_I_top15(fabric_cpu_o[47]),
        .Tile_X8Y15_O_top0(fabric_cpu_i[32]),
        .Tile_X8Y15_O_top1(fabric_cpu_i[33]),
        .Tile_X8Y15_O_top2(fabric_cpu_i[34]),
        .Tile_X8Y15_O_top3(fabric_cpu_i[35]),
        .Tile_X8Y15_O_top4(fabric_cpu_i[36]),
        .Tile_X8Y15_O_top5(fabric_cpu_i[37]),
        .Tile_X8Y15_O_top6(fabric_cpu_i[38]),
        .Tile_X8Y15_O_top7(fabric_cpu_i[39]),
        .Tile_X8Y15_O_top8(fabric_cpu_i[40]),
        .Tile_X8Y15_O_top9(fabric_cpu_i[41]),
        .Tile_X8Y15_O_top10(fabric_cpu_i[42]),
        .Tile_X8Y15_O_top11(fabric_cpu_i[43]),
        .Tile_X8Y15_O_top12(fabric_cpu_i[44]),
        .Tile_X8Y15_O_top13(fabric_cpu_i[45]),
        .Tile_X8Y15_O_top14(fabric_cpu_i[46]),
        .Tile_X8Y15_O_top15(fabric_cpu_i[47]),

        // CPU_IF 3
        .Tile_X9Y15_I_top0(fabric_cpu_o[48]),
        .Tile_X9Y15_I_top1(fabric_cpu_o[49]),
        .Tile_X9Y15_I_top2(fabric_cpu_o[50]),
        .Tile_X9Y15_I_top3(fabric_cpu_o[51]),
        .Tile_X9Y15_I_top4(fabric_cpu_o[52]),
        .Tile_X9Y15_I_top5(fabric_cpu_o[53]),
        .Tile_X9Y15_I_top6(fabric_cpu_o[54]),
        .Tile_X9Y15_I_top7(fabric_cpu_o[55]),
        .Tile_X9Y15_I_top8(fabric_cpu_o[56]),
        .Tile_X9Y15_I_top9(fabric_cpu_o[57]),
        .Tile_X9Y15_I_top10(fabric_cpu_o[58]),
        .Tile_X9Y15_I_top11(fabric_cpu_o[59]),
        .Tile_X9Y15_I_top12(fabric_cpu_o[60]),
        .Tile_X9Y15_I_top13(fabric_cpu_o[61]),
        .Tile_X9Y15_I_top14(fabric_cpu_o[62]),
        .Tile_X9Y15_I_top15(fabric_cpu_o[63]),
        .Tile_X9Y15_O_top0(fabric_cpu_i[48]),
        .Tile_X9Y15_O_top1(fabric_cpu_i[49]),
        .Tile_X9Y15_O_top2(fabric_cpu_i[50]),
        .Tile_X9Y15_O_top3(fabric_cpu_i[51]),
        .Tile_X9Y15_O_top4(fabric_cpu_i[52]),
        .Tile_X9Y15_O_top5(fabric_cpu_i[53]),
        .Tile_X9Y15_O_top6(fabric_cpu_i[54]),
        .Tile_X9Y15_O_top7(fabric_cpu_i[55]),
        .Tile_X9Y15_O_top8(fabric_cpu_i[56]),
        .Tile_X9Y15_O_top9(fabric_cpu_i[57]),
        .Tile_X9Y15_O_top10(fabric_cpu_i[58]),
        .Tile_X9Y15_O_top11(fabric_cpu_i[59]),
        .Tile_X9Y15_O_top12(fabric_cpu_i[60]),
        .Tile_X9Y15_O_top13(fabric_cpu_i[61]),
        .Tile_X9Y15_O_top14(fabric_cpu_i[62]),
        .Tile_X9Y15_O_top15(fabric_cpu_i[63]),

        // SRAM 0
        .Tile_X10Y2_DOUT_SRAM0(fabric_sram0_dout_i[0]),
        .Tile_X10Y2_DOUT_SRAM1(fabric_sram0_dout_i[1]),
        .Tile_X10Y2_DOUT_SRAM2(fabric_sram0_dout_i[2]),
        .Tile_X10Y2_DOUT_SRAM3(fabric_sram0_dout_i[3]),
        .Tile_X10Y2_DOUT_SRAM4(fabric_sram0_dout_i[4]),
        .Tile_X10Y2_DOUT_SRAM5(fabric_sram0_dout_i[5]),
        .Tile_X10Y2_DOUT_SRAM6(fabric_sram0_dout_i[6]),
        .Tile_X10Y2_DOUT_SRAM7(fabric_sram0_dout_i[7]),
        .Tile_X10Y2_DOUT_SRAM8(fabric_sram0_dout_i[8]),
        .Tile_X10Y2_DOUT_SRAM9(fabric_sram0_dout_i[9]),
        .Tile_X10Y2_DOUT_SRAM10(fabric_sram0_dout_i[10]),
        .Tile_X10Y2_DOUT_SRAM11(fabric_sram0_dout_i[11]),
        .Tile_X10Y2_DOUT_SRAM12(fabric_sram0_dout_i[12]),
        .Tile_X10Y2_DOUT_SRAM13(fabric_sram0_dout_i[13]),
        .Tile_X10Y2_DOUT_SRAM14(fabric_sram0_dout_i[14]),
        .Tile_X10Y2_DOUT_SRAM15(fabric_sram0_dout_i[15]),
        .Tile_X10Y2_DOUT_SRAM16(fabric_sram0_dout_i[16]),
        .Tile_X10Y2_DOUT_SRAM17(fabric_sram0_dout_i[17]),
        .Tile_X10Y2_DOUT_SRAM18(fabric_sram0_dout_i[18]),
        .Tile_X10Y2_DOUT_SRAM19(fabric_sram0_dout_i[19]),
        .Tile_X10Y2_DOUT_SRAM20(fabric_sram0_dout_i[20]),
        .Tile_X10Y2_DOUT_SRAM21(fabric_sram0_dout_i[21]),
        .Tile_X10Y2_DOUT_SRAM22(fabric_sram0_dout_i[22]),
        .Tile_X10Y2_DOUT_SRAM23(fabric_sram0_dout_i[23]),
        .Tile_X10Y2_DOUT_SRAM24(fabric_sram0_dout_i[24]),
        .Tile_X10Y2_DOUT_SRAM25(fabric_sram0_dout_i[25]),
        .Tile_X10Y2_DOUT_SRAM26(fabric_sram0_dout_i[26]),
        .Tile_X10Y2_DOUT_SRAM27(fabric_sram0_dout_i[27]),
        .Tile_X10Y2_DOUT_SRAM28(fabric_sram0_dout_i[28]),
        .Tile_X10Y2_DOUT_SRAM29(fabric_sram0_dout_i[29]),
        .Tile_X10Y2_DOUT_SRAM30(fabric_sram0_dout_i[30]),
        .Tile_X10Y2_DOUT_SRAM31(fabric_sram0_dout_i[31]),
        .Tile_X10Y2_ADDR_SRAM0(fabric_sram0_addr_o[0]),
        .Tile_X10Y2_ADDR_SRAM1(fabric_sram0_addr_o[1]),
        .Tile_X10Y2_ADDR_SRAM2(fabric_sram0_addr_o[2]),
        .Tile_X10Y2_ADDR_SRAM3(fabric_sram0_addr_o[3]),
        .Tile_X10Y2_ADDR_SRAM4(fabric_sram0_addr_o[4]),
        .Tile_X10Y2_ADDR_SRAM5(fabric_sram0_addr_o[5]),
        .Tile_X10Y2_ADDR_SRAM6(fabric_sram0_addr_o[6]),
        .Tile_X10Y2_ADDR_SRAM7(fabric_sram0_addr_o[7]),
        .Tile_X10Y2_ADDR_SRAM8(fabric_sram0_addr_o[8]),
        .Tile_X10Y2_ADDR_SRAM9(fabric_sram0_addr_o[9]),
        .Tile_X10Y2_BM_SRAM0(fabric_sram0_bm_o[0]),
        .Tile_X10Y2_BM_SRAM1(fabric_sram0_bm_o[1]),
        .Tile_X10Y2_BM_SRAM2(fabric_sram0_bm_o[2]),
        .Tile_X10Y2_BM_SRAM3(fabric_sram0_bm_o[3]),
        .Tile_X10Y2_BM_SRAM4(fabric_sram0_bm_o[4]),
        .Tile_X10Y2_BM_SRAM5(fabric_sram0_bm_o[5]),
        .Tile_X10Y2_BM_SRAM6(fabric_sram0_bm_o[6]),
        .Tile_X10Y2_BM_SRAM7(fabric_sram0_bm_o[7]),
        .Tile_X10Y2_BM_SRAM8(fabric_sram0_bm_o[8]),
        .Tile_X10Y2_BM_SRAM9(fabric_sram0_bm_o[9]),
        .Tile_X10Y2_BM_SRAM10(fabric_sram0_bm_o[10]),
        .Tile_X10Y2_BM_SRAM11(fabric_sram0_bm_o[11]),
        .Tile_X10Y2_BM_SRAM12(fabric_sram0_bm_o[12]),
        .Tile_X10Y2_BM_SRAM13(fabric_sram0_bm_o[13]),
        .Tile_X10Y2_BM_SRAM14(fabric_sram0_bm_o[14]),
        .Tile_X10Y2_BM_SRAM15(fabric_sram0_bm_o[15]),
        .Tile_X10Y2_BM_SRAM16(fabric_sram0_bm_o[16]),
        .Tile_X10Y2_BM_SRAM17(fabric_sram0_bm_o[17]),
        .Tile_X10Y2_BM_SRAM18(fabric_sram0_bm_o[18]),
        .Tile_X10Y2_BM_SRAM19(fabric_sram0_bm_o[19]),
        .Tile_X10Y2_BM_SRAM20(fabric_sram0_bm_o[20]),
        .Tile_X10Y2_BM_SRAM21(fabric_sram0_bm_o[21]),
        .Tile_X10Y2_BM_SRAM22(fabric_sram0_bm_o[22]),
        .Tile_X10Y2_BM_SRAM23(fabric_sram0_bm_o[23]),
        .Tile_X10Y2_BM_SRAM24(fabric_sram0_bm_o[24]),
        .Tile_X10Y2_BM_SRAM25(fabric_sram0_bm_o[25]),
        .Tile_X10Y2_BM_SRAM26(fabric_sram0_bm_o[26]),
        .Tile_X10Y2_BM_SRAM27(fabric_sram0_bm_o[27]),
        .Tile_X10Y2_BM_SRAM28(fabric_sram0_bm_o[28]),
        .Tile_X10Y2_BM_SRAM29(fabric_sram0_bm_o[29]),
        .Tile_X10Y2_BM_SRAM30(fabric_sram0_bm_o[30]),
        .Tile_X10Y2_BM_SRAM31(fabric_sram0_bm_o[31]),
        .Tile_X10Y2_DIN_SRAM0(fabric_sram0_din_o[0]),
        .Tile_X10Y2_DIN_SRAM1(fabric_sram0_din_o[1]),
        .Tile_X10Y2_DIN_SRAM2(fabric_sram0_din_o[2]),
        .Tile_X10Y2_DIN_SRAM3(fabric_sram0_din_o[3]),
        .Tile_X10Y2_DIN_SRAM4(fabric_sram0_din_o[4]),
        .Tile_X10Y2_DIN_SRAM5(fabric_sram0_din_o[5]),
        .Tile_X10Y2_DIN_SRAM6(fabric_sram0_din_o[6]),
        .Tile_X10Y2_DIN_SRAM7(fabric_sram0_din_o[7]),
        .Tile_X10Y2_DIN_SRAM8(fabric_sram0_din_o[8]),
        .Tile_X10Y2_DIN_SRAM9(fabric_sram0_din_o[9]),
        .Tile_X10Y2_DIN_SRAM10(fabric_sram0_din_o[10]),
        .Tile_X10Y2_DIN_SRAM11(fabric_sram0_din_o[11]),
        .Tile_X10Y2_DIN_SRAM12(fabric_sram0_din_o[12]),
        .Tile_X10Y2_DIN_SRAM13(fabric_sram0_din_o[13]),
        .Tile_X10Y2_DIN_SRAM14(fabric_sram0_din_o[14]),
        .Tile_X10Y2_DIN_SRAM15(fabric_sram0_din_o[15]),
        .Tile_X10Y2_DIN_SRAM16(fabric_sram0_din_o[16]),
        .Tile_X10Y2_DIN_SRAM17(fabric_sram0_din_o[17]),
        .Tile_X10Y2_DIN_SRAM18(fabric_sram0_din_o[18]),
        .Tile_X10Y2_DIN_SRAM19(fabric_sram0_din_o[19]),
        .Tile_X10Y2_DIN_SRAM20(fabric_sram0_din_o[20]),
        .Tile_X10Y2_DIN_SRAM21(fabric_sram0_din_o[21]),
        .Tile_X10Y2_DIN_SRAM22(fabric_sram0_din_o[22]),
        .Tile_X10Y2_DIN_SRAM23(fabric_sram0_din_o[23]),
        .Tile_X10Y2_DIN_SRAM24(fabric_sram0_din_o[24]),
        .Tile_X10Y2_DIN_SRAM25(fabric_sram0_din_o[25]),
        .Tile_X10Y2_DIN_SRAM26(fabric_sram0_din_o[26]),
        .Tile_X10Y2_DIN_SRAM27(fabric_sram0_din_o[27]),
        .Tile_X10Y2_DIN_SRAM28(fabric_sram0_din_o[28]),
        .Tile_X10Y2_DIN_SRAM29(fabric_sram0_din_o[29]),
        .Tile_X10Y2_DIN_SRAM30(fabric_sram0_din_o[30]),
        .Tile_X10Y2_DIN_SRAM31(fabric_sram0_din_o[31]),
        .Tile_X10Y2_WEN_SRAM(fabric_sram0_wen_o),
        .Tile_X10Y2_MEN_SRAM(fabric_sram0_men_o),
        .Tile_X10Y2_REN_SRAM(fabric_sram0_ren_o),
        .Tile_X10Y2_CLK_SRAM(fabric_sram0_clk_o),
        .Tile_X10Y2_TIE_HIGH_SRAM(fabric_sram0_tie_high_o),
        .Tile_X10Y2_TIE_LOW_SRAM(fabric_sram0_tie_low_o),
        .Tile_X10Y2_CONFIGURED_top(configured_i),

        // SRAM 1
        .Tile_X10Y4_DOUT_SRAM0(fabric_sram1_dout_i[0]),
        .Tile_X10Y4_DOUT_SRAM1(fabric_sram1_dout_i[1]),
        .Tile_X10Y4_DOUT_SRAM2(fabric_sram1_dout_i[2]),
        .Tile_X10Y4_DOUT_SRAM3(fabric_sram1_dout_i[3]),
        .Tile_X10Y4_DOUT_SRAM4(fabric_sram1_dout_i[4]),
        .Tile_X10Y4_DOUT_SRAM5(fabric_sram1_dout_i[5]),
        .Tile_X10Y4_DOUT_SRAM6(fabric_sram1_dout_i[6]),
        .Tile_X10Y4_DOUT_SRAM7(fabric_sram1_dout_i[7]),
        .Tile_X10Y4_DOUT_SRAM8(fabric_sram1_dout_i[8]),
        .Tile_X10Y4_DOUT_SRAM9(fabric_sram1_dout_i[9]),
        .Tile_X10Y4_DOUT_SRAM10(fabric_sram1_dout_i[10]),
        .Tile_X10Y4_DOUT_SRAM11(fabric_sram1_dout_i[11]),
        .Tile_X10Y4_DOUT_SRAM12(fabric_sram1_dout_i[12]),
        .Tile_X10Y4_DOUT_SRAM13(fabric_sram1_dout_i[13]),
        .Tile_X10Y4_DOUT_SRAM14(fabric_sram1_dout_i[14]),
        .Tile_X10Y4_DOUT_SRAM15(fabric_sram1_dout_i[15]),
        .Tile_X10Y4_DOUT_SRAM16(fabric_sram1_dout_i[16]),
        .Tile_X10Y4_DOUT_SRAM17(fabric_sram1_dout_i[17]),
        .Tile_X10Y4_DOUT_SRAM18(fabric_sram1_dout_i[18]),
        .Tile_X10Y4_DOUT_SRAM19(fabric_sram1_dout_i[19]),
        .Tile_X10Y4_DOUT_SRAM20(fabric_sram1_dout_i[20]),
        .Tile_X10Y4_DOUT_SRAM21(fabric_sram1_dout_i[21]),
        .Tile_X10Y4_DOUT_SRAM22(fabric_sram1_dout_i[22]),
        .Tile_X10Y4_DOUT_SRAM23(fabric_sram1_dout_i[23]),
        .Tile_X10Y4_DOUT_SRAM24(fabric_sram1_dout_i[24]),
        .Tile_X10Y4_DOUT_SRAM25(fabric_sram1_dout_i[25]),
        .Tile_X10Y4_DOUT_SRAM26(fabric_sram1_dout_i[26]),
        .Tile_X10Y4_DOUT_SRAM27(fabric_sram1_dout_i[27]),
        .Tile_X10Y4_DOUT_SRAM28(fabric_sram1_dout_i[28]),
        .Tile_X10Y4_DOUT_SRAM29(fabric_sram1_dout_i[29]),
        .Tile_X10Y4_DOUT_SRAM30(fabric_sram1_dout_i[30]),
        .Tile_X10Y4_DOUT_SRAM31(fabric_sram1_dout_i[31]),
        .Tile_X10Y4_ADDR_SRAM0(fabric_sram1_addr_o[0]),
        .Tile_X10Y4_ADDR_SRAM1(fabric_sram1_addr_o[1]),
        .Tile_X10Y4_ADDR_SRAM2(fabric_sram1_addr_o[2]),
        .Tile_X10Y4_ADDR_SRAM3(fabric_sram1_addr_o[3]),
        .Tile_X10Y4_ADDR_SRAM4(fabric_sram1_addr_o[4]),
        .Tile_X10Y4_ADDR_SRAM5(fabric_sram1_addr_o[5]),
        .Tile_X10Y4_ADDR_SRAM6(fabric_sram1_addr_o[6]),
        .Tile_X10Y4_ADDR_SRAM7(fabric_sram1_addr_o[7]),
        .Tile_X10Y4_ADDR_SRAM8(fabric_sram1_addr_o[8]),
        .Tile_X10Y4_ADDR_SRAM9(fabric_sram1_addr_o[9]),
        .Tile_X10Y4_BM_SRAM0(fabric_sram1_bm_o[0]),
        .Tile_X10Y4_BM_SRAM1(fabric_sram1_bm_o[1]),
        .Tile_X10Y4_BM_SRAM2(fabric_sram1_bm_o[2]),
        .Tile_X10Y4_BM_SRAM3(fabric_sram1_bm_o[3]),
        .Tile_X10Y4_BM_SRAM4(fabric_sram1_bm_o[4]),
        .Tile_X10Y4_BM_SRAM5(fabric_sram1_bm_o[5]),
        .Tile_X10Y4_BM_SRAM6(fabric_sram1_bm_o[6]),
        .Tile_X10Y4_BM_SRAM7(fabric_sram1_bm_o[7]),
        .Tile_X10Y4_BM_SRAM8(fabric_sram1_bm_o[8]),
        .Tile_X10Y4_BM_SRAM9(fabric_sram1_bm_o[9]),
        .Tile_X10Y4_BM_SRAM10(fabric_sram1_bm_o[10]),
        .Tile_X10Y4_BM_SRAM11(fabric_sram1_bm_o[11]),
        .Tile_X10Y4_BM_SRAM12(fabric_sram1_bm_o[12]),
        .Tile_X10Y4_BM_SRAM13(fabric_sram1_bm_o[13]),
        .Tile_X10Y4_BM_SRAM14(fabric_sram1_bm_o[14]),
        .Tile_X10Y4_BM_SRAM15(fabric_sram1_bm_o[15]),
        .Tile_X10Y4_BM_SRAM16(fabric_sram1_bm_o[16]),
        .Tile_X10Y4_BM_SRAM17(fabric_sram1_bm_o[17]),
        .Tile_X10Y4_BM_SRAM18(fabric_sram1_bm_o[18]),
        .Tile_X10Y4_BM_SRAM19(fabric_sram1_bm_o[19]),
        .Tile_X10Y4_BM_SRAM20(fabric_sram1_bm_o[20]),
        .Tile_X10Y4_BM_SRAM21(fabric_sram1_bm_o[21]),
        .Tile_X10Y4_BM_SRAM22(fabric_sram1_bm_o[22]),
        .Tile_X10Y4_BM_SRAM23(fabric_sram1_bm_o[23]),
        .Tile_X10Y4_BM_SRAM24(fabric_sram1_bm_o[24]),
        .Tile_X10Y4_BM_SRAM25(fabric_sram1_bm_o[25]),
        .Tile_X10Y4_BM_SRAM26(fabric_sram1_bm_o[26]),
        .Tile_X10Y4_BM_SRAM27(fabric_sram1_bm_o[27]),
        .Tile_X10Y4_BM_SRAM28(fabric_sram1_bm_o[28]),
        .Tile_X10Y4_BM_SRAM29(fabric_sram1_bm_o[29]),
        .Tile_X10Y4_BM_SRAM30(fabric_sram1_bm_o[30]),
        .Tile_X10Y4_BM_SRAM31(fabric_sram1_bm_o[31]),
        .Tile_X10Y4_DIN_SRAM0(fabric_sram1_din_o[0]),
        .Tile_X10Y4_DIN_SRAM1(fabric_sram1_din_o[1]),
        .Tile_X10Y4_DIN_SRAM2(fabric_sram1_din_o[2]),
        .Tile_X10Y4_DIN_SRAM3(fabric_sram1_din_o[3]),
        .Tile_X10Y4_DIN_SRAM4(fabric_sram1_din_o[4]),
        .Tile_X10Y4_DIN_SRAM5(fabric_sram1_din_o[5]),
        .Tile_X10Y4_DIN_SRAM6(fabric_sram1_din_o[6]),
        .Tile_X10Y4_DIN_SRAM7(fabric_sram1_din_o[7]),
        .Tile_X10Y4_DIN_SRAM8(fabric_sram1_din_o[8]),
        .Tile_X10Y4_DIN_SRAM9(fabric_sram1_din_o[9]),
        .Tile_X10Y4_DIN_SRAM10(fabric_sram1_din_o[10]),
        .Tile_X10Y4_DIN_SRAM11(fabric_sram1_din_o[11]),
        .Tile_X10Y4_DIN_SRAM12(fabric_sram1_din_o[12]),
        .Tile_X10Y4_DIN_SRAM13(fabric_sram1_din_o[13]),
        .Tile_X10Y4_DIN_SRAM14(fabric_sram1_din_o[14]),
        .Tile_X10Y4_DIN_SRAM15(fabric_sram1_din_o[15]),
        .Tile_X10Y4_DIN_SRAM16(fabric_sram1_din_o[16]),
        .Tile_X10Y4_DIN_SRAM17(fabric_sram1_din_o[17]),
        .Tile_X10Y4_DIN_SRAM18(fabric_sram1_din_o[18]),
        .Tile_X10Y4_DIN_SRAM19(fabric_sram1_din_o[19]),
        .Tile_X10Y4_DIN_SRAM20(fabric_sram1_din_o[20]),
        .Tile_X10Y4_DIN_SRAM21(fabric_sram1_din_o[21]),
        .Tile_X10Y4_DIN_SRAM22(fabric_sram1_din_o[22]),
        .Tile_X10Y4_DIN_SRAM23(fabric_sram1_din_o[23]),
        .Tile_X10Y4_DIN_SRAM24(fabric_sram1_din_o[24]),
        .Tile_X10Y4_DIN_SRAM25(fabric_sram1_din_o[25]),
        .Tile_X10Y4_DIN_SRAM26(fabric_sram1_din_o[26]),
        .Tile_X10Y4_DIN_SRAM27(fabric_sram1_din_o[27]),
        .Tile_X10Y4_DIN_SRAM28(fabric_sram1_din_o[28]),
        .Tile_X10Y4_DIN_SRAM29(fabric_sram1_din_o[29]),
        .Tile_X10Y4_DIN_SRAM30(fabric_sram1_din_o[30]),
        .Tile_X10Y4_DIN_SRAM31(fabric_sram1_din_o[31]),
        .Tile_X10Y4_WEN_SRAM(fabric_sram1_wen_o),
        .Tile_X10Y4_MEN_SRAM(fabric_sram1_men_o),
        .Tile_X10Y4_REN_SRAM(fabric_sram1_ren_o),
        .Tile_X10Y4_CLK_SRAM(fabric_sram1_clk_o),
        .Tile_X10Y4_TIE_HIGH_SRAM(fabric_sram1_tie_high_o),
        .Tile_X10Y4_TIE_LOW_SRAM(fabric_sram1_tie_low_o),
        .Tile_X10Y4_CONFIGURED_top(configured_i),

        // SRAM 2
        .Tile_X10Y6_DOUT_SRAM0(fabric_sram2_dout_i[0]),
        .Tile_X10Y6_DOUT_SRAM1(fabric_sram2_dout_i[1]),
        .Tile_X10Y6_DOUT_SRAM2(fabric_sram2_dout_i[2]),
        .Tile_X10Y6_DOUT_SRAM3(fabric_sram2_dout_i[3]),
        .Tile_X10Y6_DOUT_SRAM4(fabric_sram2_dout_i[4]),
        .Tile_X10Y6_DOUT_SRAM5(fabric_sram2_dout_i[5]),
        .Tile_X10Y6_DOUT_SRAM6(fabric_sram2_dout_i[6]),
        .Tile_X10Y6_DOUT_SRAM7(fabric_sram2_dout_i[7]),
        .Tile_X10Y6_DOUT_SRAM8(fabric_sram2_dout_i[8]),
        .Tile_X10Y6_DOUT_SRAM9(fabric_sram2_dout_i[9]),
        .Tile_X10Y6_DOUT_SRAM10(fabric_sram2_dout_i[10]),
        .Tile_X10Y6_DOUT_SRAM11(fabric_sram2_dout_i[11]),
        .Tile_X10Y6_DOUT_SRAM12(fabric_sram2_dout_i[12]),
        .Tile_X10Y6_DOUT_SRAM13(fabric_sram2_dout_i[13]),
        .Tile_X10Y6_DOUT_SRAM14(fabric_sram2_dout_i[14]),
        .Tile_X10Y6_DOUT_SRAM15(fabric_sram2_dout_i[15]),
        .Tile_X10Y6_DOUT_SRAM16(fabric_sram2_dout_i[16]),
        .Tile_X10Y6_DOUT_SRAM17(fabric_sram2_dout_i[17]),
        .Tile_X10Y6_DOUT_SRAM18(fabric_sram2_dout_i[18]),
        .Tile_X10Y6_DOUT_SRAM19(fabric_sram2_dout_i[19]),
        .Tile_X10Y6_DOUT_SRAM20(fabric_sram2_dout_i[20]),
        .Tile_X10Y6_DOUT_SRAM21(fabric_sram2_dout_i[21]),
        .Tile_X10Y6_DOUT_SRAM22(fabric_sram2_dout_i[22]),
        .Tile_X10Y6_DOUT_SRAM23(fabric_sram2_dout_i[23]),
        .Tile_X10Y6_DOUT_SRAM24(fabric_sram2_dout_i[24]),
        .Tile_X10Y6_DOUT_SRAM25(fabric_sram2_dout_i[25]),
        .Tile_X10Y6_DOUT_SRAM26(fabric_sram2_dout_i[26]),
        .Tile_X10Y6_DOUT_SRAM27(fabric_sram2_dout_i[27]),
        .Tile_X10Y6_DOUT_SRAM28(fabric_sram2_dout_i[28]),
        .Tile_X10Y6_DOUT_SRAM29(fabric_sram2_dout_i[29]),
        .Tile_X10Y6_DOUT_SRAM30(fabric_sram2_dout_i[30]),
        .Tile_X10Y6_DOUT_SRAM31(fabric_sram2_dout_i[31]),
        .Tile_X10Y6_ADDR_SRAM0(fabric_sram2_addr_o[0]),
        .Tile_X10Y6_ADDR_SRAM1(fabric_sram2_addr_o[1]),
        .Tile_X10Y6_ADDR_SRAM2(fabric_sram2_addr_o[2]),
        .Tile_X10Y6_ADDR_SRAM3(fabric_sram2_addr_o[3]),
        .Tile_X10Y6_ADDR_SRAM4(fabric_sram2_addr_o[4]),
        .Tile_X10Y6_ADDR_SRAM5(fabric_sram2_addr_o[5]),
        .Tile_X10Y6_ADDR_SRAM6(fabric_sram2_addr_o[6]),
        .Tile_X10Y6_ADDR_SRAM7(fabric_sram2_addr_o[7]),
        .Tile_X10Y6_ADDR_SRAM8(fabric_sram2_addr_o[8]),
        .Tile_X10Y6_ADDR_SRAM9(fabric_sram2_addr_o[9]),
        .Tile_X10Y6_BM_SRAM0(fabric_sram2_bm_o[0]),
        .Tile_X10Y6_BM_SRAM1(fabric_sram2_bm_o[1]),
        .Tile_X10Y6_BM_SRAM2(fabric_sram2_bm_o[2]),
        .Tile_X10Y6_BM_SRAM3(fabric_sram2_bm_o[3]),
        .Tile_X10Y6_BM_SRAM4(fabric_sram2_bm_o[4]),
        .Tile_X10Y6_BM_SRAM5(fabric_sram2_bm_o[5]),
        .Tile_X10Y6_BM_SRAM6(fabric_sram2_bm_o[6]),
        .Tile_X10Y6_BM_SRAM7(fabric_sram2_bm_o[7]),
        .Tile_X10Y6_BM_SRAM8(fabric_sram2_bm_o[8]),
        .Tile_X10Y6_BM_SRAM9(fabric_sram2_bm_o[9]),
        .Tile_X10Y6_BM_SRAM10(fabric_sram2_bm_o[10]),
        .Tile_X10Y6_BM_SRAM11(fabric_sram2_bm_o[11]),
        .Tile_X10Y6_BM_SRAM12(fabric_sram2_bm_o[12]),
        .Tile_X10Y6_BM_SRAM13(fabric_sram2_bm_o[13]),
        .Tile_X10Y6_BM_SRAM14(fabric_sram2_bm_o[14]),
        .Tile_X10Y6_BM_SRAM15(fabric_sram2_bm_o[15]),
        .Tile_X10Y6_BM_SRAM16(fabric_sram2_bm_o[16]),
        .Tile_X10Y6_BM_SRAM17(fabric_sram2_bm_o[17]),
        .Tile_X10Y6_BM_SRAM18(fabric_sram2_bm_o[18]),
        .Tile_X10Y6_BM_SRAM19(fabric_sram2_bm_o[19]),
        .Tile_X10Y6_BM_SRAM20(fabric_sram2_bm_o[20]),
        .Tile_X10Y6_BM_SRAM21(fabric_sram2_bm_o[21]),
        .Tile_X10Y6_BM_SRAM22(fabric_sram2_bm_o[22]),
        .Tile_X10Y6_BM_SRAM23(fabric_sram2_bm_o[23]),
        .Tile_X10Y6_BM_SRAM24(fabric_sram2_bm_o[24]),
        .Tile_X10Y6_BM_SRAM25(fabric_sram2_bm_o[25]),
        .Tile_X10Y6_BM_SRAM26(fabric_sram2_bm_o[26]),
        .Tile_X10Y6_BM_SRAM27(fabric_sram2_bm_o[27]),
        .Tile_X10Y6_BM_SRAM28(fabric_sram2_bm_o[28]),
        .Tile_X10Y6_BM_SRAM29(fabric_sram2_bm_o[29]),
        .Tile_X10Y6_BM_SRAM30(fabric_sram2_bm_o[30]),
        .Tile_X10Y6_BM_SRAM31(fabric_sram2_bm_o[31]),
        .Tile_X10Y6_DIN_SRAM0(fabric_sram2_din_o[0]),
        .Tile_X10Y6_DIN_SRAM1(fabric_sram2_din_o[1]),
        .Tile_X10Y6_DIN_SRAM2(fabric_sram2_din_o[2]),
        .Tile_X10Y6_DIN_SRAM3(fabric_sram2_din_o[3]),
        .Tile_X10Y6_DIN_SRAM4(fabric_sram2_din_o[4]),
        .Tile_X10Y6_DIN_SRAM5(fabric_sram2_din_o[5]),
        .Tile_X10Y6_DIN_SRAM6(fabric_sram2_din_o[6]),
        .Tile_X10Y6_DIN_SRAM7(fabric_sram2_din_o[7]),
        .Tile_X10Y6_DIN_SRAM8(fabric_sram2_din_o[8]),
        .Tile_X10Y6_DIN_SRAM9(fabric_sram2_din_o[9]),
        .Tile_X10Y6_DIN_SRAM10(fabric_sram2_din_o[10]),
        .Tile_X10Y6_DIN_SRAM11(fabric_sram2_din_o[11]),
        .Tile_X10Y6_DIN_SRAM12(fabric_sram2_din_o[12]),
        .Tile_X10Y6_DIN_SRAM13(fabric_sram2_din_o[13]),
        .Tile_X10Y6_DIN_SRAM14(fabric_sram2_din_o[14]),
        .Tile_X10Y6_DIN_SRAM15(fabric_sram2_din_o[15]),
        .Tile_X10Y6_DIN_SRAM16(fabric_sram2_din_o[16]),
        .Tile_X10Y6_DIN_SRAM17(fabric_sram2_din_o[17]),
        .Tile_X10Y6_DIN_SRAM18(fabric_sram2_din_o[18]),
        .Tile_X10Y6_DIN_SRAM19(fabric_sram2_din_o[19]),
        .Tile_X10Y6_DIN_SRAM20(fabric_sram2_din_o[20]),
        .Tile_X10Y6_DIN_SRAM21(fabric_sram2_din_o[21]),
        .Tile_X10Y6_DIN_SRAM22(fabric_sram2_din_o[22]),
        .Tile_X10Y6_DIN_SRAM23(fabric_sram2_din_o[23]),
        .Tile_X10Y6_DIN_SRAM24(fabric_sram2_din_o[24]),
        .Tile_X10Y6_DIN_SRAM25(fabric_sram2_din_o[25]),
        .Tile_X10Y6_DIN_SRAM26(fabric_sram2_din_o[26]),
        .Tile_X10Y6_DIN_SRAM27(fabric_sram2_din_o[27]),
        .Tile_X10Y6_DIN_SRAM28(fabric_sram2_din_o[28]),
        .Tile_X10Y6_DIN_SRAM29(fabric_sram2_din_o[29]),
        .Tile_X10Y6_DIN_SRAM30(fabric_sram2_din_o[30]),
        .Tile_X10Y6_DIN_SRAM31(fabric_sram2_din_o[31]),
        .Tile_X10Y6_WEN_SRAM(fabric_sram2_wen_o),
        .Tile_X10Y6_MEN_SRAM(fabric_sram2_men_o),
        .Tile_X10Y6_REN_SRAM(fabric_sram2_ren_o),
        .Tile_X10Y6_CLK_SRAM(fabric_sram2_clk_o),
        .Tile_X10Y6_TIE_HIGH_SRAM(fabric_sram2_tie_high_o),
        .Tile_X10Y6_TIE_LOW_SRAM(fabric_sram2_tie_low_o),
        .Tile_X10Y6_CONFIGURED_top(configured_i),

        // SRAM 3
        .Tile_X10Y8_DOUT_SRAM0(fabric_sram3_dout_i[0]),
        .Tile_X10Y8_DOUT_SRAM1(fabric_sram3_dout_i[1]),
        .Tile_X10Y8_DOUT_SRAM2(fabric_sram3_dout_i[2]),
        .Tile_X10Y8_DOUT_SRAM3(fabric_sram3_dout_i[3]),
        .Tile_X10Y8_DOUT_SRAM4(fabric_sram3_dout_i[4]),
        .Tile_X10Y8_DOUT_SRAM5(fabric_sram3_dout_i[5]),
        .Tile_X10Y8_DOUT_SRAM6(fabric_sram3_dout_i[6]),
        .Tile_X10Y8_DOUT_SRAM7(fabric_sram3_dout_i[7]),
        .Tile_X10Y8_DOUT_SRAM8(fabric_sram3_dout_i[8]),
        .Tile_X10Y8_DOUT_SRAM9(fabric_sram3_dout_i[9]),
        .Tile_X10Y8_DOUT_SRAM10(fabric_sram3_dout_i[10]),
        .Tile_X10Y8_DOUT_SRAM11(fabric_sram3_dout_i[11]),
        .Tile_X10Y8_DOUT_SRAM12(fabric_sram3_dout_i[12]),
        .Tile_X10Y8_DOUT_SRAM13(fabric_sram3_dout_i[13]),
        .Tile_X10Y8_DOUT_SRAM14(fabric_sram3_dout_i[14]),
        .Tile_X10Y8_DOUT_SRAM15(fabric_sram3_dout_i[15]),
        .Tile_X10Y8_DOUT_SRAM16(fabric_sram3_dout_i[16]),
        .Tile_X10Y8_DOUT_SRAM17(fabric_sram3_dout_i[17]),
        .Tile_X10Y8_DOUT_SRAM18(fabric_sram3_dout_i[18]),
        .Tile_X10Y8_DOUT_SRAM19(fabric_sram3_dout_i[19]),
        .Tile_X10Y8_DOUT_SRAM20(fabric_sram3_dout_i[20]),
        .Tile_X10Y8_DOUT_SRAM21(fabric_sram3_dout_i[21]),
        .Tile_X10Y8_DOUT_SRAM22(fabric_sram3_dout_i[22]),
        .Tile_X10Y8_DOUT_SRAM23(fabric_sram3_dout_i[23]),
        .Tile_X10Y8_DOUT_SRAM24(fabric_sram3_dout_i[24]),
        .Tile_X10Y8_DOUT_SRAM25(fabric_sram3_dout_i[25]),
        .Tile_X10Y8_DOUT_SRAM26(fabric_sram3_dout_i[26]),
        .Tile_X10Y8_DOUT_SRAM27(fabric_sram3_dout_i[27]),
        .Tile_X10Y8_DOUT_SRAM28(fabric_sram3_dout_i[28]),
        .Tile_X10Y8_DOUT_SRAM29(fabric_sram3_dout_i[29]),
        .Tile_X10Y8_DOUT_SRAM30(fabric_sram3_dout_i[30]),
        .Tile_X10Y8_DOUT_SRAM31(fabric_sram3_dout_i[31]),
        .Tile_X10Y8_ADDR_SRAM0(fabric_sram3_addr_o[0]),
        .Tile_X10Y8_ADDR_SRAM1(fabric_sram3_addr_o[1]),
        .Tile_X10Y8_ADDR_SRAM2(fabric_sram3_addr_o[2]),
        .Tile_X10Y8_ADDR_SRAM3(fabric_sram3_addr_o[3]),
        .Tile_X10Y8_ADDR_SRAM4(fabric_sram3_addr_o[4]),
        .Tile_X10Y8_ADDR_SRAM5(fabric_sram3_addr_o[5]),
        .Tile_X10Y8_ADDR_SRAM6(fabric_sram3_addr_o[6]),
        .Tile_X10Y8_ADDR_SRAM7(fabric_sram3_addr_o[7]),
        .Tile_X10Y8_ADDR_SRAM8(fabric_sram3_addr_o[8]),
        .Tile_X10Y8_ADDR_SRAM9(fabric_sram3_addr_o[9]),
        .Tile_X10Y8_BM_SRAM0(fabric_sram3_bm_o[0]),
        .Tile_X10Y8_BM_SRAM1(fabric_sram3_bm_o[1]),
        .Tile_X10Y8_BM_SRAM2(fabric_sram3_bm_o[2]),
        .Tile_X10Y8_BM_SRAM3(fabric_sram3_bm_o[3]),
        .Tile_X10Y8_BM_SRAM4(fabric_sram3_bm_o[4]),
        .Tile_X10Y8_BM_SRAM5(fabric_sram3_bm_o[5]),
        .Tile_X10Y8_BM_SRAM6(fabric_sram3_bm_o[6]),
        .Tile_X10Y8_BM_SRAM7(fabric_sram3_bm_o[7]),
        .Tile_X10Y8_BM_SRAM8(fabric_sram3_bm_o[8]),
        .Tile_X10Y8_BM_SRAM9(fabric_sram3_bm_o[9]),
        .Tile_X10Y8_BM_SRAM10(fabric_sram3_bm_o[10]),
        .Tile_X10Y8_BM_SRAM11(fabric_sram3_bm_o[11]),
        .Tile_X10Y8_BM_SRAM12(fabric_sram3_bm_o[12]),
        .Tile_X10Y8_BM_SRAM13(fabric_sram3_bm_o[13]),
        .Tile_X10Y8_BM_SRAM14(fabric_sram3_bm_o[14]),
        .Tile_X10Y8_BM_SRAM15(fabric_sram3_bm_o[15]),
        .Tile_X10Y8_BM_SRAM16(fabric_sram3_bm_o[16]),
        .Tile_X10Y8_BM_SRAM17(fabric_sram3_bm_o[17]),
        .Tile_X10Y8_BM_SRAM18(fabric_sram3_bm_o[18]),
        .Tile_X10Y8_BM_SRAM19(fabric_sram3_bm_o[19]),
        .Tile_X10Y8_BM_SRAM20(fabric_sram3_bm_o[20]),
        .Tile_X10Y8_BM_SRAM21(fabric_sram3_bm_o[21]),
        .Tile_X10Y8_BM_SRAM22(fabric_sram3_bm_o[22]),
        .Tile_X10Y8_BM_SRAM23(fabric_sram3_bm_o[23]),
        .Tile_X10Y8_BM_SRAM24(fabric_sram3_bm_o[24]),
        .Tile_X10Y8_BM_SRAM25(fabric_sram3_bm_o[25]),
        .Tile_X10Y8_BM_SRAM26(fabric_sram3_bm_o[26]),
        .Tile_X10Y8_BM_SRAM27(fabric_sram3_bm_o[27]),
        .Tile_X10Y8_BM_SRAM28(fabric_sram3_bm_o[28]),
        .Tile_X10Y8_BM_SRAM29(fabric_sram3_bm_o[29]),
        .Tile_X10Y8_BM_SRAM30(fabric_sram3_bm_o[30]),
        .Tile_X10Y8_BM_SRAM31(fabric_sram3_bm_o[31]),
        .Tile_X10Y8_DIN_SRAM0(fabric_sram3_din_o[0]),
        .Tile_X10Y8_DIN_SRAM1(fabric_sram3_din_o[1]),
        .Tile_X10Y8_DIN_SRAM2(fabric_sram3_din_o[2]),
        .Tile_X10Y8_DIN_SRAM3(fabric_sram3_din_o[3]),
        .Tile_X10Y8_DIN_SRAM4(fabric_sram3_din_o[4]),
        .Tile_X10Y8_DIN_SRAM5(fabric_sram3_din_o[5]),
        .Tile_X10Y8_DIN_SRAM6(fabric_sram3_din_o[6]),
        .Tile_X10Y8_DIN_SRAM7(fabric_sram3_din_o[7]),
        .Tile_X10Y8_DIN_SRAM8(fabric_sram3_din_o[8]),
        .Tile_X10Y8_DIN_SRAM9(fabric_sram3_din_o[9]),
        .Tile_X10Y8_DIN_SRAM10(fabric_sram3_din_o[10]),
        .Tile_X10Y8_DIN_SRAM11(fabric_sram3_din_o[11]),
        .Tile_X10Y8_DIN_SRAM12(fabric_sram3_din_o[12]),
        .Tile_X10Y8_DIN_SRAM13(fabric_sram3_din_o[13]),
        .Tile_X10Y8_DIN_SRAM14(fabric_sram3_din_o[14]),
        .Tile_X10Y8_DIN_SRAM15(fabric_sram3_din_o[15]),
        .Tile_X10Y8_DIN_SRAM16(fabric_sram3_din_o[16]),
        .Tile_X10Y8_DIN_SRAM17(fabric_sram3_din_o[17]),
        .Tile_X10Y8_DIN_SRAM18(fabric_sram3_din_o[18]),
        .Tile_X10Y8_DIN_SRAM19(fabric_sram3_din_o[19]),
        .Tile_X10Y8_DIN_SRAM20(fabric_sram3_din_o[20]),
        .Tile_X10Y8_DIN_SRAM21(fabric_sram3_din_o[21]),
        .Tile_X10Y8_DIN_SRAM22(fabric_sram3_din_o[22]),
        .Tile_X10Y8_DIN_SRAM23(fabric_sram3_din_o[23]),
        .Tile_X10Y8_DIN_SRAM24(fabric_sram3_din_o[24]),
        .Tile_X10Y8_DIN_SRAM25(fabric_sram3_din_o[25]),
        .Tile_X10Y8_DIN_SRAM26(fabric_sram3_din_o[26]),
        .Tile_X10Y8_DIN_SRAM27(fabric_sram3_din_o[27]),
        .Tile_X10Y8_DIN_SRAM28(fabric_sram3_din_o[28]),
        .Tile_X10Y8_DIN_SRAM29(fabric_sram3_din_o[29]),
        .Tile_X10Y8_DIN_SRAM30(fabric_sram3_din_o[30]),
        .Tile_X10Y8_DIN_SRAM31(fabric_sram3_din_o[31]),
        .Tile_X10Y8_WEN_SRAM(fabric_sram3_wen_o),
        .Tile_X10Y8_MEN_SRAM(fabric_sram3_men_o),
        .Tile_X10Y8_REN_SRAM(fabric_sram3_ren_o),
        .Tile_X10Y8_CLK_SRAM(fabric_sram3_clk_o),
        .Tile_X10Y8_TIE_HIGH_SRAM(fabric_sram3_tie_high_o),
        .Tile_X10Y8_TIE_LOW_SRAM(fabric_sram3_tie_low_o),
        .Tile_X10Y8_CONFIGURED_top(configured_i),

        // SRAM 4
        .Tile_X10Y10_DOUT_SRAM0(fabric_sram4_dout_i[0]),
        .Tile_X10Y10_DOUT_SRAM1(fabric_sram4_dout_i[1]),
        .Tile_X10Y10_DOUT_SRAM2(fabric_sram4_dout_i[2]),
        .Tile_X10Y10_DOUT_SRAM3(fabric_sram4_dout_i[3]),
        .Tile_X10Y10_DOUT_SRAM4(fabric_sram4_dout_i[4]),
        .Tile_X10Y10_DOUT_SRAM5(fabric_sram4_dout_i[5]),
        .Tile_X10Y10_DOUT_SRAM6(fabric_sram4_dout_i[6]),
        .Tile_X10Y10_DOUT_SRAM7(fabric_sram4_dout_i[7]),
        .Tile_X10Y10_DOUT_SRAM8(fabric_sram4_dout_i[8]),
        .Tile_X10Y10_DOUT_SRAM9(fabric_sram4_dout_i[9]),
        .Tile_X10Y10_DOUT_SRAM10(fabric_sram4_dout_i[10]),
        .Tile_X10Y10_DOUT_SRAM11(fabric_sram4_dout_i[11]),
        .Tile_X10Y10_DOUT_SRAM12(fabric_sram4_dout_i[12]),
        .Tile_X10Y10_DOUT_SRAM13(fabric_sram4_dout_i[13]),
        .Tile_X10Y10_DOUT_SRAM14(fabric_sram4_dout_i[14]),
        .Tile_X10Y10_DOUT_SRAM15(fabric_sram4_dout_i[15]),
        .Tile_X10Y10_DOUT_SRAM16(fabric_sram4_dout_i[16]),
        .Tile_X10Y10_DOUT_SRAM17(fabric_sram4_dout_i[17]),
        .Tile_X10Y10_DOUT_SRAM18(fabric_sram4_dout_i[18]),
        .Tile_X10Y10_DOUT_SRAM19(fabric_sram4_dout_i[19]),
        .Tile_X10Y10_DOUT_SRAM20(fabric_sram4_dout_i[20]),
        .Tile_X10Y10_DOUT_SRAM21(fabric_sram4_dout_i[21]),
        .Tile_X10Y10_DOUT_SRAM22(fabric_sram4_dout_i[22]),
        .Tile_X10Y10_DOUT_SRAM23(fabric_sram4_dout_i[23]),
        .Tile_X10Y10_DOUT_SRAM24(fabric_sram4_dout_i[24]),
        .Tile_X10Y10_DOUT_SRAM25(fabric_sram4_dout_i[25]),
        .Tile_X10Y10_DOUT_SRAM26(fabric_sram4_dout_i[26]),
        .Tile_X10Y10_DOUT_SRAM27(fabric_sram4_dout_i[27]),
        .Tile_X10Y10_DOUT_SRAM28(fabric_sram4_dout_i[28]),
        .Tile_X10Y10_DOUT_SRAM29(fabric_sram4_dout_i[29]),
        .Tile_X10Y10_DOUT_SRAM30(fabric_sram4_dout_i[30]),
        .Tile_X10Y10_DOUT_SRAM31(fabric_sram4_dout_i[31]),
        .Tile_X10Y10_ADDR_SRAM0(fabric_sram4_addr_o[0]),
        .Tile_X10Y10_ADDR_SRAM1(fabric_sram4_addr_o[1]),
        .Tile_X10Y10_ADDR_SRAM2(fabric_sram4_addr_o[2]),
        .Tile_X10Y10_ADDR_SRAM3(fabric_sram4_addr_o[3]),
        .Tile_X10Y10_ADDR_SRAM4(fabric_sram4_addr_o[4]),
        .Tile_X10Y10_ADDR_SRAM5(fabric_sram4_addr_o[5]),
        .Tile_X10Y10_ADDR_SRAM6(fabric_sram4_addr_o[6]),
        .Tile_X10Y10_ADDR_SRAM7(fabric_sram4_addr_o[7]),
        .Tile_X10Y10_ADDR_SRAM8(fabric_sram4_addr_o[8]),
        .Tile_X10Y10_ADDR_SRAM9(fabric_sram4_addr_o[9]),
        .Tile_X10Y10_BM_SRAM0(fabric_sram4_bm_o[0]),
        .Tile_X10Y10_BM_SRAM1(fabric_sram4_bm_o[1]),
        .Tile_X10Y10_BM_SRAM2(fabric_sram4_bm_o[2]),
        .Tile_X10Y10_BM_SRAM3(fabric_sram4_bm_o[3]),
        .Tile_X10Y10_BM_SRAM4(fabric_sram4_bm_o[4]),
        .Tile_X10Y10_BM_SRAM5(fabric_sram4_bm_o[5]),
        .Tile_X10Y10_BM_SRAM6(fabric_sram4_bm_o[6]),
        .Tile_X10Y10_BM_SRAM7(fabric_sram4_bm_o[7]),
        .Tile_X10Y10_BM_SRAM8(fabric_sram4_bm_o[8]),
        .Tile_X10Y10_BM_SRAM9(fabric_sram4_bm_o[9]),
        .Tile_X10Y10_BM_SRAM10(fabric_sram4_bm_o[10]),
        .Tile_X10Y10_BM_SRAM11(fabric_sram4_bm_o[11]),
        .Tile_X10Y10_BM_SRAM12(fabric_sram4_bm_o[12]),
        .Tile_X10Y10_BM_SRAM13(fabric_sram4_bm_o[13]),
        .Tile_X10Y10_BM_SRAM14(fabric_sram4_bm_o[14]),
        .Tile_X10Y10_BM_SRAM15(fabric_sram4_bm_o[15]),
        .Tile_X10Y10_BM_SRAM16(fabric_sram4_bm_o[16]),
        .Tile_X10Y10_BM_SRAM17(fabric_sram4_bm_o[17]),
        .Tile_X10Y10_BM_SRAM18(fabric_sram4_bm_o[18]),
        .Tile_X10Y10_BM_SRAM19(fabric_sram4_bm_o[19]),
        .Tile_X10Y10_BM_SRAM20(fabric_sram4_bm_o[20]),
        .Tile_X10Y10_BM_SRAM21(fabric_sram4_bm_o[21]),
        .Tile_X10Y10_BM_SRAM22(fabric_sram4_bm_o[22]),
        .Tile_X10Y10_BM_SRAM23(fabric_sram4_bm_o[23]),
        .Tile_X10Y10_BM_SRAM24(fabric_sram4_bm_o[24]),
        .Tile_X10Y10_BM_SRAM25(fabric_sram4_bm_o[25]),
        .Tile_X10Y10_BM_SRAM26(fabric_sram4_bm_o[26]),
        .Tile_X10Y10_BM_SRAM27(fabric_sram4_bm_o[27]),
        .Tile_X10Y10_BM_SRAM28(fabric_sram4_bm_o[28]),
        .Tile_X10Y10_BM_SRAM29(fabric_sram4_bm_o[29]),
        .Tile_X10Y10_BM_SRAM30(fabric_sram4_bm_o[30]),
        .Tile_X10Y10_BM_SRAM31(fabric_sram4_bm_o[31]),
        .Tile_X10Y10_DIN_SRAM0(fabric_sram4_din_o[0]),
        .Tile_X10Y10_DIN_SRAM1(fabric_sram4_din_o[1]),
        .Tile_X10Y10_DIN_SRAM2(fabric_sram4_din_o[2]),
        .Tile_X10Y10_DIN_SRAM3(fabric_sram4_din_o[3]),
        .Tile_X10Y10_DIN_SRAM4(fabric_sram4_din_o[4]),
        .Tile_X10Y10_DIN_SRAM5(fabric_sram4_din_o[5]),
        .Tile_X10Y10_DIN_SRAM6(fabric_sram4_din_o[6]),
        .Tile_X10Y10_DIN_SRAM7(fabric_sram4_din_o[7]),
        .Tile_X10Y10_DIN_SRAM8(fabric_sram4_din_o[8]),
        .Tile_X10Y10_DIN_SRAM9(fabric_sram4_din_o[9]),
        .Tile_X10Y10_DIN_SRAM10(fabric_sram4_din_o[10]),
        .Tile_X10Y10_DIN_SRAM11(fabric_sram4_din_o[11]),
        .Tile_X10Y10_DIN_SRAM12(fabric_sram4_din_o[12]),
        .Tile_X10Y10_DIN_SRAM13(fabric_sram4_din_o[13]),
        .Tile_X10Y10_DIN_SRAM14(fabric_sram4_din_o[14]),
        .Tile_X10Y10_DIN_SRAM15(fabric_sram4_din_o[15]),
        .Tile_X10Y10_DIN_SRAM16(fabric_sram4_din_o[16]),
        .Tile_X10Y10_DIN_SRAM17(fabric_sram4_din_o[17]),
        .Tile_X10Y10_DIN_SRAM18(fabric_sram4_din_o[18]),
        .Tile_X10Y10_DIN_SRAM19(fabric_sram4_din_o[19]),
        .Tile_X10Y10_DIN_SRAM20(fabric_sram4_din_o[20]),
        .Tile_X10Y10_DIN_SRAM21(fabric_sram4_din_o[21]),
        .Tile_X10Y10_DIN_SRAM22(fabric_sram4_din_o[22]),
        .Tile_X10Y10_DIN_SRAM23(fabric_sram4_din_o[23]),
        .Tile_X10Y10_DIN_SRAM24(fabric_sram4_din_o[24]),
        .Tile_X10Y10_DIN_SRAM25(fabric_sram4_din_o[25]),
        .Tile_X10Y10_DIN_SRAM26(fabric_sram4_din_o[26]),
        .Tile_X10Y10_DIN_SRAM27(fabric_sram4_din_o[27]),
        .Tile_X10Y10_DIN_SRAM28(fabric_sram4_din_o[28]),
        .Tile_X10Y10_DIN_SRAM29(fabric_sram4_din_o[29]),
        .Tile_X10Y10_DIN_SRAM30(fabric_sram4_din_o[30]),
        .Tile_X10Y10_DIN_SRAM31(fabric_sram4_din_o[31]),
        .Tile_X10Y10_WEN_SRAM(fabric_sram4_wen_o),
        .Tile_X10Y10_MEN_SRAM(fabric_sram4_men_o),
        .Tile_X10Y10_REN_SRAM(fabric_sram4_ren_o),
        .Tile_X10Y10_CLK_SRAM(fabric_sram4_clk_o),
        .Tile_X10Y10_TIE_HIGH_SRAM(fabric_sram4_tie_high_o),
        .Tile_X10Y10_TIE_LOW_SRAM(fabric_sram4_tie_low_o),
        .Tile_X10Y10_CONFIGURED_top(configured_i),

        // SRAM 5
        .Tile_X10Y12_DOUT_SRAM0(fabric_sram5_dout_i[0]),
        .Tile_X10Y12_DOUT_SRAM1(fabric_sram5_dout_i[1]),
        .Tile_X10Y12_DOUT_SRAM2(fabric_sram5_dout_i[2]),
        .Tile_X10Y12_DOUT_SRAM3(fabric_sram5_dout_i[3]),
        .Tile_X10Y12_DOUT_SRAM4(fabric_sram5_dout_i[4]),
        .Tile_X10Y12_DOUT_SRAM5(fabric_sram5_dout_i[5]),
        .Tile_X10Y12_DOUT_SRAM6(fabric_sram5_dout_i[6]),
        .Tile_X10Y12_DOUT_SRAM7(fabric_sram5_dout_i[7]),
        .Tile_X10Y12_DOUT_SRAM8(fabric_sram5_dout_i[8]),
        .Tile_X10Y12_DOUT_SRAM9(fabric_sram5_dout_i[9]),
        .Tile_X10Y12_DOUT_SRAM10(fabric_sram5_dout_i[10]),
        .Tile_X10Y12_DOUT_SRAM11(fabric_sram5_dout_i[11]),
        .Tile_X10Y12_DOUT_SRAM12(fabric_sram5_dout_i[12]),
        .Tile_X10Y12_DOUT_SRAM13(fabric_sram5_dout_i[13]),
        .Tile_X10Y12_DOUT_SRAM14(fabric_sram5_dout_i[14]),
        .Tile_X10Y12_DOUT_SRAM15(fabric_sram5_dout_i[15]),
        .Tile_X10Y12_DOUT_SRAM16(fabric_sram5_dout_i[16]),
        .Tile_X10Y12_DOUT_SRAM17(fabric_sram5_dout_i[17]),
        .Tile_X10Y12_DOUT_SRAM18(fabric_sram5_dout_i[18]),
        .Tile_X10Y12_DOUT_SRAM19(fabric_sram5_dout_i[19]),
        .Tile_X10Y12_DOUT_SRAM20(fabric_sram5_dout_i[20]),
        .Tile_X10Y12_DOUT_SRAM21(fabric_sram5_dout_i[21]),
        .Tile_X10Y12_DOUT_SRAM22(fabric_sram5_dout_i[22]),
        .Tile_X10Y12_DOUT_SRAM23(fabric_sram5_dout_i[23]),
        .Tile_X10Y12_DOUT_SRAM24(fabric_sram5_dout_i[24]),
        .Tile_X10Y12_DOUT_SRAM25(fabric_sram5_dout_i[25]),
        .Tile_X10Y12_DOUT_SRAM26(fabric_sram5_dout_i[26]),
        .Tile_X10Y12_DOUT_SRAM27(fabric_sram5_dout_i[27]),
        .Tile_X10Y12_DOUT_SRAM28(fabric_sram5_dout_i[28]),
        .Tile_X10Y12_DOUT_SRAM29(fabric_sram5_dout_i[29]),
        .Tile_X10Y12_DOUT_SRAM30(fabric_sram5_dout_i[30]),
        .Tile_X10Y12_DOUT_SRAM31(fabric_sram5_dout_i[31]),
        .Tile_X10Y12_ADDR_SRAM0(fabric_sram5_addr_o[0]),
        .Tile_X10Y12_ADDR_SRAM1(fabric_sram5_addr_o[1]),
        .Tile_X10Y12_ADDR_SRAM2(fabric_sram5_addr_o[2]),
        .Tile_X10Y12_ADDR_SRAM3(fabric_sram5_addr_o[3]),
        .Tile_X10Y12_ADDR_SRAM4(fabric_sram5_addr_o[4]),
        .Tile_X10Y12_ADDR_SRAM5(fabric_sram5_addr_o[5]),
        .Tile_X10Y12_ADDR_SRAM6(fabric_sram5_addr_o[6]),
        .Tile_X10Y12_ADDR_SRAM7(fabric_sram5_addr_o[7]),
        .Tile_X10Y12_ADDR_SRAM8(fabric_sram5_addr_o[8]),
        .Tile_X10Y12_ADDR_SRAM9(fabric_sram5_addr_o[9]),
        .Tile_X10Y12_BM_SRAM0(fabric_sram5_bm_o[0]),
        .Tile_X10Y12_BM_SRAM1(fabric_sram5_bm_o[1]),
        .Tile_X10Y12_BM_SRAM2(fabric_sram5_bm_o[2]),
        .Tile_X10Y12_BM_SRAM3(fabric_sram5_bm_o[3]),
        .Tile_X10Y12_BM_SRAM4(fabric_sram5_bm_o[4]),
        .Tile_X10Y12_BM_SRAM5(fabric_sram5_bm_o[5]),
        .Tile_X10Y12_BM_SRAM6(fabric_sram5_bm_o[6]),
        .Tile_X10Y12_BM_SRAM7(fabric_sram5_bm_o[7]),
        .Tile_X10Y12_BM_SRAM8(fabric_sram5_bm_o[8]),
        .Tile_X10Y12_BM_SRAM9(fabric_sram5_bm_o[9]),
        .Tile_X10Y12_BM_SRAM10(fabric_sram5_bm_o[10]),
        .Tile_X10Y12_BM_SRAM11(fabric_sram5_bm_o[11]),
        .Tile_X10Y12_BM_SRAM12(fabric_sram5_bm_o[12]),
        .Tile_X10Y12_BM_SRAM13(fabric_sram5_bm_o[13]),
        .Tile_X10Y12_BM_SRAM14(fabric_sram5_bm_o[14]),
        .Tile_X10Y12_BM_SRAM15(fabric_sram5_bm_o[15]),
        .Tile_X10Y12_BM_SRAM16(fabric_sram5_bm_o[16]),
        .Tile_X10Y12_BM_SRAM17(fabric_sram5_bm_o[17]),
        .Tile_X10Y12_BM_SRAM18(fabric_sram5_bm_o[18]),
        .Tile_X10Y12_BM_SRAM19(fabric_sram5_bm_o[19]),
        .Tile_X10Y12_BM_SRAM20(fabric_sram5_bm_o[20]),
        .Tile_X10Y12_BM_SRAM21(fabric_sram5_bm_o[21]),
        .Tile_X10Y12_BM_SRAM22(fabric_sram5_bm_o[22]),
        .Tile_X10Y12_BM_SRAM23(fabric_sram5_bm_o[23]),
        .Tile_X10Y12_BM_SRAM24(fabric_sram5_bm_o[24]),
        .Tile_X10Y12_BM_SRAM25(fabric_sram5_bm_o[25]),
        .Tile_X10Y12_BM_SRAM26(fabric_sram5_bm_o[26]),
        .Tile_X10Y12_BM_SRAM27(fabric_sram5_bm_o[27]),
        .Tile_X10Y12_BM_SRAM28(fabric_sram5_bm_o[28]),
        .Tile_X10Y12_BM_SRAM29(fabric_sram5_bm_o[29]),
        .Tile_X10Y12_BM_SRAM30(fabric_sram5_bm_o[30]),
        .Tile_X10Y12_BM_SRAM31(fabric_sram5_bm_o[31]),
        .Tile_X10Y12_DIN_SRAM0(fabric_sram5_din_o[0]),
        .Tile_X10Y12_DIN_SRAM1(fabric_sram5_din_o[1]),
        .Tile_X10Y12_DIN_SRAM2(fabric_sram5_din_o[2]),
        .Tile_X10Y12_DIN_SRAM3(fabric_sram5_din_o[3]),
        .Tile_X10Y12_DIN_SRAM4(fabric_sram5_din_o[4]),
        .Tile_X10Y12_DIN_SRAM5(fabric_sram5_din_o[5]),
        .Tile_X10Y12_DIN_SRAM6(fabric_sram5_din_o[6]),
        .Tile_X10Y12_DIN_SRAM7(fabric_sram5_din_o[7]),
        .Tile_X10Y12_DIN_SRAM8(fabric_sram5_din_o[8]),
        .Tile_X10Y12_DIN_SRAM9(fabric_sram5_din_o[9]),
        .Tile_X10Y12_DIN_SRAM10(fabric_sram5_din_o[10]),
        .Tile_X10Y12_DIN_SRAM11(fabric_sram5_din_o[11]),
        .Tile_X10Y12_DIN_SRAM12(fabric_sram5_din_o[12]),
        .Tile_X10Y12_DIN_SRAM13(fabric_sram5_din_o[13]),
        .Tile_X10Y12_DIN_SRAM14(fabric_sram5_din_o[14]),
        .Tile_X10Y12_DIN_SRAM15(fabric_sram5_din_o[15]),
        .Tile_X10Y12_DIN_SRAM16(fabric_sram5_din_o[16]),
        .Tile_X10Y12_DIN_SRAM17(fabric_sram5_din_o[17]),
        .Tile_X10Y12_DIN_SRAM18(fabric_sram5_din_o[18]),
        .Tile_X10Y12_DIN_SRAM19(fabric_sram5_din_o[19]),
        .Tile_X10Y12_DIN_SRAM20(fabric_sram5_din_o[20]),
        .Tile_X10Y12_DIN_SRAM21(fabric_sram5_din_o[21]),
        .Tile_X10Y12_DIN_SRAM22(fabric_sram5_din_o[22]),
        .Tile_X10Y12_DIN_SRAM23(fabric_sram5_din_o[23]),
        .Tile_X10Y12_DIN_SRAM24(fabric_sram5_din_o[24]),
        .Tile_X10Y12_DIN_SRAM25(fabric_sram5_din_o[25]),
        .Tile_X10Y12_DIN_SRAM26(fabric_sram5_din_o[26]),
        .Tile_X10Y12_DIN_SRAM27(fabric_sram5_din_o[27]),
        .Tile_X10Y12_DIN_SRAM28(fabric_sram5_din_o[28]),
        .Tile_X10Y12_DIN_SRAM29(fabric_sram5_din_o[29]),
        .Tile_X10Y12_DIN_SRAM30(fabric_sram5_din_o[30]),
        .Tile_X10Y12_DIN_SRAM31(fabric_sram5_din_o[31]),
        .Tile_X10Y12_WEN_SRAM(fabric_sram5_wen_o),
        .Tile_X10Y12_MEN_SRAM(fabric_sram5_men_o),
        .Tile_X10Y12_REN_SRAM(fabric_sram5_ren_o),
        .Tile_X10Y12_CLK_SRAM(fabric_sram5_clk_o),
        .Tile_X10Y12_TIE_HIGH_SRAM(fabric_sram5_tie_high_o),
        .Tile_X10Y12_TIE_LOW_SRAM(fabric_sram5_tie_low_o),
        .Tile_X10Y12_CONFIGURED_top(configured_i),

        // SRAM 6
        .Tile_X10Y14_DOUT_SRAM0(fabric_sram6_dout_i[0]),
        .Tile_X10Y14_DOUT_SRAM1(fabric_sram6_dout_i[1]),
        .Tile_X10Y14_DOUT_SRAM2(fabric_sram6_dout_i[2]),
        .Tile_X10Y14_DOUT_SRAM3(fabric_sram6_dout_i[3]),
        .Tile_X10Y14_DOUT_SRAM4(fabric_sram6_dout_i[4]),
        .Tile_X10Y14_DOUT_SRAM5(fabric_sram6_dout_i[5]),
        .Tile_X10Y14_DOUT_SRAM6(fabric_sram6_dout_i[6]),
        .Tile_X10Y14_DOUT_SRAM7(fabric_sram6_dout_i[7]),
        .Tile_X10Y14_DOUT_SRAM8(fabric_sram6_dout_i[8]),
        .Tile_X10Y14_DOUT_SRAM9(fabric_sram6_dout_i[9]),
        .Tile_X10Y14_DOUT_SRAM10(fabric_sram6_dout_i[10]),
        .Tile_X10Y14_DOUT_SRAM11(fabric_sram6_dout_i[11]),
        .Tile_X10Y14_DOUT_SRAM12(fabric_sram6_dout_i[12]),
        .Tile_X10Y14_DOUT_SRAM13(fabric_sram6_dout_i[13]),
        .Tile_X10Y14_DOUT_SRAM14(fabric_sram6_dout_i[14]),
        .Tile_X10Y14_DOUT_SRAM15(fabric_sram6_dout_i[15]),
        .Tile_X10Y14_DOUT_SRAM16(fabric_sram6_dout_i[16]),
        .Tile_X10Y14_DOUT_SRAM17(fabric_sram6_dout_i[17]),
        .Tile_X10Y14_DOUT_SRAM18(fabric_sram6_dout_i[18]),
        .Tile_X10Y14_DOUT_SRAM19(fabric_sram6_dout_i[19]),
        .Tile_X10Y14_DOUT_SRAM20(fabric_sram6_dout_i[20]),
        .Tile_X10Y14_DOUT_SRAM21(fabric_sram6_dout_i[21]),
        .Tile_X10Y14_DOUT_SRAM22(fabric_sram6_dout_i[22]),
        .Tile_X10Y14_DOUT_SRAM23(fabric_sram6_dout_i[23]),
        .Tile_X10Y14_DOUT_SRAM24(fabric_sram6_dout_i[24]),
        .Tile_X10Y14_DOUT_SRAM25(fabric_sram6_dout_i[25]),
        .Tile_X10Y14_DOUT_SRAM26(fabric_sram6_dout_i[26]),
        .Tile_X10Y14_DOUT_SRAM27(fabric_sram6_dout_i[27]),
        .Tile_X10Y14_DOUT_SRAM28(fabric_sram6_dout_i[28]),
        .Tile_X10Y14_DOUT_SRAM29(fabric_sram6_dout_i[29]),
        .Tile_X10Y14_DOUT_SRAM30(fabric_sram6_dout_i[30]),
        .Tile_X10Y14_DOUT_SRAM31(fabric_sram6_dout_i[31]),
        .Tile_X10Y14_ADDR_SRAM0(fabric_sram6_addr_o[0]),
        .Tile_X10Y14_ADDR_SRAM1(fabric_sram6_addr_o[1]),
        .Tile_X10Y14_ADDR_SRAM2(fabric_sram6_addr_o[2]),
        .Tile_X10Y14_ADDR_SRAM3(fabric_sram6_addr_o[3]),
        .Tile_X10Y14_ADDR_SRAM4(fabric_sram6_addr_o[4]),
        .Tile_X10Y14_ADDR_SRAM5(fabric_sram6_addr_o[5]),
        .Tile_X10Y14_ADDR_SRAM6(fabric_sram6_addr_o[6]),
        .Tile_X10Y14_ADDR_SRAM7(fabric_sram6_addr_o[7]),
        .Tile_X10Y14_ADDR_SRAM8(fabric_sram6_addr_o[8]),
        .Tile_X10Y14_ADDR_SRAM9(fabric_sram6_addr_o[9]),
        .Tile_X10Y14_BM_SRAM0(fabric_sram6_bm_o[0]),
        .Tile_X10Y14_BM_SRAM1(fabric_sram6_bm_o[1]),
        .Tile_X10Y14_BM_SRAM2(fabric_sram6_bm_o[2]),
        .Tile_X10Y14_BM_SRAM3(fabric_sram6_bm_o[3]),
        .Tile_X10Y14_BM_SRAM4(fabric_sram6_bm_o[4]),
        .Tile_X10Y14_BM_SRAM5(fabric_sram6_bm_o[5]),
        .Tile_X10Y14_BM_SRAM6(fabric_sram6_bm_o[6]),
        .Tile_X10Y14_BM_SRAM7(fabric_sram6_bm_o[7]),
        .Tile_X10Y14_BM_SRAM8(fabric_sram6_bm_o[8]),
        .Tile_X10Y14_BM_SRAM9(fabric_sram6_bm_o[9]),
        .Tile_X10Y14_BM_SRAM10(fabric_sram6_bm_o[10]),
        .Tile_X10Y14_BM_SRAM11(fabric_sram6_bm_o[11]),
        .Tile_X10Y14_BM_SRAM12(fabric_sram6_bm_o[12]),
        .Tile_X10Y14_BM_SRAM13(fabric_sram6_bm_o[13]),
        .Tile_X10Y14_BM_SRAM14(fabric_sram6_bm_o[14]),
        .Tile_X10Y14_BM_SRAM15(fabric_sram6_bm_o[15]),
        .Tile_X10Y14_BM_SRAM16(fabric_sram6_bm_o[16]),
        .Tile_X10Y14_BM_SRAM17(fabric_sram6_bm_o[17]),
        .Tile_X10Y14_BM_SRAM18(fabric_sram6_bm_o[18]),
        .Tile_X10Y14_BM_SRAM19(fabric_sram6_bm_o[19]),
        .Tile_X10Y14_BM_SRAM20(fabric_sram6_bm_o[20]),
        .Tile_X10Y14_BM_SRAM21(fabric_sram6_bm_o[21]),
        .Tile_X10Y14_BM_SRAM22(fabric_sram6_bm_o[22]),
        .Tile_X10Y14_BM_SRAM23(fabric_sram6_bm_o[23]),
        .Tile_X10Y14_BM_SRAM24(fabric_sram6_bm_o[24]),
        .Tile_X10Y14_BM_SRAM25(fabric_sram6_bm_o[25]),
        .Tile_X10Y14_BM_SRAM26(fabric_sram6_bm_o[26]),
        .Tile_X10Y14_BM_SRAM27(fabric_sram6_bm_o[27]),
        .Tile_X10Y14_BM_SRAM28(fabric_sram6_bm_o[28]),
        .Tile_X10Y14_BM_SRAM29(fabric_sram6_bm_o[29]),
        .Tile_X10Y14_BM_SRAM30(fabric_sram6_bm_o[30]),
        .Tile_X10Y14_BM_SRAM31(fabric_sram6_bm_o[31]),
        .Tile_X10Y14_DIN_SRAM0(fabric_sram6_din_o[0]),
        .Tile_X10Y14_DIN_SRAM1(fabric_sram6_din_o[1]),
        .Tile_X10Y14_DIN_SRAM2(fabric_sram6_din_o[2]),
        .Tile_X10Y14_DIN_SRAM3(fabric_sram6_din_o[3]),
        .Tile_X10Y14_DIN_SRAM4(fabric_sram6_din_o[4]),
        .Tile_X10Y14_DIN_SRAM5(fabric_sram6_din_o[5]),
        .Tile_X10Y14_DIN_SRAM6(fabric_sram6_din_o[6]),
        .Tile_X10Y14_DIN_SRAM7(fabric_sram6_din_o[7]),
        .Tile_X10Y14_DIN_SRAM8(fabric_sram6_din_o[8]),
        .Tile_X10Y14_DIN_SRAM9(fabric_sram6_din_o[9]),
        .Tile_X10Y14_DIN_SRAM10(fabric_sram6_din_o[10]),
        .Tile_X10Y14_DIN_SRAM11(fabric_sram6_din_o[11]),
        .Tile_X10Y14_DIN_SRAM12(fabric_sram6_din_o[12]),
        .Tile_X10Y14_DIN_SRAM13(fabric_sram6_din_o[13]),
        .Tile_X10Y14_DIN_SRAM14(fabric_sram6_din_o[14]),
        .Tile_X10Y14_DIN_SRAM15(fabric_sram6_din_o[15]),
        .Tile_X10Y14_DIN_SRAM16(fabric_sram6_din_o[16]),
        .Tile_X10Y14_DIN_SRAM17(fabric_sram6_din_o[17]),
        .Tile_X10Y14_DIN_SRAM18(fabric_sram6_din_o[18]),
        .Tile_X10Y14_DIN_SRAM19(fabric_sram6_din_o[19]),
        .Tile_X10Y14_DIN_SRAM20(fabric_sram6_din_o[20]),
        .Tile_X10Y14_DIN_SRAM21(fabric_sram6_din_o[21]),
        .Tile_X10Y14_DIN_SRAM22(fabric_sram6_din_o[22]),
        .Tile_X10Y14_DIN_SRAM23(fabric_sram6_din_o[23]),
        .Tile_X10Y14_DIN_SRAM24(fabric_sram6_din_o[24]),
        .Tile_X10Y14_DIN_SRAM25(fabric_sram6_din_o[25]),
        .Tile_X10Y14_DIN_SRAM26(fabric_sram6_din_o[26]),
        .Tile_X10Y14_DIN_SRAM27(fabric_sram6_din_o[27]),
        .Tile_X10Y14_DIN_SRAM28(fabric_sram6_din_o[28]),
        .Tile_X10Y14_DIN_SRAM29(fabric_sram6_din_o[29]),
        .Tile_X10Y14_DIN_SRAM30(fabric_sram6_din_o[30]),
        .Tile_X10Y14_DIN_SRAM31(fabric_sram6_din_o[31]),
        .Tile_X10Y14_WEN_SRAM(fabric_sram6_wen_o),
        .Tile_X10Y14_MEN_SRAM(fabric_sram6_men_o),
        .Tile_X10Y14_REN_SRAM(fabric_sram6_ren_o),
        .Tile_X10Y14_CLK_SRAM(fabric_sram6_clk_o),
        .Tile_X10Y14_TIE_HIGH_SRAM(fabric_sram6_tie_high_o),
        .Tile_X10Y14_TIE_LOW_SRAM(fabric_sram6_tie_low_o),
        .Tile_X10Y14_CONFIGURED_top(configured_i)
    );

    // SRAMs

    RM_IHPSG13_1P_1024x16_c2_bm_bist sram0_0 (
        .A_CLK      (fabric_sram0_clk_o),
        .A_MEN      (fabric_sram0_men_o),
        .A_WEN      (fabric_sram0_wen_o),
        .A_REN      (fabric_sram0_ren_o),
        .A_ADDR     (fabric_sram0_addr_o),
        .A_DIN      (fabric_sram0_din_o[15:0]),
        .A_DLY      (fabric_sram0_tie_high_o),
        .A_DOUT     (fabric_sram0_dout_i[15:0]),
        .A_BM       (fabric_sram0_bm_o[15:0]),

        .A_BIST_EN      (fabric_sram0_tie_low_o),
        .A_BIST_CLK     (fabric_sram0_tie_low_o),
        .A_BIST_MEN     (fabric_sram0_tie_low_o),
        .A_BIST_WEN     (fabric_sram0_tie_low_o),
        .A_BIST_REN     (fabric_sram0_tie_low_o),
        .A_BIST_ADDR    ({10{fabric_sram0_tie_low_o}}),
        .A_BIST_DIN     ({16{fabric_sram0_tie_low_o}}),
        .A_BIST_BM      ({16{fabric_sram0_tie_low_o}})
    );

    RM_IHPSG13_1P_1024x16_c2_bm_bist sram0_1 (
        .A_CLK      (fabric_sram0_clk_o),
        .A_MEN      (fabric_sram0_men_o),
        .A_WEN      (fabric_sram0_wen_o),
        .A_REN      (fabric_sram0_ren_o),
        .A_ADDR     (fabric_sram0_addr_o),
        .A_DIN      (fabric_sram0_din_o[31:16]),
        .A_DLY      (fabric_sram0_tie_high_o),
        .A_DOUT     (fabric_sram0_dout_i[31:16]),
        .A_BM       (fabric_sram0_bm_o[31:16]),

        .A_BIST_EN      (fabric_sram0_tie_low_o),
        .A_BIST_CLK     (fabric_sram0_tie_low_o),
        .A_BIST_MEN     (fabric_sram0_tie_low_o),
        .A_BIST_WEN     (fabric_sram0_tie_low_o),
        .A_BIST_REN     (fabric_sram0_tie_low_o),
        .A_BIST_ADDR    ({10{fabric_sram0_tie_low_o}}),
        .A_BIST_DIN     ({16{fabric_sram0_tie_low_o}}),
        .A_BIST_BM      ({16{fabric_sram0_tie_low_o}})
    );
    RM_IHPSG13_1P_1024x16_c2_bm_bist sram1_0 (
        .A_CLK      (fabric_sram1_clk_o),
        .A_MEN      (fabric_sram1_men_o),
        .A_WEN      (fabric_sram1_wen_o),
        .A_REN      (fabric_sram1_ren_o),
        .A_ADDR     (fabric_sram1_addr_o),
        .A_DIN      (fabric_sram1_din_o[15:0]),
        .A_DLY      (fabric_sram1_tie_high_o),
        .A_DOUT     (fabric_sram1_dout_i[15:0]),
        .A_BM       (fabric_sram1_bm_o[15:0]),

        .A_BIST_EN      (fabric_sram1_tie_low_o),
        .A_BIST_CLK     (fabric_sram1_tie_low_o),
        .A_BIST_MEN     (fabric_sram1_tie_low_o),
        .A_BIST_WEN     (fabric_sram1_tie_low_o),
        .A_BIST_REN     (fabric_sram1_tie_low_o),
        .A_BIST_ADDR    ({10{fabric_sram1_tie_low_o}}),
        .A_BIST_DIN     ({16{fabric_sram1_tie_low_o}}),
        .A_BIST_BM      ({16{fabric_sram1_tie_low_o}})
    );

    RM_IHPSG13_1P_1024x16_c2_bm_bist sram1_1 (
        .A_CLK      (fabric_sram1_clk_o),
        .A_MEN      (fabric_sram1_men_o),
        .A_WEN      (fabric_sram1_wen_o),
        .A_REN      (fabric_sram1_ren_o),
        .A_ADDR     (fabric_sram1_addr_o),
        .A_DIN      (fabric_sram1_din_o[31:16]),
        .A_DLY      (fabric_sram1_tie_high_o),
        .A_DOUT     (fabric_sram1_dout_i[31:16]),
        .A_BM       (fabric_sram1_bm_o[31:16]),

        .A_BIST_EN      (fabric_sram1_tie_low_o),
        .A_BIST_CLK     (fabric_sram1_tie_low_o),
        .A_BIST_MEN     (fabric_sram1_tie_low_o),
        .A_BIST_WEN     (fabric_sram1_tie_low_o),
        .A_BIST_REN     (fabric_sram1_tie_low_o),
        .A_BIST_ADDR    ({10{fabric_sram1_tie_low_o}}),
        .A_BIST_DIN     ({16{fabric_sram1_tie_low_o}}),
        .A_BIST_BM      ({16{fabric_sram1_tie_low_o}})
    );
    RM_IHPSG13_1P_1024x16_c2_bm_bist sram2_0 (
        .A_CLK      (fabric_sram2_clk_o),
        .A_MEN      (fabric_sram2_men_o),
        .A_WEN      (fabric_sram2_wen_o),
        .A_REN      (fabric_sram2_ren_o),
        .A_ADDR     (fabric_sram2_addr_o),
        .A_DIN      (fabric_sram2_din_o[15:0]),
        .A_DLY      (fabric_sram2_tie_high_o),
        .A_DOUT     (fabric_sram2_dout_i[15:0]),
        .A_BM       (fabric_sram2_bm_o[15:0]),

        .A_BIST_EN      (fabric_sram2_tie_low_o),
        .A_BIST_CLK     (fabric_sram2_tie_low_o),
        .A_BIST_MEN     (fabric_sram2_tie_low_o),
        .A_BIST_WEN     (fabric_sram2_tie_low_o),
        .A_BIST_REN     (fabric_sram2_tie_low_o),
        .A_BIST_ADDR    ({10{fabric_sram2_tie_low_o}}),
        .A_BIST_DIN     ({16{fabric_sram2_tie_low_o}}),
        .A_BIST_BM      ({16{fabric_sram2_tie_low_o}})
    );

    RM_IHPSG13_1P_1024x16_c2_bm_bist sram2_1 (
        .A_CLK      (fabric_sram2_clk_o),
        .A_MEN      (fabric_sram2_men_o),
        .A_WEN      (fabric_sram2_wen_o),
        .A_REN      (fabric_sram2_ren_o),
        .A_ADDR     (fabric_sram2_addr_o),
        .A_DIN      (fabric_sram2_din_o[31:16]),
        .A_DLY      (fabric_sram2_tie_high_o),
        .A_DOUT     (fabric_sram2_dout_i[31:16]),
        .A_BM       (fabric_sram2_bm_o[31:16]),

        .A_BIST_EN      (fabric_sram2_tie_low_o),
        .A_BIST_CLK     (fabric_sram2_tie_low_o),
        .A_BIST_MEN     (fabric_sram2_tie_low_o),
        .A_BIST_WEN     (fabric_sram2_tie_low_o),
        .A_BIST_REN     (fabric_sram2_tie_low_o),
        .A_BIST_ADDR    ({10{fabric_sram2_tie_low_o}}),
        .A_BIST_DIN     ({16{fabric_sram2_tie_low_o}}),
        .A_BIST_BM      ({16{fabric_sram2_tie_low_o}})
    );
    RM_IHPSG13_1P_1024x16_c2_bm_bist sram3_0 (
        .A_CLK      (fabric_sram3_clk_o),
        .A_MEN      (fabric_sram3_men_o),
        .A_WEN      (fabric_sram3_wen_o),
        .A_REN      (fabric_sram3_ren_o),
        .A_ADDR     (fabric_sram3_addr_o),
        .A_DIN      (fabric_sram3_din_o[15:0]),
        .A_DLY      (fabric_sram3_tie_high_o),
        .A_DOUT     (fabric_sram3_dout_i[15:0]),
        .A_BM       (fabric_sram3_bm_o[15:0]),

        .A_BIST_EN      (fabric_sram3_tie_low_o),
        .A_BIST_CLK     (fabric_sram3_tie_low_o),
        .A_BIST_MEN     (fabric_sram3_tie_low_o),
        .A_BIST_WEN     (fabric_sram3_tie_low_o),
        .A_BIST_REN     (fabric_sram3_tie_low_o),
        .A_BIST_ADDR    ({10{fabric_sram3_tie_low_o}}),
        .A_BIST_DIN     ({16{fabric_sram3_tie_low_o}}),
        .A_BIST_BM      ({16{fabric_sram3_tie_low_o}})
    );

    RM_IHPSG13_1P_1024x16_c2_bm_bist sram3_1 (
        .A_CLK      (fabric_sram3_clk_o),
        .A_MEN      (fabric_sram3_men_o),
        .A_WEN      (fabric_sram3_wen_o),
        .A_REN      (fabric_sram3_ren_o),
        .A_ADDR     (fabric_sram3_addr_o),
        .A_DIN      (fabric_sram3_din_o[31:16]),
        .A_DLY      (fabric_sram3_tie_high_o),
        .A_DOUT     (fabric_sram3_dout_i[31:16]),
        .A_BM       (fabric_sram3_bm_o[31:16]),

        .A_BIST_EN      (fabric_sram3_tie_low_o),
        .A_BIST_CLK     (fabric_sram3_tie_low_o),
        .A_BIST_MEN     (fabric_sram3_tie_low_o),
        .A_BIST_WEN     (fabric_sram3_tie_low_o),
        .A_BIST_REN     (fabric_sram3_tie_low_o),
        .A_BIST_ADDR    ({10{fabric_sram3_tie_low_o}}),
        .A_BIST_DIN     ({16{fabric_sram3_tie_low_o}}),
        .A_BIST_BM      ({16{fabric_sram3_tie_low_o}})
    );
    RM_IHPSG13_1P_1024x16_c2_bm_bist sram4_0 (
        .A_CLK      (fabric_sram4_clk_o),
        .A_MEN      (fabric_sram4_men_o),
        .A_WEN      (fabric_sram4_wen_o),
        .A_REN      (fabric_sram4_ren_o),
        .A_ADDR     (fabric_sram4_addr_o),
        .A_DIN      (fabric_sram4_din_o[15:0]),
        .A_DLY      (fabric_sram4_tie_high_o),
        .A_DOUT     (fabric_sram4_dout_i[15:0]),
        .A_BM       (fabric_sram4_bm_o[15:0]),

        .A_BIST_EN      (fabric_sram4_tie_low_o),
        .A_BIST_CLK     (fabric_sram4_tie_low_o),
        .A_BIST_MEN     (fabric_sram4_tie_low_o),
        .A_BIST_WEN     (fabric_sram4_tie_low_o),
        .A_BIST_REN     (fabric_sram4_tie_low_o),
        .A_BIST_ADDR    ({10{fabric_sram4_tie_low_o}}),
        .A_BIST_DIN     ({16{fabric_sram4_tie_low_o}}),
        .A_BIST_BM      ({16{fabric_sram4_tie_low_o}})
    );

    RM_IHPSG13_1P_1024x16_c2_bm_bist sram4_1 (
        .A_CLK      (fabric_sram4_clk_o),
        .A_MEN      (fabric_sram4_men_o),
        .A_WEN      (fabric_sram4_wen_o),
        .A_REN      (fabric_sram4_ren_o),
        .A_ADDR     (fabric_sram4_addr_o),
        .A_DIN      (fabric_sram4_din_o[31:16]),
        .A_DLY      (fabric_sram4_tie_high_o),
        .A_DOUT     (fabric_sram4_dout_i[31:16]),
        .A_BM       (fabric_sram4_bm_o[31:16]),

        .A_BIST_EN      (fabric_sram4_tie_low_o),
        .A_BIST_CLK     (fabric_sram4_tie_low_o),
        .A_BIST_MEN     (fabric_sram4_tie_low_o),
        .A_BIST_WEN     (fabric_sram4_tie_low_o),
        .A_BIST_REN     (fabric_sram4_tie_low_o),
        .A_BIST_ADDR    ({10{fabric_sram4_tie_low_o}}),
        .A_BIST_DIN     ({16{fabric_sram4_tie_low_o}}),
        .A_BIST_BM      ({16{fabric_sram4_tie_low_o}})
    );
    RM_IHPSG13_1P_1024x16_c2_bm_bist sram5_0 (
        .A_CLK      (fabric_sram5_clk_o),
        .A_MEN      (fabric_sram5_men_o),
        .A_WEN      (fabric_sram5_wen_o),
        .A_REN      (fabric_sram5_ren_o),
        .A_ADDR     (fabric_sram5_addr_o),
        .A_DIN      (fabric_sram5_din_o[15:0]),
        .A_DLY      (fabric_sram5_tie_high_o),
        .A_DOUT     (fabric_sram5_dout_i[15:0]),
        .A_BM       (fabric_sram5_bm_o[15:0]),

        .A_BIST_EN      (fabric_sram5_tie_low_o),
        .A_BIST_CLK     (fabric_sram5_tie_low_o),
        .A_BIST_MEN     (fabric_sram5_tie_low_o),
        .A_BIST_WEN     (fabric_sram5_tie_low_o),
        .A_BIST_REN     (fabric_sram5_tie_low_o),
        .A_BIST_ADDR    ({10{fabric_sram5_tie_low_o}}),
        .A_BIST_DIN     ({16{fabric_sram5_tie_low_o}}),
        .A_BIST_BM      ({16{fabric_sram5_tie_low_o}})
    );

    RM_IHPSG13_1P_1024x16_c2_bm_bist sram5_1 (
        .A_CLK      (fabric_sram5_clk_o),
        .A_MEN      (fabric_sram5_men_o),
        .A_WEN      (fabric_sram5_wen_o),
        .A_REN      (fabric_sram5_ren_o),
        .A_ADDR     (fabric_sram5_addr_o),
        .A_DIN      (fabric_sram5_din_o[31:16]),
        .A_DLY      (fabric_sram5_tie_high_o),
        .A_DOUT     (fabric_sram5_dout_i[31:16]),
        .A_BM       (fabric_sram5_bm_o[31:16]),

        .A_BIST_EN      (fabric_sram5_tie_low_o),
        .A_BIST_CLK     (fabric_sram5_tie_low_o),
        .A_BIST_MEN     (fabric_sram5_tie_low_o),
        .A_BIST_WEN     (fabric_sram5_tie_low_o),
        .A_BIST_REN     (fabric_sram5_tie_low_o),
        .A_BIST_ADDR    ({10{fabric_sram5_tie_low_o}}),
        .A_BIST_DIN     ({16{fabric_sram5_tie_low_o}}),
        .A_BIST_BM      ({16{fabric_sram5_tie_low_o}})
    );

    RM_IHPSG13_1P_1024x16_c2_bm_bist sram6_0 (
        .A_CLK      (fabric_sram6_clk_o),
        .A_MEN      (fabric_sram6_men_o),
        .A_WEN      (fabric_sram6_wen_o),
        .A_REN      (fabric_sram6_ren_o),
        .A_ADDR     (fabric_sram6_addr_o),
        .A_DIN      (fabric_sram6_din_o[15:0]),
        .A_DLY      (fabric_sram6_tie_high_o),
        .A_DOUT     (fabric_sram6_dout_i[15:0]),
        .A_BM       (fabric_sram6_bm_o[15:0]),

        .A_BIST_EN      (fabric_sram6_tie_low_o),
        .A_BIST_CLK     (fabric_sram6_tie_low_o),
        .A_BIST_MEN     (fabric_sram6_tie_low_o),
        .A_BIST_WEN     (fabric_sram6_tie_low_o),
        .A_BIST_REN     (fabric_sram6_tie_low_o),
        .A_BIST_ADDR    ({10{fabric_sram6_tie_low_o}}),
        .A_BIST_DIN     ({16{fabric_sram6_tie_low_o}}),
        .A_BIST_BM      ({16{fabric_sram6_tie_low_o}})
    );

    RM_IHPSG13_1P_1024x16_c2_bm_bist sram6_1 (
        .A_CLK      (fabric_sram6_clk_o),
        .A_MEN      (fabric_sram6_men_o),
        .A_WEN      (fabric_sram6_wen_o),
        .A_REN      (fabric_sram6_ren_o),
        .A_ADDR     (fabric_sram6_addr_o),
        .A_DIN      (fabric_sram6_din_o[31:16]),
        .A_DLY      (fabric_sram6_tie_high_o),
        .A_DOUT     (fabric_sram6_dout_i[31:16]),
        .A_BM       (fabric_sram6_bm_o[31:16]),

        .A_BIST_EN      (fabric_sram6_tie_low_o),
        .A_BIST_CLK     (fabric_sram6_tie_low_o),
        .A_BIST_MEN     (fabric_sram6_tie_low_o),
        .A_BIST_WEN     (fabric_sram6_tie_low_o),
        .A_BIST_REN     (fabric_sram6_tie_low_o),
        .A_BIST_ADDR    ({10{fabric_sram6_tie_low_o}}),
        .A_BIST_DIN     ({16{fabric_sram6_tie_low_o}}),
        .A_BIST_BM      ({16{fabric_sram6_tie_low_o}})
    );

endmodule

`default_nettype wire
