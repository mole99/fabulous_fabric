magic
tech ihp-sg13g2
magscale 1 2
timestamp 1743708635
<< metal2 >>
rect 0 701252 96 701272
rect 0 701212 13844 701252
rect 0 701192 96 701212
rect 0 700916 96 700936
rect 0 700876 13844 700916
rect 0 700856 96 700876
rect 0 700580 96 700600
rect 0 700540 13844 700580
rect 0 700520 96 700540
rect 0 700244 96 700264
rect 0 700204 13844 700244
rect 0 700184 96 700204
rect 0 699908 96 699928
rect 0 699868 13844 699908
rect 0 699848 96 699868
rect 0 699572 96 699592
rect 0 699532 13844 699572
rect 0 699512 96 699532
rect 0 699236 96 699256
rect 0 699196 13844 699236
rect 0 699176 96 699196
rect 0 698900 96 698920
rect 0 698860 13844 698900
rect 0 698840 96 698860
rect 0 698564 96 698584
rect 0 698524 13844 698564
rect 0 698504 96 698524
rect 0 698228 96 698248
rect 0 698188 13844 698228
rect 0 698168 96 698188
rect 0 697892 96 697912
rect 0 697852 13844 697892
rect 0 697832 96 697852
rect 0 697556 96 697576
rect 0 697516 13844 697556
rect 0 697496 96 697516
rect 0 697220 96 697240
rect 0 697180 13844 697220
rect 0 697160 96 697180
rect 0 696884 96 696904
rect 0 696844 13844 696884
rect 0 696824 96 696844
rect 0 696548 96 696568
rect 0 696508 13844 696548
rect 0 696488 96 696508
rect 0 696212 96 696232
rect 0 696172 13844 696212
rect 0 696152 96 696172
rect 0 695876 96 695896
rect 0 695836 13844 695876
rect 0 695816 96 695836
rect 0 695540 96 695560
rect 0 695500 13844 695540
rect 0 695480 96 695500
rect 0 695204 96 695224
rect 0 695164 13844 695204
rect 0 695144 96 695164
rect 0 694868 96 694888
rect 0 694828 13844 694868
rect 0 694808 96 694828
rect 0 694532 96 694552
rect 0 694492 13844 694532
rect 0 694472 96 694492
rect 0 694196 96 694216
rect 0 694156 13844 694196
rect 0 694136 96 694156
rect 0 693860 96 693880
rect 0 693820 13844 693860
rect 0 693800 96 693820
rect 0 693524 96 693544
rect 0 693484 13844 693524
rect 0 693464 96 693484
rect 0 693188 96 693208
rect 0 693148 13844 693188
rect 0 693128 96 693148
rect 0 692852 96 692872
rect 0 692812 13844 692852
rect 0 692792 96 692812
rect 0 692516 96 692536
rect 0 692476 13844 692516
rect 0 692456 96 692476
rect 0 692180 96 692200
rect 0 692140 13844 692180
rect 0 692120 96 692140
rect 0 691844 96 691864
rect 0 691804 13844 691844
rect 0 691784 96 691804
rect 0 691508 96 691528
rect 0 691468 13844 691508
rect 0 691448 96 691468
rect 0 691172 96 691192
rect 0 691132 13844 691172
rect 0 691112 96 691132
rect 0 690836 96 690856
rect 0 690796 13844 690836
rect 0 690776 96 690796
rect 0 688484 96 688504
rect 0 688444 116 688484
rect 0 688424 96 688444
rect 0 687476 96 687496
rect 0 687436 116 687476
rect 0 687416 96 687436
rect 0 686468 96 686488
rect 0 686428 116 686468
rect 0 686408 96 686428
rect 0 685460 96 685480
rect 0 685420 116 685460
rect 0 685400 96 685420
rect 0 684452 96 684472
rect 0 684412 116 684452
rect 0 684392 96 684412
rect 0 683444 96 683464
rect 0 683404 116 683444
rect 0 683384 96 683404
rect 0 682436 96 682456
rect 0 682396 116 682436
rect 0 682376 96 682396
rect 0 681428 96 681448
rect 0 681388 116 681428
rect 0 681368 96 681388
rect 0 680420 96 680440
rect 0 680380 116 680420
rect 0 680360 96 680380
rect 0 679412 96 679432
rect 0 679372 116 679412
rect 0 679352 96 679372
rect 0 678404 96 678424
rect 0 678364 116 678404
rect 0 678344 96 678364
rect 0 677396 96 677416
rect 0 677356 116 677396
rect 0 677336 96 677356
rect 0 676388 96 676408
rect 0 676348 116 676388
rect 0 676328 96 676348
rect 0 675380 96 675400
rect 0 675340 116 675380
rect 0 675320 96 675340
rect 0 674372 96 674392
rect 0 674332 116 674372
rect 0 674312 96 674332
rect 0 673364 96 673384
rect 0 673324 116 673364
rect 0 673304 96 673324
rect 0 672356 96 672376
rect 0 672316 116 672356
rect 0 672296 96 672316
rect 0 671348 96 671368
rect 0 671308 116 671348
rect 0 671288 96 671308
rect 0 670340 96 670360
rect 0 670300 116 670340
rect 0 670280 96 670300
rect 0 669332 96 669352
rect 0 669292 116 669332
rect 0 669272 96 669292
rect 0 668324 96 668344
rect 0 668284 116 668324
rect 0 668264 96 668284
rect 0 667316 96 667336
rect 0 667276 116 667316
rect 0 667256 96 667276
rect 0 666308 96 666328
rect 0 666268 116 666308
rect 0 666248 96 666268
rect 0 665300 96 665320
rect 0 665260 116 665300
rect 0 665240 96 665260
rect 0 664292 96 664312
rect 0 664252 116 664292
rect 0 664232 96 664252
rect 0 663284 96 663304
rect 0 663244 116 663284
rect 0 663224 96 663244
rect 0 662276 96 662296
rect 0 662236 116 662276
rect 0 662216 96 662236
rect 0 661268 96 661288
rect 0 661228 116 661268
rect 0 661208 96 661228
rect 0 660260 96 660280
rect 0 660220 116 660260
rect 0 660200 96 660220
rect 0 659252 96 659272
rect 0 659212 116 659252
rect 0 659192 96 659212
rect 0 658244 96 658264
rect 0 658204 116 658244
rect 0 658184 96 658204
rect 0 657236 96 657256
rect 0 657196 116 657236
rect 0 657176 96 657196
rect 0 656228 96 656248
rect 0 656188 116 656228
rect 0 656168 96 656188
rect 0 655220 96 655240
rect 0 655180 116 655220
rect 0 655160 96 655180
rect 0 654212 96 654232
rect 0 654172 116 654212
rect 0 654152 96 654172
rect 452544 653708 452640 653728
rect 452524 653668 452640 653708
rect 452544 653648 452640 653668
rect 0 653204 96 653224
rect 452544 653204 452640 653224
rect 0 653164 116 653204
rect 452524 653164 452640 653204
rect 0 653144 96 653164
rect 452544 653144 452640 653164
rect 452544 652700 452640 652720
rect 452524 652660 452640 652700
rect 452544 652640 452640 652660
rect 0 652196 96 652216
rect 452544 652196 452640 652216
rect 0 652156 116 652196
rect 452524 652156 452640 652196
rect 0 652136 96 652156
rect 452544 652136 452640 652156
rect 452544 651692 452640 651712
rect 452524 651652 452640 651692
rect 452544 651632 452640 651652
rect 0 651188 96 651208
rect 452544 651188 452640 651208
rect 0 651148 116 651188
rect 452524 651148 452640 651188
rect 0 651128 96 651148
rect 452544 651128 452640 651148
rect 452544 650684 452640 650704
rect 452524 650644 452640 650684
rect 452544 650624 452640 650644
rect 0 650180 96 650200
rect 452544 650180 452640 650200
rect 0 650140 116 650180
rect 452524 650140 452640 650180
rect 0 650120 96 650140
rect 452544 650120 452640 650140
rect 452544 649676 452640 649696
rect 452524 649636 452640 649676
rect 452544 649616 452640 649636
rect 0 649172 96 649192
rect 452544 649172 452640 649192
rect 0 649132 116 649172
rect 452524 649132 452640 649172
rect 0 649112 96 649132
rect 452544 649112 452640 649132
rect 452544 648668 452640 648688
rect 452524 648628 452640 648668
rect 452544 648608 452640 648628
rect 0 648164 96 648184
rect 452544 648164 452640 648184
rect 0 648124 116 648164
rect 452524 648124 452640 648164
rect 0 648104 96 648124
rect 452544 648104 452640 648124
rect 452544 647660 452640 647680
rect 452524 647620 452640 647660
rect 452544 647600 452640 647620
rect 0 647156 96 647176
rect 452544 647156 452640 647176
rect 0 647116 116 647156
rect 452524 647116 452640 647156
rect 0 647096 96 647116
rect 452544 647096 452640 647116
rect 452544 646652 452640 646672
rect 452524 646612 452640 646652
rect 452544 646592 452640 646612
rect 0 646148 96 646168
rect 452544 646148 452640 646168
rect 0 646108 116 646148
rect 452524 646108 452640 646148
rect 0 646088 96 646108
rect 452544 646088 452640 646108
rect 452544 645644 452640 645664
rect 452524 645604 452640 645644
rect 452544 645584 452640 645604
rect 0 645140 96 645160
rect 452544 645140 452640 645160
rect 0 645100 116 645140
rect 452524 645100 452640 645140
rect 0 645080 96 645100
rect 452544 645080 452640 645100
rect 452544 644636 452640 644656
rect 452524 644596 452640 644636
rect 452544 644576 452640 644596
rect 0 644132 96 644152
rect 452544 644132 452640 644152
rect 0 644092 116 644132
rect 452524 644092 452640 644132
rect 0 644072 96 644092
rect 452544 644072 452640 644092
rect 452544 643628 452640 643648
rect 452524 643588 452640 643628
rect 452544 643568 452640 643588
rect 0 643124 96 643144
rect 452544 643124 452640 643144
rect 0 643084 116 643124
rect 452524 643084 452640 643124
rect 0 643064 96 643084
rect 452544 643064 452640 643084
rect 452544 642620 452640 642640
rect 452524 642580 452640 642620
rect 452544 642560 452640 642580
rect 452544 642116 452640 642136
rect 452524 642076 452640 642116
rect 452544 642056 452640 642076
rect 452544 641612 452640 641632
rect 452524 641572 452640 641612
rect 452544 641552 452640 641572
rect 452544 641108 452640 641128
rect 452524 641068 452640 641108
rect 452544 641048 452640 641068
rect 452544 640604 452640 640624
rect 452524 640564 452640 640604
rect 452544 640544 452640 640564
rect 0 640100 96 640120
rect 452544 640100 452640 640120
rect 0 640060 116 640100
rect 452524 640060 452640 640100
rect 0 640040 96 640060
rect 452544 640040 452640 640060
rect 452544 639596 452640 639616
rect 452524 639556 452640 639596
rect 452544 639536 452640 639556
rect 0 639092 96 639112
rect 452544 639092 452640 639112
rect 0 639052 116 639092
rect 452524 639052 452640 639092
rect 0 639032 96 639052
rect 452544 639032 452640 639052
rect 452544 638588 452640 638608
rect 452524 638548 452640 638588
rect 452544 638528 452640 638548
rect 0 638084 96 638104
rect 452544 638084 452640 638104
rect 0 638044 116 638084
rect 452524 638044 452640 638084
rect 0 638024 96 638044
rect 452544 638024 452640 638044
rect 452544 637580 452640 637600
rect 452524 637540 452640 637580
rect 452544 637520 452640 637540
rect 0 637076 96 637096
rect 452544 637076 452640 637096
rect 0 637036 116 637076
rect 452524 637036 452640 637076
rect 0 637016 96 637036
rect 452544 637016 452640 637036
rect 452544 636572 452640 636592
rect 452524 636532 452640 636572
rect 452544 636512 452640 636532
rect 0 636068 96 636088
rect 452544 636068 452640 636088
rect 0 636028 116 636068
rect 452524 636028 452640 636068
rect 0 636008 96 636028
rect 452544 636008 452640 636028
rect 452544 635564 452640 635584
rect 452524 635524 452640 635564
rect 452544 635504 452640 635524
rect 0 635060 96 635080
rect 452544 635060 452640 635080
rect 0 635020 116 635060
rect 452524 635020 452640 635060
rect 0 635000 96 635020
rect 452544 635000 452640 635020
rect 452544 634556 452640 634576
rect 452524 634516 452640 634556
rect 452544 634496 452640 634516
rect 0 634052 96 634072
rect 452544 634052 452640 634072
rect 0 634012 116 634052
rect 452524 634012 452640 634052
rect 0 633992 96 634012
rect 452544 633992 452640 634012
rect 452544 633548 452640 633568
rect 452524 633508 452640 633548
rect 452544 633488 452640 633508
rect 0 633044 96 633064
rect 452544 633044 452640 633064
rect 0 633004 116 633044
rect 452524 633004 452640 633044
rect 0 632984 96 633004
rect 452544 632984 452640 633004
rect 452544 632540 452640 632560
rect 452524 632500 452640 632540
rect 452544 632480 452640 632500
rect 0 632036 96 632056
rect 452544 632036 452640 632056
rect 0 631996 116 632036
rect 452524 631996 452640 632036
rect 0 631976 96 631996
rect 452544 631976 452640 631996
rect 452544 631532 452640 631552
rect 452524 631492 452640 631532
rect 452544 631472 452640 631492
rect 0 631028 96 631048
rect 452544 631028 452640 631048
rect 0 630988 116 631028
rect 452524 630988 452640 631028
rect 0 630968 96 630988
rect 452544 630968 452640 630988
rect 452544 630524 452640 630544
rect 452524 630484 452640 630524
rect 452544 630464 452640 630484
rect 0 630020 96 630040
rect 452544 630020 452640 630040
rect 0 629980 116 630020
rect 452524 629980 452640 630020
rect 0 629960 96 629980
rect 452544 629960 452640 629980
rect 452544 629516 452640 629536
rect 452524 629476 452640 629516
rect 452544 629456 452640 629476
rect 0 629012 96 629032
rect 452544 629012 452640 629032
rect 0 628972 116 629012
rect 452524 628972 452640 629012
rect 0 628952 96 628972
rect 452544 628952 452640 628972
rect 452544 628508 452640 628528
rect 452524 628468 452640 628508
rect 452544 628448 452640 628468
rect 0 628004 96 628024
rect 452544 628004 452640 628024
rect 0 627964 116 628004
rect 452524 627964 452640 628004
rect 0 627944 96 627964
rect 452544 627944 452640 627964
rect 452544 627500 452640 627520
rect 452524 627460 452640 627500
rect 452544 627440 452640 627460
rect 0 626996 96 627016
rect 452544 626996 452640 627016
rect 0 626956 116 626996
rect 452524 626956 452640 626996
rect 0 626936 96 626956
rect 452544 626936 452640 626956
rect 452544 626492 452640 626512
rect 452524 626452 452640 626492
rect 452544 626432 452640 626452
rect 0 625988 96 626008
rect 452544 625988 452640 626008
rect 0 625948 116 625988
rect 452524 625948 452640 625988
rect 0 625928 96 625948
rect 452544 625928 452640 625948
rect 452544 625484 452640 625504
rect 452524 625444 452640 625484
rect 452544 625424 452640 625444
rect 0 624980 96 625000
rect 452544 624980 452640 625000
rect 0 624940 116 624980
rect 452524 624940 452640 624980
rect 0 624920 96 624940
rect 452544 624920 452640 624940
rect 452544 624476 452640 624496
rect 452524 624436 452640 624476
rect 452544 624416 452640 624436
rect 0 623972 96 623992
rect 452544 623972 452640 623992
rect 0 623932 116 623972
rect 452524 623932 452640 623972
rect 0 623912 96 623932
rect 452544 623912 452640 623932
rect 452544 623468 452640 623488
rect 452524 623428 452640 623468
rect 452544 623408 452640 623428
rect 0 622964 96 622984
rect 452544 622964 452640 622984
rect 0 622924 116 622964
rect 452524 622924 452640 622964
rect 0 622904 96 622924
rect 452544 622904 452640 622924
rect 452544 622460 452640 622480
rect 452524 622420 452640 622460
rect 452544 622400 452640 622420
rect 0 621956 96 621976
rect 452544 621956 452640 621976
rect 0 621916 116 621956
rect 452524 621916 452640 621956
rect 0 621896 96 621916
rect 452544 621896 452640 621916
rect 452544 621452 452640 621472
rect 452524 621412 452640 621452
rect 452544 621392 452640 621412
rect 0 620948 96 620968
rect 452544 620948 452640 620968
rect 0 620908 116 620948
rect 452524 620908 452640 620948
rect 0 620888 96 620908
rect 452544 620888 452640 620908
rect 452544 620444 452640 620464
rect 452524 620404 452640 620444
rect 452544 620384 452640 620404
rect 0 619940 96 619960
rect 452544 619940 452640 619960
rect 0 619900 116 619940
rect 452524 619900 452640 619940
rect 0 619880 96 619900
rect 452544 619880 452640 619900
rect 452544 619436 452640 619456
rect 452524 619396 452640 619436
rect 452544 619376 452640 619396
rect 0 618932 96 618952
rect 452544 618932 452640 618952
rect 0 618892 116 618932
rect 452524 618892 452640 618932
rect 0 618872 96 618892
rect 452544 618872 452640 618892
rect 452544 618428 452640 618448
rect 452524 618388 452640 618428
rect 452544 618368 452640 618388
rect 0 617924 96 617944
rect 452544 617924 452640 617944
rect 0 617884 116 617924
rect 452524 617884 452640 617924
rect 0 617864 96 617884
rect 452544 617864 452640 617884
rect 452544 617420 452640 617440
rect 452524 617380 452640 617420
rect 452544 617360 452640 617380
rect 0 616916 96 616936
rect 452544 616916 452640 616936
rect 0 616876 116 616916
rect 452524 616876 452640 616916
rect 0 616856 96 616876
rect 452544 616856 452640 616876
rect 452544 616412 452640 616432
rect 452524 616372 452640 616412
rect 452544 616352 452640 616372
rect 0 615908 96 615928
rect 452544 615908 452640 615928
rect 0 615868 116 615908
rect 452524 615868 452640 615908
rect 0 615848 96 615868
rect 452544 615848 452640 615868
rect 452544 615404 452640 615424
rect 452524 615364 452640 615404
rect 452544 615344 452640 615364
rect 0 614900 96 614920
rect 452544 614900 452640 614920
rect 0 614860 116 614900
rect 452524 614860 452640 614900
rect 0 614840 96 614860
rect 452544 614840 452640 614860
rect 452544 614396 452640 614416
rect 452524 614356 452640 614396
rect 452544 614336 452640 614356
rect 0 613892 96 613912
rect 452544 613892 452640 613912
rect 0 613852 116 613892
rect 452524 613852 452640 613892
rect 0 613832 96 613852
rect 452544 613832 452640 613852
rect 452544 613388 452640 613408
rect 452524 613348 452640 613388
rect 452544 613328 452640 613348
rect 0 612884 96 612904
rect 452544 612884 452640 612904
rect 0 612844 116 612884
rect 452524 612844 452640 612884
rect 0 612824 96 612844
rect 452544 612824 452640 612844
rect 452544 612380 452640 612400
rect 452524 612340 452640 612380
rect 452544 612320 452640 612340
rect 0 611876 96 611896
rect 452544 611876 452640 611896
rect 0 611836 116 611876
rect 452524 611836 452640 611876
rect 0 611816 96 611836
rect 452544 611816 452640 611836
rect 452544 611372 452640 611392
rect 452524 611332 452640 611372
rect 452544 611312 452640 611332
rect 0 610868 96 610888
rect 452544 610868 452640 610888
rect 0 610828 116 610868
rect 452524 610828 452640 610868
rect 0 610808 96 610828
rect 452544 610808 452640 610828
rect 452544 610364 452640 610384
rect 452524 610324 452640 610364
rect 452544 610304 452640 610324
rect 0 609860 96 609880
rect 452544 609860 452640 609880
rect 0 609820 116 609860
rect 452524 609820 452640 609860
rect 0 609800 96 609820
rect 452544 609800 452640 609820
rect 452544 609356 452640 609376
rect 452524 609316 452640 609356
rect 452544 609296 452640 609316
rect 0 608852 96 608872
rect 452544 608852 452640 608872
rect 0 608812 116 608852
rect 452524 608812 452640 608852
rect 0 608792 96 608812
rect 452544 608792 452640 608812
rect 452544 608348 452640 608368
rect 452524 608308 452640 608348
rect 452544 608288 452640 608308
rect 0 607844 96 607864
rect 452544 607844 452640 607864
rect 0 607804 116 607844
rect 452524 607804 452640 607844
rect 0 607784 96 607804
rect 452544 607784 452640 607804
rect 452544 607340 452640 607360
rect 452524 607300 452640 607340
rect 452544 607280 452640 607300
rect 0 606836 96 606856
rect 452544 606836 452640 606856
rect 0 606796 116 606836
rect 452524 606796 452640 606836
rect 0 606776 96 606796
rect 452544 606776 452640 606796
rect 452544 606332 452640 606352
rect 452524 606292 452640 606332
rect 452544 606272 452640 606292
rect 0 605828 96 605848
rect 452544 605828 452640 605848
rect 0 605788 116 605828
rect 452524 605788 452640 605828
rect 0 605768 96 605788
rect 452544 605768 452640 605788
rect 452544 605324 452640 605344
rect 452524 605284 452640 605324
rect 452544 605264 452640 605284
rect 0 604820 96 604840
rect 452544 604820 452640 604840
rect 0 604780 116 604820
rect 452524 604780 452640 604820
rect 0 604760 96 604780
rect 452544 604760 452640 604780
rect 452544 604316 452640 604336
rect 452524 604276 452640 604316
rect 452544 604256 452640 604276
rect 0 603812 96 603832
rect 452544 603812 452640 603832
rect 0 603772 116 603812
rect 452524 603772 452640 603812
rect 0 603752 96 603772
rect 452544 603752 452640 603772
rect 452544 603308 452640 603328
rect 452524 603268 452640 603308
rect 452544 603248 452640 603268
rect 0 602804 96 602824
rect 452544 602804 452640 602824
rect 0 602764 116 602804
rect 452524 602764 452640 602804
rect 0 602744 96 602764
rect 452544 602744 452640 602764
rect 452544 602300 452640 602320
rect 452524 602260 452640 602300
rect 452544 602240 452640 602260
rect 0 601796 96 601816
rect 452544 601796 452640 601816
rect 0 601756 116 601796
rect 452524 601756 452640 601796
rect 0 601736 96 601756
rect 452544 601736 452640 601756
rect 452544 601292 452640 601312
rect 452524 601252 452640 601292
rect 452544 601232 452640 601252
rect 0 600788 96 600808
rect 452544 600788 452640 600808
rect 0 600748 116 600788
rect 452524 600748 452640 600788
rect 0 600728 96 600748
rect 452544 600728 452640 600748
rect 452544 600284 452640 600304
rect 452524 600244 452640 600284
rect 452544 600224 452640 600244
rect 0 599780 96 599800
rect 452544 599780 452640 599800
rect 0 599740 116 599780
rect 452524 599740 452640 599780
rect 0 599720 96 599740
rect 452544 599720 452640 599740
rect 452544 599276 452640 599296
rect 452524 599236 452640 599276
rect 452544 599216 452640 599236
rect 0 598772 96 598792
rect 452544 598772 452640 598792
rect 0 598732 116 598772
rect 452524 598732 452640 598772
rect 0 598712 96 598732
rect 452544 598712 452640 598732
rect 452544 598268 452640 598288
rect 452524 598228 452640 598268
rect 452544 598208 452640 598228
rect 0 597764 96 597784
rect 452544 597764 452640 597784
rect 0 597724 116 597764
rect 452524 597724 452640 597764
rect 0 597704 96 597724
rect 452544 597704 452640 597724
rect 452544 597260 452640 597280
rect 452524 597220 452640 597260
rect 452544 597200 452640 597220
rect 0 596756 96 596776
rect 0 596716 116 596756
rect 0 596696 96 596716
rect 0 595748 96 595768
rect 0 595708 116 595748
rect 0 595688 96 595708
rect 0 594740 96 594760
rect 0 594700 116 594740
rect 0 594680 96 594700
rect 0 591716 96 591736
rect 0 591676 116 591716
rect 0 591656 96 591676
rect 0 590708 96 590728
rect 0 590668 116 590708
rect 0 590648 96 590668
rect 0 589700 96 589720
rect 0 589660 116 589700
rect 0 589640 96 589660
rect 0 588692 96 588712
rect 0 588652 116 588692
rect 0 588632 96 588652
rect 0 587684 96 587704
rect 0 587644 116 587684
rect 0 587624 96 587644
rect 0 586676 96 586696
rect 0 586636 116 586676
rect 0 586616 96 586636
rect 0 585668 96 585688
rect 0 585628 116 585668
rect 0 585608 96 585628
rect 0 584660 96 584680
rect 0 584620 116 584660
rect 0 584600 96 584620
rect 0 583652 96 583672
rect 0 583612 116 583652
rect 0 583592 96 583612
rect 0 582644 96 582664
rect 0 582604 116 582644
rect 0 582584 96 582604
rect 0 581636 96 581656
rect 0 581596 116 581636
rect 0 581576 96 581596
rect 0 580628 96 580648
rect 0 580588 116 580628
rect 0 580568 96 580588
rect 0 579620 96 579640
rect 0 579580 116 579620
rect 0 579560 96 579580
rect 0 578612 96 578632
rect 0 578572 116 578612
rect 0 578552 96 578572
rect 0 577604 96 577624
rect 0 577564 116 577604
rect 0 577544 96 577564
rect 0 576596 96 576616
rect 0 576556 116 576596
rect 0 576536 96 576556
rect 0 575588 96 575608
rect 0 575548 116 575588
rect 0 575528 96 575548
rect 0 574580 96 574600
rect 0 574540 116 574580
rect 0 574520 96 574540
rect 0 573572 96 573592
rect 0 573532 116 573572
rect 0 573512 96 573532
rect 0 572564 96 572584
rect 0 572524 116 572564
rect 0 572504 96 572524
rect 0 571556 96 571576
rect 0 571516 116 571556
rect 0 571496 96 571516
rect 0 570548 96 570568
rect 0 570508 116 570548
rect 0 570488 96 570508
rect 0 569540 96 569560
rect 0 569500 116 569540
rect 0 569480 96 569500
rect 0 568532 96 568552
rect 0 568492 116 568532
rect 0 568472 96 568492
rect 0 567524 96 567544
rect 0 567484 116 567524
rect 0 567464 96 567484
rect 0 566516 96 566536
rect 0 566476 116 566516
rect 0 566456 96 566476
rect 0 565508 96 565528
rect 0 565468 116 565508
rect 0 565448 96 565468
rect 0 564500 96 564520
rect 0 564460 116 564500
rect 0 564440 96 564460
rect 0 563492 96 563512
rect 0 563452 116 563492
rect 0 563432 96 563452
rect 0 562484 96 562504
rect 0 562444 116 562484
rect 0 562424 96 562444
rect 0 561476 96 561496
rect 0 561436 116 561476
rect 0 561416 96 561436
rect 0 560468 96 560488
rect 0 560428 116 560468
rect 0 560408 96 560428
rect 0 559460 96 559480
rect 0 559420 116 559460
rect 0 559400 96 559420
rect 0 558452 96 558472
rect 0 558412 116 558452
rect 0 558392 96 558412
rect 0 557444 96 557464
rect 0 557404 116 557444
rect 0 557384 96 557404
rect 452544 556940 452640 556960
rect 452524 556900 452640 556940
rect 452544 556880 452640 556900
rect 0 556436 96 556456
rect 452544 556436 452640 556456
rect 0 556396 116 556436
rect 452524 556396 452640 556436
rect 0 556376 96 556396
rect 452544 556376 452640 556396
rect 452544 555932 452640 555952
rect 452524 555892 452640 555932
rect 452544 555872 452640 555892
rect 0 555428 96 555448
rect 452544 555428 452640 555448
rect 0 555388 116 555428
rect 452524 555388 452640 555428
rect 0 555368 96 555388
rect 452544 555368 452640 555388
rect 452544 554924 452640 554944
rect 452524 554884 452640 554924
rect 452544 554864 452640 554884
rect 0 554420 96 554440
rect 452544 554420 452640 554440
rect 0 554380 116 554420
rect 452524 554380 452640 554420
rect 0 554360 96 554380
rect 452544 554360 452640 554380
rect 452544 553916 452640 553936
rect 452524 553876 452640 553916
rect 452544 553856 452640 553876
rect 0 553412 96 553432
rect 452544 553412 452640 553432
rect 0 553372 116 553412
rect 452524 553372 452640 553412
rect 0 553352 96 553372
rect 452544 553352 452640 553372
rect 452544 552908 452640 552928
rect 452524 552868 452640 552908
rect 452544 552848 452640 552868
rect 0 552404 96 552424
rect 452544 552404 452640 552424
rect 0 552364 116 552404
rect 452524 552364 452640 552404
rect 0 552344 96 552364
rect 452544 552344 452640 552364
rect 452544 551900 452640 551920
rect 452524 551860 452640 551900
rect 452544 551840 452640 551860
rect 0 551396 96 551416
rect 452544 551396 452640 551416
rect 0 551356 116 551396
rect 452524 551356 452640 551396
rect 0 551336 96 551356
rect 452544 551336 452640 551356
rect 452544 550892 452640 550912
rect 452524 550852 452640 550892
rect 452544 550832 452640 550852
rect 0 550388 96 550408
rect 452544 550388 452640 550408
rect 0 550348 116 550388
rect 452524 550348 452640 550388
rect 0 550328 96 550348
rect 452544 550328 452640 550348
rect 452544 549884 452640 549904
rect 452524 549844 452640 549884
rect 452544 549824 452640 549844
rect 0 549380 96 549400
rect 452544 549380 452640 549400
rect 0 549340 116 549380
rect 452524 549340 452640 549380
rect 0 549320 96 549340
rect 452544 549320 452640 549340
rect 452544 548876 452640 548896
rect 452524 548836 452640 548876
rect 452544 548816 452640 548836
rect 0 548372 96 548392
rect 452544 548372 452640 548392
rect 0 548332 116 548372
rect 452524 548332 452640 548372
rect 0 548312 96 548332
rect 452544 548312 452640 548332
rect 452544 547868 452640 547888
rect 452524 547828 452640 547868
rect 452544 547808 452640 547828
rect 0 547364 96 547384
rect 452544 547364 452640 547384
rect 0 547324 116 547364
rect 452524 547324 452640 547364
rect 0 547304 96 547324
rect 452544 547304 452640 547324
rect 452544 546860 452640 546880
rect 452524 546820 452640 546860
rect 452544 546800 452640 546820
rect 0 546356 96 546376
rect 452544 546356 452640 546376
rect 0 546316 116 546356
rect 452524 546316 452640 546356
rect 0 546296 96 546316
rect 452544 546296 452640 546316
rect 452544 545852 452640 545872
rect 452524 545812 452640 545852
rect 452544 545792 452640 545812
rect 452544 545348 452640 545368
rect 452524 545308 452640 545348
rect 452544 545288 452640 545308
rect 452544 544844 452640 544864
rect 452524 544804 452640 544844
rect 452544 544784 452640 544804
rect 452544 544340 452640 544360
rect 452524 544300 452640 544340
rect 452544 544280 452640 544300
rect 452544 543836 452640 543856
rect 452524 543796 452640 543836
rect 452544 543776 452640 543796
rect 0 543332 96 543352
rect 452544 543332 452640 543352
rect 0 543292 116 543332
rect 452524 543292 452640 543332
rect 0 543272 96 543292
rect 452544 543272 452640 543292
rect 452544 542828 452640 542848
rect 452524 542788 452640 542828
rect 452544 542768 452640 542788
rect 0 542324 96 542344
rect 452544 542324 452640 542344
rect 0 542284 116 542324
rect 452524 542284 452640 542324
rect 0 542264 96 542284
rect 452544 542264 452640 542284
rect 452544 541820 452640 541840
rect 452524 541780 452640 541820
rect 452544 541760 452640 541780
rect 0 541316 96 541336
rect 452544 541316 452640 541336
rect 0 541276 116 541316
rect 452524 541276 452640 541316
rect 0 541256 96 541276
rect 452544 541256 452640 541276
rect 452544 540812 452640 540832
rect 452524 540772 452640 540812
rect 452544 540752 452640 540772
rect 0 540308 96 540328
rect 452544 540308 452640 540328
rect 0 540268 116 540308
rect 452524 540268 452640 540308
rect 0 540248 96 540268
rect 452544 540248 452640 540268
rect 452544 539804 452640 539824
rect 452524 539764 452640 539804
rect 452544 539744 452640 539764
rect 0 539300 96 539320
rect 452544 539300 452640 539320
rect 0 539260 116 539300
rect 452524 539260 452640 539300
rect 0 539240 96 539260
rect 452544 539240 452640 539260
rect 452544 538796 452640 538816
rect 452524 538756 452640 538796
rect 452544 538736 452640 538756
rect 0 538292 96 538312
rect 452544 538292 452640 538312
rect 0 538252 116 538292
rect 452524 538252 452640 538292
rect 0 538232 96 538252
rect 452544 538232 452640 538252
rect 452544 537788 452640 537808
rect 452524 537748 452640 537788
rect 452544 537728 452640 537748
rect 0 537284 96 537304
rect 452544 537284 452640 537304
rect 0 537244 116 537284
rect 452524 537244 452640 537284
rect 0 537224 96 537244
rect 452544 537224 452640 537244
rect 452544 536780 452640 536800
rect 452524 536740 452640 536780
rect 452544 536720 452640 536740
rect 0 536276 96 536296
rect 452544 536276 452640 536296
rect 0 536236 116 536276
rect 452524 536236 452640 536276
rect 0 536216 96 536236
rect 452544 536216 452640 536236
rect 452544 535772 452640 535792
rect 452524 535732 452640 535772
rect 452544 535712 452640 535732
rect 0 535268 96 535288
rect 452544 535268 452640 535288
rect 0 535228 116 535268
rect 452524 535228 452640 535268
rect 0 535208 96 535228
rect 452544 535208 452640 535228
rect 452544 534764 452640 534784
rect 452524 534724 452640 534764
rect 452544 534704 452640 534724
rect 0 534260 96 534280
rect 452544 534260 452640 534280
rect 0 534220 116 534260
rect 452524 534220 452640 534260
rect 0 534200 96 534220
rect 452544 534200 452640 534220
rect 452544 533756 452640 533776
rect 452524 533716 452640 533756
rect 452544 533696 452640 533716
rect 0 533252 96 533272
rect 452544 533252 452640 533272
rect 0 533212 116 533252
rect 452524 533212 452640 533252
rect 0 533192 96 533212
rect 452544 533192 452640 533212
rect 452544 532748 452640 532768
rect 452524 532708 452640 532748
rect 452544 532688 452640 532708
rect 0 532244 96 532264
rect 452544 532244 452640 532264
rect 0 532204 116 532244
rect 452524 532204 452640 532244
rect 0 532184 96 532204
rect 452544 532184 452640 532204
rect 452544 531740 452640 531760
rect 452524 531700 452640 531740
rect 452544 531680 452640 531700
rect 0 531236 96 531256
rect 452544 531236 452640 531256
rect 0 531196 116 531236
rect 452524 531196 452640 531236
rect 0 531176 96 531196
rect 452544 531176 452640 531196
rect 452544 530732 452640 530752
rect 452524 530692 452640 530732
rect 452544 530672 452640 530692
rect 0 530228 96 530248
rect 452544 530228 452640 530248
rect 0 530188 116 530228
rect 452524 530188 452640 530228
rect 0 530168 96 530188
rect 452544 530168 452640 530188
rect 452544 529724 452640 529744
rect 452524 529684 452640 529724
rect 452544 529664 452640 529684
rect 0 529220 96 529240
rect 452544 529220 452640 529240
rect 0 529180 116 529220
rect 452524 529180 452640 529220
rect 0 529160 96 529180
rect 452544 529160 452640 529180
rect 452544 528716 452640 528736
rect 452524 528676 452640 528716
rect 452544 528656 452640 528676
rect 0 528212 96 528232
rect 452544 528212 452640 528232
rect 0 528172 116 528212
rect 452524 528172 452640 528212
rect 0 528152 96 528172
rect 452544 528152 452640 528172
rect 452544 527708 452640 527728
rect 452524 527668 452640 527708
rect 452544 527648 452640 527668
rect 0 527204 96 527224
rect 452544 527204 452640 527224
rect 0 527164 116 527204
rect 452524 527164 452640 527204
rect 0 527144 96 527164
rect 452544 527144 452640 527164
rect 452544 526700 452640 526720
rect 452524 526660 452640 526700
rect 452544 526640 452640 526660
rect 0 526196 96 526216
rect 452544 526196 452640 526216
rect 0 526156 116 526196
rect 452524 526156 452640 526196
rect 0 526136 96 526156
rect 452544 526136 452640 526156
rect 452544 525692 452640 525712
rect 452524 525652 452640 525692
rect 452544 525632 452640 525652
rect 0 525188 96 525208
rect 452544 525188 452640 525208
rect 0 525148 116 525188
rect 452524 525148 452640 525188
rect 0 525128 96 525148
rect 452544 525128 452640 525148
rect 452544 524684 452640 524704
rect 452524 524644 452640 524684
rect 452544 524624 452640 524644
rect 0 524180 96 524200
rect 452544 524180 452640 524200
rect 0 524140 116 524180
rect 452524 524140 452640 524180
rect 0 524120 96 524140
rect 452544 524120 452640 524140
rect 452544 523676 452640 523696
rect 452524 523636 452640 523676
rect 452544 523616 452640 523636
rect 0 523172 96 523192
rect 452544 523172 452640 523192
rect 0 523132 116 523172
rect 452524 523132 452640 523172
rect 0 523112 96 523132
rect 452544 523112 452640 523132
rect 452544 522668 452640 522688
rect 452524 522628 452640 522668
rect 452544 522608 452640 522628
rect 0 522164 96 522184
rect 452544 522164 452640 522184
rect 0 522124 116 522164
rect 452524 522124 452640 522164
rect 0 522104 96 522124
rect 452544 522104 452640 522124
rect 452544 521660 452640 521680
rect 452524 521620 452640 521660
rect 452544 521600 452640 521620
rect 0 521156 96 521176
rect 452544 521156 452640 521176
rect 0 521116 116 521156
rect 452524 521116 452640 521156
rect 0 521096 96 521116
rect 452544 521096 452640 521116
rect 452544 520652 452640 520672
rect 452524 520612 452640 520652
rect 452544 520592 452640 520612
rect 0 520148 96 520168
rect 452544 520148 452640 520168
rect 0 520108 116 520148
rect 452524 520108 452640 520148
rect 0 520088 96 520108
rect 452544 520088 452640 520108
rect 452544 519644 452640 519664
rect 452524 519604 452640 519644
rect 452544 519584 452640 519604
rect 0 519140 96 519160
rect 452544 519140 452640 519160
rect 0 519100 116 519140
rect 452524 519100 452640 519140
rect 0 519080 96 519100
rect 452544 519080 452640 519100
rect 452544 518636 452640 518656
rect 452524 518596 452640 518636
rect 452544 518576 452640 518596
rect 0 518132 96 518152
rect 452544 518132 452640 518152
rect 0 518092 116 518132
rect 452524 518092 452640 518132
rect 0 518072 96 518092
rect 452544 518072 452640 518092
rect 452544 517628 452640 517648
rect 452524 517588 452640 517628
rect 452544 517568 452640 517588
rect 0 517124 96 517144
rect 452544 517124 452640 517144
rect 0 517084 116 517124
rect 452524 517084 452640 517124
rect 0 517064 96 517084
rect 452544 517064 452640 517084
rect 452544 516620 452640 516640
rect 452524 516580 452640 516620
rect 452544 516560 452640 516580
rect 0 516116 96 516136
rect 452544 516116 452640 516136
rect 0 516076 116 516116
rect 452524 516076 452640 516116
rect 0 516056 96 516076
rect 452544 516056 452640 516076
rect 452544 515612 452640 515632
rect 452524 515572 452640 515612
rect 452544 515552 452640 515572
rect 0 515108 96 515128
rect 452544 515108 452640 515128
rect 0 515068 116 515108
rect 452524 515068 452640 515108
rect 0 515048 96 515068
rect 452544 515048 452640 515068
rect 452544 514604 452640 514624
rect 452524 514564 452640 514604
rect 452544 514544 452640 514564
rect 0 514100 96 514120
rect 452544 514100 452640 514120
rect 0 514060 116 514100
rect 452524 514060 452640 514100
rect 0 514040 96 514060
rect 452544 514040 452640 514060
rect 452544 513596 452640 513616
rect 452524 513556 452640 513596
rect 452544 513536 452640 513556
rect 0 513092 96 513112
rect 452544 513092 452640 513112
rect 0 513052 116 513092
rect 452524 513052 452640 513092
rect 0 513032 96 513052
rect 452544 513032 452640 513052
rect 452544 512588 452640 512608
rect 452524 512548 452640 512588
rect 452544 512528 452640 512548
rect 0 512084 96 512104
rect 452544 512084 452640 512104
rect 0 512044 116 512084
rect 452524 512044 452640 512084
rect 0 512024 96 512044
rect 452544 512024 452640 512044
rect 452544 511580 452640 511600
rect 452524 511540 452640 511580
rect 452544 511520 452640 511540
rect 0 511076 96 511096
rect 452544 511076 452640 511096
rect 0 511036 116 511076
rect 452524 511036 452640 511076
rect 0 511016 96 511036
rect 452544 511016 452640 511036
rect 452544 510572 452640 510592
rect 452524 510532 452640 510572
rect 452544 510512 452640 510532
rect 0 510068 96 510088
rect 452544 510068 452640 510088
rect 0 510028 116 510068
rect 452524 510028 452640 510068
rect 0 510008 96 510028
rect 452544 510008 452640 510028
rect 452544 509564 452640 509584
rect 452524 509524 452640 509564
rect 452544 509504 452640 509524
rect 0 509060 96 509080
rect 452544 509060 452640 509080
rect 0 509020 116 509060
rect 452524 509020 452640 509060
rect 0 509000 96 509020
rect 452544 509000 452640 509020
rect 452544 508556 452640 508576
rect 452524 508516 452640 508556
rect 452544 508496 452640 508516
rect 0 508052 96 508072
rect 452544 508052 452640 508072
rect 0 508012 116 508052
rect 452524 508012 452640 508052
rect 0 507992 96 508012
rect 452544 507992 452640 508012
rect 452544 507548 452640 507568
rect 452524 507508 452640 507548
rect 452544 507488 452640 507508
rect 0 507044 96 507064
rect 452544 507044 452640 507064
rect 0 507004 116 507044
rect 452524 507004 452640 507044
rect 0 506984 96 507004
rect 452544 506984 452640 507004
rect 452544 506540 452640 506560
rect 452524 506500 452640 506540
rect 452544 506480 452640 506500
rect 0 506036 96 506056
rect 452544 506036 452640 506056
rect 0 505996 116 506036
rect 452524 505996 452640 506036
rect 0 505976 96 505996
rect 452544 505976 452640 505996
rect 452544 505532 452640 505552
rect 452524 505492 452640 505532
rect 452544 505472 452640 505492
rect 0 505028 96 505048
rect 452544 505028 452640 505048
rect 0 504988 116 505028
rect 452524 504988 452640 505028
rect 0 504968 96 504988
rect 452544 504968 452640 504988
rect 452544 504524 452640 504544
rect 452524 504484 452640 504524
rect 452544 504464 452640 504484
rect 0 504020 96 504040
rect 452544 504020 452640 504040
rect 0 503980 116 504020
rect 452524 503980 452640 504020
rect 0 503960 96 503980
rect 452544 503960 452640 503980
rect 452544 503516 452640 503536
rect 452524 503476 452640 503516
rect 452544 503456 452640 503476
rect 0 503012 96 503032
rect 452544 503012 452640 503032
rect 0 502972 116 503012
rect 452524 502972 452640 503012
rect 0 502952 96 502972
rect 452544 502952 452640 502972
rect 452544 502508 452640 502528
rect 452524 502468 452640 502508
rect 452544 502448 452640 502468
rect 0 502004 96 502024
rect 452544 502004 452640 502024
rect 0 501964 116 502004
rect 452524 501964 452640 502004
rect 0 501944 96 501964
rect 452544 501944 452640 501964
rect 452544 501500 452640 501520
rect 452524 501460 452640 501500
rect 452544 501440 452640 501460
rect 0 500996 96 501016
rect 452544 500996 452640 501016
rect 0 500956 116 500996
rect 452524 500956 452640 500996
rect 0 500936 96 500956
rect 452544 500936 452640 500956
rect 452544 500492 452640 500512
rect 452524 500452 452640 500492
rect 452544 500432 452640 500452
rect 0 499988 96 500008
rect 0 499948 116 499988
rect 0 499928 96 499948
rect 0 498980 96 499000
rect 0 498940 116 498980
rect 0 498920 96 498940
rect 0 497972 96 497992
rect 0 497932 116 497972
rect 0 497912 96 497932
rect 0 494948 96 494968
rect 0 494908 116 494948
rect 0 494888 96 494908
rect 0 493940 96 493960
rect 0 493900 116 493940
rect 0 493880 96 493900
rect 0 492932 96 492952
rect 0 492892 116 492932
rect 0 492872 96 492892
rect 0 491924 96 491944
rect 0 491884 116 491924
rect 0 491864 96 491884
rect 0 490916 96 490936
rect 0 490876 116 490916
rect 0 490856 96 490876
rect 0 489908 96 489928
rect 0 489868 116 489908
rect 0 489848 96 489868
rect 0 488900 96 488920
rect 0 488860 116 488900
rect 0 488840 96 488860
rect 0 487892 96 487912
rect 0 487852 116 487892
rect 0 487832 96 487852
rect 0 486884 96 486904
rect 0 486844 116 486884
rect 0 486824 96 486844
rect 0 485876 96 485896
rect 0 485836 116 485876
rect 0 485816 96 485836
rect 0 484868 96 484888
rect 0 484828 116 484868
rect 0 484808 96 484828
rect 0 483860 96 483880
rect 0 483820 116 483860
rect 0 483800 96 483820
rect 0 482852 96 482872
rect 0 482812 116 482852
rect 0 482792 96 482812
rect 0 481844 96 481864
rect 0 481804 116 481844
rect 0 481784 96 481804
rect 0 480836 96 480856
rect 0 480796 116 480836
rect 0 480776 96 480796
rect 0 479828 96 479848
rect 0 479788 116 479828
rect 0 479768 96 479788
rect 0 478820 96 478840
rect 0 478780 116 478820
rect 0 478760 96 478780
rect 0 477812 96 477832
rect 0 477772 116 477812
rect 0 477752 96 477772
rect 0 476804 96 476824
rect 0 476764 116 476804
rect 0 476744 96 476764
rect 0 475796 96 475816
rect 0 475756 116 475796
rect 0 475736 96 475756
rect 0 474788 96 474808
rect 0 474748 116 474788
rect 0 474728 96 474748
rect 0 473780 96 473800
rect 0 473740 116 473780
rect 0 473720 96 473740
rect 0 472772 96 472792
rect 0 472732 116 472772
rect 0 472712 96 472732
rect 0 471764 96 471784
rect 0 471724 116 471764
rect 0 471704 96 471724
rect 0 470756 96 470776
rect 0 470716 116 470756
rect 0 470696 96 470716
rect 0 469748 96 469768
rect 0 469708 116 469748
rect 0 469688 96 469708
rect 0 468740 96 468760
rect 0 468700 116 468740
rect 0 468680 96 468700
rect 0 467732 96 467752
rect 0 467692 116 467732
rect 0 467672 96 467692
rect 0 466724 96 466744
rect 0 466684 116 466724
rect 0 466664 96 466684
rect 0 465716 96 465736
rect 0 465676 116 465716
rect 0 465656 96 465676
rect 0 464708 96 464728
rect 0 464668 116 464708
rect 0 464648 96 464668
rect 0 463700 96 463720
rect 0 463660 116 463700
rect 0 463640 96 463660
rect 0 462692 96 462712
rect 0 462652 116 462692
rect 0 462632 96 462652
rect 0 461684 96 461704
rect 0 461644 116 461684
rect 0 461624 96 461644
rect 0 460676 96 460696
rect 0 460636 116 460676
rect 0 460616 96 460636
rect 452544 460172 452640 460192
rect 452524 460132 452640 460172
rect 452544 460112 452640 460132
rect 0 459668 96 459688
rect 452544 459668 452640 459688
rect 0 459628 116 459668
rect 452524 459628 452640 459668
rect 0 459608 96 459628
rect 452544 459608 452640 459628
rect 452544 459164 452640 459184
rect 452524 459124 452640 459164
rect 452544 459104 452640 459124
rect 0 458660 96 458680
rect 452544 458660 452640 458680
rect 0 458620 116 458660
rect 452524 458620 452640 458660
rect 0 458600 96 458620
rect 452544 458600 452640 458620
rect 452544 458156 452640 458176
rect 452524 458116 452640 458156
rect 452544 458096 452640 458116
rect 0 457652 96 457672
rect 452544 457652 452640 457672
rect 0 457612 116 457652
rect 452524 457612 452640 457652
rect 0 457592 96 457612
rect 452544 457592 452640 457612
rect 452544 457148 452640 457168
rect 452524 457108 452640 457148
rect 452544 457088 452640 457108
rect 0 456644 96 456664
rect 452544 456644 452640 456664
rect 0 456604 116 456644
rect 452524 456604 452640 456644
rect 0 456584 96 456604
rect 452544 456584 452640 456604
rect 452544 456140 452640 456160
rect 452524 456100 452640 456140
rect 452544 456080 452640 456100
rect 0 455636 96 455656
rect 452544 455636 452640 455656
rect 0 455596 116 455636
rect 452524 455596 452640 455636
rect 0 455576 96 455596
rect 452544 455576 452640 455596
rect 452544 455132 452640 455152
rect 452524 455092 452640 455132
rect 452544 455072 452640 455092
rect 0 454628 96 454648
rect 452544 454628 452640 454648
rect 0 454588 116 454628
rect 452524 454588 452640 454628
rect 0 454568 96 454588
rect 452544 454568 452640 454588
rect 452544 454124 452640 454144
rect 452524 454084 452640 454124
rect 452544 454064 452640 454084
rect 0 453620 96 453640
rect 452544 453620 452640 453640
rect 0 453580 116 453620
rect 452524 453580 452640 453620
rect 0 453560 96 453580
rect 452544 453560 452640 453580
rect 452544 453116 452640 453136
rect 452524 453076 452640 453116
rect 452544 453056 452640 453076
rect 0 452612 96 452632
rect 452544 452612 452640 452632
rect 0 452572 116 452612
rect 452524 452572 452640 452612
rect 0 452552 96 452572
rect 452544 452552 452640 452572
rect 452544 452108 452640 452128
rect 452524 452068 452640 452108
rect 452544 452048 452640 452068
rect 0 451604 96 451624
rect 452544 451604 452640 451624
rect 0 451564 116 451604
rect 452524 451564 452640 451604
rect 0 451544 96 451564
rect 452544 451544 452640 451564
rect 452544 451100 452640 451120
rect 452524 451060 452640 451100
rect 452544 451040 452640 451060
rect 0 450596 96 450616
rect 452544 450596 452640 450616
rect 0 450556 116 450596
rect 452524 450556 452640 450596
rect 0 450536 96 450556
rect 452544 450536 452640 450556
rect 452544 450092 452640 450112
rect 452524 450052 452640 450092
rect 452544 450032 452640 450052
rect 0 449588 96 449608
rect 452544 449588 452640 449608
rect 0 449548 116 449588
rect 452524 449548 452640 449588
rect 0 449528 96 449548
rect 452544 449528 452640 449548
rect 452544 449084 452640 449104
rect 452524 449044 452640 449084
rect 452544 449024 452640 449044
rect 452544 448580 452640 448600
rect 452524 448540 452640 448580
rect 452544 448520 452640 448540
rect 452544 448076 452640 448096
rect 452524 448036 452640 448076
rect 452544 448016 452640 448036
rect 452544 447572 452640 447592
rect 452524 447532 452640 447572
rect 452544 447512 452640 447532
rect 452544 447068 452640 447088
rect 452524 447028 452640 447068
rect 452544 447008 452640 447028
rect 0 446564 96 446584
rect 452544 446564 452640 446584
rect 0 446524 116 446564
rect 452524 446524 452640 446564
rect 0 446504 96 446524
rect 452544 446504 452640 446524
rect 452544 446060 452640 446080
rect 452524 446020 452640 446060
rect 452544 446000 452640 446020
rect 0 445556 96 445576
rect 452544 445556 452640 445576
rect 0 445516 116 445556
rect 452524 445516 452640 445556
rect 0 445496 96 445516
rect 452544 445496 452640 445516
rect 452544 445052 452640 445072
rect 452524 445012 452640 445052
rect 452544 444992 452640 445012
rect 0 444548 96 444568
rect 452544 444548 452640 444568
rect 0 444508 116 444548
rect 452524 444508 452640 444548
rect 0 444488 96 444508
rect 452544 444488 452640 444508
rect 452544 444044 452640 444064
rect 452524 444004 452640 444044
rect 452544 443984 452640 444004
rect 0 443540 96 443560
rect 452544 443540 452640 443560
rect 0 443500 116 443540
rect 452524 443500 452640 443540
rect 0 443480 96 443500
rect 452544 443480 452640 443500
rect 452544 443036 452640 443056
rect 452524 442996 452640 443036
rect 452544 442976 452640 442996
rect 0 442532 96 442552
rect 452544 442532 452640 442552
rect 0 442492 116 442532
rect 452524 442492 452640 442532
rect 0 442472 96 442492
rect 452544 442472 452640 442492
rect 452544 442028 452640 442048
rect 452524 441988 452640 442028
rect 452544 441968 452640 441988
rect 0 441524 96 441544
rect 452544 441524 452640 441544
rect 0 441484 116 441524
rect 452524 441484 452640 441524
rect 0 441464 96 441484
rect 452544 441464 452640 441484
rect 452544 441020 452640 441040
rect 452524 440980 452640 441020
rect 452544 440960 452640 440980
rect 0 440516 96 440536
rect 452544 440516 452640 440536
rect 0 440476 116 440516
rect 452524 440476 452640 440516
rect 0 440456 96 440476
rect 452544 440456 452640 440476
rect 452544 440012 452640 440032
rect 452524 439972 452640 440012
rect 452544 439952 452640 439972
rect 0 439508 96 439528
rect 452544 439508 452640 439528
rect 0 439468 116 439508
rect 452524 439468 452640 439508
rect 0 439448 96 439468
rect 452544 439448 452640 439468
rect 452544 439004 452640 439024
rect 452524 438964 452640 439004
rect 452544 438944 452640 438964
rect 0 438500 96 438520
rect 452544 438500 452640 438520
rect 0 438460 116 438500
rect 452524 438460 452640 438500
rect 0 438440 96 438460
rect 452544 438440 452640 438460
rect 452544 437996 452640 438016
rect 452524 437956 452640 437996
rect 452544 437936 452640 437956
rect 0 437492 96 437512
rect 452544 437492 452640 437512
rect 0 437452 116 437492
rect 452524 437452 452640 437492
rect 0 437432 96 437452
rect 452544 437432 452640 437452
rect 452544 436988 452640 437008
rect 452524 436948 452640 436988
rect 452544 436928 452640 436948
rect 0 436484 96 436504
rect 452544 436484 452640 436504
rect 0 436444 116 436484
rect 452524 436444 452640 436484
rect 0 436424 96 436444
rect 452544 436424 452640 436444
rect 452544 435980 452640 436000
rect 452524 435940 452640 435980
rect 452544 435920 452640 435940
rect 0 435476 96 435496
rect 452544 435476 452640 435496
rect 0 435436 116 435476
rect 452524 435436 452640 435476
rect 0 435416 96 435436
rect 452544 435416 452640 435436
rect 452544 434972 452640 434992
rect 452524 434932 452640 434972
rect 452544 434912 452640 434932
rect 0 434468 96 434488
rect 452544 434468 452640 434488
rect 0 434428 116 434468
rect 452524 434428 452640 434468
rect 0 434408 96 434428
rect 452544 434408 452640 434428
rect 452544 433964 452640 433984
rect 452524 433924 452640 433964
rect 452544 433904 452640 433924
rect 0 433460 96 433480
rect 452544 433460 452640 433480
rect 0 433420 116 433460
rect 452524 433420 452640 433460
rect 0 433400 96 433420
rect 452544 433400 452640 433420
rect 452544 432956 452640 432976
rect 452524 432916 452640 432956
rect 452544 432896 452640 432916
rect 0 432452 96 432472
rect 452544 432452 452640 432472
rect 0 432412 116 432452
rect 452524 432412 452640 432452
rect 0 432392 96 432412
rect 452544 432392 452640 432412
rect 452544 431948 452640 431968
rect 452524 431908 452640 431948
rect 452544 431888 452640 431908
rect 0 431444 96 431464
rect 452544 431444 452640 431464
rect 0 431404 116 431444
rect 452524 431404 452640 431444
rect 0 431384 96 431404
rect 452544 431384 452640 431404
rect 452544 430940 452640 430960
rect 452524 430900 452640 430940
rect 452544 430880 452640 430900
rect 0 430436 96 430456
rect 452544 430436 452640 430456
rect 0 430396 116 430436
rect 452524 430396 452640 430436
rect 0 430376 96 430396
rect 452544 430376 452640 430396
rect 452544 429932 452640 429952
rect 452524 429892 452640 429932
rect 452544 429872 452640 429892
rect 0 429428 96 429448
rect 452544 429428 452640 429448
rect 0 429388 116 429428
rect 452524 429388 452640 429428
rect 0 429368 96 429388
rect 452544 429368 452640 429388
rect 452544 428924 452640 428944
rect 452524 428884 452640 428924
rect 452544 428864 452640 428884
rect 0 428420 96 428440
rect 452544 428420 452640 428440
rect 0 428380 116 428420
rect 452524 428380 452640 428420
rect 0 428360 96 428380
rect 452544 428360 452640 428380
rect 452544 427916 452640 427936
rect 452524 427876 452640 427916
rect 452544 427856 452640 427876
rect 0 427412 96 427432
rect 452544 427412 452640 427432
rect 0 427372 116 427412
rect 452524 427372 452640 427412
rect 0 427352 96 427372
rect 452544 427352 452640 427372
rect 452544 426908 452640 426928
rect 452524 426868 452640 426908
rect 452544 426848 452640 426868
rect 0 426404 96 426424
rect 452544 426404 452640 426424
rect 0 426364 116 426404
rect 452524 426364 452640 426404
rect 0 426344 96 426364
rect 452544 426344 452640 426364
rect 452544 425900 452640 425920
rect 452524 425860 452640 425900
rect 452544 425840 452640 425860
rect 0 425396 96 425416
rect 452544 425396 452640 425416
rect 0 425356 116 425396
rect 452524 425356 452640 425396
rect 0 425336 96 425356
rect 452544 425336 452640 425356
rect 452544 424892 452640 424912
rect 452524 424852 452640 424892
rect 452544 424832 452640 424852
rect 0 424388 96 424408
rect 452544 424388 452640 424408
rect 0 424348 116 424388
rect 452524 424348 452640 424388
rect 0 424328 96 424348
rect 452544 424328 452640 424348
rect 452544 423884 452640 423904
rect 452524 423844 452640 423884
rect 452544 423824 452640 423844
rect 0 423380 96 423400
rect 452544 423380 452640 423400
rect 0 423340 116 423380
rect 452524 423340 452640 423380
rect 0 423320 96 423340
rect 452544 423320 452640 423340
rect 452544 422876 452640 422896
rect 452524 422836 452640 422876
rect 452544 422816 452640 422836
rect 0 422372 96 422392
rect 452544 422372 452640 422392
rect 0 422332 116 422372
rect 452524 422332 452640 422372
rect 0 422312 96 422332
rect 452544 422312 452640 422332
rect 452544 421868 452640 421888
rect 452524 421828 452640 421868
rect 452544 421808 452640 421828
rect 0 421364 96 421384
rect 452544 421364 452640 421384
rect 0 421324 116 421364
rect 452524 421324 452640 421364
rect 0 421304 96 421324
rect 452544 421304 452640 421324
rect 452544 420860 452640 420880
rect 452524 420820 452640 420860
rect 452544 420800 452640 420820
rect 0 420356 96 420376
rect 452544 420356 452640 420376
rect 0 420316 116 420356
rect 452524 420316 452640 420356
rect 0 420296 96 420316
rect 452544 420296 452640 420316
rect 452544 419852 452640 419872
rect 452524 419812 452640 419852
rect 452544 419792 452640 419812
rect 0 419348 96 419368
rect 452544 419348 452640 419368
rect 0 419308 116 419348
rect 452524 419308 452640 419348
rect 0 419288 96 419308
rect 452544 419288 452640 419308
rect 452544 418844 452640 418864
rect 452524 418804 452640 418844
rect 452544 418784 452640 418804
rect 0 418340 96 418360
rect 452544 418340 452640 418360
rect 0 418300 116 418340
rect 452524 418300 452640 418340
rect 0 418280 96 418300
rect 452544 418280 452640 418300
rect 452544 417836 452640 417856
rect 452524 417796 452640 417836
rect 452544 417776 452640 417796
rect 0 417332 96 417352
rect 452544 417332 452640 417352
rect 0 417292 116 417332
rect 452524 417292 452640 417332
rect 0 417272 96 417292
rect 452544 417272 452640 417292
rect 452544 416828 452640 416848
rect 452524 416788 452640 416828
rect 452544 416768 452640 416788
rect 0 416324 96 416344
rect 452544 416324 452640 416344
rect 0 416284 116 416324
rect 452524 416284 452640 416324
rect 0 416264 96 416284
rect 452544 416264 452640 416284
rect 452544 415820 452640 415840
rect 452524 415780 452640 415820
rect 452544 415760 452640 415780
rect 0 415316 96 415336
rect 452544 415316 452640 415336
rect 0 415276 116 415316
rect 452524 415276 452640 415316
rect 0 415256 96 415276
rect 452544 415256 452640 415276
rect 452544 414812 452640 414832
rect 452524 414772 452640 414812
rect 452544 414752 452640 414772
rect 0 414308 96 414328
rect 452544 414308 452640 414328
rect 0 414268 116 414308
rect 452524 414268 452640 414308
rect 0 414248 96 414268
rect 452544 414248 452640 414268
rect 452544 413804 452640 413824
rect 452524 413764 452640 413804
rect 452544 413744 452640 413764
rect 0 413300 96 413320
rect 452544 413300 452640 413320
rect 0 413260 116 413300
rect 452524 413260 452640 413300
rect 0 413240 96 413260
rect 452544 413240 452640 413260
rect 452544 412796 452640 412816
rect 452524 412756 452640 412796
rect 452544 412736 452640 412756
rect 0 412292 96 412312
rect 452544 412292 452640 412312
rect 0 412252 116 412292
rect 452524 412252 452640 412292
rect 0 412232 96 412252
rect 452544 412232 452640 412252
rect 452544 411788 452640 411808
rect 452524 411748 452640 411788
rect 452544 411728 452640 411748
rect 0 411284 96 411304
rect 452544 411284 452640 411304
rect 0 411244 116 411284
rect 452524 411244 452640 411284
rect 0 411224 96 411244
rect 452544 411224 452640 411244
rect 452544 410780 452640 410800
rect 452524 410740 452640 410780
rect 452544 410720 452640 410740
rect 0 410276 96 410296
rect 452544 410276 452640 410296
rect 0 410236 116 410276
rect 452524 410236 452640 410276
rect 0 410216 96 410236
rect 452544 410216 452640 410236
rect 452544 409772 452640 409792
rect 452524 409732 452640 409772
rect 452544 409712 452640 409732
rect 0 409268 96 409288
rect 452544 409268 452640 409288
rect 0 409228 116 409268
rect 452524 409228 452640 409268
rect 0 409208 96 409228
rect 452544 409208 452640 409228
rect 452544 408764 452640 408784
rect 452524 408724 452640 408764
rect 452544 408704 452640 408724
rect 0 408260 96 408280
rect 452544 408260 452640 408280
rect 0 408220 116 408260
rect 452524 408220 452640 408260
rect 0 408200 96 408220
rect 452544 408200 452640 408220
rect 452544 407756 452640 407776
rect 452524 407716 452640 407756
rect 452544 407696 452640 407716
rect 0 407252 96 407272
rect 452544 407252 452640 407272
rect 0 407212 116 407252
rect 452524 407212 452640 407252
rect 0 407192 96 407212
rect 452544 407192 452640 407212
rect 452544 406748 452640 406768
rect 452524 406708 452640 406748
rect 452544 406688 452640 406708
rect 0 406244 96 406264
rect 452544 406244 452640 406264
rect 0 406204 116 406244
rect 452524 406204 452640 406244
rect 0 406184 96 406204
rect 452544 406184 452640 406204
rect 452544 405740 452640 405760
rect 452524 405700 452640 405740
rect 452544 405680 452640 405700
rect 0 405236 96 405256
rect 452544 405236 452640 405256
rect 0 405196 116 405236
rect 452524 405196 452640 405236
rect 0 405176 96 405196
rect 452544 405176 452640 405196
rect 452544 404732 452640 404752
rect 452524 404692 452640 404732
rect 452544 404672 452640 404692
rect 0 404228 96 404248
rect 452544 404228 452640 404248
rect 0 404188 116 404228
rect 452524 404188 452640 404228
rect 0 404168 96 404188
rect 452544 404168 452640 404188
rect 452544 403724 452640 403744
rect 452524 403684 452640 403724
rect 452544 403664 452640 403684
rect 0 403220 96 403240
rect 0 403180 116 403220
rect 0 403160 96 403180
rect 0 402212 96 402232
rect 0 402172 116 402212
rect 0 402152 96 402172
rect 0 401204 96 401224
rect 0 401164 116 401204
rect 0 401144 96 401164
rect 0 398180 96 398200
rect 0 398140 116 398180
rect 0 398120 96 398140
rect 0 397172 96 397192
rect 0 397132 116 397172
rect 0 397112 96 397132
rect 0 396164 96 396184
rect 0 396124 116 396164
rect 0 396104 96 396124
rect 0 395156 96 395176
rect 0 395116 116 395156
rect 0 395096 96 395116
rect 0 394148 96 394168
rect 0 394108 116 394148
rect 0 394088 96 394108
rect 0 393140 96 393160
rect 0 393100 116 393140
rect 0 393080 96 393100
rect 0 392132 96 392152
rect 0 392092 116 392132
rect 0 392072 96 392092
rect 0 391124 96 391144
rect 0 391084 116 391124
rect 0 391064 96 391084
rect 0 390116 96 390136
rect 0 390076 116 390116
rect 0 390056 96 390076
rect 0 389108 96 389128
rect 0 389068 116 389108
rect 0 389048 96 389068
rect 0 388100 96 388120
rect 0 388060 116 388100
rect 0 388040 96 388060
rect 0 387092 96 387112
rect 0 387052 116 387092
rect 0 387032 96 387052
rect 0 386084 96 386104
rect 0 386044 116 386084
rect 0 386024 96 386044
rect 0 385076 96 385096
rect 0 385036 116 385076
rect 0 385016 96 385036
rect 0 384068 96 384088
rect 0 384028 116 384068
rect 0 384008 96 384028
rect 0 383060 96 383080
rect 0 383020 116 383060
rect 0 383000 96 383020
rect 0 382052 96 382072
rect 0 382012 116 382052
rect 0 381992 96 382012
rect 0 381044 96 381064
rect 0 381004 116 381044
rect 0 380984 96 381004
rect 0 380036 96 380056
rect 0 379996 116 380036
rect 0 379976 96 379996
rect 0 379028 96 379048
rect 0 378988 116 379028
rect 0 378968 96 378988
rect 0 378020 96 378040
rect 0 377980 116 378020
rect 0 377960 96 377980
rect 0 377012 96 377032
rect 0 376972 116 377012
rect 0 376952 96 376972
rect 0 376004 96 376024
rect 0 375964 116 376004
rect 0 375944 96 375964
rect 0 374996 96 375016
rect 0 374956 116 374996
rect 0 374936 96 374956
rect 0 373988 96 374008
rect 0 373948 116 373988
rect 0 373928 96 373948
rect 0 372980 96 373000
rect 0 372940 116 372980
rect 0 372920 96 372940
rect 0 371972 96 371992
rect 0 371932 116 371972
rect 0 371912 96 371932
rect 0 370964 96 370984
rect 0 370924 116 370964
rect 0 370904 96 370924
rect 0 369956 96 369976
rect 0 369916 116 369956
rect 0 369896 96 369916
rect 0 368948 96 368968
rect 0 368908 116 368948
rect 0 368888 96 368908
rect 0 367940 96 367960
rect 0 367900 116 367940
rect 0 367880 96 367900
rect 0 366932 96 366952
rect 0 366892 116 366932
rect 0 366872 96 366892
rect 0 365924 96 365944
rect 0 365884 116 365924
rect 0 365864 96 365884
rect 0 364916 96 364936
rect 0 364876 116 364916
rect 0 364856 96 364876
rect 0 363908 96 363928
rect 0 363868 116 363908
rect 0 363848 96 363868
rect 452544 363404 452640 363424
rect 452524 363364 452640 363404
rect 452544 363344 452640 363364
rect 0 362900 96 362920
rect 452544 362900 452640 362920
rect 0 362860 116 362900
rect 452524 362860 452640 362900
rect 0 362840 96 362860
rect 452544 362840 452640 362860
rect 452544 362396 452640 362416
rect 452524 362356 452640 362396
rect 452544 362336 452640 362356
rect 0 361892 96 361912
rect 452544 361892 452640 361912
rect 0 361852 116 361892
rect 452524 361852 452640 361892
rect 0 361832 96 361852
rect 452544 361832 452640 361852
rect 452544 361388 452640 361408
rect 452524 361348 452640 361388
rect 452544 361328 452640 361348
rect 0 360884 96 360904
rect 452544 360884 452640 360904
rect 0 360844 116 360884
rect 452524 360844 452640 360884
rect 0 360824 96 360844
rect 452544 360824 452640 360844
rect 452544 360380 452640 360400
rect 452524 360340 452640 360380
rect 452544 360320 452640 360340
rect 0 359876 96 359896
rect 452544 359876 452640 359896
rect 0 359836 116 359876
rect 452524 359836 452640 359876
rect 0 359816 96 359836
rect 452544 359816 452640 359836
rect 452544 359372 452640 359392
rect 452524 359332 452640 359372
rect 452544 359312 452640 359332
rect 0 358868 96 358888
rect 452544 358868 452640 358888
rect 0 358828 116 358868
rect 452524 358828 452640 358868
rect 0 358808 96 358828
rect 452544 358808 452640 358828
rect 452544 358364 452640 358384
rect 452524 358324 452640 358364
rect 452544 358304 452640 358324
rect 0 357860 96 357880
rect 452544 357860 452640 357880
rect 0 357820 116 357860
rect 452524 357820 452640 357860
rect 0 357800 96 357820
rect 452544 357800 452640 357820
rect 452544 357356 452640 357376
rect 452524 357316 452640 357356
rect 452544 357296 452640 357316
rect 0 356852 96 356872
rect 452544 356852 452640 356872
rect 0 356812 116 356852
rect 452524 356812 452640 356852
rect 0 356792 96 356812
rect 452544 356792 452640 356812
rect 452544 356348 452640 356368
rect 452524 356308 452640 356348
rect 452544 356288 452640 356308
rect 0 355844 96 355864
rect 452544 355844 452640 355864
rect 0 355804 116 355844
rect 452524 355804 452640 355844
rect 0 355784 96 355804
rect 452544 355784 452640 355804
rect 452544 355340 452640 355360
rect 452524 355300 452640 355340
rect 452544 355280 452640 355300
rect 0 354836 96 354856
rect 452544 354836 452640 354856
rect 0 354796 116 354836
rect 452524 354796 452640 354836
rect 0 354776 96 354796
rect 452544 354776 452640 354796
rect 452544 354332 452640 354352
rect 452524 354292 452640 354332
rect 452544 354272 452640 354292
rect 0 353828 96 353848
rect 452544 353828 452640 353848
rect 0 353788 116 353828
rect 452524 353788 452640 353828
rect 0 353768 96 353788
rect 452544 353768 452640 353788
rect 452544 353324 452640 353344
rect 452524 353284 452640 353324
rect 452544 353264 452640 353284
rect 0 352820 96 352840
rect 452544 352820 452640 352840
rect 0 352780 116 352820
rect 452524 352780 452640 352820
rect 0 352760 96 352780
rect 452544 352760 452640 352780
rect 452544 352316 452640 352336
rect 452524 352276 452640 352316
rect 452544 352256 452640 352276
rect 452544 351812 452640 351832
rect 452524 351772 452640 351812
rect 452544 351752 452640 351772
rect 452544 351308 452640 351328
rect 452524 351268 452640 351308
rect 452544 351248 452640 351268
rect 452544 350804 452640 350824
rect 452524 350764 452640 350804
rect 452544 350744 452640 350764
rect 452544 350300 452640 350320
rect 452524 350260 452640 350300
rect 452544 350240 452640 350260
rect 0 349796 96 349816
rect 452544 349796 452640 349816
rect 0 349756 116 349796
rect 452524 349756 452640 349796
rect 0 349736 96 349756
rect 452544 349736 452640 349756
rect 452544 349292 452640 349312
rect 452524 349252 452640 349292
rect 452544 349232 452640 349252
rect 0 348788 96 348808
rect 452544 348788 452640 348808
rect 0 348748 116 348788
rect 452524 348748 452640 348788
rect 0 348728 96 348748
rect 452544 348728 452640 348748
rect 452544 348284 452640 348304
rect 452524 348244 452640 348284
rect 452544 348224 452640 348244
rect 0 347780 96 347800
rect 452544 347780 452640 347800
rect 0 347740 116 347780
rect 452524 347740 452640 347780
rect 0 347720 96 347740
rect 452544 347720 452640 347740
rect 452544 347276 452640 347296
rect 452524 347236 452640 347276
rect 452544 347216 452640 347236
rect 0 346772 96 346792
rect 452544 346772 452640 346792
rect 0 346732 116 346772
rect 452524 346732 452640 346772
rect 0 346712 96 346732
rect 452544 346712 452640 346732
rect 452544 346268 452640 346288
rect 452524 346228 452640 346268
rect 452544 346208 452640 346228
rect 0 345764 96 345784
rect 452544 345764 452640 345784
rect 0 345724 116 345764
rect 452524 345724 452640 345764
rect 0 345704 96 345724
rect 452544 345704 452640 345724
rect 452544 345260 452640 345280
rect 452524 345220 452640 345260
rect 452544 345200 452640 345220
rect 0 344756 96 344776
rect 452544 344756 452640 344776
rect 0 344716 116 344756
rect 452524 344716 452640 344756
rect 0 344696 96 344716
rect 452544 344696 452640 344716
rect 452544 344252 452640 344272
rect 452524 344212 452640 344252
rect 452544 344192 452640 344212
rect 0 343748 96 343768
rect 452544 343748 452640 343768
rect 0 343708 116 343748
rect 452524 343708 452640 343748
rect 0 343688 96 343708
rect 452544 343688 452640 343708
rect 452544 343244 452640 343264
rect 452524 343204 452640 343244
rect 452544 343184 452640 343204
rect 0 342740 96 342760
rect 452544 342740 452640 342760
rect 0 342700 116 342740
rect 452524 342700 452640 342740
rect 0 342680 96 342700
rect 452544 342680 452640 342700
rect 452544 342236 452640 342256
rect 452524 342196 452640 342236
rect 452544 342176 452640 342196
rect 0 341732 96 341752
rect 452544 341732 452640 341752
rect 0 341692 116 341732
rect 452524 341692 452640 341732
rect 0 341672 96 341692
rect 452544 341672 452640 341692
rect 452544 341228 452640 341248
rect 452524 341188 452640 341228
rect 452544 341168 452640 341188
rect 0 340724 96 340744
rect 452544 340724 452640 340744
rect 0 340684 116 340724
rect 452524 340684 452640 340724
rect 0 340664 96 340684
rect 452544 340664 452640 340684
rect 452544 340220 452640 340240
rect 452524 340180 452640 340220
rect 452544 340160 452640 340180
rect 0 339716 96 339736
rect 452544 339716 452640 339736
rect 0 339676 116 339716
rect 452524 339676 452640 339716
rect 0 339656 96 339676
rect 452544 339656 452640 339676
rect 452544 339212 452640 339232
rect 452524 339172 452640 339212
rect 452544 339152 452640 339172
rect 0 338708 96 338728
rect 452544 338708 452640 338728
rect 0 338668 116 338708
rect 452524 338668 452640 338708
rect 0 338648 96 338668
rect 452544 338648 452640 338668
rect 452544 338204 452640 338224
rect 452524 338164 452640 338204
rect 452544 338144 452640 338164
rect 0 337700 96 337720
rect 452544 337700 452640 337720
rect 0 337660 116 337700
rect 452524 337660 452640 337700
rect 0 337640 96 337660
rect 452544 337640 452640 337660
rect 452544 337196 452640 337216
rect 452524 337156 452640 337196
rect 452544 337136 452640 337156
rect 0 336692 96 336712
rect 452544 336692 452640 336712
rect 0 336652 116 336692
rect 452524 336652 452640 336692
rect 0 336632 96 336652
rect 452544 336632 452640 336652
rect 452544 336188 452640 336208
rect 452524 336148 452640 336188
rect 452544 336128 452640 336148
rect 0 335684 96 335704
rect 452544 335684 452640 335704
rect 0 335644 116 335684
rect 452524 335644 452640 335684
rect 0 335624 96 335644
rect 452544 335624 452640 335644
rect 452544 335180 452640 335200
rect 452524 335140 452640 335180
rect 452544 335120 452640 335140
rect 0 334676 96 334696
rect 452544 334676 452640 334696
rect 0 334636 116 334676
rect 452524 334636 452640 334676
rect 0 334616 96 334636
rect 452544 334616 452640 334636
rect 452544 334172 452640 334192
rect 452524 334132 452640 334172
rect 452544 334112 452640 334132
rect 0 333668 96 333688
rect 452544 333668 452640 333688
rect 0 333628 116 333668
rect 452524 333628 452640 333668
rect 0 333608 96 333628
rect 452544 333608 452640 333628
rect 452544 333164 452640 333184
rect 452524 333124 452640 333164
rect 452544 333104 452640 333124
rect 0 332660 96 332680
rect 452544 332660 452640 332680
rect 0 332620 116 332660
rect 452524 332620 452640 332660
rect 0 332600 96 332620
rect 452544 332600 452640 332620
rect 452544 332156 452640 332176
rect 452524 332116 452640 332156
rect 452544 332096 452640 332116
rect 0 331652 96 331672
rect 452544 331652 452640 331672
rect 0 331612 116 331652
rect 452524 331612 452640 331652
rect 0 331592 96 331612
rect 452544 331592 452640 331612
rect 452544 331148 452640 331168
rect 452524 331108 452640 331148
rect 452544 331088 452640 331108
rect 0 330644 96 330664
rect 452544 330644 452640 330664
rect 0 330604 116 330644
rect 452524 330604 452640 330644
rect 0 330584 96 330604
rect 452544 330584 452640 330604
rect 452544 330140 452640 330160
rect 452524 330100 452640 330140
rect 452544 330080 452640 330100
rect 0 329636 96 329656
rect 452544 329636 452640 329656
rect 0 329596 116 329636
rect 452524 329596 452640 329636
rect 0 329576 96 329596
rect 452544 329576 452640 329596
rect 452544 329132 452640 329152
rect 452524 329092 452640 329132
rect 452544 329072 452640 329092
rect 0 328628 96 328648
rect 452544 328628 452640 328648
rect 0 328588 116 328628
rect 452524 328588 452640 328628
rect 0 328568 96 328588
rect 452544 328568 452640 328588
rect 452544 328124 452640 328144
rect 452524 328084 452640 328124
rect 452544 328064 452640 328084
rect 0 327620 96 327640
rect 452544 327620 452640 327640
rect 0 327580 116 327620
rect 452524 327580 452640 327620
rect 0 327560 96 327580
rect 452544 327560 452640 327580
rect 452544 327116 452640 327136
rect 452524 327076 452640 327116
rect 452544 327056 452640 327076
rect 0 326612 96 326632
rect 452544 326612 452640 326632
rect 0 326572 116 326612
rect 452524 326572 452640 326612
rect 0 326552 96 326572
rect 452544 326552 452640 326572
rect 452544 326108 452640 326128
rect 452524 326068 452640 326108
rect 452544 326048 452640 326068
rect 0 325604 96 325624
rect 452544 325604 452640 325624
rect 0 325564 116 325604
rect 452524 325564 452640 325604
rect 0 325544 96 325564
rect 452544 325544 452640 325564
rect 452544 325100 452640 325120
rect 452524 325060 452640 325100
rect 452544 325040 452640 325060
rect 0 324596 96 324616
rect 452544 324596 452640 324616
rect 0 324556 116 324596
rect 452524 324556 452640 324596
rect 0 324536 96 324556
rect 452544 324536 452640 324556
rect 452544 324092 452640 324112
rect 452524 324052 452640 324092
rect 452544 324032 452640 324052
rect 0 323588 96 323608
rect 452544 323588 452640 323608
rect 0 323548 116 323588
rect 452524 323548 452640 323588
rect 0 323528 96 323548
rect 452544 323528 452640 323548
rect 452544 323084 452640 323104
rect 452524 323044 452640 323084
rect 452544 323024 452640 323044
rect 0 322580 96 322600
rect 452544 322580 452640 322600
rect 0 322540 116 322580
rect 452524 322540 452640 322580
rect 0 322520 96 322540
rect 452544 322520 452640 322540
rect 452544 322076 452640 322096
rect 452524 322036 452640 322076
rect 452544 322016 452640 322036
rect 0 321572 96 321592
rect 452544 321572 452640 321592
rect 0 321532 116 321572
rect 452524 321532 452640 321572
rect 0 321512 96 321532
rect 452544 321512 452640 321532
rect 452544 321068 452640 321088
rect 452524 321028 452640 321068
rect 452544 321008 452640 321028
rect 0 320564 96 320584
rect 452544 320564 452640 320584
rect 0 320524 116 320564
rect 452524 320524 452640 320564
rect 0 320504 96 320524
rect 452544 320504 452640 320524
rect 452544 320060 452640 320080
rect 452524 320020 452640 320060
rect 452544 320000 452640 320020
rect 0 319556 96 319576
rect 452544 319556 452640 319576
rect 0 319516 116 319556
rect 452524 319516 452640 319556
rect 0 319496 96 319516
rect 452544 319496 452640 319516
rect 452544 319052 452640 319072
rect 452524 319012 452640 319052
rect 452544 318992 452640 319012
rect 0 318548 96 318568
rect 452544 318548 452640 318568
rect 0 318508 116 318548
rect 452524 318508 452640 318548
rect 0 318488 96 318508
rect 452544 318488 452640 318508
rect 452544 318044 452640 318064
rect 452524 318004 452640 318044
rect 452544 317984 452640 318004
rect 0 317540 96 317560
rect 452544 317540 452640 317560
rect 0 317500 116 317540
rect 452524 317500 452640 317540
rect 0 317480 96 317500
rect 452544 317480 452640 317500
rect 452544 317036 452640 317056
rect 452524 316996 452640 317036
rect 452544 316976 452640 316996
rect 0 316532 96 316552
rect 452544 316532 452640 316552
rect 0 316492 116 316532
rect 452524 316492 452640 316532
rect 0 316472 96 316492
rect 452544 316472 452640 316492
rect 452544 316028 452640 316048
rect 452524 315988 452640 316028
rect 452544 315968 452640 315988
rect 0 315524 96 315544
rect 452544 315524 452640 315544
rect 0 315484 116 315524
rect 452524 315484 452640 315524
rect 0 315464 96 315484
rect 452544 315464 452640 315484
rect 452544 315020 452640 315040
rect 452524 314980 452640 315020
rect 452544 314960 452640 314980
rect 0 314516 96 314536
rect 452544 314516 452640 314536
rect 0 314476 116 314516
rect 452524 314476 452640 314516
rect 0 314456 96 314476
rect 452544 314456 452640 314476
rect 452544 314012 452640 314032
rect 452524 313972 452640 314012
rect 452544 313952 452640 313972
rect 0 313508 96 313528
rect 452544 313508 452640 313528
rect 0 313468 116 313508
rect 452524 313468 452640 313508
rect 0 313448 96 313468
rect 452544 313448 452640 313468
rect 452544 313004 452640 313024
rect 452524 312964 452640 313004
rect 452544 312944 452640 312964
rect 0 312500 96 312520
rect 452544 312500 452640 312520
rect 0 312460 116 312500
rect 452524 312460 452640 312500
rect 0 312440 96 312460
rect 452544 312440 452640 312460
rect 452544 311996 452640 312016
rect 452524 311956 452640 311996
rect 452544 311936 452640 311956
rect 0 311492 96 311512
rect 452544 311492 452640 311512
rect 0 311452 116 311492
rect 452524 311452 452640 311492
rect 0 311432 96 311452
rect 452544 311432 452640 311452
rect 452544 310988 452640 311008
rect 452524 310948 452640 310988
rect 452544 310928 452640 310948
rect 0 310484 96 310504
rect 452544 310484 452640 310504
rect 0 310444 116 310484
rect 452524 310444 452640 310484
rect 0 310424 96 310444
rect 452544 310424 452640 310444
rect 452544 309980 452640 310000
rect 452524 309940 452640 309980
rect 452544 309920 452640 309940
rect 0 309476 96 309496
rect 452544 309476 452640 309496
rect 0 309436 116 309476
rect 452524 309436 452640 309476
rect 0 309416 96 309436
rect 452544 309416 452640 309436
rect 452544 308972 452640 308992
rect 452524 308932 452640 308972
rect 452544 308912 452640 308932
rect 0 308468 96 308488
rect 452544 308468 452640 308488
rect 0 308428 116 308468
rect 452524 308428 452640 308468
rect 0 308408 96 308428
rect 452544 308408 452640 308428
rect 452544 307964 452640 307984
rect 452524 307924 452640 307964
rect 452544 307904 452640 307924
rect 0 307460 96 307480
rect 452544 307460 452640 307480
rect 0 307420 116 307460
rect 452524 307420 452640 307460
rect 0 307400 96 307420
rect 452544 307400 452640 307420
rect 452544 306956 452640 306976
rect 452524 306916 452640 306956
rect 452544 306896 452640 306916
rect 0 306452 96 306472
rect 0 306412 116 306452
rect 0 306392 96 306412
rect 0 305444 96 305464
rect 0 305404 116 305444
rect 0 305384 96 305404
rect 0 304436 96 304456
rect 0 304396 116 304436
rect 0 304376 96 304396
rect 0 301412 96 301432
rect 0 301372 116 301412
rect 0 301352 96 301372
rect 0 300404 96 300424
rect 0 300364 116 300404
rect 0 300344 96 300364
rect 0 299396 96 299416
rect 0 299356 116 299396
rect 0 299336 96 299356
rect 0 298388 96 298408
rect 0 298348 116 298388
rect 0 298328 96 298348
rect 0 297380 96 297400
rect 0 297340 116 297380
rect 0 297320 96 297340
rect 0 296372 96 296392
rect 0 296332 116 296372
rect 0 296312 96 296332
rect 0 295364 96 295384
rect 0 295324 116 295364
rect 0 295304 96 295324
rect 0 294356 96 294376
rect 0 294316 116 294356
rect 0 294296 96 294316
rect 0 293348 96 293368
rect 0 293308 116 293348
rect 0 293288 96 293308
rect 0 292340 96 292360
rect 0 292300 116 292340
rect 0 292280 96 292300
rect 0 291332 96 291352
rect 0 291292 116 291332
rect 0 291272 96 291292
rect 0 290324 96 290344
rect 0 290284 116 290324
rect 0 290264 96 290284
rect 0 289316 96 289336
rect 0 289276 116 289316
rect 0 289256 96 289276
rect 0 288308 96 288328
rect 0 288268 116 288308
rect 0 288248 96 288268
rect 0 287300 96 287320
rect 0 287260 116 287300
rect 0 287240 96 287260
rect 0 286292 96 286312
rect 0 286252 116 286292
rect 0 286232 96 286252
rect 0 285284 96 285304
rect 0 285244 116 285284
rect 0 285224 96 285244
rect 0 284276 96 284296
rect 0 284236 116 284276
rect 0 284216 96 284236
rect 0 283268 96 283288
rect 0 283228 116 283268
rect 0 283208 96 283228
rect 0 282260 96 282280
rect 0 282220 116 282260
rect 0 282200 96 282220
rect 0 281252 96 281272
rect 0 281212 116 281252
rect 0 281192 96 281212
rect 0 280244 96 280264
rect 0 280204 116 280244
rect 0 280184 96 280204
rect 0 279236 96 279256
rect 0 279196 116 279236
rect 0 279176 96 279196
rect 0 278228 96 278248
rect 0 278188 116 278228
rect 0 278168 96 278188
rect 0 277220 96 277240
rect 0 277180 116 277220
rect 0 277160 96 277180
rect 0 276212 96 276232
rect 0 276172 116 276212
rect 0 276152 96 276172
rect 0 275204 96 275224
rect 0 275164 116 275204
rect 0 275144 96 275164
rect 0 274196 96 274216
rect 0 274156 116 274196
rect 0 274136 96 274156
rect 0 273188 96 273208
rect 0 273148 116 273188
rect 0 273128 96 273148
rect 0 272180 96 272200
rect 0 272140 116 272180
rect 0 272120 96 272140
rect 0 271172 96 271192
rect 0 271132 116 271172
rect 0 271112 96 271132
rect 0 270164 96 270184
rect 0 270124 116 270164
rect 0 270104 96 270124
rect 0 269156 96 269176
rect 0 269116 116 269156
rect 0 269096 96 269116
rect 0 268148 96 268168
rect 0 268108 116 268148
rect 0 268088 96 268108
rect 0 267140 96 267160
rect 0 267100 116 267140
rect 0 267080 96 267100
rect 452544 266636 452640 266656
rect 452524 266596 452640 266636
rect 452544 266576 452640 266596
rect 0 266132 96 266152
rect 452544 266132 452640 266152
rect 0 266092 116 266132
rect 452524 266092 452640 266132
rect 0 266072 96 266092
rect 452544 266072 452640 266092
rect 452544 265628 452640 265648
rect 452524 265588 452640 265628
rect 452544 265568 452640 265588
rect 0 265124 96 265144
rect 452544 265124 452640 265144
rect 0 265084 116 265124
rect 452524 265084 452640 265124
rect 0 265064 96 265084
rect 452544 265064 452640 265084
rect 452544 264620 452640 264640
rect 452524 264580 452640 264620
rect 452544 264560 452640 264580
rect 0 264116 96 264136
rect 452544 264116 452640 264136
rect 0 264076 116 264116
rect 452524 264076 452640 264116
rect 0 264056 96 264076
rect 452544 264056 452640 264076
rect 452544 263612 452640 263632
rect 452524 263572 452640 263612
rect 452544 263552 452640 263572
rect 0 263108 96 263128
rect 452544 263108 452640 263128
rect 0 263068 116 263108
rect 452524 263068 452640 263108
rect 0 263048 96 263068
rect 452544 263048 452640 263068
rect 452544 262604 452640 262624
rect 452524 262564 452640 262604
rect 452544 262544 452640 262564
rect 0 262100 96 262120
rect 452544 262100 452640 262120
rect 0 262060 116 262100
rect 452524 262060 452640 262100
rect 0 262040 96 262060
rect 452544 262040 452640 262060
rect 452544 261596 452640 261616
rect 452524 261556 452640 261596
rect 452544 261536 452640 261556
rect 0 261092 96 261112
rect 452544 261092 452640 261112
rect 0 261052 116 261092
rect 452524 261052 452640 261092
rect 0 261032 96 261052
rect 452544 261032 452640 261052
rect 452544 260588 452640 260608
rect 452524 260548 452640 260588
rect 452544 260528 452640 260548
rect 0 260084 96 260104
rect 452544 260084 452640 260104
rect 0 260044 116 260084
rect 452524 260044 452640 260084
rect 0 260024 96 260044
rect 452544 260024 452640 260044
rect 452544 259580 452640 259600
rect 452524 259540 452640 259580
rect 452544 259520 452640 259540
rect 0 259076 96 259096
rect 452544 259076 452640 259096
rect 0 259036 116 259076
rect 452524 259036 452640 259076
rect 0 259016 96 259036
rect 452544 259016 452640 259036
rect 452544 258572 452640 258592
rect 452524 258532 452640 258572
rect 452544 258512 452640 258532
rect 0 258068 96 258088
rect 452544 258068 452640 258088
rect 0 258028 116 258068
rect 452524 258028 452640 258068
rect 0 258008 96 258028
rect 452544 258008 452640 258028
rect 452544 257564 452640 257584
rect 452524 257524 452640 257564
rect 452544 257504 452640 257524
rect 0 257060 96 257080
rect 452544 257060 452640 257080
rect 0 257020 116 257060
rect 452524 257020 452640 257060
rect 0 257000 96 257020
rect 452544 257000 452640 257020
rect 452544 256556 452640 256576
rect 452524 256516 452640 256556
rect 452544 256496 452640 256516
rect 0 256052 96 256072
rect 452544 256052 452640 256072
rect 0 256012 116 256052
rect 452524 256012 452640 256052
rect 0 255992 96 256012
rect 452544 255992 452640 256012
rect 452544 255548 452640 255568
rect 452524 255508 452640 255548
rect 452544 255488 452640 255508
rect 452544 255044 452640 255064
rect 452524 255004 452640 255044
rect 452544 254984 452640 255004
rect 452544 254540 452640 254560
rect 452524 254500 452640 254540
rect 452544 254480 452640 254500
rect 452544 254036 452640 254056
rect 452524 253996 452640 254036
rect 452544 253976 452640 253996
rect 452544 253532 452640 253552
rect 452524 253492 452640 253532
rect 452544 253472 452640 253492
rect 0 253028 96 253048
rect 452544 253028 452640 253048
rect 0 252988 116 253028
rect 452524 252988 452640 253028
rect 0 252968 96 252988
rect 452544 252968 452640 252988
rect 452544 252524 452640 252544
rect 452524 252484 452640 252524
rect 452544 252464 452640 252484
rect 0 252020 96 252040
rect 452544 252020 452640 252040
rect 0 251980 116 252020
rect 452524 251980 452640 252020
rect 0 251960 96 251980
rect 452544 251960 452640 251980
rect 452544 251516 452640 251536
rect 452524 251476 452640 251516
rect 452544 251456 452640 251476
rect 0 251012 96 251032
rect 452544 251012 452640 251032
rect 0 250972 116 251012
rect 452524 250972 452640 251012
rect 0 250952 96 250972
rect 452544 250952 452640 250972
rect 452544 250508 452640 250528
rect 452524 250468 452640 250508
rect 452544 250448 452640 250468
rect 0 250004 96 250024
rect 452544 250004 452640 250024
rect 0 249964 116 250004
rect 452524 249964 452640 250004
rect 0 249944 96 249964
rect 452544 249944 452640 249964
rect 452544 249500 452640 249520
rect 452524 249460 452640 249500
rect 452544 249440 452640 249460
rect 0 248996 96 249016
rect 452544 248996 452640 249016
rect 0 248956 116 248996
rect 452524 248956 452640 248996
rect 0 248936 96 248956
rect 452544 248936 452640 248956
rect 452544 248492 452640 248512
rect 452524 248452 452640 248492
rect 452544 248432 452640 248452
rect 0 247988 96 248008
rect 452544 247988 452640 248008
rect 0 247948 116 247988
rect 452524 247948 452640 247988
rect 0 247928 96 247948
rect 452544 247928 452640 247948
rect 452544 247484 452640 247504
rect 452524 247444 452640 247484
rect 452544 247424 452640 247444
rect 0 246980 96 247000
rect 452544 246980 452640 247000
rect 0 246940 116 246980
rect 452524 246940 452640 246980
rect 0 246920 96 246940
rect 452544 246920 452640 246940
rect 452544 246476 452640 246496
rect 452524 246436 452640 246476
rect 452544 246416 452640 246436
rect 0 245972 96 245992
rect 452544 245972 452640 245992
rect 0 245932 116 245972
rect 452524 245932 452640 245972
rect 0 245912 96 245932
rect 452544 245912 452640 245932
rect 452544 245468 452640 245488
rect 452524 245428 452640 245468
rect 452544 245408 452640 245428
rect 0 244964 96 244984
rect 452544 244964 452640 244984
rect 0 244924 116 244964
rect 452524 244924 452640 244964
rect 0 244904 96 244924
rect 452544 244904 452640 244924
rect 452544 244460 452640 244480
rect 452524 244420 452640 244460
rect 452544 244400 452640 244420
rect 0 243956 96 243976
rect 452544 243956 452640 243976
rect 0 243916 116 243956
rect 452524 243916 452640 243956
rect 0 243896 96 243916
rect 452544 243896 452640 243916
rect 452544 243452 452640 243472
rect 452524 243412 452640 243452
rect 452544 243392 452640 243412
rect 0 242948 96 242968
rect 452544 242948 452640 242968
rect 0 242908 116 242948
rect 452524 242908 452640 242948
rect 0 242888 96 242908
rect 452544 242888 452640 242908
rect 452544 242444 452640 242464
rect 452524 242404 452640 242444
rect 452544 242384 452640 242404
rect 0 241940 96 241960
rect 452544 241940 452640 241960
rect 0 241900 116 241940
rect 452524 241900 452640 241940
rect 0 241880 96 241900
rect 452544 241880 452640 241900
rect 452544 241436 452640 241456
rect 452524 241396 452640 241436
rect 452544 241376 452640 241396
rect 0 240932 96 240952
rect 452544 240932 452640 240952
rect 0 240892 116 240932
rect 452524 240892 452640 240932
rect 0 240872 96 240892
rect 452544 240872 452640 240892
rect 452544 240428 452640 240448
rect 452524 240388 452640 240428
rect 452544 240368 452640 240388
rect 0 239924 96 239944
rect 452544 239924 452640 239944
rect 0 239884 116 239924
rect 452524 239884 452640 239924
rect 0 239864 96 239884
rect 452544 239864 452640 239884
rect 452544 239420 452640 239440
rect 452524 239380 452640 239420
rect 452544 239360 452640 239380
rect 0 238916 96 238936
rect 452544 238916 452640 238936
rect 0 238876 116 238916
rect 452524 238876 452640 238916
rect 0 238856 96 238876
rect 452544 238856 452640 238876
rect 452544 238412 452640 238432
rect 452524 238372 452640 238412
rect 452544 238352 452640 238372
rect 0 237908 96 237928
rect 452544 237908 452640 237928
rect 0 237868 116 237908
rect 452524 237868 452640 237908
rect 0 237848 96 237868
rect 452544 237848 452640 237868
rect 452544 237404 452640 237424
rect 452524 237364 452640 237404
rect 452544 237344 452640 237364
rect 0 236900 96 236920
rect 452544 236900 452640 236920
rect 0 236860 116 236900
rect 452524 236860 452640 236900
rect 0 236840 96 236860
rect 452544 236840 452640 236860
rect 452544 236396 452640 236416
rect 452524 236356 452640 236396
rect 452544 236336 452640 236356
rect 0 235892 96 235912
rect 452544 235892 452640 235912
rect 0 235852 116 235892
rect 452524 235852 452640 235892
rect 0 235832 96 235852
rect 452544 235832 452640 235852
rect 452544 235388 452640 235408
rect 452524 235348 452640 235388
rect 452544 235328 452640 235348
rect 0 234884 96 234904
rect 452544 234884 452640 234904
rect 0 234844 116 234884
rect 452524 234844 452640 234884
rect 0 234824 96 234844
rect 452544 234824 452640 234844
rect 452544 234380 452640 234400
rect 452524 234340 452640 234380
rect 452544 234320 452640 234340
rect 0 233876 96 233896
rect 452544 233876 452640 233896
rect 0 233836 116 233876
rect 452524 233836 452640 233876
rect 0 233816 96 233836
rect 452544 233816 452640 233836
rect 452544 233372 452640 233392
rect 452524 233332 452640 233372
rect 452544 233312 452640 233332
rect 0 232868 96 232888
rect 452544 232868 452640 232888
rect 0 232828 116 232868
rect 452524 232828 452640 232868
rect 0 232808 96 232828
rect 452544 232808 452640 232828
rect 452544 232364 452640 232384
rect 452524 232324 452640 232364
rect 452544 232304 452640 232324
rect 0 231860 96 231880
rect 452544 231860 452640 231880
rect 0 231820 116 231860
rect 452524 231820 452640 231860
rect 0 231800 96 231820
rect 452544 231800 452640 231820
rect 452544 231356 452640 231376
rect 452524 231316 452640 231356
rect 452544 231296 452640 231316
rect 0 230852 96 230872
rect 452544 230852 452640 230872
rect 0 230812 116 230852
rect 452524 230812 452640 230852
rect 0 230792 96 230812
rect 452544 230792 452640 230812
rect 452544 230348 452640 230368
rect 452524 230308 452640 230348
rect 452544 230288 452640 230308
rect 0 229844 96 229864
rect 452544 229844 452640 229864
rect 0 229804 116 229844
rect 452524 229804 452640 229844
rect 0 229784 96 229804
rect 452544 229784 452640 229804
rect 452544 229340 452640 229360
rect 452524 229300 452640 229340
rect 452544 229280 452640 229300
rect 0 228836 96 228856
rect 452544 228836 452640 228856
rect 0 228796 116 228836
rect 452524 228796 452640 228836
rect 0 228776 96 228796
rect 452544 228776 452640 228796
rect 452544 228332 452640 228352
rect 452524 228292 452640 228332
rect 452544 228272 452640 228292
rect 0 227828 96 227848
rect 452544 227828 452640 227848
rect 0 227788 116 227828
rect 452524 227788 452640 227828
rect 0 227768 96 227788
rect 452544 227768 452640 227788
rect 452544 227324 452640 227344
rect 452524 227284 452640 227324
rect 452544 227264 452640 227284
rect 0 226820 96 226840
rect 452544 226820 452640 226840
rect 0 226780 116 226820
rect 452524 226780 452640 226820
rect 0 226760 96 226780
rect 452544 226760 452640 226780
rect 452544 226316 452640 226336
rect 452524 226276 452640 226316
rect 452544 226256 452640 226276
rect 0 225812 96 225832
rect 452544 225812 452640 225832
rect 0 225772 116 225812
rect 452524 225772 452640 225812
rect 0 225752 96 225772
rect 452544 225752 452640 225772
rect 452544 225308 452640 225328
rect 452524 225268 452640 225308
rect 452544 225248 452640 225268
rect 0 224804 96 224824
rect 452544 224804 452640 224824
rect 0 224764 116 224804
rect 452524 224764 452640 224804
rect 0 224744 96 224764
rect 452544 224744 452640 224764
rect 452544 224300 452640 224320
rect 452524 224260 452640 224300
rect 452544 224240 452640 224260
rect 0 223796 96 223816
rect 452544 223796 452640 223816
rect 0 223756 116 223796
rect 452524 223756 452640 223796
rect 0 223736 96 223756
rect 452544 223736 452640 223756
rect 452544 223292 452640 223312
rect 452524 223252 452640 223292
rect 452544 223232 452640 223252
rect 0 222788 96 222808
rect 452544 222788 452640 222808
rect 0 222748 116 222788
rect 452524 222748 452640 222788
rect 0 222728 96 222748
rect 452544 222728 452640 222748
rect 452544 222284 452640 222304
rect 452524 222244 452640 222284
rect 452544 222224 452640 222244
rect 0 221780 96 221800
rect 452544 221780 452640 221800
rect 0 221740 116 221780
rect 452524 221740 452640 221780
rect 0 221720 96 221740
rect 452544 221720 452640 221740
rect 452544 221276 452640 221296
rect 452524 221236 452640 221276
rect 452544 221216 452640 221236
rect 0 220772 96 220792
rect 452544 220772 452640 220792
rect 0 220732 116 220772
rect 452524 220732 452640 220772
rect 0 220712 96 220732
rect 452544 220712 452640 220732
rect 452544 220268 452640 220288
rect 452524 220228 452640 220268
rect 452544 220208 452640 220228
rect 0 219764 96 219784
rect 452544 219764 452640 219784
rect 0 219724 116 219764
rect 452524 219724 452640 219764
rect 0 219704 96 219724
rect 452544 219704 452640 219724
rect 452544 219260 452640 219280
rect 452524 219220 452640 219260
rect 452544 219200 452640 219220
rect 0 218756 96 218776
rect 452544 218756 452640 218776
rect 0 218716 116 218756
rect 452524 218716 452640 218756
rect 0 218696 96 218716
rect 452544 218696 452640 218716
rect 452544 218252 452640 218272
rect 452524 218212 452640 218252
rect 452544 218192 452640 218212
rect 0 217748 96 217768
rect 452544 217748 452640 217768
rect 0 217708 116 217748
rect 452524 217708 452640 217748
rect 0 217688 96 217708
rect 452544 217688 452640 217708
rect 452544 217244 452640 217264
rect 452524 217204 452640 217244
rect 452544 217184 452640 217204
rect 0 216740 96 216760
rect 452544 216740 452640 216760
rect 0 216700 116 216740
rect 452524 216700 452640 216740
rect 0 216680 96 216700
rect 452544 216680 452640 216700
rect 452544 216236 452640 216256
rect 452524 216196 452640 216236
rect 452544 216176 452640 216196
rect 0 215732 96 215752
rect 452544 215732 452640 215752
rect 0 215692 116 215732
rect 452524 215692 452640 215732
rect 0 215672 96 215692
rect 452544 215672 452640 215692
rect 452544 215228 452640 215248
rect 452524 215188 452640 215228
rect 452544 215168 452640 215188
rect 0 214724 96 214744
rect 452544 214724 452640 214744
rect 0 214684 116 214724
rect 452524 214684 452640 214724
rect 0 214664 96 214684
rect 452544 214664 452640 214684
rect 452544 214220 452640 214240
rect 452524 214180 452640 214220
rect 452544 214160 452640 214180
rect 0 213716 96 213736
rect 452544 213716 452640 213736
rect 0 213676 116 213716
rect 452524 213676 452640 213716
rect 0 213656 96 213676
rect 452544 213656 452640 213676
rect 452544 213212 452640 213232
rect 452524 213172 452640 213212
rect 452544 213152 452640 213172
rect 0 212708 96 212728
rect 452544 212708 452640 212728
rect 0 212668 116 212708
rect 452524 212668 452640 212708
rect 0 212648 96 212668
rect 452544 212648 452640 212668
rect 452544 212204 452640 212224
rect 452524 212164 452640 212204
rect 452544 212144 452640 212164
rect 0 211700 96 211720
rect 452544 211700 452640 211720
rect 0 211660 116 211700
rect 452524 211660 452640 211700
rect 0 211640 96 211660
rect 452544 211640 452640 211660
rect 452544 211196 452640 211216
rect 452524 211156 452640 211196
rect 452544 211136 452640 211156
rect 0 210692 96 210712
rect 452544 210692 452640 210712
rect 0 210652 116 210692
rect 452524 210652 452640 210692
rect 0 210632 96 210652
rect 452544 210632 452640 210652
rect 452544 210188 452640 210208
rect 452524 210148 452640 210188
rect 452544 210128 452640 210148
rect 0 209684 96 209704
rect 0 209644 116 209684
rect 0 209624 96 209644
rect 0 208676 96 208696
rect 0 208636 116 208676
rect 0 208616 96 208636
rect 0 207668 96 207688
rect 0 207628 116 207668
rect 0 207608 96 207628
rect 0 204644 96 204664
rect 0 204604 116 204644
rect 0 204584 96 204604
rect 0 203636 96 203656
rect 0 203596 116 203636
rect 0 203576 96 203596
rect 0 202628 96 202648
rect 0 202588 116 202628
rect 0 202568 96 202588
rect 0 201620 96 201640
rect 0 201580 116 201620
rect 0 201560 96 201580
rect 0 200612 96 200632
rect 0 200572 116 200612
rect 0 200552 96 200572
rect 0 199604 96 199624
rect 0 199564 116 199604
rect 0 199544 96 199564
rect 0 198596 96 198616
rect 0 198556 116 198596
rect 0 198536 96 198556
rect 0 197588 96 197608
rect 0 197548 116 197588
rect 0 197528 96 197548
rect 0 196580 96 196600
rect 0 196540 116 196580
rect 0 196520 96 196540
rect 0 195572 96 195592
rect 0 195532 116 195572
rect 0 195512 96 195532
rect 0 194564 96 194584
rect 0 194524 116 194564
rect 0 194504 96 194524
rect 0 193556 96 193576
rect 0 193516 116 193556
rect 0 193496 96 193516
rect 0 192548 96 192568
rect 0 192508 116 192548
rect 0 192488 96 192508
rect 0 191540 96 191560
rect 0 191500 116 191540
rect 0 191480 96 191500
rect 0 190532 96 190552
rect 0 190492 116 190532
rect 0 190472 96 190492
rect 0 189524 96 189544
rect 0 189484 116 189524
rect 0 189464 96 189484
rect 0 188516 96 188536
rect 0 188476 116 188516
rect 0 188456 96 188476
rect 0 187508 96 187528
rect 0 187468 116 187508
rect 0 187448 96 187468
rect 0 186500 96 186520
rect 0 186460 116 186500
rect 0 186440 96 186460
rect 0 185492 96 185512
rect 0 185452 116 185492
rect 0 185432 96 185452
rect 0 184484 96 184504
rect 0 184444 116 184484
rect 0 184424 96 184444
rect 0 183476 96 183496
rect 0 183436 116 183476
rect 0 183416 96 183436
rect 0 182468 96 182488
rect 0 182428 116 182468
rect 0 182408 96 182428
rect 0 181460 96 181480
rect 0 181420 116 181460
rect 0 181400 96 181420
rect 0 180452 96 180472
rect 0 180412 116 180452
rect 0 180392 96 180412
rect 0 179444 96 179464
rect 0 179404 116 179444
rect 0 179384 96 179404
rect 0 178436 96 178456
rect 0 178396 116 178436
rect 0 178376 96 178396
rect 0 177428 96 177448
rect 0 177388 116 177428
rect 0 177368 96 177388
rect 0 176420 96 176440
rect 0 176380 116 176420
rect 0 176360 96 176380
rect 0 175412 96 175432
rect 0 175372 116 175412
rect 0 175352 96 175372
rect 0 174404 96 174424
rect 0 174364 116 174404
rect 0 174344 96 174364
rect 0 173396 96 173416
rect 0 173356 116 173396
rect 0 173336 96 173356
rect 0 172388 96 172408
rect 0 172348 116 172388
rect 0 172328 96 172348
rect 0 171380 96 171400
rect 0 171340 116 171380
rect 0 171320 96 171340
rect 0 170372 96 170392
rect 0 170332 116 170372
rect 0 170312 96 170332
rect 452544 169868 452640 169888
rect 452524 169828 452640 169868
rect 452544 169808 452640 169828
rect 0 169364 96 169384
rect 452544 169364 452640 169384
rect 0 169324 116 169364
rect 452524 169324 452640 169364
rect 0 169304 96 169324
rect 452544 169304 452640 169324
rect 452544 168860 452640 168880
rect 452524 168820 452640 168860
rect 452544 168800 452640 168820
rect 0 168356 96 168376
rect 452544 168356 452640 168376
rect 0 168316 116 168356
rect 452524 168316 452640 168356
rect 0 168296 96 168316
rect 452544 168296 452640 168316
rect 452544 167852 452640 167872
rect 452524 167812 452640 167852
rect 452544 167792 452640 167812
rect 0 167348 96 167368
rect 452544 167348 452640 167368
rect 0 167308 116 167348
rect 452524 167308 452640 167348
rect 0 167288 96 167308
rect 452544 167288 452640 167308
rect 452544 166844 452640 166864
rect 452524 166804 452640 166844
rect 452544 166784 452640 166804
rect 0 166340 96 166360
rect 452544 166340 452640 166360
rect 0 166300 116 166340
rect 452524 166300 452640 166340
rect 0 166280 96 166300
rect 452544 166280 452640 166300
rect 452544 165836 452640 165856
rect 452524 165796 452640 165836
rect 452544 165776 452640 165796
rect 0 165332 96 165352
rect 452544 165332 452640 165352
rect 0 165292 116 165332
rect 452524 165292 452640 165332
rect 0 165272 96 165292
rect 452544 165272 452640 165292
rect 452544 164828 452640 164848
rect 452524 164788 452640 164828
rect 452544 164768 452640 164788
rect 0 164324 96 164344
rect 452544 164324 452640 164344
rect 0 164284 116 164324
rect 452524 164284 452640 164324
rect 0 164264 96 164284
rect 452544 164264 452640 164284
rect 452544 163820 452640 163840
rect 452524 163780 452640 163820
rect 452544 163760 452640 163780
rect 0 163316 96 163336
rect 452544 163316 452640 163336
rect 0 163276 116 163316
rect 452524 163276 452640 163316
rect 0 163256 96 163276
rect 452544 163256 452640 163276
rect 452544 162812 452640 162832
rect 452524 162772 452640 162812
rect 452544 162752 452640 162772
rect 0 162308 96 162328
rect 452544 162308 452640 162328
rect 0 162268 116 162308
rect 452524 162268 452640 162308
rect 0 162248 96 162268
rect 452544 162248 452640 162268
rect 452544 161804 452640 161824
rect 452524 161764 452640 161804
rect 452544 161744 452640 161764
rect 0 161300 96 161320
rect 452544 161300 452640 161320
rect 0 161260 116 161300
rect 452524 161260 452640 161300
rect 0 161240 96 161260
rect 452544 161240 452640 161260
rect 452544 160796 452640 160816
rect 452524 160756 452640 160796
rect 452544 160736 452640 160756
rect 0 160292 96 160312
rect 452544 160292 452640 160312
rect 0 160252 116 160292
rect 452524 160252 452640 160292
rect 0 160232 96 160252
rect 452544 160232 452640 160252
rect 452544 159788 452640 159808
rect 452524 159748 452640 159788
rect 452544 159728 452640 159748
rect 0 159284 96 159304
rect 452544 159284 452640 159304
rect 0 159244 116 159284
rect 452524 159244 452640 159284
rect 0 159224 96 159244
rect 452544 159224 452640 159244
rect 452544 158780 452640 158800
rect 452524 158740 452640 158780
rect 452544 158720 452640 158740
rect 452544 158276 452640 158296
rect 452524 158236 452640 158276
rect 452544 158216 452640 158236
rect 452544 157772 452640 157792
rect 452524 157732 452640 157772
rect 452544 157712 452640 157732
rect 452544 157268 452640 157288
rect 452524 157228 452640 157268
rect 452544 157208 452640 157228
rect 452544 156764 452640 156784
rect 452524 156724 452640 156764
rect 452544 156704 452640 156724
rect 0 156260 96 156280
rect 452544 156260 452640 156280
rect 0 156220 116 156260
rect 452524 156220 452640 156260
rect 0 156200 96 156220
rect 452544 156200 452640 156220
rect 452544 155756 452640 155776
rect 452524 155716 452640 155756
rect 452544 155696 452640 155716
rect 0 155252 96 155272
rect 452544 155252 452640 155272
rect 0 155212 116 155252
rect 452524 155212 452640 155252
rect 0 155192 96 155212
rect 452544 155192 452640 155212
rect 452544 154748 452640 154768
rect 452524 154708 452640 154748
rect 452544 154688 452640 154708
rect 0 154244 96 154264
rect 452544 154244 452640 154264
rect 0 154204 116 154244
rect 452524 154204 452640 154244
rect 0 154184 96 154204
rect 452544 154184 452640 154204
rect 452544 153740 452640 153760
rect 452524 153700 452640 153740
rect 452544 153680 452640 153700
rect 0 153236 96 153256
rect 452544 153236 452640 153256
rect 0 153196 116 153236
rect 452524 153196 452640 153236
rect 0 153176 96 153196
rect 452544 153176 452640 153196
rect 452544 152732 452640 152752
rect 452524 152692 452640 152732
rect 452544 152672 452640 152692
rect 0 152228 96 152248
rect 452544 152228 452640 152248
rect 0 152188 116 152228
rect 452524 152188 452640 152228
rect 0 152168 96 152188
rect 452544 152168 452640 152188
rect 452544 151724 452640 151744
rect 452524 151684 452640 151724
rect 452544 151664 452640 151684
rect 0 151220 96 151240
rect 452544 151220 452640 151240
rect 0 151180 116 151220
rect 452524 151180 452640 151220
rect 0 151160 96 151180
rect 452544 151160 452640 151180
rect 452544 150716 452640 150736
rect 452524 150676 452640 150716
rect 452544 150656 452640 150676
rect 0 150212 96 150232
rect 452544 150212 452640 150232
rect 0 150172 116 150212
rect 452524 150172 452640 150212
rect 0 150152 96 150172
rect 452544 150152 452640 150172
rect 452544 149708 452640 149728
rect 452524 149668 452640 149708
rect 452544 149648 452640 149668
rect 0 149204 96 149224
rect 452544 149204 452640 149224
rect 0 149164 116 149204
rect 452524 149164 452640 149204
rect 0 149144 96 149164
rect 452544 149144 452640 149164
rect 452544 148700 452640 148720
rect 452524 148660 452640 148700
rect 452544 148640 452640 148660
rect 0 148196 96 148216
rect 452544 148196 452640 148216
rect 0 148156 116 148196
rect 452524 148156 452640 148196
rect 0 148136 96 148156
rect 452544 148136 452640 148156
rect 452544 147692 452640 147712
rect 452524 147652 452640 147692
rect 452544 147632 452640 147652
rect 0 147188 96 147208
rect 452544 147188 452640 147208
rect 0 147148 116 147188
rect 452524 147148 452640 147188
rect 0 147128 96 147148
rect 452544 147128 452640 147148
rect 452544 146684 452640 146704
rect 452524 146644 452640 146684
rect 452544 146624 452640 146644
rect 0 146180 96 146200
rect 452544 146180 452640 146200
rect 0 146140 116 146180
rect 452524 146140 452640 146180
rect 0 146120 96 146140
rect 452544 146120 452640 146140
rect 452544 145676 452640 145696
rect 452524 145636 452640 145676
rect 452544 145616 452640 145636
rect 0 145172 96 145192
rect 452544 145172 452640 145192
rect 0 145132 116 145172
rect 452524 145132 452640 145172
rect 0 145112 96 145132
rect 452544 145112 452640 145132
rect 452544 144668 452640 144688
rect 452524 144628 452640 144668
rect 452544 144608 452640 144628
rect 0 144164 96 144184
rect 452544 144164 452640 144184
rect 0 144124 116 144164
rect 452524 144124 452640 144164
rect 0 144104 96 144124
rect 452544 144104 452640 144124
rect 452544 143660 452640 143680
rect 452524 143620 452640 143660
rect 452544 143600 452640 143620
rect 0 143156 96 143176
rect 452544 143156 452640 143176
rect 0 143116 116 143156
rect 452524 143116 452640 143156
rect 0 143096 96 143116
rect 452544 143096 452640 143116
rect 452544 142652 452640 142672
rect 452524 142612 452640 142652
rect 452544 142592 452640 142612
rect 0 142148 96 142168
rect 452544 142148 452640 142168
rect 0 142108 116 142148
rect 452524 142108 452640 142148
rect 0 142088 96 142108
rect 452544 142088 452640 142108
rect 452544 141644 452640 141664
rect 452524 141604 452640 141644
rect 452544 141584 452640 141604
rect 0 141140 96 141160
rect 452544 141140 452640 141160
rect 0 141100 116 141140
rect 452524 141100 452640 141140
rect 0 141080 96 141100
rect 452544 141080 452640 141100
rect 452544 140636 452640 140656
rect 452524 140596 452640 140636
rect 452544 140576 452640 140596
rect 0 140132 96 140152
rect 452544 140132 452640 140152
rect 0 140092 116 140132
rect 452524 140092 452640 140132
rect 0 140072 96 140092
rect 452544 140072 452640 140092
rect 452544 139628 452640 139648
rect 452524 139588 452640 139628
rect 452544 139568 452640 139588
rect 0 139124 96 139144
rect 452544 139124 452640 139144
rect 0 139084 116 139124
rect 452524 139084 452640 139124
rect 0 139064 96 139084
rect 452544 139064 452640 139084
rect 452544 138620 452640 138640
rect 452524 138580 452640 138620
rect 452544 138560 452640 138580
rect 0 138116 96 138136
rect 452544 138116 452640 138136
rect 0 138076 116 138116
rect 452524 138076 452640 138116
rect 0 138056 96 138076
rect 452544 138056 452640 138076
rect 452544 137612 452640 137632
rect 452524 137572 452640 137612
rect 452544 137552 452640 137572
rect 0 137108 96 137128
rect 452544 137108 452640 137128
rect 0 137068 116 137108
rect 452524 137068 452640 137108
rect 0 137048 96 137068
rect 452544 137048 452640 137068
rect 452544 136604 452640 136624
rect 452524 136564 452640 136604
rect 452544 136544 452640 136564
rect 0 136100 96 136120
rect 452544 136100 452640 136120
rect 0 136060 116 136100
rect 452524 136060 452640 136100
rect 0 136040 96 136060
rect 452544 136040 452640 136060
rect 452544 135596 452640 135616
rect 452524 135556 452640 135596
rect 452544 135536 452640 135556
rect 0 135092 96 135112
rect 452544 135092 452640 135112
rect 0 135052 116 135092
rect 452524 135052 452640 135092
rect 0 135032 96 135052
rect 452544 135032 452640 135052
rect 452544 134588 452640 134608
rect 452524 134548 452640 134588
rect 452544 134528 452640 134548
rect 0 134084 96 134104
rect 452544 134084 452640 134104
rect 0 134044 116 134084
rect 452524 134044 452640 134084
rect 0 134024 96 134044
rect 452544 134024 452640 134044
rect 452544 133580 452640 133600
rect 452524 133540 452640 133580
rect 452544 133520 452640 133540
rect 0 133076 96 133096
rect 452544 133076 452640 133096
rect 0 133036 116 133076
rect 452524 133036 452640 133076
rect 0 133016 96 133036
rect 452544 133016 452640 133036
rect 452544 132572 452640 132592
rect 452524 132532 452640 132572
rect 452544 132512 452640 132532
rect 0 132068 96 132088
rect 452544 132068 452640 132088
rect 0 132028 116 132068
rect 452524 132028 452640 132068
rect 0 132008 96 132028
rect 452544 132008 452640 132028
rect 452544 131564 452640 131584
rect 452524 131524 452640 131564
rect 452544 131504 452640 131524
rect 0 131060 96 131080
rect 452544 131060 452640 131080
rect 0 131020 116 131060
rect 452524 131020 452640 131060
rect 0 131000 96 131020
rect 452544 131000 452640 131020
rect 452544 130556 452640 130576
rect 452524 130516 452640 130556
rect 452544 130496 452640 130516
rect 0 130052 96 130072
rect 452544 130052 452640 130072
rect 0 130012 116 130052
rect 452524 130012 452640 130052
rect 0 129992 96 130012
rect 452544 129992 452640 130012
rect 452544 129548 452640 129568
rect 452524 129508 452640 129548
rect 452544 129488 452640 129508
rect 0 129044 96 129064
rect 452544 129044 452640 129064
rect 0 129004 116 129044
rect 452524 129004 452640 129044
rect 0 128984 96 129004
rect 452544 128984 452640 129004
rect 452544 128540 452640 128560
rect 452524 128500 452640 128540
rect 452544 128480 452640 128500
rect 0 128036 96 128056
rect 452544 128036 452640 128056
rect 0 127996 116 128036
rect 452524 127996 452640 128036
rect 0 127976 96 127996
rect 452544 127976 452640 127996
rect 452544 127532 452640 127552
rect 452524 127492 452640 127532
rect 452544 127472 452640 127492
rect 0 127028 96 127048
rect 452544 127028 452640 127048
rect 0 126988 116 127028
rect 452524 126988 452640 127028
rect 0 126968 96 126988
rect 452544 126968 452640 126988
rect 452544 126524 452640 126544
rect 452524 126484 452640 126524
rect 452544 126464 452640 126484
rect 0 126020 96 126040
rect 452544 126020 452640 126040
rect 0 125980 116 126020
rect 452524 125980 452640 126020
rect 0 125960 96 125980
rect 452544 125960 452640 125980
rect 452544 125516 452640 125536
rect 452524 125476 452640 125516
rect 452544 125456 452640 125476
rect 0 125012 96 125032
rect 452544 125012 452640 125032
rect 0 124972 116 125012
rect 452524 124972 452640 125012
rect 0 124952 96 124972
rect 452544 124952 452640 124972
rect 452544 124508 452640 124528
rect 452524 124468 452640 124508
rect 452544 124448 452640 124468
rect 0 124004 96 124024
rect 452544 124004 452640 124024
rect 0 123964 116 124004
rect 452524 123964 452640 124004
rect 0 123944 96 123964
rect 452544 123944 452640 123964
rect 452544 123500 452640 123520
rect 452524 123460 452640 123500
rect 452544 123440 452640 123460
rect 0 122996 96 123016
rect 452544 122996 452640 123016
rect 0 122956 116 122996
rect 452524 122956 452640 122996
rect 0 122936 96 122956
rect 452544 122936 452640 122956
rect 452544 122492 452640 122512
rect 452524 122452 452640 122492
rect 452544 122432 452640 122452
rect 0 121988 96 122008
rect 452544 121988 452640 122008
rect 0 121948 116 121988
rect 452524 121948 452640 121988
rect 0 121928 96 121948
rect 452544 121928 452640 121948
rect 452544 121484 452640 121504
rect 452524 121444 452640 121484
rect 452544 121424 452640 121444
rect 0 120980 96 121000
rect 452544 120980 452640 121000
rect 0 120940 116 120980
rect 452524 120940 452640 120980
rect 0 120920 96 120940
rect 452544 120920 452640 120940
rect 452544 120476 452640 120496
rect 452524 120436 452640 120476
rect 452544 120416 452640 120436
rect 0 119972 96 119992
rect 452544 119972 452640 119992
rect 0 119932 116 119972
rect 452524 119932 452640 119972
rect 0 119912 96 119932
rect 452544 119912 452640 119932
rect 452544 119468 452640 119488
rect 452524 119428 452640 119468
rect 452544 119408 452640 119428
rect 0 118964 96 118984
rect 452544 118964 452640 118984
rect 0 118924 116 118964
rect 452524 118924 452640 118964
rect 0 118904 96 118924
rect 452544 118904 452640 118924
rect 452544 118460 452640 118480
rect 452524 118420 452640 118460
rect 452544 118400 452640 118420
rect 0 117956 96 117976
rect 452544 117956 452640 117976
rect 0 117916 116 117956
rect 452524 117916 452640 117956
rect 0 117896 96 117916
rect 452544 117896 452640 117916
rect 452544 117452 452640 117472
rect 452524 117412 452640 117452
rect 452544 117392 452640 117412
rect 0 116948 96 116968
rect 452544 116948 452640 116968
rect 0 116908 116 116948
rect 452524 116908 452640 116948
rect 0 116888 96 116908
rect 452544 116888 452640 116908
rect 452544 116444 452640 116464
rect 452524 116404 452640 116444
rect 452544 116384 452640 116404
rect 0 115940 96 115960
rect 452544 115940 452640 115960
rect 0 115900 116 115940
rect 452524 115900 452640 115940
rect 0 115880 96 115900
rect 452544 115880 452640 115900
rect 452544 115436 452640 115456
rect 452524 115396 452640 115436
rect 452544 115376 452640 115396
rect 0 114932 96 114952
rect 452544 114932 452640 114952
rect 0 114892 116 114932
rect 452524 114892 452640 114932
rect 0 114872 96 114892
rect 452544 114872 452640 114892
rect 452544 114428 452640 114448
rect 452524 114388 452640 114428
rect 452544 114368 452640 114388
rect 0 113924 96 113944
rect 452544 113924 452640 113944
rect 0 113884 116 113924
rect 452524 113884 452640 113924
rect 0 113864 96 113884
rect 452544 113864 452640 113884
rect 452544 113420 452640 113440
rect 452524 113380 452640 113420
rect 452544 113360 452640 113380
rect 0 112916 96 112936
rect 0 112876 116 112916
rect 0 112856 96 112876
rect 0 111908 96 111928
rect 0 111868 116 111908
rect 0 111848 96 111868
rect 0 110900 96 110920
rect 0 110860 116 110900
rect 0 110840 96 110860
rect 0 107876 96 107896
rect 0 107836 116 107876
rect 0 107816 96 107836
rect 0 106868 96 106888
rect 0 106828 116 106868
rect 0 106808 96 106828
rect 0 105860 96 105880
rect 0 105820 116 105860
rect 0 105800 96 105820
rect 0 104852 96 104872
rect 0 104812 116 104852
rect 0 104792 96 104812
rect 0 103844 96 103864
rect 0 103804 116 103844
rect 0 103784 96 103804
rect 0 102836 96 102856
rect 0 102796 116 102836
rect 0 102776 96 102796
rect 0 101828 96 101848
rect 0 101788 116 101828
rect 0 101768 96 101788
rect 0 100820 96 100840
rect 0 100780 116 100820
rect 0 100760 96 100780
rect 0 99812 96 99832
rect 0 99772 116 99812
rect 0 99752 96 99772
rect 0 98804 96 98824
rect 0 98764 116 98804
rect 0 98744 96 98764
rect 0 97796 96 97816
rect 0 97756 116 97796
rect 0 97736 96 97756
rect 0 96788 96 96808
rect 0 96748 116 96788
rect 0 96728 96 96748
rect 0 95780 96 95800
rect 0 95740 116 95780
rect 0 95720 96 95740
rect 0 94772 96 94792
rect 0 94732 116 94772
rect 0 94712 96 94732
rect 0 93764 96 93784
rect 0 93724 116 93764
rect 0 93704 96 93724
rect 0 92756 96 92776
rect 0 92716 116 92756
rect 0 92696 96 92716
rect 0 91748 96 91768
rect 0 91708 116 91748
rect 0 91688 96 91708
rect 0 90740 96 90760
rect 0 90700 116 90740
rect 0 90680 96 90700
rect 0 89732 96 89752
rect 0 89692 116 89732
rect 0 89672 96 89692
rect 0 88724 96 88744
rect 0 88684 116 88724
rect 0 88664 96 88684
rect 0 87716 96 87736
rect 0 87676 116 87716
rect 0 87656 96 87676
rect 0 86708 96 86728
rect 0 86668 116 86708
rect 0 86648 96 86668
rect 0 85700 96 85720
rect 0 85660 116 85700
rect 0 85640 96 85660
rect 0 84692 96 84712
rect 0 84652 116 84692
rect 0 84632 96 84652
rect 0 83684 96 83704
rect 0 83644 116 83684
rect 0 83624 96 83644
rect 0 82676 96 82696
rect 0 82636 116 82676
rect 0 82616 96 82636
rect 0 81668 96 81688
rect 0 81628 116 81668
rect 0 81608 96 81628
rect 0 80660 96 80680
rect 0 80620 116 80660
rect 0 80600 96 80620
rect 0 79652 96 79672
rect 0 79612 116 79652
rect 0 79592 96 79612
rect 0 78644 96 78664
rect 0 78604 116 78644
rect 0 78584 96 78604
rect 0 77636 96 77656
rect 0 77596 116 77636
rect 0 77576 96 77596
rect 0 76628 96 76648
rect 0 76588 116 76628
rect 0 76568 96 76588
rect 0 75620 96 75640
rect 0 75580 116 75620
rect 0 75560 96 75580
rect 0 74612 96 74632
rect 0 74572 116 74612
rect 0 74552 96 74572
rect 0 73604 96 73624
rect 0 73564 116 73604
rect 0 73544 96 73564
rect 452544 73100 452640 73120
rect 452524 73060 452640 73100
rect 452544 73040 452640 73060
rect 0 72596 96 72616
rect 452544 72596 452640 72616
rect 0 72556 116 72596
rect 452524 72556 452640 72596
rect 0 72536 96 72556
rect 452544 72536 452640 72556
rect 452544 72092 452640 72112
rect 452524 72052 452640 72092
rect 452544 72032 452640 72052
rect 0 71588 96 71608
rect 452544 71588 452640 71608
rect 0 71548 116 71588
rect 452524 71548 452640 71588
rect 0 71528 96 71548
rect 452544 71528 452640 71548
rect 452544 71084 452640 71104
rect 452524 71044 452640 71084
rect 452544 71024 452640 71044
rect 0 70580 96 70600
rect 452544 70580 452640 70600
rect 0 70540 116 70580
rect 452524 70540 452640 70580
rect 0 70520 96 70540
rect 452544 70520 452640 70540
rect 452544 70076 452640 70096
rect 452524 70036 452640 70076
rect 452544 70016 452640 70036
rect 0 69572 96 69592
rect 452544 69572 452640 69592
rect 0 69532 116 69572
rect 452524 69532 452640 69572
rect 0 69512 96 69532
rect 452544 69512 452640 69532
rect 452544 69068 452640 69088
rect 452524 69028 452640 69068
rect 452544 69008 452640 69028
rect 0 68564 96 68584
rect 452544 68564 452640 68584
rect 0 68524 116 68564
rect 452524 68524 452640 68564
rect 0 68504 96 68524
rect 452544 68504 452640 68524
rect 452544 68060 452640 68080
rect 452524 68020 452640 68060
rect 452544 68000 452640 68020
rect 0 67556 96 67576
rect 452544 67556 452640 67576
rect 0 67516 116 67556
rect 452524 67516 452640 67556
rect 0 67496 96 67516
rect 452544 67496 452640 67516
rect 452544 67052 452640 67072
rect 452524 67012 452640 67052
rect 452544 66992 452640 67012
rect 0 66548 96 66568
rect 452544 66548 452640 66568
rect 0 66508 116 66548
rect 452524 66508 452640 66548
rect 0 66488 96 66508
rect 452544 66488 452640 66508
rect 452544 66044 452640 66064
rect 452524 66004 452640 66044
rect 452544 65984 452640 66004
rect 0 65540 96 65560
rect 452544 65540 452640 65560
rect 0 65500 116 65540
rect 452524 65500 452640 65540
rect 0 65480 96 65500
rect 452544 65480 452640 65500
rect 452544 65036 452640 65056
rect 452524 64996 452640 65036
rect 452544 64976 452640 64996
rect 0 64532 96 64552
rect 452544 64532 452640 64552
rect 0 64492 116 64532
rect 452524 64492 452640 64532
rect 0 64472 96 64492
rect 452544 64472 452640 64492
rect 452544 64028 452640 64048
rect 452524 63988 452640 64028
rect 452544 63968 452640 63988
rect 0 63524 96 63544
rect 452544 63524 452640 63544
rect 0 63484 116 63524
rect 452524 63484 452640 63524
rect 0 63464 96 63484
rect 452544 63464 452640 63484
rect 452544 63020 452640 63040
rect 452524 62980 452640 63020
rect 452544 62960 452640 62980
rect 0 62516 96 62536
rect 452544 62516 452640 62536
rect 0 62476 116 62516
rect 452524 62476 452640 62516
rect 0 62456 96 62476
rect 452544 62456 452640 62476
rect 452544 62012 452640 62032
rect 452524 61972 452640 62012
rect 452544 61952 452640 61972
rect 452544 61508 452640 61528
rect 452524 61468 452640 61508
rect 452544 61448 452640 61468
rect 452544 61004 452640 61024
rect 452524 60964 452640 61004
rect 452544 60944 452640 60964
rect 452544 60500 452640 60520
rect 452524 60460 452640 60500
rect 452544 60440 452640 60460
rect 452544 59996 452640 60016
rect 452524 59956 452640 59996
rect 452544 59936 452640 59956
rect 0 59492 96 59512
rect 452544 59492 452640 59512
rect 0 59452 116 59492
rect 452524 59452 452640 59492
rect 0 59432 96 59452
rect 452544 59432 452640 59452
rect 452544 58988 452640 59008
rect 452524 58948 452640 58988
rect 452544 58928 452640 58948
rect 0 58484 96 58504
rect 452544 58484 452640 58504
rect 0 58444 116 58484
rect 452524 58444 452640 58484
rect 0 58424 96 58444
rect 452544 58424 452640 58444
rect 452544 57980 452640 58000
rect 452524 57940 452640 57980
rect 452544 57920 452640 57940
rect 0 57476 96 57496
rect 452544 57476 452640 57496
rect 0 57436 116 57476
rect 452524 57436 452640 57476
rect 0 57416 96 57436
rect 452544 57416 452640 57436
rect 452544 56972 452640 56992
rect 452524 56932 452640 56972
rect 452544 56912 452640 56932
rect 0 56468 96 56488
rect 452544 56468 452640 56488
rect 0 56428 116 56468
rect 452524 56428 452640 56468
rect 0 56408 96 56428
rect 452544 56408 452640 56428
rect 452544 55964 452640 55984
rect 452524 55924 452640 55964
rect 452544 55904 452640 55924
rect 0 55460 96 55480
rect 452544 55460 452640 55480
rect 0 55420 116 55460
rect 452524 55420 452640 55460
rect 0 55400 96 55420
rect 452544 55400 452640 55420
rect 452544 54956 452640 54976
rect 452524 54916 452640 54956
rect 452544 54896 452640 54916
rect 0 54452 96 54472
rect 452544 54452 452640 54472
rect 0 54412 116 54452
rect 452524 54412 452640 54452
rect 0 54392 96 54412
rect 452544 54392 452640 54412
rect 452544 53948 452640 53968
rect 452524 53908 452640 53948
rect 452544 53888 452640 53908
rect 0 53444 96 53464
rect 452544 53444 452640 53464
rect 0 53404 116 53444
rect 452524 53404 452640 53444
rect 0 53384 96 53404
rect 452544 53384 452640 53404
rect 452544 52940 452640 52960
rect 452524 52900 452640 52940
rect 452544 52880 452640 52900
rect 0 52436 96 52456
rect 452544 52436 452640 52456
rect 0 52396 116 52436
rect 452524 52396 452640 52436
rect 0 52376 96 52396
rect 452544 52376 452640 52396
rect 452544 51932 452640 51952
rect 452524 51892 452640 51932
rect 452544 51872 452640 51892
rect 0 51428 96 51448
rect 452544 51428 452640 51448
rect 0 51388 116 51428
rect 452524 51388 452640 51428
rect 0 51368 96 51388
rect 452544 51368 452640 51388
rect 452544 50924 452640 50944
rect 452524 50884 452640 50924
rect 452544 50864 452640 50884
rect 0 50420 96 50440
rect 452544 50420 452640 50440
rect 0 50380 116 50420
rect 452524 50380 452640 50420
rect 0 50360 96 50380
rect 452544 50360 452640 50380
rect 452544 49916 452640 49936
rect 452524 49876 452640 49916
rect 452544 49856 452640 49876
rect 0 49412 96 49432
rect 452544 49412 452640 49432
rect 0 49372 116 49412
rect 452524 49372 452640 49412
rect 0 49352 96 49372
rect 452544 49352 452640 49372
rect 452544 48908 452640 48928
rect 452524 48868 452640 48908
rect 452544 48848 452640 48868
rect 0 48404 96 48424
rect 452544 48404 452640 48424
rect 0 48364 116 48404
rect 452524 48364 452640 48404
rect 0 48344 96 48364
rect 452544 48344 452640 48364
rect 452544 47900 452640 47920
rect 452524 47860 452640 47900
rect 452544 47840 452640 47860
rect 0 47396 96 47416
rect 452544 47396 452640 47416
rect 0 47356 116 47396
rect 452524 47356 452640 47396
rect 0 47336 96 47356
rect 452544 47336 452640 47356
rect 452544 46892 452640 46912
rect 452524 46852 452640 46892
rect 452544 46832 452640 46852
rect 0 46388 96 46408
rect 452544 46388 452640 46408
rect 0 46348 116 46388
rect 452524 46348 452640 46388
rect 0 46328 96 46348
rect 452544 46328 452640 46348
rect 452544 45884 452640 45904
rect 452524 45844 452640 45884
rect 452544 45824 452640 45844
rect 0 45380 96 45400
rect 452544 45380 452640 45400
rect 0 45340 116 45380
rect 452524 45340 452640 45380
rect 0 45320 96 45340
rect 452544 45320 452640 45340
rect 452544 44876 452640 44896
rect 452524 44836 452640 44876
rect 452544 44816 452640 44836
rect 0 44372 96 44392
rect 452544 44372 452640 44392
rect 0 44332 116 44372
rect 452524 44332 452640 44372
rect 0 44312 96 44332
rect 452544 44312 452640 44332
rect 452544 43868 452640 43888
rect 452524 43828 452640 43868
rect 452544 43808 452640 43828
rect 0 43364 96 43384
rect 452544 43364 452640 43384
rect 0 43324 116 43364
rect 452524 43324 452640 43364
rect 0 43304 96 43324
rect 452544 43304 452640 43324
rect 452544 42860 452640 42880
rect 452524 42820 452640 42860
rect 452544 42800 452640 42820
rect 0 42356 96 42376
rect 452544 42356 452640 42376
rect 0 42316 116 42356
rect 452524 42316 452640 42356
rect 0 42296 96 42316
rect 452544 42296 452640 42316
rect 452544 41852 452640 41872
rect 452524 41812 452640 41852
rect 452544 41792 452640 41812
rect 0 41348 96 41368
rect 452544 41348 452640 41368
rect 0 41308 116 41348
rect 452524 41308 452640 41348
rect 0 41288 96 41308
rect 452544 41288 452640 41308
rect 452544 40844 452640 40864
rect 452524 40804 452640 40844
rect 452544 40784 452640 40804
rect 0 40340 96 40360
rect 452544 40340 452640 40360
rect 0 40300 116 40340
rect 452524 40300 452640 40340
rect 0 40280 96 40300
rect 452544 40280 452640 40300
rect 452544 39836 452640 39856
rect 452524 39796 452640 39836
rect 452544 39776 452640 39796
rect 0 39332 96 39352
rect 452544 39332 452640 39352
rect 0 39292 116 39332
rect 452524 39292 452640 39332
rect 0 39272 96 39292
rect 452544 39272 452640 39292
rect 452544 38828 452640 38848
rect 452524 38788 452640 38828
rect 452544 38768 452640 38788
rect 0 38324 96 38344
rect 452544 38324 452640 38344
rect 0 38284 116 38324
rect 452524 38284 452640 38324
rect 0 38264 96 38284
rect 452544 38264 452640 38284
rect 452544 37820 452640 37840
rect 452524 37780 452640 37820
rect 452544 37760 452640 37780
rect 0 37316 96 37336
rect 452544 37316 452640 37336
rect 0 37276 116 37316
rect 452524 37276 452640 37316
rect 0 37256 96 37276
rect 452544 37256 452640 37276
rect 452544 36812 452640 36832
rect 452524 36772 452640 36812
rect 452544 36752 452640 36772
rect 0 36308 96 36328
rect 452544 36308 452640 36328
rect 0 36268 116 36308
rect 452524 36268 452640 36308
rect 0 36248 96 36268
rect 452544 36248 452640 36268
rect 452544 35804 452640 35824
rect 452524 35764 452640 35804
rect 452544 35744 452640 35764
rect 0 35300 96 35320
rect 452544 35300 452640 35320
rect 0 35260 116 35300
rect 452524 35260 452640 35300
rect 0 35240 96 35260
rect 452544 35240 452640 35260
rect 452544 34796 452640 34816
rect 452524 34756 452640 34796
rect 452544 34736 452640 34756
rect 0 34292 96 34312
rect 452544 34292 452640 34312
rect 0 34252 116 34292
rect 452524 34252 452640 34292
rect 0 34232 96 34252
rect 452544 34232 452640 34252
rect 452544 33788 452640 33808
rect 452524 33748 452640 33788
rect 452544 33728 452640 33748
rect 0 33284 96 33304
rect 452544 33284 452640 33304
rect 0 33244 116 33284
rect 452524 33244 452640 33284
rect 0 33224 96 33244
rect 452544 33224 452640 33244
rect 452544 32780 452640 32800
rect 452524 32740 452640 32780
rect 452544 32720 452640 32740
rect 0 32276 96 32296
rect 452544 32276 452640 32296
rect 0 32236 116 32276
rect 452524 32236 452640 32276
rect 0 32216 96 32236
rect 452544 32216 452640 32236
rect 452544 31772 452640 31792
rect 452524 31732 452640 31772
rect 452544 31712 452640 31732
rect 0 31268 96 31288
rect 452544 31268 452640 31288
rect 0 31228 116 31268
rect 452524 31228 452640 31268
rect 0 31208 96 31228
rect 452544 31208 452640 31228
rect 452544 30764 452640 30784
rect 452524 30724 452640 30764
rect 452544 30704 452640 30724
rect 0 30260 96 30280
rect 452544 30260 452640 30280
rect 0 30220 116 30260
rect 452524 30220 452640 30260
rect 0 30200 96 30220
rect 452544 30200 452640 30220
rect 452544 29756 452640 29776
rect 452524 29716 452640 29756
rect 452544 29696 452640 29716
rect 0 29252 96 29272
rect 452544 29252 452640 29272
rect 0 29212 116 29252
rect 452524 29212 452640 29252
rect 0 29192 96 29212
rect 452544 29192 452640 29212
rect 452544 28748 452640 28768
rect 452524 28708 452640 28748
rect 452544 28688 452640 28708
rect 0 28244 96 28264
rect 452544 28244 452640 28264
rect 0 28204 116 28244
rect 452524 28204 452640 28244
rect 0 28184 96 28204
rect 452544 28184 452640 28204
rect 452544 27740 452640 27760
rect 452524 27700 452640 27740
rect 452544 27680 452640 27700
rect 0 27236 96 27256
rect 452544 27236 452640 27256
rect 0 27196 116 27236
rect 452524 27196 452640 27236
rect 0 27176 96 27196
rect 452544 27176 452640 27196
rect 452544 26732 452640 26752
rect 452524 26692 452640 26732
rect 452544 26672 452640 26692
rect 0 26228 96 26248
rect 452544 26228 452640 26248
rect 0 26188 116 26228
rect 452524 26188 452640 26228
rect 0 26168 96 26188
rect 452544 26168 452640 26188
rect 452544 25724 452640 25744
rect 452524 25684 452640 25724
rect 452544 25664 452640 25684
rect 0 25220 96 25240
rect 452544 25220 452640 25240
rect 0 25180 116 25220
rect 452524 25180 452640 25220
rect 0 25160 96 25180
rect 452544 25160 452640 25180
rect 452544 24716 452640 24736
rect 452524 24676 452640 24716
rect 452544 24656 452640 24676
rect 0 24212 96 24232
rect 452544 24212 452640 24232
rect 0 24172 116 24212
rect 452524 24172 452640 24212
rect 0 24152 96 24172
rect 452544 24152 452640 24172
rect 452544 23708 452640 23728
rect 452524 23668 452640 23708
rect 452544 23648 452640 23668
rect 0 23204 96 23224
rect 452544 23204 452640 23224
rect 0 23164 116 23204
rect 452524 23164 452640 23204
rect 0 23144 96 23164
rect 452544 23144 452640 23164
rect 452544 22700 452640 22720
rect 452524 22660 452640 22700
rect 452544 22640 452640 22660
rect 0 22196 96 22216
rect 452544 22196 452640 22216
rect 0 22156 116 22196
rect 452524 22156 452640 22196
rect 0 22136 96 22156
rect 452544 22136 452640 22156
rect 452544 21692 452640 21712
rect 452524 21652 452640 21692
rect 452544 21632 452640 21652
rect 0 21188 96 21208
rect 452544 21188 452640 21208
rect 0 21148 116 21188
rect 452524 21148 452640 21188
rect 0 21128 96 21148
rect 452544 21128 452640 21148
rect 452544 20684 452640 20704
rect 452524 20644 452640 20684
rect 452544 20624 452640 20644
rect 0 20180 96 20200
rect 452544 20180 452640 20200
rect 0 20140 116 20180
rect 452524 20140 452640 20180
rect 0 20120 96 20140
rect 452544 20120 452640 20140
rect 452544 19676 452640 19696
rect 452524 19636 452640 19676
rect 452544 19616 452640 19636
rect 0 19172 96 19192
rect 452544 19172 452640 19192
rect 0 19132 116 19172
rect 452524 19132 452640 19172
rect 0 19112 96 19132
rect 452544 19112 452640 19132
rect 452544 18668 452640 18688
rect 452524 18628 452640 18668
rect 452544 18608 452640 18628
rect 0 18164 96 18184
rect 452544 18164 452640 18184
rect 0 18124 116 18164
rect 452524 18124 452640 18164
rect 0 18104 96 18124
rect 452544 18104 452640 18124
rect 452544 17660 452640 17680
rect 452524 17620 452640 17660
rect 452544 17600 452640 17620
rect 0 17156 96 17176
rect 452544 17156 452640 17176
rect 0 17116 116 17156
rect 452524 17116 452640 17156
rect 0 17096 96 17116
rect 452544 17096 452640 17116
rect 452544 16652 452640 16672
rect 452524 16612 452640 16652
rect 452544 16592 452640 16612
rect 0 16148 96 16168
rect 0 16108 116 16148
rect 0 16088 96 16108
rect 0 15140 96 15160
rect 0 15100 116 15140
rect 0 15080 96 15100
rect 96 13712 136 14092
rect 28 13672 136 13712
rect 28 13460 68 13672
rect 28 13420 186 13460
rect 0 13292 96 13312
rect 146 13292 186 13420
rect 0 13252 186 13292
rect 0 13232 96 13252
rect 0 11864 96 11884
rect 0 11824 13844 11864
rect 0 11804 96 11824
rect 0 11528 96 11548
rect 0 11488 13844 11528
rect 0 11468 96 11488
rect 0 11192 96 11212
rect 0 11152 13844 11192
rect 0 11132 96 11152
rect 0 10856 96 10876
rect 0 10816 13844 10856
rect 0 10796 96 10816
rect 0 10520 96 10540
rect 0 10480 13844 10520
rect 0 10460 96 10480
rect 0 10184 96 10204
rect 0 10144 13844 10184
rect 0 10124 96 10144
rect 0 9848 96 9868
rect 0 9808 13844 9848
rect 0 9788 96 9808
rect 0 9512 96 9532
rect 0 9472 13844 9512
rect 0 9452 96 9472
rect 0 9176 96 9196
rect 0 9136 13844 9176
rect 0 9116 96 9136
rect 0 8840 96 8860
rect 0 8800 13844 8840
rect 0 8780 96 8800
rect 0 8504 96 8524
rect 0 8464 13844 8504
rect 0 8444 96 8464
rect 0 8168 96 8188
rect 0 8128 13844 8168
rect 0 8108 96 8128
rect 0 7832 96 7852
rect 0 7792 13844 7832
rect 0 7772 96 7792
rect 0 7496 96 7516
rect 0 7456 13844 7496
rect 0 7436 96 7456
rect 0 7160 96 7180
rect 0 7120 13844 7160
rect 0 7100 96 7120
rect 0 6824 96 6844
rect 0 6784 13844 6824
rect 0 6764 96 6784
rect 0 6488 96 6508
rect 0 6448 13844 6488
rect 0 6428 96 6448
rect 0 6152 96 6172
rect 0 6112 13844 6152
rect 0 6092 96 6112
rect 0 5816 96 5836
rect 0 5776 13844 5816
rect 0 5756 96 5776
rect 0 5480 96 5500
rect 0 5440 13844 5480
rect 0 5420 96 5440
rect 0 5144 96 5164
rect 0 5104 13844 5144
rect 0 5084 96 5104
rect 0 4808 96 4828
rect 0 4768 13844 4808
rect 0 4748 96 4768
rect 0 4472 96 4492
rect 0 4432 13844 4472
rect 0 4412 96 4432
rect 0 4136 96 4156
rect 0 4096 13844 4136
rect 0 4076 96 4096
rect 0 3800 96 3820
rect 0 3760 13844 3800
rect 0 3740 96 3760
rect 0 3464 96 3484
rect 0 3424 13844 3464
rect 0 3404 96 3424
rect 0 3128 96 3148
rect 0 3088 13844 3128
rect 0 3068 96 3088
rect 0 2792 96 2812
rect 0 2752 13844 2792
rect 0 2732 96 2752
rect 0 2456 96 2476
rect 0 2416 13844 2456
rect 0 2396 96 2416
rect 0 2120 96 2140
rect 0 2080 13844 2120
rect 0 2060 96 2080
rect 0 1784 96 1804
rect 0 1744 13844 1784
rect 0 1724 96 1744
rect 0 1448 96 1468
rect 0 1408 13844 1448
rect 0 1388 96 1408
<< metal3 >>
rect 17336 702240 17416 702336
rect 18488 702240 18568 702336
rect 19640 702240 19720 702336
rect 20792 702240 20872 702336
rect 21944 702240 22024 702336
rect 23096 702240 23176 702336
rect 24248 702240 24328 702336
rect 25400 702240 25480 702336
rect 26552 702240 26632 702336
rect 27704 702240 27784 702336
rect 28856 702240 28936 702336
rect 30008 702240 30088 702336
rect 31160 702240 31240 702336
rect 32312 702240 32392 702336
rect 63704 702240 63784 702336
rect 64856 702240 64936 702336
rect 66008 702240 66088 702336
rect 67160 702240 67240 702336
rect 68312 702240 68392 702336
rect 69464 702240 69544 702336
rect 70616 702240 70696 702336
rect 71768 702240 71848 702336
rect 72920 702240 73000 702336
rect 74072 702240 74152 702336
rect 75224 702240 75304 702336
rect 76376 702240 76456 702336
rect 77528 702240 77608 702336
rect 78680 702240 78760 702336
rect 17356 702220 17396 702240
rect 18508 702220 18548 702240
rect 19660 702220 19700 702240
rect 20812 702220 20852 702240
rect 21964 702220 22004 702240
rect 23116 702220 23156 702240
rect 24268 702220 24308 702240
rect 25420 702220 25460 702240
rect 26572 702220 26612 702240
rect 27724 702220 27764 702240
rect 28876 702220 28916 702240
rect 30028 702220 30068 702240
rect 31180 702220 31220 702240
rect 32332 702220 32372 702240
rect 63724 702220 63764 702240
rect 64876 702220 64916 702240
rect 66028 702220 66068 702240
rect 67180 702220 67220 702240
rect 68332 702220 68372 702240
rect 69484 702220 69524 702240
rect 70636 702220 70676 702240
rect 71788 702220 71828 702240
rect 72940 702220 72980 702240
rect 74092 702220 74132 702240
rect 75244 702220 75284 702240
rect 76396 702220 76436 702240
rect 77548 702220 77588 702240
rect 78700 702220 78740 702240
rect 1132 104 1172 12704
rect 1112 64 1132 80
rect 1708 80 1748 12704
rect 2284 80 2324 12704
rect 2860 80 2900 12704
rect 3436 80 3476 12704
rect 4012 80 4052 12704
rect 4588 80 4628 12704
rect 5164 80 5204 12704
rect 5740 80 5780 12704
rect 6316 80 6356 12704
rect 6892 80 6932 12704
rect 7468 80 7508 12704
rect 8044 80 8084 12704
rect 8620 80 8660 12704
rect 9196 80 9236 12704
rect 9772 80 9812 12704
rect 10348 80 10388 12704
rect 10924 80 10964 12704
rect 11500 80 11540 12704
rect 12076 80 12116 12704
rect 12652 80 12692 12704
rect 15820 104 15860 860
rect 1172 64 1192 80
rect 1112 0 1192 64
rect 1688 0 1768 80
rect 2264 0 2344 80
rect 2840 0 2920 80
rect 3416 0 3496 80
rect 3992 0 4072 80
rect 4568 0 4648 80
rect 5144 0 5224 80
rect 5720 0 5800 80
rect 6296 0 6376 80
rect 6872 0 6952 80
rect 7448 0 7528 80
rect 8024 0 8104 80
rect 8600 0 8680 80
rect 9176 0 9256 80
rect 9752 0 9832 80
rect 10328 0 10408 80
rect 10904 0 10984 80
rect 11480 0 11560 80
rect 12056 0 12136 80
rect 12632 0 12712 80
rect 17932 96 17972 860
rect 20044 96 20084 860
rect 22156 96 22196 860
rect 24268 96 24308 860
rect 26380 96 26420 860
rect 28492 96 28532 860
rect 30604 96 30644 860
rect 32716 96 32756 860
rect 34828 96 34868 860
rect 36940 96 36980 860
rect 39052 96 39092 860
rect 41164 96 41204 860
rect 43276 96 43316 860
rect 45388 96 45428 860
rect 47500 96 47540 860
rect 49612 96 49652 860
rect 51724 96 51764 860
rect 53836 96 53876 860
rect 55948 96 55988 860
rect 58060 96 58100 860
rect 62572 96 62612 860
rect 64108 96 64148 860
rect 65644 96 65684 860
rect 67180 96 67220 860
rect 68716 96 68756 860
rect 70252 96 70292 860
rect 71788 96 71828 860
rect 73324 104 73364 860
rect 15820 55 15860 64
rect 17912 0 17992 96
rect 20024 0 20104 96
rect 22136 0 22216 96
rect 24248 0 24328 96
rect 26360 0 26440 96
rect 28472 0 28552 96
rect 30584 0 30664 96
rect 32696 0 32776 96
rect 34808 0 34888 96
rect 36920 0 37000 96
rect 39032 0 39112 96
rect 41144 0 41224 96
rect 43256 0 43336 96
rect 45368 0 45448 96
rect 47480 0 47560 96
rect 49592 0 49672 96
rect 51704 0 51784 96
rect 53816 0 53896 96
rect 55928 0 56008 96
rect 58040 0 58120 96
rect 62552 0 62632 96
rect 64088 0 64168 96
rect 65624 0 65704 96
rect 67160 0 67240 96
rect 68696 0 68776 96
rect 70232 0 70312 96
rect 71768 0 71848 96
rect 74860 96 74900 860
rect 76396 96 76436 860
rect 77932 96 77972 860
rect 79468 96 79508 860
rect 81004 96 81044 860
rect 82540 96 82580 860
rect 84076 96 84116 860
rect 85612 96 85652 860
rect 87148 96 87188 860
rect 88684 96 88724 860
rect 90220 96 90260 860
rect 91756 96 91796 860
rect 93292 96 93332 860
rect 94828 96 94868 860
rect 96364 96 96404 860
rect 97900 96 97940 860
rect 99436 96 99476 860
rect 100972 96 101012 860
rect 102508 96 102548 860
rect 104044 96 104084 860
rect 107980 96 108020 860
rect 109708 96 109748 860
rect 111436 96 111476 860
rect 113164 96 113204 860
rect 114892 96 114932 860
rect 116620 104 116660 860
rect 73324 55 73364 64
rect 74840 0 74920 96
rect 76376 0 76456 96
rect 77912 0 77992 96
rect 79448 0 79528 96
rect 80984 0 81064 96
rect 82520 0 82600 96
rect 84056 0 84136 96
rect 85592 0 85672 96
rect 87128 0 87208 96
rect 88664 0 88744 96
rect 90200 0 90280 96
rect 91736 0 91816 96
rect 93272 0 93352 96
rect 94808 0 94888 96
rect 96344 0 96424 96
rect 97880 0 97960 96
rect 99416 0 99496 96
rect 100952 0 101032 96
rect 102488 0 102568 96
rect 104024 0 104104 96
rect 107960 0 108040 96
rect 109688 0 109768 96
rect 111416 0 111496 96
rect 113144 0 113224 96
rect 114872 0 114952 96
rect 118348 96 118388 860
rect 120076 96 120116 860
rect 121804 96 121844 860
rect 123532 96 123572 860
rect 125260 96 125300 860
rect 126988 96 127028 860
rect 128716 96 128756 860
rect 130444 96 130484 860
rect 132172 96 132212 860
rect 133900 96 133940 860
rect 135628 96 135668 860
rect 137356 96 137396 860
rect 139084 96 139124 860
rect 140812 96 140852 860
rect 142540 96 142580 860
rect 144268 96 144308 860
rect 145996 96 146036 860
rect 147724 96 147764 860
rect 149452 96 149492 860
rect 151180 96 151220 860
rect 154540 104 154580 860
rect 116620 55 116660 64
rect 118328 0 118408 96
rect 120056 0 120136 96
rect 121784 0 121864 96
rect 123512 0 123592 96
rect 125240 0 125320 96
rect 126968 0 127048 96
rect 128696 0 128776 96
rect 130424 0 130504 96
rect 132152 0 132232 96
rect 133880 0 133960 96
rect 135608 0 135688 96
rect 137336 0 137416 96
rect 139064 0 139144 96
rect 140792 0 140872 96
rect 142520 0 142600 96
rect 144248 0 144328 96
rect 145976 0 146056 96
rect 147704 0 147784 96
rect 149432 0 149512 96
rect 151160 0 151240 96
rect 157036 96 157076 860
rect 159532 96 159572 860
rect 162028 96 162068 860
rect 164524 96 164564 860
rect 167020 96 167060 860
rect 169516 96 169556 860
rect 172012 96 172052 860
rect 174508 96 174548 860
rect 177004 96 177044 860
rect 179500 96 179540 860
rect 181996 96 182036 860
rect 184492 96 184532 860
rect 186988 96 187028 860
rect 189484 96 189524 860
rect 191980 96 192020 860
rect 194476 96 194516 860
rect 196972 96 197012 860
rect 199468 96 199508 860
rect 201964 96 202004 860
rect 204460 96 204500 860
rect 209356 96 209396 860
rect 210124 96 210164 860
rect 210892 96 210932 860
rect 211660 96 211700 860
rect 212428 96 212468 860
rect 213196 96 213236 860
rect 213964 96 214004 860
rect 214732 96 214772 860
rect 215500 96 215540 860
rect 216268 96 216308 860
rect 217036 96 217076 860
rect 217804 96 217844 860
rect 218572 96 218612 860
rect 219340 96 219380 860
rect 220108 96 220148 860
rect 220876 96 220916 860
rect 221644 96 221684 860
rect 222412 96 222452 860
rect 223180 96 223220 860
rect 223948 96 223988 860
rect 224716 96 224756 860
rect 225484 96 225524 860
rect 226252 96 226292 860
rect 227020 96 227060 860
rect 227788 96 227828 860
rect 228556 96 228596 860
rect 229324 96 229364 860
rect 230092 96 230132 860
rect 230860 96 230900 860
rect 231628 96 231668 860
rect 232396 96 232436 860
rect 233164 96 233204 860
rect 233932 104 233972 860
rect 154540 55 154580 64
rect 157016 0 157096 96
rect 159512 0 159592 96
rect 162008 0 162088 96
rect 164504 0 164584 96
rect 167000 0 167080 96
rect 169496 0 169576 96
rect 171992 0 172072 96
rect 174488 0 174568 96
rect 176984 0 177064 96
rect 179480 0 179560 96
rect 181976 0 182056 96
rect 184472 0 184552 96
rect 186968 0 187048 96
rect 189464 0 189544 96
rect 191960 0 192040 96
rect 194456 0 194536 96
rect 196952 0 197032 96
rect 199448 0 199528 96
rect 201944 0 202024 96
rect 204440 0 204520 96
rect 209336 0 209416 96
rect 210104 0 210184 96
rect 210872 0 210952 96
rect 211640 0 211720 96
rect 212408 0 212488 96
rect 213176 0 213256 96
rect 213944 0 214024 96
rect 214712 0 214792 96
rect 215480 0 215560 96
rect 216248 0 216328 96
rect 217016 0 217096 96
rect 217784 0 217864 96
rect 218552 0 218632 96
rect 219320 0 219400 96
rect 220088 0 220168 96
rect 220856 0 220936 96
rect 221624 0 221704 96
rect 222392 0 222472 96
rect 223160 0 223240 96
rect 223928 0 224008 96
rect 224696 0 224776 96
rect 225464 0 225544 96
rect 226232 0 226312 96
rect 227000 0 227080 96
rect 227768 0 227848 96
rect 228536 0 228616 96
rect 229304 0 229384 96
rect 230072 0 230152 96
rect 230840 0 230920 96
rect 231608 0 231688 96
rect 232376 0 232456 96
rect 233144 0 233224 96
rect 234700 96 234740 860
rect 235468 96 235508 860
rect 236236 96 236276 860
rect 237004 96 237044 860
rect 237772 96 237812 860
rect 238540 96 238580 860
rect 239308 96 239348 860
rect 240076 96 240116 860
rect 240844 96 240884 860
rect 241612 96 241652 860
rect 242380 96 242420 860
rect 243148 96 243188 860
rect 243916 96 243956 860
rect 244684 96 244724 860
rect 245452 96 245492 860
rect 246220 96 246260 860
rect 246988 96 247028 860
rect 247756 96 247796 860
rect 248524 96 248564 860
rect 249292 96 249332 860
rect 255724 96 255764 860
rect 256492 96 256532 860
rect 257260 96 257300 860
rect 258028 96 258068 860
rect 258796 96 258836 860
rect 259564 96 259604 860
rect 260332 96 260372 860
rect 261100 96 261140 860
rect 261868 96 261908 860
rect 262636 96 262676 860
rect 263404 96 263444 860
rect 264172 96 264212 860
rect 264940 96 264980 860
rect 265708 96 265748 860
rect 266476 96 266516 860
rect 267244 96 267284 860
rect 268012 96 268052 860
rect 268780 96 268820 860
rect 269548 96 269588 860
rect 270316 96 270356 860
rect 271084 96 271124 860
rect 271852 96 271892 860
rect 272620 96 272660 860
rect 273388 96 273428 860
rect 274156 96 274196 860
rect 274924 96 274964 860
rect 275692 96 275732 860
rect 276460 96 276500 860
rect 277228 96 277268 860
rect 277996 96 278036 860
rect 278764 96 278804 860
rect 279532 96 279572 860
rect 280300 104 280340 860
rect 233932 55 233972 64
rect 234680 0 234760 96
rect 235448 0 235528 96
rect 236216 0 236296 96
rect 236984 0 237064 96
rect 237752 0 237832 96
rect 238520 0 238600 96
rect 239288 0 239368 96
rect 240056 0 240136 96
rect 240824 0 240904 96
rect 241592 0 241672 96
rect 242360 0 242440 96
rect 243128 0 243208 96
rect 243896 0 243976 96
rect 244664 0 244744 96
rect 245432 0 245512 96
rect 246200 0 246280 96
rect 246968 0 247048 96
rect 247736 0 247816 96
rect 248504 0 248584 96
rect 249272 0 249352 96
rect 255704 0 255784 96
rect 256472 0 256552 96
rect 257240 0 257320 96
rect 258008 0 258088 96
rect 258776 0 258856 96
rect 259544 0 259624 96
rect 260312 0 260392 96
rect 261080 0 261160 96
rect 261848 0 261928 96
rect 262616 0 262696 96
rect 263384 0 263464 96
rect 264152 0 264232 96
rect 264920 0 265000 96
rect 265688 0 265768 96
rect 266456 0 266536 96
rect 267224 0 267304 96
rect 267992 0 268072 96
rect 268760 0 268840 96
rect 269528 0 269608 96
rect 270296 0 270376 96
rect 271064 0 271144 96
rect 271832 0 271912 96
rect 272600 0 272680 96
rect 273368 0 273448 96
rect 274136 0 274216 96
rect 274904 0 274984 96
rect 275672 0 275752 96
rect 276440 0 276520 96
rect 277208 0 277288 96
rect 277976 0 278056 96
rect 278744 0 278824 96
rect 279512 0 279592 96
rect 281068 96 281108 860
rect 281836 96 281876 860
rect 282604 96 282644 860
rect 283372 96 283412 860
rect 284140 96 284180 860
rect 284908 96 284948 860
rect 285676 96 285716 860
rect 286444 96 286484 860
rect 287212 96 287252 860
rect 287980 96 288020 860
rect 288748 96 288788 860
rect 289516 96 289556 860
rect 290284 96 290324 860
rect 291052 96 291092 860
rect 291820 96 291860 860
rect 292588 96 292628 860
rect 293356 96 293396 860
rect 294124 96 294164 860
rect 294892 96 294932 860
rect 295660 96 295700 860
rect 301132 104 301172 860
rect 280300 55 280340 64
rect 281048 0 281128 96
rect 281816 0 281896 96
rect 282584 0 282664 96
rect 283352 0 283432 96
rect 284120 0 284200 96
rect 284888 0 284968 96
rect 285656 0 285736 96
rect 286424 0 286504 96
rect 287192 0 287272 96
rect 287960 0 288040 96
rect 288728 0 288808 96
rect 289496 0 289576 96
rect 290264 0 290344 96
rect 291032 0 291112 96
rect 291800 0 291880 96
rect 292568 0 292648 96
rect 293336 0 293416 96
rect 294104 0 294184 96
rect 294872 0 294952 96
rect 295640 0 295720 96
rect 302860 96 302900 860
rect 304588 96 304628 860
rect 306316 96 306356 860
rect 308044 96 308084 860
rect 309772 96 309812 860
rect 311500 96 311540 860
rect 313228 96 313268 860
rect 314956 96 314996 860
rect 316684 96 316724 860
rect 318412 96 318452 860
rect 320140 96 320180 860
rect 321868 96 321908 860
rect 323596 96 323636 860
rect 325324 96 325364 860
rect 327052 96 327092 860
rect 328780 96 328820 860
rect 330508 96 330548 860
rect 332236 96 332276 860
rect 333964 96 334004 860
rect 335692 96 335732 860
rect 341356 96 341396 860
rect 342124 96 342164 860
rect 342892 96 342932 860
rect 343660 96 343700 860
rect 344428 96 344468 860
rect 345196 96 345236 860
rect 345964 96 346004 860
rect 346732 96 346772 860
rect 347500 96 347540 860
rect 348268 96 348308 860
rect 349036 96 349076 860
rect 349804 96 349844 860
rect 350572 96 350612 860
rect 351340 96 351380 860
rect 352108 96 352148 860
rect 352876 96 352916 860
rect 353644 96 353684 860
rect 354412 96 354452 860
rect 355180 96 355220 860
rect 355948 96 355988 860
rect 356716 96 356756 860
rect 357484 96 357524 860
rect 358252 96 358292 860
rect 359020 96 359060 860
rect 359788 96 359828 860
rect 360556 96 360596 860
rect 361324 96 361364 860
rect 362092 96 362132 860
rect 362860 96 362900 860
rect 363628 96 363668 860
rect 364396 96 364436 860
rect 365164 96 365204 860
rect 365932 104 365972 860
rect 301132 55 301172 64
rect 302840 0 302920 96
rect 304568 0 304648 96
rect 306296 0 306376 96
rect 308024 0 308104 96
rect 309752 0 309832 96
rect 311480 0 311560 96
rect 313208 0 313288 96
rect 314936 0 315016 96
rect 316664 0 316744 96
rect 318392 0 318472 96
rect 320120 0 320200 96
rect 321848 0 321928 96
rect 323576 0 323656 96
rect 325304 0 325384 96
rect 327032 0 327112 96
rect 328760 0 328840 96
rect 330488 0 330568 96
rect 332216 0 332296 96
rect 333944 0 334024 96
rect 335672 0 335752 96
rect 341336 0 341416 96
rect 342104 0 342184 96
rect 342872 0 342952 96
rect 343640 0 343720 96
rect 344408 0 344488 96
rect 345176 0 345256 96
rect 345944 0 346024 96
rect 346712 0 346792 96
rect 347480 0 347560 96
rect 348248 0 348328 96
rect 349016 0 349096 96
rect 349784 0 349864 96
rect 350552 0 350632 96
rect 351320 0 351400 96
rect 352088 0 352168 96
rect 352856 0 352936 96
rect 353624 0 353704 96
rect 354392 0 354472 96
rect 355160 0 355240 96
rect 355928 0 356008 96
rect 356696 0 356776 96
rect 357464 0 357544 96
rect 358232 0 358312 96
rect 359000 0 359080 96
rect 359768 0 359848 96
rect 360536 0 360616 96
rect 361304 0 361384 96
rect 362072 0 362152 96
rect 362840 0 362920 96
rect 363608 0 363688 96
rect 364376 0 364456 96
rect 365144 0 365224 96
rect 366700 96 366740 860
rect 367468 96 367508 860
rect 368236 96 368276 860
rect 369004 96 369044 860
rect 369772 96 369812 860
rect 370540 96 370580 860
rect 371308 96 371348 860
rect 372076 96 372116 860
rect 372844 96 372884 860
rect 373612 96 373652 860
rect 374380 96 374420 860
rect 375148 96 375188 860
rect 375916 96 375956 860
rect 376684 96 376724 860
rect 377452 96 377492 860
rect 378220 96 378260 860
rect 378988 96 379028 860
rect 379756 96 379796 860
rect 380524 96 380564 860
rect 381292 96 381332 860
rect 387724 96 387764 860
rect 388492 96 388532 860
rect 389260 96 389300 860
rect 390028 96 390068 860
rect 390796 96 390836 860
rect 391564 96 391604 860
rect 392332 96 392372 860
rect 393100 96 393140 860
rect 393868 96 393908 860
rect 394636 96 394676 860
rect 395404 96 395444 860
rect 396172 96 396212 860
rect 396940 96 396980 860
rect 397708 96 397748 860
rect 398476 96 398516 860
rect 399244 96 399284 860
rect 400012 96 400052 860
rect 400780 96 400820 860
rect 401548 96 401588 860
rect 402316 96 402356 860
rect 403084 96 403124 860
rect 403852 96 403892 860
rect 404620 96 404660 860
rect 405388 96 405428 860
rect 406156 96 406196 860
rect 406924 96 406964 860
rect 407692 96 407732 860
rect 408460 96 408500 860
rect 409228 96 409268 860
rect 409996 96 410036 860
rect 410764 96 410804 860
rect 411532 96 411572 860
rect 412300 104 412340 860
rect 365932 55 365972 64
rect 366680 0 366760 96
rect 367448 0 367528 96
rect 368216 0 368296 96
rect 368984 0 369064 96
rect 369752 0 369832 96
rect 370520 0 370600 96
rect 371288 0 371368 96
rect 372056 0 372136 96
rect 372824 0 372904 96
rect 373592 0 373672 96
rect 374360 0 374440 96
rect 375128 0 375208 96
rect 375896 0 375976 96
rect 376664 0 376744 96
rect 377432 0 377512 96
rect 378200 0 378280 96
rect 378968 0 379048 96
rect 379736 0 379816 96
rect 380504 0 380584 96
rect 381272 0 381352 96
rect 387704 0 387784 96
rect 388472 0 388552 96
rect 389240 0 389320 96
rect 390008 0 390088 96
rect 390776 0 390856 96
rect 391544 0 391624 96
rect 392312 0 392392 96
rect 393080 0 393160 96
rect 393848 0 393928 96
rect 394616 0 394696 96
rect 395384 0 395464 96
rect 396152 0 396232 96
rect 396920 0 397000 96
rect 397688 0 397768 96
rect 398456 0 398536 96
rect 399224 0 399304 96
rect 399992 0 400072 96
rect 400760 0 400840 96
rect 401528 0 401608 96
rect 402296 0 402376 96
rect 403064 0 403144 96
rect 403832 0 403912 96
rect 404600 0 404680 96
rect 405368 0 405448 96
rect 406136 0 406216 96
rect 406904 0 406984 96
rect 407672 0 407752 96
rect 408440 0 408520 96
rect 409208 0 409288 96
rect 409976 0 410056 96
rect 410744 0 410824 96
rect 411512 0 411592 96
rect 413068 96 413108 860
rect 413836 96 413876 860
rect 414604 96 414644 860
rect 415372 96 415412 860
rect 416140 96 416180 860
rect 416908 96 416948 860
rect 417676 96 417716 860
rect 418444 96 418484 860
rect 419212 96 419252 860
rect 419980 96 420020 860
rect 420748 96 420788 860
rect 421516 96 421556 860
rect 422284 96 422324 860
rect 423052 96 423092 860
rect 423820 96 423860 860
rect 424588 96 424628 860
rect 425356 96 425396 860
rect 426124 96 426164 860
rect 426892 96 426932 860
rect 427660 96 427700 860
rect 431980 104 432020 860
rect 412300 55 412340 64
rect 413048 0 413128 96
rect 413816 0 413896 96
rect 414584 0 414664 96
rect 415352 0 415432 96
rect 416120 0 416200 96
rect 416888 0 416968 96
rect 417656 0 417736 96
rect 418424 0 418504 96
rect 419192 0 419272 96
rect 419960 0 420040 96
rect 420728 0 420808 96
rect 421496 0 421576 96
rect 422264 0 422344 96
rect 423032 0 423112 96
rect 423800 0 423880 96
rect 424568 0 424648 96
rect 425336 0 425416 96
rect 426104 0 426184 96
rect 426872 0 426952 96
rect 427640 0 427720 96
rect 432940 80 432980 860
rect 433900 80 433940 860
rect 434860 80 434900 860
rect 435820 80 435860 860
rect 436780 80 436820 860
rect 437740 80 437780 860
rect 438700 80 438740 860
rect 439660 80 439700 860
rect 440620 80 440660 860
rect 441580 80 441620 860
rect 442540 80 442580 860
rect 443500 80 443540 860
rect 444460 80 444500 860
rect 445420 80 445460 860
rect 446380 80 446420 860
rect 447340 80 447380 860
rect 448300 80 448340 860
rect 449260 80 449300 860
rect 450220 80 450260 860
rect 451180 80 451220 860
rect 431980 55 432020 64
rect 432920 0 433000 80
rect 433880 0 433960 80
rect 434840 0 434920 80
rect 435800 0 435880 80
rect 436760 0 436840 80
rect 437720 0 437800 80
rect 438680 0 438760 80
rect 439640 0 439720 80
rect 440600 0 440680 80
rect 441560 0 441640 80
rect 442520 0 442600 80
rect 443480 0 443560 80
rect 444440 0 444520 80
rect 445400 0 445480 80
rect 446360 0 446440 80
rect 447320 0 447400 80
rect 448280 0 448360 80
rect 449240 0 449320 80
rect 450200 0 450280 80
rect 451160 0 451240 80
<< via3 >>
rect 1132 64 1172 104
rect 15820 64 15860 104
rect 73324 64 73364 104
rect 116620 64 116660 104
rect 154540 64 154580 104
rect 233932 64 233972 104
rect 280300 64 280340 104
rect 301132 64 301172 104
rect 365932 64 365972 104
rect 412300 64 412340 104
rect 431980 64 432020 104
<< metal4 >>
rect 1123 64 1132 104
rect 1172 64 15820 104
rect 15860 64 73324 104
rect 73364 64 116620 104
rect 116660 64 154540 104
rect 154580 64 233932 104
rect 233972 64 280300 104
rect 280340 64 301132 104
rect 301172 64 365932 104
rect 365972 64 412300 104
rect 412340 64 431980 104
rect 432020 64 432029 104
<< metal5 >>
rect 3748 840 4188 702240
rect 4988 840 5428 702240
rect 17476 840 17916 702240
rect 18716 840 19156 702240
rect 32596 840 33036 702240
rect 33836 840 34276 702240
rect 47716 840 48156 702240
rect 48956 840 49396 702240
rect 63844 840 64284 702240
rect 65084 840 65524 702240
rect 78964 840 79404 702240
rect 80204 840 80644 702240
rect 94084 840 94524 702240
rect 95324 840 95764 702240
rect 110212 840 110652 702240
rect 111452 840 111892 702240
rect 125332 840 125772 702240
rect 126572 840 127012 702240
rect 140452 840 140892 702240
rect 141692 840 142132 702240
rect 156580 840 157020 702240
rect 157820 840 158260 702240
rect 171700 840 172140 702240
rect 172940 840 173380 702240
rect 186820 840 187260 702240
rect 188060 840 188500 702240
rect 201940 840 202380 702240
rect 203180 840 203620 702240
rect 209860 840 210300 702240
rect 211100 840 211540 702240
rect 224980 840 225420 702240
rect 226220 840 226660 702240
rect 240100 840 240540 702240
rect 241340 840 241780 702240
rect 256228 840 256668 702240
rect 257468 840 257908 702240
rect 271348 840 271788 702240
rect 272588 840 273028 702240
rect 286468 840 286908 702240
rect 287708 840 288148 702240
rect 302596 840 303036 702240
rect 303836 840 304276 702240
rect 317716 840 318156 702240
rect 318956 840 319396 702240
rect 332836 840 333276 702240
rect 334076 840 334516 702240
rect 341860 840 342300 702240
rect 343100 840 343540 702240
rect 356980 840 357420 702240
rect 358220 840 358660 702240
rect 372100 840 372540 702240
rect 373340 840 373780 702240
rect 388228 840 388668 702240
rect 389468 840 389908 702240
rect 403348 840 403788 702240
rect 404588 840 405028 702240
rect 418468 840 418908 702240
rect 419708 840 420148 702240
rect 434596 840 435036 702240
rect 435836 840 436276 702240
rect 449716 840 450156 702240
use W_IO  Tile_X0Y1_W_IO
timestamp 0
transform 1 0 96 0 1 641676
box 0 0 1 1
use W_IO  Tile_X0Y2_W_IO
timestamp 0
transform 1 0 96 0 1 593292
box 0 0 1 1
use W_IO  Tile_X0Y3_W_IO
timestamp 0
transform 1 0 96 0 1 544908
box 0 0 1 1
use W_IO  Tile_X0Y4_W_IO
timestamp 0
transform 1 0 96 0 1 496524
box 0 0 1 1
use W_IO  Tile_X0Y5_W_IO
timestamp 0
transform 1 0 96 0 1 448140
box 0 0 1 1
use W_IO  Tile_X0Y6_W_IO
timestamp 0
transform 1 0 96 0 1 399756
box 0 0 1 1
use W_IO  Tile_X0Y7_W_IO
timestamp 0
transform 1 0 96 0 1 351372
box 0 0 1 1
use W_IO  Tile_X0Y8_W_IO
timestamp 0
transform 1 0 96 0 1 302988
box 0 0 1 1
use W_IO  Tile_X0Y9_W_IO
timestamp 0
transform 1 0 96 0 1 254604
box 0 0 1 1
use W_IO  Tile_X0Y10_W_IO
timestamp 0
transform 1 0 96 0 1 206220
box 0 0 1 1
use W_IO  Tile_X0Y11_W_IO
timestamp 0
transform 1 0 96 0 1 157836
box 0 0 1 1
use W_IO  Tile_X0Y12_W_IO
timestamp 0
transform 1 0 96 0 1 109452
box 0 0 1 1
use W_IO  Tile_X0Y13_W_IO
timestamp 0
transform 1 0 96 0 1 61068
box 0 0 1 1
use W_IO  Tile_X0Y14_W_IO
timestamp 0
transform 1 0 96 0 1 12684
box 0 0 1 1
use N_IO  Tile_X1Y0_N_IO
timestamp 0
transform 1 0 13824 0 1 690060
box 0 0 1 1
use LUT4AB  Tile_X1Y1_LUT4AB
timestamp 0
transform 1 0 13824 0 1 641676
box 0 0 1 1
use LUT4AB  Tile_X1Y2_LUT4AB
timestamp 0
transform 1 0 13824 0 1 593292
box 0 0 1 1
use LUT4AB  Tile_X1Y3_LUT4AB
timestamp 0
transform 1 0 13824 0 1 544908
box 0 0 1 1
use LUT4AB  Tile_X1Y4_LUT4AB
timestamp 0
transform 1 0 13824 0 1 496524
box 0 0 1 1
use LUT4AB  Tile_X1Y5_LUT4AB
timestamp 0
transform 1 0 13824 0 1 448140
box 0 0 1 1
use LUT4AB  Tile_X1Y6_LUT4AB
timestamp 0
transform 1 0 13824 0 1 399756
box 0 0 1 1
use LUT4AB  Tile_X1Y7_LUT4AB
timestamp 0
transform 1 0 13824 0 1 351372
box 0 0 1 1
use LUT4AB  Tile_X1Y8_LUT4AB
timestamp 0
transform 1 0 13824 0 1 302988
box 0 0 1 1
use LUT4AB  Tile_X1Y9_LUT4AB
timestamp 0
transform 1 0 13824 0 1 254604
box 0 0 1 1
use LUT4AB  Tile_X1Y10_LUT4AB
timestamp 0
transform 1 0 13824 0 1 206220
box 0 0 1 1
use LUT4AB  Tile_X1Y11_LUT4AB
timestamp 0
transform 1 0 13824 0 1 157836
box 0 0 1 1
use LUT4AB  Tile_X1Y12_LUT4AB
timestamp 0
transform 1 0 13824 0 1 109452
box 0 0 1 1
use LUT4AB  Tile_X1Y13_LUT4AB
timestamp 0
transform 1 0 13824 0 1 61068
box 0 0 1 1
use LUT4AB  Tile_X1Y14_LUT4AB
timestamp 0
transform 1 0 13824 0 1 12684
box 0 0 1 1
use S_term_single  Tile_X1Y15_S_term_single
timestamp 0
transform 1 0 13824 0 1 840
box 0 0 1 1
use N_IO  Tile_X2Y0_N_IO
timestamp 0
transform 1 0 60192 0 1 690060
box 0 0 1 1
use LUT4AB  Tile_X2Y1_LUT4AB
timestamp 0
transform 1 0 60192 0 1 641676
box 0 0 1 1
use LUT4AB  Tile_X2Y2_LUT4AB
timestamp 0
transform 1 0 60192 0 1 593292
box 0 0 1 1
use LUT4AB  Tile_X2Y3_LUT4AB
timestamp 0
transform 1 0 60192 0 1 544908
box 0 0 1 1
use LUT4AB  Tile_X2Y4_LUT4AB
timestamp 0
transform 1 0 60192 0 1 496524
box 0 0 1 1
use LUT4AB  Tile_X2Y5_LUT4AB
timestamp 0
transform 1 0 60192 0 1 448140
box 0 0 1 1
use LUT4AB  Tile_X2Y6_LUT4AB
timestamp 0
transform 1 0 60192 0 1 399756
box 0 0 1 1
use LUT4AB  Tile_X2Y7_LUT4AB
timestamp 0
transform 1 0 60192 0 1 351372
box 0 0 1 1
use LUT4AB  Tile_X2Y8_LUT4AB
timestamp 0
transform 1 0 60192 0 1 302988
box 0 0 1 1
use LUT4AB  Tile_X2Y9_LUT4AB
timestamp 0
transform 1 0 60192 0 1 254604
box 0 0 1 1
use LUT4AB  Tile_X2Y10_LUT4AB
timestamp 0
transform 1 0 60192 0 1 206220
box 0 0 1 1
use LUT4AB  Tile_X2Y11_LUT4AB
timestamp 0
transform 1 0 60192 0 1 157836
box 0 0 1 1
use LUT4AB  Tile_X2Y12_LUT4AB
timestamp 0
transform 1 0 60192 0 1 109452
box 0 0 1 1
use LUT4AB  Tile_X2Y13_LUT4AB
timestamp 0
transform 1 0 60192 0 1 61068
box 0 0 1 1
use LUT4AB  Tile_X2Y14_LUT4AB
timestamp 0
transform 1 0 60192 0 1 12684
box 0 0 1 1
use S_WARMBOOT  Tile_X2Y15_S_WARMBOOT
timestamp 0
transform 1 0 60192 0 1 840
box 0 0 1 1
use N_term_single  Tile_X3Y0_N_term_single
timestamp 0
transform 1 0 106560 0 1 690060
box 0 0 1 1
use LUT4AB  Tile_X3Y1_LUT4AB
timestamp 0
transform 1 0 106560 0 1 641676
box 0 0 1 1
use LUT4AB  Tile_X3Y2_LUT4AB
timestamp 0
transform 1 0 106560 0 1 593292
box 0 0 1 1
use LUT4AB  Tile_X3Y3_LUT4AB
timestamp 0
transform 1 0 106560 0 1 544908
box 0 0 1 1
use LUT4AB  Tile_X3Y4_LUT4AB
timestamp 0
transform 1 0 106560 0 1 496524
box 0 0 1 1
use LUT4AB  Tile_X3Y5_LUT4AB
timestamp 0
transform 1 0 106560 0 1 448140
box 0 0 1 1
use LUT4AB  Tile_X3Y6_LUT4AB
timestamp 0
transform 1 0 106560 0 1 399756
box 0 0 1 1
use LUT4AB  Tile_X3Y7_LUT4AB
timestamp 0
transform 1 0 106560 0 1 351372
box 0 0 1 1
use LUT4AB  Tile_X3Y8_LUT4AB
timestamp 0
transform 1 0 106560 0 1 302988
box 0 0 1 1
use LUT4AB  Tile_X3Y9_LUT4AB
timestamp 0
transform 1 0 106560 0 1 254604
box 0 0 1 1
use LUT4AB  Tile_X3Y10_LUT4AB
timestamp 0
transform 1 0 106560 0 1 206220
box 0 0 1 1
use LUT4AB  Tile_X3Y11_LUT4AB
timestamp 0
transform 1 0 106560 0 1 157836
box 0 0 1 1
use LUT4AB  Tile_X3Y12_LUT4AB
timestamp 0
transform 1 0 106560 0 1 109452
box 0 0 1 1
use LUT4AB  Tile_X3Y13_LUT4AB
timestamp 0
transform 1 0 106560 0 1 61068
box 0 0 1 1
use LUT4AB  Tile_X3Y14_LUT4AB
timestamp 0
transform 1 0 106560 0 1 12684
box 0 0 1 1
use S_CPU_IRQ  Tile_X3Y15_S_CPU_IRQ
timestamp 0
transform 1 0 106560 0 1 840
box 0 0 1 1
use N_term_single2  Tile_X4Y0_N_term_single2
timestamp 0
transform 1 0 152928 0 1 690060
box 0 0 1 1
use RegFile  Tile_X4Y1_RegFile
timestamp 0
transform 1 0 152928 0 1 641676
box 0 0 1 1
use RegFile  Tile_X4Y2_RegFile
timestamp 0
transform 1 0 152928 0 1 593292
box 0 0 1 1
use RegFile  Tile_X4Y3_RegFile
timestamp 0
transform 1 0 152928 0 1 544908
box 0 0 1 1
use RegFile  Tile_X4Y4_RegFile
timestamp 0
transform 1 0 152928 0 1 496524
box 0 0 1 1
use RegFile  Tile_X4Y5_RegFile
timestamp 0
transform 1 0 152928 0 1 448140
box 0 0 1 1
use RegFile  Tile_X4Y6_RegFile
timestamp 0
transform 1 0 152928 0 1 399756
box 0 0 1 1
use RegFile  Tile_X4Y7_RegFile
timestamp 0
transform 1 0 152928 0 1 351372
box 0 0 1 1
use RegFile  Tile_X4Y8_RegFile
timestamp 0
transform 1 0 152928 0 1 302988
box 0 0 1 1
use RegFile  Tile_X4Y9_RegFile
timestamp 0
transform 1 0 152928 0 1 254604
box 0 0 1 1
use RegFile  Tile_X4Y10_RegFile
timestamp 0
transform 1 0 152928 0 1 206220
box 0 0 1 1
use RegFile  Tile_X4Y11_RegFile
timestamp 0
transform 1 0 152928 0 1 157836
box 0 0 1 1
use RegFile  Tile_X4Y12_RegFile
timestamp 0
transform 1 0 152928 0 1 109452
box 0 0 1 1
use RegFile  Tile_X4Y13_RegFile
timestamp 0
transform 1 0 152928 0 1 61068
box 0 0 1 1
use RegFile  Tile_X4Y14_RegFile
timestamp 0
transform 1 0 152928 0 1 12684
box 0 0 1 1
use S_term_single2  Tile_X4Y15_S_term_single2
timestamp 0
transform 1 0 152928 0 1 840
box 0 0 1 1
use N_term_single  Tile_X5Y0_N_term_single
timestamp 0
transform 1 0 206208 0 1 690060
box 0 0 1 1
use LUT4AB  Tile_X5Y1_LUT4AB
timestamp 0
transform 1 0 206208 0 1 641676
box 0 0 1 1
use LUT4AB  Tile_X5Y2_LUT4AB
timestamp 0
transform 1 0 206208 0 1 593292
box 0 0 1 1
use LUT4AB  Tile_X5Y3_LUT4AB
timestamp 0
transform 1 0 206208 0 1 544908
box 0 0 1 1
use LUT4AB  Tile_X5Y4_LUT4AB
timestamp 0
transform 1 0 206208 0 1 496524
box 0 0 1 1
use LUT4AB  Tile_X5Y5_LUT4AB
timestamp 0
transform 1 0 206208 0 1 448140
box 0 0 1 1
use LUT4AB  Tile_X5Y6_LUT4AB
timestamp 0
transform 1 0 206208 0 1 399756
box 0 0 1 1
use LUT4AB  Tile_X5Y7_LUT4AB
timestamp 0
transform 1 0 206208 0 1 351372
box 0 0 1 1
use LUT4AB  Tile_X5Y8_LUT4AB
timestamp 0
transform 1 0 206208 0 1 302988
box 0 0 1 1
use LUT4AB  Tile_X5Y9_LUT4AB
timestamp 0
transform 1 0 206208 0 1 254604
box 0 0 1 1
use LUT4AB  Tile_X5Y10_LUT4AB
timestamp 0
transform 1 0 206208 0 1 206220
box 0 0 1 1
use LUT4AB  Tile_X5Y11_LUT4AB
timestamp 0
transform 1 0 206208 0 1 157836
box 0 0 1 1
use LUT4AB  Tile_X5Y12_LUT4AB
timestamp 0
transform 1 0 206208 0 1 109452
box 0 0 1 1
use LUT4AB  Tile_X5Y13_LUT4AB
timestamp 0
transform 1 0 206208 0 1 61068
box 0 0 1 1
use LUT4AB  Tile_X5Y14_LUT4AB
timestamp 0
transform 1 0 206208 0 1 12684
box 0 0 1 1
use S_CPU_IF  Tile_X5Y15_S_CPU_IF
timestamp 0
transform 1 0 206208 0 1 840
box 0 0 1 1
use N_term_single  Tile_X6Y0_N_term_single
timestamp 0
transform 1 0 252576 0 1 690060
box 0 0 1 1
use LUT4AB  Tile_X6Y1_LUT4AB
timestamp 0
transform 1 0 252576 0 1 641676
box 0 0 1 1
use LUT4AB  Tile_X6Y2_LUT4AB
timestamp 0
transform 1 0 252576 0 1 593292
box 0 0 1 1
use LUT4AB  Tile_X6Y3_LUT4AB
timestamp 0
transform 1 0 252576 0 1 544908
box 0 0 1 1
use LUT4AB  Tile_X6Y4_LUT4AB
timestamp 0
transform 1 0 252576 0 1 496524
box 0 0 1 1
use LUT4AB  Tile_X6Y5_LUT4AB
timestamp 0
transform 1 0 252576 0 1 448140
box 0 0 1 1
use LUT4AB  Tile_X6Y6_LUT4AB
timestamp 0
transform 1 0 252576 0 1 399756
box 0 0 1 1
use LUT4AB  Tile_X6Y7_LUT4AB
timestamp 0
transform 1 0 252576 0 1 351372
box 0 0 1 1
use LUT4AB  Tile_X6Y8_LUT4AB
timestamp 0
transform 1 0 252576 0 1 302988
box 0 0 1 1
use LUT4AB  Tile_X6Y9_LUT4AB
timestamp 0
transform 1 0 252576 0 1 254604
box 0 0 1 1
use LUT4AB  Tile_X6Y10_LUT4AB
timestamp 0
transform 1 0 252576 0 1 206220
box 0 0 1 1
use LUT4AB  Tile_X6Y11_LUT4AB
timestamp 0
transform 1 0 252576 0 1 157836
box 0 0 1 1
use LUT4AB  Tile_X6Y12_LUT4AB
timestamp 0
transform 1 0 252576 0 1 109452
box 0 0 1 1
use LUT4AB  Tile_X6Y13_LUT4AB
timestamp 0
transform 1 0 252576 0 1 61068
box 0 0 1 1
use LUT4AB  Tile_X6Y14_LUT4AB
timestamp 0
transform 1 0 252576 0 1 12684
box 0 0 1 1
use S_CPU_IF  Tile_X6Y15_S_CPU_IF
timestamp 0
transform 1 0 252576 0 1 840
box 0 0 1 1
use N_term_DSP  Tile_X7Y0_N_term_DSP
timestamp 0
transform 1 0 298944 0 1 690060
box 0 0 1 1
use DSP  Tile_X7Y1_DSP
timestamp 0
transform 1 0 298944 0 1 593292
box 0 0 1 1
use DSP  Tile_X7Y3_DSP
timestamp 0
transform 1 0 298944 0 1 496524
box 0 0 1 1
use DSP  Tile_X7Y5_DSP
timestamp 0
transform 1 0 298944 0 1 399756
box 0 0 1 1
use DSP  Tile_X7Y7_DSP
timestamp 0
transform 1 0 298944 0 1 302988
box 0 0 1 1
use DSP  Tile_X7Y9_DSP
timestamp 0
transform 1 0 298944 0 1 206220
box 0 0 1 1
use DSP  Tile_X7Y11_DSP
timestamp 0
transform 1 0 298944 0 1 109452
box 0 0 1 1
use DSP  Tile_X7Y13_DSP
timestamp 0
transform 1 0 298944 0 1 12684
box 0 0 1 1
use S_term_DSP  Tile_X7Y15_S_term_DSP
timestamp 0
transform 1 0 298944 0 1 840
box 0 0 1 1
use N_term_single  Tile_X8Y0_N_term_single
timestamp 0
transform 1 0 338208 0 1 690060
box 0 0 1 1
use LUT4AB  Tile_X8Y1_LUT4AB
timestamp 0
transform 1 0 338208 0 1 641676
box 0 0 1 1
use LUT4AB  Tile_X8Y2_LUT4AB
timestamp 0
transform 1 0 338208 0 1 593292
box 0 0 1 1
use LUT4AB  Tile_X8Y3_LUT4AB
timestamp 0
transform 1 0 338208 0 1 544908
box 0 0 1 1
use LUT4AB  Tile_X8Y4_LUT4AB
timestamp 0
transform 1 0 338208 0 1 496524
box 0 0 1 1
use LUT4AB  Tile_X8Y5_LUT4AB
timestamp 0
transform 1 0 338208 0 1 448140
box 0 0 1 1
use LUT4AB  Tile_X8Y6_LUT4AB
timestamp 0
transform 1 0 338208 0 1 399756
box 0 0 1 1
use LUT4AB  Tile_X8Y7_LUT4AB
timestamp 0
transform 1 0 338208 0 1 351372
box 0 0 1 1
use LUT4AB  Tile_X8Y8_LUT4AB
timestamp 0
transform 1 0 338208 0 1 302988
box 0 0 1 1
use LUT4AB  Tile_X8Y9_LUT4AB
timestamp 0
transform 1 0 338208 0 1 254604
box 0 0 1 1
use LUT4AB  Tile_X8Y10_LUT4AB
timestamp 0
transform 1 0 338208 0 1 206220
box 0 0 1 1
use LUT4AB  Tile_X8Y11_LUT4AB
timestamp 0
transform 1 0 338208 0 1 157836
box 0 0 1 1
use LUT4AB  Tile_X8Y12_LUT4AB
timestamp 0
transform 1 0 338208 0 1 109452
box 0 0 1 1
use LUT4AB  Tile_X8Y13_LUT4AB
timestamp 0
transform 1 0 338208 0 1 61068
box 0 0 1 1
use LUT4AB  Tile_X8Y14_LUT4AB
timestamp 0
transform 1 0 338208 0 1 12684
box 0 0 1 1
use S_CPU_IF  Tile_X8Y15_S_CPU_IF
timestamp 0
transform 1 0 338208 0 1 840
box 0 0 1 1
use N_term_single  Tile_X9Y0_N_term_single
timestamp 0
transform 1 0 384576 0 1 690060
box 0 0 1 1
use LUT4AB  Tile_X9Y1_LUT4AB
timestamp 0
transform 1 0 384576 0 1 641676
box 0 0 1 1
use LUT4AB  Tile_X9Y2_LUT4AB
timestamp 0
transform 1 0 384576 0 1 593292
box 0 0 1 1
use LUT4AB  Tile_X9Y3_LUT4AB
timestamp 0
transform 1 0 384576 0 1 544908
box 0 0 1 1
use LUT4AB  Tile_X9Y4_LUT4AB
timestamp 0
transform 1 0 384576 0 1 496524
box 0 0 1 1
use LUT4AB  Tile_X9Y5_LUT4AB
timestamp 0
transform 1 0 384576 0 1 448140
box 0 0 1 1
use LUT4AB  Tile_X9Y6_LUT4AB
timestamp 0
transform 1 0 384576 0 1 399756
box 0 0 1 1
use LUT4AB  Tile_X9Y7_LUT4AB
timestamp 0
transform 1 0 384576 0 1 351372
box 0 0 1 1
use LUT4AB  Tile_X9Y8_LUT4AB
timestamp 0
transform 1 0 384576 0 1 302988
box 0 0 1 1
use LUT4AB  Tile_X9Y9_LUT4AB
timestamp 0
transform 1 0 384576 0 1 254604
box 0 0 1 1
use LUT4AB  Tile_X9Y10_LUT4AB
timestamp 0
transform 1 0 384576 0 1 206220
box 0 0 1 1
use LUT4AB  Tile_X9Y11_LUT4AB
timestamp 0
transform 1 0 384576 0 1 157836
box 0 0 1 1
use LUT4AB  Tile_X9Y12_LUT4AB
timestamp 0
transform 1 0 384576 0 1 109452
box 0 0 1 1
use LUT4AB  Tile_X9Y13_LUT4AB
timestamp 0
transform 1 0 384576 0 1 61068
box 0 0 1 1
use LUT4AB  Tile_X9Y14_LUT4AB
timestamp 0
transform 1 0 384576 0 1 12684
box 0 0 1 1
use S_CPU_IF  Tile_X9Y15_S_CPU_IF
timestamp 0
transform 1 0 384576 0 1 840
box 0 0 1 1
use N_term_IHP_SRAM  Tile_X10Y0_N_term_IHP_SRAM
timestamp 0
transform 1 0 430944 0 1 690060
box 0 0 1 1
use IHP_SRAM  Tile_X10Y1_IHP_SRAM
timestamp 0
transform 1 0 430944 0 1 593292
box 0 0 1 1
use IHP_SRAM  Tile_X10Y3_IHP_SRAM
timestamp 0
transform 1 0 430944 0 1 496524
box 0 0 1 1
use IHP_SRAM  Tile_X10Y5_IHP_SRAM
timestamp 0
transform 1 0 430944 0 1 399756
box 0 0 1 1
use IHP_SRAM  Tile_X10Y7_IHP_SRAM
timestamp 0
transform 1 0 430944 0 1 302988
box 0 0 1 1
use IHP_SRAM  Tile_X10Y9_IHP_SRAM
timestamp 0
transform 1 0 430944 0 1 206220
box 0 0 1 1
use IHP_SRAM  Tile_X10Y11_IHP_SRAM
timestamp 0
transform 1 0 430944 0 1 109452
box 0 0 1 1
use IHP_SRAM  Tile_X10Y13_IHP_SRAM
timestamp 0
transform 1 0 430944 0 1 12684
box 0 0 1 1
use S_term_IHP_SRAM  Tile_X10Y15_S_term_IHP_SRAM
timestamp 0
transform 1 0 430944 0 1 840
box 0 0 1 1
<< labels >>
flabel metal2 s 0 690776 96 690856 0 FreeSans 320 0 0 0 FrameData[0]
port 0 nsew signal input
flabel metal2 s 0 564440 96 564520 0 FreeSans 320 0 0 0 FrameData[100]
port 1 nsew signal input
flabel metal2 s 0 565448 96 565528 0 FreeSans 320 0 0 0 FrameData[101]
port 2 nsew signal input
flabel metal2 s 0 566456 96 566536 0 FreeSans 320 0 0 0 FrameData[102]
port 3 nsew signal input
flabel metal2 s 0 567464 96 567544 0 FreeSans 320 0 0 0 FrameData[103]
port 4 nsew signal input
flabel metal2 s 0 568472 96 568552 0 FreeSans 320 0 0 0 FrameData[104]
port 5 nsew signal input
flabel metal2 s 0 569480 96 569560 0 FreeSans 320 0 0 0 FrameData[105]
port 6 nsew signal input
flabel metal2 s 0 570488 96 570568 0 FreeSans 320 0 0 0 FrameData[106]
port 7 nsew signal input
flabel metal2 s 0 571496 96 571576 0 FreeSans 320 0 0 0 FrameData[107]
port 8 nsew signal input
flabel metal2 s 0 572504 96 572584 0 FreeSans 320 0 0 0 FrameData[108]
port 9 nsew signal input
flabel metal2 s 0 573512 96 573592 0 FreeSans 320 0 0 0 FrameData[109]
port 10 nsew signal input
flabel metal2 s 0 694136 96 694216 0 FreeSans 320 0 0 0 FrameData[10]
port 11 nsew signal input
flabel metal2 s 0 574520 96 574600 0 FreeSans 320 0 0 0 FrameData[110]
port 12 nsew signal input
flabel metal2 s 0 575528 96 575608 0 FreeSans 320 0 0 0 FrameData[111]
port 13 nsew signal input
flabel metal2 s 0 576536 96 576616 0 FreeSans 320 0 0 0 FrameData[112]
port 14 nsew signal input
flabel metal2 s 0 577544 96 577624 0 FreeSans 320 0 0 0 FrameData[113]
port 15 nsew signal input
flabel metal2 s 0 578552 96 578632 0 FreeSans 320 0 0 0 FrameData[114]
port 16 nsew signal input
flabel metal2 s 0 579560 96 579640 0 FreeSans 320 0 0 0 FrameData[115]
port 17 nsew signal input
flabel metal2 s 0 580568 96 580648 0 FreeSans 320 0 0 0 FrameData[116]
port 18 nsew signal input
flabel metal2 s 0 581576 96 581656 0 FreeSans 320 0 0 0 FrameData[117]
port 19 nsew signal input
flabel metal2 s 0 582584 96 582664 0 FreeSans 320 0 0 0 FrameData[118]
port 20 nsew signal input
flabel metal2 s 0 583592 96 583672 0 FreeSans 320 0 0 0 FrameData[119]
port 21 nsew signal input
flabel metal2 s 0 694472 96 694552 0 FreeSans 320 0 0 0 FrameData[11]
port 22 nsew signal input
flabel metal2 s 0 584600 96 584680 0 FreeSans 320 0 0 0 FrameData[120]
port 23 nsew signal input
flabel metal2 s 0 585608 96 585688 0 FreeSans 320 0 0 0 FrameData[121]
port 24 nsew signal input
flabel metal2 s 0 586616 96 586696 0 FreeSans 320 0 0 0 FrameData[122]
port 25 nsew signal input
flabel metal2 s 0 587624 96 587704 0 FreeSans 320 0 0 0 FrameData[123]
port 26 nsew signal input
flabel metal2 s 0 588632 96 588712 0 FreeSans 320 0 0 0 FrameData[124]
port 27 nsew signal input
flabel metal2 s 0 589640 96 589720 0 FreeSans 320 0 0 0 FrameData[125]
port 28 nsew signal input
flabel metal2 s 0 590648 96 590728 0 FreeSans 320 0 0 0 FrameData[126]
port 29 nsew signal input
flabel metal2 s 0 591656 96 591736 0 FreeSans 320 0 0 0 FrameData[127]
port 30 nsew signal input
flabel metal2 s 0 512024 96 512104 0 FreeSans 320 0 0 0 FrameData[128]
port 31 nsew signal input
flabel metal2 s 0 513032 96 513112 0 FreeSans 320 0 0 0 FrameData[129]
port 32 nsew signal input
flabel metal2 s 0 694808 96 694888 0 FreeSans 320 0 0 0 FrameData[12]
port 33 nsew signal input
flabel metal2 s 0 514040 96 514120 0 FreeSans 320 0 0 0 FrameData[130]
port 34 nsew signal input
flabel metal2 s 0 515048 96 515128 0 FreeSans 320 0 0 0 FrameData[131]
port 35 nsew signal input
flabel metal2 s 0 516056 96 516136 0 FreeSans 320 0 0 0 FrameData[132]
port 36 nsew signal input
flabel metal2 s 0 517064 96 517144 0 FreeSans 320 0 0 0 FrameData[133]
port 37 nsew signal input
flabel metal2 s 0 518072 96 518152 0 FreeSans 320 0 0 0 FrameData[134]
port 38 nsew signal input
flabel metal2 s 0 519080 96 519160 0 FreeSans 320 0 0 0 FrameData[135]
port 39 nsew signal input
flabel metal2 s 0 520088 96 520168 0 FreeSans 320 0 0 0 FrameData[136]
port 40 nsew signal input
flabel metal2 s 0 521096 96 521176 0 FreeSans 320 0 0 0 FrameData[137]
port 41 nsew signal input
flabel metal2 s 0 522104 96 522184 0 FreeSans 320 0 0 0 FrameData[138]
port 42 nsew signal input
flabel metal2 s 0 523112 96 523192 0 FreeSans 320 0 0 0 FrameData[139]
port 43 nsew signal input
flabel metal2 s 0 695144 96 695224 0 FreeSans 320 0 0 0 FrameData[13]
port 44 nsew signal input
flabel metal2 s 0 524120 96 524200 0 FreeSans 320 0 0 0 FrameData[140]
port 45 nsew signal input
flabel metal2 s 0 525128 96 525208 0 FreeSans 320 0 0 0 FrameData[141]
port 46 nsew signal input
flabel metal2 s 0 526136 96 526216 0 FreeSans 320 0 0 0 FrameData[142]
port 47 nsew signal input
flabel metal2 s 0 527144 96 527224 0 FreeSans 320 0 0 0 FrameData[143]
port 48 nsew signal input
flabel metal2 s 0 528152 96 528232 0 FreeSans 320 0 0 0 FrameData[144]
port 49 nsew signal input
flabel metal2 s 0 529160 96 529240 0 FreeSans 320 0 0 0 FrameData[145]
port 50 nsew signal input
flabel metal2 s 0 530168 96 530248 0 FreeSans 320 0 0 0 FrameData[146]
port 51 nsew signal input
flabel metal2 s 0 531176 96 531256 0 FreeSans 320 0 0 0 FrameData[147]
port 52 nsew signal input
flabel metal2 s 0 532184 96 532264 0 FreeSans 320 0 0 0 FrameData[148]
port 53 nsew signal input
flabel metal2 s 0 533192 96 533272 0 FreeSans 320 0 0 0 FrameData[149]
port 54 nsew signal input
flabel metal2 s 0 695480 96 695560 0 FreeSans 320 0 0 0 FrameData[14]
port 55 nsew signal input
flabel metal2 s 0 534200 96 534280 0 FreeSans 320 0 0 0 FrameData[150]
port 56 nsew signal input
flabel metal2 s 0 535208 96 535288 0 FreeSans 320 0 0 0 FrameData[151]
port 57 nsew signal input
flabel metal2 s 0 536216 96 536296 0 FreeSans 320 0 0 0 FrameData[152]
port 58 nsew signal input
flabel metal2 s 0 537224 96 537304 0 FreeSans 320 0 0 0 FrameData[153]
port 59 nsew signal input
flabel metal2 s 0 538232 96 538312 0 FreeSans 320 0 0 0 FrameData[154]
port 60 nsew signal input
flabel metal2 s 0 539240 96 539320 0 FreeSans 320 0 0 0 FrameData[155]
port 61 nsew signal input
flabel metal2 s 0 540248 96 540328 0 FreeSans 320 0 0 0 FrameData[156]
port 62 nsew signal input
flabel metal2 s 0 541256 96 541336 0 FreeSans 320 0 0 0 FrameData[157]
port 63 nsew signal input
flabel metal2 s 0 542264 96 542344 0 FreeSans 320 0 0 0 FrameData[158]
port 64 nsew signal input
flabel metal2 s 0 543272 96 543352 0 FreeSans 320 0 0 0 FrameData[159]
port 65 nsew signal input
flabel metal2 s 0 695816 96 695896 0 FreeSans 320 0 0 0 FrameData[15]
port 66 nsew signal input
flabel metal2 s 0 463640 96 463720 0 FreeSans 320 0 0 0 FrameData[160]
port 67 nsew signal input
flabel metal2 s 0 464648 96 464728 0 FreeSans 320 0 0 0 FrameData[161]
port 68 nsew signal input
flabel metal2 s 0 465656 96 465736 0 FreeSans 320 0 0 0 FrameData[162]
port 69 nsew signal input
flabel metal2 s 0 466664 96 466744 0 FreeSans 320 0 0 0 FrameData[163]
port 70 nsew signal input
flabel metal2 s 0 467672 96 467752 0 FreeSans 320 0 0 0 FrameData[164]
port 71 nsew signal input
flabel metal2 s 0 468680 96 468760 0 FreeSans 320 0 0 0 FrameData[165]
port 72 nsew signal input
flabel metal2 s 0 469688 96 469768 0 FreeSans 320 0 0 0 FrameData[166]
port 73 nsew signal input
flabel metal2 s 0 470696 96 470776 0 FreeSans 320 0 0 0 FrameData[167]
port 74 nsew signal input
flabel metal2 s 0 471704 96 471784 0 FreeSans 320 0 0 0 FrameData[168]
port 75 nsew signal input
flabel metal2 s 0 472712 96 472792 0 FreeSans 320 0 0 0 FrameData[169]
port 76 nsew signal input
flabel metal2 s 0 696152 96 696232 0 FreeSans 320 0 0 0 FrameData[16]
port 77 nsew signal input
flabel metal2 s 0 473720 96 473800 0 FreeSans 320 0 0 0 FrameData[170]
port 78 nsew signal input
flabel metal2 s 0 474728 96 474808 0 FreeSans 320 0 0 0 FrameData[171]
port 79 nsew signal input
flabel metal2 s 0 475736 96 475816 0 FreeSans 320 0 0 0 FrameData[172]
port 80 nsew signal input
flabel metal2 s 0 476744 96 476824 0 FreeSans 320 0 0 0 FrameData[173]
port 81 nsew signal input
flabel metal2 s 0 477752 96 477832 0 FreeSans 320 0 0 0 FrameData[174]
port 82 nsew signal input
flabel metal2 s 0 478760 96 478840 0 FreeSans 320 0 0 0 FrameData[175]
port 83 nsew signal input
flabel metal2 s 0 479768 96 479848 0 FreeSans 320 0 0 0 FrameData[176]
port 84 nsew signal input
flabel metal2 s 0 480776 96 480856 0 FreeSans 320 0 0 0 FrameData[177]
port 85 nsew signal input
flabel metal2 s 0 481784 96 481864 0 FreeSans 320 0 0 0 FrameData[178]
port 86 nsew signal input
flabel metal2 s 0 482792 96 482872 0 FreeSans 320 0 0 0 FrameData[179]
port 87 nsew signal input
flabel metal2 s 0 696488 96 696568 0 FreeSans 320 0 0 0 FrameData[17]
port 88 nsew signal input
flabel metal2 s 0 483800 96 483880 0 FreeSans 320 0 0 0 FrameData[180]
port 89 nsew signal input
flabel metal2 s 0 484808 96 484888 0 FreeSans 320 0 0 0 FrameData[181]
port 90 nsew signal input
flabel metal2 s 0 485816 96 485896 0 FreeSans 320 0 0 0 FrameData[182]
port 91 nsew signal input
flabel metal2 s 0 486824 96 486904 0 FreeSans 320 0 0 0 FrameData[183]
port 92 nsew signal input
flabel metal2 s 0 487832 96 487912 0 FreeSans 320 0 0 0 FrameData[184]
port 93 nsew signal input
flabel metal2 s 0 488840 96 488920 0 FreeSans 320 0 0 0 FrameData[185]
port 94 nsew signal input
flabel metal2 s 0 489848 96 489928 0 FreeSans 320 0 0 0 FrameData[186]
port 95 nsew signal input
flabel metal2 s 0 490856 96 490936 0 FreeSans 320 0 0 0 FrameData[187]
port 96 nsew signal input
flabel metal2 s 0 491864 96 491944 0 FreeSans 320 0 0 0 FrameData[188]
port 97 nsew signal input
flabel metal2 s 0 492872 96 492952 0 FreeSans 320 0 0 0 FrameData[189]
port 98 nsew signal input
flabel metal2 s 0 696824 96 696904 0 FreeSans 320 0 0 0 FrameData[18]
port 99 nsew signal input
flabel metal2 s 0 493880 96 493960 0 FreeSans 320 0 0 0 FrameData[190]
port 100 nsew signal input
flabel metal2 s 0 494888 96 494968 0 FreeSans 320 0 0 0 FrameData[191]
port 101 nsew signal input
flabel metal2 s 0 415256 96 415336 0 FreeSans 320 0 0 0 FrameData[192]
port 102 nsew signal input
flabel metal2 s 0 416264 96 416344 0 FreeSans 320 0 0 0 FrameData[193]
port 103 nsew signal input
flabel metal2 s 0 417272 96 417352 0 FreeSans 320 0 0 0 FrameData[194]
port 104 nsew signal input
flabel metal2 s 0 418280 96 418360 0 FreeSans 320 0 0 0 FrameData[195]
port 105 nsew signal input
flabel metal2 s 0 419288 96 419368 0 FreeSans 320 0 0 0 FrameData[196]
port 106 nsew signal input
flabel metal2 s 0 420296 96 420376 0 FreeSans 320 0 0 0 FrameData[197]
port 107 nsew signal input
flabel metal2 s 0 421304 96 421384 0 FreeSans 320 0 0 0 FrameData[198]
port 108 nsew signal input
flabel metal2 s 0 422312 96 422392 0 FreeSans 320 0 0 0 FrameData[199]
port 109 nsew signal input
flabel metal2 s 0 697160 96 697240 0 FreeSans 320 0 0 0 FrameData[19]
port 110 nsew signal input
flabel metal2 s 0 691112 96 691192 0 FreeSans 320 0 0 0 FrameData[1]
port 111 nsew signal input
flabel metal2 s 0 423320 96 423400 0 FreeSans 320 0 0 0 FrameData[200]
port 112 nsew signal input
flabel metal2 s 0 424328 96 424408 0 FreeSans 320 0 0 0 FrameData[201]
port 113 nsew signal input
flabel metal2 s 0 425336 96 425416 0 FreeSans 320 0 0 0 FrameData[202]
port 114 nsew signal input
flabel metal2 s 0 426344 96 426424 0 FreeSans 320 0 0 0 FrameData[203]
port 115 nsew signal input
flabel metal2 s 0 427352 96 427432 0 FreeSans 320 0 0 0 FrameData[204]
port 116 nsew signal input
flabel metal2 s 0 428360 96 428440 0 FreeSans 320 0 0 0 FrameData[205]
port 117 nsew signal input
flabel metal2 s 0 429368 96 429448 0 FreeSans 320 0 0 0 FrameData[206]
port 118 nsew signal input
flabel metal2 s 0 430376 96 430456 0 FreeSans 320 0 0 0 FrameData[207]
port 119 nsew signal input
flabel metal2 s 0 431384 96 431464 0 FreeSans 320 0 0 0 FrameData[208]
port 120 nsew signal input
flabel metal2 s 0 432392 96 432472 0 FreeSans 320 0 0 0 FrameData[209]
port 121 nsew signal input
flabel metal2 s 0 697496 96 697576 0 FreeSans 320 0 0 0 FrameData[20]
port 122 nsew signal input
flabel metal2 s 0 433400 96 433480 0 FreeSans 320 0 0 0 FrameData[210]
port 123 nsew signal input
flabel metal2 s 0 434408 96 434488 0 FreeSans 320 0 0 0 FrameData[211]
port 124 nsew signal input
flabel metal2 s 0 435416 96 435496 0 FreeSans 320 0 0 0 FrameData[212]
port 125 nsew signal input
flabel metal2 s 0 436424 96 436504 0 FreeSans 320 0 0 0 FrameData[213]
port 126 nsew signal input
flabel metal2 s 0 437432 96 437512 0 FreeSans 320 0 0 0 FrameData[214]
port 127 nsew signal input
flabel metal2 s 0 438440 96 438520 0 FreeSans 320 0 0 0 FrameData[215]
port 128 nsew signal input
flabel metal2 s 0 439448 96 439528 0 FreeSans 320 0 0 0 FrameData[216]
port 129 nsew signal input
flabel metal2 s 0 440456 96 440536 0 FreeSans 320 0 0 0 FrameData[217]
port 130 nsew signal input
flabel metal2 s 0 441464 96 441544 0 FreeSans 320 0 0 0 FrameData[218]
port 131 nsew signal input
flabel metal2 s 0 442472 96 442552 0 FreeSans 320 0 0 0 FrameData[219]
port 132 nsew signal input
flabel metal2 s 0 697832 96 697912 0 FreeSans 320 0 0 0 FrameData[21]
port 133 nsew signal input
flabel metal2 s 0 443480 96 443560 0 FreeSans 320 0 0 0 FrameData[220]
port 134 nsew signal input
flabel metal2 s 0 444488 96 444568 0 FreeSans 320 0 0 0 FrameData[221]
port 135 nsew signal input
flabel metal2 s 0 445496 96 445576 0 FreeSans 320 0 0 0 FrameData[222]
port 136 nsew signal input
flabel metal2 s 0 446504 96 446584 0 FreeSans 320 0 0 0 FrameData[223]
port 137 nsew signal input
flabel metal2 s 0 366872 96 366952 0 FreeSans 320 0 0 0 FrameData[224]
port 138 nsew signal input
flabel metal2 s 0 367880 96 367960 0 FreeSans 320 0 0 0 FrameData[225]
port 139 nsew signal input
flabel metal2 s 0 368888 96 368968 0 FreeSans 320 0 0 0 FrameData[226]
port 140 nsew signal input
flabel metal2 s 0 369896 96 369976 0 FreeSans 320 0 0 0 FrameData[227]
port 141 nsew signal input
flabel metal2 s 0 370904 96 370984 0 FreeSans 320 0 0 0 FrameData[228]
port 142 nsew signal input
flabel metal2 s 0 371912 96 371992 0 FreeSans 320 0 0 0 FrameData[229]
port 143 nsew signal input
flabel metal2 s 0 698168 96 698248 0 FreeSans 320 0 0 0 FrameData[22]
port 144 nsew signal input
flabel metal2 s 0 372920 96 373000 0 FreeSans 320 0 0 0 FrameData[230]
port 145 nsew signal input
flabel metal2 s 0 373928 96 374008 0 FreeSans 320 0 0 0 FrameData[231]
port 146 nsew signal input
flabel metal2 s 0 374936 96 375016 0 FreeSans 320 0 0 0 FrameData[232]
port 147 nsew signal input
flabel metal2 s 0 375944 96 376024 0 FreeSans 320 0 0 0 FrameData[233]
port 148 nsew signal input
flabel metal2 s 0 376952 96 377032 0 FreeSans 320 0 0 0 FrameData[234]
port 149 nsew signal input
flabel metal2 s 0 377960 96 378040 0 FreeSans 320 0 0 0 FrameData[235]
port 150 nsew signal input
flabel metal2 s 0 378968 96 379048 0 FreeSans 320 0 0 0 FrameData[236]
port 151 nsew signal input
flabel metal2 s 0 379976 96 380056 0 FreeSans 320 0 0 0 FrameData[237]
port 152 nsew signal input
flabel metal2 s 0 380984 96 381064 0 FreeSans 320 0 0 0 FrameData[238]
port 153 nsew signal input
flabel metal2 s 0 381992 96 382072 0 FreeSans 320 0 0 0 FrameData[239]
port 154 nsew signal input
flabel metal2 s 0 698504 96 698584 0 FreeSans 320 0 0 0 FrameData[23]
port 155 nsew signal input
flabel metal2 s 0 383000 96 383080 0 FreeSans 320 0 0 0 FrameData[240]
port 156 nsew signal input
flabel metal2 s 0 384008 96 384088 0 FreeSans 320 0 0 0 FrameData[241]
port 157 nsew signal input
flabel metal2 s 0 385016 96 385096 0 FreeSans 320 0 0 0 FrameData[242]
port 158 nsew signal input
flabel metal2 s 0 386024 96 386104 0 FreeSans 320 0 0 0 FrameData[243]
port 159 nsew signal input
flabel metal2 s 0 387032 96 387112 0 FreeSans 320 0 0 0 FrameData[244]
port 160 nsew signal input
flabel metal2 s 0 388040 96 388120 0 FreeSans 320 0 0 0 FrameData[245]
port 161 nsew signal input
flabel metal2 s 0 389048 96 389128 0 FreeSans 320 0 0 0 FrameData[246]
port 162 nsew signal input
flabel metal2 s 0 390056 96 390136 0 FreeSans 320 0 0 0 FrameData[247]
port 163 nsew signal input
flabel metal2 s 0 391064 96 391144 0 FreeSans 320 0 0 0 FrameData[248]
port 164 nsew signal input
flabel metal2 s 0 392072 96 392152 0 FreeSans 320 0 0 0 FrameData[249]
port 165 nsew signal input
flabel metal2 s 0 698840 96 698920 0 FreeSans 320 0 0 0 FrameData[24]
port 166 nsew signal input
flabel metal2 s 0 393080 96 393160 0 FreeSans 320 0 0 0 FrameData[250]
port 167 nsew signal input
flabel metal2 s 0 394088 96 394168 0 FreeSans 320 0 0 0 FrameData[251]
port 168 nsew signal input
flabel metal2 s 0 395096 96 395176 0 FreeSans 320 0 0 0 FrameData[252]
port 169 nsew signal input
flabel metal2 s 0 396104 96 396184 0 FreeSans 320 0 0 0 FrameData[253]
port 170 nsew signal input
flabel metal2 s 0 397112 96 397192 0 FreeSans 320 0 0 0 FrameData[254]
port 171 nsew signal input
flabel metal2 s 0 398120 96 398200 0 FreeSans 320 0 0 0 FrameData[255]
port 172 nsew signal input
flabel metal2 s 0 318488 96 318568 0 FreeSans 320 0 0 0 FrameData[256]
port 173 nsew signal input
flabel metal2 s 0 319496 96 319576 0 FreeSans 320 0 0 0 FrameData[257]
port 174 nsew signal input
flabel metal2 s 0 320504 96 320584 0 FreeSans 320 0 0 0 FrameData[258]
port 175 nsew signal input
flabel metal2 s 0 321512 96 321592 0 FreeSans 320 0 0 0 FrameData[259]
port 176 nsew signal input
flabel metal2 s 0 699176 96 699256 0 FreeSans 320 0 0 0 FrameData[25]
port 177 nsew signal input
flabel metal2 s 0 322520 96 322600 0 FreeSans 320 0 0 0 FrameData[260]
port 178 nsew signal input
flabel metal2 s 0 323528 96 323608 0 FreeSans 320 0 0 0 FrameData[261]
port 179 nsew signal input
flabel metal2 s 0 324536 96 324616 0 FreeSans 320 0 0 0 FrameData[262]
port 180 nsew signal input
flabel metal2 s 0 325544 96 325624 0 FreeSans 320 0 0 0 FrameData[263]
port 181 nsew signal input
flabel metal2 s 0 326552 96 326632 0 FreeSans 320 0 0 0 FrameData[264]
port 182 nsew signal input
flabel metal2 s 0 327560 96 327640 0 FreeSans 320 0 0 0 FrameData[265]
port 183 nsew signal input
flabel metal2 s 0 328568 96 328648 0 FreeSans 320 0 0 0 FrameData[266]
port 184 nsew signal input
flabel metal2 s 0 329576 96 329656 0 FreeSans 320 0 0 0 FrameData[267]
port 185 nsew signal input
flabel metal2 s 0 330584 96 330664 0 FreeSans 320 0 0 0 FrameData[268]
port 186 nsew signal input
flabel metal2 s 0 331592 96 331672 0 FreeSans 320 0 0 0 FrameData[269]
port 187 nsew signal input
flabel metal2 s 0 699512 96 699592 0 FreeSans 320 0 0 0 FrameData[26]
port 188 nsew signal input
flabel metal2 s 0 332600 96 332680 0 FreeSans 320 0 0 0 FrameData[270]
port 189 nsew signal input
flabel metal2 s 0 333608 96 333688 0 FreeSans 320 0 0 0 FrameData[271]
port 190 nsew signal input
flabel metal2 s 0 334616 96 334696 0 FreeSans 320 0 0 0 FrameData[272]
port 191 nsew signal input
flabel metal2 s 0 335624 96 335704 0 FreeSans 320 0 0 0 FrameData[273]
port 192 nsew signal input
flabel metal2 s 0 336632 96 336712 0 FreeSans 320 0 0 0 FrameData[274]
port 193 nsew signal input
flabel metal2 s 0 337640 96 337720 0 FreeSans 320 0 0 0 FrameData[275]
port 194 nsew signal input
flabel metal2 s 0 338648 96 338728 0 FreeSans 320 0 0 0 FrameData[276]
port 195 nsew signal input
flabel metal2 s 0 339656 96 339736 0 FreeSans 320 0 0 0 FrameData[277]
port 196 nsew signal input
flabel metal2 s 0 340664 96 340744 0 FreeSans 320 0 0 0 FrameData[278]
port 197 nsew signal input
flabel metal2 s 0 341672 96 341752 0 FreeSans 320 0 0 0 FrameData[279]
port 198 nsew signal input
flabel metal2 s 0 699848 96 699928 0 FreeSans 320 0 0 0 FrameData[27]
port 199 nsew signal input
flabel metal2 s 0 342680 96 342760 0 FreeSans 320 0 0 0 FrameData[280]
port 200 nsew signal input
flabel metal2 s 0 343688 96 343768 0 FreeSans 320 0 0 0 FrameData[281]
port 201 nsew signal input
flabel metal2 s 0 344696 96 344776 0 FreeSans 320 0 0 0 FrameData[282]
port 202 nsew signal input
flabel metal2 s 0 345704 96 345784 0 FreeSans 320 0 0 0 FrameData[283]
port 203 nsew signal input
flabel metal2 s 0 346712 96 346792 0 FreeSans 320 0 0 0 FrameData[284]
port 204 nsew signal input
flabel metal2 s 0 347720 96 347800 0 FreeSans 320 0 0 0 FrameData[285]
port 205 nsew signal input
flabel metal2 s 0 348728 96 348808 0 FreeSans 320 0 0 0 FrameData[286]
port 206 nsew signal input
flabel metal2 s 0 349736 96 349816 0 FreeSans 320 0 0 0 FrameData[287]
port 207 nsew signal input
flabel metal2 s 0 270104 96 270184 0 FreeSans 320 0 0 0 FrameData[288]
port 208 nsew signal input
flabel metal2 s 0 271112 96 271192 0 FreeSans 320 0 0 0 FrameData[289]
port 209 nsew signal input
flabel metal2 s 0 700184 96 700264 0 FreeSans 320 0 0 0 FrameData[28]
port 210 nsew signal input
flabel metal2 s 0 272120 96 272200 0 FreeSans 320 0 0 0 FrameData[290]
port 211 nsew signal input
flabel metal2 s 0 273128 96 273208 0 FreeSans 320 0 0 0 FrameData[291]
port 212 nsew signal input
flabel metal2 s 0 274136 96 274216 0 FreeSans 320 0 0 0 FrameData[292]
port 213 nsew signal input
flabel metal2 s 0 275144 96 275224 0 FreeSans 320 0 0 0 FrameData[293]
port 214 nsew signal input
flabel metal2 s 0 276152 96 276232 0 FreeSans 320 0 0 0 FrameData[294]
port 215 nsew signal input
flabel metal2 s 0 277160 96 277240 0 FreeSans 320 0 0 0 FrameData[295]
port 216 nsew signal input
flabel metal2 s 0 278168 96 278248 0 FreeSans 320 0 0 0 FrameData[296]
port 217 nsew signal input
flabel metal2 s 0 279176 96 279256 0 FreeSans 320 0 0 0 FrameData[297]
port 218 nsew signal input
flabel metal2 s 0 280184 96 280264 0 FreeSans 320 0 0 0 FrameData[298]
port 219 nsew signal input
flabel metal2 s 0 281192 96 281272 0 FreeSans 320 0 0 0 FrameData[299]
port 220 nsew signal input
flabel metal2 s 0 700520 96 700600 0 FreeSans 320 0 0 0 FrameData[29]
port 221 nsew signal input
flabel metal2 s 0 691448 96 691528 0 FreeSans 320 0 0 0 FrameData[2]
port 222 nsew signal input
flabel metal2 s 0 282200 96 282280 0 FreeSans 320 0 0 0 FrameData[300]
port 223 nsew signal input
flabel metal2 s 0 283208 96 283288 0 FreeSans 320 0 0 0 FrameData[301]
port 224 nsew signal input
flabel metal2 s 0 284216 96 284296 0 FreeSans 320 0 0 0 FrameData[302]
port 225 nsew signal input
flabel metal2 s 0 285224 96 285304 0 FreeSans 320 0 0 0 FrameData[303]
port 226 nsew signal input
flabel metal2 s 0 286232 96 286312 0 FreeSans 320 0 0 0 FrameData[304]
port 227 nsew signal input
flabel metal2 s 0 287240 96 287320 0 FreeSans 320 0 0 0 FrameData[305]
port 228 nsew signal input
flabel metal2 s 0 288248 96 288328 0 FreeSans 320 0 0 0 FrameData[306]
port 229 nsew signal input
flabel metal2 s 0 289256 96 289336 0 FreeSans 320 0 0 0 FrameData[307]
port 230 nsew signal input
flabel metal2 s 0 290264 96 290344 0 FreeSans 320 0 0 0 FrameData[308]
port 231 nsew signal input
flabel metal2 s 0 291272 96 291352 0 FreeSans 320 0 0 0 FrameData[309]
port 232 nsew signal input
flabel metal2 s 0 700856 96 700936 0 FreeSans 320 0 0 0 FrameData[30]
port 233 nsew signal input
flabel metal2 s 0 292280 96 292360 0 FreeSans 320 0 0 0 FrameData[310]
port 234 nsew signal input
flabel metal2 s 0 293288 96 293368 0 FreeSans 320 0 0 0 FrameData[311]
port 235 nsew signal input
flabel metal2 s 0 294296 96 294376 0 FreeSans 320 0 0 0 FrameData[312]
port 236 nsew signal input
flabel metal2 s 0 295304 96 295384 0 FreeSans 320 0 0 0 FrameData[313]
port 237 nsew signal input
flabel metal2 s 0 296312 96 296392 0 FreeSans 320 0 0 0 FrameData[314]
port 238 nsew signal input
flabel metal2 s 0 297320 96 297400 0 FreeSans 320 0 0 0 FrameData[315]
port 239 nsew signal input
flabel metal2 s 0 298328 96 298408 0 FreeSans 320 0 0 0 FrameData[316]
port 240 nsew signal input
flabel metal2 s 0 299336 96 299416 0 FreeSans 320 0 0 0 FrameData[317]
port 241 nsew signal input
flabel metal2 s 0 300344 96 300424 0 FreeSans 320 0 0 0 FrameData[318]
port 242 nsew signal input
flabel metal2 s 0 301352 96 301432 0 FreeSans 320 0 0 0 FrameData[319]
port 243 nsew signal input
flabel metal2 s 0 701192 96 701272 0 FreeSans 320 0 0 0 FrameData[31]
port 244 nsew signal input
flabel metal2 s 0 221720 96 221800 0 FreeSans 320 0 0 0 FrameData[320]
port 245 nsew signal input
flabel metal2 s 0 222728 96 222808 0 FreeSans 320 0 0 0 FrameData[321]
port 246 nsew signal input
flabel metal2 s 0 223736 96 223816 0 FreeSans 320 0 0 0 FrameData[322]
port 247 nsew signal input
flabel metal2 s 0 224744 96 224824 0 FreeSans 320 0 0 0 FrameData[323]
port 248 nsew signal input
flabel metal2 s 0 225752 96 225832 0 FreeSans 320 0 0 0 FrameData[324]
port 249 nsew signal input
flabel metal2 s 0 226760 96 226840 0 FreeSans 320 0 0 0 FrameData[325]
port 250 nsew signal input
flabel metal2 s 0 227768 96 227848 0 FreeSans 320 0 0 0 FrameData[326]
port 251 nsew signal input
flabel metal2 s 0 228776 96 228856 0 FreeSans 320 0 0 0 FrameData[327]
port 252 nsew signal input
flabel metal2 s 0 229784 96 229864 0 FreeSans 320 0 0 0 FrameData[328]
port 253 nsew signal input
flabel metal2 s 0 230792 96 230872 0 FreeSans 320 0 0 0 FrameData[329]
port 254 nsew signal input
flabel metal2 s 0 657176 96 657256 0 FreeSans 320 0 0 0 FrameData[32]
port 255 nsew signal input
flabel metal2 s 0 231800 96 231880 0 FreeSans 320 0 0 0 FrameData[330]
port 256 nsew signal input
flabel metal2 s 0 232808 96 232888 0 FreeSans 320 0 0 0 FrameData[331]
port 257 nsew signal input
flabel metal2 s 0 233816 96 233896 0 FreeSans 320 0 0 0 FrameData[332]
port 258 nsew signal input
flabel metal2 s 0 234824 96 234904 0 FreeSans 320 0 0 0 FrameData[333]
port 259 nsew signal input
flabel metal2 s 0 235832 96 235912 0 FreeSans 320 0 0 0 FrameData[334]
port 260 nsew signal input
flabel metal2 s 0 236840 96 236920 0 FreeSans 320 0 0 0 FrameData[335]
port 261 nsew signal input
flabel metal2 s 0 237848 96 237928 0 FreeSans 320 0 0 0 FrameData[336]
port 262 nsew signal input
flabel metal2 s 0 238856 96 238936 0 FreeSans 320 0 0 0 FrameData[337]
port 263 nsew signal input
flabel metal2 s 0 239864 96 239944 0 FreeSans 320 0 0 0 FrameData[338]
port 264 nsew signal input
flabel metal2 s 0 240872 96 240952 0 FreeSans 320 0 0 0 FrameData[339]
port 265 nsew signal input
flabel metal2 s 0 658184 96 658264 0 FreeSans 320 0 0 0 FrameData[33]
port 266 nsew signal input
flabel metal2 s 0 241880 96 241960 0 FreeSans 320 0 0 0 FrameData[340]
port 267 nsew signal input
flabel metal2 s 0 242888 96 242968 0 FreeSans 320 0 0 0 FrameData[341]
port 268 nsew signal input
flabel metal2 s 0 243896 96 243976 0 FreeSans 320 0 0 0 FrameData[342]
port 269 nsew signal input
flabel metal2 s 0 244904 96 244984 0 FreeSans 320 0 0 0 FrameData[343]
port 270 nsew signal input
flabel metal2 s 0 245912 96 245992 0 FreeSans 320 0 0 0 FrameData[344]
port 271 nsew signal input
flabel metal2 s 0 246920 96 247000 0 FreeSans 320 0 0 0 FrameData[345]
port 272 nsew signal input
flabel metal2 s 0 247928 96 248008 0 FreeSans 320 0 0 0 FrameData[346]
port 273 nsew signal input
flabel metal2 s 0 248936 96 249016 0 FreeSans 320 0 0 0 FrameData[347]
port 274 nsew signal input
flabel metal2 s 0 249944 96 250024 0 FreeSans 320 0 0 0 FrameData[348]
port 275 nsew signal input
flabel metal2 s 0 250952 96 251032 0 FreeSans 320 0 0 0 FrameData[349]
port 276 nsew signal input
flabel metal2 s 0 659192 96 659272 0 FreeSans 320 0 0 0 FrameData[34]
port 277 nsew signal input
flabel metal2 s 0 251960 96 252040 0 FreeSans 320 0 0 0 FrameData[350]
port 278 nsew signal input
flabel metal2 s 0 252968 96 253048 0 FreeSans 320 0 0 0 FrameData[351]
port 279 nsew signal input
flabel metal2 s 0 173336 96 173416 0 FreeSans 320 0 0 0 FrameData[352]
port 280 nsew signal input
flabel metal2 s 0 174344 96 174424 0 FreeSans 320 0 0 0 FrameData[353]
port 281 nsew signal input
flabel metal2 s 0 175352 96 175432 0 FreeSans 320 0 0 0 FrameData[354]
port 282 nsew signal input
flabel metal2 s 0 176360 96 176440 0 FreeSans 320 0 0 0 FrameData[355]
port 283 nsew signal input
flabel metal2 s 0 177368 96 177448 0 FreeSans 320 0 0 0 FrameData[356]
port 284 nsew signal input
flabel metal2 s 0 178376 96 178456 0 FreeSans 320 0 0 0 FrameData[357]
port 285 nsew signal input
flabel metal2 s 0 179384 96 179464 0 FreeSans 320 0 0 0 FrameData[358]
port 286 nsew signal input
flabel metal2 s 0 180392 96 180472 0 FreeSans 320 0 0 0 FrameData[359]
port 287 nsew signal input
flabel metal2 s 0 660200 96 660280 0 FreeSans 320 0 0 0 FrameData[35]
port 288 nsew signal input
flabel metal2 s 0 181400 96 181480 0 FreeSans 320 0 0 0 FrameData[360]
port 289 nsew signal input
flabel metal2 s 0 182408 96 182488 0 FreeSans 320 0 0 0 FrameData[361]
port 290 nsew signal input
flabel metal2 s 0 183416 96 183496 0 FreeSans 320 0 0 0 FrameData[362]
port 291 nsew signal input
flabel metal2 s 0 184424 96 184504 0 FreeSans 320 0 0 0 FrameData[363]
port 292 nsew signal input
flabel metal2 s 0 185432 96 185512 0 FreeSans 320 0 0 0 FrameData[364]
port 293 nsew signal input
flabel metal2 s 0 186440 96 186520 0 FreeSans 320 0 0 0 FrameData[365]
port 294 nsew signal input
flabel metal2 s 0 187448 96 187528 0 FreeSans 320 0 0 0 FrameData[366]
port 295 nsew signal input
flabel metal2 s 0 188456 96 188536 0 FreeSans 320 0 0 0 FrameData[367]
port 296 nsew signal input
flabel metal2 s 0 189464 96 189544 0 FreeSans 320 0 0 0 FrameData[368]
port 297 nsew signal input
flabel metal2 s 0 190472 96 190552 0 FreeSans 320 0 0 0 FrameData[369]
port 298 nsew signal input
flabel metal2 s 0 661208 96 661288 0 FreeSans 320 0 0 0 FrameData[36]
port 299 nsew signal input
flabel metal2 s 0 191480 96 191560 0 FreeSans 320 0 0 0 FrameData[370]
port 300 nsew signal input
flabel metal2 s 0 192488 96 192568 0 FreeSans 320 0 0 0 FrameData[371]
port 301 nsew signal input
flabel metal2 s 0 193496 96 193576 0 FreeSans 320 0 0 0 FrameData[372]
port 302 nsew signal input
flabel metal2 s 0 194504 96 194584 0 FreeSans 320 0 0 0 FrameData[373]
port 303 nsew signal input
flabel metal2 s 0 195512 96 195592 0 FreeSans 320 0 0 0 FrameData[374]
port 304 nsew signal input
flabel metal2 s 0 196520 96 196600 0 FreeSans 320 0 0 0 FrameData[375]
port 305 nsew signal input
flabel metal2 s 0 197528 96 197608 0 FreeSans 320 0 0 0 FrameData[376]
port 306 nsew signal input
flabel metal2 s 0 198536 96 198616 0 FreeSans 320 0 0 0 FrameData[377]
port 307 nsew signal input
flabel metal2 s 0 199544 96 199624 0 FreeSans 320 0 0 0 FrameData[378]
port 308 nsew signal input
flabel metal2 s 0 200552 96 200632 0 FreeSans 320 0 0 0 FrameData[379]
port 309 nsew signal input
flabel metal2 s 0 662216 96 662296 0 FreeSans 320 0 0 0 FrameData[37]
port 310 nsew signal input
flabel metal2 s 0 201560 96 201640 0 FreeSans 320 0 0 0 FrameData[380]
port 311 nsew signal input
flabel metal2 s 0 202568 96 202648 0 FreeSans 320 0 0 0 FrameData[381]
port 312 nsew signal input
flabel metal2 s 0 203576 96 203656 0 FreeSans 320 0 0 0 FrameData[382]
port 313 nsew signal input
flabel metal2 s 0 204584 96 204664 0 FreeSans 320 0 0 0 FrameData[383]
port 314 nsew signal input
flabel metal2 s 0 124952 96 125032 0 FreeSans 320 0 0 0 FrameData[384]
port 315 nsew signal input
flabel metal2 s 0 125960 96 126040 0 FreeSans 320 0 0 0 FrameData[385]
port 316 nsew signal input
flabel metal2 s 0 126968 96 127048 0 FreeSans 320 0 0 0 FrameData[386]
port 317 nsew signal input
flabel metal2 s 0 127976 96 128056 0 FreeSans 320 0 0 0 FrameData[387]
port 318 nsew signal input
flabel metal2 s 0 128984 96 129064 0 FreeSans 320 0 0 0 FrameData[388]
port 319 nsew signal input
flabel metal2 s 0 129992 96 130072 0 FreeSans 320 0 0 0 FrameData[389]
port 320 nsew signal input
flabel metal2 s 0 663224 96 663304 0 FreeSans 320 0 0 0 FrameData[38]
port 321 nsew signal input
flabel metal2 s 0 131000 96 131080 0 FreeSans 320 0 0 0 FrameData[390]
port 322 nsew signal input
flabel metal2 s 0 132008 96 132088 0 FreeSans 320 0 0 0 FrameData[391]
port 323 nsew signal input
flabel metal2 s 0 133016 96 133096 0 FreeSans 320 0 0 0 FrameData[392]
port 324 nsew signal input
flabel metal2 s 0 134024 96 134104 0 FreeSans 320 0 0 0 FrameData[393]
port 325 nsew signal input
flabel metal2 s 0 135032 96 135112 0 FreeSans 320 0 0 0 FrameData[394]
port 326 nsew signal input
flabel metal2 s 0 136040 96 136120 0 FreeSans 320 0 0 0 FrameData[395]
port 327 nsew signal input
flabel metal2 s 0 137048 96 137128 0 FreeSans 320 0 0 0 FrameData[396]
port 328 nsew signal input
flabel metal2 s 0 138056 96 138136 0 FreeSans 320 0 0 0 FrameData[397]
port 329 nsew signal input
flabel metal2 s 0 139064 96 139144 0 FreeSans 320 0 0 0 FrameData[398]
port 330 nsew signal input
flabel metal2 s 0 140072 96 140152 0 FreeSans 320 0 0 0 FrameData[399]
port 331 nsew signal input
flabel metal2 s 0 664232 96 664312 0 FreeSans 320 0 0 0 FrameData[39]
port 332 nsew signal input
flabel metal2 s 0 691784 96 691864 0 FreeSans 320 0 0 0 FrameData[3]
port 333 nsew signal input
flabel metal2 s 0 141080 96 141160 0 FreeSans 320 0 0 0 FrameData[400]
port 334 nsew signal input
flabel metal2 s 0 142088 96 142168 0 FreeSans 320 0 0 0 FrameData[401]
port 335 nsew signal input
flabel metal2 s 0 143096 96 143176 0 FreeSans 320 0 0 0 FrameData[402]
port 336 nsew signal input
flabel metal2 s 0 144104 96 144184 0 FreeSans 320 0 0 0 FrameData[403]
port 337 nsew signal input
flabel metal2 s 0 145112 96 145192 0 FreeSans 320 0 0 0 FrameData[404]
port 338 nsew signal input
flabel metal2 s 0 146120 96 146200 0 FreeSans 320 0 0 0 FrameData[405]
port 339 nsew signal input
flabel metal2 s 0 147128 96 147208 0 FreeSans 320 0 0 0 FrameData[406]
port 340 nsew signal input
flabel metal2 s 0 148136 96 148216 0 FreeSans 320 0 0 0 FrameData[407]
port 341 nsew signal input
flabel metal2 s 0 149144 96 149224 0 FreeSans 320 0 0 0 FrameData[408]
port 342 nsew signal input
flabel metal2 s 0 150152 96 150232 0 FreeSans 320 0 0 0 FrameData[409]
port 343 nsew signal input
flabel metal2 s 0 665240 96 665320 0 FreeSans 320 0 0 0 FrameData[40]
port 344 nsew signal input
flabel metal2 s 0 151160 96 151240 0 FreeSans 320 0 0 0 FrameData[410]
port 345 nsew signal input
flabel metal2 s 0 152168 96 152248 0 FreeSans 320 0 0 0 FrameData[411]
port 346 nsew signal input
flabel metal2 s 0 153176 96 153256 0 FreeSans 320 0 0 0 FrameData[412]
port 347 nsew signal input
flabel metal2 s 0 154184 96 154264 0 FreeSans 320 0 0 0 FrameData[413]
port 348 nsew signal input
flabel metal2 s 0 155192 96 155272 0 FreeSans 320 0 0 0 FrameData[414]
port 349 nsew signal input
flabel metal2 s 0 156200 96 156280 0 FreeSans 320 0 0 0 FrameData[415]
port 350 nsew signal input
flabel metal2 s 0 76568 96 76648 0 FreeSans 320 0 0 0 FrameData[416]
port 351 nsew signal input
flabel metal2 s 0 77576 96 77656 0 FreeSans 320 0 0 0 FrameData[417]
port 352 nsew signal input
flabel metal2 s 0 78584 96 78664 0 FreeSans 320 0 0 0 FrameData[418]
port 353 nsew signal input
flabel metal2 s 0 79592 96 79672 0 FreeSans 320 0 0 0 FrameData[419]
port 354 nsew signal input
flabel metal2 s 0 666248 96 666328 0 FreeSans 320 0 0 0 FrameData[41]
port 355 nsew signal input
flabel metal2 s 0 80600 96 80680 0 FreeSans 320 0 0 0 FrameData[420]
port 356 nsew signal input
flabel metal2 s 0 81608 96 81688 0 FreeSans 320 0 0 0 FrameData[421]
port 357 nsew signal input
flabel metal2 s 0 82616 96 82696 0 FreeSans 320 0 0 0 FrameData[422]
port 358 nsew signal input
flabel metal2 s 0 83624 96 83704 0 FreeSans 320 0 0 0 FrameData[423]
port 359 nsew signal input
flabel metal2 s 0 84632 96 84712 0 FreeSans 320 0 0 0 FrameData[424]
port 360 nsew signal input
flabel metal2 s 0 85640 96 85720 0 FreeSans 320 0 0 0 FrameData[425]
port 361 nsew signal input
flabel metal2 s 0 86648 96 86728 0 FreeSans 320 0 0 0 FrameData[426]
port 362 nsew signal input
flabel metal2 s 0 87656 96 87736 0 FreeSans 320 0 0 0 FrameData[427]
port 363 nsew signal input
flabel metal2 s 0 88664 96 88744 0 FreeSans 320 0 0 0 FrameData[428]
port 364 nsew signal input
flabel metal2 s 0 89672 96 89752 0 FreeSans 320 0 0 0 FrameData[429]
port 365 nsew signal input
flabel metal2 s 0 667256 96 667336 0 FreeSans 320 0 0 0 FrameData[42]
port 366 nsew signal input
flabel metal2 s 0 90680 96 90760 0 FreeSans 320 0 0 0 FrameData[430]
port 367 nsew signal input
flabel metal2 s 0 91688 96 91768 0 FreeSans 320 0 0 0 FrameData[431]
port 368 nsew signal input
flabel metal2 s 0 92696 96 92776 0 FreeSans 320 0 0 0 FrameData[432]
port 369 nsew signal input
flabel metal2 s 0 93704 96 93784 0 FreeSans 320 0 0 0 FrameData[433]
port 370 nsew signal input
flabel metal2 s 0 94712 96 94792 0 FreeSans 320 0 0 0 FrameData[434]
port 371 nsew signal input
flabel metal2 s 0 95720 96 95800 0 FreeSans 320 0 0 0 FrameData[435]
port 372 nsew signal input
flabel metal2 s 0 96728 96 96808 0 FreeSans 320 0 0 0 FrameData[436]
port 373 nsew signal input
flabel metal2 s 0 97736 96 97816 0 FreeSans 320 0 0 0 FrameData[437]
port 374 nsew signal input
flabel metal2 s 0 98744 96 98824 0 FreeSans 320 0 0 0 FrameData[438]
port 375 nsew signal input
flabel metal2 s 0 99752 96 99832 0 FreeSans 320 0 0 0 FrameData[439]
port 376 nsew signal input
flabel metal2 s 0 668264 96 668344 0 FreeSans 320 0 0 0 FrameData[43]
port 377 nsew signal input
flabel metal2 s 0 100760 96 100840 0 FreeSans 320 0 0 0 FrameData[440]
port 378 nsew signal input
flabel metal2 s 0 101768 96 101848 0 FreeSans 320 0 0 0 FrameData[441]
port 379 nsew signal input
flabel metal2 s 0 102776 96 102856 0 FreeSans 320 0 0 0 FrameData[442]
port 380 nsew signal input
flabel metal2 s 0 103784 96 103864 0 FreeSans 320 0 0 0 FrameData[443]
port 381 nsew signal input
flabel metal2 s 0 104792 96 104872 0 FreeSans 320 0 0 0 FrameData[444]
port 382 nsew signal input
flabel metal2 s 0 105800 96 105880 0 FreeSans 320 0 0 0 FrameData[445]
port 383 nsew signal input
flabel metal2 s 0 106808 96 106888 0 FreeSans 320 0 0 0 FrameData[446]
port 384 nsew signal input
flabel metal2 s 0 107816 96 107896 0 FreeSans 320 0 0 0 FrameData[447]
port 385 nsew signal input
flabel metal2 s 0 28184 96 28264 0 FreeSans 320 0 0 0 FrameData[448]
port 386 nsew signal input
flabel metal2 s 0 29192 96 29272 0 FreeSans 320 0 0 0 FrameData[449]
port 387 nsew signal input
flabel metal2 s 0 669272 96 669352 0 FreeSans 320 0 0 0 FrameData[44]
port 388 nsew signal input
flabel metal2 s 0 30200 96 30280 0 FreeSans 320 0 0 0 FrameData[450]
port 389 nsew signal input
flabel metal2 s 0 31208 96 31288 0 FreeSans 320 0 0 0 FrameData[451]
port 390 nsew signal input
flabel metal2 s 0 32216 96 32296 0 FreeSans 320 0 0 0 FrameData[452]
port 391 nsew signal input
flabel metal2 s 0 33224 96 33304 0 FreeSans 320 0 0 0 FrameData[453]
port 392 nsew signal input
flabel metal2 s 0 34232 96 34312 0 FreeSans 320 0 0 0 FrameData[454]
port 393 nsew signal input
flabel metal2 s 0 35240 96 35320 0 FreeSans 320 0 0 0 FrameData[455]
port 394 nsew signal input
flabel metal2 s 0 36248 96 36328 0 FreeSans 320 0 0 0 FrameData[456]
port 395 nsew signal input
flabel metal2 s 0 37256 96 37336 0 FreeSans 320 0 0 0 FrameData[457]
port 396 nsew signal input
flabel metal2 s 0 38264 96 38344 0 FreeSans 320 0 0 0 FrameData[458]
port 397 nsew signal input
flabel metal2 s 0 39272 96 39352 0 FreeSans 320 0 0 0 FrameData[459]
port 398 nsew signal input
flabel metal2 s 0 670280 96 670360 0 FreeSans 320 0 0 0 FrameData[45]
port 399 nsew signal input
flabel metal2 s 0 40280 96 40360 0 FreeSans 320 0 0 0 FrameData[460]
port 400 nsew signal input
flabel metal2 s 0 41288 96 41368 0 FreeSans 320 0 0 0 FrameData[461]
port 401 nsew signal input
flabel metal2 s 0 42296 96 42376 0 FreeSans 320 0 0 0 FrameData[462]
port 402 nsew signal input
flabel metal2 s 0 43304 96 43384 0 FreeSans 320 0 0 0 FrameData[463]
port 403 nsew signal input
flabel metal2 s 0 44312 96 44392 0 FreeSans 320 0 0 0 FrameData[464]
port 404 nsew signal input
flabel metal2 s 0 45320 96 45400 0 FreeSans 320 0 0 0 FrameData[465]
port 405 nsew signal input
flabel metal2 s 0 46328 96 46408 0 FreeSans 320 0 0 0 FrameData[466]
port 406 nsew signal input
flabel metal2 s 0 47336 96 47416 0 FreeSans 320 0 0 0 FrameData[467]
port 407 nsew signal input
flabel metal2 s 0 48344 96 48424 0 FreeSans 320 0 0 0 FrameData[468]
port 408 nsew signal input
flabel metal2 s 0 49352 96 49432 0 FreeSans 320 0 0 0 FrameData[469]
port 409 nsew signal input
flabel metal2 s 0 671288 96 671368 0 FreeSans 320 0 0 0 FrameData[46]
port 410 nsew signal input
flabel metal2 s 0 50360 96 50440 0 FreeSans 320 0 0 0 FrameData[470]
port 411 nsew signal input
flabel metal2 s 0 51368 96 51448 0 FreeSans 320 0 0 0 FrameData[471]
port 412 nsew signal input
flabel metal2 s 0 52376 96 52456 0 FreeSans 320 0 0 0 FrameData[472]
port 413 nsew signal input
flabel metal2 s 0 53384 96 53464 0 FreeSans 320 0 0 0 FrameData[473]
port 414 nsew signal input
flabel metal2 s 0 54392 96 54472 0 FreeSans 320 0 0 0 FrameData[474]
port 415 nsew signal input
flabel metal2 s 0 55400 96 55480 0 FreeSans 320 0 0 0 FrameData[475]
port 416 nsew signal input
flabel metal2 s 0 56408 96 56488 0 FreeSans 320 0 0 0 FrameData[476]
port 417 nsew signal input
flabel metal2 s 0 57416 96 57496 0 FreeSans 320 0 0 0 FrameData[477]
port 418 nsew signal input
flabel metal2 s 0 58424 96 58504 0 FreeSans 320 0 0 0 FrameData[478]
port 419 nsew signal input
flabel metal2 s 0 59432 96 59512 0 FreeSans 320 0 0 0 FrameData[479]
port 420 nsew signal input
flabel metal2 s 0 672296 96 672376 0 FreeSans 320 0 0 0 FrameData[47]
port 421 nsew signal input
flabel metal2 s 0 1388 96 1468 0 FreeSans 320 0 0 0 FrameData[480]
port 422 nsew signal input
flabel metal2 s 0 1724 96 1804 0 FreeSans 320 0 0 0 FrameData[481]
port 423 nsew signal input
flabel metal2 s 0 2060 96 2140 0 FreeSans 320 0 0 0 FrameData[482]
port 424 nsew signal input
flabel metal2 s 0 2396 96 2476 0 FreeSans 320 0 0 0 FrameData[483]
port 425 nsew signal input
flabel metal2 s 0 2732 96 2812 0 FreeSans 320 0 0 0 FrameData[484]
port 426 nsew signal input
flabel metal2 s 0 3068 96 3148 0 FreeSans 320 0 0 0 FrameData[485]
port 427 nsew signal input
flabel metal2 s 0 3404 96 3484 0 FreeSans 320 0 0 0 FrameData[486]
port 428 nsew signal input
flabel metal2 s 0 3740 96 3820 0 FreeSans 320 0 0 0 FrameData[487]
port 429 nsew signal input
flabel metal2 s 0 4076 96 4156 0 FreeSans 320 0 0 0 FrameData[488]
port 430 nsew signal input
flabel metal2 s 0 4412 96 4492 0 FreeSans 320 0 0 0 FrameData[489]
port 431 nsew signal input
flabel metal2 s 0 673304 96 673384 0 FreeSans 320 0 0 0 FrameData[48]
port 432 nsew signal input
flabel metal2 s 0 4748 96 4828 0 FreeSans 320 0 0 0 FrameData[490]
port 433 nsew signal input
flabel metal2 s 0 5084 96 5164 0 FreeSans 320 0 0 0 FrameData[491]
port 434 nsew signal input
flabel metal2 s 0 5420 96 5500 0 FreeSans 320 0 0 0 FrameData[492]
port 435 nsew signal input
flabel metal2 s 0 5756 96 5836 0 FreeSans 320 0 0 0 FrameData[493]
port 436 nsew signal input
flabel metal2 s 0 6092 96 6172 0 FreeSans 320 0 0 0 FrameData[494]
port 437 nsew signal input
flabel metal2 s 0 6428 96 6508 0 FreeSans 320 0 0 0 FrameData[495]
port 438 nsew signal input
flabel metal2 s 0 6764 96 6844 0 FreeSans 320 0 0 0 FrameData[496]
port 439 nsew signal input
flabel metal2 s 0 7100 96 7180 0 FreeSans 320 0 0 0 FrameData[497]
port 440 nsew signal input
flabel metal2 s 0 7436 96 7516 0 FreeSans 320 0 0 0 FrameData[498]
port 441 nsew signal input
flabel metal2 s 0 7772 96 7852 0 FreeSans 320 0 0 0 FrameData[499]
port 442 nsew signal input
flabel metal2 s 0 674312 96 674392 0 FreeSans 320 0 0 0 FrameData[49]
port 443 nsew signal input
flabel metal2 s 0 692120 96 692200 0 FreeSans 320 0 0 0 FrameData[4]
port 444 nsew signal input
flabel metal2 s 0 8108 96 8188 0 FreeSans 320 0 0 0 FrameData[500]
port 445 nsew signal input
flabel metal2 s 0 8444 96 8524 0 FreeSans 320 0 0 0 FrameData[501]
port 446 nsew signal input
flabel metal2 s 0 8780 96 8860 0 FreeSans 320 0 0 0 FrameData[502]
port 447 nsew signal input
flabel metal2 s 0 9116 96 9196 0 FreeSans 320 0 0 0 FrameData[503]
port 448 nsew signal input
flabel metal2 s 0 9452 96 9532 0 FreeSans 320 0 0 0 FrameData[504]
port 449 nsew signal input
flabel metal2 s 0 9788 96 9868 0 FreeSans 320 0 0 0 FrameData[505]
port 450 nsew signal input
flabel metal2 s 0 10124 96 10204 0 FreeSans 320 0 0 0 FrameData[506]
port 451 nsew signal input
flabel metal2 s 0 10460 96 10540 0 FreeSans 320 0 0 0 FrameData[507]
port 452 nsew signal input
flabel metal2 s 0 10796 96 10876 0 FreeSans 320 0 0 0 FrameData[508]
port 453 nsew signal input
flabel metal2 s 0 11132 96 11212 0 FreeSans 320 0 0 0 FrameData[509]
port 454 nsew signal input
flabel metal2 s 0 675320 96 675400 0 FreeSans 320 0 0 0 FrameData[50]
port 455 nsew signal input
flabel metal2 s 0 11468 96 11548 0 FreeSans 320 0 0 0 FrameData[510]
port 456 nsew signal input
flabel metal2 s 0 11804 96 11884 0 FreeSans 320 0 0 0 FrameData[511]
port 457 nsew signal input
flabel metal2 s 0 676328 96 676408 0 FreeSans 320 0 0 0 FrameData[51]
port 458 nsew signal input
flabel metal2 s 0 677336 96 677416 0 FreeSans 320 0 0 0 FrameData[52]
port 459 nsew signal input
flabel metal2 s 0 678344 96 678424 0 FreeSans 320 0 0 0 FrameData[53]
port 460 nsew signal input
flabel metal2 s 0 679352 96 679432 0 FreeSans 320 0 0 0 FrameData[54]
port 461 nsew signal input
flabel metal2 s 0 680360 96 680440 0 FreeSans 320 0 0 0 FrameData[55]
port 462 nsew signal input
flabel metal2 s 0 681368 96 681448 0 FreeSans 320 0 0 0 FrameData[56]
port 463 nsew signal input
flabel metal2 s 0 682376 96 682456 0 FreeSans 320 0 0 0 FrameData[57]
port 464 nsew signal input
flabel metal2 s 0 683384 96 683464 0 FreeSans 320 0 0 0 FrameData[58]
port 465 nsew signal input
flabel metal2 s 0 684392 96 684472 0 FreeSans 320 0 0 0 FrameData[59]
port 466 nsew signal input
flabel metal2 s 0 692456 96 692536 0 FreeSans 320 0 0 0 FrameData[5]
port 467 nsew signal input
flabel metal2 s 0 685400 96 685480 0 FreeSans 320 0 0 0 FrameData[60]
port 468 nsew signal input
flabel metal2 s 0 686408 96 686488 0 FreeSans 320 0 0 0 FrameData[61]
port 469 nsew signal input
flabel metal2 s 0 687416 96 687496 0 FreeSans 320 0 0 0 FrameData[62]
port 470 nsew signal input
flabel metal2 s 0 688424 96 688504 0 FreeSans 320 0 0 0 FrameData[63]
port 471 nsew signal input
flabel metal2 s 0 608792 96 608872 0 FreeSans 320 0 0 0 FrameData[64]
port 472 nsew signal input
flabel metal2 s 0 609800 96 609880 0 FreeSans 320 0 0 0 FrameData[65]
port 473 nsew signal input
flabel metal2 s 0 610808 96 610888 0 FreeSans 320 0 0 0 FrameData[66]
port 474 nsew signal input
flabel metal2 s 0 611816 96 611896 0 FreeSans 320 0 0 0 FrameData[67]
port 475 nsew signal input
flabel metal2 s 0 612824 96 612904 0 FreeSans 320 0 0 0 FrameData[68]
port 476 nsew signal input
flabel metal2 s 0 613832 96 613912 0 FreeSans 320 0 0 0 FrameData[69]
port 477 nsew signal input
flabel metal2 s 0 692792 96 692872 0 FreeSans 320 0 0 0 FrameData[6]
port 478 nsew signal input
flabel metal2 s 0 614840 96 614920 0 FreeSans 320 0 0 0 FrameData[70]
port 479 nsew signal input
flabel metal2 s 0 615848 96 615928 0 FreeSans 320 0 0 0 FrameData[71]
port 480 nsew signal input
flabel metal2 s 0 616856 96 616936 0 FreeSans 320 0 0 0 FrameData[72]
port 481 nsew signal input
flabel metal2 s 0 617864 96 617944 0 FreeSans 320 0 0 0 FrameData[73]
port 482 nsew signal input
flabel metal2 s 0 618872 96 618952 0 FreeSans 320 0 0 0 FrameData[74]
port 483 nsew signal input
flabel metal2 s 0 619880 96 619960 0 FreeSans 320 0 0 0 FrameData[75]
port 484 nsew signal input
flabel metal2 s 0 620888 96 620968 0 FreeSans 320 0 0 0 FrameData[76]
port 485 nsew signal input
flabel metal2 s 0 621896 96 621976 0 FreeSans 320 0 0 0 FrameData[77]
port 486 nsew signal input
flabel metal2 s 0 622904 96 622984 0 FreeSans 320 0 0 0 FrameData[78]
port 487 nsew signal input
flabel metal2 s 0 623912 96 623992 0 FreeSans 320 0 0 0 FrameData[79]
port 488 nsew signal input
flabel metal2 s 0 693128 96 693208 0 FreeSans 320 0 0 0 FrameData[7]
port 489 nsew signal input
flabel metal2 s 0 624920 96 625000 0 FreeSans 320 0 0 0 FrameData[80]
port 490 nsew signal input
flabel metal2 s 0 625928 96 626008 0 FreeSans 320 0 0 0 FrameData[81]
port 491 nsew signal input
flabel metal2 s 0 626936 96 627016 0 FreeSans 320 0 0 0 FrameData[82]
port 492 nsew signal input
flabel metal2 s 0 627944 96 628024 0 FreeSans 320 0 0 0 FrameData[83]
port 493 nsew signal input
flabel metal2 s 0 628952 96 629032 0 FreeSans 320 0 0 0 FrameData[84]
port 494 nsew signal input
flabel metal2 s 0 629960 96 630040 0 FreeSans 320 0 0 0 FrameData[85]
port 495 nsew signal input
flabel metal2 s 0 630968 96 631048 0 FreeSans 320 0 0 0 FrameData[86]
port 496 nsew signal input
flabel metal2 s 0 631976 96 632056 0 FreeSans 320 0 0 0 FrameData[87]
port 497 nsew signal input
flabel metal2 s 0 632984 96 633064 0 FreeSans 320 0 0 0 FrameData[88]
port 498 nsew signal input
flabel metal2 s 0 633992 96 634072 0 FreeSans 320 0 0 0 FrameData[89]
port 499 nsew signal input
flabel metal2 s 0 693464 96 693544 0 FreeSans 320 0 0 0 FrameData[8]
port 500 nsew signal input
flabel metal2 s 0 635000 96 635080 0 FreeSans 320 0 0 0 FrameData[90]
port 501 nsew signal input
flabel metal2 s 0 636008 96 636088 0 FreeSans 320 0 0 0 FrameData[91]
port 502 nsew signal input
flabel metal2 s 0 637016 96 637096 0 FreeSans 320 0 0 0 FrameData[92]
port 503 nsew signal input
flabel metal2 s 0 638024 96 638104 0 FreeSans 320 0 0 0 FrameData[93]
port 504 nsew signal input
flabel metal2 s 0 639032 96 639112 0 FreeSans 320 0 0 0 FrameData[94]
port 505 nsew signal input
flabel metal2 s 0 640040 96 640120 0 FreeSans 320 0 0 0 FrameData[95]
port 506 nsew signal input
flabel metal2 s 0 560408 96 560488 0 FreeSans 320 0 0 0 FrameData[96]
port 507 nsew signal input
flabel metal2 s 0 561416 96 561496 0 FreeSans 320 0 0 0 FrameData[97]
port 508 nsew signal input
flabel metal2 s 0 562424 96 562504 0 FreeSans 320 0 0 0 FrameData[98]
port 509 nsew signal input
flabel metal2 s 0 563432 96 563512 0 FreeSans 320 0 0 0 FrameData[99]
port 510 nsew signal input
flabel metal2 s 0 693800 96 693880 0 FreeSans 320 0 0 0 FrameData[9]
port 511 nsew signal input
flabel metal3 s 1688 0 1768 80 0 FreeSans 320 0 0 0 FrameStrobe[0]
port 512 nsew signal input
flabel metal3 s 234680 0 234760 96 0 FreeSans 640 0 0 0 FrameStrobe[100]
port 513 nsew signal input
flabel metal3 s 235448 0 235528 96 0 FreeSans 640 0 0 0 FrameStrobe[101]
port 514 nsew signal input
flabel metal3 s 236216 0 236296 96 0 FreeSans 640 0 0 0 FrameStrobe[102]
port 515 nsew signal input
flabel metal3 s 236984 0 237064 96 0 FreeSans 640 0 0 0 FrameStrobe[103]
port 516 nsew signal input
flabel metal3 s 237752 0 237832 96 0 FreeSans 640 0 0 0 FrameStrobe[104]
port 517 nsew signal input
flabel metal3 s 238520 0 238600 96 0 FreeSans 640 0 0 0 FrameStrobe[105]
port 518 nsew signal input
flabel metal3 s 239288 0 239368 96 0 FreeSans 640 0 0 0 FrameStrobe[106]
port 519 nsew signal input
flabel metal3 s 240056 0 240136 96 0 FreeSans 640 0 0 0 FrameStrobe[107]
port 520 nsew signal input
flabel metal3 s 240824 0 240904 96 0 FreeSans 640 0 0 0 FrameStrobe[108]
port 521 nsew signal input
flabel metal3 s 241592 0 241672 96 0 FreeSans 640 0 0 0 FrameStrobe[109]
port 522 nsew signal input
flabel metal3 s 7448 0 7528 80 0 FreeSans 320 0 0 0 FrameStrobe[10]
port 523 nsew signal input
flabel metal3 s 242360 0 242440 96 0 FreeSans 640 0 0 0 FrameStrobe[110]
port 524 nsew signal input
flabel metal3 s 243128 0 243208 96 0 FreeSans 640 0 0 0 FrameStrobe[111]
port 525 nsew signal input
flabel metal3 s 243896 0 243976 96 0 FreeSans 640 0 0 0 FrameStrobe[112]
port 526 nsew signal input
flabel metal3 s 244664 0 244744 96 0 FreeSans 640 0 0 0 FrameStrobe[113]
port 527 nsew signal input
flabel metal3 s 245432 0 245512 96 0 FreeSans 640 0 0 0 FrameStrobe[114]
port 528 nsew signal input
flabel metal3 s 246200 0 246280 96 0 FreeSans 640 0 0 0 FrameStrobe[115]
port 529 nsew signal input
flabel metal3 s 246968 0 247048 96 0 FreeSans 640 0 0 0 FrameStrobe[116]
port 530 nsew signal input
flabel metal3 s 247736 0 247816 96 0 FreeSans 640 0 0 0 FrameStrobe[117]
port 531 nsew signal input
flabel metal3 s 248504 0 248584 96 0 FreeSans 640 0 0 0 FrameStrobe[118]
port 532 nsew signal input
flabel metal3 s 249272 0 249352 96 0 FreeSans 640 0 0 0 FrameStrobe[119]
port 533 nsew signal input
flabel metal3 s 8024 0 8104 80 0 FreeSans 320 0 0 0 FrameStrobe[11]
port 534 nsew signal input
flabel metal3 s 281048 0 281128 96 0 FreeSans 640 0 0 0 FrameStrobe[120]
port 535 nsew signal input
flabel metal3 s 281816 0 281896 96 0 FreeSans 640 0 0 0 FrameStrobe[121]
port 536 nsew signal input
flabel metal3 s 282584 0 282664 96 0 FreeSans 640 0 0 0 FrameStrobe[122]
port 537 nsew signal input
flabel metal3 s 283352 0 283432 96 0 FreeSans 640 0 0 0 FrameStrobe[123]
port 538 nsew signal input
flabel metal3 s 284120 0 284200 96 0 FreeSans 640 0 0 0 FrameStrobe[124]
port 539 nsew signal input
flabel metal3 s 284888 0 284968 96 0 FreeSans 640 0 0 0 FrameStrobe[125]
port 540 nsew signal input
flabel metal3 s 285656 0 285736 96 0 FreeSans 640 0 0 0 FrameStrobe[126]
port 541 nsew signal input
flabel metal3 s 286424 0 286504 96 0 FreeSans 640 0 0 0 FrameStrobe[127]
port 542 nsew signal input
flabel metal3 s 287192 0 287272 96 0 FreeSans 640 0 0 0 FrameStrobe[128]
port 543 nsew signal input
flabel metal3 s 287960 0 288040 96 0 FreeSans 640 0 0 0 FrameStrobe[129]
port 544 nsew signal input
flabel metal3 s 8600 0 8680 80 0 FreeSans 320 0 0 0 FrameStrobe[12]
port 545 nsew signal input
flabel metal3 s 288728 0 288808 96 0 FreeSans 640 0 0 0 FrameStrobe[130]
port 546 nsew signal input
flabel metal3 s 289496 0 289576 96 0 FreeSans 640 0 0 0 FrameStrobe[131]
port 547 nsew signal input
flabel metal3 s 290264 0 290344 96 0 FreeSans 640 0 0 0 FrameStrobe[132]
port 548 nsew signal input
flabel metal3 s 291032 0 291112 96 0 FreeSans 640 0 0 0 FrameStrobe[133]
port 549 nsew signal input
flabel metal3 s 291800 0 291880 96 0 FreeSans 640 0 0 0 FrameStrobe[134]
port 550 nsew signal input
flabel metal3 s 292568 0 292648 96 0 FreeSans 640 0 0 0 FrameStrobe[135]
port 551 nsew signal input
flabel metal3 s 293336 0 293416 96 0 FreeSans 640 0 0 0 FrameStrobe[136]
port 552 nsew signal input
flabel metal3 s 294104 0 294184 96 0 FreeSans 640 0 0 0 FrameStrobe[137]
port 553 nsew signal input
flabel metal3 s 294872 0 294952 96 0 FreeSans 640 0 0 0 FrameStrobe[138]
port 554 nsew signal input
flabel metal3 s 295640 0 295720 96 0 FreeSans 640 0 0 0 FrameStrobe[139]
port 555 nsew signal input
flabel metal3 s 9176 0 9256 80 0 FreeSans 320 0 0 0 FrameStrobe[13]
port 556 nsew signal input
flabel metal3 s 302840 0 302920 96 0 FreeSans 640 0 0 0 FrameStrobe[140]
port 557 nsew signal input
flabel metal3 s 304568 0 304648 96 0 FreeSans 640 0 0 0 FrameStrobe[141]
port 558 nsew signal input
flabel metal3 s 306296 0 306376 96 0 FreeSans 640 0 0 0 FrameStrobe[142]
port 559 nsew signal input
flabel metal3 s 308024 0 308104 96 0 FreeSans 640 0 0 0 FrameStrobe[143]
port 560 nsew signal input
flabel metal3 s 309752 0 309832 96 0 FreeSans 640 0 0 0 FrameStrobe[144]
port 561 nsew signal input
flabel metal3 s 311480 0 311560 96 0 FreeSans 640 0 0 0 FrameStrobe[145]
port 562 nsew signal input
flabel metal3 s 313208 0 313288 96 0 FreeSans 640 0 0 0 FrameStrobe[146]
port 563 nsew signal input
flabel metal3 s 314936 0 315016 96 0 FreeSans 640 0 0 0 FrameStrobe[147]
port 564 nsew signal input
flabel metal3 s 316664 0 316744 96 0 FreeSans 640 0 0 0 FrameStrobe[148]
port 565 nsew signal input
flabel metal3 s 318392 0 318472 96 0 FreeSans 640 0 0 0 FrameStrobe[149]
port 566 nsew signal input
flabel metal3 s 9752 0 9832 80 0 FreeSans 320 0 0 0 FrameStrobe[14]
port 567 nsew signal input
flabel metal3 s 320120 0 320200 96 0 FreeSans 640 0 0 0 FrameStrobe[150]
port 568 nsew signal input
flabel metal3 s 321848 0 321928 96 0 FreeSans 640 0 0 0 FrameStrobe[151]
port 569 nsew signal input
flabel metal3 s 323576 0 323656 96 0 FreeSans 640 0 0 0 FrameStrobe[152]
port 570 nsew signal input
flabel metal3 s 325304 0 325384 96 0 FreeSans 640 0 0 0 FrameStrobe[153]
port 571 nsew signal input
flabel metal3 s 327032 0 327112 96 0 FreeSans 640 0 0 0 FrameStrobe[154]
port 572 nsew signal input
flabel metal3 s 328760 0 328840 96 0 FreeSans 640 0 0 0 FrameStrobe[155]
port 573 nsew signal input
flabel metal3 s 330488 0 330568 96 0 FreeSans 640 0 0 0 FrameStrobe[156]
port 574 nsew signal input
flabel metal3 s 332216 0 332296 96 0 FreeSans 640 0 0 0 FrameStrobe[157]
port 575 nsew signal input
flabel metal3 s 333944 0 334024 96 0 FreeSans 640 0 0 0 FrameStrobe[158]
port 576 nsew signal input
flabel metal3 s 335672 0 335752 96 0 FreeSans 640 0 0 0 FrameStrobe[159]
port 577 nsew signal input
flabel metal3 s 10328 0 10408 80 0 FreeSans 320 0 0 0 FrameStrobe[15]
port 578 nsew signal input
flabel metal3 s 366680 0 366760 96 0 FreeSans 640 0 0 0 FrameStrobe[160]
port 579 nsew signal input
flabel metal3 s 367448 0 367528 96 0 FreeSans 640 0 0 0 FrameStrobe[161]
port 580 nsew signal input
flabel metal3 s 368216 0 368296 96 0 FreeSans 640 0 0 0 FrameStrobe[162]
port 581 nsew signal input
flabel metal3 s 368984 0 369064 96 0 FreeSans 640 0 0 0 FrameStrobe[163]
port 582 nsew signal input
flabel metal3 s 369752 0 369832 96 0 FreeSans 640 0 0 0 FrameStrobe[164]
port 583 nsew signal input
flabel metal3 s 370520 0 370600 96 0 FreeSans 640 0 0 0 FrameStrobe[165]
port 584 nsew signal input
flabel metal3 s 371288 0 371368 96 0 FreeSans 640 0 0 0 FrameStrobe[166]
port 585 nsew signal input
flabel metal3 s 372056 0 372136 96 0 FreeSans 640 0 0 0 FrameStrobe[167]
port 586 nsew signal input
flabel metal3 s 372824 0 372904 96 0 FreeSans 640 0 0 0 FrameStrobe[168]
port 587 nsew signal input
flabel metal3 s 373592 0 373672 96 0 FreeSans 640 0 0 0 FrameStrobe[169]
port 588 nsew signal input
flabel metal3 s 10904 0 10984 80 0 FreeSans 320 0 0 0 FrameStrobe[16]
port 589 nsew signal input
flabel metal3 s 374360 0 374440 96 0 FreeSans 640 0 0 0 FrameStrobe[170]
port 590 nsew signal input
flabel metal3 s 375128 0 375208 96 0 FreeSans 640 0 0 0 FrameStrobe[171]
port 591 nsew signal input
flabel metal3 s 375896 0 375976 96 0 FreeSans 640 0 0 0 FrameStrobe[172]
port 592 nsew signal input
flabel metal3 s 376664 0 376744 96 0 FreeSans 640 0 0 0 FrameStrobe[173]
port 593 nsew signal input
flabel metal3 s 377432 0 377512 96 0 FreeSans 640 0 0 0 FrameStrobe[174]
port 594 nsew signal input
flabel metal3 s 378200 0 378280 96 0 FreeSans 640 0 0 0 FrameStrobe[175]
port 595 nsew signal input
flabel metal3 s 378968 0 379048 96 0 FreeSans 640 0 0 0 FrameStrobe[176]
port 596 nsew signal input
flabel metal3 s 379736 0 379816 96 0 FreeSans 640 0 0 0 FrameStrobe[177]
port 597 nsew signal input
flabel metal3 s 380504 0 380584 96 0 FreeSans 640 0 0 0 FrameStrobe[178]
port 598 nsew signal input
flabel metal3 s 381272 0 381352 96 0 FreeSans 640 0 0 0 FrameStrobe[179]
port 599 nsew signal input
flabel metal3 s 11480 0 11560 80 0 FreeSans 320 0 0 0 FrameStrobe[17]
port 600 nsew signal input
flabel metal3 s 413048 0 413128 96 0 FreeSans 640 0 0 0 FrameStrobe[180]
port 601 nsew signal input
flabel metal3 s 413816 0 413896 96 0 FreeSans 640 0 0 0 FrameStrobe[181]
port 602 nsew signal input
flabel metal3 s 414584 0 414664 96 0 FreeSans 640 0 0 0 FrameStrobe[182]
port 603 nsew signal input
flabel metal3 s 415352 0 415432 96 0 FreeSans 640 0 0 0 FrameStrobe[183]
port 604 nsew signal input
flabel metal3 s 416120 0 416200 96 0 FreeSans 640 0 0 0 FrameStrobe[184]
port 605 nsew signal input
flabel metal3 s 416888 0 416968 96 0 FreeSans 640 0 0 0 FrameStrobe[185]
port 606 nsew signal input
flabel metal3 s 417656 0 417736 96 0 FreeSans 640 0 0 0 FrameStrobe[186]
port 607 nsew signal input
flabel metal3 s 418424 0 418504 96 0 FreeSans 640 0 0 0 FrameStrobe[187]
port 608 nsew signal input
flabel metal3 s 419192 0 419272 96 0 FreeSans 640 0 0 0 FrameStrobe[188]
port 609 nsew signal input
flabel metal3 s 419960 0 420040 96 0 FreeSans 640 0 0 0 FrameStrobe[189]
port 610 nsew signal input
flabel metal3 s 12056 0 12136 80 0 FreeSans 320 0 0 0 FrameStrobe[18]
port 611 nsew signal input
flabel metal3 s 420728 0 420808 96 0 FreeSans 640 0 0 0 FrameStrobe[190]
port 612 nsew signal input
flabel metal3 s 421496 0 421576 96 0 FreeSans 640 0 0 0 FrameStrobe[191]
port 613 nsew signal input
flabel metal3 s 422264 0 422344 96 0 FreeSans 640 0 0 0 FrameStrobe[192]
port 614 nsew signal input
flabel metal3 s 423032 0 423112 96 0 FreeSans 640 0 0 0 FrameStrobe[193]
port 615 nsew signal input
flabel metal3 s 423800 0 423880 96 0 FreeSans 640 0 0 0 FrameStrobe[194]
port 616 nsew signal input
flabel metal3 s 424568 0 424648 96 0 FreeSans 640 0 0 0 FrameStrobe[195]
port 617 nsew signal input
flabel metal3 s 425336 0 425416 96 0 FreeSans 640 0 0 0 FrameStrobe[196]
port 618 nsew signal input
flabel metal3 s 426104 0 426184 96 0 FreeSans 640 0 0 0 FrameStrobe[197]
port 619 nsew signal input
flabel metal3 s 426872 0 426952 96 0 FreeSans 640 0 0 0 FrameStrobe[198]
port 620 nsew signal input
flabel metal3 s 427640 0 427720 96 0 FreeSans 640 0 0 0 FrameStrobe[199]
port 621 nsew signal input
flabel metal3 s 12632 0 12712 80 0 FreeSans 320 0 0 0 FrameStrobe[19]
port 622 nsew signal input
flabel metal3 s 2264 0 2344 80 0 FreeSans 320 0 0 0 FrameStrobe[1]
port 623 nsew signal input
flabel metal3 s 432920 0 433000 80 0 FreeSans 320 0 0 0 FrameStrobe[200]
port 624 nsew signal input
flabel metal3 s 433880 0 433960 80 0 FreeSans 320 0 0 0 FrameStrobe[201]
port 625 nsew signal input
flabel metal3 s 434840 0 434920 80 0 FreeSans 320 0 0 0 FrameStrobe[202]
port 626 nsew signal input
flabel metal3 s 435800 0 435880 80 0 FreeSans 320 0 0 0 FrameStrobe[203]
port 627 nsew signal input
flabel metal3 s 436760 0 436840 80 0 FreeSans 320 0 0 0 FrameStrobe[204]
port 628 nsew signal input
flabel metal3 s 437720 0 437800 80 0 FreeSans 320 0 0 0 FrameStrobe[205]
port 629 nsew signal input
flabel metal3 s 438680 0 438760 80 0 FreeSans 320 0 0 0 FrameStrobe[206]
port 630 nsew signal input
flabel metal3 s 439640 0 439720 80 0 FreeSans 320 0 0 0 FrameStrobe[207]
port 631 nsew signal input
flabel metal3 s 440600 0 440680 80 0 FreeSans 320 0 0 0 FrameStrobe[208]
port 632 nsew signal input
flabel metal3 s 441560 0 441640 80 0 FreeSans 320 0 0 0 FrameStrobe[209]
port 633 nsew signal input
flabel metal3 s 17912 0 17992 96 0 FreeSans 640 0 0 0 FrameStrobe[20]
port 634 nsew signal input
flabel metal3 s 442520 0 442600 80 0 FreeSans 320 0 0 0 FrameStrobe[210]
port 635 nsew signal input
flabel metal3 s 443480 0 443560 80 0 FreeSans 320 0 0 0 FrameStrobe[211]
port 636 nsew signal input
flabel metal3 s 444440 0 444520 80 0 FreeSans 320 0 0 0 FrameStrobe[212]
port 637 nsew signal input
flabel metal3 s 445400 0 445480 80 0 FreeSans 320 0 0 0 FrameStrobe[213]
port 638 nsew signal input
flabel metal3 s 446360 0 446440 80 0 FreeSans 320 0 0 0 FrameStrobe[214]
port 639 nsew signal input
flabel metal3 s 447320 0 447400 80 0 FreeSans 320 0 0 0 FrameStrobe[215]
port 640 nsew signal input
flabel metal3 s 448280 0 448360 80 0 FreeSans 320 0 0 0 FrameStrobe[216]
port 641 nsew signal input
flabel metal3 s 449240 0 449320 80 0 FreeSans 320 0 0 0 FrameStrobe[217]
port 642 nsew signal input
flabel metal3 s 450200 0 450280 80 0 FreeSans 320 0 0 0 FrameStrobe[218]
port 643 nsew signal input
flabel metal3 s 451160 0 451240 80 0 FreeSans 320 0 0 0 FrameStrobe[219]
port 644 nsew signal input
flabel metal3 s 20024 0 20104 96 0 FreeSans 640 0 0 0 FrameStrobe[21]
port 645 nsew signal input
flabel metal3 s 22136 0 22216 96 0 FreeSans 640 0 0 0 FrameStrobe[22]
port 646 nsew signal input
flabel metal3 s 24248 0 24328 96 0 FreeSans 640 0 0 0 FrameStrobe[23]
port 647 nsew signal input
flabel metal3 s 26360 0 26440 96 0 FreeSans 640 0 0 0 FrameStrobe[24]
port 648 nsew signal input
flabel metal3 s 28472 0 28552 96 0 FreeSans 640 0 0 0 FrameStrobe[25]
port 649 nsew signal input
flabel metal3 s 30584 0 30664 96 0 FreeSans 640 0 0 0 FrameStrobe[26]
port 650 nsew signal input
flabel metal3 s 32696 0 32776 96 0 FreeSans 640 0 0 0 FrameStrobe[27]
port 651 nsew signal input
flabel metal3 s 34808 0 34888 96 0 FreeSans 640 0 0 0 FrameStrobe[28]
port 652 nsew signal input
flabel metal3 s 36920 0 37000 96 0 FreeSans 640 0 0 0 FrameStrobe[29]
port 653 nsew signal input
flabel metal3 s 2840 0 2920 80 0 FreeSans 320 0 0 0 FrameStrobe[2]
port 654 nsew signal input
flabel metal3 s 39032 0 39112 96 0 FreeSans 640 0 0 0 FrameStrobe[30]
port 655 nsew signal input
flabel metal3 s 41144 0 41224 96 0 FreeSans 640 0 0 0 FrameStrobe[31]
port 656 nsew signal input
flabel metal3 s 43256 0 43336 96 0 FreeSans 640 0 0 0 FrameStrobe[32]
port 657 nsew signal input
flabel metal3 s 45368 0 45448 96 0 FreeSans 640 0 0 0 FrameStrobe[33]
port 658 nsew signal input
flabel metal3 s 47480 0 47560 96 0 FreeSans 640 0 0 0 FrameStrobe[34]
port 659 nsew signal input
flabel metal3 s 49592 0 49672 96 0 FreeSans 640 0 0 0 FrameStrobe[35]
port 660 nsew signal input
flabel metal3 s 51704 0 51784 96 0 FreeSans 640 0 0 0 FrameStrobe[36]
port 661 nsew signal input
flabel metal3 s 53816 0 53896 96 0 FreeSans 640 0 0 0 FrameStrobe[37]
port 662 nsew signal input
flabel metal3 s 55928 0 56008 96 0 FreeSans 640 0 0 0 FrameStrobe[38]
port 663 nsew signal input
flabel metal3 s 58040 0 58120 96 0 FreeSans 640 0 0 0 FrameStrobe[39]
port 664 nsew signal input
flabel metal3 s 3416 0 3496 80 0 FreeSans 320 0 0 0 FrameStrobe[3]
port 665 nsew signal input
flabel metal3 s 74840 0 74920 96 0 FreeSans 640 0 0 0 FrameStrobe[40]
port 666 nsew signal input
flabel metal3 s 76376 0 76456 96 0 FreeSans 640 0 0 0 FrameStrobe[41]
port 667 nsew signal input
flabel metal3 s 77912 0 77992 96 0 FreeSans 640 0 0 0 FrameStrobe[42]
port 668 nsew signal input
flabel metal3 s 79448 0 79528 96 0 FreeSans 640 0 0 0 FrameStrobe[43]
port 669 nsew signal input
flabel metal3 s 80984 0 81064 96 0 FreeSans 640 0 0 0 FrameStrobe[44]
port 670 nsew signal input
flabel metal3 s 82520 0 82600 96 0 FreeSans 640 0 0 0 FrameStrobe[45]
port 671 nsew signal input
flabel metal3 s 84056 0 84136 96 0 FreeSans 640 0 0 0 FrameStrobe[46]
port 672 nsew signal input
flabel metal3 s 85592 0 85672 96 0 FreeSans 640 0 0 0 FrameStrobe[47]
port 673 nsew signal input
flabel metal3 s 87128 0 87208 96 0 FreeSans 640 0 0 0 FrameStrobe[48]
port 674 nsew signal input
flabel metal3 s 88664 0 88744 96 0 FreeSans 640 0 0 0 FrameStrobe[49]
port 675 nsew signal input
flabel metal3 s 3992 0 4072 80 0 FreeSans 320 0 0 0 FrameStrobe[4]
port 676 nsew signal input
flabel metal3 s 90200 0 90280 96 0 FreeSans 640 0 0 0 FrameStrobe[50]
port 677 nsew signal input
flabel metal3 s 91736 0 91816 96 0 FreeSans 640 0 0 0 FrameStrobe[51]
port 678 nsew signal input
flabel metal3 s 93272 0 93352 96 0 FreeSans 640 0 0 0 FrameStrobe[52]
port 679 nsew signal input
flabel metal3 s 94808 0 94888 96 0 FreeSans 640 0 0 0 FrameStrobe[53]
port 680 nsew signal input
flabel metal3 s 96344 0 96424 96 0 FreeSans 640 0 0 0 FrameStrobe[54]
port 681 nsew signal input
flabel metal3 s 97880 0 97960 96 0 FreeSans 640 0 0 0 FrameStrobe[55]
port 682 nsew signal input
flabel metal3 s 99416 0 99496 96 0 FreeSans 640 0 0 0 FrameStrobe[56]
port 683 nsew signal input
flabel metal3 s 100952 0 101032 96 0 FreeSans 640 0 0 0 FrameStrobe[57]
port 684 nsew signal input
flabel metal3 s 102488 0 102568 96 0 FreeSans 640 0 0 0 FrameStrobe[58]
port 685 nsew signal input
flabel metal3 s 104024 0 104104 96 0 FreeSans 640 0 0 0 FrameStrobe[59]
port 686 nsew signal input
flabel metal3 s 4568 0 4648 80 0 FreeSans 320 0 0 0 FrameStrobe[5]
port 687 nsew signal input
flabel metal3 s 118328 0 118408 96 0 FreeSans 640 0 0 0 FrameStrobe[60]
port 688 nsew signal input
flabel metal3 s 120056 0 120136 96 0 FreeSans 640 0 0 0 FrameStrobe[61]
port 689 nsew signal input
flabel metal3 s 121784 0 121864 96 0 FreeSans 640 0 0 0 FrameStrobe[62]
port 690 nsew signal input
flabel metal3 s 123512 0 123592 96 0 FreeSans 640 0 0 0 FrameStrobe[63]
port 691 nsew signal input
flabel metal3 s 125240 0 125320 96 0 FreeSans 640 0 0 0 FrameStrobe[64]
port 692 nsew signal input
flabel metal3 s 126968 0 127048 96 0 FreeSans 640 0 0 0 FrameStrobe[65]
port 693 nsew signal input
flabel metal3 s 128696 0 128776 96 0 FreeSans 640 0 0 0 FrameStrobe[66]
port 694 nsew signal input
flabel metal3 s 130424 0 130504 96 0 FreeSans 640 0 0 0 FrameStrobe[67]
port 695 nsew signal input
flabel metal3 s 132152 0 132232 96 0 FreeSans 640 0 0 0 FrameStrobe[68]
port 696 nsew signal input
flabel metal3 s 133880 0 133960 96 0 FreeSans 640 0 0 0 FrameStrobe[69]
port 697 nsew signal input
flabel metal3 s 5144 0 5224 80 0 FreeSans 320 0 0 0 FrameStrobe[6]
port 698 nsew signal input
flabel metal3 s 135608 0 135688 96 0 FreeSans 640 0 0 0 FrameStrobe[70]
port 699 nsew signal input
flabel metal3 s 137336 0 137416 96 0 FreeSans 640 0 0 0 FrameStrobe[71]
port 700 nsew signal input
flabel metal3 s 139064 0 139144 96 0 FreeSans 640 0 0 0 FrameStrobe[72]
port 701 nsew signal input
flabel metal3 s 140792 0 140872 96 0 FreeSans 640 0 0 0 FrameStrobe[73]
port 702 nsew signal input
flabel metal3 s 142520 0 142600 96 0 FreeSans 640 0 0 0 FrameStrobe[74]
port 703 nsew signal input
flabel metal3 s 144248 0 144328 96 0 FreeSans 640 0 0 0 FrameStrobe[75]
port 704 nsew signal input
flabel metal3 s 145976 0 146056 96 0 FreeSans 640 0 0 0 FrameStrobe[76]
port 705 nsew signal input
flabel metal3 s 147704 0 147784 96 0 FreeSans 640 0 0 0 FrameStrobe[77]
port 706 nsew signal input
flabel metal3 s 149432 0 149512 96 0 FreeSans 640 0 0 0 FrameStrobe[78]
port 707 nsew signal input
flabel metal3 s 151160 0 151240 96 0 FreeSans 640 0 0 0 FrameStrobe[79]
port 708 nsew signal input
flabel metal3 s 5720 0 5800 80 0 FreeSans 320 0 0 0 FrameStrobe[7]
port 709 nsew signal input
flabel metal3 s 157016 0 157096 96 0 FreeSans 640 0 0 0 FrameStrobe[80]
port 710 nsew signal input
flabel metal3 s 159512 0 159592 96 0 FreeSans 640 0 0 0 FrameStrobe[81]
port 711 nsew signal input
flabel metal3 s 162008 0 162088 96 0 FreeSans 640 0 0 0 FrameStrobe[82]
port 712 nsew signal input
flabel metal3 s 164504 0 164584 96 0 FreeSans 640 0 0 0 FrameStrobe[83]
port 713 nsew signal input
flabel metal3 s 167000 0 167080 96 0 FreeSans 640 0 0 0 FrameStrobe[84]
port 714 nsew signal input
flabel metal3 s 169496 0 169576 96 0 FreeSans 640 0 0 0 FrameStrobe[85]
port 715 nsew signal input
flabel metal3 s 171992 0 172072 96 0 FreeSans 640 0 0 0 FrameStrobe[86]
port 716 nsew signal input
flabel metal3 s 174488 0 174568 96 0 FreeSans 640 0 0 0 FrameStrobe[87]
port 717 nsew signal input
flabel metal3 s 176984 0 177064 96 0 FreeSans 640 0 0 0 FrameStrobe[88]
port 718 nsew signal input
flabel metal3 s 179480 0 179560 96 0 FreeSans 640 0 0 0 FrameStrobe[89]
port 719 nsew signal input
flabel metal3 s 6296 0 6376 80 0 FreeSans 320 0 0 0 FrameStrobe[8]
port 720 nsew signal input
flabel metal3 s 181976 0 182056 96 0 FreeSans 640 0 0 0 FrameStrobe[90]
port 721 nsew signal input
flabel metal3 s 184472 0 184552 96 0 FreeSans 640 0 0 0 FrameStrobe[91]
port 722 nsew signal input
flabel metal3 s 186968 0 187048 96 0 FreeSans 640 0 0 0 FrameStrobe[92]
port 723 nsew signal input
flabel metal3 s 189464 0 189544 96 0 FreeSans 640 0 0 0 FrameStrobe[93]
port 724 nsew signal input
flabel metal3 s 191960 0 192040 96 0 FreeSans 640 0 0 0 FrameStrobe[94]
port 725 nsew signal input
flabel metal3 s 194456 0 194536 96 0 FreeSans 640 0 0 0 FrameStrobe[95]
port 726 nsew signal input
flabel metal3 s 196952 0 197032 96 0 FreeSans 640 0 0 0 FrameStrobe[96]
port 727 nsew signal input
flabel metal3 s 199448 0 199528 96 0 FreeSans 640 0 0 0 FrameStrobe[97]
port 728 nsew signal input
flabel metal3 s 201944 0 202024 96 0 FreeSans 640 0 0 0 FrameStrobe[98]
port 729 nsew signal input
flabel metal3 s 204440 0 204520 96 0 FreeSans 640 0 0 0 FrameStrobe[99]
port 730 nsew signal input
flabel metal3 s 6872 0 6952 80 0 FreeSans 320 0 0 0 FrameStrobe[9]
port 731 nsew signal input
flabel metal2 s 0 208616 96 208696 0 FreeSans 320 0 0 0 Tile_X0Y10_A_I_top
port 732 nsew signal output
flabel metal2 s 0 207608 96 207688 0 FreeSans 320 0 0 0 Tile_X0Y10_A_O_top
port 733 nsew signal input
flabel metal2 s 0 209624 96 209704 0 FreeSans 320 0 0 0 Tile_X0Y10_A_T_top
port 734 nsew signal output
flabel metal2 s 0 213656 96 213736 0 FreeSans 320 0 0 0 Tile_X0Y10_A_config_C_bit0
port 735 nsew signal output
flabel metal2 s 0 214664 96 214744 0 FreeSans 320 0 0 0 Tile_X0Y10_A_config_C_bit1
port 736 nsew signal output
flabel metal2 s 0 215672 96 215752 0 FreeSans 320 0 0 0 Tile_X0Y10_A_config_C_bit2
port 737 nsew signal output
flabel metal2 s 0 216680 96 216760 0 FreeSans 320 0 0 0 Tile_X0Y10_A_config_C_bit3
port 738 nsew signal output
flabel metal2 s 0 211640 96 211720 0 FreeSans 320 0 0 0 Tile_X0Y10_B_I_top
port 739 nsew signal output
flabel metal2 s 0 210632 96 210712 0 FreeSans 320 0 0 0 Tile_X0Y10_B_O_top
port 740 nsew signal input
flabel metal2 s 0 212648 96 212728 0 FreeSans 320 0 0 0 Tile_X0Y10_B_T_top
port 741 nsew signal output
flabel metal2 s 0 217688 96 217768 0 FreeSans 320 0 0 0 Tile_X0Y10_B_config_C_bit0
port 742 nsew signal output
flabel metal2 s 0 218696 96 218776 0 FreeSans 320 0 0 0 Tile_X0Y10_B_config_C_bit1
port 743 nsew signal output
flabel metal2 s 0 219704 96 219784 0 FreeSans 320 0 0 0 Tile_X0Y10_B_config_C_bit2
port 744 nsew signal output
flabel metal2 s 0 220712 96 220792 0 FreeSans 320 0 0 0 Tile_X0Y10_B_config_C_bit3
port 745 nsew signal output
flabel metal2 s 0 160232 96 160312 0 FreeSans 320 0 0 0 Tile_X0Y11_A_I_top
port 746 nsew signal output
flabel metal2 s 0 159224 96 159304 0 FreeSans 320 0 0 0 Tile_X0Y11_A_O_top
port 747 nsew signal input
flabel metal2 s 0 161240 96 161320 0 FreeSans 320 0 0 0 Tile_X0Y11_A_T_top
port 748 nsew signal output
flabel metal2 s 0 165272 96 165352 0 FreeSans 320 0 0 0 Tile_X0Y11_A_config_C_bit0
port 749 nsew signal output
flabel metal2 s 0 166280 96 166360 0 FreeSans 320 0 0 0 Tile_X0Y11_A_config_C_bit1
port 750 nsew signal output
flabel metal2 s 0 167288 96 167368 0 FreeSans 320 0 0 0 Tile_X0Y11_A_config_C_bit2
port 751 nsew signal output
flabel metal2 s 0 168296 96 168376 0 FreeSans 320 0 0 0 Tile_X0Y11_A_config_C_bit3
port 752 nsew signal output
flabel metal2 s 0 163256 96 163336 0 FreeSans 320 0 0 0 Tile_X0Y11_B_I_top
port 753 nsew signal output
flabel metal2 s 0 162248 96 162328 0 FreeSans 320 0 0 0 Tile_X0Y11_B_O_top
port 754 nsew signal input
flabel metal2 s 0 164264 96 164344 0 FreeSans 320 0 0 0 Tile_X0Y11_B_T_top
port 755 nsew signal output
flabel metal2 s 0 169304 96 169384 0 FreeSans 320 0 0 0 Tile_X0Y11_B_config_C_bit0
port 756 nsew signal output
flabel metal2 s 0 170312 96 170392 0 FreeSans 320 0 0 0 Tile_X0Y11_B_config_C_bit1
port 757 nsew signal output
flabel metal2 s 0 171320 96 171400 0 FreeSans 320 0 0 0 Tile_X0Y11_B_config_C_bit2
port 758 nsew signal output
flabel metal2 s 0 172328 96 172408 0 FreeSans 320 0 0 0 Tile_X0Y11_B_config_C_bit3
port 759 nsew signal output
flabel metal2 s 0 111848 96 111928 0 FreeSans 320 0 0 0 Tile_X0Y12_A_I_top
port 760 nsew signal output
flabel metal2 s 0 110840 96 110920 0 FreeSans 320 0 0 0 Tile_X0Y12_A_O_top
port 761 nsew signal input
flabel metal2 s 0 112856 96 112936 0 FreeSans 320 0 0 0 Tile_X0Y12_A_T_top
port 762 nsew signal output
flabel metal2 s 0 116888 96 116968 0 FreeSans 320 0 0 0 Tile_X0Y12_A_config_C_bit0
port 763 nsew signal output
flabel metal2 s 0 117896 96 117976 0 FreeSans 320 0 0 0 Tile_X0Y12_A_config_C_bit1
port 764 nsew signal output
flabel metal2 s 0 118904 96 118984 0 FreeSans 320 0 0 0 Tile_X0Y12_A_config_C_bit2
port 765 nsew signal output
flabel metal2 s 0 119912 96 119992 0 FreeSans 320 0 0 0 Tile_X0Y12_A_config_C_bit3
port 766 nsew signal output
flabel metal2 s 0 114872 96 114952 0 FreeSans 320 0 0 0 Tile_X0Y12_B_I_top
port 767 nsew signal output
flabel metal2 s 0 113864 96 113944 0 FreeSans 320 0 0 0 Tile_X0Y12_B_O_top
port 768 nsew signal input
flabel metal2 s 0 115880 96 115960 0 FreeSans 320 0 0 0 Tile_X0Y12_B_T_top
port 769 nsew signal output
flabel metal2 s 0 120920 96 121000 0 FreeSans 320 0 0 0 Tile_X0Y12_B_config_C_bit0
port 770 nsew signal output
flabel metal2 s 0 121928 96 122008 0 FreeSans 320 0 0 0 Tile_X0Y12_B_config_C_bit1
port 771 nsew signal output
flabel metal2 s 0 122936 96 123016 0 FreeSans 320 0 0 0 Tile_X0Y12_B_config_C_bit2
port 772 nsew signal output
flabel metal2 s 0 123944 96 124024 0 FreeSans 320 0 0 0 Tile_X0Y12_B_config_C_bit3
port 773 nsew signal output
flabel metal2 s 0 63464 96 63544 0 FreeSans 320 0 0 0 Tile_X0Y13_A_I_top
port 774 nsew signal output
flabel metal2 s 0 62456 96 62536 0 FreeSans 320 0 0 0 Tile_X0Y13_A_O_top
port 775 nsew signal input
flabel metal2 s 0 64472 96 64552 0 FreeSans 320 0 0 0 Tile_X0Y13_A_T_top
port 776 nsew signal output
flabel metal2 s 0 68504 96 68584 0 FreeSans 320 0 0 0 Tile_X0Y13_A_config_C_bit0
port 777 nsew signal output
flabel metal2 s 0 69512 96 69592 0 FreeSans 320 0 0 0 Tile_X0Y13_A_config_C_bit1
port 778 nsew signal output
flabel metal2 s 0 70520 96 70600 0 FreeSans 320 0 0 0 Tile_X0Y13_A_config_C_bit2
port 779 nsew signal output
flabel metal2 s 0 71528 96 71608 0 FreeSans 320 0 0 0 Tile_X0Y13_A_config_C_bit3
port 780 nsew signal output
flabel metal2 s 0 66488 96 66568 0 FreeSans 320 0 0 0 Tile_X0Y13_B_I_top
port 781 nsew signal output
flabel metal2 s 0 65480 96 65560 0 FreeSans 320 0 0 0 Tile_X0Y13_B_O_top
port 782 nsew signal input
flabel metal2 s 0 67496 96 67576 0 FreeSans 320 0 0 0 Tile_X0Y13_B_T_top
port 783 nsew signal output
flabel metal2 s 0 72536 96 72616 0 FreeSans 320 0 0 0 Tile_X0Y13_B_config_C_bit0
port 784 nsew signal output
flabel metal2 s 0 73544 96 73624 0 FreeSans 320 0 0 0 Tile_X0Y13_B_config_C_bit1
port 785 nsew signal output
flabel metal2 s 0 74552 96 74632 0 FreeSans 320 0 0 0 Tile_X0Y13_B_config_C_bit2
port 786 nsew signal output
flabel metal2 s 0 75560 96 75640 0 FreeSans 320 0 0 0 Tile_X0Y13_B_config_C_bit3
port 787 nsew signal output
flabel metal2 s 0 15080 96 15160 0 FreeSans 320 0 0 0 Tile_X0Y14_A_I_top
port 788 nsew signal output
flabel metal2 s 0 13232 96 13312 0 FreeSans 320 0 0 0 Tile_X0Y14_A_O_top
port 789 nsew signal input
flabel metal2 s 0 16088 96 16168 0 FreeSans 320 0 0 0 Tile_X0Y14_A_T_top
port 790 nsew signal output
flabel metal2 s 0 20120 96 20200 0 FreeSans 320 0 0 0 Tile_X0Y14_A_config_C_bit0
port 791 nsew signal output
flabel metal2 s 0 21128 96 21208 0 FreeSans 320 0 0 0 Tile_X0Y14_A_config_C_bit1
port 792 nsew signal output
flabel metal2 s 0 22136 96 22216 0 FreeSans 320 0 0 0 Tile_X0Y14_A_config_C_bit2
port 793 nsew signal output
flabel metal2 s 0 23144 96 23224 0 FreeSans 320 0 0 0 Tile_X0Y14_A_config_C_bit3
port 794 nsew signal output
flabel metal2 s 0 18104 96 18184 0 FreeSans 320 0 0 0 Tile_X0Y14_B_I_top
port 795 nsew signal output
flabel metal2 s 0 17096 96 17176 0 FreeSans 320 0 0 0 Tile_X0Y14_B_O_top
port 796 nsew signal input
flabel metal2 s 0 19112 96 19192 0 FreeSans 320 0 0 0 Tile_X0Y14_B_T_top
port 797 nsew signal output
flabel metal2 s 0 24152 96 24232 0 FreeSans 320 0 0 0 Tile_X0Y14_B_config_C_bit0
port 798 nsew signal output
flabel metal2 s 0 25160 96 25240 0 FreeSans 320 0 0 0 Tile_X0Y14_B_config_C_bit1
port 799 nsew signal output
flabel metal2 s 0 26168 96 26248 0 FreeSans 320 0 0 0 Tile_X0Y14_B_config_C_bit2
port 800 nsew signal output
flabel metal2 s 0 27176 96 27256 0 FreeSans 320 0 0 0 Tile_X0Y14_B_config_C_bit3
port 801 nsew signal output
flabel metal2 s 0 644072 96 644152 0 FreeSans 320 0 0 0 Tile_X0Y1_A_I_top
port 802 nsew signal output
flabel metal2 s 0 643064 96 643144 0 FreeSans 320 0 0 0 Tile_X0Y1_A_O_top
port 803 nsew signal input
flabel metal2 s 0 645080 96 645160 0 FreeSans 320 0 0 0 Tile_X0Y1_A_T_top
port 804 nsew signal output
flabel metal2 s 0 649112 96 649192 0 FreeSans 320 0 0 0 Tile_X0Y1_A_config_C_bit0
port 805 nsew signal output
flabel metal2 s 0 650120 96 650200 0 FreeSans 320 0 0 0 Tile_X0Y1_A_config_C_bit1
port 806 nsew signal output
flabel metal2 s 0 651128 96 651208 0 FreeSans 320 0 0 0 Tile_X0Y1_A_config_C_bit2
port 807 nsew signal output
flabel metal2 s 0 652136 96 652216 0 FreeSans 320 0 0 0 Tile_X0Y1_A_config_C_bit3
port 808 nsew signal output
flabel metal2 s 0 647096 96 647176 0 FreeSans 320 0 0 0 Tile_X0Y1_B_I_top
port 809 nsew signal output
flabel metal2 s 0 646088 96 646168 0 FreeSans 320 0 0 0 Tile_X0Y1_B_O_top
port 810 nsew signal input
flabel metal2 s 0 648104 96 648184 0 FreeSans 320 0 0 0 Tile_X0Y1_B_T_top
port 811 nsew signal output
flabel metal2 s 0 653144 96 653224 0 FreeSans 320 0 0 0 Tile_X0Y1_B_config_C_bit0
port 812 nsew signal output
flabel metal2 s 0 654152 96 654232 0 FreeSans 320 0 0 0 Tile_X0Y1_B_config_C_bit1
port 813 nsew signal output
flabel metal2 s 0 655160 96 655240 0 FreeSans 320 0 0 0 Tile_X0Y1_B_config_C_bit2
port 814 nsew signal output
flabel metal2 s 0 656168 96 656248 0 FreeSans 320 0 0 0 Tile_X0Y1_B_config_C_bit3
port 815 nsew signal output
flabel metal2 s 0 595688 96 595768 0 FreeSans 320 0 0 0 Tile_X0Y2_A_I_top
port 816 nsew signal output
flabel metal2 s 0 594680 96 594760 0 FreeSans 320 0 0 0 Tile_X0Y2_A_O_top
port 817 nsew signal input
flabel metal2 s 0 596696 96 596776 0 FreeSans 320 0 0 0 Tile_X0Y2_A_T_top
port 818 nsew signal output
flabel metal2 s 0 600728 96 600808 0 FreeSans 320 0 0 0 Tile_X0Y2_A_config_C_bit0
port 819 nsew signal output
flabel metal2 s 0 601736 96 601816 0 FreeSans 320 0 0 0 Tile_X0Y2_A_config_C_bit1
port 820 nsew signal output
flabel metal2 s 0 602744 96 602824 0 FreeSans 320 0 0 0 Tile_X0Y2_A_config_C_bit2
port 821 nsew signal output
flabel metal2 s 0 603752 96 603832 0 FreeSans 320 0 0 0 Tile_X0Y2_A_config_C_bit3
port 822 nsew signal output
flabel metal2 s 0 598712 96 598792 0 FreeSans 320 0 0 0 Tile_X0Y2_B_I_top
port 823 nsew signal output
flabel metal2 s 0 597704 96 597784 0 FreeSans 320 0 0 0 Tile_X0Y2_B_O_top
port 824 nsew signal input
flabel metal2 s 0 599720 96 599800 0 FreeSans 320 0 0 0 Tile_X0Y2_B_T_top
port 825 nsew signal output
flabel metal2 s 0 604760 96 604840 0 FreeSans 320 0 0 0 Tile_X0Y2_B_config_C_bit0
port 826 nsew signal output
flabel metal2 s 0 605768 96 605848 0 FreeSans 320 0 0 0 Tile_X0Y2_B_config_C_bit1
port 827 nsew signal output
flabel metal2 s 0 606776 96 606856 0 FreeSans 320 0 0 0 Tile_X0Y2_B_config_C_bit2
port 828 nsew signal output
flabel metal2 s 0 607784 96 607864 0 FreeSans 320 0 0 0 Tile_X0Y2_B_config_C_bit3
port 829 nsew signal output
flabel metal2 s 0 547304 96 547384 0 FreeSans 320 0 0 0 Tile_X0Y3_A_I_top
port 830 nsew signal output
flabel metal2 s 0 546296 96 546376 0 FreeSans 320 0 0 0 Tile_X0Y3_A_O_top
port 831 nsew signal input
flabel metal2 s 0 548312 96 548392 0 FreeSans 320 0 0 0 Tile_X0Y3_A_T_top
port 832 nsew signal output
flabel metal2 s 0 552344 96 552424 0 FreeSans 320 0 0 0 Tile_X0Y3_A_config_C_bit0
port 833 nsew signal output
flabel metal2 s 0 553352 96 553432 0 FreeSans 320 0 0 0 Tile_X0Y3_A_config_C_bit1
port 834 nsew signal output
flabel metal2 s 0 554360 96 554440 0 FreeSans 320 0 0 0 Tile_X0Y3_A_config_C_bit2
port 835 nsew signal output
flabel metal2 s 0 555368 96 555448 0 FreeSans 320 0 0 0 Tile_X0Y3_A_config_C_bit3
port 836 nsew signal output
flabel metal2 s 0 550328 96 550408 0 FreeSans 320 0 0 0 Tile_X0Y3_B_I_top
port 837 nsew signal output
flabel metal2 s 0 549320 96 549400 0 FreeSans 320 0 0 0 Tile_X0Y3_B_O_top
port 838 nsew signal input
flabel metal2 s 0 551336 96 551416 0 FreeSans 320 0 0 0 Tile_X0Y3_B_T_top
port 839 nsew signal output
flabel metal2 s 0 556376 96 556456 0 FreeSans 320 0 0 0 Tile_X0Y3_B_config_C_bit0
port 840 nsew signal output
flabel metal2 s 0 557384 96 557464 0 FreeSans 320 0 0 0 Tile_X0Y3_B_config_C_bit1
port 841 nsew signal output
flabel metal2 s 0 558392 96 558472 0 FreeSans 320 0 0 0 Tile_X0Y3_B_config_C_bit2
port 842 nsew signal output
flabel metal2 s 0 559400 96 559480 0 FreeSans 320 0 0 0 Tile_X0Y3_B_config_C_bit3
port 843 nsew signal output
flabel metal2 s 0 498920 96 499000 0 FreeSans 320 0 0 0 Tile_X0Y4_A_I_top
port 844 nsew signal output
flabel metal2 s 0 497912 96 497992 0 FreeSans 320 0 0 0 Tile_X0Y4_A_O_top
port 845 nsew signal input
flabel metal2 s 0 499928 96 500008 0 FreeSans 320 0 0 0 Tile_X0Y4_A_T_top
port 846 nsew signal output
flabel metal2 s 0 503960 96 504040 0 FreeSans 320 0 0 0 Tile_X0Y4_A_config_C_bit0
port 847 nsew signal output
flabel metal2 s 0 504968 96 505048 0 FreeSans 320 0 0 0 Tile_X0Y4_A_config_C_bit1
port 848 nsew signal output
flabel metal2 s 0 505976 96 506056 0 FreeSans 320 0 0 0 Tile_X0Y4_A_config_C_bit2
port 849 nsew signal output
flabel metal2 s 0 506984 96 507064 0 FreeSans 320 0 0 0 Tile_X0Y4_A_config_C_bit3
port 850 nsew signal output
flabel metal2 s 0 501944 96 502024 0 FreeSans 320 0 0 0 Tile_X0Y4_B_I_top
port 851 nsew signal output
flabel metal2 s 0 500936 96 501016 0 FreeSans 320 0 0 0 Tile_X0Y4_B_O_top
port 852 nsew signal input
flabel metal2 s 0 502952 96 503032 0 FreeSans 320 0 0 0 Tile_X0Y4_B_T_top
port 853 nsew signal output
flabel metal2 s 0 507992 96 508072 0 FreeSans 320 0 0 0 Tile_X0Y4_B_config_C_bit0
port 854 nsew signal output
flabel metal2 s 0 509000 96 509080 0 FreeSans 320 0 0 0 Tile_X0Y4_B_config_C_bit1
port 855 nsew signal output
flabel metal2 s 0 510008 96 510088 0 FreeSans 320 0 0 0 Tile_X0Y4_B_config_C_bit2
port 856 nsew signal output
flabel metal2 s 0 511016 96 511096 0 FreeSans 320 0 0 0 Tile_X0Y4_B_config_C_bit3
port 857 nsew signal output
flabel metal2 s 0 450536 96 450616 0 FreeSans 320 0 0 0 Tile_X0Y5_A_I_top
port 858 nsew signal output
flabel metal2 s 0 449528 96 449608 0 FreeSans 320 0 0 0 Tile_X0Y5_A_O_top
port 859 nsew signal input
flabel metal2 s 0 451544 96 451624 0 FreeSans 320 0 0 0 Tile_X0Y5_A_T_top
port 860 nsew signal output
flabel metal2 s 0 455576 96 455656 0 FreeSans 320 0 0 0 Tile_X0Y5_A_config_C_bit0
port 861 nsew signal output
flabel metal2 s 0 456584 96 456664 0 FreeSans 320 0 0 0 Tile_X0Y5_A_config_C_bit1
port 862 nsew signal output
flabel metal2 s 0 457592 96 457672 0 FreeSans 320 0 0 0 Tile_X0Y5_A_config_C_bit2
port 863 nsew signal output
flabel metal2 s 0 458600 96 458680 0 FreeSans 320 0 0 0 Tile_X0Y5_A_config_C_bit3
port 864 nsew signal output
flabel metal2 s 0 453560 96 453640 0 FreeSans 320 0 0 0 Tile_X0Y5_B_I_top
port 865 nsew signal output
flabel metal2 s 0 452552 96 452632 0 FreeSans 320 0 0 0 Tile_X0Y5_B_O_top
port 866 nsew signal input
flabel metal2 s 0 454568 96 454648 0 FreeSans 320 0 0 0 Tile_X0Y5_B_T_top
port 867 nsew signal output
flabel metal2 s 0 459608 96 459688 0 FreeSans 320 0 0 0 Tile_X0Y5_B_config_C_bit0
port 868 nsew signal output
flabel metal2 s 0 460616 96 460696 0 FreeSans 320 0 0 0 Tile_X0Y5_B_config_C_bit1
port 869 nsew signal output
flabel metal2 s 0 461624 96 461704 0 FreeSans 320 0 0 0 Tile_X0Y5_B_config_C_bit2
port 870 nsew signal output
flabel metal2 s 0 462632 96 462712 0 FreeSans 320 0 0 0 Tile_X0Y5_B_config_C_bit3
port 871 nsew signal output
flabel metal2 s 0 402152 96 402232 0 FreeSans 320 0 0 0 Tile_X0Y6_A_I_top
port 872 nsew signal output
flabel metal2 s 0 401144 96 401224 0 FreeSans 320 0 0 0 Tile_X0Y6_A_O_top
port 873 nsew signal input
flabel metal2 s 0 403160 96 403240 0 FreeSans 320 0 0 0 Tile_X0Y6_A_T_top
port 874 nsew signal output
flabel metal2 s 0 407192 96 407272 0 FreeSans 320 0 0 0 Tile_X0Y6_A_config_C_bit0
port 875 nsew signal output
flabel metal2 s 0 408200 96 408280 0 FreeSans 320 0 0 0 Tile_X0Y6_A_config_C_bit1
port 876 nsew signal output
flabel metal2 s 0 409208 96 409288 0 FreeSans 320 0 0 0 Tile_X0Y6_A_config_C_bit2
port 877 nsew signal output
flabel metal2 s 0 410216 96 410296 0 FreeSans 320 0 0 0 Tile_X0Y6_A_config_C_bit3
port 878 nsew signal output
flabel metal2 s 0 405176 96 405256 0 FreeSans 320 0 0 0 Tile_X0Y6_B_I_top
port 879 nsew signal output
flabel metal2 s 0 404168 96 404248 0 FreeSans 320 0 0 0 Tile_X0Y6_B_O_top
port 880 nsew signal input
flabel metal2 s 0 406184 96 406264 0 FreeSans 320 0 0 0 Tile_X0Y6_B_T_top
port 881 nsew signal output
flabel metal2 s 0 411224 96 411304 0 FreeSans 320 0 0 0 Tile_X0Y6_B_config_C_bit0
port 882 nsew signal output
flabel metal2 s 0 412232 96 412312 0 FreeSans 320 0 0 0 Tile_X0Y6_B_config_C_bit1
port 883 nsew signal output
flabel metal2 s 0 413240 96 413320 0 FreeSans 320 0 0 0 Tile_X0Y6_B_config_C_bit2
port 884 nsew signal output
flabel metal2 s 0 414248 96 414328 0 FreeSans 320 0 0 0 Tile_X0Y6_B_config_C_bit3
port 885 nsew signal output
flabel metal2 s 0 353768 96 353848 0 FreeSans 320 0 0 0 Tile_X0Y7_A_I_top
port 886 nsew signal output
flabel metal2 s 0 352760 96 352840 0 FreeSans 320 0 0 0 Tile_X0Y7_A_O_top
port 887 nsew signal input
flabel metal2 s 0 354776 96 354856 0 FreeSans 320 0 0 0 Tile_X0Y7_A_T_top
port 888 nsew signal output
flabel metal2 s 0 358808 96 358888 0 FreeSans 320 0 0 0 Tile_X0Y7_A_config_C_bit0
port 889 nsew signal output
flabel metal2 s 0 359816 96 359896 0 FreeSans 320 0 0 0 Tile_X0Y7_A_config_C_bit1
port 890 nsew signal output
flabel metal2 s 0 360824 96 360904 0 FreeSans 320 0 0 0 Tile_X0Y7_A_config_C_bit2
port 891 nsew signal output
flabel metal2 s 0 361832 96 361912 0 FreeSans 320 0 0 0 Tile_X0Y7_A_config_C_bit3
port 892 nsew signal output
flabel metal2 s 0 356792 96 356872 0 FreeSans 320 0 0 0 Tile_X0Y7_B_I_top
port 893 nsew signal output
flabel metal2 s 0 355784 96 355864 0 FreeSans 320 0 0 0 Tile_X0Y7_B_O_top
port 894 nsew signal input
flabel metal2 s 0 357800 96 357880 0 FreeSans 320 0 0 0 Tile_X0Y7_B_T_top
port 895 nsew signal output
flabel metal2 s 0 362840 96 362920 0 FreeSans 320 0 0 0 Tile_X0Y7_B_config_C_bit0
port 896 nsew signal output
flabel metal2 s 0 363848 96 363928 0 FreeSans 320 0 0 0 Tile_X0Y7_B_config_C_bit1
port 897 nsew signal output
flabel metal2 s 0 364856 96 364936 0 FreeSans 320 0 0 0 Tile_X0Y7_B_config_C_bit2
port 898 nsew signal output
flabel metal2 s 0 365864 96 365944 0 FreeSans 320 0 0 0 Tile_X0Y7_B_config_C_bit3
port 899 nsew signal output
flabel metal2 s 0 305384 96 305464 0 FreeSans 320 0 0 0 Tile_X0Y8_A_I_top
port 900 nsew signal output
flabel metal2 s 0 304376 96 304456 0 FreeSans 320 0 0 0 Tile_X0Y8_A_O_top
port 901 nsew signal input
flabel metal2 s 0 306392 96 306472 0 FreeSans 320 0 0 0 Tile_X0Y8_A_T_top
port 902 nsew signal output
flabel metal2 s 0 310424 96 310504 0 FreeSans 320 0 0 0 Tile_X0Y8_A_config_C_bit0
port 903 nsew signal output
flabel metal2 s 0 311432 96 311512 0 FreeSans 320 0 0 0 Tile_X0Y8_A_config_C_bit1
port 904 nsew signal output
flabel metal2 s 0 312440 96 312520 0 FreeSans 320 0 0 0 Tile_X0Y8_A_config_C_bit2
port 905 nsew signal output
flabel metal2 s 0 313448 96 313528 0 FreeSans 320 0 0 0 Tile_X0Y8_A_config_C_bit3
port 906 nsew signal output
flabel metal2 s 0 308408 96 308488 0 FreeSans 320 0 0 0 Tile_X0Y8_B_I_top
port 907 nsew signal output
flabel metal2 s 0 307400 96 307480 0 FreeSans 320 0 0 0 Tile_X0Y8_B_O_top
port 908 nsew signal input
flabel metal2 s 0 309416 96 309496 0 FreeSans 320 0 0 0 Tile_X0Y8_B_T_top
port 909 nsew signal output
flabel metal2 s 0 314456 96 314536 0 FreeSans 320 0 0 0 Tile_X0Y8_B_config_C_bit0
port 910 nsew signal output
flabel metal2 s 0 315464 96 315544 0 FreeSans 320 0 0 0 Tile_X0Y8_B_config_C_bit1
port 911 nsew signal output
flabel metal2 s 0 316472 96 316552 0 FreeSans 320 0 0 0 Tile_X0Y8_B_config_C_bit2
port 912 nsew signal output
flabel metal2 s 0 317480 96 317560 0 FreeSans 320 0 0 0 Tile_X0Y8_B_config_C_bit3
port 913 nsew signal output
flabel metal2 s 0 257000 96 257080 0 FreeSans 320 0 0 0 Tile_X0Y9_A_I_top
port 914 nsew signal output
flabel metal2 s 0 255992 96 256072 0 FreeSans 320 0 0 0 Tile_X0Y9_A_O_top
port 915 nsew signal input
flabel metal2 s 0 258008 96 258088 0 FreeSans 320 0 0 0 Tile_X0Y9_A_T_top
port 916 nsew signal output
flabel metal2 s 0 262040 96 262120 0 FreeSans 320 0 0 0 Tile_X0Y9_A_config_C_bit0
port 917 nsew signal output
flabel metal2 s 0 263048 96 263128 0 FreeSans 320 0 0 0 Tile_X0Y9_A_config_C_bit1
port 918 nsew signal output
flabel metal2 s 0 264056 96 264136 0 FreeSans 320 0 0 0 Tile_X0Y9_A_config_C_bit2
port 919 nsew signal output
flabel metal2 s 0 265064 96 265144 0 FreeSans 320 0 0 0 Tile_X0Y9_A_config_C_bit3
port 920 nsew signal output
flabel metal2 s 0 260024 96 260104 0 FreeSans 320 0 0 0 Tile_X0Y9_B_I_top
port 921 nsew signal output
flabel metal2 s 0 259016 96 259096 0 FreeSans 320 0 0 0 Tile_X0Y9_B_O_top
port 922 nsew signal input
flabel metal2 s 0 261032 96 261112 0 FreeSans 320 0 0 0 Tile_X0Y9_B_T_top
port 923 nsew signal output
flabel metal2 s 0 266072 96 266152 0 FreeSans 320 0 0 0 Tile_X0Y9_B_config_C_bit0
port 924 nsew signal output
flabel metal2 s 0 267080 96 267160 0 FreeSans 320 0 0 0 Tile_X0Y9_B_config_C_bit1
port 925 nsew signal output
flabel metal2 s 0 268088 96 268168 0 FreeSans 320 0 0 0 Tile_X0Y9_B_config_C_bit2
port 926 nsew signal output
flabel metal2 s 0 269096 96 269176 0 FreeSans 320 0 0 0 Tile_X0Y9_B_config_C_bit3
port 927 nsew signal output
flabel metal2 s 452544 226760 452640 226840 0 FreeSans 320 0 0 0 Tile_X10Y10_ADDR_SRAM0
port 928 nsew signal output
flabel metal2 s 452544 227264 452640 227344 0 FreeSans 320 0 0 0 Tile_X10Y10_ADDR_SRAM1
port 929 nsew signal output
flabel metal2 s 452544 227768 452640 227848 0 FreeSans 320 0 0 0 Tile_X10Y10_ADDR_SRAM2
port 930 nsew signal output
flabel metal2 s 452544 228272 452640 228352 0 FreeSans 320 0 0 0 Tile_X10Y10_ADDR_SRAM3
port 931 nsew signal output
flabel metal2 s 452544 228776 452640 228856 0 FreeSans 320 0 0 0 Tile_X10Y10_ADDR_SRAM4
port 932 nsew signal output
flabel metal2 s 452544 229280 452640 229360 0 FreeSans 320 0 0 0 Tile_X10Y10_ADDR_SRAM5
port 933 nsew signal output
flabel metal2 s 452544 229784 452640 229864 0 FreeSans 320 0 0 0 Tile_X10Y10_ADDR_SRAM6
port 934 nsew signal output
flabel metal2 s 452544 230288 452640 230368 0 FreeSans 320 0 0 0 Tile_X10Y10_ADDR_SRAM7
port 935 nsew signal output
flabel metal2 s 452544 230792 452640 230872 0 FreeSans 320 0 0 0 Tile_X10Y10_ADDR_SRAM8
port 936 nsew signal output
flabel metal2 s 452544 231296 452640 231376 0 FreeSans 320 0 0 0 Tile_X10Y10_ADDR_SRAM9
port 937 nsew signal output
flabel metal2 s 452544 231800 452640 231880 0 FreeSans 320 0 0 0 Tile_X10Y10_BM_SRAM0
port 938 nsew signal output
flabel metal2 s 452544 232304 452640 232384 0 FreeSans 320 0 0 0 Tile_X10Y10_BM_SRAM1
port 939 nsew signal output
flabel metal2 s 452544 236840 452640 236920 0 FreeSans 320 0 0 0 Tile_X10Y10_BM_SRAM10
port 940 nsew signal output
flabel metal2 s 452544 237344 452640 237424 0 FreeSans 320 0 0 0 Tile_X10Y10_BM_SRAM11
port 941 nsew signal output
flabel metal2 s 452544 237848 452640 237928 0 FreeSans 320 0 0 0 Tile_X10Y10_BM_SRAM12
port 942 nsew signal output
flabel metal2 s 452544 238352 452640 238432 0 FreeSans 320 0 0 0 Tile_X10Y10_BM_SRAM13
port 943 nsew signal output
flabel metal2 s 452544 238856 452640 238936 0 FreeSans 320 0 0 0 Tile_X10Y10_BM_SRAM14
port 944 nsew signal output
flabel metal2 s 452544 239360 452640 239440 0 FreeSans 320 0 0 0 Tile_X10Y10_BM_SRAM15
port 945 nsew signal output
flabel metal2 s 452544 239864 452640 239944 0 FreeSans 320 0 0 0 Tile_X10Y10_BM_SRAM16
port 946 nsew signal output
flabel metal2 s 452544 240368 452640 240448 0 FreeSans 320 0 0 0 Tile_X10Y10_BM_SRAM17
port 947 nsew signal output
flabel metal2 s 452544 240872 452640 240952 0 FreeSans 320 0 0 0 Tile_X10Y10_BM_SRAM18
port 948 nsew signal output
flabel metal2 s 452544 241376 452640 241456 0 FreeSans 320 0 0 0 Tile_X10Y10_BM_SRAM19
port 949 nsew signal output
flabel metal2 s 452544 232808 452640 232888 0 FreeSans 320 0 0 0 Tile_X10Y10_BM_SRAM2
port 950 nsew signal output
flabel metal2 s 452544 241880 452640 241960 0 FreeSans 320 0 0 0 Tile_X10Y10_BM_SRAM20
port 951 nsew signal output
flabel metal2 s 452544 242384 452640 242464 0 FreeSans 320 0 0 0 Tile_X10Y10_BM_SRAM21
port 952 nsew signal output
flabel metal2 s 452544 242888 452640 242968 0 FreeSans 320 0 0 0 Tile_X10Y10_BM_SRAM22
port 953 nsew signal output
flabel metal2 s 452544 243392 452640 243472 0 FreeSans 320 0 0 0 Tile_X10Y10_BM_SRAM23
port 954 nsew signal output
flabel metal2 s 452544 243896 452640 243976 0 FreeSans 320 0 0 0 Tile_X10Y10_BM_SRAM24
port 955 nsew signal output
flabel metal2 s 452544 244400 452640 244480 0 FreeSans 320 0 0 0 Tile_X10Y10_BM_SRAM25
port 956 nsew signal output
flabel metal2 s 452544 244904 452640 244984 0 FreeSans 320 0 0 0 Tile_X10Y10_BM_SRAM26
port 957 nsew signal output
flabel metal2 s 452544 245408 452640 245488 0 FreeSans 320 0 0 0 Tile_X10Y10_BM_SRAM27
port 958 nsew signal output
flabel metal2 s 452544 245912 452640 245992 0 FreeSans 320 0 0 0 Tile_X10Y10_BM_SRAM28
port 959 nsew signal output
flabel metal2 s 452544 246416 452640 246496 0 FreeSans 320 0 0 0 Tile_X10Y10_BM_SRAM29
port 960 nsew signal output
flabel metal2 s 452544 233312 452640 233392 0 FreeSans 320 0 0 0 Tile_X10Y10_BM_SRAM3
port 961 nsew signal output
flabel metal2 s 452544 246920 452640 247000 0 FreeSans 320 0 0 0 Tile_X10Y10_BM_SRAM30
port 962 nsew signal output
flabel metal2 s 452544 247424 452640 247504 0 FreeSans 320 0 0 0 Tile_X10Y10_BM_SRAM31
port 963 nsew signal output
flabel metal2 s 452544 233816 452640 233896 0 FreeSans 320 0 0 0 Tile_X10Y10_BM_SRAM4
port 964 nsew signal output
flabel metal2 s 452544 234320 452640 234400 0 FreeSans 320 0 0 0 Tile_X10Y10_BM_SRAM5
port 965 nsew signal output
flabel metal2 s 452544 234824 452640 234904 0 FreeSans 320 0 0 0 Tile_X10Y10_BM_SRAM6
port 966 nsew signal output
flabel metal2 s 452544 235328 452640 235408 0 FreeSans 320 0 0 0 Tile_X10Y10_BM_SRAM7
port 967 nsew signal output
flabel metal2 s 452544 235832 452640 235912 0 FreeSans 320 0 0 0 Tile_X10Y10_BM_SRAM8
port 968 nsew signal output
flabel metal2 s 452544 236336 452640 236416 0 FreeSans 320 0 0 0 Tile_X10Y10_BM_SRAM9
port 969 nsew signal output
flabel metal2 s 452544 247928 452640 248008 0 FreeSans 320 0 0 0 Tile_X10Y10_CLK_SRAM
port 970 nsew signal output
flabel metal2 s 452544 210128 452640 210208 0 FreeSans 320 0 0 0 Tile_X10Y10_CONFIGURED_top
port 971 nsew signal input
flabel metal2 s 452544 248432 452640 248512 0 FreeSans 320 0 0 0 Tile_X10Y10_DIN_SRAM0
port 972 nsew signal output
flabel metal2 s 452544 248936 452640 249016 0 FreeSans 320 0 0 0 Tile_X10Y10_DIN_SRAM1
port 973 nsew signal output
flabel metal2 s 452544 253472 452640 253552 0 FreeSans 320 0 0 0 Tile_X10Y10_DIN_SRAM10
port 974 nsew signal output
flabel metal2 s 452544 253976 452640 254056 0 FreeSans 320 0 0 0 Tile_X10Y10_DIN_SRAM11
port 975 nsew signal output
flabel metal2 s 452544 254480 452640 254560 0 FreeSans 320 0 0 0 Tile_X10Y10_DIN_SRAM12
port 976 nsew signal output
flabel metal2 s 452544 254984 452640 255064 0 FreeSans 320 0 0 0 Tile_X10Y10_DIN_SRAM13
port 977 nsew signal output
flabel metal2 s 452544 255488 452640 255568 0 FreeSans 320 0 0 0 Tile_X10Y10_DIN_SRAM14
port 978 nsew signal output
flabel metal2 s 452544 255992 452640 256072 0 FreeSans 320 0 0 0 Tile_X10Y10_DIN_SRAM15
port 979 nsew signal output
flabel metal2 s 452544 256496 452640 256576 0 FreeSans 320 0 0 0 Tile_X10Y10_DIN_SRAM16
port 980 nsew signal output
flabel metal2 s 452544 257000 452640 257080 0 FreeSans 320 0 0 0 Tile_X10Y10_DIN_SRAM17
port 981 nsew signal output
flabel metal2 s 452544 257504 452640 257584 0 FreeSans 320 0 0 0 Tile_X10Y10_DIN_SRAM18
port 982 nsew signal output
flabel metal2 s 452544 258008 452640 258088 0 FreeSans 320 0 0 0 Tile_X10Y10_DIN_SRAM19
port 983 nsew signal output
flabel metal2 s 452544 249440 452640 249520 0 FreeSans 320 0 0 0 Tile_X10Y10_DIN_SRAM2
port 984 nsew signal output
flabel metal2 s 452544 258512 452640 258592 0 FreeSans 320 0 0 0 Tile_X10Y10_DIN_SRAM20
port 985 nsew signal output
flabel metal2 s 452544 259016 452640 259096 0 FreeSans 320 0 0 0 Tile_X10Y10_DIN_SRAM21
port 986 nsew signal output
flabel metal2 s 452544 259520 452640 259600 0 FreeSans 320 0 0 0 Tile_X10Y10_DIN_SRAM22
port 987 nsew signal output
flabel metal2 s 452544 260024 452640 260104 0 FreeSans 320 0 0 0 Tile_X10Y10_DIN_SRAM23
port 988 nsew signal output
flabel metal2 s 452544 260528 452640 260608 0 FreeSans 320 0 0 0 Tile_X10Y10_DIN_SRAM24
port 989 nsew signal output
flabel metal2 s 452544 261032 452640 261112 0 FreeSans 320 0 0 0 Tile_X10Y10_DIN_SRAM25
port 990 nsew signal output
flabel metal2 s 452544 261536 452640 261616 0 FreeSans 320 0 0 0 Tile_X10Y10_DIN_SRAM26
port 991 nsew signal output
flabel metal2 s 452544 262040 452640 262120 0 FreeSans 320 0 0 0 Tile_X10Y10_DIN_SRAM27
port 992 nsew signal output
flabel metal2 s 452544 262544 452640 262624 0 FreeSans 320 0 0 0 Tile_X10Y10_DIN_SRAM28
port 993 nsew signal output
flabel metal2 s 452544 263048 452640 263128 0 FreeSans 320 0 0 0 Tile_X10Y10_DIN_SRAM29
port 994 nsew signal output
flabel metal2 s 452544 249944 452640 250024 0 FreeSans 320 0 0 0 Tile_X10Y10_DIN_SRAM3
port 995 nsew signal output
flabel metal2 s 452544 263552 452640 263632 0 FreeSans 320 0 0 0 Tile_X10Y10_DIN_SRAM30
port 996 nsew signal output
flabel metal2 s 452544 264056 452640 264136 0 FreeSans 320 0 0 0 Tile_X10Y10_DIN_SRAM31
port 997 nsew signal output
flabel metal2 s 452544 250448 452640 250528 0 FreeSans 320 0 0 0 Tile_X10Y10_DIN_SRAM4
port 998 nsew signal output
flabel metal2 s 452544 250952 452640 251032 0 FreeSans 320 0 0 0 Tile_X10Y10_DIN_SRAM5
port 999 nsew signal output
flabel metal2 s 452544 251456 452640 251536 0 FreeSans 320 0 0 0 Tile_X10Y10_DIN_SRAM6
port 1000 nsew signal output
flabel metal2 s 452544 251960 452640 252040 0 FreeSans 320 0 0 0 Tile_X10Y10_DIN_SRAM7
port 1001 nsew signal output
flabel metal2 s 452544 252464 452640 252544 0 FreeSans 320 0 0 0 Tile_X10Y10_DIN_SRAM8
port 1002 nsew signal output
flabel metal2 s 452544 252968 452640 253048 0 FreeSans 320 0 0 0 Tile_X10Y10_DIN_SRAM9
port 1003 nsew signal output
flabel metal2 s 452544 210632 452640 210712 0 FreeSans 320 0 0 0 Tile_X10Y10_DOUT_SRAM0
port 1004 nsew signal input
flabel metal2 s 452544 211136 452640 211216 0 FreeSans 320 0 0 0 Tile_X10Y10_DOUT_SRAM1
port 1005 nsew signal input
flabel metal2 s 452544 215672 452640 215752 0 FreeSans 320 0 0 0 Tile_X10Y10_DOUT_SRAM10
port 1006 nsew signal input
flabel metal2 s 452544 216176 452640 216256 0 FreeSans 320 0 0 0 Tile_X10Y10_DOUT_SRAM11
port 1007 nsew signal input
flabel metal2 s 452544 216680 452640 216760 0 FreeSans 320 0 0 0 Tile_X10Y10_DOUT_SRAM12
port 1008 nsew signal input
flabel metal2 s 452544 217184 452640 217264 0 FreeSans 320 0 0 0 Tile_X10Y10_DOUT_SRAM13
port 1009 nsew signal input
flabel metal2 s 452544 217688 452640 217768 0 FreeSans 320 0 0 0 Tile_X10Y10_DOUT_SRAM14
port 1010 nsew signal input
flabel metal2 s 452544 218192 452640 218272 0 FreeSans 320 0 0 0 Tile_X10Y10_DOUT_SRAM15
port 1011 nsew signal input
flabel metal2 s 452544 218696 452640 218776 0 FreeSans 320 0 0 0 Tile_X10Y10_DOUT_SRAM16
port 1012 nsew signal input
flabel metal2 s 452544 219200 452640 219280 0 FreeSans 320 0 0 0 Tile_X10Y10_DOUT_SRAM17
port 1013 nsew signal input
flabel metal2 s 452544 219704 452640 219784 0 FreeSans 320 0 0 0 Tile_X10Y10_DOUT_SRAM18
port 1014 nsew signal input
flabel metal2 s 452544 220208 452640 220288 0 FreeSans 320 0 0 0 Tile_X10Y10_DOUT_SRAM19
port 1015 nsew signal input
flabel metal2 s 452544 211640 452640 211720 0 FreeSans 320 0 0 0 Tile_X10Y10_DOUT_SRAM2
port 1016 nsew signal input
flabel metal2 s 452544 220712 452640 220792 0 FreeSans 320 0 0 0 Tile_X10Y10_DOUT_SRAM20
port 1017 nsew signal input
flabel metal2 s 452544 221216 452640 221296 0 FreeSans 320 0 0 0 Tile_X10Y10_DOUT_SRAM21
port 1018 nsew signal input
flabel metal2 s 452544 221720 452640 221800 0 FreeSans 320 0 0 0 Tile_X10Y10_DOUT_SRAM22
port 1019 nsew signal input
flabel metal2 s 452544 222224 452640 222304 0 FreeSans 320 0 0 0 Tile_X10Y10_DOUT_SRAM23
port 1020 nsew signal input
flabel metal2 s 452544 222728 452640 222808 0 FreeSans 320 0 0 0 Tile_X10Y10_DOUT_SRAM24
port 1021 nsew signal input
flabel metal2 s 452544 223232 452640 223312 0 FreeSans 320 0 0 0 Tile_X10Y10_DOUT_SRAM25
port 1022 nsew signal input
flabel metal2 s 452544 223736 452640 223816 0 FreeSans 320 0 0 0 Tile_X10Y10_DOUT_SRAM26
port 1023 nsew signal input
flabel metal2 s 452544 224240 452640 224320 0 FreeSans 320 0 0 0 Tile_X10Y10_DOUT_SRAM27
port 1024 nsew signal input
flabel metal2 s 452544 224744 452640 224824 0 FreeSans 320 0 0 0 Tile_X10Y10_DOUT_SRAM28
port 1025 nsew signal input
flabel metal2 s 452544 225248 452640 225328 0 FreeSans 320 0 0 0 Tile_X10Y10_DOUT_SRAM29
port 1026 nsew signal input
flabel metal2 s 452544 212144 452640 212224 0 FreeSans 320 0 0 0 Tile_X10Y10_DOUT_SRAM3
port 1027 nsew signal input
flabel metal2 s 452544 225752 452640 225832 0 FreeSans 320 0 0 0 Tile_X10Y10_DOUT_SRAM30
port 1028 nsew signal input
flabel metal2 s 452544 226256 452640 226336 0 FreeSans 320 0 0 0 Tile_X10Y10_DOUT_SRAM31
port 1029 nsew signal input
flabel metal2 s 452544 212648 452640 212728 0 FreeSans 320 0 0 0 Tile_X10Y10_DOUT_SRAM4
port 1030 nsew signal input
flabel metal2 s 452544 213152 452640 213232 0 FreeSans 320 0 0 0 Tile_X10Y10_DOUT_SRAM5
port 1031 nsew signal input
flabel metal2 s 452544 213656 452640 213736 0 FreeSans 320 0 0 0 Tile_X10Y10_DOUT_SRAM6
port 1032 nsew signal input
flabel metal2 s 452544 214160 452640 214240 0 FreeSans 320 0 0 0 Tile_X10Y10_DOUT_SRAM7
port 1033 nsew signal input
flabel metal2 s 452544 214664 452640 214744 0 FreeSans 320 0 0 0 Tile_X10Y10_DOUT_SRAM8
port 1034 nsew signal input
flabel metal2 s 452544 215168 452640 215248 0 FreeSans 320 0 0 0 Tile_X10Y10_DOUT_SRAM9
port 1035 nsew signal input
flabel metal2 s 452544 264560 452640 264640 0 FreeSans 320 0 0 0 Tile_X10Y10_MEN_SRAM
port 1036 nsew signal output
flabel metal2 s 452544 265064 452640 265144 0 FreeSans 320 0 0 0 Tile_X10Y10_REN_SRAM
port 1037 nsew signal output
flabel metal2 s 452544 265568 452640 265648 0 FreeSans 320 0 0 0 Tile_X10Y10_TIE_HIGH_SRAM
port 1038 nsew signal output
flabel metal2 s 452544 266072 452640 266152 0 FreeSans 320 0 0 0 Tile_X10Y10_TIE_LOW_SRAM
port 1039 nsew signal output
flabel metal2 s 452544 266576 452640 266656 0 FreeSans 320 0 0 0 Tile_X10Y10_WEN_SRAM
port 1040 nsew signal output
flabel metal2 s 452544 129992 452640 130072 0 FreeSans 320 0 0 0 Tile_X10Y12_ADDR_SRAM0
port 1041 nsew signal output
flabel metal2 s 452544 130496 452640 130576 0 FreeSans 320 0 0 0 Tile_X10Y12_ADDR_SRAM1
port 1042 nsew signal output
flabel metal2 s 452544 131000 452640 131080 0 FreeSans 320 0 0 0 Tile_X10Y12_ADDR_SRAM2
port 1043 nsew signal output
flabel metal2 s 452544 131504 452640 131584 0 FreeSans 320 0 0 0 Tile_X10Y12_ADDR_SRAM3
port 1044 nsew signal output
flabel metal2 s 452544 132008 452640 132088 0 FreeSans 320 0 0 0 Tile_X10Y12_ADDR_SRAM4
port 1045 nsew signal output
flabel metal2 s 452544 132512 452640 132592 0 FreeSans 320 0 0 0 Tile_X10Y12_ADDR_SRAM5
port 1046 nsew signal output
flabel metal2 s 452544 133016 452640 133096 0 FreeSans 320 0 0 0 Tile_X10Y12_ADDR_SRAM6
port 1047 nsew signal output
flabel metal2 s 452544 133520 452640 133600 0 FreeSans 320 0 0 0 Tile_X10Y12_ADDR_SRAM7
port 1048 nsew signal output
flabel metal2 s 452544 134024 452640 134104 0 FreeSans 320 0 0 0 Tile_X10Y12_ADDR_SRAM8
port 1049 nsew signal output
flabel metal2 s 452544 134528 452640 134608 0 FreeSans 320 0 0 0 Tile_X10Y12_ADDR_SRAM9
port 1050 nsew signal output
flabel metal2 s 452544 135032 452640 135112 0 FreeSans 320 0 0 0 Tile_X10Y12_BM_SRAM0
port 1051 nsew signal output
flabel metal2 s 452544 135536 452640 135616 0 FreeSans 320 0 0 0 Tile_X10Y12_BM_SRAM1
port 1052 nsew signal output
flabel metal2 s 452544 140072 452640 140152 0 FreeSans 320 0 0 0 Tile_X10Y12_BM_SRAM10
port 1053 nsew signal output
flabel metal2 s 452544 140576 452640 140656 0 FreeSans 320 0 0 0 Tile_X10Y12_BM_SRAM11
port 1054 nsew signal output
flabel metal2 s 452544 141080 452640 141160 0 FreeSans 320 0 0 0 Tile_X10Y12_BM_SRAM12
port 1055 nsew signal output
flabel metal2 s 452544 141584 452640 141664 0 FreeSans 320 0 0 0 Tile_X10Y12_BM_SRAM13
port 1056 nsew signal output
flabel metal2 s 452544 142088 452640 142168 0 FreeSans 320 0 0 0 Tile_X10Y12_BM_SRAM14
port 1057 nsew signal output
flabel metal2 s 452544 142592 452640 142672 0 FreeSans 320 0 0 0 Tile_X10Y12_BM_SRAM15
port 1058 nsew signal output
flabel metal2 s 452544 143096 452640 143176 0 FreeSans 320 0 0 0 Tile_X10Y12_BM_SRAM16
port 1059 nsew signal output
flabel metal2 s 452544 143600 452640 143680 0 FreeSans 320 0 0 0 Tile_X10Y12_BM_SRAM17
port 1060 nsew signal output
flabel metal2 s 452544 144104 452640 144184 0 FreeSans 320 0 0 0 Tile_X10Y12_BM_SRAM18
port 1061 nsew signal output
flabel metal2 s 452544 144608 452640 144688 0 FreeSans 320 0 0 0 Tile_X10Y12_BM_SRAM19
port 1062 nsew signal output
flabel metal2 s 452544 136040 452640 136120 0 FreeSans 320 0 0 0 Tile_X10Y12_BM_SRAM2
port 1063 nsew signal output
flabel metal2 s 452544 145112 452640 145192 0 FreeSans 320 0 0 0 Tile_X10Y12_BM_SRAM20
port 1064 nsew signal output
flabel metal2 s 452544 145616 452640 145696 0 FreeSans 320 0 0 0 Tile_X10Y12_BM_SRAM21
port 1065 nsew signal output
flabel metal2 s 452544 146120 452640 146200 0 FreeSans 320 0 0 0 Tile_X10Y12_BM_SRAM22
port 1066 nsew signal output
flabel metal2 s 452544 146624 452640 146704 0 FreeSans 320 0 0 0 Tile_X10Y12_BM_SRAM23
port 1067 nsew signal output
flabel metal2 s 452544 147128 452640 147208 0 FreeSans 320 0 0 0 Tile_X10Y12_BM_SRAM24
port 1068 nsew signal output
flabel metal2 s 452544 147632 452640 147712 0 FreeSans 320 0 0 0 Tile_X10Y12_BM_SRAM25
port 1069 nsew signal output
flabel metal2 s 452544 148136 452640 148216 0 FreeSans 320 0 0 0 Tile_X10Y12_BM_SRAM26
port 1070 nsew signal output
flabel metal2 s 452544 148640 452640 148720 0 FreeSans 320 0 0 0 Tile_X10Y12_BM_SRAM27
port 1071 nsew signal output
flabel metal2 s 452544 149144 452640 149224 0 FreeSans 320 0 0 0 Tile_X10Y12_BM_SRAM28
port 1072 nsew signal output
flabel metal2 s 452544 149648 452640 149728 0 FreeSans 320 0 0 0 Tile_X10Y12_BM_SRAM29
port 1073 nsew signal output
flabel metal2 s 452544 136544 452640 136624 0 FreeSans 320 0 0 0 Tile_X10Y12_BM_SRAM3
port 1074 nsew signal output
flabel metal2 s 452544 150152 452640 150232 0 FreeSans 320 0 0 0 Tile_X10Y12_BM_SRAM30
port 1075 nsew signal output
flabel metal2 s 452544 150656 452640 150736 0 FreeSans 320 0 0 0 Tile_X10Y12_BM_SRAM31
port 1076 nsew signal output
flabel metal2 s 452544 137048 452640 137128 0 FreeSans 320 0 0 0 Tile_X10Y12_BM_SRAM4
port 1077 nsew signal output
flabel metal2 s 452544 137552 452640 137632 0 FreeSans 320 0 0 0 Tile_X10Y12_BM_SRAM5
port 1078 nsew signal output
flabel metal2 s 452544 138056 452640 138136 0 FreeSans 320 0 0 0 Tile_X10Y12_BM_SRAM6
port 1079 nsew signal output
flabel metal2 s 452544 138560 452640 138640 0 FreeSans 320 0 0 0 Tile_X10Y12_BM_SRAM7
port 1080 nsew signal output
flabel metal2 s 452544 139064 452640 139144 0 FreeSans 320 0 0 0 Tile_X10Y12_BM_SRAM8
port 1081 nsew signal output
flabel metal2 s 452544 139568 452640 139648 0 FreeSans 320 0 0 0 Tile_X10Y12_BM_SRAM9
port 1082 nsew signal output
flabel metal2 s 452544 151160 452640 151240 0 FreeSans 320 0 0 0 Tile_X10Y12_CLK_SRAM
port 1083 nsew signal output
flabel metal2 s 452544 113360 452640 113440 0 FreeSans 320 0 0 0 Tile_X10Y12_CONFIGURED_top
port 1084 nsew signal input
flabel metal2 s 452544 151664 452640 151744 0 FreeSans 320 0 0 0 Tile_X10Y12_DIN_SRAM0
port 1085 nsew signal output
flabel metal2 s 452544 152168 452640 152248 0 FreeSans 320 0 0 0 Tile_X10Y12_DIN_SRAM1
port 1086 nsew signal output
flabel metal2 s 452544 156704 452640 156784 0 FreeSans 320 0 0 0 Tile_X10Y12_DIN_SRAM10
port 1087 nsew signal output
flabel metal2 s 452544 157208 452640 157288 0 FreeSans 320 0 0 0 Tile_X10Y12_DIN_SRAM11
port 1088 nsew signal output
flabel metal2 s 452544 157712 452640 157792 0 FreeSans 320 0 0 0 Tile_X10Y12_DIN_SRAM12
port 1089 nsew signal output
flabel metal2 s 452544 158216 452640 158296 0 FreeSans 320 0 0 0 Tile_X10Y12_DIN_SRAM13
port 1090 nsew signal output
flabel metal2 s 452544 158720 452640 158800 0 FreeSans 320 0 0 0 Tile_X10Y12_DIN_SRAM14
port 1091 nsew signal output
flabel metal2 s 452544 159224 452640 159304 0 FreeSans 320 0 0 0 Tile_X10Y12_DIN_SRAM15
port 1092 nsew signal output
flabel metal2 s 452544 159728 452640 159808 0 FreeSans 320 0 0 0 Tile_X10Y12_DIN_SRAM16
port 1093 nsew signal output
flabel metal2 s 452544 160232 452640 160312 0 FreeSans 320 0 0 0 Tile_X10Y12_DIN_SRAM17
port 1094 nsew signal output
flabel metal2 s 452544 160736 452640 160816 0 FreeSans 320 0 0 0 Tile_X10Y12_DIN_SRAM18
port 1095 nsew signal output
flabel metal2 s 452544 161240 452640 161320 0 FreeSans 320 0 0 0 Tile_X10Y12_DIN_SRAM19
port 1096 nsew signal output
flabel metal2 s 452544 152672 452640 152752 0 FreeSans 320 0 0 0 Tile_X10Y12_DIN_SRAM2
port 1097 nsew signal output
flabel metal2 s 452544 161744 452640 161824 0 FreeSans 320 0 0 0 Tile_X10Y12_DIN_SRAM20
port 1098 nsew signal output
flabel metal2 s 452544 162248 452640 162328 0 FreeSans 320 0 0 0 Tile_X10Y12_DIN_SRAM21
port 1099 nsew signal output
flabel metal2 s 452544 162752 452640 162832 0 FreeSans 320 0 0 0 Tile_X10Y12_DIN_SRAM22
port 1100 nsew signal output
flabel metal2 s 452544 163256 452640 163336 0 FreeSans 320 0 0 0 Tile_X10Y12_DIN_SRAM23
port 1101 nsew signal output
flabel metal2 s 452544 163760 452640 163840 0 FreeSans 320 0 0 0 Tile_X10Y12_DIN_SRAM24
port 1102 nsew signal output
flabel metal2 s 452544 164264 452640 164344 0 FreeSans 320 0 0 0 Tile_X10Y12_DIN_SRAM25
port 1103 nsew signal output
flabel metal2 s 452544 164768 452640 164848 0 FreeSans 320 0 0 0 Tile_X10Y12_DIN_SRAM26
port 1104 nsew signal output
flabel metal2 s 452544 165272 452640 165352 0 FreeSans 320 0 0 0 Tile_X10Y12_DIN_SRAM27
port 1105 nsew signal output
flabel metal2 s 452544 165776 452640 165856 0 FreeSans 320 0 0 0 Tile_X10Y12_DIN_SRAM28
port 1106 nsew signal output
flabel metal2 s 452544 166280 452640 166360 0 FreeSans 320 0 0 0 Tile_X10Y12_DIN_SRAM29
port 1107 nsew signal output
flabel metal2 s 452544 153176 452640 153256 0 FreeSans 320 0 0 0 Tile_X10Y12_DIN_SRAM3
port 1108 nsew signal output
flabel metal2 s 452544 166784 452640 166864 0 FreeSans 320 0 0 0 Tile_X10Y12_DIN_SRAM30
port 1109 nsew signal output
flabel metal2 s 452544 167288 452640 167368 0 FreeSans 320 0 0 0 Tile_X10Y12_DIN_SRAM31
port 1110 nsew signal output
flabel metal2 s 452544 153680 452640 153760 0 FreeSans 320 0 0 0 Tile_X10Y12_DIN_SRAM4
port 1111 nsew signal output
flabel metal2 s 452544 154184 452640 154264 0 FreeSans 320 0 0 0 Tile_X10Y12_DIN_SRAM5
port 1112 nsew signal output
flabel metal2 s 452544 154688 452640 154768 0 FreeSans 320 0 0 0 Tile_X10Y12_DIN_SRAM6
port 1113 nsew signal output
flabel metal2 s 452544 155192 452640 155272 0 FreeSans 320 0 0 0 Tile_X10Y12_DIN_SRAM7
port 1114 nsew signal output
flabel metal2 s 452544 155696 452640 155776 0 FreeSans 320 0 0 0 Tile_X10Y12_DIN_SRAM8
port 1115 nsew signal output
flabel metal2 s 452544 156200 452640 156280 0 FreeSans 320 0 0 0 Tile_X10Y12_DIN_SRAM9
port 1116 nsew signal output
flabel metal2 s 452544 113864 452640 113944 0 FreeSans 320 0 0 0 Tile_X10Y12_DOUT_SRAM0
port 1117 nsew signal input
flabel metal2 s 452544 114368 452640 114448 0 FreeSans 320 0 0 0 Tile_X10Y12_DOUT_SRAM1
port 1118 nsew signal input
flabel metal2 s 452544 118904 452640 118984 0 FreeSans 320 0 0 0 Tile_X10Y12_DOUT_SRAM10
port 1119 nsew signal input
flabel metal2 s 452544 119408 452640 119488 0 FreeSans 320 0 0 0 Tile_X10Y12_DOUT_SRAM11
port 1120 nsew signal input
flabel metal2 s 452544 119912 452640 119992 0 FreeSans 320 0 0 0 Tile_X10Y12_DOUT_SRAM12
port 1121 nsew signal input
flabel metal2 s 452544 120416 452640 120496 0 FreeSans 320 0 0 0 Tile_X10Y12_DOUT_SRAM13
port 1122 nsew signal input
flabel metal2 s 452544 120920 452640 121000 0 FreeSans 320 0 0 0 Tile_X10Y12_DOUT_SRAM14
port 1123 nsew signal input
flabel metal2 s 452544 121424 452640 121504 0 FreeSans 320 0 0 0 Tile_X10Y12_DOUT_SRAM15
port 1124 nsew signal input
flabel metal2 s 452544 121928 452640 122008 0 FreeSans 320 0 0 0 Tile_X10Y12_DOUT_SRAM16
port 1125 nsew signal input
flabel metal2 s 452544 122432 452640 122512 0 FreeSans 320 0 0 0 Tile_X10Y12_DOUT_SRAM17
port 1126 nsew signal input
flabel metal2 s 452544 122936 452640 123016 0 FreeSans 320 0 0 0 Tile_X10Y12_DOUT_SRAM18
port 1127 nsew signal input
flabel metal2 s 452544 123440 452640 123520 0 FreeSans 320 0 0 0 Tile_X10Y12_DOUT_SRAM19
port 1128 nsew signal input
flabel metal2 s 452544 114872 452640 114952 0 FreeSans 320 0 0 0 Tile_X10Y12_DOUT_SRAM2
port 1129 nsew signal input
flabel metal2 s 452544 123944 452640 124024 0 FreeSans 320 0 0 0 Tile_X10Y12_DOUT_SRAM20
port 1130 nsew signal input
flabel metal2 s 452544 124448 452640 124528 0 FreeSans 320 0 0 0 Tile_X10Y12_DOUT_SRAM21
port 1131 nsew signal input
flabel metal2 s 452544 124952 452640 125032 0 FreeSans 320 0 0 0 Tile_X10Y12_DOUT_SRAM22
port 1132 nsew signal input
flabel metal2 s 452544 125456 452640 125536 0 FreeSans 320 0 0 0 Tile_X10Y12_DOUT_SRAM23
port 1133 nsew signal input
flabel metal2 s 452544 125960 452640 126040 0 FreeSans 320 0 0 0 Tile_X10Y12_DOUT_SRAM24
port 1134 nsew signal input
flabel metal2 s 452544 126464 452640 126544 0 FreeSans 320 0 0 0 Tile_X10Y12_DOUT_SRAM25
port 1135 nsew signal input
flabel metal2 s 452544 126968 452640 127048 0 FreeSans 320 0 0 0 Tile_X10Y12_DOUT_SRAM26
port 1136 nsew signal input
flabel metal2 s 452544 127472 452640 127552 0 FreeSans 320 0 0 0 Tile_X10Y12_DOUT_SRAM27
port 1137 nsew signal input
flabel metal2 s 452544 127976 452640 128056 0 FreeSans 320 0 0 0 Tile_X10Y12_DOUT_SRAM28
port 1138 nsew signal input
flabel metal2 s 452544 128480 452640 128560 0 FreeSans 320 0 0 0 Tile_X10Y12_DOUT_SRAM29
port 1139 nsew signal input
flabel metal2 s 452544 115376 452640 115456 0 FreeSans 320 0 0 0 Tile_X10Y12_DOUT_SRAM3
port 1140 nsew signal input
flabel metal2 s 452544 128984 452640 129064 0 FreeSans 320 0 0 0 Tile_X10Y12_DOUT_SRAM30
port 1141 nsew signal input
flabel metal2 s 452544 129488 452640 129568 0 FreeSans 320 0 0 0 Tile_X10Y12_DOUT_SRAM31
port 1142 nsew signal input
flabel metal2 s 452544 115880 452640 115960 0 FreeSans 320 0 0 0 Tile_X10Y12_DOUT_SRAM4
port 1143 nsew signal input
flabel metal2 s 452544 116384 452640 116464 0 FreeSans 320 0 0 0 Tile_X10Y12_DOUT_SRAM5
port 1144 nsew signal input
flabel metal2 s 452544 116888 452640 116968 0 FreeSans 320 0 0 0 Tile_X10Y12_DOUT_SRAM6
port 1145 nsew signal input
flabel metal2 s 452544 117392 452640 117472 0 FreeSans 320 0 0 0 Tile_X10Y12_DOUT_SRAM7
port 1146 nsew signal input
flabel metal2 s 452544 117896 452640 117976 0 FreeSans 320 0 0 0 Tile_X10Y12_DOUT_SRAM8
port 1147 nsew signal input
flabel metal2 s 452544 118400 452640 118480 0 FreeSans 320 0 0 0 Tile_X10Y12_DOUT_SRAM9
port 1148 nsew signal input
flabel metal2 s 452544 167792 452640 167872 0 FreeSans 320 0 0 0 Tile_X10Y12_MEN_SRAM
port 1149 nsew signal output
flabel metal2 s 452544 168296 452640 168376 0 FreeSans 320 0 0 0 Tile_X10Y12_REN_SRAM
port 1150 nsew signal output
flabel metal2 s 452544 168800 452640 168880 0 FreeSans 320 0 0 0 Tile_X10Y12_TIE_HIGH_SRAM
port 1151 nsew signal output
flabel metal2 s 452544 169304 452640 169384 0 FreeSans 320 0 0 0 Tile_X10Y12_TIE_LOW_SRAM
port 1152 nsew signal output
flabel metal2 s 452544 169808 452640 169888 0 FreeSans 320 0 0 0 Tile_X10Y12_WEN_SRAM
port 1153 nsew signal output
flabel metal2 s 452544 33224 452640 33304 0 FreeSans 320 0 0 0 Tile_X10Y14_ADDR_SRAM0
port 1154 nsew signal output
flabel metal2 s 452544 33728 452640 33808 0 FreeSans 320 0 0 0 Tile_X10Y14_ADDR_SRAM1
port 1155 nsew signal output
flabel metal2 s 452544 34232 452640 34312 0 FreeSans 320 0 0 0 Tile_X10Y14_ADDR_SRAM2
port 1156 nsew signal output
flabel metal2 s 452544 34736 452640 34816 0 FreeSans 320 0 0 0 Tile_X10Y14_ADDR_SRAM3
port 1157 nsew signal output
flabel metal2 s 452544 35240 452640 35320 0 FreeSans 320 0 0 0 Tile_X10Y14_ADDR_SRAM4
port 1158 nsew signal output
flabel metal2 s 452544 35744 452640 35824 0 FreeSans 320 0 0 0 Tile_X10Y14_ADDR_SRAM5
port 1159 nsew signal output
flabel metal2 s 452544 36248 452640 36328 0 FreeSans 320 0 0 0 Tile_X10Y14_ADDR_SRAM6
port 1160 nsew signal output
flabel metal2 s 452544 36752 452640 36832 0 FreeSans 320 0 0 0 Tile_X10Y14_ADDR_SRAM7
port 1161 nsew signal output
flabel metal2 s 452544 37256 452640 37336 0 FreeSans 320 0 0 0 Tile_X10Y14_ADDR_SRAM8
port 1162 nsew signal output
flabel metal2 s 452544 37760 452640 37840 0 FreeSans 320 0 0 0 Tile_X10Y14_ADDR_SRAM9
port 1163 nsew signal output
flabel metal2 s 452544 38264 452640 38344 0 FreeSans 320 0 0 0 Tile_X10Y14_BM_SRAM0
port 1164 nsew signal output
flabel metal2 s 452544 38768 452640 38848 0 FreeSans 320 0 0 0 Tile_X10Y14_BM_SRAM1
port 1165 nsew signal output
flabel metal2 s 452544 43304 452640 43384 0 FreeSans 320 0 0 0 Tile_X10Y14_BM_SRAM10
port 1166 nsew signal output
flabel metal2 s 452544 43808 452640 43888 0 FreeSans 320 0 0 0 Tile_X10Y14_BM_SRAM11
port 1167 nsew signal output
flabel metal2 s 452544 44312 452640 44392 0 FreeSans 320 0 0 0 Tile_X10Y14_BM_SRAM12
port 1168 nsew signal output
flabel metal2 s 452544 44816 452640 44896 0 FreeSans 320 0 0 0 Tile_X10Y14_BM_SRAM13
port 1169 nsew signal output
flabel metal2 s 452544 45320 452640 45400 0 FreeSans 320 0 0 0 Tile_X10Y14_BM_SRAM14
port 1170 nsew signal output
flabel metal2 s 452544 45824 452640 45904 0 FreeSans 320 0 0 0 Tile_X10Y14_BM_SRAM15
port 1171 nsew signal output
flabel metal2 s 452544 46328 452640 46408 0 FreeSans 320 0 0 0 Tile_X10Y14_BM_SRAM16
port 1172 nsew signal output
flabel metal2 s 452544 46832 452640 46912 0 FreeSans 320 0 0 0 Tile_X10Y14_BM_SRAM17
port 1173 nsew signal output
flabel metal2 s 452544 47336 452640 47416 0 FreeSans 320 0 0 0 Tile_X10Y14_BM_SRAM18
port 1174 nsew signal output
flabel metal2 s 452544 47840 452640 47920 0 FreeSans 320 0 0 0 Tile_X10Y14_BM_SRAM19
port 1175 nsew signal output
flabel metal2 s 452544 39272 452640 39352 0 FreeSans 320 0 0 0 Tile_X10Y14_BM_SRAM2
port 1176 nsew signal output
flabel metal2 s 452544 48344 452640 48424 0 FreeSans 320 0 0 0 Tile_X10Y14_BM_SRAM20
port 1177 nsew signal output
flabel metal2 s 452544 48848 452640 48928 0 FreeSans 320 0 0 0 Tile_X10Y14_BM_SRAM21
port 1178 nsew signal output
flabel metal2 s 452544 49352 452640 49432 0 FreeSans 320 0 0 0 Tile_X10Y14_BM_SRAM22
port 1179 nsew signal output
flabel metal2 s 452544 49856 452640 49936 0 FreeSans 320 0 0 0 Tile_X10Y14_BM_SRAM23
port 1180 nsew signal output
flabel metal2 s 452544 50360 452640 50440 0 FreeSans 320 0 0 0 Tile_X10Y14_BM_SRAM24
port 1181 nsew signal output
flabel metal2 s 452544 50864 452640 50944 0 FreeSans 320 0 0 0 Tile_X10Y14_BM_SRAM25
port 1182 nsew signal output
flabel metal2 s 452544 51368 452640 51448 0 FreeSans 320 0 0 0 Tile_X10Y14_BM_SRAM26
port 1183 nsew signal output
flabel metal2 s 452544 51872 452640 51952 0 FreeSans 320 0 0 0 Tile_X10Y14_BM_SRAM27
port 1184 nsew signal output
flabel metal2 s 452544 52376 452640 52456 0 FreeSans 320 0 0 0 Tile_X10Y14_BM_SRAM28
port 1185 nsew signal output
flabel metal2 s 452544 52880 452640 52960 0 FreeSans 320 0 0 0 Tile_X10Y14_BM_SRAM29
port 1186 nsew signal output
flabel metal2 s 452544 39776 452640 39856 0 FreeSans 320 0 0 0 Tile_X10Y14_BM_SRAM3
port 1187 nsew signal output
flabel metal2 s 452544 53384 452640 53464 0 FreeSans 320 0 0 0 Tile_X10Y14_BM_SRAM30
port 1188 nsew signal output
flabel metal2 s 452544 53888 452640 53968 0 FreeSans 320 0 0 0 Tile_X10Y14_BM_SRAM31
port 1189 nsew signal output
flabel metal2 s 452544 40280 452640 40360 0 FreeSans 320 0 0 0 Tile_X10Y14_BM_SRAM4
port 1190 nsew signal output
flabel metal2 s 452544 40784 452640 40864 0 FreeSans 320 0 0 0 Tile_X10Y14_BM_SRAM5
port 1191 nsew signal output
flabel metal2 s 452544 41288 452640 41368 0 FreeSans 320 0 0 0 Tile_X10Y14_BM_SRAM6
port 1192 nsew signal output
flabel metal2 s 452544 41792 452640 41872 0 FreeSans 320 0 0 0 Tile_X10Y14_BM_SRAM7
port 1193 nsew signal output
flabel metal2 s 452544 42296 452640 42376 0 FreeSans 320 0 0 0 Tile_X10Y14_BM_SRAM8
port 1194 nsew signal output
flabel metal2 s 452544 42800 452640 42880 0 FreeSans 320 0 0 0 Tile_X10Y14_BM_SRAM9
port 1195 nsew signal output
flabel metal2 s 452544 54392 452640 54472 0 FreeSans 320 0 0 0 Tile_X10Y14_CLK_SRAM
port 1196 nsew signal output
flabel metal2 s 452544 16592 452640 16672 0 FreeSans 320 0 0 0 Tile_X10Y14_CONFIGURED_top
port 1197 nsew signal input
flabel metal2 s 452544 54896 452640 54976 0 FreeSans 320 0 0 0 Tile_X10Y14_DIN_SRAM0
port 1198 nsew signal output
flabel metal2 s 452544 55400 452640 55480 0 FreeSans 320 0 0 0 Tile_X10Y14_DIN_SRAM1
port 1199 nsew signal output
flabel metal2 s 452544 59936 452640 60016 0 FreeSans 320 0 0 0 Tile_X10Y14_DIN_SRAM10
port 1200 nsew signal output
flabel metal2 s 452544 60440 452640 60520 0 FreeSans 320 0 0 0 Tile_X10Y14_DIN_SRAM11
port 1201 nsew signal output
flabel metal2 s 452544 60944 452640 61024 0 FreeSans 320 0 0 0 Tile_X10Y14_DIN_SRAM12
port 1202 nsew signal output
flabel metal2 s 452544 61448 452640 61528 0 FreeSans 320 0 0 0 Tile_X10Y14_DIN_SRAM13
port 1203 nsew signal output
flabel metal2 s 452544 61952 452640 62032 0 FreeSans 320 0 0 0 Tile_X10Y14_DIN_SRAM14
port 1204 nsew signal output
flabel metal2 s 452544 62456 452640 62536 0 FreeSans 320 0 0 0 Tile_X10Y14_DIN_SRAM15
port 1205 nsew signal output
flabel metal2 s 452544 62960 452640 63040 0 FreeSans 320 0 0 0 Tile_X10Y14_DIN_SRAM16
port 1206 nsew signal output
flabel metal2 s 452544 63464 452640 63544 0 FreeSans 320 0 0 0 Tile_X10Y14_DIN_SRAM17
port 1207 nsew signal output
flabel metal2 s 452544 63968 452640 64048 0 FreeSans 320 0 0 0 Tile_X10Y14_DIN_SRAM18
port 1208 nsew signal output
flabel metal2 s 452544 64472 452640 64552 0 FreeSans 320 0 0 0 Tile_X10Y14_DIN_SRAM19
port 1209 nsew signal output
flabel metal2 s 452544 55904 452640 55984 0 FreeSans 320 0 0 0 Tile_X10Y14_DIN_SRAM2
port 1210 nsew signal output
flabel metal2 s 452544 64976 452640 65056 0 FreeSans 320 0 0 0 Tile_X10Y14_DIN_SRAM20
port 1211 nsew signal output
flabel metal2 s 452544 65480 452640 65560 0 FreeSans 320 0 0 0 Tile_X10Y14_DIN_SRAM21
port 1212 nsew signal output
flabel metal2 s 452544 65984 452640 66064 0 FreeSans 320 0 0 0 Tile_X10Y14_DIN_SRAM22
port 1213 nsew signal output
flabel metal2 s 452544 66488 452640 66568 0 FreeSans 320 0 0 0 Tile_X10Y14_DIN_SRAM23
port 1214 nsew signal output
flabel metal2 s 452544 66992 452640 67072 0 FreeSans 320 0 0 0 Tile_X10Y14_DIN_SRAM24
port 1215 nsew signal output
flabel metal2 s 452544 67496 452640 67576 0 FreeSans 320 0 0 0 Tile_X10Y14_DIN_SRAM25
port 1216 nsew signal output
flabel metal2 s 452544 68000 452640 68080 0 FreeSans 320 0 0 0 Tile_X10Y14_DIN_SRAM26
port 1217 nsew signal output
flabel metal2 s 452544 68504 452640 68584 0 FreeSans 320 0 0 0 Tile_X10Y14_DIN_SRAM27
port 1218 nsew signal output
flabel metal2 s 452544 69008 452640 69088 0 FreeSans 320 0 0 0 Tile_X10Y14_DIN_SRAM28
port 1219 nsew signal output
flabel metal2 s 452544 69512 452640 69592 0 FreeSans 320 0 0 0 Tile_X10Y14_DIN_SRAM29
port 1220 nsew signal output
flabel metal2 s 452544 56408 452640 56488 0 FreeSans 320 0 0 0 Tile_X10Y14_DIN_SRAM3
port 1221 nsew signal output
flabel metal2 s 452544 70016 452640 70096 0 FreeSans 320 0 0 0 Tile_X10Y14_DIN_SRAM30
port 1222 nsew signal output
flabel metal2 s 452544 70520 452640 70600 0 FreeSans 320 0 0 0 Tile_X10Y14_DIN_SRAM31
port 1223 nsew signal output
flabel metal2 s 452544 56912 452640 56992 0 FreeSans 320 0 0 0 Tile_X10Y14_DIN_SRAM4
port 1224 nsew signal output
flabel metal2 s 452544 57416 452640 57496 0 FreeSans 320 0 0 0 Tile_X10Y14_DIN_SRAM5
port 1225 nsew signal output
flabel metal2 s 452544 57920 452640 58000 0 FreeSans 320 0 0 0 Tile_X10Y14_DIN_SRAM6
port 1226 nsew signal output
flabel metal2 s 452544 58424 452640 58504 0 FreeSans 320 0 0 0 Tile_X10Y14_DIN_SRAM7
port 1227 nsew signal output
flabel metal2 s 452544 58928 452640 59008 0 FreeSans 320 0 0 0 Tile_X10Y14_DIN_SRAM8
port 1228 nsew signal output
flabel metal2 s 452544 59432 452640 59512 0 FreeSans 320 0 0 0 Tile_X10Y14_DIN_SRAM9
port 1229 nsew signal output
flabel metal2 s 452544 17096 452640 17176 0 FreeSans 320 0 0 0 Tile_X10Y14_DOUT_SRAM0
port 1230 nsew signal input
flabel metal2 s 452544 17600 452640 17680 0 FreeSans 320 0 0 0 Tile_X10Y14_DOUT_SRAM1
port 1231 nsew signal input
flabel metal2 s 452544 22136 452640 22216 0 FreeSans 320 0 0 0 Tile_X10Y14_DOUT_SRAM10
port 1232 nsew signal input
flabel metal2 s 452544 22640 452640 22720 0 FreeSans 320 0 0 0 Tile_X10Y14_DOUT_SRAM11
port 1233 nsew signal input
flabel metal2 s 452544 23144 452640 23224 0 FreeSans 320 0 0 0 Tile_X10Y14_DOUT_SRAM12
port 1234 nsew signal input
flabel metal2 s 452544 23648 452640 23728 0 FreeSans 320 0 0 0 Tile_X10Y14_DOUT_SRAM13
port 1235 nsew signal input
flabel metal2 s 452544 24152 452640 24232 0 FreeSans 320 0 0 0 Tile_X10Y14_DOUT_SRAM14
port 1236 nsew signal input
flabel metal2 s 452544 24656 452640 24736 0 FreeSans 320 0 0 0 Tile_X10Y14_DOUT_SRAM15
port 1237 nsew signal input
flabel metal2 s 452544 25160 452640 25240 0 FreeSans 320 0 0 0 Tile_X10Y14_DOUT_SRAM16
port 1238 nsew signal input
flabel metal2 s 452544 25664 452640 25744 0 FreeSans 320 0 0 0 Tile_X10Y14_DOUT_SRAM17
port 1239 nsew signal input
flabel metal2 s 452544 26168 452640 26248 0 FreeSans 320 0 0 0 Tile_X10Y14_DOUT_SRAM18
port 1240 nsew signal input
flabel metal2 s 452544 26672 452640 26752 0 FreeSans 320 0 0 0 Tile_X10Y14_DOUT_SRAM19
port 1241 nsew signal input
flabel metal2 s 452544 18104 452640 18184 0 FreeSans 320 0 0 0 Tile_X10Y14_DOUT_SRAM2
port 1242 nsew signal input
flabel metal2 s 452544 27176 452640 27256 0 FreeSans 320 0 0 0 Tile_X10Y14_DOUT_SRAM20
port 1243 nsew signal input
flabel metal2 s 452544 27680 452640 27760 0 FreeSans 320 0 0 0 Tile_X10Y14_DOUT_SRAM21
port 1244 nsew signal input
flabel metal2 s 452544 28184 452640 28264 0 FreeSans 320 0 0 0 Tile_X10Y14_DOUT_SRAM22
port 1245 nsew signal input
flabel metal2 s 452544 28688 452640 28768 0 FreeSans 320 0 0 0 Tile_X10Y14_DOUT_SRAM23
port 1246 nsew signal input
flabel metal2 s 452544 29192 452640 29272 0 FreeSans 320 0 0 0 Tile_X10Y14_DOUT_SRAM24
port 1247 nsew signal input
flabel metal2 s 452544 29696 452640 29776 0 FreeSans 320 0 0 0 Tile_X10Y14_DOUT_SRAM25
port 1248 nsew signal input
flabel metal2 s 452544 30200 452640 30280 0 FreeSans 320 0 0 0 Tile_X10Y14_DOUT_SRAM26
port 1249 nsew signal input
flabel metal2 s 452544 30704 452640 30784 0 FreeSans 320 0 0 0 Tile_X10Y14_DOUT_SRAM27
port 1250 nsew signal input
flabel metal2 s 452544 31208 452640 31288 0 FreeSans 320 0 0 0 Tile_X10Y14_DOUT_SRAM28
port 1251 nsew signal input
flabel metal2 s 452544 31712 452640 31792 0 FreeSans 320 0 0 0 Tile_X10Y14_DOUT_SRAM29
port 1252 nsew signal input
flabel metal2 s 452544 18608 452640 18688 0 FreeSans 320 0 0 0 Tile_X10Y14_DOUT_SRAM3
port 1253 nsew signal input
flabel metal2 s 452544 32216 452640 32296 0 FreeSans 320 0 0 0 Tile_X10Y14_DOUT_SRAM30
port 1254 nsew signal input
flabel metal2 s 452544 32720 452640 32800 0 FreeSans 320 0 0 0 Tile_X10Y14_DOUT_SRAM31
port 1255 nsew signal input
flabel metal2 s 452544 19112 452640 19192 0 FreeSans 320 0 0 0 Tile_X10Y14_DOUT_SRAM4
port 1256 nsew signal input
flabel metal2 s 452544 19616 452640 19696 0 FreeSans 320 0 0 0 Tile_X10Y14_DOUT_SRAM5
port 1257 nsew signal input
flabel metal2 s 452544 20120 452640 20200 0 FreeSans 320 0 0 0 Tile_X10Y14_DOUT_SRAM6
port 1258 nsew signal input
flabel metal2 s 452544 20624 452640 20704 0 FreeSans 320 0 0 0 Tile_X10Y14_DOUT_SRAM7
port 1259 nsew signal input
flabel metal2 s 452544 21128 452640 21208 0 FreeSans 320 0 0 0 Tile_X10Y14_DOUT_SRAM8
port 1260 nsew signal input
flabel metal2 s 452544 21632 452640 21712 0 FreeSans 320 0 0 0 Tile_X10Y14_DOUT_SRAM9
port 1261 nsew signal input
flabel metal2 s 452544 71024 452640 71104 0 FreeSans 320 0 0 0 Tile_X10Y14_MEN_SRAM
port 1262 nsew signal output
flabel metal2 s 452544 71528 452640 71608 0 FreeSans 320 0 0 0 Tile_X10Y14_REN_SRAM
port 1263 nsew signal output
flabel metal2 s 452544 72032 452640 72112 0 FreeSans 320 0 0 0 Tile_X10Y14_TIE_HIGH_SRAM
port 1264 nsew signal output
flabel metal2 s 452544 72536 452640 72616 0 FreeSans 320 0 0 0 Tile_X10Y14_TIE_LOW_SRAM
port 1265 nsew signal output
flabel metal2 s 452544 73040 452640 73120 0 FreeSans 320 0 0 0 Tile_X10Y14_WEN_SRAM
port 1266 nsew signal output
flabel metal2 s 452544 613832 452640 613912 0 FreeSans 320 0 0 0 Tile_X10Y2_ADDR_SRAM0
port 1267 nsew signal output
flabel metal2 s 452544 614336 452640 614416 0 FreeSans 320 0 0 0 Tile_X10Y2_ADDR_SRAM1
port 1268 nsew signal output
flabel metal2 s 452544 614840 452640 614920 0 FreeSans 320 0 0 0 Tile_X10Y2_ADDR_SRAM2
port 1269 nsew signal output
flabel metal2 s 452544 615344 452640 615424 0 FreeSans 320 0 0 0 Tile_X10Y2_ADDR_SRAM3
port 1270 nsew signal output
flabel metal2 s 452544 615848 452640 615928 0 FreeSans 320 0 0 0 Tile_X10Y2_ADDR_SRAM4
port 1271 nsew signal output
flabel metal2 s 452544 616352 452640 616432 0 FreeSans 320 0 0 0 Tile_X10Y2_ADDR_SRAM5
port 1272 nsew signal output
flabel metal2 s 452544 616856 452640 616936 0 FreeSans 320 0 0 0 Tile_X10Y2_ADDR_SRAM6
port 1273 nsew signal output
flabel metal2 s 452544 617360 452640 617440 0 FreeSans 320 0 0 0 Tile_X10Y2_ADDR_SRAM7
port 1274 nsew signal output
flabel metal2 s 452544 617864 452640 617944 0 FreeSans 320 0 0 0 Tile_X10Y2_ADDR_SRAM8
port 1275 nsew signal output
flabel metal2 s 452544 618368 452640 618448 0 FreeSans 320 0 0 0 Tile_X10Y2_ADDR_SRAM9
port 1276 nsew signal output
flabel metal2 s 452544 618872 452640 618952 0 FreeSans 320 0 0 0 Tile_X10Y2_BM_SRAM0
port 1277 nsew signal output
flabel metal2 s 452544 619376 452640 619456 0 FreeSans 320 0 0 0 Tile_X10Y2_BM_SRAM1
port 1278 nsew signal output
flabel metal2 s 452544 623912 452640 623992 0 FreeSans 320 0 0 0 Tile_X10Y2_BM_SRAM10
port 1279 nsew signal output
flabel metal2 s 452544 624416 452640 624496 0 FreeSans 320 0 0 0 Tile_X10Y2_BM_SRAM11
port 1280 nsew signal output
flabel metal2 s 452544 624920 452640 625000 0 FreeSans 320 0 0 0 Tile_X10Y2_BM_SRAM12
port 1281 nsew signal output
flabel metal2 s 452544 625424 452640 625504 0 FreeSans 320 0 0 0 Tile_X10Y2_BM_SRAM13
port 1282 nsew signal output
flabel metal2 s 452544 625928 452640 626008 0 FreeSans 320 0 0 0 Tile_X10Y2_BM_SRAM14
port 1283 nsew signal output
flabel metal2 s 452544 626432 452640 626512 0 FreeSans 320 0 0 0 Tile_X10Y2_BM_SRAM15
port 1284 nsew signal output
flabel metal2 s 452544 626936 452640 627016 0 FreeSans 320 0 0 0 Tile_X10Y2_BM_SRAM16
port 1285 nsew signal output
flabel metal2 s 452544 627440 452640 627520 0 FreeSans 320 0 0 0 Tile_X10Y2_BM_SRAM17
port 1286 nsew signal output
flabel metal2 s 452544 627944 452640 628024 0 FreeSans 320 0 0 0 Tile_X10Y2_BM_SRAM18
port 1287 nsew signal output
flabel metal2 s 452544 628448 452640 628528 0 FreeSans 320 0 0 0 Tile_X10Y2_BM_SRAM19
port 1288 nsew signal output
flabel metal2 s 452544 619880 452640 619960 0 FreeSans 320 0 0 0 Tile_X10Y2_BM_SRAM2
port 1289 nsew signal output
flabel metal2 s 452544 628952 452640 629032 0 FreeSans 320 0 0 0 Tile_X10Y2_BM_SRAM20
port 1290 nsew signal output
flabel metal2 s 452544 629456 452640 629536 0 FreeSans 320 0 0 0 Tile_X10Y2_BM_SRAM21
port 1291 nsew signal output
flabel metal2 s 452544 629960 452640 630040 0 FreeSans 320 0 0 0 Tile_X10Y2_BM_SRAM22
port 1292 nsew signal output
flabel metal2 s 452544 630464 452640 630544 0 FreeSans 320 0 0 0 Tile_X10Y2_BM_SRAM23
port 1293 nsew signal output
flabel metal2 s 452544 630968 452640 631048 0 FreeSans 320 0 0 0 Tile_X10Y2_BM_SRAM24
port 1294 nsew signal output
flabel metal2 s 452544 631472 452640 631552 0 FreeSans 320 0 0 0 Tile_X10Y2_BM_SRAM25
port 1295 nsew signal output
flabel metal2 s 452544 631976 452640 632056 0 FreeSans 320 0 0 0 Tile_X10Y2_BM_SRAM26
port 1296 nsew signal output
flabel metal2 s 452544 632480 452640 632560 0 FreeSans 320 0 0 0 Tile_X10Y2_BM_SRAM27
port 1297 nsew signal output
flabel metal2 s 452544 632984 452640 633064 0 FreeSans 320 0 0 0 Tile_X10Y2_BM_SRAM28
port 1298 nsew signal output
flabel metal2 s 452544 633488 452640 633568 0 FreeSans 320 0 0 0 Tile_X10Y2_BM_SRAM29
port 1299 nsew signal output
flabel metal2 s 452544 620384 452640 620464 0 FreeSans 320 0 0 0 Tile_X10Y2_BM_SRAM3
port 1300 nsew signal output
flabel metal2 s 452544 633992 452640 634072 0 FreeSans 320 0 0 0 Tile_X10Y2_BM_SRAM30
port 1301 nsew signal output
flabel metal2 s 452544 634496 452640 634576 0 FreeSans 320 0 0 0 Tile_X10Y2_BM_SRAM31
port 1302 nsew signal output
flabel metal2 s 452544 620888 452640 620968 0 FreeSans 320 0 0 0 Tile_X10Y2_BM_SRAM4
port 1303 nsew signal output
flabel metal2 s 452544 621392 452640 621472 0 FreeSans 320 0 0 0 Tile_X10Y2_BM_SRAM5
port 1304 nsew signal output
flabel metal2 s 452544 621896 452640 621976 0 FreeSans 320 0 0 0 Tile_X10Y2_BM_SRAM6
port 1305 nsew signal output
flabel metal2 s 452544 622400 452640 622480 0 FreeSans 320 0 0 0 Tile_X10Y2_BM_SRAM7
port 1306 nsew signal output
flabel metal2 s 452544 622904 452640 622984 0 FreeSans 320 0 0 0 Tile_X10Y2_BM_SRAM8
port 1307 nsew signal output
flabel metal2 s 452544 623408 452640 623488 0 FreeSans 320 0 0 0 Tile_X10Y2_BM_SRAM9
port 1308 nsew signal output
flabel metal2 s 452544 635000 452640 635080 0 FreeSans 320 0 0 0 Tile_X10Y2_CLK_SRAM
port 1309 nsew signal output
flabel metal2 s 452544 597200 452640 597280 0 FreeSans 320 0 0 0 Tile_X10Y2_CONFIGURED_top
port 1310 nsew signal input
flabel metal2 s 452544 635504 452640 635584 0 FreeSans 320 0 0 0 Tile_X10Y2_DIN_SRAM0
port 1311 nsew signal output
flabel metal2 s 452544 636008 452640 636088 0 FreeSans 320 0 0 0 Tile_X10Y2_DIN_SRAM1
port 1312 nsew signal output
flabel metal2 s 452544 640544 452640 640624 0 FreeSans 320 0 0 0 Tile_X10Y2_DIN_SRAM10
port 1313 nsew signal output
flabel metal2 s 452544 641048 452640 641128 0 FreeSans 320 0 0 0 Tile_X10Y2_DIN_SRAM11
port 1314 nsew signal output
flabel metal2 s 452544 641552 452640 641632 0 FreeSans 320 0 0 0 Tile_X10Y2_DIN_SRAM12
port 1315 nsew signal output
flabel metal2 s 452544 642056 452640 642136 0 FreeSans 320 0 0 0 Tile_X10Y2_DIN_SRAM13
port 1316 nsew signal output
flabel metal2 s 452544 642560 452640 642640 0 FreeSans 320 0 0 0 Tile_X10Y2_DIN_SRAM14
port 1317 nsew signal output
flabel metal2 s 452544 643064 452640 643144 0 FreeSans 320 0 0 0 Tile_X10Y2_DIN_SRAM15
port 1318 nsew signal output
flabel metal2 s 452544 643568 452640 643648 0 FreeSans 320 0 0 0 Tile_X10Y2_DIN_SRAM16
port 1319 nsew signal output
flabel metal2 s 452544 644072 452640 644152 0 FreeSans 320 0 0 0 Tile_X10Y2_DIN_SRAM17
port 1320 nsew signal output
flabel metal2 s 452544 644576 452640 644656 0 FreeSans 320 0 0 0 Tile_X10Y2_DIN_SRAM18
port 1321 nsew signal output
flabel metal2 s 452544 645080 452640 645160 0 FreeSans 320 0 0 0 Tile_X10Y2_DIN_SRAM19
port 1322 nsew signal output
flabel metal2 s 452544 636512 452640 636592 0 FreeSans 320 0 0 0 Tile_X10Y2_DIN_SRAM2
port 1323 nsew signal output
flabel metal2 s 452544 645584 452640 645664 0 FreeSans 320 0 0 0 Tile_X10Y2_DIN_SRAM20
port 1324 nsew signal output
flabel metal2 s 452544 646088 452640 646168 0 FreeSans 320 0 0 0 Tile_X10Y2_DIN_SRAM21
port 1325 nsew signal output
flabel metal2 s 452544 646592 452640 646672 0 FreeSans 320 0 0 0 Tile_X10Y2_DIN_SRAM22
port 1326 nsew signal output
flabel metal2 s 452544 647096 452640 647176 0 FreeSans 320 0 0 0 Tile_X10Y2_DIN_SRAM23
port 1327 nsew signal output
flabel metal2 s 452544 647600 452640 647680 0 FreeSans 320 0 0 0 Tile_X10Y2_DIN_SRAM24
port 1328 nsew signal output
flabel metal2 s 452544 648104 452640 648184 0 FreeSans 320 0 0 0 Tile_X10Y2_DIN_SRAM25
port 1329 nsew signal output
flabel metal2 s 452544 648608 452640 648688 0 FreeSans 320 0 0 0 Tile_X10Y2_DIN_SRAM26
port 1330 nsew signal output
flabel metal2 s 452544 649112 452640 649192 0 FreeSans 320 0 0 0 Tile_X10Y2_DIN_SRAM27
port 1331 nsew signal output
flabel metal2 s 452544 649616 452640 649696 0 FreeSans 320 0 0 0 Tile_X10Y2_DIN_SRAM28
port 1332 nsew signal output
flabel metal2 s 452544 650120 452640 650200 0 FreeSans 320 0 0 0 Tile_X10Y2_DIN_SRAM29
port 1333 nsew signal output
flabel metal2 s 452544 637016 452640 637096 0 FreeSans 320 0 0 0 Tile_X10Y2_DIN_SRAM3
port 1334 nsew signal output
flabel metal2 s 452544 650624 452640 650704 0 FreeSans 320 0 0 0 Tile_X10Y2_DIN_SRAM30
port 1335 nsew signal output
flabel metal2 s 452544 651128 452640 651208 0 FreeSans 320 0 0 0 Tile_X10Y2_DIN_SRAM31
port 1336 nsew signal output
flabel metal2 s 452544 637520 452640 637600 0 FreeSans 320 0 0 0 Tile_X10Y2_DIN_SRAM4
port 1337 nsew signal output
flabel metal2 s 452544 638024 452640 638104 0 FreeSans 320 0 0 0 Tile_X10Y2_DIN_SRAM5
port 1338 nsew signal output
flabel metal2 s 452544 638528 452640 638608 0 FreeSans 320 0 0 0 Tile_X10Y2_DIN_SRAM6
port 1339 nsew signal output
flabel metal2 s 452544 639032 452640 639112 0 FreeSans 320 0 0 0 Tile_X10Y2_DIN_SRAM7
port 1340 nsew signal output
flabel metal2 s 452544 639536 452640 639616 0 FreeSans 320 0 0 0 Tile_X10Y2_DIN_SRAM8
port 1341 nsew signal output
flabel metal2 s 452544 640040 452640 640120 0 FreeSans 320 0 0 0 Tile_X10Y2_DIN_SRAM9
port 1342 nsew signal output
flabel metal2 s 452544 597704 452640 597784 0 FreeSans 320 0 0 0 Tile_X10Y2_DOUT_SRAM0
port 1343 nsew signal input
flabel metal2 s 452544 598208 452640 598288 0 FreeSans 320 0 0 0 Tile_X10Y2_DOUT_SRAM1
port 1344 nsew signal input
flabel metal2 s 452544 602744 452640 602824 0 FreeSans 320 0 0 0 Tile_X10Y2_DOUT_SRAM10
port 1345 nsew signal input
flabel metal2 s 452544 603248 452640 603328 0 FreeSans 320 0 0 0 Tile_X10Y2_DOUT_SRAM11
port 1346 nsew signal input
flabel metal2 s 452544 603752 452640 603832 0 FreeSans 320 0 0 0 Tile_X10Y2_DOUT_SRAM12
port 1347 nsew signal input
flabel metal2 s 452544 604256 452640 604336 0 FreeSans 320 0 0 0 Tile_X10Y2_DOUT_SRAM13
port 1348 nsew signal input
flabel metal2 s 452544 604760 452640 604840 0 FreeSans 320 0 0 0 Tile_X10Y2_DOUT_SRAM14
port 1349 nsew signal input
flabel metal2 s 452544 605264 452640 605344 0 FreeSans 320 0 0 0 Tile_X10Y2_DOUT_SRAM15
port 1350 nsew signal input
flabel metal2 s 452544 605768 452640 605848 0 FreeSans 320 0 0 0 Tile_X10Y2_DOUT_SRAM16
port 1351 nsew signal input
flabel metal2 s 452544 606272 452640 606352 0 FreeSans 320 0 0 0 Tile_X10Y2_DOUT_SRAM17
port 1352 nsew signal input
flabel metal2 s 452544 606776 452640 606856 0 FreeSans 320 0 0 0 Tile_X10Y2_DOUT_SRAM18
port 1353 nsew signal input
flabel metal2 s 452544 607280 452640 607360 0 FreeSans 320 0 0 0 Tile_X10Y2_DOUT_SRAM19
port 1354 nsew signal input
flabel metal2 s 452544 598712 452640 598792 0 FreeSans 320 0 0 0 Tile_X10Y2_DOUT_SRAM2
port 1355 nsew signal input
flabel metal2 s 452544 607784 452640 607864 0 FreeSans 320 0 0 0 Tile_X10Y2_DOUT_SRAM20
port 1356 nsew signal input
flabel metal2 s 452544 608288 452640 608368 0 FreeSans 320 0 0 0 Tile_X10Y2_DOUT_SRAM21
port 1357 nsew signal input
flabel metal2 s 452544 608792 452640 608872 0 FreeSans 320 0 0 0 Tile_X10Y2_DOUT_SRAM22
port 1358 nsew signal input
flabel metal2 s 452544 609296 452640 609376 0 FreeSans 320 0 0 0 Tile_X10Y2_DOUT_SRAM23
port 1359 nsew signal input
flabel metal2 s 452544 609800 452640 609880 0 FreeSans 320 0 0 0 Tile_X10Y2_DOUT_SRAM24
port 1360 nsew signal input
flabel metal2 s 452544 610304 452640 610384 0 FreeSans 320 0 0 0 Tile_X10Y2_DOUT_SRAM25
port 1361 nsew signal input
flabel metal2 s 452544 610808 452640 610888 0 FreeSans 320 0 0 0 Tile_X10Y2_DOUT_SRAM26
port 1362 nsew signal input
flabel metal2 s 452544 611312 452640 611392 0 FreeSans 320 0 0 0 Tile_X10Y2_DOUT_SRAM27
port 1363 nsew signal input
flabel metal2 s 452544 611816 452640 611896 0 FreeSans 320 0 0 0 Tile_X10Y2_DOUT_SRAM28
port 1364 nsew signal input
flabel metal2 s 452544 612320 452640 612400 0 FreeSans 320 0 0 0 Tile_X10Y2_DOUT_SRAM29
port 1365 nsew signal input
flabel metal2 s 452544 599216 452640 599296 0 FreeSans 320 0 0 0 Tile_X10Y2_DOUT_SRAM3
port 1366 nsew signal input
flabel metal2 s 452544 612824 452640 612904 0 FreeSans 320 0 0 0 Tile_X10Y2_DOUT_SRAM30
port 1367 nsew signal input
flabel metal2 s 452544 613328 452640 613408 0 FreeSans 320 0 0 0 Tile_X10Y2_DOUT_SRAM31
port 1368 nsew signal input
flabel metal2 s 452544 599720 452640 599800 0 FreeSans 320 0 0 0 Tile_X10Y2_DOUT_SRAM4
port 1369 nsew signal input
flabel metal2 s 452544 600224 452640 600304 0 FreeSans 320 0 0 0 Tile_X10Y2_DOUT_SRAM5
port 1370 nsew signal input
flabel metal2 s 452544 600728 452640 600808 0 FreeSans 320 0 0 0 Tile_X10Y2_DOUT_SRAM6
port 1371 nsew signal input
flabel metal2 s 452544 601232 452640 601312 0 FreeSans 320 0 0 0 Tile_X10Y2_DOUT_SRAM7
port 1372 nsew signal input
flabel metal2 s 452544 601736 452640 601816 0 FreeSans 320 0 0 0 Tile_X10Y2_DOUT_SRAM8
port 1373 nsew signal input
flabel metal2 s 452544 602240 452640 602320 0 FreeSans 320 0 0 0 Tile_X10Y2_DOUT_SRAM9
port 1374 nsew signal input
flabel metal2 s 452544 651632 452640 651712 0 FreeSans 320 0 0 0 Tile_X10Y2_MEN_SRAM
port 1375 nsew signal output
flabel metal2 s 452544 652136 452640 652216 0 FreeSans 320 0 0 0 Tile_X10Y2_REN_SRAM
port 1376 nsew signal output
flabel metal2 s 452544 652640 452640 652720 0 FreeSans 320 0 0 0 Tile_X10Y2_TIE_HIGH_SRAM
port 1377 nsew signal output
flabel metal2 s 452544 653144 452640 653224 0 FreeSans 320 0 0 0 Tile_X10Y2_TIE_LOW_SRAM
port 1378 nsew signal output
flabel metal2 s 452544 653648 452640 653728 0 FreeSans 320 0 0 0 Tile_X10Y2_WEN_SRAM
port 1379 nsew signal output
flabel metal2 s 452544 517064 452640 517144 0 FreeSans 320 0 0 0 Tile_X10Y4_ADDR_SRAM0
port 1380 nsew signal output
flabel metal2 s 452544 517568 452640 517648 0 FreeSans 320 0 0 0 Tile_X10Y4_ADDR_SRAM1
port 1381 nsew signal output
flabel metal2 s 452544 518072 452640 518152 0 FreeSans 320 0 0 0 Tile_X10Y4_ADDR_SRAM2
port 1382 nsew signal output
flabel metal2 s 452544 518576 452640 518656 0 FreeSans 320 0 0 0 Tile_X10Y4_ADDR_SRAM3
port 1383 nsew signal output
flabel metal2 s 452544 519080 452640 519160 0 FreeSans 320 0 0 0 Tile_X10Y4_ADDR_SRAM4
port 1384 nsew signal output
flabel metal2 s 452544 519584 452640 519664 0 FreeSans 320 0 0 0 Tile_X10Y4_ADDR_SRAM5
port 1385 nsew signal output
flabel metal2 s 452544 520088 452640 520168 0 FreeSans 320 0 0 0 Tile_X10Y4_ADDR_SRAM6
port 1386 nsew signal output
flabel metal2 s 452544 520592 452640 520672 0 FreeSans 320 0 0 0 Tile_X10Y4_ADDR_SRAM7
port 1387 nsew signal output
flabel metal2 s 452544 521096 452640 521176 0 FreeSans 320 0 0 0 Tile_X10Y4_ADDR_SRAM8
port 1388 nsew signal output
flabel metal2 s 452544 521600 452640 521680 0 FreeSans 320 0 0 0 Tile_X10Y4_ADDR_SRAM9
port 1389 nsew signal output
flabel metal2 s 452544 522104 452640 522184 0 FreeSans 320 0 0 0 Tile_X10Y4_BM_SRAM0
port 1390 nsew signal output
flabel metal2 s 452544 522608 452640 522688 0 FreeSans 320 0 0 0 Tile_X10Y4_BM_SRAM1
port 1391 nsew signal output
flabel metal2 s 452544 527144 452640 527224 0 FreeSans 320 0 0 0 Tile_X10Y4_BM_SRAM10
port 1392 nsew signal output
flabel metal2 s 452544 527648 452640 527728 0 FreeSans 320 0 0 0 Tile_X10Y4_BM_SRAM11
port 1393 nsew signal output
flabel metal2 s 452544 528152 452640 528232 0 FreeSans 320 0 0 0 Tile_X10Y4_BM_SRAM12
port 1394 nsew signal output
flabel metal2 s 452544 528656 452640 528736 0 FreeSans 320 0 0 0 Tile_X10Y4_BM_SRAM13
port 1395 nsew signal output
flabel metal2 s 452544 529160 452640 529240 0 FreeSans 320 0 0 0 Tile_X10Y4_BM_SRAM14
port 1396 nsew signal output
flabel metal2 s 452544 529664 452640 529744 0 FreeSans 320 0 0 0 Tile_X10Y4_BM_SRAM15
port 1397 nsew signal output
flabel metal2 s 452544 530168 452640 530248 0 FreeSans 320 0 0 0 Tile_X10Y4_BM_SRAM16
port 1398 nsew signal output
flabel metal2 s 452544 530672 452640 530752 0 FreeSans 320 0 0 0 Tile_X10Y4_BM_SRAM17
port 1399 nsew signal output
flabel metal2 s 452544 531176 452640 531256 0 FreeSans 320 0 0 0 Tile_X10Y4_BM_SRAM18
port 1400 nsew signal output
flabel metal2 s 452544 531680 452640 531760 0 FreeSans 320 0 0 0 Tile_X10Y4_BM_SRAM19
port 1401 nsew signal output
flabel metal2 s 452544 523112 452640 523192 0 FreeSans 320 0 0 0 Tile_X10Y4_BM_SRAM2
port 1402 nsew signal output
flabel metal2 s 452544 532184 452640 532264 0 FreeSans 320 0 0 0 Tile_X10Y4_BM_SRAM20
port 1403 nsew signal output
flabel metal2 s 452544 532688 452640 532768 0 FreeSans 320 0 0 0 Tile_X10Y4_BM_SRAM21
port 1404 nsew signal output
flabel metal2 s 452544 533192 452640 533272 0 FreeSans 320 0 0 0 Tile_X10Y4_BM_SRAM22
port 1405 nsew signal output
flabel metal2 s 452544 533696 452640 533776 0 FreeSans 320 0 0 0 Tile_X10Y4_BM_SRAM23
port 1406 nsew signal output
flabel metal2 s 452544 534200 452640 534280 0 FreeSans 320 0 0 0 Tile_X10Y4_BM_SRAM24
port 1407 nsew signal output
flabel metal2 s 452544 534704 452640 534784 0 FreeSans 320 0 0 0 Tile_X10Y4_BM_SRAM25
port 1408 nsew signal output
flabel metal2 s 452544 535208 452640 535288 0 FreeSans 320 0 0 0 Tile_X10Y4_BM_SRAM26
port 1409 nsew signal output
flabel metal2 s 452544 535712 452640 535792 0 FreeSans 320 0 0 0 Tile_X10Y4_BM_SRAM27
port 1410 nsew signal output
flabel metal2 s 452544 536216 452640 536296 0 FreeSans 320 0 0 0 Tile_X10Y4_BM_SRAM28
port 1411 nsew signal output
flabel metal2 s 452544 536720 452640 536800 0 FreeSans 320 0 0 0 Tile_X10Y4_BM_SRAM29
port 1412 nsew signal output
flabel metal2 s 452544 523616 452640 523696 0 FreeSans 320 0 0 0 Tile_X10Y4_BM_SRAM3
port 1413 nsew signal output
flabel metal2 s 452544 537224 452640 537304 0 FreeSans 320 0 0 0 Tile_X10Y4_BM_SRAM30
port 1414 nsew signal output
flabel metal2 s 452544 537728 452640 537808 0 FreeSans 320 0 0 0 Tile_X10Y4_BM_SRAM31
port 1415 nsew signal output
flabel metal2 s 452544 524120 452640 524200 0 FreeSans 320 0 0 0 Tile_X10Y4_BM_SRAM4
port 1416 nsew signal output
flabel metal2 s 452544 524624 452640 524704 0 FreeSans 320 0 0 0 Tile_X10Y4_BM_SRAM5
port 1417 nsew signal output
flabel metal2 s 452544 525128 452640 525208 0 FreeSans 320 0 0 0 Tile_X10Y4_BM_SRAM6
port 1418 nsew signal output
flabel metal2 s 452544 525632 452640 525712 0 FreeSans 320 0 0 0 Tile_X10Y4_BM_SRAM7
port 1419 nsew signal output
flabel metal2 s 452544 526136 452640 526216 0 FreeSans 320 0 0 0 Tile_X10Y4_BM_SRAM8
port 1420 nsew signal output
flabel metal2 s 452544 526640 452640 526720 0 FreeSans 320 0 0 0 Tile_X10Y4_BM_SRAM9
port 1421 nsew signal output
flabel metal2 s 452544 538232 452640 538312 0 FreeSans 320 0 0 0 Tile_X10Y4_CLK_SRAM
port 1422 nsew signal output
flabel metal2 s 452544 500432 452640 500512 0 FreeSans 320 0 0 0 Tile_X10Y4_CONFIGURED_top
port 1423 nsew signal input
flabel metal2 s 452544 538736 452640 538816 0 FreeSans 320 0 0 0 Tile_X10Y4_DIN_SRAM0
port 1424 nsew signal output
flabel metal2 s 452544 539240 452640 539320 0 FreeSans 320 0 0 0 Tile_X10Y4_DIN_SRAM1
port 1425 nsew signal output
flabel metal2 s 452544 543776 452640 543856 0 FreeSans 320 0 0 0 Tile_X10Y4_DIN_SRAM10
port 1426 nsew signal output
flabel metal2 s 452544 544280 452640 544360 0 FreeSans 320 0 0 0 Tile_X10Y4_DIN_SRAM11
port 1427 nsew signal output
flabel metal2 s 452544 544784 452640 544864 0 FreeSans 320 0 0 0 Tile_X10Y4_DIN_SRAM12
port 1428 nsew signal output
flabel metal2 s 452544 545288 452640 545368 0 FreeSans 320 0 0 0 Tile_X10Y4_DIN_SRAM13
port 1429 nsew signal output
flabel metal2 s 452544 545792 452640 545872 0 FreeSans 320 0 0 0 Tile_X10Y4_DIN_SRAM14
port 1430 nsew signal output
flabel metal2 s 452544 546296 452640 546376 0 FreeSans 320 0 0 0 Tile_X10Y4_DIN_SRAM15
port 1431 nsew signal output
flabel metal2 s 452544 546800 452640 546880 0 FreeSans 320 0 0 0 Tile_X10Y4_DIN_SRAM16
port 1432 nsew signal output
flabel metal2 s 452544 547304 452640 547384 0 FreeSans 320 0 0 0 Tile_X10Y4_DIN_SRAM17
port 1433 nsew signal output
flabel metal2 s 452544 547808 452640 547888 0 FreeSans 320 0 0 0 Tile_X10Y4_DIN_SRAM18
port 1434 nsew signal output
flabel metal2 s 452544 548312 452640 548392 0 FreeSans 320 0 0 0 Tile_X10Y4_DIN_SRAM19
port 1435 nsew signal output
flabel metal2 s 452544 539744 452640 539824 0 FreeSans 320 0 0 0 Tile_X10Y4_DIN_SRAM2
port 1436 nsew signal output
flabel metal2 s 452544 548816 452640 548896 0 FreeSans 320 0 0 0 Tile_X10Y4_DIN_SRAM20
port 1437 nsew signal output
flabel metal2 s 452544 549320 452640 549400 0 FreeSans 320 0 0 0 Tile_X10Y4_DIN_SRAM21
port 1438 nsew signal output
flabel metal2 s 452544 549824 452640 549904 0 FreeSans 320 0 0 0 Tile_X10Y4_DIN_SRAM22
port 1439 nsew signal output
flabel metal2 s 452544 550328 452640 550408 0 FreeSans 320 0 0 0 Tile_X10Y4_DIN_SRAM23
port 1440 nsew signal output
flabel metal2 s 452544 550832 452640 550912 0 FreeSans 320 0 0 0 Tile_X10Y4_DIN_SRAM24
port 1441 nsew signal output
flabel metal2 s 452544 551336 452640 551416 0 FreeSans 320 0 0 0 Tile_X10Y4_DIN_SRAM25
port 1442 nsew signal output
flabel metal2 s 452544 551840 452640 551920 0 FreeSans 320 0 0 0 Tile_X10Y4_DIN_SRAM26
port 1443 nsew signal output
flabel metal2 s 452544 552344 452640 552424 0 FreeSans 320 0 0 0 Tile_X10Y4_DIN_SRAM27
port 1444 nsew signal output
flabel metal2 s 452544 552848 452640 552928 0 FreeSans 320 0 0 0 Tile_X10Y4_DIN_SRAM28
port 1445 nsew signal output
flabel metal2 s 452544 553352 452640 553432 0 FreeSans 320 0 0 0 Tile_X10Y4_DIN_SRAM29
port 1446 nsew signal output
flabel metal2 s 452544 540248 452640 540328 0 FreeSans 320 0 0 0 Tile_X10Y4_DIN_SRAM3
port 1447 nsew signal output
flabel metal2 s 452544 553856 452640 553936 0 FreeSans 320 0 0 0 Tile_X10Y4_DIN_SRAM30
port 1448 nsew signal output
flabel metal2 s 452544 554360 452640 554440 0 FreeSans 320 0 0 0 Tile_X10Y4_DIN_SRAM31
port 1449 nsew signal output
flabel metal2 s 452544 540752 452640 540832 0 FreeSans 320 0 0 0 Tile_X10Y4_DIN_SRAM4
port 1450 nsew signal output
flabel metal2 s 452544 541256 452640 541336 0 FreeSans 320 0 0 0 Tile_X10Y4_DIN_SRAM5
port 1451 nsew signal output
flabel metal2 s 452544 541760 452640 541840 0 FreeSans 320 0 0 0 Tile_X10Y4_DIN_SRAM6
port 1452 nsew signal output
flabel metal2 s 452544 542264 452640 542344 0 FreeSans 320 0 0 0 Tile_X10Y4_DIN_SRAM7
port 1453 nsew signal output
flabel metal2 s 452544 542768 452640 542848 0 FreeSans 320 0 0 0 Tile_X10Y4_DIN_SRAM8
port 1454 nsew signal output
flabel metal2 s 452544 543272 452640 543352 0 FreeSans 320 0 0 0 Tile_X10Y4_DIN_SRAM9
port 1455 nsew signal output
flabel metal2 s 452544 500936 452640 501016 0 FreeSans 320 0 0 0 Tile_X10Y4_DOUT_SRAM0
port 1456 nsew signal input
flabel metal2 s 452544 501440 452640 501520 0 FreeSans 320 0 0 0 Tile_X10Y4_DOUT_SRAM1
port 1457 nsew signal input
flabel metal2 s 452544 505976 452640 506056 0 FreeSans 320 0 0 0 Tile_X10Y4_DOUT_SRAM10
port 1458 nsew signal input
flabel metal2 s 452544 506480 452640 506560 0 FreeSans 320 0 0 0 Tile_X10Y4_DOUT_SRAM11
port 1459 nsew signal input
flabel metal2 s 452544 506984 452640 507064 0 FreeSans 320 0 0 0 Tile_X10Y4_DOUT_SRAM12
port 1460 nsew signal input
flabel metal2 s 452544 507488 452640 507568 0 FreeSans 320 0 0 0 Tile_X10Y4_DOUT_SRAM13
port 1461 nsew signal input
flabel metal2 s 452544 507992 452640 508072 0 FreeSans 320 0 0 0 Tile_X10Y4_DOUT_SRAM14
port 1462 nsew signal input
flabel metal2 s 452544 508496 452640 508576 0 FreeSans 320 0 0 0 Tile_X10Y4_DOUT_SRAM15
port 1463 nsew signal input
flabel metal2 s 452544 509000 452640 509080 0 FreeSans 320 0 0 0 Tile_X10Y4_DOUT_SRAM16
port 1464 nsew signal input
flabel metal2 s 452544 509504 452640 509584 0 FreeSans 320 0 0 0 Tile_X10Y4_DOUT_SRAM17
port 1465 nsew signal input
flabel metal2 s 452544 510008 452640 510088 0 FreeSans 320 0 0 0 Tile_X10Y4_DOUT_SRAM18
port 1466 nsew signal input
flabel metal2 s 452544 510512 452640 510592 0 FreeSans 320 0 0 0 Tile_X10Y4_DOUT_SRAM19
port 1467 nsew signal input
flabel metal2 s 452544 501944 452640 502024 0 FreeSans 320 0 0 0 Tile_X10Y4_DOUT_SRAM2
port 1468 nsew signal input
flabel metal2 s 452544 511016 452640 511096 0 FreeSans 320 0 0 0 Tile_X10Y4_DOUT_SRAM20
port 1469 nsew signal input
flabel metal2 s 452544 511520 452640 511600 0 FreeSans 320 0 0 0 Tile_X10Y4_DOUT_SRAM21
port 1470 nsew signal input
flabel metal2 s 452544 512024 452640 512104 0 FreeSans 320 0 0 0 Tile_X10Y4_DOUT_SRAM22
port 1471 nsew signal input
flabel metal2 s 452544 512528 452640 512608 0 FreeSans 320 0 0 0 Tile_X10Y4_DOUT_SRAM23
port 1472 nsew signal input
flabel metal2 s 452544 513032 452640 513112 0 FreeSans 320 0 0 0 Tile_X10Y4_DOUT_SRAM24
port 1473 nsew signal input
flabel metal2 s 452544 513536 452640 513616 0 FreeSans 320 0 0 0 Tile_X10Y4_DOUT_SRAM25
port 1474 nsew signal input
flabel metal2 s 452544 514040 452640 514120 0 FreeSans 320 0 0 0 Tile_X10Y4_DOUT_SRAM26
port 1475 nsew signal input
flabel metal2 s 452544 514544 452640 514624 0 FreeSans 320 0 0 0 Tile_X10Y4_DOUT_SRAM27
port 1476 nsew signal input
flabel metal2 s 452544 515048 452640 515128 0 FreeSans 320 0 0 0 Tile_X10Y4_DOUT_SRAM28
port 1477 nsew signal input
flabel metal2 s 452544 515552 452640 515632 0 FreeSans 320 0 0 0 Tile_X10Y4_DOUT_SRAM29
port 1478 nsew signal input
flabel metal2 s 452544 502448 452640 502528 0 FreeSans 320 0 0 0 Tile_X10Y4_DOUT_SRAM3
port 1479 nsew signal input
flabel metal2 s 452544 516056 452640 516136 0 FreeSans 320 0 0 0 Tile_X10Y4_DOUT_SRAM30
port 1480 nsew signal input
flabel metal2 s 452544 516560 452640 516640 0 FreeSans 320 0 0 0 Tile_X10Y4_DOUT_SRAM31
port 1481 nsew signal input
flabel metal2 s 452544 502952 452640 503032 0 FreeSans 320 0 0 0 Tile_X10Y4_DOUT_SRAM4
port 1482 nsew signal input
flabel metal2 s 452544 503456 452640 503536 0 FreeSans 320 0 0 0 Tile_X10Y4_DOUT_SRAM5
port 1483 nsew signal input
flabel metal2 s 452544 503960 452640 504040 0 FreeSans 320 0 0 0 Tile_X10Y4_DOUT_SRAM6
port 1484 nsew signal input
flabel metal2 s 452544 504464 452640 504544 0 FreeSans 320 0 0 0 Tile_X10Y4_DOUT_SRAM7
port 1485 nsew signal input
flabel metal2 s 452544 504968 452640 505048 0 FreeSans 320 0 0 0 Tile_X10Y4_DOUT_SRAM8
port 1486 nsew signal input
flabel metal2 s 452544 505472 452640 505552 0 FreeSans 320 0 0 0 Tile_X10Y4_DOUT_SRAM9
port 1487 nsew signal input
flabel metal2 s 452544 554864 452640 554944 0 FreeSans 320 0 0 0 Tile_X10Y4_MEN_SRAM
port 1488 nsew signal output
flabel metal2 s 452544 555368 452640 555448 0 FreeSans 320 0 0 0 Tile_X10Y4_REN_SRAM
port 1489 nsew signal output
flabel metal2 s 452544 555872 452640 555952 0 FreeSans 320 0 0 0 Tile_X10Y4_TIE_HIGH_SRAM
port 1490 nsew signal output
flabel metal2 s 452544 556376 452640 556456 0 FreeSans 320 0 0 0 Tile_X10Y4_TIE_LOW_SRAM
port 1491 nsew signal output
flabel metal2 s 452544 556880 452640 556960 0 FreeSans 320 0 0 0 Tile_X10Y4_WEN_SRAM
port 1492 nsew signal output
flabel metal2 s 452544 420296 452640 420376 0 FreeSans 320 0 0 0 Tile_X10Y6_ADDR_SRAM0
port 1493 nsew signal output
flabel metal2 s 452544 420800 452640 420880 0 FreeSans 320 0 0 0 Tile_X10Y6_ADDR_SRAM1
port 1494 nsew signal output
flabel metal2 s 452544 421304 452640 421384 0 FreeSans 320 0 0 0 Tile_X10Y6_ADDR_SRAM2
port 1495 nsew signal output
flabel metal2 s 452544 421808 452640 421888 0 FreeSans 320 0 0 0 Tile_X10Y6_ADDR_SRAM3
port 1496 nsew signal output
flabel metal2 s 452544 422312 452640 422392 0 FreeSans 320 0 0 0 Tile_X10Y6_ADDR_SRAM4
port 1497 nsew signal output
flabel metal2 s 452544 422816 452640 422896 0 FreeSans 320 0 0 0 Tile_X10Y6_ADDR_SRAM5
port 1498 nsew signal output
flabel metal2 s 452544 423320 452640 423400 0 FreeSans 320 0 0 0 Tile_X10Y6_ADDR_SRAM6
port 1499 nsew signal output
flabel metal2 s 452544 423824 452640 423904 0 FreeSans 320 0 0 0 Tile_X10Y6_ADDR_SRAM7
port 1500 nsew signal output
flabel metal2 s 452544 424328 452640 424408 0 FreeSans 320 0 0 0 Tile_X10Y6_ADDR_SRAM8
port 1501 nsew signal output
flabel metal2 s 452544 424832 452640 424912 0 FreeSans 320 0 0 0 Tile_X10Y6_ADDR_SRAM9
port 1502 nsew signal output
flabel metal2 s 452544 425336 452640 425416 0 FreeSans 320 0 0 0 Tile_X10Y6_BM_SRAM0
port 1503 nsew signal output
flabel metal2 s 452544 425840 452640 425920 0 FreeSans 320 0 0 0 Tile_X10Y6_BM_SRAM1
port 1504 nsew signal output
flabel metal2 s 452544 430376 452640 430456 0 FreeSans 320 0 0 0 Tile_X10Y6_BM_SRAM10
port 1505 nsew signal output
flabel metal2 s 452544 430880 452640 430960 0 FreeSans 320 0 0 0 Tile_X10Y6_BM_SRAM11
port 1506 nsew signal output
flabel metal2 s 452544 431384 452640 431464 0 FreeSans 320 0 0 0 Tile_X10Y6_BM_SRAM12
port 1507 nsew signal output
flabel metal2 s 452544 431888 452640 431968 0 FreeSans 320 0 0 0 Tile_X10Y6_BM_SRAM13
port 1508 nsew signal output
flabel metal2 s 452544 432392 452640 432472 0 FreeSans 320 0 0 0 Tile_X10Y6_BM_SRAM14
port 1509 nsew signal output
flabel metal2 s 452544 432896 452640 432976 0 FreeSans 320 0 0 0 Tile_X10Y6_BM_SRAM15
port 1510 nsew signal output
flabel metal2 s 452544 433400 452640 433480 0 FreeSans 320 0 0 0 Tile_X10Y6_BM_SRAM16
port 1511 nsew signal output
flabel metal2 s 452544 433904 452640 433984 0 FreeSans 320 0 0 0 Tile_X10Y6_BM_SRAM17
port 1512 nsew signal output
flabel metal2 s 452544 434408 452640 434488 0 FreeSans 320 0 0 0 Tile_X10Y6_BM_SRAM18
port 1513 nsew signal output
flabel metal2 s 452544 434912 452640 434992 0 FreeSans 320 0 0 0 Tile_X10Y6_BM_SRAM19
port 1514 nsew signal output
flabel metal2 s 452544 426344 452640 426424 0 FreeSans 320 0 0 0 Tile_X10Y6_BM_SRAM2
port 1515 nsew signal output
flabel metal2 s 452544 435416 452640 435496 0 FreeSans 320 0 0 0 Tile_X10Y6_BM_SRAM20
port 1516 nsew signal output
flabel metal2 s 452544 435920 452640 436000 0 FreeSans 320 0 0 0 Tile_X10Y6_BM_SRAM21
port 1517 nsew signal output
flabel metal2 s 452544 436424 452640 436504 0 FreeSans 320 0 0 0 Tile_X10Y6_BM_SRAM22
port 1518 nsew signal output
flabel metal2 s 452544 436928 452640 437008 0 FreeSans 320 0 0 0 Tile_X10Y6_BM_SRAM23
port 1519 nsew signal output
flabel metal2 s 452544 437432 452640 437512 0 FreeSans 320 0 0 0 Tile_X10Y6_BM_SRAM24
port 1520 nsew signal output
flabel metal2 s 452544 437936 452640 438016 0 FreeSans 320 0 0 0 Tile_X10Y6_BM_SRAM25
port 1521 nsew signal output
flabel metal2 s 452544 438440 452640 438520 0 FreeSans 320 0 0 0 Tile_X10Y6_BM_SRAM26
port 1522 nsew signal output
flabel metal2 s 452544 438944 452640 439024 0 FreeSans 320 0 0 0 Tile_X10Y6_BM_SRAM27
port 1523 nsew signal output
flabel metal2 s 452544 439448 452640 439528 0 FreeSans 320 0 0 0 Tile_X10Y6_BM_SRAM28
port 1524 nsew signal output
flabel metal2 s 452544 439952 452640 440032 0 FreeSans 320 0 0 0 Tile_X10Y6_BM_SRAM29
port 1525 nsew signal output
flabel metal2 s 452544 426848 452640 426928 0 FreeSans 320 0 0 0 Tile_X10Y6_BM_SRAM3
port 1526 nsew signal output
flabel metal2 s 452544 440456 452640 440536 0 FreeSans 320 0 0 0 Tile_X10Y6_BM_SRAM30
port 1527 nsew signal output
flabel metal2 s 452544 440960 452640 441040 0 FreeSans 320 0 0 0 Tile_X10Y6_BM_SRAM31
port 1528 nsew signal output
flabel metal2 s 452544 427352 452640 427432 0 FreeSans 320 0 0 0 Tile_X10Y6_BM_SRAM4
port 1529 nsew signal output
flabel metal2 s 452544 427856 452640 427936 0 FreeSans 320 0 0 0 Tile_X10Y6_BM_SRAM5
port 1530 nsew signal output
flabel metal2 s 452544 428360 452640 428440 0 FreeSans 320 0 0 0 Tile_X10Y6_BM_SRAM6
port 1531 nsew signal output
flabel metal2 s 452544 428864 452640 428944 0 FreeSans 320 0 0 0 Tile_X10Y6_BM_SRAM7
port 1532 nsew signal output
flabel metal2 s 452544 429368 452640 429448 0 FreeSans 320 0 0 0 Tile_X10Y6_BM_SRAM8
port 1533 nsew signal output
flabel metal2 s 452544 429872 452640 429952 0 FreeSans 320 0 0 0 Tile_X10Y6_BM_SRAM9
port 1534 nsew signal output
flabel metal2 s 452544 441464 452640 441544 0 FreeSans 320 0 0 0 Tile_X10Y6_CLK_SRAM
port 1535 nsew signal output
flabel metal2 s 452544 403664 452640 403744 0 FreeSans 320 0 0 0 Tile_X10Y6_CONFIGURED_top
port 1536 nsew signal input
flabel metal2 s 452544 441968 452640 442048 0 FreeSans 320 0 0 0 Tile_X10Y6_DIN_SRAM0
port 1537 nsew signal output
flabel metal2 s 452544 442472 452640 442552 0 FreeSans 320 0 0 0 Tile_X10Y6_DIN_SRAM1
port 1538 nsew signal output
flabel metal2 s 452544 447008 452640 447088 0 FreeSans 320 0 0 0 Tile_X10Y6_DIN_SRAM10
port 1539 nsew signal output
flabel metal2 s 452544 447512 452640 447592 0 FreeSans 320 0 0 0 Tile_X10Y6_DIN_SRAM11
port 1540 nsew signal output
flabel metal2 s 452544 448016 452640 448096 0 FreeSans 320 0 0 0 Tile_X10Y6_DIN_SRAM12
port 1541 nsew signal output
flabel metal2 s 452544 448520 452640 448600 0 FreeSans 320 0 0 0 Tile_X10Y6_DIN_SRAM13
port 1542 nsew signal output
flabel metal2 s 452544 449024 452640 449104 0 FreeSans 320 0 0 0 Tile_X10Y6_DIN_SRAM14
port 1543 nsew signal output
flabel metal2 s 452544 449528 452640 449608 0 FreeSans 320 0 0 0 Tile_X10Y6_DIN_SRAM15
port 1544 nsew signal output
flabel metal2 s 452544 450032 452640 450112 0 FreeSans 320 0 0 0 Tile_X10Y6_DIN_SRAM16
port 1545 nsew signal output
flabel metal2 s 452544 450536 452640 450616 0 FreeSans 320 0 0 0 Tile_X10Y6_DIN_SRAM17
port 1546 nsew signal output
flabel metal2 s 452544 451040 452640 451120 0 FreeSans 320 0 0 0 Tile_X10Y6_DIN_SRAM18
port 1547 nsew signal output
flabel metal2 s 452544 451544 452640 451624 0 FreeSans 320 0 0 0 Tile_X10Y6_DIN_SRAM19
port 1548 nsew signal output
flabel metal2 s 452544 442976 452640 443056 0 FreeSans 320 0 0 0 Tile_X10Y6_DIN_SRAM2
port 1549 nsew signal output
flabel metal2 s 452544 452048 452640 452128 0 FreeSans 320 0 0 0 Tile_X10Y6_DIN_SRAM20
port 1550 nsew signal output
flabel metal2 s 452544 452552 452640 452632 0 FreeSans 320 0 0 0 Tile_X10Y6_DIN_SRAM21
port 1551 nsew signal output
flabel metal2 s 452544 453056 452640 453136 0 FreeSans 320 0 0 0 Tile_X10Y6_DIN_SRAM22
port 1552 nsew signal output
flabel metal2 s 452544 453560 452640 453640 0 FreeSans 320 0 0 0 Tile_X10Y6_DIN_SRAM23
port 1553 nsew signal output
flabel metal2 s 452544 454064 452640 454144 0 FreeSans 320 0 0 0 Tile_X10Y6_DIN_SRAM24
port 1554 nsew signal output
flabel metal2 s 452544 454568 452640 454648 0 FreeSans 320 0 0 0 Tile_X10Y6_DIN_SRAM25
port 1555 nsew signal output
flabel metal2 s 452544 455072 452640 455152 0 FreeSans 320 0 0 0 Tile_X10Y6_DIN_SRAM26
port 1556 nsew signal output
flabel metal2 s 452544 455576 452640 455656 0 FreeSans 320 0 0 0 Tile_X10Y6_DIN_SRAM27
port 1557 nsew signal output
flabel metal2 s 452544 456080 452640 456160 0 FreeSans 320 0 0 0 Tile_X10Y6_DIN_SRAM28
port 1558 nsew signal output
flabel metal2 s 452544 456584 452640 456664 0 FreeSans 320 0 0 0 Tile_X10Y6_DIN_SRAM29
port 1559 nsew signal output
flabel metal2 s 452544 443480 452640 443560 0 FreeSans 320 0 0 0 Tile_X10Y6_DIN_SRAM3
port 1560 nsew signal output
flabel metal2 s 452544 457088 452640 457168 0 FreeSans 320 0 0 0 Tile_X10Y6_DIN_SRAM30
port 1561 nsew signal output
flabel metal2 s 452544 457592 452640 457672 0 FreeSans 320 0 0 0 Tile_X10Y6_DIN_SRAM31
port 1562 nsew signal output
flabel metal2 s 452544 443984 452640 444064 0 FreeSans 320 0 0 0 Tile_X10Y6_DIN_SRAM4
port 1563 nsew signal output
flabel metal2 s 452544 444488 452640 444568 0 FreeSans 320 0 0 0 Tile_X10Y6_DIN_SRAM5
port 1564 nsew signal output
flabel metal2 s 452544 444992 452640 445072 0 FreeSans 320 0 0 0 Tile_X10Y6_DIN_SRAM6
port 1565 nsew signal output
flabel metal2 s 452544 445496 452640 445576 0 FreeSans 320 0 0 0 Tile_X10Y6_DIN_SRAM7
port 1566 nsew signal output
flabel metal2 s 452544 446000 452640 446080 0 FreeSans 320 0 0 0 Tile_X10Y6_DIN_SRAM8
port 1567 nsew signal output
flabel metal2 s 452544 446504 452640 446584 0 FreeSans 320 0 0 0 Tile_X10Y6_DIN_SRAM9
port 1568 nsew signal output
flabel metal2 s 452544 404168 452640 404248 0 FreeSans 320 0 0 0 Tile_X10Y6_DOUT_SRAM0
port 1569 nsew signal input
flabel metal2 s 452544 404672 452640 404752 0 FreeSans 320 0 0 0 Tile_X10Y6_DOUT_SRAM1
port 1570 nsew signal input
flabel metal2 s 452544 409208 452640 409288 0 FreeSans 320 0 0 0 Tile_X10Y6_DOUT_SRAM10
port 1571 nsew signal input
flabel metal2 s 452544 409712 452640 409792 0 FreeSans 320 0 0 0 Tile_X10Y6_DOUT_SRAM11
port 1572 nsew signal input
flabel metal2 s 452544 410216 452640 410296 0 FreeSans 320 0 0 0 Tile_X10Y6_DOUT_SRAM12
port 1573 nsew signal input
flabel metal2 s 452544 410720 452640 410800 0 FreeSans 320 0 0 0 Tile_X10Y6_DOUT_SRAM13
port 1574 nsew signal input
flabel metal2 s 452544 411224 452640 411304 0 FreeSans 320 0 0 0 Tile_X10Y6_DOUT_SRAM14
port 1575 nsew signal input
flabel metal2 s 452544 411728 452640 411808 0 FreeSans 320 0 0 0 Tile_X10Y6_DOUT_SRAM15
port 1576 nsew signal input
flabel metal2 s 452544 412232 452640 412312 0 FreeSans 320 0 0 0 Tile_X10Y6_DOUT_SRAM16
port 1577 nsew signal input
flabel metal2 s 452544 412736 452640 412816 0 FreeSans 320 0 0 0 Tile_X10Y6_DOUT_SRAM17
port 1578 nsew signal input
flabel metal2 s 452544 413240 452640 413320 0 FreeSans 320 0 0 0 Tile_X10Y6_DOUT_SRAM18
port 1579 nsew signal input
flabel metal2 s 452544 413744 452640 413824 0 FreeSans 320 0 0 0 Tile_X10Y6_DOUT_SRAM19
port 1580 nsew signal input
flabel metal2 s 452544 405176 452640 405256 0 FreeSans 320 0 0 0 Tile_X10Y6_DOUT_SRAM2
port 1581 nsew signal input
flabel metal2 s 452544 414248 452640 414328 0 FreeSans 320 0 0 0 Tile_X10Y6_DOUT_SRAM20
port 1582 nsew signal input
flabel metal2 s 452544 414752 452640 414832 0 FreeSans 320 0 0 0 Tile_X10Y6_DOUT_SRAM21
port 1583 nsew signal input
flabel metal2 s 452544 415256 452640 415336 0 FreeSans 320 0 0 0 Tile_X10Y6_DOUT_SRAM22
port 1584 nsew signal input
flabel metal2 s 452544 415760 452640 415840 0 FreeSans 320 0 0 0 Tile_X10Y6_DOUT_SRAM23
port 1585 nsew signal input
flabel metal2 s 452544 416264 452640 416344 0 FreeSans 320 0 0 0 Tile_X10Y6_DOUT_SRAM24
port 1586 nsew signal input
flabel metal2 s 452544 416768 452640 416848 0 FreeSans 320 0 0 0 Tile_X10Y6_DOUT_SRAM25
port 1587 nsew signal input
flabel metal2 s 452544 417272 452640 417352 0 FreeSans 320 0 0 0 Tile_X10Y6_DOUT_SRAM26
port 1588 nsew signal input
flabel metal2 s 452544 417776 452640 417856 0 FreeSans 320 0 0 0 Tile_X10Y6_DOUT_SRAM27
port 1589 nsew signal input
flabel metal2 s 452544 418280 452640 418360 0 FreeSans 320 0 0 0 Tile_X10Y6_DOUT_SRAM28
port 1590 nsew signal input
flabel metal2 s 452544 418784 452640 418864 0 FreeSans 320 0 0 0 Tile_X10Y6_DOUT_SRAM29
port 1591 nsew signal input
flabel metal2 s 452544 405680 452640 405760 0 FreeSans 320 0 0 0 Tile_X10Y6_DOUT_SRAM3
port 1592 nsew signal input
flabel metal2 s 452544 419288 452640 419368 0 FreeSans 320 0 0 0 Tile_X10Y6_DOUT_SRAM30
port 1593 nsew signal input
flabel metal2 s 452544 419792 452640 419872 0 FreeSans 320 0 0 0 Tile_X10Y6_DOUT_SRAM31
port 1594 nsew signal input
flabel metal2 s 452544 406184 452640 406264 0 FreeSans 320 0 0 0 Tile_X10Y6_DOUT_SRAM4
port 1595 nsew signal input
flabel metal2 s 452544 406688 452640 406768 0 FreeSans 320 0 0 0 Tile_X10Y6_DOUT_SRAM5
port 1596 nsew signal input
flabel metal2 s 452544 407192 452640 407272 0 FreeSans 320 0 0 0 Tile_X10Y6_DOUT_SRAM6
port 1597 nsew signal input
flabel metal2 s 452544 407696 452640 407776 0 FreeSans 320 0 0 0 Tile_X10Y6_DOUT_SRAM7
port 1598 nsew signal input
flabel metal2 s 452544 408200 452640 408280 0 FreeSans 320 0 0 0 Tile_X10Y6_DOUT_SRAM8
port 1599 nsew signal input
flabel metal2 s 452544 408704 452640 408784 0 FreeSans 320 0 0 0 Tile_X10Y6_DOUT_SRAM9
port 1600 nsew signal input
flabel metal2 s 452544 458096 452640 458176 0 FreeSans 320 0 0 0 Tile_X10Y6_MEN_SRAM
port 1601 nsew signal output
flabel metal2 s 452544 458600 452640 458680 0 FreeSans 320 0 0 0 Tile_X10Y6_REN_SRAM
port 1602 nsew signal output
flabel metal2 s 452544 459104 452640 459184 0 FreeSans 320 0 0 0 Tile_X10Y6_TIE_HIGH_SRAM
port 1603 nsew signal output
flabel metal2 s 452544 459608 452640 459688 0 FreeSans 320 0 0 0 Tile_X10Y6_TIE_LOW_SRAM
port 1604 nsew signal output
flabel metal2 s 452544 460112 452640 460192 0 FreeSans 320 0 0 0 Tile_X10Y6_WEN_SRAM
port 1605 nsew signal output
flabel metal2 s 452544 323528 452640 323608 0 FreeSans 320 0 0 0 Tile_X10Y8_ADDR_SRAM0
port 1606 nsew signal output
flabel metal2 s 452544 324032 452640 324112 0 FreeSans 320 0 0 0 Tile_X10Y8_ADDR_SRAM1
port 1607 nsew signal output
flabel metal2 s 452544 324536 452640 324616 0 FreeSans 320 0 0 0 Tile_X10Y8_ADDR_SRAM2
port 1608 nsew signal output
flabel metal2 s 452544 325040 452640 325120 0 FreeSans 320 0 0 0 Tile_X10Y8_ADDR_SRAM3
port 1609 nsew signal output
flabel metal2 s 452544 325544 452640 325624 0 FreeSans 320 0 0 0 Tile_X10Y8_ADDR_SRAM4
port 1610 nsew signal output
flabel metal2 s 452544 326048 452640 326128 0 FreeSans 320 0 0 0 Tile_X10Y8_ADDR_SRAM5
port 1611 nsew signal output
flabel metal2 s 452544 326552 452640 326632 0 FreeSans 320 0 0 0 Tile_X10Y8_ADDR_SRAM6
port 1612 nsew signal output
flabel metal2 s 452544 327056 452640 327136 0 FreeSans 320 0 0 0 Tile_X10Y8_ADDR_SRAM7
port 1613 nsew signal output
flabel metal2 s 452544 327560 452640 327640 0 FreeSans 320 0 0 0 Tile_X10Y8_ADDR_SRAM8
port 1614 nsew signal output
flabel metal2 s 452544 328064 452640 328144 0 FreeSans 320 0 0 0 Tile_X10Y8_ADDR_SRAM9
port 1615 nsew signal output
flabel metal2 s 452544 328568 452640 328648 0 FreeSans 320 0 0 0 Tile_X10Y8_BM_SRAM0
port 1616 nsew signal output
flabel metal2 s 452544 329072 452640 329152 0 FreeSans 320 0 0 0 Tile_X10Y8_BM_SRAM1
port 1617 nsew signal output
flabel metal2 s 452544 333608 452640 333688 0 FreeSans 320 0 0 0 Tile_X10Y8_BM_SRAM10
port 1618 nsew signal output
flabel metal2 s 452544 334112 452640 334192 0 FreeSans 320 0 0 0 Tile_X10Y8_BM_SRAM11
port 1619 nsew signal output
flabel metal2 s 452544 334616 452640 334696 0 FreeSans 320 0 0 0 Tile_X10Y8_BM_SRAM12
port 1620 nsew signal output
flabel metal2 s 452544 335120 452640 335200 0 FreeSans 320 0 0 0 Tile_X10Y8_BM_SRAM13
port 1621 nsew signal output
flabel metal2 s 452544 335624 452640 335704 0 FreeSans 320 0 0 0 Tile_X10Y8_BM_SRAM14
port 1622 nsew signal output
flabel metal2 s 452544 336128 452640 336208 0 FreeSans 320 0 0 0 Tile_X10Y8_BM_SRAM15
port 1623 nsew signal output
flabel metal2 s 452544 336632 452640 336712 0 FreeSans 320 0 0 0 Tile_X10Y8_BM_SRAM16
port 1624 nsew signal output
flabel metal2 s 452544 337136 452640 337216 0 FreeSans 320 0 0 0 Tile_X10Y8_BM_SRAM17
port 1625 nsew signal output
flabel metal2 s 452544 337640 452640 337720 0 FreeSans 320 0 0 0 Tile_X10Y8_BM_SRAM18
port 1626 nsew signal output
flabel metal2 s 452544 338144 452640 338224 0 FreeSans 320 0 0 0 Tile_X10Y8_BM_SRAM19
port 1627 nsew signal output
flabel metal2 s 452544 329576 452640 329656 0 FreeSans 320 0 0 0 Tile_X10Y8_BM_SRAM2
port 1628 nsew signal output
flabel metal2 s 452544 338648 452640 338728 0 FreeSans 320 0 0 0 Tile_X10Y8_BM_SRAM20
port 1629 nsew signal output
flabel metal2 s 452544 339152 452640 339232 0 FreeSans 320 0 0 0 Tile_X10Y8_BM_SRAM21
port 1630 nsew signal output
flabel metal2 s 452544 339656 452640 339736 0 FreeSans 320 0 0 0 Tile_X10Y8_BM_SRAM22
port 1631 nsew signal output
flabel metal2 s 452544 340160 452640 340240 0 FreeSans 320 0 0 0 Tile_X10Y8_BM_SRAM23
port 1632 nsew signal output
flabel metal2 s 452544 340664 452640 340744 0 FreeSans 320 0 0 0 Tile_X10Y8_BM_SRAM24
port 1633 nsew signal output
flabel metal2 s 452544 341168 452640 341248 0 FreeSans 320 0 0 0 Tile_X10Y8_BM_SRAM25
port 1634 nsew signal output
flabel metal2 s 452544 341672 452640 341752 0 FreeSans 320 0 0 0 Tile_X10Y8_BM_SRAM26
port 1635 nsew signal output
flabel metal2 s 452544 342176 452640 342256 0 FreeSans 320 0 0 0 Tile_X10Y8_BM_SRAM27
port 1636 nsew signal output
flabel metal2 s 452544 342680 452640 342760 0 FreeSans 320 0 0 0 Tile_X10Y8_BM_SRAM28
port 1637 nsew signal output
flabel metal2 s 452544 343184 452640 343264 0 FreeSans 320 0 0 0 Tile_X10Y8_BM_SRAM29
port 1638 nsew signal output
flabel metal2 s 452544 330080 452640 330160 0 FreeSans 320 0 0 0 Tile_X10Y8_BM_SRAM3
port 1639 nsew signal output
flabel metal2 s 452544 343688 452640 343768 0 FreeSans 320 0 0 0 Tile_X10Y8_BM_SRAM30
port 1640 nsew signal output
flabel metal2 s 452544 344192 452640 344272 0 FreeSans 320 0 0 0 Tile_X10Y8_BM_SRAM31
port 1641 nsew signal output
flabel metal2 s 452544 330584 452640 330664 0 FreeSans 320 0 0 0 Tile_X10Y8_BM_SRAM4
port 1642 nsew signal output
flabel metal2 s 452544 331088 452640 331168 0 FreeSans 320 0 0 0 Tile_X10Y8_BM_SRAM5
port 1643 nsew signal output
flabel metal2 s 452544 331592 452640 331672 0 FreeSans 320 0 0 0 Tile_X10Y8_BM_SRAM6
port 1644 nsew signal output
flabel metal2 s 452544 332096 452640 332176 0 FreeSans 320 0 0 0 Tile_X10Y8_BM_SRAM7
port 1645 nsew signal output
flabel metal2 s 452544 332600 452640 332680 0 FreeSans 320 0 0 0 Tile_X10Y8_BM_SRAM8
port 1646 nsew signal output
flabel metal2 s 452544 333104 452640 333184 0 FreeSans 320 0 0 0 Tile_X10Y8_BM_SRAM9
port 1647 nsew signal output
flabel metal2 s 452544 344696 452640 344776 0 FreeSans 320 0 0 0 Tile_X10Y8_CLK_SRAM
port 1648 nsew signal output
flabel metal2 s 452544 306896 452640 306976 0 FreeSans 320 0 0 0 Tile_X10Y8_CONFIGURED_top
port 1649 nsew signal input
flabel metal2 s 452544 345200 452640 345280 0 FreeSans 320 0 0 0 Tile_X10Y8_DIN_SRAM0
port 1650 nsew signal output
flabel metal2 s 452544 345704 452640 345784 0 FreeSans 320 0 0 0 Tile_X10Y8_DIN_SRAM1
port 1651 nsew signal output
flabel metal2 s 452544 350240 452640 350320 0 FreeSans 320 0 0 0 Tile_X10Y8_DIN_SRAM10
port 1652 nsew signal output
flabel metal2 s 452544 350744 452640 350824 0 FreeSans 320 0 0 0 Tile_X10Y8_DIN_SRAM11
port 1653 nsew signal output
flabel metal2 s 452544 351248 452640 351328 0 FreeSans 320 0 0 0 Tile_X10Y8_DIN_SRAM12
port 1654 nsew signal output
flabel metal2 s 452544 351752 452640 351832 0 FreeSans 320 0 0 0 Tile_X10Y8_DIN_SRAM13
port 1655 nsew signal output
flabel metal2 s 452544 352256 452640 352336 0 FreeSans 320 0 0 0 Tile_X10Y8_DIN_SRAM14
port 1656 nsew signal output
flabel metal2 s 452544 352760 452640 352840 0 FreeSans 320 0 0 0 Tile_X10Y8_DIN_SRAM15
port 1657 nsew signal output
flabel metal2 s 452544 353264 452640 353344 0 FreeSans 320 0 0 0 Tile_X10Y8_DIN_SRAM16
port 1658 nsew signal output
flabel metal2 s 452544 353768 452640 353848 0 FreeSans 320 0 0 0 Tile_X10Y8_DIN_SRAM17
port 1659 nsew signal output
flabel metal2 s 452544 354272 452640 354352 0 FreeSans 320 0 0 0 Tile_X10Y8_DIN_SRAM18
port 1660 nsew signal output
flabel metal2 s 452544 354776 452640 354856 0 FreeSans 320 0 0 0 Tile_X10Y8_DIN_SRAM19
port 1661 nsew signal output
flabel metal2 s 452544 346208 452640 346288 0 FreeSans 320 0 0 0 Tile_X10Y8_DIN_SRAM2
port 1662 nsew signal output
flabel metal2 s 452544 355280 452640 355360 0 FreeSans 320 0 0 0 Tile_X10Y8_DIN_SRAM20
port 1663 nsew signal output
flabel metal2 s 452544 355784 452640 355864 0 FreeSans 320 0 0 0 Tile_X10Y8_DIN_SRAM21
port 1664 nsew signal output
flabel metal2 s 452544 356288 452640 356368 0 FreeSans 320 0 0 0 Tile_X10Y8_DIN_SRAM22
port 1665 nsew signal output
flabel metal2 s 452544 356792 452640 356872 0 FreeSans 320 0 0 0 Tile_X10Y8_DIN_SRAM23
port 1666 nsew signal output
flabel metal2 s 452544 357296 452640 357376 0 FreeSans 320 0 0 0 Tile_X10Y8_DIN_SRAM24
port 1667 nsew signal output
flabel metal2 s 452544 357800 452640 357880 0 FreeSans 320 0 0 0 Tile_X10Y8_DIN_SRAM25
port 1668 nsew signal output
flabel metal2 s 452544 358304 452640 358384 0 FreeSans 320 0 0 0 Tile_X10Y8_DIN_SRAM26
port 1669 nsew signal output
flabel metal2 s 452544 358808 452640 358888 0 FreeSans 320 0 0 0 Tile_X10Y8_DIN_SRAM27
port 1670 nsew signal output
flabel metal2 s 452544 359312 452640 359392 0 FreeSans 320 0 0 0 Tile_X10Y8_DIN_SRAM28
port 1671 nsew signal output
flabel metal2 s 452544 359816 452640 359896 0 FreeSans 320 0 0 0 Tile_X10Y8_DIN_SRAM29
port 1672 nsew signal output
flabel metal2 s 452544 346712 452640 346792 0 FreeSans 320 0 0 0 Tile_X10Y8_DIN_SRAM3
port 1673 nsew signal output
flabel metal2 s 452544 360320 452640 360400 0 FreeSans 320 0 0 0 Tile_X10Y8_DIN_SRAM30
port 1674 nsew signal output
flabel metal2 s 452544 360824 452640 360904 0 FreeSans 320 0 0 0 Tile_X10Y8_DIN_SRAM31
port 1675 nsew signal output
flabel metal2 s 452544 347216 452640 347296 0 FreeSans 320 0 0 0 Tile_X10Y8_DIN_SRAM4
port 1676 nsew signal output
flabel metal2 s 452544 347720 452640 347800 0 FreeSans 320 0 0 0 Tile_X10Y8_DIN_SRAM5
port 1677 nsew signal output
flabel metal2 s 452544 348224 452640 348304 0 FreeSans 320 0 0 0 Tile_X10Y8_DIN_SRAM6
port 1678 nsew signal output
flabel metal2 s 452544 348728 452640 348808 0 FreeSans 320 0 0 0 Tile_X10Y8_DIN_SRAM7
port 1679 nsew signal output
flabel metal2 s 452544 349232 452640 349312 0 FreeSans 320 0 0 0 Tile_X10Y8_DIN_SRAM8
port 1680 nsew signal output
flabel metal2 s 452544 349736 452640 349816 0 FreeSans 320 0 0 0 Tile_X10Y8_DIN_SRAM9
port 1681 nsew signal output
flabel metal2 s 452544 307400 452640 307480 0 FreeSans 320 0 0 0 Tile_X10Y8_DOUT_SRAM0
port 1682 nsew signal input
flabel metal2 s 452544 307904 452640 307984 0 FreeSans 320 0 0 0 Tile_X10Y8_DOUT_SRAM1
port 1683 nsew signal input
flabel metal2 s 452544 312440 452640 312520 0 FreeSans 320 0 0 0 Tile_X10Y8_DOUT_SRAM10
port 1684 nsew signal input
flabel metal2 s 452544 312944 452640 313024 0 FreeSans 320 0 0 0 Tile_X10Y8_DOUT_SRAM11
port 1685 nsew signal input
flabel metal2 s 452544 313448 452640 313528 0 FreeSans 320 0 0 0 Tile_X10Y8_DOUT_SRAM12
port 1686 nsew signal input
flabel metal2 s 452544 313952 452640 314032 0 FreeSans 320 0 0 0 Tile_X10Y8_DOUT_SRAM13
port 1687 nsew signal input
flabel metal2 s 452544 314456 452640 314536 0 FreeSans 320 0 0 0 Tile_X10Y8_DOUT_SRAM14
port 1688 nsew signal input
flabel metal2 s 452544 314960 452640 315040 0 FreeSans 320 0 0 0 Tile_X10Y8_DOUT_SRAM15
port 1689 nsew signal input
flabel metal2 s 452544 315464 452640 315544 0 FreeSans 320 0 0 0 Tile_X10Y8_DOUT_SRAM16
port 1690 nsew signal input
flabel metal2 s 452544 315968 452640 316048 0 FreeSans 320 0 0 0 Tile_X10Y8_DOUT_SRAM17
port 1691 nsew signal input
flabel metal2 s 452544 316472 452640 316552 0 FreeSans 320 0 0 0 Tile_X10Y8_DOUT_SRAM18
port 1692 nsew signal input
flabel metal2 s 452544 316976 452640 317056 0 FreeSans 320 0 0 0 Tile_X10Y8_DOUT_SRAM19
port 1693 nsew signal input
flabel metal2 s 452544 308408 452640 308488 0 FreeSans 320 0 0 0 Tile_X10Y8_DOUT_SRAM2
port 1694 nsew signal input
flabel metal2 s 452544 317480 452640 317560 0 FreeSans 320 0 0 0 Tile_X10Y8_DOUT_SRAM20
port 1695 nsew signal input
flabel metal2 s 452544 317984 452640 318064 0 FreeSans 320 0 0 0 Tile_X10Y8_DOUT_SRAM21
port 1696 nsew signal input
flabel metal2 s 452544 318488 452640 318568 0 FreeSans 320 0 0 0 Tile_X10Y8_DOUT_SRAM22
port 1697 nsew signal input
flabel metal2 s 452544 318992 452640 319072 0 FreeSans 320 0 0 0 Tile_X10Y8_DOUT_SRAM23
port 1698 nsew signal input
flabel metal2 s 452544 319496 452640 319576 0 FreeSans 320 0 0 0 Tile_X10Y8_DOUT_SRAM24
port 1699 nsew signal input
flabel metal2 s 452544 320000 452640 320080 0 FreeSans 320 0 0 0 Tile_X10Y8_DOUT_SRAM25
port 1700 nsew signal input
flabel metal2 s 452544 320504 452640 320584 0 FreeSans 320 0 0 0 Tile_X10Y8_DOUT_SRAM26
port 1701 nsew signal input
flabel metal2 s 452544 321008 452640 321088 0 FreeSans 320 0 0 0 Tile_X10Y8_DOUT_SRAM27
port 1702 nsew signal input
flabel metal2 s 452544 321512 452640 321592 0 FreeSans 320 0 0 0 Tile_X10Y8_DOUT_SRAM28
port 1703 nsew signal input
flabel metal2 s 452544 322016 452640 322096 0 FreeSans 320 0 0 0 Tile_X10Y8_DOUT_SRAM29
port 1704 nsew signal input
flabel metal2 s 452544 308912 452640 308992 0 FreeSans 320 0 0 0 Tile_X10Y8_DOUT_SRAM3
port 1705 nsew signal input
flabel metal2 s 452544 322520 452640 322600 0 FreeSans 320 0 0 0 Tile_X10Y8_DOUT_SRAM30
port 1706 nsew signal input
flabel metal2 s 452544 323024 452640 323104 0 FreeSans 320 0 0 0 Tile_X10Y8_DOUT_SRAM31
port 1707 nsew signal input
flabel metal2 s 452544 309416 452640 309496 0 FreeSans 320 0 0 0 Tile_X10Y8_DOUT_SRAM4
port 1708 nsew signal input
flabel metal2 s 452544 309920 452640 310000 0 FreeSans 320 0 0 0 Tile_X10Y8_DOUT_SRAM5
port 1709 nsew signal input
flabel metal2 s 452544 310424 452640 310504 0 FreeSans 320 0 0 0 Tile_X10Y8_DOUT_SRAM6
port 1710 nsew signal input
flabel metal2 s 452544 310928 452640 311008 0 FreeSans 320 0 0 0 Tile_X10Y8_DOUT_SRAM7
port 1711 nsew signal input
flabel metal2 s 452544 311432 452640 311512 0 FreeSans 320 0 0 0 Tile_X10Y8_DOUT_SRAM8
port 1712 nsew signal input
flabel metal2 s 452544 311936 452640 312016 0 FreeSans 320 0 0 0 Tile_X10Y8_DOUT_SRAM9
port 1713 nsew signal input
flabel metal2 s 452544 361328 452640 361408 0 FreeSans 320 0 0 0 Tile_X10Y8_MEN_SRAM
port 1714 nsew signal output
flabel metal2 s 452544 361832 452640 361912 0 FreeSans 320 0 0 0 Tile_X10Y8_REN_SRAM
port 1715 nsew signal output
flabel metal2 s 452544 362336 452640 362416 0 FreeSans 320 0 0 0 Tile_X10Y8_TIE_HIGH_SRAM
port 1716 nsew signal output
flabel metal2 s 452544 362840 452640 362920 0 FreeSans 320 0 0 0 Tile_X10Y8_TIE_LOW_SRAM
port 1717 nsew signal output
flabel metal2 s 452544 363344 452640 363424 0 FreeSans 320 0 0 0 Tile_X10Y8_WEN_SRAM
port 1718 nsew signal output
flabel metal3 s 18488 702240 18568 702336 0 FreeSans 640 0 0 0 Tile_X1Y0_A_I_top
port 1719 nsew signal output
flabel metal3 s 17336 702240 17416 702336 0 FreeSans 640 0 0 0 Tile_X1Y0_A_O_top
port 1720 nsew signal input
flabel metal3 s 19640 702240 19720 702336 0 FreeSans 640 0 0 0 Tile_X1Y0_A_T_top
port 1721 nsew signal output
flabel metal3 s 24248 702240 24328 702336 0 FreeSans 640 0 0 0 Tile_X1Y0_A_config_C_bit0
port 1722 nsew signal output
flabel metal3 s 25400 702240 25480 702336 0 FreeSans 640 0 0 0 Tile_X1Y0_A_config_C_bit1
port 1723 nsew signal output
flabel metal3 s 26552 702240 26632 702336 0 FreeSans 640 0 0 0 Tile_X1Y0_A_config_C_bit2
port 1724 nsew signal output
flabel metal3 s 27704 702240 27784 702336 0 FreeSans 640 0 0 0 Tile_X1Y0_A_config_C_bit3
port 1725 nsew signal output
flabel metal3 s 21944 702240 22024 702336 0 FreeSans 640 0 0 0 Tile_X1Y0_B_I_top
port 1726 nsew signal output
flabel metal3 s 20792 702240 20872 702336 0 FreeSans 640 0 0 0 Tile_X1Y0_B_O_top
port 1727 nsew signal input
flabel metal3 s 23096 702240 23176 702336 0 FreeSans 640 0 0 0 Tile_X1Y0_B_T_top
port 1728 nsew signal output
flabel metal3 s 28856 702240 28936 702336 0 FreeSans 640 0 0 0 Tile_X1Y0_B_config_C_bit0
port 1729 nsew signal output
flabel metal3 s 30008 702240 30088 702336 0 FreeSans 640 0 0 0 Tile_X1Y0_B_config_C_bit1
port 1730 nsew signal output
flabel metal3 s 31160 702240 31240 702336 0 FreeSans 640 0 0 0 Tile_X1Y0_B_config_C_bit2
port 1731 nsew signal output
flabel metal3 s 32312 702240 32392 702336 0 FreeSans 640 0 0 0 Tile_X1Y0_B_config_C_bit3
port 1732 nsew signal output
flabel metal3 s 64856 702240 64936 702336 0 FreeSans 640 0 0 0 Tile_X2Y0_A_I_top
port 1733 nsew signal output
flabel metal3 s 63704 702240 63784 702336 0 FreeSans 640 0 0 0 Tile_X2Y0_A_O_top
port 1734 nsew signal input
flabel metal3 s 66008 702240 66088 702336 0 FreeSans 640 0 0 0 Tile_X2Y0_A_T_top
port 1735 nsew signal output
flabel metal3 s 70616 702240 70696 702336 0 FreeSans 640 0 0 0 Tile_X2Y0_A_config_C_bit0
port 1736 nsew signal output
flabel metal3 s 71768 702240 71848 702336 0 FreeSans 640 0 0 0 Tile_X2Y0_A_config_C_bit1
port 1737 nsew signal output
flabel metal3 s 72920 702240 73000 702336 0 FreeSans 640 0 0 0 Tile_X2Y0_A_config_C_bit2
port 1738 nsew signal output
flabel metal3 s 74072 702240 74152 702336 0 FreeSans 640 0 0 0 Tile_X2Y0_A_config_C_bit3
port 1739 nsew signal output
flabel metal3 s 68312 702240 68392 702336 0 FreeSans 640 0 0 0 Tile_X2Y0_B_I_top
port 1740 nsew signal output
flabel metal3 s 67160 702240 67240 702336 0 FreeSans 640 0 0 0 Tile_X2Y0_B_O_top
port 1741 nsew signal input
flabel metal3 s 69464 702240 69544 702336 0 FreeSans 640 0 0 0 Tile_X2Y0_B_T_top
port 1742 nsew signal output
flabel metal3 s 75224 702240 75304 702336 0 FreeSans 640 0 0 0 Tile_X2Y0_B_config_C_bit0
port 1743 nsew signal output
flabel metal3 s 76376 702240 76456 702336 0 FreeSans 640 0 0 0 Tile_X2Y0_B_config_C_bit1
port 1744 nsew signal output
flabel metal3 s 77528 702240 77608 702336 0 FreeSans 640 0 0 0 Tile_X2Y0_B_config_C_bit2
port 1745 nsew signal output
flabel metal3 s 78680 702240 78760 702336 0 FreeSans 640 0 0 0 Tile_X2Y0_B_config_C_bit3
port 1746 nsew signal output
flabel metal3 s 65624 0 65704 96 0 FreeSans 640 0 0 0 Tile_X2Y15_BOOT_top
port 1747 nsew signal output
flabel metal3 s 62552 0 62632 96 0 FreeSans 640 0 0 0 Tile_X2Y15_CONFIGURED_top
port 1748 nsew signal input
flabel metal3 s 64088 0 64168 96 0 FreeSans 640 0 0 0 Tile_X2Y15_RESET_top
port 1749 nsew signal input
flabel metal3 s 67160 0 67240 96 0 FreeSans 640 0 0 0 Tile_X2Y15_SLOT_top0
port 1750 nsew signal output
flabel metal3 s 68696 0 68776 96 0 FreeSans 640 0 0 0 Tile_X2Y15_SLOT_top1
port 1751 nsew signal output
flabel metal3 s 70232 0 70312 96 0 FreeSans 640 0 0 0 Tile_X2Y15_SLOT_top2
port 1752 nsew signal output
flabel metal3 s 71768 0 71848 96 0 FreeSans 640 0 0 0 Tile_X2Y15_SLOT_top3
port 1753 nsew signal output
flabel metal3 s 107960 0 108040 96 0 FreeSans 640 0 0 0 Tile_X3Y15_CONFIGURED_top
port 1754 nsew signal input
flabel metal3 s 109688 0 109768 96 0 FreeSans 640 0 0 0 Tile_X3Y15_IRQ_top0
port 1755 nsew signal output
flabel metal3 s 111416 0 111496 96 0 FreeSans 640 0 0 0 Tile_X3Y15_IRQ_top1
port 1756 nsew signal output
flabel metal3 s 113144 0 113224 96 0 FreeSans 640 0 0 0 Tile_X3Y15_IRQ_top2
port 1757 nsew signal output
flabel metal3 s 114872 0 114952 96 0 FreeSans 640 0 0 0 Tile_X3Y15_IRQ_top3
port 1758 nsew signal output
flabel metal3 s 221624 0 221704 96 0 FreeSans 640 0 0 0 Tile_X5Y15_I_top0
port 1759 nsew signal output
flabel metal3 s 222392 0 222472 96 0 FreeSans 640 0 0 0 Tile_X5Y15_I_top1
port 1760 nsew signal output
flabel metal3 s 229304 0 229384 96 0 FreeSans 640 0 0 0 Tile_X5Y15_I_top10
port 1761 nsew signal output
flabel metal3 s 230072 0 230152 96 0 FreeSans 640 0 0 0 Tile_X5Y15_I_top11
port 1762 nsew signal output
flabel metal3 s 230840 0 230920 96 0 FreeSans 640 0 0 0 Tile_X5Y15_I_top12
port 1763 nsew signal output
flabel metal3 s 231608 0 231688 96 0 FreeSans 640 0 0 0 Tile_X5Y15_I_top13
port 1764 nsew signal output
flabel metal3 s 232376 0 232456 96 0 FreeSans 640 0 0 0 Tile_X5Y15_I_top14
port 1765 nsew signal output
flabel metal3 s 233144 0 233224 96 0 FreeSans 640 0 0 0 Tile_X5Y15_I_top15
port 1766 nsew signal output
flabel metal3 s 223160 0 223240 96 0 FreeSans 640 0 0 0 Tile_X5Y15_I_top2
port 1767 nsew signal output
flabel metal3 s 223928 0 224008 96 0 FreeSans 640 0 0 0 Tile_X5Y15_I_top3
port 1768 nsew signal output
flabel metal3 s 224696 0 224776 96 0 FreeSans 640 0 0 0 Tile_X5Y15_I_top4
port 1769 nsew signal output
flabel metal3 s 225464 0 225544 96 0 FreeSans 640 0 0 0 Tile_X5Y15_I_top5
port 1770 nsew signal output
flabel metal3 s 226232 0 226312 96 0 FreeSans 640 0 0 0 Tile_X5Y15_I_top6
port 1771 nsew signal output
flabel metal3 s 227000 0 227080 96 0 FreeSans 640 0 0 0 Tile_X5Y15_I_top7
port 1772 nsew signal output
flabel metal3 s 227768 0 227848 96 0 FreeSans 640 0 0 0 Tile_X5Y15_I_top8
port 1773 nsew signal output
flabel metal3 s 228536 0 228616 96 0 FreeSans 640 0 0 0 Tile_X5Y15_I_top9
port 1774 nsew signal output
flabel metal3 s 209336 0 209416 96 0 FreeSans 640 0 0 0 Tile_X5Y15_O_top0
port 1775 nsew signal input
flabel metal3 s 210104 0 210184 96 0 FreeSans 640 0 0 0 Tile_X5Y15_O_top1
port 1776 nsew signal input
flabel metal3 s 217016 0 217096 96 0 FreeSans 640 0 0 0 Tile_X5Y15_O_top10
port 1777 nsew signal input
flabel metal3 s 217784 0 217864 96 0 FreeSans 640 0 0 0 Tile_X5Y15_O_top11
port 1778 nsew signal input
flabel metal3 s 218552 0 218632 96 0 FreeSans 640 0 0 0 Tile_X5Y15_O_top12
port 1779 nsew signal input
flabel metal3 s 219320 0 219400 96 0 FreeSans 640 0 0 0 Tile_X5Y15_O_top13
port 1780 nsew signal input
flabel metal3 s 220088 0 220168 96 0 FreeSans 640 0 0 0 Tile_X5Y15_O_top14
port 1781 nsew signal input
flabel metal3 s 220856 0 220936 96 0 FreeSans 640 0 0 0 Tile_X5Y15_O_top15
port 1782 nsew signal input
flabel metal3 s 210872 0 210952 96 0 FreeSans 640 0 0 0 Tile_X5Y15_O_top2
port 1783 nsew signal input
flabel metal3 s 211640 0 211720 96 0 FreeSans 640 0 0 0 Tile_X5Y15_O_top3
port 1784 nsew signal input
flabel metal3 s 212408 0 212488 96 0 FreeSans 640 0 0 0 Tile_X5Y15_O_top4
port 1785 nsew signal input
flabel metal3 s 213176 0 213256 96 0 FreeSans 640 0 0 0 Tile_X5Y15_O_top5
port 1786 nsew signal input
flabel metal3 s 213944 0 214024 96 0 FreeSans 640 0 0 0 Tile_X5Y15_O_top6
port 1787 nsew signal input
flabel metal3 s 214712 0 214792 96 0 FreeSans 640 0 0 0 Tile_X5Y15_O_top7
port 1788 nsew signal input
flabel metal3 s 215480 0 215560 96 0 FreeSans 640 0 0 0 Tile_X5Y15_O_top8
port 1789 nsew signal input
flabel metal3 s 216248 0 216328 96 0 FreeSans 640 0 0 0 Tile_X5Y15_O_top9
port 1790 nsew signal input
flabel metal3 s 267992 0 268072 96 0 FreeSans 640 0 0 0 Tile_X6Y15_I_top0
port 1791 nsew signal output
flabel metal3 s 268760 0 268840 96 0 FreeSans 640 0 0 0 Tile_X6Y15_I_top1
port 1792 nsew signal output
flabel metal3 s 275672 0 275752 96 0 FreeSans 640 0 0 0 Tile_X6Y15_I_top10
port 1793 nsew signal output
flabel metal3 s 276440 0 276520 96 0 FreeSans 640 0 0 0 Tile_X6Y15_I_top11
port 1794 nsew signal output
flabel metal3 s 277208 0 277288 96 0 FreeSans 640 0 0 0 Tile_X6Y15_I_top12
port 1795 nsew signal output
flabel metal3 s 277976 0 278056 96 0 FreeSans 640 0 0 0 Tile_X6Y15_I_top13
port 1796 nsew signal output
flabel metal3 s 278744 0 278824 96 0 FreeSans 640 0 0 0 Tile_X6Y15_I_top14
port 1797 nsew signal output
flabel metal3 s 279512 0 279592 96 0 FreeSans 640 0 0 0 Tile_X6Y15_I_top15
port 1798 nsew signal output
flabel metal3 s 269528 0 269608 96 0 FreeSans 640 0 0 0 Tile_X6Y15_I_top2
port 1799 nsew signal output
flabel metal3 s 270296 0 270376 96 0 FreeSans 640 0 0 0 Tile_X6Y15_I_top3
port 1800 nsew signal output
flabel metal3 s 271064 0 271144 96 0 FreeSans 640 0 0 0 Tile_X6Y15_I_top4
port 1801 nsew signal output
flabel metal3 s 271832 0 271912 96 0 FreeSans 640 0 0 0 Tile_X6Y15_I_top5
port 1802 nsew signal output
flabel metal3 s 272600 0 272680 96 0 FreeSans 640 0 0 0 Tile_X6Y15_I_top6
port 1803 nsew signal output
flabel metal3 s 273368 0 273448 96 0 FreeSans 640 0 0 0 Tile_X6Y15_I_top7
port 1804 nsew signal output
flabel metal3 s 274136 0 274216 96 0 FreeSans 640 0 0 0 Tile_X6Y15_I_top8
port 1805 nsew signal output
flabel metal3 s 274904 0 274984 96 0 FreeSans 640 0 0 0 Tile_X6Y15_I_top9
port 1806 nsew signal output
flabel metal3 s 255704 0 255784 96 0 FreeSans 640 0 0 0 Tile_X6Y15_O_top0
port 1807 nsew signal input
flabel metal3 s 256472 0 256552 96 0 FreeSans 640 0 0 0 Tile_X6Y15_O_top1
port 1808 nsew signal input
flabel metal3 s 263384 0 263464 96 0 FreeSans 640 0 0 0 Tile_X6Y15_O_top10
port 1809 nsew signal input
flabel metal3 s 264152 0 264232 96 0 FreeSans 640 0 0 0 Tile_X6Y15_O_top11
port 1810 nsew signal input
flabel metal3 s 264920 0 265000 96 0 FreeSans 640 0 0 0 Tile_X6Y15_O_top12
port 1811 nsew signal input
flabel metal3 s 265688 0 265768 96 0 FreeSans 640 0 0 0 Tile_X6Y15_O_top13
port 1812 nsew signal input
flabel metal3 s 266456 0 266536 96 0 FreeSans 640 0 0 0 Tile_X6Y15_O_top14
port 1813 nsew signal input
flabel metal3 s 267224 0 267304 96 0 FreeSans 640 0 0 0 Tile_X6Y15_O_top15
port 1814 nsew signal input
flabel metal3 s 257240 0 257320 96 0 FreeSans 640 0 0 0 Tile_X6Y15_O_top2
port 1815 nsew signal input
flabel metal3 s 258008 0 258088 96 0 FreeSans 640 0 0 0 Tile_X6Y15_O_top3
port 1816 nsew signal input
flabel metal3 s 258776 0 258856 96 0 FreeSans 640 0 0 0 Tile_X6Y15_O_top4
port 1817 nsew signal input
flabel metal3 s 259544 0 259624 96 0 FreeSans 640 0 0 0 Tile_X6Y15_O_top5
port 1818 nsew signal input
flabel metal3 s 260312 0 260392 96 0 FreeSans 640 0 0 0 Tile_X6Y15_O_top6
port 1819 nsew signal input
flabel metal3 s 261080 0 261160 96 0 FreeSans 640 0 0 0 Tile_X6Y15_O_top7
port 1820 nsew signal input
flabel metal3 s 261848 0 261928 96 0 FreeSans 640 0 0 0 Tile_X6Y15_O_top8
port 1821 nsew signal input
flabel metal3 s 262616 0 262696 96 0 FreeSans 640 0 0 0 Tile_X6Y15_O_top9
port 1822 nsew signal input
flabel metal3 s 353624 0 353704 96 0 FreeSans 640 0 0 0 Tile_X8Y15_I_top0
port 1823 nsew signal output
flabel metal3 s 354392 0 354472 96 0 FreeSans 640 0 0 0 Tile_X8Y15_I_top1
port 1824 nsew signal output
flabel metal3 s 361304 0 361384 96 0 FreeSans 640 0 0 0 Tile_X8Y15_I_top10
port 1825 nsew signal output
flabel metal3 s 362072 0 362152 96 0 FreeSans 640 0 0 0 Tile_X8Y15_I_top11
port 1826 nsew signal output
flabel metal3 s 362840 0 362920 96 0 FreeSans 640 0 0 0 Tile_X8Y15_I_top12
port 1827 nsew signal output
flabel metal3 s 363608 0 363688 96 0 FreeSans 640 0 0 0 Tile_X8Y15_I_top13
port 1828 nsew signal output
flabel metal3 s 364376 0 364456 96 0 FreeSans 640 0 0 0 Tile_X8Y15_I_top14
port 1829 nsew signal output
flabel metal3 s 365144 0 365224 96 0 FreeSans 640 0 0 0 Tile_X8Y15_I_top15
port 1830 nsew signal output
flabel metal3 s 355160 0 355240 96 0 FreeSans 640 0 0 0 Tile_X8Y15_I_top2
port 1831 nsew signal output
flabel metal3 s 355928 0 356008 96 0 FreeSans 640 0 0 0 Tile_X8Y15_I_top3
port 1832 nsew signal output
flabel metal3 s 356696 0 356776 96 0 FreeSans 640 0 0 0 Tile_X8Y15_I_top4
port 1833 nsew signal output
flabel metal3 s 357464 0 357544 96 0 FreeSans 640 0 0 0 Tile_X8Y15_I_top5
port 1834 nsew signal output
flabel metal3 s 358232 0 358312 96 0 FreeSans 640 0 0 0 Tile_X8Y15_I_top6
port 1835 nsew signal output
flabel metal3 s 359000 0 359080 96 0 FreeSans 640 0 0 0 Tile_X8Y15_I_top7
port 1836 nsew signal output
flabel metal3 s 359768 0 359848 96 0 FreeSans 640 0 0 0 Tile_X8Y15_I_top8
port 1837 nsew signal output
flabel metal3 s 360536 0 360616 96 0 FreeSans 640 0 0 0 Tile_X8Y15_I_top9
port 1838 nsew signal output
flabel metal3 s 341336 0 341416 96 0 FreeSans 640 0 0 0 Tile_X8Y15_O_top0
port 1839 nsew signal input
flabel metal3 s 342104 0 342184 96 0 FreeSans 640 0 0 0 Tile_X8Y15_O_top1
port 1840 nsew signal input
flabel metal3 s 349016 0 349096 96 0 FreeSans 640 0 0 0 Tile_X8Y15_O_top10
port 1841 nsew signal input
flabel metal3 s 349784 0 349864 96 0 FreeSans 640 0 0 0 Tile_X8Y15_O_top11
port 1842 nsew signal input
flabel metal3 s 350552 0 350632 96 0 FreeSans 640 0 0 0 Tile_X8Y15_O_top12
port 1843 nsew signal input
flabel metal3 s 351320 0 351400 96 0 FreeSans 640 0 0 0 Tile_X8Y15_O_top13
port 1844 nsew signal input
flabel metal3 s 352088 0 352168 96 0 FreeSans 640 0 0 0 Tile_X8Y15_O_top14
port 1845 nsew signal input
flabel metal3 s 352856 0 352936 96 0 FreeSans 640 0 0 0 Tile_X8Y15_O_top15
port 1846 nsew signal input
flabel metal3 s 342872 0 342952 96 0 FreeSans 640 0 0 0 Tile_X8Y15_O_top2
port 1847 nsew signal input
flabel metal3 s 343640 0 343720 96 0 FreeSans 640 0 0 0 Tile_X8Y15_O_top3
port 1848 nsew signal input
flabel metal3 s 344408 0 344488 96 0 FreeSans 640 0 0 0 Tile_X8Y15_O_top4
port 1849 nsew signal input
flabel metal3 s 345176 0 345256 96 0 FreeSans 640 0 0 0 Tile_X8Y15_O_top5
port 1850 nsew signal input
flabel metal3 s 345944 0 346024 96 0 FreeSans 640 0 0 0 Tile_X8Y15_O_top6
port 1851 nsew signal input
flabel metal3 s 346712 0 346792 96 0 FreeSans 640 0 0 0 Tile_X8Y15_O_top7
port 1852 nsew signal input
flabel metal3 s 347480 0 347560 96 0 FreeSans 640 0 0 0 Tile_X8Y15_O_top8
port 1853 nsew signal input
flabel metal3 s 348248 0 348328 96 0 FreeSans 640 0 0 0 Tile_X8Y15_O_top9
port 1854 nsew signal input
flabel metal3 s 399992 0 400072 96 0 FreeSans 640 0 0 0 Tile_X9Y15_I_top0
port 1855 nsew signal output
flabel metal3 s 400760 0 400840 96 0 FreeSans 640 0 0 0 Tile_X9Y15_I_top1
port 1856 nsew signal output
flabel metal3 s 407672 0 407752 96 0 FreeSans 640 0 0 0 Tile_X9Y15_I_top10
port 1857 nsew signal output
flabel metal3 s 408440 0 408520 96 0 FreeSans 640 0 0 0 Tile_X9Y15_I_top11
port 1858 nsew signal output
flabel metal3 s 409208 0 409288 96 0 FreeSans 640 0 0 0 Tile_X9Y15_I_top12
port 1859 nsew signal output
flabel metal3 s 409976 0 410056 96 0 FreeSans 640 0 0 0 Tile_X9Y15_I_top13
port 1860 nsew signal output
flabel metal3 s 410744 0 410824 96 0 FreeSans 640 0 0 0 Tile_X9Y15_I_top14
port 1861 nsew signal output
flabel metal3 s 411512 0 411592 96 0 FreeSans 640 0 0 0 Tile_X9Y15_I_top15
port 1862 nsew signal output
flabel metal3 s 401528 0 401608 96 0 FreeSans 640 0 0 0 Tile_X9Y15_I_top2
port 1863 nsew signal output
flabel metal3 s 402296 0 402376 96 0 FreeSans 640 0 0 0 Tile_X9Y15_I_top3
port 1864 nsew signal output
flabel metal3 s 403064 0 403144 96 0 FreeSans 640 0 0 0 Tile_X9Y15_I_top4
port 1865 nsew signal output
flabel metal3 s 403832 0 403912 96 0 FreeSans 640 0 0 0 Tile_X9Y15_I_top5
port 1866 nsew signal output
flabel metal3 s 404600 0 404680 96 0 FreeSans 640 0 0 0 Tile_X9Y15_I_top6
port 1867 nsew signal output
flabel metal3 s 405368 0 405448 96 0 FreeSans 640 0 0 0 Tile_X9Y15_I_top7
port 1868 nsew signal output
flabel metal3 s 406136 0 406216 96 0 FreeSans 640 0 0 0 Tile_X9Y15_I_top8
port 1869 nsew signal output
flabel metal3 s 406904 0 406984 96 0 FreeSans 640 0 0 0 Tile_X9Y15_I_top9
port 1870 nsew signal output
flabel metal3 s 387704 0 387784 96 0 FreeSans 640 0 0 0 Tile_X9Y15_O_top0
port 1871 nsew signal input
flabel metal3 s 388472 0 388552 96 0 FreeSans 640 0 0 0 Tile_X9Y15_O_top1
port 1872 nsew signal input
flabel metal3 s 395384 0 395464 96 0 FreeSans 640 0 0 0 Tile_X9Y15_O_top10
port 1873 nsew signal input
flabel metal3 s 396152 0 396232 96 0 FreeSans 640 0 0 0 Tile_X9Y15_O_top11
port 1874 nsew signal input
flabel metal3 s 396920 0 397000 96 0 FreeSans 640 0 0 0 Tile_X9Y15_O_top12
port 1875 nsew signal input
flabel metal3 s 397688 0 397768 96 0 FreeSans 640 0 0 0 Tile_X9Y15_O_top13
port 1876 nsew signal input
flabel metal3 s 398456 0 398536 96 0 FreeSans 640 0 0 0 Tile_X9Y15_O_top14
port 1877 nsew signal input
flabel metal3 s 399224 0 399304 96 0 FreeSans 640 0 0 0 Tile_X9Y15_O_top15
port 1878 nsew signal input
flabel metal3 s 389240 0 389320 96 0 FreeSans 640 0 0 0 Tile_X9Y15_O_top2
port 1879 nsew signal input
flabel metal3 s 390008 0 390088 96 0 FreeSans 640 0 0 0 Tile_X9Y15_O_top3
port 1880 nsew signal input
flabel metal3 s 390776 0 390856 96 0 FreeSans 640 0 0 0 Tile_X9Y15_O_top4
port 1881 nsew signal input
flabel metal3 s 391544 0 391624 96 0 FreeSans 640 0 0 0 Tile_X9Y15_O_top5
port 1882 nsew signal input
flabel metal3 s 392312 0 392392 96 0 FreeSans 640 0 0 0 Tile_X9Y15_O_top6
port 1883 nsew signal input
flabel metal3 s 393080 0 393160 96 0 FreeSans 640 0 0 0 Tile_X9Y15_O_top7
port 1884 nsew signal input
flabel metal3 s 393848 0 393928 96 0 FreeSans 640 0 0 0 Tile_X9Y15_O_top8
port 1885 nsew signal input
flabel metal3 s 394616 0 394696 96 0 FreeSans 640 0 0 0 Tile_X9Y15_O_top9
port 1886 nsew signal input
flabel metal3 s 1112 0 1192 80 0 FreeSans 320 0 0 0 UserCLK
port 1887 nsew signal input
flabel metal5 s 4988 840 5428 702240 0 FreeSans 2560 90 0 0 VGND
port 1888 nsew ground bidirectional
flabel metal5 s 18716 840 19156 702240 0 FreeSans 2560 90 0 0 VGND
port 1888 nsew ground bidirectional
flabel metal5 s 33836 840 34276 702240 0 FreeSans 2560 90 0 0 VGND
port 1888 nsew ground bidirectional
flabel metal5 s 48956 840 49396 702240 0 FreeSans 2560 90 0 0 VGND
port 1888 nsew ground bidirectional
flabel metal5 s 65084 840 65524 702240 0 FreeSans 2560 90 0 0 VGND
port 1888 nsew ground bidirectional
flabel metal5 s 80204 840 80644 702240 0 FreeSans 2560 90 0 0 VGND
port 1888 nsew ground bidirectional
flabel metal5 s 95324 840 95764 702240 0 FreeSans 2560 90 0 0 VGND
port 1888 nsew ground bidirectional
flabel metal5 s 111452 840 111892 702240 0 FreeSans 2560 90 0 0 VGND
port 1888 nsew ground bidirectional
flabel metal5 s 126572 840 127012 702240 0 FreeSans 2560 90 0 0 VGND
port 1888 nsew ground bidirectional
flabel metal5 s 141692 840 142132 702240 0 FreeSans 2560 90 0 0 VGND
port 1888 nsew ground bidirectional
flabel metal5 s 157820 840 158260 702240 0 FreeSans 2560 90 0 0 VGND
port 1888 nsew ground bidirectional
flabel metal5 s 172940 840 173380 702240 0 FreeSans 2560 90 0 0 VGND
port 1888 nsew ground bidirectional
flabel metal5 s 188060 840 188500 702240 0 FreeSans 2560 90 0 0 VGND
port 1888 nsew ground bidirectional
flabel metal5 s 203180 840 203620 702240 0 FreeSans 2560 90 0 0 VGND
port 1888 nsew ground bidirectional
flabel metal5 s 211100 840 211540 702240 0 FreeSans 2560 90 0 0 VGND
port 1888 nsew ground bidirectional
flabel metal5 s 226220 840 226660 702240 0 FreeSans 2560 90 0 0 VGND
port 1888 nsew ground bidirectional
flabel metal5 s 241340 840 241780 702240 0 FreeSans 2560 90 0 0 VGND
port 1888 nsew ground bidirectional
flabel metal5 s 257468 840 257908 702240 0 FreeSans 2560 90 0 0 VGND
port 1888 nsew ground bidirectional
flabel metal5 s 272588 840 273028 702240 0 FreeSans 2560 90 0 0 VGND
port 1888 nsew ground bidirectional
flabel metal5 s 287708 840 288148 702240 0 FreeSans 2560 90 0 0 VGND
port 1888 nsew ground bidirectional
flabel metal5 s 303836 840 304276 702240 0 FreeSans 2560 90 0 0 VGND
port 1888 nsew ground bidirectional
flabel metal5 s 318956 840 319396 702240 0 FreeSans 2560 90 0 0 VGND
port 1888 nsew ground bidirectional
flabel metal5 s 334076 840 334516 702240 0 FreeSans 2560 90 0 0 VGND
port 1888 nsew ground bidirectional
flabel metal5 s 343100 840 343540 702240 0 FreeSans 2560 90 0 0 VGND
port 1888 nsew ground bidirectional
flabel metal5 s 358220 840 358660 702240 0 FreeSans 2560 90 0 0 VGND
port 1888 nsew ground bidirectional
flabel metal5 s 373340 840 373780 702240 0 FreeSans 2560 90 0 0 VGND
port 1888 nsew ground bidirectional
flabel metal5 s 389468 840 389908 702240 0 FreeSans 2560 90 0 0 VGND
port 1888 nsew ground bidirectional
flabel metal5 s 404588 840 405028 702240 0 FreeSans 2560 90 0 0 VGND
port 1888 nsew ground bidirectional
flabel metal5 s 419708 840 420148 702240 0 FreeSans 2560 90 0 0 VGND
port 1888 nsew ground bidirectional
flabel metal5 s 435836 840 436276 702240 0 FreeSans 2560 90 0 0 VGND
port 1888 nsew ground bidirectional
flabel metal5 s 3748 840 4188 702240 0 FreeSans 2560 90 0 0 VPWR
port 1889 nsew power bidirectional
flabel metal5 s 17476 840 17916 702240 0 FreeSans 2560 90 0 0 VPWR
port 1889 nsew power bidirectional
flabel metal5 s 32596 840 33036 702240 0 FreeSans 2560 90 0 0 VPWR
port 1889 nsew power bidirectional
flabel metal5 s 47716 840 48156 702240 0 FreeSans 2560 90 0 0 VPWR
port 1889 nsew power bidirectional
flabel metal5 s 63844 840 64284 702240 0 FreeSans 2560 90 0 0 VPWR
port 1889 nsew power bidirectional
flabel metal5 s 78964 840 79404 702240 0 FreeSans 2560 90 0 0 VPWR
port 1889 nsew power bidirectional
flabel metal5 s 94084 840 94524 702240 0 FreeSans 2560 90 0 0 VPWR
port 1889 nsew power bidirectional
flabel metal5 s 110212 840 110652 702240 0 FreeSans 2560 90 0 0 VPWR
port 1889 nsew power bidirectional
flabel metal5 s 125332 840 125772 702240 0 FreeSans 2560 90 0 0 VPWR
port 1889 nsew power bidirectional
flabel metal5 s 140452 840 140892 702240 0 FreeSans 2560 90 0 0 VPWR
port 1889 nsew power bidirectional
flabel metal5 s 156580 840 157020 702240 0 FreeSans 2560 90 0 0 VPWR
port 1889 nsew power bidirectional
flabel metal5 s 171700 840 172140 702240 0 FreeSans 2560 90 0 0 VPWR
port 1889 nsew power bidirectional
flabel metal5 s 186820 840 187260 702240 0 FreeSans 2560 90 0 0 VPWR
port 1889 nsew power bidirectional
flabel metal5 s 201940 840 202380 702240 0 FreeSans 2560 90 0 0 VPWR
port 1889 nsew power bidirectional
flabel metal5 s 209860 840 210300 702240 0 FreeSans 2560 90 0 0 VPWR
port 1889 nsew power bidirectional
flabel metal5 s 224980 840 225420 702240 0 FreeSans 2560 90 0 0 VPWR
port 1889 nsew power bidirectional
flabel metal5 s 240100 840 240540 702240 0 FreeSans 2560 90 0 0 VPWR
port 1889 nsew power bidirectional
flabel metal5 s 256228 840 256668 702240 0 FreeSans 2560 90 0 0 VPWR
port 1889 nsew power bidirectional
flabel metal5 s 271348 840 271788 702240 0 FreeSans 2560 90 0 0 VPWR
port 1889 nsew power bidirectional
flabel metal5 s 286468 840 286908 702240 0 FreeSans 2560 90 0 0 VPWR
port 1889 nsew power bidirectional
flabel metal5 s 302596 840 303036 702240 0 FreeSans 2560 90 0 0 VPWR
port 1889 nsew power bidirectional
flabel metal5 s 317716 840 318156 702240 0 FreeSans 2560 90 0 0 VPWR
port 1889 nsew power bidirectional
flabel metal5 s 332836 840 333276 702240 0 FreeSans 2560 90 0 0 VPWR
port 1889 nsew power bidirectional
flabel metal5 s 341860 840 342300 702240 0 FreeSans 2560 90 0 0 VPWR
port 1889 nsew power bidirectional
flabel metal5 s 356980 840 357420 702240 0 FreeSans 2560 90 0 0 VPWR
port 1889 nsew power bidirectional
flabel metal5 s 372100 840 372540 702240 0 FreeSans 2560 90 0 0 VPWR
port 1889 nsew power bidirectional
flabel metal5 s 388228 840 388668 702240 0 FreeSans 2560 90 0 0 VPWR
port 1889 nsew power bidirectional
flabel metal5 s 403348 840 403788 702240 0 FreeSans 2560 90 0 0 VPWR
port 1889 nsew power bidirectional
flabel metal5 s 418468 840 418908 702240 0 FreeSans 2560 90 0 0 VPWR
port 1889 nsew power bidirectional
flabel metal5 s 434596 840 435036 702240 0 FreeSans 2560 90 0 0 VPWR
port 1889 nsew power bidirectional
flabel metal5 s 449716 840 450156 702240 0 FreeSans 2560 90 0 0 VPWR
port 1889 nsew power bidirectional
rlabel metal5 436056 351540 436056 351540 0 VGND
rlabel metal5 449936 351540 449936 351540 0 VPWR
rlabel metal2 6946 690816 6946 690816 0 FrameData[0]
rlabel metal2 82 564480 82 564480 0 FrameData[100]
rlabel metal2 82 565488 82 565488 0 FrameData[101]
rlabel metal2 82 566496 82 566496 0 FrameData[102]
rlabel metal2 82 567504 82 567504 0 FrameData[103]
rlabel metal2 82 568512 82 568512 0 FrameData[104]
rlabel metal2 82 569520 82 569520 0 FrameData[105]
rlabel metal2 82 570528 82 570528 0 FrameData[106]
rlabel metal2 82 571536 82 571536 0 FrameData[107]
rlabel metal2 82 572544 82 572544 0 FrameData[108]
rlabel metal2 82 573552 82 573552 0 FrameData[109]
rlabel metal2 6946 694176 6946 694176 0 FrameData[10]
rlabel metal2 82 574560 82 574560 0 FrameData[110]
rlabel metal2 82 575568 82 575568 0 FrameData[111]
rlabel metal2 82 576576 82 576576 0 FrameData[112]
rlabel metal2 82 577584 82 577584 0 FrameData[113]
rlabel metal2 82 578592 82 578592 0 FrameData[114]
rlabel metal2 82 579600 82 579600 0 FrameData[115]
rlabel metal2 82 580608 82 580608 0 FrameData[116]
rlabel metal2 82 581616 82 581616 0 FrameData[117]
rlabel metal2 82 582624 82 582624 0 FrameData[118]
rlabel metal2 82 583632 82 583632 0 FrameData[119]
rlabel metal2 6946 694512 6946 694512 0 FrameData[11]
rlabel metal2 82 584640 82 584640 0 FrameData[120]
rlabel metal2 82 585648 82 585648 0 FrameData[121]
rlabel metal2 82 586656 82 586656 0 FrameData[122]
rlabel metal2 82 587664 82 587664 0 FrameData[123]
rlabel metal2 82 588672 82 588672 0 FrameData[124]
rlabel metal2 82 589680 82 589680 0 FrameData[125]
rlabel metal2 82 590688 82 590688 0 FrameData[126]
rlabel metal2 82 591696 82 591696 0 FrameData[127]
rlabel metal2 82 512064 82 512064 0 FrameData[128]
rlabel metal2 82 513072 82 513072 0 FrameData[129]
rlabel metal2 6946 694848 6946 694848 0 FrameData[12]
rlabel metal2 82 514080 82 514080 0 FrameData[130]
rlabel metal2 82 515088 82 515088 0 FrameData[131]
rlabel metal2 82 516096 82 516096 0 FrameData[132]
rlabel metal2 82 517104 82 517104 0 FrameData[133]
rlabel metal2 82 518112 82 518112 0 FrameData[134]
rlabel metal2 82 519120 82 519120 0 FrameData[135]
rlabel metal2 82 520128 82 520128 0 FrameData[136]
rlabel metal2 82 521136 82 521136 0 FrameData[137]
rlabel metal2 82 522144 82 522144 0 FrameData[138]
rlabel metal2 82 523152 82 523152 0 FrameData[139]
rlabel metal2 6946 695184 6946 695184 0 FrameData[13]
rlabel metal2 82 524160 82 524160 0 FrameData[140]
rlabel metal2 82 525168 82 525168 0 FrameData[141]
rlabel metal2 82 526176 82 526176 0 FrameData[142]
rlabel metal2 82 527184 82 527184 0 FrameData[143]
rlabel metal2 82 528192 82 528192 0 FrameData[144]
rlabel metal2 82 529200 82 529200 0 FrameData[145]
rlabel metal2 82 530208 82 530208 0 FrameData[146]
rlabel metal2 82 531216 82 531216 0 FrameData[147]
rlabel metal2 82 532224 82 532224 0 FrameData[148]
rlabel metal2 82 533232 82 533232 0 FrameData[149]
rlabel metal2 6946 695520 6946 695520 0 FrameData[14]
rlabel metal2 82 534240 82 534240 0 FrameData[150]
rlabel metal2 82 535248 82 535248 0 FrameData[151]
rlabel metal2 82 536256 82 536256 0 FrameData[152]
rlabel metal2 82 537264 82 537264 0 FrameData[153]
rlabel metal2 82 538272 82 538272 0 FrameData[154]
rlabel metal2 82 539280 82 539280 0 FrameData[155]
rlabel metal2 82 540288 82 540288 0 FrameData[156]
rlabel metal2 82 541296 82 541296 0 FrameData[157]
rlabel metal2 82 542304 82 542304 0 FrameData[158]
rlabel metal2 82 543312 82 543312 0 FrameData[159]
rlabel metal2 6946 695856 6946 695856 0 FrameData[15]
rlabel metal2 82 463680 82 463680 0 FrameData[160]
rlabel metal2 82 464688 82 464688 0 FrameData[161]
rlabel metal2 82 465696 82 465696 0 FrameData[162]
rlabel metal2 82 466704 82 466704 0 FrameData[163]
rlabel metal2 82 467712 82 467712 0 FrameData[164]
rlabel metal2 82 468720 82 468720 0 FrameData[165]
rlabel metal2 82 469728 82 469728 0 FrameData[166]
rlabel metal2 82 470736 82 470736 0 FrameData[167]
rlabel metal2 82 471744 82 471744 0 FrameData[168]
rlabel metal2 82 472752 82 472752 0 FrameData[169]
rlabel metal2 6946 696192 6946 696192 0 FrameData[16]
rlabel metal2 82 473760 82 473760 0 FrameData[170]
rlabel metal2 82 474768 82 474768 0 FrameData[171]
rlabel metal2 82 475776 82 475776 0 FrameData[172]
rlabel metal2 82 476784 82 476784 0 FrameData[173]
rlabel metal2 82 477792 82 477792 0 FrameData[174]
rlabel metal2 82 478800 82 478800 0 FrameData[175]
rlabel metal2 82 479808 82 479808 0 FrameData[176]
rlabel metal2 82 480816 82 480816 0 FrameData[177]
rlabel metal2 82 481824 82 481824 0 FrameData[178]
rlabel metal2 82 482832 82 482832 0 FrameData[179]
rlabel metal2 6946 696528 6946 696528 0 FrameData[17]
rlabel metal2 82 483840 82 483840 0 FrameData[180]
rlabel metal2 82 484848 82 484848 0 FrameData[181]
rlabel metal2 82 485856 82 485856 0 FrameData[182]
rlabel metal2 82 486864 82 486864 0 FrameData[183]
rlabel metal2 82 487872 82 487872 0 FrameData[184]
rlabel metal2 82 488880 82 488880 0 FrameData[185]
rlabel metal2 82 489888 82 489888 0 FrameData[186]
rlabel metal2 82 490896 82 490896 0 FrameData[187]
rlabel metal2 82 491904 82 491904 0 FrameData[188]
rlabel metal2 82 492912 82 492912 0 FrameData[189]
rlabel metal2 6946 696864 6946 696864 0 FrameData[18]
rlabel metal2 82 493920 82 493920 0 FrameData[190]
rlabel metal2 82 494928 82 494928 0 FrameData[191]
rlabel metal2 82 415296 82 415296 0 FrameData[192]
rlabel metal2 82 416304 82 416304 0 FrameData[193]
rlabel metal2 82 417312 82 417312 0 FrameData[194]
rlabel metal2 82 418320 82 418320 0 FrameData[195]
rlabel metal2 82 419328 82 419328 0 FrameData[196]
rlabel metal2 82 420336 82 420336 0 FrameData[197]
rlabel metal2 82 421344 82 421344 0 FrameData[198]
rlabel metal2 82 422352 82 422352 0 FrameData[199]
rlabel metal2 6946 697200 6946 697200 0 FrameData[19]
rlabel metal2 6946 691152 6946 691152 0 FrameData[1]
rlabel metal2 82 423360 82 423360 0 FrameData[200]
rlabel metal2 82 424368 82 424368 0 FrameData[201]
rlabel metal2 82 425376 82 425376 0 FrameData[202]
rlabel metal2 82 426384 82 426384 0 FrameData[203]
rlabel metal2 82 427392 82 427392 0 FrameData[204]
rlabel metal2 82 428400 82 428400 0 FrameData[205]
rlabel metal2 82 429408 82 429408 0 FrameData[206]
rlabel metal2 82 430416 82 430416 0 FrameData[207]
rlabel metal2 82 431424 82 431424 0 FrameData[208]
rlabel metal2 82 432432 82 432432 0 FrameData[209]
rlabel metal2 6946 697536 6946 697536 0 FrameData[20]
rlabel metal2 82 433440 82 433440 0 FrameData[210]
rlabel metal2 82 434448 82 434448 0 FrameData[211]
rlabel metal2 82 435456 82 435456 0 FrameData[212]
rlabel metal2 82 436464 82 436464 0 FrameData[213]
rlabel metal2 82 437472 82 437472 0 FrameData[214]
rlabel metal2 82 438480 82 438480 0 FrameData[215]
rlabel metal2 82 439488 82 439488 0 FrameData[216]
rlabel metal2 82 440496 82 440496 0 FrameData[217]
rlabel metal2 82 441504 82 441504 0 FrameData[218]
rlabel metal2 82 442512 82 442512 0 FrameData[219]
rlabel metal2 6946 697872 6946 697872 0 FrameData[21]
rlabel metal2 82 443520 82 443520 0 FrameData[220]
rlabel metal2 82 444528 82 444528 0 FrameData[221]
rlabel metal2 82 445536 82 445536 0 FrameData[222]
rlabel metal2 82 446544 82 446544 0 FrameData[223]
rlabel metal2 82 366912 82 366912 0 FrameData[224]
rlabel metal2 82 367920 82 367920 0 FrameData[225]
rlabel metal2 82 368928 82 368928 0 FrameData[226]
rlabel metal2 82 369936 82 369936 0 FrameData[227]
rlabel metal2 82 370944 82 370944 0 FrameData[228]
rlabel metal2 82 371952 82 371952 0 FrameData[229]
rlabel metal2 6946 698208 6946 698208 0 FrameData[22]
rlabel metal2 82 372960 82 372960 0 FrameData[230]
rlabel metal2 82 373968 82 373968 0 FrameData[231]
rlabel metal2 82 374976 82 374976 0 FrameData[232]
rlabel metal2 82 375984 82 375984 0 FrameData[233]
rlabel metal2 82 376992 82 376992 0 FrameData[234]
rlabel metal2 82 378000 82 378000 0 FrameData[235]
rlabel metal2 82 379008 82 379008 0 FrameData[236]
rlabel metal2 82 380016 82 380016 0 FrameData[237]
rlabel metal2 82 381024 82 381024 0 FrameData[238]
rlabel metal2 82 382032 82 382032 0 FrameData[239]
rlabel metal2 6946 698544 6946 698544 0 FrameData[23]
rlabel metal2 82 383040 82 383040 0 FrameData[240]
rlabel metal2 82 384048 82 384048 0 FrameData[241]
rlabel metal2 82 385056 82 385056 0 FrameData[242]
rlabel metal2 82 386064 82 386064 0 FrameData[243]
rlabel metal2 82 387072 82 387072 0 FrameData[244]
rlabel metal2 82 388080 82 388080 0 FrameData[245]
rlabel metal2 82 389088 82 389088 0 FrameData[246]
rlabel metal2 82 390096 82 390096 0 FrameData[247]
rlabel metal2 82 391104 82 391104 0 FrameData[248]
rlabel metal2 82 392112 82 392112 0 FrameData[249]
rlabel metal2 6946 698880 6946 698880 0 FrameData[24]
rlabel metal2 82 393120 82 393120 0 FrameData[250]
rlabel metal2 82 394128 82 394128 0 FrameData[251]
rlabel metal2 82 395136 82 395136 0 FrameData[252]
rlabel metal2 82 396144 82 396144 0 FrameData[253]
rlabel metal2 82 397152 82 397152 0 FrameData[254]
rlabel metal2 82 398160 82 398160 0 FrameData[255]
rlabel metal2 82 318528 82 318528 0 FrameData[256]
rlabel metal2 82 319536 82 319536 0 FrameData[257]
rlabel metal2 82 320544 82 320544 0 FrameData[258]
rlabel metal2 82 321552 82 321552 0 FrameData[259]
rlabel metal2 6946 699216 6946 699216 0 FrameData[25]
rlabel metal2 82 322560 82 322560 0 FrameData[260]
rlabel metal2 82 323568 82 323568 0 FrameData[261]
rlabel metal2 82 324576 82 324576 0 FrameData[262]
rlabel metal2 82 325584 82 325584 0 FrameData[263]
rlabel metal2 82 326592 82 326592 0 FrameData[264]
rlabel metal2 82 327600 82 327600 0 FrameData[265]
rlabel metal2 82 328608 82 328608 0 FrameData[266]
rlabel metal2 82 329616 82 329616 0 FrameData[267]
rlabel metal2 82 330624 82 330624 0 FrameData[268]
rlabel metal2 82 331632 82 331632 0 FrameData[269]
rlabel metal2 6946 699552 6946 699552 0 FrameData[26]
rlabel metal2 82 332640 82 332640 0 FrameData[270]
rlabel metal2 82 333648 82 333648 0 FrameData[271]
rlabel metal2 82 334656 82 334656 0 FrameData[272]
rlabel metal2 82 335664 82 335664 0 FrameData[273]
rlabel metal2 82 336672 82 336672 0 FrameData[274]
rlabel metal2 82 337680 82 337680 0 FrameData[275]
rlabel metal2 82 338688 82 338688 0 FrameData[276]
rlabel metal2 82 339696 82 339696 0 FrameData[277]
rlabel metal2 82 340704 82 340704 0 FrameData[278]
rlabel metal2 82 341712 82 341712 0 FrameData[279]
rlabel metal2 6946 699888 6946 699888 0 FrameData[27]
rlabel metal2 82 342720 82 342720 0 FrameData[280]
rlabel metal2 82 343728 82 343728 0 FrameData[281]
rlabel metal2 82 344736 82 344736 0 FrameData[282]
rlabel metal2 82 345744 82 345744 0 FrameData[283]
rlabel metal2 82 346752 82 346752 0 FrameData[284]
rlabel metal2 82 347760 82 347760 0 FrameData[285]
rlabel metal2 82 348768 82 348768 0 FrameData[286]
rlabel metal2 82 349776 82 349776 0 FrameData[287]
rlabel metal2 82 270144 82 270144 0 FrameData[288]
rlabel metal2 82 271152 82 271152 0 FrameData[289]
rlabel metal2 6946 700224 6946 700224 0 FrameData[28]
rlabel metal2 82 272160 82 272160 0 FrameData[290]
rlabel metal2 82 273168 82 273168 0 FrameData[291]
rlabel metal2 82 274176 82 274176 0 FrameData[292]
rlabel metal2 82 275184 82 275184 0 FrameData[293]
rlabel metal2 82 276192 82 276192 0 FrameData[294]
rlabel metal2 82 277200 82 277200 0 FrameData[295]
rlabel metal2 82 278208 82 278208 0 FrameData[296]
rlabel metal2 82 279216 82 279216 0 FrameData[297]
rlabel metal2 82 280224 82 280224 0 FrameData[298]
rlabel metal2 82 281232 82 281232 0 FrameData[299]
rlabel metal2 6946 700560 6946 700560 0 FrameData[29]
rlabel metal2 6946 691488 6946 691488 0 FrameData[2]
rlabel metal2 82 282240 82 282240 0 FrameData[300]
rlabel metal2 82 283248 82 283248 0 FrameData[301]
rlabel metal2 82 284256 82 284256 0 FrameData[302]
rlabel metal2 82 285264 82 285264 0 FrameData[303]
rlabel metal2 82 286272 82 286272 0 FrameData[304]
rlabel metal2 82 287280 82 287280 0 FrameData[305]
rlabel metal2 82 288288 82 288288 0 FrameData[306]
rlabel metal2 82 289296 82 289296 0 FrameData[307]
rlabel metal2 82 290304 82 290304 0 FrameData[308]
rlabel metal2 82 291312 82 291312 0 FrameData[309]
rlabel metal2 6946 700896 6946 700896 0 FrameData[30]
rlabel metal2 82 292320 82 292320 0 FrameData[310]
rlabel metal2 82 293328 82 293328 0 FrameData[311]
rlabel metal2 82 294336 82 294336 0 FrameData[312]
rlabel metal2 82 295344 82 295344 0 FrameData[313]
rlabel metal2 82 296352 82 296352 0 FrameData[314]
rlabel metal2 82 297360 82 297360 0 FrameData[315]
rlabel metal2 82 298368 82 298368 0 FrameData[316]
rlabel metal2 82 299376 82 299376 0 FrameData[317]
rlabel metal2 82 300384 82 300384 0 FrameData[318]
rlabel metal2 82 301392 82 301392 0 FrameData[319]
rlabel metal2 6946 701232 6946 701232 0 FrameData[31]
rlabel metal2 82 221760 82 221760 0 FrameData[320]
rlabel metal2 82 222768 82 222768 0 FrameData[321]
rlabel metal2 82 223776 82 223776 0 FrameData[322]
rlabel metal2 82 224784 82 224784 0 FrameData[323]
rlabel metal2 82 225792 82 225792 0 FrameData[324]
rlabel metal2 82 226800 82 226800 0 FrameData[325]
rlabel metal2 82 227808 82 227808 0 FrameData[326]
rlabel metal2 82 228816 82 228816 0 FrameData[327]
rlabel metal2 82 229824 82 229824 0 FrameData[328]
rlabel metal2 82 230832 82 230832 0 FrameData[329]
rlabel metal2 82 657216 82 657216 0 FrameData[32]
rlabel metal2 82 231840 82 231840 0 FrameData[330]
rlabel metal2 82 232848 82 232848 0 FrameData[331]
rlabel metal2 82 233856 82 233856 0 FrameData[332]
rlabel metal2 82 234864 82 234864 0 FrameData[333]
rlabel metal2 82 235872 82 235872 0 FrameData[334]
rlabel metal2 82 236880 82 236880 0 FrameData[335]
rlabel metal2 82 237888 82 237888 0 FrameData[336]
rlabel metal2 82 238896 82 238896 0 FrameData[337]
rlabel metal2 82 239904 82 239904 0 FrameData[338]
rlabel metal2 82 240912 82 240912 0 FrameData[339]
rlabel metal2 82 658224 82 658224 0 FrameData[33]
rlabel metal2 82 241920 82 241920 0 FrameData[340]
rlabel metal2 82 242928 82 242928 0 FrameData[341]
rlabel metal2 82 243936 82 243936 0 FrameData[342]
rlabel metal2 82 244944 82 244944 0 FrameData[343]
rlabel metal2 82 245952 82 245952 0 FrameData[344]
rlabel metal2 82 246960 82 246960 0 FrameData[345]
rlabel metal2 82 247968 82 247968 0 FrameData[346]
rlabel metal2 82 248976 82 248976 0 FrameData[347]
rlabel metal2 82 249984 82 249984 0 FrameData[348]
rlabel metal2 82 250992 82 250992 0 FrameData[349]
rlabel metal2 82 659232 82 659232 0 FrameData[34]
rlabel metal2 82 252000 82 252000 0 FrameData[350]
rlabel metal2 82 253008 82 253008 0 FrameData[351]
rlabel metal2 82 173376 82 173376 0 FrameData[352]
rlabel metal2 82 174384 82 174384 0 FrameData[353]
rlabel metal2 82 175392 82 175392 0 FrameData[354]
rlabel metal2 82 176400 82 176400 0 FrameData[355]
rlabel metal2 82 177408 82 177408 0 FrameData[356]
rlabel metal2 82 178416 82 178416 0 FrameData[357]
rlabel metal2 82 179424 82 179424 0 FrameData[358]
rlabel metal2 82 180432 82 180432 0 FrameData[359]
rlabel metal2 82 660240 82 660240 0 FrameData[35]
rlabel metal2 82 181440 82 181440 0 FrameData[360]
rlabel metal2 82 182448 82 182448 0 FrameData[361]
rlabel metal2 82 183456 82 183456 0 FrameData[362]
rlabel metal2 82 184464 82 184464 0 FrameData[363]
rlabel metal2 82 185472 82 185472 0 FrameData[364]
rlabel metal2 82 186480 82 186480 0 FrameData[365]
rlabel metal2 82 187488 82 187488 0 FrameData[366]
rlabel metal2 82 188496 82 188496 0 FrameData[367]
rlabel metal2 82 189504 82 189504 0 FrameData[368]
rlabel metal2 82 190512 82 190512 0 FrameData[369]
rlabel metal2 82 661248 82 661248 0 FrameData[36]
rlabel metal2 82 191520 82 191520 0 FrameData[370]
rlabel metal2 82 192528 82 192528 0 FrameData[371]
rlabel metal2 82 193536 82 193536 0 FrameData[372]
rlabel metal2 82 194544 82 194544 0 FrameData[373]
rlabel metal2 82 195552 82 195552 0 FrameData[374]
rlabel metal2 82 196560 82 196560 0 FrameData[375]
rlabel metal2 82 197568 82 197568 0 FrameData[376]
rlabel metal2 82 198576 82 198576 0 FrameData[377]
rlabel metal2 82 199584 82 199584 0 FrameData[378]
rlabel metal2 82 200592 82 200592 0 FrameData[379]
rlabel metal2 82 662256 82 662256 0 FrameData[37]
rlabel metal2 82 201600 82 201600 0 FrameData[380]
rlabel metal2 82 202608 82 202608 0 FrameData[381]
rlabel metal2 82 203616 82 203616 0 FrameData[382]
rlabel metal2 82 204624 82 204624 0 FrameData[383]
rlabel metal2 82 124992 82 124992 0 FrameData[384]
rlabel metal2 82 126000 82 126000 0 FrameData[385]
rlabel metal2 82 127008 82 127008 0 FrameData[386]
rlabel metal2 82 128016 82 128016 0 FrameData[387]
rlabel metal2 82 129024 82 129024 0 FrameData[388]
rlabel metal2 82 130032 82 130032 0 FrameData[389]
rlabel metal2 82 663264 82 663264 0 FrameData[38]
rlabel metal2 82 131040 82 131040 0 FrameData[390]
rlabel metal2 82 132048 82 132048 0 FrameData[391]
rlabel metal2 82 133056 82 133056 0 FrameData[392]
rlabel metal2 82 134064 82 134064 0 FrameData[393]
rlabel metal2 82 135072 82 135072 0 FrameData[394]
rlabel metal2 82 136080 82 136080 0 FrameData[395]
rlabel metal2 82 137088 82 137088 0 FrameData[396]
rlabel metal2 82 138096 82 138096 0 FrameData[397]
rlabel metal2 82 139104 82 139104 0 FrameData[398]
rlabel metal2 82 140112 82 140112 0 FrameData[399]
rlabel metal2 82 664272 82 664272 0 FrameData[39]
rlabel metal2 6946 691824 6946 691824 0 FrameData[3]
rlabel metal2 82 141120 82 141120 0 FrameData[400]
rlabel metal2 82 142128 82 142128 0 FrameData[401]
rlabel metal2 82 143136 82 143136 0 FrameData[402]
rlabel metal2 82 144144 82 144144 0 FrameData[403]
rlabel metal2 82 145152 82 145152 0 FrameData[404]
rlabel metal2 82 146160 82 146160 0 FrameData[405]
rlabel metal2 82 147168 82 147168 0 FrameData[406]
rlabel metal2 82 148176 82 148176 0 FrameData[407]
rlabel metal2 82 149184 82 149184 0 FrameData[408]
rlabel metal2 82 150192 82 150192 0 FrameData[409]
rlabel metal2 82 665280 82 665280 0 FrameData[40]
rlabel metal2 82 151200 82 151200 0 FrameData[410]
rlabel metal2 82 152208 82 152208 0 FrameData[411]
rlabel metal2 82 153216 82 153216 0 FrameData[412]
rlabel metal2 82 154224 82 154224 0 FrameData[413]
rlabel metal2 82 155232 82 155232 0 FrameData[414]
rlabel metal2 82 156240 82 156240 0 FrameData[415]
rlabel metal2 82 76608 82 76608 0 FrameData[416]
rlabel metal2 82 77616 82 77616 0 FrameData[417]
rlabel metal2 82 78624 82 78624 0 FrameData[418]
rlabel metal2 82 79632 82 79632 0 FrameData[419]
rlabel metal2 82 666288 82 666288 0 FrameData[41]
rlabel metal2 82 80640 82 80640 0 FrameData[420]
rlabel metal2 82 81648 82 81648 0 FrameData[421]
rlabel metal2 82 82656 82 82656 0 FrameData[422]
rlabel metal2 82 83664 82 83664 0 FrameData[423]
rlabel metal2 82 84672 82 84672 0 FrameData[424]
rlabel metal2 82 85680 82 85680 0 FrameData[425]
rlabel metal2 82 86688 82 86688 0 FrameData[426]
rlabel metal2 82 87696 82 87696 0 FrameData[427]
rlabel metal2 82 88704 82 88704 0 FrameData[428]
rlabel metal2 82 89712 82 89712 0 FrameData[429]
rlabel metal2 82 667296 82 667296 0 FrameData[42]
rlabel metal2 82 90720 82 90720 0 FrameData[430]
rlabel metal2 82 91728 82 91728 0 FrameData[431]
rlabel metal2 82 92736 82 92736 0 FrameData[432]
rlabel metal2 82 93744 82 93744 0 FrameData[433]
rlabel metal2 82 94752 82 94752 0 FrameData[434]
rlabel metal2 82 95760 82 95760 0 FrameData[435]
rlabel metal2 82 96768 82 96768 0 FrameData[436]
rlabel metal2 82 97776 82 97776 0 FrameData[437]
rlabel metal2 82 98784 82 98784 0 FrameData[438]
rlabel metal2 82 99792 82 99792 0 FrameData[439]
rlabel metal2 82 668304 82 668304 0 FrameData[43]
rlabel metal2 82 100800 82 100800 0 FrameData[440]
rlabel metal2 82 101808 82 101808 0 FrameData[441]
rlabel metal2 82 102816 82 102816 0 FrameData[442]
rlabel metal2 82 103824 82 103824 0 FrameData[443]
rlabel metal2 82 104832 82 104832 0 FrameData[444]
rlabel metal2 82 105840 82 105840 0 FrameData[445]
rlabel metal2 82 106848 82 106848 0 FrameData[446]
rlabel metal2 82 107856 82 107856 0 FrameData[447]
rlabel metal2 82 28224 82 28224 0 FrameData[448]
rlabel metal2 82 29232 82 29232 0 FrameData[449]
rlabel metal2 82 669312 82 669312 0 FrameData[44]
rlabel metal2 82 30240 82 30240 0 FrameData[450]
rlabel metal2 82 31248 82 31248 0 FrameData[451]
rlabel metal2 82 32256 82 32256 0 FrameData[452]
rlabel metal2 82 33264 82 33264 0 FrameData[453]
rlabel metal2 82 34272 82 34272 0 FrameData[454]
rlabel metal2 82 35280 82 35280 0 FrameData[455]
rlabel metal2 82 36288 82 36288 0 FrameData[456]
rlabel metal2 82 37296 82 37296 0 FrameData[457]
rlabel metal2 82 38304 82 38304 0 FrameData[458]
rlabel metal2 82 39312 82 39312 0 FrameData[459]
rlabel metal2 82 670320 82 670320 0 FrameData[45]
rlabel metal2 82 40320 82 40320 0 FrameData[460]
rlabel metal2 82 41328 82 41328 0 FrameData[461]
rlabel metal2 82 42336 82 42336 0 FrameData[462]
rlabel metal2 82 43344 82 43344 0 FrameData[463]
rlabel metal2 82 44352 82 44352 0 FrameData[464]
rlabel metal2 82 45360 82 45360 0 FrameData[465]
rlabel metal2 82 46368 82 46368 0 FrameData[466]
rlabel metal2 82 47376 82 47376 0 FrameData[467]
rlabel metal2 82 48384 82 48384 0 FrameData[468]
rlabel metal2 82 49392 82 49392 0 FrameData[469]
rlabel metal2 82 671328 82 671328 0 FrameData[46]
rlabel metal2 82 50400 82 50400 0 FrameData[470]
rlabel metal2 82 51408 82 51408 0 FrameData[471]
rlabel metal2 82 52416 82 52416 0 FrameData[472]
rlabel metal2 82 53424 82 53424 0 FrameData[473]
rlabel metal2 82 54432 82 54432 0 FrameData[474]
rlabel metal2 82 55440 82 55440 0 FrameData[475]
rlabel metal2 82 56448 82 56448 0 FrameData[476]
rlabel metal2 82 57456 82 57456 0 FrameData[477]
rlabel metal2 82 58464 82 58464 0 FrameData[478]
rlabel metal2 82 59472 82 59472 0 FrameData[479]
rlabel metal2 82 672336 82 672336 0 FrameData[47]
rlabel metal2 6946 1428 6946 1428 0 FrameData[480]
rlabel metal2 6946 1764 6946 1764 0 FrameData[481]
rlabel metal2 6946 2100 6946 2100 0 FrameData[482]
rlabel metal2 6946 2436 6946 2436 0 FrameData[483]
rlabel metal2 6946 2772 6946 2772 0 FrameData[484]
rlabel metal2 6946 3108 6946 3108 0 FrameData[485]
rlabel metal2 6946 3444 6946 3444 0 FrameData[486]
rlabel metal2 6946 3780 6946 3780 0 FrameData[487]
rlabel metal2 6946 4116 6946 4116 0 FrameData[488]
rlabel metal2 6946 4452 6946 4452 0 FrameData[489]
rlabel metal2 82 673344 82 673344 0 FrameData[48]
rlabel metal2 6946 4788 6946 4788 0 FrameData[490]
rlabel metal2 6946 5124 6946 5124 0 FrameData[491]
rlabel metal2 6946 5460 6946 5460 0 FrameData[492]
rlabel metal2 6946 5796 6946 5796 0 FrameData[493]
rlabel metal2 6946 6132 6946 6132 0 FrameData[494]
rlabel metal2 6946 6468 6946 6468 0 FrameData[495]
rlabel metal2 6946 6804 6946 6804 0 FrameData[496]
rlabel metal2 6946 7140 6946 7140 0 FrameData[497]
rlabel metal2 6946 7476 6946 7476 0 FrameData[498]
rlabel metal2 6946 7812 6946 7812 0 FrameData[499]
rlabel metal2 82 674352 82 674352 0 FrameData[49]
rlabel metal2 6946 692160 6946 692160 0 FrameData[4]
rlabel metal2 6946 8148 6946 8148 0 FrameData[500]
rlabel metal2 6946 8484 6946 8484 0 FrameData[501]
rlabel metal2 6946 8820 6946 8820 0 FrameData[502]
rlabel metal2 6946 9156 6946 9156 0 FrameData[503]
rlabel metal2 6946 9492 6946 9492 0 FrameData[504]
rlabel metal2 6946 9828 6946 9828 0 FrameData[505]
rlabel metal2 6946 10164 6946 10164 0 FrameData[506]
rlabel metal2 6946 10500 6946 10500 0 FrameData[507]
rlabel metal2 6946 10836 6946 10836 0 FrameData[508]
rlabel metal2 6946 11172 6946 11172 0 FrameData[509]
rlabel metal2 82 675360 82 675360 0 FrameData[50]
rlabel metal2 6946 11508 6946 11508 0 FrameData[510]
rlabel metal2 6946 11844 6946 11844 0 FrameData[511]
rlabel metal2 82 676368 82 676368 0 FrameData[51]
rlabel metal2 82 677376 82 677376 0 FrameData[52]
rlabel metal2 82 678384 82 678384 0 FrameData[53]
rlabel metal2 82 679392 82 679392 0 FrameData[54]
rlabel metal2 82 680400 82 680400 0 FrameData[55]
rlabel metal2 82 681408 82 681408 0 FrameData[56]
rlabel metal2 82 682416 82 682416 0 FrameData[57]
rlabel metal2 82 683424 82 683424 0 FrameData[58]
rlabel metal2 82 684432 82 684432 0 FrameData[59]
rlabel metal2 6946 692496 6946 692496 0 FrameData[5]
rlabel metal2 82 685440 82 685440 0 FrameData[60]
rlabel metal2 82 686448 82 686448 0 FrameData[61]
rlabel metal2 82 687456 82 687456 0 FrameData[62]
rlabel metal2 82 688464 82 688464 0 FrameData[63]
rlabel metal2 82 608832 82 608832 0 FrameData[64]
rlabel metal2 82 609840 82 609840 0 FrameData[65]
rlabel metal2 82 610848 82 610848 0 FrameData[66]
rlabel metal2 82 611856 82 611856 0 FrameData[67]
rlabel metal2 82 612864 82 612864 0 FrameData[68]
rlabel metal2 82 613872 82 613872 0 FrameData[69]
rlabel metal2 6946 692832 6946 692832 0 FrameData[6]
rlabel metal2 82 614880 82 614880 0 FrameData[70]
rlabel metal2 82 615888 82 615888 0 FrameData[71]
rlabel metal2 82 616896 82 616896 0 FrameData[72]
rlabel metal2 82 617904 82 617904 0 FrameData[73]
rlabel metal2 82 618912 82 618912 0 FrameData[74]
rlabel metal2 82 619920 82 619920 0 FrameData[75]
rlabel metal2 82 620928 82 620928 0 FrameData[76]
rlabel metal2 82 621936 82 621936 0 FrameData[77]
rlabel metal2 82 622944 82 622944 0 FrameData[78]
rlabel metal2 82 623952 82 623952 0 FrameData[79]
rlabel metal2 6946 693168 6946 693168 0 FrameData[7]
rlabel metal2 82 624960 82 624960 0 FrameData[80]
rlabel metal2 82 625968 82 625968 0 FrameData[81]
rlabel metal2 82 626976 82 626976 0 FrameData[82]
rlabel metal2 82 627984 82 627984 0 FrameData[83]
rlabel metal2 82 628992 82 628992 0 FrameData[84]
rlabel metal2 82 630000 82 630000 0 FrameData[85]
rlabel metal2 82 631008 82 631008 0 FrameData[86]
rlabel metal2 82 632016 82 632016 0 FrameData[87]
rlabel metal2 82 633024 82 633024 0 FrameData[88]
rlabel metal2 82 634032 82 634032 0 FrameData[89]
rlabel metal2 6946 693504 6946 693504 0 FrameData[8]
rlabel metal2 82 635040 82 635040 0 FrameData[90]
rlabel metal2 82 636048 82 636048 0 FrameData[91]
rlabel metal2 82 637056 82 637056 0 FrameData[92]
rlabel metal2 82 638064 82 638064 0 FrameData[93]
rlabel metal2 82 639072 82 639072 0 FrameData[94]
rlabel metal2 82 640080 82 640080 0 FrameData[95]
rlabel metal2 82 560448 82 560448 0 FrameData[96]
rlabel metal2 82 561456 82 561456 0 FrameData[97]
rlabel metal2 82 562464 82 562464 0 FrameData[98]
rlabel metal2 82 563472 82 563472 0 FrameData[99]
rlabel metal2 6946 693840 6946 693840 0 FrameData[9]
rlabel metal3 1728 6372 1728 6372 0 FrameStrobe[0]
rlabel metal3 234720 454 234720 454 0 FrameStrobe[100]
rlabel metal3 235488 454 235488 454 0 FrameStrobe[101]
rlabel metal3 236256 454 236256 454 0 FrameStrobe[102]
rlabel metal3 237024 454 237024 454 0 FrameStrobe[103]
rlabel metal3 237792 454 237792 454 0 FrameStrobe[104]
rlabel metal3 238560 454 238560 454 0 FrameStrobe[105]
rlabel metal3 239328 454 239328 454 0 FrameStrobe[106]
rlabel metal3 240096 454 240096 454 0 FrameStrobe[107]
rlabel metal3 240864 454 240864 454 0 FrameStrobe[108]
rlabel metal3 241632 454 241632 454 0 FrameStrobe[109]
rlabel metal3 7488 6372 7488 6372 0 FrameStrobe[10]
rlabel metal3 242400 454 242400 454 0 FrameStrobe[110]
rlabel metal3 243168 454 243168 454 0 FrameStrobe[111]
rlabel metal3 243936 454 243936 454 0 FrameStrobe[112]
rlabel metal3 244704 454 244704 454 0 FrameStrobe[113]
rlabel metal3 245472 454 245472 454 0 FrameStrobe[114]
rlabel metal3 246240 454 246240 454 0 FrameStrobe[115]
rlabel metal3 247008 454 247008 454 0 FrameStrobe[116]
rlabel metal3 247776 454 247776 454 0 FrameStrobe[117]
rlabel metal3 248544 454 248544 454 0 FrameStrobe[118]
rlabel metal3 249312 454 249312 454 0 FrameStrobe[119]
rlabel metal3 8064 6372 8064 6372 0 FrameStrobe[11]
rlabel metal3 281088 454 281088 454 0 FrameStrobe[120]
rlabel metal3 281856 454 281856 454 0 FrameStrobe[121]
rlabel metal3 282624 454 282624 454 0 FrameStrobe[122]
rlabel metal3 283392 454 283392 454 0 FrameStrobe[123]
rlabel metal3 284160 454 284160 454 0 FrameStrobe[124]
rlabel metal3 284928 454 284928 454 0 FrameStrobe[125]
rlabel metal3 285696 454 285696 454 0 FrameStrobe[126]
rlabel metal3 286464 454 286464 454 0 FrameStrobe[127]
rlabel metal3 287232 454 287232 454 0 FrameStrobe[128]
rlabel metal3 288000 454 288000 454 0 FrameStrobe[129]
rlabel metal3 8640 6372 8640 6372 0 FrameStrobe[12]
rlabel metal3 288768 454 288768 454 0 FrameStrobe[130]
rlabel metal3 289536 454 289536 454 0 FrameStrobe[131]
rlabel metal3 290304 454 290304 454 0 FrameStrobe[132]
rlabel metal3 291072 454 291072 454 0 FrameStrobe[133]
rlabel metal3 291840 454 291840 454 0 FrameStrobe[134]
rlabel metal3 292608 454 292608 454 0 FrameStrobe[135]
rlabel metal3 293376 454 293376 454 0 FrameStrobe[136]
rlabel metal3 294144 454 294144 454 0 FrameStrobe[137]
rlabel metal3 294912 454 294912 454 0 FrameStrobe[138]
rlabel metal3 295680 454 295680 454 0 FrameStrobe[139]
rlabel metal3 9216 6372 9216 6372 0 FrameStrobe[13]
rlabel metal3 302880 454 302880 454 0 FrameStrobe[140]
rlabel metal3 304608 454 304608 454 0 FrameStrobe[141]
rlabel metal3 306336 454 306336 454 0 FrameStrobe[142]
rlabel metal3 308064 454 308064 454 0 FrameStrobe[143]
rlabel metal3 309792 454 309792 454 0 FrameStrobe[144]
rlabel metal3 311520 454 311520 454 0 FrameStrobe[145]
rlabel metal3 313248 454 313248 454 0 FrameStrobe[146]
rlabel metal3 314976 454 314976 454 0 FrameStrobe[147]
rlabel metal3 316704 454 316704 454 0 FrameStrobe[148]
rlabel metal3 318432 454 318432 454 0 FrameStrobe[149]
rlabel metal3 9792 6372 9792 6372 0 FrameStrobe[14]
rlabel metal3 320160 454 320160 454 0 FrameStrobe[150]
rlabel metal3 321888 454 321888 454 0 FrameStrobe[151]
rlabel metal3 323616 454 323616 454 0 FrameStrobe[152]
rlabel metal3 325344 454 325344 454 0 FrameStrobe[153]
rlabel metal3 327072 454 327072 454 0 FrameStrobe[154]
rlabel metal3 328800 454 328800 454 0 FrameStrobe[155]
rlabel metal3 330528 454 330528 454 0 FrameStrobe[156]
rlabel metal3 332256 454 332256 454 0 FrameStrobe[157]
rlabel metal3 333984 454 333984 454 0 FrameStrobe[158]
rlabel metal3 335712 454 335712 454 0 FrameStrobe[159]
rlabel metal3 10368 6372 10368 6372 0 FrameStrobe[15]
rlabel metal3 366720 454 366720 454 0 FrameStrobe[160]
rlabel metal3 367488 454 367488 454 0 FrameStrobe[161]
rlabel metal3 368256 454 368256 454 0 FrameStrobe[162]
rlabel metal3 369024 454 369024 454 0 FrameStrobe[163]
rlabel metal3 369792 454 369792 454 0 FrameStrobe[164]
rlabel metal3 370560 454 370560 454 0 FrameStrobe[165]
rlabel metal3 371328 454 371328 454 0 FrameStrobe[166]
rlabel metal3 372096 454 372096 454 0 FrameStrobe[167]
rlabel metal3 372864 454 372864 454 0 FrameStrobe[168]
rlabel metal3 373632 454 373632 454 0 FrameStrobe[169]
rlabel metal3 10944 6372 10944 6372 0 FrameStrobe[16]
rlabel metal3 374400 454 374400 454 0 FrameStrobe[170]
rlabel metal3 375168 454 375168 454 0 FrameStrobe[171]
rlabel metal3 375936 454 375936 454 0 FrameStrobe[172]
rlabel metal3 376704 454 376704 454 0 FrameStrobe[173]
rlabel metal3 377472 454 377472 454 0 FrameStrobe[174]
rlabel metal3 378240 454 378240 454 0 FrameStrobe[175]
rlabel metal3 379008 454 379008 454 0 FrameStrobe[176]
rlabel metal3 379776 454 379776 454 0 FrameStrobe[177]
rlabel metal3 380544 454 380544 454 0 FrameStrobe[178]
rlabel metal3 381312 454 381312 454 0 FrameStrobe[179]
rlabel metal3 11520 6372 11520 6372 0 FrameStrobe[17]
rlabel metal3 413088 454 413088 454 0 FrameStrobe[180]
rlabel metal3 413856 454 413856 454 0 FrameStrobe[181]
rlabel metal3 414624 454 414624 454 0 FrameStrobe[182]
rlabel metal3 415392 454 415392 454 0 FrameStrobe[183]
rlabel metal3 416160 454 416160 454 0 FrameStrobe[184]
rlabel metal3 416928 454 416928 454 0 FrameStrobe[185]
rlabel metal3 417696 454 417696 454 0 FrameStrobe[186]
rlabel metal3 418464 454 418464 454 0 FrameStrobe[187]
rlabel metal3 419232 454 419232 454 0 FrameStrobe[188]
rlabel metal3 420000 454 420000 454 0 FrameStrobe[189]
rlabel metal3 12096 6372 12096 6372 0 FrameStrobe[18]
rlabel metal3 420768 454 420768 454 0 FrameStrobe[190]
rlabel metal3 421536 454 421536 454 0 FrameStrobe[191]
rlabel metal3 422304 454 422304 454 0 FrameStrobe[192]
rlabel metal3 423072 454 423072 454 0 FrameStrobe[193]
rlabel metal3 423840 454 423840 454 0 FrameStrobe[194]
rlabel metal3 424608 454 424608 454 0 FrameStrobe[195]
rlabel metal3 425376 454 425376 454 0 FrameStrobe[196]
rlabel metal3 426144 454 426144 454 0 FrameStrobe[197]
rlabel metal3 426912 454 426912 454 0 FrameStrobe[198]
rlabel metal3 427680 454 427680 454 0 FrameStrobe[199]
rlabel metal3 12672 6372 12672 6372 0 FrameStrobe[19]
rlabel metal3 2304 6372 2304 6372 0 FrameStrobe[1]
rlabel metal3 432960 450 432960 450 0 FrameStrobe[200]
rlabel metal3 433920 450 433920 450 0 FrameStrobe[201]
rlabel metal3 434880 450 434880 450 0 FrameStrobe[202]
rlabel metal3 435840 450 435840 450 0 FrameStrobe[203]
rlabel metal3 436800 450 436800 450 0 FrameStrobe[204]
rlabel metal3 437760 450 437760 450 0 FrameStrobe[205]
rlabel metal3 438720 450 438720 450 0 FrameStrobe[206]
rlabel metal3 439680 450 439680 450 0 FrameStrobe[207]
rlabel metal3 440640 450 440640 450 0 FrameStrobe[208]
rlabel metal3 441600 450 441600 450 0 FrameStrobe[209]
rlabel metal3 17952 454 17952 454 0 FrameStrobe[20]
rlabel metal3 442560 450 442560 450 0 FrameStrobe[210]
rlabel metal3 443520 450 443520 450 0 FrameStrobe[211]
rlabel metal3 444480 450 444480 450 0 FrameStrobe[212]
rlabel metal3 445440 450 445440 450 0 FrameStrobe[213]
rlabel metal3 446400 450 446400 450 0 FrameStrobe[214]
rlabel metal3 447360 450 447360 450 0 FrameStrobe[215]
rlabel metal3 448320 450 448320 450 0 FrameStrobe[216]
rlabel metal3 449280 450 449280 450 0 FrameStrobe[217]
rlabel metal3 450240 450 450240 450 0 FrameStrobe[218]
rlabel metal3 451200 450 451200 450 0 FrameStrobe[219]
rlabel metal3 20064 454 20064 454 0 FrameStrobe[21]
rlabel metal3 22176 454 22176 454 0 FrameStrobe[22]
rlabel metal3 24288 454 24288 454 0 FrameStrobe[23]
rlabel metal3 26400 454 26400 454 0 FrameStrobe[24]
rlabel metal3 28512 454 28512 454 0 FrameStrobe[25]
rlabel metal3 30624 454 30624 454 0 FrameStrobe[26]
rlabel metal3 32736 454 32736 454 0 FrameStrobe[27]
rlabel metal3 34848 454 34848 454 0 FrameStrobe[28]
rlabel metal3 36960 454 36960 454 0 FrameStrobe[29]
rlabel metal3 2880 6372 2880 6372 0 FrameStrobe[2]
rlabel metal3 39072 454 39072 454 0 FrameStrobe[30]
rlabel metal3 41184 454 41184 454 0 FrameStrobe[31]
rlabel metal3 43296 454 43296 454 0 FrameStrobe[32]
rlabel metal3 45408 454 45408 454 0 FrameStrobe[33]
rlabel metal3 47520 454 47520 454 0 FrameStrobe[34]
rlabel metal3 49632 454 49632 454 0 FrameStrobe[35]
rlabel metal3 51744 454 51744 454 0 FrameStrobe[36]
rlabel metal3 53856 454 53856 454 0 FrameStrobe[37]
rlabel metal3 55968 454 55968 454 0 FrameStrobe[38]
rlabel metal3 58080 454 58080 454 0 FrameStrobe[39]
rlabel metal3 3456 6372 3456 6372 0 FrameStrobe[3]
rlabel metal3 74880 454 74880 454 0 FrameStrobe[40]
rlabel metal3 76416 454 76416 454 0 FrameStrobe[41]
rlabel metal3 77952 454 77952 454 0 FrameStrobe[42]
rlabel metal3 79488 454 79488 454 0 FrameStrobe[43]
rlabel metal3 81024 454 81024 454 0 FrameStrobe[44]
rlabel metal3 82560 454 82560 454 0 FrameStrobe[45]
rlabel metal3 84096 454 84096 454 0 FrameStrobe[46]
rlabel metal3 85632 454 85632 454 0 FrameStrobe[47]
rlabel metal3 87168 454 87168 454 0 FrameStrobe[48]
rlabel metal3 88704 454 88704 454 0 FrameStrobe[49]
rlabel metal3 4032 6372 4032 6372 0 FrameStrobe[4]
rlabel metal3 90240 454 90240 454 0 FrameStrobe[50]
rlabel metal3 91776 454 91776 454 0 FrameStrobe[51]
rlabel metal3 93312 454 93312 454 0 FrameStrobe[52]
rlabel metal3 94848 454 94848 454 0 FrameStrobe[53]
rlabel metal3 96384 454 96384 454 0 FrameStrobe[54]
rlabel metal3 97920 454 97920 454 0 FrameStrobe[55]
rlabel metal3 99456 454 99456 454 0 FrameStrobe[56]
rlabel metal3 100992 454 100992 454 0 FrameStrobe[57]
rlabel metal3 102528 454 102528 454 0 FrameStrobe[58]
rlabel metal3 104064 454 104064 454 0 FrameStrobe[59]
rlabel metal3 4608 6372 4608 6372 0 FrameStrobe[5]
rlabel metal3 118368 454 118368 454 0 FrameStrobe[60]
rlabel metal3 120096 454 120096 454 0 FrameStrobe[61]
rlabel metal3 121824 454 121824 454 0 FrameStrobe[62]
rlabel metal3 123552 454 123552 454 0 FrameStrobe[63]
rlabel metal3 125280 454 125280 454 0 FrameStrobe[64]
rlabel metal3 127008 454 127008 454 0 FrameStrobe[65]
rlabel metal3 128736 454 128736 454 0 FrameStrobe[66]
rlabel metal3 130464 454 130464 454 0 FrameStrobe[67]
rlabel metal3 132192 454 132192 454 0 FrameStrobe[68]
rlabel metal3 133920 454 133920 454 0 FrameStrobe[69]
rlabel metal3 5184 6372 5184 6372 0 FrameStrobe[6]
rlabel metal3 135648 454 135648 454 0 FrameStrobe[70]
rlabel metal3 137376 454 137376 454 0 FrameStrobe[71]
rlabel metal3 139104 454 139104 454 0 FrameStrobe[72]
rlabel metal3 140832 454 140832 454 0 FrameStrobe[73]
rlabel metal3 142560 454 142560 454 0 FrameStrobe[74]
rlabel metal3 144288 454 144288 454 0 FrameStrobe[75]
rlabel metal3 146016 454 146016 454 0 FrameStrobe[76]
rlabel metal3 147744 454 147744 454 0 FrameStrobe[77]
rlabel metal3 149472 454 149472 454 0 FrameStrobe[78]
rlabel metal3 151200 454 151200 454 0 FrameStrobe[79]
rlabel metal3 5760 6372 5760 6372 0 FrameStrobe[7]
rlabel metal3 157056 454 157056 454 0 FrameStrobe[80]
rlabel metal3 159552 454 159552 454 0 FrameStrobe[81]
rlabel metal3 162048 454 162048 454 0 FrameStrobe[82]
rlabel metal3 164544 454 164544 454 0 FrameStrobe[83]
rlabel metal3 167040 454 167040 454 0 FrameStrobe[84]
rlabel metal3 169536 454 169536 454 0 FrameStrobe[85]
rlabel metal3 172032 454 172032 454 0 FrameStrobe[86]
rlabel metal3 174528 454 174528 454 0 FrameStrobe[87]
rlabel metal3 177024 454 177024 454 0 FrameStrobe[88]
rlabel metal3 179520 454 179520 454 0 FrameStrobe[89]
rlabel metal3 6336 6372 6336 6372 0 FrameStrobe[8]
rlabel metal3 182016 454 182016 454 0 FrameStrobe[90]
rlabel metal3 184512 454 184512 454 0 FrameStrobe[91]
rlabel metal3 187008 454 187008 454 0 FrameStrobe[92]
rlabel metal3 189504 454 189504 454 0 FrameStrobe[93]
rlabel metal3 192000 454 192000 454 0 FrameStrobe[94]
rlabel metal3 194496 454 194496 454 0 FrameStrobe[95]
rlabel metal3 196992 454 196992 454 0 FrameStrobe[96]
rlabel metal3 199488 454 199488 454 0 FrameStrobe[97]
rlabel metal3 201984 454 201984 454 0 FrameStrobe[98]
rlabel metal3 204480 454 204480 454 0 FrameStrobe[99]
rlabel metal3 6912 6372 6912 6372 0 FrameStrobe[9]
rlabel metal2 82 208656 82 208656 0 Tile_X0Y10_A_I_top
rlabel metal2 82 207648 82 207648 0 Tile_X0Y10_A_O_top
rlabel metal2 82 209664 82 209664 0 Tile_X0Y10_A_T_top
rlabel metal2 82 213696 82 213696 0 Tile_X0Y10_A_config_C_bit0
rlabel metal2 82 214704 82 214704 0 Tile_X0Y10_A_config_C_bit1
rlabel metal2 82 215712 82 215712 0 Tile_X0Y10_A_config_C_bit2
rlabel metal2 82 216720 82 216720 0 Tile_X0Y10_A_config_C_bit3
rlabel metal2 82 211680 82 211680 0 Tile_X0Y10_B_I_top
rlabel metal2 82 210672 82 210672 0 Tile_X0Y10_B_O_top
rlabel metal2 82 212688 82 212688 0 Tile_X0Y10_B_T_top
rlabel metal2 82 217728 82 217728 0 Tile_X0Y10_B_config_C_bit0
rlabel metal2 82 218736 82 218736 0 Tile_X0Y10_B_config_C_bit1
rlabel metal2 82 219744 82 219744 0 Tile_X0Y10_B_config_C_bit2
rlabel metal2 82 220752 82 220752 0 Tile_X0Y10_B_config_C_bit3
rlabel metal2 82 160272 82 160272 0 Tile_X0Y11_A_I_top
rlabel metal2 82 159264 82 159264 0 Tile_X0Y11_A_O_top
rlabel metal2 82 161280 82 161280 0 Tile_X0Y11_A_T_top
rlabel metal2 82 165312 82 165312 0 Tile_X0Y11_A_config_C_bit0
rlabel metal2 82 166320 82 166320 0 Tile_X0Y11_A_config_C_bit1
rlabel metal2 82 167328 82 167328 0 Tile_X0Y11_A_config_C_bit2
rlabel metal2 82 168336 82 168336 0 Tile_X0Y11_A_config_C_bit3
rlabel metal2 82 163296 82 163296 0 Tile_X0Y11_B_I_top
rlabel metal2 82 162288 82 162288 0 Tile_X0Y11_B_O_top
rlabel metal2 82 164304 82 164304 0 Tile_X0Y11_B_T_top
rlabel metal2 82 169344 82 169344 0 Tile_X0Y11_B_config_C_bit0
rlabel metal2 82 170352 82 170352 0 Tile_X0Y11_B_config_C_bit1
rlabel metal2 82 171360 82 171360 0 Tile_X0Y11_B_config_C_bit2
rlabel metal2 82 172368 82 172368 0 Tile_X0Y11_B_config_C_bit3
rlabel metal2 82 111888 82 111888 0 Tile_X0Y12_A_I_top
rlabel metal2 82 110880 82 110880 0 Tile_X0Y12_A_O_top
rlabel metal2 82 112896 82 112896 0 Tile_X0Y12_A_T_top
rlabel metal2 82 116928 82 116928 0 Tile_X0Y12_A_config_C_bit0
rlabel metal2 82 117936 82 117936 0 Tile_X0Y12_A_config_C_bit1
rlabel metal2 82 118944 82 118944 0 Tile_X0Y12_A_config_C_bit2
rlabel metal2 82 119952 82 119952 0 Tile_X0Y12_A_config_C_bit3
rlabel metal2 82 114912 82 114912 0 Tile_X0Y12_B_I_top
rlabel metal2 82 113904 82 113904 0 Tile_X0Y12_B_O_top
rlabel metal2 82 115920 82 115920 0 Tile_X0Y12_B_T_top
rlabel metal2 82 120960 82 120960 0 Tile_X0Y12_B_config_C_bit0
rlabel metal2 82 121968 82 121968 0 Tile_X0Y12_B_config_C_bit1
rlabel metal2 82 122976 82 122976 0 Tile_X0Y12_B_config_C_bit2
rlabel metal2 82 123984 82 123984 0 Tile_X0Y12_B_config_C_bit3
rlabel metal2 82 63504 82 63504 0 Tile_X0Y13_A_I_top
rlabel metal2 82 62496 82 62496 0 Tile_X0Y13_A_O_top
rlabel metal2 82 64512 82 64512 0 Tile_X0Y13_A_T_top
rlabel metal2 82 68544 82 68544 0 Tile_X0Y13_A_config_C_bit0
rlabel metal2 82 69552 82 69552 0 Tile_X0Y13_A_config_C_bit1
rlabel metal2 82 70560 82 70560 0 Tile_X0Y13_A_config_C_bit2
rlabel metal2 82 71568 82 71568 0 Tile_X0Y13_A_config_C_bit3
rlabel metal2 82 66528 82 66528 0 Tile_X0Y13_B_I_top
rlabel metal2 82 65520 82 65520 0 Tile_X0Y13_B_O_top
rlabel metal2 82 67536 82 67536 0 Tile_X0Y13_B_T_top
rlabel metal2 82 72576 82 72576 0 Tile_X0Y13_B_config_C_bit0
rlabel metal2 82 73584 82 73584 0 Tile_X0Y13_B_config_C_bit1
rlabel metal2 82 74592 82 74592 0 Tile_X0Y13_B_config_C_bit2
rlabel metal2 82 75600 82 75600 0 Tile_X0Y13_B_config_C_bit3
rlabel metal2 82 15120 82 15120 0 Tile_X0Y14_A_I_top
rlabel metal2 117 13272 117 13272 0 Tile_X0Y14_A_O_top
rlabel metal2 82 16128 82 16128 0 Tile_X0Y14_A_T_top
rlabel metal2 82 20160 82 20160 0 Tile_X0Y14_A_config_C_bit0
rlabel metal2 82 21168 82 21168 0 Tile_X0Y14_A_config_C_bit1
rlabel metal2 82 22176 82 22176 0 Tile_X0Y14_A_config_C_bit2
rlabel metal2 82 23184 82 23184 0 Tile_X0Y14_A_config_C_bit3
rlabel metal2 82 18144 82 18144 0 Tile_X0Y14_B_I_top
rlabel metal2 82 17136 82 17136 0 Tile_X0Y14_B_O_top
rlabel metal2 82 19152 82 19152 0 Tile_X0Y14_B_T_top
rlabel metal2 82 24192 82 24192 0 Tile_X0Y14_B_config_C_bit0
rlabel metal2 82 25200 82 25200 0 Tile_X0Y14_B_config_C_bit1
rlabel metal2 82 26208 82 26208 0 Tile_X0Y14_B_config_C_bit2
rlabel metal2 82 27216 82 27216 0 Tile_X0Y14_B_config_C_bit3
rlabel metal2 82 644112 82 644112 0 Tile_X0Y1_A_I_top
rlabel metal2 82 643104 82 643104 0 Tile_X0Y1_A_O_top
rlabel metal2 82 645120 82 645120 0 Tile_X0Y1_A_T_top
rlabel metal2 82 649152 82 649152 0 Tile_X0Y1_A_config_C_bit0
rlabel metal2 82 650160 82 650160 0 Tile_X0Y1_A_config_C_bit1
rlabel metal2 82 651168 82 651168 0 Tile_X0Y1_A_config_C_bit2
rlabel metal2 82 652176 82 652176 0 Tile_X0Y1_A_config_C_bit3
rlabel metal2 82 647136 82 647136 0 Tile_X0Y1_B_I_top
rlabel metal2 82 646128 82 646128 0 Tile_X0Y1_B_O_top
rlabel metal2 82 648144 82 648144 0 Tile_X0Y1_B_T_top
rlabel metal2 82 653184 82 653184 0 Tile_X0Y1_B_config_C_bit0
rlabel metal2 82 654192 82 654192 0 Tile_X0Y1_B_config_C_bit1
rlabel metal2 82 655200 82 655200 0 Tile_X0Y1_B_config_C_bit2
rlabel metal2 82 656208 82 656208 0 Tile_X0Y1_B_config_C_bit3
rlabel metal2 82 595728 82 595728 0 Tile_X0Y2_A_I_top
rlabel metal2 82 594720 82 594720 0 Tile_X0Y2_A_O_top
rlabel metal2 82 596736 82 596736 0 Tile_X0Y2_A_T_top
rlabel metal2 82 600768 82 600768 0 Tile_X0Y2_A_config_C_bit0
rlabel metal2 82 601776 82 601776 0 Tile_X0Y2_A_config_C_bit1
rlabel metal2 82 602784 82 602784 0 Tile_X0Y2_A_config_C_bit2
rlabel metal2 82 603792 82 603792 0 Tile_X0Y2_A_config_C_bit3
rlabel metal2 82 598752 82 598752 0 Tile_X0Y2_B_I_top
rlabel metal2 82 597744 82 597744 0 Tile_X0Y2_B_O_top
rlabel metal2 82 599760 82 599760 0 Tile_X0Y2_B_T_top
rlabel metal2 82 604800 82 604800 0 Tile_X0Y2_B_config_C_bit0
rlabel metal2 82 605808 82 605808 0 Tile_X0Y2_B_config_C_bit1
rlabel metal2 82 606816 82 606816 0 Tile_X0Y2_B_config_C_bit2
rlabel metal2 82 607824 82 607824 0 Tile_X0Y2_B_config_C_bit3
rlabel metal2 82 547344 82 547344 0 Tile_X0Y3_A_I_top
rlabel metal2 82 546336 82 546336 0 Tile_X0Y3_A_O_top
rlabel metal2 82 548352 82 548352 0 Tile_X0Y3_A_T_top
rlabel metal2 82 552384 82 552384 0 Tile_X0Y3_A_config_C_bit0
rlabel metal2 82 553392 82 553392 0 Tile_X0Y3_A_config_C_bit1
rlabel metal2 82 554400 82 554400 0 Tile_X0Y3_A_config_C_bit2
rlabel metal2 82 555408 82 555408 0 Tile_X0Y3_A_config_C_bit3
rlabel metal2 82 550368 82 550368 0 Tile_X0Y3_B_I_top
rlabel metal2 82 549360 82 549360 0 Tile_X0Y3_B_O_top
rlabel metal2 82 551376 82 551376 0 Tile_X0Y3_B_T_top
rlabel metal2 82 556416 82 556416 0 Tile_X0Y3_B_config_C_bit0
rlabel metal2 82 557424 82 557424 0 Tile_X0Y3_B_config_C_bit1
rlabel metal2 82 558432 82 558432 0 Tile_X0Y3_B_config_C_bit2
rlabel metal2 82 559440 82 559440 0 Tile_X0Y3_B_config_C_bit3
rlabel metal2 82 498960 82 498960 0 Tile_X0Y4_A_I_top
rlabel metal2 82 497952 82 497952 0 Tile_X0Y4_A_O_top
rlabel metal2 82 499968 82 499968 0 Tile_X0Y4_A_T_top
rlabel metal2 82 504000 82 504000 0 Tile_X0Y4_A_config_C_bit0
rlabel metal2 82 505008 82 505008 0 Tile_X0Y4_A_config_C_bit1
rlabel metal2 82 506016 82 506016 0 Tile_X0Y4_A_config_C_bit2
rlabel metal2 82 507024 82 507024 0 Tile_X0Y4_A_config_C_bit3
rlabel metal2 82 501984 82 501984 0 Tile_X0Y4_B_I_top
rlabel metal2 82 500976 82 500976 0 Tile_X0Y4_B_O_top
rlabel metal2 82 502992 82 502992 0 Tile_X0Y4_B_T_top
rlabel metal2 82 508032 82 508032 0 Tile_X0Y4_B_config_C_bit0
rlabel metal2 82 509040 82 509040 0 Tile_X0Y4_B_config_C_bit1
rlabel metal2 82 510048 82 510048 0 Tile_X0Y4_B_config_C_bit2
rlabel metal2 82 511056 82 511056 0 Tile_X0Y4_B_config_C_bit3
rlabel metal2 82 450576 82 450576 0 Tile_X0Y5_A_I_top
rlabel metal2 82 449568 82 449568 0 Tile_X0Y5_A_O_top
rlabel metal2 82 451584 82 451584 0 Tile_X0Y5_A_T_top
rlabel metal2 82 455616 82 455616 0 Tile_X0Y5_A_config_C_bit0
rlabel metal2 82 456624 82 456624 0 Tile_X0Y5_A_config_C_bit1
rlabel metal2 82 457632 82 457632 0 Tile_X0Y5_A_config_C_bit2
rlabel metal2 82 458640 82 458640 0 Tile_X0Y5_A_config_C_bit3
rlabel metal2 82 453600 82 453600 0 Tile_X0Y5_B_I_top
rlabel metal2 82 452592 82 452592 0 Tile_X0Y5_B_O_top
rlabel metal2 82 454608 82 454608 0 Tile_X0Y5_B_T_top
rlabel metal2 82 459648 82 459648 0 Tile_X0Y5_B_config_C_bit0
rlabel metal2 82 460656 82 460656 0 Tile_X0Y5_B_config_C_bit1
rlabel metal2 82 461664 82 461664 0 Tile_X0Y5_B_config_C_bit2
rlabel metal2 82 462672 82 462672 0 Tile_X0Y5_B_config_C_bit3
rlabel metal2 82 402192 82 402192 0 Tile_X0Y6_A_I_top
rlabel metal2 82 401184 82 401184 0 Tile_X0Y6_A_O_top
rlabel metal2 82 403200 82 403200 0 Tile_X0Y6_A_T_top
rlabel metal2 82 407232 82 407232 0 Tile_X0Y6_A_config_C_bit0
rlabel metal2 82 408240 82 408240 0 Tile_X0Y6_A_config_C_bit1
rlabel metal2 82 409248 82 409248 0 Tile_X0Y6_A_config_C_bit2
rlabel metal2 82 410256 82 410256 0 Tile_X0Y6_A_config_C_bit3
rlabel metal2 82 405216 82 405216 0 Tile_X0Y6_B_I_top
rlabel metal2 82 404208 82 404208 0 Tile_X0Y6_B_O_top
rlabel metal2 82 406224 82 406224 0 Tile_X0Y6_B_T_top
rlabel metal2 82 411264 82 411264 0 Tile_X0Y6_B_config_C_bit0
rlabel metal2 82 412272 82 412272 0 Tile_X0Y6_B_config_C_bit1
rlabel metal2 82 413280 82 413280 0 Tile_X0Y6_B_config_C_bit2
rlabel metal2 82 414288 82 414288 0 Tile_X0Y6_B_config_C_bit3
rlabel metal2 82 353808 82 353808 0 Tile_X0Y7_A_I_top
rlabel metal2 82 352800 82 352800 0 Tile_X0Y7_A_O_top
rlabel metal2 82 354816 82 354816 0 Tile_X0Y7_A_T_top
rlabel metal2 82 358848 82 358848 0 Tile_X0Y7_A_config_C_bit0
rlabel metal2 82 359856 82 359856 0 Tile_X0Y7_A_config_C_bit1
rlabel metal2 82 360864 82 360864 0 Tile_X0Y7_A_config_C_bit2
rlabel metal2 82 361872 82 361872 0 Tile_X0Y7_A_config_C_bit3
rlabel metal2 82 356832 82 356832 0 Tile_X0Y7_B_I_top
rlabel metal2 82 355824 82 355824 0 Tile_X0Y7_B_O_top
rlabel metal2 82 357840 82 357840 0 Tile_X0Y7_B_T_top
rlabel metal2 82 362880 82 362880 0 Tile_X0Y7_B_config_C_bit0
rlabel metal2 82 363888 82 363888 0 Tile_X0Y7_B_config_C_bit1
rlabel metal2 82 364896 82 364896 0 Tile_X0Y7_B_config_C_bit2
rlabel metal2 82 365904 82 365904 0 Tile_X0Y7_B_config_C_bit3
rlabel metal2 82 305424 82 305424 0 Tile_X0Y8_A_I_top
rlabel metal2 82 304416 82 304416 0 Tile_X0Y8_A_O_top
rlabel metal2 82 306432 82 306432 0 Tile_X0Y8_A_T_top
rlabel metal2 82 310464 82 310464 0 Tile_X0Y8_A_config_C_bit0
rlabel metal2 82 311472 82 311472 0 Tile_X0Y8_A_config_C_bit1
rlabel metal2 82 312480 82 312480 0 Tile_X0Y8_A_config_C_bit2
rlabel metal2 82 313488 82 313488 0 Tile_X0Y8_A_config_C_bit3
rlabel metal2 82 308448 82 308448 0 Tile_X0Y8_B_I_top
rlabel metal2 82 307440 82 307440 0 Tile_X0Y8_B_O_top
rlabel metal2 82 309456 82 309456 0 Tile_X0Y8_B_T_top
rlabel metal2 82 314496 82 314496 0 Tile_X0Y8_B_config_C_bit0
rlabel metal2 82 315504 82 315504 0 Tile_X0Y8_B_config_C_bit1
rlabel metal2 82 316512 82 316512 0 Tile_X0Y8_B_config_C_bit2
rlabel metal2 82 317520 82 317520 0 Tile_X0Y8_B_config_C_bit3
rlabel metal2 82 257040 82 257040 0 Tile_X0Y9_A_I_top
rlabel metal2 82 256032 82 256032 0 Tile_X0Y9_A_O_top
rlabel metal2 82 258048 82 258048 0 Tile_X0Y9_A_T_top
rlabel metal2 82 262080 82 262080 0 Tile_X0Y9_A_config_C_bit0
rlabel metal2 82 263088 82 263088 0 Tile_X0Y9_A_config_C_bit1
rlabel metal2 82 264096 82 264096 0 Tile_X0Y9_A_config_C_bit2
rlabel metal2 82 265104 82 265104 0 Tile_X0Y9_A_config_C_bit3
rlabel metal2 82 260064 82 260064 0 Tile_X0Y9_B_I_top
rlabel metal2 82 259056 82 259056 0 Tile_X0Y9_B_O_top
rlabel metal2 82 261072 82 261072 0 Tile_X0Y9_B_T_top
rlabel metal2 82 266112 82 266112 0 Tile_X0Y9_B_config_C_bit0
rlabel metal2 82 267120 82 267120 0 Tile_X0Y9_B_config_C_bit1
rlabel metal2 82 268128 82 268128 0 Tile_X0Y9_B_config_C_bit2
rlabel metal2 82 269136 82 269136 0 Tile_X0Y9_B_config_C_bit3
rlabel metal2 452558 226800 452558 226800 0 Tile_X10Y10_ADDR_SRAM0
rlabel metal2 452558 227304 452558 227304 0 Tile_X10Y10_ADDR_SRAM1
rlabel metal2 452558 227808 452558 227808 0 Tile_X10Y10_ADDR_SRAM2
rlabel metal2 452558 228312 452558 228312 0 Tile_X10Y10_ADDR_SRAM3
rlabel metal2 452558 228816 452558 228816 0 Tile_X10Y10_ADDR_SRAM4
rlabel metal2 452558 229320 452558 229320 0 Tile_X10Y10_ADDR_SRAM5
rlabel metal2 452558 229824 452558 229824 0 Tile_X10Y10_ADDR_SRAM6
rlabel metal2 452558 230328 452558 230328 0 Tile_X10Y10_ADDR_SRAM7
rlabel metal2 452558 230832 452558 230832 0 Tile_X10Y10_ADDR_SRAM8
rlabel metal2 452558 231336 452558 231336 0 Tile_X10Y10_ADDR_SRAM9
rlabel metal2 452558 231840 452558 231840 0 Tile_X10Y10_BM_SRAM0
rlabel metal2 452558 232344 452558 232344 0 Tile_X10Y10_BM_SRAM1
rlabel metal2 452558 236880 452558 236880 0 Tile_X10Y10_BM_SRAM10
rlabel metal2 452558 237384 452558 237384 0 Tile_X10Y10_BM_SRAM11
rlabel metal2 452558 237888 452558 237888 0 Tile_X10Y10_BM_SRAM12
rlabel metal2 452558 238392 452558 238392 0 Tile_X10Y10_BM_SRAM13
rlabel metal2 452558 238896 452558 238896 0 Tile_X10Y10_BM_SRAM14
rlabel metal2 452558 239400 452558 239400 0 Tile_X10Y10_BM_SRAM15
rlabel metal2 452558 239904 452558 239904 0 Tile_X10Y10_BM_SRAM16
rlabel metal2 452558 240408 452558 240408 0 Tile_X10Y10_BM_SRAM17
rlabel metal2 452558 240912 452558 240912 0 Tile_X10Y10_BM_SRAM18
rlabel metal2 452558 241416 452558 241416 0 Tile_X10Y10_BM_SRAM19
rlabel metal2 452558 232848 452558 232848 0 Tile_X10Y10_BM_SRAM2
rlabel metal2 452558 241920 452558 241920 0 Tile_X10Y10_BM_SRAM20
rlabel metal2 452558 242424 452558 242424 0 Tile_X10Y10_BM_SRAM21
rlabel metal2 452558 242928 452558 242928 0 Tile_X10Y10_BM_SRAM22
rlabel metal2 452558 243432 452558 243432 0 Tile_X10Y10_BM_SRAM23
rlabel metal2 452558 243936 452558 243936 0 Tile_X10Y10_BM_SRAM24
rlabel metal2 452558 244440 452558 244440 0 Tile_X10Y10_BM_SRAM25
rlabel metal2 452558 244944 452558 244944 0 Tile_X10Y10_BM_SRAM26
rlabel metal2 452558 245448 452558 245448 0 Tile_X10Y10_BM_SRAM27
rlabel metal2 452558 245952 452558 245952 0 Tile_X10Y10_BM_SRAM28
rlabel metal2 452558 246456 452558 246456 0 Tile_X10Y10_BM_SRAM29
rlabel metal2 452558 233352 452558 233352 0 Tile_X10Y10_BM_SRAM3
rlabel metal2 452558 246960 452558 246960 0 Tile_X10Y10_BM_SRAM30
rlabel metal2 452558 247464 452558 247464 0 Tile_X10Y10_BM_SRAM31
rlabel metal2 452558 233856 452558 233856 0 Tile_X10Y10_BM_SRAM4
rlabel metal2 452558 234360 452558 234360 0 Tile_X10Y10_BM_SRAM5
rlabel metal2 452558 234864 452558 234864 0 Tile_X10Y10_BM_SRAM6
rlabel metal2 452558 235368 452558 235368 0 Tile_X10Y10_BM_SRAM7
rlabel metal2 452558 235872 452558 235872 0 Tile_X10Y10_BM_SRAM8
rlabel metal2 452558 236376 452558 236376 0 Tile_X10Y10_BM_SRAM9
rlabel metal2 452558 247968 452558 247968 0 Tile_X10Y10_CLK_SRAM
rlabel metal2 452558 210168 452558 210168 0 Tile_X10Y10_CONFIGURED_top
rlabel metal2 452558 248472 452558 248472 0 Tile_X10Y10_DIN_SRAM0
rlabel metal2 452558 248976 452558 248976 0 Tile_X10Y10_DIN_SRAM1
rlabel metal2 452558 253512 452558 253512 0 Tile_X10Y10_DIN_SRAM10
rlabel metal2 452558 254016 452558 254016 0 Tile_X10Y10_DIN_SRAM11
rlabel metal2 452558 254520 452558 254520 0 Tile_X10Y10_DIN_SRAM12
rlabel metal2 452558 255024 452558 255024 0 Tile_X10Y10_DIN_SRAM13
rlabel metal2 452558 255528 452558 255528 0 Tile_X10Y10_DIN_SRAM14
rlabel metal2 452558 256032 452558 256032 0 Tile_X10Y10_DIN_SRAM15
rlabel metal2 452558 256536 452558 256536 0 Tile_X10Y10_DIN_SRAM16
rlabel metal2 452558 257040 452558 257040 0 Tile_X10Y10_DIN_SRAM17
rlabel metal2 452558 257544 452558 257544 0 Tile_X10Y10_DIN_SRAM18
rlabel metal2 452558 258048 452558 258048 0 Tile_X10Y10_DIN_SRAM19
rlabel metal2 452558 249480 452558 249480 0 Tile_X10Y10_DIN_SRAM2
rlabel metal2 452558 258552 452558 258552 0 Tile_X10Y10_DIN_SRAM20
rlabel metal2 452558 259056 452558 259056 0 Tile_X10Y10_DIN_SRAM21
rlabel metal2 452558 259560 452558 259560 0 Tile_X10Y10_DIN_SRAM22
rlabel metal2 452558 260064 452558 260064 0 Tile_X10Y10_DIN_SRAM23
rlabel metal2 452558 260568 452558 260568 0 Tile_X10Y10_DIN_SRAM24
rlabel metal2 452558 261072 452558 261072 0 Tile_X10Y10_DIN_SRAM25
rlabel metal2 452558 261576 452558 261576 0 Tile_X10Y10_DIN_SRAM26
rlabel metal2 452558 262080 452558 262080 0 Tile_X10Y10_DIN_SRAM27
rlabel metal2 452558 262584 452558 262584 0 Tile_X10Y10_DIN_SRAM28
rlabel metal2 452558 263088 452558 263088 0 Tile_X10Y10_DIN_SRAM29
rlabel metal2 452558 249984 452558 249984 0 Tile_X10Y10_DIN_SRAM3
rlabel metal2 452558 263592 452558 263592 0 Tile_X10Y10_DIN_SRAM30
rlabel metal2 452558 264096 452558 264096 0 Tile_X10Y10_DIN_SRAM31
rlabel metal2 452558 250488 452558 250488 0 Tile_X10Y10_DIN_SRAM4
rlabel metal2 452558 250992 452558 250992 0 Tile_X10Y10_DIN_SRAM5
rlabel metal2 452558 251496 452558 251496 0 Tile_X10Y10_DIN_SRAM6
rlabel metal2 452558 252000 452558 252000 0 Tile_X10Y10_DIN_SRAM7
rlabel metal2 452558 252504 452558 252504 0 Tile_X10Y10_DIN_SRAM8
rlabel metal2 452558 253008 452558 253008 0 Tile_X10Y10_DIN_SRAM9
rlabel metal2 452558 210672 452558 210672 0 Tile_X10Y10_DOUT_SRAM0
rlabel metal2 452558 211176 452558 211176 0 Tile_X10Y10_DOUT_SRAM1
rlabel metal2 452558 215712 452558 215712 0 Tile_X10Y10_DOUT_SRAM10
rlabel metal2 452558 216216 452558 216216 0 Tile_X10Y10_DOUT_SRAM11
rlabel metal2 452558 216720 452558 216720 0 Tile_X10Y10_DOUT_SRAM12
rlabel metal2 452558 217224 452558 217224 0 Tile_X10Y10_DOUT_SRAM13
rlabel metal2 452558 217728 452558 217728 0 Tile_X10Y10_DOUT_SRAM14
rlabel metal2 452558 218232 452558 218232 0 Tile_X10Y10_DOUT_SRAM15
rlabel metal2 452558 218736 452558 218736 0 Tile_X10Y10_DOUT_SRAM16
rlabel metal2 452558 219240 452558 219240 0 Tile_X10Y10_DOUT_SRAM17
rlabel metal2 452558 219744 452558 219744 0 Tile_X10Y10_DOUT_SRAM18
rlabel metal2 452558 220248 452558 220248 0 Tile_X10Y10_DOUT_SRAM19
rlabel metal2 452558 211680 452558 211680 0 Tile_X10Y10_DOUT_SRAM2
rlabel metal2 452558 220752 452558 220752 0 Tile_X10Y10_DOUT_SRAM20
rlabel metal2 452558 221256 452558 221256 0 Tile_X10Y10_DOUT_SRAM21
rlabel metal2 452558 221760 452558 221760 0 Tile_X10Y10_DOUT_SRAM22
rlabel metal2 452558 222264 452558 222264 0 Tile_X10Y10_DOUT_SRAM23
rlabel metal2 452558 222768 452558 222768 0 Tile_X10Y10_DOUT_SRAM24
rlabel metal2 452558 223272 452558 223272 0 Tile_X10Y10_DOUT_SRAM25
rlabel metal2 452558 223776 452558 223776 0 Tile_X10Y10_DOUT_SRAM26
rlabel metal2 452558 224280 452558 224280 0 Tile_X10Y10_DOUT_SRAM27
rlabel metal2 452558 224784 452558 224784 0 Tile_X10Y10_DOUT_SRAM28
rlabel metal2 452558 225288 452558 225288 0 Tile_X10Y10_DOUT_SRAM29
rlabel metal2 452558 212184 452558 212184 0 Tile_X10Y10_DOUT_SRAM3
rlabel metal2 452558 225792 452558 225792 0 Tile_X10Y10_DOUT_SRAM30
rlabel metal2 452558 226296 452558 226296 0 Tile_X10Y10_DOUT_SRAM31
rlabel metal2 452558 212688 452558 212688 0 Tile_X10Y10_DOUT_SRAM4
rlabel metal2 452558 213192 452558 213192 0 Tile_X10Y10_DOUT_SRAM5
rlabel metal2 452558 213696 452558 213696 0 Tile_X10Y10_DOUT_SRAM6
rlabel metal2 452558 214200 452558 214200 0 Tile_X10Y10_DOUT_SRAM7
rlabel metal2 452558 214704 452558 214704 0 Tile_X10Y10_DOUT_SRAM8
rlabel metal2 452558 215208 452558 215208 0 Tile_X10Y10_DOUT_SRAM9
rlabel metal2 452558 264600 452558 264600 0 Tile_X10Y10_MEN_SRAM
rlabel metal2 452558 265104 452558 265104 0 Tile_X10Y10_REN_SRAM
rlabel metal2 452558 265608 452558 265608 0 Tile_X10Y10_TIE_HIGH_SRAM
rlabel metal2 452558 266112 452558 266112 0 Tile_X10Y10_TIE_LOW_SRAM
rlabel metal2 452558 266616 452558 266616 0 Tile_X10Y10_WEN_SRAM
rlabel metal2 452558 130032 452558 130032 0 Tile_X10Y12_ADDR_SRAM0
rlabel metal2 452558 130536 452558 130536 0 Tile_X10Y12_ADDR_SRAM1
rlabel metal2 452558 131040 452558 131040 0 Tile_X10Y12_ADDR_SRAM2
rlabel metal2 452558 131544 452558 131544 0 Tile_X10Y12_ADDR_SRAM3
rlabel metal2 452558 132048 452558 132048 0 Tile_X10Y12_ADDR_SRAM4
rlabel metal2 452558 132552 452558 132552 0 Tile_X10Y12_ADDR_SRAM5
rlabel metal2 452558 133056 452558 133056 0 Tile_X10Y12_ADDR_SRAM6
rlabel metal2 452558 133560 452558 133560 0 Tile_X10Y12_ADDR_SRAM7
rlabel metal2 452558 134064 452558 134064 0 Tile_X10Y12_ADDR_SRAM8
rlabel metal2 452558 134568 452558 134568 0 Tile_X10Y12_ADDR_SRAM9
rlabel metal2 452558 135072 452558 135072 0 Tile_X10Y12_BM_SRAM0
rlabel metal2 452558 135576 452558 135576 0 Tile_X10Y12_BM_SRAM1
rlabel metal2 452558 140112 452558 140112 0 Tile_X10Y12_BM_SRAM10
rlabel metal2 452558 140616 452558 140616 0 Tile_X10Y12_BM_SRAM11
rlabel metal2 452558 141120 452558 141120 0 Tile_X10Y12_BM_SRAM12
rlabel metal2 452558 141624 452558 141624 0 Tile_X10Y12_BM_SRAM13
rlabel metal2 452558 142128 452558 142128 0 Tile_X10Y12_BM_SRAM14
rlabel metal2 452558 142632 452558 142632 0 Tile_X10Y12_BM_SRAM15
rlabel metal2 452558 143136 452558 143136 0 Tile_X10Y12_BM_SRAM16
rlabel metal2 452558 143640 452558 143640 0 Tile_X10Y12_BM_SRAM17
rlabel metal2 452558 144144 452558 144144 0 Tile_X10Y12_BM_SRAM18
rlabel metal2 452558 144648 452558 144648 0 Tile_X10Y12_BM_SRAM19
rlabel metal2 452558 136080 452558 136080 0 Tile_X10Y12_BM_SRAM2
rlabel metal2 452558 145152 452558 145152 0 Tile_X10Y12_BM_SRAM20
rlabel metal2 452558 145656 452558 145656 0 Tile_X10Y12_BM_SRAM21
rlabel metal2 452558 146160 452558 146160 0 Tile_X10Y12_BM_SRAM22
rlabel metal2 452558 146664 452558 146664 0 Tile_X10Y12_BM_SRAM23
rlabel metal2 452558 147168 452558 147168 0 Tile_X10Y12_BM_SRAM24
rlabel metal2 452558 147672 452558 147672 0 Tile_X10Y12_BM_SRAM25
rlabel metal2 452558 148176 452558 148176 0 Tile_X10Y12_BM_SRAM26
rlabel metal2 452558 148680 452558 148680 0 Tile_X10Y12_BM_SRAM27
rlabel metal2 452558 149184 452558 149184 0 Tile_X10Y12_BM_SRAM28
rlabel metal2 452558 149688 452558 149688 0 Tile_X10Y12_BM_SRAM29
rlabel metal2 452558 136584 452558 136584 0 Tile_X10Y12_BM_SRAM3
rlabel metal2 452558 150192 452558 150192 0 Tile_X10Y12_BM_SRAM30
rlabel metal2 452558 150696 452558 150696 0 Tile_X10Y12_BM_SRAM31
rlabel metal2 452558 137088 452558 137088 0 Tile_X10Y12_BM_SRAM4
rlabel metal2 452558 137592 452558 137592 0 Tile_X10Y12_BM_SRAM5
rlabel metal2 452558 138096 452558 138096 0 Tile_X10Y12_BM_SRAM6
rlabel metal2 452558 138600 452558 138600 0 Tile_X10Y12_BM_SRAM7
rlabel metal2 452558 139104 452558 139104 0 Tile_X10Y12_BM_SRAM8
rlabel metal2 452558 139608 452558 139608 0 Tile_X10Y12_BM_SRAM9
rlabel metal2 452558 151200 452558 151200 0 Tile_X10Y12_CLK_SRAM
rlabel metal2 452558 113400 452558 113400 0 Tile_X10Y12_CONFIGURED_top
rlabel metal2 452558 151704 452558 151704 0 Tile_X10Y12_DIN_SRAM0
rlabel metal2 452558 152208 452558 152208 0 Tile_X10Y12_DIN_SRAM1
rlabel metal2 452558 156744 452558 156744 0 Tile_X10Y12_DIN_SRAM10
rlabel metal2 452558 157248 452558 157248 0 Tile_X10Y12_DIN_SRAM11
rlabel metal2 452558 157752 452558 157752 0 Tile_X10Y12_DIN_SRAM12
rlabel metal2 452558 158256 452558 158256 0 Tile_X10Y12_DIN_SRAM13
rlabel metal2 452558 158760 452558 158760 0 Tile_X10Y12_DIN_SRAM14
rlabel metal2 452558 159264 452558 159264 0 Tile_X10Y12_DIN_SRAM15
rlabel metal2 452558 159768 452558 159768 0 Tile_X10Y12_DIN_SRAM16
rlabel metal2 452558 160272 452558 160272 0 Tile_X10Y12_DIN_SRAM17
rlabel metal2 452558 160776 452558 160776 0 Tile_X10Y12_DIN_SRAM18
rlabel metal2 452558 161280 452558 161280 0 Tile_X10Y12_DIN_SRAM19
rlabel metal2 452558 152712 452558 152712 0 Tile_X10Y12_DIN_SRAM2
rlabel metal2 452558 161784 452558 161784 0 Tile_X10Y12_DIN_SRAM20
rlabel metal2 452558 162288 452558 162288 0 Tile_X10Y12_DIN_SRAM21
rlabel metal2 452558 162792 452558 162792 0 Tile_X10Y12_DIN_SRAM22
rlabel metal2 452558 163296 452558 163296 0 Tile_X10Y12_DIN_SRAM23
rlabel metal2 452558 163800 452558 163800 0 Tile_X10Y12_DIN_SRAM24
rlabel metal2 452558 164304 452558 164304 0 Tile_X10Y12_DIN_SRAM25
rlabel metal2 452558 164808 452558 164808 0 Tile_X10Y12_DIN_SRAM26
rlabel metal2 452558 165312 452558 165312 0 Tile_X10Y12_DIN_SRAM27
rlabel metal2 452558 165816 452558 165816 0 Tile_X10Y12_DIN_SRAM28
rlabel metal2 452558 166320 452558 166320 0 Tile_X10Y12_DIN_SRAM29
rlabel metal2 452558 153216 452558 153216 0 Tile_X10Y12_DIN_SRAM3
rlabel metal2 452558 166824 452558 166824 0 Tile_X10Y12_DIN_SRAM30
rlabel metal2 452558 167328 452558 167328 0 Tile_X10Y12_DIN_SRAM31
rlabel metal2 452558 153720 452558 153720 0 Tile_X10Y12_DIN_SRAM4
rlabel metal2 452558 154224 452558 154224 0 Tile_X10Y12_DIN_SRAM5
rlabel metal2 452558 154728 452558 154728 0 Tile_X10Y12_DIN_SRAM6
rlabel metal2 452558 155232 452558 155232 0 Tile_X10Y12_DIN_SRAM7
rlabel metal2 452558 155736 452558 155736 0 Tile_X10Y12_DIN_SRAM8
rlabel metal2 452558 156240 452558 156240 0 Tile_X10Y12_DIN_SRAM9
rlabel metal2 452558 113904 452558 113904 0 Tile_X10Y12_DOUT_SRAM0
rlabel metal2 452558 114408 452558 114408 0 Tile_X10Y12_DOUT_SRAM1
rlabel metal2 452558 118944 452558 118944 0 Tile_X10Y12_DOUT_SRAM10
rlabel metal2 452558 119448 452558 119448 0 Tile_X10Y12_DOUT_SRAM11
rlabel metal2 452558 119952 452558 119952 0 Tile_X10Y12_DOUT_SRAM12
rlabel metal2 452558 120456 452558 120456 0 Tile_X10Y12_DOUT_SRAM13
rlabel metal2 452558 120960 452558 120960 0 Tile_X10Y12_DOUT_SRAM14
rlabel metal2 452558 121464 452558 121464 0 Tile_X10Y12_DOUT_SRAM15
rlabel metal2 452558 121968 452558 121968 0 Tile_X10Y12_DOUT_SRAM16
rlabel metal2 452558 122472 452558 122472 0 Tile_X10Y12_DOUT_SRAM17
rlabel metal2 452558 122976 452558 122976 0 Tile_X10Y12_DOUT_SRAM18
rlabel metal2 452558 123480 452558 123480 0 Tile_X10Y12_DOUT_SRAM19
rlabel metal2 452558 114912 452558 114912 0 Tile_X10Y12_DOUT_SRAM2
rlabel metal2 452558 123984 452558 123984 0 Tile_X10Y12_DOUT_SRAM20
rlabel metal2 452558 124488 452558 124488 0 Tile_X10Y12_DOUT_SRAM21
rlabel metal2 452558 124992 452558 124992 0 Tile_X10Y12_DOUT_SRAM22
rlabel metal2 452558 125496 452558 125496 0 Tile_X10Y12_DOUT_SRAM23
rlabel metal2 452558 126000 452558 126000 0 Tile_X10Y12_DOUT_SRAM24
rlabel metal2 452558 126504 452558 126504 0 Tile_X10Y12_DOUT_SRAM25
rlabel metal2 452558 127008 452558 127008 0 Tile_X10Y12_DOUT_SRAM26
rlabel metal2 452558 127512 452558 127512 0 Tile_X10Y12_DOUT_SRAM27
rlabel metal2 452558 128016 452558 128016 0 Tile_X10Y12_DOUT_SRAM28
rlabel metal2 452558 128520 452558 128520 0 Tile_X10Y12_DOUT_SRAM29
rlabel metal2 452558 115416 452558 115416 0 Tile_X10Y12_DOUT_SRAM3
rlabel metal2 452558 129024 452558 129024 0 Tile_X10Y12_DOUT_SRAM30
rlabel metal2 452558 129528 452558 129528 0 Tile_X10Y12_DOUT_SRAM31
rlabel metal2 452558 115920 452558 115920 0 Tile_X10Y12_DOUT_SRAM4
rlabel metal2 452558 116424 452558 116424 0 Tile_X10Y12_DOUT_SRAM5
rlabel metal2 452558 116928 452558 116928 0 Tile_X10Y12_DOUT_SRAM6
rlabel metal2 452558 117432 452558 117432 0 Tile_X10Y12_DOUT_SRAM7
rlabel metal2 452558 117936 452558 117936 0 Tile_X10Y12_DOUT_SRAM8
rlabel metal2 452558 118440 452558 118440 0 Tile_X10Y12_DOUT_SRAM9
rlabel metal2 452558 167832 452558 167832 0 Tile_X10Y12_MEN_SRAM
rlabel metal2 452558 168336 452558 168336 0 Tile_X10Y12_REN_SRAM
rlabel metal2 452558 168840 452558 168840 0 Tile_X10Y12_TIE_HIGH_SRAM
rlabel metal2 452558 169344 452558 169344 0 Tile_X10Y12_TIE_LOW_SRAM
rlabel metal2 452558 169848 452558 169848 0 Tile_X10Y12_WEN_SRAM
rlabel metal2 452558 33264 452558 33264 0 Tile_X10Y14_ADDR_SRAM0
rlabel metal2 452558 33768 452558 33768 0 Tile_X10Y14_ADDR_SRAM1
rlabel metal2 452558 34272 452558 34272 0 Tile_X10Y14_ADDR_SRAM2
rlabel metal2 452558 34776 452558 34776 0 Tile_X10Y14_ADDR_SRAM3
rlabel metal2 452558 35280 452558 35280 0 Tile_X10Y14_ADDR_SRAM4
rlabel metal2 452558 35784 452558 35784 0 Tile_X10Y14_ADDR_SRAM5
rlabel metal2 452558 36288 452558 36288 0 Tile_X10Y14_ADDR_SRAM6
rlabel metal2 452558 36792 452558 36792 0 Tile_X10Y14_ADDR_SRAM7
rlabel metal2 452558 37296 452558 37296 0 Tile_X10Y14_ADDR_SRAM8
rlabel metal2 452558 37800 452558 37800 0 Tile_X10Y14_ADDR_SRAM9
rlabel metal2 452558 38304 452558 38304 0 Tile_X10Y14_BM_SRAM0
rlabel metal2 452558 38808 452558 38808 0 Tile_X10Y14_BM_SRAM1
rlabel metal2 452558 43344 452558 43344 0 Tile_X10Y14_BM_SRAM10
rlabel metal2 452558 43848 452558 43848 0 Tile_X10Y14_BM_SRAM11
rlabel metal2 452558 44352 452558 44352 0 Tile_X10Y14_BM_SRAM12
rlabel metal2 452558 44856 452558 44856 0 Tile_X10Y14_BM_SRAM13
rlabel metal2 452558 45360 452558 45360 0 Tile_X10Y14_BM_SRAM14
rlabel metal2 452558 45864 452558 45864 0 Tile_X10Y14_BM_SRAM15
rlabel metal2 452558 46368 452558 46368 0 Tile_X10Y14_BM_SRAM16
rlabel metal2 452558 46872 452558 46872 0 Tile_X10Y14_BM_SRAM17
rlabel metal2 452558 47376 452558 47376 0 Tile_X10Y14_BM_SRAM18
rlabel metal2 452558 47880 452558 47880 0 Tile_X10Y14_BM_SRAM19
rlabel metal2 452558 39312 452558 39312 0 Tile_X10Y14_BM_SRAM2
rlabel metal2 452558 48384 452558 48384 0 Tile_X10Y14_BM_SRAM20
rlabel metal2 452558 48888 452558 48888 0 Tile_X10Y14_BM_SRAM21
rlabel metal2 452558 49392 452558 49392 0 Tile_X10Y14_BM_SRAM22
rlabel metal2 452558 49896 452558 49896 0 Tile_X10Y14_BM_SRAM23
rlabel metal2 452558 50400 452558 50400 0 Tile_X10Y14_BM_SRAM24
rlabel metal2 452558 50904 452558 50904 0 Tile_X10Y14_BM_SRAM25
rlabel metal2 452558 51408 452558 51408 0 Tile_X10Y14_BM_SRAM26
rlabel metal2 452558 51912 452558 51912 0 Tile_X10Y14_BM_SRAM27
rlabel metal2 452558 52416 452558 52416 0 Tile_X10Y14_BM_SRAM28
rlabel metal2 452558 52920 452558 52920 0 Tile_X10Y14_BM_SRAM29
rlabel metal2 452558 39816 452558 39816 0 Tile_X10Y14_BM_SRAM3
rlabel metal2 452558 53424 452558 53424 0 Tile_X10Y14_BM_SRAM30
rlabel metal2 452558 53928 452558 53928 0 Tile_X10Y14_BM_SRAM31
rlabel metal2 452558 40320 452558 40320 0 Tile_X10Y14_BM_SRAM4
rlabel metal2 452558 40824 452558 40824 0 Tile_X10Y14_BM_SRAM5
rlabel metal2 452558 41328 452558 41328 0 Tile_X10Y14_BM_SRAM6
rlabel metal2 452558 41832 452558 41832 0 Tile_X10Y14_BM_SRAM7
rlabel metal2 452558 42336 452558 42336 0 Tile_X10Y14_BM_SRAM8
rlabel metal2 452558 42840 452558 42840 0 Tile_X10Y14_BM_SRAM9
rlabel metal2 452558 54432 452558 54432 0 Tile_X10Y14_CLK_SRAM
rlabel metal2 452558 16632 452558 16632 0 Tile_X10Y14_CONFIGURED_top
rlabel metal2 452558 54936 452558 54936 0 Tile_X10Y14_DIN_SRAM0
rlabel metal2 452558 55440 452558 55440 0 Tile_X10Y14_DIN_SRAM1
rlabel metal2 452558 59976 452558 59976 0 Tile_X10Y14_DIN_SRAM10
rlabel metal2 452558 60480 452558 60480 0 Tile_X10Y14_DIN_SRAM11
rlabel metal2 452558 60984 452558 60984 0 Tile_X10Y14_DIN_SRAM12
rlabel metal2 452558 61488 452558 61488 0 Tile_X10Y14_DIN_SRAM13
rlabel metal2 452558 61992 452558 61992 0 Tile_X10Y14_DIN_SRAM14
rlabel metal2 452558 62496 452558 62496 0 Tile_X10Y14_DIN_SRAM15
rlabel metal2 452558 63000 452558 63000 0 Tile_X10Y14_DIN_SRAM16
rlabel metal2 452558 63504 452558 63504 0 Tile_X10Y14_DIN_SRAM17
rlabel metal2 452558 64008 452558 64008 0 Tile_X10Y14_DIN_SRAM18
rlabel metal2 452558 64512 452558 64512 0 Tile_X10Y14_DIN_SRAM19
rlabel metal2 452558 55944 452558 55944 0 Tile_X10Y14_DIN_SRAM2
rlabel metal2 452558 65016 452558 65016 0 Tile_X10Y14_DIN_SRAM20
rlabel metal2 452558 65520 452558 65520 0 Tile_X10Y14_DIN_SRAM21
rlabel metal2 452558 66024 452558 66024 0 Tile_X10Y14_DIN_SRAM22
rlabel metal2 452558 66528 452558 66528 0 Tile_X10Y14_DIN_SRAM23
rlabel metal2 452558 67032 452558 67032 0 Tile_X10Y14_DIN_SRAM24
rlabel metal2 452558 67536 452558 67536 0 Tile_X10Y14_DIN_SRAM25
rlabel metal2 452558 68040 452558 68040 0 Tile_X10Y14_DIN_SRAM26
rlabel metal2 452558 68544 452558 68544 0 Tile_X10Y14_DIN_SRAM27
rlabel metal2 452558 69048 452558 69048 0 Tile_X10Y14_DIN_SRAM28
rlabel metal2 452558 69552 452558 69552 0 Tile_X10Y14_DIN_SRAM29
rlabel metal2 452558 56448 452558 56448 0 Tile_X10Y14_DIN_SRAM3
rlabel metal2 452558 70056 452558 70056 0 Tile_X10Y14_DIN_SRAM30
rlabel metal2 452558 70560 452558 70560 0 Tile_X10Y14_DIN_SRAM31
rlabel metal2 452558 56952 452558 56952 0 Tile_X10Y14_DIN_SRAM4
rlabel metal2 452558 57456 452558 57456 0 Tile_X10Y14_DIN_SRAM5
rlabel metal2 452558 57960 452558 57960 0 Tile_X10Y14_DIN_SRAM6
rlabel metal2 452558 58464 452558 58464 0 Tile_X10Y14_DIN_SRAM7
rlabel metal2 452558 58968 452558 58968 0 Tile_X10Y14_DIN_SRAM8
rlabel metal2 452558 59472 452558 59472 0 Tile_X10Y14_DIN_SRAM9
rlabel metal2 452558 17136 452558 17136 0 Tile_X10Y14_DOUT_SRAM0
rlabel metal2 452558 17640 452558 17640 0 Tile_X10Y14_DOUT_SRAM1
rlabel metal2 452558 22176 452558 22176 0 Tile_X10Y14_DOUT_SRAM10
rlabel metal2 452558 22680 452558 22680 0 Tile_X10Y14_DOUT_SRAM11
rlabel metal2 452558 23184 452558 23184 0 Tile_X10Y14_DOUT_SRAM12
rlabel metal2 452558 23688 452558 23688 0 Tile_X10Y14_DOUT_SRAM13
rlabel metal2 452558 24192 452558 24192 0 Tile_X10Y14_DOUT_SRAM14
rlabel metal2 452558 24696 452558 24696 0 Tile_X10Y14_DOUT_SRAM15
rlabel metal2 452558 25200 452558 25200 0 Tile_X10Y14_DOUT_SRAM16
rlabel metal2 452558 25704 452558 25704 0 Tile_X10Y14_DOUT_SRAM17
rlabel metal2 452558 26208 452558 26208 0 Tile_X10Y14_DOUT_SRAM18
rlabel metal2 452558 26712 452558 26712 0 Tile_X10Y14_DOUT_SRAM19
rlabel metal2 452558 18144 452558 18144 0 Tile_X10Y14_DOUT_SRAM2
rlabel metal2 452558 27216 452558 27216 0 Tile_X10Y14_DOUT_SRAM20
rlabel metal2 452558 27720 452558 27720 0 Tile_X10Y14_DOUT_SRAM21
rlabel metal2 452558 28224 452558 28224 0 Tile_X10Y14_DOUT_SRAM22
rlabel metal2 452558 28728 452558 28728 0 Tile_X10Y14_DOUT_SRAM23
rlabel metal2 452558 29232 452558 29232 0 Tile_X10Y14_DOUT_SRAM24
rlabel metal2 452558 29736 452558 29736 0 Tile_X10Y14_DOUT_SRAM25
rlabel metal2 452558 30240 452558 30240 0 Tile_X10Y14_DOUT_SRAM26
rlabel metal2 452558 30744 452558 30744 0 Tile_X10Y14_DOUT_SRAM27
rlabel metal2 452558 31248 452558 31248 0 Tile_X10Y14_DOUT_SRAM28
rlabel metal2 452558 31752 452558 31752 0 Tile_X10Y14_DOUT_SRAM29
rlabel metal2 452558 18648 452558 18648 0 Tile_X10Y14_DOUT_SRAM3
rlabel metal2 452558 32256 452558 32256 0 Tile_X10Y14_DOUT_SRAM30
rlabel metal2 452558 32760 452558 32760 0 Tile_X10Y14_DOUT_SRAM31
rlabel metal2 452558 19152 452558 19152 0 Tile_X10Y14_DOUT_SRAM4
rlabel metal2 452558 19656 452558 19656 0 Tile_X10Y14_DOUT_SRAM5
rlabel metal2 452558 20160 452558 20160 0 Tile_X10Y14_DOUT_SRAM6
rlabel metal2 452558 20664 452558 20664 0 Tile_X10Y14_DOUT_SRAM7
rlabel metal2 452558 21168 452558 21168 0 Tile_X10Y14_DOUT_SRAM8
rlabel metal2 452558 21672 452558 21672 0 Tile_X10Y14_DOUT_SRAM9
rlabel metal2 452558 71064 452558 71064 0 Tile_X10Y14_MEN_SRAM
rlabel metal2 452558 71568 452558 71568 0 Tile_X10Y14_REN_SRAM
rlabel metal2 452558 72072 452558 72072 0 Tile_X10Y14_TIE_HIGH_SRAM
rlabel metal2 452558 72576 452558 72576 0 Tile_X10Y14_TIE_LOW_SRAM
rlabel metal2 452558 73080 452558 73080 0 Tile_X10Y14_WEN_SRAM
rlabel metal2 452558 613872 452558 613872 0 Tile_X10Y2_ADDR_SRAM0
rlabel metal2 452558 614376 452558 614376 0 Tile_X10Y2_ADDR_SRAM1
rlabel metal2 452558 614880 452558 614880 0 Tile_X10Y2_ADDR_SRAM2
rlabel metal2 452558 615384 452558 615384 0 Tile_X10Y2_ADDR_SRAM3
rlabel metal2 452558 615888 452558 615888 0 Tile_X10Y2_ADDR_SRAM4
rlabel metal2 452558 616392 452558 616392 0 Tile_X10Y2_ADDR_SRAM5
rlabel metal2 452558 616896 452558 616896 0 Tile_X10Y2_ADDR_SRAM6
rlabel metal2 452558 617400 452558 617400 0 Tile_X10Y2_ADDR_SRAM7
rlabel metal2 452558 617904 452558 617904 0 Tile_X10Y2_ADDR_SRAM8
rlabel metal2 452558 618408 452558 618408 0 Tile_X10Y2_ADDR_SRAM9
rlabel metal2 452558 618912 452558 618912 0 Tile_X10Y2_BM_SRAM0
rlabel metal2 452558 619416 452558 619416 0 Tile_X10Y2_BM_SRAM1
rlabel metal2 452558 623952 452558 623952 0 Tile_X10Y2_BM_SRAM10
rlabel metal2 452558 624456 452558 624456 0 Tile_X10Y2_BM_SRAM11
rlabel metal2 452558 624960 452558 624960 0 Tile_X10Y2_BM_SRAM12
rlabel metal2 452558 625464 452558 625464 0 Tile_X10Y2_BM_SRAM13
rlabel metal2 452558 625968 452558 625968 0 Tile_X10Y2_BM_SRAM14
rlabel metal2 452558 626472 452558 626472 0 Tile_X10Y2_BM_SRAM15
rlabel metal2 452558 626976 452558 626976 0 Tile_X10Y2_BM_SRAM16
rlabel metal2 452558 627480 452558 627480 0 Tile_X10Y2_BM_SRAM17
rlabel metal2 452558 627984 452558 627984 0 Tile_X10Y2_BM_SRAM18
rlabel metal2 452558 628488 452558 628488 0 Tile_X10Y2_BM_SRAM19
rlabel metal2 452558 619920 452558 619920 0 Tile_X10Y2_BM_SRAM2
rlabel metal2 452558 628992 452558 628992 0 Tile_X10Y2_BM_SRAM20
rlabel metal2 452558 629496 452558 629496 0 Tile_X10Y2_BM_SRAM21
rlabel metal2 452558 630000 452558 630000 0 Tile_X10Y2_BM_SRAM22
rlabel metal2 452558 630504 452558 630504 0 Tile_X10Y2_BM_SRAM23
rlabel metal2 452558 631008 452558 631008 0 Tile_X10Y2_BM_SRAM24
rlabel metal2 452558 631512 452558 631512 0 Tile_X10Y2_BM_SRAM25
rlabel metal2 452558 632016 452558 632016 0 Tile_X10Y2_BM_SRAM26
rlabel metal2 452558 632520 452558 632520 0 Tile_X10Y2_BM_SRAM27
rlabel metal2 452558 633024 452558 633024 0 Tile_X10Y2_BM_SRAM28
rlabel metal2 452558 633528 452558 633528 0 Tile_X10Y2_BM_SRAM29
rlabel metal2 452558 620424 452558 620424 0 Tile_X10Y2_BM_SRAM3
rlabel metal2 452558 634032 452558 634032 0 Tile_X10Y2_BM_SRAM30
rlabel metal2 452558 634536 452558 634536 0 Tile_X10Y2_BM_SRAM31
rlabel metal2 452558 620928 452558 620928 0 Tile_X10Y2_BM_SRAM4
rlabel metal2 452558 621432 452558 621432 0 Tile_X10Y2_BM_SRAM5
rlabel metal2 452558 621936 452558 621936 0 Tile_X10Y2_BM_SRAM6
rlabel metal2 452558 622440 452558 622440 0 Tile_X10Y2_BM_SRAM7
rlabel metal2 452558 622944 452558 622944 0 Tile_X10Y2_BM_SRAM8
rlabel metal2 452558 623448 452558 623448 0 Tile_X10Y2_BM_SRAM9
rlabel metal2 452558 635040 452558 635040 0 Tile_X10Y2_CLK_SRAM
rlabel metal2 452558 597240 452558 597240 0 Tile_X10Y2_CONFIGURED_top
rlabel metal2 452558 635544 452558 635544 0 Tile_X10Y2_DIN_SRAM0
rlabel metal2 452558 636048 452558 636048 0 Tile_X10Y2_DIN_SRAM1
rlabel metal2 452558 640584 452558 640584 0 Tile_X10Y2_DIN_SRAM10
rlabel metal2 452558 641088 452558 641088 0 Tile_X10Y2_DIN_SRAM11
rlabel metal2 452558 641592 452558 641592 0 Tile_X10Y2_DIN_SRAM12
rlabel metal2 452558 642096 452558 642096 0 Tile_X10Y2_DIN_SRAM13
rlabel metal2 452558 642600 452558 642600 0 Tile_X10Y2_DIN_SRAM14
rlabel metal2 452558 643104 452558 643104 0 Tile_X10Y2_DIN_SRAM15
rlabel metal2 452558 643608 452558 643608 0 Tile_X10Y2_DIN_SRAM16
rlabel metal2 452558 644112 452558 644112 0 Tile_X10Y2_DIN_SRAM17
rlabel metal2 452558 644616 452558 644616 0 Tile_X10Y2_DIN_SRAM18
rlabel metal2 452558 645120 452558 645120 0 Tile_X10Y2_DIN_SRAM19
rlabel metal2 452558 636552 452558 636552 0 Tile_X10Y2_DIN_SRAM2
rlabel metal2 452558 645624 452558 645624 0 Tile_X10Y2_DIN_SRAM20
rlabel metal2 452558 646128 452558 646128 0 Tile_X10Y2_DIN_SRAM21
rlabel metal2 452558 646632 452558 646632 0 Tile_X10Y2_DIN_SRAM22
rlabel metal2 452558 647136 452558 647136 0 Tile_X10Y2_DIN_SRAM23
rlabel metal2 452558 647640 452558 647640 0 Tile_X10Y2_DIN_SRAM24
rlabel metal2 452558 648144 452558 648144 0 Tile_X10Y2_DIN_SRAM25
rlabel metal2 452558 648648 452558 648648 0 Tile_X10Y2_DIN_SRAM26
rlabel metal2 452558 649152 452558 649152 0 Tile_X10Y2_DIN_SRAM27
rlabel metal2 452558 649656 452558 649656 0 Tile_X10Y2_DIN_SRAM28
rlabel metal2 452558 650160 452558 650160 0 Tile_X10Y2_DIN_SRAM29
rlabel metal2 452558 637056 452558 637056 0 Tile_X10Y2_DIN_SRAM3
rlabel metal2 452558 650664 452558 650664 0 Tile_X10Y2_DIN_SRAM30
rlabel metal2 452558 651168 452558 651168 0 Tile_X10Y2_DIN_SRAM31
rlabel metal2 452558 637560 452558 637560 0 Tile_X10Y2_DIN_SRAM4
rlabel metal2 452558 638064 452558 638064 0 Tile_X10Y2_DIN_SRAM5
rlabel metal2 452558 638568 452558 638568 0 Tile_X10Y2_DIN_SRAM6
rlabel metal2 452558 639072 452558 639072 0 Tile_X10Y2_DIN_SRAM7
rlabel metal2 452558 639576 452558 639576 0 Tile_X10Y2_DIN_SRAM8
rlabel metal2 452558 640080 452558 640080 0 Tile_X10Y2_DIN_SRAM9
rlabel metal2 452558 597744 452558 597744 0 Tile_X10Y2_DOUT_SRAM0
rlabel metal2 452558 598248 452558 598248 0 Tile_X10Y2_DOUT_SRAM1
rlabel metal2 452558 602784 452558 602784 0 Tile_X10Y2_DOUT_SRAM10
rlabel metal2 452558 603288 452558 603288 0 Tile_X10Y2_DOUT_SRAM11
rlabel metal2 452558 603792 452558 603792 0 Tile_X10Y2_DOUT_SRAM12
rlabel metal2 452558 604296 452558 604296 0 Tile_X10Y2_DOUT_SRAM13
rlabel metal2 452558 604800 452558 604800 0 Tile_X10Y2_DOUT_SRAM14
rlabel metal2 452558 605304 452558 605304 0 Tile_X10Y2_DOUT_SRAM15
rlabel metal2 452558 605808 452558 605808 0 Tile_X10Y2_DOUT_SRAM16
rlabel metal2 452558 606312 452558 606312 0 Tile_X10Y2_DOUT_SRAM17
rlabel metal2 452558 606816 452558 606816 0 Tile_X10Y2_DOUT_SRAM18
rlabel metal2 452558 607320 452558 607320 0 Tile_X10Y2_DOUT_SRAM19
rlabel metal2 452558 598752 452558 598752 0 Tile_X10Y2_DOUT_SRAM2
rlabel metal2 452558 607824 452558 607824 0 Tile_X10Y2_DOUT_SRAM20
rlabel metal2 452558 608328 452558 608328 0 Tile_X10Y2_DOUT_SRAM21
rlabel metal2 452558 608832 452558 608832 0 Tile_X10Y2_DOUT_SRAM22
rlabel metal2 452558 609336 452558 609336 0 Tile_X10Y2_DOUT_SRAM23
rlabel metal2 452558 609840 452558 609840 0 Tile_X10Y2_DOUT_SRAM24
rlabel metal2 452558 610344 452558 610344 0 Tile_X10Y2_DOUT_SRAM25
rlabel metal2 452558 610848 452558 610848 0 Tile_X10Y2_DOUT_SRAM26
rlabel metal2 452558 611352 452558 611352 0 Tile_X10Y2_DOUT_SRAM27
rlabel metal2 452558 611856 452558 611856 0 Tile_X10Y2_DOUT_SRAM28
rlabel metal2 452558 612360 452558 612360 0 Tile_X10Y2_DOUT_SRAM29
rlabel metal2 452558 599256 452558 599256 0 Tile_X10Y2_DOUT_SRAM3
rlabel metal2 452558 612864 452558 612864 0 Tile_X10Y2_DOUT_SRAM30
rlabel metal2 452558 613368 452558 613368 0 Tile_X10Y2_DOUT_SRAM31
rlabel metal2 452558 599760 452558 599760 0 Tile_X10Y2_DOUT_SRAM4
rlabel metal2 452558 600264 452558 600264 0 Tile_X10Y2_DOUT_SRAM5
rlabel metal2 452558 600768 452558 600768 0 Tile_X10Y2_DOUT_SRAM6
rlabel metal2 452558 601272 452558 601272 0 Tile_X10Y2_DOUT_SRAM7
rlabel metal2 452558 601776 452558 601776 0 Tile_X10Y2_DOUT_SRAM8
rlabel metal2 452558 602280 452558 602280 0 Tile_X10Y2_DOUT_SRAM9
rlabel metal2 452558 651672 452558 651672 0 Tile_X10Y2_MEN_SRAM
rlabel metal2 452558 652176 452558 652176 0 Tile_X10Y2_REN_SRAM
rlabel metal2 452558 652680 452558 652680 0 Tile_X10Y2_TIE_HIGH_SRAM
rlabel metal2 452558 653184 452558 653184 0 Tile_X10Y2_TIE_LOW_SRAM
rlabel metal2 452558 653688 452558 653688 0 Tile_X10Y2_WEN_SRAM
rlabel metal2 452558 517104 452558 517104 0 Tile_X10Y4_ADDR_SRAM0
rlabel metal2 452558 517608 452558 517608 0 Tile_X10Y4_ADDR_SRAM1
rlabel metal2 452558 518112 452558 518112 0 Tile_X10Y4_ADDR_SRAM2
rlabel metal2 452558 518616 452558 518616 0 Tile_X10Y4_ADDR_SRAM3
rlabel metal2 452558 519120 452558 519120 0 Tile_X10Y4_ADDR_SRAM4
rlabel metal2 452558 519624 452558 519624 0 Tile_X10Y4_ADDR_SRAM5
rlabel metal2 452558 520128 452558 520128 0 Tile_X10Y4_ADDR_SRAM6
rlabel metal2 452558 520632 452558 520632 0 Tile_X10Y4_ADDR_SRAM7
rlabel metal2 452558 521136 452558 521136 0 Tile_X10Y4_ADDR_SRAM8
rlabel metal2 452558 521640 452558 521640 0 Tile_X10Y4_ADDR_SRAM9
rlabel metal2 452558 522144 452558 522144 0 Tile_X10Y4_BM_SRAM0
rlabel metal2 452558 522648 452558 522648 0 Tile_X10Y4_BM_SRAM1
rlabel metal2 452558 527184 452558 527184 0 Tile_X10Y4_BM_SRAM10
rlabel metal2 452558 527688 452558 527688 0 Tile_X10Y4_BM_SRAM11
rlabel metal2 452558 528192 452558 528192 0 Tile_X10Y4_BM_SRAM12
rlabel metal2 452558 528696 452558 528696 0 Tile_X10Y4_BM_SRAM13
rlabel metal2 452558 529200 452558 529200 0 Tile_X10Y4_BM_SRAM14
rlabel metal2 452558 529704 452558 529704 0 Tile_X10Y4_BM_SRAM15
rlabel metal2 452558 530208 452558 530208 0 Tile_X10Y4_BM_SRAM16
rlabel metal2 452558 530712 452558 530712 0 Tile_X10Y4_BM_SRAM17
rlabel metal2 452558 531216 452558 531216 0 Tile_X10Y4_BM_SRAM18
rlabel metal2 452558 531720 452558 531720 0 Tile_X10Y4_BM_SRAM19
rlabel metal2 452558 523152 452558 523152 0 Tile_X10Y4_BM_SRAM2
rlabel metal2 452558 532224 452558 532224 0 Tile_X10Y4_BM_SRAM20
rlabel metal2 452558 532728 452558 532728 0 Tile_X10Y4_BM_SRAM21
rlabel metal2 452558 533232 452558 533232 0 Tile_X10Y4_BM_SRAM22
rlabel metal2 452558 533736 452558 533736 0 Tile_X10Y4_BM_SRAM23
rlabel metal2 452558 534240 452558 534240 0 Tile_X10Y4_BM_SRAM24
rlabel metal2 452558 534744 452558 534744 0 Tile_X10Y4_BM_SRAM25
rlabel metal2 452558 535248 452558 535248 0 Tile_X10Y4_BM_SRAM26
rlabel metal2 452558 535752 452558 535752 0 Tile_X10Y4_BM_SRAM27
rlabel metal2 452558 536256 452558 536256 0 Tile_X10Y4_BM_SRAM28
rlabel metal2 452558 536760 452558 536760 0 Tile_X10Y4_BM_SRAM29
rlabel metal2 452558 523656 452558 523656 0 Tile_X10Y4_BM_SRAM3
rlabel metal2 452558 537264 452558 537264 0 Tile_X10Y4_BM_SRAM30
rlabel metal2 452558 537768 452558 537768 0 Tile_X10Y4_BM_SRAM31
rlabel metal2 452558 524160 452558 524160 0 Tile_X10Y4_BM_SRAM4
rlabel metal2 452558 524664 452558 524664 0 Tile_X10Y4_BM_SRAM5
rlabel metal2 452558 525168 452558 525168 0 Tile_X10Y4_BM_SRAM6
rlabel metal2 452558 525672 452558 525672 0 Tile_X10Y4_BM_SRAM7
rlabel metal2 452558 526176 452558 526176 0 Tile_X10Y4_BM_SRAM8
rlabel metal2 452558 526680 452558 526680 0 Tile_X10Y4_BM_SRAM9
rlabel metal2 452558 538272 452558 538272 0 Tile_X10Y4_CLK_SRAM
rlabel metal2 452558 500472 452558 500472 0 Tile_X10Y4_CONFIGURED_top
rlabel metal2 452558 538776 452558 538776 0 Tile_X10Y4_DIN_SRAM0
rlabel metal2 452558 539280 452558 539280 0 Tile_X10Y4_DIN_SRAM1
rlabel metal2 452558 543816 452558 543816 0 Tile_X10Y4_DIN_SRAM10
rlabel metal2 452558 544320 452558 544320 0 Tile_X10Y4_DIN_SRAM11
rlabel metal2 452558 544824 452558 544824 0 Tile_X10Y4_DIN_SRAM12
rlabel metal2 452558 545328 452558 545328 0 Tile_X10Y4_DIN_SRAM13
rlabel metal2 452558 545832 452558 545832 0 Tile_X10Y4_DIN_SRAM14
rlabel metal2 452558 546336 452558 546336 0 Tile_X10Y4_DIN_SRAM15
rlabel metal2 452558 546840 452558 546840 0 Tile_X10Y4_DIN_SRAM16
rlabel metal2 452558 547344 452558 547344 0 Tile_X10Y4_DIN_SRAM17
rlabel metal2 452558 547848 452558 547848 0 Tile_X10Y4_DIN_SRAM18
rlabel metal2 452558 548352 452558 548352 0 Tile_X10Y4_DIN_SRAM19
rlabel metal2 452558 539784 452558 539784 0 Tile_X10Y4_DIN_SRAM2
rlabel metal2 452558 548856 452558 548856 0 Tile_X10Y4_DIN_SRAM20
rlabel metal2 452558 549360 452558 549360 0 Tile_X10Y4_DIN_SRAM21
rlabel metal2 452558 549864 452558 549864 0 Tile_X10Y4_DIN_SRAM22
rlabel metal2 452558 550368 452558 550368 0 Tile_X10Y4_DIN_SRAM23
rlabel metal2 452558 550872 452558 550872 0 Tile_X10Y4_DIN_SRAM24
rlabel metal2 452558 551376 452558 551376 0 Tile_X10Y4_DIN_SRAM25
rlabel metal2 452558 551880 452558 551880 0 Tile_X10Y4_DIN_SRAM26
rlabel metal2 452558 552384 452558 552384 0 Tile_X10Y4_DIN_SRAM27
rlabel metal2 452558 552888 452558 552888 0 Tile_X10Y4_DIN_SRAM28
rlabel metal2 452558 553392 452558 553392 0 Tile_X10Y4_DIN_SRAM29
rlabel metal2 452558 540288 452558 540288 0 Tile_X10Y4_DIN_SRAM3
rlabel metal2 452558 553896 452558 553896 0 Tile_X10Y4_DIN_SRAM30
rlabel metal2 452558 554400 452558 554400 0 Tile_X10Y4_DIN_SRAM31
rlabel metal2 452558 540792 452558 540792 0 Tile_X10Y4_DIN_SRAM4
rlabel metal2 452558 541296 452558 541296 0 Tile_X10Y4_DIN_SRAM5
rlabel metal2 452558 541800 452558 541800 0 Tile_X10Y4_DIN_SRAM6
rlabel metal2 452558 542304 452558 542304 0 Tile_X10Y4_DIN_SRAM7
rlabel metal2 452558 542808 452558 542808 0 Tile_X10Y4_DIN_SRAM8
rlabel metal2 452558 543312 452558 543312 0 Tile_X10Y4_DIN_SRAM9
rlabel metal2 452558 500976 452558 500976 0 Tile_X10Y4_DOUT_SRAM0
rlabel metal2 452558 501480 452558 501480 0 Tile_X10Y4_DOUT_SRAM1
rlabel metal2 452558 506016 452558 506016 0 Tile_X10Y4_DOUT_SRAM10
rlabel metal2 452558 506520 452558 506520 0 Tile_X10Y4_DOUT_SRAM11
rlabel metal2 452558 507024 452558 507024 0 Tile_X10Y4_DOUT_SRAM12
rlabel metal2 452558 507528 452558 507528 0 Tile_X10Y4_DOUT_SRAM13
rlabel metal2 452558 508032 452558 508032 0 Tile_X10Y4_DOUT_SRAM14
rlabel metal2 452558 508536 452558 508536 0 Tile_X10Y4_DOUT_SRAM15
rlabel metal2 452558 509040 452558 509040 0 Tile_X10Y4_DOUT_SRAM16
rlabel metal2 452558 509544 452558 509544 0 Tile_X10Y4_DOUT_SRAM17
rlabel metal2 452558 510048 452558 510048 0 Tile_X10Y4_DOUT_SRAM18
rlabel metal2 452558 510552 452558 510552 0 Tile_X10Y4_DOUT_SRAM19
rlabel metal2 452558 501984 452558 501984 0 Tile_X10Y4_DOUT_SRAM2
rlabel metal2 452558 511056 452558 511056 0 Tile_X10Y4_DOUT_SRAM20
rlabel metal2 452558 511560 452558 511560 0 Tile_X10Y4_DOUT_SRAM21
rlabel metal2 452558 512064 452558 512064 0 Tile_X10Y4_DOUT_SRAM22
rlabel metal2 452558 512568 452558 512568 0 Tile_X10Y4_DOUT_SRAM23
rlabel metal2 452558 513072 452558 513072 0 Tile_X10Y4_DOUT_SRAM24
rlabel metal2 452558 513576 452558 513576 0 Tile_X10Y4_DOUT_SRAM25
rlabel metal2 452558 514080 452558 514080 0 Tile_X10Y4_DOUT_SRAM26
rlabel metal2 452558 514584 452558 514584 0 Tile_X10Y4_DOUT_SRAM27
rlabel metal2 452558 515088 452558 515088 0 Tile_X10Y4_DOUT_SRAM28
rlabel metal2 452558 515592 452558 515592 0 Tile_X10Y4_DOUT_SRAM29
rlabel metal2 452558 502488 452558 502488 0 Tile_X10Y4_DOUT_SRAM3
rlabel metal2 452558 516096 452558 516096 0 Tile_X10Y4_DOUT_SRAM30
rlabel metal2 452558 516600 452558 516600 0 Tile_X10Y4_DOUT_SRAM31
rlabel metal2 452558 502992 452558 502992 0 Tile_X10Y4_DOUT_SRAM4
rlabel metal2 452558 503496 452558 503496 0 Tile_X10Y4_DOUT_SRAM5
rlabel metal2 452558 504000 452558 504000 0 Tile_X10Y4_DOUT_SRAM6
rlabel metal2 452558 504504 452558 504504 0 Tile_X10Y4_DOUT_SRAM7
rlabel metal2 452558 505008 452558 505008 0 Tile_X10Y4_DOUT_SRAM8
rlabel metal2 452558 505512 452558 505512 0 Tile_X10Y4_DOUT_SRAM9
rlabel metal2 452558 554904 452558 554904 0 Tile_X10Y4_MEN_SRAM
rlabel metal2 452558 555408 452558 555408 0 Tile_X10Y4_REN_SRAM
rlabel metal2 452558 555912 452558 555912 0 Tile_X10Y4_TIE_HIGH_SRAM
rlabel metal2 452558 556416 452558 556416 0 Tile_X10Y4_TIE_LOW_SRAM
rlabel metal2 452558 556920 452558 556920 0 Tile_X10Y4_WEN_SRAM
rlabel metal2 452558 420336 452558 420336 0 Tile_X10Y6_ADDR_SRAM0
rlabel metal2 452558 420840 452558 420840 0 Tile_X10Y6_ADDR_SRAM1
rlabel metal2 452558 421344 452558 421344 0 Tile_X10Y6_ADDR_SRAM2
rlabel metal2 452558 421848 452558 421848 0 Tile_X10Y6_ADDR_SRAM3
rlabel metal2 452558 422352 452558 422352 0 Tile_X10Y6_ADDR_SRAM4
rlabel metal2 452558 422856 452558 422856 0 Tile_X10Y6_ADDR_SRAM5
rlabel metal2 452558 423360 452558 423360 0 Tile_X10Y6_ADDR_SRAM6
rlabel metal2 452558 423864 452558 423864 0 Tile_X10Y6_ADDR_SRAM7
rlabel metal2 452558 424368 452558 424368 0 Tile_X10Y6_ADDR_SRAM8
rlabel metal2 452558 424872 452558 424872 0 Tile_X10Y6_ADDR_SRAM9
rlabel metal2 452558 425376 452558 425376 0 Tile_X10Y6_BM_SRAM0
rlabel metal2 452558 425880 452558 425880 0 Tile_X10Y6_BM_SRAM1
rlabel metal2 452558 430416 452558 430416 0 Tile_X10Y6_BM_SRAM10
rlabel metal2 452558 430920 452558 430920 0 Tile_X10Y6_BM_SRAM11
rlabel metal2 452558 431424 452558 431424 0 Tile_X10Y6_BM_SRAM12
rlabel metal2 452558 431928 452558 431928 0 Tile_X10Y6_BM_SRAM13
rlabel metal2 452558 432432 452558 432432 0 Tile_X10Y6_BM_SRAM14
rlabel metal2 452558 432936 452558 432936 0 Tile_X10Y6_BM_SRAM15
rlabel metal2 452558 433440 452558 433440 0 Tile_X10Y6_BM_SRAM16
rlabel metal2 452558 433944 452558 433944 0 Tile_X10Y6_BM_SRAM17
rlabel metal2 452558 434448 452558 434448 0 Tile_X10Y6_BM_SRAM18
rlabel metal2 452558 434952 452558 434952 0 Tile_X10Y6_BM_SRAM19
rlabel metal2 452558 426384 452558 426384 0 Tile_X10Y6_BM_SRAM2
rlabel metal2 452558 435456 452558 435456 0 Tile_X10Y6_BM_SRAM20
rlabel metal2 452558 435960 452558 435960 0 Tile_X10Y6_BM_SRAM21
rlabel metal2 452558 436464 452558 436464 0 Tile_X10Y6_BM_SRAM22
rlabel metal2 452558 436968 452558 436968 0 Tile_X10Y6_BM_SRAM23
rlabel metal2 452558 437472 452558 437472 0 Tile_X10Y6_BM_SRAM24
rlabel metal2 452558 437976 452558 437976 0 Tile_X10Y6_BM_SRAM25
rlabel metal2 452558 438480 452558 438480 0 Tile_X10Y6_BM_SRAM26
rlabel metal2 452558 438984 452558 438984 0 Tile_X10Y6_BM_SRAM27
rlabel metal2 452558 439488 452558 439488 0 Tile_X10Y6_BM_SRAM28
rlabel metal2 452558 439992 452558 439992 0 Tile_X10Y6_BM_SRAM29
rlabel metal2 452558 426888 452558 426888 0 Tile_X10Y6_BM_SRAM3
rlabel metal2 452558 440496 452558 440496 0 Tile_X10Y6_BM_SRAM30
rlabel metal2 452558 441000 452558 441000 0 Tile_X10Y6_BM_SRAM31
rlabel metal2 452558 427392 452558 427392 0 Tile_X10Y6_BM_SRAM4
rlabel metal2 452558 427896 452558 427896 0 Tile_X10Y6_BM_SRAM5
rlabel metal2 452558 428400 452558 428400 0 Tile_X10Y6_BM_SRAM6
rlabel metal2 452558 428904 452558 428904 0 Tile_X10Y6_BM_SRAM7
rlabel metal2 452558 429408 452558 429408 0 Tile_X10Y6_BM_SRAM8
rlabel metal2 452558 429912 452558 429912 0 Tile_X10Y6_BM_SRAM9
rlabel metal2 452558 441504 452558 441504 0 Tile_X10Y6_CLK_SRAM
rlabel metal2 452558 403704 452558 403704 0 Tile_X10Y6_CONFIGURED_top
rlabel metal2 452558 442008 452558 442008 0 Tile_X10Y6_DIN_SRAM0
rlabel metal2 452558 442512 452558 442512 0 Tile_X10Y6_DIN_SRAM1
rlabel metal2 452558 447048 452558 447048 0 Tile_X10Y6_DIN_SRAM10
rlabel metal2 452558 447552 452558 447552 0 Tile_X10Y6_DIN_SRAM11
rlabel metal2 452558 448056 452558 448056 0 Tile_X10Y6_DIN_SRAM12
rlabel metal2 452558 448560 452558 448560 0 Tile_X10Y6_DIN_SRAM13
rlabel metal2 452558 449064 452558 449064 0 Tile_X10Y6_DIN_SRAM14
rlabel metal2 452558 449568 452558 449568 0 Tile_X10Y6_DIN_SRAM15
rlabel metal2 452558 450072 452558 450072 0 Tile_X10Y6_DIN_SRAM16
rlabel metal2 452558 450576 452558 450576 0 Tile_X10Y6_DIN_SRAM17
rlabel metal2 452558 451080 452558 451080 0 Tile_X10Y6_DIN_SRAM18
rlabel metal2 452558 451584 452558 451584 0 Tile_X10Y6_DIN_SRAM19
rlabel metal2 452558 443016 452558 443016 0 Tile_X10Y6_DIN_SRAM2
rlabel metal2 452558 452088 452558 452088 0 Tile_X10Y6_DIN_SRAM20
rlabel metal2 452558 452592 452558 452592 0 Tile_X10Y6_DIN_SRAM21
rlabel metal2 452558 453096 452558 453096 0 Tile_X10Y6_DIN_SRAM22
rlabel metal2 452558 453600 452558 453600 0 Tile_X10Y6_DIN_SRAM23
rlabel metal2 452558 454104 452558 454104 0 Tile_X10Y6_DIN_SRAM24
rlabel metal2 452558 454608 452558 454608 0 Tile_X10Y6_DIN_SRAM25
rlabel metal2 452558 455112 452558 455112 0 Tile_X10Y6_DIN_SRAM26
rlabel metal2 452558 455616 452558 455616 0 Tile_X10Y6_DIN_SRAM27
rlabel metal2 452558 456120 452558 456120 0 Tile_X10Y6_DIN_SRAM28
rlabel metal2 452558 456624 452558 456624 0 Tile_X10Y6_DIN_SRAM29
rlabel metal2 452558 443520 452558 443520 0 Tile_X10Y6_DIN_SRAM3
rlabel metal2 452558 457128 452558 457128 0 Tile_X10Y6_DIN_SRAM30
rlabel metal2 452558 457632 452558 457632 0 Tile_X10Y6_DIN_SRAM31
rlabel metal2 452558 444024 452558 444024 0 Tile_X10Y6_DIN_SRAM4
rlabel metal2 452558 444528 452558 444528 0 Tile_X10Y6_DIN_SRAM5
rlabel metal2 452558 445032 452558 445032 0 Tile_X10Y6_DIN_SRAM6
rlabel metal2 452558 445536 452558 445536 0 Tile_X10Y6_DIN_SRAM7
rlabel metal2 452558 446040 452558 446040 0 Tile_X10Y6_DIN_SRAM8
rlabel metal2 452558 446544 452558 446544 0 Tile_X10Y6_DIN_SRAM9
rlabel metal2 452558 404208 452558 404208 0 Tile_X10Y6_DOUT_SRAM0
rlabel metal2 452558 404712 452558 404712 0 Tile_X10Y6_DOUT_SRAM1
rlabel metal2 452558 409248 452558 409248 0 Tile_X10Y6_DOUT_SRAM10
rlabel metal2 452558 409752 452558 409752 0 Tile_X10Y6_DOUT_SRAM11
rlabel metal2 452558 410256 452558 410256 0 Tile_X10Y6_DOUT_SRAM12
rlabel metal2 452558 410760 452558 410760 0 Tile_X10Y6_DOUT_SRAM13
rlabel metal2 452558 411264 452558 411264 0 Tile_X10Y6_DOUT_SRAM14
rlabel metal2 452558 411768 452558 411768 0 Tile_X10Y6_DOUT_SRAM15
rlabel metal2 452558 412272 452558 412272 0 Tile_X10Y6_DOUT_SRAM16
rlabel metal2 452558 412776 452558 412776 0 Tile_X10Y6_DOUT_SRAM17
rlabel metal2 452558 413280 452558 413280 0 Tile_X10Y6_DOUT_SRAM18
rlabel metal2 452558 413784 452558 413784 0 Tile_X10Y6_DOUT_SRAM19
rlabel metal2 452558 405216 452558 405216 0 Tile_X10Y6_DOUT_SRAM2
rlabel metal2 452558 414288 452558 414288 0 Tile_X10Y6_DOUT_SRAM20
rlabel metal2 452558 414792 452558 414792 0 Tile_X10Y6_DOUT_SRAM21
rlabel metal2 452558 415296 452558 415296 0 Tile_X10Y6_DOUT_SRAM22
rlabel metal2 452558 415800 452558 415800 0 Tile_X10Y6_DOUT_SRAM23
rlabel metal2 452558 416304 452558 416304 0 Tile_X10Y6_DOUT_SRAM24
rlabel metal2 452558 416808 452558 416808 0 Tile_X10Y6_DOUT_SRAM25
rlabel metal2 452558 417312 452558 417312 0 Tile_X10Y6_DOUT_SRAM26
rlabel metal2 452558 417816 452558 417816 0 Tile_X10Y6_DOUT_SRAM27
rlabel metal2 452558 418320 452558 418320 0 Tile_X10Y6_DOUT_SRAM28
rlabel metal2 452558 418824 452558 418824 0 Tile_X10Y6_DOUT_SRAM29
rlabel metal2 452558 405720 452558 405720 0 Tile_X10Y6_DOUT_SRAM3
rlabel metal2 452558 419328 452558 419328 0 Tile_X10Y6_DOUT_SRAM30
rlabel metal2 452558 419832 452558 419832 0 Tile_X10Y6_DOUT_SRAM31
rlabel metal2 452558 406224 452558 406224 0 Tile_X10Y6_DOUT_SRAM4
rlabel metal2 452558 406728 452558 406728 0 Tile_X10Y6_DOUT_SRAM5
rlabel metal2 452558 407232 452558 407232 0 Tile_X10Y6_DOUT_SRAM6
rlabel metal2 452558 407736 452558 407736 0 Tile_X10Y6_DOUT_SRAM7
rlabel metal2 452558 408240 452558 408240 0 Tile_X10Y6_DOUT_SRAM8
rlabel metal2 452558 408744 452558 408744 0 Tile_X10Y6_DOUT_SRAM9
rlabel metal2 452558 458136 452558 458136 0 Tile_X10Y6_MEN_SRAM
rlabel metal2 452558 458640 452558 458640 0 Tile_X10Y6_REN_SRAM
rlabel metal2 452558 459144 452558 459144 0 Tile_X10Y6_TIE_HIGH_SRAM
rlabel metal2 452558 459648 452558 459648 0 Tile_X10Y6_TIE_LOW_SRAM
rlabel metal2 452558 460152 452558 460152 0 Tile_X10Y6_WEN_SRAM
rlabel metal2 452558 323568 452558 323568 0 Tile_X10Y8_ADDR_SRAM0
rlabel metal2 452558 324072 452558 324072 0 Tile_X10Y8_ADDR_SRAM1
rlabel metal2 452558 324576 452558 324576 0 Tile_X10Y8_ADDR_SRAM2
rlabel metal2 452558 325080 452558 325080 0 Tile_X10Y8_ADDR_SRAM3
rlabel metal2 452558 325584 452558 325584 0 Tile_X10Y8_ADDR_SRAM4
rlabel metal2 452558 326088 452558 326088 0 Tile_X10Y8_ADDR_SRAM5
rlabel metal2 452558 326592 452558 326592 0 Tile_X10Y8_ADDR_SRAM6
rlabel metal2 452558 327096 452558 327096 0 Tile_X10Y8_ADDR_SRAM7
rlabel metal2 452558 327600 452558 327600 0 Tile_X10Y8_ADDR_SRAM8
rlabel metal2 452558 328104 452558 328104 0 Tile_X10Y8_ADDR_SRAM9
rlabel metal2 452558 328608 452558 328608 0 Tile_X10Y8_BM_SRAM0
rlabel metal2 452558 329112 452558 329112 0 Tile_X10Y8_BM_SRAM1
rlabel metal2 452558 333648 452558 333648 0 Tile_X10Y8_BM_SRAM10
rlabel metal2 452558 334152 452558 334152 0 Tile_X10Y8_BM_SRAM11
rlabel metal2 452558 334656 452558 334656 0 Tile_X10Y8_BM_SRAM12
rlabel metal2 452558 335160 452558 335160 0 Tile_X10Y8_BM_SRAM13
rlabel metal2 452558 335664 452558 335664 0 Tile_X10Y8_BM_SRAM14
rlabel metal2 452558 336168 452558 336168 0 Tile_X10Y8_BM_SRAM15
rlabel metal2 452558 336672 452558 336672 0 Tile_X10Y8_BM_SRAM16
rlabel metal2 452558 337176 452558 337176 0 Tile_X10Y8_BM_SRAM17
rlabel metal2 452558 337680 452558 337680 0 Tile_X10Y8_BM_SRAM18
rlabel metal2 452558 338184 452558 338184 0 Tile_X10Y8_BM_SRAM19
rlabel metal2 452558 329616 452558 329616 0 Tile_X10Y8_BM_SRAM2
rlabel metal2 452558 338688 452558 338688 0 Tile_X10Y8_BM_SRAM20
rlabel metal2 452558 339192 452558 339192 0 Tile_X10Y8_BM_SRAM21
rlabel metal2 452558 339696 452558 339696 0 Tile_X10Y8_BM_SRAM22
rlabel metal2 452558 340200 452558 340200 0 Tile_X10Y8_BM_SRAM23
rlabel metal2 452558 340704 452558 340704 0 Tile_X10Y8_BM_SRAM24
rlabel metal2 452558 341208 452558 341208 0 Tile_X10Y8_BM_SRAM25
rlabel metal2 452558 341712 452558 341712 0 Tile_X10Y8_BM_SRAM26
rlabel metal2 452558 342216 452558 342216 0 Tile_X10Y8_BM_SRAM27
rlabel metal2 452558 342720 452558 342720 0 Tile_X10Y8_BM_SRAM28
rlabel metal2 452558 343224 452558 343224 0 Tile_X10Y8_BM_SRAM29
rlabel metal2 452558 330120 452558 330120 0 Tile_X10Y8_BM_SRAM3
rlabel metal2 452558 343728 452558 343728 0 Tile_X10Y8_BM_SRAM30
rlabel metal2 452558 344232 452558 344232 0 Tile_X10Y8_BM_SRAM31
rlabel metal2 452558 330624 452558 330624 0 Tile_X10Y8_BM_SRAM4
rlabel metal2 452558 331128 452558 331128 0 Tile_X10Y8_BM_SRAM5
rlabel metal2 452558 331632 452558 331632 0 Tile_X10Y8_BM_SRAM6
rlabel metal2 452558 332136 452558 332136 0 Tile_X10Y8_BM_SRAM7
rlabel metal2 452558 332640 452558 332640 0 Tile_X10Y8_BM_SRAM8
rlabel metal2 452558 333144 452558 333144 0 Tile_X10Y8_BM_SRAM9
rlabel metal2 452558 344736 452558 344736 0 Tile_X10Y8_CLK_SRAM
rlabel metal2 452558 306936 452558 306936 0 Tile_X10Y8_CONFIGURED_top
rlabel metal2 452558 345240 452558 345240 0 Tile_X10Y8_DIN_SRAM0
rlabel metal2 452558 345744 452558 345744 0 Tile_X10Y8_DIN_SRAM1
rlabel metal2 452558 350280 452558 350280 0 Tile_X10Y8_DIN_SRAM10
rlabel metal2 452558 350784 452558 350784 0 Tile_X10Y8_DIN_SRAM11
rlabel metal2 452558 351288 452558 351288 0 Tile_X10Y8_DIN_SRAM12
rlabel metal2 452558 351792 452558 351792 0 Tile_X10Y8_DIN_SRAM13
rlabel metal2 452558 352296 452558 352296 0 Tile_X10Y8_DIN_SRAM14
rlabel metal2 452558 352800 452558 352800 0 Tile_X10Y8_DIN_SRAM15
rlabel metal2 452558 353304 452558 353304 0 Tile_X10Y8_DIN_SRAM16
rlabel metal2 452558 353808 452558 353808 0 Tile_X10Y8_DIN_SRAM17
rlabel metal2 452558 354312 452558 354312 0 Tile_X10Y8_DIN_SRAM18
rlabel metal2 452558 354816 452558 354816 0 Tile_X10Y8_DIN_SRAM19
rlabel metal2 452558 346248 452558 346248 0 Tile_X10Y8_DIN_SRAM2
rlabel metal2 452558 355320 452558 355320 0 Tile_X10Y8_DIN_SRAM20
rlabel metal2 452558 355824 452558 355824 0 Tile_X10Y8_DIN_SRAM21
rlabel metal2 452558 356328 452558 356328 0 Tile_X10Y8_DIN_SRAM22
rlabel metal2 452558 356832 452558 356832 0 Tile_X10Y8_DIN_SRAM23
rlabel metal2 452558 357336 452558 357336 0 Tile_X10Y8_DIN_SRAM24
rlabel metal2 452558 357840 452558 357840 0 Tile_X10Y8_DIN_SRAM25
rlabel metal2 452558 358344 452558 358344 0 Tile_X10Y8_DIN_SRAM26
rlabel metal2 452558 358848 452558 358848 0 Tile_X10Y8_DIN_SRAM27
rlabel metal2 452558 359352 452558 359352 0 Tile_X10Y8_DIN_SRAM28
rlabel metal2 452558 359856 452558 359856 0 Tile_X10Y8_DIN_SRAM29
rlabel metal2 452558 346752 452558 346752 0 Tile_X10Y8_DIN_SRAM3
rlabel metal2 452558 360360 452558 360360 0 Tile_X10Y8_DIN_SRAM30
rlabel metal2 452558 360864 452558 360864 0 Tile_X10Y8_DIN_SRAM31
rlabel metal2 452558 347256 452558 347256 0 Tile_X10Y8_DIN_SRAM4
rlabel metal2 452558 347760 452558 347760 0 Tile_X10Y8_DIN_SRAM5
rlabel metal2 452558 348264 452558 348264 0 Tile_X10Y8_DIN_SRAM6
rlabel metal2 452558 348768 452558 348768 0 Tile_X10Y8_DIN_SRAM7
rlabel metal2 452558 349272 452558 349272 0 Tile_X10Y8_DIN_SRAM8
rlabel metal2 452558 349776 452558 349776 0 Tile_X10Y8_DIN_SRAM9
rlabel metal2 452558 307440 452558 307440 0 Tile_X10Y8_DOUT_SRAM0
rlabel metal2 452558 307944 452558 307944 0 Tile_X10Y8_DOUT_SRAM1
rlabel metal2 452558 312480 452558 312480 0 Tile_X10Y8_DOUT_SRAM10
rlabel metal2 452558 312984 452558 312984 0 Tile_X10Y8_DOUT_SRAM11
rlabel metal2 452558 313488 452558 313488 0 Tile_X10Y8_DOUT_SRAM12
rlabel metal2 452558 313992 452558 313992 0 Tile_X10Y8_DOUT_SRAM13
rlabel metal2 452558 314496 452558 314496 0 Tile_X10Y8_DOUT_SRAM14
rlabel metal2 452558 315000 452558 315000 0 Tile_X10Y8_DOUT_SRAM15
rlabel metal2 452558 315504 452558 315504 0 Tile_X10Y8_DOUT_SRAM16
rlabel metal2 452558 316008 452558 316008 0 Tile_X10Y8_DOUT_SRAM17
rlabel metal2 452558 316512 452558 316512 0 Tile_X10Y8_DOUT_SRAM18
rlabel metal2 452558 317016 452558 317016 0 Tile_X10Y8_DOUT_SRAM19
rlabel metal2 452558 308448 452558 308448 0 Tile_X10Y8_DOUT_SRAM2
rlabel metal2 452558 317520 452558 317520 0 Tile_X10Y8_DOUT_SRAM20
rlabel metal2 452558 318024 452558 318024 0 Tile_X10Y8_DOUT_SRAM21
rlabel metal2 452558 318528 452558 318528 0 Tile_X10Y8_DOUT_SRAM22
rlabel metal2 452558 319032 452558 319032 0 Tile_X10Y8_DOUT_SRAM23
rlabel metal2 452558 319536 452558 319536 0 Tile_X10Y8_DOUT_SRAM24
rlabel metal2 452558 320040 452558 320040 0 Tile_X10Y8_DOUT_SRAM25
rlabel metal2 452558 320544 452558 320544 0 Tile_X10Y8_DOUT_SRAM26
rlabel metal2 452558 321048 452558 321048 0 Tile_X10Y8_DOUT_SRAM27
rlabel metal2 452558 321552 452558 321552 0 Tile_X10Y8_DOUT_SRAM28
rlabel metal2 452558 322056 452558 322056 0 Tile_X10Y8_DOUT_SRAM29
rlabel metal2 452558 308952 452558 308952 0 Tile_X10Y8_DOUT_SRAM3
rlabel metal2 452558 322560 452558 322560 0 Tile_X10Y8_DOUT_SRAM30
rlabel metal2 452558 323064 452558 323064 0 Tile_X10Y8_DOUT_SRAM31
rlabel metal2 452558 309456 452558 309456 0 Tile_X10Y8_DOUT_SRAM4
rlabel metal2 452558 309960 452558 309960 0 Tile_X10Y8_DOUT_SRAM5
rlabel metal2 452558 310464 452558 310464 0 Tile_X10Y8_DOUT_SRAM6
rlabel metal2 452558 310968 452558 310968 0 Tile_X10Y8_DOUT_SRAM7
rlabel metal2 452558 311472 452558 311472 0 Tile_X10Y8_DOUT_SRAM8
rlabel metal2 452558 311976 452558 311976 0 Tile_X10Y8_DOUT_SRAM9
rlabel metal2 452558 361368 452558 361368 0 Tile_X10Y8_MEN_SRAM
rlabel metal2 452558 361872 452558 361872 0 Tile_X10Y8_REN_SRAM
rlabel metal2 452558 362376 452558 362376 0 Tile_X10Y8_TIE_HIGH_SRAM
rlabel metal2 452558 362880 452558 362880 0 Tile_X10Y8_TIE_LOW_SRAM
rlabel metal2 452558 363384 452558 363384 0 Tile_X10Y8_WEN_SRAM
rlabel metal3 18528 702254 18528 702254 0 Tile_X1Y0_A_I_top
rlabel metal3 17376 702254 17376 702254 0 Tile_X1Y0_A_O_top
rlabel metal3 19680 702254 19680 702254 0 Tile_X1Y0_A_T_top
rlabel metal3 24288 702254 24288 702254 0 Tile_X1Y0_A_config_C_bit0
rlabel metal3 25440 702254 25440 702254 0 Tile_X1Y0_A_config_C_bit1
rlabel metal3 26592 702254 26592 702254 0 Tile_X1Y0_A_config_C_bit2
rlabel metal3 27744 702254 27744 702254 0 Tile_X1Y0_A_config_C_bit3
rlabel metal3 21984 702254 21984 702254 0 Tile_X1Y0_B_I_top
rlabel metal3 20832 702254 20832 702254 0 Tile_X1Y0_B_O_top
rlabel metal3 23136 702254 23136 702254 0 Tile_X1Y0_B_T_top
rlabel metal3 28896 702254 28896 702254 0 Tile_X1Y0_B_config_C_bit0
rlabel metal3 30048 702254 30048 702254 0 Tile_X1Y0_B_config_C_bit1
rlabel metal3 31200 702254 31200 702254 0 Tile_X1Y0_B_config_C_bit2
rlabel metal3 32352 702254 32352 702254 0 Tile_X1Y0_B_config_C_bit3
rlabel metal3 64896 702254 64896 702254 0 Tile_X2Y0_A_I_top
rlabel metal3 63744 702254 63744 702254 0 Tile_X2Y0_A_O_top
rlabel metal3 66048 702254 66048 702254 0 Tile_X2Y0_A_T_top
rlabel metal3 70656 702254 70656 702254 0 Tile_X2Y0_A_config_C_bit0
rlabel metal3 71808 702254 71808 702254 0 Tile_X2Y0_A_config_C_bit1
rlabel metal3 72960 702254 72960 702254 0 Tile_X2Y0_A_config_C_bit2
rlabel metal3 74112 702254 74112 702254 0 Tile_X2Y0_A_config_C_bit3
rlabel metal3 68352 702254 68352 702254 0 Tile_X2Y0_B_I_top
rlabel metal3 67200 702254 67200 702254 0 Tile_X2Y0_B_O_top
rlabel metal3 69504 702254 69504 702254 0 Tile_X2Y0_B_T_top
rlabel metal3 75264 702254 75264 702254 0 Tile_X2Y0_B_config_C_bit0
rlabel metal3 76416 702254 76416 702254 0 Tile_X2Y0_B_config_C_bit1
rlabel metal3 77568 702254 77568 702254 0 Tile_X2Y0_B_config_C_bit2
rlabel metal3 78720 702254 78720 702254 0 Tile_X2Y0_B_config_C_bit3
rlabel metal3 65664 454 65664 454 0 Tile_X2Y15_BOOT_top
rlabel metal3 62592 454 62592 454 0 Tile_X2Y15_CONFIGURED_top
rlabel metal3 64128 454 64128 454 0 Tile_X2Y15_RESET_top
rlabel metal3 67200 454 67200 454 0 Tile_X2Y15_SLOT_top0
rlabel metal3 68736 454 68736 454 0 Tile_X2Y15_SLOT_top1
rlabel metal3 70272 454 70272 454 0 Tile_X2Y15_SLOT_top2
rlabel metal3 71808 454 71808 454 0 Tile_X2Y15_SLOT_top3
rlabel metal3 108000 454 108000 454 0 Tile_X3Y15_CONFIGURED_top
rlabel metal3 109728 454 109728 454 0 Tile_X3Y15_IRQ_top0
rlabel metal3 111456 454 111456 454 0 Tile_X3Y15_IRQ_top1
rlabel metal3 113184 454 113184 454 0 Tile_X3Y15_IRQ_top2
rlabel metal3 114912 454 114912 454 0 Tile_X3Y15_IRQ_top3
rlabel metal3 221664 454 221664 454 0 Tile_X5Y15_I_top0
rlabel metal3 222432 454 222432 454 0 Tile_X5Y15_I_top1
rlabel metal3 229344 454 229344 454 0 Tile_X5Y15_I_top10
rlabel metal3 230112 454 230112 454 0 Tile_X5Y15_I_top11
rlabel metal3 230880 454 230880 454 0 Tile_X5Y15_I_top12
rlabel metal3 231648 454 231648 454 0 Tile_X5Y15_I_top13
rlabel metal3 232416 454 232416 454 0 Tile_X5Y15_I_top14
rlabel metal3 233184 454 233184 454 0 Tile_X5Y15_I_top15
rlabel metal3 223200 454 223200 454 0 Tile_X5Y15_I_top2
rlabel metal3 223968 454 223968 454 0 Tile_X5Y15_I_top3
rlabel metal3 224736 454 224736 454 0 Tile_X5Y15_I_top4
rlabel metal3 225504 454 225504 454 0 Tile_X5Y15_I_top5
rlabel metal3 226272 454 226272 454 0 Tile_X5Y15_I_top6
rlabel metal3 227040 454 227040 454 0 Tile_X5Y15_I_top7
rlabel metal3 227808 454 227808 454 0 Tile_X5Y15_I_top8
rlabel metal3 228576 454 228576 454 0 Tile_X5Y15_I_top9
rlabel metal3 209376 454 209376 454 0 Tile_X5Y15_O_top0
rlabel metal3 210144 454 210144 454 0 Tile_X5Y15_O_top1
rlabel metal3 217056 454 217056 454 0 Tile_X5Y15_O_top10
rlabel metal3 217824 454 217824 454 0 Tile_X5Y15_O_top11
rlabel metal3 218592 454 218592 454 0 Tile_X5Y15_O_top12
rlabel metal3 219360 454 219360 454 0 Tile_X5Y15_O_top13
rlabel metal3 220128 454 220128 454 0 Tile_X5Y15_O_top14
rlabel metal3 220896 454 220896 454 0 Tile_X5Y15_O_top15
rlabel metal3 210912 454 210912 454 0 Tile_X5Y15_O_top2
rlabel metal3 211680 454 211680 454 0 Tile_X5Y15_O_top3
rlabel metal3 212448 454 212448 454 0 Tile_X5Y15_O_top4
rlabel metal3 213216 454 213216 454 0 Tile_X5Y15_O_top5
rlabel metal3 213984 454 213984 454 0 Tile_X5Y15_O_top6
rlabel metal3 214752 454 214752 454 0 Tile_X5Y15_O_top7
rlabel metal3 215520 454 215520 454 0 Tile_X5Y15_O_top8
rlabel metal3 216288 454 216288 454 0 Tile_X5Y15_O_top9
rlabel metal3 268032 454 268032 454 0 Tile_X6Y15_I_top0
rlabel metal3 268800 454 268800 454 0 Tile_X6Y15_I_top1
rlabel metal3 275712 454 275712 454 0 Tile_X6Y15_I_top10
rlabel metal3 276480 454 276480 454 0 Tile_X6Y15_I_top11
rlabel metal3 277248 454 277248 454 0 Tile_X6Y15_I_top12
rlabel metal3 278016 454 278016 454 0 Tile_X6Y15_I_top13
rlabel metal3 278784 454 278784 454 0 Tile_X6Y15_I_top14
rlabel metal3 279552 454 279552 454 0 Tile_X6Y15_I_top15
rlabel metal3 269568 454 269568 454 0 Tile_X6Y15_I_top2
rlabel metal3 270336 454 270336 454 0 Tile_X6Y15_I_top3
rlabel metal3 271104 454 271104 454 0 Tile_X6Y15_I_top4
rlabel metal3 271872 454 271872 454 0 Tile_X6Y15_I_top5
rlabel metal3 272640 454 272640 454 0 Tile_X6Y15_I_top6
rlabel metal3 273408 454 273408 454 0 Tile_X6Y15_I_top7
rlabel metal3 274176 454 274176 454 0 Tile_X6Y15_I_top8
rlabel metal3 274944 454 274944 454 0 Tile_X6Y15_I_top9
rlabel metal3 255744 454 255744 454 0 Tile_X6Y15_O_top0
rlabel metal3 256512 454 256512 454 0 Tile_X6Y15_O_top1
rlabel metal3 263424 454 263424 454 0 Tile_X6Y15_O_top10
rlabel metal3 264192 454 264192 454 0 Tile_X6Y15_O_top11
rlabel metal3 264960 454 264960 454 0 Tile_X6Y15_O_top12
rlabel metal3 265728 454 265728 454 0 Tile_X6Y15_O_top13
rlabel metal3 266496 454 266496 454 0 Tile_X6Y15_O_top14
rlabel metal3 267264 454 267264 454 0 Tile_X6Y15_O_top15
rlabel metal3 257280 454 257280 454 0 Tile_X6Y15_O_top2
rlabel metal3 258048 454 258048 454 0 Tile_X6Y15_O_top3
rlabel metal3 258816 454 258816 454 0 Tile_X6Y15_O_top4
rlabel metal3 259584 454 259584 454 0 Tile_X6Y15_O_top5
rlabel metal3 260352 454 260352 454 0 Tile_X6Y15_O_top6
rlabel metal3 261120 454 261120 454 0 Tile_X6Y15_O_top7
rlabel metal3 261888 454 261888 454 0 Tile_X6Y15_O_top8
rlabel metal3 262656 454 262656 454 0 Tile_X6Y15_O_top9
rlabel metal3 353664 454 353664 454 0 Tile_X8Y15_I_top0
rlabel metal3 354432 454 354432 454 0 Tile_X8Y15_I_top1
rlabel metal3 361344 454 361344 454 0 Tile_X8Y15_I_top10
rlabel metal3 362112 454 362112 454 0 Tile_X8Y15_I_top11
rlabel metal3 362880 454 362880 454 0 Tile_X8Y15_I_top12
rlabel metal3 363648 454 363648 454 0 Tile_X8Y15_I_top13
rlabel metal3 364416 454 364416 454 0 Tile_X8Y15_I_top14
rlabel metal3 365184 454 365184 454 0 Tile_X8Y15_I_top15
rlabel metal3 355200 454 355200 454 0 Tile_X8Y15_I_top2
rlabel metal3 355968 454 355968 454 0 Tile_X8Y15_I_top3
rlabel metal3 356736 454 356736 454 0 Tile_X8Y15_I_top4
rlabel metal3 357504 454 357504 454 0 Tile_X8Y15_I_top5
rlabel metal3 358272 454 358272 454 0 Tile_X8Y15_I_top6
rlabel metal3 359040 454 359040 454 0 Tile_X8Y15_I_top7
rlabel metal3 359808 454 359808 454 0 Tile_X8Y15_I_top8
rlabel metal3 360576 454 360576 454 0 Tile_X8Y15_I_top9
rlabel metal3 341376 454 341376 454 0 Tile_X8Y15_O_top0
rlabel metal3 342144 454 342144 454 0 Tile_X8Y15_O_top1
rlabel metal3 349056 454 349056 454 0 Tile_X8Y15_O_top10
rlabel metal3 349824 454 349824 454 0 Tile_X8Y15_O_top11
rlabel metal3 350592 454 350592 454 0 Tile_X8Y15_O_top12
rlabel metal3 351360 454 351360 454 0 Tile_X8Y15_O_top13
rlabel metal3 352128 454 352128 454 0 Tile_X8Y15_O_top14
rlabel metal3 352896 454 352896 454 0 Tile_X8Y15_O_top15
rlabel metal3 342912 454 342912 454 0 Tile_X8Y15_O_top2
rlabel metal3 343680 454 343680 454 0 Tile_X8Y15_O_top3
rlabel metal3 344448 454 344448 454 0 Tile_X8Y15_O_top4
rlabel metal3 345216 454 345216 454 0 Tile_X8Y15_O_top5
rlabel metal3 345984 454 345984 454 0 Tile_X8Y15_O_top6
rlabel metal3 346752 454 346752 454 0 Tile_X8Y15_O_top7
rlabel metal3 347520 454 347520 454 0 Tile_X8Y15_O_top8
rlabel metal3 348288 454 348288 454 0 Tile_X8Y15_O_top9
rlabel metal3 400032 454 400032 454 0 Tile_X9Y15_I_top0
rlabel metal3 400800 454 400800 454 0 Tile_X9Y15_I_top1
rlabel metal3 407712 454 407712 454 0 Tile_X9Y15_I_top10
rlabel metal3 408480 454 408480 454 0 Tile_X9Y15_I_top11
rlabel metal3 409248 454 409248 454 0 Tile_X9Y15_I_top12
rlabel metal3 410016 454 410016 454 0 Tile_X9Y15_I_top13
rlabel metal3 410784 454 410784 454 0 Tile_X9Y15_I_top14
rlabel metal3 411552 454 411552 454 0 Tile_X9Y15_I_top15
rlabel metal3 401568 454 401568 454 0 Tile_X9Y15_I_top2
rlabel metal3 402336 454 402336 454 0 Tile_X9Y15_I_top3
rlabel metal3 403104 454 403104 454 0 Tile_X9Y15_I_top4
rlabel metal3 403872 454 403872 454 0 Tile_X9Y15_I_top5
rlabel metal3 404640 454 404640 454 0 Tile_X9Y15_I_top6
rlabel metal3 405408 454 405408 454 0 Tile_X9Y15_I_top7
rlabel metal3 406176 454 406176 454 0 Tile_X9Y15_I_top8
rlabel metal3 406944 454 406944 454 0 Tile_X9Y15_I_top9
rlabel metal3 387744 454 387744 454 0 Tile_X9Y15_O_top0
rlabel metal3 388512 454 388512 454 0 Tile_X9Y15_O_top1
rlabel metal3 395424 454 395424 454 0 Tile_X9Y15_O_top10
rlabel metal3 396192 454 396192 454 0 Tile_X9Y15_O_top11
rlabel metal3 396960 454 396960 454 0 Tile_X9Y15_O_top12
rlabel metal3 397728 454 397728 454 0 Tile_X9Y15_O_top13
rlabel metal3 398496 454 398496 454 0 Tile_X9Y15_O_top14
rlabel metal3 399264 454 399264 454 0 Tile_X9Y15_O_top15
rlabel metal3 389280 454 389280 454 0 Tile_X9Y15_O_top2
rlabel metal3 390048 454 390048 454 0 Tile_X9Y15_O_top3
rlabel metal3 390816 454 390816 454 0 Tile_X9Y15_O_top4
rlabel metal3 391584 454 391584 454 0 Tile_X9Y15_O_top5
rlabel metal3 392352 454 392352 454 0 Tile_X9Y15_O_top6
rlabel metal3 393120 454 393120 454 0 Tile_X9Y15_O_top7
rlabel metal3 393888 454 393888 454 0 Tile_X9Y15_O_top8
rlabel metal3 394656 454 394656 454 0 Tile_X9Y15_O_top9
rlabel metal3 280320 462 280320 462 0 UserCLK
<< properties >>
string FIXED_BBOX 0 0 452640 702336
<< end >>
