* NGSPICE file created from eFPGA.ext - technology: ihp-sg13g2

* Black-box entry subcircuit for N_IO abstract view
.subckt N_IO A_I_top A_O_top A_T_top A_config_C_bit0 A_config_C_bit1 A_config_C_bit2
+ A_config_C_bit3 B_I_top B_O_top B_T_top B_config_C_bit0 B_config_C_bit1 B_config_C_bit2
+ B_config_C_bit3 Ci FrameData[0] FrameData[10] FrameData[11] FrameData[12] FrameData[13]
+ FrameData[14] FrameData[15] FrameData[16] FrameData[17] FrameData[18] FrameData[19]
+ FrameData[1] FrameData[20] FrameData[21] FrameData[22] FrameData[23] FrameData[24]
+ FrameData[25] FrameData[26] FrameData[27] FrameData[28] FrameData[29] FrameData[2]
+ FrameData[30] FrameData[31] FrameData[3] FrameData[4] FrameData[5] FrameData[6]
+ FrameData[7] FrameData[8] FrameData[9] FrameData_O[0] FrameData_O[10] FrameData_O[11]
+ FrameData_O[12] FrameData_O[13] FrameData_O[14] FrameData_O[15] FrameData_O[16]
+ FrameData_O[17] FrameData_O[18] FrameData_O[19] FrameData_O[1] FrameData_O[20] FrameData_O[21]
+ FrameData_O[22] FrameData_O[23] FrameData_O[24] FrameData_O[25] FrameData_O[26]
+ FrameData_O[27] FrameData_O[28] FrameData_O[29] FrameData_O[2] FrameData_O[30] FrameData_O[31]
+ FrameData_O[3] FrameData_O[4] FrameData_O[5] FrameData_O[6] FrameData_O[7] FrameData_O[8]
+ FrameData_O[9] FrameStrobe[0] FrameStrobe[10] FrameStrobe[11] FrameStrobe[12] FrameStrobe[13]
+ FrameStrobe[14] FrameStrobe[15] FrameStrobe[16] FrameStrobe[17] FrameStrobe[18]
+ FrameStrobe[19] FrameStrobe[1] FrameStrobe[2] FrameStrobe[3] FrameStrobe[4] FrameStrobe[5]
+ FrameStrobe[6] FrameStrobe[7] FrameStrobe[8] FrameStrobe[9] FrameStrobe_O[0] FrameStrobe_O[10]
+ FrameStrobe_O[11] FrameStrobe_O[12] FrameStrobe_O[13] FrameStrobe_O[14] FrameStrobe_O[15]
+ FrameStrobe_O[16] FrameStrobe_O[17] FrameStrobe_O[18] FrameStrobe_O[19] FrameStrobe_O[1]
+ FrameStrobe_O[2] FrameStrobe_O[3] FrameStrobe_O[4] FrameStrobe_O[5] FrameStrobe_O[6]
+ FrameStrobe_O[7] FrameStrobe_O[8] FrameStrobe_O[9] N1END[0] N1END[1] N1END[2] N1END[3]
+ N2END[0] N2END[1] N2END[2] N2END[3] N2END[4] N2END[5] N2END[6] N2END[7] N2MID[0]
+ N2MID[1] N2MID[2] N2MID[3] N2MID[4] N2MID[5] N2MID[6] N2MID[7] N4END[0] N4END[10]
+ N4END[11] N4END[12] N4END[13] N4END[14] N4END[15] N4END[1] N4END[2] N4END[3] N4END[4]
+ N4END[5] N4END[6] N4END[7] N4END[8] N4END[9] NN4END[0] NN4END[10] NN4END[11] NN4END[12]
+ NN4END[13] NN4END[14] NN4END[15] NN4END[1] NN4END[2] NN4END[3] NN4END[4] NN4END[5]
+ NN4END[6] NN4END[7] NN4END[8] NN4END[9] S1BEG[0] S1BEG[1] S1BEG[2] S1BEG[3] S2BEG[0]
+ S2BEG[1] S2BEG[2] S2BEG[3] S2BEG[4] S2BEG[5] S2BEG[6] S2BEG[7] S2BEGb[0] S2BEGb[1]
+ S2BEGb[2] S2BEGb[3] S2BEGb[4] S2BEGb[5] S2BEGb[6] S2BEGb[7] S4BEG[0] S4BEG[10] S4BEG[11]
+ S4BEG[12] S4BEG[13] S4BEG[14] S4BEG[15] S4BEG[1] S4BEG[2] S4BEG[3] S4BEG[4] S4BEG[5]
+ S4BEG[6] S4BEG[7] S4BEG[8] S4BEG[9] SS4BEG[0] SS4BEG[10] SS4BEG[11] SS4BEG[12] SS4BEG[13]
+ SS4BEG[14] SS4BEG[15] SS4BEG[1] SS4BEG[2] SS4BEG[3] SS4BEG[4] SS4BEG[5] SS4BEG[6]
+ SS4BEG[7] SS4BEG[8] SS4BEG[9] UserCLK UserCLKo VGND VPWR
.ends

* Black-box entry subcircuit for LUT4AB abstract view
.subckt LUT4AB Ci Co E1BEG[0] E1BEG[1] E1BEG[2] E1BEG[3] E1END[0] E1END[1] E1END[2]
+ E1END[3] E2BEG[0] E2BEG[1] E2BEG[2] E2BEG[3] E2BEG[4] E2BEG[5] E2BEG[6] E2BEG[7]
+ E2BEGb[0] E2BEGb[1] E2BEGb[2] E2BEGb[3] E2BEGb[4] E2BEGb[5] E2BEGb[6] E2BEGb[7]
+ E2END[0] E2END[1] E2END[2] E2END[3] E2END[4] E2END[5] E2END[6] E2END[7] E2MID[0]
+ E2MID[1] E2MID[2] E2MID[3] E2MID[4] E2MID[5] E2MID[6] E2MID[7] E6BEG[0] E6BEG[10]
+ E6BEG[11] E6BEG[1] E6BEG[2] E6BEG[3] E6BEG[4] E6BEG[5] E6BEG[6] E6BEG[7] E6BEG[8]
+ E6BEG[9] E6END[0] E6END[10] E6END[11] E6END[1] E6END[2] E6END[3] E6END[4] E6END[5]
+ E6END[6] E6END[7] E6END[8] E6END[9] EE4BEG[0] EE4BEG[10] EE4BEG[11] EE4BEG[12] EE4BEG[13]
+ EE4BEG[14] EE4BEG[15] EE4BEG[1] EE4BEG[2] EE4BEG[3] EE4BEG[4] EE4BEG[5] EE4BEG[6]
+ EE4BEG[7] EE4BEG[8] EE4BEG[9] EE4END[0] EE4END[10] EE4END[11] EE4END[12] EE4END[13]
+ EE4END[14] EE4END[15] EE4END[1] EE4END[2] EE4END[3] EE4END[4] EE4END[5] EE4END[6]
+ EE4END[7] EE4END[8] EE4END[9] FrameData[0] FrameData[10] FrameData[11] FrameData[12]
+ FrameData[13] FrameData[14] FrameData[15] FrameData[16] FrameData[17] FrameData[18]
+ FrameData[19] FrameData[1] FrameData[20] FrameData[21] FrameData[22] FrameData[23]
+ FrameData[24] FrameData[25] FrameData[26] FrameData[27] FrameData[28] FrameData[29]
+ FrameData[2] FrameData[30] FrameData[31] FrameData[3] FrameData[4] FrameData[5]
+ FrameData[6] FrameData[7] FrameData[8] FrameData[9] FrameData_O[0] FrameData_O[10]
+ FrameData_O[11] FrameData_O[12] FrameData_O[13] FrameData_O[14] FrameData_O[15]
+ FrameData_O[16] FrameData_O[17] FrameData_O[18] FrameData_O[19] FrameData_O[1] FrameData_O[20]
+ FrameData_O[21] FrameData_O[22] FrameData_O[23] FrameData_O[24] FrameData_O[25]
+ FrameData_O[26] FrameData_O[27] FrameData_O[28] FrameData_O[29] FrameData_O[2] FrameData_O[30]
+ FrameData_O[31] FrameData_O[3] FrameData_O[4] FrameData_O[5] FrameData_O[6] FrameData_O[7]
+ FrameData_O[8] FrameData_O[9] FrameStrobe[0] FrameStrobe[10] FrameStrobe[11] FrameStrobe[12]
+ FrameStrobe[13] FrameStrobe[14] FrameStrobe[15] FrameStrobe[16] FrameStrobe[17]
+ FrameStrobe[18] FrameStrobe[19] FrameStrobe[1] FrameStrobe[2] FrameStrobe[3] FrameStrobe[4]
+ FrameStrobe[5] FrameStrobe[6] FrameStrobe[7] FrameStrobe[8] FrameStrobe[9] FrameStrobe_O[0]
+ FrameStrobe_O[10] FrameStrobe_O[11] FrameStrobe_O[12] FrameStrobe_O[13] FrameStrobe_O[14]
+ FrameStrobe_O[15] FrameStrobe_O[16] FrameStrobe_O[17] FrameStrobe_O[18] FrameStrobe_O[19]
+ FrameStrobe_O[1] FrameStrobe_O[2] FrameStrobe_O[3] FrameStrobe_O[4] FrameStrobe_O[5]
+ FrameStrobe_O[6] FrameStrobe_O[7] FrameStrobe_O[8] FrameStrobe_O[9] N1BEG[0] N1BEG[1]
+ N1BEG[2] N1BEG[3] N1END[0] N1END[1] N1END[2] N1END[3] N2BEG[0] N2BEG[1] N2BEG[2]
+ N2BEG[3] N2BEG[4] N2BEG[5] N2BEG[6] N2BEG[7] N2BEGb[0] N2BEGb[1] N2BEGb[2] N2BEGb[3]
+ N2BEGb[4] N2BEGb[5] N2BEGb[6] N2BEGb[7] N2END[0] N2END[1] N2END[2] N2END[3] N2END[4]
+ N2END[5] N2END[6] N2END[7] N2MID[0] N2MID[1] N2MID[2] N2MID[3] N2MID[4] N2MID[5]
+ N2MID[6] N2MID[7] N4BEG[0] N4BEG[10] N4BEG[11] N4BEG[12] N4BEG[13] N4BEG[14] N4BEG[15]
+ N4BEG[1] N4BEG[2] N4BEG[3] N4BEG[4] N4BEG[5] N4BEG[6] N4BEG[7] N4BEG[8] N4BEG[9]
+ N4END[0] N4END[10] N4END[11] N4END[12] N4END[13] N4END[14] N4END[15] N4END[1] N4END[2]
+ N4END[3] N4END[4] N4END[5] N4END[6] N4END[7] N4END[8] N4END[9] NN4BEG[0] NN4BEG[10]
+ NN4BEG[11] NN4BEG[12] NN4BEG[13] NN4BEG[14] NN4BEG[15] NN4BEG[1] NN4BEG[2] NN4BEG[3]
+ NN4BEG[4] NN4BEG[5] NN4BEG[6] NN4BEG[7] NN4BEG[8] NN4BEG[9] NN4END[0] NN4END[10]
+ NN4END[11] NN4END[12] NN4END[13] NN4END[14] NN4END[15] NN4END[1] NN4END[2] NN4END[3]
+ NN4END[4] NN4END[5] NN4END[6] NN4END[7] NN4END[8] NN4END[9] S1BEG[0] S1BEG[1] S1BEG[2]
+ S1BEG[3] S1END[0] S1END[1] S1END[2] S1END[3] S2BEG[0] S2BEG[1] S2BEG[2] S2BEG[3]
+ S2BEG[4] S2BEG[5] S2BEG[6] S2BEG[7] S2BEGb[0] S2BEGb[1] S2BEGb[2] S2BEGb[3] S2BEGb[4]
+ S2BEGb[5] S2BEGb[6] S2BEGb[7] S2END[0] S2END[1] S2END[2] S2END[3] S2END[4] S2END[5]
+ S2END[6] S2END[7] S2MID[0] S2MID[1] S2MID[2] S2MID[3] S2MID[4] S2MID[5] S2MID[6]
+ S2MID[7] S4BEG[0] S4BEG[10] S4BEG[11] S4BEG[12] S4BEG[13] S4BEG[14] S4BEG[15] S4BEG[1]
+ S4BEG[2] S4BEG[3] S4BEG[4] S4BEG[5] S4BEG[6] S4BEG[7] S4BEG[8] S4BEG[9] S4END[0]
+ S4END[10] S4END[11] S4END[12] S4END[13] S4END[14] S4END[15] S4END[1] S4END[2] S4END[3]
+ S4END[4] S4END[5] S4END[6] S4END[7] S4END[8] S4END[9] SS4BEG[0] SS4BEG[10] SS4BEG[11]
+ SS4BEG[12] SS4BEG[13] SS4BEG[14] SS4BEG[15] SS4BEG[1] SS4BEG[2] SS4BEG[3] SS4BEG[4]
+ SS4BEG[5] SS4BEG[6] SS4BEG[7] SS4BEG[8] SS4BEG[9] SS4END[0] SS4END[10] SS4END[11]
+ SS4END[12] SS4END[13] SS4END[14] SS4END[15] SS4END[1] SS4END[2] SS4END[3] SS4END[4]
+ SS4END[5] SS4END[6] SS4END[7] SS4END[8] SS4END[9] UserCLK UserCLKo VGND VPWR W1BEG[0]
+ W1BEG[1] W1BEG[2] W1BEG[3] W1END[0] W1END[1] W1END[2] W1END[3] W2BEG[0] W2BEG[1]
+ W2BEG[2] W2BEG[3] W2BEG[4] W2BEG[5] W2BEG[6] W2BEG[7] W2BEGb[0] W2BEGb[1] W2BEGb[2]
+ W2BEGb[3] W2BEGb[4] W2BEGb[5] W2BEGb[6] W2BEGb[7] W2END[0] W2END[1] W2END[2] W2END[3]
+ W2END[4] W2END[5] W2END[6] W2END[7] W2MID[0] W2MID[1] W2MID[2] W2MID[3] W2MID[4]
+ W2MID[5] W2MID[6] W2MID[7] W6BEG[0] W6BEG[10] W6BEG[11] W6BEG[1] W6BEG[2] W6BEG[3]
+ W6BEG[4] W6BEG[5] W6BEG[6] W6BEG[7] W6BEG[8] W6BEG[9] W6END[0] W6END[10] W6END[11]
+ W6END[1] W6END[2] W6END[3] W6END[4] W6END[5] W6END[6] W6END[7] W6END[8] W6END[9]
+ WW4BEG[0] WW4BEG[10] WW4BEG[11] WW4BEG[12] WW4BEG[13] WW4BEG[14] WW4BEG[15] WW4BEG[1]
+ WW4BEG[2] WW4BEG[3] WW4BEG[4] WW4BEG[5] WW4BEG[6] WW4BEG[7] WW4BEG[8] WW4BEG[9]
+ WW4END[0] WW4END[10] WW4END[11] WW4END[12] WW4END[13] WW4END[14] WW4END[15] WW4END[1]
+ WW4END[2] WW4END[3] WW4END[4] WW4END[5] WW4END[6] WW4END[7] WW4END[8] WW4END[9]
.ends

* Black-box entry subcircuit for RegFile abstract view
.subckt RegFile E1BEG[0] E1BEG[1] E1BEG[2] E1BEG[3] E1END[0] E1END[1] E1END[2] E1END[3]
+ E2BEG[0] E2BEG[1] E2BEG[2] E2BEG[3] E2BEG[4] E2BEG[5] E2BEG[6] E2BEG[7] E2BEGb[0]
+ E2BEGb[1] E2BEGb[2] E2BEGb[3] E2BEGb[4] E2BEGb[5] E2BEGb[6] E2BEGb[7] E2END[0] E2END[1]
+ E2END[2] E2END[3] E2END[4] E2END[5] E2END[6] E2END[7] E2MID[0] E2MID[1] E2MID[2]
+ E2MID[3] E2MID[4] E2MID[5] E2MID[6] E2MID[7] E6BEG[0] E6BEG[10] E6BEG[11] E6BEG[1]
+ E6BEG[2] E6BEG[3] E6BEG[4] E6BEG[5] E6BEG[6] E6BEG[7] E6BEG[8] E6BEG[9] E6END[0]
+ E6END[10] E6END[11] E6END[1] E6END[2] E6END[3] E6END[4] E6END[5] E6END[6] E6END[7]
+ E6END[8] E6END[9] EE4BEG[0] EE4BEG[10] EE4BEG[11] EE4BEG[12] EE4BEG[13] EE4BEG[14]
+ EE4BEG[15] EE4BEG[1] EE4BEG[2] EE4BEG[3] EE4BEG[4] EE4BEG[5] EE4BEG[6] EE4BEG[7]
+ EE4BEG[8] EE4BEG[9] EE4END[0] EE4END[10] EE4END[11] EE4END[12] EE4END[13] EE4END[14]
+ EE4END[15] EE4END[1] EE4END[2] EE4END[3] EE4END[4] EE4END[5] EE4END[6] EE4END[7]
+ EE4END[8] EE4END[9] FrameData[0] FrameData[10] FrameData[11] FrameData[12] FrameData[13]
+ FrameData[14] FrameData[15] FrameData[16] FrameData[17] FrameData[18] FrameData[19]
+ FrameData[1] FrameData[20] FrameData[21] FrameData[22] FrameData[23] FrameData[24]
+ FrameData[25] FrameData[26] FrameData[27] FrameData[28] FrameData[29] FrameData[2]
+ FrameData[30] FrameData[31] FrameData[3] FrameData[4] FrameData[5] FrameData[6]
+ FrameData[7] FrameData[8] FrameData[9] FrameData_O[0] FrameData_O[10] FrameData_O[11]
+ FrameData_O[12] FrameData_O[13] FrameData_O[14] FrameData_O[15] FrameData_O[16]
+ FrameData_O[17] FrameData_O[18] FrameData_O[19] FrameData_O[1] FrameData_O[20] FrameData_O[21]
+ FrameData_O[22] FrameData_O[23] FrameData_O[24] FrameData_O[25] FrameData_O[26]
+ FrameData_O[27] FrameData_O[28] FrameData_O[29] FrameData_O[2] FrameData_O[30] FrameData_O[31]
+ FrameData_O[3] FrameData_O[4] FrameData_O[5] FrameData_O[6] FrameData_O[7] FrameData_O[8]
+ FrameData_O[9] FrameStrobe[0] FrameStrobe[10] FrameStrobe[11] FrameStrobe[12] FrameStrobe[13]
+ FrameStrobe[14] FrameStrobe[15] FrameStrobe[16] FrameStrobe[17] FrameStrobe[18]
+ FrameStrobe[19] FrameStrobe[1] FrameStrobe[2] FrameStrobe[3] FrameStrobe[4] FrameStrobe[5]
+ FrameStrobe[6] FrameStrobe[7] FrameStrobe[8] FrameStrobe[9] FrameStrobe_O[0] FrameStrobe_O[10]
+ FrameStrobe_O[11] FrameStrobe_O[12] FrameStrobe_O[13] FrameStrobe_O[14] FrameStrobe_O[15]
+ FrameStrobe_O[16] FrameStrobe_O[17] FrameStrobe_O[18] FrameStrobe_O[19] FrameStrobe_O[1]
+ FrameStrobe_O[2] FrameStrobe_O[3] FrameStrobe_O[4] FrameStrobe_O[5] FrameStrobe_O[6]
+ FrameStrobe_O[7] FrameStrobe_O[8] FrameStrobe_O[9] N1BEG[0] N1BEG[1] N1BEG[2] N1BEG[3]
+ N1END[0] N1END[1] N1END[2] N1END[3] N2BEG[0] N2BEG[1] N2BEG[2] N2BEG[3] N2BEG[4]
+ N2BEG[5] N2BEG[6] N2BEG[7] N2BEGb[0] N2BEGb[1] N2BEGb[2] N2BEGb[3] N2BEGb[4] N2BEGb[5]
+ N2BEGb[6] N2BEGb[7] N2END[0] N2END[1] N2END[2] N2END[3] N2END[4] N2END[5] N2END[6]
+ N2END[7] N2MID[0] N2MID[1] N2MID[2] N2MID[3] N2MID[4] N2MID[5] N2MID[6] N2MID[7]
+ N4BEG[0] N4BEG[10] N4BEG[11] N4BEG[12] N4BEG[13] N4BEG[14] N4BEG[15] N4BEG[1] N4BEG[2]
+ N4BEG[3] N4BEG[4] N4BEG[5] N4BEG[6] N4BEG[7] N4BEG[8] N4BEG[9] N4END[0] N4END[10]
+ N4END[11] N4END[12] N4END[13] N4END[14] N4END[15] N4END[1] N4END[2] N4END[3] N4END[4]
+ N4END[5] N4END[6] N4END[7] N4END[8] N4END[9] NN4BEG[0] NN4BEG[10] NN4BEG[11] NN4BEG[12]
+ NN4BEG[13] NN4BEG[14] NN4BEG[15] NN4BEG[1] NN4BEG[2] NN4BEG[3] NN4BEG[4] NN4BEG[5]
+ NN4BEG[6] NN4BEG[7] NN4BEG[8] NN4BEG[9] NN4END[0] NN4END[10] NN4END[11] NN4END[12]
+ NN4END[13] NN4END[14] NN4END[15] NN4END[1] NN4END[2] NN4END[3] NN4END[4] NN4END[5]
+ NN4END[6] NN4END[7] NN4END[8] NN4END[9] S1BEG[0] S1BEG[1] S1BEG[2] S1BEG[3] S1END[0]
+ S1END[1] S1END[2] S1END[3] S2BEG[0] S2BEG[1] S2BEG[2] S2BEG[3] S2BEG[4] S2BEG[5]
+ S2BEG[6] S2BEG[7] S2BEGb[0] S2BEGb[1] S2BEGb[2] S2BEGb[3] S2BEGb[4] S2BEGb[5] S2BEGb[6]
+ S2BEGb[7] S2END[0] S2END[1] S2END[2] S2END[3] S2END[4] S2END[5] S2END[6] S2END[7]
+ S2MID[0] S2MID[1] S2MID[2] S2MID[3] S2MID[4] S2MID[5] S2MID[6] S2MID[7] S4BEG[0]
+ S4BEG[10] S4BEG[11] S4BEG[12] S4BEG[13] S4BEG[14] S4BEG[15] S4BEG[1] S4BEG[2] S4BEG[3]
+ S4BEG[4] S4BEG[5] S4BEG[6] S4BEG[7] S4BEG[8] S4BEG[9] S4END[0] S4END[10] S4END[11]
+ S4END[12] S4END[13] S4END[14] S4END[15] S4END[1] S4END[2] S4END[3] S4END[4] S4END[5]
+ S4END[6] S4END[7] S4END[8] S4END[9] SS4BEG[0] SS4BEG[10] SS4BEG[11] SS4BEG[12] SS4BEG[13]
+ SS4BEG[14] SS4BEG[15] SS4BEG[1] SS4BEG[2] SS4BEG[3] SS4BEG[4] SS4BEG[5] SS4BEG[6]
+ SS4BEG[7] SS4BEG[8] SS4BEG[9] SS4END[0] SS4END[10] SS4END[11] SS4END[12] SS4END[13]
+ SS4END[14] SS4END[15] SS4END[1] SS4END[2] SS4END[3] SS4END[4] SS4END[5] SS4END[6]
+ SS4END[7] SS4END[8] SS4END[9] UserCLK UserCLKo VGND VPWR W1BEG[0] W1BEG[1] W1BEG[2]
+ W1BEG[3] W1END[0] W1END[1] W1END[2] W1END[3] W2BEG[0] W2BEG[1] W2BEG[2] W2BEG[3]
+ W2BEG[4] W2BEG[5] W2BEG[6] W2BEG[7] W2BEGb[0] W2BEGb[1] W2BEGb[2] W2BEGb[3] W2BEGb[4]
+ W2BEGb[5] W2BEGb[6] W2BEGb[7] W2END[0] W2END[1] W2END[2] W2END[3] W2END[4] W2END[5]
+ W2END[6] W2END[7] W2MID[0] W2MID[1] W2MID[2] W2MID[3] W2MID[4] W2MID[5] W2MID[6]
+ W2MID[7] W6BEG[0] W6BEG[10] W6BEG[11] W6BEG[1] W6BEG[2] W6BEG[3] W6BEG[4] W6BEG[5]
+ W6BEG[6] W6BEG[7] W6BEG[8] W6BEG[9] W6END[0] W6END[10] W6END[11] W6END[1] W6END[2]
+ W6END[3] W6END[4] W6END[5] W6END[6] W6END[7] W6END[8] W6END[9] WW4BEG[0] WW4BEG[10]
+ WW4BEG[11] WW4BEG[12] WW4BEG[13] WW4BEG[14] WW4BEG[15] WW4BEG[1] WW4BEG[2] WW4BEG[3]
+ WW4BEG[4] WW4BEG[5] WW4BEG[6] WW4BEG[7] WW4BEG[8] WW4BEG[9] WW4END[0] WW4END[10]
+ WW4END[11] WW4END[12] WW4END[13] WW4END[14] WW4END[15] WW4END[1] WW4END[2] WW4END[3]
+ WW4END[4] WW4END[5] WW4END[6] WW4END[7] WW4END[8] WW4END[9]
.ends

* Black-box entry subcircuit for S_term_IHP_SRAM abstract view
.subckt S_term_IHP_SRAM FrameData[0] FrameData[10] FrameData[11] FrameData[12] FrameData[13]
+ FrameData[14] FrameData[15] FrameData[16] FrameData[17] FrameData[18] FrameData[19]
+ FrameData[1] FrameData[20] FrameData[21] FrameData[22] FrameData[23] FrameData[24]
+ FrameData[25] FrameData[26] FrameData[27] FrameData[28] FrameData[29] FrameData[2]
+ FrameData[30] FrameData[31] FrameData[3] FrameData[4] FrameData[5] FrameData[6]
+ FrameData[7] FrameData[8] FrameData[9] FrameData_O[0] FrameData_O[10] FrameData_O[11]
+ FrameData_O[12] FrameData_O[13] FrameData_O[14] FrameData_O[15] FrameData_O[16]
+ FrameData_O[17] FrameData_O[18] FrameData_O[19] FrameData_O[1] FrameData_O[20] FrameData_O[21]
+ FrameData_O[22] FrameData_O[23] FrameData_O[24] FrameData_O[25] FrameData_O[26]
+ FrameData_O[27] FrameData_O[28] FrameData_O[29] FrameData_O[2] FrameData_O[30] FrameData_O[31]
+ FrameData_O[3] FrameData_O[4] FrameData_O[5] FrameData_O[6] FrameData_O[7] FrameData_O[8]
+ FrameData_O[9] FrameStrobe[0] FrameStrobe[10] FrameStrobe[11] FrameStrobe[12] FrameStrobe[13]
+ FrameStrobe[14] FrameStrobe[15] FrameStrobe[16] FrameStrobe[17] FrameStrobe[18]
+ FrameStrobe[19] FrameStrobe[1] FrameStrobe[2] FrameStrobe[3] FrameStrobe[4] FrameStrobe[5]
+ FrameStrobe[6] FrameStrobe[7] FrameStrobe[8] FrameStrobe[9] FrameStrobe_O[0] FrameStrobe_O[10]
+ FrameStrobe_O[11] FrameStrobe_O[12] FrameStrobe_O[13] FrameStrobe_O[14] FrameStrobe_O[15]
+ FrameStrobe_O[16] FrameStrobe_O[17] FrameStrobe_O[18] FrameStrobe_O[19] FrameStrobe_O[1]
+ FrameStrobe_O[2] FrameStrobe_O[3] FrameStrobe_O[4] FrameStrobe_O[5] FrameStrobe_O[6]
+ FrameStrobe_O[7] FrameStrobe_O[8] FrameStrobe_O[9] N1BEG[0] N1BEG[1] N1BEG[2] N1BEG[3]
+ N2BEG[0] N2BEG[1] N2BEG[2] N2BEG[3] N2BEG[4] N2BEG[5] N2BEG[6] N2BEG[7] N2BEGb[0]
+ N2BEGb[1] N2BEGb[2] N2BEGb[3] N2BEGb[4] N2BEGb[5] N2BEGb[6] N2BEGb[7] N4BEG[0] N4BEG[10]
+ N4BEG[11] N4BEG[12] N4BEG[13] N4BEG[14] N4BEG[15] N4BEG[1] N4BEG[2] N4BEG[3] N4BEG[4]
+ N4BEG[5] N4BEG[6] N4BEG[7] N4BEG[8] N4BEG[9] S1END[0] S1END[1] S1END[2] S1END[3]
+ S2END[0] S2END[1] S2END[2] S2END[3] S2END[4] S2END[5] S2END[6] S2END[7] S2MID[0]
+ S2MID[1] S2MID[2] S2MID[3] S2MID[4] S2MID[5] S2MID[6] S2MID[7] S4END[0] S4END[10]
+ S4END[11] S4END[12] S4END[13] S4END[14] S4END[15] S4END[1] S4END[2] S4END[3] S4END[4]
+ S4END[5] S4END[6] S4END[7] S4END[8] S4END[9] UserCLK UserCLKo VGND VPWR
.ends

* Black-box entry subcircuit for W_IO abstract view
.subckt W_IO A_I_top A_O_top A_T_top A_config_C_bit0 A_config_C_bit1 A_config_C_bit2
+ A_config_C_bit3 B_I_top B_O_top B_T_top B_config_C_bit0 B_config_C_bit1 B_config_C_bit2
+ B_config_C_bit3 E1BEG[0] E1BEG[1] E1BEG[2] E1BEG[3] E2BEG[0] E2BEG[1] E2BEG[2] E2BEG[3]
+ E2BEG[4] E2BEG[5] E2BEG[6] E2BEG[7] E2BEGb[0] E2BEGb[1] E2BEGb[2] E2BEGb[3] E2BEGb[4]
+ E2BEGb[5] E2BEGb[6] E2BEGb[7] E6BEG[0] E6BEG[10] E6BEG[11] E6BEG[1] E6BEG[2] E6BEG[3]
+ E6BEG[4] E6BEG[5] E6BEG[6] E6BEG[7] E6BEG[8] E6BEG[9] EE4BEG[0] EE4BEG[10] EE4BEG[11]
+ EE4BEG[12] EE4BEG[13] EE4BEG[14] EE4BEG[15] EE4BEG[1] EE4BEG[2] EE4BEG[3] EE4BEG[4]
+ EE4BEG[5] EE4BEG[6] EE4BEG[7] EE4BEG[8] EE4BEG[9] FrameData[0] FrameData[10] FrameData[11]
+ FrameData[12] FrameData[13] FrameData[14] FrameData[15] FrameData[16] FrameData[17]
+ FrameData[18] FrameData[19] FrameData[1] FrameData[20] FrameData[21] FrameData[22]
+ FrameData[23] FrameData[24] FrameData[25] FrameData[26] FrameData[27] FrameData[28]
+ FrameData[29] FrameData[2] FrameData[30] FrameData[31] FrameData[3] FrameData[4]
+ FrameData[5] FrameData[6] FrameData[7] FrameData[8] FrameData[9] FrameData_O[0]
+ FrameData_O[10] FrameData_O[11] FrameData_O[12] FrameData_O[13] FrameData_O[14]
+ FrameData_O[15] FrameData_O[16] FrameData_O[17] FrameData_O[18] FrameData_O[19]
+ FrameData_O[1] FrameData_O[20] FrameData_O[21] FrameData_O[22] FrameData_O[23] FrameData_O[24]
+ FrameData_O[25] FrameData_O[26] FrameData_O[27] FrameData_O[28] FrameData_O[29]
+ FrameData_O[2] FrameData_O[30] FrameData_O[31] FrameData_O[3] FrameData_O[4] FrameData_O[5]
+ FrameData_O[6] FrameData_O[7] FrameData_O[8] FrameData_O[9] FrameStrobe[0] FrameStrobe[10]
+ FrameStrobe[11] FrameStrobe[12] FrameStrobe[13] FrameStrobe[14] FrameStrobe[15]
+ FrameStrobe[16] FrameStrobe[17] FrameStrobe[18] FrameStrobe[19] FrameStrobe[1] FrameStrobe[2]
+ FrameStrobe[3] FrameStrobe[4] FrameStrobe[5] FrameStrobe[6] FrameStrobe[7] FrameStrobe[8]
+ FrameStrobe[9] FrameStrobe_O[0] FrameStrobe_O[10] FrameStrobe_O[11] FrameStrobe_O[12]
+ FrameStrobe_O[13] FrameStrobe_O[14] FrameStrobe_O[15] FrameStrobe_O[16] FrameStrobe_O[17]
+ FrameStrobe_O[18] FrameStrobe_O[19] FrameStrobe_O[1] FrameStrobe_O[2] FrameStrobe_O[3]
+ FrameStrobe_O[4] FrameStrobe_O[5] FrameStrobe_O[6] FrameStrobe_O[7] FrameStrobe_O[8]
+ FrameStrobe_O[9] UserCLK UserCLKo VGND VPWR W1END[0] W1END[1] W1END[2] W1END[3]
+ W2END[0] W2END[1] W2END[2] W2END[3] W2END[4] W2END[5] W2END[6] W2END[7] W2MID[0]
+ W2MID[1] W2MID[2] W2MID[3] W2MID[4] W2MID[5] W2MID[6] W2MID[7] W6END[0] W6END[10]
+ W6END[11] W6END[1] W6END[2] W6END[3] W6END[4] W6END[5] W6END[6] W6END[7] W6END[8]
+ W6END[9] WW4END[0] WW4END[10] WW4END[11] WW4END[12] WW4END[13] WW4END[14] WW4END[15]
+ WW4END[1] WW4END[2] WW4END[3] WW4END[4] WW4END[5] WW4END[6] WW4END[7] WW4END[8]
+ WW4END[9]
.ends

* Black-box entry subcircuit for S_term_DSP abstract view
.subckt S_term_DSP FrameData[0] FrameData[10] FrameData[11] FrameData[12] FrameData[13]
+ FrameData[14] FrameData[15] FrameData[16] FrameData[17] FrameData[18] FrameData[19]
+ FrameData[1] FrameData[20] FrameData[21] FrameData[22] FrameData[23] FrameData[24]
+ FrameData[25] FrameData[26] FrameData[27] FrameData[28] FrameData[29] FrameData[2]
+ FrameData[30] FrameData[31] FrameData[3] FrameData[4] FrameData[5] FrameData[6]
+ FrameData[7] FrameData[8] FrameData[9] FrameData_O[0] FrameData_O[10] FrameData_O[11]
+ FrameData_O[12] FrameData_O[13] FrameData_O[14] FrameData_O[15] FrameData_O[16]
+ FrameData_O[17] FrameData_O[18] FrameData_O[19] FrameData_O[1] FrameData_O[20] FrameData_O[21]
+ FrameData_O[22] FrameData_O[23] FrameData_O[24] FrameData_O[25] FrameData_O[26]
+ FrameData_O[27] FrameData_O[28] FrameData_O[29] FrameData_O[2] FrameData_O[30] FrameData_O[31]
+ FrameData_O[3] FrameData_O[4] FrameData_O[5] FrameData_O[6] FrameData_O[7] FrameData_O[8]
+ FrameData_O[9] FrameStrobe[0] FrameStrobe[10] FrameStrobe[11] FrameStrobe[12] FrameStrobe[13]
+ FrameStrobe[14] FrameStrobe[15] FrameStrobe[16] FrameStrobe[17] FrameStrobe[18]
+ FrameStrobe[19] FrameStrobe[1] FrameStrobe[2] FrameStrobe[3] FrameStrobe[4] FrameStrobe[5]
+ FrameStrobe[6] FrameStrobe[7] FrameStrobe[8] FrameStrobe[9] FrameStrobe_O[0] FrameStrobe_O[10]
+ FrameStrobe_O[11] FrameStrobe_O[12] FrameStrobe_O[13] FrameStrobe_O[14] FrameStrobe_O[15]
+ FrameStrobe_O[16] FrameStrobe_O[17] FrameStrobe_O[18] FrameStrobe_O[19] FrameStrobe_O[1]
+ FrameStrobe_O[2] FrameStrobe_O[3] FrameStrobe_O[4] FrameStrobe_O[5] FrameStrobe_O[6]
+ FrameStrobe_O[7] FrameStrobe_O[8] FrameStrobe_O[9] N1BEG[0] N1BEG[1] N1BEG[2] N1BEG[3]
+ N2BEG[0] N2BEG[1] N2BEG[2] N2BEG[3] N2BEG[4] N2BEG[5] N2BEG[6] N2BEG[7] N2BEGb[0]
+ N2BEGb[1] N2BEGb[2] N2BEGb[3] N2BEGb[4] N2BEGb[5] N2BEGb[6] N2BEGb[7] N4BEG[0] N4BEG[10]
+ N4BEG[11] N4BEG[12] N4BEG[13] N4BEG[14] N4BEG[15] N4BEG[1] N4BEG[2] N4BEG[3] N4BEG[4]
+ N4BEG[5] N4BEG[6] N4BEG[7] N4BEG[8] N4BEG[9] NN4BEG[0] NN4BEG[10] NN4BEG[11] NN4BEG[12]
+ NN4BEG[13] NN4BEG[14] NN4BEG[15] NN4BEG[1] NN4BEG[2] NN4BEG[3] NN4BEG[4] NN4BEG[5]
+ NN4BEG[6] NN4BEG[7] NN4BEG[8] NN4BEG[9] S1END[0] S1END[1] S1END[2] S1END[3] S2END[0]
+ S2END[1] S2END[2] S2END[3] S2END[4] S2END[5] S2END[6] S2END[7] S2MID[0] S2MID[1]
+ S2MID[2] S2MID[3] S2MID[4] S2MID[5] S2MID[6] S2MID[7] S4END[0] S4END[10] S4END[11]
+ S4END[12] S4END[13] S4END[14] S4END[15] S4END[1] S4END[2] S4END[3] S4END[4] S4END[5]
+ S4END[6] S4END[7] S4END[8] S4END[9] SS4END[0] SS4END[10] SS4END[11] SS4END[12] SS4END[13]
+ SS4END[14] SS4END[15] SS4END[1] SS4END[2] SS4END[3] SS4END[4] SS4END[5] SS4END[6]
+ SS4END[7] SS4END[8] SS4END[9] UserCLK UserCLKo VGND VPWR
.ends

* Black-box entry subcircuit for DSP abstract view
.subckt DSP Tile_X0Y0_E1BEG[0] Tile_X0Y0_E1BEG[1] Tile_X0Y0_E1BEG[2] Tile_X0Y0_E1BEG[3]
+ Tile_X0Y0_E1END[0] Tile_X0Y0_E1END[1] Tile_X0Y0_E1END[2] Tile_X0Y0_E1END[3] Tile_X0Y0_E2BEG[0]
+ Tile_X0Y0_E2BEG[1] Tile_X0Y0_E2BEG[2] Tile_X0Y0_E2BEG[3] Tile_X0Y0_E2BEG[4] Tile_X0Y0_E2BEG[5]
+ Tile_X0Y0_E2BEG[6] Tile_X0Y0_E2BEG[7] Tile_X0Y0_E2BEGb[0] Tile_X0Y0_E2BEGb[1] Tile_X0Y0_E2BEGb[2]
+ Tile_X0Y0_E2BEGb[3] Tile_X0Y0_E2BEGb[4] Tile_X0Y0_E2BEGb[5] Tile_X0Y0_E2BEGb[6]
+ Tile_X0Y0_E2BEGb[7] Tile_X0Y0_E2END[0] Tile_X0Y0_E2END[1] Tile_X0Y0_E2END[2] Tile_X0Y0_E2END[3]
+ Tile_X0Y0_E2END[4] Tile_X0Y0_E2END[5] Tile_X0Y0_E2END[6] Tile_X0Y0_E2END[7] Tile_X0Y0_E2MID[0]
+ Tile_X0Y0_E2MID[1] Tile_X0Y0_E2MID[2] Tile_X0Y0_E2MID[3] Tile_X0Y0_E2MID[4] Tile_X0Y0_E2MID[5]
+ Tile_X0Y0_E2MID[6] Tile_X0Y0_E2MID[7] Tile_X0Y0_E6BEG[0] Tile_X0Y0_E6BEG[10] Tile_X0Y0_E6BEG[11]
+ Tile_X0Y0_E6BEG[1] Tile_X0Y0_E6BEG[2] Tile_X0Y0_E6BEG[3] Tile_X0Y0_E6BEG[4] Tile_X0Y0_E6BEG[5]
+ Tile_X0Y0_E6BEG[6] Tile_X0Y0_E6BEG[7] Tile_X0Y0_E6BEG[8] Tile_X0Y0_E6BEG[9] Tile_X0Y0_E6END[0]
+ Tile_X0Y0_E6END[10] Tile_X0Y0_E6END[11] Tile_X0Y0_E6END[1] Tile_X0Y0_E6END[2] Tile_X0Y0_E6END[3]
+ Tile_X0Y0_E6END[4] Tile_X0Y0_E6END[5] Tile_X0Y0_E6END[6] Tile_X0Y0_E6END[7] Tile_X0Y0_E6END[8]
+ Tile_X0Y0_E6END[9] Tile_X0Y0_EE4BEG[0] Tile_X0Y0_EE4BEG[10] Tile_X0Y0_EE4BEG[11]
+ Tile_X0Y0_EE4BEG[12] Tile_X0Y0_EE4BEG[13] Tile_X0Y0_EE4BEG[14] Tile_X0Y0_EE4BEG[15]
+ Tile_X0Y0_EE4BEG[1] Tile_X0Y0_EE4BEG[2] Tile_X0Y0_EE4BEG[3] Tile_X0Y0_EE4BEG[4]
+ Tile_X0Y0_EE4BEG[5] Tile_X0Y0_EE4BEG[6] Tile_X0Y0_EE4BEG[7] Tile_X0Y0_EE4BEG[8]
+ Tile_X0Y0_EE4BEG[9] Tile_X0Y0_EE4END[0] Tile_X0Y0_EE4END[10] Tile_X0Y0_EE4END[11]
+ Tile_X0Y0_EE4END[12] Tile_X0Y0_EE4END[13] Tile_X0Y0_EE4END[14] Tile_X0Y0_EE4END[15]
+ Tile_X0Y0_EE4END[1] Tile_X0Y0_EE4END[2] Tile_X0Y0_EE4END[3] Tile_X0Y0_EE4END[4]
+ Tile_X0Y0_EE4END[5] Tile_X0Y0_EE4END[6] Tile_X0Y0_EE4END[7] Tile_X0Y0_EE4END[8]
+ Tile_X0Y0_EE4END[9] Tile_X0Y0_FrameData[0] Tile_X0Y0_FrameData[10] Tile_X0Y0_FrameData[11]
+ Tile_X0Y0_FrameData[12] Tile_X0Y0_FrameData[13] Tile_X0Y0_FrameData[14] Tile_X0Y0_FrameData[15]
+ Tile_X0Y0_FrameData[16] Tile_X0Y0_FrameData[17] Tile_X0Y0_FrameData[18] Tile_X0Y0_FrameData[19]
+ Tile_X0Y0_FrameData[1] Tile_X0Y0_FrameData[20] Tile_X0Y0_FrameData[21] Tile_X0Y0_FrameData[22]
+ Tile_X0Y0_FrameData[23] Tile_X0Y0_FrameData[24] Tile_X0Y0_FrameData[25] Tile_X0Y0_FrameData[26]
+ Tile_X0Y0_FrameData[27] Tile_X0Y0_FrameData[28] Tile_X0Y0_FrameData[29] Tile_X0Y0_FrameData[2]
+ Tile_X0Y0_FrameData[30] Tile_X0Y0_FrameData[31] Tile_X0Y0_FrameData[3] Tile_X0Y0_FrameData[4]
+ Tile_X0Y0_FrameData[5] Tile_X0Y0_FrameData[6] Tile_X0Y0_FrameData[7] Tile_X0Y0_FrameData[8]
+ Tile_X0Y0_FrameData[9] Tile_X0Y0_FrameData_O[0] Tile_X0Y0_FrameData_O[10] Tile_X0Y0_FrameData_O[11]
+ Tile_X0Y0_FrameData_O[12] Tile_X0Y0_FrameData_O[13] Tile_X0Y0_FrameData_O[14] Tile_X0Y0_FrameData_O[15]
+ Tile_X0Y0_FrameData_O[16] Tile_X0Y0_FrameData_O[17] Tile_X0Y0_FrameData_O[18] Tile_X0Y0_FrameData_O[19]
+ Tile_X0Y0_FrameData_O[1] Tile_X0Y0_FrameData_O[20] Tile_X0Y0_FrameData_O[21] Tile_X0Y0_FrameData_O[22]
+ Tile_X0Y0_FrameData_O[23] Tile_X0Y0_FrameData_O[24] Tile_X0Y0_FrameData_O[25] Tile_X0Y0_FrameData_O[26]
+ Tile_X0Y0_FrameData_O[27] Tile_X0Y0_FrameData_O[28] Tile_X0Y0_FrameData_O[29] Tile_X0Y0_FrameData_O[2]
+ Tile_X0Y0_FrameData_O[30] Tile_X0Y0_FrameData_O[31] Tile_X0Y0_FrameData_O[3] Tile_X0Y0_FrameData_O[4]
+ Tile_X0Y0_FrameData_O[5] Tile_X0Y0_FrameData_O[6] Tile_X0Y0_FrameData_O[7] Tile_X0Y0_FrameData_O[8]
+ Tile_X0Y0_FrameData_O[9] Tile_X0Y0_FrameStrobe_O[0] Tile_X0Y0_FrameStrobe_O[10]
+ Tile_X0Y0_FrameStrobe_O[11] Tile_X0Y0_FrameStrobe_O[12] Tile_X0Y0_FrameStrobe_O[13]
+ Tile_X0Y0_FrameStrobe_O[14] Tile_X0Y0_FrameStrobe_O[15] Tile_X0Y0_FrameStrobe_O[16]
+ Tile_X0Y0_FrameStrobe_O[17] Tile_X0Y0_FrameStrobe_O[18] Tile_X0Y0_FrameStrobe_O[19]
+ Tile_X0Y0_FrameStrobe_O[1] Tile_X0Y0_FrameStrobe_O[2] Tile_X0Y0_FrameStrobe_O[3]
+ Tile_X0Y0_FrameStrobe_O[4] Tile_X0Y0_FrameStrobe_O[5] Tile_X0Y0_FrameStrobe_O[6]
+ Tile_X0Y0_FrameStrobe_O[7] Tile_X0Y0_FrameStrobe_O[8] Tile_X0Y0_FrameStrobe_O[9]
+ Tile_X0Y0_N1BEG[0] Tile_X0Y0_N1BEG[1] Tile_X0Y0_N1BEG[2] Tile_X0Y0_N1BEG[3] Tile_X0Y0_N2BEG[0]
+ Tile_X0Y0_N2BEG[1] Tile_X0Y0_N2BEG[2] Tile_X0Y0_N2BEG[3] Tile_X0Y0_N2BEG[4] Tile_X0Y0_N2BEG[5]
+ Tile_X0Y0_N2BEG[6] Tile_X0Y0_N2BEG[7] Tile_X0Y0_N2BEGb[0] Tile_X0Y0_N2BEGb[1] Tile_X0Y0_N2BEGb[2]
+ Tile_X0Y0_N2BEGb[3] Tile_X0Y0_N2BEGb[4] Tile_X0Y0_N2BEGb[5] Tile_X0Y0_N2BEGb[6]
+ Tile_X0Y0_N2BEGb[7] Tile_X0Y0_N4BEG[0] Tile_X0Y0_N4BEG[10] Tile_X0Y0_N4BEG[11] Tile_X0Y0_N4BEG[12]
+ Tile_X0Y0_N4BEG[13] Tile_X0Y0_N4BEG[14] Tile_X0Y0_N4BEG[15] Tile_X0Y0_N4BEG[1] Tile_X0Y0_N4BEG[2]
+ Tile_X0Y0_N4BEG[3] Tile_X0Y0_N4BEG[4] Tile_X0Y0_N4BEG[5] Tile_X0Y0_N4BEG[6] Tile_X0Y0_N4BEG[7]
+ Tile_X0Y0_N4BEG[8] Tile_X0Y0_N4BEG[9] Tile_X0Y0_NN4BEG[0] Tile_X0Y0_NN4BEG[10] Tile_X0Y0_NN4BEG[11]
+ Tile_X0Y0_NN4BEG[12] Tile_X0Y0_NN4BEG[13] Tile_X0Y0_NN4BEG[14] Tile_X0Y0_NN4BEG[15]
+ Tile_X0Y0_NN4BEG[1] Tile_X0Y0_NN4BEG[2] Tile_X0Y0_NN4BEG[3] Tile_X0Y0_NN4BEG[4]
+ Tile_X0Y0_NN4BEG[5] Tile_X0Y0_NN4BEG[6] Tile_X0Y0_NN4BEG[7] Tile_X0Y0_NN4BEG[8]
+ Tile_X0Y0_NN4BEG[9] Tile_X0Y0_S1END[0] Tile_X0Y0_S1END[1] Tile_X0Y0_S1END[2] Tile_X0Y0_S1END[3]
+ Tile_X0Y0_S2END[0] Tile_X0Y0_S2END[1] Tile_X0Y0_S2END[2] Tile_X0Y0_S2END[3] Tile_X0Y0_S2END[4]
+ Tile_X0Y0_S2END[5] Tile_X0Y0_S2END[6] Tile_X0Y0_S2END[7] Tile_X0Y0_S2MID[0] Tile_X0Y0_S2MID[1]
+ Tile_X0Y0_S2MID[2] Tile_X0Y0_S2MID[3] Tile_X0Y0_S2MID[4] Tile_X0Y0_S2MID[5] Tile_X0Y0_S2MID[6]
+ Tile_X0Y0_S2MID[7] Tile_X0Y0_S4END[0] Tile_X0Y0_S4END[10] Tile_X0Y0_S4END[11] Tile_X0Y0_S4END[12]
+ Tile_X0Y0_S4END[13] Tile_X0Y0_S4END[14] Tile_X0Y0_S4END[15] Tile_X0Y0_S4END[1] Tile_X0Y0_S4END[2]
+ Tile_X0Y0_S4END[3] Tile_X0Y0_S4END[4] Tile_X0Y0_S4END[5] Tile_X0Y0_S4END[6] Tile_X0Y0_S4END[7]
+ Tile_X0Y0_S4END[8] Tile_X0Y0_S4END[9] Tile_X0Y0_SS4END[0] Tile_X0Y0_SS4END[10] Tile_X0Y0_SS4END[11]
+ Tile_X0Y0_SS4END[12] Tile_X0Y0_SS4END[13] Tile_X0Y0_SS4END[14] Tile_X0Y0_SS4END[15]
+ Tile_X0Y0_SS4END[1] Tile_X0Y0_SS4END[2] Tile_X0Y0_SS4END[3] Tile_X0Y0_SS4END[4]
+ Tile_X0Y0_SS4END[5] Tile_X0Y0_SS4END[6] Tile_X0Y0_SS4END[7] Tile_X0Y0_SS4END[8]
+ Tile_X0Y0_SS4END[9] Tile_X0Y0_UserCLKo Tile_X0Y0_W1BEG[0] Tile_X0Y0_W1BEG[1] Tile_X0Y0_W1BEG[2]
+ Tile_X0Y0_W1BEG[3] Tile_X0Y0_W1END[0] Tile_X0Y0_W1END[1] Tile_X0Y0_W1END[2] Tile_X0Y0_W1END[3]
+ Tile_X0Y0_W2BEG[0] Tile_X0Y0_W2BEG[1] Tile_X0Y0_W2BEG[2] Tile_X0Y0_W2BEG[3] Tile_X0Y0_W2BEG[4]
+ Tile_X0Y0_W2BEG[5] Tile_X0Y0_W2BEG[6] Tile_X0Y0_W2BEG[7] Tile_X0Y0_W2BEGb[0] Tile_X0Y0_W2BEGb[1]
+ Tile_X0Y0_W2BEGb[2] Tile_X0Y0_W2BEGb[3] Tile_X0Y0_W2BEGb[4] Tile_X0Y0_W2BEGb[5]
+ Tile_X0Y0_W2BEGb[6] Tile_X0Y0_W2BEGb[7] Tile_X0Y0_W2END[0] Tile_X0Y0_W2END[1] Tile_X0Y0_W2END[2]
+ Tile_X0Y0_W2END[3] Tile_X0Y0_W2END[4] Tile_X0Y0_W2END[5] Tile_X0Y0_W2END[6] Tile_X0Y0_W2END[7]
+ Tile_X0Y0_W2MID[0] Tile_X0Y0_W2MID[1] Tile_X0Y0_W2MID[2] Tile_X0Y0_W2MID[3] Tile_X0Y0_W2MID[4]
+ Tile_X0Y0_W2MID[5] Tile_X0Y0_W2MID[6] Tile_X0Y0_W2MID[7] Tile_X0Y0_W6BEG[0] Tile_X0Y0_W6BEG[10]
+ Tile_X0Y0_W6BEG[11] Tile_X0Y0_W6BEG[1] Tile_X0Y0_W6BEG[2] Tile_X0Y0_W6BEG[3] Tile_X0Y0_W6BEG[4]
+ Tile_X0Y0_W6BEG[5] Tile_X0Y0_W6BEG[6] Tile_X0Y0_W6BEG[7] Tile_X0Y0_W6BEG[8] Tile_X0Y0_W6BEG[9]
+ Tile_X0Y0_W6END[0] Tile_X0Y0_W6END[10] Tile_X0Y0_W6END[11] Tile_X0Y0_W6END[1] Tile_X0Y0_W6END[2]
+ Tile_X0Y0_W6END[3] Tile_X0Y0_W6END[4] Tile_X0Y0_W6END[5] Tile_X0Y0_W6END[6] Tile_X0Y0_W6END[7]
+ Tile_X0Y0_W6END[8] Tile_X0Y0_W6END[9] Tile_X0Y0_WW4BEG[0] Tile_X0Y0_WW4BEG[10] Tile_X0Y0_WW4BEG[11]
+ Tile_X0Y0_WW4BEG[12] Tile_X0Y0_WW4BEG[13] Tile_X0Y0_WW4BEG[14] Tile_X0Y0_WW4BEG[15]
+ Tile_X0Y0_WW4BEG[1] Tile_X0Y0_WW4BEG[2] Tile_X0Y0_WW4BEG[3] Tile_X0Y0_WW4BEG[4]
+ Tile_X0Y0_WW4BEG[5] Tile_X0Y0_WW4BEG[6] Tile_X0Y0_WW4BEG[7] Tile_X0Y0_WW4BEG[8]
+ Tile_X0Y0_WW4BEG[9] Tile_X0Y0_WW4END[0] Tile_X0Y0_WW4END[10] Tile_X0Y0_WW4END[11]
+ Tile_X0Y0_WW4END[12] Tile_X0Y0_WW4END[13] Tile_X0Y0_WW4END[14] Tile_X0Y0_WW4END[15]
+ Tile_X0Y0_WW4END[1] Tile_X0Y0_WW4END[2] Tile_X0Y0_WW4END[3] Tile_X0Y0_WW4END[4]
+ Tile_X0Y0_WW4END[5] Tile_X0Y0_WW4END[6] Tile_X0Y0_WW4END[7] Tile_X0Y0_WW4END[8]
+ Tile_X0Y0_WW4END[9] Tile_X0Y1_E1BEG[0] Tile_X0Y1_E1BEG[1] Tile_X0Y1_E1BEG[2] Tile_X0Y1_E1BEG[3]
+ Tile_X0Y1_E1END[0] Tile_X0Y1_E1END[1] Tile_X0Y1_E1END[2] Tile_X0Y1_E1END[3] Tile_X0Y1_E2BEG[0]
+ Tile_X0Y1_E2BEG[1] Tile_X0Y1_E2BEG[2] Tile_X0Y1_E2BEG[3] Tile_X0Y1_E2BEG[4] Tile_X0Y1_E2BEG[5]
+ Tile_X0Y1_E2BEG[6] Tile_X0Y1_E2BEG[7] Tile_X0Y1_E2BEGb[0] Tile_X0Y1_E2BEGb[1] Tile_X0Y1_E2BEGb[2]
+ Tile_X0Y1_E2BEGb[3] Tile_X0Y1_E2BEGb[4] Tile_X0Y1_E2BEGb[5] Tile_X0Y1_E2BEGb[6]
+ Tile_X0Y1_E2BEGb[7] Tile_X0Y1_E2END[0] Tile_X0Y1_E2END[1] Tile_X0Y1_E2END[2] Tile_X0Y1_E2END[3]
+ Tile_X0Y1_E2END[4] Tile_X0Y1_E2END[5] Tile_X0Y1_E2END[6] Tile_X0Y1_E2END[7] Tile_X0Y1_E2MID[0]
+ Tile_X0Y1_E2MID[1] Tile_X0Y1_E2MID[2] Tile_X0Y1_E2MID[3] Tile_X0Y1_E2MID[4] Tile_X0Y1_E2MID[5]
+ Tile_X0Y1_E2MID[6] Tile_X0Y1_E2MID[7] Tile_X0Y1_E6BEG[0] Tile_X0Y1_E6BEG[10] Tile_X0Y1_E6BEG[11]
+ Tile_X0Y1_E6BEG[1] Tile_X0Y1_E6BEG[2] Tile_X0Y1_E6BEG[3] Tile_X0Y1_E6BEG[4] Tile_X0Y1_E6BEG[5]
+ Tile_X0Y1_E6BEG[6] Tile_X0Y1_E6BEG[7] Tile_X0Y1_E6BEG[8] Tile_X0Y1_E6BEG[9] Tile_X0Y1_E6END[0]
+ Tile_X0Y1_E6END[10] Tile_X0Y1_E6END[11] Tile_X0Y1_E6END[1] Tile_X0Y1_E6END[2] Tile_X0Y1_E6END[3]
+ Tile_X0Y1_E6END[4] Tile_X0Y1_E6END[5] Tile_X0Y1_E6END[6] Tile_X0Y1_E6END[7] Tile_X0Y1_E6END[8]
+ Tile_X0Y1_E6END[9] Tile_X0Y1_EE4BEG[0] Tile_X0Y1_EE4BEG[10] Tile_X0Y1_EE4BEG[11]
+ Tile_X0Y1_EE4BEG[12] Tile_X0Y1_EE4BEG[13] Tile_X0Y1_EE4BEG[14] Tile_X0Y1_EE4BEG[15]
+ Tile_X0Y1_EE4BEG[1] Tile_X0Y1_EE4BEG[2] Tile_X0Y1_EE4BEG[3] Tile_X0Y1_EE4BEG[4]
+ Tile_X0Y1_EE4BEG[5] Tile_X0Y1_EE4BEG[6] Tile_X0Y1_EE4BEG[7] Tile_X0Y1_EE4BEG[8]
+ Tile_X0Y1_EE4BEG[9] Tile_X0Y1_EE4END[0] Tile_X0Y1_EE4END[10] Tile_X0Y1_EE4END[11]
+ Tile_X0Y1_EE4END[12] Tile_X0Y1_EE4END[13] Tile_X0Y1_EE4END[14] Tile_X0Y1_EE4END[15]
+ Tile_X0Y1_EE4END[1] Tile_X0Y1_EE4END[2] Tile_X0Y1_EE4END[3] Tile_X0Y1_EE4END[4]
+ Tile_X0Y1_EE4END[5] Tile_X0Y1_EE4END[6] Tile_X0Y1_EE4END[7] Tile_X0Y1_EE4END[8]
+ Tile_X0Y1_EE4END[9] Tile_X0Y1_FrameData[0] Tile_X0Y1_FrameData[10] Tile_X0Y1_FrameData[11]
+ Tile_X0Y1_FrameData[12] Tile_X0Y1_FrameData[13] Tile_X0Y1_FrameData[14] Tile_X0Y1_FrameData[15]
+ Tile_X0Y1_FrameData[16] Tile_X0Y1_FrameData[17] Tile_X0Y1_FrameData[18] Tile_X0Y1_FrameData[19]
+ Tile_X0Y1_FrameData[1] Tile_X0Y1_FrameData[20] Tile_X0Y1_FrameData[21] Tile_X0Y1_FrameData[22]
+ Tile_X0Y1_FrameData[23] Tile_X0Y1_FrameData[24] Tile_X0Y1_FrameData[25] Tile_X0Y1_FrameData[26]
+ Tile_X0Y1_FrameData[27] Tile_X0Y1_FrameData[28] Tile_X0Y1_FrameData[29] Tile_X0Y1_FrameData[2]
+ Tile_X0Y1_FrameData[30] Tile_X0Y1_FrameData[31] Tile_X0Y1_FrameData[3] Tile_X0Y1_FrameData[4]
+ Tile_X0Y1_FrameData[5] Tile_X0Y1_FrameData[6] Tile_X0Y1_FrameData[7] Tile_X0Y1_FrameData[8]
+ Tile_X0Y1_FrameData[9] Tile_X0Y1_FrameData_O[0] Tile_X0Y1_FrameData_O[10] Tile_X0Y1_FrameData_O[11]
+ Tile_X0Y1_FrameData_O[12] Tile_X0Y1_FrameData_O[13] Tile_X0Y1_FrameData_O[14] Tile_X0Y1_FrameData_O[15]
+ Tile_X0Y1_FrameData_O[16] Tile_X0Y1_FrameData_O[17] Tile_X0Y1_FrameData_O[18] Tile_X0Y1_FrameData_O[19]
+ Tile_X0Y1_FrameData_O[1] Tile_X0Y1_FrameData_O[20] Tile_X0Y1_FrameData_O[21] Tile_X0Y1_FrameData_O[22]
+ Tile_X0Y1_FrameData_O[23] Tile_X0Y1_FrameData_O[24] Tile_X0Y1_FrameData_O[25] Tile_X0Y1_FrameData_O[26]
+ Tile_X0Y1_FrameData_O[27] Tile_X0Y1_FrameData_O[28] Tile_X0Y1_FrameData_O[29] Tile_X0Y1_FrameData_O[2]
+ Tile_X0Y1_FrameData_O[30] Tile_X0Y1_FrameData_O[31] Tile_X0Y1_FrameData_O[3] Tile_X0Y1_FrameData_O[4]
+ Tile_X0Y1_FrameData_O[5] Tile_X0Y1_FrameData_O[6] Tile_X0Y1_FrameData_O[7] Tile_X0Y1_FrameData_O[8]
+ Tile_X0Y1_FrameData_O[9] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_FrameStrobe[10] Tile_X0Y1_FrameStrobe[11]
+ Tile_X0Y1_FrameStrobe[12] Tile_X0Y1_FrameStrobe[13] Tile_X0Y1_FrameStrobe[14] Tile_X0Y1_FrameStrobe[15]
+ Tile_X0Y1_FrameStrobe[16] Tile_X0Y1_FrameStrobe[17] Tile_X0Y1_FrameStrobe[18] Tile_X0Y1_FrameStrobe[19]
+ Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_FrameStrobe[4]
+ Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_FrameStrobe[8]
+ Tile_X0Y1_FrameStrobe[9] Tile_X0Y1_N1END[0] Tile_X0Y1_N1END[1] Tile_X0Y1_N1END[2]
+ Tile_X0Y1_N1END[3] Tile_X0Y1_N2END[0] Tile_X0Y1_N2END[1] Tile_X0Y1_N2END[2] Tile_X0Y1_N2END[3]
+ Tile_X0Y1_N2END[4] Tile_X0Y1_N2END[5] Tile_X0Y1_N2END[6] Tile_X0Y1_N2END[7] Tile_X0Y1_N2MID[0]
+ Tile_X0Y1_N2MID[1] Tile_X0Y1_N2MID[2] Tile_X0Y1_N2MID[3] Tile_X0Y1_N2MID[4] Tile_X0Y1_N2MID[5]
+ Tile_X0Y1_N2MID[6] Tile_X0Y1_N2MID[7] Tile_X0Y1_N4END[0] Tile_X0Y1_N4END[10] Tile_X0Y1_N4END[11]
+ Tile_X0Y1_N4END[12] Tile_X0Y1_N4END[13] Tile_X0Y1_N4END[14] Tile_X0Y1_N4END[15]
+ Tile_X0Y1_N4END[1] Tile_X0Y1_N4END[2] Tile_X0Y1_N4END[3] Tile_X0Y1_N4END[4] Tile_X0Y1_N4END[5]
+ Tile_X0Y1_N4END[6] Tile_X0Y1_N4END[7] Tile_X0Y1_N4END[8] Tile_X0Y1_N4END[9] Tile_X0Y1_NN4END[0]
+ Tile_X0Y1_NN4END[10] Tile_X0Y1_NN4END[11] Tile_X0Y1_NN4END[12] Tile_X0Y1_NN4END[13]
+ Tile_X0Y1_NN4END[14] Tile_X0Y1_NN4END[15] Tile_X0Y1_NN4END[1] Tile_X0Y1_NN4END[2]
+ Tile_X0Y1_NN4END[3] Tile_X0Y1_NN4END[4] Tile_X0Y1_NN4END[5] Tile_X0Y1_NN4END[6]
+ Tile_X0Y1_NN4END[7] Tile_X0Y1_NN4END[8] Tile_X0Y1_NN4END[9] Tile_X0Y1_S1BEG[0] Tile_X0Y1_S1BEG[1]
+ Tile_X0Y1_S1BEG[2] Tile_X0Y1_S1BEG[3] Tile_X0Y1_S2BEG[0] Tile_X0Y1_S2BEG[1] Tile_X0Y1_S2BEG[2]
+ Tile_X0Y1_S2BEG[3] Tile_X0Y1_S2BEG[4] Tile_X0Y1_S2BEG[5] Tile_X0Y1_S2BEG[6] Tile_X0Y1_S2BEG[7]
+ Tile_X0Y1_S2BEGb[0] Tile_X0Y1_S2BEGb[1] Tile_X0Y1_S2BEGb[2] Tile_X0Y1_S2BEGb[3]
+ Tile_X0Y1_S2BEGb[4] Tile_X0Y1_S2BEGb[5] Tile_X0Y1_S2BEGb[6] Tile_X0Y1_S2BEGb[7]
+ Tile_X0Y1_S4BEG[0] Tile_X0Y1_S4BEG[10] Tile_X0Y1_S4BEG[11] Tile_X0Y1_S4BEG[12] Tile_X0Y1_S4BEG[13]
+ Tile_X0Y1_S4BEG[14] Tile_X0Y1_S4BEG[15] Tile_X0Y1_S4BEG[1] Tile_X0Y1_S4BEG[2] Tile_X0Y1_S4BEG[3]
+ Tile_X0Y1_S4BEG[4] Tile_X0Y1_S4BEG[5] Tile_X0Y1_S4BEG[6] Tile_X0Y1_S4BEG[7] Tile_X0Y1_S4BEG[8]
+ Tile_X0Y1_S4BEG[9] Tile_X0Y1_SS4BEG[0] Tile_X0Y1_SS4BEG[10] Tile_X0Y1_SS4BEG[11]
+ Tile_X0Y1_SS4BEG[12] Tile_X0Y1_SS4BEG[13] Tile_X0Y1_SS4BEG[14] Tile_X0Y1_SS4BEG[15]
+ Tile_X0Y1_SS4BEG[1] Tile_X0Y1_SS4BEG[2] Tile_X0Y1_SS4BEG[3] Tile_X0Y1_SS4BEG[4]
+ Tile_X0Y1_SS4BEG[5] Tile_X0Y1_SS4BEG[6] Tile_X0Y1_SS4BEG[7] Tile_X0Y1_SS4BEG[8]
+ Tile_X0Y1_SS4BEG[9] Tile_X0Y1_UserCLK Tile_X0Y1_W1BEG[0] Tile_X0Y1_W1BEG[1] Tile_X0Y1_W1BEG[2]
+ Tile_X0Y1_W1BEG[3] Tile_X0Y1_W1END[0] Tile_X0Y1_W1END[1] Tile_X0Y1_W1END[2] Tile_X0Y1_W1END[3]
+ Tile_X0Y1_W2BEG[0] Tile_X0Y1_W2BEG[1] Tile_X0Y1_W2BEG[2] Tile_X0Y1_W2BEG[3] Tile_X0Y1_W2BEG[4]
+ Tile_X0Y1_W2BEG[5] Tile_X0Y1_W2BEG[6] Tile_X0Y1_W2BEG[7] Tile_X0Y1_W2BEGb[0] Tile_X0Y1_W2BEGb[1]
+ Tile_X0Y1_W2BEGb[2] Tile_X0Y1_W2BEGb[3] Tile_X0Y1_W2BEGb[4] Tile_X0Y1_W2BEGb[5]
+ Tile_X0Y1_W2BEGb[6] Tile_X0Y1_W2BEGb[7] Tile_X0Y1_W2END[0] Tile_X0Y1_W2END[1] Tile_X0Y1_W2END[2]
+ Tile_X0Y1_W2END[3] Tile_X0Y1_W2END[4] Tile_X0Y1_W2END[5] Tile_X0Y1_W2END[6] Tile_X0Y1_W2END[7]
+ Tile_X0Y1_W2MID[0] Tile_X0Y1_W2MID[1] Tile_X0Y1_W2MID[2] Tile_X0Y1_W2MID[3] Tile_X0Y1_W2MID[4]
+ Tile_X0Y1_W2MID[5] Tile_X0Y1_W2MID[6] Tile_X0Y1_W2MID[7] Tile_X0Y1_W6BEG[0] Tile_X0Y1_W6BEG[10]
+ Tile_X0Y1_W6BEG[11] Tile_X0Y1_W6BEG[1] Tile_X0Y1_W6BEG[2] Tile_X0Y1_W6BEG[3] Tile_X0Y1_W6BEG[4]
+ Tile_X0Y1_W6BEG[5] Tile_X0Y1_W6BEG[6] Tile_X0Y1_W6BEG[7] Tile_X0Y1_W6BEG[8] Tile_X0Y1_W6BEG[9]
+ Tile_X0Y1_W6END[0] Tile_X0Y1_W6END[10] Tile_X0Y1_W6END[11] Tile_X0Y1_W6END[1] Tile_X0Y1_W6END[2]
+ Tile_X0Y1_W6END[3] Tile_X0Y1_W6END[4] Tile_X0Y1_W6END[5] Tile_X0Y1_W6END[6] Tile_X0Y1_W6END[7]
+ Tile_X0Y1_W6END[8] Tile_X0Y1_W6END[9] Tile_X0Y1_WW4BEG[0] Tile_X0Y1_WW4BEG[10] Tile_X0Y1_WW4BEG[11]
+ Tile_X0Y1_WW4BEG[12] Tile_X0Y1_WW4BEG[13] Tile_X0Y1_WW4BEG[14] Tile_X0Y1_WW4BEG[15]
+ Tile_X0Y1_WW4BEG[1] Tile_X0Y1_WW4BEG[2] Tile_X0Y1_WW4BEG[3] Tile_X0Y1_WW4BEG[4]
+ Tile_X0Y1_WW4BEG[5] Tile_X0Y1_WW4BEG[6] Tile_X0Y1_WW4BEG[7] Tile_X0Y1_WW4BEG[8]
+ Tile_X0Y1_WW4BEG[9] Tile_X0Y1_WW4END[0] Tile_X0Y1_WW4END[10] Tile_X0Y1_WW4END[11]
+ Tile_X0Y1_WW4END[12] Tile_X0Y1_WW4END[13] Tile_X0Y1_WW4END[14] Tile_X0Y1_WW4END[15]
+ Tile_X0Y1_WW4END[1] Tile_X0Y1_WW4END[2] Tile_X0Y1_WW4END[3] Tile_X0Y1_WW4END[4]
+ Tile_X0Y1_WW4END[5] Tile_X0Y1_WW4END[6] Tile_X0Y1_WW4END[7] Tile_X0Y1_WW4END[8]
+ Tile_X0Y1_WW4END[9] VGND VPWR
.ends

* Black-box entry subcircuit for S_WARMBOOT abstract view
.subckt S_WARMBOOT BOOT_top CONFIGURED_top Co FrameData[0] FrameData[10] FrameData[11]
+ FrameData[12] FrameData[13] FrameData[14] FrameData[15] FrameData[16] FrameData[17]
+ FrameData[18] FrameData[19] FrameData[1] FrameData[20] FrameData[21] FrameData[22]
+ FrameData[23] FrameData[24] FrameData[25] FrameData[26] FrameData[27] FrameData[28]
+ FrameData[29] FrameData[2] FrameData[30] FrameData[31] FrameData[3] FrameData[4]
+ FrameData[5] FrameData[6] FrameData[7] FrameData[8] FrameData[9] FrameData_O[0]
+ FrameData_O[10] FrameData_O[11] FrameData_O[12] FrameData_O[13] FrameData_O[14]
+ FrameData_O[15] FrameData_O[16] FrameData_O[17] FrameData_O[18] FrameData_O[19]
+ FrameData_O[1] FrameData_O[20] FrameData_O[21] FrameData_O[22] FrameData_O[23] FrameData_O[24]
+ FrameData_O[25] FrameData_O[26] FrameData_O[27] FrameData_O[28] FrameData_O[29]
+ FrameData_O[2] FrameData_O[30] FrameData_O[31] FrameData_O[3] FrameData_O[4] FrameData_O[5]
+ FrameData_O[6] FrameData_O[7] FrameData_O[8] FrameData_O[9] FrameStrobe[0] FrameStrobe[10]
+ FrameStrobe[11] FrameStrobe[12] FrameStrobe[13] FrameStrobe[14] FrameStrobe[15]
+ FrameStrobe[16] FrameStrobe[17] FrameStrobe[18] FrameStrobe[19] FrameStrobe[1] FrameStrobe[2]
+ FrameStrobe[3] FrameStrobe[4] FrameStrobe[5] FrameStrobe[6] FrameStrobe[7] FrameStrobe[8]
+ FrameStrobe[9] FrameStrobe_O[0] FrameStrobe_O[10] FrameStrobe_O[11] FrameStrobe_O[12]
+ FrameStrobe_O[13] FrameStrobe_O[14] FrameStrobe_O[15] FrameStrobe_O[16] FrameStrobe_O[17]
+ FrameStrobe_O[18] FrameStrobe_O[19] FrameStrobe_O[1] FrameStrobe_O[2] FrameStrobe_O[3]
+ FrameStrobe_O[4] FrameStrobe_O[5] FrameStrobe_O[6] FrameStrobe_O[7] FrameStrobe_O[8]
+ FrameStrobe_O[9] N1BEG[0] N1BEG[1] N1BEG[2] N1BEG[3] N2BEG[0] N2BEG[1] N2BEG[2]
+ N2BEG[3] N2BEG[4] N2BEG[5] N2BEG[6] N2BEG[7] N2BEGb[0] N2BEGb[1] N2BEGb[2] N2BEGb[3]
+ N2BEGb[4] N2BEGb[5] N2BEGb[6] N2BEGb[7] N4BEG[0] N4BEG[10] N4BEG[11] N4BEG[12] N4BEG[13]
+ N4BEG[14] N4BEG[15] N4BEG[1] N4BEG[2] N4BEG[3] N4BEG[4] N4BEG[5] N4BEG[6] N4BEG[7]
+ N4BEG[8] N4BEG[9] NN4BEG[0] NN4BEG[10] NN4BEG[11] NN4BEG[12] NN4BEG[13] NN4BEG[14]
+ NN4BEG[15] NN4BEG[1] NN4BEG[2] NN4BEG[3] NN4BEG[4] NN4BEG[5] NN4BEG[6] NN4BEG[7]
+ NN4BEG[8] NN4BEG[9] RESET_top S1END[0] S1END[1] S1END[2] S1END[3] S2END[0] S2END[1]
+ S2END[2] S2END[3] S2END[4] S2END[5] S2END[6] S2END[7] S2MID[0] S2MID[1] S2MID[2]
+ S2MID[3] S2MID[4] S2MID[5] S2MID[6] S2MID[7] S4END[0] S4END[10] S4END[11] S4END[12]
+ S4END[13] S4END[14] S4END[15] S4END[1] S4END[2] S4END[3] S4END[4] S4END[5] S4END[6]
+ S4END[7] S4END[8] S4END[9] SLOT_top0 SLOT_top1 SLOT_top2 SLOT_top3 SS4END[0] SS4END[10]
+ SS4END[11] SS4END[12] SS4END[13] SS4END[14] SS4END[15] SS4END[1] SS4END[2] SS4END[3]
+ SS4END[4] SS4END[5] SS4END[6] SS4END[7] SS4END[8] SS4END[9] UserCLK UserCLKo VGND
+ VPWR
.ends

* Black-box entry subcircuit for IHP_SRAM abstract view
.subckt IHP_SRAM ADDR_SRAM0 ADDR_SRAM1 ADDR_SRAM2 ADDR_SRAM3 ADDR_SRAM4 ADDR_SRAM5
+ ADDR_SRAM6 ADDR_SRAM7 ADDR_SRAM8 ADDR_SRAM9 BM_SRAM0 BM_SRAM1 BM_SRAM10 BM_SRAM11
+ BM_SRAM12 BM_SRAM13 BM_SRAM14 BM_SRAM15 BM_SRAM16 BM_SRAM17 BM_SRAM18 BM_SRAM19
+ BM_SRAM2 BM_SRAM20 BM_SRAM21 BM_SRAM22 BM_SRAM23 BM_SRAM24 BM_SRAM25 BM_SRAM26 BM_SRAM27
+ BM_SRAM28 BM_SRAM29 BM_SRAM3 BM_SRAM30 BM_SRAM31 BM_SRAM4 BM_SRAM5 BM_SRAM6 BM_SRAM7
+ BM_SRAM8 BM_SRAM9 CLK_SRAM CONFIGURED_top DIN_SRAM0 DIN_SRAM1 DIN_SRAM10 DIN_SRAM11
+ DIN_SRAM12 DIN_SRAM13 DIN_SRAM14 DIN_SRAM15 DIN_SRAM16 DIN_SRAM17 DIN_SRAM18 DIN_SRAM19
+ DIN_SRAM2 DIN_SRAM20 DIN_SRAM21 DIN_SRAM22 DIN_SRAM23 DIN_SRAM24 DIN_SRAM25 DIN_SRAM26
+ DIN_SRAM27 DIN_SRAM28 DIN_SRAM29 DIN_SRAM3 DIN_SRAM30 DIN_SRAM31 DIN_SRAM4 DIN_SRAM5
+ DIN_SRAM6 DIN_SRAM7 DIN_SRAM8 DIN_SRAM9 DOUT_SRAM0 DOUT_SRAM1 DOUT_SRAM10 DOUT_SRAM11
+ DOUT_SRAM12 DOUT_SRAM13 DOUT_SRAM14 DOUT_SRAM15 DOUT_SRAM16 DOUT_SRAM17 DOUT_SRAM18
+ DOUT_SRAM19 DOUT_SRAM2 DOUT_SRAM20 DOUT_SRAM21 DOUT_SRAM22 DOUT_SRAM23 DOUT_SRAM24
+ DOUT_SRAM25 DOUT_SRAM26 DOUT_SRAM27 DOUT_SRAM28 DOUT_SRAM29 DOUT_SRAM3 DOUT_SRAM30
+ DOUT_SRAM31 DOUT_SRAM4 DOUT_SRAM5 DOUT_SRAM6 DOUT_SRAM7 DOUT_SRAM8 DOUT_SRAM9 MEN_SRAM
+ REN_SRAM TIE_HIGH_SRAM TIE_LOW_SRAM Tile_X0Y0_E1END[0] Tile_X0Y0_E1END[1] Tile_X0Y0_E1END[2]
+ Tile_X0Y0_E1END[3] Tile_X0Y0_E2END[0] Tile_X0Y0_E2END[1] Tile_X0Y0_E2END[2] Tile_X0Y0_E2END[3]
+ Tile_X0Y0_E2END[4] Tile_X0Y0_E2END[5] Tile_X0Y0_E2END[6] Tile_X0Y0_E2END[7] Tile_X0Y0_E2MID[0]
+ Tile_X0Y0_E2MID[1] Tile_X0Y0_E2MID[2] Tile_X0Y0_E2MID[3] Tile_X0Y0_E2MID[4] Tile_X0Y0_E2MID[5]
+ Tile_X0Y0_E2MID[6] Tile_X0Y0_E2MID[7] Tile_X0Y0_E6END[0] Tile_X0Y0_E6END[10] Tile_X0Y0_E6END[11]
+ Tile_X0Y0_E6END[1] Tile_X0Y0_E6END[2] Tile_X0Y0_E6END[3] Tile_X0Y0_E6END[4] Tile_X0Y0_E6END[5]
+ Tile_X0Y0_E6END[6] Tile_X0Y0_E6END[7] Tile_X0Y0_E6END[8] Tile_X0Y0_E6END[9] Tile_X0Y0_EE4END[0]
+ Tile_X0Y0_EE4END[10] Tile_X0Y0_EE4END[11] Tile_X0Y0_EE4END[12] Tile_X0Y0_EE4END[13]
+ Tile_X0Y0_EE4END[14] Tile_X0Y0_EE4END[15] Tile_X0Y0_EE4END[1] Tile_X0Y0_EE4END[2]
+ Tile_X0Y0_EE4END[3] Tile_X0Y0_EE4END[4] Tile_X0Y0_EE4END[5] Tile_X0Y0_EE4END[6]
+ Tile_X0Y0_EE4END[7] Tile_X0Y0_EE4END[8] Tile_X0Y0_EE4END[9] Tile_X0Y0_FrameData[0]
+ Tile_X0Y0_FrameData[10] Tile_X0Y0_FrameData[11] Tile_X0Y0_FrameData[12] Tile_X0Y0_FrameData[13]
+ Tile_X0Y0_FrameData[14] Tile_X0Y0_FrameData[15] Tile_X0Y0_FrameData[16] Tile_X0Y0_FrameData[17]
+ Tile_X0Y0_FrameData[18] Tile_X0Y0_FrameData[19] Tile_X0Y0_FrameData[1] Tile_X0Y0_FrameData[20]
+ Tile_X0Y0_FrameData[21] Tile_X0Y0_FrameData[22] Tile_X0Y0_FrameData[23] Tile_X0Y0_FrameData[24]
+ Tile_X0Y0_FrameData[25] Tile_X0Y0_FrameData[26] Tile_X0Y0_FrameData[27] Tile_X0Y0_FrameData[28]
+ Tile_X0Y0_FrameData[29] Tile_X0Y0_FrameData[2] Tile_X0Y0_FrameData[30] Tile_X0Y0_FrameData[31]
+ Tile_X0Y0_FrameData[3] Tile_X0Y0_FrameData[4] Tile_X0Y0_FrameData[5] Tile_X0Y0_FrameData[6]
+ Tile_X0Y0_FrameData[7] Tile_X0Y0_FrameData[8] Tile_X0Y0_FrameData[9] Tile_X0Y0_FrameData_O[0]
+ Tile_X0Y0_FrameData_O[10] Tile_X0Y0_FrameData_O[11] Tile_X0Y0_FrameData_O[12] Tile_X0Y0_FrameData_O[13]
+ Tile_X0Y0_FrameData_O[14] Tile_X0Y0_FrameData_O[15] Tile_X0Y0_FrameData_O[16] Tile_X0Y0_FrameData_O[17]
+ Tile_X0Y0_FrameData_O[18] Tile_X0Y0_FrameData_O[19] Tile_X0Y0_FrameData_O[1] Tile_X0Y0_FrameData_O[20]
+ Tile_X0Y0_FrameData_O[21] Tile_X0Y0_FrameData_O[22] Tile_X0Y0_FrameData_O[23] Tile_X0Y0_FrameData_O[24]
+ Tile_X0Y0_FrameData_O[25] Tile_X0Y0_FrameData_O[26] Tile_X0Y0_FrameData_O[27] Tile_X0Y0_FrameData_O[28]
+ Tile_X0Y0_FrameData_O[29] Tile_X0Y0_FrameData_O[2] Tile_X0Y0_FrameData_O[30] Tile_X0Y0_FrameData_O[31]
+ Tile_X0Y0_FrameData_O[3] Tile_X0Y0_FrameData_O[4] Tile_X0Y0_FrameData_O[5] Tile_X0Y0_FrameData_O[6]
+ Tile_X0Y0_FrameData_O[7] Tile_X0Y0_FrameData_O[8] Tile_X0Y0_FrameData_O[9] Tile_X0Y0_FrameStrobe_O[0]
+ Tile_X0Y0_FrameStrobe_O[10] Tile_X0Y0_FrameStrobe_O[11] Tile_X0Y0_FrameStrobe_O[12]
+ Tile_X0Y0_FrameStrobe_O[13] Tile_X0Y0_FrameStrobe_O[14] Tile_X0Y0_FrameStrobe_O[15]
+ Tile_X0Y0_FrameStrobe_O[16] Tile_X0Y0_FrameStrobe_O[17] Tile_X0Y0_FrameStrobe_O[18]
+ Tile_X0Y0_FrameStrobe_O[19] Tile_X0Y0_FrameStrobe_O[1] Tile_X0Y0_FrameStrobe_O[2]
+ Tile_X0Y0_FrameStrobe_O[3] Tile_X0Y0_FrameStrobe_O[4] Tile_X0Y0_FrameStrobe_O[5]
+ Tile_X0Y0_FrameStrobe_O[6] Tile_X0Y0_FrameStrobe_O[7] Tile_X0Y0_FrameStrobe_O[8]
+ Tile_X0Y0_FrameStrobe_O[9] Tile_X0Y0_N1BEG[0] Tile_X0Y0_N1BEG[1] Tile_X0Y0_N1BEG[2]
+ Tile_X0Y0_N1BEG[3] Tile_X0Y0_N2BEG[0] Tile_X0Y0_N2BEG[1] Tile_X0Y0_N2BEG[2] Tile_X0Y0_N2BEG[3]
+ Tile_X0Y0_N2BEG[4] Tile_X0Y0_N2BEG[5] Tile_X0Y0_N2BEG[6] Tile_X0Y0_N2BEG[7] Tile_X0Y0_N2BEGb[0]
+ Tile_X0Y0_N2BEGb[1] Tile_X0Y0_N2BEGb[2] Tile_X0Y0_N2BEGb[3] Tile_X0Y0_N2BEGb[4]
+ Tile_X0Y0_N2BEGb[5] Tile_X0Y0_N2BEGb[6] Tile_X0Y0_N2BEGb[7] Tile_X0Y0_N4BEG[0] Tile_X0Y0_N4BEG[10]
+ Tile_X0Y0_N4BEG[11] Tile_X0Y0_N4BEG[12] Tile_X0Y0_N4BEG[13] Tile_X0Y0_N4BEG[14]
+ Tile_X0Y0_N4BEG[15] Tile_X0Y0_N4BEG[1] Tile_X0Y0_N4BEG[2] Tile_X0Y0_N4BEG[3] Tile_X0Y0_N4BEG[4]
+ Tile_X0Y0_N4BEG[5] Tile_X0Y0_N4BEG[6] Tile_X0Y0_N4BEG[7] Tile_X0Y0_N4BEG[8] Tile_X0Y0_N4BEG[9]
+ Tile_X0Y0_S1END[0] Tile_X0Y0_S1END[1] Tile_X0Y0_S1END[2] Tile_X0Y0_S1END[3] Tile_X0Y0_S2END[0]
+ Tile_X0Y0_S2END[1] Tile_X0Y0_S2END[2] Tile_X0Y0_S2END[3] Tile_X0Y0_S2END[4] Tile_X0Y0_S2END[5]
+ Tile_X0Y0_S2END[6] Tile_X0Y0_S2END[7] Tile_X0Y0_S2MID[0] Tile_X0Y0_S2MID[1] Tile_X0Y0_S2MID[2]
+ Tile_X0Y0_S2MID[3] Tile_X0Y0_S2MID[4] Tile_X0Y0_S2MID[5] Tile_X0Y0_S2MID[6] Tile_X0Y0_S2MID[7]
+ Tile_X0Y0_S4END[0] Tile_X0Y0_S4END[10] Tile_X0Y0_S4END[11] Tile_X0Y0_S4END[12] Tile_X0Y0_S4END[13]
+ Tile_X0Y0_S4END[14] Tile_X0Y0_S4END[15] Tile_X0Y0_S4END[1] Tile_X0Y0_S4END[2] Tile_X0Y0_S4END[3]
+ Tile_X0Y0_S4END[4] Tile_X0Y0_S4END[5] Tile_X0Y0_S4END[6] Tile_X0Y0_S4END[7] Tile_X0Y0_S4END[8]
+ Tile_X0Y0_S4END[9] Tile_X0Y0_UserCLKo Tile_X0Y0_W1BEG[0] Tile_X0Y0_W1BEG[1] Tile_X0Y0_W1BEG[2]
+ Tile_X0Y0_W1BEG[3] Tile_X0Y0_W2BEG[0] Tile_X0Y0_W2BEG[1] Tile_X0Y0_W2BEG[2] Tile_X0Y0_W2BEG[3]
+ Tile_X0Y0_W2BEG[4] Tile_X0Y0_W2BEG[5] Tile_X0Y0_W2BEG[6] Tile_X0Y0_W2BEG[7] Tile_X0Y0_W2BEGb[0]
+ Tile_X0Y0_W2BEGb[1] Tile_X0Y0_W2BEGb[2] Tile_X0Y0_W2BEGb[3] Tile_X0Y0_W2BEGb[4]
+ Tile_X0Y0_W2BEGb[5] Tile_X0Y0_W2BEGb[6] Tile_X0Y0_W2BEGb[7] Tile_X0Y0_W6BEG[0] Tile_X0Y0_W6BEG[10]
+ Tile_X0Y0_W6BEG[11] Tile_X0Y0_W6BEG[1] Tile_X0Y0_W6BEG[2] Tile_X0Y0_W6BEG[3] Tile_X0Y0_W6BEG[4]
+ Tile_X0Y0_W6BEG[5] Tile_X0Y0_W6BEG[6] Tile_X0Y0_W6BEG[7] Tile_X0Y0_W6BEG[8] Tile_X0Y0_W6BEG[9]
+ Tile_X0Y0_WW4BEG[0] Tile_X0Y0_WW4BEG[10] Tile_X0Y0_WW4BEG[11] Tile_X0Y0_WW4BEG[12]
+ Tile_X0Y0_WW4BEG[13] Tile_X0Y0_WW4BEG[14] Tile_X0Y0_WW4BEG[15] Tile_X0Y0_WW4BEG[1]
+ Tile_X0Y0_WW4BEG[2] Tile_X0Y0_WW4BEG[3] Tile_X0Y0_WW4BEG[4] Tile_X0Y0_WW4BEG[5]
+ Tile_X0Y0_WW4BEG[6] Tile_X0Y0_WW4BEG[7] Tile_X0Y0_WW4BEG[8] Tile_X0Y0_WW4BEG[9]
+ Tile_X0Y1_E1END[0] Tile_X0Y1_E1END[1] Tile_X0Y1_E1END[2] Tile_X0Y1_E1END[3] Tile_X0Y1_E2END[0]
+ Tile_X0Y1_E2END[1] Tile_X0Y1_E2END[2] Tile_X0Y1_E2END[3] Tile_X0Y1_E2END[4] Tile_X0Y1_E2END[5]
+ Tile_X0Y1_E2END[6] Tile_X0Y1_E2END[7] Tile_X0Y1_E2MID[0] Tile_X0Y1_E2MID[1] Tile_X0Y1_E2MID[2]
+ Tile_X0Y1_E2MID[3] Tile_X0Y1_E2MID[4] Tile_X0Y1_E2MID[5] Tile_X0Y1_E2MID[6] Tile_X0Y1_E2MID[7]
+ Tile_X0Y1_E6END[0] Tile_X0Y1_E6END[10] Tile_X0Y1_E6END[11] Tile_X0Y1_E6END[1] Tile_X0Y1_E6END[2]
+ Tile_X0Y1_E6END[3] Tile_X0Y1_E6END[4] Tile_X0Y1_E6END[5] Tile_X0Y1_E6END[6] Tile_X0Y1_E6END[7]
+ Tile_X0Y1_E6END[8] Tile_X0Y1_E6END[9] Tile_X0Y1_EE4END[0] Tile_X0Y1_EE4END[10] Tile_X0Y1_EE4END[11]
+ Tile_X0Y1_EE4END[12] Tile_X0Y1_EE4END[13] Tile_X0Y1_EE4END[14] Tile_X0Y1_EE4END[15]
+ Tile_X0Y1_EE4END[1] Tile_X0Y1_EE4END[2] Tile_X0Y1_EE4END[3] Tile_X0Y1_EE4END[4]
+ Tile_X0Y1_EE4END[5] Tile_X0Y1_EE4END[6] Tile_X0Y1_EE4END[7] Tile_X0Y1_EE4END[8]
+ Tile_X0Y1_EE4END[9] Tile_X0Y1_FrameData[0] Tile_X0Y1_FrameData[10] Tile_X0Y1_FrameData[11]
+ Tile_X0Y1_FrameData[12] Tile_X0Y1_FrameData[13] Tile_X0Y1_FrameData[14] Tile_X0Y1_FrameData[15]
+ Tile_X0Y1_FrameData[16] Tile_X0Y1_FrameData[17] Tile_X0Y1_FrameData[18] Tile_X0Y1_FrameData[19]
+ Tile_X0Y1_FrameData[1] Tile_X0Y1_FrameData[20] Tile_X0Y1_FrameData[21] Tile_X0Y1_FrameData[22]
+ Tile_X0Y1_FrameData[23] Tile_X0Y1_FrameData[24] Tile_X0Y1_FrameData[25] Tile_X0Y1_FrameData[26]
+ Tile_X0Y1_FrameData[27] Tile_X0Y1_FrameData[28] Tile_X0Y1_FrameData[29] Tile_X0Y1_FrameData[2]
+ Tile_X0Y1_FrameData[30] Tile_X0Y1_FrameData[31] Tile_X0Y1_FrameData[3] Tile_X0Y1_FrameData[4]
+ Tile_X0Y1_FrameData[5] Tile_X0Y1_FrameData[6] Tile_X0Y1_FrameData[7] Tile_X0Y1_FrameData[8]
+ Tile_X0Y1_FrameData[9] Tile_X0Y1_FrameData_O[0] Tile_X0Y1_FrameData_O[10] Tile_X0Y1_FrameData_O[11]
+ Tile_X0Y1_FrameData_O[12] Tile_X0Y1_FrameData_O[13] Tile_X0Y1_FrameData_O[14] Tile_X0Y1_FrameData_O[15]
+ Tile_X0Y1_FrameData_O[16] Tile_X0Y1_FrameData_O[17] Tile_X0Y1_FrameData_O[18] Tile_X0Y1_FrameData_O[19]
+ Tile_X0Y1_FrameData_O[1] Tile_X0Y1_FrameData_O[20] Tile_X0Y1_FrameData_O[21] Tile_X0Y1_FrameData_O[22]
+ Tile_X0Y1_FrameData_O[23] Tile_X0Y1_FrameData_O[24] Tile_X0Y1_FrameData_O[25] Tile_X0Y1_FrameData_O[26]
+ Tile_X0Y1_FrameData_O[27] Tile_X0Y1_FrameData_O[28] Tile_X0Y1_FrameData_O[29] Tile_X0Y1_FrameData_O[2]
+ Tile_X0Y1_FrameData_O[30] Tile_X0Y1_FrameData_O[31] Tile_X0Y1_FrameData_O[3] Tile_X0Y1_FrameData_O[4]
+ Tile_X0Y1_FrameData_O[5] Tile_X0Y1_FrameData_O[6] Tile_X0Y1_FrameData_O[7] Tile_X0Y1_FrameData_O[8]
+ Tile_X0Y1_FrameData_O[9] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_FrameStrobe[10] Tile_X0Y1_FrameStrobe[11]
+ Tile_X0Y1_FrameStrobe[12] Tile_X0Y1_FrameStrobe[13] Tile_X0Y1_FrameStrobe[14] Tile_X0Y1_FrameStrobe[15]
+ Tile_X0Y1_FrameStrobe[16] Tile_X0Y1_FrameStrobe[17] Tile_X0Y1_FrameStrobe[18] Tile_X0Y1_FrameStrobe[19]
+ Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_FrameStrobe[4]
+ Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_FrameStrobe[8]
+ Tile_X0Y1_FrameStrobe[9] Tile_X0Y1_N1END[0] Tile_X0Y1_N1END[1] Tile_X0Y1_N1END[2]
+ Tile_X0Y1_N1END[3] Tile_X0Y1_N2END[0] Tile_X0Y1_N2END[1] Tile_X0Y1_N2END[2] Tile_X0Y1_N2END[3]
+ Tile_X0Y1_N2END[4] Tile_X0Y1_N2END[5] Tile_X0Y1_N2END[6] Tile_X0Y1_N2END[7] Tile_X0Y1_N2MID[0]
+ Tile_X0Y1_N2MID[1] Tile_X0Y1_N2MID[2] Tile_X0Y1_N2MID[3] Tile_X0Y1_N2MID[4] Tile_X0Y1_N2MID[5]
+ Tile_X0Y1_N2MID[6] Tile_X0Y1_N2MID[7] Tile_X0Y1_N4END[0] Tile_X0Y1_N4END[10] Tile_X0Y1_N4END[11]
+ Tile_X0Y1_N4END[12] Tile_X0Y1_N4END[13] Tile_X0Y1_N4END[14] Tile_X0Y1_N4END[15]
+ Tile_X0Y1_N4END[1] Tile_X0Y1_N4END[2] Tile_X0Y1_N4END[3] Tile_X0Y1_N4END[4] Tile_X0Y1_N4END[5]
+ Tile_X0Y1_N4END[6] Tile_X0Y1_N4END[7] Tile_X0Y1_N4END[8] Tile_X0Y1_N4END[9] Tile_X0Y1_S1BEG[0]
+ Tile_X0Y1_S1BEG[1] Tile_X0Y1_S1BEG[2] Tile_X0Y1_S1BEG[3] Tile_X0Y1_S2BEG[0] Tile_X0Y1_S2BEG[1]
+ Tile_X0Y1_S2BEG[2] Tile_X0Y1_S2BEG[3] Tile_X0Y1_S2BEG[4] Tile_X0Y1_S2BEG[5] Tile_X0Y1_S2BEG[6]
+ Tile_X0Y1_S2BEG[7] Tile_X0Y1_S2BEGb[0] Tile_X0Y1_S2BEGb[1] Tile_X0Y1_S2BEGb[2] Tile_X0Y1_S2BEGb[3]
+ Tile_X0Y1_S2BEGb[4] Tile_X0Y1_S2BEGb[5] Tile_X0Y1_S2BEGb[6] Tile_X0Y1_S2BEGb[7]
+ Tile_X0Y1_S4BEG[0] Tile_X0Y1_S4BEG[10] Tile_X0Y1_S4BEG[11] Tile_X0Y1_S4BEG[12] Tile_X0Y1_S4BEG[13]
+ Tile_X0Y1_S4BEG[14] Tile_X0Y1_S4BEG[15] Tile_X0Y1_S4BEG[1] Tile_X0Y1_S4BEG[2] Tile_X0Y1_S4BEG[3]
+ Tile_X0Y1_S4BEG[4] Tile_X0Y1_S4BEG[5] Tile_X0Y1_S4BEG[6] Tile_X0Y1_S4BEG[7] Tile_X0Y1_S4BEG[8]
+ Tile_X0Y1_S4BEG[9] Tile_X0Y1_UserCLK Tile_X0Y1_W1BEG[0] Tile_X0Y1_W1BEG[1] Tile_X0Y1_W1BEG[2]
+ Tile_X0Y1_W1BEG[3] Tile_X0Y1_W2BEG[0] Tile_X0Y1_W2BEG[1] Tile_X0Y1_W2BEG[2] Tile_X0Y1_W2BEG[3]
+ Tile_X0Y1_W2BEG[4] Tile_X0Y1_W2BEG[5] Tile_X0Y1_W2BEG[6] Tile_X0Y1_W2BEG[7] Tile_X0Y1_W2BEGb[0]
+ Tile_X0Y1_W2BEGb[1] Tile_X0Y1_W2BEGb[2] Tile_X0Y1_W2BEGb[3] Tile_X0Y1_W2BEGb[4]
+ Tile_X0Y1_W2BEGb[5] Tile_X0Y1_W2BEGb[6] Tile_X0Y1_W2BEGb[7] Tile_X0Y1_W6BEG[0] Tile_X0Y1_W6BEG[10]
+ Tile_X0Y1_W6BEG[11] Tile_X0Y1_W6BEG[1] Tile_X0Y1_W6BEG[2] Tile_X0Y1_W6BEG[3] Tile_X0Y1_W6BEG[4]
+ Tile_X0Y1_W6BEG[5] Tile_X0Y1_W6BEG[6] Tile_X0Y1_W6BEG[7] Tile_X0Y1_W6BEG[8] Tile_X0Y1_W6BEG[9]
+ Tile_X0Y1_WW4BEG[0] Tile_X0Y1_WW4BEG[10] Tile_X0Y1_WW4BEG[11] Tile_X0Y1_WW4BEG[12]
+ Tile_X0Y1_WW4BEG[13] Tile_X0Y1_WW4BEG[14] Tile_X0Y1_WW4BEG[15] Tile_X0Y1_WW4BEG[1]
+ Tile_X0Y1_WW4BEG[2] Tile_X0Y1_WW4BEG[3] Tile_X0Y1_WW4BEG[4] Tile_X0Y1_WW4BEG[5]
+ Tile_X0Y1_WW4BEG[6] Tile_X0Y1_WW4BEG[7] Tile_X0Y1_WW4BEG[8] Tile_X0Y1_WW4BEG[9]
+ VGND VPWR WEN_SRAM
.ends

* Black-box entry subcircuit for N_term_single abstract view
.subckt N_term_single Ci FrameData[0] FrameData[10] FrameData[11] FrameData[12] FrameData[13]
+ FrameData[14] FrameData[15] FrameData[16] FrameData[17] FrameData[18] FrameData[19]
+ FrameData[1] FrameData[20] FrameData[21] FrameData[22] FrameData[23] FrameData[24]
+ FrameData[25] FrameData[26] FrameData[27] FrameData[28] FrameData[29] FrameData[2]
+ FrameData[30] FrameData[31] FrameData[3] FrameData[4] FrameData[5] FrameData[6]
+ FrameData[7] FrameData[8] FrameData[9] FrameData_O[0] FrameData_O[10] FrameData_O[11]
+ FrameData_O[12] FrameData_O[13] FrameData_O[14] FrameData_O[15] FrameData_O[16]
+ FrameData_O[17] FrameData_O[18] FrameData_O[19] FrameData_O[1] FrameData_O[20] FrameData_O[21]
+ FrameData_O[22] FrameData_O[23] FrameData_O[24] FrameData_O[25] FrameData_O[26]
+ FrameData_O[27] FrameData_O[28] FrameData_O[29] FrameData_O[2] FrameData_O[30] FrameData_O[31]
+ FrameData_O[3] FrameData_O[4] FrameData_O[5] FrameData_O[6] FrameData_O[7] FrameData_O[8]
+ FrameData_O[9] FrameStrobe[0] FrameStrobe[10] FrameStrobe[11] FrameStrobe[12] FrameStrobe[13]
+ FrameStrobe[14] FrameStrobe[15] FrameStrobe[16] FrameStrobe[17] FrameStrobe[18]
+ FrameStrobe[19] FrameStrobe[1] FrameStrobe[2] FrameStrobe[3] FrameStrobe[4] FrameStrobe[5]
+ FrameStrobe[6] FrameStrobe[7] FrameStrobe[8] FrameStrobe[9] FrameStrobe_O[0] FrameStrobe_O[10]
+ FrameStrobe_O[11] FrameStrobe_O[12] FrameStrobe_O[13] FrameStrobe_O[14] FrameStrobe_O[15]
+ FrameStrobe_O[16] FrameStrobe_O[17] FrameStrobe_O[18] FrameStrobe_O[19] FrameStrobe_O[1]
+ FrameStrobe_O[2] FrameStrobe_O[3] FrameStrobe_O[4] FrameStrobe_O[5] FrameStrobe_O[6]
+ FrameStrobe_O[7] FrameStrobe_O[8] FrameStrobe_O[9] N1END[0] N1END[1] N1END[2] N1END[3]
+ N2END[0] N2END[1] N2END[2] N2END[3] N2END[4] N2END[5] N2END[6] N2END[7] N2MID[0]
+ N2MID[1] N2MID[2] N2MID[3] N2MID[4] N2MID[5] N2MID[6] N2MID[7] N4END[0] N4END[10]
+ N4END[11] N4END[12] N4END[13] N4END[14] N4END[15] N4END[1] N4END[2] N4END[3] N4END[4]
+ N4END[5] N4END[6] N4END[7] N4END[8] N4END[9] NN4END[0] NN4END[10] NN4END[11] NN4END[12]
+ NN4END[13] NN4END[14] NN4END[15] NN4END[1] NN4END[2] NN4END[3] NN4END[4] NN4END[5]
+ NN4END[6] NN4END[7] NN4END[8] NN4END[9] S1BEG[0] S1BEG[1] S1BEG[2] S1BEG[3] S2BEG[0]
+ S2BEG[1] S2BEG[2] S2BEG[3] S2BEG[4] S2BEG[5] S2BEG[6] S2BEG[7] S2BEGb[0] S2BEGb[1]
+ S2BEGb[2] S2BEGb[3] S2BEGb[4] S2BEGb[5] S2BEGb[6] S2BEGb[7] S4BEG[0] S4BEG[10] S4BEG[11]
+ S4BEG[12] S4BEG[13] S4BEG[14] S4BEG[15] S4BEG[1] S4BEG[2] S4BEG[3] S4BEG[4] S4BEG[5]
+ S4BEG[6] S4BEG[7] S4BEG[8] S4BEG[9] SS4BEG[0] SS4BEG[10] SS4BEG[11] SS4BEG[12] SS4BEG[13]
+ SS4BEG[14] SS4BEG[15] SS4BEG[1] SS4BEG[2] SS4BEG[3] SS4BEG[4] SS4BEG[5] SS4BEG[6]
+ SS4BEG[7] SS4BEG[8] SS4BEG[9] UserCLK UserCLKo VGND VPWR
.ends

* Black-box entry subcircuit for S_term_single2 abstract view
.subckt S_term_single2 FrameData[0] FrameData[10] FrameData[11] FrameData[12] FrameData[13]
+ FrameData[14] FrameData[15] FrameData[16] FrameData[17] FrameData[18] FrameData[19]
+ FrameData[1] FrameData[20] FrameData[21] FrameData[22] FrameData[23] FrameData[24]
+ FrameData[25] FrameData[26] FrameData[27] FrameData[28] FrameData[29] FrameData[2]
+ FrameData[30] FrameData[31] FrameData[3] FrameData[4] FrameData[5] FrameData[6]
+ FrameData[7] FrameData[8] FrameData[9] FrameData_O[0] FrameData_O[10] FrameData_O[11]
+ FrameData_O[12] FrameData_O[13] FrameData_O[14] FrameData_O[15] FrameData_O[16]
+ FrameData_O[17] FrameData_O[18] FrameData_O[19] FrameData_O[1] FrameData_O[20] FrameData_O[21]
+ FrameData_O[22] FrameData_O[23] FrameData_O[24] FrameData_O[25] FrameData_O[26]
+ FrameData_O[27] FrameData_O[28] FrameData_O[29] FrameData_O[2] FrameData_O[30] FrameData_O[31]
+ FrameData_O[3] FrameData_O[4] FrameData_O[5] FrameData_O[6] FrameData_O[7] FrameData_O[8]
+ FrameData_O[9] FrameStrobe[0] FrameStrobe[10] FrameStrobe[11] FrameStrobe[12] FrameStrobe[13]
+ FrameStrobe[14] FrameStrobe[15] FrameStrobe[16] FrameStrobe[17] FrameStrobe[18]
+ FrameStrobe[19] FrameStrobe[1] FrameStrobe[2] FrameStrobe[3] FrameStrobe[4] FrameStrobe[5]
+ FrameStrobe[6] FrameStrobe[7] FrameStrobe[8] FrameStrobe[9] FrameStrobe_O[0] FrameStrobe_O[10]
+ FrameStrobe_O[11] FrameStrobe_O[12] FrameStrobe_O[13] FrameStrobe_O[14] FrameStrobe_O[15]
+ FrameStrobe_O[16] FrameStrobe_O[17] FrameStrobe_O[18] FrameStrobe_O[19] FrameStrobe_O[1]
+ FrameStrobe_O[2] FrameStrobe_O[3] FrameStrobe_O[4] FrameStrobe_O[5] FrameStrobe_O[6]
+ FrameStrobe_O[7] FrameStrobe_O[8] FrameStrobe_O[9] N1BEG[0] N1BEG[1] N1BEG[2] N1BEG[3]
+ N2BEG[0] N2BEG[1] N2BEG[2] N2BEG[3] N2BEG[4] N2BEG[5] N2BEG[6] N2BEG[7] N2BEGb[0]
+ N2BEGb[1] N2BEGb[2] N2BEGb[3] N2BEGb[4] N2BEGb[5] N2BEGb[6] N2BEGb[7] N4BEG[0] N4BEG[10]
+ N4BEG[11] N4BEG[12] N4BEG[13] N4BEG[14] N4BEG[15] N4BEG[1] N4BEG[2] N4BEG[3] N4BEG[4]
+ N4BEG[5] N4BEG[6] N4BEG[7] N4BEG[8] N4BEG[9] NN4BEG[0] NN4BEG[10] NN4BEG[11] NN4BEG[12]
+ NN4BEG[13] NN4BEG[14] NN4BEG[15] NN4BEG[1] NN4BEG[2] NN4BEG[3] NN4BEG[4] NN4BEG[5]
+ NN4BEG[6] NN4BEG[7] NN4BEG[8] NN4BEG[9] S1END[0] S1END[1] S1END[2] S1END[3] S2END[0]
+ S2END[1] S2END[2] S2END[3] S2END[4] S2END[5] S2END[6] S2END[7] S2MID[0] S2MID[1]
+ S2MID[2] S2MID[3] S2MID[4] S2MID[5] S2MID[6] S2MID[7] S4END[0] S4END[10] S4END[11]
+ S4END[12] S4END[13] S4END[14] S4END[15] S4END[1] S4END[2] S4END[3] S4END[4] S4END[5]
+ S4END[6] S4END[7] S4END[8] S4END[9] SS4END[0] SS4END[10] SS4END[11] SS4END[12] SS4END[13]
+ SS4END[14] SS4END[15] SS4END[1] SS4END[2] SS4END[3] SS4END[4] SS4END[5] SS4END[6]
+ SS4END[7] SS4END[8] SS4END[9] UserCLK UserCLKo VGND VPWR
.ends

* Black-box entry subcircuit for S_term_single abstract view
.subckt S_term_single Co FrameData[0] FrameData[10] FrameData[11] FrameData[12] FrameData[13]
+ FrameData[14] FrameData[15] FrameData[16] FrameData[17] FrameData[18] FrameData[19]
+ FrameData[1] FrameData[20] FrameData[21] FrameData[22] FrameData[23] FrameData[24]
+ FrameData[25] FrameData[26] FrameData[27] FrameData[28] FrameData[29] FrameData[2]
+ FrameData[30] FrameData[31] FrameData[3] FrameData[4] FrameData[5] FrameData[6]
+ FrameData[7] FrameData[8] FrameData[9] FrameData_O[0] FrameData_O[10] FrameData_O[11]
+ FrameData_O[12] FrameData_O[13] FrameData_O[14] FrameData_O[15] FrameData_O[16]
+ FrameData_O[17] FrameData_O[18] FrameData_O[19] FrameData_O[1] FrameData_O[20] FrameData_O[21]
+ FrameData_O[22] FrameData_O[23] FrameData_O[24] FrameData_O[25] FrameData_O[26]
+ FrameData_O[27] FrameData_O[28] FrameData_O[29] FrameData_O[2] FrameData_O[30] FrameData_O[31]
+ FrameData_O[3] FrameData_O[4] FrameData_O[5] FrameData_O[6] FrameData_O[7] FrameData_O[8]
+ FrameData_O[9] FrameStrobe[0] FrameStrobe[10] FrameStrobe[11] FrameStrobe[12] FrameStrobe[13]
+ FrameStrobe[14] FrameStrobe[15] FrameStrobe[16] FrameStrobe[17] FrameStrobe[18]
+ FrameStrobe[19] FrameStrobe[1] FrameStrobe[2] FrameStrobe[3] FrameStrobe[4] FrameStrobe[5]
+ FrameStrobe[6] FrameStrobe[7] FrameStrobe[8] FrameStrobe[9] FrameStrobe_O[0] FrameStrobe_O[10]
+ FrameStrobe_O[11] FrameStrobe_O[12] FrameStrobe_O[13] FrameStrobe_O[14] FrameStrobe_O[15]
+ FrameStrobe_O[16] FrameStrobe_O[17] FrameStrobe_O[18] FrameStrobe_O[19] FrameStrobe_O[1]
+ FrameStrobe_O[2] FrameStrobe_O[3] FrameStrobe_O[4] FrameStrobe_O[5] FrameStrobe_O[6]
+ FrameStrobe_O[7] FrameStrobe_O[8] FrameStrobe_O[9] N1BEG[0] N1BEG[1] N1BEG[2] N1BEG[3]
+ N2BEG[0] N2BEG[1] N2BEG[2] N2BEG[3] N2BEG[4] N2BEG[5] N2BEG[6] N2BEG[7] N2BEGb[0]
+ N2BEGb[1] N2BEGb[2] N2BEGb[3] N2BEGb[4] N2BEGb[5] N2BEGb[6] N2BEGb[7] N4BEG[0] N4BEG[10]
+ N4BEG[11] N4BEG[12] N4BEG[13] N4BEG[14] N4BEG[15] N4BEG[1] N4BEG[2] N4BEG[3] N4BEG[4]
+ N4BEG[5] N4BEG[6] N4BEG[7] N4BEG[8] N4BEG[9] NN4BEG[0] NN4BEG[10] NN4BEG[11] NN4BEG[12]
+ NN4BEG[13] NN4BEG[14] NN4BEG[15] NN4BEG[1] NN4BEG[2] NN4BEG[3] NN4BEG[4] NN4BEG[5]
+ NN4BEG[6] NN4BEG[7] NN4BEG[8] NN4BEG[9] S1END[0] S1END[1] S1END[2] S1END[3] S2END[0]
+ S2END[1] S2END[2] S2END[3] S2END[4] S2END[5] S2END[6] S2END[7] S2MID[0] S2MID[1]
+ S2MID[2] S2MID[3] S2MID[4] S2MID[5] S2MID[6] S2MID[7] S4END[0] S4END[10] S4END[11]
+ S4END[12] S4END[13] S4END[14] S4END[15] S4END[1] S4END[2] S4END[3] S4END[4] S4END[5]
+ S4END[6] S4END[7] S4END[8] S4END[9] SS4END[0] SS4END[10] SS4END[11] SS4END[12] SS4END[13]
+ SS4END[14] SS4END[15] SS4END[1] SS4END[2] SS4END[3] SS4END[4] SS4END[5] SS4END[6]
+ SS4END[7] SS4END[8] SS4END[9] UserCLK UserCLKo VGND VPWR
.ends

* Black-box entry subcircuit for S_CPU_IF abstract view
.subckt S_CPU_IF Co FrameData[0] FrameData[10] FrameData[11] FrameData[12] FrameData[13]
+ FrameData[14] FrameData[15] FrameData[16] FrameData[17] FrameData[18] FrameData[19]
+ FrameData[1] FrameData[20] FrameData[21] FrameData[22] FrameData[23] FrameData[24]
+ FrameData[25] FrameData[26] FrameData[27] FrameData[28] FrameData[29] FrameData[2]
+ FrameData[30] FrameData[31] FrameData[3] FrameData[4] FrameData[5] FrameData[6]
+ FrameData[7] FrameData[8] FrameData[9] FrameData_O[0] FrameData_O[10] FrameData_O[11]
+ FrameData_O[12] FrameData_O[13] FrameData_O[14] FrameData_O[15] FrameData_O[16]
+ FrameData_O[17] FrameData_O[18] FrameData_O[19] FrameData_O[1] FrameData_O[20] FrameData_O[21]
+ FrameData_O[22] FrameData_O[23] FrameData_O[24] FrameData_O[25] FrameData_O[26]
+ FrameData_O[27] FrameData_O[28] FrameData_O[29] FrameData_O[2] FrameData_O[30] FrameData_O[31]
+ FrameData_O[3] FrameData_O[4] FrameData_O[5] FrameData_O[6] FrameData_O[7] FrameData_O[8]
+ FrameData_O[9] FrameStrobe[0] FrameStrobe[10] FrameStrobe[11] FrameStrobe[12] FrameStrobe[13]
+ FrameStrobe[14] FrameStrobe[15] FrameStrobe[16] FrameStrobe[17] FrameStrobe[18]
+ FrameStrobe[19] FrameStrobe[1] FrameStrobe[2] FrameStrobe[3] FrameStrobe[4] FrameStrobe[5]
+ FrameStrobe[6] FrameStrobe[7] FrameStrobe[8] FrameStrobe[9] FrameStrobe_O[0] FrameStrobe_O[10]
+ FrameStrobe_O[11] FrameStrobe_O[12] FrameStrobe_O[13] FrameStrobe_O[14] FrameStrobe_O[15]
+ FrameStrobe_O[16] FrameStrobe_O[17] FrameStrobe_O[18] FrameStrobe_O[19] FrameStrobe_O[1]
+ FrameStrobe_O[2] FrameStrobe_O[3] FrameStrobe_O[4] FrameStrobe_O[5] FrameStrobe_O[6]
+ FrameStrobe_O[7] FrameStrobe_O[8] FrameStrobe_O[9] I_top0 I_top1 I_top10 I_top11
+ I_top12 I_top13 I_top14 I_top15 I_top2 I_top3 I_top4 I_top5 I_top6 I_top7 I_top8
+ I_top9 N1BEG[0] N1BEG[1] N1BEG[2] N1BEG[3] N2BEG[0] N2BEG[1] N2BEG[2] N2BEG[3] N2BEG[4]
+ N2BEG[5] N2BEG[6] N2BEG[7] N2BEGb[0] N2BEGb[1] N2BEGb[2] N2BEGb[3] N2BEGb[4] N2BEGb[5]
+ N2BEGb[6] N2BEGb[7] N4BEG[0] N4BEG[10] N4BEG[11] N4BEG[12] N4BEG[13] N4BEG[14] N4BEG[15]
+ N4BEG[1] N4BEG[2] N4BEG[3] N4BEG[4] N4BEG[5] N4BEG[6] N4BEG[7] N4BEG[8] N4BEG[9]
+ NN4BEG[0] NN4BEG[10] NN4BEG[11] NN4BEG[12] NN4BEG[13] NN4BEG[14] NN4BEG[15] NN4BEG[1]
+ NN4BEG[2] NN4BEG[3] NN4BEG[4] NN4BEG[5] NN4BEG[6] NN4BEG[7] NN4BEG[8] NN4BEG[9]
+ O_top0 O_top1 O_top10 O_top11 O_top12 O_top13 O_top14 O_top15 O_top2 O_top3 O_top4
+ O_top5 O_top6 O_top7 O_top8 O_top9 S1END[0] S1END[1] S1END[2] S1END[3] S2END[0]
+ S2END[1] S2END[2] S2END[3] S2END[4] S2END[5] S2END[6] S2END[7] S2MID[0] S2MID[1]
+ S2MID[2] S2MID[3] S2MID[4] S2MID[5] S2MID[6] S2MID[7] S4END[0] S4END[10] S4END[11]
+ S4END[12] S4END[13] S4END[14] S4END[15] S4END[1] S4END[2] S4END[3] S4END[4] S4END[5]
+ S4END[6] S4END[7] S4END[8] S4END[9] SS4END[0] SS4END[10] SS4END[11] SS4END[12] SS4END[13]
+ SS4END[14] SS4END[15] SS4END[1] SS4END[2] SS4END[3] SS4END[4] SS4END[5] SS4END[6]
+ SS4END[7] SS4END[8] SS4END[9] UserCLK UserCLKo VGND VPWR
.ends

* Black-box entry subcircuit for N_term_IHP_SRAM abstract view
.subckt N_term_IHP_SRAM FrameData[0] FrameData[10] FrameData[11] FrameData[12] FrameData[13]
+ FrameData[14] FrameData[15] FrameData[16] FrameData[17] FrameData[18] FrameData[19]
+ FrameData[1] FrameData[20] FrameData[21] FrameData[22] FrameData[23] FrameData[24]
+ FrameData[25] FrameData[26] FrameData[27] FrameData[28] FrameData[29] FrameData[2]
+ FrameData[30] FrameData[31] FrameData[3] FrameData[4] FrameData[5] FrameData[6]
+ FrameData[7] FrameData[8] FrameData[9] FrameData_O[0] FrameData_O[10] FrameData_O[11]
+ FrameData_O[12] FrameData_O[13] FrameData_O[14] FrameData_O[15] FrameData_O[16]
+ FrameData_O[17] FrameData_O[18] FrameData_O[19] FrameData_O[1] FrameData_O[20] FrameData_O[21]
+ FrameData_O[22] FrameData_O[23] FrameData_O[24] FrameData_O[25] FrameData_O[26]
+ FrameData_O[27] FrameData_O[28] FrameData_O[29] FrameData_O[2] FrameData_O[30] FrameData_O[31]
+ FrameData_O[3] FrameData_O[4] FrameData_O[5] FrameData_O[6] FrameData_O[7] FrameData_O[8]
+ FrameData_O[9] FrameStrobe[0] FrameStrobe[10] FrameStrobe[11] FrameStrobe[12] FrameStrobe[13]
+ FrameStrobe[14] FrameStrobe[15] FrameStrobe[16] FrameStrobe[17] FrameStrobe[18]
+ FrameStrobe[19] FrameStrobe[1] FrameStrobe[2] FrameStrobe[3] FrameStrobe[4] FrameStrobe[5]
+ FrameStrobe[6] FrameStrobe[7] FrameStrobe[8] FrameStrobe[9] FrameStrobe_O[0] FrameStrobe_O[10]
+ FrameStrobe_O[11] FrameStrobe_O[12] FrameStrobe_O[13] FrameStrobe_O[14] FrameStrobe_O[15]
+ FrameStrobe_O[16] FrameStrobe_O[17] FrameStrobe_O[18] FrameStrobe_O[19] FrameStrobe_O[1]
+ FrameStrobe_O[2] FrameStrobe_O[3] FrameStrobe_O[4] FrameStrobe_O[5] FrameStrobe_O[6]
+ FrameStrobe_O[7] FrameStrobe_O[8] FrameStrobe_O[9] N1END[0] N1END[1] N1END[2] N1END[3]
+ N2END[0] N2END[1] N2END[2] N2END[3] N2END[4] N2END[5] N2END[6] N2END[7] N2MID[0]
+ N2MID[1] N2MID[2] N2MID[3] N2MID[4] N2MID[5] N2MID[6] N2MID[7] N4END[0] N4END[10]
+ N4END[11] N4END[12] N4END[13] N4END[14] N4END[15] N4END[1] N4END[2] N4END[3] N4END[4]
+ N4END[5] N4END[6] N4END[7] N4END[8] N4END[9] S1BEG[0] S1BEG[1] S1BEG[2] S1BEG[3]
+ S2BEG[0] S2BEG[1] S2BEG[2] S2BEG[3] S2BEG[4] S2BEG[5] S2BEG[6] S2BEG[7] S2BEGb[0]
+ S2BEGb[1] S2BEGb[2] S2BEGb[3] S2BEGb[4] S2BEGb[5] S2BEGb[6] S2BEGb[7] S4BEG[0] S4BEG[10]
+ S4BEG[11] S4BEG[12] S4BEG[13] S4BEG[14] S4BEG[15] S4BEG[1] S4BEG[2] S4BEG[3] S4BEG[4]
+ S4BEG[5] S4BEG[6] S4BEG[7] S4BEG[8] S4BEG[9] UserCLK UserCLKo VGND VPWR
.ends

* Black-box entry subcircuit for S_CPU_IRQ abstract view
.subckt S_CPU_IRQ CONFIGURED_top Co FrameData[0] FrameData[10] FrameData[11] FrameData[12]
+ FrameData[13] FrameData[14] FrameData[15] FrameData[16] FrameData[17] FrameData[18]
+ FrameData[19] FrameData[1] FrameData[20] FrameData[21] FrameData[22] FrameData[23]
+ FrameData[24] FrameData[25] FrameData[26] FrameData[27] FrameData[28] FrameData[29]
+ FrameData[2] FrameData[30] FrameData[31] FrameData[3] FrameData[4] FrameData[5]
+ FrameData[6] FrameData[7] FrameData[8] FrameData[9] FrameData_O[0] FrameData_O[10]
+ FrameData_O[11] FrameData_O[12] FrameData_O[13] FrameData_O[14] FrameData_O[15]
+ FrameData_O[16] FrameData_O[17] FrameData_O[18] FrameData_O[19] FrameData_O[1] FrameData_O[20]
+ FrameData_O[21] FrameData_O[22] FrameData_O[23] FrameData_O[24] FrameData_O[25]
+ FrameData_O[26] FrameData_O[27] FrameData_O[28] FrameData_O[29] FrameData_O[2] FrameData_O[30]
+ FrameData_O[31] FrameData_O[3] FrameData_O[4] FrameData_O[5] FrameData_O[6] FrameData_O[7]
+ FrameData_O[8] FrameData_O[9] FrameStrobe[0] FrameStrobe[10] FrameStrobe[11] FrameStrobe[12]
+ FrameStrobe[13] FrameStrobe[14] FrameStrobe[15] FrameStrobe[16] FrameStrobe[17]
+ FrameStrobe[18] FrameStrobe[19] FrameStrobe[1] FrameStrobe[2] FrameStrobe[3] FrameStrobe[4]
+ FrameStrobe[5] FrameStrobe[6] FrameStrobe[7] FrameStrobe[8] FrameStrobe[9] FrameStrobe_O[0]
+ FrameStrobe_O[10] FrameStrobe_O[11] FrameStrobe_O[12] FrameStrobe_O[13] FrameStrobe_O[14]
+ FrameStrobe_O[15] FrameStrobe_O[16] FrameStrobe_O[17] FrameStrobe_O[18] FrameStrobe_O[19]
+ FrameStrobe_O[1] FrameStrobe_O[2] FrameStrobe_O[3] FrameStrobe_O[4] FrameStrobe_O[5]
+ FrameStrobe_O[6] FrameStrobe_O[7] FrameStrobe_O[8] FrameStrobe_O[9] IRQ_top0 IRQ_top1
+ IRQ_top2 IRQ_top3 N1BEG[0] N1BEG[1] N1BEG[2] N1BEG[3] N2BEG[0] N2BEG[1] N2BEG[2]
+ N2BEG[3] N2BEG[4] N2BEG[5] N2BEG[6] N2BEG[7] N2BEGb[0] N2BEGb[1] N2BEGb[2] N2BEGb[3]
+ N2BEGb[4] N2BEGb[5] N2BEGb[6] N2BEGb[7] N4BEG[0] N4BEG[10] N4BEG[11] N4BEG[12] N4BEG[13]
+ N4BEG[14] N4BEG[15] N4BEG[1] N4BEG[2] N4BEG[3] N4BEG[4] N4BEG[5] N4BEG[6] N4BEG[7]
+ N4BEG[8] N4BEG[9] NN4BEG[0] NN4BEG[10] NN4BEG[11] NN4BEG[12] NN4BEG[13] NN4BEG[14]
+ NN4BEG[15] NN4BEG[1] NN4BEG[2] NN4BEG[3] NN4BEG[4] NN4BEG[5] NN4BEG[6] NN4BEG[7]
+ NN4BEG[8] NN4BEG[9] S1END[0] S1END[1] S1END[2] S1END[3] S2END[0] S2END[1] S2END[2]
+ S2END[3] S2END[4] S2END[5] S2END[6] S2END[7] S2MID[0] S2MID[1] S2MID[2] S2MID[3]
+ S2MID[4] S2MID[5] S2MID[6] S2MID[7] S4END[0] S4END[10] S4END[11] S4END[12] S4END[13]
+ S4END[14] S4END[15] S4END[1] S4END[2] S4END[3] S4END[4] S4END[5] S4END[6] S4END[7]
+ S4END[8] S4END[9] SS4END[0] SS4END[10] SS4END[11] SS4END[12] SS4END[13] SS4END[14]
+ SS4END[15] SS4END[1] SS4END[2] SS4END[3] SS4END[4] SS4END[5] SS4END[6] SS4END[7]
+ SS4END[8] SS4END[9] UserCLK UserCLKo VGND VPWR
.ends

* Black-box entry subcircuit for N_term_DSP abstract view
.subckt N_term_DSP FrameData[0] FrameData[10] FrameData[11] FrameData[12] FrameData[13]
+ FrameData[14] FrameData[15] FrameData[16] FrameData[17] FrameData[18] FrameData[19]
+ FrameData[1] FrameData[20] FrameData[21] FrameData[22] FrameData[23] FrameData[24]
+ FrameData[25] FrameData[26] FrameData[27] FrameData[28] FrameData[29] FrameData[2]
+ FrameData[30] FrameData[31] FrameData[3] FrameData[4] FrameData[5] FrameData[6]
+ FrameData[7] FrameData[8] FrameData[9] FrameData_O[0] FrameData_O[10] FrameData_O[11]
+ FrameData_O[12] FrameData_O[13] FrameData_O[14] FrameData_O[15] FrameData_O[16]
+ FrameData_O[17] FrameData_O[18] FrameData_O[19] FrameData_O[1] FrameData_O[20] FrameData_O[21]
+ FrameData_O[22] FrameData_O[23] FrameData_O[24] FrameData_O[25] FrameData_O[26]
+ FrameData_O[27] FrameData_O[28] FrameData_O[29] FrameData_O[2] FrameData_O[30] FrameData_O[31]
+ FrameData_O[3] FrameData_O[4] FrameData_O[5] FrameData_O[6] FrameData_O[7] FrameData_O[8]
+ FrameData_O[9] FrameStrobe[0] FrameStrobe[10] FrameStrobe[11] FrameStrobe[12] FrameStrobe[13]
+ FrameStrobe[14] FrameStrobe[15] FrameStrobe[16] FrameStrobe[17] FrameStrobe[18]
+ FrameStrobe[19] FrameStrobe[1] FrameStrobe[2] FrameStrobe[3] FrameStrobe[4] FrameStrobe[5]
+ FrameStrobe[6] FrameStrobe[7] FrameStrobe[8] FrameStrobe[9] FrameStrobe_O[0] FrameStrobe_O[10]
+ FrameStrobe_O[11] FrameStrobe_O[12] FrameStrobe_O[13] FrameStrobe_O[14] FrameStrobe_O[15]
+ FrameStrobe_O[16] FrameStrobe_O[17] FrameStrobe_O[18] FrameStrobe_O[19] FrameStrobe_O[1]
+ FrameStrobe_O[2] FrameStrobe_O[3] FrameStrobe_O[4] FrameStrobe_O[5] FrameStrobe_O[6]
+ FrameStrobe_O[7] FrameStrobe_O[8] FrameStrobe_O[9] N1END[0] N1END[1] N1END[2] N1END[3]
+ N2END[0] N2END[1] N2END[2] N2END[3] N2END[4] N2END[5] N2END[6] N2END[7] N2MID[0]
+ N2MID[1] N2MID[2] N2MID[3] N2MID[4] N2MID[5] N2MID[6] N2MID[7] N4END[0] N4END[10]
+ N4END[11] N4END[12] N4END[13] N4END[14] N4END[15] N4END[1] N4END[2] N4END[3] N4END[4]
+ N4END[5] N4END[6] N4END[7] N4END[8] N4END[9] NN4END[0] NN4END[10] NN4END[11] NN4END[12]
+ NN4END[13] NN4END[14] NN4END[15] NN4END[1] NN4END[2] NN4END[3] NN4END[4] NN4END[5]
+ NN4END[6] NN4END[7] NN4END[8] NN4END[9] S1BEG[0] S1BEG[1] S1BEG[2] S1BEG[3] S2BEG[0]
+ S2BEG[1] S2BEG[2] S2BEG[3] S2BEG[4] S2BEG[5] S2BEG[6] S2BEG[7] S2BEGb[0] S2BEGb[1]
+ S2BEGb[2] S2BEGb[3] S2BEGb[4] S2BEGb[5] S2BEGb[6] S2BEGb[7] S4BEG[0] S4BEG[10] S4BEG[11]
+ S4BEG[12] S4BEG[13] S4BEG[14] S4BEG[15] S4BEG[1] S4BEG[2] S4BEG[3] S4BEG[4] S4BEG[5]
+ S4BEG[6] S4BEG[7] S4BEG[8] S4BEG[9] SS4BEG[0] SS4BEG[10] SS4BEG[11] SS4BEG[12] SS4BEG[13]
+ SS4BEG[14] SS4BEG[15] SS4BEG[1] SS4BEG[2] SS4BEG[3] SS4BEG[4] SS4BEG[5] SS4BEG[6]
+ SS4BEG[7] SS4BEG[8] SS4BEG[9] UserCLK UserCLKo VGND VPWR
.ends

* Black-box entry subcircuit for N_term_single2 abstract view
.subckt N_term_single2 FrameData[0] FrameData[10] FrameData[11] FrameData[12] FrameData[13]
+ FrameData[14] FrameData[15] FrameData[16] FrameData[17] FrameData[18] FrameData[19]
+ FrameData[1] FrameData[20] FrameData[21] FrameData[22] FrameData[23] FrameData[24]
+ FrameData[25] FrameData[26] FrameData[27] FrameData[28] FrameData[29] FrameData[2]
+ FrameData[30] FrameData[31] FrameData[3] FrameData[4] FrameData[5] FrameData[6]
+ FrameData[7] FrameData[8] FrameData[9] FrameData_O[0] FrameData_O[10] FrameData_O[11]
+ FrameData_O[12] FrameData_O[13] FrameData_O[14] FrameData_O[15] FrameData_O[16]
+ FrameData_O[17] FrameData_O[18] FrameData_O[19] FrameData_O[1] FrameData_O[20] FrameData_O[21]
+ FrameData_O[22] FrameData_O[23] FrameData_O[24] FrameData_O[25] FrameData_O[26]
+ FrameData_O[27] FrameData_O[28] FrameData_O[29] FrameData_O[2] FrameData_O[30] FrameData_O[31]
+ FrameData_O[3] FrameData_O[4] FrameData_O[5] FrameData_O[6] FrameData_O[7] FrameData_O[8]
+ FrameData_O[9] FrameStrobe[0] FrameStrobe[10] FrameStrobe[11] FrameStrobe[12] FrameStrobe[13]
+ FrameStrobe[14] FrameStrobe[15] FrameStrobe[16] FrameStrobe[17] FrameStrobe[18]
+ FrameStrobe[19] FrameStrobe[1] FrameStrobe[2] FrameStrobe[3] FrameStrobe[4] FrameStrobe[5]
+ FrameStrobe[6] FrameStrobe[7] FrameStrobe[8] FrameStrobe[9] FrameStrobe_O[0] FrameStrobe_O[10]
+ FrameStrobe_O[11] FrameStrobe_O[12] FrameStrobe_O[13] FrameStrobe_O[14] FrameStrobe_O[15]
+ FrameStrobe_O[16] FrameStrobe_O[17] FrameStrobe_O[18] FrameStrobe_O[19] FrameStrobe_O[1]
+ FrameStrobe_O[2] FrameStrobe_O[3] FrameStrobe_O[4] FrameStrobe_O[5] FrameStrobe_O[6]
+ FrameStrobe_O[7] FrameStrobe_O[8] FrameStrobe_O[9] N1END[0] N1END[1] N1END[2] N1END[3]
+ N2END[0] N2END[1] N2END[2] N2END[3] N2END[4] N2END[5] N2END[6] N2END[7] N2MID[0]
+ N2MID[1] N2MID[2] N2MID[3] N2MID[4] N2MID[5] N2MID[6] N2MID[7] N4END[0] N4END[10]
+ N4END[11] N4END[12] N4END[13] N4END[14] N4END[15] N4END[1] N4END[2] N4END[3] N4END[4]
+ N4END[5] N4END[6] N4END[7] N4END[8] N4END[9] NN4END[0] NN4END[10] NN4END[11] NN4END[12]
+ NN4END[13] NN4END[14] NN4END[15] NN4END[1] NN4END[2] NN4END[3] NN4END[4] NN4END[5]
+ NN4END[6] NN4END[7] NN4END[8] NN4END[9] S1BEG[0] S1BEG[1] S1BEG[2] S1BEG[3] S2BEG[0]
+ S2BEG[1] S2BEG[2] S2BEG[3] S2BEG[4] S2BEG[5] S2BEG[6] S2BEG[7] S2BEGb[0] S2BEGb[1]
+ S2BEGb[2] S2BEGb[3] S2BEGb[4] S2BEGb[5] S2BEGb[6] S2BEGb[7] S4BEG[0] S4BEG[10] S4BEG[11]
+ S4BEG[12] S4BEG[13] S4BEG[14] S4BEG[15] S4BEG[1] S4BEG[2] S4BEG[3] S4BEG[4] S4BEG[5]
+ S4BEG[6] S4BEG[7] S4BEG[8] S4BEG[9] SS4BEG[0] SS4BEG[10] SS4BEG[11] SS4BEG[12] SS4BEG[13]
+ SS4BEG[14] SS4BEG[15] SS4BEG[1] SS4BEG[2] SS4BEG[3] SS4BEG[4] SS4BEG[5] SS4BEG[6]
+ SS4BEG[7] SS4BEG[8] SS4BEG[9] UserCLK UserCLKo VGND VPWR
.ends

.subckt eFPGA FrameData[0] FrameData[100] FrameData[101] FrameData[102] FrameData[103]
+ FrameData[104] FrameData[105] FrameData[106] FrameData[107] FrameData[108] FrameData[109]
+ FrameData[10] FrameData[110] FrameData[111] FrameData[112] FrameData[113] FrameData[114]
+ FrameData[115] FrameData[116] FrameData[117] FrameData[118] FrameData[119] FrameData[11]
+ FrameData[120] FrameData[121] FrameData[122] FrameData[123] FrameData[124] FrameData[125]
+ FrameData[126] FrameData[127] FrameData[128] FrameData[129] FrameData[12] FrameData[130]
+ FrameData[131] FrameData[132] FrameData[133] FrameData[134] FrameData[135] FrameData[136]
+ FrameData[137] FrameData[138] FrameData[139] FrameData[13] FrameData[140] FrameData[141]
+ FrameData[142] FrameData[143] FrameData[144] FrameData[145] FrameData[146] FrameData[147]
+ FrameData[148] FrameData[149] FrameData[14] FrameData[150] FrameData[151] FrameData[152]
+ FrameData[153] FrameData[154] FrameData[155] FrameData[156] FrameData[157] FrameData[158]
+ FrameData[159] FrameData[15] FrameData[160] FrameData[161] FrameData[162] FrameData[163]
+ FrameData[164] FrameData[165] FrameData[166] FrameData[167] FrameData[168] FrameData[169]
+ FrameData[16] FrameData[170] FrameData[171] FrameData[172] FrameData[173] FrameData[174]
+ FrameData[175] FrameData[176] FrameData[177] FrameData[178] FrameData[179] FrameData[17]
+ FrameData[180] FrameData[181] FrameData[182] FrameData[183] FrameData[184] FrameData[185]
+ FrameData[186] FrameData[187] FrameData[188] FrameData[189] FrameData[18] FrameData[190]
+ FrameData[191] FrameData[192] FrameData[193] FrameData[194] FrameData[195] FrameData[196]
+ FrameData[197] FrameData[198] FrameData[199] FrameData[19] FrameData[1] FrameData[200]
+ FrameData[201] FrameData[202] FrameData[203] FrameData[204] FrameData[205] FrameData[206]
+ FrameData[207] FrameData[208] FrameData[209] FrameData[20] FrameData[210] FrameData[211]
+ FrameData[212] FrameData[213] FrameData[214] FrameData[215] FrameData[216] FrameData[217]
+ FrameData[218] FrameData[219] FrameData[21] FrameData[220] FrameData[221] FrameData[222]
+ FrameData[223] FrameData[224] FrameData[225] FrameData[226] FrameData[227] FrameData[228]
+ FrameData[229] FrameData[22] FrameData[230] FrameData[231] FrameData[232] FrameData[233]
+ FrameData[234] FrameData[235] FrameData[236] FrameData[237] FrameData[238] FrameData[239]
+ FrameData[23] FrameData[240] FrameData[241] FrameData[242] FrameData[243] FrameData[244]
+ FrameData[245] FrameData[246] FrameData[247] FrameData[248] FrameData[249] FrameData[24]
+ FrameData[250] FrameData[251] FrameData[252] FrameData[253] FrameData[254] FrameData[255]
+ FrameData[256] FrameData[257] FrameData[258] FrameData[259] FrameData[25] FrameData[260]
+ FrameData[261] FrameData[262] FrameData[263] FrameData[264] FrameData[265] FrameData[266]
+ FrameData[267] FrameData[268] FrameData[269] FrameData[26] FrameData[270] FrameData[271]
+ FrameData[272] FrameData[273] FrameData[274] FrameData[275] FrameData[276] FrameData[277]
+ FrameData[278] FrameData[279] FrameData[27] FrameData[280] FrameData[281] FrameData[282]
+ FrameData[283] FrameData[284] FrameData[285] FrameData[286] FrameData[287] FrameData[288]
+ FrameData[289] FrameData[28] FrameData[290] FrameData[291] FrameData[292] FrameData[293]
+ FrameData[294] FrameData[295] FrameData[296] FrameData[297] FrameData[298] FrameData[299]
+ FrameData[29] FrameData[2] FrameData[300] FrameData[301] FrameData[302] FrameData[303]
+ FrameData[304] FrameData[305] FrameData[306] FrameData[307] FrameData[308] FrameData[309]
+ FrameData[30] FrameData[310] FrameData[311] FrameData[312] FrameData[313] FrameData[314]
+ FrameData[315] FrameData[316] FrameData[317] FrameData[318] FrameData[319] FrameData[31]
+ FrameData[320] FrameData[321] FrameData[322] FrameData[323] FrameData[324] FrameData[325]
+ FrameData[326] FrameData[327] FrameData[328] FrameData[329] FrameData[32] FrameData[330]
+ FrameData[331] FrameData[332] FrameData[333] FrameData[334] FrameData[335] FrameData[336]
+ FrameData[337] FrameData[338] FrameData[339] FrameData[33] FrameData[340] FrameData[341]
+ FrameData[342] FrameData[343] FrameData[344] FrameData[345] FrameData[346] FrameData[347]
+ FrameData[348] FrameData[349] FrameData[34] FrameData[350] FrameData[351] FrameData[352]
+ FrameData[353] FrameData[354] FrameData[355] FrameData[356] FrameData[357] FrameData[358]
+ FrameData[359] FrameData[35] FrameData[360] FrameData[361] FrameData[362] FrameData[363]
+ FrameData[364] FrameData[365] FrameData[366] FrameData[367] FrameData[368] FrameData[369]
+ FrameData[36] FrameData[370] FrameData[371] FrameData[372] FrameData[373] FrameData[374]
+ FrameData[375] FrameData[376] FrameData[377] FrameData[378] FrameData[379] FrameData[37]
+ FrameData[380] FrameData[381] FrameData[382] FrameData[383] FrameData[384] FrameData[385]
+ FrameData[386] FrameData[387] FrameData[388] FrameData[389] FrameData[38] FrameData[390]
+ FrameData[391] FrameData[392] FrameData[393] FrameData[394] FrameData[395] FrameData[396]
+ FrameData[397] FrameData[398] FrameData[399] FrameData[39] FrameData[3] FrameData[400]
+ FrameData[401] FrameData[402] FrameData[403] FrameData[404] FrameData[405] FrameData[406]
+ FrameData[407] FrameData[408] FrameData[409] FrameData[40] FrameData[410] FrameData[411]
+ FrameData[412] FrameData[413] FrameData[414] FrameData[415] FrameData[416] FrameData[417]
+ FrameData[418] FrameData[419] FrameData[41] FrameData[420] FrameData[421] FrameData[422]
+ FrameData[423] FrameData[424] FrameData[425] FrameData[426] FrameData[427] FrameData[428]
+ FrameData[429] FrameData[42] FrameData[430] FrameData[431] FrameData[432] FrameData[433]
+ FrameData[434] FrameData[435] FrameData[436] FrameData[437] FrameData[438] FrameData[439]
+ FrameData[43] FrameData[440] FrameData[441] FrameData[442] FrameData[443] FrameData[444]
+ FrameData[445] FrameData[446] FrameData[447] FrameData[448] FrameData[449] FrameData[44]
+ FrameData[450] FrameData[451] FrameData[452] FrameData[453] FrameData[454] FrameData[455]
+ FrameData[456] FrameData[457] FrameData[458] FrameData[459] FrameData[45] FrameData[460]
+ FrameData[461] FrameData[462] FrameData[463] FrameData[464] FrameData[465] FrameData[466]
+ FrameData[467] FrameData[468] FrameData[469] FrameData[46] FrameData[470] FrameData[471]
+ FrameData[472] FrameData[473] FrameData[474] FrameData[475] FrameData[476] FrameData[477]
+ FrameData[478] FrameData[479] FrameData[47] FrameData[480] FrameData[481] FrameData[482]
+ FrameData[483] FrameData[484] FrameData[485] FrameData[486] FrameData[487] FrameData[488]
+ FrameData[489] FrameData[48] FrameData[490] FrameData[491] FrameData[492] FrameData[493]
+ FrameData[494] FrameData[495] FrameData[496] FrameData[497] FrameData[498] FrameData[499]
+ FrameData[49] FrameData[4] FrameData[500] FrameData[501] FrameData[502] FrameData[503]
+ FrameData[504] FrameData[505] FrameData[506] FrameData[507] FrameData[508] FrameData[509]
+ FrameData[50] FrameData[510] FrameData[511] FrameData[51] FrameData[52] FrameData[53]
+ FrameData[54] FrameData[55] FrameData[56] FrameData[57] FrameData[58] FrameData[59]
+ FrameData[5] FrameData[60] FrameData[61] FrameData[62] FrameData[63] FrameData[64]
+ FrameData[65] FrameData[66] FrameData[67] FrameData[68] FrameData[69] FrameData[6]
+ FrameData[70] FrameData[71] FrameData[72] FrameData[73] FrameData[74] FrameData[75]
+ FrameData[76] FrameData[77] FrameData[78] FrameData[79] FrameData[7] FrameData[80]
+ FrameData[81] FrameData[82] FrameData[83] FrameData[84] FrameData[85] FrameData[86]
+ FrameData[87] FrameData[88] FrameData[89] FrameData[8] FrameData[90] FrameData[91]
+ FrameData[92] FrameData[93] FrameData[94] FrameData[95] FrameData[96] FrameData[97]
+ FrameData[98] FrameData[99] FrameData[9] FrameStrobe[0] FrameStrobe[100] FrameStrobe[101]
+ FrameStrobe[102] FrameStrobe[103] FrameStrobe[104] FrameStrobe[105] FrameStrobe[106]
+ FrameStrobe[107] FrameStrobe[108] FrameStrobe[109] FrameStrobe[10] FrameStrobe[110]
+ FrameStrobe[111] FrameStrobe[112] FrameStrobe[113] FrameStrobe[114] FrameStrobe[115]
+ FrameStrobe[116] FrameStrobe[117] FrameStrobe[118] FrameStrobe[119] FrameStrobe[11]
+ FrameStrobe[120] FrameStrobe[121] FrameStrobe[122] FrameStrobe[123] FrameStrobe[124]
+ FrameStrobe[125] FrameStrobe[126] FrameStrobe[127] FrameStrobe[128] FrameStrobe[129]
+ FrameStrobe[12] FrameStrobe[130] FrameStrobe[131] FrameStrobe[132] FrameStrobe[133]
+ FrameStrobe[134] FrameStrobe[135] FrameStrobe[136] FrameStrobe[137] FrameStrobe[138]
+ FrameStrobe[139] FrameStrobe[13] FrameStrobe[140] FrameStrobe[141] FrameStrobe[142]
+ FrameStrobe[143] FrameStrobe[144] FrameStrobe[145] FrameStrobe[146] FrameStrobe[147]
+ FrameStrobe[148] FrameStrobe[149] FrameStrobe[14] FrameStrobe[150] FrameStrobe[151]
+ FrameStrobe[152] FrameStrobe[153] FrameStrobe[154] FrameStrobe[155] FrameStrobe[156]
+ FrameStrobe[157] FrameStrobe[158] FrameStrobe[159] FrameStrobe[15] FrameStrobe[160]
+ FrameStrobe[161] FrameStrobe[162] FrameStrobe[163] FrameStrobe[164] FrameStrobe[165]
+ FrameStrobe[166] FrameStrobe[167] FrameStrobe[168] FrameStrobe[169] FrameStrobe[16]
+ FrameStrobe[170] FrameStrobe[171] FrameStrobe[172] FrameStrobe[173] FrameStrobe[174]
+ FrameStrobe[175] FrameStrobe[176] FrameStrobe[177] FrameStrobe[178] FrameStrobe[179]
+ FrameStrobe[17] FrameStrobe[180] FrameStrobe[181] FrameStrobe[182] FrameStrobe[183]
+ FrameStrobe[184] FrameStrobe[185] FrameStrobe[186] FrameStrobe[187] FrameStrobe[188]
+ FrameStrobe[189] FrameStrobe[18] FrameStrobe[190] FrameStrobe[191] FrameStrobe[192]
+ FrameStrobe[193] FrameStrobe[194] FrameStrobe[195] FrameStrobe[196] FrameStrobe[197]
+ FrameStrobe[198] FrameStrobe[199] FrameStrobe[19] FrameStrobe[1] FrameStrobe[200]
+ FrameStrobe[201] FrameStrobe[202] FrameStrobe[203] FrameStrobe[204] FrameStrobe[205]
+ FrameStrobe[206] FrameStrobe[207] FrameStrobe[208] FrameStrobe[209] FrameStrobe[20]
+ FrameStrobe[210] FrameStrobe[211] FrameStrobe[212] FrameStrobe[213] FrameStrobe[214]
+ FrameStrobe[215] FrameStrobe[216] FrameStrobe[217] FrameStrobe[218] FrameStrobe[219]
+ FrameStrobe[21] FrameStrobe[22] FrameStrobe[23] FrameStrobe[24] FrameStrobe[25]
+ FrameStrobe[26] FrameStrobe[27] FrameStrobe[28] FrameStrobe[29] FrameStrobe[2] FrameStrobe[30]
+ FrameStrobe[31] FrameStrobe[32] FrameStrobe[33] FrameStrobe[34] FrameStrobe[35]
+ FrameStrobe[36] FrameStrobe[37] FrameStrobe[38] FrameStrobe[39] FrameStrobe[3] FrameStrobe[40]
+ FrameStrobe[41] FrameStrobe[42] FrameStrobe[43] FrameStrobe[44] FrameStrobe[45]
+ FrameStrobe[46] FrameStrobe[47] FrameStrobe[48] FrameStrobe[49] FrameStrobe[4] FrameStrobe[50]
+ FrameStrobe[51] FrameStrobe[52] FrameStrobe[53] FrameStrobe[54] FrameStrobe[55]
+ FrameStrobe[56] FrameStrobe[57] FrameStrobe[58] FrameStrobe[59] FrameStrobe[5] FrameStrobe[60]
+ FrameStrobe[61] FrameStrobe[62] FrameStrobe[63] FrameStrobe[64] FrameStrobe[65]
+ FrameStrobe[66] FrameStrobe[67] FrameStrobe[68] FrameStrobe[69] FrameStrobe[6] FrameStrobe[70]
+ FrameStrobe[71] FrameStrobe[72] FrameStrobe[73] FrameStrobe[74] FrameStrobe[75]
+ FrameStrobe[76] FrameStrobe[77] FrameStrobe[78] FrameStrobe[79] FrameStrobe[7] FrameStrobe[80]
+ FrameStrobe[81] FrameStrobe[82] FrameStrobe[83] FrameStrobe[84] FrameStrobe[85]
+ FrameStrobe[86] FrameStrobe[87] FrameStrobe[88] FrameStrobe[89] FrameStrobe[8] FrameStrobe[90]
+ FrameStrobe[91] FrameStrobe[92] FrameStrobe[93] FrameStrobe[94] FrameStrobe[95]
+ FrameStrobe[96] FrameStrobe[97] FrameStrobe[98] FrameStrobe[99] FrameStrobe[9] Tile_X0Y10_A_I_top
+ Tile_X0Y10_A_O_top Tile_X0Y10_A_T_top Tile_X0Y10_A_config_C_bit0 Tile_X0Y10_A_config_C_bit1
+ Tile_X0Y10_A_config_C_bit2 Tile_X0Y10_A_config_C_bit3 Tile_X0Y10_B_I_top Tile_X0Y10_B_O_top
+ Tile_X0Y10_B_T_top Tile_X0Y10_B_config_C_bit0 Tile_X0Y10_B_config_C_bit1 Tile_X0Y10_B_config_C_bit2
+ Tile_X0Y10_B_config_C_bit3 Tile_X0Y11_A_I_top Tile_X0Y11_A_O_top Tile_X0Y11_A_T_top
+ Tile_X0Y11_A_config_C_bit0 Tile_X0Y11_A_config_C_bit1 Tile_X0Y11_A_config_C_bit2
+ Tile_X0Y11_A_config_C_bit3 Tile_X0Y11_B_I_top Tile_X0Y11_B_O_top Tile_X0Y11_B_T_top
+ Tile_X0Y11_B_config_C_bit0 Tile_X0Y11_B_config_C_bit1 Tile_X0Y11_B_config_C_bit2
+ Tile_X0Y11_B_config_C_bit3 Tile_X0Y12_A_I_top Tile_X0Y12_A_O_top Tile_X0Y12_A_T_top
+ Tile_X0Y12_A_config_C_bit0 Tile_X0Y12_A_config_C_bit1 Tile_X0Y12_A_config_C_bit2
+ Tile_X0Y12_A_config_C_bit3 Tile_X0Y12_B_I_top Tile_X0Y12_B_O_top Tile_X0Y12_B_T_top
+ Tile_X0Y12_B_config_C_bit0 Tile_X0Y12_B_config_C_bit1 Tile_X0Y12_B_config_C_bit2
+ Tile_X0Y12_B_config_C_bit3 Tile_X0Y13_A_I_top Tile_X0Y13_A_O_top Tile_X0Y13_A_T_top
+ Tile_X0Y13_A_config_C_bit0 Tile_X0Y13_A_config_C_bit1 Tile_X0Y13_A_config_C_bit2
+ Tile_X0Y13_A_config_C_bit3 Tile_X0Y13_B_I_top Tile_X0Y13_B_O_top Tile_X0Y13_B_T_top
+ Tile_X0Y13_B_config_C_bit0 Tile_X0Y13_B_config_C_bit1 Tile_X0Y13_B_config_C_bit2
+ Tile_X0Y13_B_config_C_bit3 Tile_X0Y14_A_I_top Tile_X0Y14_A_O_top Tile_X0Y14_A_T_top
+ Tile_X0Y14_A_config_C_bit0 Tile_X0Y14_A_config_C_bit1 Tile_X0Y14_A_config_C_bit2
+ Tile_X0Y14_A_config_C_bit3 Tile_X0Y14_B_I_top Tile_X0Y14_B_O_top Tile_X0Y14_B_T_top
+ Tile_X0Y14_B_config_C_bit0 Tile_X0Y14_B_config_C_bit1 Tile_X0Y14_B_config_C_bit2
+ Tile_X0Y14_B_config_C_bit3 Tile_X0Y1_A_I_top Tile_X0Y1_A_O_top Tile_X0Y1_A_T_top
+ Tile_X0Y1_A_config_C_bit0 Tile_X0Y1_A_config_C_bit1 Tile_X0Y1_A_config_C_bit2 Tile_X0Y1_A_config_C_bit3
+ Tile_X0Y1_B_I_top Tile_X0Y1_B_O_top Tile_X0Y1_B_T_top Tile_X0Y1_B_config_C_bit0
+ Tile_X0Y1_B_config_C_bit1 Tile_X0Y1_B_config_C_bit2 Tile_X0Y1_B_config_C_bit3 Tile_X0Y2_A_I_top
+ Tile_X0Y2_A_O_top Tile_X0Y2_A_T_top Tile_X0Y2_A_config_C_bit0 Tile_X0Y2_A_config_C_bit1
+ Tile_X0Y2_A_config_C_bit2 Tile_X0Y2_A_config_C_bit3 Tile_X0Y2_B_I_top Tile_X0Y2_B_O_top
+ Tile_X0Y2_B_T_top Tile_X0Y2_B_config_C_bit0 Tile_X0Y2_B_config_C_bit1 Tile_X0Y2_B_config_C_bit2
+ Tile_X0Y2_B_config_C_bit3 Tile_X0Y3_A_I_top Tile_X0Y3_A_O_top Tile_X0Y3_A_T_top
+ Tile_X0Y3_A_config_C_bit0 Tile_X0Y3_A_config_C_bit1 Tile_X0Y3_A_config_C_bit2 Tile_X0Y3_A_config_C_bit3
+ Tile_X0Y3_B_I_top Tile_X0Y3_B_O_top Tile_X0Y3_B_T_top Tile_X0Y3_B_config_C_bit0
+ Tile_X0Y3_B_config_C_bit1 Tile_X0Y3_B_config_C_bit2 Tile_X0Y3_B_config_C_bit3 Tile_X0Y4_A_I_top
+ Tile_X0Y4_A_O_top Tile_X0Y4_A_T_top Tile_X0Y4_A_config_C_bit0 Tile_X0Y4_A_config_C_bit1
+ Tile_X0Y4_A_config_C_bit2 Tile_X0Y4_A_config_C_bit3 Tile_X0Y4_B_I_top Tile_X0Y4_B_O_top
+ Tile_X0Y4_B_T_top Tile_X0Y4_B_config_C_bit0 Tile_X0Y4_B_config_C_bit1 Tile_X0Y4_B_config_C_bit2
+ Tile_X0Y4_B_config_C_bit3 Tile_X0Y5_A_I_top Tile_X0Y5_A_O_top Tile_X0Y5_A_T_top
+ Tile_X0Y5_A_config_C_bit0 Tile_X0Y5_A_config_C_bit1 Tile_X0Y5_A_config_C_bit2 Tile_X0Y5_A_config_C_bit3
+ Tile_X0Y5_B_I_top Tile_X0Y5_B_O_top Tile_X0Y5_B_T_top Tile_X0Y5_B_config_C_bit0
+ Tile_X0Y5_B_config_C_bit1 Tile_X0Y5_B_config_C_bit2 Tile_X0Y5_B_config_C_bit3 Tile_X0Y6_A_I_top
+ Tile_X0Y6_A_O_top Tile_X0Y6_A_T_top Tile_X0Y6_A_config_C_bit0 Tile_X0Y6_A_config_C_bit1
+ Tile_X0Y6_A_config_C_bit2 Tile_X0Y6_A_config_C_bit3 Tile_X0Y6_B_I_top Tile_X0Y6_B_O_top
+ Tile_X0Y6_B_T_top Tile_X0Y6_B_config_C_bit0 Tile_X0Y6_B_config_C_bit1 Tile_X0Y6_B_config_C_bit2
+ Tile_X0Y6_B_config_C_bit3 Tile_X0Y7_A_I_top Tile_X0Y7_A_O_top Tile_X0Y7_A_T_top
+ Tile_X0Y7_A_config_C_bit0 Tile_X0Y7_A_config_C_bit1 Tile_X0Y7_A_config_C_bit2 Tile_X0Y7_A_config_C_bit3
+ Tile_X0Y7_B_I_top Tile_X0Y7_B_O_top Tile_X0Y7_B_T_top Tile_X0Y7_B_config_C_bit0
+ Tile_X0Y7_B_config_C_bit1 Tile_X0Y7_B_config_C_bit2 Tile_X0Y7_B_config_C_bit3 Tile_X0Y8_A_I_top
+ Tile_X0Y8_A_O_top Tile_X0Y8_A_T_top Tile_X0Y8_A_config_C_bit0 Tile_X0Y8_A_config_C_bit1
+ Tile_X0Y8_A_config_C_bit2 Tile_X0Y8_A_config_C_bit3 Tile_X0Y8_B_I_top Tile_X0Y8_B_O_top
+ Tile_X0Y8_B_T_top Tile_X0Y8_B_config_C_bit0 Tile_X0Y8_B_config_C_bit1 Tile_X0Y8_B_config_C_bit2
+ Tile_X0Y8_B_config_C_bit3 Tile_X0Y9_A_I_top Tile_X0Y9_A_O_top Tile_X0Y9_A_T_top
+ Tile_X0Y9_A_config_C_bit0 Tile_X0Y9_A_config_C_bit1 Tile_X0Y9_A_config_C_bit2 Tile_X0Y9_A_config_C_bit3
+ Tile_X0Y9_B_I_top Tile_X0Y9_B_O_top Tile_X0Y9_B_T_top Tile_X0Y9_B_config_C_bit0
+ Tile_X0Y9_B_config_C_bit1 Tile_X0Y9_B_config_C_bit2 Tile_X0Y9_B_config_C_bit3 Tile_X10Y10_ADDR_SRAM0
+ Tile_X10Y10_ADDR_SRAM1 Tile_X10Y10_ADDR_SRAM2 Tile_X10Y10_ADDR_SRAM3 Tile_X10Y10_ADDR_SRAM4
+ Tile_X10Y10_ADDR_SRAM5 Tile_X10Y10_ADDR_SRAM6 Tile_X10Y10_ADDR_SRAM7 Tile_X10Y10_ADDR_SRAM8
+ Tile_X10Y10_ADDR_SRAM9 Tile_X10Y10_BM_SRAM0 Tile_X10Y10_BM_SRAM1 Tile_X10Y10_BM_SRAM10
+ Tile_X10Y10_BM_SRAM11 Tile_X10Y10_BM_SRAM12 Tile_X10Y10_BM_SRAM13 Tile_X10Y10_BM_SRAM14
+ Tile_X10Y10_BM_SRAM15 Tile_X10Y10_BM_SRAM16 Tile_X10Y10_BM_SRAM17 Tile_X10Y10_BM_SRAM18
+ Tile_X10Y10_BM_SRAM19 Tile_X10Y10_BM_SRAM2 Tile_X10Y10_BM_SRAM20 Tile_X10Y10_BM_SRAM21
+ Tile_X10Y10_BM_SRAM22 Tile_X10Y10_BM_SRAM23 Tile_X10Y10_BM_SRAM24 Tile_X10Y10_BM_SRAM25
+ Tile_X10Y10_BM_SRAM26 Tile_X10Y10_BM_SRAM27 Tile_X10Y10_BM_SRAM28 Tile_X10Y10_BM_SRAM29
+ Tile_X10Y10_BM_SRAM3 Tile_X10Y10_BM_SRAM30 Tile_X10Y10_BM_SRAM31 Tile_X10Y10_BM_SRAM4
+ Tile_X10Y10_BM_SRAM5 Tile_X10Y10_BM_SRAM6 Tile_X10Y10_BM_SRAM7 Tile_X10Y10_BM_SRAM8
+ Tile_X10Y10_BM_SRAM9 Tile_X10Y10_CLK_SRAM Tile_X10Y10_CONFIGURED_top Tile_X10Y10_DIN_SRAM0
+ Tile_X10Y10_DIN_SRAM1 Tile_X10Y10_DIN_SRAM10 Tile_X10Y10_DIN_SRAM11 Tile_X10Y10_DIN_SRAM12
+ Tile_X10Y10_DIN_SRAM13 Tile_X10Y10_DIN_SRAM14 Tile_X10Y10_DIN_SRAM15 Tile_X10Y10_DIN_SRAM16
+ Tile_X10Y10_DIN_SRAM17 Tile_X10Y10_DIN_SRAM18 Tile_X10Y10_DIN_SRAM19 Tile_X10Y10_DIN_SRAM2
+ Tile_X10Y10_DIN_SRAM20 Tile_X10Y10_DIN_SRAM21 Tile_X10Y10_DIN_SRAM22 Tile_X10Y10_DIN_SRAM23
+ Tile_X10Y10_DIN_SRAM24 Tile_X10Y10_DIN_SRAM25 Tile_X10Y10_DIN_SRAM26 Tile_X10Y10_DIN_SRAM27
+ Tile_X10Y10_DIN_SRAM28 Tile_X10Y10_DIN_SRAM29 Tile_X10Y10_DIN_SRAM3 Tile_X10Y10_DIN_SRAM30
+ Tile_X10Y10_DIN_SRAM31 Tile_X10Y10_DIN_SRAM4 Tile_X10Y10_DIN_SRAM5 Tile_X10Y10_DIN_SRAM6
+ Tile_X10Y10_DIN_SRAM7 Tile_X10Y10_DIN_SRAM8 Tile_X10Y10_DIN_SRAM9 Tile_X10Y10_DOUT_SRAM0
+ Tile_X10Y10_DOUT_SRAM1 Tile_X10Y10_DOUT_SRAM10 Tile_X10Y10_DOUT_SRAM11 Tile_X10Y10_DOUT_SRAM12
+ Tile_X10Y10_DOUT_SRAM13 Tile_X10Y10_DOUT_SRAM14 Tile_X10Y10_DOUT_SRAM15 Tile_X10Y10_DOUT_SRAM16
+ Tile_X10Y10_DOUT_SRAM17 Tile_X10Y10_DOUT_SRAM18 Tile_X10Y10_DOUT_SRAM19 Tile_X10Y10_DOUT_SRAM2
+ Tile_X10Y10_DOUT_SRAM20 Tile_X10Y10_DOUT_SRAM21 Tile_X10Y10_DOUT_SRAM22 Tile_X10Y10_DOUT_SRAM23
+ Tile_X10Y10_DOUT_SRAM24 Tile_X10Y10_DOUT_SRAM25 Tile_X10Y10_DOUT_SRAM26 Tile_X10Y10_DOUT_SRAM27
+ Tile_X10Y10_DOUT_SRAM28 Tile_X10Y10_DOUT_SRAM29 Tile_X10Y10_DOUT_SRAM3 Tile_X10Y10_DOUT_SRAM30
+ Tile_X10Y10_DOUT_SRAM31 Tile_X10Y10_DOUT_SRAM4 Tile_X10Y10_DOUT_SRAM5 Tile_X10Y10_DOUT_SRAM6
+ Tile_X10Y10_DOUT_SRAM7 Tile_X10Y10_DOUT_SRAM8 Tile_X10Y10_DOUT_SRAM9 Tile_X10Y10_MEN_SRAM
+ Tile_X10Y10_REN_SRAM Tile_X10Y10_TIE_HIGH_SRAM Tile_X10Y10_TIE_LOW_SRAM Tile_X10Y10_WEN_SRAM
+ Tile_X10Y12_ADDR_SRAM0 Tile_X10Y12_ADDR_SRAM1 Tile_X10Y12_ADDR_SRAM2 Tile_X10Y12_ADDR_SRAM3
+ Tile_X10Y12_ADDR_SRAM4 Tile_X10Y12_ADDR_SRAM5 Tile_X10Y12_ADDR_SRAM6 Tile_X10Y12_ADDR_SRAM7
+ Tile_X10Y12_ADDR_SRAM8 Tile_X10Y12_ADDR_SRAM9 Tile_X10Y12_BM_SRAM0 Tile_X10Y12_BM_SRAM1
+ Tile_X10Y12_BM_SRAM10 Tile_X10Y12_BM_SRAM11 Tile_X10Y12_BM_SRAM12 Tile_X10Y12_BM_SRAM13
+ Tile_X10Y12_BM_SRAM14 Tile_X10Y12_BM_SRAM15 Tile_X10Y12_BM_SRAM16 Tile_X10Y12_BM_SRAM17
+ Tile_X10Y12_BM_SRAM18 Tile_X10Y12_BM_SRAM19 Tile_X10Y12_BM_SRAM2 Tile_X10Y12_BM_SRAM20
+ Tile_X10Y12_BM_SRAM21 Tile_X10Y12_BM_SRAM22 Tile_X10Y12_BM_SRAM23 Tile_X10Y12_BM_SRAM24
+ Tile_X10Y12_BM_SRAM25 Tile_X10Y12_BM_SRAM26 Tile_X10Y12_BM_SRAM27 Tile_X10Y12_BM_SRAM28
+ Tile_X10Y12_BM_SRAM29 Tile_X10Y12_BM_SRAM3 Tile_X10Y12_BM_SRAM30 Tile_X10Y12_BM_SRAM31
+ Tile_X10Y12_BM_SRAM4 Tile_X10Y12_BM_SRAM5 Tile_X10Y12_BM_SRAM6 Tile_X10Y12_BM_SRAM7
+ Tile_X10Y12_BM_SRAM8 Tile_X10Y12_BM_SRAM9 Tile_X10Y12_CLK_SRAM Tile_X10Y12_CONFIGURED_top
+ Tile_X10Y12_DIN_SRAM0 Tile_X10Y12_DIN_SRAM1 Tile_X10Y12_DIN_SRAM10 Tile_X10Y12_DIN_SRAM11
+ Tile_X10Y12_DIN_SRAM12 Tile_X10Y12_DIN_SRAM13 Tile_X10Y12_DIN_SRAM14 Tile_X10Y12_DIN_SRAM15
+ Tile_X10Y12_DIN_SRAM16 Tile_X10Y12_DIN_SRAM17 Tile_X10Y12_DIN_SRAM18 Tile_X10Y12_DIN_SRAM19
+ Tile_X10Y12_DIN_SRAM2 Tile_X10Y12_DIN_SRAM20 Tile_X10Y12_DIN_SRAM21 Tile_X10Y12_DIN_SRAM22
+ Tile_X10Y12_DIN_SRAM23 Tile_X10Y12_DIN_SRAM24 Tile_X10Y12_DIN_SRAM25 Tile_X10Y12_DIN_SRAM26
+ Tile_X10Y12_DIN_SRAM27 Tile_X10Y12_DIN_SRAM28 Tile_X10Y12_DIN_SRAM29 Tile_X10Y12_DIN_SRAM3
+ Tile_X10Y12_DIN_SRAM30 Tile_X10Y12_DIN_SRAM31 Tile_X10Y12_DIN_SRAM4 Tile_X10Y12_DIN_SRAM5
+ Tile_X10Y12_DIN_SRAM6 Tile_X10Y12_DIN_SRAM7 Tile_X10Y12_DIN_SRAM8 Tile_X10Y12_DIN_SRAM9
+ Tile_X10Y12_DOUT_SRAM0 Tile_X10Y12_DOUT_SRAM1 Tile_X10Y12_DOUT_SRAM10 Tile_X10Y12_DOUT_SRAM11
+ Tile_X10Y12_DOUT_SRAM12 Tile_X10Y12_DOUT_SRAM13 Tile_X10Y12_DOUT_SRAM14 Tile_X10Y12_DOUT_SRAM15
+ Tile_X10Y12_DOUT_SRAM16 Tile_X10Y12_DOUT_SRAM17 Tile_X10Y12_DOUT_SRAM18 Tile_X10Y12_DOUT_SRAM19
+ Tile_X10Y12_DOUT_SRAM2 Tile_X10Y12_DOUT_SRAM20 Tile_X10Y12_DOUT_SRAM21 Tile_X10Y12_DOUT_SRAM22
+ Tile_X10Y12_DOUT_SRAM23 Tile_X10Y12_DOUT_SRAM24 Tile_X10Y12_DOUT_SRAM25 Tile_X10Y12_DOUT_SRAM26
+ Tile_X10Y12_DOUT_SRAM27 Tile_X10Y12_DOUT_SRAM28 Tile_X10Y12_DOUT_SRAM29 Tile_X10Y12_DOUT_SRAM3
+ Tile_X10Y12_DOUT_SRAM30 Tile_X10Y12_DOUT_SRAM31 Tile_X10Y12_DOUT_SRAM4 Tile_X10Y12_DOUT_SRAM5
+ Tile_X10Y12_DOUT_SRAM6 Tile_X10Y12_DOUT_SRAM7 Tile_X10Y12_DOUT_SRAM8 Tile_X10Y12_DOUT_SRAM9
+ Tile_X10Y12_MEN_SRAM Tile_X10Y12_REN_SRAM Tile_X10Y12_TIE_HIGH_SRAM Tile_X10Y12_TIE_LOW_SRAM
+ Tile_X10Y12_WEN_SRAM Tile_X10Y14_ADDR_SRAM0 Tile_X10Y14_ADDR_SRAM1 Tile_X10Y14_ADDR_SRAM2
+ Tile_X10Y14_ADDR_SRAM3 Tile_X10Y14_ADDR_SRAM4 Tile_X10Y14_ADDR_SRAM5 Tile_X10Y14_ADDR_SRAM6
+ Tile_X10Y14_ADDR_SRAM7 Tile_X10Y14_ADDR_SRAM8 Tile_X10Y14_ADDR_SRAM9 Tile_X10Y14_BM_SRAM0
+ Tile_X10Y14_BM_SRAM1 Tile_X10Y14_BM_SRAM10 Tile_X10Y14_BM_SRAM11 Tile_X10Y14_BM_SRAM12
+ Tile_X10Y14_BM_SRAM13 Tile_X10Y14_BM_SRAM14 Tile_X10Y14_BM_SRAM15 Tile_X10Y14_BM_SRAM16
+ Tile_X10Y14_BM_SRAM17 Tile_X10Y14_BM_SRAM18 Tile_X10Y14_BM_SRAM19 Tile_X10Y14_BM_SRAM2
+ Tile_X10Y14_BM_SRAM20 Tile_X10Y14_BM_SRAM21 Tile_X10Y14_BM_SRAM22 Tile_X10Y14_BM_SRAM23
+ Tile_X10Y14_BM_SRAM24 Tile_X10Y14_BM_SRAM25 Tile_X10Y14_BM_SRAM26 Tile_X10Y14_BM_SRAM27
+ Tile_X10Y14_BM_SRAM28 Tile_X10Y14_BM_SRAM29 Tile_X10Y14_BM_SRAM3 Tile_X10Y14_BM_SRAM30
+ Tile_X10Y14_BM_SRAM31 Tile_X10Y14_BM_SRAM4 Tile_X10Y14_BM_SRAM5 Tile_X10Y14_BM_SRAM6
+ Tile_X10Y14_BM_SRAM7 Tile_X10Y14_BM_SRAM8 Tile_X10Y14_BM_SRAM9 Tile_X10Y14_CLK_SRAM
+ Tile_X10Y14_CONFIGURED_top Tile_X10Y14_DIN_SRAM0 Tile_X10Y14_DIN_SRAM1 Tile_X10Y14_DIN_SRAM10
+ Tile_X10Y14_DIN_SRAM11 Tile_X10Y14_DIN_SRAM12 Tile_X10Y14_DIN_SRAM13 Tile_X10Y14_DIN_SRAM14
+ Tile_X10Y14_DIN_SRAM15 Tile_X10Y14_DIN_SRAM16 Tile_X10Y14_DIN_SRAM17 Tile_X10Y14_DIN_SRAM18
+ Tile_X10Y14_DIN_SRAM19 Tile_X10Y14_DIN_SRAM2 Tile_X10Y14_DIN_SRAM20 Tile_X10Y14_DIN_SRAM21
+ Tile_X10Y14_DIN_SRAM22 Tile_X10Y14_DIN_SRAM23 Tile_X10Y14_DIN_SRAM24 Tile_X10Y14_DIN_SRAM25
+ Tile_X10Y14_DIN_SRAM26 Tile_X10Y14_DIN_SRAM27 Tile_X10Y14_DIN_SRAM28 Tile_X10Y14_DIN_SRAM29
+ Tile_X10Y14_DIN_SRAM3 Tile_X10Y14_DIN_SRAM30 Tile_X10Y14_DIN_SRAM31 Tile_X10Y14_DIN_SRAM4
+ Tile_X10Y14_DIN_SRAM5 Tile_X10Y14_DIN_SRAM6 Tile_X10Y14_DIN_SRAM7 Tile_X10Y14_DIN_SRAM8
+ Tile_X10Y14_DIN_SRAM9 Tile_X10Y14_DOUT_SRAM0 Tile_X10Y14_DOUT_SRAM1 Tile_X10Y14_DOUT_SRAM10
+ Tile_X10Y14_DOUT_SRAM11 Tile_X10Y14_DOUT_SRAM12 Tile_X10Y14_DOUT_SRAM13 Tile_X10Y14_DOUT_SRAM14
+ Tile_X10Y14_DOUT_SRAM15 Tile_X10Y14_DOUT_SRAM16 Tile_X10Y14_DOUT_SRAM17 Tile_X10Y14_DOUT_SRAM18
+ Tile_X10Y14_DOUT_SRAM19 Tile_X10Y14_DOUT_SRAM2 Tile_X10Y14_DOUT_SRAM20 Tile_X10Y14_DOUT_SRAM21
+ Tile_X10Y14_DOUT_SRAM22 Tile_X10Y14_DOUT_SRAM23 Tile_X10Y14_DOUT_SRAM24 Tile_X10Y14_DOUT_SRAM25
+ Tile_X10Y14_DOUT_SRAM26 Tile_X10Y14_DOUT_SRAM27 Tile_X10Y14_DOUT_SRAM28 Tile_X10Y14_DOUT_SRAM29
+ Tile_X10Y14_DOUT_SRAM3 Tile_X10Y14_DOUT_SRAM30 Tile_X10Y14_DOUT_SRAM31 Tile_X10Y14_DOUT_SRAM4
+ Tile_X10Y14_DOUT_SRAM5 Tile_X10Y14_DOUT_SRAM6 Tile_X10Y14_DOUT_SRAM7 Tile_X10Y14_DOUT_SRAM8
+ Tile_X10Y14_DOUT_SRAM9 Tile_X10Y14_MEN_SRAM Tile_X10Y14_REN_SRAM Tile_X10Y14_TIE_HIGH_SRAM
+ Tile_X10Y14_TIE_LOW_SRAM Tile_X10Y14_WEN_SRAM Tile_X10Y2_ADDR_SRAM0 Tile_X10Y2_ADDR_SRAM1
+ Tile_X10Y2_ADDR_SRAM2 Tile_X10Y2_ADDR_SRAM3 Tile_X10Y2_ADDR_SRAM4 Tile_X10Y2_ADDR_SRAM5
+ Tile_X10Y2_ADDR_SRAM6 Tile_X10Y2_ADDR_SRAM7 Tile_X10Y2_ADDR_SRAM8 Tile_X10Y2_ADDR_SRAM9
+ Tile_X10Y2_BM_SRAM0 Tile_X10Y2_BM_SRAM1 Tile_X10Y2_BM_SRAM10 Tile_X10Y2_BM_SRAM11
+ Tile_X10Y2_BM_SRAM12 Tile_X10Y2_BM_SRAM13 Tile_X10Y2_BM_SRAM14 Tile_X10Y2_BM_SRAM15
+ Tile_X10Y2_BM_SRAM16 Tile_X10Y2_BM_SRAM17 Tile_X10Y2_BM_SRAM18 Tile_X10Y2_BM_SRAM19
+ Tile_X10Y2_BM_SRAM2 Tile_X10Y2_BM_SRAM20 Tile_X10Y2_BM_SRAM21 Tile_X10Y2_BM_SRAM22
+ Tile_X10Y2_BM_SRAM23 Tile_X10Y2_BM_SRAM24 Tile_X10Y2_BM_SRAM25 Tile_X10Y2_BM_SRAM26
+ Tile_X10Y2_BM_SRAM27 Tile_X10Y2_BM_SRAM28 Tile_X10Y2_BM_SRAM29 Tile_X10Y2_BM_SRAM3
+ Tile_X10Y2_BM_SRAM30 Tile_X10Y2_BM_SRAM31 Tile_X10Y2_BM_SRAM4 Tile_X10Y2_BM_SRAM5
+ Tile_X10Y2_BM_SRAM6 Tile_X10Y2_BM_SRAM7 Tile_X10Y2_BM_SRAM8 Tile_X10Y2_BM_SRAM9
+ Tile_X10Y2_CLK_SRAM Tile_X10Y2_CONFIGURED_top Tile_X10Y2_DIN_SRAM0 Tile_X10Y2_DIN_SRAM1
+ Tile_X10Y2_DIN_SRAM10 Tile_X10Y2_DIN_SRAM11 Tile_X10Y2_DIN_SRAM12 Tile_X10Y2_DIN_SRAM13
+ Tile_X10Y2_DIN_SRAM14 Tile_X10Y2_DIN_SRAM15 Tile_X10Y2_DIN_SRAM16 Tile_X10Y2_DIN_SRAM17
+ Tile_X10Y2_DIN_SRAM18 Tile_X10Y2_DIN_SRAM19 Tile_X10Y2_DIN_SRAM2 Tile_X10Y2_DIN_SRAM20
+ Tile_X10Y2_DIN_SRAM21 Tile_X10Y2_DIN_SRAM22 Tile_X10Y2_DIN_SRAM23 Tile_X10Y2_DIN_SRAM24
+ Tile_X10Y2_DIN_SRAM25 Tile_X10Y2_DIN_SRAM26 Tile_X10Y2_DIN_SRAM27 Tile_X10Y2_DIN_SRAM28
+ Tile_X10Y2_DIN_SRAM29 Tile_X10Y2_DIN_SRAM3 Tile_X10Y2_DIN_SRAM30 Tile_X10Y2_DIN_SRAM31
+ Tile_X10Y2_DIN_SRAM4 Tile_X10Y2_DIN_SRAM5 Tile_X10Y2_DIN_SRAM6 Tile_X10Y2_DIN_SRAM7
+ Tile_X10Y2_DIN_SRAM8 Tile_X10Y2_DIN_SRAM9 Tile_X10Y2_DOUT_SRAM0 Tile_X10Y2_DOUT_SRAM1
+ Tile_X10Y2_DOUT_SRAM10 Tile_X10Y2_DOUT_SRAM11 Tile_X10Y2_DOUT_SRAM12 Tile_X10Y2_DOUT_SRAM13
+ Tile_X10Y2_DOUT_SRAM14 Tile_X10Y2_DOUT_SRAM15 Tile_X10Y2_DOUT_SRAM16 Tile_X10Y2_DOUT_SRAM17
+ Tile_X10Y2_DOUT_SRAM18 Tile_X10Y2_DOUT_SRAM19 Tile_X10Y2_DOUT_SRAM2 Tile_X10Y2_DOUT_SRAM20
+ Tile_X10Y2_DOUT_SRAM21 Tile_X10Y2_DOUT_SRAM22 Tile_X10Y2_DOUT_SRAM23 Tile_X10Y2_DOUT_SRAM24
+ Tile_X10Y2_DOUT_SRAM25 Tile_X10Y2_DOUT_SRAM26 Tile_X10Y2_DOUT_SRAM27 Tile_X10Y2_DOUT_SRAM28
+ Tile_X10Y2_DOUT_SRAM29 Tile_X10Y2_DOUT_SRAM3 Tile_X10Y2_DOUT_SRAM30 Tile_X10Y2_DOUT_SRAM31
+ Tile_X10Y2_DOUT_SRAM4 Tile_X10Y2_DOUT_SRAM5 Tile_X10Y2_DOUT_SRAM6 Tile_X10Y2_DOUT_SRAM7
+ Tile_X10Y2_DOUT_SRAM8 Tile_X10Y2_DOUT_SRAM9 Tile_X10Y2_MEN_SRAM Tile_X10Y2_REN_SRAM
+ Tile_X10Y2_TIE_HIGH_SRAM Tile_X10Y2_TIE_LOW_SRAM Tile_X10Y2_WEN_SRAM Tile_X10Y4_ADDR_SRAM0
+ Tile_X10Y4_ADDR_SRAM1 Tile_X10Y4_ADDR_SRAM2 Tile_X10Y4_ADDR_SRAM3 Tile_X10Y4_ADDR_SRAM4
+ Tile_X10Y4_ADDR_SRAM5 Tile_X10Y4_ADDR_SRAM6 Tile_X10Y4_ADDR_SRAM7 Tile_X10Y4_ADDR_SRAM8
+ Tile_X10Y4_ADDR_SRAM9 Tile_X10Y4_BM_SRAM0 Tile_X10Y4_BM_SRAM1 Tile_X10Y4_BM_SRAM10
+ Tile_X10Y4_BM_SRAM11 Tile_X10Y4_BM_SRAM12 Tile_X10Y4_BM_SRAM13 Tile_X10Y4_BM_SRAM14
+ Tile_X10Y4_BM_SRAM15 Tile_X10Y4_BM_SRAM16 Tile_X10Y4_BM_SRAM17 Tile_X10Y4_BM_SRAM18
+ Tile_X10Y4_BM_SRAM19 Tile_X10Y4_BM_SRAM2 Tile_X10Y4_BM_SRAM20 Tile_X10Y4_BM_SRAM21
+ Tile_X10Y4_BM_SRAM22 Tile_X10Y4_BM_SRAM23 Tile_X10Y4_BM_SRAM24 Tile_X10Y4_BM_SRAM25
+ Tile_X10Y4_BM_SRAM26 Tile_X10Y4_BM_SRAM27 Tile_X10Y4_BM_SRAM28 Tile_X10Y4_BM_SRAM29
+ Tile_X10Y4_BM_SRAM3 Tile_X10Y4_BM_SRAM30 Tile_X10Y4_BM_SRAM31 Tile_X10Y4_BM_SRAM4
+ Tile_X10Y4_BM_SRAM5 Tile_X10Y4_BM_SRAM6 Tile_X10Y4_BM_SRAM7 Tile_X10Y4_BM_SRAM8
+ Tile_X10Y4_BM_SRAM9 Tile_X10Y4_CLK_SRAM Tile_X10Y4_CONFIGURED_top Tile_X10Y4_DIN_SRAM0
+ Tile_X10Y4_DIN_SRAM1 Tile_X10Y4_DIN_SRAM10 Tile_X10Y4_DIN_SRAM11 Tile_X10Y4_DIN_SRAM12
+ Tile_X10Y4_DIN_SRAM13 Tile_X10Y4_DIN_SRAM14 Tile_X10Y4_DIN_SRAM15 Tile_X10Y4_DIN_SRAM16
+ Tile_X10Y4_DIN_SRAM17 Tile_X10Y4_DIN_SRAM18 Tile_X10Y4_DIN_SRAM19 Tile_X10Y4_DIN_SRAM2
+ Tile_X10Y4_DIN_SRAM20 Tile_X10Y4_DIN_SRAM21 Tile_X10Y4_DIN_SRAM22 Tile_X10Y4_DIN_SRAM23
+ Tile_X10Y4_DIN_SRAM24 Tile_X10Y4_DIN_SRAM25 Tile_X10Y4_DIN_SRAM26 Tile_X10Y4_DIN_SRAM27
+ Tile_X10Y4_DIN_SRAM28 Tile_X10Y4_DIN_SRAM29 Tile_X10Y4_DIN_SRAM3 Tile_X10Y4_DIN_SRAM30
+ Tile_X10Y4_DIN_SRAM31 Tile_X10Y4_DIN_SRAM4 Tile_X10Y4_DIN_SRAM5 Tile_X10Y4_DIN_SRAM6
+ Tile_X10Y4_DIN_SRAM7 Tile_X10Y4_DIN_SRAM8 Tile_X10Y4_DIN_SRAM9 Tile_X10Y4_DOUT_SRAM0
+ Tile_X10Y4_DOUT_SRAM1 Tile_X10Y4_DOUT_SRAM10 Tile_X10Y4_DOUT_SRAM11 Tile_X10Y4_DOUT_SRAM12
+ Tile_X10Y4_DOUT_SRAM13 Tile_X10Y4_DOUT_SRAM14 Tile_X10Y4_DOUT_SRAM15 Tile_X10Y4_DOUT_SRAM16
+ Tile_X10Y4_DOUT_SRAM17 Tile_X10Y4_DOUT_SRAM18 Tile_X10Y4_DOUT_SRAM19 Tile_X10Y4_DOUT_SRAM2
+ Tile_X10Y4_DOUT_SRAM20 Tile_X10Y4_DOUT_SRAM21 Tile_X10Y4_DOUT_SRAM22 Tile_X10Y4_DOUT_SRAM23
+ Tile_X10Y4_DOUT_SRAM24 Tile_X10Y4_DOUT_SRAM25 Tile_X10Y4_DOUT_SRAM26 Tile_X10Y4_DOUT_SRAM27
+ Tile_X10Y4_DOUT_SRAM28 Tile_X10Y4_DOUT_SRAM29 Tile_X10Y4_DOUT_SRAM3 Tile_X10Y4_DOUT_SRAM30
+ Tile_X10Y4_DOUT_SRAM31 Tile_X10Y4_DOUT_SRAM4 Tile_X10Y4_DOUT_SRAM5 Tile_X10Y4_DOUT_SRAM6
+ Tile_X10Y4_DOUT_SRAM7 Tile_X10Y4_DOUT_SRAM8 Tile_X10Y4_DOUT_SRAM9 Tile_X10Y4_MEN_SRAM
+ Tile_X10Y4_REN_SRAM Tile_X10Y4_TIE_HIGH_SRAM Tile_X10Y4_TIE_LOW_SRAM Tile_X10Y4_WEN_SRAM
+ Tile_X10Y6_ADDR_SRAM0 Tile_X10Y6_ADDR_SRAM1 Tile_X10Y6_ADDR_SRAM2 Tile_X10Y6_ADDR_SRAM3
+ Tile_X10Y6_ADDR_SRAM4 Tile_X10Y6_ADDR_SRAM5 Tile_X10Y6_ADDR_SRAM6 Tile_X10Y6_ADDR_SRAM7
+ Tile_X10Y6_ADDR_SRAM8 Tile_X10Y6_ADDR_SRAM9 Tile_X10Y6_BM_SRAM0 Tile_X10Y6_BM_SRAM1
+ Tile_X10Y6_BM_SRAM10 Tile_X10Y6_BM_SRAM11 Tile_X10Y6_BM_SRAM12 Tile_X10Y6_BM_SRAM13
+ Tile_X10Y6_BM_SRAM14 Tile_X10Y6_BM_SRAM15 Tile_X10Y6_BM_SRAM16 Tile_X10Y6_BM_SRAM17
+ Tile_X10Y6_BM_SRAM18 Tile_X10Y6_BM_SRAM19 Tile_X10Y6_BM_SRAM2 Tile_X10Y6_BM_SRAM20
+ Tile_X10Y6_BM_SRAM21 Tile_X10Y6_BM_SRAM22 Tile_X10Y6_BM_SRAM23 Tile_X10Y6_BM_SRAM24
+ Tile_X10Y6_BM_SRAM25 Tile_X10Y6_BM_SRAM26 Tile_X10Y6_BM_SRAM27 Tile_X10Y6_BM_SRAM28
+ Tile_X10Y6_BM_SRAM29 Tile_X10Y6_BM_SRAM3 Tile_X10Y6_BM_SRAM30 Tile_X10Y6_BM_SRAM31
+ Tile_X10Y6_BM_SRAM4 Tile_X10Y6_BM_SRAM5 Tile_X10Y6_BM_SRAM6 Tile_X10Y6_BM_SRAM7
+ Tile_X10Y6_BM_SRAM8 Tile_X10Y6_BM_SRAM9 Tile_X10Y6_CLK_SRAM Tile_X10Y6_CONFIGURED_top
+ Tile_X10Y6_DIN_SRAM0 Tile_X10Y6_DIN_SRAM1 Tile_X10Y6_DIN_SRAM10 Tile_X10Y6_DIN_SRAM11
+ Tile_X10Y6_DIN_SRAM12 Tile_X10Y6_DIN_SRAM13 Tile_X10Y6_DIN_SRAM14 Tile_X10Y6_DIN_SRAM15
+ Tile_X10Y6_DIN_SRAM16 Tile_X10Y6_DIN_SRAM17 Tile_X10Y6_DIN_SRAM18 Tile_X10Y6_DIN_SRAM19
+ Tile_X10Y6_DIN_SRAM2 Tile_X10Y6_DIN_SRAM20 Tile_X10Y6_DIN_SRAM21 Tile_X10Y6_DIN_SRAM22
+ Tile_X10Y6_DIN_SRAM23 Tile_X10Y6_DIN_SRAM24 Tile_X10Y6_DIN_SRAM25 Tile_X10Y6_DIN_SRAM26
+ Tile_X10Y6_DIN_SRAM27 Tile_X10Y6_DIN_SRAM28 Tile_X10Y6_DIN_SRAM29 Tile_X10Y6_DIN_SRAM3
+ Tile_X10Y6_DIN_SRAM30 Tile_X10Y6_DIN_SRAM31 Tile_X10Y6_DIN_SRAM4 Tile_X10Y6_DIN_SRAM5
+ Tile_X10Y6_DIN_SRAM6 Tile_X10Y6_DIN_SRAM7 Tile_X10Y6_DIN_SRAM8 Tile_X10Y6_DIN_SRAM9
+ Tile_X10Y6_DOUT_SRAM0 Tile_X10Y6_DOUT_SRAM1 Tile_X10Y6_DOUT_SRAM10 Tile_X10Y6_DOUT_SRAM11
+ Tile_X10Y6_DOUT_SRAM12 Tile_X10Y6_DOUT_SRAM13 Tile_X10Y6_DOUT_SRAM14 Tile_X10Y6_DOUT_SRAM15
+ Tile_X10Y6_DOUT_SRAM16 Tile_X10Y6_DOUT_SRAM17 Tile_X10Y6_DOUT_SRAM18 Tile_X10Y6_DOUT_SRAM19
+ Tile_X10Y6_DOUT_SRAM2 Tile_X10Y6_DOUT_SRAM20 Tile_X10Y6_DOUT_SRAM21 Tile_X10Y6_DOUT_SRAM22
+ Tile_X10Y6_DOUT_SRAM23 Tile_X10Y6_DOUT_SRAM24 Tile_X10Y6_DOUT_SRAM25 Tile_X10Y6_DOUT_SRAM26
+ Tile_X10Y6_DOUT_SRAM27 Tile_X10Y6_DOUT_SRAM28 Tile_X10Y6_DOUT_SRAM29 Tile_X10Y6_DOUT_SRAM3
+ Tile_X10Y6_DOUT_SRAM30 Tile_X10Y6_DOUT_SRAM31 Tile_X10Y6_DOUT_SRAM4 Tile_X10Y6_DOUT_SRAM5
+ Tile_X10Y6_DOUT_SRAM6 Tile_X10Y6_DOUT_SRAM7 Tile_X10Y6_DOUT_SRAM8 Tile_X10Y6_DOUT_SRAM9
+ Tile_X10Y6_MEN_SRAM Tile_X10Y6_REN_SRAM Tile_X10Y6_TIE_HIGH_SRAM Tile_X10Y6_TIE_LOW_SRAM
+ Tile_X10Y6_WEN_SRAM Tile_X10Y8_ADDR_SRAM0 Tile_X10Y8_ADDR_SRAM1 Tile_X10Y8_ADDR_SRAM2
+ Tile_X10Y8_ADDR_SRAM3 Tile_X10Y8_ADDR_SRAM4 Tile_X10Y8_ADDR_SRAM5 Tile_X10Y8_ADDR_SRAM6
+ Tile_X10Y8_ADDR_SRAM7 Tile_X10Y8_ADDR_SRAM8 Tile_X10Y8_ADDR_SRAM9 Tile_X10Y8_BM_SRAM0
+ Tile_X10Y8_BM_SRAM1 Tile_X10Y8_BM_SRAM10 Tile_X10Y8_BM_SRAM11 Tile_X10Y8_BM_SRAM12
+ Tile_X10Y8_BM_SRAM13 Tile_X10Y8_BM_SRAM14 Tile_X10Y8_BM_SRAM15 Tile_X10Y8_BM_SRAM16
+ Tile_X10Y8_BM_SRAM17 Tile_X10Y8_BM_SRAM18 Tile_X10Y8_BM_SRAM19 Tile_X10Y8_BM_SRAM2
+ Tile_X10Y8_BM_SRAM20 Tile_X10Y8_BM_SRAM21 Tile_X10Y8_BM_SRAM22 Tile_X10Y8_BM_SRAM23
+ Tile_X10Y8_BM_SRAM24 Tile_X10Y8_BM_SRAM25 Tile_X10Y8_BM_SRAM26 Tile_X10Y8_BM_SRAM27
+ Tile_X10Y8_BM_SRAM28 Tile_X10Y8_BM_SRAM29 Tile_X10Y8_BM_SRAM3 Tile_X10Y8_BM_SRAM30
+ Tile_X10Y8_BM_SRAM31 Tile_X10Y8_BM_SRAM4 Tile_X10Y8_BM_SRAM5 Tile_X10Y8_BM_SRAM6
+ Tile_X10Y8_BM_SRAM7 Tile_X10Y8_BM_SRAM8 Tile_X10Y8_BM_SRAM9 Tile_X10Y8_CLK_SRAM
+ Tile_X10Y8_CONFIGURED_top Tile_X10Y8_DIN_SRAM0 Tile_X10Y8_DIN_SRAM1 Tile_X10Y8_DIN_SRAM10
+ Tile_X10Y8_DIN_SRAM11 Tile_X10Y8_DIN_SRAM12 Tile_X10Y8_DIN_SRAM13 Tile_X10Y8_DIN_SRAM14
+ Tile_X10Y8_DIN_SRAM15 Tile_X10Y8_DIN_SRAM16 Tile_X10Y8_DIN_SRAM17 Tile_X10Y8_DIN_SRAM18
+ Tile_X10Y8_DIN_SRAM19 Tile_X10Y8_DIN_SRAM2 Tile_X10Y8_DIN_SRAM20 Tile_X10Y8_DIN_SRAM21
+ Tile_X10Y8_DIN_SRAM22 Tile_X10Y8_DIN_SRAM23 Tile_X10Y8_DIN_SRAM24 Tile_X10Y8_DIN_SRAM25
+ Tile_X10Y8_DIN_SRAM26 Tile_X10Y8_DIN_SRAM27 Tile_X10Y8_DIN_SRAM28 Tile_X10Y8_DIN_SRAM29
+ Tile_X10Y8_DIN_SRAM3 Tile_X10Y8_DIN_SRAM30 Tile_X10Y8_DIN_SRAM31 Tile_X10Y8_DIN_SRAM4
+ Tile_X10Y8_DIN_SRAM5 Tile_X10Y8_DIN_SRAM6 Tile_X10Y8_DIN_SRAM7 Tile_X10Y8_DIN_SRAM8
+ Tile_X10Y8_DIN_SRAM9 Tile_X10Y8_DOUT_SRAM0 Tile_X10Y8_DOUT_SRAM1 Tile_X10Y8_DOUT_SRAM10
+ Tile_X10Y8_DOUT_SRAM11 Tile_X10Y8_DOUT_SRAM12 Tile_X10Y8_DOUT_SRAM13 Tile_X10Y8_DOUT_SRAM14
+ Tile_X10Y8_DOUT_SRAM15 Tile_X10Y8_DOUT_SRAM16 Tile_X10Y8_DOUT_SRAM17 Tile_X10Y8_DOUT_SRAM18
+ Tile_X10Y8_DOUT_SRAM19 Tile_X10Y8_DOUT_SRAM2 Tile_X10Y8_DOUT_SRAM20 Tile_X10Y8_DOUT_SRAM21
+ Tile_X10Y8_DOUT_SRAM22 Tile_X10Y8_DOUT_SRAM23 Tile_X10Y8_DOUT_SRAM24 Tile_X10Y8_DOUT_SRAM25
+ Tile_X10Y8_DOUT_SRAM26 Tile_X10Y8_DOUT_SRAM27 Tile_X10Y8_DOUT_SRAM28 Tile_X10Y8_DOUT_SRAM29
+ Tile_X10Y8_DOUT_SRAM3 Tile_X10Y8_DOUT_SRAM30 Tile_X10Y8_DOUT_SRAM31 Tile_X10Y8_DOUT_SRAM4
+ Tile_X10Y8_DOUT_SRAM5 Tile_X10Y8_DOUT_SRAM6 Tile_X10Y8_DOUT_SRAM7 Tile_X10Y8_DOUT_SRAM8
+ Tile_X10Y8_DOUT_SRAM9 Tile_X10Y8_MEN_SRAM Tile_X10Y8_REN_SRAM Tile_X10Y8_TIE_HIGH_SRAM
+ Tile_X10Y8_TIE_LOW_SRAM Tile_X10Y8_WEN_SRAM Tile_X1Y0_A_I_top Tile_X1Y0_A_O_top
+ Tile_X1Y0_A_T_top Tile_X1Y0_A_config_C_bit0 Tile_X1Y0_A_config_C_bit1 Tile_X1Y0_A_config_C_bit2
+ Tile_X1Y0_A_config_C_bit3 Tile_X1Y0_B_I_top Tile_X1Y0_B_O_top Tile_X1Y0_B_T_top
+ Tile_X1Y0_B_config_C_bit0 Tile_X1Y0_B_config_C_bit1 Tile_X1Y0_B_config_C_bit2 Tile_X1Y0_B_config_C_bit3
+ Tile_X2Y0_A_I_top Tile_X2Y0_A_O_top Tile_X2Y0_A_T_top Tile_X2Y0_A_config_C_bit0
+ Tile_X2Y0_A_config_C_bit1 Tile_X2Y0_A_config_C_bit2 Tile_X2Y0_A_config_C_bit3 Tile_X2Y0_B_I_top
+ Tile_X2Y0_B_O_top Tile_X2Y0_B_T_top Tile_X2Y0_B_config_C_bit0 Tile_X2Y0_B_config_C_bit1
+ Tile_X2Y0_B_config_C_bit2 Tile_X2Y0_B_config_C_bit3 Tile_X2Y15_BOOT_top Tile_X2Y15_CONFIGURED_top
+ Tile_X2Y15_RESET_top Tile_X2Y15_SLOT_top0 Tile_X2Y15_SLOT_top1 Tile_X2Y15_SLOT_top2
+ Tile_X2Y15_SLOT_top3 Tile_X3Y15_CONFIGURED_top Tile_X3Y15_IRQ_top0 Tile_X3Y15_IRQ_top1
+ Tile_X3Y15_IRQ_top2 Tile_X3Y15_IRQ_top3 Tile_X5Y15_I_top0 Tile_X5Y15_I_top1 Tile_X5Y15_I_top10
+ Tile_X5Y15_I_top11 Tile_X5Y15_I_top12 Tile_X5Y15_I_top13 Tile_X5Y15_I_top14 Tile_X5Y15_I_top15
+ Tile_X5Y15_I_top2 Tile_X5Y15_I_top3 Tile_X5Y15_I_top4 Tile_X5Y15_I_top5 Tile_X5Y15_I_top6
+ Tile_X5Y15_I_top7 Tile_X5Y15_I_top8 Tile_X5Y15_I_top9 Tile_X5Y15_O_top0 Tile_X5Y15_O_top1
+ Tile_X5Y15_O_top10 Tile_X5Y15_O_top11 Tile_X5Y15_O_top12 Tile_X5Y15_O_top13 Tile_X5Y15_O_top14
+ Tile_X5Y15_O_top15 Tile_X5Y15_O_top2 Tile_X5Y15_O_top3 Tile_X5Y15_O_top4 Tile_X5Y15_O_top5
+ Tile_X5Y15_O_top6 Tile_X5Y15_O_top7 Tile_X5Y15_O_top8 Tile_X5Y15_O_top9 Tile_X6Y15_I_top0
+ Tile_X6Y15_I_top1 Tile_X6Y15_I_top10 Tile_X6Y15_I_top11 Tile_X6Y15_I_top12 Tile_X6Y15_I_top13
+ Tile_X6Y15_I_top14 Tile_X6Y15_I_top15 Tile_X6Y15_I_top2 Tile_X6Y15_I_top3 Tile_X6Y15_I_top4
+ Tile_X6Y15_I_top5 Tile_X6Y15_I_top6 Tile_X6Y15_I_top7 Tile_X6Y15_I_top8 Tile_X6Y15_I_top9
+ Tile_X6Y15_O_top0 Tile_X6Y15_O_top1 Tile_X6Y15_O_top10 Tile_X6Y15_O_top11 Tile_X6Y15_O_top12
+ Tile_X6Y15_O_top13 Tile_X6Y15_O_top14 Tile_X6Y15_O_top15 Tile_X6Y15_O_top2 Tile_X6Y15_O_top3
+ Tile_X6Y15_O_top4 Tile_X6Y15_O_top5 Tile_X6Y15_O_top6 Tile_X6Y15_O_top7 Tile_X6Y15_O_top8
+ Tile_X6Y15_O_top9 Tile_X8Y15_I_top0 Tile_X8Y15_I_top1 Tile_X8Y15_I_top10 Tile_X8Y15_I_top11
+ Tile_X8Y15_I_top12 Tile_X8Y15_I_top13 Tile_X8Y15_I_top14 Tile_X8Y15_I_top15 Tile_X8Y15_I_top2
+ Tile_X8Y15_I_top3 Tile_X8Y15_I_top4 Tile_X8Y15_I_top5 Tile_X8Y15_I_top6 Tile_X8Y15_I_top7
+ Tile_X8Y15_I_top8 Tile_X8Y15_I_top9 Tile_X8Y15_O_top0 Tile_X8Y15_O_top1 Tile_X8Y15_O_top10
+ Tile_X8Y15_O_top11 Tile_X8Y15_O_top12 Tile_X8Y15_O_top13 Tile_X8Y15_O_top14 Tile_X8Y15_O_top15
+ Tile_X8Y15_O_top2 Tile_X8Y15_O_top3 Tile_X8Y15_O_top4 Tile_X8Y15_O_top5 Tile_X8Y15_O_top6
+ Tile_X8Y15_O_top7 Tile_X8Y15_O_top8 Tile_X8Y15_O_top9 Tile_X9Y15_I_top0 Tile_X9Y15_I_top1
+ Tile_X9Y15_I_top10 Tile_X9Y15_I_top11 Tile_X9Y15_I_top12 Tile_X9Y15_I_top13 Tile_X9Y15_I_top14
+ Tile_X9Y15_I_top15 Tile_X9Y15_I_top2 Tile_X9Y15_I_top3 Tile_X9Y15_I_top4 Tile_X9Y15_I_top5
+ Tile_X9Y15_I_top6 Tile_X9Y15_I_top7 Tile_X9Y15_I_top8 Tile_X9Y15_I_top9 Tile_X9Y15_O_top0
+ Tile_X9Y15_O_top1 Tile_X9Y15_O_top10 Tile_X9Y15_O_top11 Tile_X9Y15_O_top12 Tile_X9Y15_O_top13
+ Tile_X9Y15_O_top14 Tile_X9Y15_O_top15 Tile_X9Y15_O_top2 Tile_X9Y15_O_top3 Tile_X9Y15_O_top4
+ Tile_X9Y15_O_top5 Tile_X9Y15_O_top6 Tile_X9Y15_O_top7 Tile_X9Y15_O_top8 Tile_X9Y15_O_top9
+ UserCLK VGND VPWR
XTile_X1Y0_N_IO Tile_X1Y0_A_I_top Tile_X1Y0_A_O_top Tile_X1Y0_A_T_top Tile_X1Y0_A_config_C_bit0
+ Tile_X1Y0_A_config_C_bit1 Tile_X1Y0_A_config_C_bit2 Tile_X1Y0_A_config_C_bit3 Tile_X1Y0_B_I_top
+ Tile_X1Y0_B_O_top Tile_X1Y0_B_T_top Tile_X1Y0_B_config_C_bit0 Tile_X1Y0_B_config_C_bit1
+ Tile_X1Y0_B_config_C_bit2 Tile_X1Y0_B_config_C_bit3 Tile_X1Y0_N_IO/Ci FrameData[0]
+ FrameData[10] FrameData[11] FrameData[12] FrameData[13] FrameData[14] FrameData[15]
+ FrameData[16] FrameData[17] FrameData[18] FrameData[19] FrameData[1] FrameData[20]
+ FrameData[21] FrameData[22] FrameData[23] FrameData[24] FrameData[25] FrameData[26]
+ FrameData[27] FrameData[28] FrameData[29] FrameData[2] FrameData[30] FrameData[31]
+ FrameData[3] FrameData[4] FrameData[5] FrameData[6] FrameData[7] FrameData[8] FrameData[9]
+ Tile_X2Y0_N_IO/FrameData[0] Tile_X2Y0_N_IO/FrameData[10] Tile_X2Y0_N_IO/FrameData[11]
+ Tile_X2Y0_N_IO/FrameData[12] Tile_X2Y0_N_IO/FrameData[13] Tile_X2Y0_N_IO/FrameData[14]
+ Tile_X2Y0_N_IO/FrameData[15] Tile_X2Y0_N_IO/FrameData[16] Tile_X2Y0_N_IO/FrameData[17]
+ Tile_X2Y0_N_IO/FrameData[18] Tile_X2Y0_N_IO/FrameData[19] Tile_X2Y0_N_IO/FrameData[1]
+ Tile_X2Y0_N_IO/FrameData[20] Tile_X2Y0_N_IO/FrameData[21] Tile_X2Y0_N_IO/FrameData[22]
+ Tile_X2Y0_N_IO/FrameData[23] Tile_X2Y0_N_IO/FrameData[24] Tile_X2Y0_N_IO/FrameData[25]
+ Tile_X2Y0_N_IO/FrameData[26] Tile_X2Y0_N_IO/FrameData[27] Tile_X2Y0_N_IO/FrameData[28]
+ Tile_X2Y0_N_IO/FrameData[29] Tile_X2Y0_N_IO/FrameData[2] Tile_X2Y0_N_IO/FrameData[30]
+ Tile_X2Y0_N_IO/FrameData[31] Tile_X2Y0_N_IO/FrameData[3] Tile_X2Y0_N_IO/FrameData[4]
+ Tile_X2Y0_N_IO/FrameData[5] Tile_X2Y0_N_IO/FrameData[6] Tile_X2Y0_N_IO/FrameData[7]
+ Tile_X2Y0_N_IO/FrameData[8] Tile_X2Y0_N_IO/FrameData[9] Tile_X1Y0_N_IO/FrameStrobe[0]
+ Tile_X1Y0_N_IO/FrameStrobe[10] Tile_X1Y0_N_IO/FrameStrobe[11] Tile_X1Y0_N_IO/FrameStrobe[12]
+ Tile_X1Y0_N_IO/FrameStrobe[13] Tile_X1Y0_N_IO/FrameStrobe[14] Tile_X1Y0_N_IO/FrameStrobe[15]
+ Tile_X1Y0_N_IO/FrameStrobe[16] Tile_X1Y0_N_IO/FrameStrobe[17] Tile_X1Y0_N_IO/FrameStrobe[18]
+ Tile_X1Y0_N_IO/FrameStrobe[19] Tile_X1Y0_N_IO/FrameStrobe[1] Tile_X1Y0_N_IO/FrameStrobe[2]
+ Tile_X1Y0_N_IO/FrameStrobe[3] Tile_X1Y0_N_IO/FrameStrobe[4] Tile_X1Y0_N_IO/FrameStrobe[5]
+ Tile_X1Y0_N_IO/FrameStrobe[6] Tile_X1Y0_N_IO/FrameStrobe[7] Tile_X1Y0_N_IO/FrameStrobe[8]
+ Tile_X1Y0_N_IO/FrameStrobe[9] Tile_X1Y0_N_IO/FrameStrobe_O[0] Tile_X1Y0_N_IO/FrameStrobe_O[10]
+ Tile_X1Y0_N_IO/FrameStrobe_O[11] Tile_X1Y0_N_IO/FrameStrobe_O[12] Tile_X1Y0_N_IO/FrameStrobe_O[13]
+ Tile_X1Y0_N_IO/FrameStrobe_O[14] Tile_X1Y0_N_IO/FrameStrobe_O[15] Tile_X1Y0_N_IO/FrameStrobe_O[16]
+ Tile_X1Y0_N_IO/FrameStrobe_O[17] Tile_X1Y0_N_IO/FrameStrobe_O[18] Tile_X1Y0_N_IO/FrameStrobe_O[19]
+ Tile_X1Y0_N_IO/FrameStrobe_O[1] Tile_X1Y0_N_IO/FrameStrobe_O[2] Tile_X1Y0_N_IO/FrameStrobe_O[3]
+ Tile_X1Y0_N_IO/FrameStrobe_O[4] Tile_X1Y0_N_IO/FrameStrobe_O[5] Tile_X1Y0_N_IO/FrameStrobe_O[6]
+ Tile_X1Y0_N_IO/FrameStrobe_O[7] Tile_X1Y0_N_IO/FrameStrobe_O[8] Tile_X1Y0_N_IO/FrameStrobe_O[9]
+ Tile_X1Y0_N_IO/N1END[0] Tile_X1Y0_N_IO/N1END[1] Tile_X1Y0_N_IO/N1END[2] Tile_X1Y0_N_IO/N1END[3]
+ Tile_X1Y0_N_IO/N2END[0] Tile_X1Y0_N_IO/N2END[1] Tile_X1Y0_N_IO/N2END[2] Tile_X1Y0_N_IO/N2END[3]
+ Tile_X1Y0_N_IO/N2END[4] Tile_X1Y0_N_IO/N2END[5] Tile_X1Y0_N_IO/N2END[6] Tile_X1Y0_N_IO/N2END[7]
+ Tile_X1Y0_N_IO/N2MID[0] Tile_X1Y0_N_IO/N2MID[1] Tile_X1Y0_N_IO/N2MID[2] Tile_X1Y0_N_IO/N2MID[3]
+ Tile_X1Y0_N_IO/N2MID[4] Tile_X1Y0_N_IO/N2MID[5] Tile_X1Y0_N_IO/N2MID[6] Tile_X1Y0_N_IO/N2MID[7]
+ Tile_X1Y0_N_IO/N4END[0] Tile_X1Y0_N_IO/N4END[10] Tile_X1Y0_N_IO/N4END[11] Tile_X1Y0_N_IO/N4END[12]
+ Tile_X1Y0_N_IO/N4END[13] Tile_X1Y0_N_IO/N4END[14] Tile_X1Y0_N_IO/N4END[15] Tile_X1Y0_N_IO/N4END[1]
+ Tile_X1Y0_N_IO/N4END[2] Tile_X1Y0_N_IO/N4END[3] Tile_X1Y0_N_IO/N4END[4] Tile_X1Y0_N_IO/N4END[5]
+ Tile_X1Y0_N_IO/N4END[6] Tile_X1Y0_N_IO/N4END[7] Tile_X1Y0_N_IO/N4END[8] Tile_X1Y0_N_IO/N4END[9]
+ Tile_X1Y0_N_IO/NN4END[0] Tile_X1Y0_N_IO/NN4END[10] Tile_X1Y0_N_IO/NN4END[11] Tile_X1Y0_N_IO/NN4END[12]
+ Tile_X1Y0_N_IO/NN4END[13] Tile_X1Y0_N_IO/NN4END[14] Tile_X1Y0_N_IO/NN4END[15] Tile_X1Y0_N_IO/NN4END[1]
+ Tile_X1Y0_N_IO/NN4END[2] Tile_X1Y0_N_IO/NN4END[3] Tile_X1Y0_N_IO/NN4END[4] Tile_X1Y0_N_IO/NN4END[5]
+ Tile_X1Y0_N_IO/NN4END[6] Tile_X1Y0_N_IO/NN4END[7] Tile_X1Y0_N_IO/NN4END[8] Tile_X1Y0_N_IO/NN4END[9]
+ Tile_X1Y0_N_IO/S1BEG[0] Tile_X1Y0_N_IO/S1BEG[1] Tile_X1Y0_N_IO/S1BEG[2] Tile_X1Y0_N_IO/S1BEG[3]
+ Tile_X1Y0_N_IO/S2BEG[0] Tile_X1Y0_N_IO/S2BEG[1] Tile_X1Y0_N_IO/S2BEG[2] Tile_X1Y0_N_IO/S2BEG[3]
+ Tile_X1Y0_N_IO/S2BEG[4] Tile_X1Y0_N_IO/S2BEG[5] Tile_X1Y0_N_IO/S2BEG[6] Tile_X1Y0_N_IO/S2BEG[7]
+ Tile_X1Y0_N_IO/S2BEGb[0] Tile_X1Y0_N_IO/S2BEGb[1] Tile_X1Y0_N_IO/S2BEGb[2] Tile_X1Y0_N_IO/S2BEGb[3]
+ Tile_X1Y0_N_IO/S2BEGb[4] Tile_X1Y0_N_IO/S2BEGb[5] Tile_X1Y0_N_IO/S2BEGb[6] Tile_X1Y0_N_IO/S2BEGb[7]
+ Tile_X1Y0_N_IO/S4BEG[0] Tile_X1Y0_N_IO/S4BEG[10] Tile_X1Y0_N_IO/S4BEG[11] Tile_X1Y0_N_IO/S4BEG[12]
+ Tile_X1Y0_N_IO/S4BEG[13] Tile_X1Y0_N_IO/S4BEG[14] Tile_X1Y0_N_IO/S4BEG[15] Tile_X1Y0_N_IO/S4BEG[1]
+ Tile_X1Y0_N_IO/S4BEG[2] Tile_X1Y0_N_IO/S4BEG[3] Tile_X1Y0_N_IO/S4BEG[4] Tile_X1Y0_N_IO/S4BEG[5]
+ Tile_X1Y0_N_IO/S4BEG[6] Tile_X1Y0_N_IO/S4BEG[7] Tile_X1Y0_N_IO/S4BEG[8] Tile_X1Y0_N_IO/S4BEG[9]
+ Tile_X1Y0_N_IO/SS4BEG[0] Tile_X1Y0_N_IO/SS4BEG[10] Tile_X1Y0_N_IO/SS4BEG[11] Tile_X1Y0_N_IO/SS4BEG[12]
+ Tile_X1Y0_N_IO/SS4BEG[13] Tile_X1Y0_N_IO/SS4BEG[14] Tile_X1Y0_N_IO/SS4BEG[15] Tile_X1Y0_N_IO/SS4BEG[1]
+ Tile_X1Y0_N_IO/SS4BEG[2] Tile_X1Y0_N_IO/SS4BEG[3] Tile_X1Y0_N_IO/SS4BEG[4] Tile_X1Y0_N_IO/SS4BEG[5]
+ Tile_X1Y0_N_IO/SS4BEG[6] Tile_X1Y0_N_IO/SS4BEG[7] Tile_X1Y0_N_IO/SS4BEG[8] Tile_X1Y0_N_IO/SS4BEG[9]
+ Tile_X1Y0_N_IO/UserCLK Tile_X1Y0_N_IO/UserCLKo VGND VPWR N_IO
XTile_X3Y3_LUT4AB Tile_X3Y4_LUT4AB/Co Tile_X3Y3_LUT4AB/Co Tile_X3Y3_LUT4AB/E1BEG[0]
+ Tile_X3Y3_LUT4AB/E1BEG[1] Tile_X3Y3_LUT4AB/E1BEG[2] Tile_X3Y3_LUT4AB/E1BEG[3] Tile_X3Y3_LUT4AB/E1END[0]
+ Tile_X3Y3_LUT4AB/E1END[1] Tile_X3Y3_LUT4AB/E1END[2] Tile_X3Y3_LUT4AB/E1END[3] Tile_X3Y3_LUT4AB/E2BEG[0]
+ Tile_X3Y3_LUT4AB/E2BEG[1] Tile_X3Y3_LUT4AB/E2BEG[2] Tile_X3Y3_LUT4AB/E2BEG[3] Tile_X3Y3_LUT4AB/E2BEG[4]
+ Tile_X3Y3_LUT4AB/E2BEG[5] Tile_X3Y3_LUT4AB/E2BEG[6] Tile_X3Y3_LUT4AB/E2BEG[7] Tile_X4Y3_RegFile/E2END[0]
+ Tile_X4Y3_RegFile/E2END[1] Tile_X4Y3_RegFile/E2END[2] Tile_X4Y3_RegFile/E2END[3]
+ Tile_X4Y3_RegFile/E2END[4] Tile_X4Y3_RegFile/E2END[5] Tile_X4Y3_RegFile/E2END[6]
+ Tile_X4Y3_RegFile/E2END[7] Tile_X3Y3_LUT4AB/E2END[0] Tile_X3Y3_LUT4AB/E2END[1] Tile_X3Y3_LUT4AB/E2END[2]
+ Tile_X3Y3_LUT4AB/E2END[3] Tile_X3Y3_LUT4AB/E2END[4] Tile_X3Y3_LUT4AB/E2END[5] Tile_X3Y3_LUT4AB/E2END[6]
+ Tile_X3Y3_LUT4AB/E2END[7] Tile_X3Y3_LUT4AB/E2MID[0] Tile_X3Y3_LUT4AB/E2MID[1] Tile_X3Y3_LUT4AB/E2MID[2]
+ Tile_X3Y3_LUT4AB/E2MID[3] Tile_X3Y3_LUT4AB/E2MID[4] Tile_X3Y3_LUT4AB/E2MID[5] Tile_X3Y3_LUT4AB/E2MID[6]
+ Tile_X3Y3_LUT4AB/E2MID[7] Tile_X3Y3_LUT4AB/E6BEG[0] Tile_X3Y3_LUT4AB/E6BEG[10] Tile_X3Y3_LUT4AB/E6BEG[11]
+ Tile_X3Y3_LUT4AB/E6BEG[1] Tile_X3Y3_LUT4AB/E6BEG[2] Tile_X3Y3_LUT4AB/E6BEG[3] Tile_X3Y3_LUT4AB/E6BEG[4]
+ Tile_X3Y3_LUT4AB/E6BEG[5] Tile_X3Y3_LUT4AB/E6BEG[6] Tile_X3Y3_LUT4AB/E6BEG[7] Tile_X3Y3_LUT4AB/E6BEG[8]
+ Tile_X3Y3_LUT4AB/E6BEG[9] Tile_X3Y3_LUT4AB/E6END[0] Tile_X3Y3_LUT4AB/E6END[10] Tile_X3Y3_LUT4AB/E6END[11]
+ Tile_X3Y3_LUT4AB/E6END[1] Tile_X3Y3_LUT4AB/E6END[2] Tile_X3Y3_LUT4AB/E6END[3] Tile_X3Y3_LUT4AB/E6END[4]
+ Tile_X3Y3_LUT4AB/E6END[5] Tile_X3Y3_LUT4AB/E6END[6] Tile_X3Y3_LUT4AB/E6END[7] Tile_X3Y3_LUT4AB/E6END[8]
+ Tile_X3Y3_LUT4AB/E6END[9] Tile_X3Y3_LUT4AB/EE4BEG[0] Tile_X3Y3_LUT4AB/EE4BEG[10]
+ Tile_X3Y3_LUT4AB/EE4BEG[11] Tile_X3Y3_LUT4AB/EE4BEG[12] Tile_X3Y3_LUT4AB/EE4BEG[13]
+ Tile_X3Y3_LUT4AB/EE4BEG[14] Tile_X3Y3_LUT4AB/EE4BEG[15] Tile_X3Y3_LUT4AB/EE4BEG[1]
+ Tile_X3Y3_LUT4AB/EE4BEG[2] Tile_X3Y3_LUT4AB/EE4BEG[3] Tile_X3Y3_LUT4AB/EE4BEG[4]
+ Tile_X3Y3_LUT4AB/EE4BEG[5] Tile_X3Y3_LUT4AB/EE4BEG[6] Tile_X3Y3_LUT4AB/EE4BEG[7]
+ Tile_X3Y3_LUT4AB/EE4BEG[8] Tile_X3Y3_LUT4AB/EE4BEG[9] Tile_X3Y3_LUT4AB/EE4END[0]
+ Tile_X3Y3_LUT4AB/EE4END[10] Tile_X3Y3_LUT4AB/EE4END[11] Tile_X3Y3_LUT4AB/EE4END[12]
+ Tile_X3Y3_LUT4AB/EE4END[13] Tile_X3Y3_LUT4AB/EE4END[14] Tile_X3Y3_LUT4AB/EE4END[15]
+ Tile_X3Y3_LUT4AB/EE4END[1] Tile_X3Y3_LUT4AB/EE4END[2] Tile_X3Y3_LUT4AB/EE4END[3]
+ Tile_X3Y3_LUT4AB/EE4END[4] Tile_X3Y3_LUT4AB/EE4END[5] Tile_X3Y3_LUT4AB/EE4END[6]
+ Tile_X3Y3_LUT4AB/EE4END[7] Tile_X3Y3_LUT4AB/EE4END[8] Tile_X3Y3_LUT4AB/EE4END[9]
+ Tile_X3Y3_LUT4AB/FrameData[0] Tile_X3Y3_LUT4AB/FrameData[10] Tile_X3Y3_LUT4AB/FrameData[11]
+ Tile_X3Y3_LUT4AB/FrameData[12] Tile_X3Y3_LUT4AB/FrameData[13] Tile_X3Y3_LUT4AB/FrameData[14]
+ Tile_X3Y3_LUT4AB/FrameData[15] Tile_X3Y3_LUT4AB/FrameData[16] Tile_X3Y3_LUT4AB/FrameData[17]
+ Tile_X3Y3_LUT4AB/FrameData[18] Tile_X3Y3_LUT4AB/FrameData[19] Tile_X3Y3_LUT4AB/FrameData[1]
+ Tile_X3Y3_LUT4AB/FrameData[20] Tile_X3Y3_LUT4AB/FrameData[21] Tile_X3Y3_LUT4AB/FrameData[22]
+ Tile_X3Y3_LUT4AB/FrameData[23] Tile_X3Y3_LUT4AB/FrameData[24] Tile_X3Y3_LUT4AB/FrameData[25]
+ Tile_X3Y3_LUT4AB/FrameData[26] Tile_X3Y3_LUT4AB/FrameData[27] Tile_X3Y3_LUT4AB/FrameData[28]
+ Tile_X3Y3_LUT4AB/FrameData[29] Tile_X3Y3_LUT4AB/FrameData[2] Tile_X3Y3_LUT4AB/FrameData[30]
+ Tile_X3Y3_LUT4AB/FrameData[31] Tile_X3Y3_LUT4AB/FrameData[3] Tile_X3Y3_LUT4AB/FrameData[4]
+ Tile_X3Y3_LUT4AB/FrameData[5] Tile_X3Y3_LUT4AB/FrameData[6] Tile_X3Y3_LUT4AB/FrameData[7]
+ Tile_X3Y3_LUT4AB/FrameData[8] Tile_X3Y3_LUT4AB/FrameData[9] Tile_X4Y3_RegFile/FrameData[0]
+ Tile_X4Y3_RegFile/FrameData[10] Tile_X4Y3_RegFile/FrameData[11] Tile_X4Y3_RegFile/FrameData[12]
+ Tile_X4Y3_RegFile/FrameData[13] Tile_X4Y3_RegFile/FrameData[14] Tile_X4Y3_RegFile/FrameData[15]
+ Tile_X4Y3_RegFile/FrameData[16] Tile_X4Y3_RegFile/FrameData[17] Tile_X4Y3_RegFile/FrameData[18]
+ Tile_X4Y3_RegFile/FrameData[19] Tile_X4Y3_RegFile/FrameData[1] Tile_X4Y3_RegFile/FrameData[20]
+ Tile_X4Y3_RegFile/FrameData[21] Tile_X4Y3_RegFile/FrameData[22] Tile_X4Y3_RegFile/FrameData[23]
+ Tile_X4Y3_RegFile/FrameData[24] Tile_X4Y3_RegFile/FrameData[25] Tile_X4Y3_RegFile/FrameData[26]
+ Tile_X4Y3_RegFile/FrameData[27] Tile_X4Y3_RegFile/FrameData[28] Tile_X4Y3_RegFile/FrameData[29]
+ Tile_X4Y3_RegFile/FrameData[2] Tile_X4Y3_RegFile/FrameData[30] Tile_X4Y3_RegFile/FrameData[31]
+ Tile_X4Y3_RegFile/FrameData[3] Tile_X4Y3_RegFile/FrameData[4] Tile_X4Y3_RegFile/FrameData[5]
+ Tile_X4Y3_RegFile/FrameData[6] Tile_X4Y3_RegFile/FrameData[7] Tile_X4Y3_RegFile/FrameData[8]
+ Tile_X4Y3_RegFile/FrameData[9] Tile_X3Y3_LUT4AB/FrameStrobe[0] Tile_X3Y3_LUT4AB/FrameStrobe[10]
+ Tile_X3Y3_LUT4AB/FrameStrobe[11] Tile_X3Y3_LUT4AB/FrameStrobe[12] Tile_X3Y3_LUT4AB/FrameStrobe[13]
+ Tile_X3Y3_LUT4AB/FrameStrobe[14] Tile_X3Y3_LUT4AB/FrameStrobe[15] Tile_X3Y3_LUT4AB/FrameStrobe[16]
+ Tile_X3Y3_LUT4AB/FrameStrobe[17] Tile_X3Y3_LUT4AB/FrameStrobe[18] Tile_X3Y3_LUT4AB/FrameStrobe[19]
+ Tile_X3Y3_LUT4AB/FrameStrobe[1] Tile_X3Y3_LUT4AB/FrameStrobe[2] Tile_X3Y3_LUT4AB/FrameStrobe[3]
+ Tile_X3Y3_LUT4AB/FrameStrobe[4] Tile_X3Y3_LUT4AB/FrameStrobe[5] Tile_X3Y3_LUT4AB/FrameStrobe[6]
+ Tile_X3Y3_LUT4AB/FrameStrobe[7] Tile_X3Y3_LUT4AB/FrameStrobe[8] Tile_X3Y3_LUT4AB/FrameStrobe[9]
+ Tile_X3Y2_LUT4AB/FrameStrobe[0] Tile_X3Y2_LUT4AB/FrameStrobe[10] Tile_X3Y2_LUT4AB/FrameStrobe[11]
+ Tile_X3Y2_LUT4AB/FrameStrobe[12] Tile_X3Y2_LUT4AB/FrameStrobe[13] Tile_X3Y2_LUT4AB/FrameStrobe[14]
+ Tile_X3Y2_LUT4AB/FrameStrobe[15] Tile_X3Y2_LUT4AB/FrameStrobe[16] Tile_X3Y2_LUT4AB/FrameStrobe[17]
+ Tile_X3Y2_LUT4AB/FrameStrobe[18] Tile_X3Y2_LUT4AB/FrameStrobe[19] Tile_X3Y2_LUT4AB/FrameStrobe[1]
+ Tile_X3Y2_LUT4AB/FrameStrobe[2] Tile_X3Y2_LUT4AB/FrameStrobe[3] Tile_X3Y2_LUT4AB/FrameStrobe[4]
+ Tile_X3Y2_LUT4AB/FrameStrobe[5] Tile_X3Y2_LUT4AB/FrameStrobe[6] Tile_X3Y2_LUT4AB/FrameStrobe[7]
+ Tile_X3Y2_LUT4AB/FrameStrobe[8] Tile_X3Y2_LUT4AB/FrameStrobe[9] Tile_X3Y3_LUT4AB/N1BEG[0]
+ Tile_X3Y3_LUT4AB/N1BEG[1] Tile_X3Y3_LUT4AB/N1BEG[2] Tile_X3Y3_LUT4AB/N1BEG[3] Tile_X3Y4_LUT4AB/N1BEG[0]
+ Tile_X3Y4_LUT4AB/N1BEG[1] Tile_X3Y4_LUT4AB/N1BEG[2] Tile_X3Y4_LUT4AB/N1BEG[3] Tile_X3Y3_LUT4AB/N2BEG[0]
+ Tile_X3Y3_LUT4AB/N2BEG[1] Tile_X3Y3_LUT4AB/N2BEG[2] Tile_X3Y3_LUT4AB/N2BEG[3] Tile_X3Y3_LUT4AB/N2BEG[4]
+ Tile_X3Y3_LUT4AB/N2BEG[5] Tile_X3Y3_LUT4AB/N2BEG[6] Tile_X3Y3_LUT4AB/N2BEG[7] Tile_X3Y2_LUT4AB/N2END[0]
+ Tile_X3Y2_LUT4AB/N2END[1] Tile_X3Y2_LUT4AB/N2END[2] Tile_X3Y2_LUT4AB/N2END[3] Tile_X3Y2_LUT4AB/N2END[4]
+ Tile_X3Y2_LUT4AB/N2END[5] Tile_X3Y2_LUT4AB/N2END[6] Tile_X3Y2_LUT4AB/N2END[7] Tile_X3Y3_LUT4AB/N2END[0]
+ Tile_X3Y3_LUT4AB/N2END[1] Tile_X3Y3_LUT4AB/N2END[2] Tile_X3Y3_LUT4AB/N2END[3] Tile_X3Y3_LUT4AB/N2END[4]
+ Tile_X3Y3_LUT4AB/N2END[5] Tile_X3Y3_LUT4AB/N2END[6] Tile_X3Y3_LUT4AB/N2END[7] Tile_X3Y4_LUT4AB/N2BEG[0]
+ Tile_X3Y4_LUT4AB/N2BEG[1] Tile_X3Y4_LUT4AB/N2BEG[2] Tile_X3Y4_LUT4AB/N2BEG[3] Tile_X3Y4_LUT4AB/N2BEG[4]
+ Tile_X3Y4_LUT4AB/N2BEG[5] Tile_X3Y4_LUT4AB/N2BEG[6] Tile_X3Y4_LUT4AB/N2BEG[7] Tile_X3Y3_LUT4AB/N4BEG[0]
+ Tile_X3Y3_LUT4AB/N4BEG[10] Tile_X3Y3_LUT4AB/N4BEG[11] Tile_X3Y3_LUT4AB/N4BEG[12]
+ Tile_X3Y3_LUT4AB/N4BEG[13] Tile_X3Y3_LUT4AB/N4BEG[14] Tile_X3Y3_LUT4AB/N4BEG[15]
+ Tile_X3Y3_LUT4AB/N4BEG[1] Tile_X3Y3_LUT4AB/N4BEG[2] Tile_X3Y3_LUT4AB/N4BEG[3] Tile_X3Y3_LUT4AB/N4BEG[4]
+ Tile_X3Y3_LUT4AB/N4BEG[5] Tile_X3Y3_LUT4AB/N4BEG[6] Tile_X3Y3_LUT4AB/N4BEG[7] Tile_X3Y3_LUT4AB/N4BEG[8]
+ Tile_X3Y3_LUT4AB/N4BEG[9] Tile_X3Y4_LUT4AB/N4BEG[0] Tile_X3Y4_LUT4AB/N4BEG[10] Tile_X3Y4_LUT4AB/N4BEG[11]
+ Tile_X3Y4_LUT4AB/N4BEG[12] Tile_X3Y4_LUT4AB/N4BEG[13] Tile_X3Y4_LUT4AB/N4BEG[14]
+ Tile_X3Y4_LUT4AB/N4BEG[15] Tile_X3Y4_LUT4AB/N4BEG[1] Tile_X3Y4_LUT4AB/N4BEG[2] Tile_X3Y4_LUT4AB/N4BEG[3]
+ Tile_X3Y4_LUT4AB/N4BEG[4] Tile_X3Y4_LUT4AB/N4BEG[5] Tile_X3Y4_LUT4AB/N4BEG[6] Tile_X3Y4_LUT4AB/N4BEG[7]
+ Tile_X3Y4_LUT4AB/N4BEG[8] Tile_X3Y4_LUT4AB/N4BEG[9] Tile_X3Y3_LUT4AB/NN4BEG[0] Tile_X3Y3_LUT4AB/NN4BEG[10]
+ Tile_X3Y3_LUT4AB/NN4BEG[11] Tile_X3Y3_LUT4AB/NN4BEG[12] Tile_X3Y3_LUT4AB/NN4BEG[13]
+ Tile_X3Y3_LUT4AB/NN4BEG[14] Tile_X3Y3_LUT4AB/NN4BEG[15] Tile_X3Y3_LUT4AB/NN4BEG[1]
+ Tile_X3Y3_LUT4AB/NN4BEG[2] Tile_X3Y3_LUT4AB/NN4BEG[3] Tile_X3Y3_LUT4AB/NN4BEG[4]
+ Tile_X3Y3_LUT4AB/NN4BEG[5] Tile_X3Y3_LUT4AB/NN4BEG[6] Tile_X3Y3_LUT4AB/NN4BEG[7]
+ Tile_X3Y3_LUT4AB/NN4BEG[8] Tile_X3Y3_LUT4AB/NN4BEG[9] Tile_X3Y4_LUT4AB/NN4BEG[0]
+ Tile_X3Y4_LUT4AB/NN4BEG[10] Tile_X3Y4_LUT4AB/NN4BEG[11] Tile_X3Y4_LUT4AB/NN4BEG[12]
+ Tile_X3Y4_LUT4AB/NN4BEG[13] Tile_X3Y4_LUT4AB/NN4BEG[14] Tile_X3Y4_LUT4AB/NN4BEG[15]
+ Tile_X3Y4_LUT4AB/NN4BEG[1] Tile_X3Y4_LUT4AB/NN4BEG[2] Tile_X3Y4_LUT4AB/NN4BEG[3]
+ Tile_X3Y4_LUT4AB/NN4BEG[4] Tile_X3Y4_LUT4AB/NN4BEG[5] Tile_X3Y4_LUT4AB/NN4BEG[6]
+ Tile_X3Y4_LUT4AB/NN4BEG[7] Tile_X3Y4_LUT4AB/NN4BEG[8] Tile_X3Y4_LUT4AB/NN4BEG[9]
+ Tile_X3Y4_LUT4AB/S1END[0] Tile_X3Y4_LUT4AB/S1END[1] Tile_X3Y4_LUT4AB/S1END[2] Tile_X3Y4_LUT4AB/S1END[3]
+ Tile_X3Y3_LUT4AB/S1END[0] Tile_X3Y3_LUT4AB/S1END[1] Tile_X3Y3_LUT4AB/S1END[2] Tile_X3Y3_LUT4AB/S1END[3]
+ Tile_X3Y4_LUT4AB/S2MID[0] Tile_X3Y4_LUT4AB/S2MID[1] Tile_X3Y4_LUT4AB/S2MID[2] Tile_X3Y4_LUT4AB/S2MID[3]
+ Tile_X3Y4_LUT4AB/S2MID[4] Tile_X3Y4_LUT4AB/S2MID[5] Tile_X3Y4_LUT4AB/S2MID[6] Tile_X3Y4_LUT4AB/S2MID[7]
+ Tile_X3Y4_LUT4AB/S2END[0] Tile_X3Y4_LUT4AB/S2END[1] Tile_X3Y4_LUT4AB/S2END[2] Tile_X3Y4_LUT4AB/S2END[3]
+ Tile_X3Y4_LUT4AB/S2END[4] Tile_X3Y4_LUT4AB/S2END[5] Tile_X3Y4_LUT4AB/S2END[6] Tile_X3Y4_LUT4AB/S2END[7]
+ Tile_X3Y3_LUT4AB/S2END[0] Tile_X3Y3_LUT4AB/S2END[1] Tile_X3Y3_LUT4AB/S2END[2] Tile_X3Y3_LUT4AB/S2END[3]
+ Tile_X3Y3_LUT4AB/S2END[4] Tile_X3Y3_LUT4AB/S2END[5] Tile_X3Y3_LUT4AB/S2END[6] Tile_X3Y3_LUT4AB/S2END[7]
+ Tile_X3Y3_LUT4AB/S2MID[0] Tile_X3Y3_LUT4AB/S2MID[1] Tile_X3Y3_LUT4AB/S2MID[2] Tile_X3Y3_LUT4AB/S2MID[3]
+ Tile_X3Y3_LUT4AB/S2MID[4] Tile_X3Y3_LUT4AB/S2MID[5] Tile_X3Y3_LUT4AB/S2MID[6] Tile_X3Y3_LUT4AB/S2MID[7]
+ Tile_X3Y4_LUT4AB/S4END[0] Tile_X3Y4_LUT4AB/S4END[10] Tile_X3Y4_LUT4AB/S4END[11]
+ Tile_X3Y4_LUT4AB/S4END[12] Tile_X3Y4_LUT4AB/S4END[13] Tile_X3Y4_LUT4AB/S4END[14]
+ Tile_X3Y4_LUT4AB/S4END[15] Tile_X3Y4_LUT4AB/S4END[1] Tile_X3Y4_LUT4AB/S4END[2] Tile_X3Y4_LUT4AB/S4END[3]
+ Tile_X3Y4_LUT4AB/S4END[4] Tile_X3Y4_LUT4AB/S4END[5] Tile_X3Y4_LUT4AB/S4END[6] Tile_X3Y4_LUT4AB/S4END[7]
+ Tile_X3Y4_LUT4AB/S4END[8] Tile_X3Y4_LUT4AB/S4END[9] Tile_X3Y3_LUT4AB/S4END[0] Tile_X3Y3_LUT4AB/S4END[10]
+ Tile_X3Y3_LUT4AB/S4END[11] Tile_X3Y3_LUT4AB/S4END[12] Tile_X3Y3_LUT4AB/S4END[13]
+ Tile_X3Y3_LUT4AB/S4END[14] Tile_X3Y3_LUT4AB/S4END[15] Tile_X3Y3_LUT4AB/S4END[1]
+ Tile_X3Y3_LUT4AB/S4END[2] Tile_X3Y3_LUT4AB/S4END[3] Tile_X3Y3_LUT4AB/S4END[4] Tile_X3Y3_LUT4AB/S4END[5]
+ Tile_X3Y3_LUT4AB/S4END[6] Tile_X3Y3_LUT4AB/S4END[7] Tile_X3Y3_LUT4AB/S4END[8] Tile_X3Y3_LUT4AB/S4END[9]
+ Tile_X3Y4_LUT4AB/SS4END[0] Tile_X3Y4_LUT4AB/SS4END[10] Tile_X3Y4_LUT4AB/SS4END[11]
+ Tile_X3Y4_LUT4AB/SS4END[12] Tile_X3Y4_LUT4AB/SS4END[13] Tile_X3Y4_LUT4AB/SS4END[14]
+ Tile_X3Y4_LUT4AB/SS4END[15] Tile_X3Y4_LUT4AB/SS4END[1] Tile_X3Y4_LUT4AB/SS4END[2]
+ Tile_X3Y4_LUT4AB/SS4END[3] Tile_X3Y4_LUT4AB/SS4END[4] Tile_X3Y4_LUT4AB/SS4END[5]
+ Tile_X3Y4_LUT4AB/SS4END[6] Tile_X3Y4_LUT4AB/SS4END[7] Tile_X3Y4_LUT4AB/SS4END[8]
+ Tile_X3Y4_LUT4AB/SS4END[9] Tile_X3Y3_LUT4AB/SS4END[0] Tile_X3Y3_LUT4AB/SS4END[10]
+ Tile_X3Y3_LUT4AB/SS4END[11] Tile_X3Y3_LUT4AB/SS4END[12] Tile_X3Y3_LUT4AB/SS4END[13]
+ Tile_X3Y3_LUT4AB/SS4END[14] Tile_X3Y3_LUT4AB/SS4END[15] Tile_X3Y3_LUT4AB/SS4END[1]
+ Tile_X3Y3_LUT4AB/SS4END[2] Tile_X3Y3_LUT4AB/SS4END[3] Tile_X3Y3_LUT4AB/SS4END[4]
+ Tile_X3Y3_LUT4AB/SS4END[5] Tile_X3Y3_LUT4AB/SS4END[6] Tile_X3Y3_LUT4AB/SS4END[7]
+ Tile_X3Y3_LUT4AB/SS4END[8] Tile_X3Y3_LUT4AB/SS4END[9] Tile_X3Y3_LUT4AB/UserCLK Tile_X3Y2_LUT4AB/UserCLK
+ VGND VPWR Tile_X3Y3_LUT4AB/W1BEG[0] Tile_X3Y3_LUT4AB/W1BEG[1] Tile_X3Y3_LUT4AB/W1BEG[2]
+ Tile_X3Y3_LUT4AB/W1BEG[3] Tile_X3Y3_LUT4AB/W1END[0] Tile_X3Y3_LUT4AB/W1END[1] Tile_X3Y3_LUT4AB/W1END[2]
+ Tile_X3Y3_LUT4AB/W1END[3] Tile_X3Y3_LUT4AB/W2BEG[0] Tile_X3Y3_LUT4AB/W2BEG[1] Tile_X3Y3_LUT4AB/W2BEG[2]
+ Tile_X3Y3_LUT4AB/W2BEG[3] Tile_X3Y3_LUT4AB/W2BEG[4] Tile_X3Y3_LUT4AB/W2BEG[5] Tile_X3Y3_LUT4AB/W2BEG[6]
+ Tile_X3Y3_LUT4AB/W2BEG[7] Tile_X2Y3_LUT4AB/W2END[0] Tile_X2Y3_LUT4AB/W2END[1] Tile_X2Y3_LUT4AB/W2END[2]
+ Tile_X2Y3_LUT4AB/W2END[3] Tile_X2Y3_LUT4AB/W2END[4] Tile_X2Y3_LUT4AB/W2END[5] Tile_X2Y3_LUT4AB/W2END[6]
+ Tile_X2Y3_LUT4AB/W2END[7] Tile_X3Y3_LUT4AB/W2END[0] Tile_X3Y3_LUT4AB/W2END[1] Tile_X3Y3_LUT4AB/W2END[2]
+ Tile_X3Y3_LUT4AB/W2END[3] Tile_X3Y3_LUT4AB/W2END[4] Tile_X3Y3_LUT4AB/W2END[5] Tile_X3Y3_LUT4AB/W2END[6]
+ Tile_X3Y3_LUT4AB/W2END[7] Tile_X3Y3_LUT4AB/W2MID[0] Tile_X3Y3_LUT4AB/W2MID[1] Tile_X3Y3_LUT4AB/W2MID[2]
+ Tile_X3Y3_LUT4AB/W2MID[3] Tile_X3Y3_LUT4AB/W2MID[4] Tile_X3Y3_LUT4AB/W2MID[5] Tile_X3Y3_LUT4AB/W2MID[6]
+ Tile_X3Y3_LUT4AB/W2MID[7] Tile_X3Y3_LUT4AB/W6BEG[0] Tile_X3Y3_LUT4AB/W6BEG[10] Tile_X3Y3_LUT4AB/W6BEG[11]
+ Tile_X3Y3_LUT4AB/W6BEG[1] Tile_X3Y3_LUT4AB/W6BEG[2] Tile_X3Y3_LUT4AB/W6BEG[3] Tile_X3Y3_LUT4AB/W6BEG[4]
+ Tile_X3Y3_LUT4AB/W6BEG[5] Tile_X3Y3_LUT4AB/W6BEG[6] Tile_X3Y3_LUT4AB/W6BEG[7] Tile_X3Y3_LUT4AB/W6BEG[8]
+ Tile_X3Y3_LUT4AB/W6BEG[9] Tile_X3Y3_LUT4AB/W6END[0] Tile_X3Y3_LUT4AB/W6END[10] Tile_X3Y3_LUT4AB/W6END[11]
+ Tile_X3Y3_LUT4AB/W6END[1] Tile_X3Y3_LUT4AB/W6END[2] Tile_X3Y3_LUT4AB/W6END[3] Tile_X3Y3_LUT4AB/W6END[4]
+ Tile_X3Y3_LUT4AB/W6END[5] Tile_X3Y3_LUT4AB/W6END[6] Tile_X3Y3_LUT4AB/W6END[7] Tile_X3Y3_LUT4AB/W6END[8]
+ Tile_X3Y3_LUT4AB/W6END[9] Tile_X3Y3_LUT4AB/WW4BEG[0] Tile_X3Y3_LUT4AB/WW4BEG[10]
+ Tile_X3Y3_LUT4AB/WW4BEG[11] Tile_X3Y3_LUT4AB/WW4BEG[12] Tile_X3Y3_LUT4AB/WW4BEG[13]
+ Tile_X3Y3_LUT4AB/WW4BEG[14] Tile_X3Y3_LUT4AB/WW4BEG[15] Tile_X3Y3_LUT4AB/WW4BEG[1]
+ Tile_X3Y3_LUT4AB/WW4BEG[2] Tile_X3Y3_LUT4AB/WW4BEG[3] Tile_X3Y3_LUT4AB/WW4BEG[4]
+ Tile_X3Y3_LUT4AB/WW4BEG[5] Tile_X3Y3_LUT4AB/WW4BEG[6] Tile_X3Y3_LUT4AB/WW4BEG[7]
+ Tile_X3Y3_LUT4AB/WW4BEG[8] Tile_X3Y3_LUT4AB/WW4BEG[9] Tile_X3Y3_LUT4AB/WW4END[0]
+ Tile_X3Y3_LUT4AB/WW4END[10] Tile_X3Y3_LUT4AB/WW4END[11] Tile_X3Y3_LUT4AB/WW4END[12]
+ Tile_X3Y3_LUT4AB/WW4END[13] Tile_X3Y3_LUT4AB/WW4END[14] Tile_X3Y3_LUT4AB/WW4END[15]
+ Tile_X3Y3_LUT4AB/WW4END[1] Tile_X3Y3_LUT4AB/WW4END[2] Tile_X3Y3_LUT4AB/WW4END[3]
+ Tile_X3Y3_LUT4AB/WW4END[4] Tile_X3Y3_LUT4AB/WW4END[5] Tile_X3Y3_LUT4AB/WW4END[6]
+ Tile_X3Y3_LUT4AB/WW4END[7] Tile_X3Y3_LUT4AB/WW4END[8] Tile_X3Y3_LUT4AB/WW4END[9]
+ LUT4AB
XTile_X4Y3_RegFile Tile_X5Y3_LUT4AB/E1END[0] Tile_X5Y3_LUT4AB/E1END[1] Tile_X5Y3_LUT4AB/E1END[2]
+ Tile_X5Y3_LUT4AB/E1END[3] Tile_X3Y3_LUT4AB/E1BEG[0] Tile_X3Y3_LUT4AB/E1BEG[1] Tile_X3Y3_LUT4AB/E1BEG[2]
+ Tile_X3Y3_LUT4AB/E1BEG[3] Tile_X5Y3_LUT4AB/E2MID[0] Tile_X5Y3_LUT4AB/E2MID[1] Tile_X5Y3_LUT4AB/E2MID[2]
+ Tile_X5Y3_LUT4AB/E2MID[3] Tile_X5Y3_LUT4AB/E2MID[4] Tile_X5Y3_LUT4AB/E2MID[5] Tile_X5Y3_LUT4AB/E2MID[6]
+ Tile_X5Y3_LUT4AB/E2MID[7] Tile_X5Y3_LUT4AB/E2END[0] Tile_X5Y3_LUT4AB/E2END[1] Tile_X5Y3_LUT4AB/E2END[2]
+ Tile_X5Y3_LUT4AB/E2END[3] Tile_X5Y3_LUT4AB/E2END[4] Tile_X5Y3_LUT4AB/E2END[5] Tile_X5Y3_LUT4AB/E2END[6]
+ Tile_X5Y3_LUT4AB/E2END[7] Tile_X4Y3_RegFile/E2END[0] Tile_X4Y3_RegFile/E2END[1]
+ Tile_X4Y3_RegFile/E2END[2] Tile_X4Y3_RegFile/E2END[3] Tile_X4Y3_RegFile/E2END[4]
+ Tile_X4Y3_RegFile/E2END[5] Tile_X4Y3_RegFile/E2END[6] Tile_X4Y3_RegFile/E2END[7]
+ Tile_X3Y3_LUT4AB/E2BEG[0] Tile_X3Y3_LUT4AB/E2BEG[1] Tile_X3Y3_LUT4AB/E2BEG[2] Tile_X3Y3_LUT4AB/E2BEG[3]
+ Tile_X3Y3_LUT4AB/E2BEG[4] Tile_X3Y3_LUT4AB/E2BEG[5] Tile_X3Y3_LUT4AB/E2BEG[6] Tile_X3Y3_LUT4AB/E2BEG[7]
+ Tile_X5Y3_LUT4AB/E6END[0] Tile_X5Y3_LUT4AB/E6END[10] Tile_X5Y3_LUT4AB/E6END[11]
+ Tile_X5Y3_LUT4AB/E6END[1] Tile_X5Y3_LUT4AB/E6END[2] Tile_X5Y3_LUT4AB/E6END[3] Tile_X5Y3_LUT4AB/E6END[4]
+ Tile_X5Y3_LUT4AB/E6END[5] Tile_X5Y3_LUT4AB/E6END[6] Tile_X5Y3_LUT4AB/E6END[7] Tile_X5Y3_LUT4AB/E6END[8]
+ Tile_X5Y3_LUT4AB/E6END[9] Tile_X3Y3_LUT4AB/E6BEG[0] Tile_X3Y3_LUT4AB/E6BEG[10] Tile_X3Y3_LUT4AB/E6BEG[11]
+ Tile_X3Y3_LUT4AB/E6BEG[1] Tile_X3Y3_LUT4AB/E6BEG[2] Tile_X3Y3_LUT4AB/E6BEG[3] Tile_X3Y3_LUT4AB/E6BEG[4]
+ Tile_X3Y3_LUT4AB/E6BEG[5] Tile_X3Y3_LUT4AB/E6BEG[6] Tile_X3Y3_LUT4AB/E6BEG[7] Tile_X3Y3_LUT4AB/E6BEG[8]
+ Tile_X3Y3_LUT4AB/E6BEG[9] Tile_X5Y3_LUT4AB/EE4END[0] Tile_X5Y3_LUT4AB/EE4END[10]
+ Tile_X5Y3_LUT4AB/EE4END[11] Tile_X5Y3_LUT4AB/EE4END[12] Tile_X5Y3_LUT4AB/EE4END[13]
+ Tile_X5Y3_LUT4AB/EE4END[14] Tile_X5Y3_LUT4AB/EE4END[15] Tile_X5Y3_LUT4AB/EE4END[1]
+ Tile_X5Y3_LUT4AB/EE4END[2] Tile_X5Y3_LUT4AB/EE4END[3] Tile_X5Y3_LUT4AB/EE4END[4]
+ Tile_X5Y3_LUT4AB/EE4END[5] Tile_X5Y3_LUT4AB/EE4END[6] Tile_X5Y3_LUT4AB/EE4END[7]
+ Tile_X5Y3_LUT4AB/EE4END[8] Tile_X5Y3_LUT4AB/EE4END[9] Tile_X3Y3_LUT4AB/EE4BEG[0]
+ Tile_X3Y3_LUT4AB/EE4BEG[10] Tile_X3Y3_LUT4AB/EE4BEG[11] Tile_X3Y3_LUT4AB/EE4BEG[12]
+ Tile_X3Y3_LUT4AB/EE4BEG[13] Tile_X3Y3_LUT4AB/EE4BEG[14] Tile_X3Y3_LUT4AB/EE4BEG[15]
+ Tile_X3Y3_LUT4AB/EE4BEG[1] Tile_X3Y3_LUT4AB/EE4BEG[2] Tile_X3Y3_LUT4AB/EE4BEG[3]
+ Tile_X3Y3_LUT4AB/EE4BEG[4] Tile_X3Y3_LUT4AB/EE4BEG[5] Tile_X3Y3_LUT4AB/EE4BEG[6]
+ Tile_X3Y3_LUT4AB/EE4BEG[7] Tile_X3Y3_LUT4AB/EE4BEG[8] Tile_X3Y3_LUT4AB/EE4BEG[9]
+ Tile_X4Y3_RegFile/FrameData[0] Tile_X4Y3_RegFile/FrameData[10] Tile_X4Y3_RegFile/FrameData[11]
+ Tile_X4Y3_RegFile/FrameData[12] Tile_X4Y3_RegFile/FrameData[13] Tile_X4Y3_RegFile/FrameData[14]
+ Tile_X4Y3_RegFile/FrameData[15] Tile_X4Y3_RegFile/FrameData[16] Tile_X4Y3_RegFile/FrameData[17]
+ Tile_X4Y3_RegFile/FrameData[18] Tile_X4Y3_RegFile/FrameData[19] Tile_X4Y3_RegFile/FrameData[1]
+ Tile_X4Y3_RegFile/FrameData[20] Tile_X4Y3_RegFile/FrameData[21] Tile_X4Y3_RegFile/FrameData[22]
+ Tile_X4Y3_RegFile/FrameData[23] Tile_X4Y3_RegFile/FrameData[24] Tile_X4Y3_RegFile/FrameData[25]
+ Tile_X4Y3_RegFile/FrameData[26] Tile_X4Y3_RegFile/FrameData[27] Tile_X4Y3_RegFile/FrameData[28]
+ Tile_X4Y3_RegFile/FrameData[29] Tile_X4Y3_RegFile/FrameData[2] Tile_X4Y3_RegFile/FrameData[30]
+ Tile_X4Y3_RegFile/FrameData[31] Tile_X4Y3_RegFile/FrameData[3] Tile_X4Y3_RegFile/FrameData[4]
+ Tile_X4Y3_RegFile/FrameData[5] Tile_X4Y3_RegFile/FrameData[6] Tile_X4Y3_RegFile/FrameData[7]
+ Tile_X4Y3_RegFile/FrameData[8] Tile_X4Y3_RegFile/FrameData[9] Tile_X5Y3_LUT4AB/FrameData[0]
+ Tile_X5Y3_LUT4AB/FrameData[10] Tile_X5Y3_LUT4AB/FrameData[11] Tile_X5Y3_LUT4AB/FrameData[12]
+ Tile_X5Y3_LUT4AB/FrameData[13] Tile_X5Y3_LUT4AB/FrameData[14] Tile_X5Y3_LUT4AB/FrameData[15]
+ Tile_X5Y3_LUT4AB/FrameData[16] Tile_X5Y3_LUT4AB/FrameData[17] Tile_X5Y3_LUT4AB/FrameData[18]
+ Tile_X5Y3_LUT4AB/FrameData[19] Tile_X5Y3_LUT4AB/FrameData[1] Tile_X5Y3_LUT4AB/FrameData[20]
+ Tile_X5Y3_LUT4AB/FrameData[21] Tile_X5Y3_LUT4AB/FrameData[22] Tile_X5Y3_LUT4AB/FrameData[23]
+ Tile_X5Y3_LUT4AB/FrameData[24] Tile_X5Y3_LUT4AB/FrameData[25] Tile_X5Y3_LUT4AB/FrameData[26]
+ Tile_X5Y3_LUT4AB/FrameData[27] Tile_X5Y3_LUT4AB/FrameData[28] Tile_X5Y3_LUT4AB/FrameData[29]
+ Tile_X5Y3_LUT4AB/FrameData[2] Tile_X5Y3_LUT4AB/FrameData[30] Tile_X5Y3_LUT4AB/FrameData[31]
+ Tile_X5Y3_LUT4AB/FrameData[3] Tile_X5Y3_LUT4AB/FrameData[4] Tile_X5Y3_LUT4AB/FrameData[5]
+ Tile_X5Y3_LUT4AB/FrameData[6] Tile_X5Y3_LUT4AB/FrameData[7] Tile_X5Y3_LUT4AB/FrameData[8]
+ Tile_X5Y3_LUT4AB/FrameData[9] Tile_X4Y3_RegFile/FrameStrobe[0] Tile_X4Y3_RegFile/FrameStrobe[10]
+ Tile_X4Y3_RegFile/FrameStrobe[11] Tile_X4Y3_RegFile/FrameStrobe[12] Tile_X4Y3_RegFile/FrameStrobe[13]
+ Tile_X4Y3_RegFile/FrameStrobe[14] Tile_X4Y3_RegFile/FrameStrobe[15] Tile_X4Y3_RegFile/FrameStrobe[16]
+ Tile_X4Y3_RegFile/FrameStrobe[17] Tile_X4Y3_RegFile/FrameStrobe[18] Tile_X4Y3_RegFile/FrameStrobe[19]
+ Tile_X4Y3_RegFile/FrameStrobe[1] Tile_X4Y3_RegFile/FrameStrobe[2] Tile_X4Y3_RegFile/FrameStrobe[3]
+ Tile_X4Y3_RegFile/FrameStrobe[4] Tile_X4Y3_RegFile/FrameStrobe[5] Tile_X4Y3_RegFile/FrameStrobe[6]
+ Tile_X4Y3_RegFile/FrameStrobe[7] Tile_X4Y3_RegFile/FrameStrobe[8] Tile_X4Y3_RegFile/FrameStrobe[9]
+ Tile_X4Y2_RegFile/FrameStrobe[0] Tile_X4Y2_RegFile/FrameStrobe[10] Tile_X4Y2_RegFile/FrameStrobe[11]
+ Tile_X4Y2_RegFile/FrameStrobe[12] Tile_X4Y2_RegFile/FrameStrobe[13] Tile_X4Y2_RegFile/FrameStrobe[14]
+ Tile_X4Y2_RegFile/FrameStrobe[15] Tile_X4Y2_RegFile/FrameStrobe[16] Tile_X4Y2_RegFile/FrameStrobe[17]
+ Tile_X4Y2_RegFile/FrameStrobe[18] Tile_X4Y2_RegFile/FrameStrobe[19] Tile_X4Y2_RegFile/FrameStrobe[1]
+ Tile_X4Y2_RegFile/FrameStrobe[2] Tile_X4Y2_RegFile/FrameStrobe[3] Tile_X4Y2_RegFile/FrameStrobe[4]
+ Tile_X4Y2_RegFile/FrameStrobe[5] Tile_X4Y2_RegFile/FrameStrobe[6] Tile_X4Y2_RegFile/FrameStrobe[7]
+ Tile_X4Y2_RegFile/FrameStrobe[8] Tile_X4Y2_RegFile/FrameStrobe[9] Tile_X4Y3_RegFile/N1BEG[0]
+ Tile_X4Y3_RegFile/N1BEG[1] Tile_X4Y3_RegFile/N1BEG[2] Tile_X4Y3_RegFile/N1BEG[3]
+ Tile_X4Y4_RegFile/N1BEG[0] Tile_X4Y4_RegFile/N1BEG[1] Tile_X4Y4_RegFile/N1BEG[2]
+ Tile_X4Y4_RegFile/N1BEG[3] Tile_X4Y3_RegFile/N2BEG[0] Tile_X4Y3_RegFile/N2BEG[1]
+ Tile_X4Y3_RegFile/N2BEG[2] Tile_X4Y3_RegFile/N2BEG[3] Tile_X4Y3_RegFile/N2BEG[4]
+ Tile_X4Y3_RegFile/N2BEG[5] Tile_X4Y3_RegFile/N2BEG[6] Tile_X4Y3_RegFile/N2BEG[7]
+ Tile_X4Y2_RegFile/N2END[0] Tile_X4Y2_RegFile/N2END[1] Tile_X4Y2_RegFile/N2END[2]
+ Tile_X4Y2_RegFile/N2END[3] Tile_X4Y2_RegFile/N2END[4] Tile_X4Y2_RegFile/N2END[5]
+ Tile_X4Y2_RegFile/N2END[6] Tile_X4Y2_RegFile/N2END[7] Tile_X4Y3_RegFile/N2END[0]
+ Tile_X4Y3_RegFile/N2END[1] Tile_X4Y3_RegFile/N2END[2] Tile_X4Y3_RegFile/N2END[3]
+ Tile_X4Y3_RegFile/N2END[4] Tile_X4Y3_RegFile/N2END[5] Tile_X4Y3_RegFile/N2END[6]
+ Tile_X4Y3_RegFile/N2END[7] Tile_X4Y4_RegFile/N2BEG[0] Tile_X4Y4_RegFile/N2BEG[1]
+ Tile_X4Y4_RegFile/N2BEG[2] Tile_X4Y4_RegFile/N2BEG[3] Tile_X4Y4_RegFile/N2BEG[4]
+ Tile_X4Y4_RegFile/N2BEG[5] Tile_X4Y4_RegFile/N2BEG[6] Tile_X4Y4_RegFile/N2BEG[7]
+ Tile_X4Y3_RegFile/N4BEG[0] Tile_X4Y3_RegFile/N4BEG[10] Tile_X4Y3_RegFile/N4BEG[11]
+ Tile_X4Y3_RegFile/N4BEG[12] Tile_X4Y3_RegFile/N4BEG[13] Tile_X4Y3_RegFile/N4BEG[14]
+ Tile_X4Y3_RegFile/N4BEG[15] Tile_X4Y3_RegFile/N4BEG[1] Tile_X4Y3_RegFile/N4BEG[2]
+ Tile_X4Y3_RegFile/N4BEG[3] Tile_X4Y3_RegFile/N4BEG[4] Tile_X4Y3_RegFile/N4BEG[5]
+ Tile_X4Y3_RegFile/N4BEG[6] Tile_X4Y3_RegFile/N4BEG[7] Tile_X4Y3_RegFile/N4BEG[8]
+ Tile_X4Y3_RegFile/N4BEG[9] Tile_X4Y4_RegFile/N4BEG[0] Tile_X4Y4_RegFile/N4BEG[10]
+ Tile_X4Y4_RegFile/N4BEG[11] Tile_X4Y4_RegFile/N4BEG[12] Tile_X4Y4_RegFile/N4BEG[13]
+ Tile_X4Y4_RegFile/N4BEG[14] Tile_X4Y4_RegFile/N4BEG[15] Tile_X4Y4_RegFile/N4BEG[1]
+ Tile_X4Y4_RegFile/N4BEG[2] Tile_X4Y4_RegFile/N4BEG[3] Tile_X4Y4_RegFile/N4BEG[4]
+ Tile_X4Y4_RegFile/N4BEG[5] Tile_X4Y4_RegFile/N4BEG[6] Tile_X4Y4_RegFile/N4BEG[7]
+ Tile_X4Y4_RegFile/N4BEG[8] Tile_X4Y4_RegFile/N4BEG[9] Tile_X4Y3_RegFile/NN4BEG[0]
+ Tile_X4Y3_RegFile/NN4BEG[10] Tile_X4Y3_RegFile/NN4BEG[11] Tile_X4Y3_RegFile/NN4BEG[12]
+ Tile_X4Y3_RegFile/NN4BEG[13] Tile_X4Y3_RegFile/NN4BEG[14] Tile_X4Y3_RegFile/NN4BEG[15]
+ Tile_X4Y3_RegFile/NN4BEG[1] Tile_X4Y3_RegFile/NN4BEG[2] Tile_X4Y3_RegFile/NN4BEG[3]
+ Tile_X4Y3_RegFile/NN4BEG[4] Tile_X4Y3_RegFile/NN4BEG[5] Tile_X4Y3_RegFile/NN4BEG[6]
+ Tile_X4Y3_RegFile/NN4BEG[7] Tile_X4Y3_RegFile/NN4BEG[8] Tile_X4Y3_RegFile/NN4BEG[9]
+ Tile_X4Y4_RegFile/NN4BEG[0] Tile_X4Y4_RegFile/NN4BEG[10] Tile_X4Y4_RegFile/NN4BEG[11]
+ Tile_X4Y4_RegFile/NN4BEG[12] Tile_X4Y4_RegFile/NN4BEG[13] Tile_X4Y4_RegFile/NN4BEG[14]
+ Tile_X4Y4_RegFile/NN4BEG[15] Tile_X4Y4_RegFile/NN4BEG[1] Tile_X4Y4_RegFile/NN4BEG[2]
+ Tile_X4Y4_RegFile/NN4BEG[3] Tile_X4Y4_RegFile/NN4BEG[4] Tile_X4Y4_RegFile/NN4BEG[5]
+ Tile_X4Y4_RegFile/NN4BEG[6] Tile_X4Y4_RegFile/NN4BEG[7] Tile_X4Y4_RegFile/NN4BEG[8]
+ Tile_X4Y4_RegFile/NN4BEG[9] Tile_X4Y4_RegFile/S1END[0] Tile_X4Y4_RegFile/S1END[1]
+ Tile_X4Y4_RegFile/S1END[2] Tile_X4Y4_RegFile/S1END[3] Tile_X4Y3_RegFile/S1END[0]
+ Tile_X4Y3_RegFile/S1END[1] Tile_X4Y3_RegFile/S1END[2] Tile_X4Y3_RegFile/S1END[3]
+ Tile_X4Y4_RegFile/S2MID[0] Tile_X4Y4_RegFile/S2MID[1] Tile_X4Y4_RegFile/S2MID[2]
+ Tile_X4Y4_RegFile/S2MID[3] Tile_X4Y4_RegFile/S2MID[4] Tile_X4Y4_RegFile/S2MID[5]
+ Tile_X4Y4_RegFile/S2MID[6] Tile_X4Y4_RegFile/S2MID[7] Tile_X4Y4_RegFile/S2END[0]
+ Tile_X4Y4_RegFile/S2END[1] Tile_X4Y4_RegFile/S2END[2] Tile_X4Y4_RegFile/S2END[3]
+ Tile_X4Y4_RegFile/S2END[4] Tile_X4Y4_RegFile/S2END[5] Tile_X4Y4_RegFile/S2END[6]
+ Tile_X4Y4_RegFile/S2END[7] Tile_X4Y3_RegFile/S2END[0] Tile_X4Y3_RegFile/S2END[1]
+ Tile_X4Y3_RegFile/S2END[2] Tile_X4Y3_RegFile/S2END[3] Tile_X4Y3_RegFile/S2END[4]
+ Tile_X4Y3_RegFile/S2END[5] Tile_X4Y3_RegFile/S2END[6] Tile_X4Y3_RegFile/S2END[7]
+ Tile_X4Y3_RegFile/S2MID[0] Tile_X4Y3_RegFile/S2MID[1] Tile_X4Y3_RegFile/S2MID[2]
+ Tile_X4Y3_RegFile/S2MID[3] Tile_X4Y3_RegFile/S2MID[4] Tile_X4Y3_RegFile/S2MID[5]
+ Tile_X4Y3_RegFile/S2MID[6] Tile_X4Y3_RegFile/S2MID[7] Tile_X4Y4_RegFile/S4END[0]
+ Tile_X4Y4_RegFile/S4END[10] Tile_X4Y4_RegFile/S4END[11] Tile_X4Y4_RegFile/S4END[12]
+ Tile_X4Y4_RegFile/S4END[13] Tile_X4Y4_RegFile/S4END[14] Tile_X4Y4_RegFile/S4END[15]
+ Tile_X4Y4_RegFile/S4END[1] Tile_X4Y4_RegFile/S4END[2] Tile_X4Y4_RegFile/S4END[3]
+ Tile_X4Y4_RegFile/S4END[4] Tile_X4Y4_RegFile/S4END[5] Tile_X4Y4_RegFile/S4END[6]
+ Tile_X4Y4_RegFile/S4END[7] Tile_X4Y4_RegFile/S4END[8] Tile_X4Y4_RegFile/S4END[9]
+ Tile_X4Y3_RegFile/S4END[0] Tile_X4Y3_RegFile/S4END[10] Tile_X4Y3_RegFile/S4END[11]
+ Tile_X4Y3_RegFile/S4END[12] Tile_X4Y3_RegFile/S4END[13] Tile_X4Y3_RegFile/S4END[14]
+ Tile_X4Y3_RegFile/S4END[15] Tile_X4Y3_RegFile/S4END[1] Tile_X4Y3_RegFile/S4END[2]
+ Tile_X4Y3_RegFile/S4END[3] Tile_X4Y3_RegFile/S4END[4] Tile_X4Y3_RegFile/S4END[5]
+ Tile_X4Y3_RegFile/S4END[6] Tile_X4Y3_RegFile/S4END[7] Tile_X4Y3_RegFile/S4END[8]
+ Tile_X4Y3_RegFile/S4END[9] Tile_X4Y4_RegFile/SS4END[0] Tile_X4Y4_RegFile/SS4END[10]
+ Tile_X4Y4_RegFile/SS4END[11] Tile_X4Y4_RegFile/SS4END[12] Tile_X4Y4_RegFile/SS4END[13]
+ Tile_X4Y4_RegFile/SS4END[14] Tile_X4Y4_RegFile/SS4END[15] Tile_X4Y4_RegFile/SS4END[1]
+ Tile_X4Y4_RegFile/SS4END[2] Tile_X4Y4_RegFile/SS4END[3] Tile_X4Y4_RegFile/SS4END[4]
+ Tile_X4Y4_RegFile/SS4END[5] Tile_X4Y4_RegFile/SS4END[6] Tile_X4Y4_RegFile/SS4END[7]
+ Tile_X4Y4_RegFile/SS4END[8] Tile_X4Y4_RegFile/SS4END[9] Tile_X4Y3_RegFile/SS4END[0]
+ Tile_X4Y3_RegFile/SS4END[10] Tile_X4Y3_RegFile/SS4END[11] Tile_X4Y3_RegFile/SS4END[12]
+ Tile_X4Y3_RegFile/SS4END[13] Tile_X4Y3_RegFile/SS4END[14] Tile_X4Y3_RegFile/SS4END[15]
+ Tile_X4Y3_RegFile/SS4END[1] Tile_X4Y3_RegFile/SS4END[2] Tile_X4Y3_RegFile/SS4END[3]
+ Tile_X4Y3_RegFile/SS4END[4] Tile_X4Y3_RegFile/SS4END[5] Tile_X4Y3_RegFile/SS4END[6]
+ Tile_X4Y3_RegFile/SS4END[7] Tile_X4Y3_RegFile/SS4END[8] Tile_X4Y3_RegFile/SS4END[9]
+ Tile_X4Y3_RegFile/UserCLK Tile_X4Y2_RegFile/UserCLK VGND VPWR Tile_X3Y3_LUT4AB/W1END[0]
+ Tile_X3Y3_LUT4AB/W1END[1] Tile_X3Y3_LUT4AB/W1END[2] Tile_X3Y3_LUT4AB/W1END[3] Tile_X5Y3_LUT4AB/W1BEG[0]
+ Tile_X5Y3_LUT4AB/W1BEG[1] Tile_X5Y3_LUT4AB/W1BEG[2] Tile_X5Y3_LUT4AB/W1BEG[3] Tile_X3Y3_LUT4AB/W2MID[0]
+ Tile_X3Y3_LUT4AB/W2MID[1] Tile_X3Y3_LUT4AB/W2MID[2] Tile_X3Y3_LUT4AB/W2MID[3] Tile_X3Y3_LUT4AB/W2MID[4]
+ Tile_X3Y3_LUT4AB/W2MID[5] Tile_X3Y3_LUT4AB/W2MID[6] Tile_X3Y3_LUT4AB/W2MID[7] Tile_X3Y3_LUT4AB/W2END[0]
+ Tile_X3Y3_LUT4AB/W2END[1] Tile_X3Y3_LUT4AB/W2END[2] Tile_X3Y3_LUT4AB/W2END[3] Tile_X3Y3_LUT4AB/W2END[4]
+ Tile_X3Y3_LUT4AB/W2END[5] Tile_X3Y3_LUT4AB/W2END[6] Tile_X3Y3_LUT4AB/W2END[7] Tile_X5Y3_LUT4AB/W2BEGb[0]
+ Tile_X5Y3_LUT4AB/W2BEGb[1] Tile_X5Y3_LUT4AB/W2BEGb[2] Tile_X5Y3_LUT4AB/W2BEGb[3]
+ Tile_X5Y3_LUT4AB/W2BEGb[4] Tile_X5Y3_LUT4AB/W2BEGb[5] Tile_X5Y3_LUT4AB/W2BEGb[6]
+ Tile_X5Y3_LUT4AB/W2BEGb[7] Tile_X5Y3_LUT4AB/W2BEG[0] Tile_X5Y3_LUT4AB/W2BEG[1] Tile_X5Y3_LUT4AB/W2BEG[2]
+ Tile_X5Y3_LUT4AB/W2BEG[3] Tile_X5Y3_LUT4AB/W2BEG[4] Tile_X5Y3_LUT4AB/W2BEG[5] Tile_X5Y3_LUT4AB/W2BEG[6]
+ Tile_X5Y3_LUT4AB/W2BEG[7] Tile_X3Y3_LUT4AB/W6END[0] Tile_X3Y3_LUT4AB/W6END[10] Tile_X3Y3_LUT4AB/W6END[11]
+ Tile_X3Y3_LUT4AB/W6END[1] Tile_X3Y3_LUT4AB/W6END[2] Tile_X3Y3_LUT4AB/W6END[3] Tile_X3Y3_LUT4AB/W6END[4]
+ Tile_X3Y3_LUT4AB/W6END[5] Tile_X3Y3_LUT4AB/W6END[6] Tile_X3Y3_LUT4AB/W6END[7] Tile_X3Y3_LUT4AB/W6END[8]
+ Tile_X3Y3_LUT4AB/W6END[9] Tile_X5Y3_LUT4AB/W6BEG[0] Tile_X5Y3_LUT4AB/W6BEG[10] Tile_X5Y3_LUT4AB/W6BEG[11]
+ Tile_X5Y3_LUT4AB/W6BEG[1] Tile_X5Y3_LUT4AB/W6BEG[2] Tile_X5Y3_LUT4AB/W6BEG[3] Tile_X5Y3_LUT4AB/W6BEG[4]
+ Tile_X5Y3_LUT4AB/W6BEG[5] Tile_X5Y3_LUT4AB/W6BEG[6] Tile_X5Y3_LUT4AB/W6BEG[7] Tile_X5Y3_LUT4AB/W6BEG[8]
+ Tile_X5Y3_LUT4AB/W6BEG[9] Tile_X3Y3_LUT4AB/WW4END[0] Tile_X3Y3_LUT4AB/WW4END[10]
+ Tile_X3Y3_LUT4AB/WW4END[11] Tile_X3Y3_LUT4AB/WW4END[12] Tile_X3Y3_LUT4AB/WW4END[13]
+ Tile_X3Y3_LUT4AB/WW4END[14] Tile_X3Y3_LUT4AB/WW4END[15] Tile_X3Y3_LUT4AB/WW4END[1]
+ Tile_X3Y3_LUT4AB/WW4END[2] Tile_X3Y3_LUT4AB/WW4END[3] Tile_X3Y3_LUT4AB/WW4END[4]
+ Tile_X3Y3_LUT4AB/WW4END[5] Tile_X3Y3_LUT4AB/WW4END[6] Tile_X3Y3_LUT4AB/WW4END[7]
+ Tile_X3Y3_LUT4AB/WW4END[8] Tile_X3Y3_LUT4AB/WW4END[9] Tile_X5Y3_LUT4AB/WW4BEG[0]
+ Tile_X5Y3_LUT4AB/WW4BEG[10] Tile_X5Y3_LUT4AB/WW4BEG[11] Tile_X5Y3_LUT4AB/WW4BEG[12]
+ Tile_X5Y3_LUT4AB/WW4BEG[13] Tile_X5Y3_LUT4AB/WW4BEG[14] Tile_X5Y3_LUT4AB/WW4BEG[15]
+ Tile_X5Y3_LUT4AB/WW4BEG[1] Tile_X5Y3_LUT4AB/WW4BEG[2] Tile_X5Y3_LUT4AB/WW4BEG[3]
+ Tile_X5Y3_LUT4AB/WW4BEG[4] Tile_X5Y3_LUT4AB/WW4BEG[5] Tile_X5Y3_LUT4AB/WW4BEG[6]
+ Tile_X5Y3_LUT4AB/WW4BEG[7] Tile_X5Y3_LUT4AB/WW4BEG[8] Tile_X5Y3_LUT4AB/WW4BEG[9]
+ RegFile
XTile_X10Y15_S_term_IHP_SRAM Tile_X9Y15_S_CPU_IF/FrameData_O[0] Tile_X9Y15_S_CPU_IF/FrameData_O[10]
+ Tile_X9Y15_S_CPU_IF/FrameData_O[11] Tile_X9Y15_S_CPU_IF/FrameData_O[12] Tile_X9Y15_S_CPU_IF/FrameData_O[13]
+ Tile_X9Y15_S_CPU_IF/FrameData_O[14] Tile_X9Y15_S_CPU_IF/FrameData_O[15] Tile_X9Y15_S_CPU_IF/FrameData_O[16]
+ Tile_X9Y15_S_CPU_IF/FrameData_O[17] Tile_X9Y15_S_CPU_IF/FrameData_O[18] Tile_X9Y15_S_CPU_IF/FrameData_O[19]
+ Tile_X9Y15_S_CPU_IF/FrameData_O[1] Tile_X9Y15_S_CPU_IF/FrameData_O[20] Tile_X9Y15_S_CPU_IF/FrameData_O[21]
+ Tile_X9Y15_S_CPU_IF/FrameData_O[22] Tile_X9Y15_S_CPU_IF/FrameData_O[23] Tile_X9Y15_S_CPU_IF/FrameData_O[24]
+ Tile_X9Y15_S_CPU_IF/FrameData_O[25] Tile_X9Y15_S_CPU_IF/FrameData_O[26] Tile_X9Y15_S_CPU_IF/FrameData_O[27]
+ Tile_X9Y15_S_CPU_IF/FrameData_O[28] Tile_X9Y15_S_CPU_IF/FrameData_O[29] Tile_X9Y15_S_CPU_IF/FrameData_O[2]
+ Tile_X9Y15_S_CPU_IF/FrameData_O[30] Tile_X9Y15_S_CPU_IF/FrameData_O[31] Tile_X9Y15_S_CPU_IF/FrameData_O[3]
+ Tile_X9Y15_S_CPU_IF/FrameData_O[4] Tile_X9Y15_S_CPU_IF/FrameData_O[5] Tile_X9Y15_S_CPU_IF/FrameData_O[6]
+ Tile_X9Y15_S_CPU_IF/FrameData_O[7] Tile_X9Y15_S_CPU_IF/FrameData_O[8] Tile_X9Y15_S_CPU_IF/FrameData_O[9]
+ Tile_X10Y15_S_term_IHP_SRAM/FrameData_O[0] Tile_X10Y15_S_term_IHP_SRAM/FrameData_O[10]
+ Tile_X10Y15_S_term_IHP_SRAM/FrameData_O[11] Tile_X10Y15_S_term_IHP_SRAM/FrameData_O[12]
+ Tile_X10Y15_S_term_IHP_SRAM/FrameData_O[13] Tile_X10Y15_S_term_IHP_SRAM/FrameData_O[14]
+ Tile_X10Y15_S_term_IHP_SRAM/FrameData_O[15] Tile_X10Y15_S_term_IHP_SRAM/FrameData_O[16]
+ Tile_X10Y15_S_term_IHP_SRAM/FrameData_O[17] Tile_X10Y15_S_term_IHP_SRAM/FrameData_O[18]
+ Tile_X10Y15_S_term_IHP_SRAM/FrameData_O[19] Tile_X10Y15_S_term_IHP_SRAM/FrameData_O[1]
+ Tile_X10Y15_S_term_IHP_SRAM/FrameData_O[20] Tile_X10Y15_S_term_IHP_SRAM/FrameData_O[21]
+ Tile_X10Y15_S_term_IHP_SRAM/FrameData_O[22] Tile_X10Y15_S_term_IHP_SRAM/FrameData_O[23]
+ Tile_X10Y15_S_term_IHP_SRAM/FrameData_O[24] Tile_X10Y15_S_term_IHP_SRAM/FrameData_O[25]
+ Tile_X10Y15_S_term_IHP_SRAM/FrameData_O[26] Tile_X10Y15_S_term_IHP_SRAM/FrameData_O[27]
+ Tile_X10Y15_S_term_IHP_SRAM/FrameData_O[28] Tile_X10Y15_S_term_IHP_SRAM/FrameData_O[29]
+ Tile_X10Y15_S_term_IHP_SRAM/FrameData_O[2] Tile_X10Y15_S_term_IHP_SRAM/FrameData_O[30]
+ Tile_X10Y15_S_term_IHP_SRAM/FrameData_O[31] Tile_X10Y15_S_term_IHP_SRAM/FrameData_O[3]
+ Tile_X10Y15_S_term_IHP_SRAM/FrameData_O[4] Tile_X10Y15_S_term_IHP_SRAM/FrameData_O[5]
+ Tile_X10Y15_S_term_IHP_SRAM/FrameData_O[6] Tile_X10Y15_S_term_IHP_SRAM/FrameData_O[7]
+ Tile_X10Y15_S_term_IHP_SRAM/FrameData_O[8] Tile_X10Y15_S_term_IHP_SRAM/FrameData_O[9]
+ FrameStrobe[200] FrameStrobe[210] FrameStrobe[211] FrameStrobe[212] FrameStrobe[213]
+ FrameStrobe[214] FrameStrobe[215] FrameStrobe[216] FrameStrobe[217] FrameStrobe[218]
+ FrameStrobe[219] FrameStrobe[201] FrameStrobe[202] FrameStrobe[203] FrameStrobe[204]
+ FrameStrobe[205] FrameStrobe[206] FrameStrobe[207] FrameStrobe[208] FrameStrobe[209]
+ Tile_X10Y15_S_term_IHP_SRAM/FrameStrobe_O[0] Tile_X10Y15_S_term_IHP_SRAM/FrameStrobe_O[10]
+ Tile_X10Y15_S_term_IHP_SRAM/FrameStrobe_O[11] Tile_X10Y15_S_term_IHP_SRAM/FrameStrobe_O[12]
+ Tile_X10Y15_S_term_IHP_SRAM/FrameStrobe_O[13] Tile_X10Y15_S_term_IHP_SRAM/FrameStrobe_O[14]
+ Tile_X10Y15_S_term_IHP_SRAM/FrameStrobe_O[15] Tile_X10Y15_S_term_IHP_SRAM/FrameStrobe_O[16]
+ Tile_X10Y15_S_term_IHP_SRAM/FrameStrobe_O[17] Tile_X10Y15_S_term_IHP_SRAM/FrameStrobe_O[18]
+ Tile_X10Y15_S_term_IHP_SRAM/FrameStrobe_O[19] Tile_X10Y15_S_term_IHP_SRAM/FrameStrobe_O[1]
+ Tile_X10Y15_S_term_IHP_SRAM/FrameStrobe_O[2] Tile_X10Y15_S_term_IHP_SRAM/FrameStrobe_O[3]
+ Tile_X10Y15_S_term_IHP_SRAM/FrameStrobe_O[4] Tile_X10Y15_S_term_IHP_SRAM/FrameStrobe_O[5]
+ Tile_X10Y15_S_term_IHP_SRAM/FrameStrobe_O[6] Tile_X10Y15_S_term_IHP_SRAM/FrameStrobe_O[7]
+ Tile_X10Y15_S_term_IHP_SRAM/FrameStrobe_O[8] Tile_X10Y15_S_term_IHP_SRAM/FrameStrobe_O[9]
+ Tile_X10Y15_S_term_IHP_SRAM/N1BEG[0] Tile_X10Y15_S_term_IHP_SRAM/N1BEG[1] Tile_X10Y15_S_term_IHP_SRAM/N1BEG[2]
+ Tile_X10Y15_S_term_IHP_SRAM/N1BEG[3] Tile_X10Y15_S_term_IHP_SRAM/N2BEG[0] Tile_X10Y15_S_term_IHP_SRAM/N2BEG[1]
+ Tile_X10Y15_S_term_IHP_SRAM/N2BEG[2] Tile_X10Y15_S_term_IHP_SRAM/N2BEG[3] Tile_X10Y15_S_term_IHP_SRAM/N2BEG[4]
+ Tile_X10Y15_S_term_IHP_SRAM/N2BEG[5] Tile_X10Y15_S_term_IHP_SRAM/N2BEG[6] Tile_X10Y15_S_term_IHP_SRAM/N2BEG[7]
+ Tile_X10Y15_S_term_IHP_SRAM/N2BEGb[0] Tile_X10Y15_S_term_IHP_SRAM/N2BEGb[1] Tile_X10Y15_S_term_IHP_SRAM/N2BEGb[2]
+ Tile_X10Y15_S_term_IHP_SRAM/N2BEGb[3] Tile_X10Y15_S_term_IHP_SRAM/N2BEGb[4] Tile_X10Y15_S_term_IHP_SRAM/N2BEGb[5]
+ Tile_X10Y15_S_term_IHP_SRAM/N2BEGb[6] Tile_X10Y15_S_term_IHP_SRAM/N2BEGb[7] Tile_X10Y15_S_term_IHP_SRAM/N4BEG[0]
+ Tile_X10Y15_S_term_IHP_SRAM/N4BEG[10] Tile_X10Y15_S_term_IHP_SRAM/N4BEG[11] Tile_X10Y15_S_term_IHP_SRAM/N4BEG[12]
+ Tile_X10Y15_S_term_IHP_SRAM/N4BEG[13] Tile_X10Y15_S_term_IHP_SRAM/N4BEG[14] Tile_X10Y15_S_term_IHP_SRAM/N4BEG[15]
+ Tile_X10Y15_S_term_IHP_SRAM/N4BEG[1] Tile_X10Y15_S_term_IHP_SRAM/N4BEG[2] Tile_X10Y15_S_term_IHP_SRAM/N4BEG[3]
+ Tile_X10Y15_S_term_IHP_SRAM/N4BEG[4] Tile_X10Y15_S_term_IHP_SRAM/N4BEG[5] Tile_X10Y15_S_term_IHP_SRAM/N4BEG[6]
+ Tile_X10Y15_S_term_IHP_SRAM/N4BEG[7] Tile_X10Y15_S_term_IHP_SRAM/N4BEG[8] Tile_X10Y15_S_term_IHP_SRAM/N4BEG[9]
+ Tile_X10Y15_S_term_IHP_SRAM/S1END[0] Tile_X10Y15_S_term_IHP_SRAM/S1END[1] Tile_X10Y15_S_term_IHP_SRAM/S1END[2]
+ Tile_X10Y15_S_term_IHP_SRAM/S1END[3] Tile_X10Y15_S_term_IHP_SRAM/S2END[0] Tile_X10Y15_S_term_IHP_SRAM/S2END[1]
+ Tile_X10Y15_S_term_IHP_SRAM/S2END[2] Tile_X10Y15_S_term_IHP_SRAM/S2END[3] Tile_X10Y15_S_term_IHP_SRAM/S2END[4]
+ Tile_X10Y15_S_term_IHP_SRAM/S2END[5] Tile_X10Y15_S_term_IHP_SRAM/S2END[6] Tile_X10Y15_S_term_IHP_SRAM/S2END[7]
+ Tile_X10Y15_S_term_IHP_SRAM/S2MID[0] Tile_X10Y15_S_term_IHP_SRAM/S2MID[1] Tile_X10Y15_S_term_IHP_SRAM/S2MID[2]
+ Tile_X10Y15_S_term_IHP_SRAM/S2MID[3] Tile_X10Y15_S_term_IHP_SRAM/S2MID[4] Tile_X10Y15_S_term_IHP_SRAM/S2MID[5]
+ Tile_X10Y15_S_term_IHP_SRAM/S2MID[6] Tile_X10Y15_S_term_IHP_SRAM/S2MID[7] Tile_X10Y15_S_term_IHP_SRAM/S4END[0]
+ Tile_X10Y15_S_term_IHP_SRAM/S4END[10] Tile_X10Y15_S_term_IHP_SRAM/S4END[11] Tile_X10Y15_S_term_IHP_SRAM/S4END[12]
+ Tile_X10Y15_S_term_IHP_SRAM/S4END[13] Tile_X10Y15_S_term_IHP_SRAM/S4END[14] Tile_X10Y15_S_term_IHP_SRAM/S4END[15]
+ Tile_X10Y15_S_term_IHP_SRAM/S4END[1] Tile_X10Y15_S_term_IHP_SRAM/S4END[2] Tile_X10Y15_S_term_IHP_SRAM/S4END[3]
+ Tile_X10Y15_S_term_IHP_SRAM/S4END[4] Tile_X10Y15_S_term_IHP_SRAM/S4END[5] Tile_X10Y15_S_term_IHP_SRAM/S4END[6]
+ Tile_X10Y15_S_term_IHP_SRAM/S4END[7] Tile_X10Y15_S_term_IHP_SRAM/S4END[8] Tile_X10Y15_S_term_IHP_SRAM/S4END[9]
+ UserCLK Tile_X10Y15_S_term_IHP_SRAM/UserCLKo VGND VPWR S_term_IHP_SRAM
XTile_X2Y7_LUT4AB Tile_X2Y8_LUT4AB/Co Tile_X2Y7_LUT4AB/Co Tile_X3Y7_LUT4AB/E1END[0]
+ Tile_X3Y7_LUT4AB/E1END[1] Tile_X3Y7_LUT4AB/E1END[2] Tile_X3Y7_LUT4AB/E1END[3] Tile_X2Y7_LUT4AB/E1END[0]
+ Tile_X2Y7_LUT4AB/E1END[1] Tile_X2Y7_LUT4AB/E1END[2] Tile_X2Y7_LUT4AB/E1END[3] Tile_X3Y7_LUT4AB/E2MID[0]
+ Tile_X3Y7_LUT4AB/E2MID[1] Tile_X3Y7_LUT4AB/E2MID[2] Tile_X3Y7_LUT4AB/E2MID[3] Tile_X3Y7_LUT4AB/E2MID[4]
+ Tile_X3Y7_LUT4AB/E2MID[5] Tile_X3Y7_LUT4AB/E2MID[6] Tile_X3Y7_LUT4AB/E2MID[7] Tile_X3Y7_LUT4AB/E2END[0]
+ Tile_X3Y7_LUT4AB/E2END[1] Tile_X3Y7_LUT4AB/E2END[2] Tile_X3Y7_LUT4AB/E2END[3] Tile_X3Y7_LUT4AB/E2END[4]
+ Tile_X3Y7_LUT4AB/E2END[5] Tile_X3Y7_LUT4AB/E2END[6] Tile_X3Y7_LUT4AB/E2END[7] Tile_X2Y7_LUT4AB/E2END[0]
+ Tile_X2Y7_LUT4AB/E2END[1] Tile_X2Y7_LUT4AB/E2END[2] Tile_X2Y7_LUT4AB/E2END[3] Tile_X2Y7_LUT4AB/E2END[4]
+ Tile_X2Y7_LUT4AB/E2END[5] Tile_X2Y7_LUT4AB/E2END[6] Tile_X2Y7_LUT4AB/E2END[7] Tile_X2Y7_LUT4AB/E2MID[0]
+ Tile_X2Y7_LUT4AB/E2MID[1] Tile_X2Y7_LUT4AB/E2MID[2] Tile_X2Y7_LUT4AB/E2MID[3] Tile_X2Y7_LUT4AB/E2MID[4]
+ Tile_X2Y7_LUT4AB/E2MID[5] Tile_X2Y7_LUT4AB/E2MID[6] Tile_X2Y7_LUT4AB/E2MID[7] Tile_X3Y7_LUT4AB/E6END[0]
+ Tile_X3Y7_LUT4AB/E6END[10] Tile_X3Y7_LUT4AB/E6END[11] Tile_X3Y7_LUT4AB/E6END[1]
+ Tile_X3Y7_LUT4AB/E6END[2] Tile_X3Y7_LUT4AB/E6END[3] Tile_X3Y7_LUT4AB/E6END[4] Tile_X3Y7_LUT4AB/E6END[5]
+ Tile_X3Y7_LUT4AB/E6END[6] Tile_X3Y7_LUT4AB/E6END[7] Tile_X3Y7_LUT4AB/E6END[8] Tile_X3Y7_LUT4AB/E6END[9]
+ Tile_X2Y7_LUT4AB/E6END[0] Tile_X2Y7_LUT4AB/E6END[10] Tile_X2Y7_LUT4AB/E6END[11]
+ Tile_X2Y7_LUT4AB/E6END[1] Tile_X2Y7_LUT4AB/E6END[2] Tile_X2Y7_LUT4AB/E6END[3] Tile_X2Y7_LUT4AB/E6END[4]
+ Tile_X2Y7_LUT4AB/E6END[5] Tile_X2Y7_LUT4AB/E6END[6] Tile_X2Y7_LUT4AB/E6END[7] Tile_X2Y7_LUT4AB/E6END[8]
+ Tile_X2Y7_LUT4AB/E6END[9] Tile_X3Y7_LUT4AB/EE4END[0] Tile_X3Y7_LUT4AB/EE4END[10]
+ Tile_X3Y7_LUT4AB/EE4END[11] Tile_X3Y7_LUT4AB/EE4END[12] Tile_X3Y7_LUT4AB/EE4END[13]
+ Tile_X3Y7_LUT4AB/EE4END[14] Tile_X3Y7_LUT4AB/EE4END[15] Tile_X3Y7_LUT4AB/EE4END[1]
+ Tile_X3Y7_LUT4AB/EE4END[2] Tile_X3Y7_LUT4AB/EE4END[3] Tile_X3Y7_LUT4AB/EE4END[4]
+ Tile_X3Y7_LUT4AB/EE4END[5] Tile_X3Y7_LUT4AB/EE4END[6] Tile_X3Y7_LUT4AB/EE4END[7]
+ Tile_X3Y7_LUT4AB/EE4END[8] Tile_X3Y7_LUT4AB/EE4END[9] Tile_X2Y7_LUT4AB/EE4END[0]
+ Tile_X2Y7_LUT4AB/EE4END[10] Tile_X2Y7_LUT4AB/EE4END[11] Tile_X2Y7_LUT4AB/EE4END[12]
+ Tile_X2Y7_LUT4AB/EE4END[13] Tile_X2Y7_LUT4AB/EE4END[14] Tile_X2Y7_LUT4AB/EE4END[15]
+ Tile_X2Y7_LUT4AB/EE4END[1] Tile_X2Y7_LUT4AB/EE4END[2] Tile_X2Y7_LUT4AB/EE4END[3]
+ Tile_X2Y7_LUT4AB/EE4END[4] Tile_X2Y7_LUT4AB/EE4END[5] Tile_X2Y7_LUT4AB/EE4END[6]
+ Tile_X2Y7_LUT4AB/EE4END[7] Tile_X2Y7_LUT4AB/EE4END[8] Tile_X2Y7_LUT4AB/EE4END[9]
+ Tile_X2Y7_LUT4AB/FrameData[0] Tile_X2Y7_LUT4AB/FrameData[10] Tile_X2Y7_LUT4AB/FrameData[11]
+ Tile_X2Y7_LUT4AB/FrameData[12] Tile_X2Y7_LUT4AB/FrameData[13] Tile_X2Y7_LUT4AB/FrameData[14]
+ Tile_X2Y7_LUT4AB/FrameData[15] Tile_X2Y7_LUT4AB/FrameData[16] Tile_X2Y7_LUT4AB/FrameData[17]
+ Tile_X2Y7_LUT4AB/FrameData[18] Tile_X2Y7_LUT4AB/FrameData[19] Tile_X2Y7_LUT4AB/FrameData[1]
+ Tile_X2Y7_LUT4AB/FrameData[20] Tile_X2Y7_LUT4AB/FrameData[21] Tile_X2Y7_LUT4AB/FrameData[22]
+ Tile_X2Y7_LUT4AB/FrameData[23] Tile_X2Y7_LUT4AB/FrameData[24] Tile_X2Y7_LUT4AB/FrameData[25]
+ Tile_X2Y7_LUT4AB/FrameData[26] Tile_X2Y7_LUT4AB/FrameData[27] Tile_X2Y7_LUT4AB/FrameData[28]
+ Tile_X2Y7_LUT4AB/FrameData[29] Tile_X2Y7_LUT4AB/FrameData[2] Tile_X2Y7_LUT4AB/FrameData[30]
+ Tile_X2Y7_LUT4AB/FrameData[31] Tile_X2Y7_LUT4AB/FrameData[3] Tile_X2Y7_LUT4AB/FrameData[4]
+ Tile_X2Y7_LUT4AB/FrameData[5] Tile_X2Y7_LUT4AB/FrameData[6] Tile_X2Y7_LUT4AB/FrameData[7]
+ Tile_X2Y7_LUT4AB/FrameData[8] Tile_X2Y7_LUT4AB/FrameData[9] Tile_X3Y7_LUT4AB/FrameData[0]
+ Tile_X3Y7_LUT4AB/FrameData[10] Tile_X3Y7_LUT4AB/FrameData[11] Tile_X3Y7_LUT4AB/FrameData[12]
+ Tile_X3Y7_LUT4AB/FrameData[13] Tile_X3Y7_LUT4AB/FrameData[14] Tile_X3Y7_LUT4AB/FrameData[15]
+ Tile_X3Y7_LUT4AB/FrameData[16] Tile_X3Y7_LUT4AB/FrameData[17] Tile_X3Y7_LUT4AB/FrameData[18]
+ Tile_X3Y7_LUT4AB/FrameData[19] Tile_X3Y7_LUT4AB/FrameData[1] Tile_X3Y7_LUT4AB/FrameData[20]
+ Tile_X3Y7_LUT4AB/FrameData[21] Tile_X3Y7_LUT4AB/FrameData[22] Tile_X3Y7_LUT4AB/FrameData[23]
+ Tile_X3Y7_LUT4AB/FrameData[24] Tile_X3Y7_LUT4AB/FrameData[25] Tile_X3Y7_LUT4AB/FrameData[26]
+ Tile_X3Y7_LUT4AB/FrameData[27] Tile_X3Y7_LUT4AB/FrameData[28] Tile_X3Y7_LUT4AB/FrameData[29]
+ Tile_X3Y7_LUT4AB/FrameData[2] Tile_X3Y7_LUT4AB/FrameData[30] Tile_X3Y7_LUT4AB/FrameData[31]
+ Tile_X3Y7_LUT4AB/FrameData[3] Tile_X3Y7_LUT4AB/FrameData[4] Tile_X3Y7_LUT4AB/FrameData[5]
+ Tile_X3Y7_LUT4AB/FrameData[6] Tile_X3Y7_LUT4AB/FrameData[7] Tile_X3Y7_LUT4AB/FrameData[8]
+ Tile_X3Y7_LUT4AB/FrameData[9] Tile_X2Y7_LUT4AB/FrameStrobe[0] Tile_X2Y7_LUT4AB/FrameStrobe[10]
+ Tile_X2Y7_LUT4AB/FrameStrobe[11] Tile_X2Y7_LUT4AB/FrameStrobe[12] Tile_X2Y7_LUT4AB/FrameStrobe[13]
+ Tile_X2Y7_LUT4AB/FrameStrobe[14] Tile_X2Y7_LUT4AB/FrameStrobe[15] Tile_X2Y7_LUT4AB/FrameStrobe[16]
+ Tile_X2Y7_LUT4AB/FrameStrobe[17] Tile_X2Y7_LUT4AB/FrameStrobe[18] Tile_X2Y7_LUT4AB/FrameStrobe[19]
+ Tile_X2Y7_LUT4AB/FrameStrobe[1] Tile_X2Y7_LUT4AB/FrameStrobe[2] Tile_X2Y7_LUT4AB/FrameStrobe[3]
+ Tile_X2Y7_LUT4AB/FrameStrobe[4] Tile_X2Y7_LUT4AB/FrameStrobe[5] Tile_X2Y7_LUT4AB/FrameStrobe[6]
+ Tile_X2Y7_LUT4AB/FrameStrobe[7] Tile_X2Y7_LUT4AB/FrameStrobe[8] Tile_X2Y7_LUT4AB/FrameStrobe[9]
+ Tile_X2Y6_LUT4AB/FrameStrobe[0] Tile_X2Y6_LUT4AB/FrameStrobe[10] Tile_X2Y6_LUT4AB/FrameStrobe[11]
+ Tile_X2Y6_LUT4AB/FrameStrobe[12] Tile_X2Y6_LUT4AB/FrameStrobe[13] Tile_X2Y6_LUT4AB/FrameStrobe[14]
+ Tile_X2Y6_LUT4AB/FrameStrobe[15] Tile_X2Y6_LUT4AB/FrameStrobe[16] Tile_X2Y6_LUT4AB/FrameStrobe[17]
+ Tile_X2Y6_LUT4AB/FrameStrobe[18] Tile_X2Y6_LUT4AB/FrameStrobe[19] Tile_X2Y6_LUT4AB/FrameStrobe[1]
+ Tile_X2Y6_LUT4AB/FrameStrobe[2] Tile_X2Y6_LUT4AB/FrameStrobe[3] Tile_X2Y6_LUT4AB/FrameStrobe[4]
+ Tile_X2Y6_LUT4AB/FrameStrobe[5] Tile_X2Y6_LUT4AB/FrameStrobe[6] Tile_X2Y6_LUT4AB/FrameStrobe[7]
+ Tile_X2Y6_LUT4AB/FrameStrobe[8] Tile_X2Y6_LUT4AB/FrameStrobe[9] Tile_X2Y7_LUT4AB/N1BEG[0]
+ Tile_X2Y7_LUT4AB/N1BEG[1] Tile_X2Y7_LUT4AB/N1BEG[2] Tile_X2Y7_LUT4AB/N1BEG[3] Tile_X2Y8_LUT4AB/N1BEG[0]
+ Tile_X2Y8_LUT4AB/N1BEG[1] Tile_X2Y8_LUT4AB/N1BEG[2] Tile_X2Y8_LUT4AB/N1BEG[3] Tile_X2Y7_LUT4AB/N2BEG[0]
+ Tile_X2Y7_LUT4AB/N2BEG[1] Tile_X2Y7_LUT4AB/N2BEG[2] Tile_X2Y7_LUT4AB/N2BEG[3] Tile_X2Y7_LUT4AB/N2BEG[4]
+ Tile_X2Y7_LUT4AB/N2BEG[5] Tile_X2Y7_LUT4AB/N2BEG[6] Tile_X2Y7_LUT4AB/N2BEG[7] Tile_X2Y6_LUT4AB/N2END[0]
+ Tile_X2Y6_LUT4AB/N2END[1] Tile_X2Y6_LUT4AB/N2END[2] Tile_X2Y6_LUT4AB/N2END[3] Tile_X2Y6_LUT4AB/N2END[4]
+ Tile_X2Y6_LUT4AB/N2END[5] Tile_X2Y6_LUT4AB/N2END[6] Tile_X2Y6_LUT4AB/N2END[7] Tile_X2Y7_LUT4AB/N2END[0]
+ Tile_X2Y7_LUT4AB/N2END[1] Tile_X2Y7_LUT4AB/N2END[2] Tile_X2Y7_LUT4AB/N2END[3] Tile_X2Y7_LUT4AB/N2END[4]
+ Tile_X2Y7_LUT4AB/N2END[5] Tile_X2Y7_LUT4AB/N2END[6] Tile_X2Y7_LUT4AB/N2END[7] Tile_X2Y8_LUT4AB/N2BEG[0]
+ Tile_X2Y8_LUT4AB/N2BEG[1] Tile_X2Y8_LUT4AB/N2BEG[2] Tile_X2Y8_LUT4AB/N2BEG[3] Tile_X2Y8_LUT4AB/N2BEG[4]
+ Tile_X2Y8_LUT4AB/N2BEG[5] Tile_X2Y8_LUT4AB/N2BEG[6] Tile_X2Y8_LUT4AB/N2BEG[7] Tile_X2Y7_LUT4AB/N4BEG[0]
+ Tile_X2Y7_LUT4AB/N4BEG[10] Tile_X2Y7_LUT4AB/N4BEG[11] Tile_X2Y7_LUT4AB/N4BEG[12]
+ Tile_X2Y7_LUT4AB/N4BEG[13] Tile_X2Y7_LUT4AB/N4BEG[14] Tile_X2Y7_LUT4AB/N4BEG[15]
+ Tile_X2Y7_LUT4AB/N4BEG[1] Tile_X2Y7_LUT4AB/N4BEG[2] Tile_X2Y7_LUT4AB/N4BEG[3] Tile_X2Y7_LUT4AB/N4BEG[4]
+ Tile_X2Y7_LUT4AB/N4BEG[5] Tile_X2Y7_LUT4AB/N4BEG[6] Tile_X2Y7_LUT4AB/N4BEG[7] Tile_X2Y7_LUT4AB/N4BEG[8]
+ Tile_X2Y7_LUT4AB/N4BEG[9] Tile_X2Y8_LUT4AB/N4BEG[0] Tile_X2Y8_LUT4AB/N4BEG[10] Tile_X2Y8_LUT4AB/N4BEG[11]
+ Tile_X2Y8_LUT4AB/N4BEG[12] Tile_X2Y8_LUT4AB/N4BEG[13] Tile_X2Y8_LUT4AB/N4BEG[14]
+ Tile_X2Y8_LUT4AB/N4BEG[15] Tile_X2Y8_LUT4AB/N4BEG[1] Tile_X2Y8_LUT4AB/N4BEG[2] Tile_X2Y8_LUT4AB/N4BEG[3]
+ Tile_X2Y8_LUT4AB/N4BEG[4] Tile_X2Y8_LUT4AB/N4BEG[5] Tile_X2Y8_LUT4AB/N4BEG[6] Tile_X2Y8_LUT4AB/N4BEG[7]
+ Tile_X2Y8_LUT4AB/N4BEG[8] Tile_X2Y8_LUT4AB/N4BEG[9] Tile_X2Y7_LUT4AB/NN4BEG[0] Tile_X2Y7_LUT4AB/NN4BEG[10]
+ Tile_X2Y7_LUT4AB/NN4BEG[11] Tile_X2Y7_LUT4AB/NN4BEG[12] Tile_X2Y7_LUT4AB/NN4BEG[13]
+ Tile_X2Y7_LUT4AB/NN4BEG[14] Tile_X2Y7_LUT4AB/NN4BEG[15] Tile_X2Y7_LUT4AB/NN4BEG[1]
+ Tile_X2Y7_LUT4AB/NN4BEG[2] Tile_X2Y7_LUT4AB/NN4BEG[3] Tile_X2Y7_LUT4AB/NN4BEG[4]
+ Tile_X2Y7_LUT4AB/NN4BEG[5] Tile_X2Y7_LUT4AB/NN4BEG[6] Tile_X2Y7_LUT4AB/NN4BEG[7]
+ Tile_X2Y7_LUT4AB/NN4BEG[8] Tile_X2Y7_LUT4AB/NN4BEG[9] Tile_X2Y8_LUT4AB/NN4BEG[0]
+ Tile_X2Y8_LUT4AB/NN4BEG[10] Tile_X2Y8_LUT4AB/NN4BEG[11] Tile_X2Y8_LUT4AB/NN4BEG[12]
+ Tile_X2Y8_LUT4AB/NN4BEG[13] Tile_X2Y8_LUT4AB/NN4BEG[14] Tile_X2Y8_LUT4AB/NN4BEG[15]
+ Tile_X2Y8_LUT4AB/NN4BEG[1] Tile_X2Y8_LUT4AB/NN4BEG[2] Tile_X2Y8_LUT4AB/NN4BEG[3]
+ Tile_X2Y8_LUT4AB/NN4BEG[4] Tile_X2Y8_LUT4AB/NN4BEG[5] Tile_X2Y8_LUT4AB/NN4BEG[6]
+ Tile_X2Y8_LUT4AB/NN4BEG[7] Tile_X2Y8_LUT4AB/NN4BEG[8] Tile_X2Y8_LUT4AB/NN4BEG[9]
+ Tile_X2Y8_LUT4AB/S1END[0] Tile_X2Y8_LUT4AB/S1END[1] Tile_X2Y8_LUT4AB/S1END[2] Tile_X2Y8_LUT4AB/S1END[3]
+ Tile_X2Y7_LUT4AB/S1END[0] Tile_X2Y7_LUT4AB/S1END[1] Tile_X2Y7_LUT4AB/S1END[2] Tile_X2Y7_LUT4AB/S1END[3]
+ Tile_X2Y8_LUT4AB/S2MID[0] Tile_X2Y8_LUT4AB/S2MID[1] Tile_X2Y8_LUT4AB/S2MID[2] Tile_X2Y8_LUT4AB/S2MID[3]
+ Tile_X2Y8_LUT4AB/S2MID[4] Tile_X2Y8_LUT4AB/S2MID[5] Tile_X2Y8_LUT4AB/S2MID[6] Tile_X2Y8_LUT4AB/S2MID[7]
+ Tile_X2Y8_LUT4AB/S2END[0] Tile_X2Y8_LUT4AB/S2END[1] Tile_X2Y8_LUT4AB/S2END[2] Tile_X2Y8_LUT4AB/S2END[3]
+ Tile_X2Y8_LUT4AB/S2END[4] Tile_X2Y8_LUT4AB/S2END[5] Tile_X2Y8_LUT4AB/S2END[6] Tile_X2Y8_LUT4AB/S2END[7]
+ Tile_X2Y7_LUT4AB/S2END[0] Tile_X2Y7_LUT4AB/S2END[1] Tile_X2Y7_LUT4AB/S2END[2] Tile_X2Y7_LUT4AB/S2END[3]
+ Tile_X2Y7_LUT4AB/S2END[4] Tile_X2Y7_LUT4AB/S2END[5] Tile_X2Y7_LUT4AB/S2END[6] Tile_X2Y7_LUT4AB/S2END[7]
+ Tile_X2Y7_LUT4AB/S2MID[0] Tile_X2Y7_LUT4AB/S2MID[1] Tile_X2Y7_LUT4AB/S2MID[2] Tile_X2Y7_LUT4AB/S2MID[3]
+ Tile_X2Y7_LUT4AB/S2MID[4] Tile_X2Y7_LUT4AB/S2MID[5] Tile_X2Y7_LUT4AB/S2MID[6] Tile_X2Y7_LUT4AB/S2MID[7]
+ Tile_X2Y8_LUT4AB/S4END[0] Tile_X2Y8_LUT4AB/S4END[10] Tile_X2Y8_LUT4AB/S4END[11]
+ Tile_X2Y8_LUT4AB/S4END[12] Tile_X2Y8_LUT4AB/S4END[13] Tile_X2Y8_LUT4AB/S4END[14]
+ Tile_X2Y8_LUT4AB/S4END[15] Tile_X2Y8_LUT4AB/S4END[1] Tile_X2Y8_LUT4AB/S4END[2] Tile_X2Y8_LUT4AB/S4END[3]
+ Tile_X2Y8_LUT4AB/S4END[4] Tile_X2Y8_LUT4AB/S4END[5] Tile_X2Y8_LUT4AB/S4END[6] Tile_X2Y8_LUT4AB/S4END[7]
+ Tile_X2Y8_LUT4AB/S4END[8] Tile_X2Y8_LUT4AB/S4END[9] Tile_X2Y7_LUT4AB/S4END[0] Tile_X2Y7_LUT4AB/S4END[10]
+ Tile_X2Y7_LUT4AB/S4END[11] Tile_X2Y7_LUT4AB/S4END[12] Tile_X2Y7_LUT4AB/S4END[13]
+ Tile_X2Y7_LUT4AB/S4END[14] Tile_X2Y7_LUT4AB/S4END[15] Tile_X2Y7_LUT4AB/S4END[1]
+ Tile_X2Y7_LUT4AB/S4END[2] Tile_X2Y7_LUT4AB/S4END[3] Tile_X2Y7_LUT4AB/S4END[4] Tile_X2Y7_LUT4AB/S4END[5]
+ Tile_X2Y7_LUT4AB/S4END[6] Tile_X2Y7_LUT4AB/S4END[7] Tile_X2Y7_LUT4AB/S4END[8] Tile_X2Y7_LUT4AB/S4END[9]
+ Tile_X2Y8_LUT4AB/SS4END[0] Tile_X2Y8_LUT4AB/SS4END[10] Tile_X2Y8_LUT4AB/SS4END[11]
+ Tile_X2Y8_LUT4AB/SS4END[12] Tile_X2Y8_LUT4AB/SS4END[13] Tile_X2Y8_LUT4AB/SS4END[14]
+ Tile_X2Y8_LUT4AB/SS4END[15] Tile_X2Y8_LUT4AB/SS4END[1] Tile_X2Y8_LUT4AB/SS4END[2]
+ Tile_X2Y8_LUT4AB/SS4END[3] Tile_X2Y8_LUT4AB/SS4END[4] Tile_X2Y8_LUT4AB/SS4END[5]
+ Tile_X2Y8_LUT4AB/SS4END[6] Tile_X2Y8_LUT4AB/SS4END[7] Tile_X2Y8_LUT4AB/SS4END[8]
+ Tile_X2Y8_LUT4AB/SS4END[9] Tile_X2Y7_LUT4AB/SS4END[0] Tile_X2Y7_LUT4AB/SS4END[10]
+ Tile_X2Y7_LUT4AB/SS4END[11] Tile_X2Y7_LUT4AB/SS4END[12] Tile_X2Y7_LUT4AB/SS4END[13]
+ Tile_X2Y7_LUT4AB/SS4END[14] Tile_X2Y7_LUT4AB/SS4END[15] Tile_X2Y7_LUT4AB/SS4END[1]
+ Tile_X2Y7_LUT4AB/SS4END[2] Tile_X2Y7_LUT4AB/SS4END[3] Tile_X2Y7_LUT4AB/SS4END[4]
+ Tile_X2Y7_LUT4AB/SS4END[5] Tile_X2Y7_LUT4AB/SS4END[6] Tile_X2Y7_LUT4AB/SS4END[7]
+ Tile_X2Y7_LUT4AB/SS4END[8] Tile_X2Y7_LUT4AB/SS4END[9] Tile_X2Y7_LUT4AB/UserCLK Tile_X2Y6_LUT4AB/UserCLK
+ VGND VPWR Tile_X2Y7_LUT4AB/W1BEG[0] Tile_X2Y7_LUT4AB/W1BEG[1] Tile_X2Y7_LUT4AB/W1BEG[2]
+ Tile_X2Y7_LUT4AB/W1BEG[3] Tile_X3Y7_LUT4AB/W1BEG[0] Tile_X3Y7_LUT4AB/W1BEG[1] Tile_X3Y7_LUT4AB/W1BEG[2]
+ Tile_X3Y7_LUT4AB/W1BEG[3] Tile_X2Y7_LUT4AB/W2BEG[0] Tile_X2Y7_LUT4AB/W2BEG[1] Tile_X2Y7_LUT4AB/W2BEG[2]
+ Tile_X2Y7_LUT4AB/W2BEG[3] Tile_X2Y7_LUT4AB/W2BEG[4] Tile_X2Y7_LUT4AB/W2BEG[5] Tile_X2Y7_LUT4AB/W2BEG[6]
+ Tile_X2Y7_LUT4AB/W2BEG[7] Tile_X1Y7_LUT4AB/W2END[0] Tile_X1Y7_LUT4AB/W2END[1] Tile_X1Y7_LUT4AB/W2END[2]
+ Tile_X1Y7_LUT4AB/W2END[3] Tile_X1Y7_LUT4AB/W2END[4] Tile_X1Y7_LUT4AB/W2END[5] Tile_X1Y7_LUT4AB/W2END[6]
+ Tile_X1Y7_LUT4AB/W2END[7] Tile_X2Y7_LUT4AB/W2END[0] Tile_X2Y7_LUT4AB/W2END[1] Tile_X2Y7_LUT4AB/W2END[2]
+ Tile_X2Y7_LUT4AB/W2END[3] Tile_X2Y7_LUT4AB/W2END[4] Tile_X2Y7_LUT4AB/W2END[5] Tile_X2Y7_LUT4AB/W2END[6]
+ Tile_X2Y7_LUT4AB/W2END[7] Tile_X3Y7_LUT4AB/W2BEG[0] Tile_X3Y7_LUT4AB/W2BEG[1] Tile_X3Y7_LUT4AB/W2BEG[2]
+ Tile_X3Y7_LUT4AB/W2BEG[3] Tile_X3Y7_LUT4AB/W2BEG[4] Tile_X3Y7_LUT4AB/W2BEG[5] Tile_X3Y7_LUT4AB/W2BEG[6]
+ Tile_X3Y7_LUT4AB/W2BEG[7] Tile_X2Y7_LUT4AB/W6BEG[0] Tile_X2Y7_LUT4AB/W6BEG[10] Tile_X2Y7_LUT4AB/W6BEG[11]
+ Tile_X2Y7_LUT4AB/W6BEG[1] Tile_X2Y7_LUT4AB/W6BEG[2] Tile_X2Y7_LUT4AB/W6BEG[3] Tile_X2Y7_LUT4AB/W6BEG[4]
+ Tile_X2Y7_LUT4AB/W6BEG[5] Tile_X2Y7_LUT4AB/W6BEG[6] Tile_X2Y7_LUT4AB/W6BEG[7] Tile_X2Y7_LUT4AB/W6BEG[8]
+ Tile_X2Y7_LUT4AB/W6BEG[9] Tile_X3Y7_LUT4AB/W6BEG[0] Tile_X3Y7_LUT4AB/W6BEG[10] Tile_X3Y7_LUT4AB/W6BEG[11]
+ Tile_X3Y7_LUT4AB/W6BEG[1] Tile_X3Y7_LUT4AB/W6BEG[2] Tile_X3Y7_LUT4AB/W6BEG[3] Tile_X3Y7_LUT4AB/W6BEG[4]
+ Tile_X3Y7_LUT4AB/W6BEG[5] Tile_X3Y7_LUT4AB/W6BEG[6] Tile_X3Y7_LUT4AB/W6BEG[7] Tile_X3Y7_LUT4AB/W6BEG[8]
+ Tile_X3Y7_LUT4AB/W6BEG[9] Tile_X2Y7_LUT4AB/WW4BEG[0] Tile_X2Y7_LUT4AB/WW4BEG[10]
+ Tile_X2Y7_LUT4AB/WW4BEG[11] Tile_X2Y7_LUT4AB/WW4BEG[12] Tile_X2Y7_LUT4AB/WW4BEG[13]
+ Tile_X2Y7_LUT4AB/WW4BEG[14] Tile_X2Y7_LUT4AB/WW4BEG[15] Tile_X2Y7_LUT4AB/WW4BEG[1]
+ Tile_X2Y7_LUT4AB/WW4BEG[2] Tile_X2Y7_LUT4AB/WW4BEG[3] Tile_X2Y7_LUT4AB/WW4BEG[4]
+ Tile_X2Y7_LUT4AB/WW4BEG[5] Tile_X2Y7_LUT4AB/WW4BEG[6] Tile_X2Y7_LUT4AB/WW4BEG[7]
+ Tile_X2Y7_LUT4AB/WW4BEG[8] Tile_X2Y7_LUT4AB/WW4BEG[9] Tile_X3Y7_LUT4AB/WW4BEG[0]
+ Tile_X3Y7_LUT4AB/WW4BEG[10] Tile_X3Y7_LUT4AB/WW4BEG[11] Tile_X3Y7_LUT4AB/WW4BEG[12]
+ Tile_X3Y7_LUT4AB/WW4BEG[13] Tile_X3Y7_LUT4AB/WW4BEG[14] Tile_X3Y7_LUT4AB/WW4BEG[15]
+ Tile_X3Y7_LUT4AB/WW4BEG[1] Tile_X3Y7_LUT4AB/WW4BEG[2] Tile_X3Y7_LUT4AB/WW4BEG[3]
+ Tile_X3Y7_LUT4AB/WW4BEG[4] Tile_X3Y7_LUT4AB/WW4BEG[5] Tile_X3Y7_LUT4AB/WW4BEG[6]
+ Tile_X3Y7_LUT4AB/WW4BEG[7] Tile_X3Y7_LUT4AB/WW4BEG[8] Tile_X3Y7_LUT4AB/WW4BEG[9]
+ LUT4AB
XTile_X9Y2_LUT4AB Tile_X9Y3_LUT4AB/Co Tile_X9Y2_LUT4AB/Co Tile_X9Y2_LUT4AB/E1BEG[0]
+ Tile_X9Y2_LUT4AB/E1BEG[1] Tile_X9Y2_LUT4AB/E1BEG[2] Tile_X9Y2_LUT4AB/E1BEG[3] Tile_X9Y2_LUT4AB/E1END[0]
+ Tile_X9Y2_LUT4AB/E1END[1] Tile_X9Y2_LUT4AB/E1END[2] Tile_X9Y2_LUT4AB/E1END[3] Tile_X9Y2_LUT4AB/E2BEG[0]
+ Tile_X9Y2_LUT4AB/E2BEG[1] Tile_X9Y2_LUT4AB/E2BEG[2] Tile_X9Y2_LUT4AB/E2BEG[3] Tile_X9Y2_LUT4AB/E2BEG[4]
+ Tile_X9Y2_LUT4AB/E2BEG[5] Tile_X9Y2_LUT4AB/E2BEG[6] Tile_X9Y2_LUT4AB/E2BEG[7] Tile_X9Y2_LUT4AB/E2BEGb[0]
+ Tile_X9Y2_LUT4AB/E2BEGb[1] Tile_X9Y2_LUT4AB/E2BEGb[2] Tile_X9Y2_LUT4AB/E2BEGb[3]
+ Tile_X9Y2_LUT4AB/E2BEGb[4] Tile_X9Y2_LUT4AB/E2BEGb[5] Tile_X9Y2_LUT4AB/E2BEGb[6]
+ Tile_X9Y2_LUT4AB/E2BEGb[7] Tile_X9Y2_LUT4AB/E2END[0] Tile_X9Y2_LUT4AB/E2END[1] Tile_X9Y2_LUT4AB/E2END[2]
+ Tile_X9Y2_LUT4AB/E2END[3] Tile_X9Y2_LUT4AB/E2END[4] Tile_X9Y2_LUT4AB/E2END[5] Tile_X9Y2_LUT4AB/E2END[6]
+ Tile_X9Y2_LUT4AB/E2END[7] Tile_X9Y2_LUT4AB/E2MID[0] Tile_X9Y2_LUT4AB/E2MID[1] Tile_X9Y2_LUT4AB/E2MID[2]
+ Tile_X9Y2_LUT4AB/E2MID[3] Tile_X9Y2_LUT4AB/E2MID[4] Tile_X9Y2_LUT4AB/E2MID[5] Tile_X9Y2_LUT4AB/E2MID[6]
+ Tile_X9Y2_LUT4AB/E2MID[7] Tile_X9Y2_LUT4AB/E6BEG[0] Tile_X9Y2_LUT4AB/E6BEG[10] Tile_X9Y2_LUT4AB/E6BEG[11]
+ Tile_X9Y2_LUT4AB/E6BEG[1] Tile_X9Y2_LUT4AB/E6BEG[2] Tile_X9Y2_LUT4AB/E6BEG[3] Tile_X9Y2_LUT4AB/E6BEG[4]
+ Tile_X9Y2_LUT4AB/E6BEG[5] Tile_X9Y2_LUT4AB/E6BEG[6] Tile_X9Y2_LUT4AB/E6BEG[7] Tile_X9Y2_LUT4AB/E6BEG[8]
+ Tile_X9Y2_LUT4AB/E6BEG[9] Tile_X9Y2_LUT4AB/E6END[0] Tile_X9Y2_LUT4AB/E6END[10] Tile_X9Y2_LUT4AB/E6END[11]
+ Tile_X9Y2_LUT4AB/E6END[1] Tile_X9Y2_LUT4AB/E6END[2] Tile_X9Y2_LUT4AB/E6END[3] Tile_X9Y2_LUT4AB/E6END[4]
+ Tile_X9Y2_LUT4AB/E6END[5] Tile_X9Y2_LUT4AB/E6END[6] Tile_X9Y2_LUT4AB/E6END[7] Tile_X9Y2_LUT4AB/E6END[8]
+ Tile_X9Y2_LUT4AB/E6END[9] Tile_X9Y2_LUT4AB/EE4BEG[0] Tile_X9Y2_LUT4AB/EE4BEG[10]
+ Tile_X9Y2_LUT4AB/EE4BEG[11] Tile_X9Y2_LUT4AB/EE4BEG[12] Tile_X9Y2_LUT4AB/EE4BEG[13]
+ Tile_X9Y2_LUT4AB/EE4BEG[14] Tile_X9Y2_LUT4AB/EE4BEG[15] Tile_X9Y2_LUT4AB/EE4BEG[1]
+ Tile_X9Y2_LUT4AB/EE4BEG[2] Tile_X9Y2_LUT4AB/EE4BEG[3] Tile_X9Y2_LUT4AB/EE4BEG[4]
+ Tile_X9Y2_LUT4AB/EE4BEG[5] Tile_X9Y2_LUT4AB/EE4BEG[6] Tile_X9Y2_LUT4AB/EE4BEG[7]
+ Tile_X9Y2_LUT4AB/EE4BEG[8] Tile_X9Y2_LUT4AB/EE4BEG[9] Tile_X9Y2_LUT4AB/EE4END[0]
+ Tile_X9Y2_LUT4AB/EE4END[10] Tile_X9Y2_LUT4AB/EE4END[11] Tile_X9Y2_LUT4AB/EE4END[12]
+ Tile_X9Y2_LUT4AB/EE4END[13] Tile_X9Y2_LUT4AB/EE4END[14] Tile_X9Y2_LUT4AB/EE4END[15]
+ Tile_X9Y2_LUT4AB/EE4END[1] Tile_X9Y2_LUT4AB/EE4END[2] Tile_X9Y2_LUT4AB/EE4END[3]
+ Tile_X9Y2_LUT4AB/EE4END[4] Tile_X9Y2_LUT4AB/EE4END[5] Tile_X9Y2_LUT4AB/EE4END[6]
+ Tile_X9Y2_LUT4AB/EE4END[7] Tile_X9Y2_LUT4AB/EE4END[8] Tile_X9Y2_LUT4AB/EE4END[9]
+ Tile_X9Y2_LUT4AB/FrameData[0] Tile_X9Y2_LUT4AB/FrameData[10] Tile_X9Y2_LUT4AB/FrameData[11]
+ Tile_X9Y2_LUT4AB/FrameData[12] Tile_X9Y2_LUT4AB/FrameData[13] Tile_X9Y2_LUT4AB/FrameData[14]
+ Tile_X9Y2_LUT4AB/FrameData[15] Tile_X9Y2_LUT4AB/FrameData[16] Tile_X9Y2_LUT4AB/FrameData[17]
+ Tile_X9Y2_LUT4AB/FrameData[18] Tile_X9Y2_LUT4AB/FrameData[19] Tile_X9Y2_LUT4AB/FrameData[1]
+ Tile_X9Y2_LUT4AB/FrameData[20] Tile_X9Y2_LUT4AB/FrameData[21] Tile_X9Y2_LUT4AB/FrameData[22]
+ Tile_X9Y2_LUT4AB/FrameData[23] Tile_X9Y2_LUT4AB/FrameData[24] Tile_X9Y2_LUT4AB/FrameData[25]
+ Tile_X9Y2_LUT4AB/FrameData[26] Tile_X9Y2_LUT4AB/FrameData[27] Tile_X9Y2_LUT4AB/FrameData[28]
+ Tile_X9Y2_LUT4AB/FrameData[29] Tile_X9Y2_LUT4AB/FrameData[2] Tile_X9Y2_LUT4AB/FrameData[30]
+ Tile_X9Y2_LUT4AB/FrameData[31] Tile_X9Y2_LUT4AB/FrameData[3] Tile_X9Y2_LUT4AB/FrameData[4]
+ Tile_X9Y2_LUT4AB/FrameData[5] Tile_X9Y2_LUT4AB/FrameData[6] Tile_X9Y2_LUT4AB/FrameData[7]
+ Tile_X9Y2_LUT4AB/FrameData[8] Tile_X9Y2_LUT4AB/FrameData[9] Tile_X9Y2_LUT4AB/FrameData_O[0]
+ Tile_X9Y2_LUT4AB/FrameData_O[10] Tile_X9Y2_LUT4AB/FrameData_O[11] Tile_X9Y2_LUT4AB/FrameData_O[12]
+ Tile_X9Y2_LUT4AB/FrameData_O[13] Tile_X9Y2_LUT4AB/FrameData_O[14] Tile_X9Y2_LUT4AB/FrameData_O[15]
+ Tile_X9Y2_LUT4AB/FrameData_O[16] Tile_X9Y2_LUT4AB/FrameData_O[17] Tile_X9Y2_LUT4AB/FrameData_O[18]
+ Tile_X9Y2_LUT4AB/FrameData_O[19] Tile_X9Y2_LUT4AB/FrameData_O[1] Tile_X9Y2_LUT4AB/FrameData_O[20]
+ Tile_X9Y2_LUT4AB/FrameData_O[21] Tile_X9Y2_LUT4AB/FrameData_O[22] Tile_X9Y2_LUT4AB/FrameData_O[23]
+ Tile_X9Y2_LUT4AB/FrameData_O[24] Tile_X9Y2_LUT4AB/FrameData_O[25] Tile_X9Y2_LUT4AB/FrameData_O[26]
+ Tile_X9Y2_LUT4AB/FrameData_O[27] Tile_X9Y2_LUT4AB/FrameData_O[28] Tile_X9Y2_LUT4AB/FrameData_O[29]
+ Tile_X9Y2_LUT4AB/FrameData_O[2] Tile_X9Y2_LUT4AB/FrameData_O[30] Tile_X9Y2_LUT4AB/FrameData_O[31]
+ Tile_X9Y2_LUT4AB/FrameData_O[3] Tile_X9Y2_LUT4AB/FrameData_O[4] Tile_X9Y2_LUT4AB/FrameData_O[5]
+ Tile_X9Y2_LUT4AB/FrameData_O[6] Tile_X9Y2_LUT4AB/FrameData_O[7] Tile_X9Y2_LUT4AB/FrameData_O[8]
+ Tile_X9Y2_LUT4AB/FrameData_O[9] Tile_X9Y2_LUT4AB/FrameStrobe[0] Tile_X9Y2_LUT4AB/FrameStrobe[10]
+ Tile_X9Y2_LUT4AB/FrameStrobe[11] Tile_X9Y2_LUT4AB/FrameStrobe[12] Tile_X9Y2_LUT4AB/FrameStrobe[13]
+ Tile_X9Y2_LUT4AB/FrameStrobe[14] Tile_X9Y2_LUT4AB/FrameStrobe[15] Tile_X9Y2_LUT4AB/FrameStrobe[16]
+ Tile_X9Y2_LUT4AB/FrameStrobe[17] Tile_X9Y2_LUT4AB/FrameStrobe[18] Tile_X9Y2_LUT4AB/FrameStrobe[19]
+ Tile_X9Y2_LUT4AB/FrameStrobe[1] Tile_X9Y2_LUT4AB/FrameStrobe[2] Tile_X9Y2_LUT4AB/FrameStrobe[3]
+ Tile_X9Y2_LUT4AB/FrameStrobe[4] Tile_X9Y2_LUT4AB/FrameStrobe[5] Tile_X9Y2_LUT4AB/FrameStrobe[6]
+ Tile_X9Y2_LUT4AB/FrameStrobe[7] Tile_X9Y2_LUT4AB/FrameStrobe[8] Tile_X9Y2_LUT4AB/FrameStrobe[9]
+ Tile_X9Y1_LUT4AB/FrameStrobe[0] Tile_X9Y1_LUT4AB/FrameStrobe[10] Tile_X9Y1_LUT4AB/FrameStrobe[11]
+ Tile_X9Y1_LUT4AB/FrameStrobe[12] Tile_X9Y1_LUT4AB/FrameStrobe[13] Tile_X9Y1_LUT4AB/FrameStrobe[14]
+ Tile_X9Y1_LUT4AB/FrameStrobe[15] Tile_X9Y1_LUT4AB/FrameStrobe[16] Tile_X9Y1_LUT4AB/FrameStrobe[17]
+ Tile_X9Y1_LUT4AB/FrameStrobe[18] Tile_X9Y1_LUT4AB/FrameStrobe[19] Tile_X9Y1_LUT4AB/FrameStrobe[1]
+ Tile_X9Y1_LUT4AB/FrameStrobe[2] Tile_X9Y1_LUT4AB/FrameStrobe[3] Tile_X9Y1_LUT4AB/FrameStrobe[4]
+ Tile_X9Y1_LUT4AB/FrameStrobe[5] Tile_X9Y1_LUT4AB/FrameStrobe[6] Tile_X9Y1_LUT4AB/FrameStrobe[7]
+ Tile_X9Y1_LUT4AB/FrameStrobe[8] Tile_X9Y1_LUT4AB/FrameStrobe[9] Tile_X9Y2_LUT4AB/N1BEG[0]
+ Tile_X9Y2_LUT4AB/N1BEG[1] Tile_X9Y2_LUT4AB/N1BEG[2] Tile_X9Y2_LUT4AB/N1BEG[3] Tile_X9Y3_LUT4AB/N1BEG[0]
+ Tile_X9Y3_LUT4AB/N1BEG[1] Tile_X9Y3_LUT4AB/N1BEG[2] Tile_X9Y3_LUT4AB/N1BEG[3] Tile_X9Y2_LUT4AB/N2BEG[0]
+ Tile_X9Y2_LUT4AB/N2BEG[1] Tile_X9Y2_LUT4AB/N2BEG[2] Tile_X9Y2_LUT4AB/N2BEG[3] Tile_X9Y2_LUT4AB/N2BEG[4]
+ Tile_X9Y2_LUT4AB/N2BEG[5] Tile_X9Y2_LUT4AB/N2BEG[6] Tile_X9Y2_LUT4AB/N2BEG[7] Tile_X9Y1_LUT4AB/N2END[0]
+ Tile_X9Y1_LUT4AB/N2END[1] Tile_X9Y1_LUT4AB/N2END[2] Tile_X9Y1_LUT4AB/N2END[3] Tile_X9Y1_LUT4AB/N2END[4]
+ Tile_X9Y1_LUT4AB/N2END[5] Tile_X9Y1_LUT4AB/N2END[6] Tile_X9Y1_LUT4AB/N2END[7] Tile_X9Y2_LUT4AB/N2END[0]
+ Tile_X9Y2_LUT4AB/N2END[1] Tile_X9Y2_LUT4AB/N2END[2] Tile_X9Y2_LUT4AB/N2END[3] Tile_X9Y2_LUT4AB/N2END[4]
+ Tile_X9Y2_LUT4AB/N2END[5] Tile_X9Y2_LUT4AB/N2END[6] Tile_X9Y2_LUT4AB/N2END[7] Tile_X9Y3_LUT4AB/N2BEG[0]
+ Tile_X9Y3_LUT4AB/N2BEG[1] Tile_X9Y3_LUT4AB/N2BEG[2] Tile_X9Y3_LUT4AB/N2BEG[3] Tile_X9Y3_LUT4AB/N2BEG[4]
+ Tile_X9Y3_LUT4AB/N2BEG[5] Tile_X9Y3_LUT4AB/N2BEG[6] Tile_X9Y3_LUT4AB/N2BEG[7] Tile_X9Y2_LUT4AB/N4BEG[0]
+ Tile_X9Y2_LUT4AB/N4BEG[10] Tile_X9Y2_LUT4AB/N4BEG[11] Tile_X9Y2_LUT4AB/N4BEG[12]
+ Tile_X9Y2_LUT4AB/N4BEG[13] Tile_X9Y2_LUT4AB/N4BEG[14] Tile_X9Y2_LUT4AB/N4BEG[15]
+ Tile_X9Y2_LUT4AB/N4BEG[1] Tile_X9Y2_LUT4AB/N4BEG[2] Tile_X9Y2_LUT4AB/N4BEG[3] Tile_X9Y2_LUT4AB/N4BEG[4]
+ Tile_X9Y2_LUT4AB/N4BEG[5] Tile_X9Y2_LUT4AB/N4BEG[6] Tile_X9Y2_LUT4AB/N4BEG[7] Tile_X9Y2_LUT4AB/N4BEG[8]
+ Tile_X9Y2_LUT4AB/N4BEG[9] Tile_X9Y3_LUT4AB/N4BEG[0] Tile_X9Y3_LUT4AB/N4BEG[10] Tile_X9Y3_LUT4AB/N4BEG[11]
+ Tile_X9Y3_LUT4AB/N4BEG[12] Tile_X9Y3_LUT4AB/N4BEG[13] Tile_X9Y3_LUT4AB/N4BEG[14]
+ Tile_X9Y3_LUT4AB/N4BEG[15] Tile_X9Y3_LUT4AB/N4BEG[1] Tile_X9Y3_LUT4AB/N4BEG[2] Tile_X9Y3_LUT4AB/N4BEG[3]
+ Tile_X9Y3_LUT4AB/N4BEG[4] Tile_X9Y3_LUT4AB/N4BEG[5] Tile_X9Y3_LUT4AB/N4BEG[6] Tile_X9Y3_LUT4AB/N4BEG[7]
+ Tile_X9Y3_LUT4AB/N4BEG[8] Tile_X9Y3_LUT4AB/N4BEG[9] Tile_X9Y2_LUT4AB/NN4BEG[0] Tile_X9Y2_LUT4AB/NN4BEG[10]
+ Tile_X9Y2_LUT4AB/NN4BEG[11] Tile_X9Y2_LUT4AB/NN4BEG[12] Tile_X9Y2_LUT4AB/NN4BEG[13]
+ Tile_X9Y2_LUT4AB/NN4BEG[14] Tile_X9Y2_LUT4AB/NN4BEG[15] Tile_X9Y2_LUT4AB/NN4BEG[1]
+ Tile_X9Y2_LUT4AB/NN4BEG[2] Tile_X9Y2_LUT4AB/NN4BEG[3] Tile_X9Y2_LUT4AB/NN4BEG[4]
+ Tile_X9Y2_LUT4AB/NN4BEG[5] Tile_X9Y2_LUT4AB/NN4BEG[6] Tile_X9Y2_LUT4AB/NN4BEG[7]
+ Tile_X9Y2_LUT4AB/NN4BEG[8] Tile_X9Y2_LUT4AB/NN4BEG[9] Tile_X9Y3_LUT4AB/NN4BEG[0]
+ Tile_X9Y3_LUT4AB/NN4BEG[10] Tile_X9Y3_LUT4AB/NN4BEG[11] Tile_X9Y3_LUT4AB/NN4BEG[12]
+ Tile_X9Y3_LUT4AB/NN4BEG[13] Tile_X9Y3_LUT4AB/NN4BEG[14] Tile_X9Y3_LUT4AB/NN4BEG[15]
+ Tile_X9Y3_LUT4AB/NN4BEG[1] Tile_X9Y3_LUT4AB/NN4BEG[2] Tile_X9Y3_LUT4AB/NN4BEG[3]
+ Tile_X9Y3_LUT4AB/NN4BEG[4] Tile_X9Y3_LUT4AB/NN4BEG[5] Tile_X9Y3_LUT4AB/NN4BEG[6]
+ Tile_X9Y3_LUT4AB/NN4BEG[7] Tile_X9Y3_LUT4AB/NN4BEG[8] Tile_X9Y3_LUT4AB/NN4BEG[9]
+ Tile_X9Y3_LUT4AB/S1END[0] Tile_X9Y3_LUT4AB/S1END[1] Tile_X9Y3_LUT4AB/S1END[2] Tile_X9Y3_LUT4AB/S1END[3]
+ Tile_X9Y2_LUT4AB/S1END[0] Tile_X9Y2_LUT4AB/S1END[1] Tile_X9Y2_LUT4AB/S1END[2] Tile_X9Y2_LUT4AB/S1END[3]
+ Tile_X9Y3_LUT4AB/S2MID[0] Tile_X9Y3_LUT4AB/S2MID[1] Tile_X9Y3_LUT4AB/S2MID[2] Tile_X9Y3_LUT4AB/S2MID[3]
+ Tile_X9Y3_LUT4AB/S2MID[4] Tile_X9Y3_LUT4AB/S2MID[5] Tile_X9Y3_LUT4AB/S2MID[6] Tile_X9Y3_LUT4AB/S2MID[7]
+ Tile_X9Y3_LUT4AB/S2END[0] Tile_X9Y3_LUT4AB/S2END[1] Tile_X9Y3_LUT4AB/S2END[2] Tile_X9Y3_LUT4AB/S2END[3]
+ Tile_X9Y3_LUT4AB/S2END[4] Tile_X9Y3_LUT4AB/S2END[5] Tile_X9Y3_LUT4AB/S2END[6] Tile_X9Y3_LUT4AB/S2END[7]
+ Tile_X9Y2_LUT4AB/S2END[0] Tile_X9Y2_LUT4AB/S2END[1] Tile_X9Y2_LUT4AB/S2END[2] Tile_X9Y2_LUT4AB/S2END[3]
+ Tile_X9Y2_LUT4AB/S2END[4] Tile_X9Y2_LUT4AB/S2END[5] Tile_X9Y2_LUT4AB/S2END[6] Tile_X9Y2_LUT4AB/S2END[7]
+ Tile_X9Y2_LUT4AB/S2MID[0] Tile_X9Y2_LUT4AB/S2MID[1] Tile_X9Y2_LUT4AB/S2MID[2] Tile_X9Y2_LUT4AB/S2MID[3]
+ Tile_X9Y2_LUT4AB/S2MID[4] Tile_X9Y2_LUT4AB/S2MID[5] Tile_X9Y2_LUT4AB/S2MID[6] Tile_X9Y2_LUT4AB/S2MID[7]
+ Tile_X9Y3_LUT4AB/S4END[0] Tile_X9Y3_LUT4AB/S4END[10] Tile_X9Y3_LUT4AB/S4END[11]
+ Tile_X9Y3_LUT4AB/S4END[12] Tile_X9Y3_LUT4AB/S4END[13] Tile_X9Y3_LUT4AB/S4END[14]
+ Tile_X9Y3_LUT4AB/S4END[15] Tile_X9Y3_LUT4AB/S4END[1] Tile_X9Y3_LUT4AB/S4END[2] Tile_X9Y3_LUT4AB/S4END[3]
+ Tile_X9Y3_LUT4AB/S4END[4] Tile_X9Y3_LUT4AB/S4END[5] Tile_X9Y3_LUT4AB/S4END[6] Tile_X9Y3_LUT4AB/S4END[7]
+ Tile_X9Y3_LUT4AB/S4END[8] Tile_X9Y3_LUT4AB/S4END[9] Tile_X9Y2_LUT4AB/S4END[0] Tile_X9Y2_LUT4AB/S4END[10]
+ Tile_X9Y2_LUT4AB/S4END[11] Tile_X9Y2_LUT4AB/S4END[12] Tile_X9Y2_LUT4AB/S4END[13]
+ Tile_X9Y2_LUT4AB/S4END[14] Tile_X9Y2_LUT4AB/S4END[15] Tile_X9Y2_LUT4AB/S4END[1]
+ Tile_X9Y2_LUT4AB/S4END[2] Tile_X9Y2_LUT4AB/S4END[3] Tile_X9Y2_LUT4AB/S4END[4] Tile_X9Y2_LUT4AB/S4END[5]
+ Tile_X9Y2_LUT4AB/S4END[6] Tile_X9Y2_LUT4AB/S4END[7] Tile_X9Y2_LUT4AB/S4END[8] Tile_X9Y2_LUT4AB/S4END[9]
+ Tile_X9Y3_LUT4AB/SS4END[0] Tile_X9Y3_LUT4AB/SS4END[10] Tile_X9Y3_LUT4AB/SS4END[11]
+ Tile_X9Y3_LUT4AB/SS4END[12] Tile_X9Y3_LUT4AB/SS4END[13] Tile_X9Y3_LUT4AB/SS4END[14]
+ Tile_X9Y3_LUT4AB/SS4END[15] Tile_X9Y3_LUT4AB/SS4END[1] Tile_X9Y3_LUT4AB/SS4END[2]
+ Tile_X9Y3_LUT4AB/SS4END[3] Tile_X9Y3_LUT4AB/SS4END[4] Tile_X9Y3_LUT4AB/SS4END[5]
+ Tile_X9Y3_LUT4AB/SS4END[6] Tile_X9Y3_LUT4AB/SS4END[7] Tile_X9Y3_LUT4AB/SS4END[8]
+ Tile_X9Y3_LUT4AB/SS4END[9] Tile_X9Y2_LUT4AB/SS4END[0] Tile_X9Y2_LUT4AB/SS4END[10]
+ Tile_X9Y2_LUT4AB/SS4END[11] Tile_X9Y2_LUT4AB/SS4END[12] Tile_X9Y2_LUT4AB/SS4END[13]
+ Tile_X9Y2_LUT4AB/SS4END[14] Tile_X9Y2_LUT4AB/SS4END[15] Tile_X9Y2_LUT4AB/SS4END[1]
+ Tile_X9Y2_LUT4AB/SS4END[2] Tile_X9Y2_LUT4AB/SS4END[3] Tile_X9Y2_LUT4AB/SS4END[4]
+ Tile_X9Y2_LUT4AB/SS4END[5] Tile_X9Y2_LUT4AB/SS4END[6] Tile_X9Y2_LUT4AB/SS4END[7]
+ Tile_X9Y2_LUT4AB/SS4END[8] Tile_X9Y2_LUT4AB/SS4END[9] Tile_X9Y2_LUT4AB/UserCLK Tile_X9Y1_LUT4AB/UserCLK
+ VGND VPWR Tile_X9Y2_LUT4AB/W1BEG[0] Tile_X9Y2_LUT4AB/W1BEG[1] Tile_X9Y2_LUT4AB/W1BEG[2]
+ Tile_X9Y2_LUT4AB/W1BEG[3] Tile_X9Y2_LUT4AB/W1END[0] Tile_X9Y2_LUT4AB/W1END[1] Tile_X9Y2_LUT4AB/W1END[2]
+ Tile_X9Y2_LUT4AB/W1END[3] Tile_X9Y2_LUT4AB/W2BEG[0] Tile_X9Y2_LUT4AB/W2BEG[1] Tile_X9Y2_LUT4AB/W2BEG[2]
+ Tile_X9Y2_LUT4AB/W2BEG[3] Tile_X9Y2_LUT4AB/W2BEG[4] Tile_X9Y2_LUT4AB/W2BEG[5] Tile_X9Y2_LUT4AB/W2BEG[6]
+ Tile_X9Y2_LUT4AB/W2BEG[7] Tile_X8Y2_LUT4AB/W2END[0] Tile_X8Y2_LUT4AB/W2END[1] Tile_X8Y2_LUT4AB/W2END[2]
+ Tile_X8Y2_LUT4AB/W2END[3] Tile_X8Y2_LUT4AB/W2END[4] Tile_X8Y2_LUT4AB/W2END[5] Tile_X8Y2_LUT4AB/W2END[6]
+ Tile_X8Y2_LUT4AB/W2END[7] Tile_X9Y2_LUT4AB/W2END[0] Tile_X9Y2_LUT4AB/W2END[1] Tile_X9Y2_LUT4AB/W2END[2]
+ Tile_X9Y2_LUT4AB/W2END[3] Tile_X9Y2_LUT4AB/W2END[4] Tile_X9Y2_LUT4AB/W2END[5] Tile_X9Y2_LUT4AB/W2END[6]
+ Tile_X9Y2_LUT4AB/W2END[7] Tile_X9Y2_LUT4AB/W2MID[0] Tile_X9Y2_LUT4AB/W2MID[1] Tile_X9Y2_LUT4AB/W2MID[2]
+ Tile_X9Y2_LUT4AB/W2MID[3] Tile_X9Y2_LUT4AB/W2MID[4] Tile_X9Y2_LUT4AB/W2MID[5] Tile_X9Y2_LUT4AB/W2MID[6]
+ Tile_X9Y2_LUT4AB/W2MID[7] Tile_X9Y2_LUT4AB/W6BEG[0] Tile_X9Y2_LUT4AB/W6BEG[10] Tile_X9Y2_LUT4AB/W6BEG[11]
+ Tile_X9Y2_LUT4AB/W6BEG[1] Tile_X9Y2_LUT4AB/W6BEG[2] Tile_X9Y2_LUT4AB/W6BEG[3] Tile_X9Y2_LUT4AB/W6BEG[4]
+ Tile_X9Y2_LUT4AB/W6BEG[5] Tile_X9Y2_LUT4AB/W6BEG[6] Tile_X9Y2_LUT4AB/W6BEG[7] Tile_X9Y2_LUT4AB/W6BEG[8]
+ Tile_X9Y2_LUT4AB/W6BEG[9] Tile_X9Y2_LUT4AB/W6END[0] Tile_X9Y2_LUT4AB/W6END[10] Tile_X9Y2_LUT4AB/W6END[11]
+ Tile_X9Y2_LUT4AB/W6END[1] Tile_X9Y2_LUT4AB/W6END[2] Tile_X9Y2_LUT4AB/W6END[3] Tile_X9Y2_LUT4AB/W6END[4]
+ Tile_X9Y2_LUT4AB/W6END[5] Tile_X9Y2_LUT4AB/W6END[6] Tile_X9Y2_LUT4AB/W6END[7] Tile_X9Y2_LUT4AB/W6END[8]
+ Tile_X9Y2_LUT4AB/W6END[9] Tile_X9Y2_LUT4AB/WW4BEG[0] Tile_X9Y2_LUT4AB/WW4BEG[10]
+ Tile_X9Y2_LUT4AB/WW4BEG[11] Tile_X9Y2_LUT4AB/WW4BEG[12] Tile_X9Y2_LUT4AB/WW4BEG[13]
+ Tile_X9Y2_LUT4AB/WW4BEG[14] Tile_X9Y2_LUT4AB/WW4BEG[15] Tile_X9Y2_LUT4AB/WW4BEG[1]
+ Tile_X9Y2_LUT4AB/WW4BEG[2] Tile_X9Y2_LUT4AB/WW4BEG[3] Tile_X9Y2_LUT4AB/WW4BEG[4]
+ Tile_X9Y2_LUT4AB/WW4BEG[5] Tile_X9Y2_LUT4AB/WW4BEG[6] Tile_X9Y2_LUT4AB/WW4BEG[7]
+ Tile_X9Y2_LUT4AB/WW4BEG[8] Tile_X9Y2_LUT4AB/WW4BEG[9] Tile_X9Y2_LUT4AB/WW4END[0]
+ Tile_X9Y2_LUT4AB/WW4END[10] Tile_X9Y2_LUT4AB/WW4END[11] Tile_X9Y2_LUT4AB/WW4END[12]
+ Tile_X9Y2_LUT4AB/WW4END[13] Tile_X9Y2_LUT4AB/WW4END[14] Tile_X9Y2_LUT4AB/WW4END[15]
+ Tile_X9Y2_LUT4AB/WW4END[1] Tile_X9Y2_LUT4AB/WW4END[2] Tile_X9Y2_LUT4AB/WW4END[3]
+ Tile_X9Y2_LUT4AB/WW4END[4] Tile_X9Y2_LUT4AB/WW4END[5] Tile_X9Y2_LUT4AB/WW4END[6]
+ Tile_X9Y2_LUT4AB/WW4END[7] Tile_X9Y2_LUT4AB/WW4END[8] Tile_X9Y2_LUT4AB/WW4END[9]
+ LUT4AB
XTile_X5Y13_LUT4AB Tile_X5Y14_LUT4AB/Co Tile_X5Y13_LUT4AB/Co Tile_X6Y13_LUT4AB/E1END[0]
+ Tile_X6Y13_LUT4AB/E1END[1] Tile_X6Y13_LUT4AB/E1END[2] Tile_X6Y13_LUT4AB/E1END[3]
+ Tile_X5Y13_LUT4AB/E1END[0] Tile_X5Y13_LUT4AB/E1END[1] Tile_X5Y13_LUT4AB/E1END[2]
+ Tile_X5Y13_LUT4AB/E1END[3] Tile_X6Y13_LUT4AB/E2MID[0] Tile_X6Y13_LUT4AB/E2MID[1]
+ Tile_X6Y13_LUT4AB/E2MID[2] Tile_X6Y13_LUT4AB/E2MID[3] Tile_X6Y13_LUT4AB/E2MID[4]
+ Tile_X6Y13_LUT4AB/E2MID[5] Tile_X6Y13_LUT4AB/E2MID[6] Tile_X6Y13_LUT4AB/E2MID[7]
+ Tile_X6Y13_LUT4AB/E2END[0] Tile_X6Y13_LUT4AB/E2END[1] Tile_X6Y13_LUT4AB/E2END[2]
+ Tile_X6Y13_LUT4AB/E2END[3] Tile_X6Y13_LUT4AB/E2END[4] Tile_X6Y13_LUT4AB/E2END[5]
+ Tile_X6Y13_LUT4AB/E2END[6] Tile_X6Y13_LUT4AB/E2END[7] Tile_X5Y13_LUT4AB/E2END[0]
+ Tile_X5Y13_LUT4AB/E2END[1] Tile_X5Y13_LUT4AB/E2END[2] Tile_X5Y13_LUT4AB/E2END[3]
+ Tile_X5Y13_LUT4AB/E2END[4] Tile_X5Y13_LUT4AB/E2END[5] Tile_X5Y13_LUT4AB/E2END[6]
+ Tile_X5Y13_LUT4AB/E2END[7] Tile_X5Y13_LUT4AB/E2MID[0] Tile_X5Y13_LUT4AB/E2MID[1]
+ Tile_X5Y13_LUT4AB/E2MID[2] Tile_X5Y13_LUT4AB/E2MID[3] Tile_X5Y13_LUT4AB/E2MID[4]
+ Tile_X5Y13_LUT4AB/E2MID[5] Tile_X5Y13_LUT4AB/E2MID[6] Tile_X5Y13_LUT4AB/E2MID[7]
+ Tile_X6Y13_LUT4AB/E6END[0] Tile_X6Y13_LUT4AB/E6END[10] Tile_X6Y13_LUT4AB/E6END[11]
+ Tile_X6Y13_LUT4AB/E6END[1] Tile_X6Y13_LUT4AB/E6END[2] Tile_X6Y13_LUT4AB/E6END[3]
+ Tile_X6Y13_LUT4AB/E6END[4] Tile_X6Y13_LUT4AB/E6END[5] Tile_X6Y13_LUT4AB/E6END[6]
+ Tile_X6Y13_LUT4AB/E6END[7] Tile_X6Y13_LUT4AB/E6END[8] Tile_X6Y13_LUT4AB/E6END[9]
+ Tile_X5Y13_LUT4AB/E6END[0] Tile_X5Y13_LUT4AB/E6END[10] Tile_X5Y13_LUT4AB/E6END[11]
+ Tile_X5Y13_LUT4AB/E6END[1] Tile_X5Y13_LUT4AB/E6END[2] Tile_X5Y13_LUT4AB/E6END[3]
+ Tile_X5Y13_LUT4AB/E6END[4] Tile_X5Y13_LUT4AB/E6END[5] Tile_X5Y13_LUT4AB/E6END[6]
+ Tile_X5Y13_LUT4AB/E6END[7] Tile_X5Y13_LUT4AB/E6END[8] Tile_X5Y13_LUT4AB/E6END[9]
+ Tile_X6Y13_LUT4AB/EE4END[0] Tile_X6Y13_LUT4AB/EE4END[10] Tile_X6Y13_LUT4AB/EE4END[11]
+ Tile_X6Y13_LUT4AB/EE4END[12] Tile_X6Y13_LUT4AB/EE4END[13] Tile_X6Y13_LUT4AB/EE4END[14]
+ Tile_X6Y13_LUT4AB/EE4END[15] Tile_X6Y13_LUT4AB/EE4END[1] Tile_X6Y13_LUT4AB/EE4END[2]
+ Tile_X6Y13_LUT4AB/EE4END[3] Tile_X6Y13_LUT4AB/EE4END[4] Tile_X6Y13_LUT4AB/EE4END[5]
+ Tile_X6Y13_LUT4AB/EE4END[6] Tile_X6Y13_LUT4AB/EE4END[7] Tile_X6Y13_LUT4AB/EE4END[8]
+ Tile_X6Y13_LUT4AB/EE4END[9] Tile_X5Y13_LUT4AB/EE4END[0] Tile_X5Y13_LUT4AB/EE4END[10]
+ Tile_X5Y13_LUT4AB/EE4END[11] Tile_X5Y13_LUT4AB/EE4END[12] Tile_X5Y13_LUT4AB/EE4END[13]
+ Tile_X5Y13_LUT4AB/EE4END[14] Tile_X5Y13_LUT4AB/EE4END[15] Tile_X5Y13_LUT4AB/EE4END[1]
+ Tile_X5Y13_LUT4AB/EE4END[2] Tile_X5Y13_LUT4AB/EE4END[3] Tile_X5Y13_LUT4AB/EE4END[4]
+ Tile_X5Y13_LUT4AB/EE4END[5] Tile_X5Y13_LUT4AB/EE4END[6] Tile_X5Y13_LUT4AB/EE4END[7]
+ Tile_X5Y13_LUT4AB/EE4END[8] Tile_X5Y13_LUT4AB/EE4END[9] Tile_X5Y13_LUT4AB/FrameData[0]
+ Tile_X5Y13_LUT4AB/FrameData[10] Tile_X5Y13_LUT4AB/FrameData[11] Tile_X5Y13_LUT4AB/FrameData[12]
+ Tile_X5Y13_LUT4AB/FrameData[13] Tile_X5Y13_LUT4AB/FrameData[14] Tile_X5Y13_LUT4AB/FrameData[15]
+ Tile_X5Y13_LUT4AB/FrameData[16] Tile_X5Y13_LUT4AB/FrameData[17] Tile_X5Y13_LUT4AB/FrameData[18]
+ Tile_X5Y13_LUT4AB/FrameData[19] Tile_X5Y13_LUT4AB/FrameData[1] Tile_X5Y13_LUT4AB/FrameData[20]
+ Tile_X5Y13_LUT4AB/FrameData[21] Tile_X5Y13_LUT4AB/FrameData[22] Tile_X5Y13_LUT4AB/FrameData[23]
+ Tile_X5Y13_LUT4AB/FrameData[24] Tile_X5Y13_LUT4AB/FrameData[25] Tile_X5Y13_LUT4AB/FrameData[26]
+ Tile_X5Y13_LUT4AB/FrameData[27] Tile_X5Y13_LUT4AB/FrameData[28] Tile_X5Y13_LUT4AB/FrameData[29]
+ Tile_X5Y13_LUT4AB/FrameData[2] Tile_X5Y13_LUT4AB/FrameData[30] Tile_X5Y13_LUT4AB/FrameData[31]
+ Tile_X5Y13_LUT4AB/FrameData[3] Tile_X5Y13_LUT4AB/FrameData[4] Tile_X5Y13_LUT4AB/FrameData[5]
+ Tile_X5Y13_LUT4AB/FrameData[6] Tile_X5Y13_LUT4AB/FrameData[7] Tile_X5Y13_LUT4AB/FrameData[8]
+ Tile_X5Y13_LUT4AB/FrameData[9] Tile_X6Y13_LUT4AB/FrameData[0] Tile_X6Y13_LUT4AB/FrameData[10]
+ Tile_X6Y13_LUT4AB/FrameData[11] Tile_X6Y13_LUT4AB/FrameData[12] Tile_X6Y13_LUT4AB/FrameData[13]
+ Tile_X6Y13_LUT4AB/FrameData[14] Tile_X6Y13_LUT4AB/FrameData[15] Tile_X6Y13_LUT4AB/FrameData[16]
+ Tile_X6Y13_LUT4AB/FrameData[17] Tile_X6Y13_LUT4AB/FrameData[18] Tile_X6Y13_LUT4AB/FrameData[19]
+ Tile_X6Y13_LUT4AB/FrameData[1] Tile_X6Y13_LUT4AB/FrameData[20] Tile_X6Y13_LUT4AB/FrameData[21]
+ Tile_X6Y13_LUT4AB/FrameData[22] Tile_X6Y13_LUT4AB/FrameData[23] Tile_X6Y13_LUT4AB/FrameData[24]
+ Tile_X6Y13_LUT4AB/FrameData[25] Tile_X6Y13_LUT4AB/FrameData[26] Tile_X6Y13_LUT4AB/FrameData[27]
+ Tile_X6Y13_LUT4AB/FrameData[28] Tile_X6Y13_LUT4AB/FrameData[29] Tile_X6Y13_LUT4AB/FrameData[2]
+ Tile_X6Y13_LUT4AB/FrameData[30] Tile_X6Y13_LUT4AB/FrameData[31] Tile_X6Y13_LUT4AB/FrameData[3]
+ Tile_X6Y13_LUT4AB/FrameData[4] Tile_X6Y13_LUT4AB/FrameData[5] Tile_X6Y13_LUT4AB/FrameData[6]
+ Tile_X6Y13_LUT4AB/FrameData[7] Tile_X6Y13_LUT4AB/FrameData[8] Tile_X6Y13_LUT4AB/FrameData[9]
+ Tile_X5Y13_LUT4AB/FrameStrobe[0] Tile_X5Y13_LUT4AB/FrameStrobe[10] Tile_X5Y13_LUT4AB/FrameStrobe[11]
+ Tile_X5Y13_LUT4AB/FrameStrobe[12] Tile_X5Y13_LUT4AB/FrameStrobe[13] Tile_X5Y13_LUT4AB/FrameStrobe[14]
+ Tile_X5Y13_LUT4AB/FrameStrobe[15] Tile_X5Y13_LUT4AB/FrameStrobe[16] Tile_X5Y13_LUT4AB/FrameStrobe[17]
+ Tile_X5Y13_LUT4AB/FrameStrobe[18] Tile_X5Y13_LUT4AB/FrameStrobe[19] Tile_X5Y13_LUT4AB/FrameStrobe[1]
+ Tile_X5Y13_LUT4AB/FrameStrobe[2] Tile_X5Y13_LUT4AB/FrameStrobe[3] Tile_X5Y13_LUT4AB/FrameStrobe[4]
+ Tile_X5Y13_LUT4AB/FrameStrobe[5] Tile_X5Y13_LUT4AB/FrameStrobe[6] Tile_X5Y13_LUT4AB/FrameStrobe[7]
+ Tile_X5Y13_LUT4AB/FrameStrobe[8] Tile_X5Y13_LUT4AB/FrameStrobe[9] Tile_X5Y12_LUT4AB/FrameStrobe[0]
+ Tile_X5Y12_LUT4AB/FrameStrobe[10] Tile_X5Y12_LUT4AB/FrameStrobe[11] Tile_X5Y12_LUT4AB/FrameStrobe[12]
+ Tile_X5Y12_LUT4AB/FrameStrobe[13] Tile_X5Y12_LUT4AB/FrameStrobe[14] Tile_X5Y12_LUT4AB/FrameStrobe[15]
+ Tile_X5Y12_LUT4AB/FrameStrobe[16] Tile_X5Y12_LUT4AB/FrameStrobe[17] Tile_X5Y12_LUT4AB/FrameStrobe[18]
+ Tile_X5Y12_LUT4AB/FrameStrobe[19] Tile_X5Y12_LUT4AB/FrameStrobe[1] Tile_X5Y12_LUT4AB/FrameStrobe[2]
+ Tile_X5Y12_LUT4AB/FrameStrobe[3] Tile_X5Y12_LUT4AB/FrameStrobe[4] Tile_X5Y12_LUT4AB/FrameStrobe[5]
+ Tile_X5Y12_LUT4AB/FrameStrobe[6] Tile_X5Y12_LUT4AB/FrameStrobe[7] Tile_X5Y12_LUT4AB/FrameStrobe[8]
+ Tile_X5Y12_LUT4AB/FrameStrobe[9] Tile_X5Y13_LUT4AB/N1BEG[0] Tile_X5Y13_LUT4AB/N1BEG[1]
+ Tile_X5Y13_LUT4AB/N1BEG[2] Tile_X5Y13_LUT4AB/N1BEG[3] Tile_X5Y14_LUT4AB/N1BEG[0]
+ Tile_X5Y14_LUT4AB/N1BEG[1] Tile_X5Y14_LUT4AB/N1BEG[2] Tile_X5Y14_LUT4AB/N1BEG[3]
+ Tile_X5Y13_LUT4AB/N2BEG[0] Tile_X5Y13_LUT4AB/N2BEG[1] Tile_X5Y13_LUT4AB/N2BEG[2]
+ Tile_X5Y13_LUT4AB/N2BEG[3] Tile_X5Y13_LUT4AB/N2BEG[4] Tile_X5Y13_LUT4AB/N2BEG[5]
+ Tile_X5Y13_LUT4AB/N2BEG[6] Tile_X5Y13_LUT4AB/N2BEG[7] Tile_X5Y12_LUT4AB/N2END[0]
+ Tile_X5Y12_LUT4AB/N2END[1] Tile_X5Y12_LUT4AB/N2END[2] Tile_X5Y12_LUT4AB/N2END[3]
+ Tile_X5Y12_LUT4AB/N2END[4] Tile_X5Y12_LUT4AB/N2END[5] Tile_X5Y12_LUT4AB/N2END[6]
+ Tile_X5Y12_LUT4AB/N2END[7] Tile_X5Y13_LUT4AB/N2END[0] Tile_X5Y13_LUT4AB/N2END[1]
+ Tile_X5Y13_LUT4AB/N2END[2] Tile_X5Y13_LUT4AB/N2END[3] Tile_X5Y13_LUT4AB/N2END[4]
+ Tile_X5Y13_LUT4AB/N2END[5] Tile_X5Y13_LUT4AB/N2END[6] Tile_X5Y13_LUT4AB/N2END[7]
+ Tile_X5Y14_LUT4AB/N2BEG[0] Tile_X5Y14_LUT4AB/N2BEG[1] Tile_X5Y14_LUT4AB/N2BEG[2]
+ Tile_X5Y14_LUT4AB/N2BEG[3] Tile_X5Y14_LUT4AB/N2BEG[4] Tile_X5Y14_LUT4AB/N2BEG[5]
+ Tile_X5Y14_LUT4AB/N2BEG[6] Tile_X5Y14_LUT4AB/N2BEG[7] Tile_X5Y13_LUT4AB/N4BEG[0]
+ Tile_X5Y13_LUT4AB/N4BEG[10] Tile_X5Y13_LUT4AB/N4BEG[11] Tile_X5Y13_LUT4AB/N4BEG[12]
+ Tile_X5Y13_LUT4AB/N4BEG[13] Tile_X5Y13_LUT4AB/N4BEG[14] Tile_X5Y13_LUT4AB/N4BEG[15]
+ Tile_X5Y13_LUT4AB/N4BEG[1] Tile_X5Y13_LUT4AB/N4BEG[2] Tile_X5Y13_LUT4AB/N4BEG[3]
+ Tile_X5Y13_LUT4AB/N4BEG[4] Tile_X5Y13_LUT4AB/N4BEG[5] Tile_X5Y13_LUT4AB/N4BEG[6]
+ Tile_X5Y13_LUT4AB/N4BEG[7] Tile_X5Y13_LUT4AB/N4BEG[8] Tile_X5Y13_LUT4AB/N4BEG[9]
+ Tile_X5Y14_LUT4AB/N4BEG[0] Tile_X5Y14_LUT4AB/N4BEG[10] Tile_X5Y14_LUT4AB/N4BEG[11]
+ Tile_X5Y14_LUT4AB/N4BEG[12] Tile_X5Y14_LUT4AB/N4BEG[13] Tile_X5Y14_LUT4AB/N4BEG[14]
+ Tile_X5Y14_LUT4AB/N4BEG[15] Tile_X5Y14_LUT4AB/N4BEG[1] Tile_X5Y14_LUT4AB/N4BEG[2]
+ Tile_X5Y14_LUT4AB/N4BEG[3] Tile_X5Y14_LUT4AB/N4BEG[4] Tile_X5Y14_LUT4AB/N4BEG[5]
+ Tile_X5Y14_LUT4AB/N4BEG[6] Tile_X5Y14_LUT4AB/N4BEG[7] Tile_X5Y14_LUT4AB/N4BEG[8]
+ Tile_X5Y14_LUT4AB/N4BEG[9] Tile_X5Y13_LUT4AB/NN4BEG[0] Tile_X5Y13_LUT4AB/NN4BEG[10]
+ Tile_X5Y13_LUT4AB/NN4BEG[11] Tile_X5Y13_LUT4AB/NN4BEG[12] Tile_X5Y13_LUT4AB/NN4BEG[13]
+ Tile_X5Y13_LUT4AB/NN4BEG[14] Tile_X5Y13_LUT4AB/NN4BEG[15] Tile_X5Y13_LUT4AB/NN4BEG[1]
+ Tile_X5Y13_LUT4AB/NN4BEG[2] Tile_X5Y13_LUT4AB/NN4BEG[3] Tile_X5Y13_LUT4AB/NN4BEG[4]
+ Tile_X5Y13_LUT4AB/NN4BEG[5] Tile_X5Y13_LUT4AB/NN4BEG[6] Tile_X5Y13_LUT4AB/NN4BEG[7]
+ Tile_X5Y13_LUT4AB/NN4BEG[8] Tile_X5Y13_LUT4AB/NN4BEG[9] Tile_X5Y14_LUT4AB/NN4BEG[0]
+ Tile_X5Y14_LUT4AB/NN4BEG[10] Tile_X5Y14_LUT4AB/NN4BEG[11] Tile_X5Y14_LUT4AB/NN4BEG[12]
+ Tile_X5Y14_LUT4AB/NN4BEG[13] Tile_X5Y14_LUT4AB/NN4BEG[14] Tile_X5Y14_LUT4AB/NN4BEG[15]
+ Tile_X5Y14_LUT4AB/NN4BEG[1] Tile_X5Y14_LUT4AB/NN4BEG[2] Tile_X5Y14_LUT4AB/NN4BEG[3]
+ Tile_X5Y14_LUT4AB/NN4BEG[4] Tile_X5Y14_LUT4AB/NN4BEG[5] Tile_X5Y14_LUT4AB/NN4BEG[6]
+ Tile_X5Y14_LUT4AB/NN4BEG[7] Tile_X5Y14_LUT4AB/NN4BEG[8] Tile_X5Y14_LUT4AB/NN4BEG[9]
+ Tile_X5Y14_LUT4AB/S1END[0] Tile_X5Y14_LUT4AB/S1END[1] Tile_X5Y14_LUT4AB/S1END[2]
+ Tile_X5Y14_LUT4AB/S1END[3] Tile_X5Y13_LUT4AB/S1END[0] Tile_X5Y13_LUT4AB/S1END[1]
+ Tile_X5Y13_LUT4AB/S1END[2] Tile_X5Y13_LUT4AB/S1END[3] Tile_X5Y14_LUT4AB/S2MID[0]
+ Tile_X5Y14_LUT4AB/S2MID[1] Tile_X5Y14_LUT4AB/S2MID[2] Tile_X5Y14_LUT4AB/S2MID[3]
+ Tile_X5Y14_LUT4AB/S2MID[4] Tile_X5Y14_LUT4AB/S2MID[5] Tile_X5Y14_LUT4AB/S2MID[6]
+ Tile_X5Y14_LUT4AB/S2MID[7] Tile_X5Y14_LUT4AB/S2END[0] Tile_X5Y14_LUT4AB/S2END[1]
+ Tile_X5Y14_LUT4AB/S2END[2] Tile_X5Y14_LUT4AB/S2END[3] Tile_X5Y14_LUT4AB/S2END[4]
+ Tile_X5Y14_LUT4AB/S2END[5] Tile_X5Y14_LUT4AB/S2END[6] Tile_X5Y14_LUT4AB/S2END[7]
+ Tile_X5Y13_LUT4AB/S2END[0] Tile_X5Y13_LUT4AB/S2END[1] Tile_X5Y13_LUT4AB/S2END[2]
+ Tile_X5Y13_LUT4AB/S2END[3] Tile_X5Y13_LUT4AB/S2END[4] Tile_X5Y13_LUT4AB/S2END[5]
+ Tile_X5Y13_LUT4AB/S2END[6] Tile_X5Y13_LUT4AB/S2END[7] Tile_X5Y13_LUT4AB/S2MID[0]
+ Tile_X5Y13_LUT4AB/S2MID[1] Tile_X5Y13_LUT4AB/S2MID[2] Tile_X5Y13_LUT4AB/S2MID[3]
+ Tile_X5Y13_LUT4AB/S2MID[4] Tile_X5Y13_LUT4AB/S2MID[5] Tile_X5Y13_LUT4AB/S2MID[6]
+ Tile_X5Y13_LUT4AB/S2MID[7] Tile_X5Y14_LUT4AB/S4END[0] Tile_X5Y14_LUT4AB/S4END[10]
+ Tile_X5Y14_LUT4AB/S4END[11] Tile_X5Y14_LUT4AB/S4END[12] Tile_X5Y14_LUT4AB/S4END[13]
+ Tile_X5Y14_LUT4AB/S4END[14] Tile_X5Y14_LUT4AB/S4END[15] Tile_X5Y14_LUT4AB/S4END[1]
+ Tile_X5Y14_LUT4AB/S4END[2] Tile_X5Y14_LUT4AB/S4END[3] Tile_X5Y14_LUT4AB/S4END[4]
+ Tile_X5Y14_LUT4AB/S4END[5] Tile_X5Y14_LUT4AB/S4END[6] Tile_X5Y14_LUT4AB/S4END[7]
+ Tile_X5Y14_LUT4AB/S4END[8] Tile_X5Y14_LUT4AB/S4END[9] Tile_X5Y13_LUT4AB/S4END[0]
+ Tile_X5Y13_LUT4AB/S4END[10] Tile_X5Y13_LUT4AB/S4END[11] Tile_X5Y13_LUT4AB/S4END[12]
+ Tile_X5Y13_LUT4AB/S4END[13] Tile_X5Y13_LUT4AB/S4END[14] Tile_X5Y13_LUT4AB/S4END[15]
+ Tile_X5Y13_LUT4AB/S4END[1] Tile_X5Y13_LUT4AB/S4END[2] Tile_X5Y13_LUT4AB/S4END[3]
+ Tile_X5Y13_LUT4AB/S4END[4] Tile_X5Y13_LUT4AB/S4END[5] Tile_X5Y13_LUT4AB/S4END[6]
+ Tile_X5Y13_LUT4AB/S4END[7] Tile_X5Y13_LUT4AB/S4END[8] Tile_X5Y13_LUT4AB/S4END[9]
+ Tile_X5Y14_LUT4AB/SS4END[0] Tile_X5Y14_LUT4AB/SS4END[10] Tile_X5Y14_LUT4AB/SS4END[11]
+ Tile_X5Y14_LUT4AB/SS4END[12] Tile_X5Y14_LUT4AB/SS4END[13] Tile_X5Y14_LUT4AB/SS4END[14]
+ Tile_X5Y14_LUT4AB/SS4END[15] Tile_X5Y14_LUT4AB/SS4END[1] Tile_X5Y14_LUT4AB/SS4END[2]
+ Tile_X5Y14_LUT4AB/SS4END[3] Tile_X5Y14_LUT4AB/SS4END[4] Tile_X5Y14_LUT4AB/SS4END[5]
+ Tile_X5Y14_LUT4AB/SS4END[6] Tile_X5Y14_LUT4AB/SS4END[7] Tile_X5Y14_LUT4AB/SS4END[8]
+ Tile_X5Y14_LUT4AB/SS4END[9] Tile_X5Y13_LUT4AB/SS4END[0] Tile_X5Y13_LUT4AB/SS4END[10]
+ Tile_X5Y13_LUT4AB/SS4END[11] Tile_X5Y13_LUT4AB/SS4END[12] Tile_X5Y13_LUT4AB/SS4END[13]
+ Tile_X5Y13_LUT4AB/SS4END[14] Tile_X5Y13_LUT4AB/SS4END[15] Tile_X5Y13_LUT4AB/SS4END[1]
+ Tile_X5Y13_LUT4AB/SS4END[2] Tile_X5Y13_LUT4AB/SS4END[3] Tile_X5Y13_LUT4AB/SS4END[4]
+ Tile_X5Y13_LUT4AB/SS4END[5] Tile_X5Y13_LUT4AB/SS4END[6] Tile_X5Y13_LUT4AB/SS4END[7]
+ Tile_X5Y13_LUT4AB/SS4END[8] Tile_X5Y13_LUT4AB/SS4END[9] Tile_X5Y13_LUT4AB/UserCLK
+ Tile_X5Y12_LUT4AB/UserCLK VGND VPWR Tile_X5Y13_LUT4AB/W1BEG[0] Tile_X5Y13_LUT4AB/W1BEG[1]
+ Tile_X5Y13_LUT4AB/W1BEG[2] Tile_X5Y13_LUT4AB/W1BEG[3] Tile_X6Y13_LUT4AB/W1BEG[0]
+ Tile_X6Y13_LUT4AB/W1BEG[1] Tile_X6Y13_LUT4AB/W1BEG[2] Tile_X6Y13_LUT4AB/W1BEG[3]
+ Tile_X5Y13_LUT4AB/W2BEG[0] Tile_X5Y13_LUT4AB/W2BEG[1] Tile_X5Y13_LUT4AB/W2BEG[2]
+ Tile_X5Y13_LUT4AB/W2BEG[3] Tile_X5Y13_LUT4AB/W2BEG[4] Tile_X5Y13_LUT4AB/W2BEG[5]
+ Tile_X5Y13_LUT4AB/W2BEG[6] Tile_X5Y13_LUT4AB/W2BEG[7] Tile_X5Y13_LUT4AB/W2BEGb[0]
+ Tile_X5Y13_LUT4AB/W2BEGb[1] Tile_X5Y13_LUT4AB/W2BEGb[2] Tile_X5Y13_LUT4AB/W2BEGb[3]
+ Tile_X5Y13_LUT4AB/W2BEGb[4] Tile_X5Y13_LUT4AB/W2BEGb[5] Tile_X5Y13_LUT4AB/W2BEGb[6]
+ Tile_X5Y13_LUT4AB/W2BEGb[7] Tile_X5Y13_LUT4AB/W2END[0] Tile_X5Y13_LUT4AB/W2END[1]
+ Tile_X5Y13_LUT4AB/W2END[2] Tile_X5Y13_LUT4AB/W2END[3] Tile_X5Y13_LUT4AB/W2END[4]
+ Tile_X5Y13_LUT4AB/W2END[5] Tile_X5Y13_LUT4AB/W2END[6] Tile_X5Y13_LUT4AB/W2END[7]
+ Tile_X6Y13_LUT4AB/W2BEG[0] Tile_X6Y13_LUT4AB/W2BEG[1] Tile_X6Y13_LUT4AB/W2BEG[2]
+ Tile_X6Y13_LUT4AB/W2BEG[3] Tile_X6Y13_LUT4AB/W2BEG[4] Tile_X6Y13_LUT4AB/W2BEG[5]
+ Tile_X6Y13_LUT4AB/W2BEG[6] Tile_X6Y13_LUT4AB/W2BEG[7] Tile_X5Y13_LUT4AB/W6BEG[0]
+ Tile_X5Y13_LUT4AB/W6BEG[10] Tile_X5Y13_LUT4AB/W6BEG[11] Tile_X5Y13_LUT4AB/W6BEG[1]
+ Tile_X5Y13_LUT4AB/W6BEG[2] Tile_X5Y13_LUT4AB/W6BEG[3] Tile_X5Y13_LUT4AB/W6BEG[4]
+ Tile_X5Y13_LUT4AB/W6BEG[5] Tile_X5Y13_LUT4AB/W6BEG[6] Tile_X5Y13_LUT4AB/W6BEG[7]
+ Tile_X5Y13_LUT4AB/W6BEG[8] Tile_X5Y13_LUT4AB/W6BEG[9] Tile_X6Y13_LUT4AB/W6BEG[0]
+ Tile_X6Y13_LUT4AB/W6BEG[10] Tile_X6Y13_LUT4AB/W6BEG[11] Tile_X6Y13_LUT4AB/W6BEG[1]
+ Tile_X6Y13_LUT4AB/W6BEG[2] Tile_X6Y13_LUT4AB/W6BEG[3] Tile_X6Y13_LUT4AB/W6BEG[4]
+ Tile_X6Y13_LUT4AB/W6BEG[5] Tile_X6Y13_LUT4AB/W6BEG[6] Tile_X6Y13_LUT4AB/W6BEG[7]
+ Tile_X6Y13_LUT4AB/W6BEG[8] Tile_X6Y13_LUT4AB/W6BEG[9] Tile_X5Y13_LUT4AB/WW4BEG[0]
+ Tile_X5Y13_LUT4AB/WW4BEG[10] Tile_X5Y13_LUT4AB/WW4BEG[11] Tile_X5Y13_LUT4AB/WW4BEG[12]
+ Tile_X5Y13_LUT4AB/WW4BEG[13] Tile_X5Y13_LUT4AB/WW4BEG[14] Tile_X5Y13_LUT4AB/WW4BEG[15]
+ Tile_X5Y13_LUT4AB/WW4BEG[1] Tile_X5Y13_LUT4AB/WW4BEG[2] Tile_X5Y13_LUT4AB/WW4BEG[3]
+ Tile_X5Y13_LUT4AB/WW4BEG[4] Tile_X5Y13_LUT4AB/WW4BEG[5] Tile_X5Y13_LUT4AB/WW4BEG[6]
+ Tile_X5Y13_LUT4AB/WW4BEG[7] Tile_X5Y13_LUT4AB/WW4BEG[8] Tile_X5Y13_LUT4AB/WW4BEG[9]
+ Tile_X6Y13_LUT4AB/WW4BEG[0] Tile_X6Y13_LUT4AB/WW4BEG[10] Tile_X6Y13_LUT4AB/WW4BEG[11]
+ Tile_X6Y13_LUT4AB/WW4BEG[12] Tile_X6Y13_LUT4AB/WW4BEG[13] Tile_X6Y13_LUT4AB/WW4BEG[14]
+ Tile_X6Y13_LUT4AB/WW4BEG[15] Tile_X6Y13_LUT4AB/WW4BEG[1] Tile_X6Y13_LUT4AB/WW4BEG[2]
+ Tile_X6Y13_LUT4AB/WW4BEG[3] Tile_X6Y13_LUT4AB/WW4BEG[4] Tile_X6Y13_LUT4AB/WW4BEG[5]
+ Tile_X6Y13_LUT4AB/WW4BEG[6] Tile_X6Y13_LUT4AB/WW4BEG[7] Tile_X6Y13_LUT4AB/WW4BEG[8]
+ Tile_X6Y13_LUT4AB/WW4BEG[9] LUT4AB
XTile_X0Y6_W_IO Tile_X0Y6_A_I_top Tile_X0Y6_A_O_top Tile_X0Y6_A_T_top Tile_X0Y6_A_config_C_bit0
+ Tile_X0Y6_A_config_C_bit1 Tile_X0Y6_A_config_C_bit2 Tile_X0Y6_A_config_C_bit3 Tile_X0Y6_B_I_top
+ Tile_X0Y6_B_O_top Tile_X0Y6_B_T_top Tile_X0Y6_B_config_C_bit0 Tile_X0Y6_B_config_C_bit1
+ Tile_X0Y6_B_config_C_bit2 Tile_X0Y6_B_config_C_bit3 Tile_X0Y6_W_IO/E1BEG[0] Tile_X0Y6_W_IO/E1BEG[1]
+ Tile_X0Y6_W_IO/E1BEG[2] Tile_X0Y6_W_IO/E1BEG[3] Tile_X0Y6_W_IO/E2BEG[0] Tile_X0Y6_W_IO/E2BEG[1]
+ Tile_X0Y6_W_IO/E2BEG[2] Tile_X0Y6_W_IO/E2BEG[3] Tile_X0Y6_W_IO/E2BEG[4] Tile_X0Y6_W_IO/E2BEG[5]
+ Tile_X0Y6_W_IO/E2BEG[6] Tile_X0Y6_W_IO/E2BEG[7] Tile_X0Y6_W_IO/E2BEGb[0] Tile_X0Y6_W_IO/E2BEGb[1]
+ Tile_X0Y6_W_IO/E2BEGb[2] Tile_X0Y6_W_IO/E2BEGb[3] Tile_X0Y6_W_IO/E2BEGb[4] Tile_X0Y6_W_IO/E2BEGb[5]
+ Tile_X0Y6_W_IO/E2BEGb[6] Tile_X0Y6_W_IO/E2BEGb[7] Tile_X0Y6_W_IO/E6BEG[0] Tile_X0Y6_W_IO/E6BEG[10]
+ Tile_X0Y6_W_IO/E6BEG[11] Tile_X0Y6_W_IO/E6BEG[1] Tile_X0Y6_W_IO/E6BEG[2] Tile_X0Y6_W_IO/E6BEG[3]
+ Tile_X0Y6_W_IO/E6BEG[4] Tile_X0Y6_W_IO/E6BEG[5] Tile_X0Y6_W_IO/E6BEG[6] Tile_X0Y6_W_IO/E6BEG[7]
+ Tile_X0Y6_W_IO/E6BEG[8] Tile_X0Y6_W_IO/E6BEG[9] Tile_X0Y6_W_IO/EE4BEG[0] Tile_X0Y6_W_IO/EE4BEG[10]
+ Tile_X0Y6_W_IO/EE4BEG[11] Tile_X0Y6_W_IO/EE4BEG[12] Tile_X0Y6_W_IO/EE4BEG[13] Tile_X0Y6_W_IO/EE4BEG[14]
+ Tile_X0Y6_W_IO/EE4BEG[15] Tile_X0Y6_W_IO/EE4BEG[1] Tile_X0Y6_W_IO/EE4BEG[2] Tile_X0Y6_W_IO/EE4BEG[3]
+ Tile_X0Y6_W_IO/EE4BEG[4] Tile_X0Y6_W_IO/EE4BEG[5] Tile_X0Y6_W_IO/EE4BEG[6] Tile_X0Y6_W_IO/EE4BEG[7]
+ Tile_X0Y6_W_IO/EE4BEG[8] Tile_X0Y6_W_IO/EE4BEG[9] FrameData[192] FrameData[202]
+ FrameData[203] FrameData[204] FrameData[205] FrameData[206] FrameData[207] FrameData[208]
+ FrameData[209] FrameData[210] FrameData[211] FrameData[193] FrameData[212] FrameData[213]
+ FrameData[214] FrameData[215] FrameData[216] FrameData[217] FrameData[218] FrameData[219]
+ FrameData[220] FrameData[221] FrameData[194] FrameData[222] FrameData[223] FrameData[195]
+ FrameData[196] FrameData[197] FrameData[198] FrameData[199] FrameData[200] FrameData[201]
+ Tile_X1Y6_LUT4AB/FrameData[0] Tile_X1Y6_LUT4AB/FrameData[10] Tile_X1Y6_LUT4AB/FrameData[11]
+ Tile_X1Y6_LUT4AB/FrameData[12] Tile_X1Y6_LUT4AB/FrameData[13] Tile_X1Y6_LUT4AB/FrameData[14]
+ Tile_X1Y6_LUT4AB/FrameData[15] Tile_X1Y6_LUT4AB/FrameData[16] Tile_X1Y6_LUT4AB/FrameData[17]
+ Tile_X1Y6_LUT4AB/FrameData[18] Tile_X1Y6_LUT4AB/FrameData[19] Tile_X1Y6_LUT4AB/FrameData[1]
+ Tile_X1Y6_LUT4AB/FrameData[20] Tile_X1Y6_LUT4AB/FrameData[21] Tile_X1Y6_LUT4AB/FrameData[22]
+ Tile_X1Y6_LUT4AB/FrameData[23] Tile_X1Y6_LUT4AB/FrameData[24] Tile_X1Y6_LUT4AB/FrameData[25]
+ Tile_X1Y6_LUT4AB/FrameData[26] Tile_X1Y6_LUT4AB/FrameData[27] Tile_X1Y6_LUT4AB/FrameData[28]
+ Tile_X1Y6_LUT4AB/FrameData[29] Tile_X1Y6_LUT4AB/FrameData[2] Tile_X1Y6_LUT4AB/FrameData[30]
+ Tile_X1Y6_LUT4AB/FrameData[31] Tile_X1Y6_LUT4AB/FrameData[3] Tile_X1Y6_LUT4AB/FrameData[4]
+ Tile_X1Y6_LUT4AB/FrameData[5] Tile_X1Y6_LUT4AB/FrameData[6] Tile_X1Y6_LUT4AB/FrameData[7]
+ Tile_X1Y6_LUT4AB/FrameData[8] Tile_X1Y6_LUT4AB/FrameData[9] Tile_X0Y6_W_IO/FrameStrobe[0]
+ Tile_X0Y6_W_IO/FrameStrobe[10] Tile_X0Y6_W_IO/FrameStrobe[11] Tile_X0Y6_W_IO/FrameStrobe[12]
+ Tile_X0Y6_W_IO/FrameStrobe[13] Tile_X0Y6_W_IO/FrameStrobe[14] Tile_X0Y6_W_IO/FrameStrobe[15]
+ Tile_X0Y6_W_IO/FrameStrobe[16] Tile_X0Y6_W_IO/FrameStrobe[17] Tile_X0Y6_W_IO/FrameStrobe[18]
+ Tile_X0Y6_W_IO/FrameStrobe[19] Tile_X0Y6_W_IO/FrameStrobe[1] Tile_X0Y6_W_IO/FrameStrobe[2]
+ Tile_X0Y6_W_IO/FrameStrobe[3] Tile_X0Y6_W_IO/FrameStrobe[4] Tile_X0Y6_W_IO/FrameStrobe[5]
+ Tile_X0Y6_W_IO/FrameStrobe[6] Tile_X0Y6_W_IO/FrameStrobe[7] Tile_X0Y6_W_IO/FrameStrobe[8]
+ Tile_X0Y6_W_IO/FrameStrobe[9] Tile_X0Y5_W_IO/FrameStrobe[0] Tile_X0Y5_W_IO/FrameStrobe[10]
+ Tile_X0Y5_W_IO/FrameStrobe[11] Tile_X0Y5_W_IO/FrameStrobe[12] Tile_X0Y5_W_IO/FrameStrobe[13]
+ Tile_X0Y5_W_IO/FrameStrobe[14] Tile_X0Y5_W_IO/FrameStrobe[15] Tile_X0Y5_W_IO/FrameStrobe[16]
+ Tile_X0Y5_W_IO/FrameStrobe[17] Tile_X0Y5_W_IO/FrameStrobe[18] Tile_X0Y5_W_IO/FrameStrobe[19]
+ Tile_X0Y5_W_IO/FrameStrobe[1] Tile_X0Y5_W_IO/FrameStrobe[2] Tile_X0Y5_W_IO/FrameStrobe[3]
+ Tile_X0Y5_W_IO/FrameStrobe[4] Tile_X0Y5_W_IO/FrameStrobe[5] Tile_X0Y5_W_IO/FrameStrobe[6]
+ Tile_X0Y5_W_IO/FrameStrobe[7] Tile_X0Y5_W_IO/FrameStrobe[8] Tile_X0Y5_W_IO/FrameStrobe[9]
+ Tile_X0Y6_W_IO/UserCLK Tile_X0Y5_W_IO/UserCLK VGND VPWR Tile_X0Y6_W_IO/W1END[0]
+ Tile_X0Y6_W_IO/W1END[1] Tile_X0Y6_W_IO/W1END[2] Tile_X0Y6_W_IO/W1END[3] Tile_X0Y6_W_IO/W2END[0]
+ Tile_X0Y6_W_IO/W2END[1] Tile_X0Y6_W_IO/W2END[2] Tile_X0Y6_W_IO/W2END[3] Tile_X0Y6_W_IO/W2END[4]
+ Tile_X0Y6_W_IO/W2END[5] Tile_X0Y6_W_IO/W2END[6] Tile_X0Y6_W_IO/W2END[7] Tile_X0Y6_W_IO/W2MID[0]
+ Tile_X0Y6_W_IO/W2MID[1] Tile_X0Y6_W_IO/W2MID[2] Tile_X0Y6_W_IO/W2MID[3] Tile_X0Y6_W_IO/W2MID[4]
+ Tile_X0Y6_W_IO/W2MID[5] Tile_X0Y6_W_IO/W2MID[6] Tile_X0Y6_W_IO/W2MID[7] Tile_X0Y6_W_IO/W6END[0]
+ Tile_X0Y6_W_IO/W6END[10] Tile_X0Y6_W_IO/W6END[11] Tile_X0Y6_W_IO/W6END[1] Tile_X0Y6_W_IO/W6END[2]
+ Tile_X0Y6_W_IO/W6END[3] Tile_X0Y6_W_IO/W6END[4] Tile_X0Y6_W_IO/W6END[5] Tile_X0Y6_W_IO/W6END[6]
+ Tile_X0Y6_W_IO/W6END[7] Tile_X0Y6_W_IO/W6END[8] Tile_X0Y6_W_IO/W6END[9] Tile_X0Y6_W_IO/WW4END[0]
+ Tile_X0Y6_W_IO/WW4END[10] Tile_X0Y6_W_IO/WW4END[11] Tile_X0Y6_W_IO/WW4END[12] Tile_X0Y6_W_IO/WW4END[13]
+ Tile_X0Y6_W_IO/WW4END[14] Tile_X0Y6_W_IO/WW4END[15] Tile_X0Y6_W_IO/WW4END[1] Tile_X0Y6_W_IO/WW4END[2]
+ Tile_X0Y6_W_IO/WW4END[3] Tile_X0Y6_W_IO/WW4END[4] Tile_X0Y6_W_IO/WW4END[5] Tile_X0Y6_W_IO/WW4END[6]
+ Tile_X0Y6_W_IO/WW4END[7] Tile_X0Y6_W_IO/WW4END[8] Tile_X0Y6_W_IO/WW4END[9] W_IO
XTile_X8Y6_LUT4AB Tile_X8Y7_LUT4AB/Co Tile_X8Y6_LUT4AB/Co Tile_X9Y6_LUT4AB/E1END[0]
+ Tile_X9Y6_LUT4AB/E1END[1] Tile_X9Y6_LUT4AB/E1END[2] Tile_X9Y6_LUT4AB/E1END[3] Tile_X8Y6_LUT4AB/E1END[0]
+ Tile_X8Y6_LUT4AB/E1END[1] Tile_X8Y6_LUT4AB/E1END[2] Tile_X8Y6_LUT4AB/E1END[3] Tile_X9Y6_LUT4AB/E2MID[0]
+ Tile_X9Y6_LUT4AB/E2MID[1] Tile_X9Y6_LUT4AB/E2MID[2] Tile_X9Y6_LUT4AB/E2MID[3] Tile_X9Y6_LUT4AB/E2MID[4]
+ Tile_X9Y6_LUT4AB/E2MID[5] Tile_X9Y6_LUT4AB/E2MID[6] Tile_X9Y6_LUT4AB/E2MID[7] Tile_X9Y6_LUT4AB/E2END[0]
+ Tile_X9Y6_LUT4AB/E2END[1] Tile_X9Y6_LUT4AB/E2END[2] Tile_X9Y6_LUT4AB/E2END[3] Tile_X9Y6_LUT4AB/E2END[4]
+ Tile_X9Y6_LUT4AB/E2END[5] Tile_X9Y6_LUT4AB/E2END[6] Tile_X9Y6_LUT4AB/E2END[7] Tile_X8Y6_LUT4AB/E2END[0]
+ Tile_X8Y6_LUT4AB/E2END[1] Tile_X8Y6_LUT4AB/E2END[2] Tile_X8Y6_LUT4AB/E2END[3] Tile_X8Y6_LUT4AB/E2END[4]
+ Tile_X8Y6_LUT4AB/E2END[5] Tile_X8Y6_LUT4AB/E2END[6] Tile_X8Y6_LUT4AB/E2END[7] Tile_X8Y6_LUT4AB/E2MID[0]
+ Tile_X8Y6_LUT4AB/E2MID[1] Tile_X8Y6_LUT4AB/E2MID[2] Tile_X8Y6_LUT4AB/E2MID[3] Tile_X8Y6_LUT4AB/E2MID[4]
+ Tile_X8Y6_LUT4AB/E2MID[5] Tile_X8Y6_LUT4AB/E2MID[6] Tile_X8Y6_LUT4AB/E2MID[7] Tile_X9Y6_LUT4AB/E6END[0]
+ Tile_X9Y6_LUT4AB/E6END[10] Tile_X9Y6_LUT4AB/E6END[11] Tile_X9Y6_LUT4AB/E6END[1]
+ Tile_X9Y6_LUT4AB/E6END[2] Tile_X9Y6_LUT4AB/E6END[3] Tile_X9Y6_LUT4AB/E6END[4] Tile_X9Y6_LUT4AB/E6END[5]
+ Tile_X9Y6_LUT4AB/E6END[6] Tile_X9Y6_LUT4AB/E6END[7] Tile_X9Y6_LUT4AB/E6END[8] Tile_X9Y6_LUT4AB/E6END[9]
+ Tile_X8Y6_LUT4AB/E6END[0] Tile_X8Y6_LUT4AB/E6END[10] Tile_X8Y6_LUT4AB/E6END[11]
+ Tile_X8Y6_LUT4AB/E6END[1] Tile_X8Y6_LUT4AB/E6END[2] Tile_X8Y6_LUT4AB/E6END[3] Tile_X8Y6_LUT4AB/E6END[4]
+ Tile_X8Y6_LUT4AB/E6END[5] Tile_X8Y6_LUT4AB/E6END[6] Tile_X8Y6_LUT4AB/E6END[7] Tile_X8Y6_LUT4AB/E6END[8]
+ Tile_X8Y6_LUT4AB/E6END[9] Tile_X9Y6_LUT4AB/EE4END[0] Tile_X9Y6_LUT4AB/EE4END[10]
+ Tile_X9Y6_LUT4AB/EE4END[11] Tile_X9Y6_LUT4AB/EE4END[12] Tile_X9Y6_LUT4AB/EE4END[13]
+ Tile_X9Y6_LUT4AB/EE4END[14] Tile_X9Y6_LUT4AB/EE4END[15] Tile_X9Y6_LUT4AB/EE4END[1]
+ Tile_X9Y6_LUT4AB/EE4END[2] Tile_X9Y6_LUT4AB/EE4END[3] Tile_X9Y6_LUT4AB/EE4END[4]
+ Tile_X9Y6_LUT4AB/EE4END[5] Tile_X9Y6_LUT4AB/EE4END[6] Tile_X9Y6_LUT4AB/EE4END[7]
+ Tile_X9Y6_LUT4AB/EE4END[8] Tile_X9Y6_LUT4AB/EE4END[9] Tile_X8Y6_LUT4AB/EE4END[0]
+ Tile_X8Y6_LUT4AB/EE4END[10] Tile_X8Y6_LUT4AB/EE4END[11] Tile_X8Y6_LUT4AB/EE4END[12]
+ Tile_X8Y6_LUT4AB/EE4END[13] Tile_X8Y6_LUT4AB/EE4END[14] Tile_X8Y6_LUT4AB/EE4END[15]
+ Tile_X8Y6_LUT4AB/EE4END[1] Tile_X8Y6_LUT4AB/EE4END[2] Tile_X8Y6_LUT4AB/EE4END[3]
+ Tile_X8Y6_LUT4AB/EE4END[4] Tile_X8Y6_LUT4AB/EE4END[5] Tile_X8Y6_LUT4AB/EE4END[6]
+ Tile_X8Y6_LUT4AB/EE4END[7] Tile_X8Y6_LUT4AB/EE4END[8] Tile_X8Y6_LUT4AB/EE4END[9]
+ Tile_X8Y6_LUT4AB/FrameData[0] Tile_X8Y6_LUT4AB/FrameData[10] Tile_X8Y6_LUT4AB/FrameData[11]
+ Tile_X8Y6_LUT4AB/FrameData[12] Tile_X8Y6_LUT4AB/FrameData[13] Tile_X8Y6_LUT4AB/FrameData[14]
+ Tile_X8Y6_LUT4AB/FrameData[15] Tile_X8Y6_LUT4AB/FrameData[16] Tile_X8Y6_LUT4AB/FrameData[17]
+ Tile_X8Y6_LUT4AB/FrameData[18] Tile_X8Y6_LUT4AB/FrameData[19] Tile_X8Y6_LUT4AB/FrameData[1]
+ Tile_X8Y6_LUT4AB/FrameData[20] Tile_X8Y6_LUT4AB/FrameData[21] Tile_X8Y6_LUT4AB/FrameData[22]
+ Tile_X8Y6_LUT4AB/FrameData[23] Tile_X8Y6_LUT4AB/FrameData[24] Tile_X8Y6_LUT4AB/FrameData[25]
+ Tile_X8Y6_LUT4AB/FrameData[26] Tile_X8Y6_LUT4AB/FrameData[27] Tile_X8Y6_LUT4AB/FrameData[28]
+ Tile_X8Y6_LUT4AB/FrameData[29] Tile_X8Y6_LUT4AB/FrameData[2] Tile_X8Y6_LUT4AB/FrameData[30]
+ Tile_X8Y6_LUT4AB/FrameData[31] Tile_X8Y6_LUT4AB/FrameData[3] Tile_X8Y6_LUT4AB/FrameData[4]
+ Tile_X8Y6_LUT4AB/FrameData[5] Tile_X8Y6_LUT4AB/FrameData[6] Tile_X8Y6_LUT4AB/FrameData[7]
+ Tile_X8Y6_LUT4AB/FrameData[8] Tile_X8Y6_LUT4AB/FrameData[9] Tile_X9Y6_LUT4AB/FrameData[0]
+ Tile_X9Y6_LUT4AB/FrameData[10] Tile_X9Y6_LUT4AB/FrameData[11] Tile_X9Y6_LUT4AB/FrameData[12]
+ Tile_X9Y6_LUT4AB/FrameData[13] Tile_X9Y6_LUT4AB/FrameData[14] Tile_X9Y6_LUT4AB/FrameData[15]
+ Tile_X9Y6_LUT4AB/FrameData[16] Tile_X9Y6_LUT4AB/FrameData[17] Tile_X9Y6_LUT4AB/FrameData[18]
+ Tile_X9Y6_LUT4AB/FrameData[19] Tile_X9Y6_LUT4AB/FrameData[1] Tile_X9Y6_LUT4AB/FrameData[20]
+ Tile_X9Y6_LUT4AB/FrameData[21] Tile_X9Y6_LUT4AB/FrameData[22] Tile_X9Y6_LUT4AB/FrameData[23]
+ Tile_X9Y6_LUT4AB/FrameData[24] Tile_X9Y6_LUT4AB/FrameData[25] Tile_X9Y6_LUT4AB/FrameData[26]
+ Tile_X9Y6_LUT4AB/FrameData[27] Tile_X9Y6_LUT4AB/FrameData[28] Tile_X9Y6_LUT4AB/FrameData[29]
+ Tile_X9Y6_LUT4AB/FrameData[2] Tile_X9Y6_LUT4AB/FrameData[30] Tile_X9Y6_LUT4AB/FrameData[31]
+ Tile_X9Y6_LUT4AB/FrameData[3] Tile_X9Y6_LUT4AB/FrameData[4] Tile_X9Y6_LUT4AB/FrameData[5]
+ Tile_X9Y6_LUT4AB/FrameData[6] Tile_X9Y6_LUT4AB/FrameData[7] Tile_X9Y6_LUT4AB/FrameData[8]
+ Tile_X9Y6_LUT4AB/FrameData[9] Tile_X8Y6_LUT4AB/FrameStrobe[0] Tile_X8Y6_LUT4AB/FrameStrobe[10]
+ Tile_X8Y6_LUT4AB/FrameStrobe[11] Tile_X8Y6_LUT4AB/FrameStrobe[12] Tile_X8Y6_LUT4AB/FrameStrobe[13]
+ Tile_X8Y6_LUT4AB/FrameStrobe[14] Tile_X8Y6_LUT4AB/FrameStrobe[15] Tile_X8Y6_LUT4AB/FrameStrobe[16]
+ Tile_X8Y6_LUT4AB/FrameStrobe[17] Tile_X8Y6_LUT4AB/FrameStrobe[18] Tile_X8Y6_LUT4AB/FrameStrobe[19]
+ Tile_X8Y6_LUT4AB/FrameStrobe[1] Tile_X8Y6_LUT4AB/FrameStrobe[2] Tile_X8Y6_LUT4AB/FrameStrobe[3]
+ Tile_X8Y6_LUT4AB/FrameStrobe[4] Tile_X8Y6_LUT4AB/FrameStrobe[5] Tile_X8Y6_LUT4AB/FrameStrobe[6]
+ Tile_X8Y6_LUT4AB/FrameStrobe[7] Tile_X8Y6_LUT4AB/FrameStrobe[8] Tile_X8Y6_LUT4AB/FrameStrobe[9]
+ Tile_X8Y5_LUT4AB/FrameStrobe[0] Tile_X8Y5_LUT4AB/FrameStrobe[10] Tile_X8Y5_LUT4AB/FrameStrobe[11]
+ Tile_X8Y5_LUT4AB/FrameStrobe[12] Tile_X8Y5_LUT4AB/FrameStrobe[13] Tile_X8Y5_LUT4AB/FrameStrobe[14]
+ Tile_X8Y5_LUT4AB/FrameStrobe[15] Tile_X8Y5_LUT4AB/FrameStrobe[16] Tile_X8Y5_LUT4AB/FrameStrobe[17]
+ Tile_X8Y5_LUT4AB/FrameStrobe[18] Tile_X8Y5_LUT4AB/FrameStrobe[19] Tile_X8Y5_LUT4AB/FrameStrobe[1]
+ Tile_X8Y5_LUT4AB/FrameStrobe[2] Tile_X8Y5_LUT4AB/FrameStrobe[3] Tile_X8Y5_LUT4AB/FrameStrobe[4]
+ Tile_X8Y5_LUT4AB/FrameStrobe[5] Tile_X8Y5_LUT4AB/FrameStrobe[6] Tile_X8Y5_LUT4AB/FrameStrobe[7]
+ Tile_X8Y5_LUT4AB/FrameStrobe[8] Tile_X8Y5_LUT4AB/FrameStrobe[9] Tile_X8Y6_LUT4AB/N1BEG[0]
+ Tile_X8Y6_LUT4AB/N1BEG[1] Tile_X8Y6_LUT4AB/N1BEG[2] Tile_X8Y6_LUT4AB/N1BEG[3] Tile_X8Y7_LUT4AB/N1BEG[0]
+ Tile_X8Y7_LUT4AB/N1BEG[1] Tile_X8Y7_LUT4AB/N1BEG[2] Tile_X8Y7_LUT4AB/N1BEG[3] Tile_X8Y6_LUT4AB/N2BEG[0]
+ Tile_X8Y6_LUT4AB/N2BEG[1] Tile_X8Y6_LUT4AB/N2BEG[2] Tile_X8Y6_LUT4AB/N2BEG[3] Tile_X8Y6_LUT4AB/N2BEG[4]
+ Tile_X8Y6_LUT4AB/N2BEG[5] Tile_X8Y6_LUT4AB/N2BEG[6] Tile_X8Y6_LUT4AB/N2BEG[7] Tile_X8Y5_LUT4AB/N2END[0]
+ Tile_X8Y5_LUT4AB/N2END[1] Tile_X8Y5_LUT4AB/N2END[2] Tile_X8Y5_LUT4AB/N2END[3] Tile_X8Y5_LUT4AB/N2END[4]
+ Tile_X8Y5_LUT4AB/N2END[5] Tile_X8Y5_LUT4AB/N2END[6] Tile_X8Y5_LUT4AB/N2END[7] Tile_X8Y6_LUT4AB/N2END[0]
+ Tile_X8Y6_LUT4AB/N2END[1] Tile_X8Y6_LUT4AB/N2END[2] Tile_X8Y6_LUT4AB/N2END[3] Tile_X8Y6_LUT4AB/N2END[4]
+ Tile_X8Y6_LUT4AB/N2END[5] Tile_X8Y6_LUT4AB/N2END[6] Tile_X8Y6_LUT4AB/N2END[7] Tile_X8Y7_LUT4AB/N2BEG[0]
+ Tile_X8Y7_LUT4AB/N2BEG[1] Tile_X8Y7_LUT4AB/N2BEG[2] Tile_X8Y7_LUT4AB/N2BEG[3] Tile_X8Y7_LUT4AB/N2BEG[4]
+ Tile_X8Y7_LUT4AB/N2BEG[5] Tile_X8Y7_LUT4AB/N2BEG[6] Tile_X8Y7_LUT4AB/N2BEG[7] Tile_X8Y6_LUT4AB/N4BEG[0]
+ Tile_X8Y6_LUT4AB/N4BEG[10] Tile_X8Y6_LUT4AB/N4BEG[11] Tile_X8Y6_LUT4AB/N4BEG[12]
+ Tile_X8Y6_LUT4AB/N4BEG[13] Tile_X8Y6_LUT4AB/N4BEG[14] Tile_X8Y6_LUT4AB/N4BEG[15]
+ Tile_X8Y6_LUT4AB/N4BEG[1] Tile_X8Y6_LUT4AB/N4BEG[2] Tile_X8Y6_LUT4AB/N4BEG[3] Tile_X8Y6_LUT4AB/N4BEG[4]
+ Tile_X8Y6_LUT4AB/N4BEG[5] Tile_X8Y6_LUT4AB/N4BEG[6] Tile_X8Y6_LUT4AB/N4BEG[7] Tile_X8Y6_LUT4AB/N4BEG[8]
+ Tile_X8Y6_LUT4AB/N4BEG[9] Tile_X8Y7_LUT4AB/N4BEG[0] Tile_X8Y7_LUT4AB/N4BEG[10] Tile_X8Y7_LUT4AB/N4BEG[11]
+ Tile_X8Y7_LUT4AB/N4BEG[12] Tile_X8Y7_LUT4AB/N4BEG[13] Tile_X8Y7_LUT4AB/N4BEG[14]
+ Tile_X8Y7_LUT4AB/N4BEG[15] Tile_X8Y7_LUT4AB/N4BEG[1] Tile_X8Y7_LUT4AB/N4BEG[2] Tile_X8Y7_LUT4AB/N4BEG[3]
+ Tile_X8Y7_LUT4AB/N4BEG[4] Tile_X8Y7_LUT4AB/N4BEG[5] Tile_X8Y7_LUT4AB/N4BEG[6] Tile_X8Y7_LUT4AB/N4BEG[7]
+ Tile_X8Y7_LUT4AB/N4BEG[8] Tile_X8Y7_LUT4AB/N4BEG[9] Tile_X8Y6_LUT4AB/NN4BEG[0] Tile_X8Y6_LUT4AB/NN4BEG[10]
+ Tile_X8Y6_LUT4AB/NN4BEG[11] Tile_X8Y6_LUT4AB/NN4BEG[12] Tile_X8Y6_LUT4AB/NN4BEG[13]
+ Tile_X8Y6_LUT4AB/NN4BEG[14] Tile_X8Y6_LUT4AB/NN4BEG[15] Tile_X8Y6_LUT4AB/NN4BEG[1]
+ Tile_X8Y6_LUT4AB/NN4BEG[2] Tile_X8Y6_LUT4AB/NN4BEG[3] Tile_X8Y6_LUT4AB/NN4BEG[4]
+ Tile_X8Y6_LUT4AB/NN4BEG[5] Tile_X8Y6_LUT4AB/NN4BEG[6] Tile_X8Y6_LUT4AB/NN4BEG[7]
+ Tile_X8Y6_LUT4AB/NN4BEG[8] Tile_X8Y6_LUT4AB/NN4BEG[9] Tile_X8Y7_LUT4AB/NN4BEG[0]
+ Tile_X8Y7_LUT4AB/NN4BEG[10] Tile_X8Y7_LUT4AB/NN4BEG[11] Tile_X8Y7_LUT4AB/NN4BEG[12]
+ Tile_X8Y7_LUT4AB/NN4BEG[13] Tile_X8Y7_LUT4AB/NN4BEG[14] Tile_X8Y7_LUT4AB/NN4BEG[15]
+ Tile_X8Y7_LUT4AB/NN4BEG[1] Tile_X8Y7_LUT4AB/NN4BEG[2] Tile_X8Y7_LUT4AB/NN4BEG[3]
+ Tile_X8Y7_LUT4AB/NN4BEG[4] Tile_X8Y7_LUT4AB/NN4BEG[5] Tile_X8Y7_LUT4AB/NN4BEG[6]
+ Tile_X8Y7_LUT4AB/NN4BEG[7] Tile_X8Y7_LUT4AB/NN4BEG[8] Tile_X8Y7_LUT4AB/NN4BEG[9]
+ Tile_X8Y7_LUT4AB/S1END[0] Tile_X8Y7_LUT4AB/S1END[1] Tile_X8Y7_LUT4AB/S1END[2] Tile_X8Y7_LUT4AB/S1END[3]
+ Tile_X8Y6_LUT4AB/S1END[0] Tile_X8Y6_LUT4AB/S1END[1] Tile_X8Y6_LUT4AB/S1END[2] Tile_X8Y6_LUT4AB/S1END[3]
+ Tile_X8Y7_LUT4AB/S2MID[0] Tile_X8Y7_LUT4AB/S2MID[1] Tile_X8Y7_LUT4AB/S2MID[2] Tile_X8Y7_LUT4AB/S2MID[3]
+ Tile_X8Y7_LUT4AB/S2MID[4] Tile_X8Y7_LUT4AB/S2MID[5] Tile_X8Y7_LUT4AB/S2MID[6] Tile_X8Y7_LUT4AB/S2MID[7]
+ Tile_X8Y7_LUT4AB/S2END[0] Tile_X8Y7_LUT4AB/S2END[1] Tile_X8Y7_LUT4AB/S2END[2] Tile_X8Y7_LUT4AB/S2END[3]
+ Tile_X8Y7_LUT4AB/S2END[4] Tile_X8Y7_LUT4AB/S2END[5] Tile_X8Y7_LUT4AB/S2END[6] Tile_X8Y7_LUT4AB/S2END[7]
+ Tile_X8Y6_LUT4AB/S2END[0] Tile_X8Y6_LUT4AB/S2END[1] Tile_X8Y6_LUT4AB/S2END[2] Tile_X8Y6_LUT4AB/S2END[3]
+ Tile_X8Y6_LUT4AB/S2END[4] Tile_X8Y6_LUT4AB/S2END[5] Tile_X8Y6_LUT4AB/S2END[6] Tile_X8Y6_LUT4AB/S2END[7]
+ Tile_X8Y6_LUT4AB/S2MID[0] Tile_X8Y6_LUT4AB/S2MID[1] Tile_X8Y6_LUT4AB/S2MID[2] Tile_X8Y6_LUT4AB/S2MID[3]
+ Tile_X8Y6_LUT4AB/S2MID[4] Tile_X8Y6_LUT4AB/S2MID[5] Tile_X8Y6_LUT4AB/S2MID[6] Tile_X8Y6_LUT4AB/S2MID[7]
+ Tile_X8Y7_LUT4AB/S4END[0] Tile_X8Y7_LUT4AB/S4END[10] Tile_X8Y7_LUT4AB/S4END[11]
+ Tile_X8Y7_LUT4AB/S4END[12] Tile_X8Y7_LUT4AB/S4END[13] Tile_X8Y7_LUT4AB/S4END[14]
+ Tile_X8Y7_LUT4AB/S4END[15] Tile_X8Y7_LUT4AB/S4END[1] Tile_X8Y7_LUT4AB/S4END[2] Tile_X8Y7_LUT4AB/S4END[3]
+ Tile_X8Y7_LUT4AB/S4END[4] Tile_X8Y7_LUT4AB/S4END[5] Tile_X8Y7_LUT4AB/S4END[6] Tile_X8Y7_LUT4AB/S4END[7]
+ Tile_X8Y7_LUT4AB/S4END[8] Tile_X8Y7_LUT4AB/S4END[9] Tile_X8Y6_LUT4AB/S4END[0] Tile_X8Y6_LUT4AB/S4END[10]
+ Tile_X8Y6_LUT4AB/S4END[11] Tile_X8Y6_LUT4AB/S4END[12] Tile_X8Y6_LUT4AB/S4END[13]
+ Tile_X8Y6_LUT4AB/S4END[14] Tile_X8Y6_LUT4AB/S4END[15] Tile_X8Y6_LUT4AB/S4END[1]
+ Tile_X8Y6_LUT4AB/S4END[2] Tile_X8Y6_LUT4AB/S4END[3] Tile_X8Y6_LUT4AB/S4END[4] Tile_X8Y6_LUT4AB/S4END[5]
+ Tile_X8Y6_LUT4AB/S4END[6] Tile_X8Y6_LUT4AB/S4END[7] Tile_X8Y6_LUT4AB/S4END[8] Tile_X8Y6_LUT4AB/S4END[9]
+ Tile_X8Y7_LUT4AB/SS4END[0] Tile_X8Y7_LUT4AB/SS4END[10] Tile_X8Y7_LUT4AB/SS4END[11]
+ Tile_X8Y7_LUT4AB/SS4END[12] Tile_X8Y7_LUT4AB/SS4END[13] Tile_X8Y7_LUT4AB/SS4END[14]
+ Tile_X8Y7_LUT4AB/SS4END[15] Tile_X8Y7_LUT4AB/SS4END[1] Tile_X8Y7_LUT4AB/SS4END[2]
+ Tile_X8Y7_LUT4AB/SS4END[3] Tile_X8Y7_LUT4AB/SS4END[4] Tile_X8Y7_LUT4AB/SS4END[5]
+ Tile_X8Y7_LUT4AB/SS4END[6] Tile_X8Y7_LUT4AB/SS4END[7] Tile_X8Y7_LUT4AB/SS4END[8]
+ Tile_X8Y7_LUT4AB/SS4END[9] Tile_X8Y6_LUT4AB/SS4END[0] Tile_X8Y6_LUT4AB/SS4END[10]
+ Tile_X8Y6_LUT4AB/SS4END[11] Tile_X8Y6_LUT4AB/SS4END[12] Tile_X8Y6_LUT4AB/SS4END[13]
+ Tile_X8Y6_LUT4AB/SS4END[14] Tile_X8Y6_LUT4AB/SS4END[15] Tile_X8Y6_LUT4AB/SS4END[1]
+ Tile_X8Y6_LUT4AB/SS4END[2] Tile_X8Y6_LUT4AB/SS4END[3] Tile_X8Y6_LUT4AB/SS4END[4]
+ Tile_X8Y6_LUT4AB/SS4END[5] Tile_X8Y6_LUT4AB/SS4END[6] Tile_X8Y6_LUT4AB/SS4END[7]
+ Tile_X8Y6_LUT4AB/SS4END[8] Tile_X8Y6_LUT4AB/SS4END[9] Tile_X8Y6_LUT4AB/UserCLK Tile_X8Y5_LUT4AB/UserCLK
+ VGND VPWR Tile_X8Y6_LUT4AB/W1BEG[0] Tile_X8Y6_LUT4AB/W1BEG[1] Tile_X8Y6_LUT4AB/W1BEG[2]
+ Tile_X8Y6_LUT4AB/W1BEG[3] Tile_X9Y6_LUT4AB/W1BEG[0] Tile_X9Y6_LUT4AB/W1BEG[1] Tile_X9Y6_LUT4AB/W1BEG[2]
+ Tile_X9Y6_LUT4AB/W1BEG[3] Tile_X8Y6_LUT4AB/W2BEG[0] Tile_X8Y6_LUT4AB/W2BEG[1] Tile_X8Y6_LUT4AB/W2BEG[2]
+ Tile_X8Y6_LUT4AB/W2BEG[3] Tile_X8Y6_LUT4AB/W2BEG[4] Tile_X8Y6_LUT4AB/W2BEG[5] Tile_X8Y6_LUT4AB/W2BEG[6]
+ Tile_X8Y6_LUT4AB/W2BEG[7] Tile_X8Y6_LUT4AB/W2BEGb[0] Tile_X8Y6_LUT4AB/W2BEGb[1]
+ Tile_X8Y6_LUT4AB/W2BEGb[2] Tile_X8Y6_LUT4AB/W2BEGb[3] Tile_X8Y6_LUT4AB/W2BEGb[4]
+ Tile_X8Y6_LUT4AB/W2BEGb[5] Tile_X8Y6_LUT4AB/W2BEGb[6] Tile_X8Y6_LUT4AB/W2BEGb[7]
+ Tile_X8Y6_LUT4AB/W2END[0] Tile_X8Y6_LUT4AB/W2END[1] Tile_X8Y6_LUT4AB/W2END[2] Tile_X8Y6_LUT4AB/W2END[3]
+ Tile_X8Y6_LUT4AB/W2END[4] Tile_X8Y6_LUT4AB/W2END[5] Tile_X8Y6_LUT4AB/W2END[6] Tile_X8Y6_LUT4AB/W2END[7]
+ Tile_X9Y6_LUT4AB/W2BEG[0] Tile_X9Y6_LUT4AB/W2BEG[1] Tile_X9Y6_LUT4AB/W2BEG[2] Tile_X9Y6_LUT4AB/W2BEG[3]
+ Tile_X9Y6_LUT4AB/W2BEG[4] Tile_X9Y6_LUT4AB/W2BEG[5] Tile_X9Y6_LUT4AB/W2BEG[6] Tile_X9Y6_LUT4AB/W2BEG[7]
+ Tile_X8Y6_LUT4AB/W6BEG[0] Tile_X8Y6_LUT4AB/W6BEG[10] Tile_X8Y6_LUT4AB/W6BEG[11]
+ Tile_X8Y6_LUT4AB/W6BEG[1] Tile_X8Y6_LUT4AB/W6BEG[2] Tile_X8Y6_LUT4AB/W6BEG[3] Tile_X8Y6_LUT4AB/W6BEG[4]
+ Tile_X8Y6_LUT4AB/W6BEG[5] Tile_X8Y6_LUT4AB/W6BEG[6] Tile_X8Y6_LUT4AB/W6BEG[7] Tile_X8Y6_LUT4AB/W6BEG[8]
+ Tile_X8Y6_LUT4AB/W6BEG[9] Tile_X9Y6_LUT4AB/W6BEG[0] Tile_X9Y6_LUT4AB/W6BEG[10] Tile_X9Y6_LUT4AB/W6BEG[11]
+ Tile_X9Y6_LUT4AB/W6BEG[1] Tile_X9Y6_LUT4AB/W6BEG[2] Tile_X9Y6_LUT4AB/W6BEG[3] Tile_X9Y6_LUT4AB/W6BEG[4]
+ Tile_X9Y6_LUT4AB/W6BEG[5] Tile_X9Y6_LUT4AB/W6BEG[6] Tile_X9Y6_LUT4AB/W6BEG[7] Tile_X9Y6_LUT4AB/W6BEG[8]
+ Tile_X9Y6_LUT4AB/W6BEG[9] Tile_X8Y6_LUT4AB/WW4BEG[0] Tile_X8Y6_LUT4AB/WW4BEG[10]
+ Tile_X8Y6_LUT4AB/WW4BEG[11] Tile_X8Y6_LUT4AB/WW4BEG[12] Tile_X8Y6_LUT4AB/WW4BEG[13]
+ Tile_X8Y6_LUT4AB/WW4BEG[14] Tile_X8Y6_LUT4AB/WW4BEG[15] Tile_X8Y6_LUT4AB/WW4BEG[1]
+ Tile_X8Y6_LUT4AB/WW4BEG[2] Tile_X8Y6_LUT4AB/WW4BEG[3] Tile_X8Y6_LUT4AB/WW4BEG[4]
+ Tile_X8Y6_LUT4AB/WW4BEG[5] Tile_X8Y6_LUT4AB/WW4BEG[6] Tile_X8Y6_LUT4AB/WW4BEG[7]
+ Tile_X8Y6_LUT4AB/WW4BEG[8] Tile_X8Y6_LUT4AB/WW4BEG[9] Tile_X9Y6_LUT4AB/WW4BEG[0]
+ Tile_X9Y6_LUT4AB/WW4BEG[10] Tile_X9Y6_LUT4AB/WW4BEG[11] Tile_X9Y6_LUT4AB/WW4BEG[12]
+ Tile_X9Y6_LUT4AB/WW4BEG[13] Tile_X9Y6_LUT4AB/WW4BEG[14] Tile_X9Y6_LUT4AB/WW4BEG[15]
+ Tile_X9Y6_LUT4AB/WW4BEG[1] Tile_X9Y6_LUT4AB/WW4BEG[2] Tile_X9Y6_LUT4AB/WW4BEG[3]
+ Tile_X9Y6_LUT4AB/WW4BEG[4] Tile_X9Y6_LUT4AB/WW4BEG[5] Tile_X9Y6_LUT4AB/WW4BEG[6]
+ Tile_X9Y6_LUT4AB/WW4BEG[7] Tile_X9Y6_LUT4AB/WW4BEG[8] Tile_X9Y6_LUT4AB/WW4BEG[9]
+ LUT4AB
XTile_X5Y1_LUT4AB Tile_X5Y2_LUT4AB/Co Tile_X5Y1_LUT4AB/Co Tile_X6Y1_LUT4AB/E1END[0]
+ Tile_X6Y1_LUT4AB/E1END[1] Tile_X6Y1_LUT4AB/E1END[2] Tile_X6Y1_LUT4AB/E1END[3] Tile_X5Y1_LUT4AB/E1END[0]
+ Tile_X5Y1_LUT4AB/E1END[1] Tile_X5Y1_LUT4AB/E1END[2] Tile_X5Y1_LUT4AB/E1END[3] Tile_X6Y1_LUT4AB/E2MID[0]
+ Tile_X6Y1_LUT4AB/E2MID[1] Tile_X6Y1_LUT4AB/E2MID[2] Tile_X6Y1_LUT4AB/E2MID[3] Tile_X6Y1_LUT4AB/E2MID[4]
+ Tile_X6Y1_LUT4AB/E2MID[5] Tile_X6Y1_LUT4AB/E2MID[6] Tile_X6Y1_LUT4AB/E2MID[7] Tile_X6Y1_LUT4AB/E2END[0]
+ Tile_X6Y1_LUT4AB/E2END[1] Tile_X6Y1_LUT4AB/E2END[2] Tile_X6Y1_LUT4AB/E2END[3] Tile_X6Y1_LUT4AB/E2END[4]
+ Tile_X6Y1_LUT4AB/E2END[5] Tile_X6Y1_LUT4AB/E2END[6] Tile_X6Y1_LUT4AB/E2END[7] Tile_X5Y1_LUT4AB/E2END[0]
+ Tile_X5Y1_LUT4AB/E2END[1] Tile_X5Y1_LUT4AB/E2END[2] Tile_X5Y1_LUT4AB/E2END[3] Tile_X5Y1_LUT4AB/E2END[4]
+ Tile_X5Y1_LUT4AB/E2END[5] Tile_X5Y1_LUT4AB/E2END[6] Tile_X5Y1_LUT4AB/E2END[7] Tile_X5Y1_LUT4AB/E2MID[0]
+ Tile_X5Y1_LUT4AB/E2MID[1] Tile_X5Y1_LUT4AB/E2MID[2] Tile_X5Y1_LUT4AB/E2MID[3] Tile_X5Y1_LUT4AB/E2MID[4]
+ Tile_X5Y1_LUT4AB/E2MID[5] Tile_X5Y1_LUT4AB/E2MID[6] Tile_X5Y1_LUT4AB/E2MID[7] Tile_X6Y1_LUT4AB/E6END[0]
+ Tile_X6Y1_LUT4AB/E6END[10] Tile_X6Y1_LUT4AB/E6END[11] Tile_X6Y1_LUT4AB/E6END[1]
+ Tile_X6Y1_LUT4AB/E6END[2] Tile_X6Y1_LUT4AB/E6END[3] Tile_X6Y1_LUT4AB/E6END[4] Tile_X6Y1_LUT4AB/E6END[5]
+ Tile_X6Y1_LUT4AB/E6END[6] Tile_X6Y1_LUT4AB/E6END[7] Tile_X6Y1_LUT4AB/E6END[8] Tile_X6Y1_LUT4AB/E6END[9]
+ Tile_X5Y1_LUT4AB/E6END[0] Tile_X5Y1_LUT4AB/E6END[10] Tile_X5Y1_LUT4AB/E6END[11]
+ Tile_X5Y1_LUT4AB/E6END[1] Tile_X5Y1_LUT4AB/E6END[2] Tile_X5Y1_LUT4AB/E6END[3] Tile_X5Y1_LUT4AB/E6END[4]
+ Tile_X5Y1_LUT4AB/E6END[5] Tile_X5Y1_LUT4AB/E6END[6] Tile_X5Y1_LUT4AB/E6END[7] Tile_X5Y1_LUT4AB/E6END[8]
+ Tile_X5Y1_LUT4AB/E6END[9] Tile_X6Y1_LUT4AB/EE4END[0] Tile_X6Y1_LUT4AB/EE4END[10]
+ Tile_X6Y1_LUT4AB/EE4END[11] Tile_X6Y1_LUT4AB/EE4END[12] Tile_X6Y1_LUT4AB/EE4END[13]
+ Tile_X6Y1_LUT4AB/EE4END[14] Tile_X6Y1_LUT4AB/EE4END[15] Tile_X6Y1_LUT4AB/EE4END[1]
+ Tile_X6Y1_LUT4AB/EE4END[2] Tile_X6Y1_LUT4AB/EE4END[3] Tile_X6Y1_LUT4AB/EE4END[4]
+ Tile_X6Y1_LUT4AB/EE4END[5] Tile_X6Y1_LUT4AB/EE4END[6] Tile_X6Y1_LUT4AB/EE4END[7]
+ Tile_X6Y1_LUT4AB/EE4END[8] Tile_X6Y1_LUT4AB/EE4END[9] Tile_X5Y1_LUT4AB/EE4END[0]
+ Tile_X5Y1_LUT4AB/EE4END[10] Tile_X5Y1_LUT4AB/EE4END[11] Tile_X5Y1_LUT4AB/EE4END[12]
+ Tile_X5Y1_LUT4AB/EE4END[13] Tile_X5Y1_LUT4AB/EE4END[14] Tile_X5Y1_LUT4AB/EE4END[15]
+ Tile_X5Y1_LUT4AB/EE4END[1] Tile_X5Y1_LUT4AB/EE4END[2] Tile_X5Y1_LUT4AB/EE4END[3]
+ Tile_X5Y1_LUT4AB/EE4END[4] Tile_X5Y1_LUT4AB/EE4END[5] Tile_X5Y1_LUT4AB/EE4END[6]
+ Tile_X5Y1_LUT4AB/EE4END[7] Tile_X5Y1_LUT4AB/EE4END[8] Tile_X5Y1_LUT4AB/EE4END[9]
+ Tile_X5Y1_LUT4AB/FrameData[0] Tile_X5Y1_LUT4AB/FrameData[10] Tile_X5Y1_LUT4AB/FrameData[11]
+ Tile_X5Y1_LUT4AB/FrameData[12] Tile_X5Y1_LUT4AB/FrameData[13] Tile_X5Y1_LUT4AB/FrameData[14]
+ Tile_X5Y1_LUT4AB/FrameData[15] Tile_X5Y1_LUT4AB/FrameData[16] Tile_X5Y1_LUT4AB/FrameData[17]
+ Tile_X5Y1_LUT4AB/FrameData[18] Tile_X5Y1_LUT4AB/FrameData[19] Tile_X5Y1_LUT4AB/FrameData[1]
+ Tile_X5Y1_LUT4AB/FrameData[20] Tile_X5Y1_LUT4AB/FrameData[21] Tile_X5Y1_LUT4AB/FrameData[22]
+ Tile_X5Y1_LUT4AB/FrameData[23] Tile_X5Y1_LUT4AB/FrameData[24] Tile_X5Y1_LUT4AB/FrameData[25]
+ Tile_X5Y1_LUT4AB/FrameData[26] Tile_X5Y1_LUT4AB/FrameData[27] Tile_X5Y1_LUT4AB/FrameData[28]
+ Tile_X5Y1_LUT4AB/FrameData[29] Tile_X5Y1_LUT4AB/FrameData[2] Tile_X5Y1_LUT4AB/FrameData[30]
+ Tile_X5Y1_LUT4AB/FrameData[31] Tile_X5Y1_LUT4AB/FrameData[3] Tile_X5Y1_LUT4AB/FrameData[4]
+ Tile_X5Y1_LUT4AB/FrameData[5] Tile_X5Y1_LUT4AB/FrameData[6] Tile_X5Y1_LUT4AB/FrameData[7]
+ Tile_X5Y1_LUT4AB/FrameData[8] Tile_X5Y1_LUT4AB/FrameData[9] Tile_X6Y1_LUT4AB/FrameData[0]
+ Tile_X6Y1_LUT4AB/FrameData[10] Tile_X6Y1_LUT4AB/FrameData[11] Tile_X6Y1_LUT4AB/FrameData[12]
+ Tile_X6Y1_LUT4AB/FrameData[13] Tile_X6Y1_LUT4AB/FrameData[14] Tile_X6Y1_LUT4AB/FrameData[15]
+ Tile_X6Y1_LUT4AB/FrameData[16] Tile_X6Y1_LUT4AB/FrameData[17] Tile_X6Y1_LUT4AB/FrameData[18]
+ Tile_X6Y1_LUT4AB/FrameData[19] Tile_X6Y1_LUT4AB/FrameData[1] Tile_X6Y1_LUT4AB/FrameData[20]
+ Tile_X6Y1_LUT4AB/FrameData[21] Tile_X6Y1_LUT4AB/FrameData[22] Tile_X6Y1_LUT4AB/FrameData[23]
+ Tile_X6Y1_LUT4AB/FrameData[24] Tile_X6Y1_LUT4AB/FrameData[25] Tile_X6Y1_LUT4AB/FrameData[26]
+ Tile_X6Y1_LUT4AB/FrameData[27] Tile_X6Y1_LUT4AB/FrameData[28] Tile_X6Y1_LUT4AB/FrameData[29]
+ Tile_X6Y1_LUT4AB/FrameData[2] Tile_X6Y1_LUT4AB/FrameData[30] Tile_X6Y1_LUT4AB/FrameData[31]
+ Tile_X6Y1_LUT4AB/FrameData[3] Tile_X6Y1_LUT4AB/FrameData[4] Tile_X6Y1_LUT4AB/FrameData[5]
+ Tile_X6Y1_LUT4AB/FrameData[6] Tile_X6Y1_LUT4AB/FrameData[7] Tile_X6Y1_LUT4AB/FrameData[8]
+ Tile_X6Y1_LUT4AB/FrameData[9] Tile_X5Y1_LUT4AB/FrameStrobe[0] Tile_X5Y1_LUT4AB/FrameStrobe[10]
+ Tile_X5Y1_LUT4AB/FrameStrobe[11] Tile_X5Y1_LUT4AB/FrameStrobe[12] Tile_X5Y1_LUT4AB/FrameStrobe[13]
+ Tile_X5Y1_LUT4AB/FrameStrobe[14] Tile_X5Y1_LUT4AB/FrameStrobe[15] Tile_X5Y1_LUT4AB/FrameStrobe[16]
+ Tile_X5Y1_LUT4AB/FrameStrobe[17] Tile_X5Y1_LUT4AB/FrameStrobe[18] Tile_X5Y1_LUT4AB/FrameStrobe[19]
+ Tile_X5Y1_LUT4AB/FrameStrobe[1] Tile_X5Y1_LUT4AB/FrameStrobe[2] Tile_X5Y1_LUT4AB/FrameStrobe[3]
+ Tile_X5Y1_LUT4AB/FrameStrobe[4] Tile_X5Y1_LUT4AB/FrameStrobe[5] Tile_X5Y1_LUT4AB/FrameStrobe[6]
+ Tile_X5Y1_LUT4AB/FrameStrobe[7] Tile_X5Y1_LUT4AB/FrameStrobe[8] Tile_X5Y1_LUT4AB/FrameStrobe[9]
+ Tile_X5Y1_LUT4AB/FrameStrobe_O[0] Tile_X5Y1_LUT4AB/FrameStrobe_O[10] Tile_X5Y1_LUT4AB/FrameStrobe_O[11]
+ Tile_X5Y1_LUT4AB/FrameStrobe_O[12] Tile_X5Y1_LUT4AB/FrameStrobe_O[13] Tile_X5Y1_LUT4AB/FrameStrobe_O[14]
+ Tile_X5Y1_LUT4AB/FrameStrobe_O[15] Tile_X5Y1_LUT4AB/FrameStrobe_O[16] Tile_X5Y1_LUT4AB/FrameStrobe_O[17]
+ Tile_X5Y1_LUT4AB/FrameStrobe_O[18] Tile_X5Y1_LUT4AB/FrameStrobe_O[19] Tile_X5Y1_LUT4AB/FrameStrobe_O[1]
+ Tile_X5Y1_LUT4AB/FrameStrobe_O[2] Tile_X5Y1_LUT4AB/FrameStrobe_O[3] Tile_X5Y1_LUT4AB/FrameStrobe_O[4]
+ Tile_X5Y1_LUT4AB/FrameStrobe_O[5] Tile_X5Y1_LUT4AB/FrameStrobe_O[6] Tile_X5Y1_LUT4AB/FrameStrobe_O[7]
+ Tile_X5Y1_LUT4AB/FrameStrobe_O[8] Tile_X5Y1_LUT4AB/FrameStrobe_O[9] Tile_X5Y1_LUT4AB/N1BEG[0]
+ Tile_X5Y1_LUT4AB/N1BEG[1] Tile_X5Y1_LUT4AB/N1BEG[2] Tile_X5Y1_LUT4AB/N1BEG[3] Tile_X5Y2_LUT4AB/N1BEG[0]
+ Tile_X5Y2_LUT4AB/N1BEG[1] Tile_X5Y2_LUT4AB/N1BEG[2] Tile_X5Y2_LUT4AB/N1BEG[3] Tile_X5Y1_LUT4AB/N2BEG[0]
+ Tile_X5Y1_LUT4AB/N2BEG[1] Tile_X5Y1_LUT4AB/N2BEG[2] Tile_X5Y1_LUT4AB/N2BEG[3] Tile_X5Y1_LUT4AB/N2BEG[4]
+ Tile_X5Y1_LUT4AB/N2BEG[5] Tile_X5Y1_LUT4AB/N2BEG[6] Tile_X5Y1_LUT4AB/N2BEG[7] Tile_X5Y1_LUT4AB/N2BEGb[0]
+ Tile_X5Y1_LUT4AB/N2BEGb[1] Tile_X5Y1_LUT4AB/N2BEGb[2] Tile_X5Y1_LUT4AB/N2BEGb[3]
+ Tile_X5Y1_LUT4AB/N2BEGb[4] Tile_X5Y1_LUT4AB/N2BEGb[5] Tile_X5Y1_LUT4AB/N2BEGb[6]
+ Tile_X5Y1_LUT4AB/N2BEGb[7] Tile_X5Y1_LUT4AB/N2END[0] Tile_X5Y1_LUT4AB/N2END[1] Tile_X5Y1_LUT4AB/N2END[2]
+ Tile_X5Y1_LUT4AB/N2END[3] Tile_X5Y1_LUT4AB/N2END[4] Tile_X5Y1_LUT4AB/N2END[5] Tile_X5Y1_LUT4AB/N2END[6]
+ Tile_X5Y1_LUT4AB/N2END[7] Tile_X5Y2_LUT4AB/N2BEG[0] Tile_X5Y2_LUT4AB/N2BEG[1] Tile_X5Y2_LUT4AB/N2BEG[2]
+ Tile_X5Y2_LUT4AB/N2BEG[3] Tile_X5Y2_LUT4AB/N2BEG[4] Tile_X5Y2_LUT4AB/N2BEG[5] Tile_X5Y2_LUT4AB/N2BEG[6]
+ Tile_X5Y2_LUT4AB/N2BEG[7] Tile_X5Y1_LUT4AB/N4BEG[0] Tile_X5Y1_LUT4AB/N4BEG[10] Tile_X5Y1_LUT4AB/N4BEG[11]
+ Tile_X5Y1_LUT4AB/N4BEG[12] Tile_X5Y1_LUT4AB/N4BEG[13] Tile_X5Y1_LUT4AB/N4BEG[14]
+ Tile_X5Y1_LUT4AB/N4BEG[15] Tile_X5Y1_LUT4AB/N4BEG[1] Tile_X5Y1_LUT4AB/N4BEG[2] Tile_X5Y1_LUT4AB/N4BEG[3]
+ Tile_X5Y1_LUT4AB/N4BEG[4] Tile_X5Y1_LUT4AB/N4BEG[5] Tile_X5Y1_LUT4AB/N4BEG[6] Tile_X5Y1_LUT4AB/N4BEG[7]
+ Tile_X5Y1_LUT4AB/N4BEG[8] Tile_X5Y1_LUT4AB/N4BEG[9] Tile_X5Y2_LUT4AB/N4BEG[0] Tile_X5Y2_LUT4AB/N4BEG[10]
+ Tile_X5Y2_LUT4AB/N4BEG[11] Tile_X5Y2_LUT4AB/N4BEG[12] Tile_X5Y2_LUT4AB/N4BEG[13]
+ Tile_X5Y2_LUT4AB/N4BEG[14] Tile_X5Y2_LUT4AB/N4BEG[15] Tile_X5Y2_LUT4AB/N4BEG[1]
+ Tile_X5Y2_LUT4AB/N4BEG[2] Tile_X5Y2_LUT4AB/N4BEG[3] Tile_X5Y2_LUT4AB/N4BEG[4] Tile_X5Y2_LUT4AB/N4BEG[5]
+ Tile_X5Y2_LUT4AB/N4BEG[6] Tile_X5Y2_LUT4AB/N4BEG[7] Tile_X5Y2_LUT4AB/N4BEG[8] Tile_X5Y2_LUT4AB/N4BEG[9]
+ Tile_X5Y1_LUT4AB/NN4BEG[0] Tile_X5Y1_LUT4AB/NN4BEG[10] Tile_X5Y1_LUT4AB/NN4BEG[11]
+ Tile_X5Y1_LUT4AB/NN4BEG[12] Tile_X5Y1_LUT4AB/NN4BEG[13] Tile_X5Y1_LUT4AB/NN4BEG[14]
+ Tile_X5Y1_LUT4AB/NN4BEG[15] Tile_X5Y1_LUT4AB/NN4BEG[1] Tile_X5Y1_LUT4AB/NN4BEG[2]
+ Tile_X5Y1_LUT4AB/NN4BEG[3] Tile_X5Y1_LUT4AB/NN4BEG[4] Tile_X5Y1_LUT4AB/NN4BEG[5]
+ Tile_X5Y1_LUT4AB/NN4BEG[6] Tile_X5Y1_LUT4AB/NN4BEG[7] Tile_X5Y1_LUT4AB/NN4BEG[8]
+ Tile_X5Y1_LUT4AB/NN4BEG[9] Tile_X5Y2_LUT4AB/NN4BEG[0] Tile_X5Y2_LUT4AB/NN4BEG[10]
+ Tile_X5Y2_LUT4AB/NN4BEG[11] Tile_X5Y2_LUT4AB/NN4BEG[12] Tile_X5Y2_LUT4AB/NN4BEG[13]
+ Tile_X5Y2_LUT4AB/NN4BEG[14] Tile_X5Y2_LUT4AB/NN4BEG[15] Tile_X5Y2_LUT4AB/NN4BEG[1]
+ Tile_X5Y2_LUT4AB/NN4BEG[2] Tile_X5Y2_LUT4AB/NN4BEG[3] Tile_X5Y2_LUT4AB/NN4BEG[4]
+ Tile_X5Y2_LUT4AB/NN4BEG[5] Tile_X5Y2_LUT4AB/NN4BEG[6] Tile_X5Y2_LUT4AB/NN4BEG[7]
+ Tile_X5Y2_LUT4AB/NN4BEG[8] Tile_X5Y2_LUT4AB/NN4BEG[9] Tile_X5Y2_LUT4AB/S1END[0]
+ Tile_X5Y2_LUT4AB/S1END[1] Tile_X5Y2_LUT4AB/S1END[2] Tile_X5Y2_LUT4AB/S1END[3] Tile_X5Y1_LUT4AB/S1END[0]
+ Tile_X5Y1_LUT4AB/S1END[1] Tile_X5Y1_LUT4AB/S1END[2] Tile_X5Y1_LUT4AB/S1END[3] Tile_X5Y2_LUT4AB/S2MID[0]
+ Tile_X5Y2_LUT4AB/S2MID[1] Tile_X5Y2_LUT4AB/S2MID[2] Tile_X5Y2_LUT4AB/S2MID[3] Tile_X5Y2_LUT4AB/S2MID[4]
+ Tile_X5Y2_LUT4AB/S2MID[5] Tile_X5Y2_LUT4AB/S2MID[6] Tile_X5Y2_LUT4AB/S2MID[7] Tile_X5Y2_LUT4AB/S2END[0]
+ Tile_X5Y2_LUT4AB/S2END[1] Tile_X5Y2_LUT4AB/S2END[2] Tile_X5Y2_LUT4AB/S2END[3] Tile_X5Y2_LUT4AB/S2END[4]
+ Tile_X5Y2_LUT4AB/S2END[5] Tile_X5Y2_LUT4AB/S2END[6] Tile_X5Y2_LUT4AB/S2END[7] Tile_X5Y1_LUT4AB/S2END[0]
+ Tile_X5Y1_LUT4AB/S2END[1] Tile_X5Y1_LUT4AB/S2END[2] Tile_X5Y1_LUT4AB/S2END[3] Tile_X5Y1_LUT4AB/S2END[4]
+ Tile_X5Y1_LUT4AB/S2END[5] Tile_X5Y1_LUT4AB/S2END[6] Tile_X5Y1_LUT4AB/S2END[7] Tile_X5Y1_LUT4AB/S2MID[0]
+ Tile_X5Y1_LUT4AB/S2MID[1] Tile_X5Y1_LUT4AB/S2MID[2] Tile_X5Y1_LUT4AB/S2MID[3] Tile_X5Y1_LUT4AB/S2MID[4]
+ Tile_X5Y1_LUT4AB/S2MID[5] Tile_X5Y1_LUT4AB/S2MID[6] Tile_X5Y1_LUT4AB/S2MID[7] Tile_X5Y2_LUT4AB/S4END[0]
+ Tile_X5Y2_LUT4AB/S4END[10] Tile_X5Y2_LUT4AB/S4END[11] Tile_X5Y2_LUT4AB/S4END[12]
+ Tile_X5Y2_LUT4AB/S4END[13] Tile_X5Y2_LUT4AB/S4END[14] Tile_X5Y2_LUT4AB/S4END[15]
+ Tile_X5Y2_LUT4AB/S4END[1] Tile_X5Y2_LUT4AB/S4END[2] Tile_X5Y2_LUT4AB/S4END[3] Tile_X5Y2_LUT4AB/S4END[4]
+ Tile_X5Y2_LUT4AB/S4END[5] Tile_X5Y2_LUT4AB/S4END[6] Tile_X5Y2_LUT4AB/S4END[7] Tile_X5Y2_LUT4AB/S4END[8]
+ Tile_X5Y2_LUT4AB/S4END[9] Tile_X5Y1_LUT4AB/S4END[0] Tile_X5Y1_LUT4AB/S4END[10] Tile_X5Y1_LUT4AB/S4END[11]
+ Tile_X5Y1_LUT4AB/S4END[12] Tile_X5Y1_LUT4AB/S4END[13] Tile_X5Y1_LUT4AB/S4END[14]
+ Tile_X5Y1_LUT4AB/S4END[15] Tile_X5Y1_LUT4AB/S4END[1] Tile_X5Y1_LUT4AB/S4END[2] Tile_X5Y1_LUT4AB/S4END[3]
+ Tile_X5Y1_LUT4AB/S4END[4] Tile_X5Y1_LUT4AB/S4END[5] Tile_X5Y1_LUT4AB/S4END[6] Tile_X5Y1_LUT4AB/S4END[7]
+ Tile_X5Y1_LUT4AB/S4END[8] Tile_X5Y1_LUT4AB/S4END[9] Tile_X5Y2_LUT4AB/SS4END[0] Tile_X5Y2_LUT4AB/SS4END[10]
+ Tile_X5Y2_LUT4AB/SS4END[11] Tile_X5Y2_LUT4AB/SS4END[12] Tile_X5Y2_LUT4AB/SS4END[13]
+ Tile_X5Y2_LUT4AB/SS4END[14] Tile_X5Y2_LUT4AB/SS4END[15] Tile_X5Y2_LUT4AB/SS4END[1]
+ Tile_X5Y2_LUT4AB/SS4END[2] Tile_X5Y2_LUT4AB/SS4END[3] Tile_X5Y2_LUT4AB/SS4END[4]
+ Tile_X5Y2_LUT4AB/SS4END[5] Tile_X5Y2_LUT4AB/SS4END[6] Tile_X5Y2_LUT4AB/SS4END[7]
+ Tile_X5Y2_LUT4AB/SS4END[8] Tile_X5Y2_LUT4AB/SS4END[9] Tile_X5Y1_LUT4AB/SS4END[0]
+ Tile_X5Y1_LUT4AB/SS4END[10] Tile_X5Y1_LUT4AB/SS4END[11] Tile_X5Y1_LUT4AB/SS4END[12]
+ Tile_X5Y1_LUT4AB/SS4END[13] Tile_X5Y1_LUT4AB/SS4END[14] Tile_X5Y1_LUT4AB/SS4END[15]
+ Tile_X5Y1_LUT4AB/SS4END[1] Tile_X5Y1_LUT4AB/SS4END[2] Tile_X5Y1_LUT4AB/SS4END[3]
+ Tile_X5Y1_LUT4AB/SS4END[4] Tile_X5Y1_LUT4AB/SS4END[5] Tile_X5Y1_LUT4AB/SS4END[6]
+ Tile_X5Y1_LUT4AB/SS4END[7] Tile_X5Y1_LUT4AB/SS4END[8] Tile_X5Y1_LUT4AB/SS4END[9]
+ Tile_X5Y1_LUT4AB/UserCLK Tile_X5Y1_LUT4AB/UserCLKo VGND VPWR Tile_X5Y1_LUT4AB/W1BEG[0]
+ Tile_X5Y1_LUT4AB/W1BEG[1] Tile_X5Y1_LUT4AB/W1BEG[2] Tile_X5Y1_LUT4AB/W1BEG[3] Tile_X6Y1_LUT4AB/W1BEG[0]
+ Tile_X6Y1_LUT4AB/W1BEG[1] Tile_X6Y1_LUT4AB/W1BEG[2] Tile_X6Y1_LUT4AB/W1BEG[3] Tile_X5Y1_LUT4AB/W2BEG[0]
+ Tile_X5Y1_LUT4AB/W2BEG[1] Tile_X5Y1_LUT4AB/W2BEG[2] Tile_X5Y1_LUT4AB/W2BEG[3] Tile_X5Y1_LUT4AB/W2BEG[4]
+ Tile_X5Y1_LUT4AB/W2BEG[5] Tile_X5Y1_LUT4AB/W2BEG[6] Tile_X5Y1_LUT4AB/W2BEG[7] Tile_X5Y1_LUT4AB/W2BEGb[0]
+ Tile_X5Y1_LUT4AB/W2BEGb[1] Tile_X5Y1_LUT4AB/W2BEGb[2] Tile_X5Y1_LUT4AB/W2BEGb[3]
+ Tile_X5Y1_LUT4AB/W2BEGb[4] Tile_X5Y1_LUT4AB/W2BEGb[5] Tile_X5Y1_LUT4AB/W2BEGb[6]
+ Tile_X5Y1_LUT4AB/W2BEGb[7] Tile_X5Y1_LUT4AB/W2END[0] Tile_X5Y1_LUT4AB/W2END[1] Tile_X5Y1_LUT4AB/W2END[2]
+ Tile_X5Y1_LUT4AB/W2END[3] Tile_X5Y1_LUT4AB/W2END[4] Tile_X5Y1_LUT4AB/W2END[5] Tile_X5Y1_LUT4AB/W2END[6]
+ Tile_X5Y1_LUT4AB/W2END[7] Tile_X6Y1_LUT4AB/W2BEG[0] Tile_X6Y1_LUT4AB/W2BEG[1] Tile_X6Y1_LUT4AB/W2BEG[2]
+ Tile_X6Y1_LUT4AB/W2BEG[3] Tile_X6Y1_LUT4AB/W2BEG[4] Tile_X6Y1_LUT4AB/W2BEG[5] Tile_X6Y1_LUT4AB/W2BEG[6]
+ Tile_X6Y1_LUT4AB/W2BEG[7] Tile_X5Y1_LUT4AB/W6BEG[0] Tile_X5Y1_LUT4AB/W6BEG[10] Tile_X5Y1_LUT4AB/W6BEG[11]
+ Tile_X5Y1_LUT4AB/W6BEG[1] Tile_X5Y1_LUT4AB/W6BEG[2] Tile_X5Y1_LUT4AB/W6BEG[3] Tile_X5Y1_LUT4AB/W6BEG[4]
+ Tile_X5Y1_LUT4AB/W6BEG[5] Tile_X5Y1_LUT4AB/W6BEG[6] Tile_X5Y1_LUT4AB/W6BEG[7] Tile_X5Y1_LUT4AB/W6BEG[8]
+ Tile_X5Y1_LUT4AB/W6BEG[9] Tile_X6Y1_LUT4AB/W6BEG[0] Tile_X6Y1_LUT4AB/W6BEG[10] Tile_X6Y1_LUT4AB/W6BEG[11]
+ Tile_X6Y1_LUT4AB/W6BEG[1] Tile_X6Y1_LUT4AB/W6BEG[2] Tile_X6Y1_LUT4AB/W6BEG[3] Tile_X6Y1_LUT4AB/W6BEG[4]
+ Tile_X6Y1_LUT4AB/W6BEG[5] Tile_X6Y1_LUT4AB/W6BEG[6] Tile_X6Y1_LUT4AB/W6BEG[7] Tile_X6Y1_LUT4AB/W6BEG[8]
+ Tile_X6Y1_LUT4AB/W6BEG[9] Tile_X5Y1_LUT4AB/WW4BEG[0] Tile_X5Y1_LUT4AB/WW4BEG[10]
+ Tile_X5Y1_LUT4AB/WW4BEG[11] Tile_X5Y1_LUT4AB/WW4BEG[12] Tile_X5Y1_LUT4AB/WW4BEG[13]
+ Tile_X5Y1_LUT4AB/WW4BEG[14] Tile_X5Y1_LUT4AB/WW4BEG[15] Tile_X5Y1_LUT4AB/WW4BEG[1]
+ Tile_X5Y1_LUT4AB/WW4BEG[2] Tile_X5Y1_LUT4AB/WW4BEG[3] Tile_X5Y1_LUT4AB/WW4BEG[4]
+ Tile_X5Y1_LUT4AB/WW4BEG[5] Tile_X5Y1_LUT4AB/WW4BEG[6] Tile_X5Y1_LUT4AB/WW4BEG[7]
+ Tile_X5Y1_LUT4AB/WW4BEG[8] Tile_X5Y1_LUT4AB/WW4BEG[9] Tile_X6Y1_LUT4AB/WW4BEG[0]
+ Tile_X6Y1_LUT4AB/WW4BEG[10] Tile_X6Y1_LUT4AB/WW4BEG[11] Tile_X6Y1_LUT4AB/WW4BEG[12]
+ Tile_X6Y1_LUT4AB/WW4BEG[13] Tile_X6Y1_LUT4AB/WW4BEG[14] Tile_X6Y1_LUT4AB/WW4BEG[15]
+ Tile_X6Y1_LUT4AB/WW4BEG[1] Tile_X6Y1_LUT4AB/WW4BEG[2] Tile_X6Y1_LUT4AB/WW4BEG[3]
+ Tile_X6Y1_LUT4AB/WW4BEG[4] Tile_X6Y1_LUT4AB/WW4BEG[5] Tile_X6Y1_LUT4AB/WW4BEG[6]
+ Tile_X6Y1_LUT4AB/WW4BEG[7] Tile_X6Y1_LUT4AB/WW4BEG[8] Tile_X6Y1_LUT4AB/WW4BEG[9]
+ LUT4AB
XTile_X9Y13_LUT4AB Tile_X9Y14_LUT4AB/Co Tile_X9Y13_LUT4AB/Co Tile_X9Y13_LUT4AB/E1BEG[0]
+ Tile_X9Y13_LUT4AB/E1BEG[1] Tile_X9Y13_LUT4AB/E1BEG[2] Tile_X9Y13_LUT4AB/E1BEG[3]
+ Tile_X9Y13_LUT4AB/E1END[0] Tile_X9Y13_LUT4AB/E1END[1] Tile_X9Y13_LUT4AB/E1END[2]
+ Tile_X9Y13_LUT4AB/E1END[3] Tile_X9Y13_LUT4AB/E2BEG[0] Tile_X9Y13_LUT4AB/E2BEG[1]
+ Tile_X9Y13_LUT4AB/E2BEG[2] Tile_X9Y13_LUT4AB/E2BEG[3] Tile_X9Y13_LUT4AB/E2BEG[4]
+ Tile_X9Y13_LUT4AB/E2BEG[5] Tile_X9Y13_LUT4AB/E2BEG[6] Tile_X9Y13_LUT4AB/E2BEG[7]
+ Tile_X9Y13_LUT4AB/E2BEGb[0] Tile_X9Y13_LUT4AB/E2BEGb[1] Tile_X9Y13_LUT4AB/E2BEGb[2]
+ Tile_X9Y13_LUT4AB/E2BEGb[3] Tile_X9Y13_LUT4AB/E2BEGb[4] Tile_X9Y13_LUT4AB/E2BEGb[5]
+ Tile_X9Y13_LUT4AB/E2BEGb[6] Tile_X9Y13_LUT4AB/E2BEGb[7] Tile_X9Y13_LUT4AB/E2END[0]
+ Tile_X9Y13_LUT4AB/E2END[1] Tile_X9Y13_LUT4AB/E2END[2] Tile_X9Y13_LUT4AB/E2END[3]
+ Tile_X9Y13_LUT4AB/E2END[4] Tile_X9Y13_LUT4AB/E2END[5] Tile_X9Y13_LUT4AB/E2END[6]
+ Tile_X9Y13_LUT4AB/E2END[7] Tile_X9Y13_LUT4AB/E2MID[0] Tile_X9Y13_LUT4AB/E2MID[1]
+ Tile_X9Y13_LUT4AB/E2MID[2] Tile_X9Y13_LUT4AB/E2MID[3] Tile_X9Y13_LUT4AB/E2MID[4]
+ Tile_X9Y13_LUT4AB/E2MID[5] Tile_X9Y13_LUT4AB/E2MID[6] Tile_X9Y13_LUT4AB/E2MID[7]
+ Tile_X9Y13_LUT4AB/E6BEG[0] Tile_X9Y13_LUT4AB/E6BEG[10] Tile_X9Y13_LUT4AB/E6BEG[11]
+ Tile_X9Y13_LUT4AB/E6BEG[1] Tile_X9Y13_LUT4AB/E6BEG[2] Tile_X9Y13_LUT4AB/E6BEG[3]
+ Tile_X9Y13_LUT4AB/E6BEG[4] Tile_X9Y13_LUT4AB/E6BEG[5] Tile_X9Y13_LUT4AB/E6BEG[6]
+ Tile_X9Y13_LUT4AB/E6BEG[7] Tile_X9Y13_LUT4AB/E6BEG[8] Tile_X9Y13_LUT4AB/E6BEG[9]
+ Tile_X9Y13_LUT4AB/E6END[0] Tile_X9Y13_LUT4AB/E6END[10] Tile_X9Y13_LUT4AB/E6END[11]
+ Tile_X9Y13_LUT4AB/E6END[1] Tile_X9Y13_LUT4AB/E6END[2] Tile_X9Y13_LUT4AB/E6END[3]
+ Tile_X9Y13_LUT4AB/E6END[4] Tile_X9Y13_LUT4AB/E6END[5] Tile_X9Y13_LUT4AB/E6END[6]
+ Tile_X9Y13_LUT4AB/E6END[7] Tile_X9Y13_LUT4AB/E6END[8] Tile_X9Y13_LUT4AB/E6END[9]
+ Tile_X9Y13_LUT4AB/EE4BEG[0] Tile_X9Y13_LUT4AB/EE4BEG[10] Tile_X9Y13_LUT4AB/EE4BEG[11]
+ Tile_X9Y13_LUT4AB/EE4BEG[12] Tile_X9Y13_LUT4AB/EE4BEG[13] Tile_X9Y13_LUT4AB/EE4BEG[14]
+ Tile_X9Y13_LUT4AB/EE4BEG[15] Tile_X9Y13_LUT4AB/EE4BEG[1] Tile_X9Y13_LUT4AB/EE4BEG[2]
+ Tile_X9Y13_LUT4AB/EE4BEG[3] Tile_X9Y13_LUT4AB/EE4BEG[4] Tile_X9Y13_LUT4AB/EE4BEG[5]
+ Tile_X9Y13_LUT4AB/EE4BEG[6] Tile_X9Y13_LUT4AB/EE4BEG[7] Tile_X9Y13_LUT4AB/EE4BEG[8]
+ Tile_X9Y13_LUT4AB/EE4BEG[9] Tile_X9Y13_LUT4AB/EE4END[0] Tile_X9Y13_LUT4AB/EE4END[10]
+ Tile_X9Y13_LUT4AB/EE4END[11] Tile_X9Y13_LUT4AB/EE4END[12] Tile_X9Y13_LUT4AB/EE4END[13]
+ Tile_X9Y13_LUT4AB/EE4END[14] Tile_X9Y13_LUT4AB/EE4END[15] Tile_X9Y13_LUT4AB/EE4END[1]
+ Tile_X9Y13_LUT4AB/EE4END[2] Tile_X9Y13_LUT4AB/EE4END[3] Tile_X9Y13_LUT4AB/EE4END[4]
+ Tile_X9Y13_LUT4AB/EE4END[5] Tile_X9Y13_LUT4AB/EE4END[6] Tile_X9Y13_LUT4AB/EE4END[7]
+ Tile_X9Y13_LUT4AB/EE4END[8] Tile_X9Y13_LUT4AB/EE4END[9] Tile_X9Y13_LUT4AB/FrameData[0]
+ Tile_X9Y13_LUT4AB/FrameData[10] Tile_X9Y13_LUT4AB/FrameData[11] Tile_X9Y13_LUT4AB/FrameData[12]
+ Tile_X9Y13_LUT4AB/FrameData[13] Tile_X9Y13_LUT4AB/FrameData[14] Tile_X9Y13_LUT4AB/FrameData[15]
+ Tile_X9Y13_LUT4AB/FrameData[16] Tile_X9Y13_LUT4AB/FrameData[17] Tile_X9Y13_LUT4AB/FrameData[18]
+ Tile_X9Y13_LUT4AB/FrameData[19] Tile_X9Y13_LUT4AB/FrameData[1] Tile_X9Y13_LUT4AB/FrameData[20]
+ Tile_X9Y13_LUT4AB/FrameData[21] Tile_X9Y13_LUT4AB/FrameData[22] Tile_X9Y13_LUT4AB/FrameData[23]
+ Tile_X9Y13_LUT4AB/FrameData[24] Tile_X9Y13_LUT4AB/FrameData[25] Tile_X9Y13_LUT4AB/FrameData[26]
+ Tile_X9Y13_LUT4AB/FrameData[27] Tile_X9Y13_LUT4AB/FrameData[28] Tile_X9Y13_LUT4AB/FrameData[29]
+ Tile_X9Y13_LUT4AB/FrameData[2] Tile_X9Y13_LUT4AB/FrameData[30] Tile_X9Y13_LUT4AB/FrameData[31]
+ Tile_X9Y13_LUT4AB/FrameData[3] Tile_X9Y13_LUT4AB/FrameData[4] Tile_X9Y13_LUT4AB/FrameData[5]
+ Tile_X9Y13_LUT4AB/FrameData[6] Tile_X9Y13_LUT4AB/FrameData[7] Tile_X9Y13_LUT4AB/FrameData[8]
+ Tile_X9Y13_LUT4AB/FrameData[9] Tile_X9Y13_LUT4AB/FrameData_O[0] Tile_X9Y13_LUT4AB/FrameData_O[10]
+ Tile_X9Y13_LUT4AB/FrameData_O[11] Tile_X9Y13_LUT4AB/FrameData_O[12] Tile_X9Y13_LUT4AB/FrameData_O[13]
+ Tile_X9Y13_LUT4AB/FrameData_O[14] Tile_X9Y13_LUT4AB/FrameData_O[15] Tile_X9Y13_LUT4AB/FrameData_O[16]
+ Tile_X9Y13_LUT4AB/FrameData_O[17] Tile_X9Y13_LUT4AB/FrameData_O[18] Tile_X9Y13_LUT4AB/FrameData_O[19]
+ Tile_X9Y13_LUT4AB/FrameData_O[1] Tile_X9Y13_LUT4AB/FrameData_O[20] Tile_X9Y13_LUT4AB/FrameData_O[21]
+ Tile_X9Y13_LUT4AB/FrameData_O[22] Tile_X9Y13_LUT4AB/FrameData_O[23] Tile_X9Y13_LUT4AB/FrameData_O[24]
+ Tile_X9Y13_LUT4AB/FrameData_O[25] Tile_X9Y13_LUT4AB/FrameData_O[26] Tile_X9Y13_LUT4AB/FrameData_O[27]
+ Tile_X9Y13_LUT4AB/FrameData_O[28] Tile_X9Y13_LUT4AB/FrameData_O[29] Tile_X9Y13_LUT4AB/FrameData_O[2]
+ Tile_X9Y13_LUT4AB/FrameData_O[30] Tile_X9Y13_LUT4AB/FrameData_O[31] Tile_X9Y13_LUT4AB/FrameData_O[3]
+ Tile_X9Y13_LUT4AB/FrameData_O[4] Tile_X9Y13_LUT4AB/FrameData_O[5] Tile_X9Y13_LUT4AB/FrameData_O[6]
+ Tile_X9Y13_LUT4AB/FrameData_O[7] Tile_X9Y13_LUT4AB/FrameData_O[8] Tile_X9Y13_LUT4AB/FrameData_O[9]
+ Tile_X9Y13_LUT4AB/FrameStrobe[0] Tile_X9Y13_LUT4AB/FrameStrobe[10] Tile_X9Y13_LUT4AB/FrameStrobe[11]
+ Tile_X9Y13_LUT4AB/FrameStrobe[12] Tile_X9Y13_LUT4AB/FrameStrobe[13] Tile_X9Y13_LUT4AB/FrameStrobe[14]
+ Tile_X9Y13_LUT4AB/FrameStrobe[15] Tile_X9Y13_LUT4AB/FrameStrobe[16] Tile_X9Y13_LUT4AB/FrameStrobe[17]
+ Tile_X9Y13_LUT4AB/FrameStrobe[18] Tile_X9Y13_LUT4AB/FrameStrobe[19] Tile_X9Y13_LUT4AB/FrameStrobe[1]
+ Tile_X9Y13_LUT4AB/FrameStrobe[2] Tile_X9Y13_LUT4AB/FrameStrobe[3] Tile_X9Y13_LUT4AB/FrameStrobe[4]
+ Tile_X9Y13_LUT4AB/FrameStrobe[5] Tile_X9Y13_LUT4AB/FrameStrobe[6] Tile_X9Y13_LUT4AB/FrameStrobe[7]
+ Tile_X9Y13_LUT4AB/FrameStrobe[8] Tile_X9Y13_LUT4AB/FrameStrobe[9] Tile_X9Y12_LUT4AB/FrameStrobe[0]
+ Tile_X9Y12_LUT4AB/FrameStrobe[10] Tile_X9Y12_LUT4AB/FrameStrobe[11] Tile_X9Y12_LUT4AB/FrameStrobe[12]
+ Tile_X9Y12_LUT4AB/FrameStrobe[13] Tile_X9Y12_LUT4AB/FrameStrobe[14] Tile_X9Y12_LUT4AB/FrameStrobe[15]
+ Tile_X9Y12_LUT4AB/FrameStrobe[16] Tile_X9Y12_LUT4AB/FrameStrobe[17] Tile_X9Y12_LUT4AB/FrameStrobe[18]
+ Tile_X9Y12_LUT4AB/FrameStrobe[19] Tile_X9Y12_LUT4AB/FrameStrobe[1] Tile_X9Y12_LUT4AB/FrameStrobe[2]
+ Tile_X9Y12_LUT4AB/FrameStrobe[3] Tile_X9Y12_LUT4AB/FrameStrobe[4] Tile_X9Y12_LUT4AB/FrameStrobe[5]
+ Tile_X9Y12_LUT4AB/FrameStrobe[6] Tile_X9Y12_LUT4AB/FrameStrobe[7] Tile_X9Y12_LUT4AB/FrameStrobe[8]
+ Tile_X9Y12_LUT4AB/FrameStrobe[9] Tile_X9Y13_LUT4AB/N1BEG[0] Tile_X9Y13_LUT4AB/N1BEG[1]
+ Tile_X9Y13_LUT4AB/N1BEG[2] Tile_X9Y13_LUT4AB/N1BEG[3] Tile_X9Y14_LUT4AB/N1BEG[0]
+ Tile_X9Y14_LUT4AB/N1BEG[1] Tile_X9Y14_LUT4AB/N1BEG[2] Tile_X9Y14_LUT4AB/N1BEG[3]
+ Tile_X9Y13_LUT4AB/N2BEG[0] Tile_X9Y13_LUT4AB/N2BEG[1] Tile_X9Y13_LUT4AB/N2BEG[2]
+ Tile_X9Y13_LUT4AB/N2BEG[3] Tile_X9Y13_LUT4AB/N2BEG[4] Tile_X9Y13_LUT4AB/N2BEG[5]
+ Tile_X9Y13_LUT4AB/N2BEG[6] Tile_X9Y13_LUT4AB/N2BEG[7] Tile_X9Y12_LUT4AB/N2END[0]
+ Tile_X9Y12_LUT4AB/N2END[1] Tile_X9Y12_LUT4AB/N2END[2] Tile_X9Y12_LUT4AB/N2END[3]
+ Tile_X9Y12_LUT4AB/N2END[4] Tile_X9Y12_LUT4AB/N2END[5] Tile_X9Y12_LUT4AB/N2END[6]
+ Tile_X9Y12_LUT4AB/N2END[7] Tile_X9Y13_LUT4AB/N2END[0] Tile_X9Y13_LUT4AB/N2END[1]
+ Tile_X9Y13_LUT4AB/N2END[2] Tile_X9Y13_LUT4AB/N2END[3] Tile_X9Y13_LUT4AB/N2END[4]
+ Tile_X9Y13_LUT4AB/N2END[5] Tile_X9Y13_LUT4AB/N2END[6] Tile_X9Y13_LUT4AB/N2END[7]
+ Tile_X9Y14_LUT4AB/N2BEG[0] Tile_X9Y14_LUT4AB/N2BEG[1] Tile_X9Y14_LUT4AB/N2BEG[2]
+ Tile_X9Y14_LUT4AB/N2BEG[3] Tile_X9Y14_LUT4AB/N2BEG[4] Tile_X9Y14_LUT4AB/N2BEG[5]
+ Tile_X9Y14_LUT4AB/N2BEG[6] Tile_X9Y14_LUT4AB/N2BEG[7] Tile_X9Y13_LUT4AB/N4BEG[0]
+ Tile_X9Y13_LUT4AB/N4BEG[10] Tile_X9Y13_LUT4AB/N4BEG[11] Tile_X9Y13_LUT4AB/N4BEG[12]
+ Tile_X9Y13_LUT4AB/N4BEG[13] Tile_X9Y13_LUT4AB/N4BEG[14] Tile_X9Y13_LUT4AB/N4BEG[15]
+ Tile_X9Y13_LUT4AB/N4BEG[1] Tile_X9Y13_LUT4AB/N4BEG[2] Tile_X9Y13_LUT4AB/N4BEG[3]
+ Tile_X9Y13_LUT4AB/N4BEG[4] Tile_X9Y13_LUT4AB/N4BEG[5] Tile_X9Y13_LUT4AB/N4BEG[6]
+ Tile_X9Y13_LUT4AB/N4BEG[7] Tile_X9Y13_LUT4AB/N4BEG[8] Tile_X9Y13_LUT4AB/N4BEG[9]
+ Tile_X9Y14_LUT4AB/N4BEG[0] Tile_X9Y14_LUT4AB/N4BEG[10] Tile_X9Y14_LUT4AB/N4BEG[11]
+ Tile_X9Y14_LUT4AB/N4BEG[12] Tile_X9Y14_LUT4AB/N4BEG[13] Tile_X9Y14_LUT4AB/N4BEG[14]
+ Tile_X9Y14_LUT4AB/N4BEG[15] Tile_X9Y14_LUT4AB/N4BEG[1] Tile_X9Y14_LUT4AB/N4BEG[2]
+ Tile_X9Y14_LUT4AB/N4BEG[3] Tile_X9Y14_LUT4AB/N4BEG[4] Tile_X9Y14_LUT4AB/N4BEG[5]
+ Tile_X9Y14_LUT4AB/N4BEG[6] Tile_X9Y14_LUT4AB/N4BEG[7] Tile_X9Y14_LUT4AB/N4BEG[8]
+ Tile_X9Y14_LUT4AB/N4BEG[9] Tile_X9Y13_LUT4AB/NN4BEG[0] Tile_X9Y13_LUT4AB/NN4BEG[10]
+ Tile_X9Y13_LUT4AB/NN4BEG[11] Tile_X9Y13_LUT4AB/NN4BEG[12] Tile_X9Y13_LUT4AB/NN4BEG[13]
+ Tile_X9Y13_LUT4AB/NN4BEG[14] Tile_X9Y13_LUT4AB/NN4BEG[15] Tile_X9Y13_LUT4AB/NN4BEG[1]
+ Tile_X9Y13_LUT4AB/NN4BEG[2] Tile_X9Y13_LUT4AB/NN4BEG[3] Tile_X9Y13_LUT4AB/NN4BEG[4]
+ Tile_X9Y13_LUT4AB/NN4BEG[5] Tile_X9Y13_LUT4AB/NN4BEG[6] Tile_X9Y13_LUT4AB/NN4BEG[7]
+ Tile_X9Y13_LUT4AB/NN4BEG[8] Tile_X9Y13_LUT4AB/NN4BEG[9] Tile_X9Y14_LUT4AB/NN4BEG[0]
+ Tile_X9Y14_LUT4AB/NN4BEG[10] Tile_X9Y14_LUT4AB/NN4BEG[11] Tile_X9Y14_LUT4AB/NN4BEG[12]
+ Tile_X9Y14_LUT4AB/NN4BEG[13] Tile_X9Y14_LUT4AB/NN4BEG[14] Tile_X9Y14_LUT4AB/NN4BEG[15]
+ Tile_X9Y14_LUT4AB/NN4BEG[1] Tile_X9Y14_LUT4AB/NN4BEG[2] Tile_X9Y14_LUT4AB/NN4BEG[3]
+ Tile_X9Y14_LUT4AB/NN4BEG[4] Tile_X9Y14_LUT4AB/NN4BEG[5] Tile_X9Y14_LUT4AB/NN4BEG[6]
+ Tile_X9Y14_LUT4AB/NN4BEG[7] Tile_X9Y14_LUT4AB/NN4BEG[8] Tile_X9Y14_LUT4AB/NN4BEG[9]
+ Tile_X9Y14_LUT4AB/S1END[0] Tile_X9Y14_LUT4AB/S1END[1] Tile_X9Y14_LUT4AB/S1END[2]
+ Tile_X9Y14_LUT4AB/S1END[3] Tile_X9Y13_LUT4AB/S1END[0] Tile_X9Y13_LUT4AB/S1END[1]
+ Tile_X9Y13_LUT4AB/S1END[2] Tile_X9Y13_LUT4AB/S1END[3] Tile_X9Y14_LUT4AB/S2MID[0]
+ Tile_X9Y14_LUT4AB/S2MID[1] Tile_X9Y14_LUT4AB/S2MID[2] Tile_X9Y14_LUT4AB/S2MID[3]
+ Tile_X9Y14_LUT4AB/S2MID[4] Tile_X9Y14_LUT4AB/S2MID[5] Tile_X9Y14_LUT4AB/S2MID[6]
+ Tile_X9Y14_LUT4AB/S2MID[7] Tile_X9Y14_LUT4AB/S2END[0] Tile_X9Y14_LUT4AB/S2END[1]
+ Tile_X9Y14_LUT4AB/S2END[2] Tile_X9Y14_LUT4AB/S2END[3] Tile_X9Y14_LUT4AB/S2END[4]
+ Tile_X9Y14_LUT4AB/S2END[5] Tile_X9Y14_LUT4AB/S2END[6] Tile_X9Y14_LUT4AB/S2END[7]
+ Tile_X9Y13_LUT4AB/S2END[0] Tile_X9Y13_LUT4AB/S2END[1] Tile_X9Y13_LUT4AB/S2END[2]
+ Tile_X9Y13_LUT4AB/S2END[3] Tile_X9Y13_LUT4AB/S2END[4] Tile_X9Y13_LUT4AB/S2END[5]
+ Tile_X9Y13_LUT4AB/S2END[6] Tile_X9Y13_LUT4AB/S2END[7] Tile_X9Y13_LUT4AB/S2MID[0]
+ Tile_X9Y13_LUT4AB/S2MID[1] Tile_X9Y13_LUT4AB/S2MID[2] Tile_X9Y13_LUT4AB/S2MID[3]
+ Tile_X9Y13_LUT4AB/S2MID[4] Tile_X9Y13_LUT4AB/S2MID[5] Tile_X9Y13_LUT4AB/S2MID[6]
+ Tile_X9Y13_LUT4AB/S2MID[7] Tile_X9Y14_LUT4AB/S4END[0] Tile_X9Y14_LUT4AB/S4END[10]
+ Tile_X9Y14_LUT4AB/S4END[11] Tile_X9Y14_LUT4AB/S4END[12] Tile_X9Y14_LUT4AB/S4END[13]
+ Tile_X9Y14_LUT4AB/S4END[14] Tile_X9Y14_LUT4AB/S4END[15] Tile_X9Y14_LUT4AB/S4END[1]
+ Tile_X9Y14_LUT4AB/S4END[2] Tile_X9Y14_LUT4AB/S4END[3] Tile_X9Y14_LUT4AB/S4END[4]
+ Tile_X9Y14_LUT4AB/S4END[5] Tile_X9Y14_LUT4AB/S4END[6] Tile_X9Y14_LUT4AB/S4END[7]
+ Tile_X9Y14_LUT4AB/S4END[8] Tile_X9Y14_LUT4AB/S4END[9] Tile_X9Y13_LUT4AB/S4END[0]
+ Tile_X9Y13_LUT4AB/S4END[10] Tile_X9Y13_LUT4AB/S4END[11] Tile_X9Y13_LUT4AB/S4END[12]
+ Tile_X9Y13_LUT4AB/S4END[13] Tile_X9Y13_LUT4AB/S4END[14] Tile_X9Y13_LUT4AB/S4END[15]
+ Tile_X9Y13_LUT4AB/S4END[1] Tile_X9Y13_LUT4AB/S4END[2] Tile_X9Y13_LUT4AB/S4END[3]
+ Tile_X9Y13_LUT4AB/S4END[4] Tile_X9Y13_LUT4AB/S4END[5] Tile_X9Y13_LUT4AB/S4END[6]
+ Tile_X9Y13_LUT4AB/S4END[7] Tile_X9Y13_LUT4AB/S4END[8] Tile_X9Y13_LUT4AB/S4END[9]
+ Tile_X9Y14_LUT4AB/SS4END[0] Tile_X9Y14_LUT4AB/SS4END[10] Tile_X9Y14_LUT4AB/SS4END[11]
+ Tile_X9Y14_LUT4AB/SS4END[12] Tile_X9Y14_LUT4AB/SS4END[13] Tile_X9Y14_LUT4AB/SS4END[14]
+ Tile_X9Y14_LUT4AB/SS4END[15] Tile_X9Y14_LUT4AB/SS4END[1] Tile_X9Y14_LUT4AB/SS4END[2]
+ Tile_X9Y14_LUT4AB/SS4END[3] Tile_X9Y14_LUT4AB/SS4END[4] Tile_X9Y14_LUT4AB/SS4END[5]
+ Tile_X9Y14_LUT4AB/SS4END[6] Tile_X9Y14_LUT4AB/SS4END[7] Tile_X9Y14_LUT4AB/SS4END[8]
+ Tile_X9Y14_LUT4AB/SS4END[9] Tile_X9Y13_LUT4AB/SS4END[0] Tile_X9Y13_LUT4AB/SS4END[10]
+ Tile_X9Y13_LUT4AB/SS4END[11] Tile_X9Y13_LUT4AB/SS4END[12] Tile_X9Y13_LUT4AB/SS4END[13]
+ Tile_X9Y13_LUT4AB/SS4END[14] Tile_X9Y13_LUT4AB/SS4END[15] Tile_X9Y13_LUT4AB/SS4END[1]
+ Tile_X9Y13_LUT4AB/SS4END[2] Tile_X9Y13_LUT4AB/SS4END[3] Tile_X9Y13_LUT4AB/SS4END[4]
+ Tile_X9Y13_LUT4AB/SS4END[5] Tile_X9Y13_LUT4AB/SS4END[6] Tile_X9Y13_LUT4AB/SS4END[7]
+ Tile_X9Y13_LUT4AB/SS4END[8] Tile_X9Y13_LUT4AB/SS4END[9] Tile_X9Y13_LUT4AB/UserCLK
+ Tile_X9Y12_LUT4AB/UserCLK VGND VPWR Tile_X9Y13_LUT4AB/W1BEG[0] Tile_X9Y13_LUT4AB/W1BEG[1]
+ Tile_X9Y13_LUT4AB/W1BEG[2] Tile_X9Y13_LUT4AB/W1BEG[3] Tile_X9Y13_LUT4AB/W1END[0]
+ Tile_X9Y13_LUT4AB/W1END[1] Tile_X9Y13_LUT4AB/W1END[2] Tile_X9Y13_LUT4AB/W1END[3]
+ Tile_X9Y13_LUT4AB/W2BEG[0] Tile_X9Y13_LUT4AB/W2BEG[1] Tile_X9Y13_LUT4AB/W2BEG[2]
+ Tile_X9Y13_LUT4AB/W2BEG[3] Tile_X9Y13_LUT4AB/W2BEG[4] Tile_X9Y13_LUT4AB/W2BEG[5]
+ Tile_X9Y13_LUT4AB/W2BEG[6] Tile_X9Y13_LUT4AB/W2BEG[7] Tile_X8Y13_LUT4AB/W2END[0]
+ Tile_X8Y13_LUT4AB/W2END[1] Tile_X8Y13_LUT4AB/W2END[2] Tile_X8Y13_LUT4AB/W2END[3]
+ Tile_X8Y13_LUT4AB/W2END[4] Tile_X8Y13_LUT4AB/W2END[5] Tile_X8Y13_LUT4AB/W2END[6]
+ Tile_X8Y13_LUT4AB/W2END[7] Tile_X9Y13_LUT4AB/W2END[0] Tile_X9Y13_LUT4AB/W2END[1]
+ Tile_X9Y13_LUT4AB/W2END[2] Tile_X9Y13_LUT4AB/W2END[3] Tile_X9Y13_LUT4AB/W2END[4]
+ Tile_X9Y13_LUT4AB/W2END[5] Tile_X9Y13_LUT4AB/W2END[6] Tile_X9Y13_LUT4AB/W2END[7]
+ Tile_X9Y13_LUT4AB/W2MID[0] Tile_X9Y13_LUT4AB/W2MID[1] Tile_X9Y13_LUT4AB/W2MID[2]
+ Tile_X9Y13_LUT4AB/W2MID[3] Tile_X9Y13_LUT4AB/W2MID[4] Tile_X9Y13_LUT4AB/W2MID[5]
+ Tile_X9Y13_LUT4AB/W2MID[6] Tile_X9Y13_LUT4AB/W2MID[7] Tile_X9Y13_LUT4AB/W6BEG[0]
+ Tile_X9Y13_LUT4AB/W6BEG[10] Tile_X9Y13_LUT4AB/W6BEG[11] Tile_X9Y13_LUT4AB/W6BEG[1]
+ Tile_X9Y13_LUT4AB/W6BEG[2] Tile_X9Y13_LUT4AB/W6BEG[3] Tile_X9Y13_LUT4AB/W6BEG[4]
+ Tile_X9Y13_LUT4AB/W6BEG[5] Tile_X9Y13_LUT4AB/W6BEG[6] Tile_X9Y13_LUT4AB/W6BEG[7]
+ Tile_X9Y13_LUT4AB/W6BEG[8] Tile_X9Y13_LUT4AB/W6BEG[9] Tile_X9Y13_LUT4AB/W6END[0]
+ Tile_X9Y13_LUT4AB/W6END[10] Tile_X9Y13_LUT4AB/W6END[11] Tile_X9Y13_LUT4AB/W6END[1]
+ Tile_X9Y13_LUT4AB/W6END[2] Tile_X9Y13_LUT4AB/W6END[3] Tile_X9Y13_LUT4AB/W6END[4]
+ Tile_X9Y13_LUT4AB/W6END[5] Tile_X9Y13_LUT4AB/W6END[6] Tile_X9Y13_LUT4AB/W6END[7]
+ Tile_X9Y13_LUT4AB/W6END[8] Tile_X9Y13_LUT4AB/W6END[9] Tile_X9Y13_LUT4AB/WW4BEG[0]
+ Tile_X9Y13_LUT4AB/WW4BEG[10] Tile_X9Y13_LUT4AB/WW4BEG[11] Tile_X9Y13_LUT4AB/WW4BEG[12]
+ Tile_X9Y13_LUT4AB/WW4BEG[13] Tile_X9Y13_LUT4AB/WW4BEG[14] Tile_X9Y13_LUT4AB/WW4BEG[15]
+ Tile_X9Y13_LUT4AB/WW4BEG[1] Tile_X9Y13_LUT4AB/WW4BEG[2] Tile_X9Y13_LUT4AB/WW4BEG[3]
+ Tile_X9Y13_LUT4AB/WW4BEG[4] Tile_X9Y13_LUT4AB/WW4BEG[5] Tile_X9Y13_LUT4AB/WW4BEG[6]
+ Tile_X9Y13_LUT4AB/WW4BEG[7] Tile_X9Y13_LUT4AB/WW4BEG[8] Tile_X9Y13_LUT4AB/WW4BEG[9]
+ Tile_X9Y13_LUT4AB/WW4END[0] Tile_X9Y13_LUT4AB/WW4END[10] Tile_X9Y13_LUT4AB/WW4END[11]
+ Tile_X9Y13_LUT4AB/WW4END[12] Tile_X9Y13_LUT4AB/WW4END[13] Tile_X9Y13_LUT4AB/WW4END[14]
+ Tile_X9Y13_LUT4AB/WW4END[15] Tile_X9Y13_LUT4AB/WW4END[1] Tile_X9Y13_LUT4AB/WW4END[2]
+ Tile_X9Y13_LUT4AB/WW4END[3] Tile_X9Y13_LUT4AB/WW4END[4] Tile_X9Y13_LUT4AB/WW4END[5]
+ Tile_X9Y13_LUT4AB/WW4END[6] Tile_X9Y13_LUT4AB/WW4END[7] Tile_X9Y13_LUT4AB/WW4END[8]
+ Tile_X9Y13_LUT4AB/WW4END[9] LUT4AB
XTile_X4Y12_RegFile Tile_X5Y12_LUT4AB/E1END[0] Tile_X5Y12_LUT4AB/E1END[1] Tile_X5Y12_LUT4AB/E1END[2]
+ Tile_X5Y12_LUT4AB/E1END[3] Tile_X3Y12_LUT4AB/E1BEG[0] Tile_X3Y12_LUT4AB/E1BEG[1]
+ Tile_X3Y12_LUT4AB/E1BEG[2] Tile_X3Y12_LUT4AB/E1BEG[3] Tile_X5Y12_LUT4AB/E2MID[0]
+ Tile_X5Y12_LUT4AB/E2MID[1] Tile_X5Y12_LUT4AB/E2MID[2] Tile_X5Y12_LUT4AB/E2MID[3]
+ Tile_X5Y12_LUT4AB/E2MID[4] Tile_X5Y12_LUT4AB/E2MID[5] Tile_X5Y12_LUT4AB/E2MID[6]
+ Tile_X5Y12_LUT4AB/E2MID[7] Tile_X5Y12_LUT4AB/E2END[0] Tile_X5Y12_LUT4AB/E2END[1]
+ Tile_X5Y12_LUT4AB/E2END[2] Tile_X5Y12_LUT4AB/E2END[3] Tile_X5Y12_LUT4AB/E2END[4]
+ Tile_X5Y12_LUT4AB/E2END[5] Tile_X5Y12_LUT4AB/E2END[6] Tile_X5Y12_LUT4AB/E2END[7]
+ Tile_X4Y12_RegFile/E2END[0] Tile_X4Y12_RegFile/E2END[1] Tile_X4Y12_RegFile/E2END[2]
+ Tile_X4Y12_RegFile/E2END[3] Tile_X4Y12_RegFile/E2END[4] Tile_X4Y12_RegFile/E2END[5]
+ Tile_X4Y12_RegFile/E2END[6] Tile_X4Y12_RegFile/E2END[7] Tile_X3Y12_LUT4AB/E2BEG[0]
+ Tile_X3Y12_LUT4AB/E2BEG[1] Tile_X3Y12_LUT4AB/E2BEG[2] Tile_X3Y12_LUT4AB/E2BEG[3]
+ Tile_X3Y12_LUT4AB/E2BEG[4] Tile_X3Y12_LUT4AB/E2BEG[5] Tile_X3Y12_LUT4AB/E2BEG[6]
+ Tile_X3Y12_LUT4AB/E2BEG[7] Tile_X5Y12_LUT4AB/E6END[0] Tile_X5Y12_LUT4AB/E6END[10]
+ Tile_X5Y12_LUT4AB/E6END[11] Tile_X5Y12_LUT4AB/E6END[1] Tile_X5Y12_LUT4AB/E6END[2]
+ Tile_X5Y12_LUT4AB/E6END[3] Tile_X5Y12_LUT4AB/E6END[4] Tile_X5Y12_LUT4AB/E6END[5]
+ Tile_X5Y12_LUT4AB/E6END[6] Tile_X5Y12_LUT4AB/E6END[7] Tile_X5Y12_LUT4AB/E6END[8]
+ Tile_X5Y12_LUT4AB/E6END[9] Tile_X3Y12_LUT4AB/E6BEG[0] Tile_X3Y12_LUT4AB/E6BEG[10]
+ Tile_X3Y12_LUT4AB/E6BEG[11] Tile_X3Y12_LUT4AB/E6BEG[1] Tile_X3Y12_LUT4AB/E6BEG[2]
+ Tile_X3Y12_LUT4AB/E6BEG[3] Tile_X3Y12_LUT4AB/E6BEG[4] Tile_X3Y12_LUT4AB/E6BEG[5]
+ Tile_X3Y12_LUT4AB/E6BEG[6] Tile_X3Y12_LUT4AB/E6BEG[7] Tile_X3Y12_LUT4AB/E6BEG[8]
+ Tile_X3Y12_LUT4AB/E6BEG[9] Tile_X5Y12_LUT4AB/EE4END[0] Tile_X5Y12_LUT4AB/EE4END[10]
+ Tile_X5Y12_LUT4AB/EE4END[11] Tile_X5Y12_LUT4AB/EE4END[12] Tile_X5Y12_LUT4AB/EE4END[13]
+ Tile_X5Y12_LUT4AB/EE4END[14] Tile_X5Y12_LUT4AB/EE4END[15] Tile_X5Y12_LUT4AB/EE4END[1]
+ Tile_X5Y12_LUT4AB/EE4END[2] Tile_X5Y12_LUT4AB/EE4END[3] Tile_X5Y12_LUT4AB/EE4END[4]
+ Tile_X5Y12_LUT4AB/EE4END[5] Tile_X5Y12_LUT4AB/EE4END[6] Tile_X5Y12_LUT4AB/EE4END[7]
+ Tile_X5Y12_LUT4AB/EE4END[8] Tile_X5Y12_LUT4AB/EE4END[9] Tile_X3Y12_LUT4AB/EE4BEG[0]
+ Tile_X3Y12_LUT4AB/EE4BEG[10] Tile_X3Y12_LUT4AB/EE4BEG[11] Tile_X3Y12_LUT4AB/EE4BEG[12]
+ Tile_X3Y12_LUT4AB/EE4BEG[13] Tile_X3Y12_LUT4AB/EE4BEG[14] Tile_X3Y12_LUT4AB/EE4BEG[15]
+ Tile_X3Y12_LUT4AB/EE4BEG[1] Tile_X3Y12_LUT4AB/EE4BEG[2] Tile_X3Y12_LUT4AB/EE4BEG[3]
+ Tile_X3Y12_LUT4AB/EE4BEG[4] Tile_X3Y12_LUT4AB/EE4BEG[5] Tile_X3Y12_LUT4AB/EE4BEG[6]
+ Tile_X3Y12_LUT4AB/EE4BEG[7] Tile_X3Y12_LUT4AB/EE4BEG[8] Tile_X3Y12_LUT4AB/EE4BEG[9]
+ Tile_X4Y12_RegFile/FrameData[0] Tile_X4Y12_RegFile/FrameData[10] Tile_X4Y12_RegFile/FrameData[11]
+ Tile_X4Y12_RegFile/FrameData[12] Tile_X4Y12_RegFile/FrameData[13] Tile_X4Y12_RegFile/FrameData[14]
+ Tile_X4Y12_RegFile/FrameData[15] Tile_X4Y12_RegFile/FrameData[16] Tile_X4Y12_RegFile/FrameData[17]
+ Tile_X4Y12_RegFile/FrameData[18] Tile_X4Y12_RegFile/FrameData[19] Tile_X4Y12_RegFile/FrameData[1]
+ Tile_X4Y12_RegFile/FrameData[20] Tile_X4Y12_RegFile/FrameData[21] Tile_X4Y12_RegFile/FrameData[22]
+ Tile_X4Y12_RegFile/FrameData[23] Tile_X4Y12_RegFile/FrameData[24] Tile_X4Y12_RegFile/FrameData[25]
+ Tile_X4Y12_RegFile/FrameData[26] Tile_X4Y12_RegFile/FrameData[27] Tile_X4Y12_RegFile/FrameData[28]
+ Tile_X4Y12_RegFile/FrameData[29] Tile_X4Y12_RegFile/FrameData[2] Tile_X4Y12_RegFile/FrameData[30]
+ Tile_X4Y12_RegFile/FrameData[31] Tile_X4Y12_RegFile/FrameData[3] Tile_X4Y12_RegFile/FrameData[4]
+ Tile_X4Y12_RegFile/FrameData[5] Tile_X4Y12_RegFile/FrameData[6] Tile_X4Y12_RegFile/FrameData[7]
+ Tile_X4Y12_RegFile/FrameData[8] Tile_X4Y12_RegFile/FrameData[9] Tile_X5Y12_LUT4AB/FrameData[0]
+ Tile_X5Y12_LUT4AB/FrameData[10] Tile_X5Y12_LUT4AB/FrameData[11] Tile_X5Y12_LUT4AB/FrameData[12]
+ Tile_X5Y12_LUT4AB/FrameData[13] Tile_X5Y12_LUT4AB/FrameData[14] Tile_X5Y12_LUT4AB/FrameData[15]
+ Tile_X5Y12_LUT4AB/FrameData[16] Tile_X5Y12_LUT4AB/FrameData[17] Tile_X5Y12_LUT4AB/FrameData[18]
+ Tile_X5Y12_LUT4AB/FrameData[19] Tile_X5Y12_LUT4AB/FrameData[1] Tile_X5Y12_LUT4AB/FrameData[20]
+ Tile_X5Y12_LUT4AB/FrameData[21] Tile_X5Y12_LUT4AB/FrameData[22] Tile_X5Y12_LUT4AB/FrameData[23]
+ Tile_X5Y12_LUT4AB/FrameData[24] Tile_X5Y12_LUT4AB/FrameData[25] Tile_X5Y12_LUT4AB/FrameData[26]
+ Tile_X5Y12_LUT4AB/FrameData[27] Tile_X5Y12_LUT4AB/FrameData[28] Tile_X5Y12_LUT4AB/FrameData[29]
+ Tile_X5Y12_LUT4AB/FrameData[2] Tile_X5Y12_LUT4AB/FrameData[30] Tile_X5Y12_LUT4AB/FrameData[31]
+ Tile_X5Y12_LUT4AB/FrameData[3] Tile_X5Y12_LUT4AB/FrameData[4] Tile_X5Y12_LUT4AB/FrameData[5]
+ Tile_X5Y12_LUT4AB/FrameData[6] Tile_X5Y12_LUT4AB/FrameData[7] Tile_X5Y12_LUT4AB/FrameData[8]
+ Tile_X5Y12_LUT4AB/FrameData[9] Tile_X4Y12_RegFile/FrameStrobe[0] Tile_X4Y12_RegFile/FrameStrobe[10]
+ Tile_X4Y12_RegFile/FrameStrobe[11] Tile_X4Y12_RegFile/FrameStrobe[12] Tile_X4Y12_RegFile/FrameStrobe[13]
+ Tile_X4Y12_RegFile/FrameStrobe[14] Tile_X4Y12_RegFile/FrameStrobe[15] Tile_X4Y12_RegFile/FrameStrobe[16]
+ Tile_X4Y12_RegFile/FrameStrobe[17] Tile_X4Y12_RegFile/FrameStrobe[18] Tile_X4Y12_RegFile/FrameStrobe[19]
+ Tile_X4Y12_RegFile/FrameStrobe[1] Tile_X4Y12_RegFile/FrameStrobe[2] Tile_X4Y12_RegFile/FrameStrobe[3]
+ Tile_X4Y12_RegFile/FrameStrobe[4] Tile_X4Y12_RegFile/FrameStrobe[5] Tile_X4Y12_RegFile/FrameStrobe[6]
+ Tile_X4Y12_RegFile/FrameStrobe[7] Tile_X4Y12_RegFile/FrameStrobe[8] Tile_X4Y12_RegFile/FrameStrobe[9]
+ Tile_X4Y11_RegFile/FrameStrobe[0] Tile_X4Y11_RegFile/FrameStrobe[10] Tile_X4Y11_RegFile/FrameStrobe[11]
+ Tile_X4Y11_RegFile/FrameStrobe[12] Tile_X4Y11_RegFile/FrameStrobe[13] Tile_X4Y11_RegFile/FrameStrobe[14]
+ Tile_X4Y11_RegFile/FrameStrobe[15] Tile_X4Y11_RegFile/FrameStrobe[16] Tile_X4Y11_RegFile/FrameStrobe[17]
+ Tile_X4Y11_RegFile/FrameStrobe[18] Tile_X4Y11_RegFile/FrameStrobe[19] Tile_X4Y11_RegFile/FrameStrobe[1]
+ Tile_X4Y11_RegFile/FrameStrobe[2] Tile_X4Y11_RegFile/FrameStrobe[3] Tile_X4Y11_RegFile/FrameStrobe[4]
+ Tile_X4Y11_RegFile/FrameStrobe[5] Tile_X4Y11_RegFile/FrameStrobe[6] Tile_X4Y11_RegFile/FrameStrobe[7]
+ Tile_X4Y11_RegFile/FrameStrobe[8] Tile_X4Y11_RegFile/FrameStrobe[9] Tile_X4Y12_RegFile/N1BEG[0]
+ Tile_X4Y12_RegFile/N1BEG[1] Tile_X4Y12_RegFile/N1BEG[2] Tile_X4Y12_RegFile/N1BEG[3]
+ Tile_X4Y13_RegFile/N1BEG[0] Tile_X4Y13_RegFile/N1BEG[1] Tile_X4Y13_RegFile/N1BEG[2]
+ Tile_X4Y13_RegFile/N1BEG[3] Tile_X4Y12_RegFile/N2BEG[0] Tile_X4Y12_RegFile/N2BEG[1]
+ Tile_X4Y12_RegFile/N2BEG[2] Tile_X4Y12_RegFile/N2BEG[3] Tile_X4Y12_RegFile/N2BEG[4]
+ Tile_X4Y12_RegFile/N2BEG[5] Tile_X4Y12_RegFile/N2BEG[6] Tile_X4Y12_RegFile/N2BEG[7]
+ Tile_X4Y11_RegFile/N2END[0] Tile_X4Y11_RegFile/N2END[1] Tile_X4Y11_RegFile/N2END[2]
+ Tile_X4Y11_RegFile/N2END[3] Tile_X4Y11_RegFile/N2END[4] Tile_X4Y11_RegFile/N2END[5]
+ Tile_X4Y11_RegFile/N2END[6] Tile_X4Y11_RegFile/N2END[7] Tile_X4Y12_RegFile/N2END[0]
+ Tile_X4Y12_RegFile/N2END[1] Tile_X4Y12_RegFile/N2END[2] Tile_X4Y12_RegFile/N2END[3]
+ Tile_X4Y12_RegFile/N2END[4] Tile_X4Y12_RegFile/N2END[5] Tile_X4Y12_RegFile/N2END[6]
+ Tile_X4Y12_RegFile/N2END[7] Tile_X4Y13_RegFile/N2BEG[0] Tile_X4Y13_RegFile/N2BEG[1]
+ Tile_X4Y13_RegFile/N2BEG[2] Tile_X4Y13_RegFile/N2BEG[3] Tile_X4Y13_RegFile/N2BEG[4]
+ Tile_X4Y13_RegFile/N2BEG[5] Tile_X4Y13_RegFile/N2BEG[6] Tile_X4Y13_RegFile/N2BEG[7]
+ Tile_X4Y12_RegFile/N4BEG[0] Tile_X4Y12_RegFile/N4BEG[10] Tile_X4Y12_RegFile/N4BEG[11]
+ Tile_X4Y12_RegFile/N4BEG[12] Tile_X4Y12_RegFile/N4BEG[13] Tile_X4Y12_RegFile/N4BEG[14]
+ Tile_X4Y12_RegFile/N4BEG[15] Tile_X4Y12_RegFile/N4BEG[1] Tile_X4Y12_RegFile/N4BEG[2]
+ Tile_X4Y12_RegFile/N4BEG[3] Tile_X4Y12_RegFile/N4BEG[4] Tile_X4Y12_RegFile/N4BEG[5]
+ Tile_X4Y12_RegFile/N4BEG[6] Tile_X4Y12_RegFile/N4BEG[7] Tile_X4Y12_RegFile/N4BEG[8]
+ Tile_X4Y12_RegFile/N4BEG[9] Tile_X4Y13_RegFile/N4BEG[0] Tile_X4Y13_RegFile/N4BEG[10]
+ Tile_X4Y13_RegFile/N4BEG[11] Tile_X4Y13_RegFile/N4BEG[12] Tile_X4Y13_RegFile/N4BEG[13]
+ Tile_X4Y13_RegFile/N4BEG[14] Tile_X4Y13_RegFile/N4BEG[15] Tile_X4Y13_RegFile/N4BEG[1]
+ Tile_X4Y13_RegFile/N4BEG[2] Tile_X4Y13_RegFile/N4BEG[3] Tile_X4Y13_RegFile/N4BEG[4]
+ Tile_X4Y13_RegFile/N4BEG[5] Tile_X4Y13_RegFile/N4BEG[6] Tile_X4Y13_RegFile/N4BEG[7]
+ Tile_X4Y13_RegFile/N4BEG[8] Tile_X4Y13_RegFile/N4BEG[9] Tile_X4Y12_RegFile/NN4BEG[0]
+ Tile_X4Y12_RegFile/NN4BEG[10] Tile_X4Y12_RegFile/NN4BEG[11] Tile_X4Y12_RegFile/NN4BEG[12]
+ Tile_X4Y12_RegFile/NN4BEG[13] Tile_X4Y12_RegFile/NN4BEG[14] Tile_X4Y12_RegFile/NN4BEG[15]
+ Tile_X4Y12_RegFile/NN4BEG[1] Tile_X4Y12_RegFile/NN4BEG[2] Tile_X4Y12_RegFile/NN4BEG[3]
+ Tile_X4Y12_RegFile/NN4BEG[4] Tile_X4Y12_RegFile/NN4BEG[5] Tile_X4Y12_RegFile/NN4BEG[6]
+ Tile_X4Y12_RegFile/NN4BEG[7] Tile_X4Y12_RegFile/NN4BEG[8] Tile_X4Y12_RegFile/NN4BEG[9]
+ Tile_X4Y13_RegFile/NN4BEG[0] Tile_X4Y13_RegFile/NN4BEG[10] Tile_X4Y13_RegFile/NN4BEG[11]
+ Tile_X4Y13_RegFile/NN4BEG[12] Tile_X4Y13_RegFile/NN4BEG[13] Tile_X4Y13_RegFile/NN4BEG[14]
+ Tile_X4Y13_RegFile/NN4BEG[15] Tile_X4Y13_RegFile/NN4BEG[1] Tile_X4Y13_RegFile/NN4BEG[2]
+ Tile_X4Y13_RegFile/NN4BEG[3] Tile_X4Y13_RegFile/NN4BEG[4] Tile_X4Y13_RegFile/NN4BEG[5]
+ Tile_X4Y13_RegFile/NN4BEG[6] Tile_X4Y13_RegFile/NN4BEG[7] Tile_X4Y13_RegFile/NN4BEG[8]
+ Tile_X4Y13_RegFile/NN4BEG[9] Tile_X4Y13_RegFile/S1END[0] Tile_X4Y13_RegFile/S1END[1]
+ Tile_X4Y13_RegFile/S1END[2] Tile_X4Y13_RegFile/S1END[3] Tile_X4Y12_RegFile/S1END[0]
+ Tile_X4Y12_RegFile/S1END[1] Tile_X4Y12_RegFile/S1END[2] Tile_X4Y12_RegFile/S1END[3]
+ Tile_X4Y13_RegFile/S2MID[0] Tile_X4Y13_RegFile/S2MID[1] Tile_X4Y13_RegFile/S2MID[2]
+ Tile_X4Y13_RegFile/S2MID[3] Tile_X4Y13_RegFile/S2MID[4] Tile_X4Y13_RegFile/S2MID[5]
+ Tile_X4Y13_RegFile/S2MID[6] Tile_X4Y13_RegFile/S2MID[7] Tile_X4Y13_RegFile/S2END[0]
+ Tile_X4Y13_RegFile/S2END[1] Tile_X4Y13_RegFile/S2END[2] Tile_X4Y13_RegFile/S2END[3]
+ Tile_X4Y13_RegFile/S2END[4] Tile_X4Y13_RegFile/S2END[5] Tile_X4Y13_RegFile/S2END[6]
+ Tile_X4Y13_RegFile/S2END[7] Tile_X4Y12_RegFile/S2END[0] Tile_X4Y12_RegFile/S2END[1]
+ Tile_X4Y12_RegFile/S2END[2] Tile_X4Y12_RegFile/S2END[3] Tile_X4Y12_RegFile/S2END[4]
+ Tile_X4Y12_RegFile/S2END[5] Tile_X4Y12_RegFile/S2END[6] Tile_X4Y12_RegFile/S2END[7]
+ Tile_X4Y12_RegFile/S2MID[0] Tile_X4Y12_RegFile/S2MID[1] Tile_X4Y12_RegFile/S2MID[2]
+ Tile_X4Y12_RegFile/S2MID[3] Tile_X4Y12_RegFile/S2MID[4] Tile_X4Y12_RegFile/S2MID[5]
+ Tile_X4Y12_RegFile/S2MID[6] Tile_X4Y12_RegFile/S2MID[7] Tile_X4Y13_RegFile/S4END[0]
+ Tile_X4Y13_RegFile/S4END[10] Tile_X4Y13_RegFile/S4END[11] Tile_X4Y13_RegFile/S4END[12]
+ Tile_X4Y13_RegFile/S4END[13] Tile_X4Y13_RegFile/S4END[14] Tile_X4Y13_RegFile/S4END[15]
+ Tile_X4Y13_RegFile/S4END[1] Tile_X4Y13_RegFile/S4END[2] Tile_X4Y13_RegFile/S4END[3]
+ Tile_X4Y13_RegFile/S4END[4] Tile_X4Y13_RegFile/S4END[5] Tile_X4Y13_RegFile/S4END[6]
+ Tile_X4Y13_RegFile/S4END[7] Tile_X4Y13_RegFile/S4END[8] Tile_X4Y13_RegFile/S4END[9]
+ Tile_X4Y12_RegFile/S4END[0] Tile_X4Y12_RegFile/S4END[10] Tile_X4Y12_RegFile/S4END[11]
+ Tile_X4Y12_RegFile/S4END[12] Tile_X4Y12_RegFile/S4END[13] Tile_X4Y12_RegFile/S4END[14]
+ Tile_X4Y12_RegFile/S4END[15] Tile_X4Y12_RegFile/S4END[1] Tile_X4Y12_RegFile/S4END[2]
+ Tile_X4Y12_RegFile/S4END[3] Tile_X4Y12_RegFile/S4END[4] Tile_X4Y12_RegFile/S4END[5]
+ Tile_X4Y12_RegFile/S4END[6] Tile_X4Y12_RegFile/S4END[7] Tile_X4Y12_RegFile/S4END[8]
+ Tile_X4Y12_RegFile/S4END[9] Tile_X4Y13_RegFile/SS4END[0] Tile_X4Y13_RegFile/SS4END[10]
+ Tile_X4Y13_RegFile/SS4END[11] Tile_X4Y13_RegFile/SS4END[12] Tile_X4Y13_RegFile/SS4END[13]
+ Tile_X4Y13_RegFile/SS4END[14] Tile_X4Y13_RegFile/SS4END[15] Tile_X4Y13_RegFile/SS4END[1]
+ Tile_X4Y13_RegFile/SS4END[2] Tile_X4Y13_RegFile/SS4END[3] Tile_X4Y13_RegFile/SS4END[4]
+ Tile_X4Y13_RegFile/SS4END[5] Tile_X4Y13_RegFile/SS4END[6] Tile_X4Y13_RegFile/SS4END[7]
+ Tile_X4Y13_RegFile/SS4END[8] Tile_X4Y13_RegFile/SS4END[9] Tile_X4Y12_RegFile/SS4END[0]
+ Tile_X4Y12_RegFile/SS4END[10] Tile_X4Y12_RegFile/SS4END[11] Tile_X4Y12_RegFile/SS4END[12]
+ Tile_X4Y12_RegFile/SS4END[13] Tile_X4Y12_RegFile/SS4END[14] Tile_X4Y12_RegFile/SS4END[15]
+ Tile_X4Y12_RegFile/SS4END[1] Tile_X4Y12_RegFile/SS4END[2] Tile_X4Y12_RegFile/SS4END[3]
+ Tile_X4Y12_RegFile/SS4END[4] Tile_X4Y12_RegFile/SS4END[5] Tile_X4Y12_RegFile/SS4END[6]
+ Tile_X4Y12_RegFile/SS4END[7] Tile_X4Y12_RegFile/SS4END[8] Tile_X4Y12_RegFile/SS4END[9]
+ Tile_X4Y12_RegFile/UserCLK Tile_X4Y11_RegFile/UserCLK VGND VPWR Tile_X3Y12_LUT4AB/W1END[0]
+ Tile_X3Y12_LUT4AB/W1END[1] Tile_X3Y12_LUT4AB/W1END[2] Tile_X3Y12_LUT4AB/W1END[3]
+ Tile_X5Y12_LUT4AB/W1BEG[0] Tile_X5Y12_LUT4AB/W1BEG[1] Tile_X5Y12_LUT4AB/W1BEG[2]
+ Tile_X5Y12_LUT4AB/W1BEG[3] Tile_X3Y12_LUT4AB/W2MID[0] Tile_X3Y12_LUT4AB/W2MID[1]
+ Tile_X3Y12_LUT4AB/W2MID[2] Tile_X3Y12_LUT4AB/W2MID[3] Tile_X3Y12_LUT4AB/W2MID[4]
+ Tile_X3Y12_LUT4AB/W2MID[5] Tile_X3Y12_LUT4AB/W2MID[6] Tile_X3Y12_LUT4AB/W2MID[7]
+ Tile_X3Y12_LUT4AB/W2END[0] Tile_X3Y12_LUT4AB/W2END[1] Tile_X3Y12_LUT4AB/W2END[2]
+ Tile_X3Y12_LUT4AB/W2END[3] Tile_X3Y12_LUT4AB/W2END[4] Tile_X3Y12_LUT4AB/W2END[5]
+ Tile_X3Y12_LUT4AB/W2END[6] Tile_X3Y12_LUT4AB/W2END[7] Tile_X5Y12_LUT4AB/W2BEGb[0]
+ Tile_X5Y12_LUT4AB/W2BEGb[1] Tile_X5Y12_LUT4AB/W2BEGb[2] Tile_X5Y12_LUT4AB/W2BEGb[3]
+ Tile_X5Y12_LUT4AB/W2BEGb[4] Tile_X5Y12_LUT4AB/W2BEGb[5] Tile_X5Y12_LUT4AB/W2BEGb[6]
+ Tile_X5Y12_LUT4AB/W2BEGb[7] Tile_X5Y12_LUT4AB/W2BEG[0] Tile_X5Y12_LUT4AB/W2BEG[1]
+ Tile_X5Y12_LUT4AB/W2BEG[2] Tile_X5Y12_LUT4AB/W2BEG[3] Tile_X5Y12_LUT4AB/W2BEG[4]
+ Tile_X5Y12_LUT4AB/W2BEG[5] Tile_X5Y12_LUT4AB/W2BEG[6] Tile_X5Y12_LUT4AB/W2BEG[7]
+ Tile_X3Y12_LUT4AB/W6END[0] Tile_X3Y12_LUT4AB/W6END[10] Tile_X3Y12_LUT4AB/W6END[11]
+ Tile_X3Y12_LUT4AB/W6END[1] Tile_X3Y12_LUT4AB/W6END[2] Tile_X3Y12_LUT4AB/W6END[3]
+ Tile_X3Y12_LUT4AB/W6END[4] Tile_X3Y12_LUT4AB/W6END[5] Tile_X3Y12_LUT4AB/W6END[6]
+ Tile_X3Y12_LUT4AB/W6END[7] Tile_X3Y12_LUT4AB/W6END[8] Tile_X3Y12_LUT4AB/W6END[9]
+ Tile_X5Y12_LUT4AB/W6BEG[0] Tile_X5Y12_LUT4AB/W6BEG[10] Tile_X5Y12_LUT4AB/W6BEG[11]
+ Tile_X5Y12_LUT4AB/W6BEG[1] Tile_X5Y12_LUT4AB/W6BEG[2] Tile_X5Y12_LUT4AB/W6BEG[3]
+ Tile_X5Y12_LUT4AB/W6BEG[4] Tile_X5Y12_LUT4AB/W6BEG[5] Tile_X5Y12_LUT4AB/W6BEG[6]
+ Tile_X5Y12_LUT4AB/W6BEG[7] Tile_X5Y12_LUT4AB/W6BEG[8] Tile_X5Y12_LUT4AB/W6BEG[9]
+ Tile_X3Y12_LUT4AB/WW4END[0] Tile_X3Y12_LUT4AB/WW4END[10] Tile_X3Y12_LUT4AB/WW4END[11]
+ Tile_X3Y12_LUT4AB/WW4END[12] Tile_X3Y12_LUT4AB/WW4END[13] Tile_X3Y12_LUT4AB/WW4END[14]
+ Tile_X3Y12_LUT4AB/WW4END[15] Tile_X3Y12_LUT4AB/WW4END[1] Tile_X3Y12_LUT4AB/WW4END[2]
+ Tile_X3Y12_LUT4AB/WW4END[3] Tile_X3Y12_LUT4AB/WW4END[4] Tile_X3Y12_LUT4AB/WW4END[5]
+ Tile_X3Y12_LUT4AB/WW4END[6] Tile_X3Y12_LUT4AB/WW4END[7] Tile_X3Y12_LUT4AB/WW4END[8]
+ Tile_X3Y12_LUT4AB/WW4END[9] Tile_X5Y12_LUT4AB/WW4BEG[0] Tile_X5Y12_LUT4AB/WW4BEG[10]
+ Tile_X5Y12_LUT4AB/WW4BEG[11] Tile_X5Y12_LUT4AB/WW4BEG[12] Tile_X5Y12_LUT4AB/WW4BEG[13]
+ Tile_X5Y12_LUT4AB/WW4BEG[14] Tile_X5Y12_LUT4AB/WW4BEG[15] Tile_X5Y12_LUT4AB/WW4BEG[1]
+ Tile_X5Y12_LUT4AB/WW4BEG[2] Tile_X5Y12_LUT4AB/WW4BEG[3] Tile_X5Y12_LUT4AB/WW4BEG[4]
+ Tile_X5Y12_LUT4AB/WW4BEG[5] Tile_X5Y12_LUT4AB/WW4BEG[6] Tile_X5Y12_LUT4AB/WW4BEG[7]
+ Tile_X5Y12_LUT4AB/WW4BEG[8] Tile_X5Y12_LUT4AB/WW4BEG[9] RegFile
XTile_X7Y15_S_term_DSP Tile_X7Y15_S_term_DSP/FrameData[0] Tile_X7Y15_S_term_DSP/FrameData[10]
+ Tile_X7Y15_S_term_DSP/FrameData[11] Tile_X7Y15_S_term_DSP/FrameData[12] Tile_X7Y15_S_term_DSP/FrameData[13]
+ Tile_X7Y15_S_term_DSP/FrameData[14] Tile_X7Y15_S_term_DSP/FrameData[15] Tile_X7Y15_S_term_DSP/FrameData[16]
+ Tile_X7Y15_S_term_DSP/FrameData[17] Tile_X7Y15_S_term_DSP/FrameData[18] Tile_X7Y15_S_term_DSP/FrameData[19]
+ Tile_X7Y15_S_term_DSP/FrameData[1] Tile_X7Y15_S_term_DSP/FrameData[20] Tile_X7Y15_S_term_DSP/FrameData[21]
+ Tile_X7Y15_S_term_DSP/FrameData[22] Tile_X7Y15_S_term_DSP/FrameData[23] Tile_X7Y15_S_term_DSP/FrameData[24]
+ Tile_X7Y15_S_term_DSP/FrameData[25] Tile_X7Y15_S_term_DSP/FrameData[26] Tile_X7Y15_S_term_DSP/FrameData[27]
+ Tile_X7Y15_S_term_DSP/FrameData[28] Tile_X7Y15_S_term_DSP/FrameData[29] Tile_X7Y15_S_term_DSP/FrameData[2]
+ Tile_X7Y15_S_term_DSP/FrameData[30] Tile_X7Y15_S_term_DSP/FrameData[31] Tile_X7Y15_S_term_DSP/FrameData[3]
+ Tile_X7Y15_S_term_DSP/FrameData[4] Tile_X7Y15_S_term_DSP/FrameData[5] Tile_X7Y15_S_term_DSP/FrameData[6]
+ Tile_X7Y15_S_term_DSP/FrameData[7] Tile_X7Y15_S_term_DSP/FrameData[8] Tile_X7Y15_S_term_DSP/FrameData[9]
+ Tile_X8Y15_S_CPU_IF/FrameData[0] Tile_X8Y15_S_CPU_IF/FrameData[10] Tile_X8Y15_S_CPU_IF/FrameData[11]
+ Tile_X8Y15_S_CPU_IF/FrameData[12] Tile_X8Y15_S_CPU_IF/FrameData[13] Tile_X8Y15_S_CPU_IF/FrameData[14]
+ Tile_X8Y15_S_CPU_IF/FrameData[15] Tile_X8Y15_S_CPU_IF/FrameData[16] Tile_X8Y15_S_CPU_IF/FrameData[17]
+ Tile_X8Y15_S_CPU_IF/FrameData[18] Tile_X8Y15_S_CPU_IF/FrameData[19] Tile_X8Y15_S_CPU_IF/FrameData[1]
+ Tile_X8Y15_S_CPU_IF/FrameData[20] Tile_X8Y15_S_CPU_IF/FrameData[21] Tile_X8Y15_S_CPU_IF/FrameData[22]
+ Tile_X8Y15_S_CPU_IF/FrameData[23] Tile_X8Y15_S_CPU_IF/FrameData[24] Tile_X8Y15_S_CPU_IF/FrameData[25]
+ Tile_X8Y15_S_CPU_IF/FrameData[26] Tile_X8Y15_S_CPU_IF/FrameData[27] Tile_X8Y15_S_CPU_IF/FrameData[28]
+ Tile_X8Y15_S_CPU_IF/FrameData[29] Tile_X8Y15_S_CPU_IF/FrameData[2] Tile_X8Y15_S_CPU_IF/FrameData[30]
+ Tile_X8Y15_S_CPU_IF/FrameData[31] Tile_X8Y15_S_CPU_IF/FrameData[3] Tile_X8Y15_S_CPU_IF/FrameData[4]
+ Tile_X8Y15_S_CPU_IF/FrameData[5] Tile_X8Y15_S_CPU_IF/FrameData[6] Tile_X8Y15_S_CPU_IF/FrameData[7]
+ Tile_X8Y15_S_CPU_IF/FrameData[8] Tile_X8Y15_S_CPU_IF/FrameData[9] FrameStrobe[140]
+ FrameStrobe[150] FrameStrobe[151] FrameStrobe[152] FrameStrobe[153] FrameStrobe[154]
+ FrameStrobe[155] FrameStrobe[156] FrameStrobe[157] FrameStrobe[158] FrameStrobe[159]
+ FrameStrobe[141] FrameStrobe[142] FrameStrobe[143] FrameStrobe[144] FrameStrobe[145]
+ FrameStrobe[146] FrameStrobe[147] FrameStrobe[148] FrameStrobe[149] Tile_X7Y15_S_term_DSP/FrameStrobe_O[0]
+ Tile_X7Y15_S_term_DSP/FrameStrobe_O[10] Tile_X7Y15_S_term_DSP/FrameStrobe_O[11]
+ Tile_X7Y15_S_term_DSP/FrameStrobe_O[12] Tile_X7Y15_S_term_DSP/FrameStrobe_O[13]
+ Tile_X7Y15_S_term_DSP/FrameStrobe_O[14] Tile_X7Y15_S_term_DSP/FrameStrobe_O[15]
+ Tile_X7Y15_S_term_DSP/FrameStrobe_O[16] Tile_X7Y15_S_term_DSP/FrameStrobe_O[17]
+ Tile_X7Y15_S_term_DSP/FrameStrobe_O[18] Tile_X7Y15_S_term_DSP/FrameStrobe_O[19]
+ Tile_X7Y15_S_term_DSP/FrameStrobe_O[1] Tile_X7Y15_S_term_DSP/FrameStrobe_O[2] Tile_X7Y15_S_term_DSP/FrameStrobe_O[3]
+ Tile_X7Y15_S_term_DSP/FrameStrobe_O[4] Tile_X7Y15_S_term_DSP/FrameStrobe_O[5] Tile_X7Y15_S_term_DSP/FrameStrobe_O[6]
+ Tile_X7Y15_S_term_DSP/FrameStrobe_O[7] Tile_X7Y15_S_term_DSP/FrameStrobe_O[8] Tile_X7Y15_S_term_DSP/FrameStrobe_O[9]
+ Tile_X7Y15_S_term_DSP/N1BEG[0] Tile_X7Y15_S_term_DSP/N1BEG[1] Tile_X7Y15_S_term_DSP/N1BEG[2]
+ Tile_X7Y15_S_term_DSP/N1BEG[3] Tile_X7Y15_S_term_DSP/N2BEG[0] Tile_X7Y15_S_term_DSP/N2BEG[1]
+ Tile_X7Y15_S_term_DSP/N2BEG[2] Tile_X7Y15_S_term_DSP/N2BEG[3] Tile_X7Y15_S_term_DSP/N2BEG[4]
+ Tile_X7Y15_S_term_DSP/N2BEG[5] Tile_X7Y15_S_term_DSP/N2BEG[6] Tile_X7Y15_S_term_DSP/N2BEG[7]
+ Tile_X7Y15_S_term_DSP/N2BEGb[0] Tile_X7Y15_S_term_DSP/N2BEGb[1] Tile_X7Y15_S_term_DSP/N2BEGb[2]
+ Tile_X7Y15_S_term_DSP/N2BEGb[3] Tile_X7Y15_S_term_DSP/N2BEGb[4] Tile_X7Y15_S_term_DSP/N2BEGb[5]
+ Tile_X7Y15_S_term_DSP/N2BEGb[6] Tile_X7Y15_S_term_DSP/N2BEGb[7] Tile_X7Y15_S_term_DSP/N4BEG[0]
+ Tile_X7Y15_S_term_DSP/N4BEG[10] Tile_X7Y15_S_term_DSP/N4BEG[11] Tile_X7Y15_S_term_DSP/N4BEG[12]
+ Tile_X7Y15_S_term_DSP/N4BEG[13] Tile_X7Y15_S_term_DSP/N4BEG[14] Tile_X7Y15_S_term_DSP/N4BEG[15]
+ Tile_X7Y15_S_term_DSP/N4BEG[1] Tile_X7Y15_S_term_DSP/N4BEG[2] Tile_X7Y15_S_term_DSP/N4BEG[3]
+ Tile_X7Y15_S_term_DSP/N4BEG[4] Tile_X7Y15_S_term_DSP/N4BEG[5] Tile_X7Y15_S_term_DSP/N4BEG[6]
+ Tile_X7Y15_S_term_DSP/N4BEG[7] Tile_X7Y15_S_term_DSP/N4BEG[8] Tile_X7Y15_S_term_DSP/N4BEG[9]
+ Tile_X7Y15_S_term_DSP/NN4BEG[0] Tile_X7Y15_S_term_DSP/NN4BEG[10] Tile_X7Y15_S_term_DSP/NN4BEG[11]
+ Tile_X7Y15_S_term_DSP/NN4BEG[12] Tile_X7Y15_S_term_DSP/NN4BEG[13] Tile_X7Y15_S_term_DSP/NN4BEG[14]
+ Tile_X7Y15_S_term_DSP/NN4BEG[15] Tile_X7Y15_S_term_DSP/NN4BEG[1] Tile_X7Y15_S_term_DSP/NN4BEG[2]
+ Tile_X7Y15_S_term_DSP/NN4BEG[3] Tile_X7Y15_S_term_DSP/NN4BEG[4] Tile_X7Y15_S_term_DSP/NN4BEG[5]
+ Tile_X7Y15_S_term_DSP/NN4BEG[6] Tile_X7Y15_S_term_DSP/NN4BEG[7] Tile_X7Y15_S_term_DSP/NN4BEG[8]
+ Tile_X7Y15_S_term_DSP/NN4BEG[9] Tile_X7Y15_S_term_DSP/S1END[0] Tile_X7Y15_S_term_DSP/S1END[1]
+ Tile_X7Y15_S_term_DSP/S1END[2] Tile_X7Y15_S_term_DSP/S1END[3] Tile_X7Y15_S_term_DSP/S2END[0]
+ Tile_X7Y15_S_term_DSP/S2END[1] Tile_X7Y15_S_term_DSP/S2END[2] Tile_X7Y15_S_term_DSP/S2END[3]
+ Tile_X7Y15_S_term_DSP/S2END[4] Tile_X7Y15_S_term_DSP/S2END[5] Tile_X7Y15_S_term_DSP/S2END[6]
+ Tile_X7Y15_S_term_DSP/S2END[7] Tile_X7Y15_S_term_DSP/S2MID[0] Tile_X7Y15_S_term_DSP/S2MID[1]
+ Tile_X7Y15_S_term_DSP/S2MID[2] Tile_X7Y15_S_term_DSP/S2MID[3] Tile_X7Y15_S_term_DSP/S2MID[4]
+ Tile_X7Y15_S_term_DSP/S2MID[5] Tile_X7Y15_S_term_DSP/S2MID[6] Tile_X7Y15_S_term_DSP/S2MID[7]
+ Tile_X7Y15_S_term_DSP/S4END[0] Tile_X7Y15_S_term_DSP/S4END[10] Tile_X7Y15_S_term_DSP/S4END[11]
+ Tile_X7Y15_S_term_DSP/S4END[12] Tile_X7Y15_S_term_DSP/S4END[13] Tile_X7Y15_S_term_DSP/S4END[14]
+ Tile_X7Y15_S_term_DSP/S4END[15] Tile_X7Y15_S_term_DSP/S4END[1] Tile_X7Y15_S_term_DSP/S4END[2]
+ Tile_X7Y15_S_term_DSP/S4END[3] Tile_X7Y15_S_term_DSP/S4END[4] Tile_X7Y15_S_term_DSP/S4END[5]
+ Tile_X7Y15_S_term_DSP/S4END[6] Tile_X7Y15_S_term_DSP/S4END[7] Tile_X7Y15_S_term_DSP/S4END[8]
+ Tile_X7Y15_S_term_DSP/S4END[9] Tile_X7Y15_S_term_DSP/SS4END[0] Tile_X7Y15_S_term_DSP/SS4END[10]
+ Tile_X7Y15_S_term_DSP/SS4END[11] Tile_X7Y15_S_term_DSP/SS4END[12] Tile_X7Y15_S_term_DSP/SS4END[13]
+ Tile_X7Y15_S_term_DSP/SS4END[14] Tile_X7Y15_S_term_DSP/SS4END[15] Tile_X7Y15_S_term_DSP/SS4END[1]
+ Tile_X7Y15_S_term_DSP/SS4END[2] Tile_X7Y15_S_term_DSP/SS4END[3] Tile_X7Y15_S_term_DSP/SS4END[4]
+ Tile_X7Y15_S_term_DSP/SS4END[5] Tile_X7Y15_S_term_DSP/SS4END[6] Tile_X7Y15_S_term_DSP/SS4END[7]
+ Tile_X7Y15_S_term_DSP/SS4END[8] Tile_X7Y15_S_term_DSP/SS4END[9] UserCLK Tile_X7Y15_S_term_DSP/UserCLKo
+ VGND VPWR S_term_DSP
XTile_X3Y9_LUT4AB Tile_X3Y9_LUT4AB/Ci Tile_X3Y9_LUT4AB/Co Tile_X3Y9_LUT4AB/E1BEG[0]
+ Tile_X3Y9_LUT4AB/E1BEG[1] Tile_X3Y9_LUT4AB/E1BEG[2] Tile_X3Y9_LUT4AB/E1BEG[3] Tile_X3Y9_LUT4AB/E1END[0]
+ Tile_X3Y9_LUT4AB/E1END[1] Tile_X3Y9_LUT4AB/E1END[2] Tile_X3Y9_LUT4AB/E1END[3] Tile_X3Y9_LUT4AB/E2BEG[0]
+ Tile_X3Y9_LUT4AB/E2BEG[1] Tile_X3Y9_LUT4AB/E2BEG[2] Tile_X3Y9_LUT4AB/E2BEG[3] Tile_X3Y9_LUT4AB/E2BEG[4]
+ Tile_X3Y9_LUT4AB/E2BEG[5] Tile_X3Y9_LUT4AB/E2BEG[6] Tile_X3Y9_LUT4AB/E2BEG[7] Tile_X4Y9_RegFile/E2END[0]
+ Tile_X4Y9_RegFile/E2END[1] Tile_X4Y9_RegFile/E2END[2] Tile_X4Y9_RegFile/E2END[3]
+ Tile_X4Y9_RegFile/E2END[4] Tile_X4Y9_RegFile/E2END[5] Tile_X4Y9_RegFile/E2END[6]
+ Tile_X4Y9_RegFile/E2END[7] Tile_X3Y9_LUT4AB/E2END[0] Tile_X3Y9_LUT4AB/E2END[1] Tile_X3Y9_LUT4AB/E2END[2]
+ Tile_X3Y9_LUT4AB/E2END[3] Tile_X3Y9_LUT4AB/E2END[4] Tile_X3Y9_LUT4AB/E2END[5] Tile_X3Y9_LUT4AB/E2END[6]
+ Tile_X3Y9_LUT4AB/E2END[7] Tile_X3Y9_LUT4AB/E2MID[0] Tile_X3Y9_LUT4AB/E2MID[1] Tile_X3Y9_LUT4AB/E2MID[2]
+ Tile_X3Y9_LUT4AB/E2MID[3] Tile_X3Y9_LUT4AB/E2MID[4] Tile_X3Y9_LUT4AB/E2MID[5] Tile_X3Y9_LUT4AB/E2MID[6]
+ Tile_X3Y9_LUT4AB/E2MID[7] Tile_X3Y9_LUT4AB/E6BEG[0] Tile_X3Y9_LUT4AB/E6BEG[10] Tile_X3Y9_LUT4AB/E6BEG[11]
+ Tile_X3Y9_LUT4AB/E6BEG[1] Tile_X3Y9_LUT4AB/E6BEG[2] Tile_X3Y9_LUT4AB/E6BEG[3] Tile_X3Y9_LUT4AB/E6BEG[4]
+ Tile_X3Y9_LUT4AB/E6BEG[5] Tile_X3Y9_LUT4AB/E6BEG[6] Tile_X3Y9_LUT4AB/E6BEG[7] Tile_X3Y9_LUT4AB/E6BEG[8]
+ Tile_X3Y9_LUT4AB/E6BEG[9] Tile_X3Y9_LUT4AB/E6END[0] Tile_X3Y9_LUT4AB/E6END[10] Tile_X3Y9_LUT4AB/E6END[11]
+ Tile_X3Y9_LUT4AB/E6END[1] Tile_X3Y9_LUT4AB/E6END[2] Tile_X3Y9_LUT4AB/E6END[3] Tile_X3Y9_LUT4AB/E6END[4]
+ Tile_X3Y9_LUT4AB/E6END[5] Tile_X3Y9_LUT4AB/E6END[6] Tile_X3Y9_LUT4AB/E6END[7] Tile_X3Y9_LUT4AB/E6END[8]
+ Tile_X3Y9_LUT4AB/E6END[9] Tile_X3Y9_LUT4AB/EE4BEG[0] Tile_X3Y9_LUT4AB/EE4BEG[10]
+ Tile_X3Y9_LUT4AB/EE4BEG[11] Tile_X3Y9_LUT4AB/EE4BEG[12] Tile_X3Y9_LUT4AB/EE4BEG[13]
+ Tile_X3Y9_LUT4AB/EE4BEG[14] Tile_X3Y9_LUT4AB/EE4BEG[15] Tile_X3Y9_LUT4AB/EE4BEG[1]
+ Tile_X3Y9_LUT4AB/EE4BEG[2] Tile_X3Y9_LUT4AB/EE4BEG[3] Tile_X3Y9_LUT4AB/EE4BEG[4]
+ Tile_X3Y9_LUT4AB/EE4BEG[5] Tile_X3Y9_LUT4AB/EE4BEG[6] Tile_X3Y9_LUT4AB/EE4BEG[7]
+ Tile_X3Y9_LUT4AB/EE4BEG[8] Tile_X3Y9_LUT4AB/EE4BEG[9] Tile_X3Y9_LUT4AB/EE4END[0]
+ Tile_X3Y9_LUT4AB/EE4END[10] Tile_X3Y9_LUT4AB/EE4END[11] Tile_X3Y9_LUT4AB/EE4END[12]
+ Tile_X3Y9_LUT4AB/EE4END[13] Tile_X3Y9_LUT4AB/EE4END[14] Tile_X3Y9_LUT4AB/EE4END[15]
+ Tile_X3Y9_LUT4AB/EE4END[1] Tile_X3Y9_LUT4AB/EE4END[2] Tile_X3Y9_LUT4AB/EE4END[3]
+ Tile_X3Y9_LUT4AB/EE4END[4] Tile_X3Y9_LUT4AB/EE4END[5] Tile_X3Y9_LUT4AB/EE4END[6]
+ Tile_X3Y9_LUT4AB/EE4END[7] Tile_X3Y9_LUT4AB/EE4END[8] Tile_X3Y9_LUT4AB/EE4END[9]
+ Tile_X3Y9_LUT4AB/FrameData[0] Tile_X3Y9_LUT4AB/FrameData[10] Tile_X3Y9_LUT4AB/FrameData[11]
+ Tile_X3Y9_LUT4AB/FrameData[12] Tile_X3Y9_LUT4AB/FrameData[13] Tile_X3Y9_LUT4AB/FrameData[14]
+ Tile_X3Y9_LUT4AB/FrameData[15] Tile_X3Y9_LUT4AB/FrameData[16] Tile_X3Y9_LUT4AB/FrameData[17]
+ Tile_X3Y9_LUT4AB/FrameData[18] Tile_X3Y9_LUT4AB/FrameData[19] Tile_X3Y9_LUT4AB/FrameData[1]
+ Tile_X3Y9_LUT4AB/FrameData[20] Tile_X3Y9_LUT4AB/FrameData[21] Tile_X3Y9_LUT4AB/FrameData[22]
+ Tile_X3Y9_LUT4AB/FrameData[23] Tile_X3Y9_LUT4AB/FrameData[24] Tile_X3Y9_LUT4AB/FrameData[25]
+ Tile_X3Y9_LUT4AB/FrameData[26] Tile_X3Y9_LUT4AB/FrameData[27] Tile_X3Y9_LUT4AB/FrameData[28]
+ Tile_X3Y9_LUT4AB/FrameData[29] Tile_X3Y9_LUT4AB/FrameData[2] Tile_X3Y9_LUT4AB/FrameData[30]
+ Tile_X3Y9_LUT4AB/FrameData[31] Tile_X3Y9_LUT4AB/FrameData[3] Tile_X3Y9_LUT4AB/FrameData[4]
+ Tile_X3Y9_LUT4AB/FrameData[5] Tile_X3Y9_LUT4AB/FrameData[6] Tile_X3Y9_LUT4AB/FrameData[7]
+ Tile_X3Y9_LUT4AB/FrameData[8] Tile_X3Y9_LUT4AB/FrameData[9] Tile_X4Y9_RegFile/FrameData[0]
+ Tile_X4Y9_RegFile/FrameData[10] Tile_X4Y9_RegFile/FrameData[11] Tile_X4Y9_RegFile/FrameData[12]
+ Tile_X4Y9_RegFile/FrameData[13] Tile_X4Y9_RegFile/FrameData[14] Tile_X4Y9_RegFile/FrameData[15]
+ Tile_X4Y9_RegFile/FrameData[16] Tile_X4Y9_RegFile/FrameData[17] Tile_X4Y9_RegFile/FrameData[18]
+ Tile_X4Y9_RegFile/FrameData[19] Tile_X4Y9_RegFile/FrameData[1] Tile_X4Y9_RegFile/FrameData[20]
+ Tile_X4Y9_RegFile/FrameData[21] Tile_X4Y9_RegFile/FrameData[22] Tile_X4Y9_RegFile/FrameData[23]
+ Tile_X4Y9_RegFile/FrameData[24] Tile_X4Y9_RegFile/FrameData[25] Tile_X4Y9_RegFile/FrameData[26]
+ Tile_X4Y9_RegFile/FrameData[27] Tile_X4Y9_RegFile/FrameData[28] Tile_X4Y9_RegFile/FrameData[29]
+ Tile_X4Y9_RegFile/FrameData[2] Tile_X4Y9_RegFile/FrameData[30] Tile_X4Y9_RegFile/FrameData[31]
+ Tile_X4Y9_RegFile/FrameData[3] Tile_X4Y9_RegFile/FrameData[4] Tile_X4Y9_RegFile/FrameData[5]
+ Tile_X4Y9_RegFile/FrameData[6] Tile_X4Y9_RegFile/FrameData[7] Tile_X4Y9_RegFile/FrameData[8]
+ Tile_X4Y9_RegFile/FrameData[9] Tile_X3Y9_LUT4AB/FrameStrobe[0] Tile_X3Y9_LUT4AB/FrameStrobe[10]
+ Tile_X3Y9_LUT4AB/FrameStrobe[11] Tile_X3Y9_LUT4AB/FrameStrobe[12] Tile_X3Y9_LUT4AB/FrameStrobe[13]
+ Tile_X3Y9_LUT4AB/FrameStrobe[14] Tile_X3Y9_LUT4AB/FrameStrobe[15] Tile_X3Y9_LUT4AB/FrameStrobe[16]
+ Tile_X3Y9_LUT4AB/FrameStrobe[17] Tile_X3Y9_LUT4AB/FrameStrobe[18] Tile_X3Y9_LUT4AB/FrameStrobe[19]
+ Tile_X3Y9_LUT4AB/FrameStrobe[1] Tile_X3Y9_LUT4AB/FrameStrobe[2] Tile_X3Y9_LUT4AB/FrameStrobe[3]
+ Tile_X3Y9_LUT4AB/FrameStrobe[4] Tile_X3Y9_LUT4AB/FrameStrobe[5] Tile_X3Y9_LUT4AB/FrameStrobe[6]
+ Tile_X3Y9_LUT4AB/FrameStrobe[7] Tile_X3Y9_LUT4AB/FrameStrobe[8] Tile_X3Y9_LUT4AB/FrameStrobe[9]
+ Tile_X3Y8_LUT4AB/FrameStrobe[0] Tile_X3Y8_LUT4AB/FrameStrobe[10] Tile_X3Y8_LUT4AB/FrameStrobe[11]
+ Tile_X3Y8_LUT4AB/FrameStrobe[12] Tile_X3Y8_LUT4AB/FrameStrobe[13] Tile_X3Y8_LUT4AB/FrameStrobe[14]
+ Tile_X3Y8_LUT4AB/FrameStrobe[15] Tile_X3Y8_LUT4AB/FrameStrobe[16] Tile_X3Y8_LUT4AB/FrameStrobe[17]
+ Tile_X3Y8_LUT4AB/FrameStrobe[18] Tile_X3Y8_LUT4AB/FrameStrobe[19] Tile_X3Y8_LUT4AB/FrameStrobe[1]
+ Tile_X3Y8_LUT4AB/FrameStrobe[2] Tile_X3Y8_LUT4AB/FrameStrobe[3] Tile_X3Y8_LUT4AB/FrameStrobe[4]
+ Tile_X3Y8_LUT4AB/FrameStrobe[5] Tile_X3Y8_LUT4AB/FrameStrobe[6] Tile_X3Y8_LUT4AB/FrameStrobe[7]
+ Tile_X3Y8_LUT4AB/FrameStrobe[8] Tile_X3Y8_LUT4AB/FrameStrobe[9] Tile_X3Y9_LUT4AB/N1BEG[0]
+ Tile_X3Y9_LUT4AB/N1BEG[1] Tile_X3Y9_LUT4AB/N1BEG[2] Tile_X3Y9_LUT4AB/N1BEG[3] Tile_X3Y9_LUT4AB/N1END[0]
+ Tile_X3Y9_LUT4AB/N1END[1] Tile_X3Y9_LUT4AB/N1END[2] Tile_X3Y9_LUT4AB/N1END[3] Tile_X3Y9_LUT4AB/N2BEG[0]
+ Tile_X3Y9_LUT4AB/N2BEG[1] Tile_X3Y9_LUT4AB/N2BEG[2] Tile_X3Y9_LUT4AB/N2BEG[3] Tile_X3Y9_LUT4AB/N2BEG[4]
+ Tile_X3Y9_LUT4AB/N2BEG[5] Tile_X3Y9_LUT4AB/N2BEG[6] Tile_X3Y9_LUT4AB/N2BEG[7] Tile_X3Y8_LUT4AB/N2END[0]
+ Tile_X3Y8_LUT4AB/N2END[1] Tile_X3Y8_LUT4AB/N2END[2] Tile_X3Y8_LUT4AB/N2END[3] Tile_X3Y8_LUT4AB/N2END[4]
+ Tile_X3Y8_LUT4AB/N2END[5] Tile_X3Y8_LUT4AB/N2END[6] Tile_X3Y8_LUT4AB/N2END[7] Tile_X3Y9_LUT4AB/N2END[0]
+ Tile_X3Y9_LUT4AB/N2END[1] Tile_X3Y9_LUT4AB/N2END[2] Tile_X3Y9_LUT4AB/N2END[3] Tile_X3Y9_LUT4AB/N2END[4]
+ Tile_X3Y9_LUT4AB/N2END[5] Tile_X3Y9_LUT4AB/N2END[6] Tile_X3Y9_LUT4AB/N2END[7] Tile_X3Y9_LUT4AB/N2MID[0]
+ Tile_X3Y9_LUT4AB/N2MID[1] Tile_X3Y9_LUT4AB/N2MID[2] Tile_X3Y9_LUT4AB/N2MID[3] Tile_X3Y9_LUT4AB/N2MID[4]
+ Tile_X3Y9_LUT4AB/N2MID[5] Tile_X3Y9_LUT4AB/N2MID[6] Tile_X3Y9_LUT4AB/N2MID[7] Tile_X3Y9_LUT4AB/N4BEG[0]
+ Tile_X3Y9_LUT4AB/N4BEG[10] Tile_X3Y9_LUT4AB/N4BEG[11] Tile_X3Y9_LUT4AB/N4BEG[12]
+ Tile_X3Y9_LUT4AB/N4BEG[13] Tile_X3Y9_LUT4AB/N4BEG[14] Tile_X3Y9_LUT4AB/N4BEG[15]
+ Tile_X3Y9_LUT4AB/N4BEG[1] Tile_X3Y9_LUT4AB/N4BEG[2] Tile_X3Y9_LUT4AB/N4BEG[3] Tile_X3Y9_LUT4AB/N4BEG[4]
+ Tile_X3Y9_LUT4AB/N4BEG[5] Tile_X3Y9_LUT4AB/N4BEG[6] Tile_X3Y9_LUT4AB/N4BEG[7] Tile_X3Y9_LUT4AB/N4BEG[8]
+ Tile_X3Y9_LUT4AB/N4BEG[9] Tile_X3Y9_LUT4AB/N4END[0] Tile_X3Y9_LUT4AB/N4END[10] Tile_X3Y9_LUT4AB/N4END[11]
+ Tile_X3Y9_LUT4AB/N4END[12] Tile_X3Y9_LUT4AB/N4END[13] Tile_X3Y9_LUT4AB/N4END[14]
+ Tile_X3Y9_LUT4AB/N4END[15] Tile_X3Y9_LUT4AB/N4END[1] Tile_X3Y9_LUT4AB/N4END[2] Tile_X3Y9_LUT4AB/N4END[3]
+ Tile_X3Y9_LUT4AB/N4END[4] Tile_X3Y9_LUT4AB/N4END[5] Tile_X3Y9_LUT4AB/N4END[6] Tile_X3Y9_LUT4AB/N4END[7]
+ Tile_X3Y9_LUT4AB/N4END[8] Tile_X3Y9_LUT4AB/N4END[9] Tile_X3Y9_LUT4AB/NN4BEG[0] Tile_X3Y9_LUT4AB/NN4BEG[10]
+ Tile_X3Y9_LUT4AB/NN4BEG[11] Tile_X3Y9_LUT4AB/NN4BEG[12] Tile_X3Y9_LUT4AB/NN4BEG[13]
+ Tile_X3Y9_LUT4AB/NN4BEG[14] Tile_X3Y9_LUT4AB/NN4BEG[15] Tile_X3Y9_LUT4AB/NN4BEG[1]
+ Tile_X3Y9_LUT4AB/NN4BEG[2] Tile_X3Y9_LUT4AB/NN4BEG[3] Tile_X3Y9_LUT4AB/NN4BEG[4]
+ Tile_X3Y9_LUT4AB/NN4BEG[5] Tile_X3Y9_LUT4AB/NN4BEG[6] Tile_X3Y9_LUT4AB/NN4BEG[7]
+ Tile_X3Y9_LUT4AB/NN4BEG[8] Tile_X3Y9_LUT4AB/NN4BEG[9] Tile_X3Y9_LUT4AB/NN4END[0]
+ Tile_X3Y9_LUT4AB/NN4END[10] Tile_X3Y9_LUT4AB/NN4END[11] Tile_X3Y9_LUT4AB/NN4END[12]
+ Tile_X3Y9_LUT4AB/NN4END[13] Tile_X3Y9_LUT4AB/NN4END[14] Tile_X3Y9_LUT4AB/NN4END[15]
+ Tile_X3Y9_LUT4AB/NN4END[1] Tile_X3Y9_LUT4AB/NN4END[2] Tile_X3Y9_LUT4AB/NN4END[3]
+ Tile_X3Y9_LUT4AB/NN4END[4] Tile_X3Y9_LUT4AB/NN4END[5] Tile_X3Y9_LUT4AB/NN4END[6]
+ Tile_X3Y9_LUT4AB/NN4END[7] Tile_X3Y9_LUT4AB/NN4END[8] Tile_X3Y9_LUT4AB/NN4END[9]
+ Tile_X3Y9_LUT4AB/S1BEG[0] Tile_X3Y9_LUT4AB/S1BEG[1] Tile_X3Y9_LUT4AB/S1BEG[2] Tile_X3Y9_LUT4AB/S1BEG[3]
+ Tile_X3Y9_LUT4AB/S1END[0] Tile_X3Y9_LUT4AB/S1END[1] Tile_X3Y9_LUT4AB/S1END[2] Tile_X3Y9_LUT4AB/S1END[3]
+ Tile_X3Y9_LUT4AB/S2BEG[0] Tile_X3Y9_LUT4AB/S2BEG[1] Tile_X3Y9_LUT4AB/S2BEG[2] Tile_X3Y9_LUT4AB/S2BEG[3]
+ Tile_X3Y9_LUT4AB/S2BEG[4] Tile_X3Y9_LUT4AB/S2BEG[5] Tile_X3Y9_LUT4AB/S2BEG[6] Tile_X3Y9_LUT4AB/S2BEG[7]
+ Tile_X3Y9_LUT4AB/S2BEGb[0] Tile_X3Y9_LUT4AB/S2BEGb[1] Tile_X3Y9_LUT4AB/S2BEGb[2]
+ Tile_X3Y9_LUT4AB/S2BEGb[3] Tile_X3Y9_LUT4AB/S2BEGb[4] Tile_X3Y9_LUT4AB/S2BEGb[5]
+ Tile_X3Y9_LUT4AB/S2BEGb[6] Tile_X3Y9_LUT4AB/S2BEGb[7] Tile_X3Y9_LUT4AB/S2END[0]
+ Tile_X3Y9_LUT4AB/S2END[1] Tile_X3Y9_LUT4AB/S2END[2] Tile_X3Y9_LUT4AB/S2END[3] Tile_X3Y9_LUT4AB/S2END[4]
+ Tile_X3Y9_LUT4AB/S2END[5] Tile_X3Y9_LUT4AB/S2END[6] Tile_X3Y9_LUT4AB/S2END[7] Tile_X3Y9_LUT4AB/S2MID[0]
+ Tile_X3Y9_LUT4AB/S2MID[1] Tile_X3Y9_LUT4AB/S2MID[2] Tile_X3Y9_LUT4AB/S2MID[3] Tile_X3Y9_LUT4AB/S2MID[4]
+ Tile_X3Y9_LUT4AB/S2MID[5] Tile_X3Y9_LUT4AB/S2MID[6] Tile_X3Y9_LUT4AB/S2MID[7] Tile_X3Y9_LUT4AB/S4BEG[0]
+ Tile_X3Y9_LUT4AB/S4BEG[10] Tile_X3Y9_LUT4AB/S4BEG[11] Tile_X3Y9_LUT4AB/S4BEG[12]
+ Tile_X3Y9_LUT4AB/S4BEG[13] Tile_X3Y9_LUT4AB/S4BEG[14] Tile_X3Y9_LUT4AB/S4BEG[15]
+ Tile_X3Y9_LUT4AB/S4BEG[1] Tile_X3Y9_LUT4AB/S4BEG[2] Tile_X3Y9_LUT4AB/S4BEG[3] Tile_X3Y9_LUT4AB/S4BEG[4]
+ Tile_X3Y9_LUT4AB/S4BEG[5] Tile_X3Y9_LUT4AB/S4BEG[6] Tile_X3Y9_LUT4AB/S4BEG[7] Tile_X3Y9_LUT4AB/S4BEG[8]
+ Tile_X3Y9_LUT4AB/S4BEG[9] Tile_X3Y9_LUT4AB/S4END[0] Tile_X3Y9_LUT4AB/S4END[10] Tile_X3Y9_LUT4AB/S4END[11]
+ Tile_X3Y9_LUT4AB/S4END[12] Tile_X3Y9_LUT4AB/S4END[13] Tile_X3Y9_LUT4AB/S4END[14]
+ Tile_X3Y9_LUT4AB/S4END[15] Tile_X3Y9_LUT4AB/S4END[1] Tile_X3Y9_LUT4AB/S4END[2] Tile_X3Y9_LUT4AB/S4END[3]
+ Tile_X3Y9_LUT4AB/S4END[4] Tile_X3Y9_LUT4AB/S4END[5] Tile_X3Y9_LUT4AB/S4END[6] Tile_X3Y9_LUT4AB/S4END[7]
+ Tile_X3Y9_LUT4AB/S4END[8] Tile_X3Y9_LUT4AB/S4END[9] Tile_X3Y9_LUT4AB/SS4BEG[0] Tile_X3Y9_LUT4AB/SS4BEG[10]
+ Tile_X3Y9_LUT4AB/SS4BEG[11] Tile_X3Y9_LUT4AB/SS4BEG[12] Tile_X3Y9_LUT4AB/SS4BEG[13]
+ Tile_X3Y9_LUT4AB/SS4BEG[14] Tile_X3Y9_LUT4AB/SS4BEG[15] Tile_X3Y9_LUT4AB/SS4BEG[1]
+ Tile_X3Y9_LUT4AB/SS4BEG[2] Tile_X3Y9_LUT4AB/SS4BEG[3] Tile_X3Y9_LUT4AB/SS4BEG[4]
+ Tile_X3Y9_LUT4AB/SS4BEG[5] Tile_X3Y9_LUT4AB/SS4BEG[6] Tile_X3Y9_LUT4AB/SS4BEG[7]
+ Tile_X3Y9_LUT4AB/SS4BEG[8] Tile_X3Y9_LUT4AB/SS4BEG[9] Tile_X3Y9_LUT4AB/SS4END[0]
+ Tile_X3Y9_LUT4AB/SS4END[10] Tile_X3Y9_LUT4AB/SS4END[11] Tile_X3Y9_LUT4AB/SS4END[12]
+ Tile_X3Y9_LUT4AB/SS4END[13] Tile_X3Y9_LUT4AB/SS4END[14] Tile_X3Y9_LUT4AB/SS4END[15]
+ Tile_X3Y9_LUT4AB/SS4END[1] Tile_X3Y9_LUT4AB/SS4END[2] Tile_X3Y9_LUT4AB/SS4END[3]
+ Tile_X3Y9_LUT4AB/SS4END[4] Tile_X3Y9_LUT4AB/SS4END[5] Tile_X3Y9_LUT4AB/SS4END[6]
+ Tile_X3Y9_LUT4AB/SS4END[7] Tile_X3Y9_LUT4AB/SS4END[8] Tile_X3Y9_LUT4AB/SS4END[9]
+ Tile_X3Y9_LUT4AB/UserCLK Tile_X3Y8_LUT4AB/UserCLK VGND VPWR Tile_X3Y9_LUT4AB/W1BEG[0]
+ Tile_X3Y9_LUT4AB/W1BEG[1] Tile_X3Y9_LUT4AB/W1BEG[2] Tile_X3Y9_LUT4AB/W1BEG[3] Tile_X3Y9_LUT4AB/W1END[0]
+ Tile_X3Y9_LUT4AB/W1END[1] Tile_X3Y9_LUT4AB/W1END[2] Tile_X3Y9_LUT4AB/W1END[3] Tile_X3Y9_LUT4AB/W2BEG[0]
+ Tile_X3Y9_LUT4AB/W2BEG[1] Tile_X3Y9_LUT4AB/W2BEG[2] Tile_X3Y9_LUT4AB/W2BEG[3] Tile_X3Y9_LUT4AB/W2BEG[4]
+ Tile_X3Y9_LUT4AB/W2BEG[5] Tile_X3Y9_LUT4AB/W2BEG[6] Tile_X3Y9_LUT4AB/W2BEG[7] Tile_X2Y9_LUT4AB/W2END[0]
+ Tile_X2Y9_LUT4AB/W2END[1] Tile_X2Y9_LUT4AB/W2END[2] Tile_X2Y9_LUT4AB/W2END[3] Tile_X2Y9_LUT4AB/W2END[4]
+ Tile_X2Y9_LUT4AB/W2END[5] Tile_X2Y9_LUT4AB/W2END[6] Tile_X2Y9_LUT4AB/W2END[7] Tile_X3Y9_LUT4AB/W2END[0]
+ Tile_X3Y9_LUT4AB/W2END[1] Tile_X3Y9_LUT4AB/W2END[2] Tile_X3Y9_LUT4AB/W2END[3] Tile_X3Y9_LUT4AB/W2END[4]
+ Tile_X3Y9_LUT4AB/W2END[5] Tile_X3Y9_LUT4AB/W2END[6] Tile_X3Y9_LUT4AB/W2END[7] Tile_X3Y9_LUT4AB/W2MID[0]
+ Tile_X3Y9_LUT4AB/W2MID[1] Tile_X3Y9_LUT4AB/W2MID[2] Tile_X3Y9_LUT4AB/W2MID[3] Tile_X3Y9_LUT4AB/W2MID[4]
+ Tile_X3Y9_LUT4AB/W2MID[5] Tile_X3Y9_LUT4AB/W2MID[6] Tile_X3Y9_LUT4AB/W2MID[7] Tile_X3Y9_LUT4AB/W6BEG[0]
+ Tile_X3Y9_LUT4AB/W6BEG[10] Tile_X3Y9_LUT4AB/W6BEG[11] Tile_X3Y9_LUT4AB/W6BEG[1]
+ Tile_X3Y9_LUT4AB/W6BEG[2] Tile_X3Y9_LUT4AB/W6BEG[3] Tile_X3Y9_LUT4AB/W6BEG[4] Tile_X3Y9_LUT4AB/W6BEG[5]
+ Tile_X3Y9_LUT4AB/W6BEG[6] Tile_X3Y9_LUT4AB/W6BEG[7] Tile_X3Y9_LUT4AB/W6BEG[8] Tile_X3Y9_LUT4AB/W6BEG[9]
+ Tile_X3Y9_LUT4AB/W6END[0] Tile_X3Y9_LUT4AB/W6END[10] Tile_X3Y9_LUT4AB/W6END[11]
+ Tile_X3Y9_LUT4AB/W6END[1] Tile_X3Y9_LUT4AB/W6END[2] Tile_X3Y9_LUT4AB/W6END[3] Tile_X3Y9_LUT4AB/W6END[4]
+ Tile_X3Y9_LUT4AB/W6END[5] Tile_X3Y9_LUT4AB/W6END[6] Tile_X3Y9_LUT4AB/W6END[7] Tile_X3Y9_LUT4AB/W6END[8]
+ Tile_X3Y9_LUT4AB/W6END[9] Tile_X3Y9_LUT4AB/WW4BEG[0] Tile_X3Y9_LUT4AB/WW4BEG[10]
+ Tile_X3Y9_LUT4AB/WW4BEG[11] Tile_X3Y9_LUT4AB/WW4BEG[12] Tile_X3Y9_LUT4AB/WW4BEG[13]
+ Tile_X3Y9_LUT4AB/WW4BEG[14] Tile_X3Y9_LUT4AB/WW4BEG[15] Tile_X3Y9_LUT4AB/WW4BEG[1]
+ Tile_X3Y9_LUT4AB/WW4BEG[2] Tile_X3Y9_LUT4AB/WW4BEG[3] Tile_X3Y9_LUT4AB/WW4BEG[4]
+ Tile_X3Y9_LUT4AB/WW4BEG[5] Tile_X3Y9_LUT4AB/WW4BEG[6] Tile_X3Y9_LUT4AB/WW4BEG[7]
+ Tile_X3Y9_LUT4AB/WW4BEG[8] Tile_X3Y9_LUT4AB/WW4BEG[9] Tile_X3Y9_LUT4AB/WW4END[0]
+ Tile_X3Y9_LUT4AB/WW4END[10] Tile_X3Y9_LUT4AB/WW4END[11] Tile_X3Y9_LUT4AB/WW4END[12]
+ Tile_X3Y9_LUT4AB/WW4END[13] Tile_X3Y9_LUT4AB/WW4END[14] Tile_X3Y9_LUT4AB/WW4END[15]
+ Tile_X3Y9_LUT4AB/WW4END[1] Tile_X3Y9_LUT4AB/WW4END[2] Tile_X3Y9_LUT4AB/WW4END[3]
+ Tile_X3Y9_LUT4AB/WW4END[4] Tile_X3Y9_LUT4AB/WW4END[5] Tile_X3Y9_LUT4AB/WW4END[6]
+ Tile_X3Y9_LUT4AB/WW4END[7] Tile_X3Y9_LUT4AB/WW4END[8] Tile_X3Y9_LUT4AB/WW4END[9]
+ LUT4AB
XTile_X7Y11_DSP Tile_X8Y11_LUT4AB/E1END[0] Tile_X8Y11_LUT4AB/E1END[1] Tile_X8Y11_LUT4AB/E1END[2]
+ Tile_X8Y11_LUT4AB/E1END[3] Tile_X6Y11_LUT4AB/E1BEG[0] Tile_X6Y11_LUT4AB/E1BEG[1]
+ Tile_X6Y11_LUT4AB/E1BEG[2] Tile_X6Y11_LUT4AB/E1BEG[3] Tile_X8Y11_LUT4AB/E2MID[0]
+ Tile_X8Y11_LUT4AB/E2MID[1] Tile_X8Y11_LUT4AB/E2MID[2] Tile_X8Y11_LUT4AB/E2MID[3]
+ Tile_X8Y11_LUT4AB/E2MID[4] Tile_X8Y11_LUT4AB/E2MID[5] Tile_X8Y11_LUT4AB/E2MID[6]
+ Tile_X8Y11_LUT4AB/E2MID[7] Tile_X8Y11_LUT4AB/E2END[0] Tile_X8Y11_LUT4AB/E2END[1]
+ Tile_X8Y11_LUT4AB/E2END[2] Tile_X8Y11_LUT4AB/E2END[3] Tile_X8Y11_LUT4AB/E2END[4]
+ Tile_X8Y11_LUT4AB/E2END[5] Tile_X8Y11_LUT4AB/E2END[6] Tile_X8Y11_LUT4AB/E2END[7]
+ Tile_X6Y11_LUT4AB/E2BEGb[0] Tile_X6Y11_LUT4AB/E2BEGb[1] Tile_X6Y11_LUT4AB/E2BEGb[2]
+ Tile_X6Y11_LUT4AB/E2BEGb[3] Tile_X6Y11_LUT4AB/E2BEGb[4] Tile_X6Y11_LUT4AB/E2BEGb[5]
+ Tile_X6Y11_LUT4AB/E2BEGb[6] Tile_X6Y11_LUT4AB/E2BEGb[7] Tile_X6Y11_LUT4AB/E2BEG[0]
+ Tile_X6Y11_LUT4AB/E2BEG[1] Tile_X6Y11_LUT4AB/E2BEG[2] Tile_X6Y11_LUT4AB/E2BEG[3]
+ Tile_X6Y11_LUT4AB/E2BEG[4] Tile_X6Y11_LUT4AB/E2BEG[5] Tile_X6Y11_LUT4AB/E2BEG[6]
+ Tile_X6Y11_LUT4AB/E2BEG[7] Tile_X8Y11_LUT4AB/E6END[0] Tile_X8Y11_LUT4AB/E6END[10]
+ Tile_X8Y11_LUT4AB/E6END[11] Tile_X8Y11_LUT4AB/E6END[1] Tile_X8Y11_LUT4AB/E6END[2]
+ Tile_X8Y11_LUT4AB/E6END[3] Tile_X8Y11_LUT4AB/E6END[4] Tile_X8Y11_LUT4AB/E6END[5]
+ Tile_X8Y11_LUT4AB/E6END[6] Tile_X8Y11_LUT4AB/E6END[7] Tile_X8Y11_LUT4AB/E6END[8]
+ Tile_X8Y11_LUT4AB/E6END[9] Tile_X6Y11_LUT4AB/E6BEG[0] Tile_X6Y11_LUT4AB/E6BEG[10]
+ Tile_X6Y11_LUT4AB/E6BEG[11] Tile_X6Y11_LUT4AB/E6BEG[1] Tile_X6Y11_LUT4AB/E6BEG[2]
+ Tile_X6Y11_LUT4AB/E6BEG[3] Tile_X6Y11_LUT4AB/E6BEG[4] Tile_X6Y11_LUT4AB/E6BEG[5]
+ Tile_X6Y11_LUT4AB/E6BEG[6] Tile_X6Y11_LUT4AB/E6BEG[7] Tile_X6Y11_LUT4AB/E6BEG[8]
+ Tile_X6Y11_LUT4AB/E6BEG[9] Tile_X8Y11_LUT4AB/EE4END[0] Tile_X8Y11_LUT4AB/EE4END[10]
+ Tile_X8Y11_LUT4AB/EE4END[11] Tile_X8Y11_LUT4AB/EE4END[12] Tile_X8Y11_LUT4AB/EE4END[13]
+ Tile_X8Y11_LUT4AB/EE4END[14] Tile_X8Y11_LUT4AB/EE4END[15] Tile_X8Y11_LUT4AB/EE4END[1]
+ Tile_X8Y11_LUT4AB/EE4END[2] Tile_X8Y11_LUT4AB/EE4END[3] Tile_X8Y11_LUT4AB/EE4END[4]
+ Tile_X8Y11_LUT4AB/EE4END[5] Tile_X8Y11_LUT4AB/EE4END[6] Tile_X8Y11_LUT4AB/EE4END[7]
+ Tile_X8Y11_LUT4AB/EE4END[8] Tile_X8Y11_LUT4AB/EE4END[9] Tile_X6Y11_LUT4AB/EE4BEG[0]
+ Tile_X6Y11_LUT4AB/EE4BEG[10] Tile_X6Y11_LUT4AB/EE4BEG[11] Tile_X6Y11_LUT4AB/EE4BEG[12]
+ Tile_X6Y11_LUT4AB/EE4BEG[13] Tile_X6Y11_LUT4AB/EE4BEG[14] Tile_X6Y11_LUT4AB/EE4BEG[15]
+ Tile_X6Y11_LUT4AB/EE4BEG[1] Tile_X6Y11_LUT4AB/EE4BEG[2] Tile_X6Y11_LUT4AB/EE4BEG[3]
+ Tile_X6Y11_LUT4AB/EE4BEG[4] Tile_X6Y11_LUT4AB/EE4BEG[5] Tile_X6Y11_LUT4AB/EE4BEG[6]
+ Tile_X6Y11_LUT4AB/EE4BEG[7] Tile_X6Y11_LUT4AB/EE4BEG[8] Tile_X6Y11_LUT4AB/EE4BEG[9]
+ Tile_X6Y11_LUT4AB/FrameData_O[0] Tile_X6Y11_LUT4AB/FrameData_O[10] Tile_X6Y11_LUT4AB/FrameData_O[11]
+ Tile_X6Y11_LUT4AB/FrameData_O[12] Tile_X6Y11_LUT4AB/FrameData_O[13] Tile_X6Y11_LUT4AB/FrameData_O[14]
+ Tile_X6Y11_LUT4AB/FrameData_O[15] Tile_X6Y11_LUT4AB/FrameData_O[16] Tile_X6Y11_LUT4AB/FrameData_O[17]
+ Tile_X6Y11_LUT4AB/FrameData_O[18] Tile_X6Y11_LUT4AB/FrameData_O[19] Tile_X6Y11_LUT4AB/FrameData_O[1]
+ Tile_X6Y11_LUT4AB/FrameData_O[20] Tile_X6Y11_LUT4AB/FrameData_O[21] Tile_X6Y11_LUT4AB/FrameData_O[22]
+ Tile_X6Y11_LUT4AB/FrameData_O[23] Tile_X6Y11_LUT4AB/FrameData_O[24] Tile_X6Y11_LUT4AB/FrameData_O[25]
+ Tile_X6Y11_LUT4AB/FrameData_O[26] Tile_X6Y11_LUT4AB/FrameData_O[27] Tile_X6Y11_LUT4AB/FrameData_O[28]
+ Tile_X6Y11_LUT4AB/FrameData_O[29] Tile_X6Y11_LUT4AB/FrameData_O[2] Tile_X6Y11_LUT4AB/FrameData_O[30]
+ Tile_X6Y11_LUT4AB/FrameData_O[31] Tile_X6Y11_LUT4AB/FrameData_O[3] Tile_X6Y11_LUT4AB/FrameData_O[4]
+ Tile_X6Y11_LUT4AB/FrameData_O[5] Tile_X6Y11_LUT4AB/FrameData_O[6] Tile_X6Y11_LUT4AB/FrameData_O[7]
+ Tile_X6Y11_LUT4AB/FrameData_O[8] Tile_X6Y11_LUT4AB/FrameData_O[9] Tile_X8Y11_LUT4AB/FrameData[0]
+ Tile_X8Y11_LUT4AB/FrameData[10] Tile_X8Y11_LUT4AB/FrameData[11] Tile_X8Y11_LUT4AB/FrameData[12]
+ Tile_X8Y11_LUT4AB/FrameData[13] Tile_X8Y11_LUT4AB/FrameData[14] Tile_X8Y11_LUT4AB/FrameData[15]
+ Tile_X8Y11_LUT4AB/FrameData[16] Tile_X8Y11_LUT4AB/FrameData[17] Tile_X8Y11_LUT4AB/FrameData[18]
+ Tile_X8Y11_LUT4AB/FrameData[19] Tile_X8Y11_LUT4AB/FrameData[1] Tile_X8Y11_LUT4AB/FrameData[20]
+ Tile_X8Y11_LUT4AB/FrameData[21] Tile_X8Y11_LUT4AB/FrameData[22] Tile_X8Y11_LUT4AB/FrameData[23]
+ Tile_X8Y11_LUT4AB/FrameData[24] Tile_X8Y11_LUT4AB/FrameData[25] Tile_X8Y11_LUT4AB/FrameData[26]
+ Tile_X8Y11_LUT4AB/FrameData[27] Tile_X8Y11_LUT4AB/FrameData[28] Tile_X8Y11_LUT4AB/FrameData[29]
+ Tile_X8Y11_LUT4AB/FrameData[2] Tile_X8Y11_LUT4AB/FrameData[30] Tile_X8Y11_LUT4AB/FrameData[31]
+ Tile_X8Y11_LUT4AB/FrameData[3] Tile_X8Y11_LUT4AB/FrameData[4] Tile_X8Y11_LUT4AB/FrameData[5]
+ Tile_X8Y11_LUT4AB/FrameData[6] Tile_X8Y11_LUT4AB/FrameData[7] Tile_X8Y11_LUT4AB/FrameData[8]
+ Tile_X8Y11_LUT4AB/FrameData[9] Tile_X7Y9_DSP/Tile_X0Y1_FrameStrobe[0] Tile_X7Y9_DSP/Tile_X0Y1_FrameStrobe[10]
+ Tile_X7Y9_DSP/Tile_X0Y1_FrameStrobe[11] Tile_X7Y9_DSP/Tile_X0Y1_FrameStrobe[12]
+ Tile_X7Y9_DSP/Tile_X0Y1_FrameStrobe[13] Tile_X7Y9_DSP/Tile_X0Y1_FrameStrobe[14]
+ Tile_X7Y9_DSP/Tile_X0Y1_FrameStrobe[15] Tile_X7Y9_DSP/Tile_X0Y1_FrameStrobe[16]
+ Tile_X7Y9_DSP/Tile_X0Y1_FrameStrobe[17] Tile_X7Y9_DSP/Tile_X0Y1_FrameStrobe[18]
+ Tile_X7Y9_DSP/Tile_X0Y1_FrameStrobe[19] Tile_X7Y9_DSP/Tile_X0Y1_FrameStrobe[1] Tile_X7Y9_DSP/Tile_X0Y1_FrameStrobe[2]
+ Tile_X7Y9_DSP/Tile_X0Y1_FrameStrobe[3] Tile_X7Y9_DSP/Tile_X0Y1_FrameStrobe[4] Tile_X7Y9_DSP/Tile_X0Y1_FrameStrobe[5]
+ Tile_X7Y9_DSP/Tile_X0Y1_FrameStrobe[6] Tile_X7Y9_DSP/Tile_X0Y1_FrameStrobe[7] Tile_X7Y9_DSP/Tile_X0Y1_FrameStrobe[8]
+ Tile_X7Y9_DSP/Tile_X0Y1_FrameStrobe[9] Tile_X7Y9_DSP/Tile_X0Y1_N1END[0] Tile_X7Y9_DSP/Tile_X0Y1_N1END[1]
+ Tile_X7Y9_DSP/Tile_X0Y1_N1END[2] Tile_X7Y9_DSP/Tile_X0Y1_N1END[3] Tile_X7Y9_DSP/Tile_X0Y1_N2MID[0]
+ Tile_X7Y9_DSP/Tile_X0Y1_N2MID[1] Tile_X7Y9_DSP/Tile_X0Y1_N2MID[2] Tile_X7Y9_DSP/Tile_X0Y1_N2MID[3]
+ Tile_X7Y9_DSP/Tile_X0Y1_N2MID[4] Tile_X7Y9_DSP/Tile_X0Y1_N2MID[5] Tile_X7Y9_DSP/Tile_X0Y1_N2MID[6]
+ Tile_X7Y9_DSP/Tile_X0Y1_N2MID[7] Tile_X7Y9_DSP/Tile_X0Y1_N2END[0] Tile_X7Y9_DSP/Tile_X0Y1_N2END[1]
+ Tile_X7Y9_DSP/Tile_X0Y1_N2END[2] Tile_X7Y9_DSP/Tile_X0Y1_N2END[3] Tile_X7Y9_DSP/Tile_X0Y1_N2END[4]
+ Tile_X7Y9_DSP/Tile_X0Y1_N2END[5] Tile_X7Y9_DSP/Tile_X0Y1_N2END[6] Tile_X7Y9_DSP/Tile_X0Y1_N2END[7]
+ Tile_X7Y9_DSP/Tile_X0Y1_N4END[0] Tile_X7Y9_DSP/Tile_X0Y1_N4END[10] Tile_X7Y9_DSP/Tile_X0Y1_N4END[11]
+ Tile_X7Y9_DSP/Tile_X0Y1_N4END[12] Tile_X7Y9_DSP/Tile_X0Y1_N4END[13] Tile_X7Y9_DSP/Tile_X0Y1_N4END[14]
+ Tile_X7Y9_DSP/Tile_X0Y1_N4END[15] Tile_X7Y9_DSP/Tile_X0Y1_N4END[1] Tile_X7Y9_DSP/Tile_X0Y1_N4END[2]
+ Tile_X7Y9_DSP/Tile_X0Y1_N4END[3] Tile_X7Y9_DSP/Tile_X0Y1_N4END[4] Tile_X7Y9_DSP/Tile_X0Y1_N4END[5]
+ Tile_X7Y9_DSP/Tile_X0Y1_N4END[6] Tile_X7Y9_DSP/Tile_X0Y1_N4END[7] Tile_X7Y9_DSP/Tile_X0Y1_N4END[8]
+ Tile_X7Y9_DSP/Tile_X0Y1_N4END[9] Tile_X7Y9_DSP/Tile_X0Y1_NN4END[0] Tile_X7Y9_DSP/Tile_X0Y1_NN4END[10]
+ Tile_X7Y9_DSP/Tile_X0Y1_NN4END[11] Tile_X7Y9_DSP/Tile_X0Y1_NN4END[12] Tile_X7Y9_DSP/Tile_X0Y1_NN4END[13]
+ Tile_X7Y9_DSP/Tile_X0Y1_NN4END[14] Tile_X7Y9_DSP/Tile_X0Y1_NN4END[15] Tile_X7Y9_DSP/Tile_X0Y1_NN4END[1]
+ Tile_X7Y9_DSP/Tile_X0Y1_NN4END[2] Tile_X7Y9_DSP/Tile_X0Y1_NN4END[3] Tile_X7Y9_DSP/Tile_X0Y1_NN4END[4]
+ Tile_X7Y9_DSP/Tile_X0Y1_NN4END[5] Tile_X7Y9_DSP/Tile_X0Y1_NN4END[6] Tile_X7Y9_DSP/Tile_X0Y1_NN4END[7]
+ Tile_X7Y9_DSP/Tile_X0Y1_NN4END[8] Tile_X7Y9_DSP/Tile_X0Y1_NN4END[9] Tile_X7Y9_DSP/Tile_X0Y1_S1BEG[0]
+ Tile_X7Y9_DSP/Tile_X0Y1_S1BEG[1] Tile_X7Y9_DSP/Tile_X0Y1_S1BEG[2] Tile_X7Y9_DSP/Tile_X0Y1_S1BEG[3]
+ Tile_X7Y9_DSP/Tile_X0Y1_S2BEGb[0] Tile_X7Y9_DSP/Tile_X0Y1_S2BEGb[1] Tile_X7Y9_DSP/Tile_X0Y1_S2BEGb[2]
+ Tile_X7Y9_DSP/Tile_X0Y1_S2BEGb[3] Tile_X7Y9_DSP/Tile_X0Y1_S2BEGb[4] Tile_X7Y9_DSP/Tile_X0Y1_S2BEGb[5]
+ Tile_X7Y9_DSP/Tile_X0Y1_S2BEGb[6] Tile_X7Y9_DSP/Tile_X0Y1_S2BEGb[7] Tile_X7Y9_DSP/Tile_X0Y1_S2BEG[0]
+ Tile_X7Y9_DSP/Tile_X0Y1_S2BEG[1] Tile_X7Y9_DSP/Tile_X0Y1_S2BEG[2] Tile_X7Y9_DSP/Tile_X0Y1_S2BEG[3]
+ Tile_X7Y9_DSP/Tile_X0Y1_S2BEG[4] Tile_X7Y9_DSP/Tile_X0Y1_S2BEG[5] Tile_X7Y9_DSP/Tile_X0Y1_S2BEG[6]
+ Tile_X7Y9_DSP/Tile_X0Y1_S2BEG[7] Tile_X7Y9_DSP/Tile_X0Y1_S4BEG[0] Tile_X7Y9_DSP/Tile_X0Y1_S4BEG[10]
+ Tile_X7Y9_DSP/Tile_X0Y1_S4BEG[11] Tile_X7Y9_DSP/Tile_X0Y1_S4BEG[12] Tile_X7Y9_DSP/Tile_X0Y1_S4BEG[13]
+ Tile_X7Y9_DSP/Tile_X0Y1_S4BEG[14] Tile_X7Y9_DSP/Tile_X0Y1_S4BEG[15] Tile_X7Y9_DSP/Tile_X0Y1_S4BEG[1]
+ Tile_X7Y9_DSP/Tile_X0Y1_S4BEG[2] Tile_X7Y9_DSP/Tile_X0Y1_S4BEG[3] Tile_X7Y9_DSP/Tile_X0Y1_S4BEG[4]
+ Tile_X7Y9_DSP/Tile_X0Y1_S4BEG[5] Tile_X7Y9_DSP/Tile_X0Y1_S4BEG[6] Tile_X7Y9_DSP/Tile_X0Y1_S4BEG[7]
+ Tile_X7Y9_DSP/Tile_X0Y1_S4BEG[8] Tile_X7Y9_DSP/Tile_X0Y1_S4BEG[9] Tile_X7Y9_DSP/Tile_X0Y1_SS4BEG[0]
+ Tile_X7Y9_DSP/Tile_X0Y1_SS4BEG[10] Tile_X7Y9_DSP/Tile_X0Y1_SS4BEG[11] Tile_X7Y9_DSP/Tile_X0Y1_SS4BEG[12]
+ Tile_X7Y9_DSP/Tile_X0Y1_SS4BEG[13] Tile_X7Y9_DSP/Tile_X0Y1_SS4BEG[14] Tile_X7Y9_DSP/Tile_X0Y1_SS4BEG[15]
+ Tile_X7Y9_DSP/Tile_X0Y1_SS4BEG[1] Tile_X7Y9_DSP/Tile_X0Y1_SS4BEG[2] Tile_X7Y9_DSP/Tile_X0Y1_SS4BEG[3]
+ Tile_X7Y9_DSP/Tile_X0Y1_SS4BEG[4] Tile_X7Y9_DSP/Tile_X0Y1_SS4BEG[5] Tile_X7Y9_DSP/Tile_X0Y1_SS4BEG[6]
+ Tile_X7Y9_DSP/Tile_X0Y1_SS4BEG[7] Tile_X7Y9_DSP/Tile_X0Y1_SS4BEG[8] Tile_X7Y9_DSP/Tile_X0Y1_SS4BEG[9]
+ Tile_X7Y9_DSP/Tile_X0Y1_UserCLK Tile_X6Y11_LUT4AB/W1END[0] Tile_X6Y11_LUT4AB/W1END[1]
+ Tile_X6Y11_LUT4AB/W1END[2] Tile_X6Y11_LUT4AB/W1END[3] Tile_X8Y11_LUT4AB/W1BEG[0]
+ Tile_X8Y11_LUT4AB/W1BEG[1] Tile_X8Y11_LUT4AB/W1BEG[2] Tile_X8Y11_LUT4AB/W1BEG[3]
+ Tile_X6Y11_LUT4AB/W2MID[0] Tile_X6Y11_LUT4AB/W2MID[1] Tile_X6Y11_LUT4AB/W2MID[2]
+ Tile_X6Y11_LUT4AB/W2MID[3] Tile_X6Y11_LUT4AB/W2MID[4] Tile_X6Y11_LUT4AB/W2MID[5]
+ Tile_X6Y11_LUT4AB/W2MID[6] Tile_X6Y11_LUT4AB/W2MID[7] Tile_X6Y11_LUT4AB/W2END[0]
+ Tile_X6Y11_LUT4AB/W2END[1] Tile_X6Y11_LUT4AB/W2END[2] Tile_X6Y11_LUT4AB/W2END[3]
+ Tile_X6Y11_LUT4AB/W2END[4] Tile_X6Y11_LUT4AB/W2END[5] Tile_X6Y11_LUT4AB/W2END[6]
+ Tile_X6Y11_LUT4AB/W2END[7] Tile_X8Y11_LUT4AB/W2BEGb[0] Tile_X8Y11_LUT4AB/W2BEGb[1]
+ Tile_X8Y11_LUT4AB/W2BEGb[2] Tile_X8Y11_LUT4AB/W2BEGb[3] Tile_X8Y11_LUT4AB/W2BEGb[4]
+ Tile_X8Y11_LUT4AB/W2BEGb[5] Tile_X8Y11_LUT4AB/W2BEGb[6] Tile_X8Y11_LUT4AB/W2BEGb[7]
+ Tile_X8Y11_LUT4AB/W2BEG[0] Tile_X8Y11_LUT4AB/W2BEG[1] Tile_X8Y11_LUT4AB/W2BEG[2]
+ Tile_X8Y11_LUT4AB/W2BEG[3] Tile_X8Y11_LUT4AB/W2BEG[4] Tile_X8Y11_LUT4AB/W2BEG[5]
+ Tile_X8Y11_LUT4AB/W2BEG[6] Tile_X8Y11_LUT4AB/W2BEG[7] Tile_X6Y11_LUT4AB/W6END[0]
+ Tile_X6Y11_LUT4AB/W6END[10] Tile_X6Y11_LUT4AB/W6END[11] Tile_X6Y11_LUT4AB/W6END[1]
+ Tile_X6Y11_LUT4AB/W6END[2] Tile_X6Y11_LUT4AB/W6END[3] Tile_X6Y11_LUT4AB/W6END[4]
+ Tile_X6Y11_LUT4AB/W6END[5] Tile_X6Y11_LUT4AB/W6END[6] Tile_X6Y11_LUT4AB/W6END[7]
+ Tile_X6Y11_LUT4AB/W6END[8] Tile_X6Y11_LUT4AB/W6END[9] Tile_X8Y11_LUT4AB/W6BEG[0]
+ Tile_X8Y11_LUT4AB/W6BEG[10] Tile_X8Y11_LUT4AB/W6BEG[11] Tile_X8Y11_LUT4AB/W6BEG[1]
+ Tile_X8Y11_LUT4AB/W6BEG[2] Tile_X8Y11_LUT4AB/W6BEG[3] Tile_X8Y11_LUT4AB/W6BEG[4]
+ Tile_X8Y11_LUT4AB/W6BEG[5] Tile_X8Y11_LUT4AB/W6BEG[6] Tile_X8Y11_LUT4AB/W6BEG[7]
+ Tile_X8Y11_LUT4AB/W6BEG[8] Tile_X8Y11_LUT4AB/W6BEG[9] Tile_X6Y11_LUT4AB/WW4END[0]
+ Tile_X6Y11_LUT4AB/WW4END[10] Tile_X6Y11_LUT4AB/WW4END[11] Tile_X6Y11_LUT4AB/WW4END[12]
+ Tile_X6Y11_LUT4AB/WW4END[13] Tile_X6Y11_LUT4AB/WW4END[14] Tile_X6Y11_LUT4AB/WW4END[15]
+ Tile_X6Y11_LUT4AB/WW4END[1] Tile_X6Y11_LUT4AB/WW4END[2] Tile_X6Y11_LUT4AB/WW4END[3]
+ Tile_X6Y11_LUT4AB/WW4END[4] Tile_X6Y11_LUT4AB/WW4END[5] Tile_X6Y11_LUT4AB/WW4END[6]
+ Tile_X6Y11_LUT4AB/WW4END[7] Tile_X6Y11_LUT4AB/WW4END[8] Tile_X6Y11_LUT4AB/WW4END[9]
+ Tile_X8Y11_LUT4AB/WW4BEG[0] Tile_X8Y11_LUT4AB/WW4BEG[10] Tile_X8Y11_LUT4AB/WW4BEG[11]
+ Tile_X8Y11_LUT4AB/WW4BEG[12] Tile_X8Y11_LUT4AB/WW4BEG[13] Tile_X8Y11_LUT4AB/WW4BEG[14]
+ Tile_X8Y11_LUT4AB/WW4BEG[15] Tile_X8Y11_LUT4AB/WW4BEG[1] Tile_X8Y11_LUT4AB/WW4BEG[2]
+ Tile_X8Y11_LUT4AB/WW4BEG[3] Tile_X8Y11_LUT4AB/WW4BEG[4] Tile_X8Y11_LUT4AB/WW4BEG[5]
+ Tile_X8Y11_LUT4AB/WW4BEG[6] Tile_X8Y11_LUT4AB/WW4BEG[7] Tile_X8Y11_LUT4AB/WW4BEG[8]
+ Tile_X8Y11_LUT4AB/WW4BEG[9] Tile_X8Y12_LUT4AB/E1END[0] Tile_X8Y12_LUT4AB/E1END[1]
+ Tile_X8Y12_LUT4AB/E1END[2] Tile_X8Y12_LUT4AB/E1END[3] Tile_X6Y12_LUT4AB/E1BEG[0]
+ Tile_X6Y12_LUT4AB/E1BEG[1] Tile_X6Y12_LUT4AB/E1BEG[2] Tile_X6Y12_LUT4AB/E1BEG[3]
+ Tile_X8Y12_LUT4AB/E2MID[0] Tile_X8Y12_LUT4AB/E2MID[1] Tile_X8Y12_LUT4AB/E2MID[2]
+ Tile_X8Y12_LUT4AB/E2MID[3] Tile_X8Y12_LUT4AB/E2MID[4] Tile_X8Y12_LUT4AB/E2MID[5]
+ Tile_X8Y12_LUT4AB/E2MID[6] Tile_X8Y12_LUT4AB/E2MID[7] Tile_X8Y12_LUT4AB/E2END[0]
+ Tile_X8Y12_LUT4AB/E2END[1] Tile_X8Y12_LUT4AB/E2END[2] Tile_X8Y12_LUT4AB/E2END[3]
+ Tile_X8Y12_LUT4AB/E2END[4] Tile_X8Y12_LUT4AB/E2END[5] Tile_X8Y12_LUT4AB/E2END[6]
+ Tile_X8Y12_LUT4AB/E2END[7] Tile_X6Y12_LUT4AB/E2BEGb[0] Tile_X6Y12_LUT4AB/E2BEGb[1]
+ Tile_X6Y12_LUT4AB/E2BEGb[2] Tile_X6Y12_LUT4AB/E2BEGb[3] Tile_X6Y12_LUT4AB/E2BEGb[4]
+ Tile_X6Y12_LUT4AB/E2BEGb[5] Tile_X6Y12_LUT4AB/E2BEGb[6] Tile_X6Y12_LUT4AB/E2BEGb[7]
+ Tile_X6Y12_LUT4AB/E2BEG[0] Tile_X6Y12_LUT4AB/E2BEG[1] Tile_X6Y12_LUT4AB/E2BEG[2]
+ Tile_X6Y12_LUT4AB/E2BEG[3] Tile_X6Y12_LUT4AB/E2BEG[4] Tile_X6Y12_LUT4AB/E2BEG[5]
+ Tile_X6Y12_LUT4AB/E2BEG[6] Tile_X6Y12_LUT4AB/E2BEG[7] Tile_X8Y12_LUT4AB/E6END[0]
+ Tile_X8Y12_LUT4AB/E6END[10] Tile_X8Y12_LUT4AB/E6END[11] Tile_X8Y12_LUT4AB/E6END[1]
+ Tile_X8Y12_LUT4AB/E6END[2] Tile_X8Y12_LUT4AB/E6END[3] Tile_X8Y12_LUT4AB/E6END[4]
+ Tile_X8Y12_LUT4AB/E6END[5] Tile_X8Y12_LUT4AB/E6END[6] Tile_X8Y12_LUT4AB/E6END[7]
+ Tile_X8Y12_LUT4AB/E6END[8] Tile_X8Y12_LUT4AB/E6END[9] Tile_X6Y12_LUT4AB/E6BEG[0]
+ Tile_X6Y12_LUT4AB/E6BEG[10] Tile_X6Y12_LUT4AB/E6BEG[11] Tile_X6Y12_LUT4AB/E6BEG[1]
+ Tile_X6Y12_LUT4AB/E6BEG[2] Tile_X6Y12_LUT4AB/E6BEG[3] Tile_X6Y12_LUT4AB/E6BEG[4]
+ Tile_X6Y12_LUT4AB/E6BEG[5] Tile_X6Y12_LUT4AB/E6BEG[6] Tile_X6Y12_LUT4AB/E6BEG[7]
+ Tile_X6Y12_LUT4AB/E6BEG[8] Tile_X6Y12_LUT4AB/E6BEG[9] Tile_X8Y12_LUT4AB/EE4END[0]
+ Tile_X8Y12_LUT4AB/EE4END[10] Tile_X8Y12_LUT4AB/EE4END[11] Tile_X8Y12_LUT4AB/EE4END[12]
+ Tile_X8Y12_LUT4AB/EE4END[13] Tile_X8Y12_LUT4AB/EE4END[14] Tile_X8Y12_LUT4AB/EE4END[15]
+ Tile_X8Y12_LUT4AB/EE4END[1] Tile_X8Y12_LUT4AB/EE4END[2] Tile_X8Y12_LUT4AB/EE4END[3]
+ Tile_X8Y12_LUT4AB/EE4END[4] Tile_X8Y12_LUT4AB/EE4END[5] Tile_X8Y12_LUT4AB/EE4END[6]
+ Tile_X8Y12_LUT4AB/EE4END[7] Tile_X8Y12_LUT4AB/EE4END[8] Tile_X8Y12_LUT4AB/EE4END[9]
+ Tile_X6Y12_LUT4AB/EE4BEG[0] Tile_X6Y12_LUT4AB/EE4BEG[10] Tile_X6Y12_LUT4AB/EE4BEG[11]
+ Tile_X6Y12_LUT4AB/EE4BEG[12] Tile_X6Y12_LUT4AB/EE4BEG[13] Tile_X6Y12_LUT4AB/EE4BEG[14]
+ Tile_X6Y12_LUT4AB/EE4BEG[15] Tile_X6Y12_LUT4AB/EE4BEG[1] Tile_X6Y12_LUT4AB/EE4BEG[2]
+ Tile_X6Y12_LUT4AB/EE4BEG[3] Tile_X6Y12_LUT4AB/EE4BEG[4] Tile_X6Y12_LUT4AB/EE4BEG[5]
+ Tile_X6Y12_LUT4AB/EE4BEG[6] Tile_X6Y12_LUT4AB/EE4BEG[7] Tile_X6Y12_LUT4AB/EE4BEG[8]
+ Tile_X6Y12_LUT4AB/EE4BEG[9] Tile_X6Y12_LUT4AB/FrameData_O[0] Tile_X6Y12_LUT4AB/FrameData_O[10]
+ Tile_X6Y12_LUT4AB/FrameData_O[11] Tile_X6Y12_LUT4AB/FrameData_O[12] Tile_X6Y12_LUT4AB/FrameData_O[13]
+ Tile_X6Y12_LUT4AB/FrameData_O[14] Tile_X6Y12_LUT4AB/FrameData_O[15] Tile_X6Y12_LUT4AB/FrameData_O[16]
+ Tile_X6Y12_LUT4AB/FrameData_O[17] Tile_X6Y12_LUT4AB/FrameData_O[18] Tile_X6Y12_LUT4AB/FrameData_O[19]
+ Tile_X6Y12_LUT4AB/FrameData_O[1] Tile_X6Y12_LUT4AB/FrameData_O[20] Tile_X6Y12_LUT4AB/FrameData_O[21]
+ Tile_X6Y12_LUT4AB/FrameData_O[22] Tile_X6Y12_LUT4AB/FrameData_O[23] Tile_X6Y12_LUT4AB/FrameData_O[24]
+ Tile_X6Y12_LUT4AB/FrameData_O[25] Tile_X6Y12_LUT4AB/FrameData_O[26] Tile_X6Y12_LUT4AB/FrameData_O[27]
+ Tile_X6Y12_LUT4AB/FrameData_O[28] Tile_X6Y12_LUT4AB/FrameData_O[29] Tile_X6Y12_LUT4AB/FrameData_O[2]
+ Tile_X6Y12_LUT4AB/FrameData_O[30] Tile_X6Y12_LUT4AB/FrameData_O[31] Tile_X6Y12_LUT4AB/FrameData_O[3]
+ Tile_X6Y12_LUT4AB/FrameData_O[4] Tile_X6Y12_LUT4AB/FrameData_O[5] Tile_X6Y12_LUT4AB/FrameData_O[6]
+ Tile_X6Y12_LUT4AB/FrameData_O[7] Tile_X6Y12_LUT4AB/FrameData_O[8] Tile_X6Y12_LUT4AB/FrameData_O[9]
+ Tile_X8Y12_LUT4AB/FrameData[0] Tile_X8Y12_LUT4AB/FrameData[10] Tile_X8Y12_LUT4AB/FrameData[11]
+ Tile_X8Y12_LUT4AB/FrameData[12] Tile_X8Y12_LUT4AB/FrameData[13] Tile_X8Y12_LUT4AB/FrameData[14]
+ Tile_X8Y12_LUT4AB/FrameData[15] Tile_X8Y12_LUT4AB/FrameData[16] Tile_X8Y12_LUT4AB/FrameData[17]
+ Tile_X8Y12_LUT4AB/FrameData[18] Tile_X8Y12_LUT4AB/FrameData[19] Tile_X8Y12_LUT4AB/FrameData[1]
+ Tile_X8Y12_LUT4AB/FrameData[20] Tile_X8Y12_LUT4AB/FrameData[21] Tile_X8Y12_LUT4AB/FrameData[22]
+ Tile_X8Y12_LUT4AB/FrameData[23] Tile_X8Y12_LUT4AB/FrameData[24] Tile_X8Y12_LUT4AB/FrameData[25]
+ Tile_X8Y12_LUT4AB/FrameData[26] Tile_X8Y12_LUT4AB/FrameData[27] Tile_X8Y12_LUT4AB/FrameData[28]
+ Tile_X8Y12_LUT4AB/FrameData[29] Tile_X8Y12_LUT4AB/FrameData[2] Tile_X8Y12_LUT4AB/FrameData[30]
+ Tile_X8Y12_LUT4AB/FrameData[31] Tile_X8Y12_LUT4AB/FrameData[3] Tile_X8Y12_LUT4AB/FrameData[4]
+ Tile_X8Y12_LUT4AB/FrameData[5] Tile_X8Y12_LUT4AB/FrameData[6] Tile_X8Y12_LUT4AB/FrameData[7]
+ Tile_X8Y12_LUT4AB/FrameData[8] Tile_X8Y12_LUT4AB/FrameData[9] Tile_X7Y11_DSP/Tile_X0Y1_FrameStrobe[0]
+ Tile_X7Y11_DSP/Tile_X0Y1_FrameStrobe[10] Tile_X7Y11_DSP/Tile_X0Y1_FrameStrobe[11]
+ Tile_X7Y11_DSP/Tile_X0Y1_FrameStrobe[12] Tile_X7Y11_DSP/Tile_X0Y1_FrameStrobe[13]
+ Tile_X7Y11_DSP/Tile_X0Y1_FrameStrobe[14] Tile_X7Y11_DSP/Tile_X0Y1_FrameStrobe[15]
+ Tile_X7Y11_DSP/Tile_X0Y1_FrameStrobe[16] Tile_X7Y11_DSP/Tile_X0Y1_FrameStrobe[17]
+ Tile_X7Y11_DSP/Tile_X0Y1_FrameStrobe[18] Tile_X7Y11_DSP/Tile_X0Y1_FrameStrobe[19]
+ Tile_X7Y11_DSP/Tile_X0Y1_FrameStrobe[1] Tile_X7Y11_DSP/Tile_X0Y1_FrameStrobe[2]
+ Tile_X7Y11_DSP/Tile_X0Y1_FrameStrobe[3] Tile_X7Y11_DSP/Tile_X0Y1_FrameStrobe[4]
+ Tile_X7Y11_DSP/Tile_X0Y1_FrameStrobe[5] Tile_X7Y11_DSP/Tile_X0Y1_FrameStrobe[6]
+ Tile_X7Y11_DSP/Tile_X0Y1_FrameStrobe[7] Tile_X7Y11_DSP/Tile_X0Y1_FrameStrobe[8]
+ Tile_X7Y11_DSP/Tile_X0Y1_FrameStrobe[9] Tile_X7Y13_DSP/Tile_X0Y0_N1BEG[0] Tile_X7Y13_DSP/Tile_X0Y0_N1BEG[1]
+ Tile_X7Y13_DSP/Tile_X0Y0_N1BEG[2] Tile_X7Y13_DSP/Tile_X0Y0_N1BEG[3] Tile_X7Y11_DSP/Tile_X0Y1_N2END[0]
+ Tile_X7Y11_DSP/Tile_X0Y1_N2END[1] Tile_X7Y11_DSP/Tile_X0Y1_N2END[2] Tile_X7Y11_DSP/Tile_X0Y1_N2END[3]
+ Tile_X7Y11_DSP/Tile_X0Y1_N2END[4] Tile_X7Y11_DSP/Tile_X0Y1_N2END[5] Tile_X7Y11_DSP/Tile_X0Y1_N2END[6]
+ Tile_X7Y11_DSP/Tile_X0Y1_N2END[7] Tile_X7Y13_DSP/Tile_X0Y0_N2BEG[0] Tile_X7Y13_DSP/Tile_X0Y0_N2BEG[1]
+ Tile_X7Y13_DSP/Tile_X0Y0_N2BEG[2] Tile_X7Y13_DSP/Tile_X0Y0_N2BEG[3] Tile_X7Y13_DSP/Tile_X0Y0_N2BEG[4]
+ Tile_X7Y13_DSP/Tile_X0Y0_N2BEG[5] Tile_X7Y13_DSP/Tile_X0Y0_N2BEG[6] Tile_X7Y13_DSP/Tile_X0Y0_N2BEG[7]
+ Tile_X7Y13_DSP/Tile_X0Y0_N4BEG[0] Tile_X7Y13_DSP/Tile_X0Y0_N4BEG[10] Tile_X7Y13_DSP/Tile_X0Y0_N4BEG[11]
+ Tile_X7Y13_DSP/Tile_X0Y0_N4BEG[12] Tile_X7Y13_DSP/Tile_X0Y0_N4BEG[13] Tile_X7Y13_DSP/Tile_X0Y0_N4BEG[14]
+ Tile_X7Y13_DSP/Tile_X0Y0_N4BEG[15] Tile_X7Y13_DSP/Tile_X0Y0_N4BEG[1] Tile_X7Y13_DSP/Tile_X0Y0_N4BEG[2]
+ Tile_X7Y13_DSP/Tile_X0Y0_N4BEG[3] Tile_X7Y13_DSP/Tile_X0Y0_N4BEG[4] Tile_X7Y13_DSP/Tile_X0Y0_N4BEG[5]
+ Tile_X7Y13_DSP/Tile_X0Y0_N4BEG[6] Tile_X7Y13_DSP/Tile_X0Y0_N4BEG[7] Tile_X7Y13_DSP/Tile_X0Y0_N4BEG[8]
+ Tile_X7Y13_DSP/Tile_X0Y0_N4BEG[9] Tile_X7Y13_DSP/Tile_X0Y0_NN4BEG[0] Tile_X7Y13_DSP/Tile_X0Y0_NN4BEG[10]
+ Tile_X7Y13_DSP/Tile_X0Y0_NN4BEG[11] Tile_X7Y13_DSP/Tile_X0Y0_NN4BEG[12] Tile_X7Y13_DSP/Tile_X0Y0_NN4BEG[13]
+ Tile_X7Y13_DSP/Tile_X0Y0_NN4BEG[14] Tile_X7Y13_DSP/Tile_X0Y0_NN4BEG[15] Tile_X7Y13_DSP/Tile_X0Y0_NN4BEG[1]
+ Tile_X7Y13_DSP/Tile_X0Y0_NN4BEG[2] Tile_X7Y13_DSP/Tile_X0Y0_NN4BEG[3] Tile_X7Y13_DSP/Tile_X0Y0_NN4BEG[4]
+ Tile_X7Y13_DSP/Tile_X0Y0_NN4BEG[5] Tile_X7Y13_DSP/Tile_X0Y0_NN4BEG[6] Tile_X7Y13_DSP/Tile_X0Y0_NN4BEG[7]
+ Tile_X7Y13_DSP/Tile_X0Y0_NN4BEG[8] Tile_X7Y13_DSP/Tile_X0Y0_NN4BEG[9] Tile_X7Y13_DSP/Tile_X0Y0_S1END[0]
+ Tile_X7Y13_DSP/Tile_X0Y0_S1END[1] Tile_X7Y13_DSP/Tile_X0Y0_S1END[2] Tile_X7Y13_DSP/Tile_X0Y0_S1END[3]
+ Tile_X7Y13_DSP/Tile_X0Y0_S2MID[0] Tile_X7Y13_DSP/Tile_X0Y0_S2MID[1] Tile_X7Y13_DSP/Tile_X0Y0_S2MID[2]
+ Tile_X7Y13_DSP/Tile_X0Y0_S2MID[3] Tile_X7Y13_DSP/Tile_X0Y0_S2MID[4] Tile_X7Y13_DSP/Tile_X0Y0_S2MID[5]
+ Tile_X7Y13_DSP/Tile_X0Y0_S2MID[6] Tile_X7Y13_DSP/Tile_X0Y0_S2MID[7] Tile_X7Y13_DSP/Tile_X0Y0_S2END[0]
+ Tile_X7Y13_DSP/Tile_X0Y0_S2END[1] Tile_X7Y13_DSP/Tile_X0Y0_S2END[2] Tile_X7Y13_DSP/Tile_X0Y0_S2END[3]
+ Tile_X7Y13_DSP/Tile_X0Y0_S2END[4] Tile_X7Y13_DSP/Tile_X0Y0_S2END[5] Tile_X7Y13_DSP/Tile_X0Y0_S2END[6]
+ Tile_X7Y13_DSP/Tile_X0Y0_S2END[7] Tile_X7Y13_DSP/Tile_X0Y0_S4END[0] Tile_X7Y13_DSP/Tile_X0Y0_S4END[10]
+ Tile_X7Y13_DSP/Tile_X0Y0_S4END[11] Tile_X7Y13_DSP/Tile_X0Y0_S4END[12] Tile_X7Y13_DSP/Tile_X0Y0_S4END[13]
+ Tile_X7Y13_DSP/Tile_X0Y0_S4END[14] Tile_X7Y13_DSP/Tile_X0Y0_S4END[15] Tile_X7Y13_DSP/Tile_X0Y0_S4END[1]
+ Tile_X7Y13_DSP/Tile_X0Y0_S4END[2] Tile_X7Y13_DSP/Tile_X0Y0_S4END[3] Tile_X7Y13_DSP/Tile_X0Y0_S4END[4]
+ Tile_X7Y13_DSP/Tile_X0Y0_S4END[5] Tile_X7Y13_DSP/Tile_X0Y0_S4END[6] Tile_X7Y13_DSP/Tile_X0Y0_S4END[7]
+ Tile_X7Y13_DSP/Tile_X0Y0_S4END[8] Tile_X7Y13_DSP/Tile_X0Y0_S4END[9] Tile_X7Y13_DSP/Tile_X0Y0_SS4END[0]
+ Tile_X7Y13_DSP/Tile_X0Y0_SS4END[10] Tile_X7Y13_DSP/Tile_X0Y0_SS4END[11] Tile_X7Y13_DSP/Tile_X0Y0_SS4END[12]
+ Tile_X7Y13_DSP/Tile_X0Y0_SS4END[13] Tile_X7Y13_DSP/Tile_X0Y0_SS4END[14] Tile_X7Y13_DSP/Tile_X0Y0_SS4END[15]
+ Tile_X7Y13_DSP/Tile_X0Y0_SS4END[1] Tile_X7Y13_DSP/Tile_X0Y0_SS4END[2] Tile_X7Y13_DSP/Tile_X0Y0_SS4END[3]
+ Tile_X7Y13_DSP/Tile_X0Y0_SS4END[4] Tile_X7Y13_DSP/Tile_X0Y0_SS4END[5] Tile_X7Y13_DSP/Tile_X0Y0_SS4END[6]
+ Tile_X7Y13_DSP/Tile_X0Y0_SS4END[7] Tile_X7Y13_DSP/Tile_X0Y0_SS4END[8] Tile_X7Y13_DSP/Tile_X0Y0_SS4END[9]
+ Tile_X7Y11_DSP/Tile_X0Y1_UserCLK Tile_X6Y12_LUT4AB/W1END[0] Tile_X6Y12_LUT4AB/W1END[1]
+ Tile_X6Y12_LUT4AB/W1END[2] Tile_X6Y12_LUT4AB/W1END[3] Tile_X8Y12_LUT4AB/W1BEG[0]
+ Tile_X8Y12_LUT4AB/W1BEG[1] Tile_X8Y12_LUT4AB/W1BEG[2] Tile_X8Y12_LUT4AB/W1BEG[3]
+ Tile_X6Y12_LUT4AB/W2MID[0] Tile_X6Y12_LUT4AB/W2MID[1] Tile_X6Y12_LUT4AB/W2MID[2]
+ Tile_X6Y12_LUT4AB/W2MID[3] Tile_X6Y12_LUT4AB/W2MID[4] Tile_X6Y12_LUT4AB/W2MID[5]
+ Tile_X6Y12_LUT4AB/W2MID[6] Tile_X6Y12_LUT4AB/W2MID[7] Tile_X6Y12_LUT4AB/W2END[0]
+ Tile_X6Y12_LUT4AB/W2END[1] Tile_X6Y12_LUT4AB/W2END[2] Tile_X6Y12_LUT4AB/W2END[3]
+ Tile_X6Y12_LUT4AB/W2END[4] Tile_X6Y12_LUT4AB/W2END[5] Tile_X6Y12_LUT4AB/W2END[6]
+ Tile_X6Y12_LUT4AB/W2END[7] Tile_X8Y12_LUT4AB/W2BEGb[0] Tile_X8Y12_LUT4AB/W2BEGb[1]
+ Tile_X8Y12_LUT4AB/W2BEGb[2] Tile_X8Y12_LUT4AB/W2BEGb[3] Tile_X8Y12_LUT4AB/W2BEGb[4]
+ Tile_X8Y12_LUT4AB/W2BEGb[5] Tile_X8Y12_LUT4AB/W2BEGb[6] Tile_X8Y12_LUT4AB/W2BEGb[7]
+ Tile_X8Y12_LUT4AB/W2BEG[0] Tile_X8Y12_LUT4AB/W2BEG[1] Tile_X8Y12_LUT4AB/W2BEG[2]
+ Tile_X8Y12_LUT4AB/W2BEG[3] Tile_X8Y12_LUT4AB/W2BEG[4] Tile_X8Y12_LUT4AB/W2BEG[5]
+ Tile_X8Y12_LUT4AB/W2BEG[6] Tile_X8Y12_LUT4AB/W2BEG[7] Tile_X6Y12_LUT4AB/W6END[0]
+ Tile_X6Y12_LUT4AB/W6END[10] Tile_X6Y12_LUT4AB/W6END[11] Tile_X6Y12_LUT4AB/W6END[1]
+ Tile_X6Y12_LUT4AB/W6END[2] Tile_X6Y12_LUT4AB/W6END[3] Tile_X6Y12_LUT4AB/W6END[4]
+ Tile_X6Y12_LUT4AB/W6END[5] Tile_X6Y12_LUT4AB/W6END[6] Tile_X6Y12_LUT4AB/W6END[7]
+ Tile_X6Y12_LUT4AB/W6END[8] Tile_X6Y12_LUT4AB/W6END[9] Tile_X8Y12_LUT4AB/W6BEG[0]
+ Tile_X8Y12_LUT4AB/W6BEG[10] Tile_X8Y12_LUT4AB/W6BEG[11] Tile_X8Y12_LUT4AB/W6BEG[1]
+ Tile_X8Y12_LUT4AB/W6BEG[2] Tile_X8Y12_LUT4AB/W6BEG[3] Tile_X8Y12_LUT4AB/W6BEG[4]
+ Tile_X8Y12_LUT4AB/W6BEG[5] Tile_X8Y12_LUT4AB/W6BEG[6] Tile_X8Y12_LUT4AB/W6BEG[7]
+ Tile_X8Y12_LUT4AB/W6BEG[8] Tile_X8Y12_LUT4AB/W6BEG[9] Tile_X6Y12_LUT4AB/WW4END[0]
+ Tile_X6Y12_LUT4AB/WW4END[10] Tile_X6Y12_LUT4AB/WW4END[11] Tile_X6Y12_LUT4AB/WW4END[12]
+ Tile_X6Y12_LUT4AB/WW4END[13] Tile_X6Y12_LUT4AB/WW4END[14] Tile_X6Y12_LUT4AB/WW4END[15]
+ Tile_X6Y12_LUT4AB/WW4END[1] Tile_X6Y12_LUT4AB/WW4END[2] Tile_X6Y12_LUT4AB/WW4END[3]
+ Tile_X6Y12_LUT4AB/WW4END[4] Tile_X6Y12_LUT4AB/WW4END[5] Tile_X6Y12_LUT4AB/WW4END[6]
+ Tile_X6Y12_LUT4AB/WW4END[7] Tile_X6Y12_LUT4AB/WW4END[8] Tile_X6Y12_LUT4AB/WW4END[9]
+ Tile_X8Y12_LUT4AB/WW4BEG[0] Tile_X8Y12_LUT4AB/WW4BEG[10] Tile_X8Y12_LUT4AB/WW4BEG[11]
+ Tile_X8Y12_LUT4AB/WW4BEG[12] Tile_X8Y12_LUT4AB/WW4BEG[13] Tile_X8Y12_LUT4AB/WW4BEG[14]
+ Tile_X8Y12_LUT4AB/WW4BEG[15] Tile_X8Y12_LUT4AB/WW4BEG[1] Tile_X8Y12_LUT4AB/WW4BEG[2]
+ Tile_X8Y12_LUT4AB/WW4BEG[3] Tile_X8Y12_LUT4AB/WW4BEG[4] Tile_X8Y12_LUT4AB/WW4BEG[5]
+ Tile_X8Y12_LUT4AB/WW4BEG[6] Tile_X8Y12_LUT4AB/WW4BEG[7] Tile_X8Y12_LUT4AB/WW4BEG[8]
+ Tile_X8Y12_LUT4AB/WW4BEG[9] VGND VPWR DSP
XTile_X9Y8_LUT4AB Tile_X9Y9_LUT4AB/Co Tile_X9Y8_LUT4AB/Co Tile_X9Y8_LUT4AB/E1BEG[0]
+ Tile_X9Y8_LUT4AB/E1BEG[1] Tile_X9Y8_LUT4AB/E1BEG[2] Tile_X9Y8_LUT4AB/E1BEG[3] Tile_X9Y8_LUT4AB/E1END[0]
+ Tile_X9Y8_LUT4AB/E1END[1] Tile_X9Y8_LUT4AB/E1END[2] Tile_X9Y8_LUT4AB/E1END[3] Tile_X9Y8_LUT4AB/E2BEG[0]
+ Tile_X9Y8_LUT4AB/E2BEG[1] Tile_X9Y8_LUT4AB/E2BEG[2] Tile_X9Y8_LUT4AB/E2BEG[3] Tile_X9Y8_LUT4AB/E2BEG[4]
+ Tile_X9Y8_LUT4AB/E2BEG[5] Tile_X9Y8_LUT4AB/E2BEG[6] Tile_X9Y8_LUT4AB/E2BEG[7] Tile_X9Y8_LUT4AB/E2BEGb[0]
+ Tile_X9Y8_LUT4AB/E2BEGb[1] Tile_X9Y8_LUT4AB/E2BEGb[2] Tile_X9Y8_LUT4AB/E2BEGb[3]
+ Tile_X9Y8_LUT4AB/E2BEGb[4] Tile_X9Y8_LUT4AB/E2BEGb[5] Tile_X9Y8_LUT4AB/E2BEGb[6]
+ Tile_X9Y8_LUT4AB/E2BEGb[7] Tile_X9Y8_LUT4AB/E2END[0] Tile_X9Y8_LUT4AB/E2END[1] Tile_X9Y8_LUT4AB/E2END[2]
+ Tile_X9Y8_LUT4AB/E2END[3] Tile_X9Y8_LUT4AB/E2END[4] Tile_X9Y8_LUT4AB/E2END[5] Tile_X9Y8_LUT4AB/E2END[6]
+ Tile_X9Y8_LUT4AB/E2END[7] Tile_X9Y8_LUT4AB/E2MID[0] Tile_X9Y8_LUT4AB/E2MID[1] Tile_X9Y8_LUT4AB/E2MID[2]
+ Tile_X9Y8_LUT4AB/E2MID[3] Tile_X9Y8_LUT4AB/E2MID[4] Tile_X9Y8_LUT4AB/E2MID[5] Tile_X9Y8_LUT4AB/E2MID[6]
+ Tile_X9Y8_LUT4AB/E2MID[7] Tile_X9Y8_LUT4AB/E6BEG[0] Tile_X9Y8_LUT4AB/E6BEG[10] Tile_X9Y8_LUT4AB/E6BEG[11]
+ Tile_X9Y8_LUT4AB/E6BEG[1] Tile_X9Y8_LUT4AB/E6BEG[2] Tile_X9Y8_LUT4AB/E6BEG[3] Tile_X9Y8_LUT4AB/E6BEG[4]
+ Tile_X9Y8_LUT4AB/E6BEG[5] Tile_X9Y8_LUT4AB/E6BEG[6] Tile_X9Y8_LUT4AB/E6BEG[7] Tile_X9Y8_LUT4AB/E6BEG[8]
+ Tile_X9Y8_LUT4AB/E6BEG[9] Tile_X9Y8_LUT4AB/E6END[0] Tile_X9Y8_LUT4AB/E6END[10] Tile_X9Y8_LUT4AB/E6END[11]
+ Tile_X9Y8_LUT4AB/E6END[1] Tile_X9Y8_LUT4AB/E6END[2] Tile_X9Y8_LUT4AB/E6END[3] Tile_X9Y8_LUT4AB/E6END[4]
+ Tile_X9Y8_LUT4AB/E6END[5] Tile_X9Y8_LUT4AB/E6END[6] Tile_X9Y8_LUT4AB/E6END[7] Tile_X9Y8_LUT4AB/E6END[8]
+ Tile_X9Y8_LUT4AB/E6END[9] Tile_X9Y8_LUT4AB/EE4BEG[0] Tile_X9Y8_LUT4AB/EE4BEG[10]
+ Tile_X9Y8_LUT4AB/EE4BEG[11] Tile_X9Y8_LUT4AB/EE4BEG[12] Tile_X9Y8_LUT4AB/EE4BEG[13]
+ Tile_X9Y8_LUT4AB/EE4BEG[14] Tile_X9Y8_LUT4AB/EE4BEG[15] Tile_X9Y8_LUT4AB/EE4BEG[1]
+ Tile_X9Y8_LUT4AB/EE4BEG[2] Tile_X9Y8_LUT4AB/EE4BEG[3] Tile_X9Y8_LUT4AB/EE4BEG[4]
+ Tile_X9Y8_LUT4AB/EE4BEG[5] Tile_X9Y8_LUT4AB/EE4BEG[6] Tile_X9Y8_LUT4AB/EE4BEG[7]
+ Tile_X9Y8_LUT4AB/EE4BEG[8] Tile_X9Y8_LUT4AB/EE4BEG[9] Tile_X9Y8_LUT4AB/EE4END[0]
+ Tile_X9Y8_LUT4AB/EE4END[10] Tile_X9Y8_LUT4AB/EE4END[11] Tile_X9Y8_LUT4AB/EE4END[12]
+ Tile_X9Y8_LUT4AB/EE4END[13] Tile_X9Y8_LUT4AB/EE4END[14] Tile_X9Y8_LUT4AB/EE4END[15]
+ Tile_X9Y8_LUT4AB/EE4END[1] Tile_X9Y8_LUT4AB/EE4END[2] Tile_X9Y8_LUT4AB/EE4END[3]
+ Tile_X9Y8_LUT4AB/EE4END[4] Tile_X9Y8_LUT4AB/EE4END[5] Tile_X9Y8_LUT4AB/EE4END[6]
+ Tile_X9Y8_LUT4AB/EE4END[7] Tile_X9Y8_LUT4AB/EE4END[8] Tile_X9Y8_LUT4AB/EE4END[9]
+ Tile_X9Y8_LUT4AB/FrameData[0] Tile_X9Y8_LUT4AB/FrameData[10] Tile_X9Y8_LUT4AB/FrameData[11]
+ Tile_X9Y8_LUT4AB/FrameData[12] Tile_X9Y8_LUT4AB/FrameData[13] Tile_X9Y8_LUT4AB/FrameData[14]
+ Tile_X9Y8_LUT4AB/FrameData[15] Tile_X9Y8_LUT4AB/FrameData[16] Tile_X9Y8_LUT4AB/FrameData[17]
+ Tile_X9Y8_LUT4AB/FrameData[18] Tile_X9Y8_LUT4AB/FrameData[19] Tile_X9Y8_LUT4AB/FrameData[1]
+ Tile_X9Y8_LUT4AB/FrameData[20] Tile_X9Y8_LUT4AB/FrameData[21] Tile_X9Y8_LUT4AB/FrameData[22]
+ Tile_X9Y8_LUT4AB/FrameData[23] Tile_X9Y8_LUT4AB/FrameData[24] Tile_X9Y8_LUT4AB/FrameData[25]
+ Tile_X9Y8_LUT4AB/FrameData[26] Tile_X9Y8_LUT4AB/FrameData[27] Tile_X9Y8_LUT4AB/FrameData[28]
+ Tile_X9Y8_LUT4AB/FrameData[29] Tile_X9Y8_LUT4AB/FrameData[2] Tile_X9Y8_LUT4AB/FrameData[30]
+ Tile_X9Y8_LUT4AB/FrameData[31] Tile_X9Y8_LUT4AB/FrameData[3] Tile_X9Y8_LUT4AB/FrameData[4]
+ Tile_X9Y8_LUT4AB/FrameData[5] Tile_X9Y8_LUT4AB/FrameData[6] Tile_X9Y8_LUT4AB/FrameData[7]
+ Tile_X9Y8_LUT4AB/FrameData[8] Tile_X9Y8_LUT4AB/FrameData[9] Tile_X9Y8_LUT4AB/FrameData_O[0]
+ Tile_X9Y8_LUT4AB/FrameData_O[10] Tile_X9Y8_LUT4AB/FrameData_O[11] Tile_X9Y8_LUT4AB/FrameData_O[12]
+ Tile_X9Y8_LUT4AB/FrameData_O[13] Tile_X9Y8_LUT4AB/FrameData_O[14] Tile_X9Y8_LUT4AB/FrameData_O[15]
+ Tile_X9Y8_LUT4AB/FrameData_O[16] Tile_X9Y8_LUT4AB/FrameData_O[17] Tile_X9Y8_LUT4AB/FrameData_O[18]
+ Tile_X9Y8_LUT4AB/FrameData_O[19] Tile_X9Y8_LUT4AB/FrameData_O[1] Tile_X9Y8_LUT4AB/FrameData_O[20]
+ Tile_X9Y8_LUT4AB/FrameData_O[21] Tile_X9Y8_LUT4AB/FrameData_O[22] Tile_X9Y8_LUT4AB/FrameData_O[23]
+ Tile_X9Y8_LUT4AB/FrameData_O[24] Tile_X9Y8_LUT4AB/FrameData_O[25] Tile_X9Y8_LUT4AB/FrameData_O[26]
+ Tile_X9Y8_LUT4AB/FrameData_O[27] Tile_X9Y8_LUT4AB/FrameData_O[28] Tile_X9Y8_LUT4AB/FrameData_O[29]
+ Tile_X9Y8_LUT4AB/FrameData_O[2] Tile_X9Y8_LUT4AB/FrameData_O[30] Tile_X9Y8_LUT4AB/FrameData_O[31]
+ Tile_X9Y8_LUT4AB/FrameData_O[3] Tile_X9Y8_LUT4AB/FrameData_O[4] Tile_X9Y8_LUT4AB/FrameData_O[5]
+ Tile_X9Y8_LUT4AB/FrameData_O[6] Tile_X9Y8_LUT4AB/FrameData_O[7] Tile_X9Y8_LUT4AB/FrameData_O[8]
+ Tile_X9Y8_LUT4AB/FrameData_O[9] Tile_X9Y8_LUT4AB/FrameStrobe[0] Tile_X9Y8_LUT4AB/FrameStrobe[10]
+ Tile_X9Y8_LUT4AB/FrameStrobe[11] Tile_X9Y8_LUT4AB/FrameStrobe[12] Tile_X9Y8_LUT4AB/FrameStrobe[13]
+ Tile_X9Y8_LUT4AB/FrameStrobe[14] Tile_X9Y8_LUT4AB/FrameStrobe[15] Tile_X9Y8_LUT4AB/FrameStrobe[16]
+ Tile_X9Y8_LUT4AB/FrameStrobe[17] Tile_X9Y8_LUT4AB/FrameStrobe[18] Tile_X9Y8_LUT4AB/FrameStrobe[19]
+ Tile_X9Y8_LUT4AB/FrameStrobe[1] Tile_X9Y8_LUT4AB/FrameStrobe[2] Tile_X9Y8_LUT4AB/FrameStrobe[3]
+ Tile_X9Y8_LUT4AB/FrameStrobe[4] Tile_X9Y8_LUT4AB/FrameStrobe[5] Tile_X9Y8_LUT4AB/FrameStrobe[6]
+ Tile_X9Y8_LUT4AB/FrameStrobe[7] Tile_X9Y8_LUT4AB/FrameStrobe[8] Tile_X9Y8_LUT4AB/FrameStrobe[9]
+ Tile_X9Y7_LUT4AB/FrameStrobe[0] Tile_X9Y7_LUT4AB/FrameStrobe[10] Tile_X9Y7_LUT4AB/FrameStrobe[11]
+ Tile_X9Y7_LUT4AB/FrameStrobe[12] Tile_X9Y7_LUT4AB/FrameStrobe[13] Tile_X9Y7_LUT4AB/FrameStrobe[14]
+ Tile_X9Y7_LUT4AB/FrameStrobe[15] Tile_X9Y7_LUT4AB/FrameStrobe[16] Tile_X9Y7_LUT4AB/FrameStrobe[17]
+ Tile_X9Y7_LUT4AB/FrameStrobe[18] Tile_X9Y7_LUT4AB/FrameStrobe[19] Tile_X9Y7_LUT4AB/FrameStrobe[1]
+ Tile_X9Y7_LUT4AB/FrameStrobe[2] Tile_X9Y7_LUT4AB/FrameStrobe[3] Tile_X9Y7_LUT4AB/FrameStrobe[4]
+ Tile_X9Y7_LUT4AB/FrameStrobe[5] Tile_X9Y7_LUT4AB/FrameStrobe[6] Tile_X9Y7_LUT4AB/FrameStrobe[7]
+ Tile_X9Y7_LUT4AB/FrameStrobe[8] Tile_X9Y7_LUT4AB/FrameStrobe[9] Tile_X9Y8_LUT4AB/N1BEG[0]
+ Tile_X9Y8_LUT4AB/N1BEG[1] Tile_X9Y8_LUT4AB/N1BEG[2] Tile_X9Y8_LUT4AB/N1BEG[3] Tile_X9Y9_LUT4AB/N1BEG[0]
+ Tile_X9Y9_LUT4AB/N1BEG[1] Tile_X9Y9_LUT4AB/N1BEG[2] Tile_X9Y9_LUT4AB/N1BEG[3] Tile_X9Y8_LUT4AB/N2BEG[0]
+ Tile_X9Y8_LUT4AB/N2BEG[1] Tile_X9Y8_LUT4AB/N2BEG[2] Tile_X9Y8_LUT4AB/N2BEG[3] Tile_X9Y8_LUT4AB/N2BEG[4]
+ Tile_X9Y8_LUT4AB/N2BEG[5] Tile_X9Y8_LUT4AB/N2BEG[6] Tile_X9Y8_LUT4AB/N2BEG[7] Tile_X9Y7_LUT4AB/N2END[0]
+ Tile_X9Y7_LUT4AB/N2END[1] Tile_X9Y7_LUT4AB/N2END[2] Tile_X9Y7_LUT4AB/N2END[3] Tile_X9Y7_LUT4AB/N2END[4]
+ Tile_X9Y7_LUT4AB/N2END[5] Tile_X9Y7_LUT4AB/N2END[6] Tile_X9Y7_LUT4AB/N2END[7] Tile_X9Y8_LUT4AB/N2END[0]
+ Tile_X9Y8_LUT4AB/N2END[1] Tile_X9Y8_LUT4AB/N2END[2] Tile_X9Y8_LUT4AB/N2END[3] Tile_X9Y8_LUT4AB/N2END[4]
+ Tile_X9Y8_LUT4AB/N2END[5] Tile_X9Y8_LUT4AB/N2END[6] Tile_X9Y8_LUT4AB/N2END[7] Tile_X9Y9_LUT4AB/N2BEG[0]
+ Tile_X9Y9_LUT4AB/N2BEG[1] Tile_X9Y9_LUT4AB/N2BEG[2] Tile_X9Y9_LUT4AB/N2BEG[3] Tile_X9Y9_LUT4AB/N2BEG[4]
+ Tile_X9Y9_LUT4AB/N2BEG[5] Tile_X9Y9_LUT4AB/N2BEG[6] Tile_X9Y9_LUT4AB/N2BEG[7] Tile_X9Y8_LUT4AB/N4BEG[0]
+ Tile_X9Y8_LUT4AB/N4BEG[10] Tile_X9Y8_LUT4AB/N4BEG[11] Tile_X9Y8_LUT4AB/N4BEG[12]
+ Tile_X9Y8_LUT4AB/N4BEG[13] Tile_X9Y8_LUT4AB/N4BEG[14] Tile_X9Y8_LUT4AB/N4BEG[15]
+ Tile_X9Y8_LUT4AB/N4BEG[1] Tile_X9Y8_LUT4AB/N4BEG[2] Tile_X9Y8_LUT4AB/N4BEG[3] Tile_X9Y8_LUT4AB/N4BEG[4]
+ Tile_X9Y8_LUT4AB/N4BEG[5] Tile_X9Y8_LUT4AB/N4BEG[6] Tile_X9Y8_LUT4AB/N4BEG[7] Tile_X9Y8_LUT4AB/N4BEG[8]
+ Tile_X9Y8_LUT4AB/N4BEG[9] Tile_X9Y9_LUT4AB/N4BEG[0] Tile_X9Y9_LUT4AB/N4BEG[10] Tile_X9Y9_LUT4AB/N4BEG[11]
+ Tile_X9Y9_LUT4AB/N4BEG[12] Tile_X9Y9_LUT4AB/N4BEG[13] Tile_X9Y9_LUT4AB/N4BEG[14]
+ Tile_X9Y9_LUT4AB/N4BEG[15] Tile_X9Y9_LUT4AB/N4BEG[1] Tile_X9Y9_LUT4AB/N4BEG[2] Tile_X9Y9_LUT4AB/N4BEG[3]
+ Tile_X9Y9_LUT4AB/N4BEG[4] Tile_X9Y9_LUT4AB/N4BEG[5] Tile_X9Y9_LUT4AB/N4BEG[6] Tile_X9Y9_LUT4AB/N4BEG[7]
+ Tile_X9Y9_LUT4AB/N4BEG[8] Tile_X9Y9_LUT4AB/N4BEG[9] Tile_X9Y8_LUT4AB/NN4BEG[0] Tile_X9Y8_LUT4AB/NN4BEG[10]
+ Tile_X9Y8_LUT4AB/NN4BEG[11] Tile_X9Y8_LUT4AB/NN4BEG[12] Tile_X9Y8_LUT4AB/NN4BEG[13]
+ Tile_X9Y8_LUT4AB/NN4BEG[14] Tile_X9Y8_LUT4AB/NN4BEG[15] Tile_X9Y8_LUT4AB/NN4BEG[1]
+ Tile_X9Y8_LUT4AB/NN4BEG[2] Tile_X9Y8_LUT4AB/NN4BEG[3] Tile_X9Y8_LUT4AB/NN4BEG[4]
+ Tile_X9Y8_LUT4AB/NN4BEG[5] Tile_X9Y8_LUT4AB/NN4BEG[6] Tile_X9Y8_LUT4AB/NN4BEG[7]
+ Tile_X9Y8_LUT4AB/NN4BEG[8] Tile_X9Y8_LUT4AB/NN4BEG[9] Tile_X9Y9_LUT4AB/NN4BEG[0]
+ Tile_X9Y9_LUT4AB/NN4BEG[10] Tile_X9Y9_LUT4AB/NN4BEG[11] Tile_X9Y9_LUT4AB/NN4BEG[12]
+ Tile_X9Y9_LUT4AB/NN4BEG[13] Tile_X9Y9_LUT4AB/NN4BEG[14] Tile_X9Y9_LUT4AB/NN4BEG[15]
+ Tile_X9Y9_LUT4AB/NN4BEG[1] Tile_X9Y9_LUT4AB/NN4BEG[2] Tile_X9Y9_LUT4AB/NN4BEG[3]
+ Tile_X9Y9_LUT4AB/NN4BEG[4] Tile_X9Y9_LUT4AB/NN4BEG[5] Tile_X9Y9_LUT4AB/NN4BEG[6]
+ Tile_X9Y9_LUT4AB/NN4BEG[7] Tile_X9Y9_LUT4AB/NN4BEG[8] Tile_X9Y9_LUT4AB/NN4BEG[9]
+ Tile_X9Y9_LUT4AB/S1END[0] Tile_X9Y9_LUT4AB/S1END[1] Tile_X9Y9_LUT4AB/S1END[2] Tile_X9Y9_LUT4AB/S1END[3]
+ Tile_X9Y8_LUT4AB/S1END[0] Tile_X9Y8_LUT4AB/S1END[1] Tile_X9Y8_LUT4AB/S1END[2] Tile_X9Y8_LUT4AB/S1END[3]
+ Tile_X9Y9_LUT4AB/S2MID[0] Tile_X9Y9_LUT4AB/S2MID[1] Tile_X9Y9_LUT4AB/S2MID[2] Tile_X9Y9_LUT4AB/S2MID[3]
+ Tile_X9Y9_LUT4AB/S2MID[4] Tile_X9Y9_LUT4AB/S2MID[5] Tile_X9Y9_LUT4AB/S2MID[6] Tile_X9Y9_LUT4AB/S2MID[7]
+ Tile_X9Y9_LUT4AB/S2END[0] Tile_X9Y9_LUT4AB/S2END[1] Tile_X9Y9_LUT4AB/S2END[2] Tile_X9Y9_LUT4AB/S2END[3]
+ Tile_X9Y9_LUT4AB/S2END[4] Tile_X9Y9_LUT4AB/S2END[5] Tile_X9Y9_LUT4AB/S2END[6] Tile_X9Y9_LUT4AB/S2END[7]
+ Tile_X9Y8_LUT4AB/S2END[0] Tile_X9Y8_LUT4AB/S2END[1] Tile_X9Y8_LUT4AB/S2END[2] Tile_X9Y8_LUT4AB/S2END[3]
+ Tile_X9Y8_LUT4AB/S2END[4] Tile_X9Y8_LUT4AB/S2END[5] Tile_X9Y8_LUT4AB/S2END[6] Tile_X9Y8_LUT4AB/S2END[7]
+ Tile_X9Y8_LUT4AB/S2MID[0] Tile_X9Y8_LUT4AB/S2MID[1] Tile_X9Y8_LUT4AB/S2MID[2] Tile_X9Y8_LUT4AB/S2MID[3]
+ Tile_X9Y8_LUT4AB/S2MID[4] Tile_X9Y8_LUT4AB/S2MID[5] Tile_X9Y8_LUT4AB/S2MID[6] Tile_X9Y8_LUT4AB/S2MID[7]
+ Tile_X9Y9_LUT4AB/S4END[0] Tile_X9Y9_LUT4AB/S4END[10] Tile_X9Y9_LUT4AB/S4END[11]
+ Tile_X9Y9_LUT4AB/S4END[12] Tile_X9Y9_LUT4AB/S4END[13] Tile_X9Y9_LUT4AB/S4END[14]
+ Tile_X9Y9_LUT4AB/S4END[15] Tile_X9Y9_LUT4AB/S4END[1] Tile_X9Y9_LUT4AB/S4END[2] Tile_X9Y9_LUT4AB/S4END[3]
+ Tile_X9Y9_LUT4AB/S4END[4] Tile_X9Y9_LUT4AB/S4END[5] Tile_X9Y9_LUT4AB/S4END[6] Tile_X9Y9_LUT4AB/S4END[7]
+ Tile_X9Y9_LUT4AB/S4END[8] Tile_X9Y9_LUT4AB/S4END[9] Tile_X9Y8_LUT4AB/S4END[0] Tile_X9Y8_LUT4AB/S4END[10]
+ Tile_X9Y8_LUT4AB/S4END[11] Tile_X9Y8_LUT4AB/S4END[12] Tile_X9Y8_LUT4AB/S4END[13]
+ Tile_X9Y8_LUT4AB/S4END[14] Tile_X9Y8_LUT4AB/S4END[15] Tile_X9Y8_LUT4AB/S4END[1]
+ Tile_X9Y8_LUT4AB/S4END[2] Tile_X9Y8_LUT4AB/S4END[3] Tile_X9Y8_LUT4AB/S4END[4] Tile_X9Y8_LUT4AB/S4END[5]
+ Tile_X9Y8_LUT4AB/S4END[6] Tile_X9Y8_LUT4AB/S4END[7] Tile_X9Y8_LUT4AB/S4END[8] Tile_X9Y8_LUT4AB/S4END[9]
+ Tile_X9Y9_LUT4AB/SS4END[0] Tile_X9Y9_LUT4AB/SS4END[10] Tile_X9Y9_LUT4AB/SS4END[11]
+ Tile_X9Y9_LUT4AB/SS4END[12] Tile_X9Y9_LUT4AB/SS4END[13] Tile_X9Y9_LUT4AB/SS4END[14]
+ Tile_X9Y9_LUT4AB/SS4END[15] Tile_X9Y9_LUT4AB/SS4END[1] Tile_X9Y9_LUT4AB/SS4END[2]
+ Tile_X9Y9_LUT4AB/SS4END[3] Tile_X9Y9_LUT4AB/SS4END[4] Tile_X9Y9_LUT4AB/SS4END[5]
+ Tile_X9Y9_LUT4AB/SS4END[6] Tile_X9Y9_LUT4AB/SS4END[7] Tile_X9Y9_LUT4AB/SS4END[8]
+ Tile_X9Y9_LUT4AB/SS4END[9] Tile_X9Y8_LUT4AB/SS4END[0] Tile_X9Y8_LUT4AB/SS4END[10]
+ Tile_X9Y8_LUT4AB/SS4END[11] Tile_X9Y8_LUT4AB/SS4END[12] Tile_X9Y8_LUT4AB/SS4END[13]
+ Tile_X9Y8_LUT4AB/SS4END[14] Tile_X9Y8_LUT4AB/SS4END[15] Tile_X9Y8_LUT4AB/SS4END[1]
+ Tile_X9Y8_LUT4AB/SS4END[2] Tile_X9Y8_LUT4AB/SS4END[3] Tile_X9Y8_LUT4AB/SS4END[4]
+ Tile_X9Y8_LUT4AB/SS4END[5] Tile_X9Y8_LUT4AB/SS4END[6] Tile_X9Y8_LUT4AB/SS4END[7]
+ Tile_X9Y8_LUT4AB/SS4END[8] Tile_X9Y8_LUT4AB/SS4END[9] Tile_X9Y8_LUT4AB/UserCLK Tile_X9Y7_LUT4AB/UserCLK
+ VGND VPWR Tile_X9Y8_LUT4AB/W1BEG[0] Tile_X9Y8_LUT4AB/W1BEG[1] Tile_X9Y8_LUT4AB/W1BEG[2]
+ Tile_X9Y8_LUT4AB/W1BEG[3] Tile_X9Y8_LUT4AB/W1END[0] Tile_X9Y8_LUT4AB/W1END[1] Tile_X9Y8_LUT4AB/W1END[2]
+ Tile_X9Y8_LUT4AB/W1END[3] Tile_X9Y8_LUT4AB/W2BEG[0] Tile_X9Y8_LUT4AB/W2BEG[1] Tile_X9Y8_LUT4AB/W2BEG[2]
+ Tile_X9Y8_LUT4AB/W2BEG[3] Tile_X9Y8_LUT4AB/W2BEG[4] Tile_X9Y8_LUT4AB/W2BEG[5] Tile_X9Y8_LUT4AB/W2BEG[6]
+ Tile_X9Y8_LUT4AB/W2BEG[7] Tile_X8Y8_LUT4AB/W2END[0] Tile_X8Y8_LUT4AB/W2END[1] Tile_X8Y8_LUT4AB/W2END[2]
+ Tile_X8Y8_LUT4AB/W2END[3] Tile_X8Y8_LUT4AB/W2END[4] Tile_X8Y8_LUT4AB/W2END[5] Tile_X8Y8_LUT4AB/W2END[6]
+ Tile_X8Y8_LUT4AB/W2END[7] Tile_X9Y8_LUT4AB/W2END[0] Tile_X9Y8_LUT4AB/W2END[1] Tile_X9Y8_LUT4AB/W2END[2]
+ Tile_X9Y8_LUT4AB/W2END[3] Tile_X9Y8_LUT4AB/W2END[4] Tile_X9Y8_LUT4AB/W2END[5] Tile_X9Y8_LUT4AB/W2END[6]
+ Tile_X9Y8_LUT4AB/W2END[7] Tile_X9Y8_LUT4AB/W2MID[0] Tile_X9Y8_LUT4AB/W2MID[1] Tile_X9Y8_LUT4AB/W2MID[2]
+ Tile_X9Y8_LUT4AB/W2MID[3] Tile_X9Y8_LUT4AB/W2MID[4] Tile_X9Y8_LUT4AB/W2MID[5] Tile_X9Y8_LUT4AB/W2MID[6]
+ Tile_X9Y8_LUT4AB/W2MID[7] Tile_X9Y8_LUT4AB/W6BEG[0] Tile_X9Y8_LUT4AB/W6BEG[10] Tile_X9Y8_LUT4AB/W6BEG[11]
+ Tile_X9Y8_LUT4AB/W6BEG[1] Tile_X9Y8_LUT4AB/W6BEG[2] Tile_X9Y8_LUT4AB/W6BEG[3] Tile_X9Y8_LUT4AB/W6BEG[4]
+ Tile_X9Y8_LUT4AB/W6BEG[5] Tile_X9Y8_LUT4AB/W6BEG[6] Tile_X9Y8_LUT4AB/W6BEG[7] Tile_X9Y8_LUT4AB/W6BEG[8]
+ Tile_X9Y8_LUT4AB/W6BEG[9] Tile_X9Y8_LUT4AB/W6END[0] Tile_X9Y8_LUT4AB/W6END[10] Tile_X9Y8_LUT4AB/W6END[11]
+ Tile_X9Y8_LUT4AB/W6END[1] Tile_X9Y8_LUT4AB/W6END[2] Tile_X9Y8_LUT4AB/W6END[3] Tile_X9Y8_LUT4AB/W6END[4]
+ Tile_X9Y8_LUT4AB/W6END[5] Tile_X9Y8_LUT4AB/W6END[6] Tile_X9Y8_LUT4AB/W6END[7] Tile_X9Y8_LUT4AB/W6END[8]
+ Tile_X9Y8_LUT4AB/W6END[9] Tile_X9Y8_LUT4AB/WW4BEG[0] Tile_X9Y8_LUT4AB/WW4BEG[10]
+ Tile_X9Y8_LUT4AB/WW4BEG[11] Tile_X9Y8_LUT4AB/WW4BEG[12] Tile_X9Y8_LUT4AB/WW4BEG[13]
+ Tile_X9Y8_LUT4AB/WW4BEG[14] Tile_X9Y8_LUT4AB/WW4BEG[15] Tile_X9Y8_LUT4AB/WW4BEG[1]
+ Tile_X9Y8_LUT4AB/WW4BEG[2] Tile_X9Y8_LUT4AB/WW4BEG[3] Tile_X9Y8_LUT4AB/WW4BEG[4]
+ Tile_X9Y8_LUT4AB/WW4BEG[5] Tile_X9Y8_LUT4AB/WW4BEG[6] Tile_X9Y8_LUT4AB/WW4BEG[7]
+ Tile_X9Y8_LUT4AB/WW4BEG[8] Tile_X9Y8_LUT4AB/WW4BEG[9] Tile_X9Y8_LUT4AB/WW4END[0]
+ Tile_X9Y8_LUT4AB/WW4END[10] Tile_X9Y8_LUT4AB/WW4END[11] Tile_X9Y8_LUT4AB/WW4END[12]
+ Tile_X9Y8_LUT4AB/WW4END[13] Tile_X9Y8_LUT4AB/WW4END[14] Tile_X9Y8_LUT4AB/WW4END[15]
+ Tile_X9Y8_LUT4AB/WW4END[1] Tile_X9Y8_LUT4AB/WW4END[2] Tile_X9Y8_LUT4AB/WW4END[3]
+ Tile_X9Y8_LUT4AB/WW4END[4] Tile_X9Y8_LUT4AB/WW4END[5] Tile_X9Y8_LUT4AB/WW4END[6]
+ Tile_X9Y8_LUT4AB/WW4END[7] Tile_X9Y8_LUT4AB/WW4END[8] Tile_X9Y8_LUT4AB/WW4END[9]
+ LUT4AB
XTile_X6Y3_LUT4AB Tile_X6Y4_LUT4AB/Co Tile_X6Y3_LUT4AB/Co Tile_X6Y3_LUT4AB/E1BEG[0]
+ Tile_X6Y3_LUT4AB/E1BEG[1] Tile_X6Y3_LUT4AB/E1BEG[2] Tile_X6Y3_LUT4AB/E1BEG[3] Tile_X6Y3_LUT4AB/E1END[0]
+ Tile_X6Y3_LUT4AB/E1END[1] Tile_X6Y3_LUT4AB/E1END[2] Tile_X6Y3_LUT4AB/E1END[3] Tile_X6Y3_LUT4AB/E2BEG[0]
+ Tile_X6Y3_LUT4AB/E2BEG[1] Tile_X6Y3_LUT4AB/E2BEG[2] Tile_X6Y3_LUT4AB/E2BEG[3] Tile_X6Y3_LUT4AB/E2BEG[4]
+ Tile_X6Y3_LUT4AB/E2BEG[5] Tile_X6Y3_LUT4AB/E2BEG[6] Tile_X6Y3_LUT4AB/E2BEG[7] Tile_X6Y3_LUT4AB/E2BEGb[0]
+ Tile_X6Y3_LUT4AB/E2BEGb[1] Tile_X6Y3_LUT4AB/E2BEGb[2] Tile_X6Y3_LUT4AB/E2BEGb[3]
+ Tile_X6Y3_LUT4AB/E2BEGb[4] Tile_X6Y3_LUT4AB/E2BEGb[5] Tile_X6Y3_LUT4AB/E2BEGb[6]
+ Tile_X6Y3_LUT4AB/E2BEGb[7] Tile_X6Y3_LUT4AB/E2END[0] Tile_X6Y3_LUT4AB/E2END[1] Tile_X6Y3_LUT4AB/E2END[2]
+ Tile_X6Y3_LUT4AB/E2END[3] Tile_X6Y3_LUT4AB/E2END[4] Tile_X6Y3_LUT4AB/E2END[5] Tile_X6Y3_LUT4AB/E2END[6]
+ Tile_X6Y3_LUT4AB/E2END[7] Tile_X6Y3_LUT4AB/E2MID[0] Tile_X6Y3_LUT4AB/E2MID[1] Tile_X6Y3_LUT4AB/E2MID[2]
+ Tile_X6Y3_LUT4AB/E2MID[3] Tile_X6Y3_LUT4AB/E2MID[4] Tile_X6Y3_LUT4AB/E2MID[5] Tile_X6Y3_LUT4AB/E2MID[6]
+ Tile_X6Y3_LUT4AB/E2MID[7] Tile_X6Y3_LUT4AB/E6BEG[0] Tile_X6Y3_LUT4AB/E6BEG[10] Tile_X6Y3_LUT4AB/E6BEG[11]
+ Tile_X6Y3_LUT4AB/E6BEG[1] Tile_X6Y3_LUT4AB/E6BEG[2] Tile_X6Y3_LUT4AB/E6BEG[3] Tile_X6Y3_LUT4AB/E6BEG[4]
+ Tile_X6Y3_LUT4AB/E6BEG[5] Tile_X6Y3_LUT4AB/E6BEG[6] Tile_X6Y3_LUT4AB/E6BEG[7] Tile_X6Y3_LUT4AB/E6BEG[8]
+ Tile_X6Y3_LUT4AB/E6BEG[9] Tile_X6Y3_LUT4AB/E6END[0] Tile_X6Y3_LUT4AB/E6END[10] Tile_X6Y3_LUT4AB/E6END[11]
+ Tile_X6Y3_LUT4AB/E6END[1] Tile_X6Y3_LUT4AB/E6END[2] Tile_X6Y3_LUT4AB/E6END[3] Tile_X6Y3_LUT4AB/E6END[4]
+ Tile_X6Y3_LUT4AB/E6END[5] Tile_X6Y3_LUT4AB/E6END[6] Tile_X6Y3_LUT4AB/E6END[7] Tile_X6Y3_LUT4AB/E6END[8]
+ Tile_X6Y3_LUT4AB/E6END[9] Tile_X6Y3_LUT4AB/EE4BEG[0] Tile_X6Y3_LUT4AB/EE4BEG[10]
+ Tile_X6Y3_LUT4AB/EE4BEG[11] Tile_X6Y3_LUT4AB/EE4BEG[12] Tile_X6Y3_LUT4AB/EE4BEG[13]
+ Tile_X6Y3_LUT4AB/EE4BEG[14] Tile_X6Y3_LUT4AB/EE4BEG[15] Tile_X6Y3_LUT4AB/EE4BEG[1]
+ Tile_X6Y3_LUT4AB/EE4BEG[2] Tile_X6Y3_LUT4AB/EE4BEG[3] Tile_X6Y3_LUT4AB/EE4BEG[4]
+ Tile_X6Y3_LUT4AB/EE4BEG[5] Tile_X6Y3_LUT4AB/EE4BEG[6] Tile_X6Y3_LUT4AB/EE4BEG[7]
+ Tile_X6Y3_LUT4AB/EE4BEG[8] Tile_X6Y3_LUT4AB/EE4BEG[9] Tile_X6Y3_LUT4AB/EE4END[0]
+ Tile_X6Y3_LUT4AB/EE4END[10] Tile_X6Y3_LUT4AB/EE4END[11] Tile_X6Y3_LUT4AB/EE4END[12]
+ Tile_X6Y3_LUT4AB/EE4END[13] Tile_X6Y3_LUT4AB/EE4END[14] Tile_X6Y3_LUT4AB/EE4END[15]
+ Tile_X6Y3_LUT4AB/EE4END[1] Tile_X6Y3_LUT4AB/EE4END[2] Tile_X6Y3_LUT4AB/EE4END[3]
+ Tile_X6Y3_LUT4AB/EE4END[4] Tile_X6Y3_LUT4AB/EE4END[5] Tile_X6Y3_LUT4AB/EE4END[6]
+ Tile_X6Y3_LUT4AB/EE4END[7] Tile_X6Y3_LUT4AB/EE4END[8] Tile_X6Y3_LUT4AB/EE4END[9]
+ Tile_X6Y3_LUT4AB/FrameData[0] Tile_X6Y3_LUT4AB/FrameData[10] Tile_X6Y3_LUT4AB/FrameData[11]
+ Tile_X6Y3_LUT4AB/FrameData[12] Tile_X6Y3_LUT4AB/FrameData[13] Tile_X6Y3_LUT4AB/FrameData[14]
+ Tile_X6Y3_LUT4AB/FrameData[15] Tile_X6Y3_LUT4AB/FrameData[16] Tile_X6Y3_LUT4AB/FrameData[17]
+ Tile_X6Y3_LUT4AB/FrameData[18] Tile_X6Y3_LUT4AB/FrameData[19] Tile_X6Y3_LUT4AB/FrameData[1]
+ Tile_X6Y3_LUT4AB/FrameData[20] Tile_X6Y3_LUT4AB/FrameData[21] Tile_X6Y3_LUT4AB/FrameData[22]
+ Tile_X6Y3_LUT4AB/FrameData[23] Tile_X6Y3_LUT4AB/FrameData[24] Tile_X6Y3_LUT4AB/FrameData[25]
+ Tile_X6Y3_LUT4AB/FrameData[26] Tile_X6Y3_LUT4AB/FrameData[27] Tile_X6Y3_LUT4AB/FrameData[28]
+ Tile_X6Y3_LUT4AB/FrameData[29] Tile_X6Y3_LUT4AB/FrameData[2] Tile_X6Y3_LUT4AB/FrameData[30]
+ Tile_X6Y3_LUT4AB/FrameData[31] Tile_X6Y3_LUT4AB/FrameData[3] Tile_X6Y3_LUT4AB/FrameData[4]
+ Tile_X6Y3_LUT4AB/FrameData[5] Tile_X6Y3_LUT4AB/FrameData[6] Tile_X6Y3_LUT4AB/FrameData[7]
+ Tile_X6Y3_LUT4AB/FrameData[8] Tile_X6Y3_LUT4AB/FrameData[9] Tile_X6Y3_LUT4AB/FrameData_O[0]
+ Tile_X6Y3_LUT4AB/FrameData_O[10] Tile_X6Y3_LUT4AB/FrameData_O[11] Tile_X6Y3_LUT4AB/FrameData_O[12]
+ Tile_X6Y3_LUT4AB/FrameData_O[13] Tile_X6Y3_LUT4AB/FrameData_O[14] Tile_X6Y3_LUT4AB/FrameData_O[15]
+ Tile_X6Y3_LUT4AB/FrameData_O[16] Tile_X6Y3_LUT4AB/FrameData_O[17] Tile_X6Y3_LUT4AB/FrameData_O[18]
+ Tile_X6Y3_LUT4AB/FrameData_O[19] Tile_X6Y3_LUT4AB/FrameData_O[1] Tile_X6Y3_LUT4AB/FrameData_O[20]
+ Tile_X6Y3_LUT4AB/FrameData_O[21] Tile_X6Y3_LUT4AB/FrameData_O[22] Tile_X6Y3_LUT4AB/FrameData_O[23]
+ Tile_X6Y3_LUT4AB/FrameData_O[24] Tile_X6Y3_LUT4AB/FrameData_O[25] Tile_X6Y3_LUT4AB/FrameData_O[26]
+ Tile_X6Y3_LUT4AB/FrameData_O[27] Tile_X6Y3_LUT4AB/FrameData_O[28] Tile_X6Y3_LUT4AB/FrameData_O[29]
+ Tile_X6Y3_LUT4AB/FrameData_O[2] Tile_X6Y3_LUT4AB/FrameData_O[30] Tile_X6Y3_LUT4AB/FrameData_O[31]
+ Tile_X6Y3_LUT4AB/FrameData_O[3] Tile_X6Y3_LUT4AB/FrameData_O[4] Tile_X6Y3_LUT4AB/FrameData_O[5]
+ Tile_X6Y3_LUT4AB/FrameData_O[6] Tile_X6Y3_LUT4AB/FrameData_O[7] Tile_X6Y3_LUT4AB/FrameData_O[8]
+ Tile_X6Y3_LUT4AB/FrameData_O[9] Tile_X6Y3_LUT4AB/FrameStrobe[0] Tile_X6Y3_LUT4AB/FrameStrobe[10]
+ Tile_X6Y3_LUT4AB/FrameStrobe[11] Tile_X6Y3_LUT4AB/FrameStrobe[12] Tile_X6Y3_LUT4AB/FrameStrobe[13]
+ Tile_X6Y3_LUT4AB/FrameStrobe[14] Tile_X6Y3_LUT4AB/FrameStrobe[15] Tile_X6Y3_LUT4AB/FrameStrobe[16]
+ Tile_X6Y3_LUT4AB/FrameStrobe[17] Tile_X6Y3_LUT4AB/FrameStrobe[18] Tile_X6Y3_LUT4AB/FrameStrobe[19]
+ Tile_X6Y3_LUT4AB/FrameStrobe[1] Tile_X6Y3_LUT4AB/FrameStrobe[2] Tile_X6Y3_LUT4AB/FrameStrobe[3]
+ Tile_X6Y3_LUT4AB/FrameStrobe[4] Tile_X6Y3_LUT4AB/FrameStrobe[5] Tile_X6Y3_LUT4AB/FrameStrobe[6]
+ Tile_X6Y3_LUT4AB/FrameStrobe[7] Tile_X6Y3_LUT4AB/FrameStrobe[8] Tile_X6Y3_LUT4AB/FrameStrobe[9]
+ Tile_X6Y2_LUT4AB/FrameStrobe[0] Tile_X6Y2_LUT4AB/FrameStrobe[10] Tile_X6Y2_LUT4AB/FrameStrobe[11]
+ Tile_X6Y2_LUT4AB/FrameStrobe[12] Tile_X6Y2_LUT4AB/FrameStrobe[13] Tile_X6Y2_LUT4AB/FrameStrobe[14]
+ Tile_X6Y2_LUT4AB/FrameStrobe[15] Tile_X6Y2_LUT4AB/FrameStrobe[16] Tile_X6Y2_LUT4AB/FrameStrobe[17]
+ Tile_X6Y2_LUT4AB/FrameStrobe[18] Tile_X6Y2_LUT4AB/FrameStrobe[19] Tile_X6Y2_LUT4AB/FrameStrobe[1]
+ Tile_X6Y2_LUT4AB/FrameStrobe[2] Tile_X6Y2_LUT4AB/FrameStrobe[3] Tile_X6Y2_LUT4AB/FrameStrobe[4]
+ Tile_X6Y2_LUT4AB/FrameStrobe[5] Tile_X6Y2_LUT4AB/FrameStrobe[6] Tile_X6Y2_LUT4AB/FrameStrobe[7]
+ Tile_X6Y2_LUT4AB/FrameStrobe[8] Tile_X6Y2_LUT4AB/FrameStrobe[9] Tile_X6Y3_LUT4AB/N1BEG[0]
+ Tile_X6Y3_LUT4AB/N1BEG[1] Tile_X6Y3_LUT4AB/N1BEG[2] Tile_X6Y3_LUT4AB/N1BEG[3] Tile_X6Y4_LUT4AB/N1BEG[0]
+ Tile_X6Y4_LUT4AB/N1BEG[1] Tile_X6Y4_LUT4AB/N1BEG[2] Tile_X6Y4_LUT4AB/N1BEG[3] Tile_X6Y3_LUT4AB/N2BEG[0]
+ Tile_X6Y3_LUT4AB/N2BEG[1] Tile_X6Y3_LUT4AB/N2BEG[2] Tile_X6Y3_LUT4AB/N2BEG[3] Tile_X6Y3_LUT4AB/N2BEG[4]
+ Tile_X6Y3_LUT4AB/N2BEG[5] Tile_X6Y3_LUT4AB/N2BEG[6] Tile_X6Y3_LUT4AB/N2BEG[7] Tile_X6Y2_LUT4AB/N2END[0]
+ Tile_X6Y2_LUT4AB/N2END[1] Tile_X6Y2_LUT4AB/N2END[2] Tile_X6Y2_LUT4AB/N2END[3] Tile_X6Y2_LUT4AB/N2END[4]
+ Tile_X6Y2_LUT4AB/N2END[5] Tile_X6Y2_LUT4AB/N2END[6] Tile_X6Y2_LUT4AB/N2END[7] Tile_X6Y3_LUT4AB/N2END[0]
+ Tile_X6Y3_LUT4AB/N2END[1] Tile_X6Y3_LUT4AB/N2END[2] Tile_X6Y3_LUT4AB/N2END[3] Tile_X6Y3_LUT4AB/N2END[4]
+ Tile_X6Y3_LUT4AB/N2END[5] Tile_X6Y3_LUT4AB/N2END[6] Tile_X6Y3_LUT4AB/N2END[7] Tile_X6Y4_LUT4AB/N2BEG[0]
+ Tile_X6Y4_LUT4AB/N2BEG[1] Tile_X6Y4_LUT4AB/N2BEG[2] Tile_X6Y4_LUT4AB/N2BEG[3] Tile_X6Y4_LUT4AB/N2BEG[4]
+ Tile_X6Y4_LUT4AB/N2BEG[5] Tile_X6Y4_LUT4AB/N2BEG[6] Tile_X6Y4_LUT4AB/N2BEG[7] Tile_X6Y3_LUT4AB/N4BEG[0]
+ Tile_X6Y3_LUT4AB/N4BEG[10] Tile_X6Y3_LUT4AB/N4BEG[11] Tile_X6Y3_LUT4AB/N4BEG[12]
+ Tile_X6Y3_LUT4AB/N4BEG[13] Tile_X6Y3_LUT4AB/N4BEG[14] Tile_X6Y3_LUT4AB/N4BEG[15]
+ Tile_X6Y3_LUT4AB/N4BEG[1] Tile_X6Y3_LUT4AB/N4BEG[2] Tile_X6Y3_LUT4AB/N4BEG[3] Tile_X6Y3_LUT4AB/N4BEG[4]
+ Tile_X6Y3_LUT4AB/N4BEG[5] Tile_X6Y3_LUT4AB/N4BEG[6] Tile_X6Y3_LUT4AB/N4BEG[7] Tile_X6Y3_LUT4AB/N4BEG[8]
+ Tile_X6Y3_LUT4AB/N4BEG[9] Tile_X6Y4_LUT4AB/N4BEG[0] Tile_X6Y4_LUT4AB/N4BEG[10] Tile_X6Y4_LUT4AB/N4BEG[11]
+ Tile_X6Y4_LUT4AB/N4BEG[12] Tile_X6Y4_LUT4AB/N4BEG[13] Tile_X6Y4_LUT4AB/N4BEG[14]
+ Tile_X6Y4_LUT4AB/N4BEG[15] Tile_X6Y4_LUT4AB/N4BEG[1] Tile_X6Y4_LUT4AB/N4BEG[2] Tile_X6Y4_LUT4AB/N4BEG[3]
+ Tile_X6Y4_LUT4AB/N4BEG[4] Tile_X6Y4_LUT4AB/N4BEG[5] Tile_X6Y4_LUT4AB/N4BEG[6] Tile_X6Y4_LUT4AB/N4BEG[7]
+ Tile_X6Y4_LUT4AB/N4BEG[8] Tile_X6Y4_LUT4AB/N4BEG[9] Tile_X6Y3_LUT4AB/NN4BEG[0] Tile_X6Y3_LUT4AB/NN4BEG[10]
+ Tile_X6Y3_LUT4AB/NN4BEG[11] Tile_X6Y3_LUT4AB/NN4BEG[12] Tile_X6Y3_LUT4AB/NN4BEG[13]
+ Tile_X6Y3_LUT4AB/NN4BEG[14] Tile_X6Y3_LUT4AB/NN4BEG[15] Tile_X6Y3_LUT4AB/NN4BEG[1]
+ Tile_X6Y3_LUT4AB/NN4BEG[2] Tile_X6Y3_LUT4AB/NN4BEG[3] Tile_X6Y3_LUT4AB/NN4BEG[4]
+ Tile_X6Y3_LUT4AB/NN4BEG[5] Tile_X6Y3_LUT4AB/NN4BEG[6] Tile_X6Y3_LUT4AB/NN4BEG[7]
+ Tile_X6Y3_LUT4AB/NN4BEG[8] Tile_X6Y3_LUT4AB/NN4BEG[9] Tile_X6Y4_LUT4AB/NN4BEG[0]
+ Tile_X6Y4_LUT4AB/NN4BEG[10] Tile_X6Y4_LUT4AB/NN4BEG[11] Tile_X6Y4_LUT4AB/NN4BEG[12]
+ Tile_X6Y4_LUT4AB/NN4BEG[13] Tile_X6Y4_LUT4AB/NN4BEG[14] Tile_X6Y4_LUT4AB/NN4BEG[15]
+ Tile_X6Y4_LUT4AB/NN4BEG[1] Tile_X6Y4_LUT4AB/NN4BEG[2] Tile_X6Y4_LUT4AB/NN4BEG[3]
+ Tile_X6Y4_LUT4AB/NN4BEG[4] Tile_X6Y4_LUT4AB/NN4BEG[5] Tile_X6Y4_LUT4AB/NN4BEG[6]
+ Tile_X6Y4_LUT4AB/NN4BEG[7] Tile_X6Y4_LUT4AB/NN4BEG[8] Tile_X6Y4_LUT4AB/NN4BEG[9]
+ Tile_X6Y4_LUT4AB/S1END[0] Tile_X6Y4_LUT4AB/S1END[1] Tile_X6Y4_LUT4AB/S1END[2] Tile_X6Y4_LUT4AB/S1END[3]
+ Tile_X6Y3_LUT4AB/S1END[0] Tile_X6Y3_LUT4AB/S1END[1] Tile_X6Y3_LUT4AB/S1END[2] Tile_X6Y3_LUT4AB/S1END[3]
+ Tile_X6Y4_LUT4AB/S2MID[0] Tile_X6Y4_LUT4AB/S2MID[1] Tile_X6Y4_LUT4AB/S2MID[2] Tile_X6Y4_LUT4AB/S2MID[3]
+ Tile_X6Y4_LUT4AB/S2MID[4] Tile_X6Y4_LUT4AB/S2MID[5] Tile_X6Y4_LUT4AB/S2MID[6] Tile_X6Y4_LUT4AB/S2MID[7]
+ Tile_X6Y4_LUT4AB/S2END[0] Tile_X6Y4_LUT4AB/S2END[1] Tile_X6Y4_LUT4AB/S2END[2] Tile_X6Y4_LUT4AB/S2END[3]
+ Tile_X6Y4_LUT4AB/S2END[4] Tile_X6Y4_LUT4AB/S2END[5] Tile_X6Y4_LUT4AB/S2END[6] Tile_X6Y4_LUT4AB/S2END[7]
+ Tile_X6Y3_LUT4AB/S2END[0] Tile_X6Y3_LUT4AB/S2END[1] Tile_X6Y3_LUT4AB/S2END[2] Tile_X6Y3_LUT4AB/S2END[3]
+ Tile_X6Y3_LUT4AB/S2END[4] Tile_X6Y3_LUT4AB/S2END[5] Tile_X6Y3_LUT4AB/S2END[6] Tile_X6Y3_LUT4AB/S2END[7]
+ Tile_X6Y3_LUT4AB/S2MID[0] Tile_X6Y3_LUT4AB/S2MID[1] Tile_X6Y3_LUT4AB/S2MID[2] Tile_X6Y3_LUT4AB/S2MID[3]
+ Tile_X6Y3_LUT4AB/S2MID[4] Tile_X6Y3_LUT4AB/S2MID[5] Tile_X6Y3_LUT4AB/S2MID[6] Tile_X6Y3_LUT4AB/S2MID[7]
+ Tile_X6Y4_LUT4AB/S4END[0] Tile_X6Y4_LUT4AB/S4END[10] Tile_X6Y4_LUT4AB/S4END[11]
+ Tile_X6Y4_LUT4AB/S4END[12] Tile_X6Y4_LUT4AB/S4END[13] Tile_X6Y4_LUT4AB/S4END[14]
+ Tile_X6Y4_LUT4AB/S4END[15] Tile_X6Y4_LUT4AB/S4END[1] Tile_X6Y4_LUT4AB/S4END[2] Tile_X6Y4_LUT4AB/S4END[3]
+ Tile_X6Y4_LUT4AB/S4END[4] Tile_X6Y4_LUT4AB/S4END[5] Tile_X6Y4_LUT4AB/S4END[6] Tile_X6Y4_LUT4AB/S4END[7]
+ Tile_X6Y4_LUT4AB/S4END[8] Tile_X6Y4_LUT4AB/S4END[9] Tile_X6Y3_LUT4AB/S4END[0] Tile_X6Y3_LUT4AB/S4END[10]
+ Tile_X6Y3_LUT4AB/S4END[11] Tile_X6Y3_LUT4AB/S4END[12] Tile_X6Y3_LUT4AB/S4END[13]
+ Tile_X6Y3_LUT4AB/S4END[14] Tile_X6Y3_LUT4AB/S4END[15] Tile_X6Y3_LUT4AB/S4END[1]
+ Tile_X6Y3_LUT4AB/S4END[2] Tile_X6Y3_LUT4AB/S4END[3] Tile_X6Y3_LUT4AB/S4END[4] Tile_X6Y3_LUT4AB/S4END[5]
+ Tile_X6Y3_LUT4AB/S4END[6] Tile_X6Y3_LUT4AB/S4END[7] Tile_X6Y3_LUT4AB/S4END[8] Tile_X6Y3_LUT4AB/S4END[9]
+ Tile_X6Y4_LUT4AB/SS4END[0] Tile_X6Y4_LUT4AB/SS4END[10] Tile_X6Y4_LUT4AB/SS4END[11]
+ Tile_X6Y4_LUT4AB/SS4END[12] Tile_X6Y4_LUT4AB/SS4END[13] Tile_X6Y4_LUT4AB/SS4END[14]
+ Tile_X6Y4_LUT4AB/SS4END[15] Tile_X6Y4_LUT4AB/SS4END[1] Tile_X6Y4_LUT4AB/SS4END[2]
+ Tile_X6Y4_LUT4AB/SS4END[3] Tile_X6Y4_LUT4AB/SS4END[4] Tile_X6Y4_LUT4AB/SS4END[5]
+ Tile_X6Y4_LUT4AB/SS4END[6] Tile_X6Y4_LUT4AB/SS4END[7] Tile_X6Y4_LUT4AB/SS4END[8]
+ Tile_X6Y4_LUT4AB/SS4END[9] Tile_X6Y3_LUT4AB/SS4END[0] Tile_X6Y3_LUT4AB/SS4END[10]
+ Tile_X6Y3_LUT4AB/SS4END[11] Tile_X6Y3_LUT4AB/SS4END[12] Tile_X6Y3_LUT4AB/SS4END[13]
+ Tile_X6Y3_LUT4AB/SS4END[14] Tile_X6Y3_LUT4AB/SS4END[15] Tile_X6Y3_LUT4AB/SS4END[1]
+ Tile_X6Y3_LUT4AB/SS4END[2] Tile_X6Y3_LUT4AB/SS4END[3] Tile_X6Y3_LUT4AB/SS4END[4]
+ Tile_X6Y3_LUT4AB/SS4END[5] Tile_X6Y3_LUT4AB/SS4END[6] Tile_X6Y3_LUT4AB/SS4END[7]
+ Tile_X6Y3_LUT4AB/SS4END[8] Tile_X6Y3_LUT4AB/SS4END[9] Tile_X6Y3_LUT4AB/UserCLK Tile_X6Y2_LUT4AB/UserCLK
+ VGND VPWR Tile_X6Y3_LUT4AB/W1BEG[0] Tile_X6Y3_LUT4AB/W1BEG[1] Tile_X6Y3_LUT4AB/W1BEG[2]
+ Tile_X6Y3_LUT4AB/W1BEG[3] Tile_X6Y3_LUT4AB/W1END[0] Tile_X6Y3_LUT4AB/W1END[1] Tile_X6Y3_LUT4AB/W1END[2]
+ Tile_X6Y3_LUT4AB/W1END[3] Tile_X6Y3_LUT4AB/W2BEG[0] Tile_X6Y3_LUT4AB/W2BEG[1] Tile_X6Y3_LUT4AB/W2BEG[2]
+ Tile_X6Y3_LUT4AB/W2BEG[3] Tile_X6Y3_LUT4AB/W2BEG[4] Tile_X6Y3_LUT4AB/W2BEG[5] Tile_X6Y3_LUT4AB/W2BEG[6]
+ Tile_X6Y3_LUT4AB/W2BEG[7] Tile_X5Y3_LUT4AB/W2END[0] Tile_X5Y3_LUT4AB/W2END[1] Tile_X5Y3_LUT4AB/W2END[2]
+ Tile_X5Y3_LUT4AB/W2END[3] Tile_X5Y3_LUT4AB/W2END[4] Tile_X5Y3_LUT4AB/W2END[5] Tile_X5Y3_LUT4AB/W2END[6]
+ Tile_X5Y3_LUT4AB/W2END[7] Tile_X6Y3_LUT4AB/W2END[0] Tile_X6Y3_LUT4AB/W2END[1] Tile_X6Y3_LUT4AB/W2END[2]
+ Tile_X6Y3_LUT4AB/W2END[3] Tile_X6Y3_LUT4AB/W2END[4] Tile_X6Y3_LUT4AB/W2END[5] Tile_X6Y3_LUT4AB/W2END[6]
+ Tile_X6Y3_LUT4AB/W2END[7] Tile_X6Y3_LUT4AB/W2MID[0] Tile_X6Y3_LUT4AB/W2MID[1] Tile_X6Y3_LUT4AB/W2MID[2]
+ Tile_X6Y3_LUT4AB/W2MID[3] Tile_X6Y3_LUT4AB/W2MID[4] Tile_X6Y3_LUT4AB/W2MID[5] Tile_X6Y3_LUT4AB/W2MID[6]
+ Tile_X6Y3_LUT4AB/W2MID[7] Tile_X6Y3_LUT4AB/W6BEG[0] Tile_X6Y3_LUT4AB/W6BEG[10] Tile_X6Y3_LUT4AB/W6BEG[11]
+ Tile_X6Y3_LUT4AB/W6BEG[1] Tile_X6Y3_LUT4AB/W6BEG[2] Tile_X6Y3_LUT4AB/W6BEG[3] Tile_X6Y3_LUT4AB/W6BEG[4]
+ Tile_X6Y3_LUT4AB/W6BEG[5] Tile_X6Y3_LUT4AB/W6BEG[6] Tile_X6Y3_LUT4AB/W6BEG[7] Tile_X6Y3_LUT4AB/W6BEG[8]
+ Tile_X6Y3_LUT4AB/W6BEG[9] Tile_X6Y3_LUT4AB/W6END[0] Tile_X6Y3_LUT4AB/W6END[10] Tile_X6Y3_LUT4AB/W6END[11]
+ Tile_X6Y3_LUT4AB/W6END[1] Tile_X6Y3_LUT4AB/W6END[2] Tile_X6Y3_LUT4AB/W6END[3] Tile_X6Y3_LUT4AB/W6END[4]
+ Tile_X6Y3_LUT4AB/W6END[5] Tile_X6Y3_LUT4AB/W6END[6] Tile_X6Y3_LUT4AB/W6END[7] Tile_X6Y3_LUT4AB/W6END[8]
+ Tile_X6Y3_LUT4AB/W6END[9] Tile_X6Y3_LUT4AB/WW4BEG[0] Tile_X6Y3_LUT4AB/WW4BEG[10]
+ Tile_X6Y3_LUT4AB/WW4BEG[11] Tile_X6Y3_LUT4AB/WW4BEG[12] Tile_X6Y3_LUT4AB/WW4BEG[13]
+ Tile_X6Y3_LUT4AB/WW4BEG[14] Tile_X6Y3_LUT4AB/WW4BEG[15] Tile_X6Y3_LUT4AB/WW4BEG[1]
+ Tile_X6Y3_LUT4AB/WW4BEG[2] Tile_X6Y3_LUT4AB/WW4BEG[3] Tile_X6Y3_LUT4AB/WW4BEG[4]
+ Tile_X6Y3_LUT4AB/WW4BEG[5] Tile_X6Y3_LUT4AB/WW4BEG[6] Tile_X6Y3_LUT4AB/WW4BEG[7]
+ Tile_X6Y3_LUT4AB/WW4BEG[8] Tile_X6Y3_LUT4AB/WW4BEG[9] Tile_X6Y3_LUT4AB/WW4END[0]
+ Tile_X6Y3_LUT4AB/WW4END[10] Tile_X6Y3_LUT4AB/WW4END[11] Tile_X6Y3_LUT4AB/WW4END[12]
+ Tile_X6Y3_LUT4AB/WW4END[13] Tile_X6Y3_LUT4AB/WW4END[14] Tile_X6Y3_LUT4AB/WW4END[15]
+ Tile_X6Y3_LUT4AB/WW4END[1] Tile_X6Y3_LUT4AB/WW4END[2] Tile_X6Y3_LUT4AB/WW4END[3]
+ Tile_X6Y3_LUT4AB/WW4END[4] Tile_X6Y3_LUT4AB/WW4END[5] Tile_X6Y3_LUT4AB/WW4END[6]
+ Tile_X6Y3_LUT4AB/WW4END[7] Tile_X6Y3_LUT4AB/WW4END[8] Tile_X6Y3_LUT4AB/WW4END[9]
+ LUT4AB
XTile_X0Y9_W_IO Tile_X0Y9_A_I_top Tile_X0Y9_A_O_top Tile_X0Y9_A_T_top Tile_X0Y9_A_config_C_bit0
+ Tile_X0Y9_A_config_C_bit1 Tile_X0Y9_A_config_C_bit2 Tile_X0Y9_A_config_C_bit3 Tile_X0Y9_B_I_top
+ Tile_X0Y9_B_O_top Tile_X0Y9_B_T_top Tile_X0Y9_B_config_C_bit0 Tile_X0Y9_B_config_C_bit1
+ Tile_X0Y9_B_config_C_bit2 Tile_X0Y9_B_config_C_bit3 Tile_X0Y9_W_IO/E1BEG[0] Tile_X0Y9_W_IO/E1BEG[1]
+ Tile_X0Y9_W_IO/E1BEG[2] Tile_X0Y9_W_IO/E1BEG[3] Tile_X0Y9_W_IO/E2BEG[0] Tile_X0Y9_W_IO/E2BEG[1]
+ Tile_X0Y9_W_IO/E2BEG[2] Tile_X0Y9_W_IO/E2BEG[3] Tile_X0Y9_W_IO/E2BEG[4] Tile_X0Y9_W_IO/E2BEG[5]
+ Tile_X0Y9_W_IO/E2BEG[6] Tile_X0Y9_W_IO/E2BEG[7] Tile_X0Y9_W_IO/E2BEGb[0] Tile_X0Y9_W_IO/E2BEGb[1]
+ Tile_X0Y9_W_IO/E2BEGb[2] Tile_X0Y9_W_IO/E2BEGb[3] Tile_X0Y9_W_IO/E2BEGb[4] Tile_X0Y9_W_IO/E2BEGb[5]
+ Tile_X0Y9_W_IO/E2BEGb[6] Tile_X0Y9_W_IO/E2BEGb[7] Tile_X0Y9_W_IO/E6BEG[0] Tile_X0Y9_W_IO/E6BEG[10]
+ Tile_X0Y9_W_IO/E6BEG[11] Tile_X0Y9_W_IO/E6BEG[1] Tile_X0Y9_W_IO/E6BEG[2] Tile_X0Y9_W_IO/E6BEG[3]
+ Tile_X0Y9_W_IO/E6BEG[4] Tile_X0Y9_W_IO/E6BEG[5] Tile_X0Y9_W_IO/E6BEG[6] Tile_X0Y9_W_IO/E6BEG[7]
+ Tile_X0Y9_W_IO/E6BEG[8] Tile_X0Y9_W_IO/E6BEG[9] Tile_X0Y9_W_IO/EE4BEG[0] Tile_X0Y9_W_IO/EE4BEG[10]
+ Tile_X0Y9_W_IO/EE4BEG[11] Tile_X0Y9_W_IO/EE4BEG[12] Tile_X0Y9_W_IO/EE4BEG[13] Tile_X0Y9_W_IO/EE4BEG[14]
+ Tile_X0Y9_W_IO/EE4BEG[15] Tile_X0Y9_W_IO/EE4BEG[1] Tile_X0Y9_W_IO/EE4BEG[2] Tile_X0Y9_W_IO/EE4BEG[3]
+ Tile_X0Y9_W_IO/EE4BEG[4] Tile_X0Y9_W_IO/EE4BEG[5] Tile_X0Y9_W_IO/EE4BEG[6] Tile_X0Y9_W_IO/EE4BEG[7]
+ Tile_X0Y9_W_IO/EE4BEG[8] Tile_X0Y9_W_IO/EE4BEG[9] FrameData[288] FrameData[298]
+ FrameData[299] FrameData[300] FrameData[301] FrameData[302] FrameData[303] FrameData[304]
+ FrameData[305] FrameData[306] FrameData[307] FrameData[289] FrameData[308] FrameData[309]
+ FrameData[310] FrameData[311] FrameData[312] FrameData[313] FrameData[314] FrameData[315]
+ FrameData[316] FrameData[317] FrameData[290] FrameData[318] FrameData[319] FrameData[291]
+ FrameData[292] FrameData[293] FrameData[294] FrameData[295] FrameData[296] FrameData[297]
+ Tile_X1Y9_LUT4AB/FrameData[0] Tile_X1Y9_LUT4AB/FrameData[10] Tile_X1Y9_LUT4AB/FrameData[11]
+ Tile_X1Y9_LUT4AB/FrameData[12] Tile_X1Y9_LUT4AB/FrameData[13] Tile_X1Y9_LUT4AB/FrameData[14]
+ Tile_X1Y9_LUT4AB/FrameData[15] Tile_X1Y9_LUT4AB/FrameData[16] Tile_X1Y9_LUT4AB/FrameData[17]
+ Tile_X1Y9_LUT4AB/FrameData[18] Tile_X1Y9_LUT4AB/FrameData[19] Tile_X1Y9_LUT4AB/FrameData[1]
+ Tile_X1Y9_LUT4AB/FrameData[20] Tile_X1Y9_LUT4AB/FrameData[21] Tile_X1Y9_LUT4AB/FrameData[22]
+ Tile_X1Y9_LUT4AB/FrameData[23] Tile_X1Y9_LUT4AB/FrameData[24] Tile_X1Y9_LUT4AB/FrameData[25]
+ Tile_X1Y9_LUT4AB/FrameData[26] Tile_X1Y9_LUT4AB/FrameData[27] Tile_X1Y9_LUT4AB/FrameData[28]
+ Tile_X1Y9_LUT4AB/FrameData[29] Tile_X1Y9_LUT4AB/FrameData[2] Tile_X1Y9_LUT4AB/FrameData[30]
+ Tile_X1Y9_LUT4AB/FrameData[31] Tile_X1Y9_LUT4AB/FrameData[3] Tile_X1Y9_LUT4AB/FrameData[4]
+ Tile_X1Y9_LUT4AB/FrameData[5] Tile_X1Y9_LUT4AB/FrameData[6] Tile_X1Y9_LUT4AB/FrameData[7]
+ Tile_X1Y9_LUT4AB/FrameData[8] Tile_X1Y9_LUT4AB/FrameData[9] Tile_X0Y9_W_IO/FrameStrobe[0]
+ Tile_X0Y9_W_IO/FrameStrobe[10] Tile_X0Y9_W_IO/FrameStrobe[11] Tile_X0Y9_W_IO/FrameStrobe[12]
+ Tile_X0Y9_W_IO/FrameStrobe[13] Tile_X0Y9_W_IO/FrameStrobe[14] Tile_X0Y9_W_IO/FrameStrobe[15]
+ Tile_X0Y9_W_IO/FrameStrobe[16] Tile_X0Y9_W_IO/FrameStrobe[17] Tile_X0Y9_W_IO/FrameStrobe[18]
+ Tile_X0Y9_W_IO/FrameStrobe[19] Tile_X0Y9_W_IO/FrameStrobe[1] Tile_X0Y9_W_IO/FrameStrobe[2]
+ Tile_X0Y9_W_IO/FrameStrobe[3] Tile_X0Y9_W_IO/FrameStrobe[4] Tile_X0Y9_W_IO/FrameStrobe[5]
+ Tile_X0Y9_W_IO/FrameStrobe[6] Tile_X0Y9_W_IO/FrameStrobe[7] Tile_X0Y9_W_IO/FrameStrobe[8]
+ Tile_X0Y9_W_IO/FrameStrobe[9] Tile_X0Y8_W_IO/FrameStrobe[0] Tile_X0Y8_W_IO/FrameStrobe[10]
+ Tile_X0Y8_W_IO/FrameStrobe[11] Tile_X0Y8_W_IO/FrameStrobe[12] Tile_X0Y8_W_IO/FrameStrobe[13]
+ Tile_X0Y8_W_IO/FrameStrobe[14] Tile_X0Y8_W_IO/FrameStrobe[15] Tile_X0Y8_W_IO/FrameStrobe[16]
+ Tile_X0Y8_W_IO/FrameStrobe[17] Tile_X0Y8_W_IO/FrameStrobe[18] Tile_X0Y8_W_IO/FrameStrobe[19]
+ Tile_X0Y8_W_IO/FrameStrobe[1] Tile_X0Y8_W_IO/FrameStrobe[2] Tile_X0Y8_W_IO/FrameStrobe[3]
+ Tile_X0Y8_W_IO/FrameStrobe[4] Tile_X0Y8_W_IO/FrameStrobe[5] Tile_X0Y8_W_IO/FrameStrobe[6]
+ Tile_X0Y8_W_IO/FrameStrobe[7] Tile_X0Y8_W_IO/FrameStrobe[8] Tile_X0Y8_W_IO/FrameStrobe[9]
+ Tile_X0Y9_W_IO/UserCLK Tile_X0Y8_W_IO/UserCLK VGND VPWR Tile_X0Y9_W_IO/W1END[0]
+ Tile_X0Y9_W_IO/W1END[1] Tile_X0Y9_W_IO/W1END[2] Tile_X0Y9_W_IO/W1END[3] Tile_X0Y9_W_IO/W2END[0]
+ Tile_X0Y9_W_IO/W2END[1] Tile_X0Y9_W_IO/W2END[2] Tile_X0Y9_W_IO/W2END[3] Tile_X0Y9_W_IO/W2END[4]
+ Tile_X0Y9_W_IO/W2END[5] Tile_X0Y9_W_IO/W2END[6] Tile_X0Y9_W_IO/W2END[7] Tile_X0Y9_W_IO/W2MID[0]
+ Tile_X0Y9_W_IO/W2MID[1] Tile_X0Y9_W_IO/W2MID[2] Tile_X0Y9_W_IO/W2MID[3] Tile_X0Y9_W_IO/W2MID[4]
+ Tile_X0Y9_W_IO/W2MID[5] Tile_X0Y9_W_IO/W2MID[6] Tile_X0Y9_W_IO/W2MID[7] Tile_X0Y9_W_IO/W6END[0]
+ Tile_X0Y9_W_IO/W6END[10] Tile_X0Y9_W_IO/W6END[11] Tile_X0Y9_W_IO/W6END[1] Tile_X0Y9_W_IO/W6END[2]
+ Tile_X0Y9_W_IO/W6END[3] Tile_X0Y9_W_IO/W6END[4] Tile_X0Y9_W_IO/W6END[5] Tile_X0Y9_W_IO/W6END[6]
+ Tile_X0Y9_W_IO/W6END[7] Tile_X0Y9_W_IO/W6END[8] Tile_X0Y9_W_IO/W6END[9] Tile_X0Y9_W_IO/WW4END[0]
+ Tile_X0Y9_W_IO/WW4END[10] Tile_X0Y9_W_IO/WW4END[11] Tile_X0Y9_W_IO/WW4END[12] Tile_X0Y9_W_IO/WW4END[13]
+ Tile_X0Y9_W_IO/WW4END[14] Tile_X0Y9_W_IO/WW4END[15] Tile_X0Y9_W_IO/WW4END[1] Tile_X0Y9_W_IO/WW4END[2]
+ Tile_X0Y9_W_IO/WW4END[3] Tile_X0Y9_W_IO/WW4END[4] Tile_X0Y9_W_IO/WW4END[5] Tile_X0Y9_W_IO/WW4END[6]
+ Tile_X0Y9_W_IO/WW4END[7] Tile_X0Y9_W_IO/WW4END[8] Tile_X0Y9_W_IO/WW4END[9] W_IO
XTile_X2Y15_S_WARMBOOT Tile_X2Y15_BOOT_top Tile_X2Y15_CONFIGURED_top Tile_X2Y14_LUT4AB/Ci
+ Tile_X2Y15_S_WARMBOOT/FrameData[0] Tile_X2Y15_S_WARMBOOT/FrameData[10] Tile_X2Y15_S_WARMBOOT/FrameData[11]
+ Tile_X2Y15_S_WARMBOOT/FrameData[12] Tile_X2Y15_S_WARMBOOT/FrameData[13] Tile_X2Y15_S_WARMBOOT/FrameData[14]
+ Tile_X2Y15_S_WARMBOOT/FrameData[15] Tile_X2Y15_S_WARMBOOT/FrameData[16] Tile_X2Y15_S_WARMBOOT/FrameData[17]
+ Tile_X2Y15_S_WARMBOOT/FrameData[18] Tile_X2Y15_S_WARMBOOT/FrameData[19] Tile_X2Y15_S_WARMBOOT/FrameData[1]
+ Tile_X2Y15_S_WARMBOOT/FrameData[20] Tile_X2Y15_S_WARMBOOT/FrameData[21] Tile_X2Y15_S_WARMBOOT/FrameData[22]
+ Tile_X2Y15_S_WARMBOOT/FrameData[23] Tile_X2Y15_S_WARMBOOT/FrameData[24] Tile_X2Y15_S_WARMBOOT/FrameData[25]
+ Tile_X2Y15_S_WARMBOOT/FrameData[26] Tile_X2Y15_S_WARMBOOT/FrameData[27] Tile_X2Y15_S_WARMBOOT/FrameData[28]
+ Tile_X2Y15_S_WARMBOOT/FrameData[29] Tile_X2Y15_S_WARMBOOT/FrameData[2] Tile_X2Y15_S_WARMBOOT/FrameData[30]
+ Tile_X2Y15_S_WARMBOOT/FrameData[31] Tile_X2Y15_S_WARMBOOT/FrameData[3] Tile_X2Y15_S_WARMBOOT/FrameData[4]
+ Tile_X2Y15_S_WARMBOOT/FrameData[5] Tile_X2Y15_S_WARMBOOT/FrameData[6] Tile_X2Y15_S_WARMBOOT/FrameData[7]
+ Tile_X2Y15_S_WARMBOOT/FrameData[8] Tile_X2Y15_S_WARMBOOT/FrameData[9] Tile_X3Y15_S_CPU_IRQ/FrameData[0]
+ Tile_X3Y15_S_CPU_IRQ/FrameData[10] Tile_X3Y15_S_CPU_IRQ/FrameData[11] Tile_X3Y15_S_CPU_IRQ/FrameData[12]
+ Tile_X3Y15_S_CPU_IRQ/FrameData[13] Tile_X3Y15_S_CPU_IRQ/FrameData[14] Tile_X3Y15_S_CPU_IRQ/FrameData[15]
+ Tile_X3Y15_S_CPU_IRQ/FrameData[16] Tile_X3Y15_S_CPU_IRQ/FrameData[17] Tile_X3Y15_S_CPU_IRQ/FrameData[18]
+ Tile_X3Y15_S_CPU_IRQ/FrameData[19] Tile_X3Y15_S_CPU_IRQ/FrameData[1] Tile_X3Y15_S_CPU_IRQ/FrameData[20]
+ Tile_X3Y15_S_CPU_IRQ/FrameData[21] Tile_X3Y15_S_CPU_IRQ/FrameData[22] Tile_X3Y15_S_CPU_IRQ/FrameData[23]
+ Tile_X3Y15_S_CPU_IRQ/FrameData[24] Tile_X3Y15_S_CPU_IRQ/FrameData[25] Tile_X3Y15_S_CPU_IRQ/FrameData[26]
+ Tile_X3Y15_S_CPU_IRQ/FrameData[27] Tile_X3Y15_S_CPU_IRQ/FrameData[28] Tile_X3Y15_S_CPU_IRQ/FrameData[29]
+ Tile_X3Y15_S_CPU_IRQ/FrameData[2] Tile_X3Y15_S_CPU_IRQ/FrameData[30] Tile_X3Y15_S_CPU_IRQ/FrameData[31]
+ Tile_X3Y15_S_CPU_IRQ/FrameData[3] Tile_X3Y15_S_CPU_IRQ/FrameData[4] Tile_X3Y15_S_CPU_IRQ/FrameData[5]
+ Tile_X3Y15_S_CPU_IRQ/FrameData[6] Tile_X3Y15_S_CPU_IRQ/FrameData[7] Tile_X3Y15_S_CPU_IRQ/FrameData[8]
+ Tile_X3Y15_S_CPU_IRQ/FrameData[9] FrameStrobe[40] FrameStrobe[50] FrameStrobe[51]
+ FrameStrobe[52] FrameStrobe[53] FrameStrobe[54] FrameStrobe[55] FrameStrobe[56]
+ FrameStrobe[57] FrameStrobe[58] FrameStrobe[59] FrameStrobe[41] FrameStrobe[42]
+ FrameStrobe[43] FrameStrobe[44] FrameStrobe[45] FrameStrobe[46] FrameStrobe[47]
+ FrameStrobe[48] FrameStrobe[49] Tile_X2Y14_LUT4AB/FrameStrobe[0] Tile_X2Y14_LUT4AB/FrameStrobe[10]
+ Tile_X2Y14_LUT4AB/FrameStrobe[11] Tile_X2Y14_LUT4AB/FrameStrobe[12] Tile_X2Y14_LUT4AB/FrameStrobe[13]
+ Tile_X2Y14_LUT4AB/FrameStrobe[14] Tile_X2Y14_LUT4AB/FrameStrobe[15] Tile_X2Y14_LUT4AB/FrameStrobe[16]
+ Tile_X2Y14_LUT4AB/FrameStrobe[17] Tile_X2Y14_LUT4AB/FrameStrobe[18] Tile_X2Y14_LUT4AB/FrameStrobe[19]
+ Tile_X2Y14_LUT4AB/FrameStrobe[1] Tile_X2Y14_LUT4AB/FrameStrobe[2] Tile_X2Y14_LUT4AB/FrameStrobe[3]
+ Tile_X2Y14_LUT4AB/FrameStrobe[4] Tile_X2Y14_LUT4AB/FrameStrobe[5] Tile_X2Y14_LUT4AB/FrameStrobe[6]
+ Tile_X2Y14_LUT4AB/FrameStrobe[7] Tile_X2Y14_LUT4AB/FrameStrobe[8] Tile_X2Y14_LUT4AB/FrameStrobe[9]
+ Tile_X2Y14_LUT4AB/N1END[0] Tile_X2Y14_LUT4AB/N1END[1] Tile_X2Y14_LUT4AB/N1END[2]
+ Tile_X2Y14_LUT4AB/N1END[3] Tile_X2Y14_LUT4AB/N2MID[0] Tile_X2Y14_LUT4AB/N2MID[1]
+ Tile_X2Y14_LUT4AB/N2MID[2] Tile_X2Y14_LUT4AB/N2MID[3] Tile_X2Y14_LUT4AB/N2MID[4]
+ Tile_X2Y14_LUT4AB/N2MID[5] Tile_X2Y14_LUT4AB/N2MID[6] Tile_X2Y14_LUT4AB/N2MID[7]
+ Tile_X2Y14_LUT4AB/N2END[0] Tile_X2Y14_LUT4AB/N2END[1] Tile_X2Y14_LUT4AB/N2END[2]
+ Tile_X2Y14_LUT4AB/N2END[3] Tile_X2Y14_LUT4AB/N2END[4] Tile_X2Y14_LUT4AB/N2END[5]
+ Tile_X2Y14_LUT4AB/N2END[6] Tile_X2Y14_LUT4AB/N2END[7] Tile_X2Y14_LUT4AB/N4END[0]
+ Tile_X2Y14_LUT4AB/N4END[10] Tile_X2Y14_LUT4AB/N4END[11] Tile_X2Y14_LUT4AB/N4END[12]
+ Tile_X2Y14_LUT4AB/N4END[13] Tile_X2Y14_LUT4AB/N4END[14] Tile_X2Y14_LUT4AB/N4END[15]
+ Tile_X2Y14_LUT4AB/N4END[1] Tile_X2Y14_LUT4AB/N4END[2] Tile_X2Y14_LUT4AB/N4END[3]
+ Tile_X2Y14_LUT4AB/N4END[4] Tile_X2Y14_LUT4AB/N4END[5] Tile_X2Y14_LUT4AB/N4END[6]
+ Tile_X2Y14_LUT4AB/N4END[7] Tile_X2Y14_LUT4AB/N4END[8] Tile_X2Y14_LUT4AB/N4END[9]
+ Tile_X2Y14_LUT4AB/NN4END[0] Tile_X2Y14_LUT4AB/NN4END[10] Tile_X2Y14_LUT4AB/NN4END[11]
+ Tile_X2Y14_LUT4AB/NN4END[12] Tile_X2Y14_LUT4AB/NN4END[13] Tile_X2Y14_LUT4AB/NN4END[14]
+ Tile_X2Y14_LUT4AB/NN4END[15] Tile_X2Y14_LUT4AB/NN4END[1] Tile_X2Y14_LUT4AB/NN4END[2]
+ Tile_X2Y14_LUT4AB/NN4END[3] Tile_X2Y14_LUT4AB/NN4END[4] Tile_X2Y14_LUT4AB/NN4END[5]
+ Tile_X2Y14_LUT4AB/NN4END[6] Tile_X2Y14_LUT4AB/NN4END[7] Tile_X2Y14_LUT4AB/NN4END[8]
+ Tile_X2Y14_LUT4AB/NN4END[9] Tile_X2Y15_RESET_top Tile_X2Y14_LUT4AB/S1BEG[0] Tile_X2Y14_LUT4AB/S1BEG[1]
+ Tile_X2Y14_LUT4AB/S1BEG[2] Tile_X2Y14_LUT4AB/S1BEG[3] Tile_X2Y14_LUT4AB/S2BEGb[0]
+ Tile_X2Y14_LUT4AB/S2BEGb[1] Tile_X2Y14_LUT4AB/S2BEGb[2] Tile_X2Y14_LUT4AB/S2BEGb[3]
+ Tile_X2Y14_LUT4AB/S2BEGb[4] Tile_X2Y14_LUT4AB/S2BEGb[5] Tile_X2Y14_LUT4AB/S2BEGb[6]
+ Tile_X2Y14_LUT4AB/S2BEGb[7] Tile_X2Y14_LUT4AB/S2BEG[0] Tile_X2Y14_LUT4AB/S2BEG[1]
+ Tile_X2Y14_LUT4AB/S2BEG[2] Tile_X2Y14_LUT4AB/S2BEG[3] Tile_X2Y14_LUT4AB/S2BEG[4]
+ Tile_X2Y14_LUT4AB/S2BEG[5] Tile_X2Y14_LUT4AB/S2BEG[6] Tile_X2Y14_LUT4AB/S2BEG[7]
+ Tile_X2Y14_LUT4AB/S4BEG[0] Tile_X2Y14_LUT4AB/S4BEG[10] Tile_X2Y14_LUT4AB/S4BEG[11]
+ Tile_X2Y14_LUT4AB/S4BEG[12] Tile_X2Y14_LUT4AB/S4BEG[13] Tile_X2Y14_LUT4AB/S4BEG[14]
+ Tile_X2Y14_LUT4AB/S4BEG[15] Tile_X2Y14_LUT4AB/S4BEG[1] Tile_X2Y14_LUT4AB/S4BEG[2]
+ Tile_X2Y14_LUT4AB/S4BEG[3] Tile_X2Y14_LUT4AB/S4BEG[4] Tile_X2Y14_LUT4AB/S4BEG[5]
+ Tile_X2Y14_LUT4AB/S4BEG[6] Tile_X2Y14_LUT4AB/S4BEG[7] Tile_X2Y14_LUT4AB/S4BEG[8]
+ Tile_X2Y14_LUT4AB/S4BEG[9] Tile_X2Y15_SLOT_top0 Tile_X2Y15_SLOT_top1 Tile_X2Y15_SLOT_top2
+ Tile_X2Y15_SLOT_top3 Tile_X2Y14_LUT4AB/SS4BEG[0] Tile_X2Y14_LUT4AB/SS4BEG[10] Tile_X2Y14_LUT4AB/SS4BEG[11]
+ Tile_X2Y14_LUT4AB/SS4BEG[12] Tile_X2Y14_LUT4AB/SS4BEG[13] Tile_X2Y14_LUT4AB/SS4BEG[14]
+ Tile_X2Y14_LUT4AB/SS4BEG[15] Tile_X2Y14_LUT4AB/SS4BEG[1] Tile_X2Y14_LUT4AB/SS4BEG[2]
+ Tile_X2Y14_LUT4AB/SS4BEG[3] Tile_X2Y14_LUT4AB/SS4BEG[4] Tile_X2Y14_LUT4AB/SS4BEG[5]
+ Tile_X2Y14_LUT4AB/SS4BEG[6] Tile_X2Y14_LUT4AB/SS4BEG[7] Tile_X2Y14_LUT4AB/SS4BEG[8]
+ Tile_X2Y14_LUT4AB/SS4BEG[9] UserCLK Tile_X2Y14_LUT4AB/UserCLK VGND VPWR S_WARMBOOT
XTile_X8Y12_LUT4AB Tile_X8Y13_LUT4AB/Co Tile_X8Y12_LUT4AB/Co Tile_X9Y12_LUT4AB/E1END[0]
+ Tile_X9Y12_LUT4AB/E1END[1] Tile_X9Y12_LUT4AB/E1END[2] Tile_X9Y12_LUT4AB/E1END[3]
+ Tile_X8Y12_LUT4AB/E1END[0] Tile_X8Y12_LUT4AB/E1END[1] Tile_X8Y12_LUT4AB/E1END[2]
+ Tile_X8Y12_LUT4AB/E1END[3] Tile_X9Y12_LUT4AB/E2MID[0] Tile_X9Y12_LUT4AB/E2MID[1]
+ Tile_X9Y12_LUT4AB/E2MID[2] Tile_X9Y12_LUT4AB/E2MID[3] Tile_X9Y12_LUT4AB/E2MID[4]
+ Tile_X9Y12_LUT4AB/E2MID[5] Tile_X9Y12_LUT4AB/E2MID[6] Tile_X9Y12_LUT4AB/E2MID[7]
+ Tile_X9Y12_LUT4AB/E2END[0] Tile_X9Y12_LUT4AB/E2END[1] Tile_X9Y12_LUT4AB/E2END[2]
+ Tile_X9Y12_LUT4AB/E2END[3] Tile_X9Y12_LUT4AB/E2END[4] Tile_X9Y12_LUT4AB/E2END[5]
+ Tile_X9Y12_LUT4AB/E2END[6] Tile_X9Y12_LUT4AB/E2END[7] Tile_X8Y12_LUT4AB/E2END[0]
+ Tile_X8Y12_LUT4AB/E2END[1] Tile_X8Y12_LUT4AB/E2END[2] Tile_X8Y12_LUT4AB/E2END[3]
+ Tile_X8Y12_LUT4AB/E2END[4] Tile_X8Y12_LUT4AB/E2END[5] Tile_X8Y12_LUT4AB/E2END[6]
+ Tile_X8Y12_LUT4AB/E2END[7] Tile_X8Y12_LUT4AB/E2MID[0] Tile_X8Y12_LUT4AB/E2MID[1]
+ Tile_X8Y12_LUT4AB/E2MID[2] Tile_X8Y12_LUT4AB/E2MID[3] Tile_X8Y12_LUT4AB/E2MID[4]
+ Tile_X8Y12_LUT4AB/E2MID[5] Tile_X8Y12_LUT4AB/E2MID[6] Tile_X8Y12_LUT4AB/E2MID[7]
+ Tile_X9Y12_LUT4AB/E6END[0] Tile_X9Y12_LUT4AB/E6END[10] Tile_X9Y12_LUT4AB/E6END[11]
+ Tile_X9Y12_LUT4AB/E6END[1] Tile_X9Y12_LUT4AB/E6END[2] Tile_X9Y12_LUT4AB/E6END[3]
+ Tile_X9Y12_LUT4AB/E6END[4] Tile_X9Y12_LUT4AB/E6END[5] Tile_X9Y12_LUT4AB/E6END[6]
+ Tile_X9Y12_LUT4AB/E6END[7] Tile_X9Y12_LUT4AB/E6END[8] Tile_X9Y12_LUT4AB/E6END[9]
+ Tile_X8Y12_LUT4AB/E6END[0] Tile_X8Y12_LUT4AB/E6END[10] Tile_X8Y12_LUT4AB/E6END[11]
+ Tile_X8Y12_LUT4AB/E6END[1] Tile_X8Y12_LUT4AB/E6END[2] Tile_X8Y12_LUT4AB/E6END[3]
+ Tile_X8Y12_LUT4AB/E6END[4] Tile_X8Y12_LUT4AB/E6END[5] Tile_X8Y12_LUT4AB/E6END[6]
+ Tile_X8Y12_LUT4AB/E6END[7] Tile_X8Y12_LUT4AB/E6END[8] Tile_X8Y12_LUT4AB/E6END[9]
+ Tile_X9Y12_LUT4AB/EE4END[0] Tile_X9Y12_LUT4AB/EE4END[10] Tile_X9Y12_LUT4AB/EE4END[11]
+ Tile_X9Y12_LUT4AB/EE4END[12] Tile_X9Y12_LUT4AB/EE4END[13] Tile_X9Y12_LUT4AB/EE4END[14]
+ Tile_X9Y12_LUT4AB/EE4END[15] Tile_X9Y12_LUT4AB/EE4END[1] Tile_X9Y12_LUT4AB/EE4END[2]
+ Tile_X9Y12_LUT4AB/EE4END[3] Tile_X9Y12_LUT4AB/EE4END[4] Tile_X9Y12_LUT4AB/EE4END[5]
+ Tile_X9Y12_LUT4AB/EE4END[6] Tile_X9Y12_LUT4AB/EE4END[7] Tile_X9Y12_LUT4AB/EE4END[8]
+ Tile_X9Y12_LUT4AB/EE4END[9] Tile_X8Y12_LUT4AB/EE4END[0] Tile_X8Y12_LUT4AB/EE4END[10]
+ Tile_X8Y12_LUT4AB/EE4END[11] Tile_X8Y12_LUT4AB/EE4END[12] Tile_X8Y12_LUT4AB/EE4END[13]
+ Tile_X8Y12_LUT4AB/EE4END[14] Tile_X8Y12_LUT4AB/EE4END[15] Tile_X8Y12_LUT4AB/EE4END[1]
+ Tile_X8Y12_LUT4AB/EE4END[2] Tile_X8Y12_LUT4AB/EE4END[3] Tile_X8Y12_LUT4AB/EE4END[4]
+ Tile_X8Y12_LUT4AB/EE4END[5] Tile_X8Y12_LUT4AB/EE4END[6] Tile_X8Y12_LUT4AB/EE4END[7]
+ Tile_X8Y12_LUT4AB/EE4END[8] Tile_X8Y12_LUT4AB/EE4END[9] Tile_X8Y12_LUT4AB/FrameData[0]
+ Tile_X8Y12_LUT4AB/FrameData[10] Tile_X8Y12_LUT4AB/FrameData[11] Tile_X8Y12_LUT4AB/FrameData[12]
+ Tile_X8Y12_LUT4AB/FrameData[13] Tile_X8Y12_LUT4AB/FrameData[14] Tile_X8Y12_LUT4AB/FrameData[15]
+ Tile_X8Y12_LUT4AB/FrameData[16] Tile_X8Y12_LUT4AB/FrameData[17] Tile_X8Y12_LUT4AB/FrameData[18]
+ Tile_X8Y12_LUT4AB/FrameData[19] Tile_X8Y12_LUT4AB/FrameData[1] Tile_X8Y12_LUT4AB/FrameData[20]
+ Tile_X8Y12_LUT4AB/FrameData[21] Tile_X8Y12_LUT4AB/FrameData[22] Tile_X8Y12_LUT4AB/FrameData[23]
+ Tile_X8Y12_LUT4AB/FrameData[24] Tile_X8Y12_LUT4AB/FrameData[25] Tile_X8Y12_LUT4AB/FrameData[26]
+ Tile_X8Y12_LUT4AB/FrameData[27] Tile_X8Y12_LUT4AB/FrameData[28] Tile_X8Y12_LUT4AB/FrameData[29]
+ Tile_X8Y12_LUT4AB/FrameData[2] Tile_X8Y12_LUT4AB/FrameData[30] Tile_X8Y12_LUT4AB/FrameData[31]
+ Tile_X8Y12_LUT4AB/FrameData[3] Tile_X8Y12_LUT4AB/FrameData[4] Tile_X8Y12_LUT4AB/FrameData[5]
+ Tile_X8Y12_LUT4AB/FrameData[6] Tile_X8Y12_LUT4AB/FrameData[7] Tile_X8Y12_LUT4AB/FrameData[8]
+ Tile_X8Y12_LUT4AB/FrameData[9] Tile_X9Y12_LUT4AB/FrameData[0] Tile_X9Y12_LUT4AB/FrameData[10]
+ Tile_X9Y12_LUT4AB/FrameData[11] Tile_X9Y12_LUT4AB/FrameData[12] Tile_X9Y12_LUT4AB/FrameData[13]
+ Tile_X9Y12_LUT4AB/FrameData[14] Tile_X9Y12_LUT4AB/FrameData[15] Tile_X9Y12_LUT4AB/FrameData[16]
+ Tile_X9Y12_LUT4AB/FrameData[17] Tile_X9Y12_LUT4AB/FrameData[18] Tile_X9Y12_LUT4AB/FrameData[19]
+ Tile_X9Y12_LUT4AB/FrameData[1] Tile_X9Y12_LUT4AB/FrameData[20] Tile_X9Y12_LUT4AB/FrameData[21]
+ Tile_X9Y12_LUT4AB/FrameData[22] Tile_X9Y12_LUT4AB/FrameData[23] Tile_X9Y12_LUT4AB/FrameData[24]
+ Tile_X9Y12_LUT4AB/FrameData[25] Tile_X9Y12_LUT4AB/FrameData[26] Tile_X9Y12_LUT4AB/FrameData[27]
+ Tile_X9Y12_LUT4AB/FrameData[28] Tile_X9Y12_LUT4AB/FrameData[29] Tile_X9Y12_LUT4AB/FrameData[2]
+ Tile_X9Y12_LUT4AB/FrameData[30] Tile_X9Y12_LUT4AB/FrameData[31] Tile_X9Y12_LUT4AB/FrameData[3]
+ Tile_X9Y12_LUT4AB/FrameData[4] Tile_X9Y12_LUT4AB/FrameData[5] Tile_X9Y12_LUT4AB/FrameData[6]
+ Tile_X9Y12_LUT4AB/FrameData[7] Tile_X9Y12_LUT4AB/FrameData[8] Tile_X9Y12_LUT4AB/FrameData[9]
+ Tile_X8Y12_LUT4AB/FrameStrobe[0] Tile_X8Y12_LUT4AB/FrameStrobe[10] Tile_X8Y12_LUT4AB/FrameStrobe[11]
+ Tile_X8Y12_LUT4AB/FrameStrobe[12] Tile_X8Y12_LUT4AB/FrameStrobe[13] Tile_X8Y12_LUT4AB/FrameStrobe[14]
+ Tile_X8Y12_LUT4AB/FrameStrobe[15] Tile_X8Y12_LUT4AB/FrameStrobe[16] Tile_X8Y12_LUT4AB/FrameStrobe[17]
+ Tile_X8Y12_LUT4AB/FrameStrobe[18] Tile_X8Y12_LUT4AB/FrameStrobe[19] Tile_X8Y12_LUT4AB/FrameStrobe[1]
+ Tile_X8Y12_LUT4AB/FrameStrobe[2] Tile_X8Y12_LUT4AB/FrameStrobe[3] Tile_X8Y12_LUT4AB/FrameStrobe[4]
+ Tile_X8Y12_LUT4AB/FrameStrobe[5] Tile_X8Y12_LUT4AB/FrameStrobe[6] Tile_X8Y12_LUT4AB/FrameStrobe[7]
+ Tile_X8Y12_LUT4AB/FrameStrobe[8] Tile_X8Y12_LUT4AB/FrameStrobe[9] Tile_X8Y11_LUT4AB/FrameStrobe[0]
+ Tile_X8Y11_LUT4AB/FrameStrobe[10] Tile_X8Y11_LUT4AB/FrameStrobe[11] Tile_X8Y11_LUT4AB/FrameStrobe[12]
+ Tile_X8Y11_LUT4AB/FrameStrobe[13] Tile_X8Y11_LUT4AB/FrameStrobe[14] Tile_X8Y11_LUT4AB/FrameStrobe[15]
+ Tile_X8Y11_LUT4AB/FrameStrobe[16] Tile_X8Y11_LUT4AB/FrameStrobe[17] Tile_X8Y11_LUT4AB/FrameStrobe[18]
+ Tile_X8Y11_LUT4AB/FrameStrobe[19] Tile_X8Y11_LUT4AB/FrameStrobe[1] Tile_X8Y11_LUT4AB/FrameStrobe[2]
+ Tile_X8Y11_LUT4AB/FrameStrobe[3] Tile_X8Y11_LUT4AB/FrameStrobe[4] Tile_X8Y11_LUT4AB/FrameStrobe[5]
+ Tile_X8Y11_LUT4AB/FrameStrobe[6] Tile_X8Y11_LUT4AB/FrameStrobe[7] Tile_X8Y11_LUT4AB/FrameStrobe[8]
+ Tile_X8Y11_LUT4AB/FrameStrobe[9] Tile_X8Y12_LUT4AB/N1BEG[0] Tile_X8Y12_LUT4AB/N1BEG[1]
+ Tile_X8Y12_LUT4AB/N1BEG[2] Tile_X8Y12_LUT4AB/N1BEG[3] Tile_X8Y13_LUT4AB/N1BEG[0]
+ Tile_X8Y13_LUT4AB/N1BEG[1] Tile_X8Y13_LUT4AB/N1BEG[2] Tile_X8Y13_LUT4AB/N1BEG[3]
+ Tile_X8Y12_LUT4AB/N2BEG[0] Tile_X8Y12_LUT4AB/N2BEG[1] Tile_X8Y12_LUT4AB/N2BEG[2]
+ Tile_X8Y12_LUT4AB/N2BEG[3] Tile_X8Y12_LUT4AB/N2BEG[4] Tile_X8Y12_LUT4AB/N2BEG[5]
+ Tile_X8Y12_LUT4AB/N2BEG[6] Tile_X8Y12_LUT4AB/N2BEG[7] Tile_X8Y11_LUT4AB/N2END[0]
+ Tile_X8Y11_LUT4AB/N2END[1] Tile_X8Y11_LUT4AB/N2END[2] Tile_X8Y11_LUT4AB/N2END[3]
+ Tile_X8Y11_LUT4AB/N2END[4] Tile_X8Y11_LUT4AB/N2END[5] Tile_X8Y11_LUT4AB/N2END[6]
+ Tile_X8Y11_LUT4AB/N2END[7] Tile_X8Y12_LUT4AB/N2END[0] Tile_X8Y12_LUT4AB/N2END[1]
+ Tile_X8Y12_LUT4AB/N2END[2] Tile_X8Y12_LUT4AB/N2END[3] Tile_X8Y12_LUT4AB/N2END[4]
+ Tile_X8Y12_LUT4AB/N2END[5] Tile_X8Y12_LUT4AB/N2END[6] Tile_X8Y12_LUT4AB/N2END[7]
+ Tile_X8Y13_LUT4AB/N2BEG[0] Tile_X8Y13_LUT4AB/N2BEG[1] Tile_X8Y13_LUT4AB/N2BEG[2]
+ Tile_X8Y13_LUT4AB/N2BEG[3] Tile_X8Y13_LUT4AB/N2BEG[4] Tile_X8Y13_LUT4AB/N2BEG[5]
+ Tile_X8Y13_LUT4AB/N2BEG[6] Tile_X8Y13_LUT4AB/N2BEG[7] Tile_X8Y12_LUT4AB/N4BEG[0]
+ Tile_X8Y12_LUT4AB/N4BEG[10] Tile_X8Y12_LUT4AB/N4BEG[11] Tile_X8Y12_LUT4AB/N4BEG[12]
+ Tile_X8Y12_LUT4AB/N4BEG[13] Tile_X8Y12_LUT4AB/N4BEG[14] Tile_X8Y12_LUT4AB/N4BEG[15]
+ Tile_X8Y12_LUT4AB/N4BEG[1] Tile_X8Y12_LUT4AB/N4BEG[2] Tile_X8Y12_LUT4AB/N4BEG[3]
+ Tile_X8Y12_LUT4AB/N4BEG[4] Tile_X8Y12_LUT4AB/N4BEG[5] Tile_X8Y12_LUT4AB/N4BEG[6]
+ Tile_X8Y12_LUT4AB/N4BEG[7] Tile_X8Y12_LUT4AB/N4BEG[8] Tile_X8Y12_LUT4AB/N4BEG[9]
+ Tile_X8Y13_LUT4AB/N4BEG[0] Tile_X8Y13_LUT4AB/N4BEG[10] Tile_X8Y13_LUT4AB/N4BEG[11]
+ Tile_X8Y13_LUT4AB/N4BEG[12] Tile_X8Y13_LUT4AB/N4BEG[13] Tile_X8Y13_LUT4AB/N4BEG[14]
+ Tile_X8Y13_LUT4AB/N4BEG[15] Tile_X8Y13_LUT4AB/N4BEG[1] Tile_X8Y13_LUT4AB/N4BEG[2]
+ Tile_X8Y13_LUT4AB/N4BEG[3] Tile_X8Y13_LUT4AB/N4BEG[4] Tile_X8Y13_LUT4AB/N4BEG[5]
+ Tile_X8Y13_LUT4AB/N4BEG[6] Tile_X8Y13_LUT4AB/N4BEG[7] Tile_X8Y13_LUT4AB/N4BEG[8]
+ Tile_X8Y13_LUT4AB/N4BEG[9] Tile_X8Y12_LUT4AB/NN4BEG[0] Tile_X8Y12_LUT4AB/NN4BEG[10]
+ Tile_X8Y12_LUT4AB/NN4BEG[11] Tile_X8Y12_LUT4AB/NN4BEG[12] Tile_X8Y12_LUT4AB/NN4BEG[13]
+ Tile_X8Y12_LUT4AB/NN4BEG[14] Tile_X8Y12_LUT4AB/NN4BEG[15] Tile_X8Y12_LUT4AB/NN4BEG[1]
+ Tile_X8Y12_LUT4AB/NN4BEG[2] Tile_X8Y12_LUT4AB/NN4BEG[3] Tile_X8Y12_LUT4AB/NN4BEG[4]
+ Tile_X8Y12_LUT4AB/NN4BEG[5] Tile_X8Y12_LUT4AB/NN4BEG[6] Tile_X8Y12_LUT4AB/NN4BEG[7]
+ Tile_X8Y12_LUT4AB/NN4BEG[8] Tile_X8Y12_LUT4AB/NN4BEG[9] Tile_X8Y13_LUT4AB/NN4BEG[0]
+ Tile_X8Y13_LUT4AB/NN4BEG[10] Tile_X8Y13_LUT4AB/NN4BEG[11] Tile_X8Y13_LUT4AB/NN4BEG[12]
+ Tile_X8Y13_LUT4AB/NN4BEG[13] Tile_X8Y13_LUT4AB/NN4BEG[14] Tile_X8Y13_LUT4AB/NN4BEG[15]
+ Tile_X8Y13_LUT4AB/NN4BEG[1] Tile_X8Y13_LUT4AB/NN4BEG[2] Tile_X8Y13_LUT4AB/NN4BEG[3]
+ Tile_X8Y13_LUT4AB/NN4BEG[4] Tile_X8Y13_LUT4AB/NN4BEG[5] Tile_X8Y13_LUT4AB/NN4BEG[6]
+ Tile_X8Y13_LUT4AB/NN4BEG[7] Tile_X8Y13_LUT4AB/NN4BEG[8] Tile_X8Y13_LUT4AB/NN4BEG[9]
+ Tile_X8Y13_LUT4AB/S1END[0] Tile_X8Y13_LUT4AB/S1END[1] Tile_X8Y13_LUT4AB/S1END[2]
+ Tile_X8Y13_LUT4AB/S1END[3] Tile_X8Y12_LUT4AB/S1END[0] Tile_X8Y12_LUT4AB/S1END[1]
+ Tile_X8Y12_LUT4AB/S1END[2] Tile_X8Y12_LUT4AB/S1END[3] Tile_X8Y13_LUT4AB/S2MID[0]
+ Tile_X8Y13_LUT4AB/S2MID[1] Tile_X8Y13_LUT4AB/S2MID[2] Tile_X8Y13_LUT4AB/S2MID[3]
+ Tile_X8Y13_LUT4AB/S2MID[4] Tile_X8Y13_LUT4AB/S2MID[5] Tile_X8Y13_LUT4AB/S2MID[6]
+ Tile_X8Y13_LUT4AB/S2MID[7] Tile_X8Y13_LUT4AB/S2END[0] Tile_X8Y13_LUT4AB/S2END[1]
+ Tile_X8Y13_LUT4AB/S2END[2] Tile_X8Y13_LUT4AB/S2END[3] Tile_X8Y13_LUT4AB/S2END[4]
+ Tile_X8Y13_LUT4AB/S2END[5] Tile_X8Y13_LUT4AB/S2END[6] Tile_X8Y13_LUT4AB/S2END[7]
+ Tile_X8Y12_LUT4AB/S2END[0] Tile_X8Y12_LUT4AB/S2END[1] Tile_X8Y12_LUT4AB/S2END[2]
+ Tile_X8Y12_LUT4AB/S2END[3] Tile_X8Y12_LUT4AB/S2END[4] Tile_X8Y12_LUT4AB/S2END[5]
+ Tile_X8Y12_LUT4AB/S2END[6] Tile_X8Y12_LUT4AB/S2END[7] Tile_X8Y12_LUT4AB/S2MID[0]
+ Tile_X8Y12_LUT4AB/S2MID[1] Tile_X8Y12_LUT4AB/S2MID[2] Tile_X8Y12_LUT4AB/S2MID[3]
+ Tile_X8Y12_LUT4AB/S2MID[4] Tile_X8Y12_LUT4AB/S2MID[5] Tile_X8Y12_LUT4AB/S2MID[6]
+ Tile_X8Y12_LUT4AB/S2MID[7] Tile_X8Y13_LUT4AB/S4END[0] Tile_X8Y13_LUT4AB/S4END[10]
+ Tile_X8Y13_LUT4AB/S4END[11] Tile_X8Y13_LUT4AB/S4END[12] Tile_X8Y13_LUT4AB/S4END[13]
+ Tile_X8Y13_LUT4AB/S4END[14] Tile_X8Y13_LUT4AB/S4END[15] Tile_X8Y13_LUT4AB/S4END[1]
+ Tile_X8Y13_LUT4AB/S4END[2] Tile_X8Y13_LUT4AB/S4END[3] Tile_X8Y13_LUT4AB/S4END[4]
+ Tile_X8Y13_LUT4AB/S4END[5] Tile_X8Y13_LUT4AB/S4END[6] Tile_X8Y13_LUT4AB/S4END[7]
+ Tile_X8Y13_LUT4AB/S4END[8] Tile_X8Y13_LUT4AB/S4END[9] Tile_X8Y12_LUT4AB/S4END[0]
+ Tile_X8Y12_LUT4AB/S4END[10] Tile_X8Y12_LUT4AB/S4END[11] Tile_X8Y12_LUT4AB/S4END[12]
+ Tile_X8Y12_LUT4AB/S4END[13] Tile_X8Y12_LUT4AB/S4END[14] Tile_X8Y12_LUT4AB/S4END[15]
+ Tile_X8Y12_LUT4AB/S4END[1] Tile_X8Y12_LUT4AB/S4END[2] Tile_X8Y12_LUT4AB/S4END[3]
+ Tile_X8Y12_LUT4AB/S4END[4] Tile_X8Y12_LUT4AB/S4END[5] Tile_X8Y12_LUT4AB/S4END[6]
+ Tile_X8Y12_LUT4AB/S4END[7] Tile_X8Y12_LUT4AB/S4END[8] Tile_X8Y12_LUT4AB/S4END[9]
+ Tile_X8Y13_LUT4AB/SS4END[0] Tile_X8Y13_LUT4AB/SS4END[10] Tile_X8Y13_LUT4AB/SS4END[11]
+ Tile_X8Y13_LUT4AB/SS4END[12] Tile_X8Y13_LUT4AB/SS4END[13] Tile_X8Y13_LUT4AB/SS4END[14]
+ Tile_X8Y13_LUT4AB/SS4END[15] Tile_X8Y13_LUT4AB/SS4END[1] Tile_X8Y13_LUT4AB/SS4END[2]
+ Tile_X8Y13_LUT4AB/SS4END[3] Tile_X8Y13_LUT4AB/SS4END[4] Tile_X8Y13_LUT4AB/SS4END[5]
+ Tile_X8Y13_LUT4AB/SS4END[6] Tile_X8Y13_LUT4AB/SS4END[7] Tile_X8Y13_LUT4AB/SS4END[8]
+ Tile_X8Y13_LUT4AB/SS4END[9] Tile_X8Y12_LUT4AB/SS4END[0] Tile_X8Y12_LUT4AB/SS4END[10]
+ Tile_X8Y12_LUT4AB/SS4END[11] Tile_X8Y12_LUT4AB/SS4END[12] Tile_X8Y12_LUT4AB/SS4END[13]
+ Tile_X8Y12_LUT4AB/SS4END[14] Tile_X8Y12_LUT4AB/SS4END[15] Tile_X8Y12_LUT4AB/SS4END[1]
+ Tile_X8Y12_LUT4AB/SS4END[2] Tile_X8Y12_LUT4AB/SS4END[3] Tile_X8Y12_LUT4AB/SS4END[4]
+ Tile_X8Y12_LUT4AB/SS4END[5] Tile_X8Y12_LUT4AB/SS4END[6] Tile_X8Y12_LUT4AB/SS4END[7]
+ Tile_X8Y12_LUT4AB/SS4END[8] Tile_X8Y12_LUT4AB/SS4END[9] Tile_X8Y12_LUT4AB/UserCLK
+ Tile_X8Y11_LUT4AB/UserCLK VGND VPWR Tile_X8Y12_LUT4AB/W1BEG[0] Tile_X8Y12_LUT4AB/W1BEG[1]
+ Tile_X8Y12_LUT4AB/W1BEG[2] Tile_X8Y12_LUT4AB/W1BEG[3] Tile_X9Y12_LUT4AB/W1BEG[0]
+ Tile_X9Y12_LUT4AB/W1BEG[1] Tile_X9Y12_LUT4AB/W1BEG[2] Tile_X9Y12_LUT4AB/W1BEG[3]
+ Tile_X8Y12_LUT4AB/W2BEG[0] Tile_X8Y12_LUT4AB/W2BEG[1] Tile_X8Y12_LUT4AB/W2BEG[2]
+ Tile_X8Y12_LUT4AB/W2BEG[3] Tile_X8Y12_LUT4AB/W2BEG[4] Tile_X8Y12_LUT4AB/W2BEG[5]
+ Tile_X8Y12_LUT4AB/W2BEG[6] Tile_X8Y12_LUT4AB/W2BEG[7] Tile_X8Y12_LUT4AB/W2BEGb[0]
+ Tile_X8Y12_LUT4AB/W2BEGb[1] Tile_X8Y12_LUT4AB/W2BEGb[2] Tile_X8Y12_LUT4AB/W2BEGb[3]
+ Tile_X8Y12_LUT4AB/W2BEGb[4] Tile_X8Y12_LUT4AB/W2BEGb[5] Tile_X8Y12_LUT4AB/W2BEGb[6]
+ Tile_X8Y12_LUT4AB/W2BEGb[7] Tile_X8Y12_LUT4AB/W2END[0] Tile_X8Y12_LUT4AB/W2END[1]
+ Tile_X8Y12_LUT4AB/W2END[2] Tile_X8Y12_LUT4AB/W2END[3] Tile_X8Y12_LUT4AB/W2END[4]
+ Tile_X8Y12_LUT4AB/W2END[5] Tile_X8Y12_LUT4AB/W2END[6] Tile_X8Y12_LUT4AB/W2END[7]
+ Tile_X9Y12_LUT4AB/W2BEG[0] Tile_X9Y12_LUT4AB/W2BEG[1] Tile_X9Y12_LUT4AB/W2BEG[2]
+ Tile_X9Y12_LUT4AB/W2BEG[3] Tile_X9Y12_LUT4AB/W2BEG[4] Tile_X9Y12_LUT4AB/W2BEG[5]
+ Tile_X9Y12_LUT4AB/W2BEG[6] Tile_X9Y12_LUT4AB/W2BEG[7] Tile_X8Y12_LUT4AB/W6BEG[0]
+ Tile_X8Y12_LUT4AB/W6BEG[10] Tile_X8Y12_LUT4AB/W6BEG[11] Tile_X8Y12_LUT4AB/W6BEG[1]
+ Tile_X8Y12_LUT4AB/W6BEG[2] Tile_X8Y12_LUT4AB/W6BEG[3] Tile_X8Y12_LUT4AB/W6BEG[4]
+ Tile_X8Y12_LUT4AB/W6BEG[5] Tile_X8Y12_LUT4AB/W6BEG[6] Tile_X8Y12_LUT4AB/W6BEG[7]
+ Tile_X8Y12_LUT4AB/W6BEG[8] Tile_X8Y12_LUT4AB/W6BEG[9] Tile_X9Y12_LUT4AB/W6BEG[0]
+ Tile_X9Y12_LUT4AB/W6BEG[10] Tile_X9Y12_LUT4AB/W6BEG[11] Tile_X9Y12_LUT4AB/W6BEG[1]
+ Tile_X9Y12_LUT4AB/W6BEG[2] Tile_X9Y12_LUT4AB/W6BEG[3] Tile_X9Y12_LUT4AB/W6BEG[4]
+ Tile_X9Y12_LUT4AB/W6BEG[5] Tile_X9Y12_LUT4AB/W6BEG[6] Tile_X9Y12_LUT4AB/W6BEG[7]
+ Tile_X9Y12_LUT4AB/W6BEG[8] Tile_X9Y12_LUT4AB/W6BEG[9] Tile_X8Y12_LUT4AB/WW4BEG[0]
+ Tile_X8Y12_LUT4AB/WW4BEG[10] Tile_X8Y12_LUT4AB/WW4BEG[11] Tile_X8Y12_LUT4AB/WW4BEG[12]
+ Tile_X8Y12_LUT4AB/WW4BEG[13] Tile_X8Y12_LUT4AB/WW4BEG[14] Tile_X8Y12_LUT4AB/WW4BEG[15]
+ Tile_X8Y12_LUT4AB/WW4BEG[1] Tile_X8Y12_LUT4AB/WW4BEG[2] Tile_X8Y12_LUT4AB/WW4BEG[3]
+ Tile_X8Y12_LUT4AB/WW4BEG[4] Tile_X8Y12_LUT4AB/WW4BEG[5] Tile_X8Y12_LUT4AB/WW4BEG[6]
+ Tile_X8Y12_LUT4AB/WW4BEG[7] Tile_X8Y12_LUT4AB/WW4BEG[8] Tile_X8Y12_LUT4AB/WW4BEG[9]
+ Tile_X9Y12_LUT4AB/WW4BEG[0] Tile_X9Y12_LUT4AB/WW4BEG[10] Tile_X9Y12_LUT4AB/WW4BEG[11]
+ Tile_X9Y12_LUT4AB/WW4BEG[12] Tile_X9Y12_LUT4AB/WW4BEG[13] Tile_X9Y12_LUT4AB/WW4BEG[14]
+ Tile_X9Y12_LUT4AB/WW4BEG[15] Tile_X9Y12_LUT4AB/WW4BEG[1] Tile_X9Y12_LUT4AB/WW4BEG[2]
+ Tile_X9Y12_LUT4AB/WW4BEG[3] Tile_X9Y12_LUT4AB/WW4BEG[4] Tile_X9Y12_LUT4AB/WW4BEG[5]
+ Tile_X9Y12_LUT4AB/WW4BEG[6] Tile_X9Y12_LUT4AB/WW4BEG[7] Tile_X9Y12_LUT4AB/WW4BEG[8]
+ Tile_X9Y12_LUT4AB/WW4BEG[9] LUT4AB
XTile_X2Y2_LUT4AB Tile_X2Y3_LUT4AB/Co Tile_X2Y2_LUT4AB/Co Tile_X3Y2_LUT4AB/E1END[0]
+ Tile_X3Y2_LUT4AB/E1END[1] Tile_X3Y2_LUT4AB/E1END[2] Tile_X3Y2_LUT4AB/E1END[3] Tile_X2Y2_LUT4AB/E1END[0]
+ Tile_X2Y2_LUT4AB/E1END[1] Tile_X2Y2_LUT4AB/E1END[2] Tile_X2Y2_LUT4AB/E1END[3] Tile_X3Y2_LUT4AB/E2MID[0]
+ Tile_X3Y2_LUT4AB/E2MID[1] Tile_X3Y2_LUT4AB/E2MID[2] Tile_X3Y2_LUT4AB/E2MID[3] Tile_X3Y2_LUT4AB/E2MID[4]
+ Tile_X3Y2_LUT4AB/E2MID[5] Tile_X3Y2_LUT4AB/E2MID[6] Tile_X3Y2_LUT4AB/E2MID[7] Tile_X3Y2_LUT4AB/E2END[0]
+ Tile_X3Y2_LUT4AB/E2END[1] Tile_X3Y2_LUT4AB/E2END[2] Tile_X3Y2_LUT4AB/E2END[3] Tile_X3Y2_LUT4AB/E2END[4]
+ Tile_X3Y2_LUT4AB/E2END[5] Tile_X3Y2_LUT4AB/E2END[6] Tile_X3Y2_LUT4AB/E2END[7] Tile_X2Y2_LUT4AB/E2END[0]
+ Tile_X2Y2_LUT4AB/E2END[1] Tile_X2Y2_LUT4AB/E2END[2] Tile_X2Y2_LUT4AB/E2END[3] Tile_X2Y2_LUT4AB/E2END[4]
+ Tile_X2Y2_LUT4AB/E2END[5] Tile_X2Y2_LUT4AB/E2END[6] Tile_X2Y2_LUT4AB/E2END[7] Tile_X2Y2_LUT4AB/E2MID[0]
+ Tile_X2Y2_LUT4AB/E2MID[1] Tile_X2Y2_LUT4AB/E2MID[2] Tile_X2Y2_LUT4AB/E2MID[3] Tile_X2Y2_LUT4AB/E2MID[4]
+ Tile_X2Y2_LUT4AB/E2MID[5] Tile_X2Y2_LUT4AB/E2MID[6] Tile_X2Y2_LUT4AB/E2MID[7] Tile_X3Y2_LUT4AB/E6END[0]
+ Tile_X3Y2_LUT4AB/E6END[10] Tile_X3Y2_LUT4AB/E6END[11] Tile_X3Y2_LUT4AB/E6END[1]
+ Tile_X3Y2_LUT4AB/E6END[2] Tile_X3Y2_LUT4AB/E6END[3] Tile_X3Y2_LUT4AB/E6END[4] Tile_X3Y2_LUT4AB/E6END[5]
+ Tile_X3Y2_LUT4AB/E6END[6] Tile_X3Y2_LUT4AB/E6END[7] Tile_X3Y2_LUT4AB/E6END[8] Tile_X3Y2_LUT4AB/E6END[9]
+ Tile_X2Y2_LUT4AB/E6END[0] Tile_X2Y2_LUT4AB/E6END[10] Tile_X2Y2_LUT4AB/E6END[11]
+ Tile_X2Y2_LUT4AB/E6END[1] Tile_X2Y2_LUT4AB/E6END[2] Tile_X2Y2_LUT4AB/E6END[3] Tile_X2Y2_LUT4AB/E6END[4]
+ Tile_X2Y2_LUT4AB/E6END[5] Tile_X2Y2_LUT4AB/E6END[6] Tile_X2Y2_LUT4AB/E6END[7] Tile_X2Y2_LUT4AB/E6END[8]
+ Tile_X2Y2_LUT4AB/E6END[9] Tile_X3Y2_LUT4AB/EE4END[0] Tile_X3Y2_LUT4AB/EE4END[10]
+ Tile_X3Y2_LUT4AB/EE4END[11] Tile_X3Y2_LUT4AB/EE4END[12] Tile_X3Y2_LUT4AB/EE4END[13]
+ Tile_X3Y2_LUT4AB/EE4END[14] Tile_X3Y2_LUT4AB/EE4END[15] Tile_X3Y2_LUT4AB/EE4END[1]
+ Tile_X3Y2_LUT4AB/EE4END[2] Tile_X3Y2_LUT4AB/EE4END[3] Tile_X3Y2_LUT4AB/EE4END[4]
+ Tile_X3Y2_LUT4AB/EE4END[5] Tile_X3Y2_LUT4AB/EE4END[6] Tile_X3Y2_LUT4AB/EE4END[7]
+ Tile_X3Y2_LUT4AB/EE4END[8] Tile_X3Y2_LUT4AB/EE4END[9] Tile_X2Y2_LUT4AB/EE4END[0]
+ Tile_X2Y2_LUT4AB/EE4END[10] Tile_X2Y2_LUT4AB/EE4END[11] Tile_X2Y2_LUT4AB/EE4END[12]
+ Tile_X2Y2_LUT4AB/EE4END[13] Tile_X2Y2_LUT4AB/EE4END[14] Tile_X2Y2_LUT4AB/EE4END[15]
+ Tile_X2Y2_LUT4AB/EE4END[1] Tile_X2Y2_LUT4AB/EE4END[2] Tile_X2Y2_LUT4AB/EE4END[3]
+ Tile_X2Y2_LUT4AB/EE4END[4] Tile_X2Y2_LUT4AB/EE4END[5] Tile_X2Y2_LUT4AB/EE4END[6]
+ Tile_X2Y2_LUT4AB/EE4END[7] Tile_X2Y2_LUT4AB/EE4END[8] Tile_X2Y2_LUT4AB/EE4END[9]
+ Tile_X2Y2_LUT4AB/FrameData[0] Tile_X2Y2_LUT4AB/FrameData[10] Tile_X2Y2_LUT4AB/FrameData[11]
+ Tile_X2Y2_LUT4AB/FrameData[12] Tile_X2Y2_LUT4AB/FrameData[13] Tile_X2Y2_LUT4AB/FrameData[14]
+ Tile_X2Y2_LUT4AB/FrameData[15] Tile_X2Y2_LUT4AB/FrameData[16] Tile_X2Y2_LUT4AB/FrameData[17]
+ Tile_X2Y2_LUT4AB/FrameData[18] Tile_X2Y2_LUT4AB/FrameData[19] Tile_X2Y2_LUT4AB/FrameData[1]
+ Tile_X2Y2_LUT4AB/FrameData[20] Tile_X2Y2_LUT4AB/FrameData[21] Tile_X2Y2_LUT4AB/FrameData[22]
+ Tile_X2Y2_LUT4AB/FrameData[23] Tile_X2Y2_LUT4AB/FrameData[24] Tile_X2Y2_LUT4AB/FrameData[25]
+ Tile_X2Y2_LUT4AB/FrameData[26] Tile_X2Y2_LUT4AB/FrameData[27] Tile_X2Y2_LUT4AB/FrameData[28]
+ Tile_X2Y2_LUT4AB/FrameData[29] Tile_X2Y2_LUT4AB/FrameData[2] Tile_X2Y2_LUT4AB/FrameData[30]
+ Tile_X2Y2_LUT4AB/FrameData[31] Tile_X2Y2_LUT4AB/FrameData[3] Tile_X2Y2_LUT4AB/FrameData[4]
+ Tile_X2Y2_LUT4AB/FrameData[5] Tile_X2Y2_LUT4AB/FrameData[6] Tile_X2Y2_LUT4AB/FrameData[7]
+ Tile_X2Y2_LUT4AB/FrameData[8] Tile_X2Y2_LUT4AB/FrameData[9] Tile_X3Y2_LUT4AB/FrameData[0]
+ Tile_X3Y2_LUT4AB/FrameData[10] Tile_X3Y2_LUT4AB/FrameData[11] Tile_X3Y2_LUT4AB/FrameData[12]
+ Tile_X3Y2_LUT4AB/FrameData[13] Tile_X3Y2_LUT4AB/FrameData[14] Tile_X3Y2_LUT4AB/FrameData[15]
+ Tile_X3Y2_LUT4AB/FrameData[16] Tile_X3Y2_LUT4AB/FrameData[17] Tile_X3Y2_LUT4AB/FrameData[18]
+ Tile_X3Y2_LUT4AB/FrameData[19] Tile_X3Y2_LUT4AB/FrameData[1] Tile_X3Y2_LUT4AB/FrameData[20]
+ Tile_X3Y2_LUT4AB/FrameData[21] Tile_X3Y2_LUT4AB/FrameData[22] Tile_X3Y2_LUT4AB/FrameData[23]
+ Tile_X3Y2_LUT4AB/FrameData[24] Tile_X3Y2_LUT4AB/FrameData[25] Tile_X3Y2_LUT4AB/FrameData[26]
+ Tile_X3Y2_LUT4AB/FrameData[27] Tile_X3Y2_LUT4AB/FrameData[28] Tile_X3Y2_LUT4AB/FrameData[29]
+ Tile_X3Y2_LUT4AB/FrameData[2] Tile_X3Y2_LUT4AB/FrameData[30] Tile_X3Y2_LUT4AB/FrameData[31]
+ Tile_X3Y2_LUT4AB/FrameData[3] Tile_X3Y2_LUT4AB/FrameData[4] Tile_X3Y2_LUT4AB/FrameData[5]
+ Tile_X3Y2_LUT4AB/FrameData[6] Tile_X3Y2_LUT4AB/FrameData[7] Tile_X3Y2_LUT4AB/FrameData[8]
+ Tile_X3Y2_LUT4AB/FrameData[9] Tile_X2Y2_LUT4AB/FrameStrobe[0] Tile_X2Y2_LUT4AB/FrameStrobe[10]
+ Tile_X2Y2_LUT4AB/FrameStrobe[11] Tile_X2Y2_LUT4AB/FrameStrobe[12] Tile_X2Y2_LUT4AB/FrameStrobe[13]
+ Tile_X2Y2_LUT4AB/FrameStrobe[14] Tile_X2Y2_LUT4AB/FrameStrobe[15] Tile_X2Y2_LUT4AB/FrameStrobe[16]
+ Tile_X2Y2_LUT4AB/FrameStrobe[17] Tile_X2Y2_LUT4AB/FrameStrobe[18] Tile_X2Y2_LUT4AB/FrameStrobe[19]
+ Tile_X2Y2_LUT4AB/FrameStrobe[1] Tile_X2Y2_LUT4AB/FrameStrobe[2] Tile_X2Y2_LUT4AB/FrameStrobe[3]
+ Tile_X2Y2_LUT4AB/FrameStrobe[4] Tile_X2Y2_LUT4AB/FrameStrobe[5] Tile_X2Y2_LUT4AB/FrameStrobe[6]
+ Tile_X2Y2_LUT4AB/FrameStrobe[7] Tile_X2Y2_LUT4AB/FrameStrobe[8] Tile_X2Y2_LUT4AB/FrameStrobe[9]
+ Tile_X2Y1_LUT4AB/FrameStrobe[0] Tile_X2Y1_LUT4AB/FrameStrobe[10] Tile_X2Y1_LUT4AB/FrameStrobe[11]
+ Tile_X2Y1_LUT4AB/FrameStrobe[12] Tile_X2Y1_LUT4AB/FrameStrobe[13] Tile_X2Y1_LUT4AB/FrameStrobe[14]
+ Tile_X2Y1_LUT4AB/FrameStrobe[15] Tile_X2Y1_LUT4AB/FrameStrobe[16] Tile_X2Y1_LUT4AB/FrameStrobe[17]
+ Tile_X2Y1_LUT4AB/FrameStrobe[18] Tile_X2Y1_LUT4AB/FrameStrobe[19] Tile_X2Y1_LUT4AB/FrameStrobe[1]
+ Tile_X2Y1_LUT4AB/FrameStrobe[2] Tile_X2Y1_LUT4AB/FrameStrobe[3] Tile_X2Y1_LUT4AB/FrameStrobe[4]
+ Tile_X2Y1_LUT4AB/FrameStrobe[5] Tile_X2Y1_LUT4AB/FrameStrobe[6] Tile_X2Y1_LUT4AB/FrameStrobe[7]
+ Tile_X2Y1_LUT4AB/FrameStrobe[8] Tile_X2Y1_LUT4AB/FrameStrobe[9] Tile_X2Y2_LUT4AB/N1BEG[0]
+ Tile_X2Y2_LUT4AB/N1BEG[1] Tile_X2Y2_LUT4AB/N1BEG[2] Tile_X2Y2_LUT4AB/N1BEG[3] Tile_X2Y3_LUT4AB/N1BEG[0]
+ Tile_X2Y3_LUT4AB/N1BEG[1] Tile_X2Y3_LUT4AB/N1BEG[2] Tile_X2Y3_LUT4AB/N1BEG[3] Tile_X2Y2_LUT4AB/N2BEG[0]
+ Tile_X2Y2_LUT4AB/N2BEG[1] Tile_X2Y2_LUT4AB/N2BEG[2] Tile_X2Y2_LUT4AB/N2BEG[3] Tile_X2Y2_LUT4AB/N2BEG[4]
+ Tile_X2Y2_LUT4AB/N2BEG[5] Tile_X2Y2_LUT4AB/N2BEG[6] Tile_X2Y2_LUT4AB/N2BEG[7] Tile_X2Y1_LUT4AB/N2END[0]
+ Tile_X2Y1_LUT4AB/N2END[1] Tile_X2Y1_LUT4AB/N2END[2] Tile_X2Y1_LUT4AB/N2END[3] Tile_X2Y1_LUT4AB/N2END[4]
+ Tile_X2Y1_LUT4AB/N2END[5] Tile_X2Y1_LUT4AB/N2END[6] Tile_X2Y1_LUT4AB/N2END[7] Tile_X2Y2_LUT4AB/N2END[0]
+ Tile_X2Y2_LUT4AB/N2END[1] Tile_X2Y2_LUT4AB/N2END[2] Tile_X2Y2_LUT4AB/N2END[3] Tile_X2Y2_LUT4AB/N2END[4]
+ Tile_X2Y2_LUT4AB/N2END[5] Tile_X2Y2_LUT4AB/N2END[6] Tile_X2Y2_LUT4AB/N2END[7] Tile_X2Y3_LUT4AB/N2BEG[0]
+ Tile_X2Y3_LUT4AB/N2BEG[1] Tile_X2Y3_LUT4AB/N2BEG[2] Tile_X2Y3_LUT4AB/N2BEG[3] Tile_X2Y3_LUT4AB/N2BEG[4]
+ Tile_X2Y3_LUT4AB/N2BEG[5] Tile_X2Y3_LUT4AB/N2BEG[6] Tile_X2Y3_LUT4AB/N2BEG[7] Tile_X2Y2_LUT4AB/N4BEG[0]
+ Tile_X2Y2_LUT4AB/N4BEG[10] Tile_X2Y2_LUT4AB/N4BEG[11] Tile_X2Y2_LUT4AB/N4BEG[12]
+ Tile_X2Y2_LUT4AB/N4BEG[13] Tile_X2Y2_LUT4AB/N4BEG[14] Tile_X2Y2_LUT4AB/N4BEG[15]
+ Tile_X2Y2_LUT4AB/N4BEG[1] Tile_X2Y2_LUT4AB/N4BEG[2] Tile_X2Y2_LUT4AB/N4BEG[3] Tile_X2Y2_LUT4AB/N4BEG[4]
+ Tile_X2Y2_LUT4AB/N4BEG[5] Tile_X2Y2_LUT4AB/N4BEG[6] Tile_X2Y2_LUT4AB/N4BEG[7] Tile_X2Y2_LUT4AB/N4BEG[8]
+ Tile_X2Y2_LUT4AB/N4BEG[9] Tile_X2Y3_LUT4AB/N4BEG[0] Tile_X2Y3_LUT4AB/N4BEG[10] Tile_X2Y3_LUT4AB/N4BEG[11]
+ Tile_X2Y3_LUT4AB/N4BEG[12] Tile_X2Y3_LUT4AB/N4BEG[13] Tile_X2Y3_LUT4AB/N4BEG[14]
+ Tile_X2Y3_LUT4AB/N4BEG[15] Tile_X2Y3_LUT4AB/N4BEG[1] Tile_X2Y3_LUT4AB/N4BEG[2] Tile_X2Y3_LUT4AB/N4BEG[3]
+ Tile_X2Y3_LUT4AB/N4BEG[4] Tile_X2Y3_LUT4AB/N4BEG[5] Tile_X2Y3_LUT4AB/N4BEG[6] Tile_X2Y3_LUT4AB/N4BEG[7]
+ Tile_X2Y3_LUT4AB/N4BEG[8] Tile_X2Y3_LUT4AB/N4BEG[9] Tile_X2Y2_LUT4AB/NN4BEG[0] Tile_X2Y2_LUT4AB/NN4BEG[10]
+ Tile_X2Y2_LUT4AB/NN4BEG[11] Tile_X2Y2_LUT4AB/NN4BEG[12] Tile_X2Y2_LUT4AB/NN4BEG[13]
+ Tile_X2Y2_LUT4AB/NN4BEG[14] Tile_X2Y2_LUT4AB/NN4BEG[15] Tile_X2Y2_LUT4AB/NN4BEG[1]
+ Tile_X2Y2_LUT4AB/NN4BEG[2] Tile_X2Y2_LUT4AB/NN4BEG[3] Tile_X2Y2_LUT4AB/NN4BEG[4]
+ Tile_X2Y2_LUT4AB/NN4BEG[5] Tile_X2Y2_LUT4AB/NN4BEG[6] Tile_X2Y2_LUT4AB/NN4BEG[7]
+ Tile_X2Y2_LUT4AB/NN4BEG[8] Tile_X2Y2_LUT4AB/NN4BEG[9] Tile_X2Y3_LUT4AB/NN4BEG[0]
+ Tile_X2Y3_LUT4AB/NN4BEG[10] Tile_X2Y3_LUT4AB/NN4BEG[11] Tile_X2Y3_LUT4AB/NN4BEG[12]
+ Tile_X2Y3_LUT4AB/NN4BEG[13] Tile_X2Y3_LUT4AB/NN4BEG[14] Tile_X2Y3_LUT4AB/NN4BEG[15]
+ Tile_X2Y3_LUT4AB/NN4BEG[1] Tile_X2Y3_LUT4AB/NN4BEG[2] Tile_X2Y3_LUT4AB/NN4BEG[3]
+ Tile_X2Y3_LUT4AB/NN4BEG[4] Tile_X2Y3_LUT4AB/NN4BEG[5] Tile_X2Y3_LUT4AB/NN4BEG[6]
+ Tile_X2Y3_LUT4AB/NN4BEG[7] Tile_X2Y3_LUT4AB/NN4BEG[8] Tile_X2Y3_LUT4AB/NN4BEG[9]
+ Tile_X2Y3_LUT4AB/S1END[0] Tile_X2Y3_LUT4AB/S1END[1] Tile_X2Y3_LUT4AB/S1END[2] Tile_X2Y3_LUT4AB/S1END[3]
+ Tile_X2Y2_LUT4AB/S1END[0] Tile_X2Y2_LUT4AB/S1END[1] Tile_X2Y2_LUT4AB/S1END[2] Tile_X2Y2_LUT4AB/S1END[3]
+ Tile_X2Y3_LUT4AB/S2MID[0] Tile_X2Y3_LUT4AB/S2MID[1] Tile_X2Y3_LUT4AB/S2MID[2] Tile_X2Y3_LUT4AB/S2MID[3]
+ Tile_X2Y3_LUT4AB/S2MID[4] Tile_X2Y3_LUT4AB/S2MID[5] Tile_X2Y3_LUT4AB/S2MID[6] Tile_X2Y3_LUT4AB/S2MID[7]
+ Tile_X2Y3_LUT4AB/S2END[0] Tile_X2Y3_LUT4AB/S2END[1] Tile_X2Y3_LUT4AB/S2END[2] Tile_X2Y3_LUT4AB/S2END[3]
+ Tile_X2Y3_LUT4AB/S2END[4] Tile_X2Y3_LUT4AB/S2END[5] Tile_X2Y3_LUT4AB/S2END[6] Tile_X2Y3_LUT4AB/S2END[7]
+ Tile_X2Y2_LUT4AB/S2END[0] Tile_X2Y2_LUT4AB/S2END[1] Tile_X2Y2_LUT4AB/S2END[2] Tile_X2Y2_LUT4AB/S2END[3]
+ Tile_X2Y2_LUT4AB/S2END[4] Tile_X2Y2_LUT4AB/S2END[5] Tile_X2Y2_LUT4AB/S2END[6] Tile_X2Y2_LUT4AB/S2END[7]
+ Tile_X2Y2_LUT4AB/S2MID[0] Tile_X2Y2_LUT4AB/S2MID[1] Tile_X2Y2_LUT4AB/S2MID[2] Tile_X2Y2_LUT4AB/S2MID[3]
+ Tile_X2Y2_LUT4AB/S2MID[4] Tile_X2Y2_LUT4AB/S2MID[5] Tile_X2Y2_LUT4AB/S2MID[6] Tile_X2Y2_LUT4AB/S2MID[7]
+ Tile_X2Y3_LUT4AB/S4END[0] Tile_X2Y3_LUT4AB/S4END[10] Tile_X2Y3_LUT4AB/S4END[11]
+ Tile_X2Y3_LUT4AB/S4END[12] Tile_X2Y3_LUT4AB/S4END[13] Tile_X2Y3_LUT4AB/S4END[14]
+ Tile_X2Y3_LUT4AB/S4END[15] Tile_X2Y3_LUT4AB/S4END[1] Tile_X2Y3_LUT4AB/S4END[2] Tile_X2Y3_LUT4AB/S4END[3]
+ Tile_X2Y3_LUT4AB/S4END[4] Tile_X2Y3_LUT4AB/S4END[5] Tile_X2Y3_LUT4AB/S4END[6] Tile_X2Y3_LUT4AB/S4END[7]
+ Tile_X2Y3_LUT4AB/S4END[8] Tile_X2Y3_LUT4AB/S4END[9] Tile_X2Y2_LUT4AB/S4END[0] Tile_X2Y2_LUT4AB/S4END[10]
+ Tile_X2Y2_LUT4AB/S4END[11] Tile_X2Y2_LUT4AB/S4END[12] Tile_X2Y2_LUT4AB/S4END[13]
+ Tile_X2Y2_LUT4AB/S4END[14] Tile_X2Y2_LUT4AB/S4END[15] Tile_X2Y2_LUT4AB/S4END[1]
+ Tile_X2Y2_LUT4AB/S4END[2] Tile_X2Y2_LUT4AB/S4END[3] Tile_X2Y2_LUT4AB/S4END[4] Tile_X2Y2_LUT4AB/S4END[5]
+ Tile_X2Y2_LUT4AB/S4END[6] Tile_X2Y2_LUT4AB/S4END[7] Tile_X2Y2_LUT4AB/S4END[8] Tile_X2Y2_LUT4AB/S4END[9]
+ Tile_X2Y3_LUT4AB/SS4END[0] Tile_X2Y3_LUT4AB/SS4END[10] Tile_X2Y3_LUT4AB/SS4END[11]
+ Tile_X2Y3_LUT4AB/SS4END[12] Tile_X2Y3_LUT4AB/SS4END[13] Tile_X2Y3_LUT4AB/SS4END[14]
+ Tile_X2Y3_LUT4AB/SS4END[15] Tile_X2Y3_LUT4AB/SS4END[1] Tile_X2Y3_LUT4AB/SS4END[2]
+ Tile_X2Y3_LUT4AB/SS4END[3] Tile_X2Y3_LUT4AB/SS4END[4] Tile_X2Y3_LUT4AB/SS4END[5]
+ Tile_X2Y3_LUT4AB/SS4END[6] Tile_X2Y3_LUT4AB/SS4END[7] Tile_X2Y3_LUT4AB/SS4END[8]
+ Tile_X2Y3_LUT4AB/SS4END[9] Tile_X2Y2_LUT4AB/SS4END[0] Tile_X2Y2_LUT4AB/SS4END[10]
+ Tile_X2Y2_LUT4AB/SS4END[11] Tile_X2Y2_LUT4AB/SS4END[12] Tile_X2Y2_LUT4AB/SS4END[13]
+ Tile_X2Y2_LUT4AB/SS4END[14] Tile_X2Y2_LUT4AB/SS4END[15] Tile_X2Y2_LUT4AB/SS4END[1]
+ Tile_X2Y2_LUT4AB/SS4END[2] Tile_X2Y2_LUT4AB/SS4END[3] Tile_X2Y2_LUT4AB/SS4END[4]
+ Tile_X2Y2_LUT4AB/SS4END[5] Tile_X2Y2_LUT4AB/SS4END[6] Tile_X2Y2_LUT4AB/SS4END[7]
+ Tile_X2Y2_LUT4AB/SS4END[8] Tile_X2Y2_LUT4AB/SS4END[9] Tile_X2Y2_LUT4AB/UserCLK Tile_X2Y1_LUT4AB/UserCLK
+ VGND VPWR Tile_X2Y2_LUT4AB/W1BEG[0] Tile_X2Y2_LUT4AB/W1BEG[1] Tile_X2Y2_LUT4AB/W1BEG[2]
+ Tile_X2Y2_LUT4AB/W1BEG[3] Tile_X3Y2_LUT4AB/W1BEG[0] Tile_X3Y2_LUT4AB/W1BEG[1] Tile_X3Y2_LUT4AB/W1BEG[2]
+ Tile_X3Y2_LUT4AB/W1BEG[3] Tile_X2Y2_LUT4AB/W2BEG[0] Tile_X2Y2_LUT4AB/W2BEG[1] Tile_X2Y2_LUT4AB/W2BEG[2]
+ Tile_X2Y2_LUT4AB/W2BEG[3] Tile_X2Y2_LUT4AB/W2BEG[4] Tile_X2Y2_LUT4AB/W2BEG[5] Tile_X2Y2_LUT4AB/W2BEG[6]
+ Tile_X2Y2_LUT4AB/W2BEG[7] Tile_X1Y2_LUT4AB/W2END[0] Tile_X1Y2_LUT4AB/W2END[1] Tile_X1Y2_LUT4AB/W2END[2]
+ Tile_X1Y2_LUT4AB/W2END[3] Tile_X1Y2_LUT4AB/W2END[4] Tile_X1Y2_LUT4AB/W2END[5] Tile_X1Y2_LUT4AB/W2END[6]
+ Tile_X1Y2_LUT4AB/W2END[7] Tile_X2Y2_LUT4AB/W2END[0] Tile_X2Y2_LUT4AB/W2END[1] Tile_X2Y2_LUT4AB/W2END[2]
+ Tile_X2Y2_LUT4AB/W2END[3] Tile_X2Y2_LUT4AB/W2END[4] Tile_X2Y2_LUT4AB/W2END[5] Tile_X2Y2_LUT4AB/W2END[6]
+ Tile_X2Y2_LUT4AB/W2END[7] Tile_X3Y2_LUT4AB/W2BEG[0] Tile_X3Y2_LUT4AB/W2BEG[1] Tile_X3Y2_LUT4AB/W2BEG[2]
+ Tile_X3Y2_LUT4AB/W2BEG[3] Tile_X3Y2_LUT4AB/W2BEG[4] Tile_X3Y2_LUT4AB/W2BEG[5] Tile_X3Y2_LUT4AB/W2BEG[6]
+ Tile_X3Y2_LUT4AB/W2BEG[7] Tile_X2Y2_LUT4AB/W6BEG[0] Tile_X2Y2_LUT4AB/W6BEG[10] Tile_X2Y2_LUT4AB/W6BEG[11]
+ Tile_X2Y2_LUT4AB/W6BEG[1] Tile_X2Y2_LUT4AB/W6BEG[2] Tile_X2Y2_LUT4AB/W6BEG[3] Tile_X2Y2_LUT4AB/W6BEG[4]
+ Tile_X2Y2_LUT4AB/W6BEG[5] Tile_X2Y2_LUT4AB/W6BEG[6] Tile_X2Y2_LUT4AB/W6BEG[7] Tile_X2Y2_LUT4AB/W6BEG[8]
+ Tile_X2Y2_LUT4AB/W6BEG[9] Tile_X3Y2_LUT4AB/W6BEG[0] Tile_X3Y2_LUT4AB/W6BEG[10] Tile_X3Y2_LUT4AB/W6BEG[11]
+ Tile_X3Y2_LUT4AB/W6BEG[1] Tile_X3Y2_LUT4AB/W6BEG[2] Tile_X3Y2_LUT4AB/W6BEG[3] Tile_X3Y2_LUT4AB/W6BEG[4]
+ Tile_X3Y2_LUT4AB/W6BEG[5] Tile_X3Y2_LUT4AB/W6BEG[6] Tile_X3Y2_LUT4AB/W6BEG[7] Tile_X3Y2_LUT4AB/W6BEG[8]
+ Tile_X3Y2_LUT4AB/W6BEG[9] Tile_X2Y2_LUT4AB/WW4BEG[0] Tile_X2Y2_LUT4AB/WW4BEG[10]
+ Tile_X2Y2_LUT4AB/WW4BEG[11] Tile_X2Y2_LUT4AB/WW4BEG[12] Tile_X2Y2_LUT4AB/WW4BEG[13]
+ Tile_X2Y2_LUT4AB/WW4BEG[14] Tile_X2Y2_LUT4AB/WW4BEG[15] Tile_X2Y2_LUT4AB/WW4BEG[1]
+ Tile_X2Y2_LUT4AB/WW4BEG[2] Tile_X2Y2_LUT4AB/WW4BEG[3] Tile_X2Y2_LUT4AB/WW4BEG[4]
+ Tile_X2Y2_LUT4AB/WW4BEG[5] Tile_X2Y2_LUT4AB/WW4BEG[6] Tile_X2Y2_LUT4AB/WW4BEG[7]
+ Tile_X2Y2_LUT4AB/WW4BEG[8] Tile_X2Y2_LUT4AB/WW4BEG[9] Tile_X3Y2_LUT4AB/WW4BEG[0]
+ Tile_X3Y2_LUT4AB/WW4BEG[10] Tile_X3Y2_LUT4AB/WW4BEG[11] Tile_X3Y2_LUT4AB/WW4BEG[12]
+ Tile_X3Y2_LUT4AB/WW4BEG[13] Tile_X3Y2_LUT4AB/WW4BEG[14] Tile_X3Y2_LUT4AB/WW4BEG[15]
+ Tile_X3Y2_LUT4AB/WW4BEG[1] Tile_X3Y2_LUT4AB/WW4BEG[2] Tile_X3Y2_LUT4AB/WW4BEG[3]
+ Tile_X3Y2_LUT4AB/WW4BEG[4] Tile_X3Y2_LUT4AB/WW4BEG[5] Tile_X3Y2_LUT4AB/WW4BEG[6]
+ Tile_X3Y2_LUT4AB/WW4BEG[7] Tile_X3Y2_LUT4AB/WW4BEG[8] Tile_X3Y2_LUT4AB/WW4BEG[9]
+ LUT4AB
XTile_X5Y7_LUT4AB Tile_X5Y8_LUT4AB/Co Tile_X5Y7_LUT4AB/Co Tile_X6Y7_LUT4AB/E1END[0]
+ Tile_X6Y7_LUT4AB/E1END[1] Tile_X6Y7_LUT4AB/E1END[2] Tile_X6Y7_LUT4AB/E1END[3] Tile_X5Y7_LUT4AB/E1END[0]
+ Tile_X5Y7_LUT4AB/E1END[1] Tile_X5Y7_LUT4AB/E1END[2] Tile_X5Y7_LUT4AB/E1END[3] Tile_X6Y7_LUT4AB/E2MID[0]
+ Tile_X6Y7_LUT4AB/E2MID[1] Tile_X6Y7_LUT4AB/E2MID[2] Tile_X6Y7_LUT4AB/E2MID[3] Tile_X6Y7_LUT4AB/E2MID[4]
+ Tile_X6Y7_LUT4AB/E2MID[5] Tile_X6Y7_LUT4AB/E2MID[6] Tile_X6Y7_LUT4AB/E2MID[7] Tile_X6Y7_LUT4AB/E2END[0]
+ Tile_X6Y7_LUT4AB/E2END[1] Tile_X6Y7_LUT4AB/E2END[2] Tile_X6Y7_LUT4AB/E2END[3] Tile_X6Y7_LUT4AB/E2END[4]
+ Tile_X6Y7_LUT4AB/E2END[5] Tile_X6Y7_LUT4AB/E2END[6] Tile_X6Y7_LUT4AB/E2END[7] Tile_X5Y7_LUT4AB/E2END[0]
+ Tile_X5Y7_LUT4AB/E2END[1] Tile_X5Y7_LUT4AB/E2END[2] Tile_X5Y7_LUT4AB/E2END[3] Tile_X5Y7_LUT4AB/E2END[4]
+ Tile_X5Y7_LUT4AB/E2END[5] Tile_X5Y7_LUT4AB/E2END[6] Tile_X5Y7_LUT4AB/E2END[7] Tile_X5Y7_LUT4AB/E2MID[0]
+ Tile_X5Y7_LUT4AB/E2MID[1] Tile_X5Y7_LUT4AB/E2MID[2] Tile_X5Y7_LUT4AB/E2MID[3] Tile_X5Y7_LUT4AB/E2MID[4]
+ Tile_X5Y7_LUT4AB/E2MID[5] Tile_X5Y7_LUT4AB/E2MID[6] Tile_X5Y7_LUT4AB/E2MID[7] Tile_X6Y7_LUT4AB/E6END[0]
+ Tile_X6Y7_LUT4AB/E6END[10] Tile_X6Y7_LUT4AB/E6END[11] Tile_X6Y7_LUT4AB/E6END[1]
+ Tile_X6Y7_LUT4AB/E6END[2] Tile_X6Y7_LUT4AB/E6END[3] Tile_X6Y7_LUT4AB/E6END[4] Tile_X6Y7_LUT4AB/E6END[5]
+ Tile_X6Y7_LUT4AB/E6END[6] Tile_X6Y7_LUT4AB/E6END[7] Tile_X6Y7_LUT4AB/E6END[8] Tile_X6Y7_LUT4AB/E6END[9]
+ Tile_X5Y7_LUT4AB/E6END[0] Tile_X5Y7_LUT4AB/E6END[10] Tile_X5Y7_LUT4AB/E6END[11]
+ Tile_X5Y7_LUT4AB/E6END[1] Tile_X5Y7_LUT4AB/E6END[2] Tile_X5Y7_LUT4AB/E6END[3] Tile_X5Y7_LUT4AB/E6END[4]
+ Tile_X5Y7_LUT4AB/E6END[5] Tile_X5Y7_LUT4AB/E6END[6] Tile_X5Y7_LUT4AB/E6END[7] Tile_X5Y7_LUT4AB/E6END[8]
+ Tile_X5Y7_LUT4AB/E6END[9] Tile_X6Y7_LUT4AB/EE4END[0] Tile_X6Y7_LUT4AB/EE4END[10]
+ Tile_X6Y7_LUT4AB/EE4END[11] Tile_X6Y7_LUT4AB/EE4END[12] Tile_X6Y7_LUT4AB/EE4END[13]
+ Tile_X6Y7_LUT4AB/EE4END[14] Tile_X6Y7_LUT4AB/EE4END[15] Tile_X6Y7_LUT4AB/EE4END[1]
+ Tile_X6Y7_LUT4AB/EE4END[2] Tile_X6Y7_LUT4AB/EE4END[3] Tile_X6Y7_LUT4AB/EE4END[4]
+ Tile_X6Y7_LUT4AB/EE4END[5] Tile_X6Y7_LUT4AB/EE4END[6] Tile_X6Y7_LUT4AB/EE4END[7]
+ Tile_X6Y7_LUT4AB/EE4END[8] Tile_X6Y7_LUT4AB/EE4END[9] Tile_X5Y7_LUT4AB/EE4END[0]
+ Tile_X5Y7_LUT4AB/EE4END[10] Tile_X5Y7_LUT4AB/EE4END[11] Tile_X5Y7_LUT4AB/EE4END[12]
+ Tile_X5Y7_LUT4AB/EE4END[13] Tile_X5Y7_LUT4AB/EE4END[14] Tile_X5Y7_LUT4AB/EE4END[15]
+ Tile_X5Y7_LUT4AB/EE4END[1] Tile_X5Y7_LUT4AB/EE4END[2] Tile_X5Y7_LUT4AB/EE4END[3]
+ Tile_X5Y7_LUT4AB/EE4END[4] Tile_X5Y7_LUT4AB/EE4END[5] Tile_X5Y7_LUT4AB/EE4END[6]
+ Tile_X5Y7_LUT4AB/EE4END[7] Tile_X5Y7_LUT4AB/EE4END[8] Tile_X5Y7_LUT4AB/EE4END[9]
+ Tile_X5Y7_LUT4AB/FrameData[0] Tile_X5Y7_LUT4AB/FrameData[10] Tile_X5Y7_LUT4AB/FrameData[11]
+ Tile_X5Y7_LUT4AB/FrameData[12] Tile_X5Y7_LUT4AB/FrameData[13] Tile_X5Y7_LUT4AB/FrameData[14]
+ Tile_X5Y7_LUT4AB/FrameData[15] Tile_X5Y7_LUT4AB/FrameData[16] Tile_X5Y7_LUT4AB/FrameData[17]
+ Tile_X5Y7_LUT4AB/FrameData[18] Tile_X5Y7_LUT4AB/FrameData[19] Tile_X5Y7_LUT4AB/FrameData[1]
+ Tile_X5Y7_LUT4AB/FrameData[20] Tile_X5Y7_LUT4AB/FrameData[21] Tile_X5Y7_LUT4AB/FrameData[22]
+ Tile_X5Y7_LUT4AB/FrameData[23] Tile_X5Y7_LUT4AB/FrameData[24] Tile_X5Y7_LUT4AB/FrameData[25]
+ Tile_X5Y7_LUT4AB/FrameData[26] Tile_X5Y7_LUT4AB/FrameData[27] Tile_X5Y7_LUT4AB/FrameData[28]
+ Tile_X5Y7_LUT4AB/FrameData[29] Tile_X5Y7_LUT4AB/FrameData[2] Tile_X5Y7_LUT4AB/FrameData[30]
+ Tile_X5Y7_LUT4AB/FrameData[31] Tile_X5Y7_LUT4AB/FrameData[3] Tile_X5Y7_LUT4AB/FrameData[4]
+ Tile_X5Y7_LUT4AB/FrameData[5] Tile_X5Y7_LUT4AB/FrameData[6] Tile_X5Y7_LUT4AB/FrameData[7]
+ Tile_X5Y7_LUT4AB/FrameData[8] Tile_X5Y7_LUT4AB/FrameData[9] Tile_X6Y7_LUT4AB/FrameData[0]
+ Tile_X6Y7_LUT4AB/FrameData[10] Tile_X6Y7_LUT4AB/FrameData[11] Tile_X6Y7_LUT4AB/FrameData[12]
+ Tile_X6Y7_LUT4AB/FrameData[13] Tile_X6Y7_LUT4AB/FrameData[14] Tile_X6Y7_LUT4AB/FrameData[15]
+ Tile_X6Y7_LUT4AB/FrameData[16] Tile_X6Y7_LUT4AB/FrameData[17] Tile_X6Y7_LUT4AB/FrameData[18]
+ Tile_X6Y7_LUT4AB/FrameData[19] Tile_X6Y7_LUT4AB/FrameData[1] Tile_X6Y7_LUT4AB/FrameData[20]
+ Tile_X6Y7_LUT4AB/FrameData[21] Tile_X6Y7_LUT4AB/FrameData[22] Tile_X6Y7_LUT4AB/FrameData[23]
+ Tile_X6Y7_LUT4AB/FrameData[24] Tile_X6Y7_LUT4AB/FrameData[25] Tile_X6Y7_LUT4AB/FrameData[26]
+ Tile_X6Y7_LUT4AB/FrameData[27] Tile_X6Y7_LUT4AB/FrameData[28] Tile_X6Y7_LUT4AB/FrameData[29]
+ Tile_X6Y7_LUT4AB/FrameData[2] Tile_X6Y7_LUT4AB/FrameData[30] Tile_X6Y7_LUT4AB/FrameData[31]
+ Tile_X6Y7_LUT4AB/FrameData[3] Tile_X6Y7_LUT4AB/FrameData[4] Tile_X6Y7_LUT4AB/FrameData[5]
+ Tile_X6Y7_LUT4AB/FrameData[6] Tile_X6Y7_LUT4AB/FrameData[7] Tile_X6Y7_LUT4AB/FrameData[8]
+ Tile_X6Y7_LUT4AB/FrameData[9] Tile_X5Y7_LUT4AB/FrameStrobe[0] Tile_X5Y7_LUT4AB/FrameStrobe[10]
+ Tile_X5Y7_LUT4AB/FrameStrobe[11] Tile_X5Y7_LUT4AB/FrameStrobe[12] Tile_X5Y7_LUT4AB/FrameStrobe[13]
+ Tile_X5Y7_LUT4AB/FrameStrobe[14] Tile_X5Y7_LUT4AB/FrameStrobe[15] Tile_X5Y7_LUT4AB/FrameStrobe[16]
+ Tile_X5Y7_LUT4AB/FrameStrobe[17] Tile_X5Y7_LUT4AB/FrameStrobe[18] Tile_X5Y7_LUT4AB/FrameStrobe[19]
+ Tile_X5Y7_LUT4AB/FrameStrobe[1] Tile_X5Y7_LUT4AB/FrameStrobe[2] Tile_X5Y7_LUT4AB/FrameStrobe[3]
+ Tile_X5Y7_LUT4AB/FrameStrobe[4] Tile_X5Y7_LUT4AB/FrameStrobe[5] Tile_X5Y7_LUT4AB/FrameStrobe[6]
+ Tile_X5Y7_LUT4AB/FrameStrobe[7] Tile_X5Y7_LUT4AB/FrameStrobe[8] Tile_X5Y7_LUT4AB/FrameStrobe[9]
+ Tile_X5Y6_LUT4AB/FrameStrobe[0] Tile_X5Y6_LUT4AB/FrameStrobe[10] Tile_X5Y6_LUT4AB/FrameStrobe[11]
+ Tile_X5Y6_LUT4AB/FrameStrobe[12] Tile_X5Y6_LUT4AB/FrameStrobe[13] Tile_X5Y6_LUT4AB/FrameStrobe[14]
+ Tile_X5Y6_LUT4AB/FrameStrobe[15] Tile_X5Y6_LUT4AB/FrameStrobe[16] Tile_X5Y6_LUT4AB/FrameStrobe[17]
+ Tile_X5Y6_LUT4AB/FrameStrobe[18] Tile_X5Y6_LUT4AB/FrameStrobe[19] Tile_X5Y6_LUT4AB/FrameStrobe[1]
+ Tile_X5Y6_LUT4AB/FrameStrobe[2] Tile_X5Y6_LUT4AB/FrameStrobe[3] Tile_X5Y6_LUT4AB/FrameStrobe[4]
+ Tile_X5Y6_LUT4AB/FrameStrobe[5] Tile_X5Y6_LUT4AB/FrameStrobe[6] Tile_X5Y6_LUT4AB/FrameStrobe[7]
+ Tile_X5Y6_LUT4AB/FrameStrobe[8] Tile_X5Y6_LUT4AB/FrameStrobe[9] Tile_X5Y7_LUT4AB/N1BEG[0]
+ Tile_X5Y7_LUT4AB/N1BEG[1] Tile_X5Y7_LUT4AB/N1BEG[2] Tile_X5Y7_LUT4AB/N1BEG[3] Tile_X5Y8_LUT4AB/N1BEG[0]
+ Tile_X5Y8_LUT4AB/N1BEG[1] Tile_X5Y8_LUT4AB/N1BEG[2] Tile_X5Y8_LUT4AB/N1BEG[3] Tile_X5Y7_LUT4AB/N2BEG[0]
+ Tile_X5Y7_LUT4AB/N2BEG[1] Tile_X5Y7_LUT4AB/N2BEG[2] Tile_X5Y7_LUT4AB/N2BEG[3] Tile_X5Y7_LUT4AB/N2BEG[4]
+ Tile_X5Y7_LUT4AB/N2BEG[5] Tile_X5Y7_LUT4AB/N2BEG[6] Tile_X5Y7_LUT4AB/N2BEG[7] Tile_X5Y6_LUT4AB/N2END[0]
+ Tile_X5Y6_LUT4AB/N2END[1] Tile_X5Y6_LUT4AB/N2END[2] Tile_X5Y6_LUT4AB/N2END[3] Tile_X5Y6_LUT4AB/N2END[4]
+ Tile_X5Y6_LUT4AB/N2END[5] Tile_X5Y6_LUT4AB/N2END[6] Tile_X5Y6_LUT4AB/N2END[7] Tile_X5Y7_LUT4AB/N2END[0]
+ Tile_X5Y7_LUT4AB/N2END[1] Tile_X5Y7_LUT4AB/N2END[2] Tile_X5Y7_LUT4AB/N2END[3] Tile_X5Y7_LUT4AB/N2END[4]
+ Tile_X5Y7_LUT4AB/N2END[5] Tile_X5Y7_LUT4AB/N2END[6] Tile_X5Y7_LUT4AB/N2END[7] Tile_X5Y8_LUT4AB/N2BEG[0]
+ Tile_X5Y8_LUT4AB/N2BEG[1] Tile_X5Y8_LUT4AB/N2BEG[2] Tile_X5Y8_LUT4AB/N2BEG[3] Tile_X5Y8_LUT4AB/N2BEG[4]
+ Tile_X5Y8_LUT4AB/N2BEG[5] Tile_X5Y8_LUT4AB/N2BEG[6] Tile_X5Y8_LUT4AB/N2BEG[7] Tile_X5Y7_LUT4AB/N4BEG[0]
+ Tile_X5Y7_LUT4AB/N4BEG[10] Tile_X5Y7_LUT4AB/N4BEG[11] Tile_X5Y7_LUT4AB/N4BEG[12]
+ Tile_X5Y7_LUT4AB/N4BEG[13] Tile_X5Y7_LUT4AB/N4BEG[14] Tile_X5Y7_LUT4AB/N4BEG[15]
+ Tile_X5Y7_LUT4AB/N4BEG[1] Tile_X5Y7_LUT4AB/N4BEG[2] Tile_X5Y7_LUT4AB/N4BEG[3] Tile_X5Y7_LUT4AB/N4BEG[4]
+ Tile_X5Y7_LUT4AB/N4BEG[5] Tile_X5Y7_LUT4AB/N4BEG[6] Tile_X5Y7_LUT4AB/N4BEG[7] Tile_X5Y7_LUT4AB/N4BEG[8]
+ Tile_X5Y7_LUT4AB/N4BEG[9] Tile_X5Y8_LUT4AB/N4BEG[0] Tile_X5Y8_LUT4AB/N4BEG[10] Tile_X5Y8_LUT4AB/N4BEG[11]
+ Tile_X5Y8_LUT4AB/N4BEG[12] Tile_X5Y8_LUT4AB/N4BEG[13] Tile_X5Y8_LUT4AB/N4BEG[14]
+ Tile_X5Y8_LUT4AB/N4BEG[15] Tile_X5Y8_LUT4AB/N4BEG[1] Tile_X5Y8_LUT4AB/N4BEG[2] Tile_X5Y8_LUT4AB/N4BEG[3]
+ Tile_X5Y8_LUT4AB/N4BEG[4] Tile_X5Y8_LUT4AB/N4BEG[5] Tile_X5Y8_LUT4AB/N4BEG[6] Tile_X5Y8_LUT4AB/N4BEG[7]
+ Tile_X5Y8_LUT4AB/N4BEG[8] Tile_X5Y8_LUT4AB/N4BEG[9] Tile_X5Y7_LUT4AB/NN4BEG[0] Tile_X5Y7_LUT4AB/NN4BEG[10]
+ Tile_X5Y7_LUT4AB/NN4BEG[11] Tile_X5Y7_LUT4AB/NN4BEG[12] Tile_X5Y7_LUT4AB/NN4BEG[13]
+ Tile_X5Y7_LUT4AB/NN4BEG[14] Tile_X5Y7_LUT4AB/NN4BEG[15] Tile_X5Y7_LUT4AB/NN4BEG[1]
+ Tile_X5Y7_LUT4AB/NN4BEG[2] Tile_X5Y7_LUT4AB/NN4BEG[3] Tile_X5Y7_LUT4AB/NN4BEG[4]
+ Tile_X5Y7_LUT4AB/NN4BEG[5] Tile_X5Y7_LUT4AB/NN4BEG[6] Tile_X5Y7_LUT4AB/NN4BEG[7]
+ Tile_X5Y7_LUT4AB/NN4BEG[8] Tile_X5Y7_LUT4AB/NN4BEG[9] Tile_X5Y8_LUT4AB/NN4BEG[0]
+ Tile_X5Y8_LUT4AB/NN4BEG[10] Tile_X5Y8_LUT4AB/NN4BEG[11] Tile_X5Y8_LUT4AB/NN4BEG[12]
+ Tile_X5Y8_LUT4AB/NN4BEG[13] Tile_X5Y8_LUT4AB/NN4BEG[14] Tile_X5Y8_LUT4AB/NN4BEG[15]
+ Tile_X5Y8_LUT4AB/NN4BEG[1] Tile_X5Y8_LUT4AB/NN4BEG[2] Tile_X5Y8_LUT4AB/NN4BEG[3]
+ Tile_X5Y8_LUT4AB/NN4BEG[4] Tile_X5Y8_LUT4AB/NN4BEG[5] Tile_X5Y8_LUT4AB/NN4BEG[6]
+ Tile_X5Y8_LUT4AB/NN4BEG[7] Tile_X5Y8_LUT4AB/NN4BEG[8] Tile_X5Y8_LUT4AB/NN4BEG[9]
+ Tile_X5Y8_LUT4AB/S1END[0] Tile_X5Y8_LUT4AB/S1END[1] Tile_X5Y8_LUT4AB/S1END[2] Tile_X5Y8_LUT4AB/S1END[3]
+ Tile_X5Y7_LUT4AB/S1END[0] Tile_X5Y7_LUT4AB/S1END[1] Tile_X5Y7_LUT4AB/S1END[2] Tile_X5Y7_LUT4AB/S1END[3]
+ Tile_X5Y8_LUT4AB/S2MID[0] Tile_X5Y8_LUT4AB/S2MID[1] Tile_X5Y8_LUT4AB/S2MID[2] Tile_X5Y8_LUT4AB/S2MID[3]
+ Tile_X5Y8_LUT4AB/S2MID[4] Tile_X5Y8_LUT4AB/S2MID[5] Tile_X5Y8_LUT4AB/S2MID[6] Tile_X5Y8_LUT4AB/S2MID[7]
+ Tile_X5Y8_LUT4AB/S2END[0] Tile_X5Y8_LUT4AB/S2END[1] Tile_X5Y8_LUT4AB/S2END[2] Tile_X5Y8_LUT4AB/S2END[3]
+ Tile_X5Y8_LUT4AB/S2END[4] Tile_X5Y8_LUT4AB/S2END[5] Tile_X5Y8_LUT4AB/S2END[6] Tile_X5Y8_LUT4AB/S2END[7]
+ Tile_X5Y7_LUT4AB/S2END[0] Tile_X5Y7_LUT4AB/S2END[1] Tile_X5Y7_LUT4AB/S2END[2] Tile_X5Y7_LUT4AB/S2END[3]
+ Tile_X5Y7_LUT4AB/S2END[4] Tile_X5Y7_LUT4AB/S2END[5] Tile_X5Y7_LUT4AB/S2END[6] Tile_X5Y7_LUT4AB/S2END[7]
+ Tile_X5Y7_LUT4AB/S2MID[0] Tile_X5Y7_LUT4AB/S2MID[1] Tile_X5Y7_LUT4AB/S2MID[2] Tile_X5Y7_LUT4AB/S2MID[3]
+ Tile_X5Y7_LUT4AB/S2MID[4] Tile_X5Y7_LUT4AB/S2MID[5] Tile_X5Y7_LUT4AB/S2MID[6] Tile_X5Y7_LUT4AB/S2MID[7]
+ Tile_X5Y8_LUT4AB/S4END[0] Tile_X5Y8_LUT4AB/S4END[10] Tile_X5Y8_LUT4AB/S4END[11]
+ Tile_X5Y8_LUT4AB/S4END[12] Tile_X5Y8_LUT4AB/S4END[13] Tile_X5Y8_LUT4AB/S4END[14]
+ Tile_X5Y8_LUT4AB/S4END[15] Tile_X5Y8_LUT4AB/S4END[1] Tile_X5Y8_LUT4AB/S4END[2] Tile_X5Y8_LUT4AB/S4END[3]
+ Tile_X5Y8_LUT4AB/S4END[4] Tile_X5Y8_LUT4AB/S4END[5] Tile_X5Y8_LUT4AB/S4END[6] Tile_X5Y8_LUT4AB/S4END[7]
+ Tile_X5Y8_LUT4AB/S4END[8] Tile_X5Y8_LUT4AB/S4END[9] Tile_X5Y7_LUT4AB/S4END[0] Tile_X5Y7_LUT4AB/S4END[10]
+ Tile_X5Y7_LUT4AB/S4END[11] Tile_X5Y7_LUT4AB/S4END[12] Tile_X5Y7_LUT4AB/S4END[13]
+ Tile_X5Y7_LUT4AB/S4END[14] Tile_X5Y7_LUT4AB/S4END[15] Tile_X5Y7_LUT4AB/S4END[1]
+ Tile_X5Y7_LUT4AB/S4END[2] Tile_X5Y7_LUT4AB/S4END[3] Tile_X5Y7_LUT4AB/S4END[4] Tile_X5Y7_LUT4AB/S4END[5]
+ Tile_X5Y7_LUT4AB/S4END[6] Tile_X5Y7_LUT4AB/S4END[7] Tile_X5Y7_LUT4AB/S4END[8] Tile_X5Y7_LUT4AB/S4END[9]
+ Tile_X5Y8_LUT4AB/SS4END[0] Tile_X5Y8_LUT4AB/SS4END[10] Tile_X5Y8_LUT4AB/SS4END[11]
+ Tile_X5Y8_LUT4AB/SS4END[12] Tile_X5Y8_LUT4AB/SS4END[13] Tile_X5Y8_LUT4AB/SS4END[14]
+ Tile_X5Y8_LUT4AB/SS4END[15] Tile_X5Y8_LUT4AB/SS4END[1] Tile_X5Y8_LUT4AB/SS4END[2]
+ Tile_X5Y8_LUT4AB/SS4END[3] Tile_X5Y8_LUT4AB/SS4END[4] Tile_X5Y8_LUT4AB/SS4END[5]
+ Tile_X5Y8_LUT4AB/SS4END[6] Tile_X5Y8_LUT4AB/SS4END[7] Tile_X5Y8_LUT4AB/SS4END[8]
+ Tile_X5Y8_LUT4AB/SS4END[9] Tile_X5Y7_LUT4AB/SS4END[0] Tile_X5Y7_LUT4AB/SS4END[10]
+ Tile_X5Y7_LUT4AB/SS4END[11] Tile_X5Y7_LUT4AB/SS4END[12] Tile_X5Y7_LUT4AB/SS4END[13]
+ Tile_X5Y7_LUT4AB/SS4END[14] Tile_X5Y7_LUT4AB/SS4END[15] Tile_X5Y7_LUT4AB/SS4END[1]
+ Tile_X5Y7_LUT4AB/SS4END[2] Tile_X5Y7_LUT4AB/SS4END[3] Tile_X5Y7_LUT4AB/SS4END[4]
+ Tile_X5Y7_LUT4AB/SS4END[5] Tile_X5Y7_LUT4AB/SS4END[6] Tile_X5Y7_LUT4AB/SS4END[7]
+ Tile_X5Y7_LUT4AB/SS4END[8] Tile_X5Y7_LUT4AB/SS4END[9] Tile_X5Y7_LUT4AB/UserCLK Tile_X5Y6_LUT4AB/UserCLK
+ VGND VPWR Tile_X5Y7_LUT4AB/W1BEG[0] Tile_X5Y7_LUT4AB/W1BEG[1] Tile_X5Y7_LUT4AB/W1BEG[2]
+ Tile_X5Y7_LUT4AB/W1BEG[3] Tile_X6Y7_LUT4AB/W1BEG[0] Tile_X6Y7_LUT4AB/W1BEG[1] Tile_X6Y7_LUT4AB/W1BEG[2]
+ Tile_X6Y7_LUT4AB/W1BEG[3] Tile_X5Y7_LUT4AB/W2BEG[0] Tile_X5Y7_LUT4AB/W2BEG[1] Tile_X5Y7_LUT4AB/W2BEG[2]
+ Tile_X5Y7_LUT4AB/W2BEG[3] Tile_X5Y7_LUT4AB/W2BEG[4] Tile_X5Y7_LUT4AB/W2BEG[5] Tile_X5Y7_LUT4AB/W2BEG[6]
+ Tile_X5Y7_LUT4AB/W2BEG[7] Tile_X5Y7_LUT4AB/W2BEGb[0] Tile_X5Y7_LUT4AB/W2BEGb[1]
+ Tile_X5Y7_LUT4AB/W2BEGb[2] Tile_X5Y7_LUT4AB/W2BEGb[3] Tile_X5Y7_LUT4AB/W2BEGb[4]
+ Tile_X5Y7_LUT4AB/W2BEGb[5] Tile_X5Y7_LUT4AB/W2BEGb[6] Tile_X5Y7_LUT4AB/W2BEGb[7]
+ Tile_X5Y7_LUT4AB/W2END[0] Tile_X5Y7_LUT4AB/W2END[1] Tile_X5Y7_LUT4AB/W2END[2] Tile_X5Y7_LUT4AB/W2END[3]
+ Tile_X5Y7_LUT4AB/W2END[4] Tile_X5Y7_LUT4AB/W2END[5] Tile_X5Y7_LUT4AB/W2END[6] Tile_X5Y7_LUT4AB/W2END[7]
+ Tile_X6Y7_LUT4AB/W2BEG[0] Tile_X6Y7_LUT4AB/W2BEG[1] Tile_X6Y7_LUT4AB/W2BEG[2] Tile_X6Y7_LUT4AB/W2BEG[3]
+ Tile_X6Y7_LUT4AB/W2BEG[4] Tile_X6Y7_LUT4AB/W2BEG[5] Tile_X6Y7_LUT4AB/W2BEG[6] Tile_X6Y7_LUT4AB/W2BEG[7]
+ Tile_X5Y7_LUT4AB/W6BEG[0] Tile_X5Y7_LUT4AB/W6BEG[10] Tile_X5Y7_LUT4AB/W6BEG[11]
+ Tile_X5Y7_LUT4AB/W6BEG[1] Tile_X5Y7_LUT4AB/W6BEG[2] Tile_X5Y7_LUT4AB/W6BEG[3] Tile_X5Y7_LUT4AB/W6BEG[4]
+ Tile_X5Y7_LUT4AB/W6BEG[5] Tile_X5Y7_LUT4AB/W6BEG[6] Tile_X5Y7_LUT4AB/W6BEG[7] Tile_X5Y7_LUT4AB/W6BEG[8]
+ Tile_X5Y7_LUT4AB/W6BEG[9] Tile_X6Y7_LUT4AB/W6BEG[0] Tile_X6Y7_LUT4AB/W6BEG[10] Tile_X6Y7_LUT4AB/W6BEG[11]
+ Tile_X6Y7_LUT4AB/W6BEG[1] Tile_X6Y7_LUT4AB/W6BEG[2] Tile_X6Y7_LUT4AB/W6BEG[3] Tile_X6Y7_LUT4AB/W6BEG[4]
+ Tile_X6Y7_LUT4AB/W6BEG[5] Tile_X6Y7_LUT4AB/W6BEG[6] Tile_X6Y7_LUT4AB/W6BEG[7] Tile_X6Y7_LUT4AB/W6BEG[8]
+ Tile_X6Y7_LUT4AB/W6BEG[9] Tile_X5Y7_LUT4AB/WW4BEG[0] Tile_X5Y7_LUT4AB/WW4BEG[10]
+ Tile_X5Y7_LUT4AB/WW4BEG[11] Tile_X5Y7_LUT4AB/WW4BEG[12] Tile_X5Y7_LUT4AB/WW4BEG[13]
+ Tile_X5Y7_LUT4AB/WW4BEG[14] Tile_X5Y7_LUT4AB/WW4BEG[15] Tile_X5Y7_LUT4AB/WW4BEG[1]
+ Tile_X5Y7_LUT4AB/WW4BEG[2] Tile_X5Y7_LUT4AB/WW4BEG[3] Tile_X5Y7_LUT4AB/WW4BEG[4]
+ Tile_X5Y7_LUT4AB/WW4BEG[5] Tile_X5Y7_LUT4AB/WW4BEG[6] Tile_X5Y7_LUT4AB/WW4BEG[7]
+ Tile_X5Y7_LUT4AB/WW4BEG[8] Tile_X5Y7_LUT4AB/WW4BEG[9] Tile_X6Y7_LUT4AB/WW4BEG[0]
+ Tile_X6Y7_LUT4AB/WW4BEG[10] Tile_X6Y7_LUT4AB/WW4BEG[11] Tile_X6Y7_LUT4AB/WW4BEG[12]
+ Tile_X6Y7_LUT4AB/WW4BEG[13] Tile_X6Y7_LUT4AB/WW4BEG[14] Tile_X6Y7_LUT4AB/WW4BEG[15]
+ Tile_X6Y7_LUT4AB/WW4BEG[1] Tile_X6Y7_LUT4AB/WW4BEG[2] Tile_X6Y7_LUT4AB/WW4BEG[3]
+ Tile_X6Y7_LUT4AB/WW4BEG[4] Tile_X6Y7_LUT4AB/WW4BEG[5] Tile_X6Y7_LUT4AB/WW4BEG[6]
+ Tile_X6Y7_LUT4AB/WW4BEG[7] Tile_X6Y7_LUT4AB/WW4BEG[8] Tile_X6Y7_LUT4AB/WW4BEG[9]
+ LUT4AB
XTile_X1Y6_LUT4AB Tile_X1Y7_LUT4AB/Co Tile_X1Y6_LUT4AB/Co Tile_X2Y6_LUT4AB/E1END[0]
+ Tile_X2Y6_LUT4AB/E1END[1] Tile_X2Y6_LUT4AB/E1END[2] Tile_X2Y6_LUT4AB/E1END[3] Tile_X0Y6_W_IO/E1BEG[0]
+ Tile_X0Y6_W_IO/E1BEG[1] Tile_X0Y6_W_IO/E1BEG[2] Tile_X0Y6_W_IO/E1BEG[3] Tile_X2Y6_LUT4AB/E2MID[0]
+ Tile_X2Y6_LUT4AB/E2MID[1] Tile_X2Y6_LUT4AB/E2MID[2] Tile_X2Y6_LUT4AB/E2MID[3] Tile_X2Y6_LUT4AB/E2MID[4]
+ Tile_X2Y6_LUT4AB/E2MID[5] Tile_X2Y6_LUT4AB/E2MID[6] Tile_X2Y6_LUT4AB/E2MID[7] Tile_X2Y6_LUT4AB/E2END[0]
+ Tile_X2Y6_LUT4AB/E2END[1] Tile_X2Y6_LUT4AB/E2END[2] Tile_X2Y6_LUT4AB/E2END[3] Tile_X2Y6_LUT4AB/E2END[4]
+ Tile_X2Y6_LUT4AB/E2END[5] Tile_X2Y6_LUT4AB/E2END[6] Tile_X2Y6_LUT4AB/E2END[7] Tile_X0Y6_W_IO/E2BEGb[0]
+ Tile_X0Y6_W_IO/E2BEGb[1] Tile_X0Y6_W_IO/E2BEGb[2] Tile_X0Y6_W_IO/E2BEGb[3] Tile_X0Y6_W_IO/E2BEGb[4]
+ Tile_X0Y6_W_IO/E2BEGb[5] Tile_X0Y6_W_IO/E2BEGb[6] Tile_X0Y6_W_IO/E2BEGb[7] Tile_X0Y6_W_IO/E2BEG[0]
+ Tile_X0Y6_W_IO/E2BEG[1] Tile_X0Y6_W_IO/E2BEG[2] Tile_X0Y6_W_IO/E2BEG[3] Tile_X0Y6_W_IO/E2BEG[4]
+ Tile_X0Y6_W_IO/E2BEG[5] Tile_X0Y6_W_IO/E2BEG[6] Tile_X0Y6_W_IO/E2BEG[7] Tile_X2Y6_LUT4AB/E6END[0]
+ Tile_X2Y6_LUT4AB/E6END[10] Tile_X2Y6_LUT4AB/E6END[11] Tile_X2Y6_LUT4AB/E6END[1]
+ Tile_X2Y6_LUT4AB/E6END[2] Tile_X2Y6_LUT4AB/E6END[3] Tile_X2Y6_LUT4AB/E6END[4] Tile_X2Y6_LUT4AB/E6END[5]
+ Tile_X2Y6_LUT4AB/E6END[6] Tile_X2Y6_LUT4AB/E6END[7] Tile_X2Y6_LUT4AB/E6END[8] Tile_X2Y6_LUT4AB/E6END[9]
+ Tile_X0Y6_W_IO/E6BEG[0] Tile_X0Y6_W_IO/E6BEG[10] Tile_X0Y6_W_IO/E6BEG[11] Tile_X0Y6_W_IO/E6BEG[1]
+ Tile_X0Y6_W_IO/E6BEG[2] Tile_X0Y6_W_IO/E6BEG[3] Tile_X0Y6_W_IO/E6BEG[4] Tile_X0Y6_W_IO/E6BEG[5]
+ Tile_X0Y6_W_IO/E6BEG[6] Tile_X0Y6_W_IO/E6BEG[7] Tile_X0Y6_W_IO/E6BEG[8] Tile_X0Y6_W_IO/E6BEG[9]
+ Tile_X2Y6_LUT4AB/EE4END[0] Tile_X2Y6_LUT4AB/EE4END[10] Tile_X2Y6_LUT4AB/EE4END[11]
+ Tile_X2Y6_LUT4AB/EE4END[12] Tile_X2Y6_LUT4AB/EE4END[13] Tile_X2Y6_LUT4AB/EE4END[14]
+ Tile_X2Y6_LUT4AB/EE4END[15] Tile_X2Y6_LUT4AB/EE4END[1] Tile_X2Y6_LUT4AB/EE4END[2]
+ Tile_X2Y6_LUT4AB/EE4END[3] Tile_X2Y6_LUT4AB/EE4END[4] Tile_X2Y6_LUT4AB/EE4END[5]
+ Tile_X2Y6_LUT4AB/EE4END[6] Tile_X2Y6_LUT4AB/EE4END[7] Tile_X2Y6_LUT4AB/EE4END[8]
+ Tile_X2Y6_LUT4AB/EE4END[9] Tile_X0Y6_W_IO/EE4BEG[0] Tile_X0Y6_W_IO/EE4BEG[10] Tile_X0Y6_W_IO/EE4BEG[11]
+ Tile_X0Y6_W_IO/EE4BEG[12] Tile_X0Y6_W_IO/EE4BEG[13] Tile_X0Y6_W_IO/EE4BEG[14] Tile_X0Y6_W_IO/EE4BEG[15]
+ Tile_X0Y6_W_IO/EE4BEG[1] Tile_X0Y6_W_IO/EE4BEG[2] Tile_X0Y6_W_IO/EE4BEG[3] Tile_X0Y6_W_IO/EE4BEG[4]
+ Tile_X0Y6_W_IO/EE4BEG[5] Tile_X0Y6_W_IO/EE4BEG[6] Tile_X0Y6_W_IO/EE4BEG[7] Tile_X0Y6_W_IO/EE4BEG[8]
+ Tile_X0Y6_W_IO/EE4BEG[9] Tile_X1Y6_LUT4AB/FrameData[0] Tile_X1Y6_LUT4AB/FrameData[10]
+ Tile_X1Y6_LUT4AB/FrameData[11] Tile_X1Y6_LUT4AB/FrameData[12] Tile_X1Y6_LUT4AB/FrameData[13]
+ Tile_X1Y6_LUT4AB/FrameData[14] Tile_X1Y6_LUT4AB/FrameData[15] Tile_X1Y6_LUT4AB/FrameData[16]
+ Tile_X1Y6_LUT4AB/FrameData[17] Tile_X1Y6_LUT4AB/FrameData[18] Tile_X1Y6_LUT4AB/FrameData[19]
+ Tile_X1Y6_LUT4AB/FrameData[1] Tile_X1Y6_LUT4AB/FrameData[20] Tile_X1Y6_LUT4AB/FrameData[21]
+ Tile_X1Y6_LUT4AB/FrameData[22] Tile_X1Y6_LUT4AB/FrameData[23] Tile_X1Y6_LUT4AB/FrameData[24]
+ Tile_X1Y6_LUT4AB/FrameData[25] Tile_X1Y6_LUT4AB/FrameData[26] Tile_X1Y6_LUT4AB/FrameData[27]
+ Tile_X1Y6_LUT4AB/FrameData[28] Tile_X1Y6_LUT4AB/FrameData[29] Tile_X1Y6_LUT4AB/FrameData[2]
+ Tile_X1Y6_LUT4AB/FrameData[30] Tile_X1Y6_LUT4AB/FrameData[31] Tile_X1Y6_LUT4AB/FrameData[3]
+ Tile_X1Y6_LUT4AB/FrameData[4] Tile_X1Y6_LUT4AB/FrameData[5] Tile_X1Y6_LUT4AB/FrameData[6]
+ Tile_X1Y6_LUT4AB/FrameData[7] Tile_X1Y6_LUT4AB/FrameData[8] Tile_X1Y6_LUT4AB/FrameData[9]
+ Tile_X2Y6_LUT4AB/FrameData[0] Tile_X2Y6_LUT4AB/FrameData[10] Tile_X2Y6_LUT4AB/FrameData[11]
+ Tile_X2Y6_LUT4AB/FrameData[12] Tile_X2Y6_LUT4AB/FrameData[13] Tile_X2Y6_LUT4AB/FrameData[14]
+ Tile_X2Y6_LUT4AB/FrameData[15] Tile_X2Y6_LUT4AB/FrameData[16] Tile_X2Y6_LUT4AB/FrameData[17]
+ Tile_X2Y6_LUT4AB/FrameData[18] Tile_X2Y6_LUT4AB/FrameData[19] Tile_X2Y6_LUT4AB/FrameData[1]
+ Tile_X2Y6_LUT4AB/FrameData[20] Tile_X2Y6_LUT4AB/FrameData[21] Tile_X2Y6_LUT4AB/FrameData[22]
+ Tile_X2Y6_LUT4AB/FrameData[23] Tile_X2Y6_LUT4AB/FrameData[24] Tile_X2Y6_LUT4AB/FrameData[25]
+ Tile_X2Y6_LUT4AB/FrameData[26] Tile_X2Y6_LUT4AB/FrameData[27] Tile_X2Y6_LUT4AB/FrameData[28]
+ Tile_X2Y6_LUT4AB/FrameData[29] Tile_X2Y6_LUT4AB/FrameData[2] Tile_X2Y6_LUT4AB/FrameData[30]
+ Tile_X2Y6_LUT4AB/FrameData[31] Tile_X2Y6_LUT4AB/FrameData[3] Tile_X2Y6_LUT4AB/FrameData[4]
+ Tile_X2Y6_LUT4AB/FrameData[5] Tile_X2Y6_LUT4AB/FrameData[6] Tile_X2Y6_LUT4AB/FrameData[7]
+ Tile_X2Y6_LUT4AB/FrameData[8] Tile_X2Y6_LUT4AB/FrameData[9] Tile_X1Y6_LUT4AB/FrameStrobe[0]
+ Tile_X1Y6_LUT4AB/FrameStrobe[10] Tile_X1Y6_LUT4AB/FrameStrobe[11] Tile_X1Y6_LUT4AB/FrameStrobe[12]
+ Tile_X1Y6_LUT4AB/FrameStrobe[13] Tile_X1Y6_LUT4AB/FrameStrobe[14] Tile_X1Y6_LUT4AB/FrameStrobe[15]
+ Tile_X1Y6_LUT4AB/FrameStrobe[16] Tile_X1Y6_LUT4AB/FrameStrobe[17] Tile_X1Y6_LUT4AB/FrameStrobe[18]
+ Tile_X1Y6_LUT4AB/FrameStrobe[19] Tile_X1Y6_LUT4AB/FrameStrobe[1] Tile_X1Y6_LUT4AB/FrameStrobe[2]
+ Tile_X1Y6_LUT4AB/FrameStrobe[3] Tile_X1Y6_LUT4AB/FrameStrobe[4] Tile_X1Y6_LUT4AB/FrameStrobe[5]
+ Tile_X1Y6_LUT4AB/FrameStrobe[6] Tile_X1Y6_LUT4AB/FrameStrobe[7] Tile_X1Y6_LUT4AB/FrameStrobe[8]
+ Tile_X1Y6_LUT4AB/FrameStrobe[9] Tile_X1Y5_LUT4AB/FrameStrobe[0] Tile_X1Y5_LUT4AB/FrameStrobe[10]
+ Tile_X1Y5_LUT4AB/FrameStrobe[11] Tile_X1Y5_LUT4AB/FrameStrobe[12] Tile_X1Y5_LUT4AB/FrameStrobe[13]
+ Tile_X1Y5_LUT4AB/FrameStrobe[14] Tile_X1Y5_LUT4AB/FrameStrobe[15] Tile_X1Y5_LUT4AB/FrameStrobe[16]
+ Tile_X1Y5_LUT4AB/FrameStrobe[17] Tile_X1Y5_LUT4AB/FrameStrobe[18] Tile_X1Y5_LUT4AB/FrameStrobe[19]
+ Tile_X1Y5_LUT4AB/FrameStrobe[1] Tile_X1Y5_LUT4AB/FrameStrobe[2] Tile_X1Y5_LUT4AB/FrameStrobe[3]
+ Tile_X1Y5_LUT4AB/FrameStrobe[4] Tile_X1Y5_LUT4AB/FrameStrobe[5] Tile_X1Y5_LUT4AB/FrameStrobe[6]
+ Tile_X1Y5_LUT4AB/FrameStrobe[7] Tile_X1Y5_LUT4AB/FrameStrobe[8] Tile_X1Y5_LUT4AB/FrameStrobe[9]
+ Tile_X1Y6_LUT4AB/N1BEG[0] Tile_X1Y6_LUT4AB/N1BEG[1] Tile_X1Y6_LUT4AB/N1BEG[2] Tile_X1Y6_LUT4AB/N1BEG[3]
+ Tile_X1Y7_LUT4AB/N1BEG[0] Tile_X1Y7_LUT4AB/N1BEG[1] Tile_X1Y7_LUT4AB/N1BEG[2] Tile_X1Y7_LUT4AB/N1BEG[3]
+ Tile_X1Y6_LUT4AB/N2BEG[0] Tile_X1Y6_LUT4AB/N2BEG[1] Tile_X1Y6_LUT4AB/N2BEG[2] Tile_X1Y6_LUT4AB/N2BEG[3]
+ Tile_X1Y6_LUT4AB/N2BEG[4] Tile_X1Y6_LUT4AB/N2BEG[5] Tile_X1Y6_LUT4AB/N2BEG[6] Tile_X1Y6_LUT4AB/N2BEG[7]
+ Tile_X1Y5_LUT4AB/N2END[0] Tile_X1Y5_LUT4AB/N2END[1] Tile_X1Y5_LUT4AB/N2END[2] Tile_X1Y5_LUT4AB/N2END[3]
+ Tile_X1Y5_LUT4AB/N2END[4] Tile_X1Y5_LUT4AB/N2END[5] Tile_X1Y5_LUT4AB/N2END[6] Tile_X1Y5_LUT4AB/N2END[7]
+ Tile_X1Y6_LUT4AB/N2END[0] Tile_X1Y6_LUT4AB/N2END[1] Tile_X1Y6_LUT4AB/N2END[2] Tile_X1Y6_LUT4AB/N2END[3]
+ Tile_X1Y6_LUT4AB/N2END[4] Tile_X1Y6_LUT4AB/N2END[5] Tile_X1Y6_LUT4AB/N2END[6] Tile_X1Y6_LUT4AB/N2END[7]
+ Tile_X1Y7_LUT4AB/N2BEG[0] Tile_X1Y7_LUT4AB/N2BEG[1] Tile_X1Y7_LUT4AB/N2BEG[2] Tile_X1Y7_LUT4AB/N2BEG[3]
+ Tile_X1Y7_LUT4AB/N2BEG[4] Tile_X1Y7_LUT4AB/N2BEG[5] Tile_X1Y7_LUT4AB/N2BEG[6] Tile_X1Y7_LUT4AB/N2BEG[7]
+ Tile_X1Y6_LUT4AB/N4BEG[0] Tile_X1Y6_LUT4AB/N4BEG[10] Tile_X1Y6_LUT4AB/N4BEG[11]
+ Tile_X1Y6_LUT4AB/N4BEG[12] Tile_X1Y6_LUT4AB/N4BEG[13] Tile_X1Y6_LUT4AB/N4BEG[14]
+ Tile_X1Y6_LUT4AB/N4BEG[15] Tile_X1Y6_LUT4AB/N4BEG[1] Tile_X1Y6_LUT4AB/N4BEG[2] Tile_X1Y6_LUT4AB/N4BEG[3]
+ Tile_X1Y6_LUT4AB/N4BEG[4] Tile_X1Y6_LUT4AB/N4BEG[5] Tile_X1Y6_LUT4AB/N4BEG[6] Tile_X1Y6_LUT4AB/N4BEG[7]
+ Tile_X1Y6_LUT4AB/N4BEG[8] Tile_X1Y6_LUT4AB/N4BEG[9] Tile_X1Y7_LUT4AB/N4BEG[0] Tile_X1Y7_LUT4AB/N4BEG[10]
+ Tile_X1Y7_LUT4AB/N4BEG[11] Tile_X1Y7_LUT4AB/N4BEG[12] Tile_X1Y7_LUT4AB/N4BEG[13]
+ Tile_X1Y7_LUT4AB/N4BEG[14] Tile_X1Y7_LUT4AB/N4BEG[15] Tile_X1Y7_LUT4AB/N4BEG[1]
+ Tile_X1Y7_LUT4AB/N4BEG[2] Tile_X1Y7_LUT4AB/N4BEG[3] Tile_X1Y7_LUT4AB/N4BEG[4] Tile_X1Y7_LUT4AB/N4BEG[5]
+ Tile_X1Y7_LUT4AB/N4BEG[6] Tile_X1Y7_LUT4AB/N4BEG[7] Tile_X1Y7_LUT4AB/N4BEG[8] Tile_X1Y7_LUT4AB/N4BEG[9]
+ Tile_X1Y6_LUT4AB/NN4BEG[0] Tile_X1Y6_LUT4AB/NN4BEG[10] Tile_X1Y6_LUT4AB/NN4BEG[11]
+ Tile_X1Y6_LUT4AB/NN4BEG[12] Tile_X1Y6_LUT4AB/NN4BEG[13] Tile_X1Y6_LUT4AB/NN4BEG[14]
+ Tile_X1Y6_LUT4AB/NN4BEG[15] Tile_X1Y6_LUT4AB/NN4BEG[1] Tile_X1Y6_LUT4AB/NN4BEG[2]
+ Tile_X1Y6_LUT4AB/NN4BEG[3] Tile_X1Y6_LUT4AB/NN4BEG[4] Tile_X1Y6_LUT4AB/NN4BEG[5]
+ Tile_X1Y6_LUT4AB/NN4BEG[6] Tile_X1Y6_LUT4AB/NN4BEG[7] Tile_X1Y6_LUT4AB/NN4BEG[8]
+ Tile_X1Y6_LUT4AB/NN4BEG[9] Tile_X1Y7_LUT4AB/NN4BEG[0] Tile_X1Y7_LUT4AB/NN4BEG[10]
+ Tile_X1Y7_LUT4AB/NN4BEG[11] Tile_X1Y7_LUT4AB/NN4BEG[12] Tile_X1Y7_LUT4AB/NN4BEG[13]
+ Tile_X1Y7_LUT4AB/NN4BEG[14] Tile_X1Y7_LUT4AB/NN4BEG[15] Tile_X1Y7_LUT4AB/NN4BEG[1]
+ Tile_X1Y7_LUT4AB/NN4BEG[2] Tile_X1Y7_LUT4AB/NN4BEG[3] Tile_X1Y7_LUT4AB/NN4BEG[4]
+ Tile_X1Y7_LUT4AB/NN4BEG[5] Tile_X1Y7_LUT4AB/NN4BEG[6] Tile_X1Y7_LUT4AB/NN4BEG[7]
+ Tile_X1Y7_LUT4AB/NN4BEG[8] Tile_X1Y7_LUT4AB/NN4BEG[9] Tile_X1Y7_LUT4AB/S1END[0]
+ Tile_X1Y7_LUT4AB/S1END[1] Tile_X1Y7_LUT4AB/S1END[2] Tile_X1Y7_LUT4AB/S1END[3] Tile_X1Y6_LUT4AB/S1END[0]
+ Tile_X1Y6_LUT4AB/S1END[1] Tile_X1Y6_LUT4AB/S1END[2] Tile_X1Y6_LUT4AB/S1END[3] Tile_X1Y7_LUT4AB/S2MID[0]
+ Tile_X1Y7_LUT4AB/S2MID[1] Tile_X1Y7_LUT4AB/S2MID[2] Tile_X1Y7_LUT4AB/S2MID[3] Tile_X1Y7_LUT4AB/S2MID[4]
+ Tile_X1Y7_LUT4AB/S2MID[5] Tile_X1Y7_LUT4AB/S2MID[6] Tile_X1Y7_LUT4AB/S2MID[7] Tile_X1Y7_LUT4AB/S2END[0]
+ Tile_X1Y7_LUT4AB/S2END[1] Tile_X1Y7_LUT4AB/S2END[2] Tile_X1Y7_LUT4AB/S2END[3] Tile_X1Y7_LUT4AB/S2END[4]
+ Tile_X1Y7_LUT4AB/S2END[5] Tile_X1Y7_LUT4AB/S2END[6] Tile_X1Y7_LUT4AB/S2END[7] Tile_X1Y6_LUT4AB/S2END[0]
+ Tile_X1Y6_LUT4AB/S2END[1] Tile_X1Y6_LUT4AB/S2END[2] Tile_X1Y6_LUT4AB/S2END[3] Tile_X1Y6_LUT4AB/S2END[4]
+ Tile_X1Y6_LUT4AB/S2END[5] Tile_X1Y6_LUT4AB/S2END[6] Tile_X1Y6_LUT4AB/S2END[7] Tile_X1Y6_LUT4AB/S2MID[0]
+ Tile_X1Y6_LUT4AB/S2MID[1] Tile_X1Y6_LUT4AB/S2MID[2] Tile_X1Y6_LUT4AB/S2MID[3] Tile_X1Y6_LUT4AB/S2MID[4]
+ Tile_X1Y6_LUT4AB/S2MID[5] Tile_X1Y6_LUT4AB/S2MID[6] Tile_X1Y6_LUT4AB/S2MID[7] Tile_X1Y7_LUT4AB/S4END[0]
+ Tile_X1Y7_LUT4AB/S4END[10] Tile_X1Y7_LUT4AB/S4END[11] Tile_X1Y7_LUT4AB/S4END[12]
+ Tile_X1Y7_LUT4AB/S4END[13] Tile_X1Y7_LUT4AB/S4END[14] Tile_X1Y7_LUT4AB/S4END[15]
+ Tile_X1Y7_LUT4AB/S4END[1] Tile_X1Y7_LUT4AB/S4END[2] Tile_X1Y7_LUT4AB/S4END[3] Tile_X1Y7_LUT4AB/S4END[4]
+ Tile_X1Y7_LUT4AB/S4END[5] Tile_X1Y7_LUT4AB/S4END[6] Tile_X1Y7_LUT4AB/S4END[7] Tile_X1Y7_LUT4AB/S4END[8]
+ Tile_X1Y7_LUT4AB/S4END[9] Tile_X1Y6_LUT4AB/S4END[0] Tile_X1Y6_LUT4AB/S4END[10] Tile_X1Y6_LUT4AB/S4END[11]
+ Tile_X1Y6_LUT4AB/S4END[12] Tile_X1Y6_LUT4AB/S4END[13] Tile_X1Y6_LUT4AB/S4END[14]
+ Tile_X1Y6_LUT4AB/S4END[15] Tile_X1Y6_LUT4AB/S4END[1] Tile_X1Y6_LUT4AB/S4END[2] Tile_X1Y6_LUT4AB/S4END[3]
+ Tile_X1Y6_LUT4AB/S4END[4] Tile_X1Y6_LUT4AB/S4END[5] Tile_X1Y6_LUT4AB/S4END[6] Tile_X1Y6_LUT4AB/S4END[7]
+ Tile_X1Y6_LUT4AB/S4END[8] Tile_X1Y6_LUT4AB/S4END[9] Tile_X1Y7_LUT4AB/SS4END[0] Tile_X1Y7_LUT4AB/SS4END[10]
+ Tile_X1Y7_LUT4AB/SS4END[11] Tile_X1Y7_LUT4AB/SS4END[12] Tile_X1Y7_LUT4AB/SS4END[13]
+ Tile_X1Y7_LUT4AB/SS4END[14] Tile_X1Y7_LUT4AB/SS4END[15] Tile_X1Y7_LUT4AB/SS4END[1]
+ Tile_X1Y7_LUT4AB/SS4END[2] Tile_X1Y7_LUT4AB/SS4END[3] Tile_X1Y7_LUT4AB/SS4END[4]
+ Tile_X1Y7_LUT4AB/SS4END[5] Tile_X1Y7_LUT4AB/SS4END[6] Tile_X1Y7_LUT4AB/SS4END[7]
+ Tile_X1Y7_LUT4AB/SS4END[8] Tile_X1Y7_LUT4AB/SS4END[9] Tile_X1Y6_LUT4AB/SS4END[0]
+ Tile_X1Y6_LUT4AB/SS4END[10] Tile_X1Y6_LUT4AB/SS4END[11] Tile_X1Y6_LUT4AB/SS4END[12]
+ Tile_X1Y6_LUT4AB/SS4END[13] Tile_X1Y6_LUT4AB/SS4END[14] Tile_X1Y6_LUT4AB/SS4END[15]
+ Tile_X1Y6_LUT4AB/SS4END[1] Tile_X1Y6_LUT4AB/SS4END[2] Tile_X1Y6_LUT4AB/SS4END[3]
+ Tile_X1Y6_LUT4AB/SS4END[4] Tile_X1Y6_LUT4AB/SS4END[5] Tile_X1Y6_LUT4AB/SS4END[6]
+ Tile_X1Y6_LUT4AB/SS4END[7] Tile_X1Y6_LUT4AB/SS4END[8] Tile_X1Y6_LUT4AB/SS4END[9]
+ Tile_X1Y6_LUT4AB/UserCLK Tile_X1Y5_LUT4AB/UserCLK VGND VPWR Tile_X0Y6_W_IO/W1END[0]
+ Tile_X0Y6_W_IO/W1END[1] Tile_X0Y6_W_IO/W1END[2] Tile_X0Y6_W_IO/W1END[3] Tile_X2Y6_LUT4AB/W1BEG[0]
+ Tile_X2Y6_LUT4AB/W1BEG[1] Tile_X2Y6_LUT4AB/W1BEG[2] Tile_X2Y6_LUT4AB/W1BEG[3] Tile_X0Y6_W_IO/W2MID[0]
+ Tile_X0Y6_W_IO/W2MID[1] Tile_X0Y6_W_IO/W2MID[2] Tile_X0Y6_W_IO/W2MID[3] Tile_X0Y6_W_IO/W2MID[4]
+ Tile_X0Y6_W_IO/W2MID[5] Tile_X0Y6_W_IO/W2MID[6] Tile_X0Y6_W_IO/W2MID[7] Tile_X0Y6_W_IO/W2END[0]
+ Tile_X0Y6_W_IO/W2END[1] Tile_X0Y6_W_IO/W2END[2] Tile_X0Y6_W_IO/W2END[3] Tile_X0Y6_W_IO/W2END[4]
+ Tile_X0Y6_W_IO/W2END[5] Tile_X0Y6_W_IO/W2END[6] Tile_X0Y6_W_IO/W2END[7] Tile_X1Y6_LUT4AB/W2END[0]
+ Tile_X1Y6_LUT4AB/W2END[1] Tile_X1Y6_LUT4AB/W2END[2] Tile_X1Y6_LUT4AB/W2END[3] Tile_X1Y6_LUT4AB/W2END[4]
+ Tile_X1Y6_LUT4AB/W2END[5] Tile_X1Y6_LUT4AB/W2END[6] Tile_X1Y6_LUT4AB/W2END[7] Tile_X2Y6_LUT4AB/W2BEG[0]
+ Tile_X2Y6_LUT4AB/W2BEG[1] Tile_X2Y6_LUT4AB/W2BEG[2] Tile_X2Y6_LUT4AB/W2BEG[3] Tile_X2Y6_LUT4AB/W2BEG[4]
+ Tile_X2Y6_LUT4AB/W2BEG[5] Tile_X2Y6_LUT4AB/W2BEG[6] Tile_X2Y6_LUT4AB/W2BEG[7] Tile_X0Y6_W_IO/W6END[0]
+ Tile_X0Y6_W_IO/W6END[10] Tile_X0Y6_W_IO/W6END[11] Tile_X0Y6_W_IO/W6END[1] Tile_X0Y6_W_IO/W6END[2]
+ Tile_X0Y6_W_IO/W6END[3] Tile_X0Y6_W_IO/W6END[4] Tile_X0Y6_W_IO/W6END[5] Tile_X0Y6_W_IO/W6END[6]
+ Tile_X0Y6_W_IO/W6END[7] Tile_X0Y6_W_IO/W6END[8] Tile_X0Y6_W_IO/W6END[9] Tile_X2Y6_LUT4AB/W6BEG[0]
+ Tile_X2Y6_LUT4AB/W6BEG[10] Tile_X2Y6_LUT4AB/W6BEG[11] Tile_X2Y6_LUT4AB/W6BEG[1]
+ Tile_X2Y6_LUT4AB/W6BEG[2] Tile_X2Y6_LUT4AB/W6BEG[3] Tile_X2Y6_LUT4AB/W6BEG[4] Tile_X2Y6_LUT4AB/W6BEG[5]
+ Tile_X2Y6_LUT4AB/W6BEG[6] Tile_X2Y6_LUT4AB/W6BEG[7] Tile_X2Y6_LUT4AB/W6BEG[8] Tile_X2Y6_LUT4AB/W6BEG[9]
+ Tile_X0Y6_W_IO/WW4END[0] Tile_X0Y6_W_IO/WW4END[10] Tile_X0Y6_W_IO/WW4END[11] Tile_X0Y6_W_IO/WW4END[12]
+ Tile_X0Y6_W_IO/WW4END[13] Tile_X0Y6_W_IO/WW4END[14] Tile_X0Y6_W_IO/WW4END[15] Tile_X0Y6_W_IO/WW4END[1]
+ Tile_X0Y6_W_IO/WW4END[2] Tile_X0Y6_W_IO/WW4END[3] Tile_X0Y6_W_IO/WW4END[4] Tile_X0Y6_W_IO/WW4END[5]
+ Tile_X0Y6_W_IO/WW4END[6] Tile_X0Y6_W_IO/WW4END[7] Tile_X0Y6_W_IO/WW4END[8] Tile_X0Y6_W_IO/WW4END[9]
+ Tile_X2Y6_LUT4AB/WW4BEG[0] Tile_X2Y6_LUT4AB/WW4BEG[10] Tile_X2Y6_LUT4AB/WW4BEG[11]
+ Tile_X2Y6_LUT4AB/WW4BEG[12] Tile_X2Y6_LUT4AB/WW4BEG[13] Tile_X2Y6_LUT4AB/WW4BEG[14]
+ Tile_X2Y6_LUT4AB/WW4BEG[15] Tile_X2Y6_LUT4AB/WW4BEG[1] Tile_X2Y6_LUT4AB/WW4BEG[2]
+ Tile_X2Y6_LUT4AB/WW4BEG[3] Tile_X2Y6_LUT4AB/WW4BEG[4] Tile_X2Y6_LUT4AB/WW4BEG[5]
+ Tile_X2Y6_LUT4AB/WW4BEG[6] Tile_X2Y6_LUT4AB/WW4BEG[7] Tile_X2Y6_LUT4AB/WW4BEG[8]
+ Tile_X2Y6_LUT4AB/WW4BEG[9] LUT4AB
XTile_X8Y1_LUT4AB Tile_X8Y2_LUT4AB/Co Tile_X8Y1_LUT4AB/Co Tile_X9Y1_LUT4AB/E1END[0]
+ Tile_X9Y1_LUT4AB/E1END[1] Tile_X9Y1_LUT4AB/E1END[2] Tile_X9Y1_LUT4AB/E1END[3] Tile_X8Y1_LUT4AB/E1END[0]
+ Tile_X8Y1_LUT4AB/E1END[1] Tile_X8Y1_LUT4AB/E1END[2] Tile_X8Y1_LUT4AB/E1END[3] Tile_X9Y1_LUT4AB/E2MID[0]
+ Tile_X9Y1_LUT4AB/E2MID[1] Tile_X9Y1_LUT4AB/E2MID[2] Tile_X9Y1_LUT4AB/E2MID[3] Tile_X9Y1_LUT4AB/E2MID[4]
+ Tile_X9Y1_LUT4AB/E2MID[5] Tile_X9Y1_LUT4AB/E2MID[6] Tile_X9Y1_LUT4AB/E2MID[7] Tile_X9Y1_LUT4AB/E2END[0]
+ Tile_X9Y1_LUT4AB/E2END[1] Tile_X9Y1_LUT4AB/E2END[2] Tile_X9Y1_LUT4AB/E2END[3] Tile_X9Y1_LUT4AB/E2END[4]
+ Tile_X9Y1_LUT4AB/E2END[5] Tile_X9Y1_LUT4AB/E2END[6] Tile_X9Y1_LUT4AB/E2END[7] Tile_X8Y1_LUT4AB/E2END[0]
+ Tile_X8Y1_LUT4AB/E2END[1] Tile_X8Y1_LUT4AB/E2END[2] Tile_X8Y1_LUT4AB/E2END[3] Tile_X8Y1_LUT4AB/E2END[4]
+ Tile_X8Y1_LUT4AB/E2END[5] Tile_X8Y1_LUT4AB/E2END[6] Tile_X8Y1_LUT4AB/E2END[7] Tile_X8Y1_LUT4AB/E2MID[0]
+ Tile_X8Y1_LUT4AB/E2MID[1] Tile_X8Y1_LUT4AB/E2MID[2] Tile_X8Y1_LUT4AB/E2MID[3] Tile_X8Y1_LUT4AB/E2MID[4]
+ Tile_X8Y1_LUT4AB/E2MID[5] Tile_X8Y1_LUT4AB/E2MID[6] Tile_X8Y1_LUT4AB/E2MID[7] Tile_X9Y1_LUT4AB/E6END[0]
+ Tile_X9Y1_LUT4AB/E6END[10] Tile_X9Y1_LUT4AB/E6END[11] Tile_X9Y1_LUT4AB/E6END[1]
+ Tile_X9Y1_LUT4AB/E6END[2] Tile_X9Y1_LUT4AB/E6END[3] Tile_X9Y1_LUT4AB/E6END[4] Tile_X9Y1_LUT4AB/E6END[5]
+ Tile_X9Y1_LUT4AB/E6END[6] Tile_X9Y1_LUT4AB/E6END[7] Tile_X9Y1_LUT4AB/E6END[8] Tile_X9Y1_LUT4AB/E6END[9]
+ Tile_X8Y1_LUT4AB/E6END[0] Tile_X8Y1_LUT4AB/E6END[10] Tile_X8Y1_LUT4AB/E6END[11]
+ Tile_X8Y1_LUT4AB/E6END[1] Tile_X8Y1_LUT4AB/E6END[2] Tile_X8Y1_LUT4AB/E6END[3] Tile_X8Y1_LUT4AB/E6END[4]
+ Tile_X8Y1_LUT4AB/E6END[5] Tile_X8Y1_LUT4AB/E6END[6] Tile_X8Y1_LUT4AB/E6END[7] Tile_X8Y1_LUT4AB/E6END[8]
+ Tile_X8Y1_LUT4AB/E6END[9] Tile_X9Y1_LUT4AB/EE4END[0] Tile_X9Y1_LUT4AB/EE4END[10]
+ Tile_X9Y1_LUT4AB/EE4END[11] Tile_X9Y1_LUT4AB/EE4END[12] Tile_X9Y1_LUT4AB/EE4END[13]
+ Tile_X9Y1_LUT4AB/EE4END[14] Tile_X9Y1_LUT4AB/EE4END[15] Tile_X9Y1_LUT4AB/EE4END[1]
+ Tile_X9Y1_LUT4AB/EE4END[2] Tile_X9Y1_LUT4AB/EE4END[3] Tile_X9Y1_LUT4AB/EE4END[4]
+ Tile_X9Y1_LUT4AB/EE4END[5] Tile_X9Y1_LUT4AB/EE4END[6] Tile_X9Y1_LUT4AB/EE4END[7]
+ Tile_X9Y1_LUT4AB/EE4END[8] Tile_X9Y1_LUT4AB/EE4END[9] Tile_X8Y1_LUT4AB/EE4END[0]
+ Tile_X8Y1_LUT4AB/EE4END[10] Tile_X8Y1_LUT4AB/EE4END[11] Tile_X8Y1_LUT4AB/EE4END[12]
+ Tile_X8Y1_LUT4AB/EE4END[13] Tile_X8Y1_LUT4AB/EE4END[14] Tile_X8Y1_LUT4AB/EE4END[15]
+ Tile_X8Y1_LUT4AB/EE4END[1] Tile_X8Y1_LUT4AB/EE4END[2] Tile_X8Y1_LUT4AB/EE4END[3]
+ Tile_X8Y1_LUT4AB/EE4END[4] Tile_X8Y1_LUT4AB/EE4END[5] Tile_X8Y1_LUT4AB/EE4END[6]
+ Tile_X8Y1_LUT4AB/EE4END[7] Tile_X8Y1_LUT4AB/EE4END[8] Tile_X8Y1_LUT4AB/EE4END[9]
+ Tile_X8Y1_LUT4AB/FrameData[0] Tile_X8Y1_LUT4AB/FrameData[10] Tile_X8Y1_LUT4AB/FrameData[11]
+ Tile_X8Y1_LUT4AB/FrameData[12] Tile_X8Y1_LUT4AB/FrameData[13] Tile_X8Y1_LUT4AB/FrameData[14]
+ Tile_X8Y1_LUT4AB/FrameData[15] Tile_X8Y1_LUT4AB/FrameData[16] Tile_X8Y1_LUT4AB/FrameData[17]
+ Tile_X8Y1_LUT4AB/FrameData[18] Tile_X8Y1_LUT4AB/FrameData[19] Tile_X8Y1_LUT4AB/FrameData[1]
+ Tile_X8Y1_LUT4AB/FrameData[20] Tile_X8Y1_LUT4AB/FrameData[21] Tile_X8Y1_LUT4AB/FrameData[22]
+ Tile_X8Y1_LUT4AB/FrameData[23] Tile_X8Y1_LUT4AB/FrameData[24] Tile_X8Y1_LUT4AB/FrameData[25]
+ Tile_X8Y1_LUT4AB/FrameData[26] Tile_X8Y1_LUT4AB/FrameData[27] Tile_X8Y1_LUT4AB/FrameData[28]
+ Tile_X8Y1_LUT4AB/FrameData[29] Tile_X8Y1_LUT4AB/FrameData[2] Tile_X8Y1_LUT4AB/FrameData[30]
+ Tile_X8Y1_LUT4AB/FrameData[31] Tile_X8Y1_LUT4AB/FrameData[3] Tile_X8Y1_LUT4AB/FrameData[4]
+ Tile_X8Y1_LUT4AB/FrameData[5] Tile_X8Y1_LUT4AB/FrameData[6] Tile_X8Y1_LUT4AB/FrameData[7]
+ Tile_X8Y1_LUT4AB/FrameData[8] Tile_X8Y1_LUT4AB/FrameData[9] Tile_X9Y1_LUT4AB/FrameData[0]
+ Tile_X9Y1_LUT4AB/FrameData[10] Tile_X9Y1_LUT4AB/FrameData[11] Tile_X9Y1_LUT4AB/FrameData[12]
+ Tile_X9Y1_LUT4AB/FrameData[13] Tile_X9Y1_LUT4AB/FrameData[14] Tile_X9Y1_LUT4AB/FrameData[15]
+ Tile_X9Y1_LUT4AB/FrameData[16] Tile_X9Y1_LUT4AB/FrameData[17] Tile_X9Y1_LUT4AB/FrameData[18]
+ Tile_X9Y1_LUT4AB/FrameData[19] Tile_X9Y1_LUT4AB/FrameData[1] Tile_X9Y1_LUT4AB/FrameData[20]
+ Tile_X9Y1_LUT4AB/FrameData[21] Tile_X9Y1_LUT4AB/FrameData[22] Tile_X9Y1_LUT4AB/FrameData[23]
+ Tile_X9Y1_LUT4AB/FrameData[24] Tile_X9Y1_LUT4AB/FrameData[25] Tile_X9Y1_LUT4AB/FrameData[26]
+ Tile_X9Y1_LUT4AB/FrameData[27] Tile_X9Y1_LUT4AB/FrameData[28] Tile_X9Y1_LUT4AB/FrameData[29]
+ Tile_X9Y1_LUT4AB/FrameData[2] Tile_X9Y1_LUT4AB/FrameData[30] Tile_X9Y1_LUT4AB/FrameData[31]
+ Tile_X9Y1_LUT4AB/FrameData[3] Tile_X9Y1_LUT4AB/FrameData[4] Tile_X9Y1_LUT4AB/FrameData[5]
+ Tile_X9Y1_LUT4AB/FrameData[6] Tile_X9Y1_LUT4AB/FrameData[7] Tile_X9Y1_LUT4AB/FrameData[8]
+ Tile_X9Y1_LUT4AB/FrameData[9] Tile_X8Y1_LUT4AB/FrameStrobe[0] Tile_X8Y1_LUT4AB/FrameStrobe[10]
+ Tile_X8Y1_LUT4AB/FrameStrobe[11] Tile_X8Y1_LUT4AB/FrameStrobe[12] Tile_X8Y1_LUT4AB/FrameStrobe[13]
+ Tile_X8Y1_LUT4AB/FrameStrobe[14] Tile_X8Y1_LUT4AB/FrameStrobe[15] Tile_X8Y1_LUT4AB/FrameStrobe[16]
+ Tile_X8Y1_LUT4AB/FrameStrobe[17] Tile_X8Y1_LUT4AB/FrameStrobe[18] Tile_X8Y1_LUT4AB/FrameStrobe[19]
+ Tile_X8Y1_LUT4AB/FrameStrobe[1] Tile_X8Y1_LUT4AB/FrameStrobe[2] Tile_X8Y1_LUT4AB/FrameStrobe[3]
+ Tile_X8Y1_LUT4AB/FrameStrobe[4] Tile_X8Y1_LUT4AB/FrameStrobe[5] Tile_X8Y1_LUT4AB/FrameStrobe[6]
+ Tile_X8Y1_LUT4AB/FrameStrobe[7] Tile_X8Y1_LUT4AB/FrameStrobe[8] Tile_X8Y1_LUT4AB/FrameStrobe[9]
+ Tile_X8Y1_LUT4AB/FrameStrobe_O[0] Tile_X8Y1_LUT4AB/FrameStrobe_O[10] Tile_X8Y1_LUT4AB/FrameStrobe_O[11]
+ Tile_X8Y1_LUT4AB/FrameStrobe_O[12] Tile_X8Y1_LUT4AB/FrameStrobe_O[13] Tile_X8Y1_LUT4AB/FrameStrobe_O[14]
+ Tile_X8Y1_LUT4AB/FrameStrobe_O[15] Tile_X8Y1_LUT4AB/FrameStrobe_O[16] Tile_X8Y1_LUT4AB/FrameStrobe_O[17]
+ Tile_X8Y1_LUT4AB/FrameStrobe_O[18] Tile_X8Y1_LUT4AB/FrameStrobe_O[19] Tile_X8Y1_LUT4AB/FrameStrobe_O[1]
+ Tile_X8Y1_LUT4AB/FrameStrobe_O[2] Tile_X8Y1_LUT4AB/FrameStrobe_O[3] Tile_X8Y1_LUT4AB/FrameStrobe_O[4]
+ Tile_X8Y1_LUT4AB/FrameStrobe_O[5] Tile_X8Y1_LUT4AB/FrameStrobe_O[6] Tile_X8Y1_LUT4AB/FrameStrobe_O[7]
+ Tile_X8Y1_LUT4AB/FrameStrobe_O[8] Tile_X8Y1_LUT4AB/FrameStrobe_O[9] Tile_X8Y1_LUT4AB/N1BEG[0]
+ Tile_X8Y1_LUT4AB/N1BEG[1] Tile_X8Y1_LUT4AB/N1BEG[2] Tile_X8Y1_LUT4AB/N1BEG[3] Tile_X8Y2_LUT4AB/N1BEG[0]
+ Tile_X8Y2_LUT4AB/N1BEG[1] Tile_X8Y2_LUT4AB/N1BEG[2] Tile_X8Y2_LUT4AB/N1BEG[3] Tile_X8Y1_LUT4AB/N2BEG[0]
+ Tile_X8Y1_LUT4AB/N2BEG[1] Tile_X8Y1_LUT4AB/N2BEG[2] Tile_X8Y1_LUT4AB/N2BEG[3] Tile_X8Y1_LUT4AB/N2BEG[4]
+ Tile_X8Y1_LUT4AB/N2BEG[5] Tile_X8Y1_LUT4AB/N2BEG[6] Tile_X8Y1_LUT4AB/N2BEG[7] Tile_X8Y1_LUT4AB/N2BEGb[0]
+ Tile_X8Y1_LUT4AB/N2BEGb[1] Tile_X8Y1_LUT4AB/N2BEGb[2] Tile_X8Y1_LUT4AB/N2BEGb[3]
+ Tile_X8Y1_LUT4AB/N2BEGb[4] Tile_X8Y1_LUT4AB/N2BEGb[5] Tile_X8Y1_LUT4AB/N2BEGb[6]
+ Tile_X8Y1_LUT4AB/N2BEGb[7] Tile_X8Y1_LUT4AB/N2END[0] Tile_X8Y1_LUT4AB/N2END[1] Tile_X8Y1_LUT4AB/N2END[2]
+ Tile_X8Y1_LUT4AB/N2END[3] Tile_X8Y1_LUT4AB/N2END[4] Tile_X8Y1_LUT4AB/N2END[5] Tile_X8Y1_LUT4AB/N2END[6]
+ Tile_X8Y1_LUT4AB/N2END[7] Tile_X8Y2_LUT4AB/N2BEG[0] Tile_X8Y2_LUT4AB/N2BEG[1] Tile_X8Y2_LUT4AB/N2BEG[2]
+ Tile_X8Y2_LUT4AB/N2BEG[3] Tile_X8Y2_LUT4AB/N2BEG[4] Tile_X8Y2_LUT4AB/N2BEG[5] Tile_X8Y2_LUT4AB/N2BEG[6]
+ Tile_X8Y2_LUT4AB/N2BEG[7] Tile_X8Y1_LUT4AB/N4BEG[0] Tile_X8Y1_LUT4AB/N4BEG[10] Tile_X8Y1_LUT4AB/N4BEG[11]
+ Tile_X8Y1_LUT4AB/N4BEG[12] Tile_X8Y1_LUT4AB/N4BEG[13] Tile_X8Y1_LUT4AB/N4BEG[14]
+ Tile_X8Y1_LUT4AB/N4BEG[15] Tile_X8Y1_LUT4AB/N4BEG[1] Tile_X8Y1_LUT4AB/N4BEG[2] Tile_X8Y1_LUT4AB/N4BEG[3]
+ Tile_X8Y1_LUT4AB/N4BEG[4] Tile_X8Y1_LUT4AB/N4BEG[5] Tile_X8Y1_LUT4AB/N4BEG[6] Tile_X8Y1_LUT4AB/N4BEG[7]
+ Tile_X8Y1_LUT4AB/N4BEG[8] Tile_X8Y1_LUT4AB/N4BEG[9] Tile_X8Y2_LUT4AB/N4BEG[0] Tile_X8Y2_LUT4AB/N4BEG[10]
+ Tile_X8Y2_LUT4AB/N4BEG[11] Tile_X8Y2_LUT4AB/N4BEG[12] Tile_X8Y2_LUT4AB/N4BEG[13]
+ Tile_X8Y2_LUT4AB/N4BEG[14] Tile_X8Y2_LUT4AB/N4BEG[15] Tile_X8Y2_LUT4AB/N4BEG[1]
+ Tile_X8Y2_LUT4AB/N4BEG[2] Tile_X8Y2_LUT4AB/N4BEG[3] Tile_X8Y2_LUT4AB/N4BEG[4] Tile_X8Y2_LUT4AB/N4BEG[5]
+ Tile_X8Y2_LUT4AB/N4BEG[6] Tile_X8Y2_LUT4AB/N4BEG[7] Tile_X8Y2_LUT4AB/N4BEG[8] Tile_X8Y2_LUT4AB/N4BEG[9]
+ Tile_X8Y1_LUT4AB/NN4BEG[0] Tile_X8Y1_LUT4AB/NN4BEG[10] Tile_X8Y1_LUT4AB/NN4BEG[11]
+ Tile_X8Y1_LUT4AB/NN4BEG[12] Tile_X8Y1_LUT4AB/NN4BEG[13] Tile_X8Y1_LUT4AB/NN4BEG[14]
+ Tile_X8Y1_LUT4AB/NN4BEG[15] Tile_X8Y1_LUT4AB/NN4BEG[1] Tile_X8Y1_LUT4AB/NN4BEG[2]
+ Tile_X8Y1_LUT4AB/NN4BEG[3] Tile_X8Y1_LUT4AB/NN4BEG[4] Tile_X8Y1_LUT4AB/NN4BEG[5]
+ Tile_X8Y1_LUT4AB/NN4BEG[6] Tile_X8Y1_LUT4AB/NN4BEG[7] Tile_X8Y1_LUT4AB/NN4BEG[8]
+ Tile_X8Y1_LUT4AB/NN4BEG[9] Tile_X8Y2_LUT4AB/NN4BEG[0] Tile_X8Y2_LUT4AB/NN4BEG[10]
+ Tile_X8Y2_LUT4AB/NN4BEG[11] Tile_X8Y2_LUT4AB/NN4BEG[12] Tile_X8Y2_LUT4AB/NN4BEG[13]
+ Tile_X8Y2_LUT4AB/NN4BEG[14] Tile_X8Y2_LUT4AB/NN4BEG[15] Tile_X8Y2_LUT4AB/NN4BEG[1]
+ Tile_X8Y2_LUT4AB/NN4BEG[2] Tile_X8Y2_LUT4AB/NN4BEG[3] Tile_X8Y2_LUT4AB/NN4BEG[4]
+ Tile_X8Y2_LUT4AB/NN4BEG[5] Tile_X8Y2_LUT4AB/NN4BEG[6] Tile_X8Y2_LUT4AB/NN4BEG[7]
+ Tile_X8Y2_LUT4AB/NN4BEG[8] Tile_X8Y2_LUT4AB/NN4BEG[9] Tile_X8Y2_LUT4AB/S1END[0]
+ Tile_X8Y2_LUT4AB/S1END[1] Tile_X8Y2_LUT4AB/S1END[2] Tile_X8Y2_LUT4AB/S1END[3] Tile_X8Y1_LUT4AB/S1END[0]
+ Tile_X8Y1_LUT4AB/S1END[1] Tile_X8Y1_LUT4AB/S1END[2] Tile_X8Y1_LUT4AB/S1END[3] Tile_X8Y2_LUT4AB/S2MID[0]
+ Tile_X8Y2_LUT4AB/S2MID[1] Tile_X8Y2_LUT4AB/S2MID[2] Tile_X8Y2_LUT4AB/S2MID[3] Tile_X8Y2_LUT4AB/S2MID[4]
+ Tile_X8Y2_LUT4AB/S2MID[5] Tile_X8Y2_LUT4AB/S2MID[6] Tile_X8Y2_LUT4AB/S2MID[7] Tile_X8Y2_LUT4AB/S2END[0]
+ Tile_X8Y2_LUT4AB/S2END[1] Tile_X8Y2_LUT4AB/S2END[2] Tile_X8Y2_LUT4AB/S2END[3] Tile_X8Y2_LUT4AB/S2END[4]
+ Tile_X8Y2_LUT4AB/S2END[5] Tile_X8Y2_LUT4AB/S2END[6] Tile_X8Y2_LUT4AB/S2END[7] Tile_X8Y1_LUT4AB/S2END[0]
+ Tile_X8Y1_LUT4AB/S2END[1] Tile_X8Y1_LUT4AB/S2END[2] Tile_X8Y1_LUT4AB/S2END[3] Tile_X8Y1_LUT4AB/S2END[4]
+ Tile_X8Y1_LUT4AB/S2END[5] Tile_X8Y1_LUT4AB/S2END[6] Tile_X8Y1_LUT4AB/S2END[7] Tile_X8Y1_LUT4AB/S2MID[0]
+ Tile_X8Y1_LUT4AB/S2MID[1] Tile_X8Y1_LUT4AB/S2MID[2] Tile_X8Y1_LUT4AB/S2MID[3] Tile_X8Y1_LUT4AB/S2MID[4]
+ Tile_X8Y1_LUT4AB/S2MID[5] Tile_X8Y1_LUT4AB/S2MID[6] Tile_X8Y1_LUT4AB/S2MID[7] Tile_X8Y2_LUT4AB/S4END[0]
+ Tile_X8Y2_LUT4AB/S4END[10] Tile_X8Y2_LUT4AB/S4END[11] Tile_X8Y2_LUT4AB/S4END[12]
+ Tile_X8Y2_LUT4AB/S4END[13] Tile_X8Y2_LUT4AB/S4END[14] Tile_X8Y2_LUT4AB/S4END[15]
+ Tile_X8Y2_LUT4AB/S4END[1] Tile_X8Y2_LUT4AB/S4END[2] Tile_X8Y2_LUT4AB/S4END[3] Tile_X8Y2_LUT4AB/S4END[4]
+ Tile_X8Y2_LUT4AB/S4END[5] Tile_X8Y2_LUT4AB/S4END[6] Tile_X8Y2_LUT4AB/S4END[7] Tile_X8Y2_LUT4AB/S4END[8]
+ Tile_X8Y2_LUT4AB/S4END[9] Tile_X8Y1_LUT4AB/S4END[0] Tile_X8Y1_LUT4AB/S4END[10] Tile_X8Y1_LUT4AB/S4END[11]
+ Tile_X8Y1_LUT4AB/S4END[12] Tile_X8Y1_LUT4AB/S4END[13] Tile_X8Y1_LUT4AB/S4END[14]
+ Tile_X8Y1_LUT4AB/S4END[15] Tile_X8Y1_LUT4AB/S4END[1] Tile_X8Y1_LUT4AB/S4END[2] Tile_X8Y1_LUT4AB/S4END[3]
+ Tile_X8Y1_LUT4AB/S4END[4] Tile_X8Y1_LUT4AB/S4END[5] Tile_X8Y1_LUT4AB/S4END[6] Tile_X8Y1_LUT4AB/S4END[7]
+ Tile_X8Y1_LUT4AB/S4END[8] Tile_X8Y1_LUT4AB/S4END[9] Tile_X8Y2_LUT4AB/SS4END[0] Tile_X8Y2_LUT4AB/SS4END[10]
+ Tile_X8Y2_LUT4AB/SS4END[11] Tile_X8Y2_LUT4AB/SS4END[12] Tile_X8Y2_LUT4AB/SS4END[13]
+ Tile_X8Y2_LUT4AB/SS4END[14] Tile_X8Y2_LUT4AB/SS4END[15] Tile_X8Y2_LUT4AB/SS4END[1]
+ Tile_X8Y2_LUT4AB/SS4END[2] Tile_X8Y2_LUT4AB/SS4END[3] Tile_X8Y2_LUT4AB/SS4END[4]
+ Tile_X8Y2_LUT4AB/SS4END[5] Tile_X8Y2_LUT4AB/SS4END[6] Tile_X8Y2_LUT4AB/SS4END[7]
+ Tile_X8Y2_LUT4AB/SS4END[8] Tile_X8Y2_LUT4AB/SS4END[9] Tile_X8Y1_LUT4AB/SS4END[0]
+ Tile_X8Y1_LUT4AB/SS4END[10] Tile_X8Y1_LUT4AB/SS4END[11] Tile_X8Y1_LUT4AB/SS4END[12]
+ Tile_X8Y1_LUT4AB/SS4END[13] Tile_X8Y1_LUT4AB/SS4END[14] Tile_X8Y1_LUT4AB/SS4END[15]
+ Tile_X8Y1_LUT4AB/SS4END[1] Tile_X8Y1_LUT4AB/SS4END[2] Tile_X8Y1_LUT4AB/SS4END[3]
+ Tile_X8Y1_LUT4AB/SS4END[4] Tile_X8Y1_LUT4AB/SS4END[5] Tile_X8Y1_LUT4AB/SS4END[6]
+ Tile_X8Y1_LUT4AB/SS4END[7] Tile_X8Y1_LUT4AB/SS4END[8] Tile_X8Y1_LUT4AB/SS4END[9]
+ Tile_X8Y1_LUT4AB/UserCLK Tile_X8Y1_LUT4AB/UserCLKo VGND VPWR Tile_X8Y1_LUT4AB/W1BEG[0]
+ Tile_X8Y1_LUT4AB/W1BEG[1] Tile_X8Y1_LUT4AB/W1BEG[2] Tile_X8Y1_LUT4AB/W1BEG[3] Tile_X9Y1_LUT4AB/W1BEG[0]
+ Tile_X9Y1_LUT4AB/W1BEG[1] Tile_X9Y1_LUT4AB/W1BEG[2] Tile_X9Y1_LUT4AB/W1BEG[3] Tile_X8Y1_LUT4AB/W2BEG[0]
+ Tile_X8Y1_LUT4AB/W2BEG[1] Tile_X8Y1_LUT4AB/W2BEG[2] Tile_X8Y1_LUT4AB/W2BEG[3] Tile_X8Y1_LUT4AB/W2BEG[4]
+ Tile_X8Y1_LUT4AB/W2BEG[5] Tile_X8Y1_LUT4AB/W2BEG[6] Tile_X8Y1_LUT4AB/W2BEG[7] Tile_X8Y1_LUT4AB/W2BEGb[0]
+ Tile_X8Y1_LUT4AB/W2BEGb[1] Tile_X8Y1_LUT4AB/W2BEGb[2] Tile_X8Y1_LUT4AB/W2BEGb[3]
+ Tile_X8Y1_LUT4AB/W2BEGb[4] Tile_X8Y1_LUT4AB/W2BEGb[5] Tile_X8Y1_LUT4AB/W2BEGb[6]
+ Tile_X8Y1_LUT4AB/W2BEGb[7] Tile_X8Y1_LUT4AB/W2END[0] Tile_X8Y1_LUT4AB/W2END[1] Tile_X8Y1_LUT4AB/W2END[2]
+ Tile_X8Y1_LUT4AB/W2END[3] Tile_X8Y1_LUT4AB/W2END[4] Tile_X8Y1_LUT4AB/W2END[5] Tile_X8Y1_LUT4AB/W2END[6]
+ Tile_X8Y1_LUT4AB/W2END[7] Tile_X9Y1_LUT4AB/W2BEG[0] Tile_X9Y1_LUT4AB/W2BEG[1] Tile_X9Y1_LUT4AB/W2BEG[2]
+ Tile_X9Y1_LUT4AB/W2BEG[3] Tile_X9Y1_LUT4AB/W2BEG[4] Tile_X9Y1_LUT4AB/W2BEG[5] Tile_X9Y1_LUT4AB/W2BEG[6]
+ Tile_X9Y1_LUT4AB/W2BEG[7] Tile_X8Y1_LUT4AB/W6BEG[0] Tile_X8Y1_LUT4AB/W6BEG[10] Tile_X8Y1_LUT4AB/W6BEG[11]
+ Tile_X8Y1_LUT4AB/W6BEG[1] Tile_X8Y1_LUT4AB/W6BEG[2] Tile_X8Y1_LUT4AB/W6BEG[3] Tile_X8Y1_LUT4AB/W6BEG[4]
+ Tile_X8Y1_LUT4AB/W6BEG[5] Tile_X8Y1_LUT4AB/W6BEG[6] Tile_X8Y1_LUT4AB/W6BEG[7] Tile_X8Y1_LUT4AB/W6BEG[8]
+ Tile_X8Y1_LUT4AB/W6BEG[9] Tile_X9Y1_LUT4AB/W6BEG[0] Tile_X9Y1_LUT4AB/W6BEG[10] Tile_X9Y1_LUT4AB/W6BEG[11]
+ Tile_X9Y1_LUT4AB/W6BEG[1] Tile_X9Y1_LUT4AB/W6BEG[2] Tile_X9Y1_LUT4AB/W6BEG[3] Tile_X9Y1_LUT4AB/W6BEG[4]
+ Tile_X9Y1_LUT4AB/W6BEG[5] Tile_X9Y1_LUT4AB/W6BEG[6] Tile_X9Y1_LUT4AB/W6BEG[7] Tile_X9Y1_LUT4AB/W6BEG[8]
+ Tile_X9Y1_LUT4AB/W6BEG[9] Tile_X8Y1_LUT4AB/WW4BEG[0] Tile_X8Y1_LUT4AB/WW4BEG[10]
+ Tile_X8Y1_LUT4AB/WW4BEG[11] Tile_X8Y1_LUT4AB/WW4BEG[12] Tile_X8Y1_LUT4AB/WW4BEG[13]
+ Tile_X8Y1_LUT4AB/WW4BEG[14] Tile_X8Y1_LUT4AB/WW4BEG[15] Tile_X8Y1_LUT4AB/WW4BEG[1]
+ Tile_X8Y1_LUT4AB/WW4BEG[2] Tile_X8Y1_LUT4AB/WW4BEG[3] Tile_X8Y1_LUT4AB/WW4BEG[4]
+ Tile_X8Y1_LUT4AB/WW4BEG[5] Tile_X8Y1_LUT4AB/WW4BEG[6] Tile_X8Y1_LUT4AB/WW4BEG[7]
+ Tile_X8Y1_LUT4AB/WW4BEG[8] Tile_X8Y1_LUT4AB/WW4BEG[9] Tile_X9Y1_LUT4AB/WW4BEG[0]
+ Tile_X9Y1_LUT4AB/WW4BEG[10] Tile_X9Y1_LUT4AB/WW4BEG[11] Tile_X9Y1_LUT4AB/WW4BEG[12]
+ Tile_X9Y1_LUT4AB/WW4BEG[13] Tile_X9Y1_LUT4AB/WW4BEG[14] Tile_X9Y1_LUT4AB/WW4BEG[15]
+ Tile_X9Y1_LUT4AB/WW4BEG[1] Tile_X9Y1_LUT4AB/WW4BEG[2] Tile_X9Y1_LUT4AB/WW4BEG[3]
+ Tile_X9Y1_LUT4AB/WW4BEG[4] Tile_X9Y1_LUT4AB/WW4BEG[5] Tile_X9Y1_LUT4AB/WW4BEG[6]
+ Tile_X9Y1_LUT4AB/WW4BEG[7] Tile_X9Y1_LUT4AB/WW4BEG[8] Tile_X9Y1_LUT4AB/WW4BEG[9]
+ LUT4AB
XTile_X3Y11_LUT4AB Tile_X3Y12_LUT4AB/Co Tile_X3Y11_LUT4AB/Co Tile_X3Y11_LUT4AB/E1BEG[0]
+ Tile_X3Y11_LUT4AB/E1BEG[1] Tile_X3Y11_LUT4AB/E1BEG[2] Tile_X3Y11_LUT4AB/E1BEG[3]
+ Tile_X3Y11_LUT4AB/E1END[0] Tile_X3Y11_LUT4AB/E1END[1] Tile_X3Y11_LUT4AB/E1END[2]
+ Tile_X3Y11_LUT4AB/E1END[3] Tile_X3Y11_LUT4AB/E2BEG[0] Tile_X3Y11_LUT4AB/E2BEG[1]
+ Tile_X3Y11_LUT4AB/E2BEG[2] Tile_X3Y11_LUT4AB/E2BEG[3] Tile_X3Y11_LUT4AB/E2BEG[4]
+ Tile_X3Y11_LUT4AB/E2BEG[5] Tile_X3Y11_LUT4AB/E2BEG[6] Tile_X3Y11_LUT4AB/E2BEG[7]
+ Tile_X4Y11_RegFile/E2END[0] Tile_X4Y11_RegFile/E2END[1] Tile_X4Y11_RegFile/E2END[2]
+ Tile_X4Y11_RegFile/E2END[3] Tile_X4Y11_RegFile/E2END[4] Tile_X4Y11_RegFile/E2END[5]
+ Tile_X4Y11_RegFile/E2END[6] Tile_X4Y11_RegFile/E2END[7] Tile_X3Y11_LUT4AB/E2END[0]
+ Tile_X3Y11_LUT4AB/E2END[1] Tile_X3Y11_LUT4AB/E2END[2] Tile_X3Y11_LUT4AB/E2END[3]
+ Tile_X3Y11_LUT4AB/E2END[4] Tile_X3Y11_LUT4AB/E2END[5] Tile_X3Y11_LUT4AB/E2END[6]
+ Tile_X3Y11_LUT4AB/E2END[7] Tile_X3Y11_LUT4AB/E2MID[0] Tile_X3Y11_LUT4AB/E2MID[1]
+ Tile_X3Y11_LUT4AB/E2MID[2] Tile_X3Y11_LUT4AB/E2MID[3] Tile_X3Y11_LUT4AB/E2MID[4]
+ Tile_X3Y11_LUT4AB/E2MID[5] Tile_X3Y11_LUT4AB/E2MID[6] Tile_X3Y11_LUT4AB/E2MID[7]
+ Tile_X3Y11_LUT4AB/E6BEG[0] Tile_X3Y11_LUT4AB/E6BEG[10] Tile_X3Y11_LUT4AB/E6BEG[11]
+ Tile_X3Y11_LUT4AB/E6BEG[1] Tile_X3Y11_LUT4AB/E6BEG[2] Tile_X3Y11_LUT4AB/E6BEG[3]
+ Tile_X3Y11_LUT4AB/E6BEG[4] Tile_X3Y11_LUT4AB/E6BEG[5] Tile_X3Y11_LUT4AB/E6BEG[6]
+ Tile_X3Y11_LUT4AB/E6BEG[7] Tile_X3Y11_LUT4AB/E6BEG[8] Tile_X3Y11_LUT4AB/E6BEG[9]
+ Tile_X3Y11_LUT4AB/E6END[0] Tile_X3Y11_LUT4AB/E6END[10] Tile_X3Y11_LUT4AB/E6END[11]
+ Tile_X3Y11_LUT4AB/E6END[1] Tile_X3Y11_LUT4AB/E6END[2] Tile_X3Y11_LUT4AB/E6END[3]
+ Tile_X3Y11_LUT4AB/E6END[4] Tile_X3Y11_LUT4AB/E6END[5] Tile_X3Y11_LUT4AB/E6END[6]
+ Tile_X3Y11_LUT4AB/E6END[7] Tile_X3Y11_LUT4AB/E6END[8] Tile_X3Y11_LUT4AB/E6END[9]
+ Tile_X3Y11_LUT4AB/EE4BEG[0] Tile_X3Y11_LUT4AB/EE4BEG[10] Tile_X3Y11_LUT4AB/EE4BEG[11]
+ Tile_X3Y11_LUT4AB/EE4BEG[12] Tile_X3Y11_LUT4AB/EE4BEG[13] Tile_X3Y11_LUT4AB/EE4BEG[14]
+ Tile_X3Y11_LUT4AB/EE4BEG[15] Tile_X3Y11_LUT4AB/EE4BEG[1] Tile_X3Y11_LUT4AB/EE4BEG[2]
+ Tile_X3Y11_LUT4AB/EE4BEG[3] Tile_X3Y11_LUT4AB/EE4BEG[4] Tile_X3Y11_LUT4AB/EE4BEG[5]
+ Tile_X3Y11_LUT4AB/EE4BEG[6] Tile_X3Y11_LUT4AB/EE4BEG[7] Tile_X3Y11_LUT4AB/EE4BEG[8]
+ Tile_X3Y11_LUT4AB/EE4BEG[9] Tile_X3Y11_LUT4AB/EE4END[0] Tile_X3Y11_LUT4AB/EE4END[10]
+ Tile_X3Y11_LUT4AB/EE4END[11] Tile_X3Y11_LUT4AB/EE4END[12] Tile_X3Y11_LUT4AB/EE4END[13]
+ Tile_X3Y11_LUT4AB/EE4END[14] Tile_X3Y11_LUT4AB/EE4END[15] Tile_X3Y11_LUT4AB/EE4END[1]
+ Tile_X3Y11_LUT4AB/EE4END[2] Tile_X3Y11_LUT4AB/EE4END[3] Tile_X3Y11_LUT4AB/EE4END[4]
+ Tile_X3Y11_LUT4AB/EE4END[5] Tile_X3Y11_LUT4AB/EE4END[6] Tile_X3Y11_LUT4AB/EE4END[7]
+ Tile_X3Y11_LUT4AB/EE4END[8] Tile_X3Y11_LUT4AB/EE4END[9] Tile_X3Y11_LUT4AB/FrameData[0]
+ Tile_X3Y11_LUT4AB/FrameData[10] Tile_X3Y11_LUT4AB/FrameData[11] Tile_X3Y11_LUT4AB/FrameData[12]
+ Tile_X3Y11_LUT4AB/FrameData[13] Tile_X3Y11_LUT4AB/FrameData[14] Tile_X3Y11_LUT4AB/FrameData[15]
+ Tile_X3Y11_LUT4AB/FrameData[16] Tile_X3Y11_LUT4AB/FrameData[17] Tile_X3Y11_LUT4AB/FrameData[18]
+ Tile_X3Y11_LUT4AB/FrameData[19] Tile_X3Y11_LUT4AB/FrameData[1] Tile_X3Y11_LUT4AB/FrameData[20]
+ Tile_X3Y11_LUT4AB/FrameData[21] Tile_X3Y11_LUT4AB/FrameData[22] Tile_X3Y11_LUT4AB/FrameData[23]
+ Tile_X3Y11_LUT4AB/FrameData[24] Tile_X3Y11_LUT4AB/FrameData[25] Tile_X3Y11_LUT4AB/FrameData[26]
+ Tile_X3Y11_LUT4AB/FrameData[27] Tile_X3Y11_LUT4AB/FrameData[28] Tile_X3Y11_LUT4AB/FrameData[29]
+ Tile_X3Y11_LUT4AB/FrameData[2] Tile_X3Y11_LUT4AB/FrameData[30] Tile_X3Y11_LUT4AB/FrameData[31]
+ Tile_X3Y11_LUT4AB/FrameData[3] Tile_X3Y11_LUT4AB/FrameData[4] Tile_X3Y11_LUT4AB/FrameData[5]
+ Tile_X3Y11_LUT4AB/FrameData[6] Tile_X3Y11_LUT4AB/FrameData[7] Tile_X3Y11_LUT4AB/FrameData[8]
+ Tile_X3Y11_LUT4AB/FrameData[9] Tile_X4Y11_RegFile/FrameData[0] Tile_X4Y11_RegFile/FrameData[10]
+ Tile_X4Y11_RegFile/FrameData[11] Tile_X4Y11_RegFile/FrameData[12] Tile_X4Y11_RegFile/FrameData[13]
+ Tile_X4Y11_RegFile/FrameData[14] Tile_X4Y11_RegFile/FrameData[15] Tile_X4Y11_RegFile/FrameData[16]
+ Tile_X4Y11_RegFile/FrameData[17] Tile_X4Y11_RegFile/FrameData[18] Tile_X4Y11_RegFile/FrameData[19]
+ Tile_X4Y11_RegFile/FrameData[1] Tile_X4Y11_RegFile/FrameData[20] Tile_X4Y11_RegFile/FrameData[21]
+ Tile_X4Y11_RegFile/FrameData[22] Tile_X4Y11_RegFile/FrameData[23] Tile_X4Y11_RegFile/FrameData[24]
+ Tile_X4Y11_RegFile/FrameData[25] Tile_X4Y11_RegFile/FrameData[26] Tile_X4Y11_RegFile/FrameData[27]
+ Tile_X4Y11_RegFile/FrameData[28] Tile_X4Y11_RegFile/FrameData[29] Tile_X4Y11_RegFile/FrameData[2]
+ Tile_X4Y11_RegFile/FrameData[30] Tile_X4Y11_RegFile/FrameData[31] Tile_X4Y11_RegFile/FrameData[3]
+ Tile_X4Y11_RegFile/FrameData[4] Tile_X4Y11_RegFile/FrameData[5] Tile_X4Y11_RegFile/FrameData[6]
+ Tile_X4Y11_RegFile/FrameData[7] Tile_X4Y11_RegFile/FrameData[8] Tile_X4Y11_RegFile/FrameData[9]
+ Tile_X3Y11_LUT4AB/FrameStrobe[0] Tile_X3Y11_LUT4AB/FrameStrobe[10] Tile_X3Y11_LUT4AB/FrameStrobe[11]
+ Tile_X3Y11_LUT4AB/FrameStrobe[12] Tile_X3Y11_LUT4AB/FrameStrobe[13] Tile_X3Y11_LUT4AB/FrameStrobe[14]
+ Tile_X3Y11_LUT4AB/FrameStrobe[15] Tile_X3Y11_LUT4AB/FrameStrobe[16] Tile_X3Y11_LUT4AB/FrameStrobe[17]
+ Tile_X3Y11_LUT4AB/FrameStrobe[18] Tile_X3Y11_LUT4AB/FrameStrobe[19] Tile_X3Y11_LUT4AB/FrameStrobe[1]
+ Tile_X3Y11_LUT4AB/FrameStrobe[2] Tile_X3Y11_LUT4AB/FrameStrobe[3] Tile_X3Y11_LUT4AB/FrameStrobe[4]
+ Tile_X3Y11_LUT4AB/FrameStrobe[5] Tile_X3Y11_LUT4AB/FrameStrobe[6] Tile_X3Y11_LUT4AB/FrameStrobe[7]
+ Tile_X3Y11_LUT4AB/FrameStrobe[8] Tile_X3Y11_LUT4AB/FrameStrobe[9] Tile_X3Y10_LUT4AB/FrameStrobe[0]
+ Tile_X3Y10_LUT4AB/FrameStrobe[10] Tile_X3Y10_LUT4AB/FrameStrobe[11] Tile_X3Y10_LUT4AB/FrameStrobe[12]
+ Tile_X3Y10_LUT4AB/FrameStrobe[13] Tile_X3Y10_LUT4AB/FrameStrobe[14] Tile_X3Y10_LUT4AB/FrameStrobe[15]
+ Tile_X3Y10_LUT4AB/FrameStrobe[16] Tile_X3Y10_LUT4AB/FrameStrobe[17] Tile_X3Y10_LUT4AB/FrameStrobe[18]
+ Tile_X3Y10_LUT4AB/FrameStrobe[19] Tile_X3Y10_LUT4AB/FrameStrobe[1] Tile_X3Y10_LUT4AB/FrameStrobe[2]
+ Tile_X3Y10_LUT4AB/FrameStrobe[3] Tile_X3Y10_LUT4AB/FrameStrobe[4] Tile_X3Y10_LUT4AB/FrameStrobe[5]
+ Tile_X3Y10_LUT4AB/FrameStrobe[6] Tile_X3Y10_LUT4AB/FrameStrobe[7] Tile_X3Y10_LUT4AB/FrameStrobe[8]
+ Tile_X3Y10_LUT4AB/FrameStrobe[9] Tile_X3Y11_LUT4AB/N1BEG[0] Tile_X3Y11_LUT4AB/N1BEG[1]
+ Tile_X3Y11_LUT4AB/N1BEG[2] Tile_X3Y11_LUT4AB/N1BEG[3] Tile_X3Y12_LUT4AB/N1BEG[0]
+ Tile_X3Y12_LUT4AB/N1BEG[1] Tile_X3Y12_LUT4AB/N1BEG[2] Tile_X3Y12_LUT4AB/N1BEG[3]
+ Tile_X3Y11_LUT4AB/N2BEG[0] Tile_X3Y11_LUT4AB/N2BEG[1] Tile_X3Y11_LUT4AB/N2BEG[2]
+ Tile_X3Y11_LUT4AB/N2BEG[3] Tile_X3Y11_LUT4AB/N2BEG[4] Tile_X3Y11_LUT4AB/N2BEG[5]
+ Tile_X3Y11_LUT4AB/N2BEG[6] Tile_X3Y11_LUT4AB/N2BEG[7] Tile_X3Y10_LUT4AB/N2END[0]
+ Tile_X3Y10_LUT4AB/N2END[1] Tile_X3Y10_LUT4AB/N2END[2] Tile_X3Y10_LUT4AB/N2END[3]
+ Tile_X3Y10_LUT4AB/N2END[4] Tile_X3Y10_LUT4AB/N2END[5] Tile_X3Y10_LUT4AB/N2END[6]
+ Tile_X3Y10_LUT4AB/N2END[7] Tile_X3Y11_LUT4AB/N2END[0] Tile_X3Y11_LUT4AB/N2END[1]
+ Tile_X3Y11_LUT4AB/N2END[2] Tile_X3Y11_LUT4AB/N2END[3] Tile_X3Y11_LUT4AB/N2END[4]
+ Tile_X3Y11_LUT4AB/N2END[5] Tile_X3Y11_LUT4AB/N2END[6] Tile_X3Y11_LUT4AB/N2END[7]
+ Tile_X3Y12_LUT4AB/N2BEG[0] Tile_X3Y12_LUT4AB/N2BEG[1] Tile_X3Y12_LUT4AB/N2BEG[2]
+ Tile_X3Y12_LUT4AB/N2BEG[3] Tile_X3Y12_LUT4AB/N2BEG[4] Tile_X3Y12_LUT4AB/N2BEG[5]
+ Tile_X3Y12_LUT4AB/N2BEG[6] Tile_X3Y12_LUT4AB/N2BEG[7] Tile_X3Y11_LUT4AB/N4BEG[0]
+ Tile_X3Y11_LUT4AB/N4BEG[10] Tile_X3Y11_LUT4AB/N4BEG[11] Tile_X3Y11_LUT4AB/N4BEG[12]
+ Tile_X3Y11_LUT4AB/N4BEG[13] Tile_X3Y11_LUT4AB/N4BEG[14] Tile_X3Y11_LUT4AB/N4BEG[15]
+ Tile_X3Y11_LUT4AB/N4BEG[1] Tile_X3Y11_LUT4AB/N4BEG[2] Tile_X3Y11_LUT4AB/N4BEG[3]
+ Tile_X3Y11_LUT4AB/N4BEG[4] Tile_X3Y11_LUT4AB/N4BEG[5] Tile_X3Y11_LUT4AB/N4BEG[6]
+ Tile_X3Y11_LUT4AB/N4BEG[7] Tile_X3Y11_LUT4AB/N4BEG[8] Tile_X3Y11_LUT4AB/N4BEG[9]
+ Tile_X3Y12_LUT4AB/N4BEG[0] Tile_X3Y12_LUT4AB/N4BEG[10] Tile_X3Y12_LUT4AB/N4BEG[11]
+ Tile_X3Y12_LUT4AB/N4BEG[12] Tile_X3Y12_LUT4AB/N4BEG[13] Tile_X3Y12_LUT4AB/N4BEG[14]
+ Tile_X3Y12_LUT4AB/N4BEG[15] Tile_X3Y12_LUT4AB/N4BEG[1] Tile_X3Y12_LUT4AB/N4BEG[2]
+ Tile_X3Y12_LUT4AB/N4BEG[3] Tile_X3Y12_LUT4AB/N4BEG[4] Tile_X3Y12_LUT4AB/N4BEG[5]
+ Tile_X3Y12_LUT4AB/N4BEG[6] Tile_X3Y12_LUT4AB/N4BEG[7] Tile_X3Y12_LUT4AB/N4BEG[8]
+ Tile_X3Y12_LUT4AB/N4BEG[9] Tile_X3Y11_LUT4AB/NN4BEG[0] Tile_X3Y11_LUT4AB/NN4BEG[10]
+ Tile_X3Y11_LUT4AB/NN4BEG[11] Tile_X3Y11_LUT4AB/NN4BEG[12] Tile_X3Y11_LUT4AB/NN4BEG[13]
+ Tile_X3Y11_LUT4AB/NN4BEG[14] Tile_X3Y11_LUT4AB/NN4BEG[15] Tile_X3Y11_LUT4AB/NN4BEG[1]
+ Tile_X3Y11_LUT4AB/NN4BEG[2] Tile_X3Y11_LUT4AB/NN4BEG[3] Tile_X3Y11_LUT4AB/NN4BEG[4]
+ Tile_X3Y11_LUT4AB/NN4BEG[5] Tile_X3Y11_LUT4AB/NN4BEG[6] Tile_X3Y11_LUT4AB/NN4BEG[7]
+ Tile_X3Y11_LUT4AB/NN4BEG[8] Tile_X3Y11_LUT4AB/NN4BEG[9] Tile_X3Y12_LUT4AB/NN4BEG[0]
+ Tile_X3Y12_LUT4AB/NN4BEG[10] Tile_X3Y12_LUT4AB/NN4BEG[11] Tile_X3Y12_LUT4AB/NN4BEG[12]
+ Tile_X3Y12_LUT4AB/NN4BEG[13] Tile_X3Y12_LUT4AB/NN4BEG[14] Tile_X3Y12_LUT4AB/NN4BEG[15]
+ Tile_X3Y12_LUT4AB/NN4BEG[1] Tile_X3Y12_LUT4AB/NN4BEG[2] Tile_X3Y12_LUT4AB/NN4BEG[3]
+ Tile_X3Y12_LUT4AB/NN4BEG[4] Tile_X3Y12_LUT4AB/NN4BEG[5] Tile_X3Y12_LUT4AB/NN4BEG[6]
+ Tile_X3Y12_LUT4AB/NN4BEG[7] Tile_X3Y12_LUT4AB/NN4BEG[8] Tile_X3Y12_LUT4AB/NN4BEG[9]
+ Tile_X3Y12_LUT4AB/S1END[0] Tile_X3Y12_LUT4AB/S1END[1] Tile_X3Y12_LUT4AB/S1END[2]
+ Tile_X3Y12_LUT4AB/S1END[3] Tile_X3Y11_LUT4AB/S1END[0] Tile_X3Y11_LUT4AB/S1END[1]
+ Tile_X3Y11_LUT4AB/S1END[2] Tile_X3Y11_LUT4AB/S1END[3] Tile_X3Y12_LUT4AB/S2MID[0]
+ Tile_X3Y12_LUT4AB/S2MID[1] Tile_X3Y12_LUT4AB/S2MID[2] Tile_X3Y12_LUT4AB/S2MID[3]
+ Tile_X3Y12_LUT4AB/S2MID[4] Tile_X3Y12_LUT4AB/S2MID[5] Tile_X3Y12_LUT4AB/S2MID[6]
+ Tile_X3Y12_LUT4AB/S2MID[7] Tile_X3Y12_LUT4AB/S2END[0] Tile_X3Y12_LUT4AB/S2END[1]
+ Tile_X3Y12_LUT4AB/S2END[2] Tile_X3Y12_LUT4AB/S2END[3] Tile_X3Y12_LUT4AB/S2END[4]
+ Tile_X3Y12_LUT4AB/S2END[5] Tile_X3Y12_LUT4AB/S2END[6] Tile_X3Y12_LUT4AB/S2END[7]
+ Tile_X3Y11_LUT4AB/S2END[0] Tile_X3Y11_LUT4AB/S2END[1] Tile_X3Y11_LUT4AB/S2END[2]
+ Tile_X3Y11_LUT4AB/S2END[3] Tile_X3Y11_LUT4AB/S2END[4] Tile_X3Y11_LUT4AB/S2END[5]
+ Tile_X3Y11_LUT4AB/S2END[6] Tile_X3Y11_LUT4AB/S2END[7] Tile_X3Y11_LUT4AB/S2MID[0]
+ Tile_X3Y11_LUT4AB/S2MID[1] Tile_X3Y11_LUT4AB/S2MID[2] Tile_X3Y11_LUT4AB/S2MID[3]
+ Tile_X3Y11_LUT4AB/S2MID[4] Tile_X3Y11_LUT4AB/S2MID[5] Tile_X3Y11_LUT4AB/S2MID[6]
+ Tile_X3Y11_LUT4AB/S2MID[7] Tile_X3Y12_LUT4AB/S4END[0] Tile_X3Y12_LUT4AB/S4END[10]
+ Tile_X3Y12_LUT4AB/S4END[11] Tile_X3Y12_LUT4AB/S4END[12] Tile_X3Y12_LUT4AB/S4END[13]
+ Tile_X3Y12_LUT4AB/S4END[14] Tile_X3Y12_LUT4AB/S4END[15] Tile_X3Y12_LUT4AB/S4END[1]
+ Tile_X3Y12_LUT4AB/S4END[2] Tile_X3Y12_LUT4AB/S4END[3] Tile_X3Y12_LUT4AB/S4END[4]
+ Tile_X3Y12_LUT4AB/S4END[5] Tile_X3Y12_LUT4AB/S4END[6] Tile_X3Y12_LUT4AB/S4END[7]
+ Tile_X3Y12_LUT4AB/S4END[8] Tile_X3Y12_LUT4AB/S4END[9] Tile_X3Y11_LUT4AB/S4END[0]
+ Tile_X3Y11_LUT4AB/S4END[10] Tile_X3Y11_LUT4AB/S4END[11] Tile_X3Y11_LUT4AB/S4END[12]
+ Tile_X3Y11_LUT4AB/S4END[13] Tile_X3Y11_LUT4AB/S4END[14] Tile_X3Y11_LUT4AB/S4END[15]
+ Tile_X3Y11_LUT4AB/S4END[1] Tile_X3Y11_LUT4AB/S4END[2] Tile_X3Y11_LUT4AB/S4END[3]
+ Tile_X3Y11_LUT4AB/S4END[4] Tile_X3Y11_LUT4AB/S4END[5] Tile_X3Y11_LUT4AB/S4END[6]
+ Tile_X3Y11_LUT4AB/S4END[7] Tile_X3Y11_LUT4AB/S4END[8] Tile_X3Y11_LUT4AB/S4END[9]
+ Tile_X3Y12_LUT4AB/SS4END[0] Tile_X3Y12_LUT4AB/SS4END[10] Tile_X3Y12_LUT4AB/SS4END[11]
+ Tile_X3Y12_LUT4AB/SS4END[12] Tile_X3Y12_LUT4AB/SS4END[13] Tile_X3Y12_LUT4AB/SS4END[14]
+ Tile_X3Y12_LUT4AB/SS4END[15] Tile_X3Y12_LUT4AB/SS4END[1] Tile_X3Y12_LUT4AB/SS4END[2]
+ Tile_X3Y12_LUT4AB/SS4END[3] Tile_X3Y12_LUT4AB/SS4END[4] Tile_X3Y12_LUT4AB/SS4END[5]
+ Tile_X3Y12_LUT4AB/SS4END[6] Tile_X3Y12_LUT4AB/SS4END[7] Tile_X3Y12_LUT4AB/SS4END[8]
+ Tile_X3Y12_LUT4AB/SS4END[9] Tile_X3Y11_LUT4AB/SS4END[0] Tile_X3Y11_LUT4AB/SS4END[10]
+ Tile_X3Y11_LUT4AB/SS4END[11] Tile_X3Y11_LUT4AB/SS4END[12] Tile_X3Y11_LUT4AB/SS4END[13]
+ Tile_X3Y11_LUT4AB/SS4END[14] Tile_X3Y11_LUT4AB/SS4END[15] Tile_X3Y11_LUT4AB/SS4END[1]
+ Tile_X3Y11_LUT4AB/SS4END[2] Tile_X3Y11_LUT4AB/SS4END[3] Tile_X3Y11_LUT4AB/SS4END[4]
+ Tile_X3Y11_LUT4AB/SS4END[5] Tile_X3Y11_LUT4AB/SS4END[6] Tile_X3Y11_LUT4AB/SS4END[7]
+ Tile_X3Y11_LUT4AB/SS4END[8] Tile_X3Y11_LUT4AB/SS4END[9] Tile_X3Y11_LUT4AB/UserCLK
+ Tile_X3Y10_LUT4AB/UserCLK VGND VPWR Tile_X3Y11_LUT4AB/W1BEG[0] Tile_X3Y11_LUT4AB/W1BEG[1]
+ Tile_X3Y11_LUT4AB/W1BEG[2] Tile_X3Y11_LUT4AB/W1BEG[3] Tile_X3Y11_LUT4AB/W1END[0]
+ Tile_X3Y11_LUT4AB/W1END[1] Tile_X3Y11_LUT4AB/W1END[2] Tile_X3Y11_LUT4AB/W1END[3]
+ Tile_X3Y11_LUT4AB/W2BEG[0] Tile_X3Y11_LUT4AB/W2BEG[1] Tile_X3Y11_LUT4AB/W2BEG[2]
+ Tile_X3Y11_LUT4AB/W2BEG[3] Tile_X3Y11_LUT4AB/W2BEG[4] Tile_X3Y11_LUT4AB/W2BEG[5]
+ Tile_X3Y11_LUT4AB/W2BEG[6] Tile_X3Y11_LUT4AB/W2BEG[7] Tile_X2Y11_LUT4AB/W2END[0]
+ Tile_X2Y11_LUT4AB/W2END[1] Tile_X2Y11_LUT4AB/W2END[2] Tile_X2Y11_LUT4AB/W2END[3]
+ Tile_X2Y11_LUT4AB/W2END[4] Tile_X2Y11_LUT4AB/W2END[5] Tile_X2Y11_LUT4AB/W2END[6]
+ Tile_X2Y11_LUT4AB/W2END[7] Tile_X3Y11_LUT4AB/W2END[0] Tile_X3Y11_LUT4AB/W2END[1]
+ Tile_X3Y11_LUT4AB/W2END[2] Tile_X3Y11_LUT4AB/W2END[3] Tile_X3Y11_LUT4AB/W2END[4]
+ Tile_X3Y11_LUT4AB/W2END[5] Tile_X3Y11_LUT4AB/W2END[6] Tile_X3Y11_LUT4AB/W2END[7]
+ Tile_X3Y11_LUT4AB/W2MID[0] Tile_X3Y11_LUT4AB/W2MID[1] Tile_X3Y11_LUT4AB/W2MID[2]
+ Tile_X3Y11_LUT4AB/W2MID[3] Tile_X3Y11_LUT4AB/W2MID[4] Tile_X3Y11_LUT4AB/W2MID[5]
+ Tile_X3Y11_LUT4AB/W2MID[6] Tile_X3Y11_LUT4AB/W2MID[7] Tile_X3Y11_LUT4AB/W6BEG[0]
+ Tile_X3Y11_LUT4AB/W6BEG[10] Tile_X3Y11_LUT4AB/W6BEG[11] Tile_X3Y11_LUT4AB/W6BEG[1]
+ Tile_X3Y11_LUT4AB/W6BEG[2] Tile_X3Y11_LUT4AB/W6BEG[3] Tile_X3Y11_LUT4AB/W6BEG[4]
+ Tile_X3Y11_LUT4AB/W6BEG[5] Tile_X3Y11_LUT4AB/W6BEG[6] Tile_X3Y11_LUT4AB/W6BEG[7]
+ Tile_X3Y11_LUT4AB/W6BEG[8] Tile_X3Y11_LUT4AB/W6BEG[9] Tile_X3Y11_LUT4AB/W6END[0]
+ Tile_X3Y11_LUT4AB/W6END[10] Tile_X3Y11_LUT4AB/W6END[11] Tile_X3Y11_LUT4AB/W6END[1]
+ Tile_X3Y11_LUT4AB/W6END[2] Tile_X3Y11_LUT4AB/W6END[3] Tile_X3Y11_LUT4AB/W6END[4]
+ Tile_X3Y11_LUT4AB/W6END[5] Tile_X3Y11_LUT4AB/W6END[6] Tile_X3Y11_LUT4AB/W6END[7]
+ Tile_X3Y11_LUT4AB/W6END[8] Tile_X3Y11_LUT4AB/W6END[9] Tile_X3Y11_LUT4AB/WW4BEG[0]
+ Tile_X3Y11_LUT4AB/WW4BEG[10] Tile_X3Y11_LUT4AB/WW4BEG[11] Tile_X3Y11_LUT4AB/WW4BEG[12]
+ Tile_X3Y11_LUT4AB/WW4BEG[13] Tile_X3Y11_LUT4AB/WW4BEG[14] Tile_X3Y11_LUT4AB/WW4BEG[15]
+ Tile_X3Y11_LUT4AB/WW4BEG[1] Tile_X3Y11_LUT4AB/WW4BEG[2] Tile_X3Y11_LUT4AB/WW4BEG[3]
+ Tile_X3Y11_LUT4AB/WW4BEG[4] Tile_X3Y11_LUT4AB/WW4BEG[5] Tile_X3Y11_LUT4AB/WW4BEG[6]
+ Tile_X3Y11_LUT4AB/WW4BEG[7] Tile_X3Y11_LUT4AB/WW4BEG[8] Tile_X3Y11_LUT4AB/WW4BEG[9]
+ Tile_X3Y11_LUT4AB/WW4END[0] Tile_X3Y11_LUT4AB/WW4END[10] Tile_X3Y11_LUT4AB/WW4END[11]
+ Tile_X3Y11_LUT4AB/WW4END[12] Tile_X3Y11_LUT4AB/WW4END[13] Tile_X3Y11_LUT4AB/WW4END[14]
+ Tile_X3Y11_LUT4AB/WW4END[15] Tile_X3Y11_LUT4AB/WW4END[1] Tile_X3Y11_LUT4AB/WW4END[2]
+ Tile_X3Y11_LUT4AB/WW4END[3] Tile_X3Y11_LUT4AB/WW4END[4] Tile_X3Y11_LUT4AB/WW4END[5]
+ Tile_X3Y11_LUT4AB/WW4END[6] Tile_X3Y11_LUT4AB/WW4END[7] Tile_X3Y11_LUT4AB/WW4END[8]
+ Tile_X3Y11_LUT4AB/WW4END[9] LUT4AB
XTile_X10Y5_IHP_SRAM Tile_X10Y6_ADDR_SRAM0 Tile_X10Y6_ADDR_SRAM1 Tile_X10Y6_ADDR_SRAM2
+ Tile_X10Y6_ADDR_SRAM3 Tile_X10Y6_ADDR_SRAM4 Tile_X10Y6_ADDR_SRAM5 Tile_X10Y6_ADDR_SRAM6
+ Tile_X10Y6_ADDR_SRAM7 Tile_X10Y6_ADDR_SRAM8 Tile_X10Y6_ADDR_SRAM9 Tile_X10Y6_BM_SRAM0
+ Tile_X10Y6_BM_SRAM1 Tile_X10Y6_BM_SRAM10 Tile_X10Y6_BM_SRAM11 Tile_X10Y6_BM_SRAM12
+ Tile_X10Y6_BM_SRAM13 Tile_X10Y6_BM_SRAM14 Tile_X10Y6_BM_SRAM15 Tile_X10Y6_BM_SRAM16
+ Tile_X10Y6_BM_SRAM17 Tile_X10Y6_BM_SRAM18 Tile_X10Y6_BM_SRAM19 Tile_X10Y6_BM_SRAM2
+ Tile_X10Y6_BM_SRAM20 Tile_X10Y6_BM_SRAM21 Tile_X10Y6_BM_SRAM22 Tile_X10Y6_BM_SRAM23
+ Tile_X10Y6_BM_SRAM24 Tile_X10Y6_BM_SRAM25 Tile_X10Y6_BM_SRAM26 Tile_X10Y6_BM_SRAM27
+ Tile_X10Y6_BM_SRAM28 Tile_X10Y6_BM_SRAM29 Tile_X10Y6_BM_SRAM3 Tile_X10Y6_BM_SRAM30
+ Tile_X10Y6_BM_SRAM31 Tile_X10Y6_BM_SRAM4 Tile_X10Y6_BM_SRAM5 Tile_X10Y6_BM_SRAM6
+ Tile_X10Y6_BM_SRAM7 Tile_X10Y6_BM_SRAM8 Tile_X10Y6_BM_SRAM9 Tile_X10Y6_CLK_SRAM
+ Tile_X10Y6_CONFIGURED_top Tile_X10Y6_DIN_SRAM0 Tile_X10Y6_DIN_SRAM1 Tile_X10Y6_DIN_SRAM10
+ Tile_X10Y6_DIN_SRAM11 Tile_X10Y6_DIN_SRAM12 Tile_X10Y6_DIN_SRAM13 Tile_X10Y6_DIN_SRAM14
+ Tile_X10Y6_DIN_SRAM15 Tile_X10Y6_DIN_SRAM16 Tile_X10Y6_DIN_SRAM17 Tile_X10Y6_DIN_SRAM18
+ Tile_X10Y6_DIN_SRAM19 Tile_X10Y6_DIN_SRAM2 Tile_X10Y6_DIN_SRAM20 Tile_X10Y6_DIN_SRAM21
+ Tile_X10Y6_DIN_SRAM22 Tile_X10Y6_DIN_SRAM23 Tile_X10Y6_DIN_SRAM24 Tile_X10Y6_DIN_SRAM25
+ Tile_X10Y6_DIN_SRAM26 Tile_X10Y6_DIN_SRAM27 Tile_X10Y6_DIN_SRAM28 Tile_X10Y6_DIN_SRAM29
+ Tile_X10Y6_DIN_SRAM3 Tile_X10Y6_DIN_SRAM30 Tile_X10Y6_DIN_SRAM31 Tile_X10Y6_DIN_SRAM4
+ Tile_X10Y6_DIN_SRAM5 Tile_X10Y6_DIN_SRAM6 Tile_X10Y6_DIN_SRAM7 Tile_X10Y6_DIN_SRAM8
+ Tile_X10Y6_DIN_SRAM9 Tile_X10Y6_DOUT_SRAM0 Tile_X10Y6_DOUT_SRAM1 Tile_X10Y6_DOUT_SRAM10
+ Tile_X10Y6_DOUT_SRAM11 Tile_X10Y6_DOUT_SRAM12 Tile_X10Y6_DOUT_SRAM13 Tile_X10Y6_DOUT_SRAM14
+ Tile_X10Y6_DOUT_SRAM15 Tile_X10Y6_DOUT_SRAM16 Tile_X10Y6_DOUT_SRAM17 Tile_X10Y6_DOUT_SRAM18
+ Tile_X10Y6_DOUT_SRAM19 Tile_X10Y6_DOUT_SRAM2 Tile_X10Y6_DOUT_SRAM20 Tile_X10Y6_DOUT_SRAM21
+ Tile_X10Y6_DOUT_SRAM22 Tile_X10Y6_DOUT_SRAM23 Tile_X10Y6_DOUT_SRAM24 Tile_X10Y6_DOUT_SRAM25
+ Tile_X10Y6_DOUT_SRAM26 Tile_X10Y6_DOUT_SRAM27 Tile_X10Y6_DOUT_SRAM28 Tile_X10Y6_DOUT_SRAM29
+ Tile_X10Y6_DOUT_SRAM3 Tile_X10Y6_DOUT_SRAM30 Tile_X10Y6_DOUT_SRAM31 Tile_X10Y6_DOUT_SRAM4
+ Tile_X10Y6_DOUT_SRAM5 Tile_X10Y6_DOUT_SRAM6 Tile_X10Y6_DOUT_SRAM7 Tile_X10Y6_DOUT_SRAM8
+ Tile_X10Y6_DOUT_SRAM9 Tile_X10Y6_MEN_SRAM Tile_X10Y6_REN_SRAM Tile_X10Y6_TIE_HIGH_SRAM
+ Tile_X10Y6_TIE_LOW_SRAM Tile_X9Y5_LUT4AB/E1BEG[0] Tile_X9Y5_LUT4AB/E1BEG[1] Tile_X9Y5_LUT4AB/E1BEG[2]
+ Tile_X9Y5_LUT4AB/E1BEG[3] Tile_X9Y5_LUT4AB/E2BEGb[0] Tile_X9Y5_LUT4AB/E2BEGb[1]
+ Tile_X9Y5_LUT4AB/E2BEGb[2] Tile_X9Y5_LUT4AB/E2BEGb[3] Tile_X9Y5_LUT4AB/E2BEGb[4]
+ Tile_X9Y5_LUT4AB/E2BEGb[5] Tile_X9Y5_LUT4AB/E2BEGb[6] Tile_X9Y5_LUT4AB/E2BEGb[7]
+ Tile_X9Y5_LUT4AB/E2BEG[0] Tile_X9Y5_LUT4AB/E2BEG[1] Tile_X9Y5_LUT4AB/E2BEG[2] Tile_X9Y5_LUT4AB/E2BEG[3]
+ Tile_X9Y5_LUT4AB/E2BEG[4] Tile_X9Y5_LUT4AB/E2BEG[5] Tile_X9Y5_LUT4AB/E2BEG[6] Tile_X9Y5_LUT4AB/E2BEG[7]
+ Tile_X9Y5_LUT4AB/E6BEG[0] Tile_X9Y5_LUT4AB/E6BEG[10] Tile_X9Y5_LUT4AB/E6BEG[11]
+ Tile_X9Y5_LUT4AB/E6BEG[1] Tile_X9Y5_LUT4AB/E6BEG[2] Tile_X9Y5_LUT4AB/E6BEG[3] Tile_X9Y5_LUT4AB/E6BEG[4]
+ Tile_X9Y5_LUT4AB/E6BEG[5] Tile_X9Y5_LUT4AB/E6BEG[6] Tile_X9Y5_LUT4AB/E6BEG[7] Tile_X9Y5_LUT4AB/E6BEG[8]
+ Tile_X9Y5_LUT4AB/E6BEG[9] Tile_X9Y5_LUT4AB/EE4BEG[0] Tile_X9Y5_LUT4AB/EE4BEG[10]
+ Tile_X9Y5_LUT4AB/EE4BEG[11] Tile_X9Y5_LUT4AB/EE4BEG[12] Tile_X9Y5_LUT4AB/EE4BEG[13]
+ Tile_X9Y5_LUT4AB/EE4BEG[14] Tile_X9Y5_LUT4AB/EE4BEG[15] Tile_X9Y5_LUT4AB/EE4BEG[1]
+ Tile_X9Y5_LUT4AB/EE4BEG[2] Tile_X9Y5_LUT4AB/EE4BEG[3] Tile_X9Y5_LUT4AB/EE4BEG[4]
+ Tile_X9Y5_LUT4AB/EE4BEG[5] Tile_X9Y5_LUT4AB/EE4BEG[6] Tile_X9Y5_LUT4AB/EE4BEG[7]
+ Tile_X9Y5_LUT4AB/EE4BEG[8] Tile_X9Y5_LUT4AB/EE4BEG[9] Tile_X9Y5_LUT4AB/FrameData_O[0]
+ Tile_X9Y5_LUT4AB/FrameData_O[10] Tile_X9Y5_LUT4AB/FrameData_O[11] Tile_X9Y5_LUT4AB/FrameData_O[12]
+ Tile_X9Y5_LUT4AB/FrameData_O[13] Tile_X9Y5_LUT4AB/FrameData_O[14] Tile_X9Y5_LUT4AB/FrameData_O[15]
+ Tile_X9Y5_LUT4AB/FrameData_O[16] Tile_X9Y5_LUT4AB/FrameData_O[17] Tile_X9Y5_LUT4AB/FrameData_O[18]
+ Tile_X9Y5_LUT4AB/FrameData_O[19] Tile_X9Y5_LUT4AB/FrameData_O[1] Tile_X9Y5_LUT4AB/FrameData_O[20]
+ Tile_X9Y5_LUT4AB/FrameData_O[21] Tile_X9Y5_LUT4AB/FrameData_O[22] Tile_X9Y5_LUT4AB/FrameData_O[23]
+ Tile_X9Y5_LUT4AB/FrameData_O[24] Tile_X9Y5_LUT4AB/FrameData_O[25] Tile_X9Y5_LUT4AB/FrameData_O[26]
+ Tile_X9Y5_LUT4AB/FrameData_O[27] Tile_X9Y5_LUT4AB/FrameData_O[28] Tile_X9Y5_LUT4AB/FrameData_O[29]
+ Tile_X9Y5_LUT4AB/FrameData_O[2] Tile_X9Y5_LUT4AB/FrameData_O[30] Tile_X9Y5_LUT4AB/FrameData_O[31]
+ Tile_X9Y5_LUT4AB/FrameData_O[3] Tile_X9Y5_LUT4AB/FrameData_O[4] Tile_X9Y5_LUT4AB/FrameData_O[5]
+ Tile_X9Y5_LUT4AB/FrameData_O[6] Tile_X9Y5_LUT4AB/FrameData_O[7] Tile_X9Y5_LUT4AB/FrameData_O[8]
+ Tile_X9Y5_LUT4AB/FrameData_O[9] Tile_X10Y5_IHP_SRAM/Tile_X0Y0_FrameData_O[0] Tile_X10Y5_IHP_SRAM/Tile_X0Y0_FrameData_O[10]
+ Tile_X10Y5_IHP_SRAM/Tile_X0Y0_FrameData_O[11] Tile_X10Y5_IHP_SRAM/Tile_X0Y0_FrameData_O[12]
+ Tile_X10Y5_IHP_SRAM/Tile_X0Y0_FrameData_O[13] Tile_X10Y5_IHP_SRAM/Tile_X0Y0_FrameData_O[14]
+ Tile_X10Y5_IHP_SRAM/Tile_X0Y0_FrameData_O[15] Tile_X10Y5_IHP_SRAM/Tile_X0Y0_FrameData_O[16]
+ Tile_X10Y5_IHP_SRAM/Tile_X0Y0_FrameData_O[17] Tile_X10Y5_IHP_SRAM/Tile_X0Y0_FrameData_O[18]
+ Tile_X10Y5_IHP_SRAM/Tile_X0Y0_FrameData_O[19] Tile_X10Y5_IHP_SRAM/Tile_X0Y0_FrameData_O[1]
+ Tile_X10Y5_IHP_SRAM/Tile_X0Y0_FrameData_O[20] Tile_X10Y5_IHP_SRAM/Tile_X0Y0_FrameData_O[21]
+ Tile_X10Y5_IHP_SRAM/Tile_X0Y0_FrameData_O[22] Tile_X10Y5_IHP_SRAM/Tile_X0Y0_FrameData_O[23]
+ Tile_X10Y5_IHP_SRAM/Tile_X0Y0_FrameData_O[24] Tile_X10Y5_IHP_SRAM/Tile_X0Y0_FrameData_O[25]
+ Tile_X10Y5_IHP_SRAM/Tile_X0Y0_FrameData_O[26] Tile_X10Y5_IHP_SRAM/Tile_X0Y0_FrameData_O[27]
+ Tile_X10Y5_IHP_SRAM/Tile_X0Y0_FrameData_O[28] Tile_X10Y5_IHP_SRAM/Tile_X0Y0_FrameData_O[29]
+ Tile_X10Y5_IHP_SRAM/Tile_X0Y0_FrameData_O[2] Tile_X10Y5_IHP_SRAM/Tile_X0Y0_FrameData_O[30]
+ Tile_X10Y5_IHP_SRAM/Tile_X0Y0_FrameData_O[31] Tile_X10Y5_IHP_SRAM/Tile_X0Y0_FrameData_O[3]
+ Tile_X10Y5_IHP_SRAM/Tile_X0Y0_FrameData_O[4] Tile_X10Y5_IHP_SRAM/Tile_X0Y0_FrameData_O[5]
+ Tile_X10Y5_IHP_SRAM/Tile_X0Y0_FrameData_O[6] Tile_X10Y5_IHP_SRAM/Tile_X0Y0_FrameData_O[7]
+ Tile_X10Y5_IHP_SRAM/Tile_X0Y0_FrameData_O[8] Tile_X10Y5_IHP_SRAM/Tile_X0Y0_FrameData_O[9]
+ Tile_X10Y3_IHP_SRAM/Tile_X0Y1_FrameStrobe[0] Tile_X10Y3_IHP_SRAM/Tile_X0Y1_FrameStrobe[10]
+ Tile_X10Y3_IHP_SRAM/Tile_X0Y1_FrameStrobe[11] Tile_X10Y3_IHP_SRAM/Tile_X0Y1_FrameStrobe[12]
+ Tile_X10Y3_IHP_SRAM/Tile_X0Y1_FrameStrobe[13] Tile_X10Y3_IHP_SRAM/Tile_X0Y1_FrameStrobe[14]
+ Tile_X10Y3_IHP_SRAM/Tile_X0Y1_FrameStrobe[15] Tile_X10Y3_IHP_SRAM/Tile_X0Y1_FrameStrobe[16]
+ Tile_X10Y3_IHP_SRAM/Tile_X0Y1_FrameStrobe[17] Tile_X10Y3_IHP_SRAM/Tile_X0Y1_FrameStrobe[18]
+ Tile_X10Y3_IHP_SRAM/Tile_X0Y1_FrameStrobe[19] Tile_X10Y3_IHP_SRAM/Tile_X0Y1_FrameStrobe[1]
+ Tile_X10Y3_IHP_SRAM/Tile_X0Y1_FrameStrobe[2] Tile_X10Y3_IHP_SRAM/Tile_X0Y1_FrameStrobe[3]
+ Tile_X10Y3_IHP_SRAM/Tile_X0Y1_FrameStrobe[4] Tile_X10Y3_IHP_SRAM/Tile_X0Y1_FrameStrobe[5]
+ Tile_X10Y3_IHP_SRAM/Tile_X0Y1_FrameStrobe[6] Tile_X10Y3_IHP_SRAM/Tile_X0Y1_FrameStrobe[7]
+ Tile_X10Y3_IHP_SRAM/Tile_X0Y1_FrameStrobe[8] Tile_X10Y3_IHP_SRAM/Tile_X0Y1_FrameStrobe[9]
+ Tile_X10Y5_IHP_SRAM/Tile_X0Y0_N1BEG[0] Tile_X10Y5_IHP_SRAM/Tile_X0Y0_N1BEG[1] Tile_X10Y5_IHP_SRAM/Tile_X0Y0_N1BEG[2]
+ Tile_X10Y5_IHP_SRAM/Tile_X0Y0_N1BEG[3] Tile_X10Y5_IHP_SRAM/Tile_X0Y0_N2BEG[0] Tile_X10Y5_IHP_SRAM/Tile_X0Y0_N2BEG[1]
+ Tile_X10Y5_IHP_SRAM/Tile_X0Y0_N2BEG[2] Tile_X10Y5_IHP_SRAM/Tile_X0Y0_N2BEG[3] Tile_X10Y5_IHP_SRAM/Tile_X0Y0_N2BEG[4]
+ Tile_X10Y5_IHP_SRAM/Tile_X0Y0_N2BEG[5] Tile_X10Y5_IHP_SRAM/Tile_X0Y0_N2BEG[6] Tile_X10Y5_IHP_SRAM/Tile_X0Y0_N2BEG[7]
+ Tile_X10Y3_IHP_SRAM/Tile_X0Y1_N2END[0] Tile_X10Y3_IHP_SRAM/Tile_X0Y1_N2END[1] Tile_X10Y3_IHP_SRAM/Tile_X0Y1_N2END[2]
+ Tile_X10Y3_IHP_SRAM/Tile_X0Y1_N2END[3] Tile_X10Y3_IHP_SRAM/Tile_X0Y1_N2END[4] Tile_X10Y3_IHP_SRAM/Tile_X0Y1_N2END[5]
+ Tile_X10Y3_IHP_SRAM/Tile_X0Y1_N2END[6] Tile_X10Y3_IHP_SRAM/Tile_X0Y1_N2END[7] Tile_X10Y5_IHP_SRAM/Tile_X0Y0_N4BEG[0]
+ Tile_X10Y5_IHP_SRAM/Tile_X0Y0_N4BEG[10] Tile_X10Y5_IHP_SRAM/Tile_X0Y0_N4BEG[11]
+ Tile_X10Y5_IHP_SRAM/Tile_X0Y0_N4BEG[12] Tile_X10Y5_IHP_SRAM/Tile_X0Y0_N4BEG[13]
+ Tile_X10Y5_IHP_SRAM/Tile_X0Y0_N4BEG[14] Tile_X10Y5_IHP_SRAM/Tile_X0Y0_N4BEG[15]
+ Tile_X10Y5_IHP_SRAM/Tile_X0Y0_N4BEG[1] Tile_X10Y5_IHP_SRAM/Tile_X0Y0_N4BEG[2] Tile_X10Y5_IHP_SRAM/Tile_X0Y0_N4BEG[3]
+ Tile_X10Y5_IHP_SRAM/Tile_X0Y0_N4BEG[4] Tile_X10Y5_IHP_SRAM/Tile_X0Y0_N4BEG[5] Tile_X10Y5_IHP_SRAM/Tile_X0Y0_N4BEG[6]
+ Tile_X10Y5_IHP_SRAM/Tile_X0Y0_N4BEG[7] Tile_X10Y5_IHP_SRAM/Tile_X0Y0_N4BEG[8] Tile_X10Y5_IHP_SRAM/Tile_X0Y0_N4BEG[9]
+ Tile_X10Y5_IHP_SRAM/Tile_X0Y0_S1END[0] Tile_X10Y5_IHP_SRAM/Tile_X0Y0_S1END[1] Tile_X10Y5_IHP_SRAM/Tile_X0Y0_S1END[2]
+ Tile_X10Y5_IHP_SRAM/Tile_X0Y0_S1END[3] Tile_X10Y5_IHP_SRAM/Tile_X0Y0_S2END[0] Tile_X10Y5_IHP_SRAM/Tile_X0Y0_S2END[1]
+ Tile_X10Y5_IHP_SRAM/Tile_X0Y0_S2END[2] Tile_X10Y5_IHP_SRAM/Tile_X0Y0_S2END[3] Tile_X10Y5_IHP_SRAM/Tile_X0Y0_S2END[4]
+ Tile_X10Y5_IHP_SRAM/Tile_X0Y0_S2END[5] Tile_X10Y5_IHP_SRAM/Tile_X0Y0_S2END[6] Tile_X10Y5_IHP_SRAM/Tile_X0Y0_S2END[7]
+ Tile_X10Y5_IHP_SRAM/Tile_X0Y0_S2MID[0] Tile_X10Y5_IHP_SRAM/Tile_X0Y0_S2MID[1] Tile_X10Y5_IHP_SRAM/Tile_X0Y0_S2MID[2]
+ Tile_X10Y5_IHP_SRAM/Tile_X0Y0_S2MID[3] Tile_X10Y5_IHP_SRAM/Tile_X0Y0_S2MID[4] Tile_X10Y5_IHP_SRAM/Tile_X0Y0_S2MID[5]
+ Tile_X10Y5_IHP_SRAM/Tile_X0Y0_S2MID[6] Tile_X10Y5_IHP_SRAM/Tile_X0Y0_S2MID[7] Tile_X10Y5_IHP_SRAM/Tile_X0Y0_S4END[0]
+ Tile_X10Y5_IHP_SRAM/Tile_X0Y0_S4END[10] Tile_X10Y5_IHP_SRAM/Tile_X0Y0_S4END[11]
+ Tile_X10Y5_IHP_SRAM/Tile_X0Y0_S4END[12] Tile_X10Y5_IHP_SRAM/Tile_X0Y0_S4END[13]
+ Tile_X10Y5_IHP_SRAM/Tile_X0Y0_S4END[14] Tile_X10Y5_IHP_SRAM/Tile_X0Y0_S4END[15]
+ Tile_X10Y5_IHP_SRAM/Tile_X0Y0_S4END[1] Tile_X10Y5_IHP_SRAM/Tile_X0Y0_S4END[2] Tile_X10Y5_IHP_SRAM/Tile_X0Y0_S4END[3]
+ Tile_X10Y5_IHP_SRAM/Tile_X0Y0_S4END[4] Tile_X10Y5_IHP_SRAM/Tile_X0Y0_S4END[5] Tile_X10Y5_IHP_SRAM/Tile_X0Y0_S4END[6]
+ Tile_X10Y5_IHP_SRAM/Tile_X0Y0_S4END[7] Tile_X10Y5_IHP_SRAM/Tile_X0Y0_S4END[8] Tile_X10Y5_IHP_SRAM/Tile_X0Y0_S4END[9]
+ Tile_X10Y3_IHP_SRAM/Tile_X0Y1_UserCLK Tile_X9Y5_LUT4AB/W1END[0] Tile_X9Y5_LUT4AB/W1END[1]
+ Tile_X9Y5_LUT4AB/W1END[2] Tile_X9Y5_LUT4AB/W1END[3] Tile_X9Y5_LUT4AB/W2MID[0] Tile_X9Y5_LUT4AB/W2MID[1]
+ Tile_X9Y5_LUT4AB/W2MID[2] Tile_X9Y5_LUT4AB/W2MID[3] Tile_X9Y5_LUT4AB/W2MID[4] Tile_X9Y5_LUT4AB/W2MID[5]
+ Tile_X9Y5_LUT4AB/W2MID[6] Tile_X9Y5_LUT4AB/W2MID[7] Tile_X9Y5_LUT4AB/W2END[0] Tile_X9Y5_LUT4AB/W2END[1]
+ Tile_X9Y5_LUT4AB/W2END[2] Tile_X9Y5_LUT4AB/W2END[3] Tile_X9Y5_LUT4AB/W2END[4] Tile_X9Y5_LUT4AB/W2END[5]
+ Tile_X9Y5_LUT4AB/W2END[6] Tile_X9Y5_LUT4AB/W2END[7] Tile_X9Y5_LUT4AB/W6END[0] Tile_X9Y5_LUT4AB/W6END[10]
+ Tile_X9Y5_LUT4AB/W6END[11] Tile_X9Y5_LUT4AB/W6END[1] Tile_X9Y5_LUT4AB/W6END[2] Tile_X9Y5_LUT4AB/W6END[3]
+ Tile_X9Y5_LUT4AB/W6END[4] Tile_X9Y5_LUT4AB/W6END[5] Tile_X9Y5_LUT4AB/W6END[6] Tile_X9Y5_LUT4AB/W6END[7]
+ Tile_X9Y5_LUT4AB/W6END[8] Tile_X9Y5_LUT4AB/W6END[9] Tile_X9Y5_LUT4AB/WW4END[0] Tile_X9Y5_LUT4AB/WW4END[10]
+ Tile_X9Y5_LUT4AB/WW4END[11] Tile_X9Y5_LUT4AB/WW4END[12] Tile_X9Y5_LUT4AB/WW4END[13]
+ Tile_X9Y5_LUT4AB/WW4END[14] Tile_X9Y5_LUT4AB/WW4END[15] Tile_X9Y5_LUT4AB/WW4END[1]
+ Tile_X9Y5_LUT4AB/WW4END[2] Tile_X9Y5_LUT4AB/WW4END[3] Tile_X9Y5_LUT4AB/WW4END[4]
+ Tile_X9Y5_LUT4AB/WW4END[5] Tile_X9Y5_LUT4AB/WW4END[6] Tile_X9Y5_LUT4AB/WW4END[7]
+ Tile_X9Y5_LUT4AB/WW4END[8] Tile_X9Y5_LUT4AB/WW4END[9] Tile_X9Y6_LUT4AB/E1BEG[0]
+ Tile_X9Y6_LUT4AB/E1BEG[1] Tile_X9Y6_LUT4AB/E1BEG[2] Tile_X9Y6_LUT4AB/E1BEG[3] Tile_X9Y6_LUT4AB/E2BEGb[0]
+ Tile_X9Y6_LUT4AB/E2BEGb[1] Tile_X9Y6_LUT4AB/E2BEGb[2] Tile_X9Y6_LUT4AB/E2BEGb[3]
+ Tile_X9Y6_LUT4AB/E2BEGb[4] Tile_X9Y6_LUT4AB/E2BEGb[5] Tile_X9Y6_LUT4AB/E2BEGb[6]
+ Tile_X9Y6_LUT4AB/E2BEGb[7] Tile_X9Y6_LUT4AB/E2BEG[0] Tile_X9Y6_LUT4AB/E2BEG[1] Tile_X9Y6_LUT4AB/E2BEG[2]
+ Tile_X9Y6_LUT4AB/E2BEG[3] Tile_X9Y6_LUT4AB/E2BEG[4] Tile_X9Y6_LUT4AB/E2BEG[5] Tile_X9Y6_LUT4AB/E2BEG[6]
+ Tile_X9Y6_LUT4AB/E2BEG[7] Tile_X9Y6_LUT4AB/E6BEG[0] Tile_X9Y6_LUT4AB/E6BEG[10] Tile_X9Y6_LUT4AB/E6BEG[11]
+ Tile_X9Y6_LUT4AB/E6BEG[1] Tile_X9Y6_LUT4AB/E6BEG[2] Tile_X9Y6_LUT4AB/E6BEG[3] Tile_X9Y6_LUT4AB/E6BEG[4]
+ Tile_X9Y6_LUT4AB/E6BEG[5] Tile_X9Y6_LUT4AB/E6BEG[6] Tile_X9Y6_LUT4AB/E6BEG[7] Tile_X9Y6_LUT4AB/E6BEG[8]
+ Tile_X9Y6_LUT4AB/E6BEG[9] Tile_X9Y6_LUT4AB/EE4BEG[0] Tile_X9Y6_LUT4AB/EE4BEG[10]
+ Tile_X9Y6_LUT4AB/EE4BEG[11] Tile_X9Y6_LUT4AB/EE4BEG[12] Tile_X9Y6_LUT4AB/EE4BEG[13]
+ Tile_X9Y6_LUT4AB/EE4BEG[14] Tile_X9Y6_LUT4AB/EE4BEG[15] Tile_X9Y6_LUT4AB/EE4BEG[1]
+ Tile_X9Y6_LUT4AB/EE4BEG[2] Tile_X9Y6_LUT4AB/EE4BEG[3] Tile_X9Y6_LUT4AB/EE4BEG[4]
+ Tile_X9Y6_LUT4AB/EE4BEG[5] Tile_X9Y6_LUT4AB/EE4BEG[6] Tile_X9Y6_LUT4AB/EE4BEG[7]
+ Tile_X9Y6_LUT4AB/EE4BEG[8] Tile_X9Y6_LUT4AB/EE4BEG[9] Tile_X9Y6_LUT4AB/FrameData_O[0]
+ Tile_X9Y6_LUT4AB/FrameData_O[10] Tile_X9Y6_LUT4AB/FrameData_O[11] Tile_X9Y6_LUT4AB/FrameData_O[12]
+ Tile_X9Y6_LUT4AB/FrameData_O[13] Tile_X9Y6_LUT4AB/FrameData_O[14] Tile_X9Y6_LUT4AB/FrameData_O[15]
+ Tile_X9Y6_LUT4AB/FrameData_O[16] Tile_X9Y6_LUT4AB/FrameData_O[17] Tile_X9Y6_LUT4AB/FrameData_O[18]
+ Tile_X9Y6_LUT4AB/FrameData_O[19] Tile_X9Y6_LUT4AB/FrameData_O[1] Tile_X9Y6_LUT4AB/FrameData_O[20]
+ Tile_X9Y6_LUT4AB/FrameData_O[21] Tile_X9Y6_LUT4AB/FrameData_O[22] Tile_X9Y6_LUT4AB/FrameData_O[23]
+ Tile_X9Y6_LUT4AB/FrameData_O[24] Tile_X9Y6_LUT4AB/FrameData_O[25] Tile_X9Y6_LUT4AB/FrameData_O[26]
+ Tile_X9Y6_LUT4AB/FrameData_O[27] Tile_X9Y6_LUT4AB/FrameData_O[28] Tile_X9Y6_LUT4AB/FrameData_O[29]
+ Tile_X9Y6_LUT4AB/FrameData_O[2] Tile_X9Y6_LUT4AB/FrameData_O[30] Tile_X9Y6_LUT4AB/FrameData_O[31]
+ Tile_X9Y6_LUT4AB/FrameData_O[3] Tile_X9Y6_LUT4AB/FrameData_O[4] Tile_X9Y6_LUT4AB/FrameData_O[5]
+ Tile_X9Y6_LUT4AB/FrameData_O[6] Tile_X9Y6_LUT4AB/FrameData_O[7] Tile_X9Y6_LUT4AB/FrameData_O[8]
+ Tile_X9Y6_LUT4AB/FrameData_O[9] Tile_X10Y5_IHP_SRAM/Tile_X0Y1_FrameData_O[0] Tile_X10Y5_IHP_SRAM/Tile_X0Y1_FrameData_O[10]
+ Tile_X10Y5_IHP_SRAM/Tile_X0Y1_FrameData_O[11] Tile_X10Y5_IHP_SRAM/Tile_X0Y1_FrameData_O[12]
+ Tile_X10Y5_IHP_SRAM/Tile_X0Y1_FrameData_O[13] Tile_X10Y5_IHP_SRAM/Tile_X0Y1_FrameData_O[14]
+ Tile_X10Y5_IHP_SRAM/Tile_X0Y1_FrameData_O[15] Tile_X10Y5_IHP_SRAM/Tile_X0Y1_FrameData_O[16]
+ Tile_X10Y5_IHP_SRAM/Tile_X0Y1_FrameData_O[17] Tile_X10Y5_IHP_SRAM/Tile_X0Y1_FrameData_O[18]
+ Tile_X10Y5_IHP_SRAM/Tile_X0Y1_FrameData_O[19] Tile_X10Y5_IHP_SRAM/Tile_X0Y1_FrameData_O[1]
+ Tile_X10Y5_IHP_SRAM/Tile_X0Y1_FrameData_O[20] Tile_X10Y5_IHP_SRAM/Tile_X0Y1_FrameData_O[21]
+ Tile_X10Y5_IHP_SRAM/Tile_X0Y1_FrameData_O[22] Tile_X10Y5_IHP_SRAM/Tile_X0Y1_FrameData_O[23]
+ Tile_X10Y5_IHP_SRAM/Tile_X0Y1_FrameData_O[24] Tile_X10Y5_IHP_SRAM/Tile_X0Y1_FrameData_O[25]
+ Tile_X10Y5_IHP_SRAM/Tile_X0Y1_FrameData_O[26] Tile_X10Y5_IHP_SRAM/Tile_X0Y1_FrameData_O[27]
+ Tile_X10Y5_IHP_SRAM/Tile_X0Y1_FrameData_O[28] Tile_X10Y5_IHP_SRAM/Tile_X0Y1_FrameData_O[29]
+ Tile_X10Y5_IHP_SRAM/Tile_X0Y1_FrameData_O[2] Tile_X10Y5_IHP_SRAM/Tile_X0Y1_FrameData_O[30]
+ Tile_X10Y5_IHP_SRAM/Tile_X0Y1_FrameData_O[31] Tile_X10Y5_IHP_SRAM/Tile_X0Y1_FrameData_O[3]
+ Tile_X10Y5_IHP_SRAM/Tile_X0Y1_FrameData_O[4] Tile_X10Y5_IHP_SRAM/Tile_X0Y1_FrameData_O[5]
+ Tile_X10Y5_IHP_SRAM/Tile_X0Y1_FrameData_O[6] Tile_X10Y5_IHP_SRAM/Tile_X0Y1_FrameData_O[7]
+ Tile_X10Y5_IHP_SRAM/Tile_X0Y1_FrameData_O[8] Tile_X10Y5_IHP_SRAM/Tile_X0Y1_FrameData_O[9]
+ Tile_X10Y5_IHP_SRAM/Tile_X0Y1_FrameStrobe[0] Tile_X10Y5_IHP_SRAM/Tile_X0Y1_FrameStrobe[10]
+ Tile_X10Y5_IHP_SRAM/Tile_X0Y1_FrameStrobe[11] Tile_X10Y5_IHP_SRAM/Tile_X0Y1_FrameStrobe[12]
+ Tile_X10Y5_IHP_SRAM/Tile_X0Y1_FrameStrobe[13] Tile_X10Y5_IHP_SRAM/Tile_X0Y1_FrameStrobe[14]
+ Tile_X10Y5_IHP_SRAM/Tile_X0Y1_FrameStrobe[15] Tile_X10Y5_IHP_SRAM/Tile_X0Y1_FrameStrobe[16]
+ Tile_X10Y5_IHP_SRAM/Tile_X0Y1_FrameStrobe[17] Tile_X10Y5_IHP_SRAM/Tile_X0Y1_FrameStrobe[18]
+ Tile_X10Y5_IHP_SRAM/Tile_X0Y1_FrameStrobe[19] Tile_X10Y5_IHP_SRAM/Tile_X0Y1_FrameStrobe[1]
+ Tile_X10Y5_IHP_SRAM/Tile_X0Y1_FrameStrobe[2] Tile_X10Y5_IHP_SRAM/Tile_X0Y1_FrameStrobe[3]
+ Tile_X10Y5_IHP_SRAM/Tile_X0Y1_FrameStrobe[4] Tile_X10Y5_IHP_SRAM/Tile_X0Y1_FrameStrobe[5]
+ Tile_X10Y5_IHP_SRAM/Tile_X0Y1_FrameStrobe[6] Tile_X10Y5_IHP_SRAM/Tile_X0Y1_FrameStrobe[7]
+ Tile_X10Y5_IHP_SRAM/Tile_X0Y1_FrameStrobe[8] Tile_X10Y5_IHP_SRAM/Tile_X0Y1_FrameStrobe[9]
+ Tile_X10Y7_IHP_SRAM/Tile_X0Y0_N1BEG[0] Tile_X10Y7_IHP_SRAM/Tile_X0Y0_N1BEG[1] Tile_X10Y7_IHP_SRAM/Tile_X0Y0_N1BEG[2]
+ Tile_X10Y7_IHP_SRAM/Tile_X0Y0_N1BEG[3] Tile_X10Y5_IHP_SRAM/Tile_X0Y1_N2END[0] Tile_X10Y5_IHP_SRAM/Tile_X0Y1_N2END[1]
+ Tile_X10Y5_IHP_SRAM/Tile_X0Y1_N2END[2] Tile_X10Y5_IHP_SRAM/Tile_X0Y1_N2END[3] Tile_X10Y5_IHP_SRAM/Tile_X0Y1_N2END[4]
+ Tile_X10Y5_IHP_SRAM/Tile_X0Y1_N2END[5] Tile_X10Y5_IHP_SRAM/Tile_X0Y1_N2END[6] Tile_X10Y5_IHP_SRAM/Tile_X0Y1_N2END[7]
+ Tile_X10Y7_IHP_SRAM/Tile_X0Y0_N2BEG[0] Tile_X10Y7_IHP_SRAM/Tile_X0Y0_N2BEG[1] Tile_X10Y7_IHP_SRAM/Tile_X0Y0_N2BEG[2]
+ Tile_X10Y7_IHP_SRAM/Tile_X0Y0_N2BEG[3] Tile_X10Y7_IHP_SRAM/Tile_X0Y0_N2BEG[4] Tile_X10Y7_IHP_SRAM/Tile_X0Y0_N2BEG[5]
+ Tile_X10Y7_IHP_SRAM/Tile_X0Y0_N2BEG[6] Tile_X10Y7_IHP_SRAM/Tile_X0Y0_N2BEG[7] Tile_X10Y7_IHP_SRAM/Tile_X0Y0_N4BEG[0]
+ Tile_X10Y7_IHP_SRAM/Tile_X0Y0_N4BEG[10] Tile_X10Y7_IHP_SRAM/Tile_X0Y0_N4BEG[11]
+ Tile_X10Y7_IHP_SRAM/Tile_X0Y0_N4BEG[12] Tile_X10Y7_IHP_SRAM/Tile_X0Y0_N4BEG[13]
+ Tile_X10Y7_IHP_SRAM/Tile_X0Y0_N4BEG[14] Tile_X10Y7_IHP_SRAM/Tile_X0Y0_N4BEG[15]
+ Tile_X10Y7_IHP_SRAM/Tile_X0Y0_N4BEG[1] Tile_X10Y7_IHP_SRAM/Tile_X0Y0_N4BEG[2] Tile_X10Y7_IHP_SRAM/Tile_X0Y0_N4BEG[3]
+ Tile_X10Y7_IHP_SRAM/Tile_X0Y0_N4BEG[4] Tile_X10Y7_IHP_SRAM/Tile_X0Y0_N4BEG[5] Tile_X10Y7_IHP_SRAM/Tile_X0Y0_N4BEG[6]
+ Tile_X10Y7_IHP_SRAM/Tile_X0Y0_N4BEG[7] Tile_X10Y7_IHP_SRAM/Tile_X0Y0_N4BEG[8] Tile_X10Y7_IHP_SRAM/Tile_X0Y0_N4BEG[9]
+ Tile_X10Y7_IHP_SRAM/Tile_X0Y0_S1END[0] Tile_X10Y7_IHP_SRAM/Tile_X0Y0_S1END[1] Tile_X10Y7_IHP_SRAM/Tile_X0Y0_S1END[2]
+ Tile_X10Y7_IHP_SRAM/Tile_X0Y0_S1END[3] Tile_X10Y7_IHP_SRAM/Tile_X0Y0_S2MID[0] Tile_X10Y7_IHP_SRAM/Tile_X0Y0_S2MID[1]
+ Tile_X10Y7_IHP_SRAM/Tile_X0Y0_S2MID[2] Tile_X10Y7_IHP_SRAM/Tile_X0Y0_S2MID[3] Tile_X10Y7_IHP_SRAM/Tile_X0Y0_S2MID[4]
+ Tile_X10Y7_IHP_SRAM/Tile_X0Y0_S2MID[5] Tile_X10Y7_IHP_SRAM/Tile_X0Y0_S2MID[6] Tile_X10Y7_IHP_SRAM/Tile_X0Y0_S2MID[7]
+ Tile_X10Y7_IHP_SRAM/Tile_X0Y0_S2END[0] Tile_X10Y7_IHP_SRAM/Tile_X0Y0_S2END[1] Tile_X10Y7_IHP_SRAM/Tile_X0Y0_S2END[2]
+ Tile_X10Y7_IHP_SRAM/Tile_X0Y0_S2END[3] Tile_X10Y7_IHP_SRAM/Tile_X0Y0_S2END[4] Tile_X10Y7_IHP_SRAM/Tile_X0Y0_S2END[5]
+ Tile_X10Y7_IHP_SRAM/Tile_X0Y0_S2END[6] Tile_X10Y7_IHP_SRAM/Tile_X0Y0_S2END[7] Tile_X10Y7_IHP_SRAM/Tile_X0Y0_S4END[0]
+ Tile_X10Y7_IHP_SRAM/Tile_X0Y0_S4END[10] Tile_X10Y7_IHP_SRAM/Tile_X0Y0_S4END[11]
+ Tile_X10Y7_IHP_SRAM/Tile_X0Y0_S4END[12] Tile_X10Y7_IHP_SRAM/Tile_X0Y0_S4END[13]
+ Tile_X10Y7_IHP_SRAM/Tile_X0Y0_S4END[14] Tile_X10Y7_IHP_SRAM/Tile_X0Y0_S4END[15]
+ Tile_X10Y7_IHP_SRAM/Tile_X0Y0_S4END[1] Tile_X10Y7_IHP_SRAM/Tile_X0Y0_S4END[2] Tile_X10Y7_IHP_SRAM/Tile_X0Y0_S4END[3]
+ Tile_X10Y7_IHP_SRAM/Tile_X0Y0_S4END[4] Tile_X10Y7_IHP_SRAM/Tile_X0Y0_S4END[5] Tile_X10Y7_IHP_SRAM/Tile_X0Y0_S4END[6]
+ Tile_X10Y7_IHP_SRAM/Tile_X0Y0_S4END[7] Tile_X10Y7_IHP_SRAM/Tile_X0Y0_S4END[8] Tile_X10Y7_IHP_SRAM/Tile_X0Y0_S4END[9]
+ Tile_X10Y5_IHP_SRAM/Tile_X0Y1_UserCLK Tile_X9Y6_LUT4AB/W1END[0] Tile_X9Y6_LUT4AB/W1END[1]
+ Tile_X9Y6_LUT4AB/W1END[2] Tile_X9Y6_LUT4AB/W1END[3] Tile_X9Y6_LUT4AB/W2MID[0] Tile_X9Y6_LUT4AB/W2MID[1]
+ Tile_X9Y6_LUT4AB/W2MID[2] Tile_X9Y6_LUT4AB/W2MID[3] Tile_X9Y6_LUT4AB/W2MID[4] Tile_X9Y6_LUT4AB/W2MID[5]
+ Tile_X9Y6_LUT4AB/W2MID[6] Tile_X9Y6_LUT4AB/W2MID[7] Tile_X9Y6_LUT4AB/W2END[0] Tile_X9Y6_LUT4AB/W2END[1]
+ Tile_X9Y6_LUT4AB/W2END[2] Tile_X9Y6_LUT4AB/W2END[3] Tile_X9Y6_LUT4AB/W2END[4] Tile_X9Y6_LUT4AB/W2END[5]
+ Tile_X9Y6_LUT4AB/W2END[6] Tile_X9Y6_LUT4AB/W2END[7] Tile_X9Y6_LUT4AB/W6END[0] Tile_X9Y6_LUT4AB/W6END[10]
+ Tile_X9Y6_LUT4AB/W6END[11] Tile_X9Y6_LUT4AB/W6END[1] Tile_X9Y6_LUT4AB/W6END[2] Tile_X9Y6_LUT4AB/W6END[3]
+ Tile_X9Y6_LUT4AB/W6END[4] Tile_X9Y6_LUT4AB/W6END[5] Tile_X9Y6_LUT4AB/W6END[6] Tile_X9Y6_LUT4AB/W6END[7]
+ Tile_X9Y6_LUT4AB/W6END[8] Tile_X9Y6_LUT4AB/W6END[9] Tile_X9Y6_LUT4AB/WW4END[0] Tile_X9Y6_LUT4AB/WW4END[10]
+ Tile_X9Y6_LUT4AB/WW4END[11] Tile_X9Y6_LUT4AB/WW4END[12] Tile_X9Y6_LUT4AB/WW4END[13]
+ Tile_X9Y6_LUT4AB/WW4END[14] Tile_X9Y6_LUT4AB/WW4END[15] Tile_X9Y6_LUT4AB/WW4END[1]
+ Tile_X9Y6_LUT4AB/WW4END[2] Tile_X9Y6_LUT4AB/WW4END[3] Tile_X9Y6_LUT4AB/WW4END[4]
+ Tile_X9Y6_LUT4AB/WW4END[5] Tile_X9Y6_LUT4AB/WW4END[6] Tile_X9Y6_LUT4AB/WW4END[7]
+ Tile_X9Y6_LUT4AB/WW4END[8] Tile_X9Y6_LUT4AB/WW4END[9] VGND VPWR Tile_X10Y6_WEN_SRAM
+ IHP_SRAM
XTile_X1Y14_LUT4AB Tile_X1Y14_LUT4AB/Ci Tile_X1Y14_LUT4AB/Co Tile_X2Y14_LUT4AB/E1END[0]
+ Tile_X2Y14_LUT4AB/E1END[1] Tile_X2Y14_LUT4AB/E1END[2] Tile_X2Y14_LUT4AB/E1END[3]
+ Tile_X0Y14_W_IO/E1BEG[0] Tile_X0Y14_W_IO/E1BEG[1] Tile_X0Y14_W_IO/E1BEG[2] Tile_X0Y14_W_IO/E1BEG[3]
+ Tile_X2Y14_LUT4AB/E2MID[0] Tile_X2Y14_LUT4AB/E2MID[1] Tile_X2Y14_LUT4AB/E2MID[2]
+ Tile_X2Y14_LUT4AB/E2MID[3] Tile_X2Y14_LUT4AB/E2MID[4] Tile_X2Y14_LUT4AB/E2MID[5]
+ Tile_X2Y14_LUT4AB/E2MID[6] Tile_X2Y14_LUT4AB/E2MID[7] Tile_X2Y14_LUT4AB/E2END[0]
+ Tile_X2Y14_LUT4AB/E2END[1] Tile_X2Y14_LUT4AB/E2END[2] Tile_X2Y14_LUT4AB/E2END[3]
+ Tile_X2Y14_LUT4AB/E2END[4] Tile_X2Y14_LUT4AB/E2END[5] Tile_X2Y14_LUT4AB/E2END[6]
+ Tile_X2Y14_LUT4AB/E2END[7] Tile_X0Y14_W_IO/E2BEGb[0] Tile_X0Y14_W_IO/E2BEGb[1] Tile_X0Y14_W_IO/E2BEGb[2]
+ Tile_X0Y14_W_IO/E2BEGb[3] Tile_X0Y14_W_IO/E2BEGb[4] Tile_X0Y14_W_IO/E2BEGb[5] Tile_X0Y14_W_IO/E2BEGb[6]
+ Tile_X0Y14_W_IO/E2BEGb[7] Tile_X0Y14_W_IO/E2BEG[0] Tile_X0Y14_W_IO/E2BEG[1] Tile_X0Y14_W_IO/E2BEG[2]
+ Tile_X0Y14_W_IO/E2BEG[3] Tile_X0Y14_W_IO/E2BEG[4] Tile_X0Y14_W_IO/E2BEG[5] Tile_X0Y14_W_IO/E2BEG[6]
+ Tile_X0Y14_W_IO/E2BEG[7] Tile_X2Y14_LUT4AB/E6END[0] Tile_X2Y14_LUT4AB/E6END[10]
+ Tile_X2Y14_LUT4AB/E6END[11] Tile_X2Y14_LUT4AB/E6END[1] Tile_X2Y14_LUT4AB/E6END[2]
+ Tile_X2Y14_LUT4AB/E6END[3] Tile_X2Y14_LUT4AB/E6END[4] Tile_X2Y14_LUT4AB/E6END[5]
+ Tile_X2Y14_LUT4AB/E6END[6] Tile_X2Y14_LUT4AB/E6END[7] Tile_X2Y14_LUT4AB/E6END[8]
+ Tile_X2Y14_LUT4AB/E6END[9] Tile_X0Y14_W_IO/E6BEG[0] Tile_X0Y14_W_IO/E6BEG[10] Tile_X0Y14_W_IO/E6BEG[11]
+ Tile_X0Y14_W_IO/E6BEG[1] Tile_X0Y14_W_IO/E6BEG[2] Tile_X0Y14_W_IO/E6BEG[3] Tile_X0Y14_W_IO/E6BEG[4]
+ Tile_X0Y14_W_IO/E6BEG[5] Tile_X0Y14_W_IO/E6BEG[6] Tile_X0Y14_W_IO/E6BEG[7] Tile_X0Y14_W_IO/E6BEG[8]
+ Tile_X0Y14_W_IO/E6BEG[9] Tile_X2Y14_LUT4AB/EE4END[0] Tile_X2Y14_LUT4AB/EE4END[10]
+ Tile_X2Y14_LUT4AB/EE4END[11] Tile_X2Y14_LUT4AB/EE4END[12] Tile_X2Y14_LUT4AB/EE4END[13]
+ Tile_X2Y14_LUT4AB/EE4END[14] Tile_X2Y14_LUT4AB/EE4END[15] Tile_X2Y14_LUT4AB/EE4END[1]
+ Tile_X2Y14_LUT4AB/EE4END[2] Tile_X2Y14_LUT4AB/EE4END[3] Tile_X2Y14_LUT4AB/EE4END[4]
+ Tile_X2Y14_LUT4AB/EE4END[5] Tile_X2Y14_LUT4AB/EE4END[6] Tile_X2Y14_LUT4AB/EE4END[7]
+ Tile_X2Y14_LUT4AB/EE4END[8] Tile_X2Y14_LUT4AB/EE4END[9] Tile_X0Y14_W_IO/EE4BEG[0]
+ Tile_X0Y14_W_IO/EE4BEG[10] Tile_X0Y14_W_IO/EE4BEG[11] Tile_X0Y14_W_IO/EE4BEG[12]
+ Tile_X0Y14_W_IO/EE4BEG[13] Tile_X0Y14_W_IO/EE4BEG[14] Tile_X0Y14_W_IO/EE4BEG[15]
+ Tile_X0Y14_W_IO/EE4BEG[1] Tile_X0Y14_W_IO/EE4BEG[2] Tile_X0Y14_W_IO/EE4BEG[3] Tile_X0Y14_W_IO/EE4BEG[4]
+ Tile_X0Y14_W_IO/EE4BEG[5] Tile_X0Y14_W_IO/EE4BEG[6] Tile_X0Y14_W_IO/EE4BEG[7] Tile_X0Y14_W_IO/EE4BEG[8]
+ Tile_X0Y14_W_IO/EE4BEG[9] Tile_X1Y14_LUT4AB/FrameData[0] Tile_X1Y14_LUT4AB/FrameData[10]
+ Tile_X1Y14_LUT4AB/FrameData[11] Tile_X1Y14_LUT4AB/FrameData[12] Tile_X1Y14_LUT4AB/FrameData[13]
+ Tile_X1Y14_LUT4AB/FrameData[14] Tile_X1Y14_LUT4AB/FrameData[15] Tile_X1Y14_LUT4AB/FrameData[16]
+ Tile_X1Y14_LUT4AB/FrameData[17] Tile_X1Y14_LUT4AB/FrameData[18] Tile_X1Y14_LUT4AB/FrameData[19]
+ Tile_X1Y14_LUT4AB/FrameData[1] Tile_X1Y14_LUT4AB/FrameData[20] Tile_X1Y14_LUT4AB/FrameData[21]
+ Tile_X1Y14_LUT4AB/FrameData[22] Tile_X1Y14_LUT4AB/FrameData[23] Tile_X1Y14_LUT4AB/FrameData[24]
+ Tile_X1Y14_LUT4AB/FrameData[25] Tile_X1Y14_LUT4AB/FrameData[26] Tile_X1Y14_LUT4AB/FrameData[27]
+ Tile_X1Y14_LUT4AB/FrameData[28] Tile_X1Y14_LUT4AB/FrameData[29] Tile_X1Y14_LUT4AB/FrameData[2]
+ Tile_X1Y14_LUT4AB/FrameData[30] Tile_X1Y14_LUT4AB/FrameData[31] Tile_X1Y14_LUT4AB/FrameData[3]
+ Tile_X1Y14_LUT4AB/FrameData[4] Tile_X1Y14_LUT4AB/FrameData[5] Tile_X1Y14_LUT4AB/FrameData[6]
+ Tile_X1Y14_LUT4AB/FrameData[7] Tile_X1Y14_LUT4AB/FrameData[8] Tile_X1Y14_LUT4AB/FrameData[9]
+ Tile_X2Y14_LUT4AB/FrameData[0] Tile_X2Y14_LUT4AB/FrameData[10] Tile_X2Y14_LUT4AB/FrameData[11]
+ Tile_X2Y14_LUT4AB/FrameData[12] Tile_X2Y14_LUT4AB/FrameData[13] Tile_X2Y14_LUT4AB/FrameData[14]
+ Tile_X2Y14_LUT4AB/FrameData[15] Tile_X2Y14_LUT4AB/FrameData[16] Tile_X2Y14_LUT4AB/FrameData[17]
+ Tile_X2Y14_LUT4AB/FrameData[18] Tile_X2Y14_LUT4AB/FrameData[19] Tile_X2Y14_LUT4AB/FrameData[1]
+ Tile_X2Y14_LUT4AB/FrameData[20] Tile_X2Y14_LUT4AB/FrameData[21] Tile_X2Y14_LUT4AB/FrameData[22]
+ Tile_X2Y14_LUT4AB/FrameData[23] Tile_X2Y14_LUT4AB/FrameData[24] Tile_X2Y14_LUT4AB/FrameData[25]
+ Tile_X2Y14_LUT4AB/FrameData[26] Tile_X2Y14_LUT4AB/FrameData[27] Tile_X2Y14_LUT4AB/FrameData[28]
+ Tile_X2Y14_LUT4AB/FrameData[29] Tile_X2Y14_LUT4AB/FrameData[2] Tile_X2Y14_LUT4AB/FrameData[30]
+ Tile_X2Y14_LUT4AB/FrameData[31] Tile_X2Y14_LUT4AB/FrameData[3] Tile_X2Y14_LUT4AB/FrameData[4]
+ Tile_X2Y14_LUT4AB/FrameData[5] Tile_X2Y14_LUT4AB/FrameData[6] Tile_X2Y14_LUT4AB/FrameData[7]
+ Tile_X2Y14_LUT4AB/FrameData[8] Tile_X2Y14_LUT4AB/FrameData[9] Tile_X1Y14_LUT4AB/FrameStrobe[0]
+ Tile_X1Y14_LUT4AB/FrameStrobe[10] Tile_X1Y14_LUT4AB/FrameStrobe[11] Tile_X1Y14_LUT4AB/FrameStrobe[12]
+ Tile_X1Y14_LUT4AB/FrameStrobe[13] Tile_X1Y14_LUT4AB/FrameStrobe[14] Tile_X1Y14_LUT4AB/FrameStrobe[15]
+ Tile_X1Y14_LUT4AB/FrameStrobe[16] Tile_X1Y14_LUT4AB/FrameStrobe[17] Tile_X1Y14_LUT4AB/FrameStrobe[18]
+ Tile_X1Y14_LUT4AB/FrameStrobe[19] Tile_X1Y14_LUT4AB/FrameStrobe[1] Tile_X1Y14_LUT4AB/FrameStrobe[2]
+ Tile_X1Y14_LUT4AB/FrameStrobe[3] Tile_X1Y14_LUT4AB/FrameStrobe[4] Tile_X1Y14_LUT4AB/FrameStrobe[5]
+ Tile_X1Y14_LUT4AB/FrameStrobe[6] Tile_X1Y14_LUT4AB/FrameStrobe[7] Tile_X1Y14_LUT4AB/FrameStrobe[8]
+ Tile_X1Y14_LUT4AB/FrameStrobe[9] Tile_X1Y13_LUT4AB/FrameStrobe[0] Tile_X1Y13_LUT4AB/FrameStrobe[10]
+ Tile_X1Y13_LUT4AB/FrameStrobe[11] Tile_X1Y13_LUT4AB/FrameStrobe[12] Tile_X1Y13_LUT4AB/FrameStrobe[13]
+ Tile_X1Y13_LUT4AB/FrameStrobe[14] Tile_X1Y13_LUT4AB/FrameStrobe[15] Tile_X1Y13_LUT4AB/FrameStrobe[16]
+ Tile_X1Y13_LUT4AB/FrameStrobe[17] Tile_X1Y13_LUT4AB/FrameStrobe[18] Tile_X1Y13_LUT4AB/FrameStrobe[19]
+ Tile_X1Y13_LUT4AB/FrameStrobe[1] Tile_X1Y13_LUT4AB/FrameStrobe[2] Tile_X1Y13_LUT4AB/FrameStrobe[3]
+ Tile_X1Y13_LUT4AB/FrameStrobe[4] Tile_X1Y13_LUT4AB/FrameStrobe[5] Tile_X1Y13_LUT4AB/FrameStrobe[6]
+ Tile_X1Y13_LUT4AB/FrameStrobe[7] Tile_X1Y13_LUT4AB/FrameStrobe[8] Tile_X1Y13_LUT4AB/FrameStrobe[9]
+ Tile_X1Y14_LUT4AB/N1BEG[0] Tile_X1Y14_LUT4AB/N1BEG[1] Tile_X1Y14_LUT4AB/N1BEG[2]
+ Tile_X1Y14_LUT4AB/N1BEG[3] Tile_X1Y14_LUT4AB/N1END[0] Tile_X1Y14_LUT4AB/N1END[1]
+ Tile_X1Y14_LUT4AB/N1END[2] Tile_X1Y14_LUT4AB/N1END[3] Tile_X1Y14_LUT4AB/N2BEG[0]
+ Tile_X1Y14_LUT4AB/N2BEG[1] Tile_X1Y14_LUT4AB/N2BEG[2] Tile_X1Y14_LUT4AB/N2BEG[3]
+ Tile_X1Y14_LUT4AB/N2BEG[4] Tile_X1Y14_LUT4AB/N2BEG[5] Tile_X1Y14_LUT4AB/N2BEG[6]
+ Tile_X1Y14_LUT4AB/N2BEG[7] Tile_X1Y13_LUT4AB/N2END[0] Tile_X1Y13_LUT4AB/N2END[1]
+ Tile_X1Y13_LUT4AB/N2END[2] Tile_X1Y13_LUT4AB/N2END[3] Tile_X1Y13_LUT4AB/N2END[4]
+ Tile_X1Y13_LUT4AB/N2END[5] Tile_X1Y13_LUT4AB/N2END[6] Tile_X1Y13_LUT4AB/N2END[7]
+ Tile_X1Y14_LUT4AB/N2END[0] Tile_X1Y14_LUT4AB/N2END[1] Tile_X1Y14_LUT4AB/N2END[2]
+ Tile_X1Y14_LUT4AB/N2END[3] Tile_X1Y14_LUT4AB/N2END[4] Tile_X1Y14_LUT4AB/N2END[5]
+ Tile_X1Y14_LUT4AB/N2END[6] Tile_X1Y14_LUT4AB/N2END[7] Tile_X1Y14_LUT4AB/N2MID[0]
+ Tile_X1Y14_LUT4AB/N2MID[1] Tile_X1Y14_LUT4AB/N2MID[2] Tile_X1Y14_LUT4AB/N2MID[3]
+ Tile_X1Y14_LUT4AB/N2MID[4] Tile_X1Y14_LUT4AB/N2MID[5] Tile_X1Y14_LUT4AB/N2MID[6]
+ Tile_X1Y14_LUT4AB/N2MID[7] Tile_X1Y14_LUT4AB/N4BEG[0] Tile_X1Y14_LUT4AB/N4BEG[10]
+ Tile_X1Y14_LUT4AB/N4BEG[11] Tile_X1Y14_LUT4AB/N4BEG[12] Tile_X1Y14_LUT4AB/N4BEG[13]
+ Tile_X1Y14_LUT4AB/N4BEG[14] Tile_X1Y14_LUT4AB/N4BEG[15] Tile_X1Y14_LUT4AB/N4BEG[1]
+ Tile_X1Y14_LUT4AB/N4BEG[2] Tile_X1Y14_LUT4AB/N4BEG[3] Tile_X1Y14_LUT4AB/N4BEG[4]
+ Tile_X1Y14_LUT4AB/N4BEG[5] Tile_X1Y14_LUT4AB/N4BEG[6] Tile_X1Y14_LUT4AB/N4BEG[7]
+ Tile_X1Y14_LUT4AB/N4BEG[8] Tile_X1Y14_LUT4AB/N4BEG[9] Tile_X1Y14_LUT4AB/N4END[0]
+ Tile_X1Y14_LUT4AB/N4END[10] Tile_X1Y14_LUT4AB/N4END[11] Tile_X1Y14_LUT4AB/N4END[12]
+ Tile_X1Y14_LUT4AB/N4END[13] Tile_X1Y14_LUT4AB/N4END[14] Tile_X1Y14_LUT4AB/N4END[15]
+ Tile_X1Y14_LUT4AB/N4END[1] Tile_X1Y14_LUT4AB/N4END[2] Tile_X1Y14_LUT4AB/N4END[3]
+ Tile_X1Y14_LUT4AB/N4END[4] Tile_X1Y14_LUT4AB/N4END[5] Tile_X1Y14_LUT4AB/N4END[6]
+ Tile_X1Y14_LUT4AB/N4END[7] Tile_X1Y14_LUT4AB/N4END[8] Tile_X1Y14_LUT4AB/N4END[9]
+ Tile_X1Y14_LUT4AB/NN4BEG[0] Tile_X1Y14_LUT4AB/NN4BEG[10] Tile_X1Y14_LUT4AB/NN4BEG[11]
+ Tile_X1Y14_LUT4AB/NN4BEG[12] Tile_X1Y14_LUT4AB/NN4BEG[13] Tile_X1Y14_LUT4AB/NN4BEG[14]
+ Tile_X1Y14_LUT4AB/NN4BEG[15] Tile_X1Y14_LUT4AB/NN4BEG[1] Tile_X1Y14_LUT4AB/NN4BEG[2]
+ Tile_X1Y14_LUT4AB/NN4BEG[3] Tile_X1Y14_LUT4AB/NN4BEG[4] Tile_X1Y14_LUT4AB/NN4BEG[5]
+ Tile_X1Y14_LUT4AB/NN4BEG[6] Tile_X1Y14_LUT4AB/NN4BEG[7] Tile_X1Y14_LUT4AB/NN4BEG[8]
+ Tile_X1Y14_LUT4AB/NN4BEG[9] Tile_X1Y14_LUT4AB/NN4END[0] Tile_X1Y14_LUT4AB/NN4END[10]
+ Tile_X1Y14_LUT4AB/NN4END[11] Tile_X1Y14_LUT4AB/NN4END[12] Tile_X1Y14_LUT4AB/NN4END[13]
+ Tile_X1Y14_LUT4AB/NN4END[14] Tile_X1Y14_LUT4AB/NN4END[15] Tile_X1Y14_LUT4AB/NN4END[1]
+ Tile_X1Y14_LUT4AB/NN4END[2] Tile_X1Y14_LUT4AB/NN4END[3] Tile_X1Y14_LUT4AB/NN4END[4]
+ Tile_X1Y14_LUT4AB/NN4END[5] Tile_X1Y14_LUT4AB/NN4END[6] Tile_X1Y14_LUT4AB/NN4END[7]
+ Tile_X1Y14_LUT4AB/NN4END[8] Tile_X1Y14_LUT4AB/NN4END[9] Tile_X1Y14_LUT4AB/S1BEG[0]
+ Tile_X1Y14_LUT4AB/S1BEG[1] Tile_X1Y14_LUT4AB/S1BEG[2] Tile_X1Y14_LUT4AB/S1BEG[3]
+ Tile_X1Y14_LUT4AB/S1END[0] Tile_X1Y14_LUT4AB/S1END[1] Tile_X1Y14_LUT4AB/S1END[2]
+ Tile_X1Y14_LUT4AB/S1END[3] Tile_X1Y14_LUT4AB/S2BEG[0] Tile_X1Y14_LUT4AB/S2BEG[1]
+ Tile_X1Y14_LUT4AB/S2BEG[2] Tile_X1Y14_LUT4AB/S2BEG[3] Tile_X1Y14_LUT4AB/S2BEG[4]
+ Tile_X1Y14_LUT4AB/S2BEG[5] Tile_X1Y14_LUT4AB/S2BEG[6] Tile_X1Y14_LUT4AB/S2BEG[7]
+ Tile_X1Y14_LUT4AB/S2BEGb[0] Tile_X1Y14_LUT4AB/S2BEGb[1] Tile_X1Y14_LUT4AB/S2BEGb[2]
+ Tile_X1Y14_LUT4AB/S2BEGb[3] Tile_X1Y14_LUT4AB/S2BEGb[4] Tile_X1Y14_LUT4AB/S2BEGb[5]
+ Tile_X1Y14_LUT4AB/S2BEGb[6] Tile_X1Y14_LUT4AB/S2BEGb[7] Tile_X1Y14_LUT4AB/S2END[0]
+ Tile_X1Y14_LUT4AB/S2END[1] Tile_X1Y14_LUT4AB/S2END[2] Tile_X1Y14_LUT4AB/S2END[3]
+ Tile_X1Y14_LUT4AB/S2END[4] Tile_X1Y14_LUT4AB/S2END[5] Tile_X1Y14_LUT4AB/S2END[6]
+ Tile_X1Y14_LUT4AB/S2END[7] Tile_X1Y14_LUT4AB/S2MID[0] Tile_X1Y14_LUT4AB/S2MID[1]
+ Tile_X1Y14_LUT4AB/S2MID[2] Tile_X1Y14_LUT4AB/S2MID[3] Tile_X1Y14_LUT4AB/S2MID[4]
+ Tile_X1Y14_LUT4AB/S2MID[5] Tile_X1Y14_LUT4AB/S2MID[6] Tile_X1Y14_LUT4AB/S2MID[7]
+ Tile_X1Y14_LUT4AB/S4BEG[0] Tile_X1Y14_LUT4AB/S4BEG[10] Tile_X1Y14_LUT4AB/S4BEG[11]
+ Tile_X1Y14_LUT4AB/S4BEG[12] Tile_X1Y14_LUT4AB/S4BEG[13] Tile_X1Y14_LUT4AB/S4BEG[14]
+ Tile_X1Y14_LUT4AB/S4BEG[15] Tile_X1Y14_LUT4AB/S4BEG[1] Tile_X1Y14_LUT4AB/S4BEG[2]
+ Tile_X1Y14_LUT4AB/S4BEG[3] Tile_X1Y14_LUT4AB/S4BEG[4] Tile_X1Y14_LUT4AB/S4BEG[5]
+ Tile_X1Y14_LUT4AB/S4BEG[6] Tile_X1Y14_LUT4AB/S4BEG[7] Tile_X1Y14_LUT4AB/S4BEG[8]
+ Tile_X1Y14_LUT4AB/S4BEG[9] Tile_X1Y14_LUT4AB/S4END[0] Tile_X1Y14_LUT4AB/S4END[10]
+ Tile_X1Y14_LUT4AB/S4END[11] Tile_X1Y14_LUT4AB/S4END[12] Tile_X1Y14_LUT4AB/S4END[13]
+ Tile_X1Y14_LUT4AB/S4END[14] Tile_X1Y14_LUT4AB/S4END[15] Tile_X1Y14_LUT4AB/S4END[1]
+ Tile_X1Y14_LUT4AB/S4END[2] Tile_X1Y14_LUT4AB/S4END[3] Tile_X1Y14_LUT4AB/S4END[4]
+ Tile_X1Y14_LUT4AB/S4END[5] Tile_X1Y14_LUT4AB/S4END[6] Tile_X1Y14_LUT4AB/S4END[7]
+ Tile_X1Y14_LUT4AB/S4END[8] Tile_X1Y14_LUT4AB/S4END[9] Tile_X1Y14_LUT4AB/SS4BEG[0]
+ Tile_X1Y14_LUT4AB/SS4BEG[10] Tile_X1Y14_LUT4AB/SS4BEG[11] Tile_X1Y14_LUT4AB/SS4BEG[12]
+ Tile_X1Y14_LUT4AB/SS4BEG[13] Tile_X1Y14_LUT4AB/SS4BEG[14] Tile_X1Y14_LUT4AB/SS4BEG[15]
+ Tile_X1Y14_LUT4AB/SS4BEG[1] Tile_X1Y14_LUT4AB/SS4BEG[2] Tile_X1Y14_LUT4AB/SS4BEG[3]
+ Tile_X1Y14_LUT4AB/SS4BEG[4] Tile_X1Y14_LUT4AB/SS4BEG[5] Tile_X1Y14_LUT4AB/SS4BEG[6]
+ Tile_X1Y14_LUT4AB/SS4BEG[7] Tile_X1Y14_LUT4AB/SS4BEG[8] Tile_X1Y14_LUT4AB/SS4BEG[9]
+ Tile_X1Y14_LUT4AB/SS4END[0] Tile_X1Y14_LUT4AB/SS4END[10] Tile_X1Y14_LUT4AB/SS4END[11]
+ Tile_X1Y14_LUT4AB/SS4END[12] Tile_X1Y14_LUT4AB/SS4END[13] Tile_X1Y14_LUT4AB/SS4END[14]
+ Tile_X1Y14_LUT4AB/SS4END[15] Tile_X1Y14_LUT4AB/SS4END[1] Tile_X1Y14_LUT4AB/SS4END[2]
+ Tile_X1Y14_LUT4AB/SS4END[3] Tile_X1Y14_LUT4AB/SS4END[4] Tile_X1Y14_LUT4AB/SS4END[5]
+ Tile_X1Y14_LUT4AB/SS4END[6] Tile_X1Y14_LUT4AB/SS4END[7] Tile_X1Y14_LUT4AB/SS4END[8]
+ Tile_X1Y14_LUT4AB/SS4END[9] Tile_X1Y14_LUT4AB/UserCLK Tile_X1Y13_LUT4AB/UserCLK
+ VGND VPWR Tile_X0Y14_W_IO/W1END[0] Tile_X0Y14_W_IO/W1END[1] Tile_X0Y14_W_IO/W1END[2]
+ Tile_X0Y14_W_IO/W1END[3] Tile_X2Y14_LUT4AB/W1BEG[0] Tile_X2Y14_LUT4AB/W1BEG[1] Tile_X2Y14_LUT4AB/W1BEG[2]
+ Tile_X2Y14_LUT4AB/W1BEG[3] Tile_X0Y14_W_IO/W2MID[0] Tile_X0Y14_W_IO/W2MID[1] Tile_X0Y14_W_IO/W2MID[2]
+ Tile_X0Y14_W_IO/W2MID[3] Tile_X0Y14_W_IO/W2MID[4] Tile_X0Y14_W_IO/W2MID[5] Tile_X0Y14_W_IO/W2MID[6]
+ Tile_X0Y14_W_IO/W2MID[7] Tile_X0Y14_W_IO/W2END[0] Tile_X0Y14_W_IO/W2END[1] Tile_X0Y14_W_IO/W2END[2]
+ Tile_X0Y14_W_IO/W2END[3] Tile_X0Y14_W_IO/W2END[4] Tile_X0Y14_W_IO/W2END[5] Tile_X0Y14_W_IO/W2END[6]
+ Tile_X0Y14_W_IO/W2END[7] Tile_X1Y14_LUT4AB/W2END[0] Tile_X1Y14_LUT4AB/W2END[1] Tile_X1Y14_LUT4AB/W2END[2]
+ Tile_X1Y14_LUT4AB/W2END[3] Tile_X1Y14_LUT4AB/W2END[4] Tile_X1Y14_LUT4AB/W2END[5]
+ Tile_X1Y14_LUT4AB/W2END[6] Tile_X1Y14_LUT4AB/W2END[7] Tile_X2Y14_LUT4AB/W2BEG[0]
+ Tile_X2Y14_LUT4AB/W2BEG[1] Tile_X2Y14_LUT4AB/W2BEG[2] Tile_X2Y14_LUT4AB/W2BEG[3]
+ Tile_X2Y14_LUT4AB/W2BEG[4] Tile_X2Y14_LUT4AB/W2BEG[5] Tile_X2Y14_LUT4AB/W2BEG[6]
+ Tile_X2Y14_LUT4AB/W2BEG[7] Tile_X0Y14_W_IO/W6END[0] Tile_X0Y14_W_IO/W6END[10] Tile_X0Y14_W_IO/W6END[11]
+ Tile_X0Y14_W_IO/W6END[1] Tile_X0Y14_W_IO/W6END[2] Tile_X0Y14_W_IO/W6END[3] Tile_X0Y14_W_IO/W6END[4]
+ Tile_X0Y14_W_IO/W6END[5] Tile_X0Y14_W_IO/W6END[6] Tile_X0Y14_W_IO/W6END[7] Tile_X0Y14_W_IO/W6END[8]
+ Tile_X0Y14_W_IO/W6END[9] Tile_X2Y14_LUT4AB/W6BEG[0] Tile_X2Y14_LUT4AB/W6BEG[10]
+ Tile_X2Y14_LUT4AB/W6BEG[11] Tile_X2Y14_LUT4AB/W6BEG[1] Tile_X2Y14_LUT4AB/W6BEG[2]
+ Tile_X2Y14_LUT4AB/W6BEG[3] Tile_X2Y14_LUT4AB/W6BEG[4] Tile_X2Y14_LUT4AB/W6BEG[5]
+ Tile_X2Y14_LUT4AB/W6BEG[6] Tile_X2Y14_LUT4AB/W6BEG[7] Tile_X2Y14_LUT4AB/W6BEG[8]
+ Tile_X2Y14_LUT4AB/W6BEG[9] Tile_X0Y14_W_IO/WW4END[0] Tile_X0Y14_W_IO/WW4END[10]
+ Tile_X0Y14_W_IO/WW4END[11] Tile_X0Y14_W_IO/WW4END[12] Tile_X0Y14_W_IO/WW4END[13]
+ Tile_X0Y14_W_IO/WW4END[14] Tile_X0Y14_W_IO/WW4END[15] Tile_X0Y14_W_IO/WW4END[1]
+ Tile_X0Y14_W_IO/WW4END[2] Tile_X0Y14_W_IO/WW4END[3] Tile_X0Y14_W_IO/WW4END[4] Tile_X0Y14_W_IO/WW4END[5]
+ Tile_X0Y14_W_IO/WW4END[6] Tile_X0Y14_W_IO/WW4END[7] Tile_X0Y14_W_IO/WW4END[8] Tile_X0Y14_W_IO/WW4END[9]
+ Tile_X2Y14_LUT4AB/WW4BEG[0] Tile_X2Y14_LUT4AB/WW4BEG[10] Tile_X2Y14_LUT4AB/WW4BEG[11]
+ Tile_X2Y14_LUT4AB/WW4BEG[12] Tile_X2Y14_LUT4AB/WW4BEG[13] Tile_X2Y14_LUT4AB/WW4BEG[14]
+ Tile_X2Y14_LUT4AB/WW4BEG[15] Tile_X2Y14_LUT4AB/WW4BEG[1] Tile_X2Y14_LUT4AB/WW4BEG[2]
+ Tile_X2Y14_LUT4AB/WW4BEG[3] Tile_X2Y14_LUT4AB/WW4BEG[4] Tile_X2Y14_LUT4AB/WW4BEG[5]
+ Tile_X2Y14_LUT4AB/WW4BEG[6] Tile_X2Y14_LUT4AB/WW4BEG[7] Tile_X2Y14_LUT4AB/WW4BEG[8]
+ Tile_X2Y14_LUT4AB/WW4BEG[9] LUT4AB
XTile_X6Y9_LUT4AB Tile_X6Y9_LUT4AB/Ci Tile_X6Y9_LUT4AB/Co Tile_X6Y9_LUT4AB/E1BEG[0]
+ Tile_X6Y9_LUT4AB/E1BEG[1] Tile_X6Y9_LUT4AB/E1BEG[2] Tile_X6Y9_LUT4AB/E1BEG[3] Tile_X6Y9_LUT4AB/E1END[0]
+ Tile_X6Y9_LUT4AB/E1END[1] Tile_X6Y9_LUT4AB/E1END[2] Tile_X6Y9_LUT4AB/E1END[3] Tile_X6Y9_LUT4AB/E2BEG[0]
+ Tile_X6Y9_LUT4AB/E2BEG[1] Tile_X6Y9_LUT4AB/E2BEG[2] Tile_X6Y9_LUT4AB/E2BEG[3] Tile_X6Y9_LUT4AB/E2BEG[4]
+ Tile_X6Y9_LUT4AB/E2BEG[5] Tile_X6Y9_LUT4AB/E2BEG[6] Tile_X6Y9_LUT4AB/E2BEG[7] Tile_X6Y9_LUT4AB/E2BEGb[0]
+ Tile_X6Y9_LUT4AB/E2BEGb[1] Tile_X6Y9_LUT4AB/E2BEGb[2] Tile_X6Y9_LUT4AB/E2BEGb[3]
+ Tile_X6Y9_LUT4AB/E2BEGb[4] Tile_X6Y9_LUT4AB/E2BEGb[5] Tile_X6Y9_LUT4AB/E2BEGb[6]
+ Tile_X6Y9_LUT4AB/E2BEGb[7] Tile_X6Y9_LUT4AB/E2END[0] Tile_X6Y9_LUT4AB/E2END[1] Tile_X6Y9_LUT4AB/E2END[2]
+ Tile_X6Y9_LUT4AB/E2END[3] Tile_X6Y9_LUT4AB/E2END[4] Tile_X6Y9_LUT4AB/E2END[5] Tile_X6Y9_LUT4AB/E2END[6]
+ Tile_X6Y9_LUT4AB/E2END[7] Tile_X6Y9_LUT4AB/E2MID[0] Tile_X6Y9_LUT4AB/E2MID[1] Tile_X6Y9_LUT4AB/E2MID[2]
+ Tile_X6Y9_LUT4AB/E2MID[3] Tile_X6Y9_LUT4AB/E2MID[4] Tile_X6Y9_LUT4AB/E2MID[5] Tile_X6Y9_LUT4AB/E2MID[6]
+ Tile_X6Y9_LUT4AB/E2MID[7] Tile_X6Y9_LUT4AB/E6BEG[0] Tile_X6Y9_LUT4AB/E6BEG[10] Tile_X6Y9_LUT4AB/E6BEG[11]
+ Tile_X6Y9_LUT4AB/E6BEG[1] Tile_X6Y9_LUT4AB/E6BEG[2] Tile_X6Y9_LUT4AB/E6BEG[3] Tile_X6Y9_LUT4AB/E6BEG[4]
+ Tile_X6Y9_LUT4AB/E6BEG[5] Tile_X6Y9_LUT4AB/E6BEG[6] Tile_X6Y9_LUT4AB/E6BEG[7] Tile_X6Y9_LUT4AB/E6BEG[8]
+ Tile_X6Y9_LUT4AB/E6BEG[9] Tile_X6Y9_LUT4AB/E6END[0] Tile_X6Y9_LUT4AB/E6END[10] Tile_X6Y9_LUT4AB/E6END[11]
+ Tile_X6Y9_LUT4AB/E6END[1] Tile_X6Y9_LUT4AB/E6END[2] Tile_X6Y9_LUT4AB/E6END[3] Tile_X6Y9_LUT4AB/E6END[4]
+ Tile_X6Y9_LUT4AB/E6END[5] Tile_X6Y9_LUT4AB/E6END[6] Tile_X6Y9_LUT4AB/E6END[7] Tile_X6Y9_LUT4AB/E6END[8]
+ Tile_X6Y9_LUT4AB/E6END[9] Tile_X6Y9_LUT4AB/EE4BEG[0] Tile_X6Y9_LUT4AB/EE4BEG[10]
+ Tile_X6Y9_LUT4AB/EE4BEG[11] Tile_X6Y9_LUT4AB/EE4BEG[12] Tile_X6Y9_LUT4AB/EE4BEG[13]
+ Tile_X6Y9_LUT4AB/EE4BEG[14] Tile_X6Y9_LUT4AB/EE4BEG[15] Tile_X6Y9_LUT4AB/EE4BEG[1]
+ Tile_X6Y9_LUT4AB/EE4BEG[2] Tile_X6Y9_LUT4AB/EE4BEG[3] Tile_X6Y9_LUT4AB/EE4BEG[4]
+ Tile_X6Y9_LUT4AB/EE4BEG[5] Tile_X6Y9_LUT4AB/EE4BEG[6] Tile_X6Y9_LUT4AB/EE4BEG[7]
+ Tile_X6Y9_LUT4AB/EE4BEG[8] Tile_X6Y9_LUT4AB/EE4BEG[9] Tile_X6Y9_LUT4AB/EE4END[0]
+ Tile_X6Y9_LUT4AB/EE4END[10] Tile_X6Y9_LUT4AB/EE4END[11] Tile_X6Y9_LUT4AB/EE4END[12]
+ Tile_X6Y9_LUT4AB/EE4END[13] Tile_X6Y9_LUT4AB/EE4END[14] Tile_X6Y9_LUT4AB/EE4END[15]
+ Tile_X6Y9_LUT4AB/EE4END[1] Tile_X6Y9_LUT4AB/EE4END[2] Tile_X6Y9_LUT4AB/EE4END[3]
+ Tile_X6Y9_LUT4AB/EE4END[4] Tile_X6Y9_LUT4AB/EE4END[5] Tile_X6Y9_LUT4AB/EE4END[6]
+ Tile_X6Y9_LUT4AB/EE4END[7] Tile_X6Y9_LUT4AB/EE4END[8] Tile_X6Y9_LUT4AB/EE4END[9]
+ Tile_X6Y9_LUT4AB/FrameData[0] Tile_X6Y9_LUT4AB/FrameData[10] Tile_X6Y9_LUT4AB/FrameData[11]
+ Tile_X6Y9_LUT4AB/FrameData[12] Tile_X6Y9_LUT4AB/FrameData[13] Tile_X6Y9_LUT4AB/FrameData[14]
+ Tile_X6Y9_LUT4AB/FrameData[15] Tile_X6Y9_LUT4AB/FrameData[16] Tile_X6Y9_LUT4AB/FrameData[17]
+ Tile_X6Y9_LUT4AB/FrameData[18] Tile_X6Y9_LUT4AB/FrameData[19] Tile_X6Y9_LUT4AB/FrameData[1]
+ Tile_X6Y9_LUT4AB/FrameData[20] Tile_X6Y9_LUT4AB/FrameData[21] Tile_X6Y9_LUT4AB/FrameData[22]
+ Tile_X6Y9_LUT4AB/FrameData[23] Tile_X6Y9_LUT4AB/FrameData[24] Tile_X6Y9_LUT4AB/FrameData[25]
+ Tile_X6Y9_LUT4AB/FrameData[26] Tile_X6Y9_LUT4AB/FrameData[27] Tile_X6Y9_LUT4AB/FrameData[28]
+ Tile_X6Y9_LUT4AB/FrameData[29] Tile_X6Y9_LUT4AB/FrameData[2] Tile_X6Y9_LUT4AB/FrameData[30]
+ Tile_X6Y9_LUT4AB/FrameData[31] Tile_X6Y9_LUT4AB/FrameData[3] Tile_X6Y9_LUT4AB/FrameData[4]
+ Tile_X6Y9_LUT4AB/FrameData[5] Tile_X6Y9_LUT4AB/FrameData[6] Tile_X6Y9_LUT4AB/FrameData[7]
+ Tile_X6Y9_LUT4AB/FrameData[8] Tile_X6Y9_LUT4AB/FrameData[9] Tile_X6Y9_LUT4AB/FrameData_O[0]
+ Tile_X6Y9_LUT4AB/FrameData_O[10] Tile_X6Y9_LUT4AB/FrameData_O[11] Tile_X6Y9_LUT4AB/FrameData_O[12]
+ Tile_X6Y9_LUT4AB/FrameData_O[13] Tile_X6Y9_LUT4AB/FrameData_O[14] Tile_X6Y9_LUT4AB/FrameData_O[15]
+ Tile_X6Y9_LUT4AB/FrameData_O[16] Tile_X6Y9_LUT4AB/FrameData_O[17] Tile_X6Y9_LUT4AB/FrameData_O[18]
+ Tile_X6Y9_LUT4AB/FrameData_O[19] Tile_X6Y9_LUT4AB/FrameData_O[1] Tile_X6Y9_LUT4AB/FrameData_O[20]
+ Tile_X6Y9_LUT4AB/FrameData_O[21] Tile_X6Y9_LUT4AB/FrameData_O[22] Tile_X6Y9_LUT4AB/FrameData_O[23]
+ Tile_X6Y9_LUT4AB/FrameData_O[24] Tile_X6Y9_LUT4AB/FrameData_O[25] Tile_X6Y9_LUT4AB/FrameData_O[26]
+ Tile_X6Y9_LUT4AB/FrameData_O[27] Tile_X6Y9_LUT4AB/FrameData_O[28] Tile_X6Y9_LUT4AB/FrameData_O[29]
+ Tile_X6Y9_LUT4AB/FrameData_O[2] Tile_X6Y9_LUT4AB/FrameData_O[30] Tile_X6Y9_LUT4AB/FrameData_O[31]
+ Tile_X6Y9_LUT4AB/FrameData_O[3] Tile_X6Y9_LUT4AB/FrameData_O[4] Tile_X6Y9_LUT4AB/FrameData_O[5]
+ Tile_X6Y9_LUT4AB/FrameData_O[6] Tile_X6Y9_LUT4AB/FrameData_O[7] Tile_X6Y9_LUT4AB/FrameData_O[8]
+ Tile_X6Y9_LUT4AB/FrameData_O[9] Tile_X6Y9_LUT4AB/FrameStrobe[0] Tile_X6Y9_LUT4AB/FrameStrobe[10]
+ Tile_X6Y9_LUT4AB/FrameStrobe[11] Tile_X6Y9_LUT4AB/FrameStrobe[12] Tile_X6Y9_LUT4AB/FrameStrobe[13]
+ Tile_X6Y9_LUT4AB/FrameStrobe[14] Tile_X6Y9_LUT4AB/FrameStrobe[15] Tile_X6Y9_LUT4AB/FrameStrobe[16]
+ Tile_X6Y9_LUT4AB/FrameStrobe[17] Tile_X6Y9_LUT4AB/FrameStrobe[18] Tile_X6Y9_LUT4AB/FrameStrobe[19]
+ Tile_X6Y9_LUT4AB/FrameStrobe[1] Tile_X6Y9_LUT4AB/FrameStrobe[2] Tile_X6Y9_LUT4AB/FrameStrobe[3]
+ Tile_X6Y9_LUT4AB/FrameStrobe[4] Tile_X6Y9_LUT4AB/FrameStrobe[5] Tile_X6Y9_LUT4AB/FrameStrobe[6]
+ Tile_X6Y9_LUT4AB/FrameStrobe[7] Tile_X6Y9_LUT4AB/FrameStrobe[8] Tile_X6Y9_LUT4AB/FrameStrobe[9]
+ Tile_X6Y8_LUT4AB/FrameStrobe[0] Tile_X6Y8_LUT4AB/FrameStrobe[10] Tile_X6Y8_LUT4AB/FrameStrobe[11]
+ Tile_X6Y8_LUT4AB/FrameStrobe[12] Tile_X6Y8_LUT4AB/FrameStrobe[13] Tile_X6Y8_LUT4AB/FrameStrobe[14]
+ Tile_X6Y8_LUT4AB/FrameStrobe[15] Tile_X6Y8_LUT4AB/FrameStrobe[16] Tile_X6Y8_LUT4AB/FrameStrobe[17]
+ Tile_X6Y8_LUT4AB/FrameStrobe[18] Tile_X6Y8_LUT4AB/FrameStrobe[19] Tile_X6Y8_LUT4AB/FrameStrobe[1]
+ Tile_X6Y8_LUT4AB/FrameStrobe[2] Tile_X6Y8_LUT4AB/FrameStrobe[3] Tile_X6Y8_LUT4AB/FrameStrobe[4]
+ Tile_X6Y8_LUT4AB/FrameStrobe[5] Tile_X6Y8_LUT4AB/FrameStrobe[6] Tile_X6Y8_LUT4AB/FrameStrobe[7]
+ Tile_X6Y8_LUT4AB/FrameStrobe[8] Tile_X6Y8_LUT4AB/FrameStrobe[9] Tile_X6Y9_LUT4AB/N1BEG[0]
+ Tile_X6Y9_LUT4AB/N1BEG[1] Tile_X6Y9_LUT4AB/N1BEG[2] Tile_X6Y9_LUT4AB/N1BEG[3] Tile_X6Y9_LUT4AB/N1END[0]
+ Tile_X6Y9_LUT4AB/N1END[1] Tile_X6Y9_LUT4AB/N1END[2] Tile_X6Y9_LUT4AB/N1END[3] Tile_X6Y9_LUT4AB/N2BEG[0]
+ Tile_X6Y9_LUT4AB/N2BEG[1] Tile_X6Y9_LUT4AB/N2BEG[2] Tile_X6Y9_LUT4AB/N2BEG[3] Tile_X6Y9_LUT4AB/N2BEG[4]
+ Tile_X6Y9_LUT4AB/N2BEG[5] Tile_X6Y9_LUT4AB/N2BEG[6] Tile_X6Y9_LUT4AB/N2BEG[7] Tile_X6Y8_LUT4AB/N2END[0]
+ Tile_X6Y8_LUT4AB/N2END[1] Tile_X6Y8_LUT4AB/N2END[2] Tile_X6Y8_LUT4AB/N2END[3] Tile_X6Y8_LUT4AB/N2END[4]
+ Tile_X6Y8_LUT4AB/N2END[5] Tile_X6Y8_LUT4AB/N2END[6] Tile_X6Y8_LUT4AB/N2END[7] Tile_X6Y9_LUT4AB/N2END[0]
+ Tile_X6Y9_LUT4AB/N2END[1] Tile_X6Y9_LUT4AB/N2END[2] Tile_X6Y9_LUT4AB/N2END[3] Tile_X6Y9_LUT4AB/N2END[4]
+ Tile_X6Y9_LUT4AB/N2END[5] Tile_X6Y9_LUT4AB/N2END[6] Tile_X6Y9_LUT4AB/N2END[7] Tile_X6Y9_LUT4AB/N2MID[0]
+ Tile_X6Y9_LUT4AB/N2MID[1] Tile_X6Y9_LUT4AB/N2MID[2] Tile_X6Y9_LUT4AB/N2MID[3] Tile_X6Y9_LUT4AB/N2MID[4]
+ Tile_X6Y9_LUT4AB/N2MID[5] Tile_X6Y9_LUT4AB/N2MID[6] Tile_X6Y9_LUT4AB/N2MID[7] Tile_X6Y9_LUT4AB/N4BEG[0]
+ Tile_X6Y9_LUT4AB/N4BEG[10] Tile_X6Y9_LUT4AB/N4BEG[11] Tile_X6Y9_LUT4AB/N4BEG[12]
+ Tile_X6Y9_LUT4AB/N4BEG[13] Tile_X6Y9_LUT4AB/N4BEG[14] Tile_X6Y9_LUT4AB/N4BEG[15]
+ Tile_X6Y9_LUT4AB/N4BEG[1] Tile_X6Y9_LUT4AB/N4BEG[2] Tile_X6Y9_LUT4AB/N4BEG[3] Tile_X6Y9_LUT4AB/N4BEG[4]
+ Tile_X6Y9_LUT4AB/N4BEG[5] Tile_X6Y9_LUT4AB/N4BEG[6] Tile_X6Y9_LUT4AB/N4BEG[7] Tile_X6Y9_LUT4AB/N4BEG[8]
+ Tile_X6Y9_LUT4AB/N4BEG[9] Tile_X6Y9_LUT4AB/N4END[0] Tile_X6Y9_LUT4AB/N4END[10] Tile_X6Y9_LUT4AB/N4END[11]
+ Tile_X6Y9_LUT4AB/N4END[12] Tile_X6Y9_LUT4AB/N4END[13] Tile_X6Y9_LUT4AB/N4END[14]
+ Tile_X6Y9_LUT4AB/N4END[15] Tile_X6Y9_LUT4AB/N4END[1] Tile_X6Y9_LUT4AB/N4END[2] Tile_X6Y9_LUT4AB/N4END[3]
+ Tile_X6Y9_LUT4AB/N4END[4] Tile_X6Y9_LUT4AB/N4END[5] Tile_X6Y9_LUT4AB/N4END[6] Tile_X6Y9_LUT4AB/N4END[7]
+ Tile_X6Y9_LUT4AB/N4END[8] Tile_X6Y9_LUT4AB/N4END[9] Tile_X6Y9_LUT4AB/NN4BEG[0] Tile_X6Y9_LUT4AB/NN4BEG[10]
+ Tile_X6Y9_LUT4AB/NN4BEG[11] Tile_X6Y9_LUT4AB/NN4BEG[12] Tile_X6Y9_LUT4AB/NN4BEG[13]
+ Tile_X6Y9_LUT4AB/NN4BEG[14] Tile_X6Y9_LUT4AB/NN4BEG[15] Tile_X6Y9_LUT4AB/NN4BEG[1]
+ Tile_X6Y9_LUT4AB/NN4BEG[2] Tile_X6Y9_LUT4AB/NN4BEG[3] Tile_X6Y9_LUT4AB/NN4BEG[4]
+ Tile_X6Y9_LUT4AB/NN4BEG[5] Tile_X6Y9_LUT4AB/NN4BEG[6] Tile_X6Y9_LUT4AB/NN4BEG[7]
+ Tile_X6Y9_LUT4AB/NN4BEG[8] Tile_X6Y9_LUT4AB/NN4BEG[9] Tile_X6Y9_LUT4AB/NN4END[0]
+ Tile_X6Y9_LUT4AB/NN4END[10] Tile_X6Y9_LUT4AB/NN4END[11] Tile_X6Y9_LUT4AB/NN4END[12]
+ Tile_X6Y9_LUT4AB/NN4END[13] Tile_X6Y9_LUT4AB/NN4END[14] Tile_X6Y9_LUT4AB/NN4END[15]
+ Tile_X6Y9_LUT4AB/NN4END[1] Tile_X6Y9_LUT4AB/NN4END[2] Tile_X6Y9_LUT4AB/NN4END[3]
+ Tile_X6Y9_LUT4AB/NN4END[4] Tile_X6Y9_LUT4AB/NN4END[5] Tile_X6Y9_LUT4AB/NN4END[6]
+ Tile_X6Y9_LUT4AB/NN4END[7] Tile_X6Y9_LUT4AB/NN4END[8] Tile_X6Y9_LUT4AB/NN4END[9]
+ Tile_X6Y9_LUT4AB/S1BEG[0] Tile_X6Y9_LUT4AB/S1BEG[1] Tile_X6Y9_LUT4AB/S1BEG[2] Tile_X6Y9_LUT4AB/S1BEG[3]
+ Tile_X6Y9_LUT4AB/S1END[0] Tile_X6Y9_LUT4AB/S1END[1] Tile_X6Y9_LUT4AB/S1END[2] Tile_X6Y9_LUT4AB/S1END[3]
+ Tile_X6Y9_LUT4AB/S2BEG[0] Tile_X6Y9_LUT4AB/S2BEG[1] Tile_X6Y9_LUT4AB/S2BEG[2] Tile_X6Y9_LUT4AB/S2BEG[3]
+ Tile_X6Y9_LUT4AB/S2BEG[4] Tile_X6Y9_LUT4AB/S2BEG[5] Tile_X6Y9_LUT4AB/S2BEG[6] Tile_X6Y9_LUT4AB/S2BEG[7]
+ Tile_X6Y9_LUT4AB/S2BEGb[0] Tile_X6Y9_LUT4AB/S2BEGb[1] Tile_X6Y9_LUT4AB/S2BEGb[2]
+ Tile_X6Y9_LUT4AB/S2BEGb[3] Tile_X6Y9_LUT4AB/S2BEGb[4] Tile_X6Y9_LUT4AB/S2BEGb[5]
+ Tile_X6Y9_LUT4AB/S2BEGb[6] Tile_X6Y9_LUT4AB/S2BEGb[7] Tile_X6Y9_LUT4AB/S2END[0]
+ Tile_X6Y9_LUT4AB/S2END[1] Tile_X6Y9_LUT4AB/S2END[2] Tile_X6Y9_LUT4AB/S2END[3] Tile_X6Y9_LUT4AB/S2END[4]
+ Tile_X6Y9_LUT4AB/S2END[5] Tile_X6Y9_LUT4AB/S2END[6] Tile_X6Y9_LUT4AB/S2END[7] Tile_X6Y9_LUT4AB/S2MID[0]
+ Tile_X6Y9_LUT4AB/S2MID[1] Tile_X6Y9_LUT4AB/S2MID[2] Tile_X6Y9_LUT4AB/S2MID[3] Tile_X6Y9_LUT4AB/S2MID[4]
+ Tile_X6Y9_LUT4AB/S2MID[5] Tile_X6Y9_LUT4AB/S2MID[6] Tile_X6Y9_LUT4AB/S2MID[7] Tile_X6Y9_LUT4AB/S4BEG[0]
+ Tile_X6Y9_LUT4AB/S4BEG[10] Tile_X6Y9_LUT4AB/S4BEG[11] Tile_X6Y9_LUT4AB/S4BEG[12]
+ Tile_X6Y9_LUT4AB/S4BEG[13] Tile_X6Y9_LUT4AB/S4BEG[14] Tile_X6Y9_LUT4AB/S4BEG[15]
+ Tile_X6Y9_LUT4AB/S4BEG[1] Tile_X6Y9_LUT4AB/S4BEG[2] Tile_X6Y9_LUT4AB/S4BEG[3] Tile_X6Y9_LUT4AB/S4BEG[4]
+ Tile_X6Y9_LUT4AB/S4BEG[5] Tile_X6Y9_LUT4AB/S4BEG[6] Tile_X6Y9_LUT4AB/S4BEG[7] Tile_X6Y9_LUT4AB/S4BEG[8]
+ Tile_X6Y9_LUT4AB/S4BEG[9] Tile_X6Y9_LUT4AB/S4END[0] Tile_X6Y9_LUT4AB/S4END[10] Tile_X6Y9_LUT4AB/S4END[11]
+ Tile_X6Y9_LUT4AB/S4END[12] Tile_X6Y9_LUT4AB/S4END[13] Tile_X6Y9_LUT4AB/S4END[14]
+ Tile_X6Y9_LUT4AB/S4END[15] Tile_X6Y9_LUT4AB/S4END[1] Tile_X6Y9_LUT4AB/S4END[2] Tile_X6Y9_LUT4AB/S4END[3]
+ Tile_X6Y9_LUT4AB/S4END[4] Tile_X6Y9_LUT4AB/S4END[5] Tile_X6Y9_LUT4AB/S4END[6] Tile_X6Y9_LUT4AB/S4END[7]
+ Tile_X6Y9_LUT4AB/S4END[8] Tile_X6Y9_LUT4AB/S4END[9] Tile_X6Y9_LUT4AB/SS4BEG[0] Tile_X6Y9_LUT4AB/SS4BEG[10]
+ Tile_X6Y9_LUT4AB/SS4BEG[11] Tile_X6Y9_LUT4AB/SS4BEG[12] Tile_X6Y9_LUT4AB/SS4BEG[13]
+ Tile_X6Y9_LUT4AB/SS4BEG[14] Tile_X6Y9_LUT4AB/SS4BEG[15] Tile_X6Y9_LUT4AB/SS4BEG[1]
+ Tile_X6Y9_LUT4AB/SS4BEG[2] Tile_X6Y9_LUT4AB/SS4BEG[3] Tile_X6Y9_LUT4AB/SS4BEG[4]
+ Tile_X6Y9_LUT4AB/SS4BEG[5] Tile_X6Y9_LUT4AB/SS4BEG[6] Tile_X6Y9_LUT4AB/SS4BEG[7]
+ Tile_X6Y9_LUT4AB/SS4BEG[8] Tile_X6Y9_LUT4AB/SS4BEG[9] Tile_X6Y9_LUT4AB/SS4END[0]
+ Tile_X6Y9_LUT4AB/SS4END[10] Tile_X6Y9_LUT4AB/SS4END[11] Tile_X6Y9_LUT4AB/SS4END[12]
+ Tile_X6Y9_LUT4AB/SS4END[13] Tile_X6Y9_LUT4AB/SS4END[14] Tile_X6Y9_LUT4AB/SS4END[15]
+ Tile_X6Y9_LUT4AB/SS4END[1] Tile_X6Y9_LUT4AB/SS4END[2] Tile_X6Y9_LUT4AB/SS4END[3]
+ Tile_X6Y9_LUT4AB/SS4END[4] Tile_X6Y9_LUT4AB/SS4END[5] Tile_X6Y9_LUT4AB/SS4END[6]
+ Tile_X6Y9_LUT4AB/SS4END[7] Tile_X6Y9_LUT4AB/SS4END[8] Tile_X6Y9_LUT4AB/SS4END[9]
+ Tile_X6Y9_LUT4AB/UserCLK Tile_X6Y8_LUT4AB/UserCLK VGND VPWR Tile_X6Y9_LUT4AB/W1BEG[0]
+ Tile_X6Y9_LUT4AB/W1BEG[1] Tile_X6Y9_LUT4AB/W1BEG[2] Tile_X6Y9_LUT4AB/W1BEG[3] Tile_X6Y9_LUT4AB/W1END[0]
+ Tile_X6Y9_LUT4AB/W1END[1] Tile_X6Y9_LUT4AB/W1END[2] Tile_X6Y9_LUT4AB/W1END[3] Tile_X6Y9_LUT4AB/W2BEG[0]
+ Tile_X6Y9_LUT4AB/W2BEG[1] Tile_X6Y9_LUT4AB/W2BEG[2] Tile_X6Y9_LUT4AB/W2BEG[3] Tile_X6Y9_LUT4AB/W2BEG[4]
+ Tile_X6Y9_LUT4AB/W2BEG[5] Tile_X6Y9_LUT4AB/W2BEG[6] Tile_X6Y9_LUT4AB/W2BEG[7] Tile_X5Y9_LUT4AB/W2END[0]
+ Tile_X5Y9_LUT4AB/W2END[1] Tile_X5Y9_LUT4AB/W2END[2] Tile_X5Y9_LUT4AB/W2END[3] Tile_X5Y9_LUT4AB/W2END[4]
+ Tile_X5Y9_LUT4AB/W2END[5] Tile_X5Y9_LUT4AB/W2END[6] Tile_X5Y9_LUT4AB/W2END[7] Tile_X6Y9_LUT4AB/W2END[0]
+ Tile_X6Y9_LUT4AB/W2END[1] Tile_X6Y9_LUT4AB/W2END[2] Tile_X6Y9_LUT4AB/W2END[3] Tile_X6Y9_LUT4AB/W2END[4]
+ Tile_X6Y9_LUT4AB/W2END[5] Tile_X6Y9_LUT4AB/W2END[6] Tile_X6Y9_LUT4AB/W2END[7] Tile_X6Y9_LUT4AB/W2MID[0]
+ Tile_X6Y9_LUT4AB/W2MID[1] Tile_X6Y9_LUT4AB/W2MID[2] Tile_X6Y9_LUT4AB/W2MID[3] Tile_X6Y9_LUT4AB/W2MID[4]
+ Tile_X6Y9_LUT4AB/W2MID[5] Tile_X6Y9_LUT4AB/W2MID[6] Tile_X6Y9_LUT4AB/W2MID[7] Tile_X6Y9_LUT4AB/W6BEG[0]
+ Tile_X6Y9_LUT4AB/W6BEG[10] Tile_X6Y9_LUT4AB/W6BEG[11] Tile_X6Y9_LUT4AB/W6BEG[1]
+ Tile_X6Y9_LUT4AB/W6BEG[2] Tile_X6Y9_LUT4AB/W6BEG[3] Tile_X6Y9_LUT4AB/W6BEG[4] Tile_X6Y9_LUT4AB/W6BEG[5]
+ Tile_X6Y9_LUT4AB/W6BEG[6] Tile_X6Y9_LUT4AB/W6BEG[7] Tile_X6Y9_LUT4AB/W6BEG[8] Tile_X6Y9_LUT4AB/W6BEG[9]
+ Tile_X6Y9_LUT4AB/W6END[0] Tile_X6Y9_LUT4AB/W6END[10] Tile_X6Y9_LUT4AB/W6END[11]
+ Tile_X6Y9_LUT4AB/W6END[1] Tile_X6Y9_LUT4AB/W6END[2] Tile_X6Y9_LUT4AB/W6END[3] Tile_X6Y9_LUT4AB/W6END[4]
+ Tile_X6Y9_LUT4AB/W6END[5] Tile_X6Y9_LUT4AB/W6END[6] Tile_X6Y9_LUT4AB/W6END[7] Tile_X6Y9_LUT4AB/W6END[8]
+ Tile_X6Y9_LUT4AB/W6END[9] Tile_X6Y9_LUT4AB/WW4BEG[0] Tile_X6Y9_LUT4AB/WW4BEG[10]
+ Tile_X6Y9_LUT4AB/WW4BEG[11] Tile_X6Y9_LUT4AB/WW4BEG[12] Tile_X6Y9_LUT4AB/WW4BEG[13]
+ Tile_X6Y9_LUT4AB/WW4BEG[14] Tile_X6Y9_LUT4AB/WW4BEG[15] Tile_X6Y9_LUT4AB/WW4BEG[1]
+ Tile_X6Y9_LUT4AB/WW4BEG[2] Tile_X6Y9_LUT4AB/WW4BEG[3] Tile_X6Y9_LUT4AB/WW4BEG[4]
+ Tile_X6Y9_LUT4AB/WW4BEG[5] Tile_X6Y9_LUT4AB/WW4BEG[6] Tile_X6Y9_LUT4AB/WW4BEG[7]
+ Tile_X6Y9_LUT4AB/WW4BEG[8] Tile_X6Y9_LUT4AB/WW4BEG[9] Tile_X6Y9_LUT4AB/WW4END[0]
+ Tile_X6Y9_LUT4AB/WW4END[10] Tile_X6Y9_LUT4AB/WW4END[11] Tile_X6Y9_LUT4AB/WW4END[12]
+ Tile_X6Y9_LUT4AB/WW4END[13] Tile_X6Y9_LUT4AB/WW4END[14] Tile_X6Y9_LUT4AB/WW4END[15]
+ Tile_X6Y9_LUT4AB/WW4END[1] Tile_X6Y9_LUT4AB/WW4END[2] Tile_X6Y9_LUT4AB/WW4END[3]
+ Tile_X6Y9_LUT4AB/WW4END[4] Tile_X6Y9_LUT4AB/WW4END[5] Tile_X6Y9_LUT4AB/WW4END[6]
+ Tile_X6Y9_LUT4AB/WW4END[7] Tile_X6Y9_LUT4AB/WW4END[8] Tile_X6Y9_LUT4AB/WW4END[9]
+ LUT4AB
XTile_X2Y0_N_IO Tile_X2Y0_A_I_top Tile_X2Y0_A_O_top Tile_X2Y0_A_T_top Tile_X2Y0_A_config_C_bit0
+ Tile_X2Y0_A_config_C_bit1 Tile_X2Y0_A_config_C_bit2 Tile_X2Y0_A_config_C_bit3 Tile_X2Y0_B_I_top
+ Tile_X2Y0_B_O_top Tile_X2Y0_B_T_top Tile_X2Y0_B_config_C_bit0 Tile_X2Y0_B_config_C_bit1
+ Tile_X2Y0_B_config_C_bit2 Tile_X2Y0_B_config_C_bit3 Tile_X2Y0_N_IO/Ci Tile_X2Y0_N_IO/FrameData[0]
+ Tile_X2Y0_N_IO/FrameData[10] Tile_X2Y0_N_IO/FrameData[11] Tile_X2Y0_N_IO/FrameData[12]
+ Tile_X2Y0_N_IO/FrameData[13] Tile_X2Y0_N_IO/FrameData[14] Tile_X2Y0_N_IO/FrameData[15]
+ Tile_X2Y0_N_IO/FrameData[16] Tile_X2Y0_N_IO/FrameData[17] Tile_X2Y0_N_IO/FrameData[18]
+ Tile_X2Y0_N_IO/FrameData[19] Tile_X2Y0_N_IO/FrameData[1] Tile_X2Y0_N_IO/FrameData[20]
+ Tile_X2Y0_N_IO/FrameData[21] Tile_X2Y0_N_IO/FrameData[22] Tile_X2Y0_N_IO/FrameData[23]
+ Tile_X2Y0_N_IO/FrameData[24] Tile_X2Y0_N_IO/FrameData[25] Tile_X2Y0_N_IO/FrameData[26]
+ Tile_X2Y0_N_IO/FrameData[27] Tile_X2Y0_N_IO/FrameData[28] Tile_X2Y0_N_IO/FrameData[29]
+ Tile_X2Y0_N_IO/FrameData[2] Tile_X2Y0_N_IO/FrameData[30] Tile_X2Y0_N_IO/FrameData[31]
+ Tile_X2Y0_N_IO/FrameData[3] Tile_X2Y0_N_IO/FrameData[4] Tile_X2Y0_N_IO/FrameData[5]
+ Tile_X2Y0_N_IO/FrameData[6] Tile_X2Y0_N_IO/FrameData[7] Tile_X2Y0_N_IO/FrameData[8]
+ Tile_X2Y0_N_IO/FrameData[9] Tile_X2Y0_N_IO/FrameData_O[0] Tile_X2Y0_N_IO/FrameData_O[10]
+ Tile_X2Y0_N_IO/FrameData_O[11] Tile_X2Y0_N_IO/FrameData_O[12] Tile_X2Y0_N_IO/FrameData_O[13]
+ Tile_X2Y0_N_IO/FrameData_O[14] Tile_X2Y0_N_IO/FrameData_O[15] Tile_X2Y0_N_IO/FrameData_O[16]
+ Tile_X2Y0_N_IO/FrameData_O[17] Tile_X2Y0_N_IO/FrameData_O[18] Tile_X2Y0_N_IO/FrameData_O[19]
+ Tile_X2Y0_N_IO/FrameData_O[1] Tile_X2Y0_N_IO/FrameData_O[20] Tile_X2Y0_N_IO/FrameData_O[21]
+ Tile_X2Y0_N_IO/FrameData_O[22] Tile_X2Y0_N_IO/FrameData_O[23] Tile_X2Y0_N_IO/FrameData_O[24]
+ Tile_X2Y0_N_IO/FrameData_O[25] Tile_X2Y0_N_IO/FrameData_O[26] Tile_X2Y0_N_IO/FrameData_O[27]
+ Tile_X2Y0_N_IO/FrameData_O[28] Tile_X2Y0_N_IO/FrameData_O[29] Tile_X2Y0_N_IO/FrameData_O[2]
+ Tile_X2Y0_N_IO/FrameData_O[30] Tile_X2Y0_N_IO/FrameData_O[31] Tile_X2Y0_N_IO/FrameData_O[3]
+ Tile_X2Y0_N_IO/FrameData_O[4] Tile_X2Y0_N_IO/FrameData_O[5] Tile_X2Y0_N_IO/FrameData_O[6]
+ Tile_X2Y0_N_IO/FrameData_O[7] Tile_X2Y0_N_IO/FrameData_O[8] Tile_X2Y0_N_IO/FrameData_O[9]
+ Tile_X2Y0_N_IO/FrameStrobe[0] Tile_X2Y0_N_IO/FrameStrobe[10] Tile_X2Y0_N_IO/FrameStrobe[11]
+ Tile_X2Y0_N_IO/FrameStrobe[12] Tile_X2Y0_N_IO/FrameStrobe[13] Tile_X2Y0_N_IO/FrameStrobe[14]
+ Tile_X2Y0_N_IO/FrameStrobe[15] Tile_X2Y0_N_IO/FrameStrobe[16] Tile_X2Y0_N_IO/FrameStrobe[17]
+ Tile_X2Y0_N_IO/FrameStrobe[18] Tile_X2Y0_N_IO/FrameStrobe[19] Tile_X2Y0_N_IO/FrameStrobe[1]
+ Tile_X2Y0_N_IO/FrameStrobe[2] Tile_X2Y0_N_IO/FrameStrobe[3] Tile_X2Y0_N_IO/FrameStrobe[4]
+ Tile_X2Y0_N_IO/FrameStrobe[5] Tile_X2Y0_N_IO/FrameStrobe[6] Tile_X2Y0_N_IO/FrameStrobe[7]
+ Tile_X2Y0_N_IO/FrameStrobe[8] Tile_X2Y0_N_IO/FrameStrobe[9] Tile_X2Y0_N_IO/FrameStrobe_O[0]
+ Tile_X2Y0_N_IO/FrameStrobe_O[10] Tile_X2Y0_N_IO/FrameStrobe_O[11] Tile_X2Y0_N_IO/FrameStrobe_O[12]
+ Tile_X2Y0_N_IO/FrameStrobe_O[13] Tile_X2Y0_N_IO/FrameStrobe_O[14] Tile_X2Y0_N_IO/FrameStrobe_O[15]
+ Tile_X2Y0_N_IO/FrameStrobe_O[16] Tile_X2Y0_N_IO/FrameStrobe_O[17] Tile_X2Y0_N_IO/FrameStrobe_O[18]
+ Tile_X2Y0_N_IO/FrameStrobe_O[19] Tile_X2Y0_N_IO/FrameStrobe_O[1] Tile_X2Y0_N_IO/FrameStrobe_O[2]
+ Tile_X2Y0_N_IO/FrameStrobe_O[3] Tile_X2Y0_N_IO/FrameStrobe_O[4] Tile_X2Y0_N_IO/FrameStrobe_O[5]
+ Tile_X2Y0_N_IO/FrameStrobe_O[6] Tile_X2Y0_N_IO/FrameStrobe_O[7] Tile_X2Y0_N_IO/FrameStrobe_O[8]
+ Tile_X2Y0_N_IO/FrameStrobe_O[9] Tile_X2Y0_N_IO/N1END[0] Tile_X2Y0_N_IO/N1END[1]
+ Tile_X2Y0_N_IO/N1END[2] Tile_X2Y0_N_IO/N1END[3] Tile_X2Y0_N_IO/N2END[0] Tile_X2Y0_N_IO/N2END[1]
+ Tile_X2Y0_N_IO/N2END[2] Tile_X2Y0_N_IO/N2END[3] Tile_X2Y0_N_IO/N2END[4] Tile_X2Y0_N_IO/N2END[5]
+ Tile_X2Y0_N_IO/N2END[6] Tile_X2Y0_N_IO/N2END[7] Tile_X2Y0_N_IO/N2MID[0] Tile_X2Y0_N_IO/N2MID[1]
+ Tile_X2Y0_N_IO/N2MID[2] Tile_X2Y0_N_IO/N2MID[3] Tile_X2Y0_N_IO/N2MID[4] Tile_X2Y0_N_IO/N2MID[5]
+ Tile_X2Y0_N_IO/N2MID[6] Tile_X2Y0_N_IO/N2MID[7] Tile_X2Y0_N_IO/N4END[0] Tile_X2Y0_N_IO/N4END[10]
+ Tile_X2Y0_N_IO/N4END[11] Tile_X2Y0_N_IO/N4END[12] Tile_X2Y0_N_IO/N4END[13] Tile_X2Y0_N_IO/N4END[14]
+ Tile_X2Y0_N_IO/N4END[15] Tile_X2Y0_N_IO/N4END[1] Tile_X2Y0_N_IO/N4END[2] Tile_X2Y0_N_IO/N4END[3]
+ Tile_X2Y0_N_IO/N4END[4] Tile_X2Y0_N_IO/N4END[5] Tile_X2Y0_N_IO/N4END[6] Tile_X2Y0_N_IO/N4END[7]
+ Tile_X2Y0_N_IO/N4END[8] Tile_X2Y0_N_IO/N4END[9] Tile_X2Y0_N_IO/NN4END[0] Tile_X2Y0_N_IO/NN4END[10]
+ Tile_X2Y0_N_IO/NN4END[11] Tile_X2Y0_N_IO/NN4END[12] Tile_X2Y0_N_IO/NN4END[13] Tile_X2Y0_N_IO/NN4END[14]
+ Tile_X2Y0_N_IO/NN4END[15] Tile_X2Y0_N_IO/NN4END[1] Tile_X2Y0_N_IO/NN4END[2] Tile_X2Y0_N_IO/NN4END[3]
+ Tile_X2Y0_N_IO/NN4END[4] Tile_X2Y0_N_IO/NN4END[5] Tile_X2Y0_N_IO/NN4END[6] Tile_X2Y0_N_IO/NN4END[7]
+ Tile_X2Y0_N_IO/NN4END[8] Tile_X2Y0_N_IO/NN4END[9] Tile_X2Y0_N_IO/S1BEG[0] Tile_X2Y0_N_IO/S1BEG[1]
+ Tile_X2Y0_N_IO/S1BEG[2] Tile_X2Y0_N_IO/S1BEG[3] Tile_X2Y0_N_IO/S2BEG[0] Tile_X2Y0_N_IO/S2BEG[1]
+ Tile_X2Y0_N_IO/S2BEG[2] Tile_X2Y0_N_IO/S2BEG[3] Tile_X2Y0_N_IO/S2BEG[4] Tile_X2Y0_N_IO/S2BEG[5]
+ Tile_X2Y0_N_IO/S2BEG[6] Tile_X2Y0_N_IO/S2BEG[7] Tile_X2Y0_N_IO/S2BEGb[0] Tile_X2Y0_N_IO/S2BEGb[1]
+ Tile_X2Y0_N_IO/S2BEGb[2] Tile_X2Y0_N_IO/S2BEGb[3] Tile_X2Y0_N_IO/S2BEGb[4] Tile_X2Y0_N_IO/S2BEGb[5]
+ Tile_X2Y0_N_IO/S2BEGb[6] Tile_X2Y0_N_IO/S2BEGb[7] Tile_X2Y0_N_IO/S4BEG[0] Tile_X2Y0_N_IO/S4BEG[10]
+ Tile_X2Y0_N_IO/S4BEG[11] Tile_X2Y0_N_IO/S4BEG[12] Tile_X2Y0_N_IO/S4BEG[13] Tile_X2Y0_N_IO/S4BEG[14]
+ Tile_X2Y0_N_IO/S4BEG[15] Tile_X2Y0_N_IO/S4BEG[1] Tile_X2Y0_N_IO/S4BEG[2] Tile_X2Y0_N_IO/S4BEG[3]
+ Tile_X2Y0_N_IO/S4BEG[4] Tile_X2Y0_N_IO/S4BEG[5] Tile_X2Y0_N_IO/S4BEG[6] Tile_X2Y0_N_IO/S4BEG[7]
+ Tile_X2Y0_N_IO/S4BEG[8] Tile_X2Y0_N_IO/S4BEG[9] Tile_X2Y0_N_IO/SS4BEG[0] Tile_X2Y0_N_IO/SS4BEG[10]
+ Tile_X2Y0_N_IO/SS4BEG[11] Tile_X2Y0_N_IO/SS4BEG[12] Tile_X2Y0_N_IO/SS4BEG[13] Tile_X2Y0_N_IO/SS4BEG[14]
+ Tile_X2Y0_N_IO/SS4BEG[15] Tile_X2Y0_N_IO/SS4BEG[1] Tile_X2Y0_N_IO/SS4BEG[2] Tile_X2Y0_N_IO/SS4BEG[3]
+ Tile_X2Y0_N_IO/SS4BEG[4] Tile_X2Y0_N_IO/SS4BEG[5] Tile_X2Y0_N_IO/SS4BEG[6] Tile_X2Y0_N_IO/SS4BEG[7]
+ Tile_X2Y0_N_IO/SS4BEG[8] Tile_X2Y0_N_IO/SS4BEG[9] Tile_X2Y0_N_IO/UserCLK Tile_X2Y0_N_IO/UserCLKo
+ VGND VPWR N_IO
XTile_X3Y4_LUT4AB Tile_X3Y5_LUT4AB/Co Tile_X3Y4_LUT4AB/Co Tile_X3Y4_LUT4AB/E1BEG[0]
+ Tile_X3Y4_LUT4AB/E1BEG[1] Tile_X3Y4_LUT4AB/E1BEG[2] Tile_X3Y4_LUT4AB/E1BEG[3] Tile_X3Y4_LUT4AB/E1END[0]
+ Tile_X3Y4_LUT4AB/E1END[1] Tile_X3Y4_LUT4AB/E1END[2] Tile_X3Y4_LUT4AB/E1END[3] Tile_X3Y4_LUT4AB/E2BEG[0]
+ Tile_X3Y4_LUT4AB/E2BEG[1] Tile_X3Y4_LUT4AB/E2BEG[2] Tile_X3Y4_LUT4AB/E2BEG[3] Tile_X3Y4_LUT4AB/E2BEG[4]
+ Tile_X3Y4_LUT4AB/E2BEG[5] Tile_X3Y4_LUT4AB/E2BEG[6] Tile_X3Y4_LUT4AB/E2BEG[7] Tile_X4Y4_RegFile/E2END[0]
+ Tile_X4Y4_RegFile/E2END[1] Tile_X4Y4_RegFile/E2END[2] Tile_X4Y4_RegFile/E2END[3]
+ Tile_X4Y4_RegFile/E2END[4] Tile_X4Y4_RegFile/E2END[5] Tile_X4Y4_RegFile/E2END[6]
+ Tile_X4Y4_RegFile/E2END[7] Tile_X3Y4_LUT4AB/E2END[0] Tile_X3Y4_LUT4AB/E2END[1] Tile_X3Y4_LUT4AB/E2END[2]
+ Tile_X3Y4_LUT4AB/E2END[3] Tile_X3Y4_LUT4AB/E2END[4] Tile_X3Y4_LUT4AB/E2END[5] Tile_X3Y4_LUT4AB/E2END[6]
+ Tile_X3Y4_LUT4AB/E2END[7] Tile_X3Y4_LUT4AB/E2MID[0] Tile_X3Y4_LUT4AB/E2MID[1] Tile_X3Y4_LUT4AB/E2MID[2]
+ Tile_X3Y4_LUT4AB/E2MID[3] Tile_X3Y4_LUT4AB/E2MID[4] Tile_X3Y4_LUT4AB/E2MID[5] Tile_X3Y4_LUT4AB/E2MID[6]
+ Tile_X3Y4_LUT4AB/E2MID[7] Tile_X3Y4_LUT4AB/E6BEG[0] Tile_X3Y4_LUT4AB/E6BEG[10] Tile_X3Y4_LUT4AB/E6BEG[11]
+ Tile_X3Y4_LUT4AB/E6BEG[1] Tile_X3Y4_LUT4AB/E6BEG[2] Tile_X3Y4_LUT4AB/E6BEG[3] Tile_X3Y4_LUT4AB/E6BEG[4]
+ Tile_X3Y4_LUT4AB/E6BEG[5] Tile_X3Y4_LUT4AB/E6BEG[6] Tile_X3Y4_LUT4AB/E6BEG[7] Tile_X3Y4_LUT4AB/E6BEG[8]
+ Tile_X3Y4_LUT4AB/E6BEG[9] Tile_X3Y4_LUT4AB/E6END[0] Tile_X3Y4_LUT4AB/E6END[10] Tile_X3Y4_LUT4AB/E6END[11]
+ Tile_X3Y4_LUT4AB/E6END[1] Tile_X3Y4_LUT4AB/E6END[2] Tile_X3Y4_LUT4AB/E6END[3] Tile_X3Y4_LUT4AB/E6END[4]
+ Tile_X3Y4_LUT4AB/E6END[5] Tile_X3Y4_LUT4AB/E6END[6] Tile_X3Y4_LUT4AB/E6END[7] Tile_X3Y4_LUT4AB/E6END[8]
+ Tile_X3Y4_LUT4AB/E6END[9] Tile_X3Y4_LUT4AB/EE4BEG[0] Tile_X3Y4_LUT4AB/EE4BEG[10]
+ Tile_X3Y4_LUT4AB/EE4BEG[11] Tile_X3Y4_LUT4AB/EE4BEG[12] Tile_X3Y4_LUT4AB/EE4BEG[13]
+ Tile_X3Y4_LUT4AB/EE4BEG[14] Tile_X3Y4_LUT4AB/EE4BEG[15] Tile_X3Y4_LUT4AB/EE4BEG[1]
+ Tile_X3Y4_LUT4AB/EE4BEG[2] Tile_X3Y4_LUT4AB/EE4BEG[3] Tile_X3Y4_LUT4AB/EE4BEG[4]
+ Tile_X3Y4_LUT4AB/EE4BEG[5] Tile_X3Y4_LUT4AB/EE4BEG[6] Tile_X3Y4_LUT4AB/EE4BEG[7]
+ Tile_X3Y4_LUT4AB/EE4BEG[8] Tile_X3Y4_LUT4AB/EE4BEG[9] Tile_X3Y4_LUT4AB/EE4END[0]
+ Tile_X3Y4_LUT4AB/EE4END[10] Tile_X3Y4_LUT4AB/EE4END[11] Tile_X3Y4_LUT4AB/EE4END[12]
+ Tile_X3Y4_LUT4AB/EE4END[13] Tile_X3Y4_LUT4AB/EE4END[14] Tile_X3Y4_LUT4AB/EE4END[15]
+ Tile_X3Y4_LUT4AB/EE4END[1] Tile_X3Y4_LUT4AB/EE4END[2] Tile_X3Y4_LUT4AB/EE4END[3]
+ Tile_X3Y4_LUT4AB/EE4END[4] Tile_X3Y4_LUT4AB/EE4END[5] Tile_X3Y4_LUT4AB/EE4END[6]
+ Tile_X3Y4_LUT4AB/EE4END[7] Tile_X3Y4_LUT4AB/EE4END[8] Tile_X3Y4_LUT4AB/EE4END[9]
+ Tile_X3Y4_LUT4AB/FrameData[0] Tile_X3Y4_LUT4AB/FrameData[10] Tile_X3Y4_LUT4AB/FrameData[11]
+ Tile_X3Y4_LUT4AB/FrameData[12] Tile_X3Y4_LUT4AB/FrameData[13] Tile_X3Y4_LUT4AB/FrameData[14]
+ Tile_X3Y4_LUT4AB/FrameData[15] Tile_X3Y4_LUT4AB/FrameData[16] Tile_X3Y4_LUT4AB/FrameData[17]
+ Tile_X3Y4_LUT4AB/FrameData[18] Tile_X3Y4_LUT4AB/FrameData[19] Tile_X3Y4_LUT4AB/FrameData[1]
+ Tile_X3Y4_LUT4AB/FrameData[20] Tile_X3Y4_LUT4AB/FrameData[21] Tile_X3Y4_LUT4AB/FrameData[22]
+ Tile_X3Y4_LUT4AB/FrameData[23] Tile_X3Y4_LUT4AB/FrameData[24] Tile_X3Y4_LUT4AB/FrameData[25]
+ Tile_X3Y4_LUT4AB/FrameData[26] Tile_X3Y4_LUT4AB/FrameData[27] Tile_X3Y4_LUT4AB/FrameData[28]
+ Tile_X3Y4_LUT4AB/FrameData[29] Tile_X3Y4_LUT4AB/FrameData[2] Tile_X3Y4_LUT4AB/FrameData[30]
+ Tile_X3Y4_LUT4AB/FrameData[31] Tile_X3Y4_LUT4AB/FrameData[3] Tile_X3Y4_LUT4AB/FrameData[4]
+ Tile_X3Y4_LUT4AB/FrameData[5] Tile_X3Y4_LUT4AB/FrameData[6] Tile_X3Y4_LUT4AB/FrameData[7]
+ Tile_X3Y4_LUT4AB/FrameData[8] Tile_X3Y4_LUT4AB/FrameData[9] Tile_X4Y4_RegFile/FrameData[0]
+ Tile_X4Y4_RegFile/FrameData[10] Tile_X4Y4_RegFile/FrameData[11] Tile_X4Y4_RegFile/FrameData[12]
+ Tile_X4Y4_RegFile/FrameData[13] Tile_X4Y4_RegFile/FrameData[14] Tile_X4Y4_RegFile/FrameData[15]
+ Tile_X4Y4_RegFile/FrameData[16] Tile_X4Y4_RegFile/FrameData[17] Tile_X4Y4_RegFile/FrameData[18]
+ Tile_X4Y4_RegFile/FrameData[19] Tile_X4Y4_RegFile/FrameData[1] Tile_X4Y4_RegFile/FrameData[20]
+ Tile_X4Y4_RegFile/FrameData[21] Tile_X4Y4_RegFile/FrameData[22] Tile_X4Y4_RegFile/FrameData[23]
+ Tile_X4Y4_RegFile/FrameData[24] Tile_X4Y4_RegFile/FrameData[25] Tile_X4Y4_RegFile/FrameData[26]
+ Tile_X4Y4_RegFile/FrameData[27] Tile_X4Y4_RegFile/FrameData[28] Tile_X4Y4_RegFile/FrameData[29]
+ Tile_X4Y4_RegFile/FrameData[2] Tile_X4Y4_RegFile/FrameData[30] Tile_X4Y4_RegFile/FrameData[31]
+ Tile_X4Y4_RegFile/FrameData[3] Tile_X4Y4_RegFile/FrameData[4] Tile_X4Y4_RegFile/FrameData[5]
+ Tile_X4Y4_RegFile/FrameData[6] Tile_X4Y4_RegFile/FrameData[7] Tile_X4Y4_RegFile/FrameData[8]
+ Tile_X4Y4_RegFile/FrameData[9] Tile_X3Y4_LUT4AB/FrameStrobe[0] Tile_X3Y4_LUT4AB/FrameStrobe[10]
+ Tile_X3Y4_LUT4AB/FrameStrobe[11] Tile_X3Y4_LUT4AB/FrameStrobe[12] Tile_X3Y4_LUT4AB/FrameStrobe[13]
+ Tile_X3Y4_LUT4AB/FrameStrobe[14] Tile_X3Y4_LUT4AB/FrameStrobe[15] Tile_X3Y4_LUT4AB/FrameStrobe[16]
+ Tile_X3Y4_LUT4AB/FrameStrobe[17] Tile_X3Y4_LUT4AB/FrameStrobe[18] Tile_X3Y4_LUT4AB/FrameStrobe[19]
+ Tile_X3Y4_LUT4AB/FrameStrobe[1] Tile_X3Y4_LUT4AB/FrameStrobe[2] Tile_X3Y4_LUT4AB/FrameStrobe[3]
+ Tile_X3Y4_LUT4AB/FrameStrobe[4] Tile_X3Y4_LUT4AB/FrameStrobe[5] Tile_X3Y4_LUT4AB/FrameStrobe[6]
+ Tile_X3Y4_LUT4AB/FrameStrobe[7] Tile_X3Y4_LUT4AB/FrameStrobe[8] Tile_X3Y4_LUT4AB/FrameStrobe[9]
+ Tile_X3Y3_LUT4AB/FrameStrobe[0] Tile_X3Y3_LUT4AB/FrameStrobe[10] Tile_X3Y3_LUT4AB/FrameStrobe[11]
+ Tile_X3Y3_LUT4AB/FrameStrobe[12] Tile_X3Y3_LUT4AB/FrameStrobe[13] Tile_X3Y3_LUT4AB/FrameStrobe[14]
+ Tile_X3Y3_LUT4AB/FrameStrobe[15] Tile_X3Y3_LUT4AB/FrameStrobe[16] Tile_X3Y3_LUT4AB/FrameStrobe[17]
+ Tile_X3Y3_LUT4AB/FrameStrobe[18] Tile_X3Y3_LUT4AB/FrameStrobe[19] Tile_X3Y3_LUT4AB/FrameStrobe[1]
+ Tile_X3Y3_LUT4AB/FrameStrobe[2] Tile_X3Y3_LUT4AB/FrameStrobe[3] Tile_X3Y3_LUT4AB/FrameStrobe[4]
+ Tile_X3Y3_LUT4AB/FrameStrobe[5] Tile_X3Y3_LUT4AB/FrameStrobe[6] Tile_X3Y3_LUT4AB/FrameStrobe[7]
+ Tile_X3Y3_LUT4AB/FrameStrobe[8] Tile_X3Y3_LUT4AB/FrameStrobe[9] Tile_X3Y4_LUT4AB/N1BEG[0]
+ Tile_X3Y4_LUT4AB/N1BEG[1] Tile_X3Y4_LUT4AB/N1BEG[2] Tile_X3Y4_LUT4AB/N1BEG[3] Tile_X3Y5_LUT4AB/N1BEG[0]
+ Tile_X3Y5_LUT4AB/N1BEG[1] Tile_X3Y5_LUT4AB/N1BEG[2] Tile_X3Y5_LUT4AB/N1BEG[3] Tile_X3Y4_LUT4AB/N2BEG[0]
+ Tile_X3Y4_LUT4AB/N2BEG[1] Tile_X3Y4_LUT4AB/N2BEG[2] Tile_X3Y4_LUT4AB/N2BEG[3] Tile_X3Y4_LUT4AB/N2BEG[4]
+ Tile_X3Y4_LUT4AB/N2BEG[5] Tile_X3Y4_LUT4AB/N2BEG[6] Tile_X3Y4_LUT4AB/N2BEG[7] Tile_X3Y3_LUT4AB/N2END[0]
+ Tile_X3Y3_LUT4AB/N2END[1] Tile_X3Y3_LUT4AB/N2END[2] Tile_X3Y3_LUT4AB/N2END[3] Tile_X3Y3_LUT4AB/N2END[4]
+ Tile_X3Y3_LUT4AB/N2END[5] Tile_X3Y3_LUT4AB/N2END[6] Tile_X3Y3_LUT4AB/N2END[7] Tile_X3Y4_LUT4AB/N2END[0]
+ Tile_X3Y4_LUT4AB/N2END[1] Tile_X3Y4_LUT4AB/N2END[2] Tile_X3Y4_LUT4AB/N2END[3] Tile_X3Y4_LUT4AB/N2END[4]
+ Tile_X3Y4_LUT4AB/N2END[5] Tile_X3Y4_LUT4AB/N2END[6] Tile_X3Y4_LUT4AB/N2END[7] Tile_X3Y5_LUT4AB/N2BEG[0]
+ Tile_X3Y5_LUT4AB/N2BEG[1] Tile_X3Y5_LUT4AB/N2BEG[2] Tile_X3Y5_LUT4AB/N2BEG[3] Tile_X3Y5_LUT4AB/N2BEG[4]
+ Tile_X3Y5_LUT4AB/N2BEG[5] Tile_X3Y5_LUT4AB/N2BEG[6] Tile_X3Y5_LUT4AB/N2BEG[7] Tile_X3Y4_LUT4AB/N4BEG[0]
+ Tile_X3Y4_LUT4AB/N4BEG[10] Tile_X3Y4_LUT4AB/N4BEG[11] Tile_X3Y4_LUT4AB/N4BEG[12]
+ Tile_X3Y4_LUT4AB/N4BEG[13] Tile_X3Y4_LUT4AB/N4BEG[14] Tile_X3Y4_LUT4AB/N4BEG[15]
+ Tile_X3Y4_LUT4AB/N4BEG[1] Tile_X3Y4_LUT4AB/N4BEG[2] Tile_X3Y4_LUT4AB/N4BEG[3] Tile_X3Y4_LUT4AB/N4BEG[4]
+ Tile_X3Y4_LUT4AB/N4BEG[5] Tile_X3Y4_LUT4AB/N4BEG[6] Tile_X3Y4_LUT4AB/N4BEG[7] Tile_X3Y4_LUT4AB/N4BEG[8]
+ Tile_X3Y4_LUT4AB/N4BEG[9] Tile_X3Y5_LUT4AB/N4BEG[0] Tile_X3Y5_LUT4AB/N4BEG[10] Tile_X3Y5_LUT4AB/N4BEG[11]
+ Tile_X3Y5_LUT4AB/N4BEG[12] Tile_X3Y5_LUT4AB/N4BEG[13] Tile_X3Y5_LUT4AB/N4BEG[14]
+ Tile_X3Y5_LUT4AB/N4BEG[15] Tile_X3Y5_LUT4AB/N4BEG[1] Tile_X3Y5_LUT4AB/N4BEG[2] Tile_X3Y5_LUT4AB/N4BEG[3]
+ Tile_X3Y5_LUT4AB/N4BEG[4] Tile_X3Y5_LUT4AB/N4BEG[5] Tile_X3Y5_LUT4AB/N4BEG[6] Tile_X3Y5_LUT4AB/N4BEG[7]
+ Tile_X3Y5_LUT4AB/N4BEG[8] Tile_X3Y5_LUT4AB/N4BEG[9] Tile_X3Y4_LUT4AB/NN4BEG[0] Tile_X3Y4_LUT4AB/NN4BEG[10]
+ Tile_X3Y4_LUT4AB/NN4BEG[11] Tile_X3Y4_LUT4AB/NN4BEG[12] Tile_X3Y4_LUT4AB/NN4BEG[13]
+ Tile_X3Y4_LUT4AB/NN4BEG[14] Tile_X3Y4_LUT4AB/NN4BEG[15] Tile_X3Y4_LUT4AB/NN4BEG[1]
+ Tile_X3Y4_LUT4AB/NN4BEG[2] Tile_X3Y4_LUT4AB/NN4BEG[3] Tile_X3Y4_LUT4AB/NN4BEG[4]
+ Tile_X3Y4_LUT4AB/NN4BEG[5] Tile_X3Y4_LUT4AB/NN4BEG[6] Tile_X3Y4_LUT4AB/NN4BEG[7]
+ Tile_X3Y4_LUT4AB/NN4BEG[8] Tile_X3Y4_LUT4AB/NN4BEG[9] Tile_X3Y5_LUT4AB/NN4BEG[0]
+ Tile_X3Y5_LUT4AB/NN4BEG[10] Tile_X3Y5_LUT4AB/NN4BEG[11] Tile_X3Y5_LUT4AB/NN4BEG[12]
+ Tile_X3Y5_LUT4AB/NN4BEG[13] Tile_X3Y5_LUT4AB/NN4BEG[14] Tile_X3Y5_LUT4AB/NN4BEG[15]
+ Tile_X3Y5_LUT4AB/NN4BEG[1] Tile_X3Y5_LUT4AB/NN4BEG[2] Tile_X3Y5_LUT4AB/NN4BEG[3]
+ Tile_X3Y5_LUT4AB/NN4BEG[4] Tile_X3Y5_LUT4AB/NN4BEG[5] Tile_X3Y5_LUT4AB/NN4BEG[6]
+ Tile_X3Y5_LUT4AB/NN4BEG[7] Tile_X3Y5_LUT4AB/NN4BEG[8] Tile_X3Y5_LUT4AB/NN4BEG[9]
+ Tile_X3Y5_LUT4AB/S1END[0] Tile_X3Y5_LUT4AB/S1END[1] Tile_X3Y5_LUT4AB/S1END[2] Tile_X3Y5_LUT4AB/S1END[3]
+ Tile_X3Y4_LUT4AB/S1END[0] Tile_X3Y4_LUT4AB/S1END[1] Tile_X3Y4_LUT4AB/S1END[2] Tile_X3Y4_LUT4AB/S1END[3]
+ Tile_X3Y5_LUT4AB/S2MID[0] Tile_X3Y5_LUT4AB/S2MID[1] Tile_X3Y5_LUT4AB/S2MID[2] Tile_X3Y5_LUT4AB/S2MID[3]
+ Tile_X3Y5_LUT4AB/S2MID[4] Tile_X3Y5_LUT4AB/S2MID[5] Tile_X3Y5_LUT4AB/S2MID[6] Tile_X3Y5_LUT4AB/S2MID[7]
+ Tile_X3Y5_LUT4AB/S2END[0] Tile_X3Y5_LUT4AB/S2END[1] Tile_X3Y5_LUT4AB/S2END[2] Tile_X3Y5_LUT4AB/S2END[3]
+ Tile_X3Y5_LUT4AB/S2END[4] Tile_X3Y5_LUT4AB/S2END[5] Tile_X3Y5_LUT4AB/S2END[6] Tile_X3Y5_LUT4AB/S2END[7]
+ Tile_X3Y4_LUT4AB/S2END[0] Tile_X3Y4_LUT4AB/S2END[1] Tile_X3Y4_LUT4AB/S2END[2] Tile_X3Y4_LUT4AB/S2END[3]
+ Tile_X3Y4_LUT4AB/S2END[4] Tile_X3Y4_LUT4AB/S2END[5] Tile_X3Y4_LUT4AB/S2END[6] Tile_X3Y4_LUT4AB/S2END[7]
+ Tile_X3Y4_LUT4AB/S2MID[0] Tile_X3Y4_LUT4AB/S2MID[1] Tile_X3Y4_LUT4AB/S2MID[2] Tile_X3Y4_LUT4AB/S2MID[3]
+ Tile_X3Y4_LUT4AB/S2MID[4] Tile_X3Y4_LUT4AB/S2MID[5] Tile_X3Y4_LUT4AB/S2MID[6] Tile_X3Y4_LUT4AB/S2MID[7]
+ Tile_X3Y5_LUT4AB/S4END[0] Tile_X3Y5_LUT4AB/S4END[10] Tile_X3Y5_LUT4AB/S4END[11]
+ Tile_X3Y5_LUT4AB/S4END[12] Tile_X3Y5_LUT4AB/S4END[13] Tile_X3Y5_LUT4AB/S4END[14]
+ Tile_X3Y5_LUT4AB/S4END[15] Tile_X3Y5_LUT4AB/S4END[1] Tile_X3Y5_LUT4AB/S4END[2] Tile_X3Y5_LUT4AB/S4END[3]
+ Tile_X3Y5_LUT4AB/S4END[4] Tile_X3Y5_LUT4AB/S4END[5] Tile_X3Y5_LUT4AB/S4END[6] Tile_X3Y5_LUT4AB/S4END[7]
+ Tile_X3Y5_LUT4AB/S4END[8] Tile_X3Y5_LUT4AB/S4END[9] Tile_X3Y4_LUT4AB/S4END[0] Tile_X3Y4_LUT4AB/S4END[10]
+ Tile_X3Y4_LUT4AB/S4END[11] Tile_X3Y4_LUT4AB/S4END[12] Tile_X3Y4_LUT4AB/S4END[13]
+ Tile_X3Y4_LUT4AB/S4END[14] Tile_X3Y4_LUT4AB/S4END[15] Tile_X3Y4_LUT4AB/S4END[1]
+ Tile_X3Y4_LUT4AB/S4END[2] Tile_X3Y4_LUT4AB/S4END[3] Tile_X3Y4_LUT4AB/S4END[4] Tile_X3Y4_LUT4AB/S4END[5]
+ Tile_X3Y4_LUT4AB/S4END[6] Tile_X3Y4_LUT4AB/S4END[7] Tile_X3Y4_LUT4AB/S4END[8] Tile_X3Y4_LUT4AB/S4END[9]
+ Tile_X3Y5_LUT4AB/SS4END[0] Tile_X3Y5_LUT4AB/SS4END[10] Tile_X3Y5_LUT4AB/SS4END[11]
+ Tile_X3Y5_LUT4AB/SS4END[12] Tile_X3Y5_LUT4AB/SS4END[13] Tile_X3Y5_LUT4AB/SS4END[14]
+ Tile_X3Y5_LUT4AB/SS4END[15] Tile_X3Y5_LUT4AB/SS4END[1] Tile_X3Y5_LUT4AB/SS4END[2]
+ Tile_X3Y5_LUT4AB/SS4END[3] Tile_X3Y5_LUT4AB/SS4END[4] Tile_X3Y5_LUT4AB/SS4END[5]
+ Tile_X3Y5_LUT4AB/SS4END[6] Tile_X3Y5_LUT4AB/SS4END[7] Tile_X3Y5_LUT4AB/SS4END[8]
+ Tile_X3Y5_LUT4AB/SS4END[9] Tile_X3Y4_LUT4AB/SS4END[0] Tile_X3Y4_LUT4AB/SS4END[10]
+ Tile_X3Y4_LUT4AB/SS4END[11] Tile_X3Y4_LUT4AB/SS4END[12] Tile_X3Y4_LUT4AB/SS4END[13]
+ Tile_X3Y4_LUT4AB/SS4END[14] Tile_X3Y4_LUT4AB/SS4END[15] Tile_X3Y4_LUT4AB/SS4END[1]
+ Tile_X3Y4_LUT4AB/SS4END[2] Tile_X3Y4_LUT4AB/SS4END[3] Tile_X3Y4_LUT4AB/SS4END[4]
+ Tile_X3Y4_LUT4AB/SS4END[5] Tile_X3Y4_LUT4AB/SS4END[6] Tile_X3Y4_LUT4AB/SS4END[7]
+ Tile_X3Y4_LUT4AB/SS4END[8] Tile_X3Y4_LUT4AB/SS4END[9] Tile_X3Y4_LUT4AB/UserCLK Tile_X3Y3_LUT4AB/UserCLK
+ VGND VPWR Tile_X3Y4_LUT4AB/W1BEG[0] Tile_X3Y4_LUT4AB/W1BEG[1] Tile_X3Y4_LUT4AB/W1BEG[2]
+ Tile_X3Y4_LUT4AB/W1BEG[3] Tile_X3Y4_LUT4AB/W1END[0] Tile_X3Y4_LUT4AB/W1END[1] Tile_X3Y4_LUT4AB/W1END[2]
+ Tile_X3Y4_LUT4AB/W1END[3] Tile_X3Y4_LUT4AB/W2BEG[0] Tile_X3Y4_LUT4AB/W2BEG[1] Tile_X3Y4_LUT4AB/W2BEG[2]
+ Tile_X3Y4_LUT4AB/W2BEG[3] Tile_X3Y4_LUT4AB/W2BEG[4] Tile_X3Y4_LUT4AB/W2BEG[5] Tile_X3Y4_LUT4AB/W2BEG[6]
+ Tile_X3Y4_LUT4AB/W2BEG[7] Tile_X2Y4_LUT4AB/W2END[0] Tile_X2Y4_LUT4AB/W2END[1] Tile_X2Y4_LUT4AB/W2END[2]
+ Tile_X2Y4_LUT4AB/W2END[3] Tile_X2Y4_LUT4AB/W2END[4] Tile_X2Y4_LUT4AB/W2END[5] Tile_X2Y4_LUT4AB/W2END[6]
+ Tile_X2Y4_LUT4AB/W2END[7] Tile_X3Y4_LUT4AB/W2END[0] Tile_X3Y4_LUT4AB/W2END[1] Tile_X3Y4_LUT4AB/W2END[2]
+ Tile_X3Y4_LUT4AB/W2END[3] Tile_X3Y4_LUT4AB/W2END[4] Tile_X3Y4_LUT4AB/W2END[5] Tile_X3Y4_LUT4AB/W2END[6]
+ Tile_X3Y4_LUT4AB/W2END[7] Tile_X3Y4_LUT4AB/W2MID[0] Tile_X3Y4_LUT4AB/W2MID[1] Tile_X3Y4_LUT4AB/W2MID[2]
+ Tile_X3Y4_LUT4AB/W2MID[3] Tile_X3Y4_LUT4AB/W2MID[4] Tile_X3Y4_LUT4AB/W2MID[5] Tile_X3Y4_LUT4AB/W2MID[6]
+ Tile_X3Y4_LUT4AB/W2MID[7] Tile_X3Y4_LUT4AB/W6BEG[0] Tile_X3Y4_LUT4AB/W6BEG[10] Tile_X3Y4_LUT4AB/W6BEG[11]
+ Tile_X3Y4_LUT4AB/W6BEG[1] Tile_X3Y4_LUT4AB/W6BEG[2] Tile_X3Y4_LUT4AB/W6BEG[3] Tile_X3Y4_LUT4AB/W6BEG[4]
+ Tile_X3Y4_LUT4AB/W6BEG[5] Tile_X3Y4_LUT4AB/W6BEG[6] Tile_X3Y4_LUT4AB/W6BEG[7] Tile_X3Y4_LUT4AB/W6BEG[8]
+ Tile_X3Y4_LUT4AB/W6BEG[9] Tile_X3Y4_LUT4AB/W6END[0] Tile_X3Y4_LUT4AB/W6END[10] Tile_X3Y4_LUT4AB/W6END[11]
+ Tile_X3Y4_LUT4AB/W6END[1] Tile_X3Y4_LUT4AB/W6END[2] Tile_X3Y4_LUT4AB/W6END[3] Tile_X3Y4_LUT4AB/W6END[4]
+ Tile_X3Y4_LUT4AB/W6END[5] Tile_X3Y4_LUT4AB/W6END[6] Tile_X3Y4_LUT4AB/W6END[7] Tile_X3Y4_LUT4AB/W6END[8]
+ Tile_X3Y4_LUT4AB/W6END[9] Tile_X3Y4_LUT4AB/WW4BEG[0] Tile_X3Y4_LUT4AB/WW4BEG[10]
+ Tile_X3Y4_LUT4AB/WW4BEG[11] Tile_X3Y4_LUT4AB/WW4BEG[12] Tile_X3Y4_LUT4AB/WW4BEG[13]
+ Tile_X3Y4_LUT4AB/WW4BEG[14] Tile_X3Y4_LUT4AB/WW4BEG[15] Tile_X3Y4_LUT4AB/WW4BEG[1]
+ Tile_X3Y4_LUT4AB/WW4BEG[2] Tile_X3Y4_LUT4AB/WW4BEG[3] Tile_X3Y4_LUT4AB/WW4BEG[4]
+ Tile_X3Y4_LUT4AB/WW4BEG[5] Tile_X3Y4_LUT4AB/WW4BEG[6] Tile_X3Y4_LUT4AB/WW4BEG[7]
+ Tile_X3Y4_LUT4AB/WW4BEG[8] Tile_X3Y4_LUT4AB/WW4BEG[9] Tile_X3Y4_LUT4AB/WW4END[0]
+ Tile_X3Y4_LUT4AB/WW4END[10] Tile_X3Y4_LUT4AB/WW4END[11] Tile_X3Y4_LUT4AB/WW4END[12]
+ Tile_X3Y4_LUT4AB/WW4END[13] Tile_X3Y4_LUT4AB/WW4END[14] Tile_X3Y4_LUT4AB/WW4END[15]
+ Tile_X3Y4_LUT4AB/WW4END[1] Tile_X3Y4_LUT4AB/WW4END[2] Tile_X3Y4_LUT4AB/WW4END[3]
+ Tile_X3Y4_LUT4AB/WW4END[4] Tile_X3Y4_LUT4AB/WW4END[5] Tile_X3Y4_LUT4AB/WW4END[6]
+ Tile_X3Y4_LUT4AB/WW4END[7] Tile_X3Y4_LUT4AB/WW4END[8] Tile_X3Y4_LUT4AB/WW4END[9]
+ LUT4AB
XTile_X2Y8_LUT4AB Tile_X2Y9_LUT4AB/Co Tile_X2Y8_LUT4AB/Co Tile_X3Y8_LUT4AB/E1END[0]
+ Tile_X3Y8_LUT4AB/E1END[1] Tile_X3Y8_LUT4AB/E1END[2] Tile_X3Y8_LUT4AB/E1END[3] Tile_X2Y8_LUT4AB/E1END[0]
+ Tile_X2Y8_LUT4AB/E1END[1] Tile_X2Y8_LUT4AB/E1END[2] Tile_X2Y8_LUT4AB/E1END[3] Tile_X3Y8_LUT4AB/E2MID[0]
+ Tile_X3Y8_LUT4AB/E2MID[1] Tile_X3Y8_LUT4AB/E2MID[2] Tile_X3Y8_LUT4AB/E2MID[3] Tile_X3Y8_LUT4AB/E2MID[4]
+ Tile_X3Y8_LUT4AB/E2MID[5] Tile_X3Y8_LUT4AB/E2MID[6] Tile_X3Y8_LUT4AB/E2MID[7] Tile_X3Y8_LUT4AB/E2END[0]
+ Tile_X3Y8_LUT4AB/E2END[1] Tile_X3Y8_LUT4AB/E2END[2] Tile_X3Y8_LUT4AB/E2END[3] Tile_X3Y8_LUT4AB/E2END[4]
+ Tile_X3Y8_LUT4AB/E2END[5] Tile_X3Y8_LUT4AB/E2END[6] Tile_X3Y8_LUT4AB/E2END[7] Tile_X2Y8_LUT4AB/E2END[0]
+ Tile_X2Y8_LUT4AB/E2END[1] Tile_X2Y8_LUT4AB/E2END[2] Tile_X2Y8_LUT4AB/E2END[3] Tile_X2Y8_LUT4AB/E2END[4]
+ Tile_X2Y8_LUT4AB/E2END[5] Tile_X2Y8_LUT4AB/E2END[6] Tile_X2Y8_LUT4AB/E2END[7] Tile_X2Y8_LUT4AB/E2MID[0]
+ Tile_X2Y8_LUT4AB/E2MID[1] Tile_X2Y8_LUT4AB/E2MID[2] Tile_X2Y8_LUT4AB/E2MID[3] Tile_X2Y8_LUT4AB/E2MID[4]
+ Tile_X2Y8_LUT4AB/E2MID[5] Tile_X2Y8_LUT4AB/E2MID[6] Tile_X2Y8_LUT4AB/E2MID[7] Tile_X3Y8_LUT4AB/E6END[0]
+ Tile_X3Y8_LUT4AB/E6END[10] Tile_X3Y8_LUT4AB/E6END[11] Tile_X3Y8_LUT4AB/E6END[1]
+ Tile_X3Y8_LUT4AB/E6END[2] Tile_X3Y8_LUT4AB/E6END[3] Tile_X3Y8_LUT4AB/E6END[4] Tile_X3Y8_LUT4AB/E6END[5]
+ Tile_X3Y8_LUT4AB/E6END[6] Tile_X3Y8_LUT4AB/E6END[7] Tile_X3Y8_LUT4AB/E6END[8] Tile_X3Y8_LUT4AB/E6END[9]
+ Tile_X2Y8_LUT4AB/E6END[0] Tile_X2Y8_LUT4AB/E6END[10] Tile_X2Y8_LUT4AB/E6END[11]
+ Tile_X2Y8_LUT4AB/E6END[1] Tile_X2Y8_LUT4AB/E6END[2] Tile_X2Y8_LUT4AB/E6END[3] Tile_X2Y8_LUT4AB/E6END[4]
+ Tile_X2Y8_LUT4AB/E6END[5] Tile_X2Y8_LUT4AB/E6END[6] Tile_X2Y8_LUT4AB/E6END[7] Tile_X2Y8_LUT4AB/E6END[8]
+ Tile_X2Y8_LUT4AB/E6END[9] Tile_X3Y8_LUT4AB/EE4END[0] Tile_X3Y8_LUT4AB/EE4END[10]
+ Tile_X3Y8_LUT4AB/EE4END[11] Tile_X3Y8_LUT4AB/EE4END[12] Tile_X3Y8_LUT4AB/EE4END[13]
+ Tile_X3Y8_LUT4AB/EE4END[14] Tile_X3Y8_LUT4AB/EE4END[15] Tile_X3Y8_LUT4AB/EE4END[1]
+ Tile_X3Y8_LUT4AB/EE4END[2] Tile_X3Y8_LUT4AB/EE4END[3] Tile_X3Y8_LUT4AB/EE4END[4]
+ Tile_X3Y8_LUT4AB/EE4END[5] Tile_X3Y8_LUT4AB/EE4END[6] Tile_X3Y8_LUT4AB/EE4END[7]
+ Tile_X3Y8_LUT4AB/EE4END[8] Tile_X3Y8_LUT4AB/EE4END[9] Tile_X2Y8_LUT4AB/EE4END[0]
+ Tile_X2Y8_LUT4AB/EE4END[10] Tile_X2Y8_LUT4AB/EE4END[11] Tile_X2Y8_LUT4AB/EE4END[12]
+ Tile_X2Y8_LUT4AB/EE4END[13] Tile_X2Y8_LUT4AB/EE4END[14] Tile_X2Y8_LUT4AB/EE4END[15]
+ Tile_X2Y8_LUT4AB/EE4END[1] Tile_X2Y8_LUT4AB/EE4END[2] Tile_X2Y8_LUT4AB/EE4END[3]
+ Tile_X2Y8_LUT4AB/EE4END[4] Tile_X2Y8_LUT4AB/EE4END[5] Tile_X2Y8_LUT4AB/EE4END[6]
+ Tile_X2Y8_LUT4AB/EE4END[7] Tile_X2Y8_LUT4AB/EE4END[8] Tile_X2Y8_LUT4AB/EE4END[9]
+ Tile_X2Y8_LUT4AB/FrameData[0] Tile_X2Y8_LUT4AB/FrameData[10] Tile_X2Y8_LUT4AB/FrameData[11]
+ Tile_X2Y8_LUT4AB/FrameData[12] Tile_X2Y8_LUT4AB/FrameData[13] Tile_X2Y8_LUT4AB/FrameData[14]
+ Tile_X2Y8_LUT4AB/FrameData[15] Tile_X2Y8_LUT4AB/FrameData[16] Tile_X2Y8_LUT4AB/FrameData[17]
+ Tile_X2Y8_LUT4AB/FrameData[18] Tile_X2Y8_LUT4AB/FrameData[19] Tile_X2Y8_LUT4AB/FrameData[1]
+ Tile_X2Y8_LUT4AB/FrameData[20] Tile_X2Y8_LUT4AB/FrameData[21] Tile_X2Y8_LUT4AB/FrameData[22]
+ Tile_X2Y8_LUT4AB/FrameData[23] Tile_X2Y8_LUT4AB/FrameData[24] Tile_X2Y8_LUT4AB/FrameData[25]
+ Tile_X2Y8_LUT4AB/FrameData[26] Tile_X2Y8_LUT4AB/FrameData[27] Tile_X2Y8_LUT4AB/FrameData[28]
+ Tile_X2Y8_LUT4AB/FrameData[29] Tile_X2Y8_LUT4AB/FrameData[2] Tile_X2Y8_LUT4AB/FrameData[30]
+ Tile_X2Y8_LUT4AB/FrameData[31] Tile_X2Y8_LUT4AB/FrameData[3] Tile_X2Y8_LUT4AB/FrameData[4]
+ Tile_X2Y8_LUT4AB/FrameData[5] Tile_X2Y8_LUT4AB/FrameData[6] Tile_X2Y8_LUT4AB/FrameData[7]
+ Tile_X2Y8_LUT4AB/FrameData[8] Tile_X2Y8_LUT4AB/FrameData[9] Tile_X3Y8_LUT4AB/FrameData[0]
+ Tile_X3Y8_LUT4AB/FrameData[10] Tile_X3Y8_LUT4AB/FrameData[11] Tile_X3Y8_LUT4AB/FrameData[12]
+ Tile_X3Y8_LUT4AB/FrameData[13] Tile_X3Y8_LUT4AB/FrameData[14] Tile_X3Y8_LUT4AB/FrameData[15]
+ Tile_X3Y8_LUT4AB/FrameData[16] Tile_X3Y8_LUT4AB/FrameData[17] Tile_X3Y8_LUT4AB/FrameData[18]
+ Tile_X3Y8_LUT4AB/FrameData[19] Tile_X3Y8_LUT4AB/FrameData[1] Tile_X3Y8_LUT4AB/FrameData[20]
+ Tile_X3Y8_LUT4AB/FrameData[21] Tile_X3Y8_LUT4AB/FrameData[22] Tile_X3Y8_LUT4AB/FrameData[23]
+ Tile_X3Y8_LUT4AB/FrameData[24] Tile_X3Y8_LUT4AB/FrameData[25] Tile_X3Y8_LUT4AB/FrameData[26]
+ Tile_X3Y8_LUT4AB/FrameData[27] Tile_X3Y8_LUT4AB/FrameData[28] Tile_X3Y8_LUT4AB/FrameData[29]
+ Tile_X3Y8_LUT4AB/FrameData[2] Tile_X3Y8_LUT4AB/FrameData[30] Tile_X3Y8_LUT4AB/FrameData[31]
+ Tile_X3Y8_LUT4AB/FrameData[3] Tile_X3Y8_LUT4AB/FrameData[4] Tile_X3Y8_LUT4AB/FrameData[5]
+ Tile_X3Y8_LUT4AB/FrameData[6] Tile_X3Y8_LUT4AB/FrameData[7] Tile_X3Y8_LUT4AB/FrameData[8]
+ Tile_X3Y8_LUT4AB/FrameData[9] Tile_X2Y8_LUT4AB/FrameStrobe[0] Tile_X2Y8_LUT4AB/FrameStrobe[10]
+ Tile_X2Y8_LUT4AB/FrameStrobe[11] Tile_X2Y8_LUT4AB/FrameStrobe[12] Tile_X2Y8_LUT4AB/FrameStrobe[13]
+ Tile_X2Y8_LUT4AB/FrameStrobe[14] Tile_X2Y8_LUT4AB/FrameStrobe[15] Tile_X2Y8_LUT4AB/FrameStrobe[16]
+ Tile_X2Y8_LUT4AB/FrameStrobe[17] Tile_X2Y8_LUT4AB/FrameStrobe[18] Tile_X2Y8_LUT4AB/FrameStrobe[19]
+ Tile_X2Y8_LUT4AB/FrameStrobe[1] Tile_X2Y8_LUT4AB/FrameStrobe[2] Tile_X2Y8_LUT4AB/FrameStrobe[3]
+ Tile_X2Y8_LUT4AB/FrameStrobe[4] Tile_X2Y8_LUT4AB/FrameStrobe[5] Tile_X2Y8_LUT4AB/FrameStrobe[6]
+ Tile_X2Y8_LUT4AB/FrameStrobe[7] Tile_X2Y8_LUT4AB/FrameStrobe[8] Tile_X2Y8_LUT4AB/FrameStrobe[9]
+ Tile_X2Y7_LUT4AB/FrameStrobe[0] Tile_X2Y7_LUT4AB/FrameStrobe[10] Tile_X2Y7_LUT4AB/FrameStrobe[11]
+ Tile_X2Y7_LUT4AB/FrameStrobe[12] Tile_X2Y7_LUT4AB/FrameStrobe[13] Tile_X2Y7_LUT4AB/FrameStrobe[14]
+ Tile_X2Y7_LUT4AB/FrameStrobe[15] Tile_X2Y7_LUT4AB/FrameStrobe[16] Tile_X2Y7_LUT4AB/FrameStrobe[17]
+ Tile_X2Y7_LUT4AB/FrameStrobe[18] Tile_X2Y7_LUT4AB/FrameStrobe[19] Tile_X2Y7_LUT4AB/FrameStrobe[1]
+ Tile_X2Y7_LUT4AB/FrameStrobe[2] Tile_X2Y7_LUT4AB/FrameStrobe[3] Tile_X2Y7_LUT4AB/FrameStrobe[4]
+ Tile_X2Y7_LUT4AB/FrameStrobe[5] Tile_X2Y7_LUT4AB/FrameStrobe[6] Tile_X2Y7_LUT4AB/FrameStrobe[7]
+ Tile_X2Y7_LUT4AB/FrameStrobe[8] Tile_X2Y7_LUT4AB/FrameStrobe[9] Tile_X2Y8_LUT4AB/N1BEG[0]
+ Tile_X2Y8_LUT4AB/N1BEG[1] Tile_X2Y8_LUT4AB/N1BEG[2] Tile_X2Y8_LUT4AB/N1BEG[3] Tile_X2Y9_LUT4AB/N1BEG[0]
+ Tile_X2Y9_LUT4AB/N1BEG[1] Tile_X2Y9_LUT4AB/N1BEG[2] Tile_X2Y9_LUT4AB/N1BEG[3] Tile_X2Y8_LUT4AB/N2BEG[0]
+ Tile_X2Y8_LUT4AB/N2BEG[1] Tile_X2Y8_LUT4AB/N2BEG[2] Tile_X2Y8_LUT4AB/N2BEG[3] Tile_X2Y8_LUT4AB/N2BEG[4]
+ Tile_X2Y8_LUT4AB/N2BEG[5] Tile_X2Y8_LUT4AB/N2BEG[6] Tile_X2Y8_LUT4AB/N2BEG[7] Tile_X2Y7_LUT4AB/N2END[0]
+ Tile_X2Y7_LUT4AB/N2END[1] Tile_X2Y7_LUT4AB/N2END[2] Tile_X2Y7_LUT4AB/N2END[3] Tile_X2Y7_LUT4AB/N2END[4]
+ Tile_X2Y7_LUT4AB/N2END[5] Tile_X2Y7_LUT4AB/N2END[6] Tile_X2Y7_LUT4AB/N2END[7] Tile_X2Y8_LUT4AB/N2END[0]
+ Tile_X2Y8_LUT4AB/N2END[1] Tile_X2Y8_LUT4AB/N2END[2] Tile_X2Y8_LUT4AB/N2END[3] Tile_X2Y8_LUT4AB/N2END[4]
+ Tile_X2Y8_LUT4AB/N2END[5] Tile_X2Y8_LUT4AB/N2END[6] Tile_X2Y8_LUT4AB/N2END[7] Tile_X2Y9_LUT4AB/N2BEG[0]
+ Tile_X2Y9_LUT4AB/N2BEG[1] Tile_X2Y9_LUT4AB/N2BEG[2] Tile_X2Y9_LUT4AB/N2BEG[3] Tile_X2Y9_LUT4AB/N2BEG[4]
+ Tile_X2Y9_LUT4AB/N2BEG[5] Tile_X2Y9_LUT4AB/N2BEG[6] Tile_X2Y9_LUT4AB/N2BEG[7] Tile_X2Y8_LUT4AB/N4BEG[0]
+ Tile_X2Y8_LUT4AB/N4BEG[10] Tile_X2Y8_LUT4AB/N4BEG[11] Tile_X2Y8_LUT4AB/N4BEG[12]
+ Tile_X2Y8_LUT4AB/N4BEG[13] Tile_X2Y8_LUT4AB/N4BEG[14] Tile_X2Y8_LUT4AB/N4BEG[15]
+ Tile_X2Y8_LUT4AB/N4BEG[1] Tile_X2Y8_LUT4AB/N4BEG[2] Tile_X2Y8_LUT4AB/N4BEG[3] Tile_X2Y8_LUT4AB/N4BEG[4]
+ Tile_X2Y8_LUT4AB/N4BEG[5] Tile_X2Y8_LUT4AB/N4BEG[6] Tile_X2Y8_LUT4AB/N4BEG[7] Tile_X2Y8_LUT4AB/N4BEG[8]
+ Tile_X2Y8_LUT4AB/N4BEG[9] Tile_X2Y9_LUT4AB/N4BEG[0] Tile_X2Y9_LUT4AB/N4BEG[10] Tile_X2Y9_LUT4AB/N4BEG[11]
+ Tile_X2Y9_LUT4AB/N4BEG[12] Tile_X2Y9_LUT4AB/N4BEG[13] Tile_X2Y9_LUT4AB/N4BEG[14]
+ Tile_X2Y9_LUT4AB/N4BEG[15] Tile_X2Y9_LUT4AB/N4BEG[1] Tile_X2Y9_LUT4AB/N4BEG[2] Tile_X2Y9_LUT4AB/N4BEG[3]
+ Tile_X2Y9_LUT4AB/N4BEG[4] Tile_X2Y9_LUT4AB/N4BEG[5] Tile_X2Y9_LUT4AB/N4BEG[6] Tile_X2Y9_LUT4AB/N4BEG[7]
+ Tile_X2Y9_LUT4AB/N4BEG[8] Tile_X2Y9_LUT4AB/N4BEG[9] Tile_X2Y8_LUT4AB/NN4BEG[0] Tile_X2Y8_LUT4AB/NN4BEG[10]
+ Tile_X2Y8_LUT4AB/NN4BEG[11] Tile_X2Y8_LUT4AB/NN4BEG[12] Tile_X2Y8_LUT4AB/NN4BEG[13]
+ Tile_X2Y8_LUT4AB/NN4BEG[14] Tile_X2Y8_LUT4AB/NN4BEG[15] Tile_X2Y8_LUT4AB/NN4BEG[1]
+ Tile_X2Y8_LUT4AB/NN4BEG[2] Tile_X2Y8_LUT4AB/NN4BEG[3] Tile_X2Y8_LUT4AB/NN4BEG[4]
+ Tile_X2Y8_LUT4AB/NN4BEG[5] Tile_X2Y8_LUT4AB/NN4BEG[6] Tile_X2Y8_LUT4AB/NN4BEG[7]
+ Tile_X2Y8_LUT4AB/NN4BEG[8] Tile_X2Y8_LUT4AB/NN4BEG[9] Tile_X2Y9_LUT4AB/NN4BEG[0]
+ Tile_X2Y9_LUT4AB/NN4BEG[10] Tile_X2Y9_LUT4AB/NN4BEG[11] Tile_X2Y9_LUT4AB/NN4BEG[12]
+ Tile_X2Y9_LUT4AB/NN4BEG[13] Tile_X2Y9_LUT4AB/NN4BEG[14] Tile_X2Y9_LUT4AB/NN4BEG[15]
+ Tile_X2Y9_LUT4AB/NN4BEG[1] Tile_X2Y9_LUT4AB/NN4BEG[2] Tile_X2Y9_LUT4AB/NN4BEG[3]
+ Tile_X2Y9_LUT4AB/NN4BEG[4] Tile_X2Y9_LUT4AB/NN4BEG[5] Tile_X2Y9_LUT4AB/NN4BEG[6]
+ Tile_X2Y9_LUT4AB/NN4BEG[7] Tile_X2Y9_LUT4AB/NN4BEG[8] Tile_X2Y9_LUT4AB/NN4BEG[9]
+ Tile_X2Y9_LUT4AB/S1END[0] Tile_X2Y9_LUT4AB/S1END[1] Tile_X2Y9_LUT4AB/S1END[2] Tile_X2Y9_LUT4AB/S1END[3]
+ Tile_X2Y8_LUT4AB/S1END[0] Tile_X2Y8_LUT4AB/S1END[1] Tile_X2Y8_LUT4AB/S1END[2] Tile_X2Y8_LUT4AB/S1END[3]
+ Tile_X2Y9_LUT4AB/S2MID[0] Tile_X2Y9_LUT4AB/S2MID[1] Tile_X2Y9_LUT4AB/S2MID[2] Tile_X2Y9_LUT4AB/S2MID[3]
+ Tile_X2Y9_LUT4AB/S2MID[4] Tile_X2Y9_LUT4AB/S2MID[5] Tile_X2Y9_LUT4AB/S2MID[6] Tile_X2Y9_LUT4AB/S2MID[7]
+ Tile_X2Y9_LUT4AB/S2END[0] Tile_X2Y9_LUT4AB/S2END[1] Tile_X2Y9_LUT4AB/S2END[2] Tile_X2Y9_LUT4AB/S2END[3]
+ Tile_X2Y9_LUT4AB/S2END[4] Tile_X2Y9_LUT4AB/S2END[5] Tile_X2Y9_LUT4AB/S2END[6] Tile_X2Y9_LUT4AB/S2END[7]
+ Tile_X2Y8_LUT4AB/S2END[0] Tile_X2Y8_LUT4AB/S2END[1] Tile_X2Y8_LUT4AB/S2END[2] Tile_X2Y8_LUT4AB/S2END[3]
+ Tile_X2Y8_LUT4AB/S2END[4] Tile_X2Y8_LUT4AB/S2END[5] Tile_X2Y8_LUT4AB/S2END[6] Tile_X2Y8_LUT4AB/S2END[7]
+ Tile_X2Y8_LUT4AB/S2MID[0] Tile_X2Y8_LUT4AB/S2MID[1] Tile_X2Y8_LUT4AB/S2MID[2] Tile_X2Y8_LUT4AB/S2MID[3]
+ Tile_X2Y8_LUT4AB/S2MID[4] Tile_X2Y8_LUT4AB/S2MID[5] Tile_X2Y8_LUT4AB/S2MID[6] Tile_X2Y8_LUT4AB/S2MID[7]
+ Tile_X2Y9_LUT4AB/S4END[0] Tile_X2Y9_LUT4AB/S4END[10] Tile_X2Y9_LUT4AB/S4END[11]
+ Tile_X2Y9_LUT4AB/S4END[12] Tile_X2Y9_LUT4AB/S4END[13] Tile_X2Y9_LUT4AB/S4END[14]
+ Tile_X2Y9_LUT4AB/S4END[15] Tile_X2Y9_LUT4AB/S4END[1] Tile_X2Y9_LUT4AB/S4END[2] Tile_X2Y9_LUT4AB/S4END[3]
+ Tile_X2Y9_LUT4AB/S4END[4] Tile_X2Y9_LUT4AB/S4END[5] Tile_X2Y9_LUT4AB/S4END[6] Tile_X2Y9_LUT4AB/S4END[7]
+ Tile_X2Y9_LUT4AB/S4END[8] Tile_X2Y9_LUT4AB/S4END[9] Tile_X2Y8_LUT4AB/S4END[0] Tile_X2Y8_LUT4AB/S4END[10]
+ Tile_X2Y8_LUT4AB/S4END[11] Tile_X2Y8_LUT4AB/S4END[12] Tile_X2Y8_LUT4AB/S4END[13]
+ Tile_X2Y8_LUT4AB/S4END[14] Tile_X2Y8_LUT4AB/S4END[15] Tile_X2Y8_LUT4AB/S4END[1]
+ Tile_X2Y8_LUT4AB/S4END[2] Tile_X2Y8_LUT4AB/S4END[3] Tile_X2Y8_LUT4AB/S4END[4] Tile_X2Y8_LUT4AB/S4END[5]
+ Tile_X2Y8_LUT4AB/S4END[6] Tile_X2Y8_LUT4AB/S4END[7] Tile_X2Y8_LUT4AB/S4END[8] Tile_X2Y8_LUT4AB/S4END[9]
+ Tile_X2Y9_LUT4AB/SS4END[0] Tile_X2Y9_LUT4AB/SS4END[10] Tile_X2Y9_LUT4AB/SS4END[11]
+ Tile_X2Y9_LUT4AB/SS4END[12] Tile_X2Y9_LUT4AB/SS4END[13] Tile_X2Y9_LUT4AB/SS4END[14]
+ Tile_X2Y9_LUT4AB/SS4END[15] Tile_X2Y9_LUT4AB/SS4END[1] Tile_X2Y9_LUT4AB/SS4END[2]
+ Tile_X2Y9_LUT4AB/SS4END[3] Tile_X2Y9_LUT4AB/SS4END[4] Tile_X2Y9_LUT4AB/SS4END[5]
+ Tile_X2Y9_LUT4AB/SS4END[6] Tile_X2Y9_LUT4AB/SS4END[7] Tile_X2Y9_LUT4AB/SS4END[8]
+ Tile_X2Y9_LUT4AB/SS4END[9] Tile_X2Y8_LUT4AB/SS4END[0] Tile_X2Y8_LUT4AB/SS4END[10]
+ Tile_X2Y8_LUT4AB/SS4END[11] Tile_X2Y8_LUT4AB/SS4END[12] Tile_X2Y8_LUT4AB/SS4END[13]
+ Tile_X2Y8_LUT4AB/SS4END[14] Tile_X2Y8_LUT4AB/SS4END[15] Tile_X2Y8_LUT4AB/SS4END[1]
+ Tile_X2Y8_LUT4AB/SS4END[2] Tile_X2Y8_LUT4AB/SS4END[3] Tile_X2Y8_LUT4AB/SS4END[4]
+ Tile_X2Y8_LUT4AB/SS4END[5] Tile_X2Y8_LUT4AB/SS4END[6] Tile_X2Y8_LUT4AB/SS4END[7]
+ Tile_X2Y8_LUT4AB/SS4END[8] Tile_X2Y8_LUT4AB/SS4END[9] Tile_X2Y8_LUT4AB/UserCLK Tile_X2Y7_LUT4AB/UserCLK
+ VGND VPWR Tile_X2Y8_LUT4AB/W1BEG[0] Tile_X2Y8_LUT4AB/W1BEG[1] Tile_X2Y8_LUT4AB/W1BEG[2]
+ Tile_X2Y8_LUT4AB/W1BEG[3] Tile_X3Y8_LUT4AB/W1BEG[0] Tile_X3Y8_LUT4AB/W1BEG[1] Tile_X3Y8_LUT4AB/W1BEG[2]
+ Tile_X3Y8_LUT4AB/W1BEG[3] Tile_X2Y8_LUT4AB/W2BEG[0] Tile_X2Y8_LUT4AB/W2BEG[1] Tile_X2Y8_LUT4AB/W2BEG[2]
+ Tile_X2Y8_LUT4AB/W2BEG[3] Tile_X2Y8_LUT4AB/W2BEG[4] Tile_X2Y8_LUT4AB/W2BEG[5] Tile_X2Y8_LUT4AB/W2BEG[6]
+ Tile_X2Y8_LUT4AB/W2BEG[7] Tile_X1Y8_LUT4AB/W2END[0] Tile_X1Y8_LUT4AB/W2END[1] Tile_X1Y8_LUT4AB/W2END[2]
+ Tile_X1Y8_LUT4AB/W2END[3] Tile_X1Y8_LUT4AB/W2END[4] Tile_X1Y8_LUT4AB/W2END[5] Tile_X1Y8_LUT4AB/W2END[6]
+ Tile_X1Y8_LUT4AB/W2END[7] Tile_X2Y8_LUT4AB/W2END[0] Tile_X2Y8_LUT4AB/W2END[1] Tile_X2Y8_LUT4AB/W2END[2]
+ Tile_X2Y8_LUT4AB/W2END[3] Tile_X2Y8_LUT4AB/W2END[4] Tile_X2Y8_LUT4AB/W2END[5] Tile_X2Y8_LUT4AB/W2END[6]
+ Tile_X2Y8_LUT4AB/W2END[7] Tile_X3Y8_LUT4AB/W2BEG[0] Tile_X3Y8_LUT4AB/W2BEG[1] Tile_X3Y8_LUT4AB/W2BEG[2]
+ Tile_X3Y8_LUT4AB/W2BEG[3] Tile_X3Y8_LUT4AB/W2BEG[4] Tile_X3Y8_LUT4AB/W2BEG[5] Tile_X3Y8_LUT4AB/W2BEG[6]
+ Tile_X3Y8_LUT4AB/W2BEG[7] Tile_X2Y8_LUT4AB/W6BEG[0] Tile_X2Y8_LUT4AB/W6BEG[10] Tile_X2Y8_LUT4AB/W6BEG[11]
+ Tile_X2Y8_LUT4AB/W6BEG[1] Tile_X2Y8_LUT4AB/W6BEG[2] Tile_X2Y8_LUT4AB/W6BEG[3] Tile_X2Y8_LUT4AB/W6BEG[4]
+ Tile_X2Y8_LUT4AB/W6BEG[5] Tile_X2Y8_LUT4AB/W6BEG[6] Tile_X2Y8_LUT4AB/W6BEG[7] Tile_X2Y8_LUT4AB/W6BEG[8]
+ Tile_X2Y8_LUT4AB/W6BEG[9] Tile_X3Y8_LUT4AB/W6BEG[0] Tile_X3Y8_LUT4AB/W6BEG[10] Tile_X3Y8_LUT4AB/W6BEG[11]
+ Tile_X3Y8_LUT4AB/W6BEG[1] Tile_X3Y8_LUT4AB/W6BEG[2] Tile_X3Y8_LUT4AB/W6BEG[3] Tile_X3Y8_LUT4AB/W6BEG[4]
+ Tile_X3Y8_LUT4AB/W6BEG[5] Tile_X3Y8_LUT4AB/W6BEG[6] Tile_X3Y8_LUT4AB/W6BEG[7] Tile_X3Y8_LUT4AB/W6BEG[8]
+ Tile_X3Y8_LUT4AB/W6BEG[9] Tile_X2Y8_LUT4AB/WW4BEG[0] Tile_X2Y8_LUT4AB/WW4BEG[10]
+ Tile_X2Y8_LUT4AB/WW4BEG[11] Tile_X2Y8_LUT4AB/WW4BEG[12] Tile_X2Y8_LUT4AB/WW4BEG[13]
+ Tile_X2Y8_LUT4AB/WW4BEG[14] Tile_X2Y8_LUT4AB/WW4BEG[15] Tile_X2Y8_LUT4AB/WW4BEG[1]
+ Tile_X2Y8_LUT4AB/WW4BEG[2] Tile_X2Y8_LUT4AB/WW4BEG[3] Tile_X2Y8_LUT4AB/WW4BEG[4]
+ Tile_X2Y8_LUT4AB/WW4BEG[5] Tile_X2Y8_LUT4AB/WW4BEG[6] Tile_X2Y8_LUT4AB/WW4BEG[7]
+ Tile_X2Y8_LUT4AB/WW4BEG[8] Tile_X2Y8_LUT4AB/WW4BEG[9] Tile_X3Y8_LUT4AB/WW4BEG[0]
+ Tile_X3Y8_LUT4AB/WW4BEG[10] Tile_X3Y8_LUT4AB/WW4BEG[11] Tile_X3Y8_LUT4AB/WW4BEG[12]
+ Tile_X3Y8_LUT4AB/WW4BEG[13] Tile_X3Y8_LUT4AB/WW4BEG[14] Tile_X3Y8_LUT4AB/WW4BEG[15]
+ Tile_X3Y8_LUT4AB/WW4BEG[1] Tile_X3Y8_LUT4AB/WW4BEG[2] Tile_X3Y8_LUT4AB/WW4BEG[3]
+ Tile_X3Y8_LUT4AB/WW4BEG[4] Tile_X3Y8_LUT4AB/WW4BEG[5] Tile_X3Y8_LUT4AB/WW4BEG[6]
+ Tile_X3Y8_LUT4AB/WW4BEG[7] Tile_X3Y8_LUT4AB/WW4BEG[8] Tile_X3Y8_LUT4AB/WW4BEG[9]
+ LUT4AB
XTile_X5Y14_LUT4AB Tile_X5Y14_LUT4AB/Ci Tile_X5Y14_LUT4AB/Co Tile_X6Y14_LUT4AB/E1END[0]
+ Tile_X6Y14_LUT4AB/E1END[1] Tile_X6Y14_LUT4AB/E1END[2] Tile_X6Y14_LUT4AB/E1END[3]
+ Tile_X5Y14_LUT4AB/E1END[0] Tile_X5Y14_LUT4AB/E1END[1] Tile_X5Y14_LUT4AB/E1END[2]
+ Tile_X5Y14_LUT4AB/E1END[3] Tile_X6Y14_LUT4AB/E2MID[0] Tile_X6Y14_LUT4AB/E2MID[1]
+ Tile_X6Y14_LUT4AB/E2MID[2] Tile_X6Y14_LUT4AB/E2MID[3] Tile_X6Y14_LUT4AB/E2MID[4]
+ Tile_X6Y14_LUT4AB/E2MID[5] Tile_X6Y14_LUT4AB/E2MID[6] Tile_X6Y14_LUT4AB/E2MID[7]
+ Tile_X6Y14_LUT4AB/E2END[0] Tile_X6Y14_LUT4AB/E2END[1] Tile_X6Y14_LUT4AB/E2END[2]
+ Tile_X6Y14_LUT4AB/E2END[3] Tile_X6Y14_LUT4AB/E2END[4] Tile_X6Y14_LUT4AB/E2END[5]
+ Tile_X6Y14_LUT4AB/E2END[6] Tile_X6Y14_LUT4AB/E2END[7] Tile_X5Y14_LUT4AB/E2END[0]
+ Tile_X5Y14_LUT4AB/E2END[1] Tile_X5Y14_LUT4AB/E2END[2] Tile_X5Y14_LUT4AB/E2END[3]
+ Tile_X5Y14_LUT4AB/E2END[4] Tile_X5Y14_LUT4AB/E2END[5] Tile_X5Y14_LUT4AB/E2END[6]
+ Tile_X5Y14_LUT4AB/E2END[7] Tile_X5Y14_LUT4AB/E2MID[0] Tile_X5Y14_LUT4AB/E2MID[1]
+ Tile_X5Y14_LUT4AB/E2MID[2] Tile_X5Y14_LUT4AB/E2MID[3] Tile_X5Y14_LUT4AB/E2MID[4]
+ Tile_X5Y14_LUT4AB/E2MID[5] Tile_X5Y14_LUT4AB/E2MID[6] Tile_X5Y14_LUT4AB/E2MID[7]
+ Tile_X6Y14_LUT4AB/E6END[0] Tile_X6Y14_LUT4AB/E6END[10] Tile_X6Y14_LUT4AB/E6END[11]
+ Tile_X6Y14_LUT4AB/E6END[1] Tile_X6Y14_LUT4AB/E6END[2] Tile_X6Y14_LUT4AB/E6END[3]
+ Tile_X6Y14_LUT4AB/E6END[4] Tile_X6Y14_LUT4AB/E6END[5] Tile_X6Y14_LUT4AB/E6END[6]
+ Tile_X6Y14_LUT4AB/E6END[7] Tile_X6Y14_LUT4AB/E6END[8] Tile_X6Y14_LUT4AB/E6END[9]
+ Tile_X5Y14_LUT4AB/E6END[0] Tile_X5Y14_LUT4AB/E6END[10] Tile_X5Y14_LUT4AB/E6END[11]
+ Tile_X5Y14_LUT4AB/E6END[1] Tile_X5Y14_LUT4AB/E6END[2] Tile_X5Y14_LUT4AB/E6END[3]
+ Tile_X5Y14_LUT4AB/E6END[4] Tile_X5Y14_LUT4AB/E6END[5] Tile_X5Y14_LUT4AB/E6END[6]
+ Tile_X5Y14_LUT4AB/E6END[7] Tile_X5Y14_LUT4AB/E6END[8] Tile_X5Y14_LUT4AB/E6END[9]
+ Tile_X6Y14_LUT4AB/EE4END[0] Tile_X6Y14_LUT4AB/EE4END[10] Tile_X6Y14_LUT4AB/EE4END[11]
+ Tile_X6Y14_LUT4AB/EE4END[12] Tile_X6Y14_LUT4AB/EE4END[13] Tile_X6Y14_LUT4AB/EE4END[14]
+ Tile_X6Y14_LUT4AB/EE4END[15] Tile_X6Y14_LUT4AB/EE4END[1] Tile_X6Y14_LUT4AB/EE4END[2]
+ Tile_X6Y14_LUT4AB/EE4END[3] Tile_X6Y14_LUT4AB/EE4END[4] Tile_X6Y14_LUT4AB/EE4END[5]
+ Tile_X6Y14_LUT4AB/EE4END[6] Tile_X6Y14_LUT4AB/EE4END[7] Tile_X6Y14_LUT4AB/EE4END[8]
+ Tile_X6Y14_LUT4AB/EE4END[9] Tile_X5Y14_LUT4AB/EE4END[0] Tile_X5Y14_LUT4AB/EE4END[10]
+ Tile_X5Y14_LUT4AB/EE4END[11] Tile_X5Y14_LUT4AB/EE4END[12] Tile_X5Y14_LUT4AB/EE4END[13]
+ Tile_X5Y14_LUT4AB/EE4END[14] Tile_X5Y14_LUT4AB/EE4END[15] Tile_X5Y14_LUT4AB/EE4END[1]
+ Tile_X5Y14_LUT4AB/EE4END[2] Tile_X5Y14_LUT4AB/EE4END[3] Tile_X5Y14_LUT4AB/EE4END[4]
+ Tile_X5Y14_LUT4AB/EE4END[5] Tile_X5Y14_LUT4AB/EE4END[6] Tile_X5Y14_LUT4AB/EE4END[7]
+ Tile_X5Y14_LUT4AB/EE4END[8] Tile_X5Y14_LUT4AB/EE4END[9] Tile_X5Y14_LUT4AB/FrameData[0]
+ Tile_X5Y14_LUT4AB/FrameData[10] Tile_X5Y14_LUT4AB/FrameData[11] Tile_X5Y14_LUT4AB/FrameData[12]
+ Tile_X5Y14_LUT4AB/FrameData[13] Tile_X5Y14_LUT4AB/FrameData[14] Tile_X5Y14_LUT4AB/FrameData[15]
+ Tile_X5Y14_LUT4AB/FrameData[16] Tile_X5Y14_LUT4AB/FrameData[17] Tile_X5Y14_LUT4AB/FrameData[18]
+ Tile_X5Y14_LUT4AB/FrameData[19] Tile_X5Y14_LUT4AB/FrameData[1] Tile_X5Y14_LUT4AB/FrameData[20]
+ Tile_X5Y14_LUT4AB/FrameData[21] Tile_X5Y14_LUT4AB/FrameData[22] Tile_X5Y14_LUT4AB/FrameData[23]
+ Tile_X5Y14_LUT4AB/FrameData[24] Tile_X5Y14_LUT4AB/FrameData[25] Tile_X5Y14_LUT4AB/FrameData[26]
+ Tile_X5Y14_LUT4AB/FrameData[27] Tile_X5Y14_LUT4AB/FrameData[28] Tile_X5Y14_LUT4AB/FrameData[29]
+ Tile_X5Y14_LUT4AB/FrameData[2] Tile_X5Y14_LUT4AB/FrameData[30] Tile_X5Y14_LUT4AB/FrameData[31]
+ Tile_X5Y14_LUT4AB/FrameData[3] Tile_X5Y14_LUT4AB/FrameData[4] Tile_X5Y14_LUT4AB/FrameData[5]
+ Tile_X5Y14_LUT4AB/FrameData[6] Tile_X5Y14_LUT4AB/FrameData[7] Tile_X5Y14_LUT4AB/FrameData[8]
+ Tile_X5Y14_LUT4AB/FrameData[9] Tile_X6Y14_LUT4AB/FrameData[0] Tile_X6Y14_LUT4AB/FrameData[10]
+ Tile_X6Y14_LUT4AB/FrameData[11] Tile_X6Y14_LUT4AB/FrameData[12] Tile_X6Y14_LUT4AB/FrameData[13]
+ Tile_X6Y14_LUT4AB/FrameData[14] Tile_X6Y14_LUT4AB/FrameData[15] Tile_X6Y14_LUT4AB/FrameData[16]
+ Tile_X6Y14_LUT4AB/FrameData[17] Tile_X6Y14_LUT4AB/FrameData[18] Tile_X6Y14_LUT4AB/FrameData[19]
+ Tile_X6Y14_LUT4AB/FrameData[1] Tile_X6Y14_LUT4AB/FrameData[20] Tile_X6Y14_LUT4AB/FrameData[21]
+ Tile_X6Y14_LUT4AB/FrameData[22] Tile_X6Y14_LUT4AB/FrameData[23] Tile_X6Y14_LUT4AB/FrameData[24]
+ Tile_X6Y14_LUT4AB/FrameData[25] Tile_X6Y14_LUT4AB/FrameData[26] Tile_X6Y14_LUT4AB/FrameData[27]
+ Tile_X6Y14_LUT4AB/FrameData[28] Tile_X6Y14_LUT4AB/FrameData[29] Tile_X6Y14_LUT4AB/FrameData[2]
+ Tile_X6Y14_LUT4AB/FrameData[30] Tile_X6Y14_LUT4AB/FrameData[31] Tile_X6Y14_LUT4AB/FrameData[3]
+ Tile_X6Y14_LUT4AB/FrameData[4] Tile_X6Y14_LUT4AB/FrameData[5] Tile_X6Y14_LUT4AB/FrameData[6]
+ Tile_X6Y14_LUT4AB/FrameData[7] Tile_X6Y14_LUT4AB/FrameData[8] Tile_X6Y14_LUT4AB/FrameData[9]
+ Tile_X5Y14_LUT4AB/FrameStrobe[0] Tile_X5Y14_LUT4AB/FrameStrobe[10] Tile_X5Y14_LUT4AB/FrameStrobe[11]
+ Tile_X5Y14_LUT4AB/FrameStrobe[12] Tile_X5Y14_LUT4AB/FrameStrobe[13] Tile_X5Y14_LUT4AB/FrameStrobe[14]
+ Tile_X5Y14_LUT4AB/FrameStrobe[15] Tile_X5Y14_LUT4AB/FrameStrobe[16] Tile_X5Y14_LUT4AB/FrameStrobe[17]
+ Tile_X5Y14_LUT4AB/FrameStrobe[18] Tile_X5Y14_LUT4AB/FrameStrobe[19] Tile_X5Y14_LUT4AB/FrameStrobe[1]
+ Tile_X5Y14_LUT4AB/FrameStrobe[2] Tile_X5Y14_LUT4AB/FrameStrobe[3] Tile_X5Y14_LUT4AB/FrameStrobe[4]
+ Tile_X5Y14_LUT4AB/FrameStrobe[5] Tile_X5Y14_LUT4AB/FrameStrobe[6] Tile_X5Y14_LUT4AB/FrameStrobe[7]
+ Tile_X5Y14_LUT4AB/FrameStrobe[8] Tile_X5Y14_LUT4AB/FrameStrobe[9] Tile_X5Y13_LUT4AB/FrameStrobe[0]
+ Tile_X5Y13_LUT4AB/FrameStrobe[10] Tile_X5Y13_LUT4AB/FrameStrobe[11] Tile_X5Y13_LUT4AB/FrameStrobe[12]
+ Tile_X5Y13_LUT4AB/FrameStrobe[13] Tile_X5Y13_LUT4AB/FrameStrobe[14] Tile_X5Y13_LUT4AB/FrameStrobe[15]
+ Tile_X5Y13_LUT4AB/FrameStrobe[16] Tile_X5Y13_LUT4AB/FrameStrobe[17] Tile_X5Y13_LUT4AB/FrameStrobe[18]
+ Tile_X5Y13_LUT4AB/FrameStrobe[19] Tile_X5Y13_LUT4AB/FrameStrobe[1] Tile_X5Y13_LUT4AB/FrameStrobe[2]
+ Tile_X5Y13_LUT4AB/FrameStrobe[3] Tile_X5Y13_LUT4AB/FrameStrobe[4] Tile_X5Y13_LUT4AB/FrameStrobe[5]
+ Tile_X5Y13_LUT4AB/FrameStrobe[6] Tile_X5Y13_LUT4AB/FrameStrobe[7] Tile_X5Y13_LUT4AB/FrameStrobe[8]
+ Tile_X5Y13_LUT4AB/FrameStrobe[9] Tile_X5Y14_LUT4AB/N1BEG[0] Tile_X5Y14_LUT4AB/N1BEG[1]
+ Tile_X5Y14_LUT4AB/N1BEG[2] Tile_X5Y14_LUT4AB/N1BEG[3] Tile_X5Y14_LUT4AB/N1END[0]
+ Tile_X5Y14_LUT4AB/N1END[1] Tile_X5Y14_LUT4AB/N1END[2] Tile_X5Y14_LUT4AB/N1END[3]
+ Tile_X5Y14_LUT4AB/N2BEG[0] Tile_X5Y14_LUT4AB/N2BEG[1] Tile_X5Y14_LUT4AB/N2BEG[2]
+ Tile_X5Y14_LUT4AB/N2BEG[3] Tile_X5Y14_LUT4AB/N2BEG[4] Tile_X5Y14_LUT4AB/N2BEG[5]
+ Tile_X5Y14_LUT4AB/N2BEG[6] Tile_X5Y14_LUT4AB/N2BEG[7] Tile_X5Y13_LUT4AB/N2END[0]
+ Tile_X5Y13_LUT4AB/N2END[1] Tile_X5Y13_LUT4AB/N2END[2] Tile_X5Y13_LUT4AB/N2END[3]
+ Tile_X5Y13_LUT4AB/N2END[4] Tile_X5Y13_LUT4AB/N2END[5] Tile_X5Y13_LUT4AB/N2END[6]
+ Tile_X5Y13_LUT4AB/N2END[7] Tile_X5Y14_LUT4AB/N2END[0] Tile_X5Y14_LUT4AB/N2END[1]
+ Tile_X5Y14_LUT4AB/N2END[2] Tile_X5Y14_LUT4AB/N2END[3] Tile_X5Y14_LUT4AB/N2END[4]
+ Tile_X5Y14_LUT4AB/N2END[5] Tile_X5Y14_LUT4AB/N2END[6] Tile_X5Y14_LUT4AB/N2END[7]
+ Tile_X5Y14_LUT4AB/N2MID[0] Tile_X5Y14_LUT4AB/N2MID[1] Tile_X5Y14_LUT4AB/N2MID[2]
+ Tile_X5Y14_LUT4AB/N2MID[3] Tile_X5Y14_LUT4AB/N2MID[4] Tile_X5Y14_LUT4AB/N2MID[5]
+ Tile_X5Y14_LUT4AB/N2MID[6] Tile_X5Y14_LUT4AB/N2MID[7] Tile_X5Y14_LUT4AB/N4BEG[0]
+ Tile_X5Y14_LUT4AB/N4BEG[10] Tile_X5Y14_LUT4AB/N4BEG[11] Tile_X5Y14_LUT4AB/N4BEG[12]
+ Tile_X5Y14_LUT4AB/N4BEG[13] Tile_X5Y14_LUT4AB/N4BEG[14] Tile_X5Y14_LUT4AB/N4BEG[15]
+ Tile_X5Y14_LUT4AB/N4BEG[1] Tile_X5Y14_LUT4AB/N4BEG[2] Tile_X5Y14_LUT4AB/N4BEG[3]
+ Tile_X5Y14_LUT4AB/N4BEG[4] Tile_X5Y14_LUT4AB/N4BEG[5] Tile_X5Y14_LUT4AB/N4BEG[6]
+ Tile_X5Y14_LUT4AB/N4BEG[7] Tile_X5Y14_LUT4AB/N4BEG[8] Tile_X5Y14_LUT4AB/N4BEG[9]
+ Tile_X5Y14_LUT4AB/N4END[0] Tile_X5Y14_LUT4AB/N4END[10] Tile_X5Y14_LUT4AB/N4END[11]
+ Tile_X5Y14_LUT4AB/N4END[12] Tile_X5Y14_LUT4AB/N4END[13] Tile_X5Y14_LUT4AB/N4END[14]
+ Tile_X5Y14_LUT4AB/N4END[15] Tile_X5Y14_LUT4AB/N4END[1] Tile_X5Y14_LUT4AB/N4END[2]
+ Tile_X5Y14_LUT4AB/N4END[3] Tile_X5Y14_LUT4AB/N4END[4] Tile_X5Y14_LUT4AB/N4END[5]
+ Tile_X5Y14_LUT4AB/N4END[6] Tile_X5Y14_LUT4AB/N4END[7] Tile_X5Y14_LUT4AB/N4END[8]
+ Tile_X5Y14_LUT4AB/N4END[9] Tile_X5Y14_LUT4AB/NN4BEG[0] Tile_X5Y14_LUT4AB/NN4BEG[10]
+ Tile_X5Y14_LUT4AB/NN4BEG[11] Tile_X5Y14_LUT4AB/NN4BEG[12] Tile_X5Y14_LUT4AB/NN4BEG[13]
+ Tile_X5Y14_LUT4AB/NN4BEG[14] Tile_X5Y14_LUT4AB/NN4BEG[15] Tile_X5Y14_LUT4AB/NN4BEG[1]
+ Tile_X5Y14_LUT4AB/NN4BEG[2] Tile_X5Y14_LUT4AB/NN4BEG[3] Tile_X5Y14_LUT4AB/NN4BEG[4]
+ Tile_X5Y14_LUT4AB/NN4BEG[5] Tile_X5Y14_LUT4AB/NN4BEG[6] Tile_X5Y14_LUT4AB/NN4BEG[7]
+ Tile_X5Y14_LUT4AB/NN4BEG[8] Tile_X5Y14_LUT4AB/NN4BEG[9] Tile_X5Y14_LUT4AB/NN4END[0]
+ Tile_X5Y14_LUT4AB/NN4END[10] Tile_X5Y14_LUT4AB/NN4END[11] Tile_X5Y14_LUT4AB/NN4END[12]
+ Tile_X5Y14_LUT4AB/NN4END[13] Tile_X5Y14_LUT4AB/NN4END[14] Tile_X5Y14_LUT4AB/NN4END[15]
+ Tile_X5Y14_LUT4AB/NN4END[1] Tile_X5Y14_LUT4AB/NN4END[2] Tile_X5Y14_LUT4AB/NN4END[3]
+ Tile_X5Y14_LUT4AB/NN4END[4] Tile_X5Y14_LUT4AB/NN4END[5] Tile_X5Y14_LUT4AB/NN4END[6]
+ Tile_X5Y14_LUT4AB/NN4END[7] Tile_X5Y14_LUT4AB/NN4END[8] Tile_X5Y14_LUT4AB/NN4END[9]
+ Tile_X5Y14_LUT4AB/S1BEG[0] Tile_X5Y14_LUT4AB/S1BEG[1] Tile_X5Y14_LUT4AB/S1BEG[2]
+ Tile_X5Y14_LUT4AB/S1BEG[3] Tile_X5Y14_LUT4AB/S1END[0] Tile_X5Y14_LUT4AB/S1END[1]
+ Tile_X5Y14_LUT4AB/S1END[2] Tile_X5Y14_LUT4AB/S1END[3] Tile_X5Y14_LUT4AB/S2BEG[0]
+ Tile_X5Y14_LUT4AB/S2BEG[1] Tile_X5Y14_LUT4AB/S2BEG[2] Tile_X5Y14_LUT4AB/S2BEG[3]
+ Tile_X5Y14_LUT4AB/S2BEG[4] Tile_X5Y14_LUT4AB/S2BEG[5] Tile_X5Y14_LUT4AB/S2BEG[6]
+ Tile_X5Y14_LUT4AB/S2BEG[7] Tile_X5Y14_LUT4AB/S2BEGb[0] Tile_X5Y14_LUT4AB/S2BEGb[1]
+ Tile_X5Y14_LUT4AB/S2BEGb[2] Tile_X5Y14_LUT4AB/S2BEGb[3] Tile_X5Y14_LUT4AB/S2BEGb[4]
+ Tile_X5Y14_LUT4AB/S2BEGb[5] Tile_X5Y14_LUT4AB/S2BEGb[6] Tile_X5Y14_LUT4AB/S2BEGb[7]
+ Tile_X5Y14_LUT4AB/S2END[0] Tile_X5Y14_LUT4AB/S2END[1] Tile_X5Y14_LUT4AB/S2END[2]
+ Tile_X5Y14_LUT4AB/S2END[3] Tile_X5Y14_LUT4AB/S2END[4] Tile_X5Y14_LUT4AB/S2END[5]
+ Tile_X5Y14_LUT4AB/S2END[6] Tile_X5Y14_LUT4AB/S2END[7] Tile_X5Y14_LUT4AB/S2MID[0]
+ Tile_X5Y14_LUT4AB/S2MID[1] Tile_X5Y14_LUT4AB/S2MID[2] Tile_X5Y14_LUT4AB/S2MID[3]
+ Tile_X5Y14_LUT4AB/S2MID[4] Tile_X5Y14_LUT4AB/S2MID[5] Tile_X5Y14_LUT4AB/S2MID[6]
+ Tile_X5Y14_LUT4AB/S2MID[7] Tile_X5Y14_LUT4AB/S4BEG[0] Tile_X5Y14_LUT4AB/S4BEG[10]
+ Tile_X5Y14_LUT4AB/S4BEG[11] Tile_X5Y14_LUT4AB/S4BEG[12] Tile_X5Y14_LUT4AB/S4BEG[13]
+ Tile_X5Y14_LUT4AB/S4BEG[14] Tile_X5Y14_LUT4AB/S4BEG[15] Tile_X5Y14_LUT4AB/S4BEG[1]
+ Tile_X5Y14_LUT4AB/S4BEG[2] Tile_X5Y14_LUT4AB/S4BEG[3] Tile_X5Y14_LUT4AB/S4BEG[4]
+ Tile_X5Y14_LUT4AB/S4BEG[5] Tile_X5Y14_LUT4AB/S4BEG[6] Tile_X5Y14_LUT4AB/S4BEG[7]
+ Tile_X5Y14_LUT4AB/S4BEG[8] Tile_X5Y14_LUT4AB/S4BEG[9] Tile_X5Y14_LUT4AB/S4END[0]
+ Tile_X5Y14_LUT4AB/S4END[10] Tile_X5Y14_LUT4AB/S4END[11] Tile_X5Y14_LUT4AB/S4END[12]
+ Tile_X5Y14_LUT4AB/S4END[13] Tile_X5Y14_LUT4AB/S4END[14] Tile_X5Y14_LUT4AB/S4END[15]
+ Tile_X5Y14_LUT4AB/S4END[1] Tile_X5Y14_LUT4AB/S4END[2] Tile_X5Y14_LUT4AB/S4END[3]
+ Tile_X5Y14_LUT4AB/S4END[4] Tile_X5Y14_LUT4AB/S4END[5] Tile_X5Y14_LUT4AB/S4END[6]
+ Tile_X5Y14_LUT4AB/S4END[7] Tile_X5Y14_LUT4AB/S4END[8] Tile_X5Y14_LUT4AB/S4END[9]
+ Tile_X5Y14_LUT4AB/SS4BEG[0] Tile_X5Y14_LUT4AB/SS4BEG[10] Tile_X5Y14_LUT4AB/SS4BEG[11]
+ Tile_X5Y14_LUT4AB/SS4BEG[12] Tile_X5Y14_LUT4AB/SS4BEG[13] Tile_X5Y14_LUT4AB/SS4BEG[14]
+ Tile_X5Y14_LUT4AB/SS4BEG[15] Tile_X5Y14_LUT4AB/SS4BEG[1] Tile_X5Y14_LUT4AB/SS4BEG[2]
+ Tile_X5Y14_LUT4AB/SS4BEG[3] Tile_X5Y14_LUT4AB/SS4BEG[4] Tile_X5Y14_LUT4AB/SS4BEG[5]
+ Tile_X5Y14_LUT4AB/SS4BEG[6] Tile_X5Y14_LUT4AB/SS4BEG[7] Tile_X5Y14_LUT4AB/SS4BEG[8]
+ Tile_X5Y14_LUT4AB/SS4BEG[9] Tile_X5Y14_LUT4AB/SS4END[0] Tile_X5Y14_LUT4AB/SS4END[10]
+ Tile_X5Y14_LUT4AB/SS4END[11] Tile_X5Y14_LUT4AB/SS4END[12] Tile_X5Y14_LUT4AB/SS4END[13]
+ Tile_X5Y14_LUT4AB/SS4END[14] Tile_X5Y14_LUT4AB/SS4END[15] Tile_X5Y14_LUT4AB/SS4END[1]
+ Tile_X5Y14_LUT4AB/SS4END[2] Tile_X5Y14_LUT4AB/SS4END[3] Tile_X5Y14_LUT4AB/SS4END[4]
+ Tile_X5Y14_LUT4AB/SS4END[5] Tile_X5Y14_LUT4AB/SS4END[6] Tile_X5Y14_LUT4AB/SS4END[7]
+ Tile_X5Y14_LUT4AB/SS4END[8] Tile_X5Y14_LUT4AB/SS4END[9] Tile_X5Y14_LUT4AB/UserCLK
+ Tile_X5Y13_LUT4AB/UserCLK VGND VPWR Tile_X5Y14_LUT4AB/W1BEG[0] Tile_X5Y14_LUT4AB/W1BEG[1]
+ Tile_X5Y14_LUT4AB/W1BEG[2] Tile_X5Y14_LUT4AB/W1BEG[3] Tile_X6Y14_LUT4AB/W1BEG[0]
+ Tile_X6Y14_LUT4AB/W1BEG[1] Tile_X6Y14_LUT4AB/W1BEG[2] Tile_X6Y14_LUT4AB/W1BEG[3]
+ Tile_X5Y14_LUT4AB/W2BEG[0] Tile_X5Y14_LUT4AB/W2BEG[1] Tile_X5Y14_LUT4AB/W2BEG[2]
+ Tile_X5Y14_LUT4AB/W2BEG[3] Tile_X5Y14_LUT4AB/W2BEG[4] Tile_X5Y14_LUT4AB/W2BEG[5]
+ Tile_X5Y14_LUT4AB/W2BEG[6] Tile_X5Y14_LUT4AB/W2BEG[7] Tile_X5Y14_LUT4AB/W2BEGb[0]
+ Tile_X5Y14_LUT4AB/W2BEGb[1] Tile_X5Y14_LUT4AB/W2BEGb[2] Tile_X5Y14_LUT4AB/W2BEGb[3]
+ Tile_X5Y14_LUT4AB/W2BEGb[4] Tile_X5Y14_LUT4AB/W2BEGb[5] Tile_X5Y14_LUT4AB/W2BEGb[6]
+ Tile_X5Y14_LUT4AB/W2BEGb[7] Tile_X5Y14_LUT4AB/W2END[0] Tile_X5Y14_LUT4AB/W2END[1]
+ Tile_X5Y14_LUT4AB/W2END[2] Tile_X5Y14_LUT4AB/W2END[3] Tile_X5Y14_LUT4AB/W2END[4]
+ Tile_X5Y14_LUT4AB/W2END[5] Tile_X5Y14_LUT4AB/W2END[6] Tile_X5Y14_LUT4AB/W2END[7]
+ Tile_X6Y14_LUT4AB/W2BEG[0] Tile_X6Y14_LUT4AB/W2BEG[1] Tile_X6Y14_LUT4AB/W2BEG[2]
+ Tile_X6Y14_LUT4AB/W2BEG[3] Tile_X6Y14_LUT4AB/W2BEG[4] Tile_X6Y14_LUT4AB/W2BEG[5]
+ Tile_X6Y14_LUT4AB/W2BEG[6] Tile_X6Y14_LUT4AB/W2BEG[7] Tile_X5Y14_LUT4AB/W6BEG[0]
+ Tile_X5Y14_LUT4AB/W6BEG[10] Tile_X5Y14_LUT4AB/W6BEG[11] Tile_X5Y14_LUT4AB/W6BEG[1]
+ Tile_X5Y14_LUT4AB/W6BEG[2] Tile_X5Y14_LUT4AB/W6BEG[3] Tile_X5Y14_LUT4AB/W6BEG[4]
+ Tile_X5Y14_LUT4AB/W6BEG[5] Tile_X5Y14_LUT4AB/W6BEG[6] Tile_X5Y14_LUT4AB/W6BEG[7]
+ Tile_X5Y14_LUT4AB/W6BEG[8] Tile_X5Y14_LUT4AB/W6BEG[9] Tile_X6Y14_LUT4AB/W6BEG[0]
+ Tile_X6Y14_LUT4AB/W6BEG[10] Tile_X6Y14_LUT4AB/W6BEG[11] Tile_X6Y14_LUT4AB/W6BEG[1]
+ Tile_X6Y14_LUT4AB/W6BEG[2] Tile_X6Y14_LUT4AB/W6BEG[3] Tile_X6Y14_LUT4AB/W6BEG[4]
+ Tile_X6Y14_LUT4AB/W6BEG[5] Tile_X6Y14_LUT4AB/W6BEG[6] Tile_X6Y14_LUT4AB/W6BEG[7]
+ Tile_X6Y14_LUT4AB/W6BEG[8] Tile_X6Y14_LUT4AB/W6BEG[9] Tile_X5Y14_LUT4AB/WW4BEG[0]
+ Tile_X5Y14_LUT4AB/WW4BEG[10] Tile_X5Y14_LUT4AB/WW4BEG[11] Tile_X5Y14_LUT4AB/WW4BEG[12]
+ Tile_X5Y14_LUT4AB/WW4BEG[13] Tile_X5Y14_LUT4AB/WW4BEG[14] Tile_X5Y14_LUT4AB/WW4BEG[15]
+ Tile_X5Y14_LUT4AB/WW4BEG[1] Tile_X5Y14_LUT4AB/WW4BEG[2] Tile_X5Y14_LUT4AB/WW4BEG[3]
+ Tile_X5Y14_LUT4AB/WW4BEG[4] Tile_X5Y14_LUT4AB/WW4BEG[5] Tile_X5Y14_LUT4AB/WW4BEG[6]
+ Tile_X5Y14_LUT4AB/WW4BEG[7] Tile_X5Y14_LUT4AB/WW4BEG[8] Tile_X5Y14_LUT4AB/WW4BEG[9]
+ Tile_X6Y14_LUT4AB/WW4BEG[0] Tile_X6Y14_LUT4AB/WW4BEG[10] Tile_X6Y14_LUT4AB/WW4BEG[11]
+ Tile_X6Y14_LUT4AB/WW4BEG[12] Tile_X6Y14_LUT4AB/WW4BEG[13] Tile_X6Y14_LUT4AB/WW4BEG[14]
+ Tile_X6Y14_LUT4AB/WW4BEG[15] Tile_X6Y14_LUT4AB/WW4BEG[1] Tile_X6Y14_LUT4AB/WW4BEG[2]
+ Tile_X6Y14_LUT4AB/WW4BEG[3] Tile_X6Y14_LUT4AB/WW4BEG[4] Tile_X6Y14_LUT4AB/WW4BEG[5]
+ Tile_X6Y14_LUT4AB/WW4BEG[6] Tile_X6Y14_LUT4AB/WW4BEG[7] Tile_X6Y14_LUT4AB/WW4BEG[8]
+ Tile_X6Y14_LUT4AB/WW4BEG[9] LUT4AB
XTile_X9Y3_LUT4AB Tile_X9Y4_LUT4AB/Co Tile_X9Y3_LUT4AB/Co Tile_X9Y3_LUT4AB/E1BEG[0]
+ Tile_X9Y3_LUT4AB/E1BEG[1] Tile_X9Y3_LUT4AB/E1BEG[2] Tile_X9Y3_LUT4AB/E1BEG[3] Tile_X9Y3_LUT4AB/E1END[0]
+ Tile_X9Y3_LUT4AB/E1END[1] Tile_X9Y3_LUT4AB/E1END[2] Tile_X9Y3_LUT4AB/E1END[3] Tile_X9Y3_LUT4AB/E2BEG[0]
+ Tile_X9Y3_LUT4AB/E2BEG[1] Tile_X9Y3_LUT4AB/E2BEG[2] Tile_X9Y3_LUT4AB/E2BEG[3] Tile_X9Y3_LUT4AB/E2BEG[4]
+ Tile_X9Y3_LUT4AB/E2BEG[5] Tile_X9Y3_LUT4AB/E2BEG[6] Tile_X9Y3_LUT4AB/E2BEG[7] Tile_X9Y3_LUT4AB/E2BEGb[0]
+ Tile_X9Y3_LUT4AB/E2BEGb[1] Tile_X9Y3_LUT4AB/E2BEGb[2] Tile_X9Y3_LUT4AB/E2BEGb[3]
+ Tile_X9Y3_LUT4AB/E2BEGb[4] Tile_X9Y3_LUT4AB/E2BEGb[5] Tile_X9Y3_LUT4AB/E2BEGb[6]
+ Tile_X9Y3_LUT4AB/E2BEGb[7] Tile_X9Y3_LUT4AB/E2END[0] Tile_X9Y3_LUT4AB/E2END[1] Tile_X9Y3_LUT4AB/E2END[2]
+ Tile_X9Y3_LUT4AB/E2END[3] Tile_X9Y3_LUT4AB/E2END[4] Tile_X9Y3_LUT4AB/E2END[5] Tile_X9Y3_LUT4AB/E2END[6]
+ Tile_X9Y3_LUT4AB/E2END[7] Tile_X9Y3_LUT4AB/E2MID[0] Tile_X9Y3_LUT4AB/E2MID[1] Tile_X9Y3_LUT4AB/E2MID[2]
+ Tile_X9Y3_LUT4AB/E2MID[3] Tile_X9Y3_LUT4AB/E2MID[4] Tile_X9Y3_LUT4AB/E2MID[5] Tile_X9Y3_LUT4AB/E2MID[6]
+ Tile_X9Y3_LUT4AB/E2MID[7] Tile_X9Y3_LUT4AB/E6BEG[0] Tile_X9Y3_LUT4AB/E6BEG[10] Tile_X9Y3_LUT4AB/E6BEG[11]
+ Tile_X9Y3_LUT4AB/E6BEG[1] Tile_X9Y3_LUT4AB/E6BEG[2] Tile_X9Y3_LUT4AB/E6BEG[3] Tile_X9Y3_LUT4AB/E6BEG[4]
+ Tile_X9Y3_LUT4AB/E6BEG[5] Tile_X9Y3_LUT4AB/E6BEG[6] Tile_X9Y3_LUT4AB/E6BEG[7] Tile_X9Y3_LUT4AB/E6BEG[8]
+ Tile_X9Y3_LUT4AB/E6BEG[9] Tile_X9Y3_LUT4AB/E6END[0] Tile_X9Y3_LUT4AB/E6END[10] Tile_X9Y3_LUT4AB/E6END[11]
+ Tile_X9Y3_LUT4AB/E6END[1] Tile_X9Y3_LUT4AB/E6END[2] Tile_X9Y3_LUT4AB/E6END[3] Tile_X9Y3_LUT4AB/E6END[4]
+ Tile_X9Y3_LUT4AB/E6END[5] Tile_X9Y3_LUT4AB/E6END[6] Tile_X9Y3_LUT4AB/E6END[7] Tile_X9Y3_LUT4AB/E6END[8]
+ Tile_X9Y3_LUT4AB/E6END[9] Tile_X9Y3_LUT4AB/EE4BEG[0] Tile_X9Y3_LUT4AB/EE4BEG[10]
+ Tile_X9Y3_LUT4AB/EE4BEG[11] Tile_X9Y3_LUT4AB/EE4BEG[12] Tile_X9Y3_LUT4AB/EE4BEG[13]
+ Tile_X9Y3_LUT4AB/EE4BEG[14] Tile_X9Y3_LUT4AB/EE4BEG[15] Tile_X9Y3_LUT4AB/EE4BEG[1]
+ Tile_X9Y3_LUT4AB/EE4BEG[2] Tile_X9Y3_LUT4AB/EE4BEG[3] Tile_X9Y3_LUT4AB/EE4BEG[4]
+ Tile_X9Y3_LUT4AB/EE4BEG[5] Tile_X9Y3_LUT4AB/EE4BEG[6] Tile_X9Y3_LUT4AB/EE4BEG[7]
+ Tile_X9Y3_LUT4AB/EE4BEG[8] Tile_X9Y3_LUT4AB/EE4BEG[9] Tile_X9Y3_LUT4AB/EE4END[0]
+ Tile_X9Y3_LUT4AB/EE4END[10] Tile_X9Y3_LUT4AB/EE4END[11] Tile_X9Y3_LUT4AB/EE4END[12]
+ Tile_X9Y3_LUT4AB/EE4END[13] Tile_X9Y3_LUT4AB/EE4END[14] Tile_X9Y3_LUT4AB/EE4END[15]
+ Tile_X9Y3_LUT4AB/EE4END[1] Tile_X9Y3_LUT4AB/EE4END[2] Tile_X9Y3_LUT4AB/EE4END[3]
+ Tile_X9Y3_LUT4AB/EE4END[4] Tile_X9Y3_LUT4AB/EE4END[5] Tile_X9Y3_LUT4AB/EE4END[6]
+ Tile_X9Y3_LUT4AB/EE4END[7] Tile_X9Y3_LUT4AB/EE4END[8] Tile_X9Y3_LUT4AB/EE4END[9]
+ Tile_X9Y3_LUT4AB/FrameData[0] Tile_X9Y3_LUT4AB/FrameData[10] Tile_X9Y3_LUT4AB/FrameData[11]
+ Tile_X9Y3_LUT4AB/FrameData[12] Tile_X9Y3_LUT4AB/FrameData[13] Tile_X9Y3_LUT4AB/FrameData[14]
+ Tile_X9Y3_LUT4AB/FrameData[15] Tile_X9Y3_LUT4AB/FrameData[16] Tile_X9Y3_LUT4AB/FrameData[17]
+ Tile_X9Y3_LUT4AB/FrameData[18] Tile_X9Y3_LUT4AB/FrameData[19] Tile_X9Y3_LUT4AB/FrameData[1]
+ Tile_X9Y3_LUT4AB/FrameData[20] Tile_X9Y3_LUT4AB/FrameData[21] Tile_X9Y3_LUT4AB/FrameData[22]
+ Tile_X9Y3_LUT4AB/FrameData[23] Tile_X9Y3_LUT4AB/FrameData[24] Tile_X9Y3_LUT4AB/FrameData[25]
+ Tile_X9Y3_LUT4AB/FrameData[26] Tile_X9Y3_LUT4AB/FrameData[27] Tile_X9Y3_LUT4AB/FrameData[28]
+ Tile_X9Y3_LUT4AB/FrameData[29] Tile_X9Y3_LUT4AB/FrameData[2] Tile_X9Y3_LUT4AB/FrameData[30]
+ Tile_X9Y3_LUT4AB/FrameData[31] Tile_X9Y3_LUT4AB/FrameData[3] Tile_X9Y3_LUT4AB/FrameData[4]
+ Tile_X9Y3_LUT4AB/FrameData[5] Tile_X9Y3_LUT4AB/FrameData[6] Tile_X9Y3_LUT4AB/FrameData[7]
+ Tile_X9Y3_LUT4AB/FrameData[8] Tile_X9Y3_LUT4AB/FrameData[9] Tile_X9Y3_LUT4AB/FrameData_O[0]
+ Tile_X9Y3_LUT4AB/FrameData_O[10] Tile_X9Y3_LUT4AB/FrameData_O[11] Tile_X9Y3_LUT4AB/FrameData_O[12]
+ Tile_X9Y3_LUT4AB/FrameData_O[13] Tile_X9Y3_LUT4AB/FrameData_O[14] Tile_X9Y3_LUT4AB/FrameData_O[15]
+ Tile_X9Y3_LUT4AB/FrameData_O[16] Tile_X9Y3_LUT4AB/FrameData_O[17] Tile_X9Y3_LUT4AB/FrameData_O[18]
+ Tile_X9Y3_LUT4AB/FrameData_O[19] Tile_X9Y3_LUT4AB/FrameData_O[1] Tile_X9Y3_LUT4AB/FrameData_O[20]
+ Tile_X9Y3_LUT4AB/FrameData_O[21] Tile_X9Y3_LUT4AB/FrameData_O[22] Tile_X9Y3_LUT4AB/FrameData_O[23]
+ Tile_X9Y3_LUT4AB/FrameData_O[24] Tile_X9Y3_LUT4AB/FrameData_O[25] Tile_X9Y3_LUT4AB/FrameData_O[26]
+ Tile_X9Y3_LUT4AB/FrameData_O[27] Tile_X9Y3_LUT4AB/FrameData_O[28] Tile_X9Y3_LUT4AB/FrameData_O[29]
+ Tile_X9Y3_LUT4AB/FrameData_O[2] Tile_X9Y3_LUT4AB/FrameData_O[30] Tile_X9Y3_LUT4AB/FrameData_O[31]
+ Tile_X9Y3_LUT4AB/FrameData_O[3] Tile_X9Y3_LUT4AB/FrameData_O[4] Tile_X9Y3_LUT4AB/FrameData_O[5]
+ Tile_X9Y3_LUT4AB/FrameData_O[6] Tile_X9Y3_LUT4AB/FrameData_O[7] Tile_X9Y3_LUT4AB/FrameData_O[8]
+ Tile_X9Y3_LUT4AB/FrameData_O[9] Tile_X9Y3_LUT4AB/FrameStrobe[0] Tile_X9Y3_LUT4AB/FrameStrobe[10]
+ Tile_X9Y3_LUT4AB/FrameStrobe[11] Tile_X9Y3_LUT4AB/FrameStrobe[12] Tile_X9Y3_LUT4AB/FrameStrobe[13]
+ Tile_X9Y3_LUT4AB/FrameStrobe[14] Tile_X9Y3_LUT4AB/FrameStrobe[15] Tile_X9Y3_LUT4AB/FrameStrobe[16]
+ Tile_X9Y3_LUT4AB/FrameStrobe[17] Tile_X9Y3_LUT4AB/FrameStrobe[18] Tile_X9Y3_LUT4AB/FrameStrobe[19]
+ Tile_X9Y3_LUT4AB/FrameStrobe[1] Tile_X9Y3_LUT4AB/FrameStrobe[2] Tile_X9Y3_LUT4AB/FrameStrobe[3]
+ Tile_X9Y3_LUT4AB/FrameStrobe[4] Tile_X9Y3_LUT4AB/FrameStrobe[5] Tile_X9Y3_LUT4AB/FrameStrobe[6]
+ Tile_X9Y3_LUT4AB/FrameStrobe[7] Tile_X9Y3_LUT4AB/FrameStrobe[8] Tile_X9Y3_LUT4AB/FrameStrobe[9]
+ Tile_X9Y2_LUT4AB/FrameStrobe[0] Tile_X9Y2_LUT4AB/FrameStrobe[10] Tile_X9Y2_LUT4AB/FrameStrobe[11]
+ Tile_X9Y2_LUT4AB/FrameStrobe[12] Tile_X9Y2_LUT4AB/FrameStrobe[13] Tile_X9Y2_LUT4AB/FrameStrobe[14]
+ Tile_X9Y2_LUT4AB/FrameStrobe[15] Tile_X9Y2_LUT4AB/FrameStrobe[16] Tile_X9Y2_LUT4AB/FrameStrobe[17]
+ Tile_X9Y2_LUT4AB/FrameStrobe[18] Tile_X9Y2_LUT4AB/FrameStrobe[19] Tile_X9Y2_LUT4AB/FrameStrobe[1]
+ Tile_X9Y2_LUT4AB/FrameStrobe[2] Tile_X9Y2_LUT4AB/FrameStrobe[3] Tile_X9Y2_LUT4AB/FrameStrobe[4]
+ Tile_X9Y2_LUT4AB/FrameStrobe[5] Tile_X9Y2_LUT4AB/FrameStrobe[6] Tile_X9Y2_LUT4AB/FrameStrobe[7]
+ Tile_X9Y2_LUT4AB/FrameStrobe[8] Tile_X9Y2_LUT4AB/FrameStrobe[9] Tile_X9Y3_LUT4AB/N1BEG[0]
+ Tile_X9Y3_LUT4AB/N1BEG[1] Tile_X9Y3_LUT4AB/N1BEG[2] Tile_X9Y3_LUT4AB/N1BEG[3] Tile_X9Y4_LUT4AB/N1BEG[0]
+ Tile_X9Y4_LUT4AB/N1BEG[1] Tile_X9Y4_LUT4AB/N1BEG[2] Tile_X9Y4_LUT4AB/N1BEG[3] Tile_X9Y3_LUT4AB/N2BEG[0]
+ Tile_X9Y3_LUT4AB/N2BEG[1] Tile_X9Y3_LUT4AB/N2BEG[2] Tile_X9Y3_LUT4AB/N2BEG[3] Tile_X9Y3_LUT4AB/N2BEG[4]
+ Tile_X9Y3_LUT4AB/N2BEG[5] Tile_X9Y3_LUT4AB/N2BEG[6] Tile_X9Y3_LUT4AB/N2BEG[7] Tile_X9Y2_LUT4AB/N2END[0]
+ Tile_X9Y2_LUT4AB/N2END[1] Tile_X9Y2_LUT4AB/N2END[2] Tile_X9Y2_LUT4AB/N2END[3] Tile_X9Y2_LUT4AB/N2END[4]
+ Tile_X9Y2_LUT4AB/N2END[5] Tile_X9Y2_LUT4AB/N2END[6] Tile_X9Y2_LUT4AB/N2END[7] Tile_X9Y3_LUT4AB/N2END[0]
+ Tile_X9Y3_LUT4AB/N2END[1] Tile_X9Y3_LUT4AB/N2END[2] Tile_X9Y3_LUT4AB/N2END[3] Tile_X9Y3_LUT4AB/N2END[4]
+ Tile_X9Y3_LUT4AB/N2END[5] Tile_X9Y3_LUT4AB/N2END[6] Tile_X9Y3_LUT4AB/N2END[7] Tile_X9Y4_LUT4AB/N2BEG[0]
+ Tile_X9Y4_LUT4AB/N2BEG[1] Tile_X9Y4_LUT4AB/N2BEG[2] Tile_X9Y4_LUT4AB/N2BEG[3] Tile_X9Y4_LUT4AB/N2BEG[4]
+ Tile_X9Y4_LUT4AB/N2BEG[5] Tile_X9Y4_LUT4AB/N2BEG[6] Tile_X9Y4_LUT4AB/N2BEG[7] Tile_X9Y3_LUT4AB/N4BEG[0]
+ Tile_X9Y3_LUT4AB/N4BEG[10] Tile_X9Y3_LUT4AB/N4BEG[11] Tile_X9Y3_LUT4AB/N4BEG[12]
+ Tile_X9Y3_LUT4AB/N4BEG[13] Tile_X9Y3_LUT4AB/N4BEG[14] Tile_X9Y3_LUT4AB/N4BEG[15]
+ Tile_X9Y3_LUT4AB/N4BEG[1] Tile_X9Y3_LUT4AB/N4BEG[2] Tile_X9Y3_LUT4AB/N4BEG[3] Tile_X9Y3_LUT4AB/N4BEG[4]
+ Tile_X9Y3_LUT4AB/N4BEG[5] Tile_X9Y3_LUT4AB/N4BEG[6] Tile_X9Y3_LUT4AB/N4BEG[7] Tile_X9Y3_LUT4AB/N4BEG[8]
+ Tile_X9Y3_LUT4AB/N4BEG[9] Tile_X9Y4_LUT4AB/N4BEG[0] Tile_X9Y4_LUT4AB/N4BEG[10] Tile_X9Y4_LUT4AB/N4BEG[11]
+ Tile_X9Y4_LUT4AB/N4BEG[12] Tile_X9Y4_LUT4AB/N4BEG[13] Tile_X9Y4_LUT4AB/N4BEG[14]
+ Tile_X9Y4_LUT4AB/N4BEG[15] Tile_X9Y4_LUT4AB/N4BEG[1] Tile_X9Y4_LUT4AB/N4BEG[2] Tile_X9Y4_LUT4AB/N4BEG[3]
+ Tile_X9Y4_LUT4AB/N4BEG[4] Tile_X9Y4_LUT4AB/N4BEG[5] Tile_X9Y4_LUT4AB/N4BEG[6] Tile_X9Y4_LUT4AB/N4BEG[7]
+ Tile_X9Y4_LUT4AB/N4BEG[8] Tile_X9Y4_LUT4AB/N4BEG[9] Tile_X9Y3_LUT4AB/NN4BEG[0] Tile_X9Y3_LUT4AB/NN4BEG[10]
+ Tile_X9Y3_LUT4AB/NN4BEG[11] Tile_X9Y3_LUT4AB/NN4BEG[12] Tile_X9Y3_LUT4AB/NN4BEG[13]
+ Tile_X9Y3_LUT4AB/NN4BEG[14] Tile_X9Y3_LUT4AB/NN4BEG[15] Tile_X9Y3_LUT4AB/NN4BEG[1]
+ Tile_X9Y3_LUT4AB/NN4BEG[2] Tile_X9Y3_LUT4AB/NN4BEG[3] Tile_X9Y3_LUT4AB/NN4BEG[4]
+ Tile_X9Y3_LUT4AB/NN4BEG[5] Tile_X9Y3_LUT4AB/NN4BEG[6] Tile_X9Y3_LUT4AB/NN4BEG[7]
+ Tile_X9Y3_LUT4AB/NN4BEG[8] Tile_X9Y3_LUT4AB/NN4BEG[9] Tile_X9Y4_LUT4AB/NN4BEG[0]
+ Tile_X9Y4_LUT4AB/NN4BEG[10] Tile_X9Y4_LUT4AB/NN4BEG[11] Tile_X9Y4_LUT4AB/NN4BEG[12]
+ Tile_X9Y4_LUT4AB/NN4BEG[13] Tile_X9Y4_LUT4AB/NN4BEG[14] Tile_X9Y4_LUT4AB/NN4BEG[15]
+ Tile_X9Y4_LUT4AB/NN4BEG[1] Tile_X9Y4_LUT4AB/NN4BEG[2] Tile_X9Y4_LUT4AB/NN4BEG[3]
+ Tile_X9Y4_LUT4AB/NN4BEG[4] Tile_X9Y4_LUT4AB/NN4BEG[5] Tile_X9Y4_LUT4AB/NN4BEG[6]
+ Tile_X9Y4_LUT4AB/NN4BEG[7] Tile_X9Y4_LUT4AB/NN4BEG[8] Tile_X9Y4_LUT4AB/NN4BEG[9]
+ Tile_X9Y4_LUT4AB/S1END[0] Tile_X9Y4_LUT4AB/S1END[1] Tile_X9Y4_LUT4AB/S1END[2] Tile_X9Y4_LUT4AB/S1END[3]
+ Tile_X9Y3_LUT4AB/S1END[0] Tile_X9Y3_LUT4AB/S1END[1] Tile_X9Y3_LUT4AB/S1END[2] Tile_X9Y3_LUT4AB/S1END[3]
+ Tile_X9Y4_LUT4AB/S2MID[0] Tile_X9Y4_LUT4AB/S2MID[1] Tile_X9Y4_LUT4AB/S2MID[2] Tile_X9Y4_LUT4AB/S2MID[3]
+ Tile_X9Y4_LUT4AB/S2MID[4] Tile_X9Y4_LUT4AB/S2MID[5] Tile_X9Y4_LUT4AB/S2MID[6] Tile_X9Y4_LUT4AB/S2MID[7]
+ Tile_X9Y4_LUT4AB/S2END[0] Tile_X9Y4_LUT4AB/S2END[1] Tile_X9Y4_LUT4AB/S2END[2] Tile_X9Y4_LUT4AB/S2END[3]
+ Tile_X9Y4_LUT4AB/S2END[4] Tile_X9Y4_LUT4AB/S2END[5] Tile_X9Y4_LUT4AB/S2END[6] Tile_X9Y4_LUT4AB/S2END[7]
+ Tile_X9Y3_LUT4AB/S2END[0] Tile_X9Y3_LUT4AB/S2END[1] Tile_X9Y3_LUT4AB/S2END[2] Tile_X9Y3_LUT4AB/S2END[3]
+ Tile_X9Y3_LUT4AB/S2END[4] Tile_X9Y3_LUT4AB/S2END[5] Tile_X9Y3_LUT4AB/S2END[6] Tile_X9Y3_LUT4AB/S2END[7]
+ Tile_X9Y3_LUT4AB/S2MID[0] Tile_X9Y3_LUT4AB/S2MID[1] Tile_X9Y3_LUT4AB/S2MID[2] Tile_X9Y3_LUT4AB/S2MID[3]
+ Tile_X9Y3_LUT4AB/S2MID[4] Tile_X9Y3_LUT4AB/S2MID[5] Tile_X9Y3_LUT4AB/S2MID[6] Tile_X9Y3_LUT4AB/S2MID[7]
+ Tile_X9Y4_LUT4AB/S4END[0] Tile_X9Y4_LUT4AB/S4END[10] Tile_X9Y4_LUT4AB/S4END[11]
+ Tile_X9Y4_LUT4AB/S4END[12] Tile_X9Y4_LUT4AB/S4END[13] Tile_X9Y4_LUT4AB/S4END[14]
+ Tile_X9Y4_LUT4AB/S4END[15] Tile_X9Y4_LUT4AB/S4END[1] Tile_X9Y4_LUT4AB/S4END[2] Tile_X9Y4_LUT4AB/S4END[3]
+ Tile_X9Y4_LUT4AB/S4END[4] Tile_X9Y4_LUT4AB/S4END[5] Tile_X9Y4_LUT4AB/S4END[6] Tile_X9Y4_LUT4AB/S4END[7]
+ Tile_X9Y4_LUT4AB/S4END[8] Tile_X9Y4_LUT4AB/S4END[9] Tile_X9Y3_LUT4AB/S4END[0] Tile_X9Y3_LUT4AB/S4END[10]
+ Tile_X9Y3_LUT4AB/S4END[11] Tile_X9Y3_LUT4AB/S4END[12] Tile_X9Y3_LUT4AB/S4END[13]
+ Tile_X9Y3_LUT4AB/S4END[14] Tile_X9Y3_LUT4AB/S4END[15] Tile_X9Y3_LUT4AB/S4END[1]
+ Tile_X9Y3_LUT4AB/S4END[2] Tile_X9Y3_LUT4AB/S4END[3] Tile_X9Y3_LUT4AB/S4END[4] Tile_X9Y3_LUT4AB/S4END[5]
+ Tile_X9Y3_LUT4AB/S4END[6] Tile_X9Y3_LUT4AB/S4END[7] Tile_X9Y3_LUT4AB/S4END[8] Tile_X9Y3_LUT4AB/S4END[9]
+ Tile_X9Y4_LUT4AB/SS4END[0] Tile_X9Y4_LUT4AB/SS4END[10] Tile_X9Y4_LUT4AB/SS4END[11]
+ Tile_X9Y4_LUT4AB/SS4END[12] Tile_X9Y4_LUT4AB/SS4END[13] Tile_X9Y4_LUT4AB/SS4END[14]
+ Tile_X9Y4_LUT4AB/SS4END[15] Tile_X9Y4_LUT4AB/SS4END[1] Tile_X9Y4_LUT4AB/SS4END[2]
+ Tile_X9Y4_LUT4AB/SS4END[3] Tile_X9Y4_LUT4AB/SS4END[4] Tile_X9Y4_LUT4AB/SS4END[5]
+ Tile_X9Y4_LUT4AB/SS4END[6] Tile_X9Y4_LUT4AB/SS4END[7] Tile_X9Y4_LUT4AB/SS4END[8]
+ Tile_X9Y4_LUT4AB/SS4END[9] Tile_X9Y3_LUT4AB/SS4END[0] Tile_X9Y3_LUT4AB/SS4END[10]
+ Tile_X9Y3_LUT4AB/SS4END[11] Tile_X9Y3_LUT4AB/SS4END[12] Tile_X9Y3_LUT4AB/SS4END[13]
+ Tile_X9Y3_LUT4AB/SS4END[14] Tile_X9Y3_LUT4AB/SS4END[15] Tile_X9Y3_LUT4AB/SS4END[1]
+ Tile_X9Y3_LUT4AB/SS4END[2] Tile_X9Y3_LUT4AB/SS4END[3] Tile_X9Y3_LUT4AB/SS4END[4]
+ Tile_X9Y3_LUT4AB/SS4END[5] Tile_X9Y3_LUT4AB/SS4END[6] Tile_X9Y3_LUT4AB/SS4END[7]
+ Tile_X9Y3_LUT4AB/SS4END[8] Tile_X9Y3_LUT4AB/SS4END[9] Tile_X9Y3_LUT4AB/UserCLK Tile_X9Y2_LUT4AB/UserCLK
+ VGND VPWR Tile_X9Y3_LUT4AB/W1BEG[0] Tile_X9Y3_LUT4AB/W1BEG[1] Tile_X9Y3_LUT4AB/W1BEG[2]
+ Tile_X9Y3_LUT4AB/W1BEG[3] Tile_X9Y3_LUT4AB/W1END[0] Tile_X9Y3_LUT4AB/W1END[1] Tile_X9Y3_LUT4AB/W1END[2]
+ Tile_X9Y3_LUT4AB/W1END[3] Tile_X9Y3_LUT4AB/W2BEG[0] Tile_X9Y3_LUT4AB/W2BEG[1] Tile_X9Y3_LUT4AB/W2BEG[2]
+ Tile_X9Y3_LUT4AB/W2BEG[3] Tile_X9Y3_LUT4AB/W2BEG[4] Tile_X9Y3_LUT4AB/W2BEG[5] Tile_X9Y3_LUT4AB/W2BEG[6]
+ Tile_X9Y3_LUT4AB/W2BEG[7] Tile_X8Y3_LUT4AB/W2END[0] Tile_X8Y3_LUT4AB/W2END[1] Tile_X8Y3_LUT4AB/W2END[2]
+ Tile_X8Y3_LUT4AB/W2END[3] Tile_X8Y3_LUT4AB/W2END[4] Tile_X8Y3_LUT4AB/W2END[5] Tile_X8Y3_LUT4AB/W2END[6]
+ Tile_X8Y3_LUT4AB/W2END[7] Tile_X9Y3_LUT4AB/W2END[0] Tile_X9Y3_LUT4AB/W2END[1] Tile_X9Y3_LUT4AB/W2END[2]
+ Tile_X9Y3_LUT4AB/W2END[3] Tile_X9Y3_LUT4AB/W2END[4] Tile_X9Y3_LUT4AB/W2END[5] Tile_X9Y3_LUT4AB/W2END[6]
+ Tile_X9Y3_LUT4AB/W2END[7] Tile_X9Y3_LUT4AB/W2MID[0] Tile_X9Y3_LUT4AB/W2MID[1] Tile_X9Y3_LUT4AB/W2MID[2]
+ Tile_X9Y3_LUT4AB/W2MID[3] Tile_X9Y3_LUT4AB/W2MID[4] Tile_X9Y3_LUT4AB/W2MID[5] Tile_X9Y3_LUT4AB/W2MID[6]
+ Tile_X9Y3_LUT4AB/W2MID[7] Tile_X9Y3_LUT4AB/W6BEG[0] Tile_X9Y3_LUT4AB/W6BEG[10] Tile_X9Y3_LUT4AB/W6BEG[11]
+ Tile_X9Y3_LUT4AB/W6BEG[1] Tile_X9Y3_LUT4AB/W6BEG[2] Tile_X9Y3_LUT4AB/W6BEG[3] Tile_X9Y3_LUT4AB/W6BEG[4]
+ Tile_X9Y3_LUT4AB/W6BEG[5] Tile_X9Y3_LUT4AB/W6BEG[6] Tile_X9Y3_LUT4AB/W6BEG[7] Tile_X9Y3_LUT4AB/W6BEG[8]
+ Tile_X9Y3_LUT4AB/W6BEG[9] Tile_X9Y3_LUT4AB/W6END[0] Tile_X9Y3_LUT4AB/W6END[10] Tile_X9Y3_LUT4AB/W6END[11]
+ Tile_X9Y3_LUT4AB/W6END[1] Tile_X9Y3_LUT4AB/W6END[2] Tile_X9Y3_LUT4AB/W6END[3] Tile_X9Y3_LUT4AB/W6END[4]
+ Tile_X9Y3_LUT4AB/W6END[5] Tile_X9Y3_LUT4AB/W6END[6] Tile_X9Y3_LUT4AB/W6END[7] Tile_X9Y3_LUT4AB/W6END[8]
+ Tile_X9Y3_LUT4AB/W6END[9] Tile_X9Y3_LUT4AB/WW4BEG[0] Tile_X9Y3_LUT4AB/WW4BEG[10]
+ Tile_X9Y3_LUT4AB/WW4BEG[11] Tile_X9Y3_LUT4AB/WW4BEG[12] Tile_X9Y3_LUT4AB/WW4BEG[13]
+ Tile_X9Y3_LUT4AB/WW4BEG[14] Tile_X9Y3_LUT4AB/WW4BEG[15] Tile_X9Y3_LUT4AB/WW4BEG[1]
+ Tile_X9Y3_LUT4AB/WW4BEG[2] Tile_X9Y3_LUT4AB/WW4BEG[3] Tile_X9Y3_LUT4AB/WW4BEG[4]
+ Tile_X9Y3_LUT4AB/WW4BEG[5] Tile_X9Y3_LUT4AB/WW4BEG[6] Tile_X9Y3_LUT4AB/WW4BEG[7]
+ Tile_X9Y3_LUT4AB/WW4BEG[8] Tile_X9Y3_LUT4AB/WW4BEG[9] Tile_X9Y3_LUT4AB/WW4END[0]
+ Tile_X9Y3_LUT4AB/WW4END[10] Tile_X9Y3_LUT4AB/WW4END[11] Tile_X9Y3_LUT4AB/WW4END[12]
+ Tile_X9Y3_LUT4AB/WW4END[13] Tile_X9Y3_LUT4AB/WW4END[14] Tile_X9Y3_LUT4AB/WW4END[15]
+ Tile_X9Y3_LUT4AB/WW4END[1] Tile_X9Y3_LUT4AB/WW4END[2] Tile_X9Y3_LUT4AB/WW4END[3]
+ Tile_X9Y3_LUT4AB/WW4END[4] Tile_X9Y3_LUT4AB/WW4END[5] Tile_X9Y3_LUT4AB/WW4END[6]
+ Tile_X9Y3_LUT4AB/WW4END[7] Tile_X9Y3_LUT4AB/WW4END[8] Tile_X9Y3_LUT4AB/WW4END[9]
+ LUT4AB
XTile_X0Y10_W_IO Tile_X0Y10_A_I_top Tile_X0Y10_A_O_top Tile_X0Y10_A_T_top Tile_X0Y10_A_config_C_bit0
+ Tile_X0Y10_A_config_C_bit1 Tile_X0Y10_A_config_C_bit2 Tile_X0Y10_A_config_C_bit3
+ Tile_X0Y10_B_I_top Tile_X0Y10_B_O_top Tile_X0Y10_B_T_top Tile_X0Y10_B_config_C_bit0
+ Tile_X0Y10_B_config_C_bit1 Tile_X0Y10_B_config_C_bit2 Tile_X0Y10_B_config_C_bit3
+ Tile_X0Y10_W_IO/E1BEG[0] Tile_X0Y10_W_IO/E1BEG[1] Tile_X0Y10_W_IO/E1BEG[2] Tile_X0Y10_W_IO/E1BEG[3]
+ Tile_X0Y10_W_IO/E2BEG[0] Tile_X0Y10_W_IO/E2BEG[1] Tile_X0Y10_W_IO/E2BEG[2] Tile_X0Y10_W_IO/E2BEG[3]
+ Tile_X0Y10_W_IO/E2BEG[4] Tile_X0Y10_W_IO/E2BEG[5] Tile_X0Y10_W_IO/E2BEG[6] Tile_X0Y10_W_IO/E2BEG[7]
+ Tile_X0Y10_W_IO/E2BEGb[0] Tile_X0Y10_W_IO/E2BEGb[1] Tile_X0Y10_W_IO/E2BEGb[2] Tile_X0Y10_W_IO/E2BEGb[3]
+ Tile_X0Y10_W_IO/E2BEGb[4] Tile_X0Y10_W_IO/E2BEGb[5] Tile_X0Y10_W_IO/E2BEGb[6] Tile_X0Y10_W_IO/E2BEGb[7]
+ Tile_X0Y10_W_IO/E6BEG[0] Tile_X0Y10_W_IO/E6BEG[10] Tile_X0Y10_W_IO/E6BEG[11] Tile_X0Y10_W_IO/E6BEG[1]
+ Tile_X0Y10_W_IO/E6BEG[2] Tile_X0Y10_W_IO/E6BEG[3] Tile_X0Y10_W_IO/E6BEG[4] Tile_X0Y10_W_IO/E6BEG[5]
+ Tile_X0Y10_W_IO/E6BEG[6] Tile_X0Y10_W_IO/E6BEG[7] Tile_X0Y10_W_IO/E6BEG[8] Tile_X0Y10_W_IO/E6BEG[9]
+ Tile_X0Y10_W_IO/EE4BEG[0] Tile_X0Y10_W_IO/EE4BEG[10] Tile_X0Y10_W_IO/EE4BEG[11]
+ Tile_X0Y10_W_IO/EE4BEG[12] Tile_X0Y10_W_IO/EE4BEG[13] Tile_X0Y10_W_IO/EE4BEG[14]
+ Tile_X0Y10_W_IO/EE4BEG[15] Tile_X0Y10_W_IO/EE4BEG[1] Tile_X0Y10_W_IO/EE4BEG[2] Tile_X0Y10_W_IO/EE4BEG[3]
+ Tile_X0Y10_W_IO/EE4BEG[4] Tile_X0Y10_W_IO/EE4BEG[5] Tile_X0Y10_W_IO/EE4BEG[6] Tile_X0Y10_W_IO/EE4BEG[7]
+ Tile_X0Y10_W_IO/EE4BEG[8] Tile_X0Y10_W_IO/EE4BEG[9] FrameData[320] FrameData[330]
+ FrameData[331] FrameData[332] FrameData[333] FrameData[334] FrameData[335] FrameData[336]
+ FrameData[337] FrameData[338] FrameData[339] FrameData[321] FrameData[340] FrameData[341]
+ FrameData[342] FrameData[343] FrameData[344] FrameData[345] FrameData[346] FrameData[347]
+ FrameData[348] FrameData[349] FrameData[322] FrameData[350] FrameData[351] FrameData[323]
+ FrameData[324] FrameData[325] FrameData[326] FrameData[327] FrameData[328] FrameData[329]
+ Tile_X1Y10_LUT4AB/FrameData[0] Tile_X1Y10_LUT4AB/FrameData[10] Tile_X1Y10_LUT4AB/FrameData[11]
+ Tile_X1Y10_LUT4AB/FrameData[12] Tile_X1Y10_LUT4AB/FrameData[13] Tile_X1Y10_LUT4AB/FrameData[14]
+ Tile_X1Y10_LUT4AB/FrameData[15] Tile_X1Y10_LUT4AB/FrameData[16] Tile_X1Y10_LUT4AB/FrameData[17]
+ Tile_X1Y10_LUT4AB/FrameData[18] Tile_X1Y10_LUT4AB/FrameData[19] Tile_X1Y10_LUT4AB/FrameData[1]
+ Tile_X1Y10_LUT4AB/FrameData[20] Tile_X1Y10_LUT4AB/FrameData[21] Tile_X1Y10_LUT4AB/FrameData[22]
+ Tile_X1Y10_LUT4AB/FrameData[23] Tile_X1Y10_LUT4AB/FrameData[24] Tile_X1Y10_LUT4AB/FrameData[25]
+ Tile_X1Y10_LUT4AB/FrameData[26] Tile_X1Y10_LUT4AB/FrameData[27] Tile_X1Y10_LUT4AB/FrameData[28]
+ Tile_X1Y10_LUT4AB/FrameData[29] Tile_X1Y10_LUT4AB/FrameData[2] Tile_X1Y10_LUT4AB/FrameData[30]
+ Tile_X1Y10_LUT4AB/FrameData[31] Tile_X1Y10_LUT4AB/FrameData[3] Tile_X1Y10_LUT4AB/FrameData[4]
+ Tile_X1Y10_LUT4AB/FrameData[5] Tile_X1Y10_LUT4AB/FrameData[6] Tile_X1Y10_LUT4AB/FrameData[7]
+ Tile_X1Y10_LUT4AB/FrameData[8] Tile_X1Y10_LUT4AB/FrameData[9] Tile_X0Y10_W_IO/FrameStrobe[0]
+ Tile_X0Y10_W_IO/FrameStrobe[10] Tile_X0Y10_W_IO/FrameStrobe[11] Tile_X0Y10_W_IO/FrameStrobe[12]
+ Tile_X0Y10_W_IO/FrameStrobe[13] Tile_X0Y10_W_IO/FrameStrobe[14] Tile_X0Y10_W_IO/FrameStrobe[15]
+ Tile_X0Y10_W_IO/FrameStrobe[16] Tile_X0Y10_W_IO/FrameStrobe[17] Tile_X0Y10_W_IO/FrameStrobe[18]
+ Tile_X0Y10_W_IO/FrameStrobe[19] Tile_X0Y10_W_IO/FrameStrobe[1] Tile_X0Y10_W_IO/FrameStrobe[2]
+ Tile_X0Y10_W_IO/FrameStrobe[3] Tile_X0Y10_W_IO/FrameStrobe[4] Tile_X0Y10_W_IO/FrameStrobe[5]
+ Tile_X0Y10_W_IO/FrameStrobe[6] Tile_X0Y10_W_IO/FrameStrobe[7] Tile_X0Y10_W_IO/FrameStrobe[8]
+ Tile_X0Y10_W_IO/FrameStrobe[9] Tile_X0Y9_W_IO/FrameStrobe[0] Tile_X0Y9_W_IO/FrameStrobe[10]
+ Tile_X0Y9_W_IO/FrameStrobe[11] Tile_X0Y9_W_IO/FrameStrobe[12] Tile_X0Y9_W_IO/FrameStrobe[13]
+ Tile_X0Y9_W_IO/FrameStrobe[14] Tile_X0Y9_W_IO/FrameStrobe[15] Tile_X0Y9_W_IO/FrameStrobe[16]
+ Tile_X0Y9_W_IO/FrameStrobe[17] Tile_X0Y9_W_IO/FrameStrobe[18] Tile_X0Y9_W_IO/FrameStrobe[19]
+ Tile_X0Y9_W_IO/FrameStrobe[1] Tile_X0Y9_W_IO/FrameStrobe[2] Tile_X0Y9_W_IO/FrameStrobe[3]
+ Tile_X0Y9_W_IO/FrameStrobe[4] Tile_X0Y9_W_IO/FrameStrobe[5] Tile_X0Y9_W_IO/FrameStrobe[6]
+ Tile_X0Y9_W_IO/FrameStrobe[7] Tile_X0Y9_W_IO/FrameStrobe[8] Tile_X0Y9_W_IO/FrameStrobe[9]
+ Tile_X0Y10_W_IO/UserCLK Tile_X0Y9_W_IO/UserCLK VGND VPWR Tile_X0Y10_W_IO/W1END[0]
+ Tile_X0Y10_W_IO/W1END[1] Tile_X0Y10_W_IO/W1END[2] Tile_X0Y10_W_IO/W1END[3] Tile_X0Y10_W_IO/W2END[0]
+ Tile_X0Y10_W_IO/W2END[1] Tile_X0Y10_W_IO/W2END[2] Tile_X0Y10_W_IO/W2END[3] Tile_X0Y10_W_IO/W2END[4]
+ Tile_X0Y10_W_IO/W2END[5] Tile_X0Y10_W_IO/W2END[6] Tile_X0Y10_W_IO/W2END[7] Tile_X0Y10_W_IO/W2MID[0]
+ Tile_X0Y10_W_IO/W2MID[1] Tile_X0Y10_W_IO/W2MID[2] Tile_X0Y10_W_IO/W2MID[3] Tile_X0Y10_W_IO/W2MID[4]
+ Tile_X0Y10_W_IO/W2MID[5] Tile_X0Y10_W_IO/W2MID[6] Tile_X0Y10_W_IO/W2MID[7] Tile_X0Y10_W_IO/W6END[0]
+ Tile_X0Y10_W_IO/W6END[10] Tile_X0Y10_W_IO/W6END[11] Tile_X0Y10_W_IO/W6END[1] Tile_X0Y10_W_IO/W6END[2]
+ Tile_X0Y10_W_IO/W6END[3] Tile_X0Y10_W_IO/W6END[4] Tile_X0Y10_W_IO/W6END[5] Tile_X0Y10_W_IO/W6END[6]
+ Tile_X0Y10_W_IO/W6END[7] Tile_X0Y10_W_IO/W6END[8] Tile_X0Y10_W_IO/W6END[9] Tile_X0Y10_W_IO/WW4END[0]
+ Tile_X0Y10_W_IO/WW4END[10] Tile_X0Y10_W_IO/WW4END[11] Tile_X0Y10_W_IO/WW4END[12]
+ Tile_X0Y10_W_IO/WW4END[13] Tile_X0Y10_W_IO/WW4END[14] Tile_X0Y10_W_IO/WW4END[15]
+ Tile_X0Y10_W_IO/WW4END[1] Tile_X0Y10_W_IO/WW4END[2] Tile_X0Y10_W_IO/WW4END[3] Tile_X0Y10_W_IO/WW4END[4]
+ Tile_X0Y10_W_IO/WW4END[5] Tile_X0Y10_W_IO/WW4END[6] Tile_X0Y10_W_IO/WW4END[7] Tile_X0Y10_W_IO/WW4END[8]
+ Tile_X0Y10_W_IO/WW4END[9] W_IO
XTile_X7Y1_DSP Tile_X8Y1_LUT4AB/E1END[0] Tile_X8Y1_LUT4AB/E1END[1] Tile_X8Y1_LUT4AB/E1END[2]
+ Tile_X8Y1_LUT4AB/E1END[3] Tile_X6Y1_LUT4AB/E1BEG[0] Tile_X6Y1_LUT4AB/E1BEG[1] Tile_X6Y1_LUT4AB/E1BEG[2]
+ Tile_X6Y1_LUT4AB/E1BEG[3] Tile_X8Y1_LUT4AB/E2MID[0] Tile_X8Y1_LUT4AB/E2MID[1] Tile_X8Y1_LUT4AB/E2MID[2]
+ Tile_X8Y1_LUT4AB/E2MID[3] Tile_X8Y1_LUT4AB/E2MID[4] Tile_X8Y1_LUT4AB/E2MID[5] Tile_X8Y1_LUT4AB/E2MID[6]
+ Tile_X8Y1_LUT4AB/E2MID[7] Tile_X8Y1_LUT4AB/E2END[0] Tile_X8Y1_LUT4AB/E2END[1] Tile_X8Y1_LUT4AB/E2END[2]
+ Tile_X8Y1_LUT4AB/E2END[3] Tile_X8Y1_LUT4AB/E2END[4] Tile_X8Y1_LUT4AB/E2END[5] Tile_X8Y1_LUT4AB/E2END[6]
+ Tile_X8Y1_LUT4AB/E2END[7] Tile_X6Y1_LUT4AB/E2BEGb[0] Tile_X6Y1_LUT4AB/E2BEGb[1]
+ Tile_X6Y1_LUT4AB/E2BEGb[2] Tile_X6Y1_LUT4AB/E2BEGb[3] Tile_X6Y1_LUT4AB/E2BEGb[4]
+ Tile_X6Y1_LUT4AB/E2BEGb[5] Tile_X6Y1_LUT4AB/E2BEGb[6] Tile_X6Y1_LUT4AB/E2BEGb[7]
+ Tile_X6Y1_LUT4AB/E2BEG[0] Tile_X6Y1_LUT4AB/E2BEG[1] Tile_X6Y1_LUT4AB/E2BEG[2] Tile_X6Y1_LUT4AB/E2BEG[3]
+ Tile_X6Y1_LUT4AB/E2BEG[4] Tile_X6Y1_LUT4AB/E2BEG[5] Tile_X6Y1_LUT4AB/E2BEG[6] Tile_X6Y1_LUT4AB/E2BEG[7]
+ Tile_X8Y1_LUT4AB/E6END[0] Tile_X8Y1_LUT4AB/E6END[10] Tile_X8Y1_LUT4AB/E6END[11]
+ Tile_X8Y1_LUT4AB/E6END[1] Tile_X8Y1_LUT4AB/E6END[2] Tile_X8Y1_LUT4AB/E6END[3] Tile_X8Y1_LUT4AB/E6END[4]
+ Tile_X8Y1_LUT4AB/E6END[5] Tile_X8Y1_LUT4AB/E6END[6] Tile_X8Y1_LUT4AB/E6END[7] Tile_X8Y1_LUT4AB/E6END[8]
+ Tile_X8Y1_LUT4AB/E6END[9] Tile_X6Y1_LUT4AB/E6BEG[0] Tile_X6Y1_LUT4AB/E6BEG[10] Tile_X6Y1_LUT4AB/E6BEG[11]
+ Tile_X6Y1_LUT4AB/E6BEG[1] Tile_X6Y1_LUT4AB/E6BEG[2] Tile_X6Y1_LUT4AB/E6BEG[3] Tile_X6Y1_LUT4AB/E6BEG[4]
+ Tile_X6Y1_LUT4AB/E6BEG[5] Tile_X6Y1_LUT4AB/E6BEG[6] Tile_X6Y1_LUT4AB/E6BEG[7] Tile_X6Y1_LUT4AB/E6BEG[8]
+ Tile_X6Y1_LUT4AB/E6BEG[9] Tile_X8Y1_LUT4AB/EE4END[0] Tile_X8Y1_LUT4AB/EE4END[10]
+ Tile_X8Y1_LUT4AB/EE4END[11] Tile_X8Y1_LUT4AB/EE4END[12] Tile_X8Y1_LUT4AB/EE4END[13]
+ Tile_X8Y1_LUT4AB/EE4END[14] Tile_X8Y1_LUT4AB/EE4END[15] Tile_X8Y1_LUT4AB/EE4END[1]
+ Tile_X8Y1_LUT4AB/EE4END[2] Tile_X8Y1_LUT4AB/EE4END[3] Tile_X8Y1_LUT4AB/EE4END[4]
+ Tile_X8Y1_LUT4AB/EE4END[5] Tile_X8Y1_LUT4AB/EE4END[6] Tile_X8Y1_LUT4AB/EE4END[7]
+ Tile_X8Y1_LUT4AB/EE4END[8] Tile_X8Y1_LUT4AB/EE4END[9] Tile_X6Y1_LUT4AB/EE4BEG[0]
+ Tile_X6Y1_LUT4AB/EE4BEG[10] Tile_X6Y1_LUT4AB/EE4BEG[11] Tile_X6Y1_LUT4AB/EE4BEG[12]
+ Tile_X6Y1_LUT4AB/EE4BEG[13] Tile_X6Y1_LUT4AB/EE4BEG[14] Tile_X6Y1_LUT4AB/EE4BEG[15]
+ Tile_X6Y1_LUT4AB/EE4BEG[1] Tile_X6Y1_LUT4AB/EE4BEG[2] Tile_X6Y1_LUT4AB/EE4BEG[3]
+ Tile_X6Y1_LUT4AB/EE4BEG[4] Tile_X6Y1_LUT4AB/EE4BEG[5] Tile_X6Y1_LUT4AB/EE4BEG[6]
+ Tile_X6Y1_LUT4AB/EE4BEG[7] Tile_X6Y1_LUT4AB/EE4BEG[8] Tile_X6Y1_LUT4AB/EE4BEG[9]
+ Tile_X6Y1_LUT4AB/FrameData_O[0] Tile_X6Y1_LUT4AB/FrameData_O[10] Tile_X6Y1_LUT4AB/FrameData_O[11]
+ Tile_X6Y1_LUT4AB/FrameData_O[12] Tile_X6Y1_LUT4AB/FrameData_O[13] Tile_X6Y1_LUT4AB/FrameData_O[14]
+ Tile_X6Y1_LUT4AB/FrameData_O[15] Tile_X6Y1_LUT4AB/FrameData_O[16] Tile_X6Y1_LUT4AB/FrameData_O[17]
+ Tile_X6Y1_LUT4AB/FrameData_O[18] Tile_X6Y1_LUT4AB/FrameData_O[19] Tile_X6Y1_LUT4AB/FrameData_O[1]
+ Tile_X6Y1_LUT4AB/FrameData_O[20] Tile_X6Y1_LUT4AB/FrameData_O[21] Tile_X6Y1_LUT4AB/FrameData_O[22]
+ Tile_X6Y1_LUT4AB/FrameData_O[23] Tile_X6Y1_LUT4AB/FrameData_O[24] Tile_X6Y1_LUT4AB/FrameData_O[25]
+ Tile_X6Y1_LUT4AB/FrameData_O[26] Tile_X6Y1_LUT4AB/FrameData_O[27] Tile_X6Y1_LUT4AB/FrameData_O[28]
+ Tile_X6Y1_LUT4AB/FrameData_O[29] Tile_X6Y1_LUT4AB/FrameData_O[2] Tile_X6Y1_LUT4AB/FrameData_O[30]
+ Tile_X6Y1_LUT4AB/FrameData_O[31] Tile_X6Y1_LUT4AB/FrameData_O[3] Tile_X6Y1_LUT4AB/FrameData_O[4]
+ Tile_X6Y1_LUT4AB/FrameData_O[5] Tile_X6Y1_LUT4AB/FrameData_O[6] Tile_X6Y1_LUT4AB/FrameData_O[7]
+ Tile_X6Y1_LUT4AB/FrameData_O[8] Tile_X6Y1_LUT4AB/FrameData_O[9] Tile_X8Y1_LUT4AB/FrameData[0]
+ Tile_X8Y1_LUT4AB/FrameData[10] Tile_X8Y1_LUT4AB/FrameData[11] Tile_X8Y1_LUT4AB/FrameData[12]
+ Tile_X8Y1_LUT4AB/FrameData[13] Tile_X8Y1_LUT4AB/FrameData[14] Tile_X8Y1_LUT4AB/FrameData[15]
+ Tile_X8Y1_LUT4AB/FrameData[16] Tile_X8Y1_LUT4AB/FrameData[17] Tile_X8Y1_LUT4AB/FrameData[18]
+ Tile_X8Y1_LUT4AB/FrameData[19] Tile_X8Y1_LUT4AB/FrameData[1] Tile_X8Y1_LUT4AB/FrameData[20]
+ Tile_X8Y1_LUT4AB/FrameData[21] Tile_X8Y1_LUT4AB/FrameData[22] Tile_X8Y1_LUT4AB/FrameData[23]
+ Tile_X8Y1_LUT4AB/FrameData[24] Tile_X8Y1_LUT4AB/FrameData[25] Tile_X8Y1_LUT4AB/FrameData[26]
+ Tile_X8Y1_LUT4AB/FrameData[27] Tile_X8Y1_LUT4AB/FrameData[28] Tile_X8Y1_LUT4AB/FrameData[29]
+ Tile_X8Y1_LUT4AB/FrameData[2] Tile_X8Y1_LUT4AB/FrameData[30] Tile_X8Y1_LUT4AB/FrameData[31]
+ Tile_X8Y1_LUT4AB/FrameData[3] Tile_X8Y1_LUT4AB/FrameData[4] Tile_X8Y1_LUT4AB/FrameData[5]
+ Tile_X8Y1_LUT4AB/FrameData[6] Tile_X8Y1_LUT4AB/FrameData[7] Tile_X8Y1_LUT4AB/FrameData[8]
+ Tile_X8Y1_LUT4AB/FrameData[9] Tile_X7Y0_N_term_DSP/FrameStrobe[0] Tile_X7Y0_N_term_DSP/FrameStrobe[10]
+ Tile_X7Y0_N_term_DSP/FrameStrobe[11] Tile_X7Y0_N_term_DSP/FrameStrobe[12] Tile_X7Y0_N_term_DSP/FrameStrobe[13]
+ Tile_X7Y0_N_term_DSP/FrameStrobe[14] Tile_X7Y0_N_term_DSP/FrameStrobe[15] Tile_X7Y0_N_term_DSP/FrameStrobe[16]
+ Tile_X7Y0_N_term_DSP/FrameStrobe[17] Tile_X7Y0_N_term_DSP/FrameStrobe[18] Tile_X7Y0_N_term_DSP/FrameStrobe[19]
+ Tile_X7Y0_N_term_DSP/FrameStrobe[1] Tile_X7Y0_N_term_DSP/FrameStrobe[2] Tile_X7Y0_N_term_DSP/FrameStrobe[3]
+ Tile_X7Y0_N_term_DSP/FrameStrobe[4] Tile_X7Y0_N_term_DSP/FrameStrobe[5] Tile_X7Y0_N_term_DSP/FrameStrobe[6]
+ Tile_X7Y0_N_term_DSP/FrameStrobe[7] Tile_X7Y0_N_term_DSP/FrameStrobe[8] Tile_X7Y0_N_term_DSP/FrameStrobe[9]
+ Tile_X7Y0_N_term_DSP/N1END[0] Tile_X7Y0_N_term_DSP/N1END[1] Tile_X7Y0_N_term_DSP/N1END[2]
+ Tile_X7Y0_N_term_DSP/N1END[3] Tile_X7Y0_N_term_DSP/N2MID[0] Tile_X7Y0_N_term_DSP/N2MID[1]
+ Tile_X7Y0_N_term_DSP/N2MID[2] Tile_X7Y0_N_term_DSP/N2MID[3] Tile_X7Y0_N_term_DSP/N2MID[4]
+ Tile_X7Y0_N_term_DSP/N2MID[5] Tile_X7Y0_N_term_DSP/N2MID[6] Tile_X7Y0_N_term_DSP/N2MID[7]
+ Tile_X7Y0_N_term_DSP/N2END[0] Tile_X7Y0_N_term_DSP/N2END[1] Tile_X7Y0_N_term_DSP/N2END[2]
+ Tile_X7Y0_N_term_DSP/N2END[3] Tile_X7Y0_N_term_DSP/N2END[4] Tile_X7Y0_N_term_DSP/N2END[5]
+ Tile_X7Y0_N_term_DSP/N2END[6] Tile_X7Y0_N_term_DSP/N2END[7] Tile_X7Y0_N_term_DSP/N4END[0]
+ Tile_X7Y0_N_term_DSP/N4END[10] Tile_X7Y0_N_term_DSP/N4END[11] Tile_X7Y0_N_term_DSP/N4END[12]
+ Tile_X7Y0_N_term_DSP/N4END[13] Tile_X7Y0_N_term_DSP/N4END[14] Tile_X7Y0_N_term_DSP/N4END[15]
+ Tile_X7Y0_N_term_DSP/N4END[1] Tile_X7Y0_N_term_DSP/N4END[2] Tile_X7Y0_N_term_DSP/N4END[3]
+ Tile_X7Y0_N_term_DSP/N4END[4] Tile_X7Y0_N_term_DSP/N4END[5] Tile_X7Y0_N_term_DSP/N4END[6]
+ Tile_X7Y0_N_term_DSP/N4END[7] Tile_X7Y0_N_term_DSP/N4END[8] Tile_X7Y0_N_term_DSP/N4END[9]
+ Tile_X7Y0_N_term_DSP/NN4END[0] Tile_X7Y0_N_term_DSP/NN4END[10] Tile_X7Y0_N_term_DSP/NN4END[11]
+ Tile_X7Y0_N_term_DSP/NN4END[12] Tile_X7Y0_N_term_DSP/NN4END[13] Tile_X7Y0_N_term_DSP/NN4END[14]
+ Tile_X7Y0_N_term_DSP/NN4END[15] Tile_X7Y0_N_term_DSP/NN4END[1] Tile_X7Y0_N_term_DSP/NN4END[2]
+ Tile_X7Y0_N_term_DSP/NN4END[3] Tile_X7Y0_N_term_DSP/NN4END[4] Tile_X7Y0_N_term_DSP/NN4END[5]
+ Tile_X7Y0_N_term_DSP/NN4END[6] Tile_X7Y0_N_term_DSP/NN4END[7] Tile_X7Y0_N_term_DSP/NN4END[8]
+ Tile_X7Y0_N_term_DSP/NN4END[9] Tile_X7Y0_N_term_DSP/S1BEG[0] Tile_X7Y0_N_term_DSP/S1BEG[1]
+ Tile_X7Y0_N_term_DSP/S1BEG[2] Tile_X7Y0_N_term_DSP/S1BEG[3] Tile_X7Y0_N_term_DSP/S2BEGb[0]
+ Tile_X7Y0_N_term_DSP/S2BEGb[1] Tile_X7Y0_N_term_DSP/S2BEGb[2] Tile_X7Y0_N_term_DSP/S2BEGb[3]
+ Tile_X7Y0_N_term_DSP/S2BEGb[4] Tile_X7Y0_N_term_DSP/S2BEGb[5] Tile_X7Y0_N_term_DSP/S2BEGb[6]
+ Tile_X7Y0_N_term_DSP/S2BEGb[7] Tile_X7Y0_N_term_DSP/S2BEG[0] Tile_X7Y0_N_term_DSP/S2BEG[1]
+ Tile_X7Y0_N_term_DSP/S2BEG[2] Tile_X7Y0_N_term_DSP/S2BEG[3] Tile_X7Y0_N_term_DSP/S2BEG[4]
+ Tile_X7Y0_N_term_DSP/S2BEG[5] Tile_X7Y0_N_term_DSP/S2BEG[6] Tile_X7Y0_N_term_DSP/S2BEG[7]
+ Tile_X7Y0_N_term_DSP/S4BEG[0] Tile_X7Y0_N_term_DSP/S4BEG[10] Tile_X7Y0_N_term_DSP/S4BEG[11]
+ Tile_X7Y0_N_term_DSP/S4BEG[12] Tile_X7Y0_N_term_DSP/S4BEG[13] Tile_X7Y0_N_term_DSP/S4BEG[14]
+ Tile_X7Y0_N_term_DSP/S4BEG[15] Tile_X7Y0_N_term_DSP/S4BEG[1] Tile_X7Y0_N_term_DSP/S4BEG[2]
+ Tile_X7Y0_N_term_DSP/S4BEG[3] Tile_X7Y0_N_term_DSP/S4BEG[4] Tile_X7Y0_N_term_DSP/S4BEG[5]
+ Tile_X7Y0_N_term_DSP/S4BEG[6] Tile_X7Y0_N_term_DSP/S4BEG[7] Tile_X7Y0_N_term_DSP/S4BEG[8]
+ Tile_X7Y0_N_term_DSP/S4BEG[9] Tile_X7Y0_N_term_DSP/SS4BEG[0] Tile_X7Y0_N_term_DSP/SS4BEG[10]
+ Tile_X7Y0_N_term_DSP/SS4BEG[11] Tile_X7Y0_N_term_DSP/SS4BEG[12] Tile_X7Y0_N_term_DSP/SS4BEG[13]
+ Tile_X7Y0_N_term_DSP/SS4BEG[14] Tile_X7Y0_N_term_DSP/SS4BEG[15] Tile_X7Y0_N_term_DSP/SS4BEG[1]
+ Tile_X7Y0_N_term_DSP/SS4BEG[2] Tile_X7Y0_N_term_DSP/SS4BEG[3] Tile_X7Y0_N_term_DSP/SS4BEG[4]
+ Tile_X7Y0_N_term_DSP/SS4BEG[5] Tile_X7Y0_N_term_DSP/SS4BEG[6] Tile_X7Y0_N_term_DSP/SS4BEG[7]
+ Tile_X7Y0_N_term_DSP/SS4BEG[8] Tile_X7Y0_N_term_DSP/SS4BEG[9] Tile_X7Y0_N_term_DSP/UserCLK
+ Tile_X6Y1_LUT4AB/W1END[0] Tile_X6Y1_LUT4AB/W1END[1] Tile_X6Y1_LUT4AB/W1END[2] Tile_X6Y1_LUT4AB/W1END[3]
+ Tile_X8Y1_LUT4AB/W1BEG[0] Tile_X8Y1_LUT4AB/W1BEG[1] Tile_X8Y1_LUT4AB/W1BEG[2] Tile_X8Y1_LUT4AB/W1BEG[3]
+ Tile_X6Y1_LUT4AB/W2MID[0] Tile_X6Y1_LUT4AB/W2MID[1] Tile_X6Y1_LUT4AB/W2MID[2] Tile_X6Y1_LUT4AB/W2MID[3]
+ Tile_X6Y1_LUT4AB/W2MID[4] Tile_X6Y1_LUT4AB/W2MID[5] Tile_X6Y1_LUT4AB/W2MID[6] Tile_X6Y1_LUT4AB/W2MID[7]
+ Tile_X6Y1_LUT4AB/W2END[0] Tile_X6Y1_LUT4AB/W2END[1] Tile_X6Y1_LUT4AB/W2END[2] Tile_X6Y1_LUT4AB/W2END[3]
+ Tile_X6Y1_LUT4AB/W2END[4] Tile_X6Y1_LUT4AB/W2END[5] Tile_X6Y1_LUT4AB/W2END[6] Tile_X6Y1_LUT4AB/W2END[7]
+ Tile_X8Y1_LUT4AB/W2BEGb[0] Tile_X8Y1_LUT4AB/W2BEGb[1] Tile_X8Y1_LUT4AB/W2BEGb[2]
+ Tile_X8Y1_LUT4AB/W2BEGb[3] Tile_X8Y1_LUT4AB/W2BEGb[4] Tile_X8Y1_LUT4AB/W2BEGb[5]
+ Tile_X8Y1_LUT4AB/W2BEGb[6] Tile_X8Y1_LUT4AB/W2BEGb[7] Tile_X8Y1_LUT4AB/W2BEG[0]
+ Tile_X8Y1_LUT4AB/W2BEG[1] Tile_X8Y1_LUT4AB/W2BEG[2] Tile_X8Y1_LUT4AB/W2BEG[3] Tile_X8Y1_LUT4AB/W2BEG[4]
+ Tile_X8Y1_LUT4AB/W2BEG[5] Tile_X8Y1_LUT4AB/W2BEG[6] Tile_X8Y1_LUT4AB/W2BEG[7] Tile_X6Y1_LUT4AB/W6END[0]
+ Tile_X6Y1_LUT4AB/W6END[10] Tile_X6Y1_LUT4AB/W6END[11] Tile_X6Y1_LUT4AB/W6END[1]
+ Tile_X6Y1_LUT4AB/W6END[2] Tile_X6Y1_LUT4AB/W6END[3] Tile_X6Y1_LUT4AB/W6END[4] Tile_X6Y1_LUT4AB/W6END[5]
+ Tile_X6Y1_LUT4AB/W6END[6] Tile_X6Y1_LUT4AB/W6END[7] Tile_X6Y1_LUT4AB/W6END[8] Tile_X6Y1_LUT4AB/W6END[9]
+ Tile_X8Y1_LUT4AB/W6BEG[0] Tile_X8Y1_LUT4AB/W6BEG[10] Tile_X8Y1_LUT4AB/W6BEG[11]
+ Tile_X8Y1_LUT4AB/W6BEG[1] Tile_X8Y1_LUT4AB/W6BEG[2] Tile_X8Y1_LUT4AB/W6BEG[3] Tile_X8Y1_LUT4AB/W6BEG[4]
+ Tile_X8Y1_LUT4AB/W6BEG[5] Tile_X8Y1_LUT4AB/W6BEG[6] Tile_X8Y1_LUT4AB/W6BEG[7] Tile_X8Y1_LUT4AB/W6BEG[8]
+ Tile_X8Y1_LUT4AB/W6BEG[9] Tile_X6Y1_LUT4AB/WW4END[0] Tile_X6Y1_LUT4AB/WW4END[10]
+ Tile_X6Y1_LUT4AB/WW4END[11] Tile_X6Y1_LUT4AB/WW4END[12] Tile_X6Y1_LUT4AB/WW4END[13]
+ Tile_X6Y1_LUT4AB/WW4END[14] Tile_X6Y1_LUT4AB/WW4END[15] Tile_X6Y1_LUT4AB/WW4END[1]
+ Tile_X6Y1_LUT4AB/WW4END[2] Tile_X6Y1_LUT4AB/WW4END[3] Tile_X6Y1_LUT4AB/WW4END[4]
+ Tile_X6Y1_LUT4AB/WW4END[5] Tile_X6Y1_LUT4AB/WW4END[6] Tile_X6Y1_LUT4AB/WW4END[7]
+ Tile_X6Y1_LUT4AB/WW4END[8] Tile_X6Y1_LUT4AB/WW4END[9] Tile_X8Y1_LUT4AB/WW4BEG[0]
+ Tile_X8Y1_LUT4AB/WW4BEG[10] Tile_X8Y1_LUT4AB/WW4BEG[11] Tile_X8Y1_LUT4AB/WW4BEG[12]
+ Tile_X8Y1_LUT4AB/WW4BEG[13] Tile_X8Y1_LUT4AB/WW4BEG[14] Tile_X8Y1_LUT4AB/WW4BEG[15]
+ Tile_X8Y1_LUT4AB/WW4BEG[1] Tile_X8Y1_LUT4AB/WW4BEG[2] Tile_X8Y1_LUT4AB/WW4BEG[3]
+ Tile_X8Y1_LUT4AB/WW4BEG[4] Tile_X8Y1_LUT4AB/WW4BEG[5] Tile_X8Y1_LUT4AB/WW4BEG[6]
+ Tile_X8Y1_LUT4AB/WW4BEG[7] Tile_X8Y1_LUT4AB/WW4BEG[8] Tile_X8Y1_LUT4AB/WW4BEG[9]
+ Tile_X8Y2_LUT4AB/E1END[0] Tile_X8Y2_LUT4AB/E1END[1] Tile_X8Y2_LUT4AB/E1END[2] Tile_X8Y2_LUT4AB/E1END[3]
+ Tile_X6Y2_LUT4AB/E1BEG[0] Tile_X6Y2_LUT4AB/E1BEG[1] Tile_X6Y2_LUT4AB/E1BEG[2] Tile_X6Y2_LUT4AB/E1BEG[3]
+ Tile_X8Y2_LUT4AB/E2MID[0] Tile_X8Y2_LUT4AB/E2MID[1] Tile_X8Y2_LUT4AB/E2MID[2] Tile_X8Y2_LUT4AB/E2MID[3]
+ Tile_X8Y2_LUT4AB/E2MID[4] Tile_X8Y2_LUT4AB/E2MID[5] Tile_X8Y2_LUT4AB/E2MID[6] Tile_X8Y2_LUT4AB/E2MID[7]
+ Tile_X8Y2_LUT4AB/E2END[0] Tile_X8Y2_LUT4AB/E2END[1] Tile_X8Y2_LUT4AB/E2END[2] Tile_X8Y2_LUT4AB/E2END[3]
+ Tile_X8Y2_LUT4AB/E2END[4] Tile_X8Y2_LUT4AB/E2END[5] Tile_X8Y2_LUT4AB/E2END[6] Tile_X8Y2_LUT4AB/E2END[7]
+ Tile_X6Y2_LUT4AB/E2BEGb[0] Tile_X6Y2_LUT4AB/E2BEGb[1] Tile_X6Y2_LUT4AB/E2BEGb[2]
+ Tile_X6Y2_LUT4AB/E2BEGb[3] Tile_X6Y2_LUT4AB/E2BEGb[4] Tile_X6Y2_LUT4AB/E2BEGb[5]
+ Tile_X6Y2_LUT4AB/E2BEGb[6] Tile_X6Y2_LUT4AB/E2BEGb[7] Tile_X6Y2_LUT4AB/E2BEG[0]
+ Tile_X6Y2_LUT4AB/E2BEG[1] Tile_X6Y2_LUT4AB/E2BEG[2] Tile_X6Y2_LUT4AB/E2BEG[3] Tile_X6Y2_LUT4AB/E2BEG[4]
+ Tile_X6Y2_LUT4AB/E2BEG[5] Tile_X6Y2_LUT4AB/E2BEG[6] Tile_X6Y2_LUT4AB/E2BEG[7] Tile_X8Y2_LUT4AB/E6END[0]
+ Tile_X8Y2_LUT4AB/E6END[10] Tile_X8Y2_LUT4AB/E6END[11] Tile_X8Y2_LUT4AB/E6END[1]
+ Tile_X8Y2_LUT4AB/E6END[2] Tile_X8Y2_LUT4AB/E6END[3] Tile_X8Y2_LUT4AB/E6END[4] Tile_X8Y2_LUT4AB/E6END[5]
+ Tile_X8Y2_LUT4AB/E6END[6] Tile_X8Y2_LUT4AB/E6END[7] Tile_X8Y2_LUT4AB/E6END[8] Tile_X8Y2_LUT4AB/E6END[9]
+ Tile_X6Y2_LUT4AB/E6BEG[0] Tile_X6Y2_LUT4AB/E6BEG[10] Tile_X6Y2_LUT4AB/E6BEG[11]
+ Tile_X6Y2_LUT4AB/E6BEG[1] Tile_X6Y2_LUT4AB/E6BEG[2] Tile_X6Y2_LUT4AB/E6BEG[3] Tile_X6Y2_LUT4AB/E6BEG[4]
+ Tile_X6Y2_LUT4AB/E6BEG[5] Tile_X6Y2_LUT4AB/E6BEG[6] Tile_X6Y2_LUT4AB/E6BEG[7] Tile_X6Y2_LUT4AB/E6BEG[8]
+ Tile_X6Y2_LUT4AB/E6BEG[9] Tile_X8Y2_LUT4AB/EE4END[0] Tile_X8Y2_LUT4AB/EE4END[10]
+ Tile_X8Y2_LUT4AB/EE4END[11] Tile_X8Y2_LUT4AB/EE4END[12] Tile_X8Y2_LUT4AB/EE4END[13]
+ Tile_X8Y2_LUT4AB/EE4END[14] Tile_X8Y2_LUT4AB/EE4END[15] Tile_X8Y2_LUT4AB/EE4END[1]
+ Tile_X8Y2_LUT4AB/EE4END[2] Tile_X8Y2_LUT4AB/EE4END[3] Tile_X8Y2_LUT4AB/EE4END[4]
+ Tile_X8Y2_LUT4AB/EE4END[5] Tile_X8Y2_LUT4AB/EE4END[6] Tile_X8Y2_LUT4AB/EE4END[7]
+ Tile_X8Y2_LUT4AB/EE4END[8] Tile_X8Y2_LUT4AB/EE4END[9] Tile_X6Y2_LUT4AB/EE4BEG[0]
+ Tile_X6Y2_LUT4AB/EE4BEG[10] Tile_X6Y2_LUT4AB/EE4BEG[11] Tile_X6Y2_LUT4AB/EE4BEG[12]
+ Tile_X6Y2_LUT4AB/EE4BEG[13] Tile_X6Y2_LUT4AB/EE4BEG[14] Tile_X6Y2_LUT4AB/EE4BEG[15]
+ Tile_X6Y2_LUT4AB/EE4BEG[1] Tile_X6Y2_LUT4AB/EE4BEG[2] Tile_X6Y2_LUT4AB/EE4BEG[3]
+ Tile_X6Y2_LUT4AB/EE4BEG[4] Tile_X6Y2_LUT4AB/EE4BEG[5] Tile_X6Y2_LUT4AB/EE4BEG[6]
+ Tile_X6Y2_LUT4AB/EE4BEG[7] Tile_X6Y2_LUT4AB/EE4BEG[8] Tile_X6Y2_LUT4AB/EE4BEG[9]
+ Tile_X6Y2_LUT4AB/FrameData_O[0] Tile_X6Y2_LUT4AB/FrameData_O[10] Tile_X6Y2_LUT4AB/FrameData_O[11]
+ Tile_X6Y2_LUT4AB/FrameData_O[12] Tile_X6Y2_LUT4AB/FrameData_O[13] Tile_X6Y2_LUT4AB/FrameData_O[14]
+ Tile_X6Y2_LUT4AB/FrameData_O[15] Tile_X6Y2_LUT4AB/FrameData_O[16] Tile_X6Y2_LUT4AB/FrameData_O[17]
+ Tile_X6Y2_LUT4AB/FrameData_O[18] Tile_X6Y2_LUT4AB/FrameData_O[19] Tile_X6Y2_LUT4AB/FrameData_O[1]
+ Tile_X6Y2_LUT4AB/FrameData_O[20] Tile_X6Y2_LUT4AB/FrameData_O[21] Tile_X6Y2_LUT4AB/FrameData_O[22]
+ Tile_X6Y2_LUT4AB/FrameData_O[23] Tile_X6Y2_LUT4AB/FrameData_O[24] Tile_X6Y2_LUT4AB/FrameData_O[25]
+ Tile_X6Y2_LUT4AB/FrameData_O[26] Tile_X6Y2_LUT4AB/FrameData_O[27] Tile_X6Y2_LUT4AB/FrameData_O[28]
+ Tile_X6Y2_LUT4AB/FrameData_O[29] Tile_X6Y2_LUT4AB/FrameData_O[2] Tile_X6Y2_LUT4AB/FrameData_O[30]
+ Tile_X6Y2_LUT4AB/FrameData_O[31] Tile_X6Y2_LUT4AB/FrameData_O[3] Tile_X6Y2_LUT4AB/FrameData_O[4]
+ Tile_X6Y2_LUT4AB/FrameData_O[5] Tile_X6Y2_LUT4AB/FrameData_O[6] Tile_X6Y2_LUT4AB/FrameData_O[7]
+ Tile_X6Y2_LUT4AB/FrameData_O[8] Tile_X6Y2_LUT4AB/FrameData_O[9] Tile_X8Y2_LUT4AB/FrameData[0]
+ Tile_X8Y2_LUT4AB/FrameData[10] Tile_X8Y2_LUT4AB/FrameData[11] Tile_X8Y2_LUT4AB/FrameData[12]
+ Tile_X8Y2_LUT4AB/FrameData[13] Tile_X8Y2_LUT4AB/FrameData[14] Tile_X8Y2_LUT4AB/FrameData[15]
+ Tile_X8Y2_LUT4AB/FrameData[16] Tile_X8Y2_LUT4AB/FrameData[17] Tile_X8Y2_LUT4AB/FrameData[18]
+ Tile_X8Y2_LUT4AB/FrameData[19] Tile_X8Y2_LUT4AB/FrameData[1] Tile_X8Y2_LUT4AB/FrameData[20]
+ Tile_X8Y2_LUT4AB/FrameData[21] Tile_X8Y2_LUT4AB/FrameData[22] Tile_X8Y2_LUT4AB/FrameData[23]
+ Tile_X8Y2_LUT4AB/FrameData[24] Tile_X8Y2_LUT4AB/FrameData[25] Tile_X8Y2_LUT4AB/FrameData[26]
+ Tile_X8Y2_LUT4AB/FrameData[27] Tile_X8Y2_LUT4AB/FrameData[28] Tile_X8Y2_LUT4AB/FrameData[29]
+ Tile_X8Y2_LUT4AB/FrameData[2] Tile_X8Y2_LUT4AB/FrameData[30] Tile_X8Y2_LUT4AB/FrameData[31]
+ Tile_X8Y2_LUT4AB/FrameData[3] Tile_X8Y2_LUT4AB/FrameData[4] Tile_X8Y2_LUT4AB/FrameData[5]
+ Tile_X8Y2_LUT4AB/FrameData[6] Tile_X8Y2_LUT4AB/FrameData[7] Tile_X8Y2_LUT4AB/FrameData[8]
+ Tile_X8Y2_LUT4AB/FrameData[9] Tile_X7Y1_DSP/Tile_X0Y1_FrameStrobe[0] Tile_X7Y1_DSP/Tile_X0Y1_FrameStrobe[10]
+ Tile_X7Y1_DSP/Tile_X0Y1_FrameStrobe[11] Tile_X7Y1_DSP/Tile_X0Y1_FrameStrobe[12]
+ Tile_X7Y1_DSP/Tile_X0Y1_FrameStrobe[13] Tile_X7Y1_DSP/Tile_X0Y1_FrameStrobe[14]
+ Tile_X7Y1_DSP/Tile_X0Y1_FrameStrobe[15] Tile_X7Y1_DSP/Tile_X0Y1_FrameStrobe[16]
+ Tile_X7Y1_DSP/Tile_X0Y1_FrameStrobe[17] Tile_X7Y1_DSP/Tile_X0Y1_FrameStrobe[18]
+ Tile_X7Y1_DSP/Tile_X0Y1_FrameStrobe[19] Tile_X7Y1_DSP/Tile_X0Y1_FrameStrobe[1] Tile_X7Y1_DSP/Tile_X0Y1_FrameStrobe[2]
+ Tile_X7Y1_DSP/Tile_X0Y1_FrameStrobe[3] Tile_X7Y1_DSP/Tile_X0Y1_FrameStrobe[4] Tile_X7Y1_DSP/Tile_X0Y1_FrameStrobe[5]
+ Tile_X7Y1_DSP/Tile_X0Y1_FrameStrobe[6] Tile_X7Y1_DSP/Tile_X0Y1_FrameStrobe[7] Tile_X7Y1_DSP/Tile_X0Y1_FrameStrobe[8]
+ Tile_X7Y1_DSP/Tile_X0Y1_FrameStrobe[9] Tile_X7Y3_DSP/Tile_X0Y0_N1BEG[0] Tile_X7Y3_DSP/Tile_X0Y0_N1BEG[1]
+ Tile_X7Y3_DSP/Tile_X0Y0_N1BEG[2] Tile_X7Y3_DSP/Tile_X0Y0_N1BEG[3] Tile_X7Y1_DSP/Tile_X0Y1_N2END[0]
+ Tile_X7Y1_DSP/Tile_X0Y1_N2END[1] Tile_X7Y1_DSP/Tile_X0Y1_N2END[2] Tile_X7Y1_DSP/Tile_X0Y1_N2END[3]
+ Tile_X7Y1_DSP/Tile_X0Y1_N2END[4] Tile_X7Y1_DSP/Tile_X0Y1_N2END[5] Tile_X7Y1_DSP/Tile_X0Y1_N2END[6]
+ Tile_X7Y1_DSP/Tile_X0Y1_N2END[7] Tile_X7Y3_DSP/Tile_X0Y0_N2BEG[0] Tile_X7Y3_DSP/Tile_X0Y0_N2BEG[1]
+ Tile_X7Y3_DSP/Tile_X0Y0_N2BEG[2] Tile_X7Y3_DSP/Tile_X0Y0_N2BEG[3] Tile_X7Y3_DSP/Tile_X0Y0_N2BEG[4]
+ Tile_X7Y3_DSP/Tile_X0Y0_N2BEG[5] Tile_X7Y3_DSP/Tile_X0Y0_N2BEG[6] Tile_X7Y3_DSP/Tile_X0Y0_N2BEG[7]
+ Tile_X7Y3_DSP/Tile_X0Y0_N4BEG[0] Tile_X7Y3_DSP/Tile_X0Y0_N4BEG[10] Tile_X7Y3_DSP/Tile_X0Y0_N4BEG[11]
+ Tile_X7Y3_DSP/Tile_X0Y0_N4BEG[12] Tile_X7Y3_DSP/Tile_X0Y0_N4BEG[13] Tile_X7Y3_DSP/Tile_X0Y0_N4BEG[14]
+ Tile_X7Y3_DSP/Tile_X0Y0_N4BEG[15] Tile_X7Y3_DSP/Tile_X0Y0_N4BEG[1] Tile_X7Y3_DSP/Tile_X0Y0_N4BEG[2]
+ Tile_X7Y3_DSP/Tile_X0Y0_N4BEG[3] Tile_X7Y3_DSP/Tile_X0Y0_N4BEG[4] Tile_X7Y3_DSP/Tile_X0Y0_N4BEG[5]
+ Tile_X7Y3_DSP/Tile_X0Y0_N4BEG[6] Tile_X7Y3_DSP/Tile_X0Y0_N4BEG[7] Tile_X7Y3_DSP/Tile_X0Y0_N4BEG[8]
+ Tile_X7Y3_DSP/Tile_X0Y0_N4BEG[9] Tile_X7Y3_DSP/Tile_X0Y0_NN4BEG[0] Tile_X7Y3_DSP/Tile_X0Y0_NN4BEG[10]
+ Tile_X7Y3_DSP/Tile_X0Y0_NN4BEG[11] Tile_X7Y3_DSP/Tile_X0Y0_NN4BEG[12] Tile_X7Y3_DSP/Tile_X0Y0_NN4BEG[13]
+ Tile_X7Y3_DSP/Tile_X0Y0_NN4BEG[14] Tile_X7Y3_DSP/Tile_X0Y0_NN4BEG[15] Tile_X7Y3_DSP/Tile_X0Y0_NN4BEG[1]
+ Tile_X7Y3_DSP/Tile_X0Y0_NN4BEG[2] Tile_X7Y3_DSP/Tile_X0Y0_NN4BEG[3] Tile_X7Y3_DSP/Tile_X0Y0_NN4BEG[4]
+ Tile_X7Y3_DSP/Tile_X0Y0_NN4BEG[5] Tile_X7Y3_DSP/Tile_X0Y0_NN4BEG[6] Tile_X7Y3_DSP/Tile_X0Y0_NN4BEG[7]
+ Tile_X7Y3_DSP/Tile_X0Y0_NN4BEG[8] Tile_X7Y3_DSP/Tile_X0Y0_NN4BEG[9] Tile_X7Y3_DSP/Tile_X0Y0_S1END[0]
+ Tile_X7Y3_DSP/Tile_X0Y0_S1END[1] Tile_X7Y3_DSP/Tile_X0Y0_S1END[2] Tile_X7Y3_DSP/Tile_X0Y0_S1END[3]
+ Tile_X7Y3_DSP/Tile_X0Y0_S2MID[0] Tile_X7Y3_DSP/Tile_X0Y0_S2MID[1] Tile_X7Y3_DSP/Tile_X0Y0_S2MID[2]
+ Tile_X7Y3_DSP/Tile_X0Y0_S2MID[3] Tile_X7Y3_DSP/Tile_X0Y0_S2MID[4] Tile_X7Y3_DSP/Tile_X0Y0_S2MID[5]
+ Tile_X7Y3_DSP/Tile_X0Y0_S2MID[6] Tile_X7Y3_DSP/Tile_X0Y0_S2MID[7] Tile_X7Y3_DSP/Tile_X0Y0_S2END[0]
+ Tile_X7Y3_DSP/Tile_X0Y0_S2END[1] Tile_X7Y3_DSP/Tile_X0Y0_S2END[2] Tile_X7Y3_DSP/Tile_X0Y0_S2END[3]
+ Tile_X7Y3_DSP/Tile_X0Y0_S2END[4] Tile_X7Y3_DSP/Tile_X0Y0_S2END[5] Tile_X7Y3_DSP/Tile_X0Y0_S2END[6]
+ Tile_X7Y3_DSP/Tile_X0Y0_S2END[7] Tile_X7Y3_DSP/Tile_X0Y0_S4END[0] Tile_X7Y3_DSP/Tile_X0Y0_S4END[10]
+ Tile_X7Y3_DSP/Tile_X0Y0_S4END[11] Tile_X7Y3_DSP/Tile_X0Y0_S4END[12] Tile_X7Y3_DSP/Tile_X0Y0_S4END[13]
+ Tile_X7Y3_DSP/Tile_X0Y0_S4END[14] Tile_X7Y3_DSP/Tile_X0Y0_S4END[15] Tile_X7Y3_DSP/Tile_X0Y0_S4END[1]
+ Tile_X7Y3_DSP/Tile_X0Y0_S4END[2] Tile_X7Y3_DSP/Tile_X0Y0_S4END[3] Tile_X7Y3_DSP/Tile_X0Y0_S4END[4]
+ Tile_X7Y3_DSP/Tile_X0Y0_S4END[5] Tile_X7Y3_DSP/Tile_X0Y0_S4END[6] Tile_X7Y3_DSP/Tile_X0Y0_S4END[7]
+ Tile_X7Y3_DSP/Tile_X0Y0_S4END[8] Tile_X7Y3_DSP/Tile_X0Y0_S4END[9] Tile_X7Y3_DSP/Tile_X0Y0_SS4END[0]
+ Tile_X7Y3_DSP/Tile_X0Y0_SS4END[10] Tile_X7Y3_DSP/Tile_X0Y0_SS4END[11] Tile_X7Y3_DSP/Tile_X0Y0_SS4END[12]
+ Tile_X7Y3_DSP/Tile_X0Y0_SS4END[13] Tile_X7Y3_DSP/Tile_X0Y0_SS4END[14] Tile_X7Y3_DSP/Tile_X0Y0_SS4END[15]
+ Tile_X7Y3_DSP/Tile_X0Y0_SS4END[1] Tile_X7Y3_DSP/Tile_X0Y0_SS4END[2] Tile_X7Y3_DSP/Tile_X0Y0_SS4END[3]
+ Tile_X7Y3_DSP/Tile_X0Y0_SS4END[4] Tile_X7Y3_DSP/Tile_X0Y0_SS4END[5] Tile_X7Y3_DSP/Tile_X0Y0_SS4END[6]
+ Tile_X7Y3_DSP/Tile_X0Y0_SS4END[7] Tile_X7Y3_DSP/Tile_X0Y0_SS4END[8] Tile_X7Y3_DSP/Tile_X0Y0_SS4END[9]
+ Tile_X7Y1_DSP/Tile_X0Y1_UserCLK Tile_X6Y2_LUT4AB/W1END[0] Tile_X6Y2_LUT4AB/W1END[1]
+ Tile_X6Y2_LUT4AB/W1END[2] Tile_X6Y2_LUT4AB/W1END[3] Tile_X8Y2_LUT4AB/W1BEG[0] Tile_X8Y2_LUT4AB/W1BEG[1]
+ Tile_X8Y2_LUT4AB/W1BEG[2] Tile_X8Y2_LUT4AB/W1BEG[3] Tile_X6Y2_LUT4AB/W2MID[0] Tile_X6Y2_LUT4AB/W2MID[1]
+ Tile_X6Y2_LUT4AB/W2MID[2] Tile_X6Y2_LUT4AB/W2MID[3] Tile_X6Y2_LUT4AB/W2MID[4] Tile_X6Y2_LUT4AB/W2MID[5]
+ Tile_X6Y2_LUT4AB/W2MID[6] Tile_X6Y2_LUT4AB/W2MID[7] Tile_X6Y2_LUT4AB/W2END[0] Tile_X6Y2_LUT4AB/W2END[1]
+ Tile_X6Y2_LUT4AB/W2END[2] Tile_X6Y2_LUT4AB/W2END[3] Tile_X6Y2_LUT4AB/W2END[4] Tile_X6Y2_LUT4AB/W2END[5]
+ Tile_X6Y2_LUT4AB/W2END[6] Tile_X6Y2_LUT4AB/W2END[7] Tile_X8Y2_LUT4AB/W2BEGb[0] Tile_X8Y2_LUT4AB/W2BEGb[1]
+ Tile_X8Y2_LUT4AB/W2BEGb[2] Tile_X8Y2_LUT4AB/W2BEGb[3] Tile_X8Y2_LUT4AB/W2BEGb[4]
+ Tile_X8Y2_LUT4AB/W2BEGb[5] Tile_X8Y2_LUT4AB/W2BEGb[6] Tile_X8Y2_LUT4AB/W2BEGb[7]
+ Tile_X8Y2_LUT4AB/W2BEG[0] Tile_X8Y2_LUT4AB/W2BEG[1] Tile_X8Y2_LUT4AB/W2BEG[2] Tile_X8Y2_LUT4AB/W2BEG[3]
+ Tile_X8Y2_LUT4AB/W2BEG[4] Tile_X8Y2_LUT4AB/W2BEG[5] Tile_X8Y2_LUT4AB/W2BEG[6] Tile_X8Y2_LUT4AB/W2BEG[7]
+ Tile_X6Y2_LUT4AB/W6END[0] Tile_X6Y2_LUT4AB/W6END[10] Tile_X6Y2_LUT4AB/W6END[11]
+ Tile_X6Y2_LUT4AB/W6END[1] Tile_X6Y2_LUT4AB/W6END[2] Tile_X6Y2_LUT4AB/W6END[3] Tile_X6Y2_LUT4AB/W6END[4]
+ Tile_X6Y2_LUT4AB/W6END[5] Tile_X6Y2_LUT4AB/W6END[6] Tile_X6Y2_LUT4AB/W6END[7] Tile_X6Y2_LUT4AB/W6END[8]
+ Tile_X6Y2_LUT4AB/W6END[9] Tile_X8Y2_LUT4AB/W6BEG[0] Tile_X8Y2_LUT4AB/W6BEG[10] Tile_X8Y2_LUT4AB/W6BEG[11]
+ Tile_X8Y2_LUT4AB/W6BEG[1] Tile_X8Y2_LUT4AB/W6BEG[2] Tile_X8Y2_LUT4AB/W6BEG[3] Tile_X8Y2_LUT4AB/W6BEG[4]
+ Tile_X8Y2_LUT4AB/W6BEG[5] Tile_X8Y2_LUT4AB/W6BEG[6] Tile_X8Y2_LUT4AB/W6BEG[7] Tile_X8Y2_LUT4AB/W6BEG[8]
+ Tile_X8Y2_LUT4AB/W6BEG[9] Tile_X6Y2_LUT4AB/WW4END[0] Tile_X6Y2_LUT4AB/WW4END[10]
+ Tile_X6Y2_LUT4AB/WW4END[11] Tile_X6Y2_LUT4AB/WW4END[12] Tile_X6Y2_LUT4AB/WW4END[13]
+ Tile_X6Y2_LUT4AB/WW4END[14] Tile_X6Y2_LUT4AB/WW4END[15] Tile_X6Y2_LUT4AB/WW4END[1]
+ Tile_X6Y2_LUT4AB/WW4END[2] Tile_X6Y2_LUT4AB/WW4END[3] Tile_X6Y2_LUT4AB/WW4END[4]
+ Tile_X6Y2_LUT4AB/WW4END[5] Tile_X6Y2_LUT4AB/WW4END[6] Tile_X6Y2_LUT4AB/WW4END[7]
+ Tile_X6Y2_LUT4AB/WW4END[8] Tile_X6Y2_LUT4AB/WW4END[9] Tile_X8Y2_LUT4AB/WW4BEG[0]
+ Tile_X8Y2_LUT4AB/WW4BEG[10] Tile_X8Y2_LUT4AB/WW4BEG[11] Tile_X8Y2_LUT4AB/WW4BEG[12]
+ Tile_X8Y2_LUT4AB/WW4BEG[13] Tile_X8Y2_LUT4AB/WW4BEG[14] Tile_X8Y2_LUT4AB/WW4BEG[15]
+ Tile_X8Y2_LUT4AB/WW4BEG[1] Tile_X8Y2_LUT4AB/WW4BEG[2] Tile_X8Y2_LUT4AB/WW4BEG[3]
+ Tile_X8Y2_LUT4AB/WW4BEG[4] Tile_X8Y2_LUT4AB/WW4BEG[5] Tile_X8Y2_LUT4AB/WW4BEG[6]
+ Tile_X8Y2_LUT4AB/WW4BEG[7] Tile_X8Y2_LUT4AB/WW4BEG[8] Tile_X8Y2_LUT4AB/WW4BEG[9]
+ VGND VPWR DSP
XTile_X2Y10_LUT4AB Tile_X2Y11_LUT4AB/Co Tile_X2Y9_LUT4AB/Ci Tile_X3Y10_LUT4AB/E1END[0]
+ Tile_X3Y10_LUT4AB/E1END[1] Tile_X3Y10_LUT4AB/E1END[2] Tile_X3Y10_LUT4AB/E1END[3]
+ Tile_X2Y10_LUT4AB/E1END[0] Tile_X2Y10_LUT4AB/E1END[1] Tile_X2Y10_LUT4AB/E1END[2]
+ Tile_X2Y10_LUT4AB/E1END[3] Tile_X3Y10_LUT4AB/E2MID[0] Tile_X3Y10_LUT4AB/E2MID[1]
+ Tile_X3Y10_LUT4AB/E2MID[2] Tile_X3Y10_LUT4AB/E2MID[3] Tile_X3Y10_LUT4AB/E2MID[4]
+ Tile_X3Y10_LUT4AB/E2MID[5] Tile_X3Y10_LUT4AB/E2MID[6] Tile_X3Y10_LUT4AB/E2MID[7]
+ Tile_X3Y10_LUT4AB/E2END[0] Tile_X3Y10_LUT4AB/E2END[1] Tile_X3Y10_LUT4AB/E2END[2]
+ Tile_X3Y10_LUT4AB/E2END[3] Tile_X3Y10_LUT4AB/E2END[4] Tile_X3Y10_LUT4AB/E2END[5]
+ Tile_X3Y10_LUT4AB/E2END[6] Tile_X3Y10_LUT4AB/E2END[7] Tile_X2Y10_LUT4AB/E2END[0]
+ Tile_X2Y10_LUT4AB/E2END[1] Tile_X2Y10_LUT4AB/E2END[2] Tile_X2Y10_LUT4AB/E2END[3]
+ Tile_X2Y10_LUT4AB/E2END[4] Tile_X2Y10_LUT4AB/E2END[5] Tile_X2Y10_LUT4AB/E2END[6]
+ Tile_X2Y10_LUT4AB/E2END[7] Tile_X2Y10_LUT4AB/E2MID[0] Tile_X2Y10_LUT4AB/E2MID[1]
+ Tile_X2Y10_LUT4AB/E2MID[2] Tile_X2Y10_LUT4AB/E2MID[3] Tile_X2Y10_LUT4AB/E2MID[4]
+ Tile_X2Y10_LUT4AB/E2MID[5] Tile_X2Y10_LUT4AB/E2MID[6] Tile_X2Y10_LUT4AB/E2MID[7]
+ Tile_X3Y10_LUT4AB/E6END[0] Tile_X3Y10_LUT4AB/E6END[10] Tile_X3Y10_LUT4AB/E6END[11]
+ Tile_X3Y10_LUT4AB/E6END[1] Tile_X3Y10_LUT4AB/E6END[2] Tile_X3Y10_LUT4AB/E6END[3]
+ Tile_X3Y10_LUT4AB/E6END[4] Tile_X3Y10_LUT4AB/E6END[5] Tile_X3Y10_LUT4AB/E6END[6]
+ Tile_X3Y10_LUT4AB/E6END[7] Tile_X3Y10_LUT4AB/E6END[8] Tile_X3Y10_LUT4AB/E6END[9]
+ Tile_X2Y10_LUT4AB/E6END[0] Tile_X2Y10_LUT4AB/E6END[10] Tile_X2Y10_LUT4AB/E6END[11]
+ Tile_X2Y10_LUT4AB/E6END[1] Tile_X2Y10_LUT4AB/E6END[2] Tile_X2Y10_LUT4AB/E6END[3]
+ Tile_X2Y10_LUT4AB/E6END[4] Tile_X2Y10_LUT4AB/E6END[5] Tile_X2Y10_LUT4AB/E6END[6]
+ Tile_X2Y10_LUT4AB/E6END[7] Tile_X2Y10_LUT4AB/E6END[8] Tile_X2Y10_LUT4AB/E6END[9]
+ Tile_X3Y10_LUT4AB/EE4END[0] Tile_X3Y10_LUT4AB/EE4END[10] Tile_X3Y10_LUT4AB/EE4END[11]
+ Tile_X3Y10_LUT4AB/EE4END[12] Tile_X3Y10_LUT4AB/EE4END[13] Tile_X3Y10_LUT4AB/EE4END[14]
+ Tile_X3Y10_LUT4AB/EE4END[15] Tile_X3Y10_LUT4AB/EE4END[1] Tile_X3Y10_LUT4AB/EE4END[2]
+ Tile_X3Y10_LUT4AB/EE4END[3] Tile_X3Y10_LUT4AB/EE4END[4] Tile_X3Y10_LUT4AB/EE4END[5]
+ Tile_X3Y10_LUT4AB/EE4END[6] Tile_X3Y10_LUT4AB/EE4END[7] Tile_X3Y10_LUT4AB/EE4END[8]
+ Tile_X3Y10_LUT4AB/EE4END[9] Tile_X2Y10_LUT4AB/EE4END[0] Tile_X2Y10_LUT4AB/EE4END[10]
+ Tile_X2Y10_LUT4AB/EE4END[11] Tile_X2Y10_LUT4AB/EE4END[12] Tile_X2Y10_LUT4AB/EE4END[13]
+ Tile_X2Y10_LUT4AB/EE4END[14] Tile_X2Y10_LUT4AB/EE4END[15] Tile_X2Y10_LUT4AB/EE4END[1]
+ Tile_X2Y10_LUT4AB/EE4END[2] Tile_X2Y10_LUT4AB/EE4END[3] Tile_X2Y10_LUT4AB/EE4END[4]
+ Tile_X2Y10_LUT4AB/EE4END[5] Tile_X2Y10_LUT4AB/EE4END[6] Tile_X2Y10_LUT4AB/EE4END[7]
+ Tile_X2Y10_LUT4AB/EE4END[8] Tile_X2Y10_LUT4AB/EE4END[9] Tile_X2Y10_LUT4AB/FrameData[0]
+ Tile_X2Y10_LUT4AB/FrameData[10] Tile_X2Y10_LUT4AB/FrameData[11] Tile_X2Y10_LUT4AB/FrameData[12]
+ Tile_X2Y10_LUT4AB/FrameData[13] Tile_X2Y10_LUT4AB/FrameData[14] Tile_X2Y10_LUT4AB/FrameData[15]
+ Tile_X2Y10_LUT4AB/FrameData[16] Tile_X2Y10_LUT4AB/FrameData[17] Tile_X2Y10_LUT4AB/FrameData[18]
+ Tile_X2Y10_LUT4AB/FrameData[19] Tile_X2Y10_LUT4AB/FrameData[1] Tile_X2Y10_LUT4AB/FrameData[20]
+ Tile_X2Y10_LUT4AB/FrameData[21] Tile_X2Y10_LUT4AB/FrameData[22] Tile_X2Y10_LUT4AB/FrameData[23]
+ Tile_X2Y10_LUT4AB/FrameData[24] Tile_X2Y10_LUT4AB/FrameData[25] Tile_X2Y10_LUT4AB/FrameData[26]
+ Tile_X2Y10_LUT4AB/FrameData[27] Tile_X2Y10_LUT4AB/FrameData[28] Tile_X2Y10_LUT4AB/FrameData[29]
+ Tile_X2Y10_LUT4AB/FrameData[2] Tile_X2Y10_LUT4AB/FrameData[30] Tile_X2Y10_LUT4AB/FrameData[31]
+ Tile_X2Y10_LUT4AB/FrameData[3] Tile_X2Y10_LUT4AB/FrameData[4] Tile_X2Y10_LUT4AB/FrameData[5]
+ Tile_X2Y10_LUT4AB/FrameData[6] Tile_X2Y10_LUT4AB/FrameData[7] Tile_X2Y10_LUT4AB/FrameData[8]
+ Tile_X2Y10_LUT4AB/FrameData[9] Tile_X3Y10_LUT4AB/FrameData[0] Tile_X3Y10_LUT4AB/FrameData[10]
+ Tile_X3Y10_LUT4AB/FrameData[11] Tile_X3Y10_LUT4AB/FrameData[12] Tile_X3Y10_LUT4AB/FrameData[13]
+ Tile_X3Y10_LUT4AB/FrameData[14] Tile_X3Y10_LUT4AB/FrameData[15] Tile_X3Y10_LUT4AB/FrameData[16]
+ Tile_X3Y10_LUT4AB/FrameData[17] Tile_X3Y10_LUT4AB/FrameData[18] Tile_X3Y10_LUT4AB/FrameData[19]
+ Tile_X3Y10_LUT4AB/FrameData[1] Tile_X3Y10_LUT4AB/FrameData[20] Tile_X3Y10_LUT4AB/FrameData[21]
+ Tile_X3Y10_LUT4AB/FrameData[22] Tile_X3Y10_LUT4AB/FrameData[23] Tile_X3Y10_LUT4AB/FrameData[24]
+ Tile_X3Y10_LUT4AB/FrameData[25] Tile_X3Y10_LUT4AB/FrameData[26] Tile_X3Y10_LUT4AB/FrameData[27]
+ Tile_X3Y10_LUT4AB/FrameData[28] Tile_X3Y10_LUT4AB/FrameData[29] Tile_X3Y10_LUT4AB/FrameData[2]
+ Tile_X3Y10_LUT4AB/FrameData[30] Tile_X3Y10_LUT4AB/FrameData[31] Tile_X3Y10_LUT4AB/FrameData[3]
+ Tile_X3Y10_LUT4AB/FrameData[4] Tile_X3Y10_LUT4AB/FrameData[5] Tile_X3Y10_LUT4AB/FrameData[6]
+ Tile_X3Y10_LUT4AB/FrameData[7] Tile_X3Y10_LUT4AB/FrameData[8] Tile_X3Y10_LUT4AB/FrameData[9]
+ Tile_X2Y10_LUT4AB/FrameStrobe[0] Tile_X2Y10_LUT4AB/FrameStrobe[10] Tile_X2Y10_LUT4AB/FrameStrobe[11]
+ Tile_X2Y10_LUT4AB/FrameStrobe[12] Tile_X2Y10_LUT4AB/FrameStrobe[13] Tile_X2Y10_LUT4AB/FrameStrobe[14]
+ Tile_X2Y10_LUT4AB/FrameStrobe[15] Tile_X2Y10_LUT4AB/FrameStrobe[16] Tile_X2Y10_LUT4AB/FrameStrobe[17]
+ Tile_X2Y10_LUT4AB/FrameStrobe[18] Tile_X2Y10_LUT4AB/FrameStrobe[19] Tile_X2Y10_LUT4AB/FrameStrobe[1]
+ Tile_X2Y10_LUT4AB/FrameStrobe[2] Tile_X2Y10_LUT4AB/FrameStrobe[3] Tile_X2Y10_LUT4AB/FrameStrobe[4]
+ Tile_X2Y10_LUT4AB/FrameStrobe[5] Tile_X2Y10_LUT4AB/FrameStrobe[6] Tile_X2Y10_LUT4AB/FrameStrobe[7]
+ Tile_X2Y10_LUT4AB/FrameStrobe[8] Tile_X2Y10_LUT4AB/FrameStrobe[9] Tile_X2Y9_LUT4AB/FrameStrobe[0]
+ Tile_X2Y9_LUT4AB/FrameStrobe[10] Tile_X2Y9_LUT4AB/FrameStrobe[11] Tile_X2Y9_LUT4AB/FrameStrobe[12]
+ Tile_X2Y9_LUT4AB/FrameStrobe[13] Tile_X2Y9_LUT4AB/FrameStrobe[14] Tile_X2Y9_LUT4AB/FrameStrobe[15]
+ Tile_X2Y9_LUT4AB/FrameStrobe[16] Tile_X2Y9_LUT4AB/FrameStrobe[17] Tile_X2Y9_LUT4AB/FrameStrobe[18]
+ Tile_X2Y9_LUT4AB/FrameStrobe[19] Tile_X2Y9_LUT4AB/FrameStrobe[1] Tile_X2Y9_LUT4AB/FrameStrobe[2]
+ Tile_X2Y9_LUT4AB/FrameStrobe[3] Tile_X2Y9_LUT4AB/FrameStrobe[4] Tile_X2Y9_LUT4AB/FrameStrobe[5]
+ Tile_X2Y9_LUT4AB/FrameStrobe[6] Tile_X2Y9_LUT4AB/FrameStrobe[7] Tile_X2Y9_LUT4AB/FrameStrobe[8]
+ Tile_X2Y9_LUT4AB/FrameStrobe[9] Tile_X2Y9_LUT4AB/N1END[0] Tile_X2Y9_LUT4AB/N1END[1]
+ Tile_X2Y9_LUT4AB/N1END[2] Tile_X2Y9_LUT4AB/N1END[3] Tile_X2Y11_LUT4AB/N1BEG[0] Tile_X2Y11_LUT4AB/N1BEG[1]
+ Tile_X2Y11_LUT4AB/N1BEG[2] Tile_X2Y11_LUT4AB/N1BEG[3] Tile_X2Y9_LUT4AB/N2MID[0]
+ Tile_X2Y9_LUT4AB/N2MID[1] Tile_X2Y9_LUT4AB/N2MID[2] Tile_X2Y9_LUT4AB/N2MID[3] Tile_X2Y9_LUT4AB/N2MID[4]
+ Tile_X2Y9_LUT4AB/N2MID[5] Tile_X2Y9_LUT4AB/N2MID[6] Tile_X2Y9_LUT4AB/N2MID[7] Tile_X2Y9_LUT4AB/N2END[0]
+ Tile_X2Y9_LUT4AB/N2END[1] Tile_X2Y9_LUT4AB/N2END[2] Tile_X2Y9_LUT4AB/N2END[3] Tile_X2Y9_LUT4AB/N2END[4]
+ Tile_X2Y9_LUT4AB/N2END[5] Tile_X2Y9_LUT4AB/N2END[6] Tile_X2Y9_LUT4AB/N2END[7] Tile_X2Y10_LUT4AB/N2END[0]
+ Tile_X2Y10_LUT4AB/N2END[1] Tile_X2Y10_LUT4AB/N2END[2] Tile_X2Y10_LUT4AB/N2END[3]
+ Tile_X2Y10_LUT4AB/N2END[4] Tile_X2Y10_LUT4AB/N2END[5] Tile_X2Y10_LUT4AB/N2END[6]
+ Tile_X2Y10_LUT4AB/N2END[7] Tile_X2Y11_LUT4AB/N2BEG[0] Tile_X2Y11_LUT4AB/N2BEG[1]
+ Tile_X2Y11_LUT4AB/N2BEG[2] Tile_X2Y11_LUT4AB/N2BEG[3] Tile_X2Y11_LUT4AB/N2BEG[4]
+ Tile_X2Y11_LUT4AB/N2BEG[5] Tile_X2Y11_LUT4AB/N2BEG[6] Tile_X2Y11_LUT4AB/N2BEG[7]
+ Tile_X2Y9_LUT4AB/N4END[0] Tile_X2Y9_LUT4AB/N4END[10] Tile_X2Y9_LUT4AB/N4END[11]
+ Tile_X2Y9_LUT4AB/N4END[12] Tile_X2Y9_LUT4AB/N4END[13] Tile_X2Y9_LUT4AB/N4END[14]
+ Tile_X2Y9_LUT4AB/N4END[15] Tile_X2Y9_LUT4AB/N4END[1] Tile_X2Y9_LUT4AB/N4END[2] Tile_X2Y9_LUT4AB/N4END[3]
+ Tile_X2Y9_LUT4AB/N4END[4] Tile_X2Y9_LUT4AB/N4END[5] Tile_X2Y9_LUT4AB/N4END[6] Tile_X2Y9_LUT4AB/N4END[7]
+ Tile_X2Y9_LUT4AB/N4END[8] Tile_X2Y9_LUT4AB/N4END[9] Tile_X2Y11_LUT4AB/N4BEG[0] Tile_X2Y11_LUT4AB/N4BEG[10]
+ Tile_X2Y11_LUT4AB/N4BEG[11] Tile_X2Y11_LUT4AB/N4BEG[12] Tile_X2Y11_LUT4AB/N4BEG[13]
+ Tile_X2Y11_LUT4AB/N4BEG[14] Tile_X2Y11_LUT4AB/N4BEG[15] Tile_X2Y11_LUT4AB/N4BEG[1]
+ Tile_X2Y11_LUT4AB/N4BEG[2] Tile_X2Y11_LUT4AB/N4BEG[3] Tile_X2Y11_LUT4AB/N4BEG[4]
+ Tile_X2Y11_LUT4AB/N4BEG[5] Tile_X2Y11_LUT4AB/N4BEG[6] Tile_X2Y11_LUT4AB/N4BEG[7]
+ Tile_X2Y11_LUT4AB/N4BEG[8] Tile_X2Y11_LUT4AB/N4BEG[9] Tile_X2Y9_LUT4AB/NN4END[0]
+ Tile_X2Y9_LUT4AB/NN4END[10] Tile_X2Y9_LUT4AB/NN4END[11] Tile_X2Y9_LUT4AB/NN4END[12]
+ Tile_X2Y9_LUT4AB/NN4END[13] Tile_X2Y9_LUT4AB/NN4END[14] Tile_X2Y9_LUT4AB/NN4END[15]
+ Tile_X2Y9_LUT4AB/NN4END[1] Tile_X2Y9_LUT4AB/NN4END[2] Tile_X2Y9_LUT4AB/NN4END[3]
+ Tile_X2Y9_LUT4AB/NN4END[4] Tile_X2Y9_LUT4AB/NN4END[5] Tile_X2Y9_LUT4AB/NN4END[6]
+ Tile_X2Y9_LUT4AB/NN4END[7] Tile_X2Y9_LUT4AB/NN4END[8] Tile_X2Y9_LUT4AB/NN4END[9]
+ Tile_X2Y11_LUT4AB/NN4BEG[0] Tile_X2Y11_LUT4AB/NN4BEG[10] Tile_X2Y11_LUT4AB/NN4BEG[11]
+ Tile_X2Y11_LUT4AB/NN4BEG[12] Tile_X2Y11_LUT4AB/NN4BEG[13] Tile_X2Y11_LUT4AB/NN4BEG[14]
+ Tile_X2Y11_LUT4AB/NN4BEG[15] Tile_X2Y11_LUT4AB/NN4BEG[1] Tile_X2Y11_LUT4AB/NN4BEG[2]
+ Tile_X2Y11_LUT4AB/NN4BEG[3] Tile_X2Y11_LUT4AB/NN4BEG[4] Tile_X2Y11_LUT4AB/NN4BEG[5]
+ Tile_X2Y11_LUT4AB/NN4BEG[6] Tile_X2Y11_LUT4AB/NN4BEG[7] Tile_X2Y11_LUT4AB/NN4BEG[8]
+ Tile_X2Y11_LUT4AB/NN4BEG[9] Tile_X2Y11_LUT4AB/S1END[0] Tile_X2Y11_LUT4AB/S1END[1]
+ Tile_X2Y11_LUT4AB/S1END[2] Tile_X2Y11_LUT4AB/S1END[3] Tile_X2Y9_LUT4AB/S1BEG[0]
+ Tile_X2Y9_LUT4AB/S1BEG[1] Tile_X2Y9_LUT4AB/S1BEG[2] Tile_X2Y9_LUT4AB/S1BEG[3] Tile_X2Y11_LUT4AB/S2MID[0]
+ Tile_X2Y11_LUT4AB/S2MID[1] Tile_X2Y11_LUT4AB/S2MID[2] Tile_X2Y11_LUT4AB/S2MID[3]
+ Tile_X2Y11_LUT4AB/S2MID[4] Tile_X2Y11_LUT4AB/S2MID[5] Tile_X2Y11_LUT4AB/S2MID[6]
+ Tile_X2Y11_LUT4AB/S2MID[7] Tile_X2Y11_LUT4AB/S2END[0] Tile_X2Y11_LUT4AB/S2END[1]
+ Tile_X2Y11_LUT4AB/S2END[2] Tile_X2Y11_LUT4AB/S2END[3] Tile_X2Y11_LUT4AB/S2END[4]
+ Tile_X2Y11_LUT4AB/S2END[5] Tile_X2Y11_LUT4AB/S2END[6] Tile_X2Y11_LUT4AB/S2END[7]
+ Tile_X2Y9_LUT4AB/S2BEGb[0] Tile_X2Y9_LUT4AB/S2BEGb[1] Tile_X2Y9_LUT4AB/S2BEGb[2]
+ Tile_X2Y9_LUT4AB/S2BEGb[3] Tile_X2Y9_LUT4AB/S2BEGb[4] Tile_X2Y9_LUT4AB/S2BEGb[5]
+ Tile_X2Y9_LUT4AB/S2BEGb[6] Tile_X2Y9_LUT4AB/S2BEGb[7] Tile_X2Y9_LUT4AB/S2BEG[0]
+ Tile_X2Y9_LUT4AB/S2BEG[1] Tile_X2Y9_LUT4AB/S2BEG[2] Tile_X2Y9_LUT4AB/S2BEG[3] Tile_X2Y9_LUT4AB/S2BEG[4]
+ Tile_X2Y9_LUT4AB/S2BEG[5] Tile_X2Y9_LUT4AB/S2BEG[6] Tile_X2Y9_LUT4AB/S2BEG[7] Tile_X2Y11_LUT4AB/S4END[0]
+ Tile_X2Y11_LUT4AB/S4END[10] Tile_X2Y11_LUT4AB/S4END[11] Tile_X2Y11_LUT4AB/S4END[12]
+ Tile_X2Y11_LUT4AB/S4END[13] Tile_X2Y11_LUT4AB/S4END[14] Tile_X2Y11_LUT4AB/S4END[15]
+ Tile_X2Y11_LUT4AB/S4END[1] Tile_X2Y11_LUT4AB/S4END[2] Tile_X2Y11_LUT4AB/S4END[3]
+ Tile_X2Y11_LUT4AB/S4END[4] Tile_X2Y11_LUT4AB/S4END[5] Tile_X2Y11_LUT4AB/S4END[6]
+ Tile_X2Y11_LUT4AB/S4END[7] Tile_X2Y11_LUT4AB/S4END[8] Tile_X2Y11_LUT4AB/S4END[9]
+ Tile_X2Y9_LUT4AB/S4BEG[0] Tile_X2Y9_LUT4AB/S4BEG[10] Tile_X2Y9_LUT4AB/S4BEG[11]
+ Tile_X2Y9_LUT4AB/S4BEG[12] Tile_X2Y9_LUT4AB/S4BEG[13] Tile_X2Y9_LUT4AB/S4BEG[14]
+ Tile_X2Y9_LUT4AB/S4BEG[15] Tile_X2Y9_LUT4AB/S4BEG[1] Tile_X2Y9_LUT4AB/S4BEG[2] Tile_X2Y9_LUT4AB/S4BEG[3]
+ Tile_X2Y9_LUT4AB/S4BEG[4] Tile_X2Y9_LUT4AB/S4BEG[5] Tile_X2Y9_LUT4AB/S4BEG[6] Tile_X2Y9_LUT4AB/S4BEG[7]
+ Tile_X2Y9_LUT4AB/S4BEG[8] Tile_X2Y9_LUT4AB/S4BEG[9] Tile_X2Y11_LUT4AB/SS4END[0]
+ Tile_X2Y11_LUT4AB/SS4END[10] Tile_X2Y11_LUT4AB/SS4END[11] Tile_X2Y11_LUT4AB/SS4END[12]
+ Tile_X2Y11_LUT4AB/SS4END[13] Tile_X2Y11_LUT4AB/SS4END[14] Tile_X2Y11_LUT4AB/SS4END[15]
+ Tile_X2Y11_LUT4AB/SS4END[1] Tile_X2Y11_LUT4AB/SS4END[2] Tile_X2Y11_LUT4AB/SS4END[3]
+ Tile_X2Y11_LUT4AB/SS4END[4] Tile_X2Y11_LUT4AB/SS4END[5] Tile_X2Y11_LUT4AB/SS4END[6]
+ Tile_X2Y11_LUT4AB/SS4END[7] Tile_X2Y11_LUT4AB/SS4END[8] Tile_X2Y11_LUT4AB/SS4END[9]
+ Tile_X2Y9_LUT4AB/SS4BEG[0] Tile_X2Y9_LUT4AB/SS4BEG[10] Tile_X2Y9_LUT4AB/SS4BEG[11]
+ Tile_X2Y9_LUT4AB/SS4BEG[12] Tile_X2Y9_LUT4AB/SS4BEG[13] Tile_X2Y9_LUT4AB/SS4BEG[14]
+ Tile_X2Y9_LUT4AB/SS4BEG[15] Tile_X2Y9_LUT4AB/SS4BEG[1] Tile_X2Y9_LUT4AB/SS4BEG[2]
+ Tile_X2Y9_LUT4AB/SS4BEG[3] Tile_X2Y9_LUT4AB/SS4BEG[4] Tile_X2Y9_LUT4AB/SS4BEG[5]
+ Tile_X2Y9_LUT4AB/SS4BEG[6] Tile_X2Y9_LUT4AB/SS4BEG[7] Tile_X2Y9_LUT4AB/SS4BEG[8]
+ Tile_X2Y9_LUT4AB/SS4BEG[9] Tile_X2Y10_LUT4AB/UserCLK Tile_X2Y9_LUT4AB/UserCLK VGND
+ VPWR Tile_X2Y10_LUT4AB/W1BEG[0] Tile_X2Y10_LUT4AB/W1BEG[1] Tile_X2Y10_LUT4AB/W1BEG[2]
+ Tile_X2Y10_LUT4AB/W1BEG[3] Tile_X3Y10_LUT4AB/W1BEG[0] Tile_X3Y10_LUT4AB/W1BEG[1]
+ Tile_X3Y10_LUT4AB/W1BEG[2] Tile_X3Y10_LUT4AB/W1BEG[3] Tile_X2Y10_LUT4AB/W2BEG[0]
+ Tile_X2Y10_LUT4AB/W2BEG[1] Tile_X2Y10_LUT4AB/W2BEG[2] Tile_X2Y10_LUT4AB/W2BEG[3]
+ Tile_X2Y10_LUT4AB/W2BEG[4] Tile_X2Y10_LUT4AB/W2BEG[5] Tile_X2Y10_LUT4AB/W2BEG[6]
+ Tile_X2Y10_LUT4AB/W2BEG[7] Tile_X1Y10_LUT4AB/W2END[0] Tile_X1Y10_LUT4AB/W2END[1]
+ Tile_X1Y10_LUT4AB/W2END[2] Tile_X1Y10_LUT4AB/W2END[3] Tile_X1Y10_LUT4AB/W2END[4]
+ Tile_X1Y10_LUT4AB/W2END[5] Tile_X1Y10_LUT4AB/W2END[6] Tile_X1Y10_LUT4AB/W2END[7]
+ Tile_X2Y10_LUT4AB/W2END[0] Tile_X2Y10_LUT4AB/W2END[1] Tile_X2Y10_LUT4AB/W2END[2]
+ Tile_X2Y10_LUT4AB/W2END[3] Tile_X2Y10_LUT4AB/W2END[4] Tile_X2Y10_LUT4AB/W2END[5]
+ Tile_X2Y10_LUT4AB/W2END[6] Tile_X2Y10_LUT4AB/W2END[7] Tile_X3Y10_LUT4AB/W2BEG[0]
+ Tile_X3Y10_LUT4AB/W2BEG[1] Tile_X3Y10_LUT4AB/W2BEG[2] Tile_X3Y10_LUT4AB/W2BEG[3]
+ Tile_X3Y10_LUT4AB/W2BEG[4] Tile_X3Y10_LUT4AB/W2BEG[5] Tile_X3Y10_LUT4AB/W2BEG[6]
+ Tile_X3Y10_LUT4AB/W2BEG[7] Tile_X2Y10_LUT4AB/W6BEG[0] Tile_X2Y10_LUT4AB/W6BEG[10]
+ Tile_X2Y10_LUT4AB/W6BEG[11] Tile_X2Y10_LUT4AB/W6BEG[1] Tile_X2Y10_LUT4AB/W6BEG[2]
+ Tile_X2Y10_LUT4AB/W6BEG[3] Tile_X2Y10_LUT4AB/W6BEG[4] Tile_X2Y10_LUT4AB/W6BEG[5]
+ Tile_X2Y10_LUT4AB/W6BEG[6] Tile_X2Y10_LUT4AB/W6BEG[7] Tile_X2Y10_LUT4AB/W6BEG[8]
+ Tile_X2Y10_LUT4AB/W6BEG[9] Tile_X3Y10_LUT4AB/W6BEG[0] Tile_X3Y10_LUT4AB/W6BEG[10]
+ Tile_X3Y10_LUT4AB/W6BEG[11] Tile_X3Y10_LUT4AB/W6BEG[1] Tile_X3Y10_LUT4AB/W6BEG[2]
+ Tile_X3Y10_LUT4AB/W6BEG[3] Tile_X3Y10_LUT4AB/W6BEG[4] Tile_X3Y10_LUT4AB/W6BEG[5]
+ Tile_X3Y10_LUT4AB/W6BEG[6] Tile_X3Y10_LUT4AB/W6BEG[7] Tile_X3Y10_LUT4AB/W6BEG[8]
+ Tile_X3Y10_LUT4AB/W6BEG[9] Tile_X2Y10_LUT4AB/WW4BEG[0] Tile_X2Y10_LUT4AB/WW4BEG[10]
+ Tile_X2Y10_LUT4AB/WW4BEG[11] Tile_X2Y10_LUT4AB/WW4BEG[12] Tile_X2Y10_LUT4AB/WW4BEG[13]
+ Tile_X2Y10_LUT4AB/WW4BEG[14] Tile_X2Y10_LUT4AB/WW4BEG[15] Tile_X2Y10_LUT4AB/WW4BEG[1]
+ Tile_X2Y10_LUT4AB/WW4BEG[2] Tile_X2Y10_LUT4AB/WW4BEG[3] Tile_X2Y10_LUT4AB/WW4BEG[4]
+ Tile_X2Y10_LUT4AB/WW4BEG[5] Tile_X2Y10_LUT4AB/WW4BEG[6] Tile_X2Y10_LUT4AB/WW4BEG[7]
+ Tile_X2Y10_LUT4AB/WW4BEG[8] Tile_X2Y10_LUT4AB/WW4BEG[9] Tile_X3Y10_LUT4AB/WW4BEG[0]
+ Tile_X3Y10_LUT4AB/WW4BEG[10] Tile_X3Y10_LUT4AB/WW4BEG[11] Tile_X3Y10_LUT4AB/WW4BEG[12]
+ Tile_X3Y10_LUT4AB/WW4BEG[13] Tile_X3Y10_LUT4AB/WW4BEG[14] Tile_X3Y10_LUT4AB/WW4BEG[15]
+ Tile_X3Y10_LUT4AB/WW4BEG[1] Tile_X3Y10_LUT4AB/WW4BEG[2] Tile_X3Y10_LUT4AB/WW4BEG[3]
+ Tile_X3Y10_LUT4AB/WW4BEG[4] Tile_X3Y10_LUT4AB/WW4BEG[5] Tile_X3Y10_LUT4AB/WW4BEG[6]
+ Tile_X3Y10_LUT4AB/WW4BEG[7] Tile_X3Y10_LUT4AB/WW4BEG[8] Tile_X3Y10_LUT4AB/WW4BEG[9]
+ LUT4AB
XTile_X8Y7_LUT4AB Tile_X8Y8_LUT4AB/Co Tile_X8Y7_LUT4AB/Co Tile_X9Y7_LUT4AB/E1END[0]
+ Tile_X9Y7_LUT4AB/E1END[1] Tile_X9Y7_LUT4AB/E1END[2] Tile_X9Y7_LUT4AB/E1END[3] Tile_X8Y7_LUT4AB/E1END[0]
+ Tile_X8Y7_LUT4AB/E1END[1] Tile_X8Y7_LUT4AB/E1END[2] Tile_X8Y7_LUT4AB/E1END[3] Tile_X9Y7_LUT4AB/E2MID[0]
+ Tile_X9Y7_LUT4AB/E2MID[1] Tile_X9Y7_LUT4AB/E2MID[2] Tile_X9Y7_LUT4AB/E2MID[3] Tile_X9Y7_LUT4AB/E2MID[4]
+ Tile_X9Y7_LUT4AB/E2MID[5] Tile_X9Y7_LUT4AB/E2MID[6] Tile_X9Y7_LUT4AB/E2MID[7] Tile_X9Y7_LUT4AB/E2END[0]
+ Tile_X9Y7_LUT4AB/E2END[1] Tile_X9Y7_LUT4AB/E2END[2] Tile_X9Y7_LUT4AB/E2END[3] Tile_X9Y7_LUT4AB/E2END[4]
+ Tile_X9Y7_LUT4AB/E2END[5] Tile_X9Y7_LUT4AB/E2END[6] Tile_X9Y7_LUT4AB/E2END[7] Tile_X8Y7_LUT4AB/E2END[0]
+ Tile_X8Y7_LUT4AB/E2END[1] Tile_X8Y7_LUT4AB/E2END[2] Tile_X8Y7_LUT4AB/E2END[3] Tile_X8Y7_LUT4AB/E2END[4]
+ Tile_X8Y7_LUT4AB/E2END[5] Tile_X8Y7_LUT4AB/E2END[6] Tile_X8Y7_LUT4AB/E2END[7] Tile_X8Y7_LUT4AB/E2MID[0]
+ Tile_X8Y7_LUT4AB/E2MID[1] Tile_X8Y7_LUT4AB/E2MID[2] Tile_X8Y7_LUT4AB/E2MID[3] Tile_X8Y7_LUT4AB/E2MID[4]
+ Tile_X8Y7_LUT4AB/E2MID[5] Tile_X8Y7_LUT4AB/E2MID[6] Tile_X8Y7_LUT4AB/E2MID[7] Tile_X9Y7_LUT4AB/E6END[0]
+ Tile_X9Y7_LUT4AB/E6END[10] Tile_X9Y7_LUT4AB/E6END[11] Tile_X9Y7_LUT4AB/E6END[1]
+ Tile_X9Y7_LUT4AB/E6END[2] Tile_X9Y7_LUT4AB/E6END[3] Tile_X9Y7_LUT4AB/E6END[4] Tile_X9Y7_LUT4AB/E6END[5]
+ Tile_X9Y7_LUT4AB/E6END[6] Tile_X9Y7_LUT4AB/E6END[7] Tile_X9Y7_LUT4AB/E6END[8] Tile_X9Y7_LUT4AB/E6END[9]
+ Tile_X8Y7_LUT4AB/E6END[0] Tile_X8Y7_LUT4AB/E6END[10] Tile_X8Y7_LUT4AB/E6END[11]
+ Tile_X8Y7_LUT4AB/E6END[1] Tile_X8Y7_LUT4AB/E6END[2] Tile_X8Y7_LUT4AB/E6END[3] Tile_X8Y7_LUT4AB/E6END[4]
+ Tile_X8Y7_LUT4AB/E6END[5] Tile_X8Y7_LUT4AB/E6END[6] Tile_X8Y7_LUT4AB/E6END[7] Tile_X8Y7_LUT4AB/E6END[8]
+ Tile_X8Y7_LUT4AB/E6END[9] Tile_X9Y7_LUT4AB/EE4END[0] Tile_X9Y7_LUT4AB/EE4END[10]
+ Tile_X9Y7_LUT4AB/EE4END[11] Tile_X9Y7_LUT4AB/EE4END[12] Tile_X9Y7_LUT4AB/EE4END[13]
+ Tile_X9Y7_LUT4AB/EE4END[14] Tile_X9Y7_LUT4AB/EE4END[15] Tile_X9Y7_LUT4AB/EE4END[1]
+ Tile_X9Y7_LUT4AB/EE4END[2] Tile_X9Y7_LUT4AB/EE4END[3] Tile_X9Y7_LUT4AB/EE4END[4]
+ Tile_X9Y7_LUT4AB/EE4END[5] Tile_X9Y7_LUT4AB/EE4END[6] Tile_X9Y7_LUT4AB/EE4END[7]
+ Tile_X9Y7_LUT4AB/EE4END[8] Tile_X9Y7_LUT4AB/EE4END[9] Tile_X8Y7_LUT4AB/EE4END[0]
+ Tile_X8Y7_LUT4AB/EE4END[10] Tile_X8Y7_LUT4AB/EE4END[11] Tile_X8Y7_LUT4AB/EE4END[12]
+ Tile_X8Y7_LUT4AB/EE4END[13] Tile_X8Y7_LUT4AB/EE4END[14] Tile_X8Y7_LUT4AB/EE4END[15]
+ Tile_X8Y7_LUT4AB/EE4END[1] Tile_X8Y7_LUT4AB/EE4END[2] Tile_X8Y7_LUT4AB/EE4END[3]
+ Tile_X8Y7_LUT4AB/EE4END[4] Tile_X8Y7_LUT4AB/EE4END[5] Tile_X8Y7_LUT4AB/EE4END[6]
+ Tile_X8Y7_LUT4AB/EE4END[7] Tile_X8Y7_LUT4AB/EE4END[8] Tile_X8Y7_LUT4AB/EE4END[9]
+ Tile_X8Y7_LUT4AB/FrameData[0] Tile_X8Y7_LUT4AB/FrameData[10] Tile_X8Y7_LUT4AB/FrameData[11]
+ Tile_X8Y7_LUT4AB/FrameData[12] Tile_X8Y7_LUT4AB/FrameData[13] Tile_X8Y7_LUT4AB/FrameData[14]
+ Tile_X8Y7_LUT4AB/FrameData[15] Tile_X8Y7_LUT4AB/FrameData[16] Tile_X8Y7_LUT4AB/FrameData[17]
+ Tile_X8Y7_LUT4AB/FrameData[18] Tile_X8Y7_LUT4AB/FrameData[19] Tile_X8Y7_LUT4AB/FrameData[1]
+ Tile_X8Y7_LUT4AB/FrameData[20] Tile_X8Y7_LUT4AB/FrameData[21] Tile_X8Y7_LUT4AB/FrameData[22]
+ Tile_X8Y7_LUT4AB/FrameData[23] Tile_X8Y7_LUT4AB/FrameData[24] Tile_X8Y7_LUT4AB/FrameData[25]
+ Tile_X8Y7_LUT4AB/FrameData[26] Tile_X8Y7_LUT4AB/FrameData[27] Tile_X8Y7_LUT4AB/FrameData[28]
+ Tile_X8Y7_LUT4AB/FrameData[29] Tile_X8Y7_LUT4AB/FrameData[2] Tile_X8Y7_LUT4AB/FrameData[30]
+ Tile_X8Y7_LUT4AB/FrameData[31] Tile_X8Y7_LUT4AB/FrameData[3] Tile_X8Y7_LUT4AB/FrameData[4]
+ Tile_X8Y7_LUT4AB/FrameData[5] Tile_X8Y7_LUT4AB/FrameData[6] Tile_X8Y7_LUT4AB/FrameData[7]
+ Tile_X8Y7_LUT4AB/FrameData[8] Tile_X8Y7_LUT4AB/FrameData[9] Tile_X9Y7_LUT4AB/FrameData[0]
+ Tile_X9Y7_LUT4AB/FrameData[10] Tile_X9Y7_LUT4AB/FrameData[11] Tile_X9Y7_LUT4AB/FrameData[12]
+ Tile_X9Y7_LUT4AB/FrameData[13] Tile_X9Y7_LUT4AB/FrameData[14] Tile_X9Y7_LUT4AB/FrameData[15]
+ Tile_X9Y7_LUT4AB/FrameData[16] Tile_X9Y7_LUT4AB/FrameData[17] Tile_X9Y7_LUT4AB/FrameData[18]
+ Tile_X9Y7_LUT4AB/FrameData[19] Tile_X9Y7_LUT4AB/FrameData[1] Tile_X9Y7_LUT4AB/FrameData[20]
+ Tile_X9Y7_LUT4AB/FrameData[21] Tile_X9Y7_LUT4AB/FrameData[22] Tile_X9Y7_LUT4AB/FrameData[23]
+ Tile_X9Y7_LUT4AB/FrameData[24] Tile_X9Y7_LUT4AB/FrameData[25] Tile_X9Y7_LUT4AB/FrameData[26]
+ Tile_X9Y7_LUT4AB/FrameData[27] Tile_X9Y7_LUT4AB/FrameData[28] Tile_X9Y7_LUT4AB/FrameData[29]
+ Tile_X9Y7_LUT4AB/FrameData[2] Tile_X9Y7_LUT4AB/FrameData[30] Tile_X9Y7_LUT4AB/FrameData[31]
+ Tile_X9Y7_LUT4AB/FrameData[3] Tile_X9Y7_LUT4AB/FrameData[4] Tile_X9Y7_LUT4AB/FrameData[5]
+ Tile_X9Y7_LUT4AB/FrameData[6] Tile_X9Y7_LUT4AB/FrameData[7] Tile_X9Y7_LUT4AB/FrameData[8]
+ Tile_X9Y7_LUT4AB/FrameData[9] Tile_X8Y7_LUT4AB/FrameStrobe[0] Tile_X8Y7_LUT4AB/FrameStrobe[10]
+ Tile_X8Y7_LUT4AB/FrameStrobe[11] Tile_X8Y7_LUT4AB/FrameStrobe[12] Tile_X8Y7_LUT4AB/FrameStrobe[13]
+ Tile_X8Y7_LUT4AB/FrameStrobe[14] Tile_X8Y7_LUT4AB/FrameStrobe[15] Tile_X8Y7_LUT4AB/FrameStrobe[16]
+ Tile_X8Y7_LUT4AB/FrameStrobe[17] Tile_X8Y7_LUT4AB/FrameStrobe[18] Tile_X8Y7_LUT4AB/FrameStrobe[19]
+ Tile_X8Y7_LUT4AB/FrameStrobe[1] Tile_X8Y7_LUT4AB/FrameStrobe[2] Tile_X8Y7_LUT4AB/FrameStrobe[3]
+ Tile_X8Y7_LUT4AB/FrameStrobe[4] Tile_X8Y7_LUT4AB/FrameStrobe[5] Tile_X8Y7_LUT4AB/FrameStrobe[6]
+ Tile_X8Y7_LUT4AB/FrameStrobe[7] Tile_X8Y7_LUT4AB/FrameStrobe[8] Tile_X8Y7_LUT4AB/FrameStrobe[9]
+ Tile_X8Y6_LUT4AB/FrameStrobe[0] Tile_X8Y6_LUT4AB/FrameStrobe[10] Tile_X8Y6_LUT4AB/FrameStrobe[11]
+ Tile_X8Y6_LUT4AB/FrameStrobe[12] Tile_X8Y6_LUT4AB/FrameStrobe[13] Tile_X8Y6_LUT4AB/FrameStrobe[14]
+ Tile_X8Y6_LUT4AB/FrameStrobe[15] Tile_X8Y6_LUT4AB/FrameStrobe[16] Tile_X8Y6_LUT4AB/FrameStrobe[17]
+ Tile_X8Y6_LUT4AB/FrameStrobe[18] Tile_X8Y6_LUT4AB/FrameStrobe[19] Tile_X8Y6_LUT4AB/FrameStrobe[1]
+ Tile_X8Y6_LUT4AB/FrameStrobe[2] Tile_X8Y6_LUT4AB/FrameStrobe[3] Tile_X8Y6_LUT4AB/FrameStrobe[4]
+ Tile_X8Y6_LUT4AB/FrameStrobe[5] Tile_X8Y6_LUT4AB/FrameStrobe[6] Tile_X8Y6_LUT4AB/FrameStrobe[7]
+ Tile_X8Y6_LUT4AB/FrameStrobe[8] Tile_X8Y6_LUT4AB/FrameStrobe[9] Tile_X8Y7_LUT4AB/N1BEG[0]
+ Tile_X8Y7_LUT4AB/N1BEG[1] Tile_X8Y7_LUT4AB/N1BEG[2] Tile_X8Y7_LUT4AB/N1BEG[3] Tile_X8Y8_LUT4AB/N1BEG[0]
+ Tile_X8Y8_LUT4AB/N1BEG[1] Tile_X8Y8_LUT4AB/N1BEG[2] Tile_X8Y8_LUT4AB/N1BEG[3] Tile_X8Y7_LUT4AB/N2BEG[0]
+ Tile_X8Y7_LUT4AB/N2BEG[1] Tile_X8Y7_LUT4AB/N2BEG[2] Tile_X8Y7_LUT4AB/N2BEG[3] Tile_X8Y7_LUT4AB/N2BEG[4]
+ Tile_X8Y7_LUT4AB/N2BEG[5] Tile_X8Y7_LUT4AB/N2BEG[6] Tile_X8Y7_LUT4AB/N2BEG[7] Tile_X8Y6_LUT4AB/N2END[0]
+ Tile_X8Y6_LUT4AB/N2END[1] Tile_X8Y6_LUT4AB/N2END[2] Tile_X8Y6_LUT4AB/N2END[3] Tile_X8Y6_LUT4AB/N2END[4]
+ Tile_X8Y6_LUT4AB/N2END[5] Tile_X8Y6_LUT4AB/N2END[6] Tile_X8Y6_LUT4AB/N2END[7] Tile_X8Y7_LUT4AB/N2END[0]
+ Tile_X8Y7_LUT4AB/N2END[1] Tile_X8Y7_LUT4AB/N2END[2] Tile_X8Y7_LUT4AB/N2END[3] Tile_X8Y7_LUT4AB/N2END[4]
+ Tile_X8Y7_LUT4AB/N2END[5] Tile_X8Y7_LUT4AB/N2END[6] Tile_X8Y7_LUT4AB/N2END[7] Tile_X8Y8_LUT4AB/N2BEG[0]
+ Tile_X8Y8_LUT4AB/N2BEG[1] Tile_X8Y8_LUT4AB/N2BEG[2] Tile_X8Y8_LUT4AB/N2BEG[3] Tile_X8Y8_LUT4AB/N2BEG[4]
+ Tile_X8Y8_LUT4AB/N2BEG[5] Tile_X8Y8_LUT4AB/N2BEG[6] Tile_X8Y8_LUT4AB/N2BEG[7] Tile_X8Y7_LUT4AB/N4BEG[0]
+ Tile_X8Y7_LUT4AB/N4BEG[10] Tile_X8Y7_LUT4AB/N4BEG[11] Tile_X8Y7_LUT4AB/N4BEG[12]
+ Tile_X8Y7_LUT4AB/N4BEG[13] Tile_X8Y7_LUT4AB/N4BEG[14] Tile_X8Y7_LUT4AB/N4BEG[15]
+ Tile_X8Y7_LUT4AB/N4BEG[1] Tile_X8Y7_LUT4AB/N4BEG[2] Tile_X8Y7_LUT4AB/N4BEG[3] Tile_X8Y7_LUT4AB/N4BEG[4]
+ Tile_X8Y7_LUT4AB/N4BEG[5] Tile_X8Y7_LUT4AB/N4BEG[6] Tile_X8Y7_LUT4AB/N4BEG[7] Tile_X8Y7_LUT4AB/N4BEG[8]
+ Tile_X8Y7_LUT4AB/N4BEG[9] Tile_X8Y8_LUT4AB/N4BEG[0] Tile_X8Y8_LUT4AB/N4BEG[10] Tile_X8Y8_LUT4AB/N4BEG[11]
+ Tile_X8Y8_LUT4AB/N4BEG[12] Tile_X8Y8_LUT4AB/N4BEG[13] Tile_X8Y8_LUT4AB/N4BEG[14]
+ Tile_X8Y8_LUT4AB/N4BEG[15] Tile_X8Y8_LUT4AB/N4BEG[1] Tile_X8Y8_LUT4AB/N4BEG[2] Tile_X8Y8_LUT4AB/N4BEG[3]
+ Tile_X8Y8_LUT4AB/N4BEG[4] Tile_X8Y8_LUT4AB/N4BEG[5] Tile_X8Y8_LUT4AB/N4BEG[6] Tile_X8Y8_LUT4AB/N4BEG[7]
+ Tile_X8Y8_LUT4AB/N4BEG[8] Tile_X8Y8_LUT4AB/N4BEG[9] Tile_X8Y7_LUT4AB/NN4BEG[0] Tile_X8Y7_LUT4AB/NN4BEG[10]
+ Tile_X8Y7_LUT4AB/NN4BEG[11] Tile_X8Y7_LUT4AB/NN4BEG[12] Tile_X8Y7_LUT4AB/NN4BEG[13]
+ Tile_X8Y7_LUT4AB/NN4BEG[14] Tile_X8Y7_LUT4AB/NN4BEG[15] Tile_X8Y7_LUT4AB/NN4BEG[1]
+ Tile_X8Y7_LUT4AB/NN4BEG[2] Tile_X8Y7_LUT4AB/NN4BEG[3] Tile_X8Y7_LUT4AB/NN4BEG[4]
+ Tile_X8Y7_LUT4AB/NN4BEG[5] Tile_X8Y7_LUT4AB/NN4BEG[6] Tile_X8Y7_LUT4AB/NN4BEG[7]
+ Tile_X8Y7_LUT4AB/NN4BEG[8] Tile_X8Y7_LUT4AB/NN4BEG[9] Tile_X8Y8_LUT4AB/NN4BEG[0]
+ Tile_X8Y8_LUT4AB/NN4BEG[10] Tile_X8Y8_LUT4AB/NN4BEG[11] Tile_X8Y8_LUT4AB/NN4BEG[12]
+ Tile_X8Y8_LUT4AB/NN4BEG[13] Tile_X8Y8_LUT4AB/NN4BEG[14] Tile_X8Y8_LUT4AB/NN4BEG[15]
+ Tile_X8Y8_LUT4AB/NN4BEG[1] Tile_X8Y8_LUT4AB/NN4BEG[2] Tile_X8Y8_LUT4AB/NN4BEG[3]
+ Tile_X8Y8_LUT4AB/NN4BEG[4] Tile_X8Y8_LUT4AB/NN4BEG[5] Tile_X8Y8_LUT4AB/NN4BEG[6]
+ Tile_X8Y8_LUT4AB/NN4BEG[7] Tile_X8Y8_LUT4AB/NN4BEG[8] Tile_X8Y8_LUT4AB/NN4BEG[9]
+ Tile_X8Y8_LUT4AB/S1END[0] Tile_X8Y8_LUT4AB/S1END[1] Tile_X8Y8_LUT4AB/S1END[2] Tile_X8Y8_LUT4AB/S1END[3]
+ Tile_X8Y7_LUT4AB/S1END[0] Tile_X8Y7_LUT4AB/S1END[1] Tile_X8Y7_LUT4AB/S1END[2] Tile_X8Y7_LUT4AB/S1END[3]
+ Tile_X8Y8_LUT4AB/S2MID[0] Tile_X8Y8_LUT4AB/S2MID[1] Tile_X8Y8_LUT4AB/S2MID[2] Tile_X8Y8_LUT4AB/S2MID[3]
+ Tile_X8Y8_LUT4AB/S2MID[4] Tile_X8Y8_LUT4AB/S2MID[5] Tile_X8Y8_LUT4AB/S2MID[6] Tile_X8Y8_LUT4AB/S2MID[7]
+ Tile_X8Y8_LUT4AB/S2END[0] Tile_X8Y8_LUT4AB/S2END[1] Tile_X8Y8_LUT4AB/S2END[2] Tile_X8Y8_LUT4AB/S2END[3]
+ Tile_X8Y8_LUT4AB/S2END[4] Tile_X8Y8_LUT4AB/S2END[5] Tile_X8Y8_LUT4AB/S2END[6] Tile_X8Y8_LUT4AB/S2END[7]
+ Tile_X8Y7_LUT4AB/S2END[0] Tile_X8Y7_LUT4AB/S2END[1] Tile_X8Y7_LUT4AB/S2END[2] Tile_X8Y7_LUT4AB/S2END[3]
+ Tile_X8Y7_LUT4AB/S2END[4] Tile_X8Y7_LUT4AB/S2END[5] Tile_X8Y7_LUT4AB/S2END[6] Tile_X8Y7_LUT4AB/S2END[7]
+ Tile_X8Y7_LUT4AB/S2MID[0] Tile_X8Y7_LUT4AB/S2MID[1] Tile_X8Y7_LUT4AB/S2MID[2] Tile_X8Y7_LUT4AB/S2MID[3]
+ Tile_X8Y7_LUT4AB/S2MID[4] Tile_X8Y7_LUT4AB/S2MID[5] Tile_X8Y7_LUT4AB/S2MID[6] Tile_X8Y7_LUT4AB/S2MID[7]
+ Tile_X8Y8_LUT4AB/S4END[0] Tile_X8Y8_LUT4AB/S4END[10] Tile_X8Y8_LUT4AB/S4END[11]
+ Tile_X8Y8_LUT4AB/S4END[12] Tile_X8Y8_LUT4AB/S4END[13] Tile_X8Y8_LUT4AB/S4END[14]
+ Tile_X8Y8_LUT4AB/S4END[15] Tile_X8Y8_LUT4AB/S4END[1] Tile_X8Y8_LUT4AB/S4END[2] Tile_X8Y8_LUT4AB/S4END[3]
+ Tile_X8Y8_LUT4AB/S4END[4] Tile_X8Y8_LUT4AB/S4END[5] Tile_X8Y8_LUT4AB/S4END[6] Tile_X8Y8_LUT4AB/S4END[7]
+ Tile_X8Y8_LUT4AB/S4END[8] Tile_X8Y8_LUT4AB/S4END[9] Tile_X8Y7_LUT4AB/S4END[0] Tile_X8Y7_LUT4AB/S4END[10]
+ Tile_X8Y7_LUT4AB/S4END[11] Tile_X8Y7_LUT4AB/S4END[12] Tile_X8Y7_LUT4AB/S4END[13]
+ Tile_X8Y7_LUT4AB/S4END[14] Tile_X8Y7_LUT4AB/S4END[15] Tile_X8Y7_LUT4AB/S4END[1]
+ Tile_X8Y7_LUT4AB/S4END[2] Tile_X8Y7_LUT4AB/S4END[3] Tile_X8Y7_LUT4AB/S4END[4] Tile_X8Y7_LUT4AB/S4END[5]
+ Tile_X8Y7_LUT4AB/S4END[6] Tile_X8Y7_LUT4AB/S4END[7] Tile_X8Y7_LUT4AB/S4END[8] Tile_X8Y7_LUT4AB/S4END[9]
+ Tile_X8Y8_LUT4AB/SS4END[0] Tile_X8Y8_LUT4AB/SS4END[10] Tile_X8Y8_LUT4AB/SS4END[11]
+ Tile_X8Y8_LUT4AB/SS4END[12] Tile_X8Y8_LUT4AB/SS4END[13] Tile_X8Y8_LUT4AB/SS4END[14]
+ Tile_X8Y8_LUT4AB/SS4END[15] Tile_X8Y8_LUT4AB/SS4END[1] Tile_X8Y8_LUT4AB/SS4END[2]
+ Tile_X8Y8_LUT4AB/SS4END[3] Tile_X8Y8_LUT4AB/SS4END[4] Tile_X8Y8_LUT4AB/SS4END[5]
+ Tile_X8Y8_LUT4AB/SS4END[6] Tile_X8Y8_LUT4AB/SS4END[7] Tile_X8Y8_LUT4AB/SS4END[8]
+ Tile_X8Y8_LUT4AB/SS4END[9] Tile_X8Y7_LUT4AB/SS4END[0] Tile_X8Y7_LUT4AB/SS4END[10]
+ Tile_X8Y7_LUT4AB/SS4END[11] Tile_X8Y7_LUT4AB/SS4END[12] Tile_X8Y7_LUT4AB/SS4END[13]
+ Tile_X8Y7_LUT4AB/SS4END[14] Tile_X8Y7_LUT4AB/SS4END[15] Tile_X8Y7_LUT4AB/SS4END[1]
+ Tile_X8Y7_LUT4AB/SS4END[2] Tile_X8Y7_LUT4AB/SS4END[3] Tile_X8Y7_LUT4AB/SS4END[4]
+ Tile_X8Y7_LUT4AB/SS4END[5] Tile_X8Y7_LUT4AB/SS4END[6] Tile_X8Y7_LUT4AB/SS4END[7]
+ Tile_X8Y7_LUT4AB/SS4END[8] Tile_X8Y7_LUT4AB/SS4END[9] Tile_X8Y7_LUT4AB/UserCLK Tile_X8Y6_LUT4AB/UserCLK
+ VGND VPWR Tile_X8Y7_LUT4AB/W1BEG[0] Tile_X8Y7_LUT4AB/W1BEG[1] Tile_X8Y7_LUT4AB/W1BEG[2]
+ Tile_X8Y7_LUT4AB/W1BEG[3] Tile_X9Y7_LUT4AB/W1BEG[0] Tile_X9Y7_LUT4AB/W1BEG[1] Tile_X9Y7_LUT4AB/W1BEG[2]
+ Tile_X9Y7_LUT4AB/W1BEG[3] Tile_X8Y7_LUT4AB/W2BEG[0] Tile_X8Y7_LUT4AB/W2BEG[1] Tile_X8Y7_LUT4AB/W2BEG[2]
+ Tile_X8Y7_LUT4AB/W2BEG[3] Tile_X8Y7_LUT4AB/W2BEG[4] Tile_X8Y7_LUT4AB/W2BEG[5] Tile_X8Y7_LUT4AB/W2BEG[6]
+ Tile_X8Y7_LUT4AB/W2BEG[7] Tile_X8Y7_LUT4AB/W2BEGb[0] Tile_X8Y7_LUT4AB/W2BEGb[1]
+ Tile_X8Y7_LUT4AB/W2BEGb[2] Tile_X8Y7_LUT4AB/W2BEGb[3] Tile_X8Y7_LUT4AB/W2BEGb[4]
+ Tile_X8Y7_LUT4AB/W2BEGb[5] Tile_X8Y7_LUT4AB/W2BEGb[6] Tile_X8Y7_LUT4AB/W2BEGb[7]
+ Tile_X8Y7_LUT4AB/W2END[0] Tile_X8Y7_LUT4AB/W2END[1] Tile_X8Y7_LUT4AB/W2END[2] Tile_X8Y7_LUT4AB/W2END[3]
+ Tile_X8Y7_LUT4AB/W2END[4] Tile_X8Y7_LUT4AB/W2END[5] Tile_X8Y7_LUT4AB/W2END[6] Tile_X8Y7_LUT4AB/W2END[7]
+ Tile_X9Y7_LUT4AB/W2BEG[0] Tile_X9Y7_LUT4AB/W2BEG[1] Tile_X9Y7_LUT4AB/W2BEG[2] Tile_X9Y7_LUT4AB/W2BEG[3]
+ Tile_X9Y7_LUT4AB/W2BEG[4] Tile_X9Y7_LUT4AB/W2BEG[5] Tile_X9Y7_LUT4AB/W2BEG[6] Tile_X9Y7_LUT4AB/W2BEG[7]
+ Tile_X8Y7_LUT4AB/W6BEG[0] Tile_X8Y7_LUT4AB/W6BEG[10] Tile_X8Y7_LUT4AB/W6BEG[11]
+ Tile_X8Y7_LUT4AB/W6BEG[1] Tile_X8Y7_LUT4AB/W6BEG[2] Tile_X8Y7_LUT4AB/W6BEG[3] Tile_X8Y7_LUT4AB/W6BEG[4]
+ Tile_X8Y7_LUT4AB/W6BEG[5] Tile_X8Y7_LUT4AB/W6BEG[6] Tile_X8Y7_LUT4AB/W6BEG[7] Tile_X8Y7_LUT4AB/W6BEG[8]
+ Tile_X8Y7_LUT4AB/W6BEG[9] Tile_X9Y7_LUT4AB/W6BEG[0] Tile_X9Y7_LUT4AB/W6BEG[10] Tile_X9Y7_LUT4AB/W6BEG[11]
+ Tile_X9Y7_LUT4AB/W6BEG[1] Tile_X9Y7_LUT4AB/W6BEG[2] Tile_X9Y7_LUT4AB/W6BEG[3] Tile_X9Y7_LUT4AB/W6BEG[4]
+ Tile_X9Y7_LUT4AB/W6BEG[5] Tile_X9Y7_LUT4AB/W6BEG[6] Tile_X9Y7_LUT4AB/W6BEG[7] Tile_X9Y7_LUT4AB/W6BEG[8]
+ Tile_X9Y7_LUT4AB/W6BEG[9] Tile_X8Y7_LUT4AB/WW4BEG[0] Tile_X8Y7_LUT4AB/WW4BEG[10]
+ Tile_X8Y7_LUT4AB/WW4BEG[11] Tile_X8Y7_LUT4AB/WW4BEG[12] Tile_X8Y7_LUT4AB/WW4BEG[13]
+ Tile_X8Y7_LUT4AB/WW4BEG[14] Tile_X8Y7_LUT4AB/WW4BEG[15] Tile_X8Y7_LUT4AB/WW4BEG[1]
+ Tile_X8Y7_LUT4AB/WW4BEG[2] Tile_X8Y7_LUT4AB/WW4BEG[3] Tile_X8Y7_LUT4AB/WW4BEG[4]
+ Tile_X8Y7_LUT4AB/WW4BEG[5] Tile_X8Y7_LUT4AB/WW4BEG[6] Tile_X8Y7_LUT4AB/WW4BEG[7]
+ Tile_X8Y7_LUT4AB/WW4BEG[8] Tile_X8Y7_LUT4AB/WW4BEG[9] Tile_X9Y7_LUT4AB/WW4BEG[0]
+ Tile_X9Y7_LUT4AB/WW4BEG[10] Tile_X9Y7_LUT4AB/WW4BEG[11] Tile_X9Y7_LUT4AB/WW4BEG[12]
+ Tile_X9Y7_LUT4AB/WW4BEG[13] Tile_X9Y7_LUT4AB/WW4BEG[14] Tile_X9Y7_LUT4AB/WW4BEG[15]
+ Tile_X9Y7_LUT4AB/WW4BEG[1] Tile_X9Y7_LUT4AB/WW4BEG[2] Tile_X9Y7_LUT4AB/WW4BEG[3]
+ Tile_X9Y7_LUT4AB/WW4BEG[4] Tile_X9Y7_LUT4AB/WW4BEG[5] Tile_X9Y7_LUT4AB/WW4BEG[6]
+ Tile_X9Y7_LUT4AB/WW4BEG[7] Tile_X9Y7_LUT4AB/WW4BEG[8] Tile_X9Y7_LUT4AB/WW4BEG[9]
+ LUT4AB
XTile_X5Y2_LUT4AB Tile_X5Y3_LUT4AB/Co Tile_X5Y2_LUT4AB/Co Tile_X6Y2_LUT4AB/E1END[0]
+ Tile_X6Y2_LUT4AB/E1END[1] Tile_X6Y2_LUT4AB/E1END[2] Tile_X6Y2_LUT4AB/E1END[3] Tile_X5Y2_LUT4AB/E1END[0]
+ Tile_X5Y2_LUT4AB/E1END[1] Tile_X5Y2_LUT4AB/E1END[2] Tile_X5Y2_LUT4AB/E1END[3] Tile_X6Y2_LUT4AB/E2MID[0]
+ Tile_X6Y2_LUT4AB/E2MID[1] Tile_X6Y2_LUT4AB/E2MID[2] Tile_X6Y2_LUT4AB/E2MID[3] Tile_X6Y2_LUT4AB/E2MID[4]
+ Tile_X6Y2_LUT4AB/E2MID[5] Tile_X6Y2_LUT4AB/E2MID[6] Tile_X6Y2_LUT4AB/E2MID[7] Tile_X6Y2_LUT4AB/E2END[0]
+ Tile_X6Y2_LUT4AB/E2END[1] Tile_X6Y2_LUT4AB/E2END[2] Tile_X6Y2_LUT4AB/E2END[3] Tile_X6Y2_LUT4AB/E2END[4]
+ Tile_X6Y2_LUT4AB/E2END[5] Tile_X6Y2_LUT4AB/E2END[6] Tile_X6Y2_LUT4AB/E2END[7] Tile_X5Y2_LUT4AB/E2END[0]
+ Tile_X5Y2_LUT4AB/E2END[1] Tile_X5Y2_LUT4AB/E2END[2] Tile_X5Y2_LUT4AB/E2END[3] Tile_X5Y2_LUT4AB/E2END[4]
+ Tile_X5Y2_LUT4AB/E2END[5] Tile_X5Y2_LUT4AB/E2END[6] Tile_X5Y2_LUT4AB/E2END[7] Tile_X5Y2_LUT4AB/E2MID[0]
+ Tile_X5Y2_LUT4AB/E2MID[1] Tile_X5Y2_LUT4AB/E2MID[2] Tile_X5Y2_LUT4AB/E2MID[3] Tile_X5Y2_LUT4AB/E2MID[4]
+ Tile_X5Y2_LUT4AB/E2MID[5] Tile_X5Y2_LUT4AB/E2MID[6] Tile_X5Y2_LUT4AB/E2MID[7] Tile_X6Y2_LUT4AB/E6END[0]
+ Tile_X6Y2_LUT4AB/E6END[10] Tile_X6Y2_LUT4AB/E6END[11] Tile_X6Y2_LUT4AB/E6END[1]
+ Tile_X6Y2_LUT4AB/E6END[2] Tile_X6Y2_LUT4AB/E6END[3] Tile_X6Y2_LUT4AB/E6END[4] Tile_X6Y2_LUT4AB/E6END[5]
+ Tile_X6Y2_LUT4AB/E6END[6] Tile_X6Y2_LUT4AB/E6END[7] Tile_X6Y2_LUT4AB/E6END[8] Tile_X6Y2_LUT4AB/E6END[9]
+ Tile_X5Y2_LUT4AB/E6END[0] Tile_X5Y2_LUT4AB/E6END[10] Tile_X5Y2_LUT4AB/E6END[11]
+ Tile_X5Y2_LUT4AB/E6END[1] Tile_X5Y2_LUT4AB/E6END[2] Tile_X5Y2_LUT4AB/E6END[3] Tile_X5Y2_LUT4AB/E6END[4]
+ Tile_X5Y2_LUT4AB/E6END[5] Tile_X5Y2_LUT4AB/E6END[6] Tile_X5Y2_LUT4AB/E6END[7] Tile_X5Y2_LUT4AB/E6END[8]
+ Tile_X5Y2_LUT4AB/E6END[9] Tile_X6Y2_LUT4AB/EE4END[0] Tile_X6Y2_LUT4AB/EE4END[10]
+ Tile_X6Y2_LUT4AB/EE4END[11] Tile_X6Y2_LUT4AB/EE4END[12] Tile_X6Y2_LUT4AB/EE4END[13]
+ Tile_X6Y2_LUT4AB/EE4END[14] Tile_X6Y2_LUT4AB/EE4END[15] Tile_X6Y2_LUT4AB/EE4END[1]
+ Tile_X6Y2_LUT4AB/EE4END[2] Tile_X6Y2_LUT4AB/EE4END[3] Tile_X6Y2_LUT4AB/EE4END[4]
+ Tile_X6Y2_LUT4AB/EE4END[5] Tile_X6Y2_LUT4AB/EE4END[6] Tile_X6Y2_LUT4AB/EE4END[7]
+ Tile_X6Y2_LUT4AB/EE4END[8] Tile_X6Y2_LUT4AB/EE4END[9] Tile_X5Y2_LUT4AB/EE4END[0]
+ Tile_X5Y2_LUT4AB/EE4END[10] Tile_X5Y2_LUT4AB/EE4END[11] Tile_X5Y2_LUT4AB/EE4END[12]
+ Tile_X5Y2_LUT4AB/EE4END[13] Tile_X5Y2_LUT4AB/EE4END[14] Tile_X5Y2_LUT4AB/EE4END[15]
+ Tile_X5Y2_LUT4AB/EE4END[1] Tile_X5Y2_LUT4AB/EE4END[2] Tile_X5Y2_LUT4AB/EE4END[3]
+ Tile_X5Y2_LUT4AB/EE4END[4] Tile_X5Y2_LUT4AB/EE4END[5] Tile_X5Y2_LUT4AB/EE4END[6]
+ Tile_X5Y2_LUT4AB/EE4END[7] Tile_X5Y2_LUT4AB/EE4END[8] Tile_X5Y2_LUT4AB/EE4END[9]
+ Tile_X5Y2_LUT4AB/FrameData[0] Tile_X5Y2_LUT4AB/FrameData[10] Tile_X5Y2_LUT4AB/FrameData[11]
+ Tile_X5Y2_LUT4AB/FrameData[12] Tile_X5Y2_LUT4AB/FrameData[13] Tile_X5Y2_LUT4AB/FrameData[14]
+ Tile_X5Y2_LUT4AB/FrameData[15] Tile_X5Y2_LUT4AB/FrameData[16] Tile_X5Y2_LUT4AB/FrameData[17]
+ Tile_X5Y2_LUT4AB/FrameData[18] Tile_X5Y2_LUT4AB/FrameData[19] Tile_X5Y2_LUT4AB/FrameData[1]
+ Tile_X5Y2_LUT4AB/FrameData[20] Tile_X5Y2_LUT4AB/FrameData[21] Tile_X5Y2_LUT4AB/FrameData[22]
+ Tile_X5Y2_LUT4AB/FrameData[23] Tile_X5Y2_LUT4AB/FrameData[24] Tile_X5Y2_LUT4AB/FrameData[25]
+ Tile_X5Y2_LUT4AB/FrameData[26] Tile_X5Y2_LUT4AB/FrameData[27] Tile_X5Y2_LUT4AB/FrameData[28]
+ Tile_X5Y2_LUT4AB/FrameData[29] Tile_X5Y2_LUT4AB/FrameData[2] Tile_X5Y2_LUT4AB/FrameData[30]
+ Tile_X5Y2_LUT4AB/FrameData[31] Tile_X5Y2_LUT4AB/FrameData[3] Tile_X5Y2_LUT4AB/FrameData[4]
+ Tile_X5Y2_LUT4AB/FrameData[5] Tile_X5Y2_LUT4AB/FrameData[6] Tile_X5Y2_LUT4AB/FrameData[7]
+ Tile_X5Y2_LUT4AB/FrameData[8] Tile_X5Y2_LUT4AB/FrameData[9] Tile_X6Y2_LUT4AB/FrameData[0]
+ Tile_X6Y2_LUT4AB/FrameData[10] Tile_X6Y2_LUT4AB/FrameData[11] Tile_X6Y2_LUT4AB/FrameData[12]
+ Tile_X6Y2_LUT4AB/FrameData[13] Tile_X6Y2_LUT4AB/FrameData[14] Tile_X6Y2_LUT4AB/FrameData[15]
+ Tile_X6Y2_LUT4AB/FrameData[16] Tile_X6Y2_LUT4AB/FrameData[17] Tile_X6Y2_LUT4AB/FrameData[18]
+ Tile_X6Y2_LUT4AB/FrameData[19] Tile_X6Y2_LUT4AB/FrameData[1] Tile_X6Y2_LUT4AB/FrameData[20]
+ Tile_X6Y2_LUT4AB/FrameData[21] Tile_X6Y2_LUT4AB/FrameData[22] Tile_X6Y2_LUT4AB/FrameData[23]
+ Tile_X6Y2_LUT4AB/FrameData[24] Tile_X6Y2_LUT4AB/FrameData[25] Tile_X6Y2_LUT4AB/FrameData[26]
+ Tile_X6Y2_LUT4AB/FrameData[27] Tile_X6Y2_LUT4AB/FrameData[28] Tile_X6Y2_LUT4AB/FrameData[29]
+ Tile_X6Y2_LUT4AB/FrameData[2] Tile_X6Y2_LUT4AB/FrameData[30] Tile_X6Y2_LUT4AB/FrameData[31]
+ Tile_X6Y2_LUT4AB/FrameData[3] Tile_X6Y2_LUT4AB/FrameData[4] Tile_X6Y2_LUT4AB/FrameData[5]
+ Tile_X6Y2_LUT4AB/FrameData[6] Tile_X6Y2_LUT4AB/FrameData[7] Tile_X6Y2_LUT4AB/FrameData[8]
+ Tile_X6Y2_LUT4AB/FrameData[9] Tile_X5Y2_LUT4AB/FrameStrobe[0] Tile_X5Y2_LUT4AB/FrameStrobe[10]
+ Tile_X5Y2_LUT4AB/FrameStrobe[11] Tile_X5Y2_LUT4AB/FrameStrobe[12] Tile_X5Y2_LUT4AB/FrameStrobe[13]
+ Tile_X5Y2_LUT4AB/FrameStrobe[14] Tile_X5Y2_LUT4AB/FrameStrobe[15] Tile_X5Y2_LUT4AB/FrameStrobe[16]
+ Tile_X5Y2_LUT4AB/FrameStrobe[17] Tile_X5Y2_LUT4AB/FrameStrobe[18] Tile_X5Y2_LUT4AB/FrameStrobe[19]
+ Tile_X5Y2_LUT4AB/FrameStrobe[1] Tile_X5Y2_LUT4AB/FrameStrobe[2] Tile_X5Y2_LUT4AB/FrameStrobe[3]
+ Tile_X5Y2_LUT4AB/FrameStrobe[4] Tile_X5Y2_LUT4AB/FrameStrobe[5] Tile_X5Y2_LUT4AB/FrameStrobe[6]
+ Tile_X5Y2_LUT4AB/FrameStrobe[7] Tile_X5Y2_LUT4AB/FrameStrobe[8] Tile_X5Y2_LUT4AB/FrameStrobe[9]
+ Tile_X5Y1_LUT4AB/FrameStrobe[0] Tile_X5Y1_LUT4AB/FrameStrobe[10] Tile_X5Y1_LUT4AB/FrameStrobe[11]
+ Tile_X5Y1_LUT4AB/FrameStrobe[12] Tile_X5Y1_LUT4AB/FrameStrobe[13] Tile_X5Y1_LUT4AB/FrameStrobe[14]
+ Tile_X5Y1_LUT4AB/FrameStrobe[15] Tile_X5Y1_LUT4AB/FrameStrobe[16] Tile_X5Y1_LUT4AB/FrameStrobe[17]
+ Tile_X5Y1_LUT4AB/FrameStrobe[18] Tile_X5Y1_LUT4AB/FrameStrobe[19] Tile_X5Y1_LUT4AB/FrameStrobe[1]
+ Tile_X5Y1_LUT4AB/FrameStrobe[2] Tile_X5Y1_LUT4AB/FrameStrobe[3] Tile_X5Y1_LUT4AB/FrameStrobe[4]
+ Tile_X5Y1_LUT4AB/FrameStrobe[5] Tile_X5Y1_LUT4AB/FrameStrobe[6] Tile_X5Y1_LUT4AB/FrameStrobe[7]
+ Tile_X5Y1_LUT4AB/FrameStrobe[8] Tile_X5Y1_LUT4AB/FrameStrobe[9] Tile_X5Y2_LUT4AB/N1BEG[0]
+ Tile_X5Y2_LUT4AB/N1BEG[1] Tile_X5Y2_LUT4AB/N1BEG[2] Tile_X5Y2_LUT4AB/N1BEG[3] Tile_X5Y3_LUT4AB/N1BEG[0]
+ Tile_X5Y3_LUT4AB/N1BEG[1] Tile_X5Y3_LUT4AB/N1BEG[2] Tile_X5Y3_LUT4AB/N1BEG[3] Tile_X5Y2_LUT4AB/N2BEG[0]
+ Tile_X5Y2_LUT4AB/N2BEG[1] Tile_X5Y2_LUT4AB/N2BEG[2] Tile_X5Y2_LUT4AB/N2BEG[3] Tile_X5Y2_LUT4AB/N2BEG[4]
+ Tile_X5Y2_LUT4AB/N2BEG[5] Tile_X5Y2_LUT4AB/N2BEG[6] Tile_X5Y2_LUT4AB/N2BEG[7] Tile_X5Y1_LUT4AB/N2END[0]
+ Tile_X5Y1_LUT4AB/N2END[1] Tile_X5Y1_LUT4AB/N2END[2] Tile_X5Y1_LUT4AB/N2END[3] Tile_X5Y1_LUT4AB/N2END[4]
+ Tile_X5Y1_LUT4AB/N2END[5] Tile_X5Y1_LUT4AB/N2END[6] Tile_X5Y1_LUT4AB/N2END[7] Tile_X5Y2_LUT4AB/N2END[0]
+ Tile_X5Y2_LUT4AB/N2END[1] Tile_X5Y2_LUT4AB/N2END[2] Tile_X5Y2_LUT4AB/N2END[3] Tile_X5Y2_LUT4AB/N2END[4]
+ Tile_X5Y2_LUT4AB/N2END[5] Tile_X5Y2_LUT4AB/N2END[6] Tile_X5Y2_LUT4AB/N2END[7] Tile_X5Y3_LUT4AB/N2BEG[0]
+ Tile_X5Y3_LUT4AB/N2BEG[1] Tile_X5Y3_LUT4AB/N2BEG[2] Tile_X5Y3_LUT4AB/N2BEG[3] Tile_X5Y3_LUT4AB/N2BEG[4]
+ Tile_X5Y3_LUT4AB/N2BEG[5] Tile_X5Y3_LUT4AB/N2BEG[6] Tile_X5Y3_LUT4AB/N2BEG[7] Tile_X5Y2_LUT4AB/N4BEG[0]
+ Tile_X5Y2_LUT4AB/N4BEG[10] Tile_X5Y2_LUT4AB/N4BEG[11] Tile_X5Y2_LUT4AB/N4BEG[12]
+ Tile_X5Y2_LUT4AB/N4BEG[13] Tile_X5Y2_LUT4AB/N4BEG[14] Tile_X5Y2_LUT4AB/N4BEG[15]
+ Tile_X5Y2_LUT4AB/N4BEG[1] Tile_X5Y2_LUT4AB/N4BEG[2] Tile_X5Y2_LUT4AB/N4BEG[3] Tile_X5Y2_LUT4AB/N4BEG[4]
+ Tile_X5Y2_LUT4AB/N4BEG[5] Tile_X5Y2_LUT4AB/N4BEG[6] Tile_X5Y2_LUT4AB/N4BEG[7] Tile_X5Y2_LUT4AB/N4BEG[8]
+ Tile_X5Y2_LUT4AB/N4BEG[9] Tile_X5Y3_LUT4AB/N4BEG[0] Tile_X5Y3_LUT4AB/N4BEG[10] Tile_X5Y3_LUT4AB/N4BEG[11]
+ Tile_X5Y3_LUT4AB/N4BEG[12] Tile_X5Y3_LUT4AB/N4BEG[13] Tile_X5Y3_LUT4AB/N4BEG[14]
+ Tile_X5Y3_LUT4AB/N4BEG[15] Tile_X5Y3_LUT4AB/N4BEG[1] Tile_X5Y3_LUT4AB/N4BEG[2] Tile_X5Y3_LUT4AB/N4BEG[3]
+ Tile_X5Y3_LUT4AB/N4BEG[4] Tile_X5Y3_LUT4AB/N4BEG[5] Tile_X5Y3_LUT4AB/N4BEG[6] Tile_X5Y3_LUT4AB/N4BEG[7]
+ Tile_X5Y3_LUT4AB/N4BEG[8] Tile_X5Y3_LUT4AB/N4BEG[9] Tile_X5Y2_LUT4AB/NN4BEG[0] Tile_X5Y2_LUT4AB/NN4BEG[10]
+ Tile_X5Y2_LUT4AB/NN4BEG[11] Tile_X5Y2_LUT4AB/NN4BEG[12] Tile_X5Y2_LUT4AB/NN4BEG[13]
+ Tile_X5Y2_LUT4AB/NN4BEG[14] Tile_X5Y2_LUT4AB/NN4BEG[15] Tile_X5Y2_LUT4AB/NN4BEG[1]
+ Tile_X5Y2_LUT4AB/NN4BEG[2] Tile_X5Y2_LUT4AB/NN4BEG[3] Tile_X5Y2_LUT4AB/NN4BEG[4]
+ Tile_X5Y2_LUT4AB/NN4BEG[5] Tile_X5Y2_LUT4AB/NN4BEG[6] Tile_X5Y2_LUT4AB/NN4BEG[7]
+ Tile_X5Y2_LUT4AB/NN4BEG[8] Tile_X5Y2_LUT4AB/NN4BEG[9] Tile_X5Y3_LUT4AB/NN4BEG[0]
+ Tile_X5Y3_LUT4AB/NN4BEG[10] Tile_X5Y3_LUT4AB/NN4BEG[11] Tile_X5Y3_LUT4AB/NN4BEG[12]
+ Tile_X5Y3_LUT4AB/NN4BEG[13] Tile_X5Y3_LUT4AB/NN4BEG[14] Tile_X5Y3_LUT4AB/NN4BEG[15]
+ Tile_X5Y3_LUT4AB/NN4BEG[1] Tile_X5Y3_LUT4AB/NN4BEG[2] Tile_X5Y3_LUT4AB/NN4BEG[3]
+ Tile_X5Y3_LUT4AB/NN4BEG[4] Tile_X5Y3_LUT4AB/NN4BEG[5] Tile_X5Y3_LUT4AB/NN4BEG[6]
+ Tile_X5Y3_LUT4AB/NN4BEG[7] Tile_X5Y3_LUT4AB/NN4BEG[8] Tile_X5Y3_LUT4AB/NN4BEG[9]
+ Tile_X5Y3_LUT4AB/S1END[0] Tile_X5Y3_LUT4AB/S1END[1] Tile_X5Y3_LUT4AB/S1END[2] Tile_X5Y3_LUT4AB/S1END[3]
+ Tile_X5Y2_LUT4AB/S1END[0] Tile_X5Y2_LUT4AB/S1END[1] Tile_X5Y2_LUT4AB/S1END[2] Tile_X5Y2_LUT4AB/S1END[3]
+ Tile_X5Y3_LUT4AB/S2MID[0] Tile_X5Y3_LUT4AB/S2MID[1] Tile_X5Y3_LUT4AB/S2MID[2] Tile_X5Y3_LUT4AB/S2MID[3]
+ Tile_X5Y3_LUT4AB/S2MID[4] Tile_X5Y3_LUT4AB/S2MID[5] Tile_X5Y3_LUT4AB/S2MID[6] Tile_X5Y3_LUT4AB/S2MID[7]
+ Tile_X5Y3_LUT4AB/S2END[0] Tile_X5Y3_LUT4AB/S2END[1] Tile_X5Y3_LUT4AB/S2END[2] Tile_X5Y3_LUT4AB/S2END[3]
+ Tile_X5Y3_LUT4AB/S2END[4] Tile_X5Y3_LUT4AB/S2END[5] Tile_X5Y3_LUT4AB/S2END[6] Tile_X5Y3_LUT4AB/S2END[7]
+ Tile_X5Y2_LUT4AB/S2END[0] Tile_X5Y2_LUT4AB/S2END[1] Tile_X5Y2_LUT4AB/S2END[2] Tile_X5Y2_LUT4AB/S2END[3]
+ Tile_X5Y2_LUT4AB/S2END[4] Tile_X5Y2_LUT4AB/S2END[5] Tile_X5Y2_LUT4AB/S2END[6] Tile_X5Y2_LUT4AB/S2END[7]
+ Tile_X5Y2_LUT4AB/S2MID[0] Tile_X5Y2_LUT4AB/S2MID[1] Tile_X5Y2_LUT4AB/S2MID[2] Tile_X5Y2_LUT4AB/S2MID[3]
+ Tile_X5Y2_LUT4AB/S2MID[4] Tile_X5Y2_LUT4AB/S2MID[5] Tile_X5Y2_LUT4AB/S2MID[6] Tile_X5Y2_LUT4AB/S2MID[7]
+ Tile_X5Y3_LUT4AB/S4END[0] Tile_X5Y3_LUT4AB/S4END[10] Tile_X5Y3_LUT4AB/S4END[11]
+ Tile_X5Y3_LUT4AB/S4END[12] Tile_X5Y3_LUT4AB/S4END[13] Tile_X5Y3_LUT4AB/S4END[14]
+ Tile_X5Y3_LUT4AB/S4END[15] Tile_X5Y3_LUT4AB/S4END[1] Tile_X5Y3_LUT4AB/S4END[2] Tile_X5Y3_LUT4AB/S4END[3]
+ Tile_X5Y3_LUT4AB/S4END[4] Tile_X5Y3_LUT4AB/S4END[5] Tile_X5Y3_LUT4AB/S4END[6] Tile_X5Y3_LUT4AB/S4END[7]
+ Tile_X5Y3_LUT4AB/S4END[8] Tile_X5Y3_LUT4AB/S4END[9] Tile_X5Y2_LUT4AB/S4END[0] Tile_X5Y2_LUT4AB/S4END[10]
+ Tile_X5Y2_LUT4AB/S4END[11] Tile_X5Y2_LUT4AB/S4END[12] Tile_X5Y2_LUT4AB/S4END[13]
+ Tile_X5Y2_LUT4AB/S4END[14] Tile_X5Y2_LUT4AB/S4END[15] Tile_X5Y2_LUT4AB/S4END[1]
+ Tile_X5Y2_LUT4AB/S4END[2] Tile_X5Y2_LUT4AB/S4END[3] Tile_X5Y2_LUT4AB/S4END[4] Tile_X5Y2_LUT4AB/S4END[5]
+ Tile_X5Y2_LUT4AB/S4END[6] Tile_X5Y2_LUT4AB/S4END[7] Tile_X5Y2_LUT4AB/S4END[8] Tile_X5Y2_LUT4AB/S4END[9]
+ Tile_X5Y3_LUT4AB/SS4END[0] Tile_X5Y3_LUT4AB/SS4END[10] Tile_X5Y3_LUT4AB/SS4END[11]
+ Tile_X5Y3_LUT4AB/SS4END[12] Tile_X5Y3_LUT4AB/SS4END[13] Tile_X5Y3_LUT4AB/SS4END[14]
+ Tile_X5Y3_LUT4AB/SS4END[15] Tile_X5Y3_LUT4AB/SS4END[1] Tile_X5Y3_LUT4AB/SS4END[2]
+ Tile_X5Y3_LUT4AB/SS4END[3] Tile_X5Y3_LUT4AB/SS4END[4] Tile_X5Y3_LUT4AB/SS4END[5]
+ Tile_X5Y3_LUT4AB/SS4END[6] Tile_X5Y3_LUT4AB/SS4END[7] Tile_X5Y3_LUT4AB/SS4END[8]
+ Tile_X5Y3_LUT4AB/SS4END[9] Tile_X5Y2_LUT4AB/SS4END[0] Tile_X5Y2_LUT4AB/SS4END[10]
+ Tile_X5Y2_LUT4AB/SS4END[11] Tile_X5Y2_LUT4AB/SS4END[12] Tile_X5Y2_LUT4AB/SS4END[13]
+ Tile_X5Y2_LUT4AB/SS4END[14] Tile_X5Y2_LUT4AB/SS4END[15] Tile_X5Y2_LUT4AB/SS4END[1]
+ Tile_X5Y2_LUT4AB/SS4END[2] Tile_X5Y2_LUT4AB/SS4END[3] Tile_X5Y2_LUT4AB/SS4END[4]
+ Tile_X5Y2_LUT4AB/SS4END[5] Tile_X5Y2_LUT4AB/SS4END[6] Tile_X5Y2_LUT4AB/SS4END[7]
+ Tile_X5Y2_LUT4AB/SS4END[8] Tile_X5Y2_LUT4AB/SS4END[9] Tile_X5Y2_LUT4AB/UserCLK Tile_X5Y1_LUT4AB/UserCLK
+ VGND VPWR Tile_X5Y2_LUT4AB/W1BEG[0] Tile_X5Y2_LUT4AB/W1BEG[1] Tile_X5Y2_LUT4AB/W1BEG[2]
+ Tile_X5Y2_LUT4AB/W1BEG[3] Tile_X6Y2_LUT4AB/W1BEG[0] Tile_X6Y2_LUT4AB/W1BEG[1] Tile_X6Y2_LUT4AB/W1BEG[2]
+ Tile_X6Y2_LUT4AB/W1BEG[3] Tile_X5Y2_LUT4AB/W2BEG[0] Tile_X5Y2_LUT4AB/W2BEG[1] Tile_X5Y2_LUT4AB/W2BEG[2]
+ Tile_X5Y2_LUT4AB/W2BEG[3] Tile_X5Y2_LUT4AB/W2BEG[4] Tile_X5Y2_LUT4AB/W2BEG[5] Tile_X5Y2_LUT4AB/W2BEG[6]
+ Tile_X5Y2_LUT4AB/W2BEG[7] Tile_X5Y2_LUT4AB/W2BEGb[0] Tile_X5Y2_LUT4AB/W2BEGb[1]
+ Tile_X5Y2_LUT4AB/W2BEGb[2] Tile_X5Y2_LUT4AB/W2BEGb[3] Tile_X5Y2_LUT4AB/W2BEGb[4]
+ Tile_X5Y2_LUT4AB/W2BEGb[5] Tile_X5Y2_LUT4AB/W2BEGb[6] Tile_X5Y2_LUT4AB/W2BEGb[7]
+ Tile_X5Y2_LUT4AB/W2END[0] Tile_X5Y2_LUT4AB/W2END[1] Tile_X5Y2_LUT4AB/W2END[2] Tile_X5Y2_LUT4AB/W2END[3]
+ Tile_X5Y2_LUT4AB/W2END[4] Tile_X5Y2_LUT4AB/W2END[5] Tile_X5Y2_LUT4AB/W2END[6] Tile_X5Y2_LUT4AB/W2END[7]
+ Tile_X6Y2_LUT4AB/W2BEG[0] Tile_X6Y2_LUT4AB/W2BEG[1] Tile_X6Y2_LUT4AB/W2BEG[2] Tile_X6Y2_LUT4AB/W2BEG[3]
+ Tile_X6Y2_LUT4AB/W2BEG[4] Tile_X6Y2_LUT4AB/W2BEG[5] Tile_X6Y2_LUT4AB/W2BEG[6] Tile_X6Y2_LUT4AB/W2BEG[7]
+ Tile_X5Y2_LUT4AB/W6BEG[0] Tile_X5Y2_LUT4AB/W6BEG[10] Tile_X5Y2_LUT4AB/W6BEG[11]
+ Tile_X5Y2_LUT4AB/W6BEG[1] Tile_X5Y2_LUT4AB/W6BEG[2] Tile_X5Y2_LUT4AB/W6BEG[3] Tile_X5Y2_LUT4AB/W6BEG[4]
+ Tile_X5Y2_LUT4AB/W6BEG[5] Tile_X5Y2_LUT4AB/W6BEG[6] Tile_X5Y2_LUT4AB/W6BEG[7] Tile_X5Y2_LUT4AB/W6BEG[8]
+ Tile_X5Y2_LUT4AB/W6BEG[9] Tile_X6Y2_LUT4AB/W6BEG[0] Tile_X6Y2_LUT4AB/W6BEG[10] Tile_X6Y2_LUT4AB/W6BEG[11]
+ Tile_X6Y2_LUT4AB/W6BEG[1] Tile_X6Y2_LUT4AB/W6BEG[2] Tile_X6Y2_LUT4AB/W6BEG[3] Tile_X6Y2_LUT4AB/W6BEG[4]
+ Tile_X6Y2_LUT4AB/W6BEG[5] Tile_X6Y2_LUT4AB/W6BEG[6] Tile_X6Y2_LUT4AB/W6BEG[7] Tile_X6Y2_LUT4AB/W6BEG[8]
+ Tile_X6Y2_LUT4AB/W6BEG[9] Tile_X5Y2_LUT4AB/WW4BEG[0] Tile_X5Y2_LUT4AB/WW4BEG[10]
+ Tile_X5Y2_LUT4AB/WW4BEG[11] Tile_X5Y2_LUT4AB/WW4BEG[12] Tile_X5Y2_LUT4AB/WW4BEG[13]
+ Tile_X5Y2_LUT4AB/WW4BEG[14] Tile_X5Y2_LUT4AB/WW4BEG[15] Tile_X5Y2_LUT4AB/WW4BEG[1]
+ Tile_X5Y2_LUT4AB/WW4BEG[2] Tile_X5Y2_LUT4AB/WW4BEG[3] Tile_X5Y2_LUT4AB/WW4BEG[4]
+ Tile_X5Y2_LUT4AB/WW4BEG[5] Tile_X5Y2_LUT4AB/WW4BEG[6] Tile_X5Y2_LUT4AB/WW4BEG[7]
+ Tile_X5Y2_LUT4AB/WW4BEG[8] Tile_X5Y2_LUT4AB/WW4BEG[9] Tile_X6Y2_LUT4AB/WW4BEG[0]
+ Tile_X6Y2_LUT4AB/WW4BEG[10] Tile_X6Y2_LUT4AB/WW4BEG[11] Tile_X6Y2_LUT4AB/WW4BEG[12]
+ Tile_X6Y2_LUT4AB/WW4BEG[13] Tile_X6Y2_LUT4AB/WW4BEG[14] Tile_X6Y2_LUT4AB/WW4BEG[15]
+ Tile_X6Y2_LUT4AB/WW4BEG[1] Tile_X6Y2_LUT4AB/WW4BEG[2] Tile_X6Y2_LUT4AB/WW4BEG[3]
+ Tile_X6Y2_LUT4AB/WW4BEG[4] Tile_X6Y2_LUT4AB/WW4BEG[5] Tile_X6Y2_LUT4AB/WW4BEG[6]
+ Tile_X6Y2_LUT4AB/WW4BEG[7] Tile_X6Y2_LUT4AB/WW4BEG[8] Tile_X6Y2_LUT4AB/WW4BEG[9]
+ LUT4AB
XTile_X9Y14_LUT4AB Tile_X9Y14_LUT4AB/Ci Tile_X9Y14_LUT4AB/Co Tile_X9Y14_LUT4AB/E1BEG[0]
+ Tile_X9Y14_LUT4AB/E1BEG[1] Tile_X9Y14_LUT4AB/E1BEG[2] Tile_X9Y14_LUT4AB/E1BEG[3]
+ Tile_X9Y14_LUT4AB/E1END[0] Tile_X9Y14_LUT4AB/E1END[1] Tile_X9Y14_LUT4AB/E1END[2]
+ Tile_X9Y14_LUT4AB/E1END[3] Tile_X9Y14_LUT4AB/E2BEG[0] Tile_X9Y14_LUT4AB/E2BEG[1]
+ Tile_X9Y14_LUT4AB/E2BEG[2] Tile_X9Y14_LUT4AB/E2BEG[3] Tile_X9Y14_LUT4AB/E2BEG[4]
+ Tile_X9Y14_LUT4AB/E2BEG[5] Tile_X9Y14_LUT4AB/E2BEG[6] Tile_X9Y14_LUT4AB/E2BEG[7]
+ Tile_X9Y14_LUT4AB/E2BEGb[0] Tile_X9Y14_LUT4AB/E2BEGb[1] Tile_X9Y14_LUT4AB/E2BEGb[2]
+ Tile_X9Y14_LUT4AB/E2BEGb[3] Tile_X9Y14_LUT4AB/E2BEGb[4] Tile_X9Y14_LUT4AB/E2BEGb[5]
+ Tile_X9Y14_LUT4AB/E2BEGb[6] Tile_X9Y14_LUT4AB/E2BEGb[7] Tile_X9Y14_LUT4AB/E2END[0]
+ Tile_X9Y14_LUT4AB/E2END[1] Tile_X9Y14_LUT4AB/E2END[2] Tile_X9Y14_LUT4AB/E2END[3]
+ Tile_X9Y14_LUT4AB/E2END[4] Tile_X9Y14_LUT4AB/E2END[5] Tile_X9Y14_LUT4AB/E2END[6]
+ Tile_X9Y14_LUT4AB/E2END[7] Tile_X9Y14_LUT4AB/E2MID[0] Tile_X9Y14_LUT4AB/E2MID[1]
+ Tile_X9Y14_LUT4AB/E2MID[2] Tile_X9Y14_LUT4AB/E2MID[3] Tile_X9Y14_LUT4AB/E2MID[4]
+ Tile_X9Y14_LUT4AB/E2MID[5] Tile_X9Y14_LUT4AB/E2MID[6] Tile_X9Y14_LUT4AB/E2MID[7]
+ Tile_X9Y14_LUT4AB/E6BEG[0] Tile_X9Y14_LUT4AB/E6BEG[10] Tile_X9Y14_LUT4AB/E6BEG[11]
+ Tile_X9Y14_LUT4AB/E6BEG[1] Tile_X9Y14_LUT4AB/E6BEG[2] Tile_X9Y14_LUT4AB/E6BEG[3]
+ Tile_X9Y14_LUT4AB/E6BEG[4] Tile_X9Y14_LUT4AB/E6BEG[5] Tile_X9Y14_LUT4AB/E6BEG[6]
+ Tile_X9Y14_LUT4AB/E6BEG[7] Tile_X9Y14_LUT4AB/E6BEG[8] Tile_X9Y14_LUT4AB/E6BEG[9]
+ Tile_X9Y14_LUT4AB/E6END[0] Tile_X9Y14_LUT4AB/E6END[10] Tile_X9Y14_LUT4AB/E6END[11]
+ Tile_X9Y14_LUT4AB/E6END[1] Tile_X9Y14_LUT4AB/E6END[2] Tile_X9Y14_LUT4AB/E6END[3]
+ Tile_X9Y14_LUT4AB/E6END[4] Tile_X9Y14_LUT4AB/E6END[5] Tile_X9Y14_LUT4AB/E6END[6]
+ Tile_X9Y14_LUT4AB/E6END[7] Tile_X9Y14_LUT4AB/E6END[8] Tile_X9Y14_LUT4AB/E6END[9]
+ Tile_X9Y14_LUT4AB/EE4BEG[0] Tile_X9Y14_LUT4AB/EE4BEG[10] Tile_X9Y14_LUT4AB/EE4BEG[11]
+ Tile_X9Y14_LUT4AB/EE4BEG[12] Tile_X9Y14_LUT4AB/EE4BEG[13] Tile_X9Y14_LUT4AB/EE4BEG[14]
+ Tile_X9Y14_LUT4AB/EE4BEG[15] Tile_X9Y14_LUT4AB/EE4BEG[1] Tile_X9Y14_LUT4AB/EE4BEG[2]
+ Tile_X9Y14_LUT4AB/EE4BEG[3] Tile_X9Y14_LUT4AB/EE4BEG[4] Tile_X9Y14_LUT4AB/EE4BEG[5]
+ Tile_X9Y14_LUT4AB/EE4BEG[6] Tile_X9Y14_LUT4AB/EE4BEG[7] Tile_X9Y14_LUT4AB/EE4BEG[8]
+ Tile_X9Y14_LUT4AB/EE4BEG[9] Tile_X9Y14_LUT4AB/EE4END[0] Tile_X9Y14_LUT4AB/EE4END[10]
+ Tile_X9Y14_LUT4AB/EE4END[11] Tile_X9Y14_LUT4AB/EE4END[12] Tile_X9Y14_LUT4AB/EE4END[13]
+ Tile_X9Y14_LUT4AB/EE4END[14] Tile_X9Y14_LUT4AB/EE4END[15] Tile_X9Y14_LUT4AB/EE4END[1]
+ Tile_X9Y14_LUT4AB/EE4END[2] Tile_X9Y14_LUT4AB/EE4END[3] Tile_X9Y14_LUT4AB/EE4END[4]
+ Tile_X9Y14_LUT4AB/EE4END[5] Tile_X9Y14_LUT4AB/EE4END[6] Tile_X9Y14_LUT4AB/EE4END[7]
+ Tile_X9Y14_LUT4AB/EE4END[8] Tile_X9Y14_LUT4AB/EE4END[9] Tile_X9Y14_LUT4AB/FrameData[0]
+ Tile_X9Y14_LUT4AB/FrameData[10] Tile_X9Y14_LUT4AB/FrameData[11] Tile_X9Y14_LUT4AB/FrameData[12]
+ Tile_X9Y14_LUT4AB/FrameData[13] Tile_X9Y14_LUT4AB/FrameData[14] Tile_X9Y14_LUT4AB/FrameData[15]
+ Tile_X9Y14_LUT4AB/FrameData[16] Tile_X9Y14_LUT4AB/FrameData[17] Tile_X9Y14_LUT4AB/FrameData[18]
+ Tile_X9Y14_LUT4AB/FrameData[19] Tile_X9Y14_LUT4AB/FrameData[1] Tile_X9Y14_LUT4AB/FrameData[20]
+ Tile_X9Y14_LUT4AB/FrameData[21] Tile_X9Y14_LUT4AB/FrameData[22] Tile_X9Y14_LUT4AB/FrameData[23]
+ Tile_X9Y14_LUT4AB/FrameData[24] Tile_X9Y14_LUT4AB/FrameData[25] Tile_X9Y14_LUT4AB/FrameData[26]
+ Tile_X9Y14_LUT4AB/FrameData[27] Tile_X9Y14_LUT4AB/FrameData[28] Tile_X9Y14_LUT4AB/FrameData[29]
+ Tile_X9Y14_LUT4AB/FrameData[2] Tile_X9Y14_LUT4AB/FrameData[30] Tile_X9Y14_LUT4AB/FrameData[31]
+ Tile_X9Y14_LUT4AB/FrameData[3] Tile_X9Y14_LUT4AB/FrameData[4] Tile_X9Y14_LUT4AB/FrameData[5]
+ Tile_X9Y14_LUT4AB/FrameData[6] Tile_X9Y14_LUT4AB/FrameData[7] Tile_X9Y14_LUT4AB/FrameData[8]
+ Tile_X9Y14_LUT4AB/FrameData[9] Tile_X9Y14_LUT4AB/FrameData_O[0] Tile_X9Y14_LUT4AB/FrameData_O[10]
+ Tile_X9Y14_LUT4AB/FrameData_O[11] Tile_X9Y14_LUT4AB/FrameData_O[12] Tile_X9Y14_LUT4AB/FrameData_O[13]
+ Tile_X9Y14_LUT4AB/FrameData_O[14] Tile_X9Y14_LUT4AB/FrameData_O[15] Tile_X9Y14_LUT4AB/FrameData_O[16]
+ Tile_X9Y14_LUT4AB/FrameData_O[17] Tile_X9Y14_LUT4AB/FrameData_O[18] Tile_X9Y14_LUT4AB/FrameData_O[19]
+ Tile_X9Y14_LUT4AB/FrameData_O[1] Tile_X9Y14_LUT4AB/FrameData_O[20] Tile_X9Y14_LUT4AB/FrameData_O[21]
+ Tile_X9Y14_LUT4AB/FrameData_O[22] Tile_X9Y14_LUT4AB/FrameData_O[23] Tile_X9Y14_LUT4AB/FrameData_O[24]
+ Tile_X9Y14_LUT4AB/FrameData_O[25] Tile_X9Y14_LUT4AB/FrameData_O[26] Tile_X9Y14_LUT4AB/FrameData_O[27]
+ Tile_X9Y14_LUT4AB/FrameData_O[28] Tile_X9Y14_LUT4AB/FrameData_O[29] Tile_X9Y14_LUT4AB/FrameData_O[2]
+ Tile_X9Y14_LUT4AB/FrameData_O[30] Tile_X9Y14_LUT4AB/FrameData_O[31] Tile_X9Y14_LUT4AB/FrameData_O[3]
+ Tile_X9Y14_LUT4AB/FrameData_O[4] Tile_X9Y14_LUT4AB/FrameData_O[5] Tile_X9Y14_LUT4AB/FrameData_O[6]
+ Tile_X9Y14_LUT4AB/FrameData_O[7] Tile_X9Y14_LUT4AB/FrameData_O[8] Tile_X9Y14_LUT4AB/FrameData_O[9]
+ Tile_X9Y14_LUT4AB/FrameStrobe[0] Tile_X9Y14_LUT4AB/FrameStrobe[10] Tile_X9Y14_LUT4AB/FrameStrobe[11]
+ Tile_X9Y14_LUT4AB/FrameStrobe[12] Tile_X9Y14_LUT4AB/FrameStrobe[13] Tile_X9Y14_LUT4AB/FrameStrobe[14]
+ Tile_X9Y14_LUT4AB/FrameStrobe[15] Tile_X9Y14_LUT4AB/FrameStrobe[16] Tile_X9Y14_LUT4AB/FrameStrobe[17]
+ Tile_X9Y14_LUT4AB/FrameStrobe[18] Tile_X9Y14_LUT4AB/FrameStrobe[19] Tile_X9Y14_LUT4AB/FrameStrobe[1]
+ Tile_X9Y14_LUT4AB/FrameStrobe[2] Tile_X9Y14_LUT4AB/FrameStrobe[3] Tile_X9Y14_LUT4AB/FrameStrobe[4]
+ Tile_X9Y14_LUT4AB/FrameStrobe[5] Tile_X9Y14_LUT4AB/FrameStrobe[6] Tile_X9Y14_LUT4AB/FrameStrobe[7]
+ Tile_X9Y14_LUT4AB/FrameStrobe[8] Tile_X9Y14_LUT4AB/FrameStrobe[9] Tile_X9Y13_LUT4AB/FrameStrobe[0]
+ Tile_X9Y13_LUT4AB/FrameStrobe[10] Tile_X9Y13_LUT4AB/FrameStrobe[11] Tile_X9Y13_LUT4AB/FrameStrobe[12]
+ Tile_X9Y13_LUT4AB/FrameStrobe[13] Tile_X9Y13_LUT4AB/FrameStrobe[14] Tile_X9Y13_LUT4AB/FrameStrobe[15]
+ Tile_X9Y13_LUT4AB/FrameStrobe[16] Tile_X9Y13_LUT4AB/FrameStrobe[17] Tile_X9Y13_LUT4AB/FrameStrobe[18]
+ Tile_X9Y13_LUT4AB/FrameStrobe[19] Tile_X9Y13_LUT4AB/FrameStrobe[1] Tile_X9Y13_LUT4AB/FrameStrobe[2]
+ Tile_X9Y13_LUT4AB/FrameStrobe[3] Tile_X9Y13_LUT4AB/FrameStrobe[4] Tile_X9Y13_LUT4AB/FrameStrobe[5]
+ Tile_X9Y13_LUT4AB/FrameStrobe[6] Tile_X9Y13_LUT4AB/FrameStrobe[7] Tile_X9Y13_LUT4AB/FrameStrobe[8]
+ Tile_X9Y13_LUT4AB/FrameStrobe[9] Tile_X9Y14_LUT4AB/N1BEG[0] Tile_X9Y14_LUT4AB/N1BEG[1]
+ Tile_X9Y14_LUT4AB/N1BEG[2] Tile_X9Y14_LUT4AB/N1BEG[3] Tile_X9Y14_LUT4AB/N1END[0]
+ Tile_X9Y14_LUT4AB/N1END[1] Tile_X9Y14_LUT4AB/N1END[2] Tile_X9Y14_LUT4AB/N1END[3]
+ Tile_X9Y14_LUT4AB/N2BEG[0] Tile_X9Y14_LUT4AB/N2BEG[1] Tile_X9Y14_LUT4AB/N2BEG[2]
+ Tile_X9Y14_LUT4AB/N2BEG[3] Tile_X9Y14_LUT4AB/N2BEG[4] Tile_X9Y14_LUT4AB/N2BEG[5]
+ Tile_X9Y14_LUT4AB/N2BEG[6] Tile_X9Y14_LUT4AB/N2BEG[7] Tile_X9Y13_LUT4AB/N2END[0]
+ Tile_X9Y13_LUT4AB/N2END[1] Tile_X9Y13_LUT4AB/N2END[2] Tile_X9Y13_LUT4AB/N2END[3]
+ Tile_X9Y13_LUT4AB/N2END[4] Tile_X9Y13_LUT4AB/N2END[5] Tile_X9Y13_LUT4AB/N2END[6]
+ Tile_X9Y13_LUT4AB/N2END[7] Tile_X9Y14_LUT4AB/N2END[0] Tile_X9Y14_LUT4AB/N2END[1]
+ Tile_X9Y14_LUT4AB/N2END[2] Tile_X9Y14_LUT4AB/N2END[3] Tile_X9Y14_LUT4AB/N2END[4]
+ Tile_X9Y14_LUT4AB/N2END[5] Tile_X9Y14_LUT4AB/N2END[6] Tile_X9Y14_LUT4AB/N2END[7]
+ Tile_X9Y14_LUT4AB/N2MID[0] Tile_X9Y14_LUT4AB/N2MID[1] Tile_X9Y14_LUT4AB/N2MID[2]
+ Tile_X9Y14_LUT4AB/N2MID[3] Tile_X9Y14_LUT4AB/N2MID[4] Tile_X9Y14_LUT4AB/N2MID[5]
+ Tile_X9Y14_LUT4AB/N2MID[6] Tile_X9Y14_LUT4AB/N2MID[7] Tile_X9Y14_LUT4AB/N4BEG[0]
+ Tile_X9Y14_LUT4AB/N4BEG[10] Tile_X9Y14_LUT4AB/N4BEG[11] Tile_X9Y14_LUT4AB/N4BEG[12]
+ Tile_X9Y14_LUT4AB/N4BEG[13] Tile_X9Y14_LUT4AB/N4BEG[14] Tile_X9Y14_LUT4AB/N4BEG[15]
+ Tile_X9Y14_LUT4AB/N4BEG[1] Tile_X9Y14_LUT4AB/N4BEG[2] Tile_X9Y14_LUT4AB/N4BEG[3]
+ Tile_X9Y14_LUT4AB/N4BEG[4] Tile_X9Y14_LUT4AB/N4BEG[5] Tile_X9Y14_LUT4AB/N4BEG[6]
+ Tile_X9Y14_LUT4AB/N4BEG[7] Tile_X9Y14_LUT4AB/N4BEG[8] Tile_X9Y14_LUT4AB/N4BEG[9]
+ Tile_X9Y14_LUT4AB/N4END[0] Tile_X9Y14_LUT4AB/N4END[10] Tile_X9Y14_LUT4AB/N4END[11]
+ Tile_X9Y14_LUT4AB/N4END[12] Tile_X9Y14_LUT4AB/N4END[13] Tile_X9Y14_LUT4AB/N4END[14]
+ Tile_X9Y14_LUT4AB/N4END[15] Tile_X9Y14_LUT4AB/N4END[1] Tile_X9Y14_LUT4AB/N4END[2]
+ Tile_X9Y14_LUT4AB/N4END[3] Tile_X9Y14_LUT4AB/N4END[4] Tile_X9Y14_LUT4AB/N4END[5]
+ Tile_X9Y14_LUT4AB/N4END[6] Tile_X9Y14_LUT4AB/N4END[7] Tile_X9Y14_LUT4AB/N4END[8]
+ Tile_X9Y14_LUT4AB/N4END[9] Tile_X9Y14_LUT4AB/NN4BEG[0] Tile_X9Y14_LUT4AB/NN4BEG[10]
+ Tile_X9Y14_LUT4AB/NN4BEG[11] Tile_X9Y14_LUT4AB/NN4BEG[12] Tile_X9Y14_LUT4AB/NN4BEG[13]
+ Tile_X9Y14_LUT4AB/NN4BEG[14] Tile_X9Y14_LUT4AB/NN4BEG[15] Tile_X9Y14_LUT4AB/NN4BEG[1]
+ Tile_X9Y14_LUT4AB/NN4BEG[2] Tile_X9Y14_LUT4AB/NN4BEG[3] Tile_X9Y14_LUT4AB/NN4BEG[4]
+ Tile_X9Y14_LUT4AB/NN4BEG[5] Tile_X9Y14_LUT4AB/NN4BEG[6] Tile_X9Y14_LUT4AB/NN4BEG[7]
+ Tile_X9Y14_LUT4AB/NN4BEG[8] Tile_X9Y14_LUT4AB/NN4BEG[9] Tile_X9Y14_LUT4AB/NN4END[0]
+ Tile_X9Y14_LUT4AB/NN4END[10] Tile_X9Y14_LUT4AB/NN4END[11] Tile_X9Y14_LUT4AB/NN4END[12]
+ Tile_X9Y14_LUT4AB/NN4END[13] Tile_X9Y14_LUT4AB/NN4END[14] Tile_X9Y14_LUT4AB/NN4END[15]
+ Tile_X9Y14_LUT4AB/NN4END[1] Tile_X9Y14_LUT4AB/NN4END[2] Tile_X9Y14_LUT4AB/NN4END[3]
+ Tile_X9Y14_LUT4AB/NN4END[4] Tile_X9Y14_LUT4AB/NN4END[5] Tile_X9Y14_LUT4AB/NN4END[6]
+ Tile_X9Y14_LUT4AB/NN4END[7] Tile_X9Y14_LUT4AB/NN4END[8] Tile_X9Y14_LUT4AB/NN4END[9]
+ Tile_X9Y14_LUT4AB/S1BEG[0] Tile_X9Y14_LUT4AB/S1BEG[1] Tile_X9Y14_LUT4AB/S1BEG[2]
+ Tile_X9Y14_LUT4AB/S1BEG[3] Tile_X9Y14_LUT4AB/S1END[0] Tile_X9Y14_LUT4AB/S1END[1]
+ Tile_X9Y14_LUT4AB/S1END[2] Tile_X9Y14_LUT4AB/S1END[3] Tile_X9Y14_LUT4AB/S2BEG[0]
+ Tile_X9Y14_LUT4AB/S2BEG[1] Tile_X9Y14_LUT4AB/S2BEG[2] Tile_X9Y14_LUT4AB/S2BEG[3]
+ Tile_X9Y14_LUT4AB/S2BEG[4] Tile_X9Y14_LUT4AB/S2BEG[5] Tile_X9Y14_LUT4AB/S2BEG[6]
+ Tile_X9Y14_LUT4AB/S2BEG[7] Tile_X9Y14_LUT4AB/S2BEGb[0] Tile_X9Y14_LUT4AB/S2BEGb[1]
+ Tile_X9Y14_LUT4AB/S2BEGb[2] Tile_X9Y14_LUT4AB/S2BEGb[3] Tile_X9Y14_LUT4AB/S2BEGb[4]
+ Tile_X9Y14_LUT4AB/S2BEGb[5] Tile_X9Y14_LUT4AB/S2BEGb[6] Tile_X9Y14_LUT4AB/S2BEGb[7]
+ Tile_X9Y14_LUT4AB/S2END[0] Tile_X9Y14_LUT4AB/S2END[1] Tile_X9Y14_LUT4AB/S2END[2]
+ Tile_X9Y14_LUT4AB/S2END[3] Tile_X9Y14_LUT4AB/S2END[4] Tile_X9Y14_LUT4AB/S2END[5]
+ Tile_X9Y14_LUT4AB/S2END[6] Tile_X9Y14_LUT4AB/S2END[7] Tile_X9Y14_LUT4AB/S2MID[0]
+ Tile_X9Y14_LUT4AB/S2MID[1] Tile_X9Y14_LUT4AB/S2MID[2] Tile_X9Y14_LUT4AB/S2MID[3]
+ Tile_X9Y14_LUT4AB/S2MID[4] Tile_X9Y14_LUT4AB/S2MID[5] Tile_X9Y14_LUT4AB/S2MID[6]
+ Tile_X9Y14_LUT4AB/S2MID[7] Tile_X9Y14_LUT4AB/S4BEG[0] Tile_X9Y14_LUT4AB/S4BEG[10]
+ Tile_X9Y14_LUT4AB/S4BEG[11] Tile_X9Y14_LUT4AB/S4BEG[12] Tile_X9Y14_LUT4AB/S4BEG[13]
+ Tile_X9Y14_LUT4AB/S4BEG[14] Tile_X9Y14_LUT4AB/S4BEG[15] Tile_X9Y14_LUT4AB/S4BEG[1]
+ Tile_X9Y14_LUT4AB/S4BEG[2] Tile_X9Y14_LUT4AB/S4BEG[3] Tile_X9Y14_LUT4AB/S4BEG[4]
+ Tile_X9Y14_LUT4AB/S4BEG[5] Tile_X9Y14_LUT4AB/S4BEG[6] Tile_X9Y14_LUT4AB/S4BEG[7]
+ Tile_X9Y14_LUT4AB/S4BEG[8] Tile_X9Y14_LUT4AB/S4BEG[9] Tile_X9Y14_LUT4AB/S4END[0]
+ Tile_X9Y14_LUT4AB/S4END[10] Tile_X9Y14_LUT4AB/S4END[11] Tile_X9Y14_LUT4AB/S4END[12]
+ Tile_X9Y14_LUT4AB/S4END[13] Tile_X9Y14_LUT4AB/S4END[14] Tile_X9Y14_LUT4AB/S4END[15]
+ Tile_X9Y14_LUT4AB/S4END[1] Tile_X9Y14_LUT4AB/S4END[2] Tile_X9Y14_LUT4AB/S4END[3]
+ Tile_X9Y14_LUT4AB/S4END[4] Tile_X9Y14_LUT4AB/S4END[5] Tile_X9Y14_LUT4AB/S4END[6]
+ Tile_X9Y14_LUT4AB/S4END[7] Tile_X9Y14_LUT4AB/S4END[8] Tile_X9Y14_LUT4AB/S4END[9]
+ Tile_X9Y14_LUT4AB/SS4BEG[0] Tile_X9Y14_LUT4AB/SS4BEG[10] Tile_X9Y14_LUT4AB/SS4BEG[11]
+ Tile_X9Y14_LUT4AB/SS4BEG[12] Tile_X9Y14_LUT4AB/SS4BEG[13] Tile_X9Y14_LUT4AB/SS4BEG[14]
+ Tile_X9Y14_LUT4AB/SS4BEG[15] Tile_X9Y14_LUT4AB/SS4BEG[1] Tile_X9Y14_LUT4AB/SS4BEG[2]
+ Tile_X9Y14_LUT4AB/SS4BEG[3] Tile_X9Y14_LUT4AB/SS4BEG[4] Tile_X9Y14_LUT4AB/SS4BEG[5]
+ Tile_X9Y14_LUT4AB/SS4BEG[6] Tile_X9Y14_LUT4AB/SS4BEG[7] Tile_X9Y14_LUT4AB/SS4BEG[8]
+ Tile_X9Y14_LUT4AB/SS4BEG[9] Tile_X9Y14_LUT4AB/SS4END[0] Tile_X9Y14_LUT4AB/SS4END[10]
+ Tile_X9Y14_LUT4AB/SS4END[11] Tile_X9Y14_LUT4AB/SS4END[12] Tile_X9Y14_LUT4AB/SS4END[13]
+ Tile_X9Y14_LUT4AB/SS4END[14] Tile_X9Y14_LUT4AB/SS4END[15] Tile_X9Y14_LUT4AB/SS4END[1]
+ Tile_X9Y14_LUT4AB/SS4END[2] Tile_X9Y14_LUT4AB/SS4END[3] Tile_X9Y14_LUT4AB/SS4END[4]
+ Tile_X9Y14_LUT4AB/SS4END[5] Tile_X9Y14_LUT4AB/SS4END[6] Tile_X9Y14_LUT4AB/SS4END[7]
+ Tile_X9Y14_LUT4AB/SS4END[8] Tile_X9Y14_LUT4AB/SS4END[9] Tile_X9Y14_LUT4AB/UserCLK
+ Tile_X9Y13_LUT4AB/UserCLK VGND VPWR Tile_X9Y14_LUT4AB/W1BEG[0] Tile_X9Y14_LUT4AB/W1BEG[1]
+ Tile_X9Y14_LUT4AB/W1BEG[2] Tile_X9Y14_LUT4AB/W1BEG[3] Tile_X9Y14_LUT4AB/W1END[0]
+ Tile_X9Y14_LUT4AB/W1END[1] Tile_X9Y14_LUT4AB/W1END[2] Tile_X9Y14_LUT4AB/W1END[3]
+ Tile_X9Y14_LUT4AB/W2BEG[0] Tile_X9Y14_LUT4AB/W2BEG[1] Tile_X9Y14_LUT4AB/W2BEG[2]
+ Tile_X9Y14_LUT4AB/W2BEG[3] Tile_X9Y14_LUT4AB/W2BEG[4] Tile_X9Y14_LUT4AB/W2BEG[5]
+ Tile_X9Y14_LUT4AB/W2BEG[6] Tile_X9Y14_LUT4AB/W2BEG[7] Tile_X8Y14_LUT4AB/W2END[0]
+ Tile_X8Y14_LUT4AB/W2END[1] Tile_X8Y14_LUT4AB/W2END[2] Tile_X8Y14_LUT4AB/W2END[3]
+ Tile_X8Y14_LUT4AB/W2END[4] Tile_X8Y14_LUT4AB/W2END[5] Tile_X8Y14_LUT4AB/W2END[6]
+ Tile_X8Y14_LUT4AB/W2END[7] Tile_X9Y14_LUT4AB/W2END[0] Tile_X9Y14_LUT4AB/W2END[1]
+ Tile_X9Y14_LUT4AB/W2END[2] Tile_X9Y14_LUT4AB/W2END[3] Tile_X9Y14_LUT4AB/W2END[4]
+ Tile_X9Y14_LUT4AB/W2END[5] Tile_X9Y14_LUT4AB/W2END[6] Tile_X9Y14_LUT4AB/W2END[7]
+ Tile_X9Y14_LUT4AB/W2MID[0] Tile_X9Y14_LUT4AB/W2MID[1] Tile_X9Y14_LUT4AB/W2MID[2]
+ Tile_X9Y14_LUT4AB/W2MID[3] Tile_X9Y14_LUT4AB/W2MID[4] Tile_X9Y14_LUT4AB/W2MID[5]
+ Tile_X9Y14_LUT4AB/W2MID[6] Tile_X9Y14_LUT4AB/W2MID[7] Tile_X9Y14_LUT4AB/W6BEG[0]
+ Tile_X9Y14_LUT4AB/W6BEG[10] Tile_X9Y14_LUT4AB/W6BEG[11] Tile_X9Y14_LUT4AB/W6BEG[1]
+ Tile_X9Y14_LUT4AB/W6BEG[2] Tile_X9Y14_LUT4AB/W6BEG[3] Tile_X9Y14_LUT4AB/W6BEG[4]
+ Tile_X9Y14_LUT4AB/W6BEG[5] Tile_X9Y14_LUT4AB/W6BEG[6] Tile_X9Y14_LUT4AB/W6BEG[7]
+ Tile_X9Y14_LUT4AB/W6BEG[8] Tile_X9Y14_LUT4AB/W6BEG[9] Tile_X9Y14_LUT4AB/W6END[0]
+ Tile_X9Y14_LUT4AB/W6END[10] Tile_X9Y14_LUT4AB/W6END[11] Tile_X9Y14_LUT4AB/W6END[1]
+ Tile_X9Y14_LUT4AB/W6END[2] Tile_X9Y14_LUT4AB/W6END[3] Tile_X9Y14_LUT4AB/W6END[4]
+ Tile_X9Y14_LUT4AB/W6END[5] Tile_X9Y14_LUT4AB/W6END[6] Tile_X9Y14_LUT4AB/W6END[7]
+ Tile_X9Y14_LUT4AB/W6END[8] Tile_X9Y14_LUT4AB/W6END[9] Tile_X9Y14_LUT4AB/WW4BEG[0]
+ Tile_X9Y14_LUT4AB/WW4BEG[10] Tile_X9Y14_LUT4AB/WW4BEG[11] Tile_X9Y14_LUT4AB/WW4BEG[12]
+ Tile_X9Y14_LUT4AB/WW4BEG[13] Tile_X9Y14_LUT4AB/WW4BEG[14] Tile_X9Y14_LUT4AB/WW4BEG[15]
+ Tile_X9Y14_LUT4AB/WW4BEG[1] Tile_X9Y14_LUT4AB/WW4BEG[2] Tile_X9Y14_LUT4AB/WW4BEG[3]
+ Tile_X9Y14_LUT4AB/WW4BEG[4] Tile_X9Y14_LUT4AB/WW4BEG[5] Tile_X9Y14_LUT4AB/WW4BEG[6]
+ Tile_X9Y14_LUT4AB/WW4BEG[7] Tile_X9Y14_LUT4AB/WW4BEG[8] Tile_X9Y14_LUT4AB/WW4BEG[9]
+ Tile_X9Y14_LUT4AB/WW4END[0] Tile_X9Y14_LUT4AB/WW4END[10] Tile_X9Y14_LUT4AB/WW4END[11]
+ Tile_X9Y14_LUT4AB/WW4END[12] Tile_X9Y14_LUT4AB/WW4END[13] Tile_X9Y14_LUT4AB/WW4END[14]
+ Tile_X9Y14_LUT4AB/WW4END[15] Tile_X9Y14_LUT4AB/WW4END[1] Tile_X9Y14_LUT4AB/WW4END[2]
+ Tile_X9Y14_LUT4AB/WW4END[3] Tile_X9Y14_LUT4AB/WW4END[4] Tile_X9Y14_LUT4AB/WW4END[5]
+ Tile_X9Y14_LUT4AB/WW4END[6] Tile_X9Y14_LUT4AB/WW4END[7] Tile_X9Y14_LUT4AB/WW4END[8]
+ Tile_X9Y14_LUT4AB/WW4END[9] LUT4AB
XTile_X1Y1_LUT4AB Tile_X1Y2_LUT4AB/Co Tile_X1Y0_N_IO/Ci Tile_X2Y1_LUT4AB/E1END[0]
+ Tile_X2Y1_LUT4AB/E1END[1] Tile_X2Y1_LUT4AB/E1END[2] Tile_X2Y1_LUT4AB/E1END[3] Tile_X0Y1_W_IO/E1BEG[0]
+ Tile_X0Y1_W_IO/E1BEG[1] Tile_X0Y1_W_IO/E1BEG[2] Tile_X0Y1_W_IO/E1BEG[3] Tile_X2Y1_LUT4AB/E2MID[0]
+ Tile_X2Y1_LUT4AB/E2MID[1] Tile_X2Y1_LUT4AB/E2MID[2] Tile_X2Y1_LUT4AB/E2MID[3] Tile_X2Y1_LUT4AB/E2MID[4]
+ Tile_X2Y1_LUT4AB/E2MID[5] Tile_X2Y1_LUT4AB/E2MID[6] Tile_X2Y1_LUT4AB/E2MID[7] Tile_X2Y1_LUT4AB/E2END[0]
+ Tile_X2Y1_LUT4AB/E2END[1] Tile_X2Y1_LUT4AB/E2END[2] Tile_X2Y1_LUT4AB/E2END[3] Tile_X2Y1_LUT4AB/E2END[4]
+ Tile_X2Y1_LUT4AB/E2END[5] Tile_X2Y1_LUT4AB/E2END[6] Tile_X2Y1_LUT4AB/E2END[7] Tile_X0Y1_W_IO/E2BEGb[0]
+ Tile_X0Y1_W_IO/E2BEGb[1] Tile_X0Y1_W_IO/E2BEGb[2] Tile_X0Y1_W_IO/E2BEGb[3] Tile_X0Y1_W_IO/E2BEGb[4]
+ Tile_X0Y1_W_IO/E2BEGb[5] Tile_X0Y1_W_IO/E2BEGb[6] Tile_X0Y1_W_IO/E2BEGb[7] Tile_X0Y1_W_IO/E2BEG[0]
+ Tile_X0Y1_W_IO/E2BEG[1] Tile_X0Y1_W_IO/E2BEG[2] Tile_X0Y1_W_IO/E2BEG[3] Tile_X0Y1_W_IO/E2BEG[4]
+ Tile_X0Y1_W_IO/E2BEG[5] Tile_X0Y1_W_IO/E2BEG[6] Tile_X0Y1_W_IO/E2BEG[7] Tile_X2Y1_LUT4AB/E6END[0]
+ Tile_X2Y1_LUT4AB/E6END[10] Tile_X2Y1_LUT4AB/E6END[11] Tile_X2Y1_LUT4AB/E6END[1]
+ Tile_X2Y1_LUT4AB/E6END[2] Tile_X2Y1_LUT4AB/E6END[3] Tile_X2Y1_LUT4AB/E6END[4] Tile_X2Y1_LUT4AB/E6END[5]
+ Tile_X2Y1_LUT4AB/E6END[6] Tile_X2Y1_LUT4AB/E6END[7] Tile_X2Y1_LUT4AB/E6END[8] Tile_X2Y1_LUT4AB/E6END[9]
+ Tile_X0Y1_W_IO/E6BEG[0] Tile_X0Y1_W_IO/E6BEG[10] Tile_X0Y1_W_IO/E6BEG[11] Tile_X0Y1_W_IO/E6BEG[1]
+ Tile_X0Y1_W_IO/E6BEG[2] Tile_X0Y1_W_IO/E6BEG[3] Tile_X0Y1_W_IO/E6BEG[4] Tile_X0Y1_W_IO/E6BEG[5]
+ Tile_X0Y1_W_IO/E6BEG[6] Tile_X0Y1_W_IO/E6BEG[7] Tile_X0Y1_W_IO/E6BEG[8] Tile_X0Y1_W_IO/E6BEG[9]
+ Tile_X2Y1_LUT4AB/EE4END[0] Tile_X2Y1_LUT4AB/EE4END[10] Tile_X2Y1_LUT4AB/EE4END[11]
+ Tile_X2Y1_LUT4AB/EE4END[12] Tile_X2Y1_LUT4AB/EE4END[13] Tile_X2Y1_LUT4AB/EE4END[14]
+ Tile_X2Y1_LUT4AB/EE4END[15] Tile_X2Y1_LUT4AB/EE4END[1] Tile_X2Y1_LUT4AB/EE4END[2]
+ Tile_X2Y1_LUT4AB/EE4END[3] Tile_X2Y1_LUT4AB/EE4END[4] Tile_X2Y1_LUT4AB/EE4END[5]
+ Tile_X2Y1_LUT4AB/EE4END[6] Tile_X2Y1_LUT4AB/EE4END[7] Tile_X2Y1_LUT4AB/EE4END[8]
+ Tile_X2Y1_LUT4AB/EE4END[9] Tile_X0Y1_W_IO/EE4BEG[0] Tile_X0Y1_W_IO/EE4BEG[10] Tile_X0Y1_W_IO/EE4BEG[11]
+ Tile_X0Y1_W_IO/EE4BEG[12] Tile_X0Y1_W_IO/EE4BEG[13] Tile_X0Y1_W_IO/EE4BEG[14] Tile_X0Y1_W_IO/EE4BEG[15]
+ Tile_X0Y1_W_IO/EE4BEG[1] Tile_X0Y1_W_IO/EE4BEG[2] Tile_X0Y1_W_IO/EE4BEG[3] Tile_X0Y1_W_IO/EE4BEG[4]
+ Tile_X0Y1_W_IO/EE4BEG[5] Tile_X0Y1_W_IO/EE4BEG[6] Tile_X0Y1_W_IO/EE4BEG[7] Tile_X0Y1_W_IO/EE4BEG[8]
+ Tile_X0Y1_W_IO/EE4BEG[9] Tile_X1Y1_LUT4AB/FrameData[0] Tile_X1Y1_LUT4AB/FrameData[10]
+ Tile_X1Y1_LUT4AB/FrameData[11] Tile_X1Y1_LUT4AB/FrameData[12] Tile_X1Y1_LUT4AB/FrameData[13]
+ Tile_X1Y1_LUT4AB/FrameData[14] Tile_X1Y1_LUT4AB/FrameData[15] Tile_X1Y1_LUT4AB/FrameData[16]
+ Tile_X1Y1_LUT4AB/FrameData[17] Tile_X1Y1_LUT4AB/FrameData[18] Tile_X1Y1_LUT4AB/FrameData[19]
+ Tile_X1Y1_LUT4AB/FrameData[1] Tile_X1Y1_LUT4AB/FrameData[20] Tile_X1Y1_LUT4AB/FrameData[21]
+ Tile_X1Y1_LUT4AB/FrameData[22] Tile_X1Y1_LUT4AB/FrameData[23] Tile_X1Y1_LUT4AB/FrameData[24]
+ Tile_X1Y1_LUT4AB/FrameData[25] Tile_X1Y1_LUT4AB/FrameData[26] Tile_X1Y1_LUT4AB/FrameData[27]
+ Tile_X1Y1_LUT4AB/FrameData[28] Tile_X1Y1_LUT4AB/FrameData[29] Tile_X1Y1_LUT4AB/FrameData[2]
+ Tile_X1Y1_LUT4AB/FrameData[30] Tile_X1Y1_LUT4AB/FrameData[31] Tile_X1Y1_LUT4AB/FrameData[3]
+ Tile_X1Y1_LUT4AB/FrameData[4] Tile_X1Y1_LUT4AB/FrameData[5] Tile_X1Y1_LUT4AB/FrameData[6]
+ Tile_X1Y1_LUT4AB/FrameData[7] Tile_X1Y1_LUT4AB/FrameData[8] Tile_X1Y1_LUT4AB/FrameData[9]
+ Tile_X2Y1_LUT4AB/FrameData[0] Tile_X2Y1_LUT4AB/FrameData[10] Tile_X2Y1_LUT4AB/FrameData[11]
+ Tile_X2Y1_LUT4AB/FrameData[12] Tile_X2Y1_LUT4AB/FrameData[13] Tile_X2Y1_LUT4AB/FrameData[14]
+ Tile_X2Y1_LUT4AB/FrameData[15] Tile_X2Y1_LUT4AB/FrameData[16] Tile_X2Y1_LUT4AB/FrameData[17]
+ Tile_X2Y1_LUT4AB/FrameData[18] Tile_X2Y1_LUT4AB/FrameData[19] Tile_X2Y1_LUT4AB/FrameData[1]
+ Tile_X2Y1_LUT4AB/FrameData[20] Tile_X2Y1_LUT4AB/FrameData[21] Tile_X2Y1_LUT4AB/FrameData[22]
+ Tile_X2Y1_LUT4AB/FrameData[23] Tile_X2Y1_LUT4AB/FrameData[24] Tile_X2Y1_LUT4AB/FrameData[25]
+ Tile_X2Y1_LUT4AB/FrameData[26] Tile_X2Y1_LUT4AB/FrameData[27] Tile_X2Y1_LUT4AB/FrameData[28]
+ Tile_X2Y1_LUT4AB/FrameData[29] Tile_X2Y1_LUT4AB/FrameData[2] Tile_X2Y1_LUT4AB/FrameData[30]
+ Tile_X2Y1_LUT4AB/FrameData[31] Tile_X2Y1_LUT4AB/FrameData[3] Tile_X2Y1_LUT4AB/FrameData[4]
+ Tile_X2Y1_LUT4AB/FrameData[5] Tile_X2Y1_LUT4AB/FrameData[6] Tile_X2Y1_LUT4AB/FrameData[7]
+ Tile_X2Y1_LUT4AB/FrameData[8] Tile_X2Y1_LUT4AB/FrameData[9] Tile_X1Y1_LUT4AB/FrameStrobe[0]
+ Tile_X1Y1_LUT4AB/FrameStrobe[10] Tile_X1Y1_LUT4AB/FrameStrobe[11] Tile_X1Y1_LUT4AB/FrameStrobe[12]
+ Tile_X1Y1_LUT4AB/FrameStrobe[13] Tile_X1Y1_LUT4AB/FrameStrobe[14] Tile_X1Y1_LUT4AB/FrameStrobe[15]
+ Tile_X1Y1_LUT4AB/FrameStrobe[16] Tile_X1Y1_LUT4AB/FrameStrobe[17] Tile_X1Y1_LUT4AB/FrameStrobe[18]
+ Tile_X1Y1_LUT4AB/FrameStrobe[19] Tile_X1Y1_LUT4AB/FrameStrobe[1] Tile_X1Y1_LUT4AB/FrameStrobe[2]
+ Tile_X1Y1_LUT4AB/FrameStrobe[3] Tile_X1Y1_LUT4AB/FrameStrobe[4] Tile_X1Y1_LUT4AB/FrameStrobe[5]
+ Tile_X1Y1_LUT4AB/FrameStrobe[6] Tile_X1Y1_LUT4AB/FrameStrobe[7] Tile_X1Y1_LUT4AB/FrameStrobe[8]
+ Tile_X1Y1_LUT4AB/FrameStrobe[9] Tile_X1Y0_N_IO/FrameStrobe[0] Tile_X1Y0_N_IO/FrameStrobe[10]
+ Tile_X1Y0_N_IO/FrameStrobe[11] Tile_X1Y0_N_IO/FrameStrobe[12] Tile_X1Y0_N_IO/FrameStrobe[13]
+ Tile_X1Y0_N_IO/FrameStrobe[14] Tile_X1Y0_N_IO/FrameStrobe[15] Tile_X1Y0_N_IO/FrameStrobe[16]
+ Tile_X1Y0_N_IO/FrameStrobe[17] Tile_X1Y0_N_IO/FrameStrobe[18] Tile_X1Y0_N_IO/FrameStrobe[19]
+ Tile_X1Y0_N_IO/FrameStrobe[1] Tile_X1Y0_N_IO/FrameStrobe[2] Tile_X1Y0_N_IO/FrameStrobe[3]
+ Tile_X1Y0_N_IO/FrameStrobe[4] Tile_X1Y0_N_IO/FrameStrobe[5] Tile_X1Y0_N_IO/FrameStrobe[6]
+ Tile_X1Y0_N_IO/FrameStrobe[7] Tile_X1Y0_N_IO/FrameStrobe[8] Tile_X1Y0_N_IO/FrameStrobe[9]
+ Tile_X1Y0_N_IO/N1END[0] Tile_X1Y0_N_IO/N1END[1] Tile_X1Y0_N_IO/N1END[2] Tile_X1Y0_N_IO/N1END[3]
+ Tile_X1Y2_LUT4AB/N1BEG[0] Tile_X1Y2_LUT4AB/N1BEG[1] Tile_X1Y2_LUT4AB/N1BEG[2] Tile_X1Y2_LUT4AB/N1BEG[3]
+ Tile_X1Y0_N_IO/N2MID[0] Tile_X1Y0_N_IO/N2MID[1] Tile_X1Y0_N_IO/N2MID[2] Tile_X1Y0_N_IO/N2MID[3]
+ Tile_X1Y0_N_IO/N2MID[4] Tile_X1Y0_N_IO/N2MID[5] Tile_X1Y0_N_IO/N2MID[6] Tile_X1Y0_N_IO/N2MID[7]
+ Tile_X1Y0_N_IO/N2END[0] Tile_X1Y0_N_IO/N2END[1] Tile_X1Y0_N_IO/N2END[2] Tile_X1Y0_N_IO/N2END[3]
+ Tile_X1Y0_N_IO/N2END[4] Tile_X1Y0_N_IO/N2END[5] Tile_X1Y0_N_IO/N2END[6] Tile_X1Y0_N_IO/N2END[7]
+ Tile_X1Y1_LUT4AB/N2END[0] Tile_X1Y1_LUT4AB/N2END[1] Tile_X1Y1_LUT4AB/N2END[2] Tile_X1Y1_LUT4AB/N2END[3]
+ Tile_X1Y1_LUT4AB/N2END[4] Tile_X1Y1_LUT4AB/N2END[5] Tile_X1Y1_LUT4AB/N2END[6] Tile_X1Y1_LUT4AB/N2END[7]
+ Tile_X1Y2_LUT4AB/N2BEG[0] Tile_X1Y2_LUT4AB/N2BEG[1] Tile_X1Y2_LUT4AB/N2BEG[2] Tile_X1Y2_LUT4AB/N2BEG[3]
+ Tile_X1Y2_LUT4AB/N2BEG[4] Tile_X1Y2_LUT4AB/N2BEG[5] Tile_X1Y2_LUT4AB/N2BEG[6] Tile_X1Y2_LUT4AB/N2BEG[7]
+ Tile_X1Y0_N_IO/N4END[0] Tile_X1Y0_N_IO/N4END[10] Tile_X1Y0_N_IO/N4END[11] Tile_X1Y0_N_IO/N4END[12]
+ Tile_X1Y0_N_IO/N4END[13] Tile_X1Y0_N_IO/N4END[14] Tile_X1Y0_N_IO/N4END[15] Tile_X1Y0_N_IO/N4END[1]
+ Tile_X1Y0_N_IO/N4END[2] Tile_X1Y0_N_IO/N4END[3] Tile_X1Y0_N_IO/N4END[4] Tile_X1Y0_N_IO/N4END[5]
+ Tile_X1Y0_N_IO/N4END[6] Tile_X1Y0_N_IO/N4END[7] Tile_X1Y0_N_IO/N4END[8] Tile_X1Y0_N_IO/N4END[9]
+ Tile_X1Y2_LUT4AB/N4BEG[0] Tile_X1Y2_LUT4AB/N4BEG[10] Tile_X1Y2_LUT4AB/N4BEG[11]
+ Tile_X1Y2_LUT4AB/N4BEG[12] Tile_X1Y2_LUT4AB/N4BEG[13] Tile_X1Y2_LUT4AB/N4BEG[14]
+ Tile_X1Y2_LUT4AB/N4BEG[15] Tile_X1Y2_LUT4AB/N4BEG[1] Tile_X1Y2_LUT4AB/N4BEG[2] Tile_X1Y2_LUT4AB/N4BEG[3]
+ Tile_X1Y2_LUT4AB/N4BEG[4] Tile_X1Y2_LUT4AB/N4BEG[5] Tile_X1Y2_LUT4AB/N4BEG[6] Tile_X1Y2_LUT4AB/N4BEG[7]
+ Tile_X1Y2_LUT4AB/N4BEG[8] Tile_X1Y2_LUT4AB/N4BEG[9] Tile_X1Y0_N_IO/NN4END[0] Tile_X1Y0_N_IO/NN4END[10]
+ Tile_X1Y0_N_IO/NN4END[11] Tile_X1Y0_N_IO/NN4END[12] Tile_X1Y0_N_IO/NN4END[13] Tile_X1Y0_N_IO/NN4END[14]
+ Tile_X1Y0_N_IO/NN4END[15] Tile_X1Y0_N_IO/NN4END[1] Tile_X1Y0_N_IO/NN4END[2] Tile_X1Y0_N_IO/NN4END[3]
+ Tile_X1Y0_N_IO/NN4END[4] Tile_X1Y0_N_IO/NN4END[5] Tile_X1Y0_N_IO/NN4END[6] Tile_X1Y0_N_IO/NN4END[7]
+ Tile_X1Y0_N_IO/NN4END[8] Tile_X1Y0_N_IO/NN4END[9] Tile_X1Y2_LUT4AB/NN4BEG[0] Tile_X1Y2_LUT4AB/NN4BEG[10]
+ Tile_X1Y2_LUT4AB/NN4BEG[11] Tile_X1Y2_LUT4AB/NN4BEG[12] Tile_X1Y2_LUT4AB/NN4BEG[13]
+ Tile_X1Y2_LUT4AB/NN4BEG[14] Tile_X1Y2_LUT4AB/NN4BEG[15] Tile_X1Y2_LUT4AB/NN4BEG[1]
+ Tile_X1Y2_LUT4AB/NN4BEG[2] Tile_X1Y2_LUT4AB/NN4BEG[3] Tile_X1Y2_LUT4AB/NN4BEG[4]
+ Tile_X1Y2_LUT4AB/NN4BEG[5] Tile_X1Y2_LUT4AB/NN4BEG[6] Tile_X1Y2_LUT4AB/NN4BEG[7]
+ Tile_X1Y2_LUT4AB/NN4BEG[8] Tile_X1Y2_LUT4AB/NN4BEG[9] Tile_X1Y2_LUT4AB/S1END[0]
+ Tile_X1Y2_LUT4AB/S1END[1] Tile_X1Y2_LUT4AB/S1END[2] Tile_X1Y2_LUT4AB/S1END[3] Tile_X1Y0_N_IO/S1BEG[0]
+ Tile_X1Y0_N_IO/S1BEG[1] Tile_X1Y0_N_IO/S1BEG[2] Tile_X1Y0_N_IO/S1BEG[3] Tile_X1Y2_LUT4AB/S2MID[0]
+ Tile_X1Y2_LUT4AB/S2MID[1] Tile_X1Y2_LUT4AB/S2MID[2] Tile_X1Y2_LUT4AB/S2MID[3] Tile_X1Y2_LUT4AB/S2MID[4]
+ Tile_X1Y2_LUT4AB/S2MID[5] Tile_X1Y2_LUT4AB/S2MID[6] Tile_X1Y2_LUT4AB/S2MID[7] Tile_X1Y2_LUT4AB/S2END[0]
+ Tile_X1Y2_LUT4AB/S2END[1] Tile_X1Y2_LUT4AB/S2END[2] Tile_X1Y2_LUT4AB/S2END[3] Tile_X1Y2_LUT4AB/S2END[4]
+ Tile_X1Y2_LUT4AB/S2END[5] Tile_X1Y2_LUT4AB/S2END[6] Tile_X1Y2_LUT4AB/S2END[7] Tile_X1Y0_N_IO/S2BEGb[0]
+ Tile_X1Y0_N_IO/S2BEGb[1] Tile_X1Y0_N_IO/S2BEGb[2] Tile_X1Y0_N_IO/S2BEGb[3] Tile_X1Y0_N_IO/S2BEGb[4]
+ Tile_X1Y0_N_IO/S2BEGb[5] Tile_X1Y0_N_IO/S2BEGb[6] Tile_X1Y0_N_IO/S2BEGb[7] Tile_X1Y0_N_IO/S2BEG[0]
+ Tile_X1Y0_N_IO/S2BEG[1] Tile_X1Y0_N_IO/S2BEG[2] Tile_X1Y0_N_IO/S2BEG[3] Tile_X1Y0_N_IO/S2BEG[4]
+ Tile_X1Y0_N_IO/S2BEG[5] Tile_X1Y0_N_IO/S2BEG[6] Tile_X1Y0_N_IO/S2BEG[7] Tile_X1Y2_LUT4AB/S4END[0]
+ Tile_X1Y2_LUT4AB/S4END[10] Tile_X1Y2_LUT4AB/S4END[11] Tile_X1Y2_LUT4AB/S4END[12]
+ Tile_X1Y2_LUT4AB/S4END[13] Tile_X1Y2_LUT4AB/S4END[14] Tile_X1Y2_LUT4AB/S4END[15]
+ Tile_X1Y2_LUT4AB/S4END[1] Tile_X1Y2_LUT4AB/S4END[2] Tile_X1Y2_LUT4AB/S4END[3] Tile_X1Y2_LUT4AB/S4END[4]
+ Tile_X1Y2_LUT4AB/S4END[5] Tile_X1Y2_LUT4AB/S4END[6] Tile_X1Y2_LUT4AB/S4END[7] Tile_X1Y2_LUT4AB/S4END[8]
+ Tile_X1Y2_LUT4AB/S4END[9] Tile_X1Y0_N_IO/S4BEG[0] Tile_X1Y0_N_IO/S4BEG[10] Tile_X1Y0_N_IO/S4BEG[11]
+ Tile_X1Y0_N_IO/S4BEG[12] Tile_X1Y0_N_IO/S4BEG[13] Tile_X1Y0_N_IO/S4BEG[14] Tile_X1Y0_N_IO/S4BEG[15]
+ Tile_X1Y0_N_IO/S4BEG[1] Tile_X1Y0_N_IO/S4BEG[2] Tile_X1Y0_N_IO/S4BEG[3] Tile_X1Y0_N_IO/S4BEG[4]
+ Tile_X1Y0_N_IO/S4BEG[5] Tile_X1Y0_N_IO/S4BEG[6] Tile_X1Y0_N_IO/S4BEG[7] Tile_X1Y0_N_IO/S4BEG[8]
+ Tile_X1Y0_N_IO/S4BEG[9] Tile_X1Y2_LUT4AB/SS4END[0] Tile_X1Y2_LUT4AB/SS4END[10] Tile_X1Y2_LUT4AB/SS4END[11]
+ Tile_X1Y2_LUT4AB/SS4END[12] Tile_X1Y2_LUT4AB/SS4END[13] Tile_X1Y2_LUT4AB/SS4END[14]
+ Tile_X1Y2_LUT4AB/SS4END[15] Tile_X1Y2_LUT4AB/SS4END[1] Tile_X1Y2_LUT4AB/SS4END[2]
+ Tile_X1Y2_LUT4AB/SS4END[3] Tile_X1Y2_LUT4AB/SS4END[4] Tile_X1Y2_LUT4AB/SS4END[5]
+ Tile_X1Y2_LUT4AB/SS4END[6] Tile_X1Y2_LUT4AB/SS4END[7] Tile_X1Y2_LUT4AB/SS4END[8]
+ Tile_X1Y2_LUT4AB/SS4END[9] Tile_X1Y0_N_IO/SS4BEG[0] Tile_X1Y0_N_IO/SS4BEG[10] Tile_X1Y0_N_IO/SS4BEG[11]
+ Tile_X1Y0_N_IO/SS4BEG[12] Tile_X1Y0_N_IO/SS4BEG[13] Tile_X1Y0_N_IO/SS4BEG[14] Tile_X1Y0_N_IO/SS4BEG[15]
+ Tile_X1Y0_N_IO/SS4BEG[1] Tile_X1Y0_N_IO/SS4BEG[2] Tile_X1Y0_N_IO/SS4BEG[3] Tile_X1Y0_N_IO/SS4BEG[4]
+ Tile_X1Y0_N_IO/SS4BEG[5] Tile_X1Y0_N_IO/SS4BEG[6] Tile_X1Y0_N_IO/SS4BEG[7] Tile_X1Y0_N_IO/SS4BEG[8]
+ Tile_X1Y0_N_IO/SS4BEG[9] Tile_X1Y1_LUT4AB/UserCLK Tile_X1Y0_N_IO/UserCLK VGND VPWR
+ Tile_X0Y1_W_IO/W1END[0] Tile_X0Y1_W_IO/W1END[1] Tile_X0Y1_W_IO/W1END[2] Tile_X0Y1_W_IO/W1END[3]
+ Tile_X2Y1_LUT4AB/W1BEG[0] Tile_X2Y1_LUT4AB/W1BEG[1] Tile_X2Y1_LUT4AB/W1BEG[2] Tile_X2Y1_LUT4AB/W1BEG[3]
+ Tile_X0Y1_W_IO/W2MID[0] Tile_X0Y1_W_IO/W2MID[1] Tile_X0Y1_W_IO/W2MID[2] Tile_X0Y1_W_IO/W2MID[3]
+ Tile_X0Y1_W_IO/W2MID[4] Tile_X0Y1_W_IO/W2MID[5] Tile_X0Y1_W_IO/W2MID[6] Tile_X0Y1_W_IO/W2MID[7]
+ Tile_X0Y1_W_IO/W2END[0] Tile_X0Y1_W_IO/W2END[1] Tile_X0Y1_W_IO/W2END[2] Tile_X0Y1_W_IO/W2END[3]
+ Tile_X0Y1_W_IO/W2END[4] Tile_X0Y1_W_IO/W2END[5] Tile_X0Y1_W_IO/W2END[6] Tile_X0Y1_W_IO/W2END[7]
+ Tile_X1Y1_LUT4AB/W2END[0] Tile_X1Y1_LUT4AB/W2END[1] Tile_X1Y1_LUT4AB/W2END[2] Tile_X1Y1_LUT4AB/W2END[3]
+ Tile_X1Y1_LUT4AB/W2END[4] Tile_X1Y1_LUT4AB/W2END[5] Tile_X1Y1_LUT4AB/W2END[6] Tile_X1Y1_LUT4AB/W2END[7]
+ Tile_X2Y1_LUT4AB/W2BEG[0] Tile_X2Y1_LUT4AB/W2BEG[1] Tile_X2Y1_LUT4AB/W2BEG[2] Tile_X2Y1_LUT4AB/W2BEG[3]
+ Tile_X2Y1_LUT4AB/W2BEG[4] Tile_X2Y1_LUT4AB/W2BEG[5] Tile_X2Y1_LUT4AB/W2BEG[6] Tile_X2Y1_LUT4AB/W2BEG[7]
+ Tile_X0Y1_W_IO/W6END[0] Tile_X0Y1_W_IO/W6END[10] Tile_X0Y1_W_IO/W6END[11] Tile_X0Y1_W_IO/W6END[1]
+ Tile_X0Y1_W_IO/W6END[2] Tile_X0Y1_W_IO/W6END[3] Tile_X0Y1_W_IO/W6END[4] Tile_X0Y1_W_IO/W6END[5]
+ Tile_X0Y1_W_IO/W6END[6] Tile_X0Y1_W_IO/W6END[7] Tile_X0Y1_W_IO/W6END[8] Tile_X0Y1_W_IO/W6END[9]
+ Tile_X2Y1_LUT4AB/W6BEG[0] Tile_X2Y1_LUT4AB/W6BEG[10] Tile_X2Y1_LUT4AB/W6BEG[11]
+ Tile_X2Y1_LUT4AB/W6BEG[1] Tile_X2Y1_LUT4AB/W6BEG[2] Tile_X2Y1_LUT4AB/W6BEG[3] Tile_X2Y1_LUT4AB/W6BEG[4]
+ Tile_X2Y1_LUT4AB/W6BEG[5] Tile_X2Y1_LUT4AB/W6BEG[6] Tile_X2Y1_LUT4AB/W6BEG[7] Tile_X2Y1_LUT4AB/W6BEG[8]
+ Tile_X2Y1_LUT4AB/W6BEG[9] Tile_X0Y1_W_IO/WW4END[0] Tile_X0Y1_W_IO/WW4END[10] Tile_X0Y1_W_IO/WW4END[11]
+ Tile_X0Y1_W_IO/WW4END[12] Tile_X0Y1_W_IO/WW4END[13] Tile_X0Y1_W_IO/WW4END[14] Tile_X0Y1_W_IO/WW4END[15]
+ Tile_X0Y1_W_IO/WW4END[1] Tile_X0Y1_W_IO/WW4END[2] Tile_X0Y1_W_IO/WW4END[3] Tile_X0Y1_W_IO/WW4END[4]
+ Tile_X0Y1_W_IO/WW4END[5] Tile_X0Y1_W_IO/WW4END[6] Tile_X0Y1_W_IO/WW4END[7] Tile_X0Y1_W_IO/WW4END[8]
+ Tile_X0Y1_W_IO/WW4END[9] Tile_X2Y1_LUT4AB/WW4BEG[0] Tile_X2Y1_LUT4AB/WW4BEG[10]
+ Tile_X2Y1_LUT4AB/WW4BEG[11] Tile_X2Y1_LUT4AB/WW4BEG[12] Tile_X2Y1_LUT4AB/WW4BEG[13]
+ Tile_X2Y1_LUT4AB/WW4BEG[14] Tile_X2Y1_LUT4AB/WW4BEG[15] Tile_X2Y1_LUT4AB/WW4BEG[1]
+ Tile_X2Y1_LUT4AB/WW4BEG[2] Tile_X2Y1_LUT4AB/WW4BEG[3] Tile_X2Y1_LUT4AB/WW4BEG[4]
+ Tile_X2Y1_LUT4AB/WW4BEG[5] Tile_X2Y1_LUT4AB/WW4BEG[6] Tile_X2Y1_LUT4AB/WW4BEG[7]
+ Tile_X2Y1_LUT4AB/WW4BEG[8] Tile_X2Y1_LUT4AB/WW4BEG[9] LUT4AB
XTile_X4Y6_RegFile Tile_X5Y6_LUT4AB/E1END[0] Tile_X5Y6_LUT4AB/E1END[1] Tile_X5Y6_LUT4AB/E1END[2]
+ Tile_X5Y6_LUT4AB/E1END[3] Tile_X3Y6_LUT4AB/E1BEG[0] Tile_X3Y6_LUT4AB/E1BEG[1] Tile_X3Y6_LUT4AB/E1BEG[2]
+ Tile_X3Y6_LUT4AB/E1BEG[3] Tile_X5Y6_LUT4AB/E2MID[0] Tile_X5Y6_LUT4AB/E2MID[1] Tile_X5Y6_LUT4AB/E2MID[2]
+ Tile_X5Y6_LUT4AB/E2MID[3] Tile_X5Y6_LUT4AB/E2MID[4] Tile_X5Y6_LUT4AB/E2MID[5] Tile_X5Y6_LUT4AB/E2MID[6]
+ Tile_X5Y6_LUT4AB/E2MID[7] Tile_X5Y6_LUT4AB/E2END[0] Tile_X5Y6_LUT4AB/E2END[1] Tile_X5Y6_LUT4AB/E2END[2]
+ Tile_X5Y6_LUT4AB/E2END[3] Tile_X5Y6_LUT4AB/E2END[4] Tile_X5Y6_LUT4AB/E2END[5] Tile_X5Y6_LUT4AB/E2END[6]
+ Tile_X5Y6_LUT4AB/E2END[7] Tile_X4Y6_RegFile/E2END[0] Tile_X4Y6_RegFile/E2END[1]
+ Tile_X4Y6_RegFile/E2END[2] Tile_X4Y6_RegFile/E2END[3] Tile_X4Y6_RegFile/E2END[4]
+ Tile_X4Y6_RegFile/E2END[5] Tile_X4Y6_RegFile/E2END[6] Tile_X4Y6_RegFile/E2END[7]
+ Tile_X3Y6_LUT4AB/E2BEG[0] Tile_X3Y6_LUT4AB/E2BEG[1] Tile_X3Y6_LUT4AB/E2BEG[2] Tile_X3Y6_LUT4AB/E2BEG[3]
+ Tile_X3Y6_LUT4AB/E2BEG[4] Tile_X3Y6_LUT4AB/E2BEG[5] Tile_X3Y6_LUT4AB/E2BEG[6] Tile_X3Y6_LUT4AB/E2BEG[7]
+ Tile_X5Y6_LUT4AB/E6END[0] Tile_X5Y6_LUT4AB/E6END[10] Tile_X5Y6_LUT4AB/E6END[11]
+ Tile_X5Y6_LUT4AB/E6END[1] Tile_X5Y6_LUT4AB/E6END[2] Tile_X5Y6_LUT4AB/E6END[3] Tile_X5Y6_LUT4AB/E6END[4]
+ Tile_X5Y6_LUT4AB/E6END[5] Tile_X5Y6_LUT4AB/E6END[6] Tile_X5Y6_LUT4AB/E6END[7] Tile_X5Y6_LUT4AB/E6END[8]
+ Tile_X5Y6_LUT4AB/E6END[9] Tile_X3Y6_LUT4AB/E6BEG[0] Tile_X3Y6_LUT4AB/E6BEG[10] Tile_X3Y6_LUT4AB/E6BEG[11]
+ Tile_X3Y6_LUT4AB/E6BEG[1] Tile_X3Y6_LUT4AB/E6BEG[2] Tile_X3Y6_LUT4AB/E6BEG[3] Tile_X3Y6_LUT4AB/E6BEG[4]
+ Tile_X3Y6_LUT4AB/E6BEG[5] Tile_X3Y6_LUT4AB/E6BEG[6] Tile_X3Y6_LUT4AB/E6BEG[7] Tile_X3Y6_LUT4AB/E6BEG[8]
+ Tile_X3Y6_LUT4AB/E6BEG[9] Tile_X5Y6_LUT4AB/EE4END[0] Tile_X5Y6_LUT4AB/EE4END[10]
+ Tile_X5Y6_LUT4AB/EE4END[11] Tile_X5Y6_LUT4AB/EE4END[12] Tile_X5Y6_LUT4AB/EE4END[13]
+ Tile_X5Y6_LUT4AB/EE4END[14] Tile_X5Y6_LUT4AB/EE4END[15] Tile_X5Y6_LUT4AB/EE4END[1]
+ Tile_X5Y6_LUT4AB/EE4END[2] Tile_X5Y6_LUT4AB/EE4END[3] Tile_X5Y6_LUT4AB/EE4END[4]
+ Tile_X5Y6_LUT4AB/EE4END[5] Tile_X5Y6_LUT4AB/EE4END[6] Tile_X5Y6_LUT4AB/EE4END[7]
+ Tile_X5Y6_LUT4AB/EE4END[8] Tile_X5Y6_LUT4AB/EE4END[9] Tile_X3Y6_LUT4AB/EE4BEG[0]
+ Tile_X3Y6_LUT4AB/EE4BEG[10] Tile_X3Y6_LUT4AB/EE4BEG[11] Tile_X3Y6_LUT4AB/EE4BEG[12]
+ Tile_X3Y6_LUT4AB/EE4BEG[13] Tile_X3Y6_LUT4AB/EE4BEG[14] Tile_X3Y6_LUT4AB/EE4BEG[15]
+ Tile_X3Y6_LUT4AB/EE4BEG[1] Tile_X3Y6_LUT4AB/EE4BEG[2] Tile_X3Y6_LUT4AB/EE4BEG[3]
+ Tile_X3Y6_LUT4AB/EE4BEG[4] Tile_X3Y6_LUT4AB/EE4BEG[5] Tile_X3Y6_LUT4AB/EE4BEG[6]
+ Tile_X3Y6_LUT4AB/EE4BEG[7] Tile_X3Y6_LUT4AB/EE4BEG[8] Tile_X3Y6_LUT4AB/EE4BEG[9]
+ Tile_X4Y6_RegFile/FrameData[0] Tile_X4Y6_RegFile/FrameData[10] Tile_X4Y6_RegFile/FrameData[11]
+ Tile_X4Y6_RegFile/FrameData[12] Tile_X4Y6_RegFile/FrameData[13] Tile_X4Y6_RegFile/FrameData[14]
+ Tile_X4Y6_RegFile/FrameData[15] Tile_X4Y6_RegFile/FrameData[16] Tile_X4Y6_RegFile/FrameData[17]
+ Tile_X4Y6_RegFile/FrameData[18] Tile_X4Y6_RegFile/FrameData[19] Tile_X4Y6_RegFile/FrameData[1]
+ Tile_X4Y6_RegFile/FrameData[20] Tile_X4Y6_RegFile/FrameData[21] Tile_X4Y6_RegFile/FrameData[22]
+ Tile_X4Y6_RegFile/FrameData[23] Tile_X4Y6_RegFile/FrameData[24] Tile_X4Y6_RegFile/FrameData[25]
+ Tile_X4Y6_RegFile/FrameData[26] Tile_X4Y6_RegFile/FrameData[27] Tile_X4Y6_RegFile/FrameData[28]
+ Tile_X4Y6_RegFile/FrameData[29] Tile_X4Y6_RegFile/FrameData[2] Tile_X4Y6_RegFile/FrameData[30]
+ Tile_X4Y6_RegFile/FrameData[31] Tile_X4Y6_RegFile/FrameData[3] Tile_X4Y6_RegFile/FrameData[4]
+ Tile_X4Y6_RegFile/FrameData[5] Tile_X4Y6_RegFile/FrameData[6] Tile_X4Y6_RegFile/FrameData[7]
+ Tile_X4Y6_RegFile/FrameData[8] Tile_X4Y6_RegFile/FrameData[9] Tile_X5Y6_LUT4AB/FrameData[0]
+ Tile_X5Y6_LUT4AB/FrameData[10] Tile_X5Y6_LUT4AB/FrameData[11] Tile_X5Y6_LUT4AB/FrameData[12]
+ Tile_X5Y6_LUT4AB/FrameData[13] Tile_X5Y6_LUT4AB/FrameData[14] Tile_X5Y6_LUT4AB/FrameData[15]
+ Tile_X5Y6_LUT4AB/FrameData[16] Tile_X5Y6_LUT4AB/FrameData[17] Tile_X5Y6_LUT4AB/FrameData[18]
+ Tile_X5Y6_LUT4AB/FrameData[19] Tile_X5Y6_LUT4AB/FrameData[1] Tile_X5Y6_LUT4AB/FrameData[20]
+ Tile_X5Y6_LUT4AB/FrameData[21] Tile_X5Y6_LUT4AB/FrameData[22] Tile_X5Y6_LUT4AB/FrameData[23]
+ Tile_X5Y6_LUT4AB/FrameData[24] Tile_X5Y6_LUT4AB/FrameData[25] Tile_X5Y6_LUT4AB/FrameData[26]
+ Tile_X5Y6_LUT4AB/FrameData[27] Tile_X5Y6_LUT4AB/FrameData[28] Tile_X5Y6_LUT4AB/FrameData[29]
+ Tile_X5Y6_LUT4AB/FrameData[2] Tile_X5Y6_LUT4AB/FrameData[30] Tile_X5Y6_LUT4AB/FrameData[31]
+ Tile_X5Y6_LUT4AB/FrameData[3] Tile_X5Y6_LUT4AB/FrameData[4] Tile_X5Y6_LUT4AB/FrameData[5]
+ Tile_X5Y6_LUT4AB/FrameData[6] Tile_X5Y6_LUT4AB/FrameData[7] Tile_X5Y6_LUT4AB/FrameData[8]
+ Tile_X5Y6_LUT4AB/FrameData[9] Tile_X4Y6_RegFile/FrameStrobe[0] Tile_X4Y6_RegFile/FrameStrobe[10]
+ Tile_X4Y6_RegFile/FrameStrobe[11] Tile_X4Y6_RegFile/FrameStrobe[12] Tile_X4Y6_RegFile/FrameStrobe[13]
+ Tile_X4Y6_RegFile/FrameStrobe[14] Tile_X4Y6_RegFile/FrameStrobe[15] Tile_X4Y6_RegFile/FrameStrobe[16]
+ Tile_X4Y6_RegFile/FrameStrobe[17] Tile_X4Y6_RegFile/FrameStrobe[18] Tile_X4Y6_RegFile/FrameStrobe[19]
+ Tile_X4Y6_RegFile/FrameStrobe[1] Tile_X4Y6_RegFile/FrameStrobe[2] Tile_X4Y6_RegFile/FrameStrobe[3]
+ Tile_X4Y6_RegFile/FrameStrobe[4] Tile_X4Y6_RegFile/FrameStrobe[5] Tile_X4Y6_RegFile/FrameStrobe[6]
+ Tile_X4Y6_RegFile/FrameStrobe[7] Tile_X4Y6_RegFile/FrameStrobe[8] Tile_X4Y6_RegFile/FrameStrobe[9]
+ Tile_X4Y5_RegFile/FrameStrobe[0] Tile_X4Y5_RegFile/FrameStrobe[10] Tile_X4Y5_RegFile/FrameStrobe[11]
+ Tile_X4Y5_RegFile/FrameStrobe[12] Tile_X4Y5_RegFile/FrameStrobe[13] Tile_X4Y5_RegFile/FrameStrobe[14]
+ Tile_X4Y5_RegFile/FrameStrobe[15] Tile_X4Y5_RegFile/FrameStrobe[16] Tile_X4Y5_RegFile/FrameStrobe[17]
+ Tile_X4Y5_RegFile/FrameStrobe[18] Tile_X4Y5_RegFile/FrameStrobe[19] Tile_X4Y5_RegFile/FrameStrobe[1]
+ Tile_X4Y5_RegFile/FrameStrobe[2] Tile_X4Y5_RegFile/FrameStrobe[3] Tile_X4Y5_RegFile/FrameStrobe[4]
+ Tile_X4Y5_RegFile/FrameStrobe[5] Tile_X4Y5_RegFile/FrameStrobe[6] Tile_X4Y5_RegFile/FrameStrobe[7]
+ Tile_X4Y5_RegFile/FrameStrobe[8] Tile_X4Y5_RegFile/FrameStrobe[9] Tile_X4Y6_RegFile/N1BEG[0]
+ Tile_X4Y6_RegFile/N1BEG[1] Tile_X4Y6_RegFile/N1BEG[2] Tile_X4Y6_RegFile/N1BEG[3]
+ Tile_X4Y7_RegFile/N1BEG[0] Tile_X4Y7_RegFile/N1BEG[1] Tile_X4Y7_RegFile/N1BEG[2]
+ Tile_X4Y7_RegFile/N1BEG[3] Tile_X4Y6_RegFile/N2BEG[0] Tile_X4Y6_RegFile/N2BEG[1]
+ Tile_X4Y6_RegFile/N2BEG[2] Tile_X4Y6_RegFile/N2BEG[3] Tile_X4Y6_RegFile/N2BEG[4]
+ Tile_X4Y6_RegFile/N2BEG[5] Tile_X4Y6_RegFile/N2BEG[6] Tile_X4Y6_RegFile/N2BEG[7]
+ Tile_X4Y5_RegFile/N2END[0] Tile_X4Y5_RegFile/N2END[1] Tile_X4Y5_RegFile/N2END[2]
+ Tile_X4Y5_RegFile/N2END[3] Tile_X4Y5_RegFile/N2END[4] Tile_X4Y5_RegFile/N2END[5]
+ Tile_X4Y5_RegFile/N2END[6] Tile_X4Y5_RegFile/N2END[7] Tile_X4Y6_RegFile/N2END[0]
+ Tile_X4Y6_RegFile/N2END[1] Tile_X4Y6_RegFile/N2END[2] Tile_X4Y6_RegFile/N2END[3]
+ Tile_X4Y6_RegFile/N2END[4] Tile_X4Y6_RegFile/N2END[5] Tile_X4Y6_RegFile/N2END[6]
+ Tile_X4Y6_RegFile/N2END[7] Tile_X4Y7_RegFile/N2BEG[0] Tile_X4Y7_RegFile/N2BEG[1]
+ Tile_X4Y7_RegFile/N2BEG[2] Tile_X4Y7_RegFile/N2BEG[3] Tile_X4Y7_RegFile/N2BEG[4]
+ Tile_X4Y7_RegFile/N2BEG[5] Tile_X4Y7_RegFile/N2BEG[6] Tile_X4Y7_RegFile/N2BEG[7]
+ Tile_X4Y6_RegFile/N4BEG[0] Tile_X4Y6_RegFile/N4BEG[10] Tile_X4Y6_RegFile/N4BEG[11]
+ Tile_X4Y6_RegFile/N4BEG[12] Tile_X4Y6_RegFile/N4BEG[13] Tile_X4Y6_RegFile/N4BEG[14]
+ Tile_X4Y6_RegFile/N4BEG[15] Tile_X4Y6_RegFile/N4BEG[1] Tile_X4Y6_RegFile/N4BEG[2]
+ Tile_X4Y6_RegFile/N4BEG[3] Tile_X4Y6_RegFile/N4BEG[4] Tile_X4Y6_RegFile/N4BEG[5]
+ Tile_X4Y6_RegFile/N4BEG[6] Tile_X4Y6_RegFile/N4BEG[7] Tile_X4Y6_RegFile/N4BEG[8]
+ Tile_X4Y6_RegFile/N4BEG[9] Tile_X4Y7_RegFile/N4BEG[0] Tile_X4Y7_RegFile/N4BEG[10]
+ Tile_X4Y7_RegFile/N4BEG[11] Tile_X4Y7_RegFile/N4BEG[12] Tile_X4Y7_RegFile/N4BEG[13]
+ Tile_X4Y7_RegFile/N4BEG[14] Tile_X4Y7_RegFile/N4BEG[15] Tile_X4Y7_RegFile/N4BEG[1]
+ Tile_X4Y7_RegFile/N4BEG[2] Tile_X4Y7_RegFile/N4BEG[3] Tile_X4Y7_RegFile/N4BEG[4]
+ Tile_X4Y7_RegFile/N4BEG[5] Tile_X4Y7_RegFile/N4BEG[6] Tile_X4Y7_RegFile/N4BEG[7]
+ Tile_X4Y7_RegFile/N4BEG[8] Tile_X4Y7_RegFile/N4BEG[9] Tile_X4Y6_RegFile/NN4BEG[0]
+ Tile_X4Y6_RegFile/NN4BEG[10] Tile_X4Y6_RegFile/NN4BEG[11] Tile_X4Y6_RegFile/NN4BEG[12]
+ Tile_X4Y6_RegFile/NN4BEG[13] Tile_X4Y6_RegFile/NN4BEG[14] Tile_X4Y6_RegFile/NN4BEG[15]
+ Tile_X4Y6_RegFile/NN4BEG[1] Tile_X4Y6_RegFile/NN4BEG[2] Tile_X4Y6_RegFile/NN4BEG[3]
+ Tile_X4Y6_RegFile/NN4BEG[4] Tile_X4Y6_RegFile/NN4BEG[5] Tile_X4Y6_RegFile/NN4BEG[6]
+ Tile_X4Y6_RegFile/NN4BEG[7] Tile_X4Y6_RegFile/NN4BEG[8] Tile_X4Y6_RegFile/NN4BEG[9]
+ Tile_X4Y7_RegFile/NN4BEG[0] Tile_X4Y7_RegFile/NN4BEG[10] Tile_X4Y7_RegFile/NN4BEG[11]
+ Tile_X4Y7_RegFile/NN4BEG[12] Tile_X4Y7_RegFile/NN4BEG[13] Tile_X4Y7_RegFile/NN4BEG[14]
+ Tile_X4Y7_RegFile/NN4BEG[15] Tile_X4Y7_RegFile/NN4BEG[1] Tile_X4Y7_RegFile/NN4BEG[2]
+ Tile_X4Y7_RegFile/NN4BEG[3] Tile_X4Y7_RegFile/NN4BEG[4] Tile_X4Y7_RegFile/NN4BEG[5]
+ Tile_X4Y7_RegFile/NN4BEG[6] Tile_X4Y7_RegFile/NN4BEG[7] Tile_X4Y7_RegFile/NN4BEG[8]
+ Tile_X4Y7_RegFile/NN4BEG[9] Tile_X4Y7_RegFile/S1END[0] Tile_X4Y7_RegFile/S1END[1]
+ Tile_X4Y7_RegFile/S1END[2] Tile_X4Y7_RegFile/S1END[3] Tile_X4Y6_RegFile/S1END[0]
+ Tile_X4Y6_RegFile/S1END[1] Tile_X4Y6_RegFile/S1END[2] Tile_X4Y6_RegFile/S1END[3]
+ Tile_X4Y7_RegFile/S2MID[0] Tile_X4Y7_RegFile/S2MID[1] Tile_X4Y7_RegFile/S2MID[2]
+ Tile_X4Y7_RegFile/S2MID[3] Tile_X4Y7_RegFile/S2MID[4] Tile_X4Y7_RegFile/S2MID[5]
+ Tile_X4Y7_RegFile/S2MID[6] Tile_X4Y7_RegFile/S2MID[7] Tile_X4Y7_RegFile/S2END[0]
+ Tile_X4Y7_RegFile/S2END[1] Tile_X4Y7_RegFile/S2END[2] Tile_X4Y7_RegFile/S2END[3]
+ Tile_X4Y7_RegFile/S2END[4] Tile_X4Y7_RegFile/S2END[5] Tile_X4Y7_RegFile/S2END[6]
+ Tile_X4Y7_RegFile/S2END[7] Tile_X4Y6_RegFile/S2END[0] Tile_X4Y6_RegFile/S2END[1]
+ Tile_X4Y6_RegFile/S2END[2] Tile_X4Y6_RegFile/S2END[3] Tile_X4Y6_RegFile/S2END[4]
+ Tile_X4Y6_RegFile/S2END[5] Tile_X4Y6_RegFile/S2END[6] Tile_X4Y6_RegFile/S2END[7]
+ Tile_X4Y6_RegFile/S2MID[0] Tile_X4Y6_RegFile/S2MID[1] Tile_X4Y6_RegFile/S2MID[2]
+ Tile_X4Y6_RegFile/S2MID[3] Tile_X4Y6_RegFile/S2MID[4] Tile_X4Y6_RegFile/S2MID[5]
+ Tile_X4Y6_RegFile/S2MID[6] Tile_X4Y6_RegFile/S2MID[7] Tile_X4Y7_RegFile/S4END[0]
+ Tile_X4Y7_RegFile/S4END[10] Tile_X4Y7_RegFile/S4END[11] Tile_X4Y7_RegFile/S4END[12]
+ Tile_X4Y7_RegFile/S4END[13] Tile_X4Y7_RegFile/S4END[14] Tile_X4Y7_RegFile/S4END[15]
+ Tile_X4Y7_RegFile/S4END[1] Tile_X4Y7_RegFile/S4END[2] Tile_X4Y7_RegFile/S4END[3]
+ Tile_X4Y7_RegFile/S4END[4] Tile_X4Y7_RegFile/S4END[5] Tile_X4Y7_RegFile/S4END[6]
+ Tile_X4Y7_RegFile/S4END[7] Tile_X4Y7_RegFile/S4END[8] Tile_X4Y7_RegFile/S4END[9]
+ Tile_X4Y6_RegFile/S4END[0] Tile_X4Y6_RegFile/S4END[10] Tile_X4Y6_RegFile/S4END[11]
+ Tile_X4Y6_RegFile/S4END[12] Tile_X4Y6_RegFile/S4END[13] Tile_X4Y6_RegFile/S4END[14]
+ Tile_X4Y6_RegFile/S4END[15] Tile_X4Y6_RegFile/S4END[1] Tile_X4Y6_RegFile/S4END[2]
+ Tile_X4Y6_RegFile/S4END[3] Tile_X4Y6_RegFile/S4END[4] Tile_X4Y6_RegFile/S4END[5]
+ Tile_X4Y6_RegFile/S4END[6] Tile_X4Y6_RegFile/S4END[7] Tile_X4Y6_RegFile/S4END[8]
+ Tile_X4Y6_RegFile/S4END[9] Tile_X4Y7_RegFile/SS4END[0] Tile_X4Y7_RegFile/SS4END[10]
+ Tile_X4Y7_RegFile/SS4END[11] Tile_X4Y7_RegFile/SS4END[12] Tile_X4Y7_RegFile/SS4END[13]
+ Tile_X4Y7_RegFile/SS4END[14] Tile_X4Y7_RegFile/SS4END[15] Tile_X4Y7_RegFile/SS4END[1]
+ Tile_X4Y7_RegFile/SS4END[2] Tile_X4Y7_RegFile/SS4END[3] Tile_X4Y7_RegFile/SS4END[4]
+ Tile_X4Y7_RegFile/SS4END[5] Tile_X4Y7_RegFile/SS4END[6] Tile_X4Y7_RegFile/SS4END[7]
+ Tile_X4Y7_RegFile/SS4END[8] Tile_X4Y7_RegFile/SS4END[9] Tile_X4Y6_RegFile/SS4END[0]
+ Tile_X4Y6_RegFile/SS4END[10] Tile_X4Y6_RegFile/SS4END[11] Tile_X4Y6_RegFile/SS4END[12]
+ Tile_X4Y6_RegFile/SS4END[13] Tile_X4Y6_RegFile/SS4END[14] Tile_X4Y6_RegFile/SS4END[15]
+ Tile_X4Y6_RegFile/SS4END[1] Tile_X4Y6_RegFile/SS4END[2] Tile_X4Y6_RegFile/SS4END[3]
+ Tile_X4Y6_RegFile/SS4END[4] Tile_X4Y6_RegFile/SS4END[5] Tile_X4Y6_RegFile/SS4END[6]
+ Tile_X4Y6_RegFile/SS4END[7] Tile_X4Y6_RegFile/SS4END[8] Tile_X4Y6_RegFile/SS4END[9]
+ Tile_X4Y6_RegFile/UserCLK Tile_X4Y5_RegFile/UserCLK VGND VPWR Tile_X3Y6_LUT4AB/W1END[0]
+ Tile_X3Y6_LUT4AB/W1END[1] Tile_X3Y6_LUT4AB/W1END[2] Tile_X3Y6_LUT4AB/W1END[3] Tile_X5Y6_LUT4AB/W1BEG[0]
+ Tile_X5Y6_LUT4AB/W1BEG[1] Tile_X5Y6_LUT4AB/W1BEG[2] Tile_X5Y6_LUT4AB/W1BEG[3] Tile_X3Y6_LUT4AB/W2MID[0]
+ Tile_X3Y6_LUT4AB/W2MID[1] Tile_X3Y6_LUT4AB/W2MID[2] Tile_X3Y6_LUT4AB/W2MID[3] Tile_X3Y6_LUT4AB/W2MID[4]
+ Tile_X3Y6_LUT4AB/W2MID[5] Tile_X3Y6_LUT4AB/W2MID[6] Tile_X3Y6_LUT4AB/W2MID[7] Tile_X3Y6_LUT4AB/W2END[0]
+ Tile_X3Y6_LUT4AB/W2END[1] Tile_X3Y6_LUT4AB/W2END[2] Tile_X3Y6_LUT4AB/W2END[3] Tile_X3Y6_LUT4AB/W2END[4]
+ Tile_X3Y6_LUT4AB/W2END[5] Tile_X3Y6_LUT4AB/W2END[6] Tile_X3Y6_LUT4AB/W2END[7] Tile_X5Y6_LUT4AB/W2BEGb[0]
+ Tile_X5Y6_LUT4AB/W2BEGb[1] Tile_X5Y6_LUT4AB/W2BEGb[2] Tile_X5Y6_LUT4AB/W2BEGb[3]
+ Tile_X5Y6_LUT4AB/W2BEGb[4] Tile_X5Y6_LUT4AB/W2BEGb[5] Tile_X5Y6_LUT4AB/W2BEGb[6]
+ Tile_X5Y6_LUT4AB/W2BEGb[7] Tile_X5Y6_LUT4AB/W2BEG[0] Tile_X5Y6_LUT4AB/W2BEG[1] Tile_X5Y6_LUT4AB/W2BEG[2]
+ Tile_X5Y6_LUT4AB/W2BEG[3] Tile_X5Y6_LUT4AB/W2BEG[4] Tile_X5Y6_LUT4AB/W2BEG[5] Tile_X5Y6_LUT4AB/W2BEG[6]
+ Tile_X5Y6_LUT4AB/W2BEG[7] Tile_X3Y6_LUT4AB/W6END[0] Tile_X3Y6_LUT4AB/W6END[10] Tile_X3Y6_LUT4AB/W6END[11]
+ Tile_X3Y6_LUT4AB/W6END[1] Tile_X3Y6_LUT4AB/W6END[2] Tile_X3Y6_LUT4AB/W6END[3] Tile_X3Y6_LUT4AB/W6END[4]
+ Tile_X3Y6_LUT4AB/W6END[5] Tile_X3Y6_LUT4AB/W6END[6] Tile_X3Y6_LUT4AB/W6END[7] Tile_X3Y6_LUT4AB/W6END[8]
+ Tile_X3Y6_LUT4AB/W6END[9] Tile_X5Y6_LUT4AB/W6BEG[0] Tile_X5Y6_LUT4AB/W6BEG[10] Tile_X5Y6_LUT4AB/W6BEG[11]
+ Tile_X5Y6_LUT4AB/W6BEG[1] Tile_X5Y6_LUT4AB/W6BEG[2] Tile_X5Y6_LUT4AB/W6BEG[3] Tile_X5Y6_LUT4AB/W6BEG[4]
+ Tile_X5Y6_LUT4AB/W6BEG[5] Tile_X5Y6_LUT4AB/W6BEG[6] Tile_X5Y6_LUT4AB/W6BEG[7] Tile_X5Y6_LUT4AB/W6BEG[8]
+ Tile_X5Y6_LUT4AB/W6BEG[9] Tile_X3Y6_LUT4AB/WW4END[0] Tile_X3Y6_LUT4AB/WW4END[10]
+ Tile_X3Y6_LUT4AB/WW4END[11] Tile_X3Y6_LUT4AB/WW4END[12] Tile_X3Y6_LUT4AB/WW4END[13]
+ Tile_X3Y6_LUT4AB/WW4END[14] Tile_X3Y6_LUT4AB/WW4END[15] Tile_X3Y6_LUT4AB/WW4END[1]
+ Tile_X3Y6_LUT4AB/WW4END[2] Tile_X3Y6_LUT4AB/WW4END[3] Tile_X3Y6_LUT4AB/WW4END[4]
+ Tile_X3Y6_LUT4AB/WW4END[5] Tile_X3Y6_LUT4AB/WW4END[6] Tile_X3Y6_LUT4AB/WW4END[7]
+ Tile_X3Y6_LUT4AB/WW4END[8] Tile_X3Y6_LUT4AB/WW4END[9] Tile_X5Y6_LUT4AB/WW4BEG[0]
+ Tile_X5Y6_LUT4AB/WW4BEG[10] Tile_X5Y6_LUT4AB/WW4BEG[11] Tile_X5Y6_LUT4AB/WW4BEG[12]
+ Tile_X5Y6_LUT4AB/WW4BEG[13] Tile_X5Y6_LUT4AB/WW4BEG[14] Tile_X5Y6_LUT4AB/WW4BEG[15]
+ Tile_X5Y6_LUT4AB/WW4BEG[1] Tile_X5Y6_LUT4AB/WW4BEG[2] Tile_X5Y6_LUT4AB/WW4BEG[3]
+ Tile_X5Y6_LUT4AB/WW4BEG[4] Tile_X5Y6_LUT4AB/WW4BEG[5] Tile_X5Y6_LUT4AB/WW4BEG[6]
+ Tile_X5Y6_LUT4AB/WW4BEG[7] Tile_X5Y6_LUT4AB/WW4BEG[8] Tile_X5Y6_LUT4AB/WW4BEG[9]
+ RegFile
XTile_X6Y10_LUT4AB Tile_X6Y11_LUT4AB/Co Tile_X6Y9_LUT4AB/Ci Tile_X6Y10_LUT4AB/E1BEG[0]
+ Tile_X6Y10_LUT4AB/E1BEG[1] Tile_X6Y10_LUT4AB/E1BEG[2] Tile_X6Y10_LUT4AB/E1BEG[3]
+ Tile_X6Y10_LUT4AB/E1END[0] Tile_X6Y10_LUT4AB/E1END[1] Tile_X6Y10_LUT4AB/E1END[2]
+ Tile_X6Y10_LUT4AB/E1END[3] Tile_X6Y10_LUT4AB/E2BEG[0] Tile_X6Y10_LUT4AB/E2BEG[1]
+ Tile_X6Y10_LUT4AB/E2BEG[2] Tile_X6Y10_LUT4AB/E2BEG[3] Tile_X6Y10_LUT4AB/E2BEG[4]
+ Tile_X6Y10_LUT4AB/E2BEG[5] Tile_X6Y10_LUT4AB/E2BEG[6] Tile_X6Y10_LUT4AB/E2BEG[7]
+ Tile_X6Y10_LUT4AB/E2BEGb[0] Tile_X6Y10_LUT4AB/E2BEGb[1] Tile_X6Y10_LUT4AB/E2BEGb[2]
+ Tile_X6Y10_LUT4AB/E2BEGb[3] Tile_X6Y10_LUT4AB/E2BEGb[4] Tile_X6Y10_LUT4AB/E2BEGb[5]
+ Tile_X6Y10_LUT4AB/E2BEGb[6] Tile_X6Y10_LUT4AB/E2BEGb[7] Tile_X6Y10_LUT4AB/E2END[0]
+ Tile_X6Y10_LUT4AB/E2END[1] Tile_X6Y10_LUT4AB/E2END[2] Tile_X6Y10_LUT4AB/E2END[3]
+ Tile_X6Y10_LUT4AB/E2END[4] Tile_X6Y10_LUT4AB/E2END[5] Tile_X6Y10_LUT4AB/E2END[6]
+ Tile_X6Y10_LUT4AB/E2END[7] Tile_X6Y10_LUT4AB/E2MID[0] Tile_X6Y10_LUT4AB/E2MID[1]
+ Tile_X6Y10_LUT4AB/E2MID[2] Tile_X6Y10_LUT4AB/E2MID[3] Tile_X6Y10_LUT4AB/E2MID[4]
+ Tile_X6Y10_LUT4AB/E2MID[5] Tile_X6Y10_LUT4AB/E2MID[6] Tile_X6Y10_LUT4AB/E2MID[7]
+ Tile_X6Y10_LUT4AB/E6BEG[0] Tile_X6Y10_LUT4AB/E6BEG[10] Tile_X6Y10_LUT4AB/E6BEG[11]
+ Tile_X6Y10_LUT4AB/E6BEG[1] Tile_X6Y10_LUT4AB/E6BEG[2] Tile_X6Y10_LUT4AB/E6BEG[3]
+ Tile_X6Y10_LUT4AB/E6BEG[4] Tile_X6Y10_LUT4AB/E6BEG[5] Tile_X6Y10_LUT4AB/E6BEG[6]
+ Tile_X6Y10_LUT4AB/E6BEG[7] Tile_X6Y10_LUT4AB/E6BEG[8] Tile_X6Y10_LUT4AB/E6BEG[9]
+ Tile_X6Y10_LUT4AB/E6END[0] Tile_X6Y10_LUT4AB/E6END[10] Tile_X6Y10_LUT4AB/E6END[11]
+ Tile_X6Y10_LUT4AB/E6END[1] Tile_X6Y10_LUT4AB/E6END[2] Tile_X6Y10_LUT4AB/E6END[3]
+ Tile_X6Y10_LUT4AB/E6END[4] Tile_X6Y10_LUT4AB/E6END[5] Tile_X6Y10_LUT4AB/E6END[6]
+ Tile_X6Y10_LUT4AB/E6END[7] Tile_X6Y10_LUT4AB/E6END[8] Tile_X6Y10_LUT4AB/E6END[9]
+ Tile_X6Y10_LUT4AB/EE4BEG[0] Tile_X6Y10_LUT4AB/EE4BEG[10] Tile_X6Y10_LUT4AB/EE4BEG[11]
+ Tile_X6Y10_LUT4AB/EE4BEG[12] Tile_X6Y10_LUT4AB/EE4BEG[13] Tile_X6Y10_LUT4AB/EE4BEG[14]
+ Tile_X6Y10_LUT4AB/EE4BEG[15] Tile_X6Y10_LUT4AB/EE4BEG[1] Tile_X6Y10_LUT4AB/EE4BEG[2]
+ Tile_X6Y10_LUT4AB/EE4BEG[3] Tile_X6Y10_LUT4AB/EE4BEG[4] Tile_X6Y10_LUT4AB/EE4BEG[5]
+ Tile_X6Y10_LUT4AB/EE4BEG[6] Tile_X6Y10_LUT4AB/EE4BEG[7] Tile_X6Y10_LUT4AB/EE4BEG[8]
+ Tile_X6Y10_LUT4AB/EE4BEG[9] Tile_X6Y10_LUT4AB/EE4END[0] Tile_X6Y10_LUT4AB/EE4END[10]
+ Tile_X6Y10_LUT4AB/EE4END[11] Tile_X6Y10_LUT4AB/EE4END[12] Tile_X6Y10_LUT4AB/EE4END[13]
+ Tile_X6Y10_LUT4AB/EE4END[14] Tile_X6Y10_LUT4AB/EE4END[15] Tile_X6Y10_LUT4AB/EE4END[1]
+ Tile_X6Y10_LUT4AB/EE4END[2] Tile_X6Y10_LUT4AB/EE4END[3] Tile_X6Y10_LUT4AB/EE4END[4]
+ Tile_X6Y10_LUT4AB/EE4END[5] Tile_X6Y10_LUT4AB/EE4END[6] Tile_X6Y10_LUT4AB/EE4END[7]
+ Tile_X6Y10_LUT4AB/EE4END[8] Tile_X6Y10_LUT4AB/EE4END[9] Tile_X6Y10_LUT4AB/FrameData[0]
+ Tile_X6Y10_LUT4AB/FrameData[10] Tile_X6Y10_LUT4AB/FrameData[11] Tile_X6Y10_LUT4AB/FrameData[12]
+ Tile_X6Y10_LUT4AB/FrameData[13] Tile_X6Y10_LUT4AB/FrameData[14] Tile_X6Y10_LUT4AB/FrameData[15]
+ Tile_X6Y10_LUT4AB/FrameData[16] Tile_X6Y10_LUT4AB/FrameData[17] Tile_X6Y10_LUT4AB/FrameData[18]
+ Tile_X6Y10_LUT4AB/FrameData[19] Tile_X6Y10_LUT4AB/FrameData[1] Tile_X6Y10_LUT4AB/FrameData[20]
+ Tile_X6Y10_LUT4AB/FrameData[21] Tile_X6Y10_LUT4AB/FrameData[22] Tile_X6Y10_LUT4AB/FrameData[23]
+ Tile_X6Y10_LUT4AB/FrameData[24] Tile_X6Y10_LUT4AB/FrameData[25] Tile_X6Y10_LUT4AB/FrameData[26]
+ Tile_X6Y10_LUT4AB/FrameData[27] Tile_X6Y10_LUT4AB/FrameData[28] Tile_X6Y10_LUT4AB/FrameData[29]
+ Tile_X6Y10_LUT4AB/FrameData[2] Tile_X6Y10_LUT4AB/FrameData[30] Tile_X6Y10_LUT4AB/FrameData[31]
+ Tile_X6Y10_LUT4AB/FrameData[3] Tile_X6Y10_LUT4AB/FrameData[4] Tile_X6Y10_LUT4AB/FrameData[5]
+ Tile_X6Y10_LUT4AB/FrameData[6] Tile_X6Y10_LUT4AB/FrameData[7] Tile_X6Y10_LUT4AB/FrameData[8]
+ Tile_X6Y10_LUT4AB/FrameData[9] Tile_X6Y10_LUT4AB/FrameData_O[0] Tile_X6Y10_LUT4AB/FrameData_O[10]
+ Tile_X6Y10_LUT4AB/FrameData_O[11] Tile_X6Y10_LUT4AB/FrameData_O[12] Tile_X6Y10_LUT4AB/FrameData_O[13]
+ Tile_X6Y10_LUT4AB/FrameData_O[14] Tile_X6Y10_LUT4AB/FrameData_O[15] Tile_X6Y10_LUT4AB/FrameData_O[16]
+ Tile_X6Y10_LUT4AB/FrameData_O[17] Tile_X6Y10_LUT4AB/FrameData_O[18] Tile_X6Y10_LUT4AB/FrameData_O[19]
+ Tile_X6Y10_LUT4AB/FrameData_O[1] Tile_X6Y10_LUT4AB/FrameData_O[20] Tile_X6Y10_LUT4AB/FrameData_O[21]
+ Tile_X6Y10_LUT4AB/FrameData_O[22] Tile_X6Y10_LUT4AB/FrameData_O[23] Tile_X6Y10_LUT4AB/FrameData_O[24]
+ Tile_X6Y10_LUT4AB/FrameData_O[25] Tile_X6Y10_LUT4AB/FrameData_O[26] Tile_X6Y10_LUT4AB/FrameData_O[27]
+ Tile_X6Y10_LUT4AB/FrameData_O[28] Tile_X6Y10_LUT4AB/FrameData_O[29] Tile_X6Y10_LUT4AB/FrameData_O[2]
+ Tile_X6Y10_LUT4AB/FrameData_O[30] Tile_X6Y10_LUT4AB/FrameData_O[31] Tile_X6Y10_LUT4AB/FrameData_O[3]
+ Tile_X6Y10_LUT4AB/FrameData_O[4] Tile_X6Y10_LUT4AB/FrameData_O[5] Tile_X6Y10_LUT4AB/FrameData_O[6]
+ Tile_X6Y10_LUT4AB/FrameData_O[7] Tile_X6Y10_LUT4AB/FrameData_O[8] Tile_X6Y10_LUT4AB/FrameData_O[9]
+ Tile_X6Y10_LUT4AB/FrameStrobe[0] Tile_X6Y10_LUT4AB/FrameStrobe[10] Tile_X6Y10_LUT4AB/FrameStrobe[11]
+ Tile_X6Y10_LUT4AB/FrameStrobe[12] Tile_X6Y10_LUT4AB/FrameStrobe[13] Tile_X6Y10_LUT4AB/FrameStrobe[14]
+ Tile_X6Y10_LUT4AB/FrameStrobe[15] Tile_X6Y10_LUT4AB/FrameStrobe[16] Tile_X6Y10_LUT4AB/FrameStrobe[17]
+ Tile_X6Y10_LUT4AB/FrameStrobe[18] Tile_X6Y10_LUT4AB/FrameStrobe[19] Tile_X6Y10_LUT4AB/FrameStrobe[1]
+ Tile_X6Y10_LUT4AB/FrameStrobe[2] Tile_X6Y10_LUT4AB/FrameStrobe[3] Tile_X6Y10_LUT4AB/FrameStrobe[4]
+ Tile_X6Y10_LUT4AB/FrameStrobe[5] Tile_X6Y10_LUT4AB/FrameStrobe[6] Tile_X6Y10_LUT4AB/FrameStrobe[7]
+ Tile_X6Y10_LUT4AB/FrameStrobe[8] Tile_X6Y10_LUT4AB/FrameStrobe[9] Tile_X6Y9_LUT4AB/FrameStrobe[0]
+ Tile_X6Y9_LUT4AB/FrameStrobe[10] Tile_X6Y9_LUT4AB/FrameStrobe[11] Tile_X6Y9_LUT4AB/FrameStrobe[12]
+ Tile_X6Y9_LUT4AB/FrameStrobe[13] Tile_X6Y9_LUT4AB/FrameStrobe[14] Tile_X6Y9_LUT4AB/FrameStrobe[15]
+ Tile_X6Y9_LUT4AB/FrameStrobe[16] Tile_X6Y9_LUT4AB/FrameStrobe[17] Tile_X6Y9_LUT4AB/FrameStrobe[18]
+ Tile_X6Y9_LUT4AB/FrameStrobe[19] Tile_X6Y9_LUT4AB/FrameStrobe[1] Tile_X6Y9_LUT4AB/FrameStrobe[2]
+ Tile_X6Y9_LUT4AB/FrameStrobe[3] Tile_X6Y9_LUT4AB/FrameStrobe[4] Tile_X6Y9_LUT4AB/FrameStrobe[5]
+ Tile_X6Y9_LUT4AB/FrameStrobe[6] Tile_X6Y9_LUT4AB/FrameStrobe[7] Tile_X6Y9_LUT4AB/FrameStrobe[8]
+ Tile_X6Y9_LUT4AB/FrameStrobe[9] Tile_X6Y9_LUT4AB/N1END[0] Tile_X6Y9_LUT4AB/N1END[1]
+ Tile_X6Y9_LUT4AB/N1END[2] Tile_X6Y9_LUT4AB/N1END[3] Tile_X6Y11_LUT4AB/N1BEG[0] Tile_X6Y11_LUT4AB/N1BEG[1]
+ Tile_X6Y11_LUT4AB/N1BEG[2] Tile_X6Y11_LUT4AB/N1BEG[3] Tile_X6Y9_LUT4AB/N2MID[0]
+ Tile_X6Y9_LUT4AB/N2MID[1] Tile_X6Y9_LUT4AB/N2MID[2] Tile_X6Y9_LUT4AB/N2MID[3] Tile_X6Y9_LUT4AB/N2MID[4]
+ Tile_X6Y9_LUT4AB/N2MID[5] Tile_X6Y9_LUT4AB/N2MID[6] Tile_X6Y9_LUT4AB/N2MID[7] Tile_X6Y9_LUT4AB/N2END[0]
+ Tile_X6Y9_LUT4AB/N2END[1] Tile_X6Y9_LUT4AB/N2END[2] Tile_X6Y9_LUT4AB/N2END[3] Tile_X6Y9_LUT4AB/N2END[4]
+ Tile_X6Y9_LUT4AB/N2END[5] Tile_X6Y9_LUT4AB/N2END[6] Tile_X6Y9_LUT4AB/N2END[7] Tile_X6Y10_LUT4AB/N2END[0]
+ Tile_X6Y10_LUT4AB/N2END[1] Tile_X6Y10_LUT4AB/N2END[2] Tile_X6Y10_LUT4AB/N2END[3]
+ Tile_X6Y10_LUT4AB/N2END[4] Tile_X6Y10_LUT4AB/N2END[5] Tile_X6Y10_LUT4AB/N2END[6]
+ Tile_X6Y10_LUT4AB/N2END[7] Tile_X6Y11_LUT4AB/N2BEG[0] Tile_X6Y11_LUT4AB/N2BEG[1]
+ Tile_X6Y11_LUT4AB/N2BEG[2] Tile_X6Y11_LUT4AB/N2BEG[3] Tile_X6Y11_LUT4AB/N2BEG[4]
+ Tile_X6Y11_LUT4AB/N2BEG[5] Tile_X6Y11_LUT4AB/N2BEG[6] Tile_X6Y11_LUT4AB/N2BEG[7]
+ Tile_X6Y9_LUT4AB/N4END[0] Tile_X6Y9_LUT4AB/N4END[10] Tile_X6Y9_LUT4AB/N4END[11]
+ Tile_X6Y9_LUT4AB/N4END[12] Tile_X6Y9_LUT4AB/N4END[13] Tile_X6Y9_LUT4AB/N4END[14]
+ Tile_X6Y9_LUT4AB/N4END[15] Tile_X6Y9_LUT4AB/N4END[1] Tile_X6Y9_LUT4AB/N4END[2] Tile_X6Y9_LUT4AB/N4END[3]
+ Tile_X6Y9_LUT4AB/N4END[4] Tile_X6Y9_LUT4AB/N4END[5] Tile_X6Y9_LUT4AB/N4END[6] Tile_X6Y9_LUT4AB/N4END[7]
+ Tile_X6Y9_LUT4AB/N4END[8] Tile_X6Y9_LUT4AB/N4END[9] Tile_X6Y11_LUT4AB/N4BEG[0] Tile_X6Y11_LUT4AB/N4BEG[10]
+ Tile_X6Y11_LUT4AB/N4BEG[11] Tile_X6Y11_LUT4AB/N4BEG[12] Tile_X6Y11_LUT4AB/N4BEG[13]
+ Tile_X6Y11_LUT4AB/N4BEG[14] Tile_X6Y11_LUT4AB/N4BEG[15] Tile_X6Y11_LUT4AB/N4BEG[1]
+ Tile_X6Y11_LUT4AB/N4BEG[2] Tile_X6Y11_LUT4AB/N4BEG[3] Tile_X6Y11_LUT4AB/N4BEG[4]
+ Tile_X6Y11_LUT4AB/N4BEG[5] Tile_X6Y11_LUT4AB/N4BEG[6] Tile_X6Y11_LUT4AB/N4BEG[7]
+ Tile_X6Y11_LUT4AB/N4BEG[8] Tile_X6Y11_LUT4AB/N4BEG[9] Tile_X6Y9_LUT4AB/NN4END[0]
+ Tile_X6Y9_LUT4AB/NN4END[10] Tile_X6Y9_LUT4AB/NN4END[11] Tile_X6Y9_LUT4AB/NN4END[12]
+ Tile_X6Y9_LUT4AB/NN4END[13] Tile_X6Y9_LUT4AB/NN4END[14] Tile_X6Y9_LUT4AB/NN4END[15]
+ Tile_X6Y9_LUT4AB/NN4END[1] Tile_X6Y9_LUT4AB/NN4END[2] Tile_X6Y9_LUT4AB/NN4END[3]
+ Tile_X6Y9_LUT4AB/NN4END[4] Tile_X6Y9_LUT4AB/NN4END[5] Tile_X6Y9_LUT4AB/NN4END[6]
+ Tile_X6Y9_LUT4AB/NN4END[7] Tile_X6Y9_LUT4AB/NN4END[8] Tile_X6Y9_LUT4AB/NN4END[9]
+ Tile_X6Y11_LUT4AB/NN4BEG[0] Tile_X6Y11_LUT4AB/NN4BEG[10] Tile_X6Y11_LUT4AB/NN4BEG[11]
+ Tile_X6Y11_LUT4AB/NN4BEG[12] Tile_X6Y11_LUT4AB/NN4BEG[13] Tile_X6Y11_LUT4AB/NN4BEG[14]
+ Tile_X6Y11_LUT4AB/NN4BEG[15] Tile_X6Y11_LUT4AB/NN4BEG[1] Tile_X6Y11_LUT4AB/NN4BEG[2]
+ Tile_X6Y11_LUT4AB/NN4BEG[3] Tile_X6Y11_LUT4AB/NN4BEG[4] Tile_X6Y11_LUT4AB/NN4BEG[5]
+ Tile_X6Y11_LUT4AB/NN4BEG[6] Tile_X6Y11_LUT4AB/NN4BEG[7] Tile_X6Y11_LUT4AB/NN4BEG[8]
+ Tile_X6Y11_LUT4AB/NN4BEG[9] Tile_X6Y11_LUT4AB/S1END[0] Tile_X6Y11_LUT4AB/S1END[1]
+ Tile_X6Y11_LUT4AB/S1END[2] Tile_X6Y11_LUT4AB/S1END[3] Tile_X6Y9_LUT4AB/S1BEG[0]
+ Tile_X6Y9_LUT4AB/S1BEG[1] Tile_X6Y9_LUT4AB/S1BEG[2] Tile_X6Y9_LUT4AB/S1BEG[3] Tile_X6Y11_LUT4AB/S2MID[0]
+ Tile_X6Y11_LUT4AB/S2MID[1] Tile_X6Y11_LUT4AB/S2MID[2] Tile_X6Y11_LUT4AB/S2MID[3]
+ Tile_X6Y11_LUT4AB/S2MID[4] Tile_X6Y11_LUT4AB/S2MID[5] Tile_X6Y11_LUT4AB/S2MID[6]
+ Tile_X6Y11_LUT4AB/S2MID[7] Tile_X6Y11_LUT4AB/S2END[0] Tile_X6Y11_LUT4AB/S2END[1]
+ Tile_X6Y11_LUT4AB/S2END[2] Tile_X6Y11_LUT4AB/S2END[3] Tile_X6Y11_LUT4AB/S2END[4]
+ Tile_X6Y11_LUT4AB/S2END[5] Tile_X6Y11_LUT4AB/S2END[6] Tile_X6Y11_LUT4AB/S2END[7]
+ Tile_X6Y9_LUT4AB/S2BEGb[0] Tile_X6Y9_LUT4AB/S2BEGb[1] Tile_X6Y9_LUT4AB/S2BEGb[2]
+ Tile_X6Y9_LUT4AB/S2BEGb[3] Tile_X6Y9_LUT4AB/S2BEGb[4] Tile_X6Y9_LUT4AB/S2BEGb[5]
+ Tile_X6Y9_LUT4AB/S2BEGb[6] Tile_X6Y9_LUT4AB/S2BEGb[7] Tile_X6Y9_LUT4AB/S2BEG[0]
+ Tile_X6Y9_LUT4AB/S2BEG[1] Tile_X6Y9_LUT4AB/S2BEG[2] Tile_X6Y9_LUT4AB/S2BEG[3] Tile_X6Y9_LUT4AB/S2BEG[4]
+ Tile_X6Y9_LUT4AB/S2BEG[5] Tile_X6Y9_LUT4AB/S2BEG[6] Tile_X6Y9_LUT4AB/S2BEG[7] Tile_X6Y11_LUT4AB/S4END[0]
+ Tile_X6Y11_LUT4AB/S4END[10] Tile_X6Y11_LUT4AB/S4END[11] Tile_X6Y11_LUT4AB/S4END[12]
+ Tile_X6Y11_LUT4AB/S4END[13] Tile_X6Y11_LUT4AB/S4END[14] Tile_X6Y11_LUT4AB/S4END[15]
+ Tile_X6Y11_LUT4AB/S4END[1] Tile_X6Y11_LUT4AB/S4END[2] Tile_X6Y11_LUT4AB/S4END[3]
+ Tile_X6Y11_LUT4AB/S4END[4] Tile_X6Y11_LUT4AB/S4END[5] Tile_X6Y11_LUT4AB/S4END[6]
+ Tile_X6Y11_LUT4AB/S4END[7] Tile_X6Y11_LUT4AB/S4END[8] Tile_X6Y11_LUT4AB/S4END[9]
+ Tile_X6Y9_LUT4AB/S4BEG[0] Tile_X6Y9_LUT4AB/S4BEG[10] Tile_X6Y9_LUT4AB/S4BEG[11]
+ Tile_X6Y9_LUT4AB/S4BEG[12] Tile_X6Y9_LUT4AB/S4BEG[13] Tile_X6Y9_LUT4AB/S4BEG[14]
+ Tile_X6Y9_LUT4AB/S4BEG[15] Tile_X6Y9_LUT4AB/S4BEG[1] Tile_X6Y9_LUT4AB/S4BEG[2] Tile_X6Y9_LUT4AB/S4BEG[3]
+ Tile_X6Y9_LUT4AB/S4BEG[4] Tile_X6Y9_LUT4AB/S4BEG[5] Tile_X6Y9_LUT4AB/S4BEG[6] Tile_X6Y9_LUT4AB/S4BEG[7]
+ Tile_X6Y9_LUT4AB/S4BEG[8] Tile_X6Y9_LUT4AB/S4BEG[9] Tile_X6Y11_LUT4AB/SS4END[0]
+ Tile_X6Y11_LUT4AB/SS4END[10] Tile_X6Y11_LUT4AB/SS4END[11] Tile_X6Y11_LUT4AB/SS4END[12]
+ Tile_X6Y11_LUT4AB/SS4END[13] Tile_X6Y11_LUT4AB/SS4END[14] Tile_X6Y11_LUT4AB/SS4END[15]
+ Tile_X6Y11_LUT4AB/SS4END[1] Tile_X6Y11_LUT4AB/SS4END[2] Tile_X6Y11_LUT4AB/SS4END[3]
+ Tile_X6Y11_LUT4AB/SS4END[4] Tile_X6Y11_LUT4AB/SS4END[5] Tile_X6Y11_LUT4AB/SS4END[6]
+ Tile_X6Y11_LUT4AB/SS4END[7] Tile_X6Y11_LUT4AB/SS4END[8] Tile_X6Y11_LUT4AB/SS4END[9]
+ Tile_X6Y9_LUT4AB/SS4BEG[0] Tile_X6Y9_LUT4AB/SS4BEG[10] Tile_X6Y9_LUT4AB/SS4BEG[11]
+ Tile_X6Y9_LUT4AB/SS4BEG[12] Tile_X6Y9_LUT4AB/SS4BEG[13] Tile_X6Y9_LUT4AB/SS4BEG[14]
+ Tile_X6Y9_LUT4AB/SS4BEG[15] Tile_X6Y9_LUT4AB/SS4BEG[1] Tile_X6Y9_LUT4AB/SS4BEG[2]
+ Tile_X6Y9_LUT4AB/SS4BEG[3] Tile_X6Y9_LUT4AB/SS4BEG[4] Tile_X6Y9_LUT4AB/SS4BEG[5]
+ Tile_X6Y9_LUT4AB/SS4BEG[6] Tile_X6Y9_LUT4AB/SS4BEG[7] Tile_X6Y9_LUT4AB/SS4BEG[8]
+ Tile_X6Y9_LUT4AB/SS4BEG[9] Tile_X6Y10_LUT4AB/UserCLK Tile_X6Y9_LUT4AB/UserCLK VGND
+ VPWR Tile_X6Y10_LUT4AB/W1BEG[0] Tile_X6Y10_LUT4AB/W1BEG[1] Tile_X6Y10_LUT4AB/W1BEG[2]
+ Tile_X6Y10_LUT4AB/W1BEG[3] Tile_X6Y10_LUT4AB/W1END[0] Tile_X6Y10_LUT4AB/W1END[1]
+ Tile_X6Y10_LUT4AB/W1END[2] Tile_X6Y10_LUT4AB/W1END[3] Tile_X6Y10_LUT4AB/W2BEG[0]
+ Tile_X6Y10_LUT4AB/W2BEG[1] Tile_X6Y10_LUT4AB/W2BEG[2] Tile_X6Y10_LUT4AB/W2BEG[3]
+ Tile_X6Y10_LUT4AB/W2BEG[4] Tile_X6Y10_LUT4AB/W2BEG[5] Tile_X6Y10_LUT4AB/W2BEG[6]
+ Tile_X6Y10_LUT4AB/W2BEG[7] Tile_X5Y10_LUT4AB/W2END[0] Tile_X5Y10_LUT4AB/W2END[1]
+ Tile_X5Y10_LUT4AB/W2END[2] Tile_X5Y10_LUT4AB/W2END[3] Tile_X5Y10_LUT4AB/W2END[4]
+ Tile_X5Y10_LUT4AB/W2END[5] Tile_X5Y10_LUT4AB/W2END[6] Tile_X5Y10_LUT4AB/W2END[7]
+ Tile_X6Y10_LUT4AB/W2END[0] Tile_X6Y10_LUT4AB/W2END[1] Tile_X6Y10_LUT4AB/W2END[2]
+ Tile_X6Y10_LUT4AB/W2END[3] Tile_X6Y10_LUT4AB/W2END[4] Tile_X6Y10_LUT4AB/W2END[5]
+ Tile_X6Y10_LUT4AB/W2END[6] Tile_X6Y10_LUT4AB/W2END[7] Tile_X6Y10_LUT4AB/W2MID[0]
+ Tile_X6Y10_LUT4AB/W2MID[1] Tile_X6Y10_LUT4AB/W2MID[2] Tile_X6Y10_LUT4AB/W2MID[3]
+ Tile_X6Y10_LUT4AB/W2MID[4] Tile_X6Y10_LUT4AB/W2MID[5] Tile_X6Y10_LUT4AB/W2MID[6]
+ Tile_X6Y10_LUT4AB/W2MID[7] Tile_X6Y10_LUT4AB/W6BEG[0] Tile_X6Y10_LUT4AB/W6BEG[10]
+ Tile_X6Y10_LUT4AB/W6BEG[11] Tile_X6Y10_LUT4AB/W6BEG[1] Tile_X6Y10_LUT4AB/W6BEG[2]
+ Tile_X6Y10_LUT4AB/W6BEG[3] Tile_X6Y10_LUT4AB/W6BEG[4] Tile_X6Y10_LUT4AB/W6BEG[5]
+ Tile_X6Y10_LUT4AB/W6BEG[6] Tile_X6Y10_LUT4AB/W6BEG[7] Tile_X6Y10_LUT4AB/W6BEG[8]
+ Tile_X6Y10_LUT4AB/W6BEG[9] Tile_X6Y10_LUT4AB/W6END[0] Tile_X6Y10_LUT4AB/W6END[10]
+ Tile_X6Y10_LUT4AB/W6END[11] Tile_X6Y10_LUT4AB/W6END[1] Tile_X6Y10_LUT4AB/W6END[2]
+ Tile_X6Y10_LUT4AB/W6END[3] Tile_X6Y10_LUT4AB/W6END[4] Tile_X6Y10_LUT4AB/W6END[5]
+ Tile_X6Y10_LUT4AB/W6END[6] Tile_X6Y10_LUT4AB/W6END[7] Tile_X6Y10_LUT4AB/W6END[8]
+ Tile_X6Y10_LUT4AB/W6END[9] Tile_X6Y10_LUT4AB/WW4BEG[0] Tile_X6Y10_LUT4AB/WW4BEG[10]
+ Tile_X6Y10_LUT4AB/WW4BEG[11] Tile_X6Y10_LUT4AB/WW4BEG[12] Tile_X6Y10_LUT4AB/WW4BEG[13]
+ Tile_X6Y10_LUT4AB/WW4BEG[14] Tile_X6Y10_LUT4AB/WW4BEG[15] Tile_X6Y10_LUT4AB/WW4BEG[1]
+ Tile_X6Y10_LUT4AB/WW4BEG[2] Tile_X6Y10_LUT4AB/WW4BEG[3] Tile_X6Y10_LUT4AB/WW4BEG[4]
+ Tile_X6Y10_LUT4AB/WW4BEG[5] Tile_X6Y10_LUT4AB/WW4BEG[6] Tile_X6Y10_LUT4AB/WW4BEG[7]
+ Tile_X6Y10_LUT4AB/WW4BEG[8] Tile_X6Y10_LUT4AB/WW4BEG[9] Tile_X6Y10_LUT4AB/WW4END[0]
+ Tile_X6Y10_LUT4AB/WW4END[10] Tile_X6Y10_LUT4AB/WW4END[11] Tile_X6Y10_LUT4AB/WW4END[12]
+ Tile_X6Y10_LUT4AB/WW4END[13] Tile_X6Y10_LUT4AB/WW4END[14] Tile_X6Y10_LUT4AB/WW4END[15]
+ Tile_X6Y10_LUT4AB/WW4END[1] Tile_X6Y10_LUT4AB/WW4END[2] Tile_X6Y10_LUT4AB/WW4END[3]
+ Tile_X6Y10_LUT4AB/WW4END[4] Tile_X6Y10_LUT4AB/WW4END[5] Tile_X6Y10_LUT4AB/WW4END[6]
+ Tile_X6Y10_LUT4AB/WW4END[7] Tile_X6Y10_LUT4AB/WW4END[8] Tile_X6Y10_LUT4AB/WW4END[9]
+ LUT4AB
XTile_X0Y2_W_IO Tile_X0Y2_A_I_top Tile_X0Y2_A_O_top Tile_X0Y2_A_T_top Tile_X0Y2_A_config_C_bit0
+ Tile_X0Y2_A_config_C_bit1 Tile_X0Y2_A_config_C_bit2 Tile_X0Y2_A_config_C_bit3 Tile_X0Y2_B_I_top
+ Tile_X0Y2_B_O_top Tile_X0Y2_B_T_top Tile_X0Y2_B_config_C_bit0 Tile_X0Y2_B_config_C_bit1
+ Tile_X0Y2_B_config_C_bit2 Tile_X0Y2_B_config_C_bit3 Tile_X0Y2_W_IO/E1BEG[0] Tile_X0Y2_W_IO/E1BEG[1]
+ Tile_X0Y2_W_IO/E1BEG[2] Tile_X0Y2_W_IO/E1BEG[3] Tile_X0Y2_W_IO/E2BEG[0] Tile_X0Y2_W_IO/E2BEG[1]
+ Tile_X0Y2_W_IO/E2BEG[2] Tile_X0Y2_W_IO/E2BEG[3] Tile_X0Y2_W_IO/E2BEG[4] Tile_X0Y2_W_IO/E2BEG[5]
+ Tile_X0Y2_W_IO/E2BEG[6] Tile_X0Y2_W_IO/E2BEG[7] Tile_X0Y2_W_IO/E2BEGb[0] Tile_X0Y2_W_IO/E2BEGb[1]
+ Tile_X0Y2_W_IO/E2BEGb[2] Tile_X0Y2_W_IO/E2BEGb[3] Tile_X0Y2_W_IO/E2BEGb[4] Tile_X0Y2_W_IO/E2BEGb[5]
+ Tile_X0Y2_W_IO/E2BEGb[6] Tile_X0Y2_W_IO/E2BEGb[7] Tile_X0Y2_W_IO/E6BEG[0] Tile_X0Y2_W_IO/E6BEG[10]
+ Tile_X0Y2_W_IO/E6BEG[11] Tile_X0Y2_W_IO/E6BEG[1] Tile_X0Y2_W_IO/E6BEG[2] Tile_X0Y2_W_IO/E6BEG[3]
+ Tile_X0Y2_W_IO/E6BEG[4] Tile_X0Y2_W_IO/E6BEG[5] Tile_X0Y2_W_IO/E6BEG[6] Tile_X0Y2_W_IO/E6BEG[7]
+ Tile_X0Y2_W_IO/E6BEG[8] Tile_X0Y2_W_IO/E6BEG[9] Tile_X0Y2_W_IO/EE4BEG[0] Tile_X0Y2_W_IO/EE4BEG[10]
+ Tile_X0Y2_W_IO/EE4BEG[11] Tile_X0Y2_W_IO/EE4BEG[12] Tile_X0Y2_W_IO/EE4BEG[13] Tile_X0Y2_W_IO/EE4BEG[14]
+ Tile_X0Y2_W_IO/EE4BEG[15] Tile_X0Y2_W_IO/EE4BEG[1] Tile_X0Y2_W_IO/EE4BEG[2] Tile_X0Y2_W_IO/EE4BEG[3]
+ Tile_X0Y2_W_IO/EE4BEG[4] Tile_X0Y2_W_IO/EE4BEG[5] Tile_X0Y2_W_IO/EE4BEG[6] Tile_X0Y2_W_IO/EE4BEG[7]
+ Tile_X0Y2_W_IO/EE4BEG[8] Tile_X0Y2_W_IO/EE4BEG[9] FrameData[64] FrameData[74] FrameData[75]
+ FrameData[76] FrameData[77] FrameData[78] FrameData[79] FrameData[80] FrameData[81]
+ FrameData[82] FrameData[83] FrameData[65] FrameData[84] FrameData[85] FrameData[86]
+ FrameData[87] FrameData[88] FrameData[89] FrameData[90] FrameData[91] FrameData[92]
+ FrameData[93] FrameData[66] FrameData[94] FrameData[95] FrameData[67] FrameData[68]
+ FrameData[69] FrameData[70] FrameData[71] FrameData[72] FrameData[73] Tile_X1Y2_LUT4AB/FrameData[0]
+ Tile_X1Y2_LUT4AB/FrameData[10] Tile_X1Y2_LUT4AB/FrameData[11] Tile_X1Y2_LUT4AB/FrameData[12]
+ Tile_X1Y2_LUT4AB/FrameData[13] Tile_X1Y2_LUT4AB/FrameData[14] Tile_X1Y2_LUT4AB/FrameData[15]
+ Tile_X1Y2_LUT4AB/FrameData[16] Tile_X1Y2_LUT4AB/FrameData[17] Tile_X1Y2_LUT4AB/FrameData[18]
+ Tile_X1Y2_LUT4AB/FrameData[19] Tile_X1Y2_LUT4AB/FrameData[1] Tile_X1Y2_LUT4AB/FrameData[20]
+ Tile_X1Y2_LUT4AB/FrameData[21] Tile_X1Y2_LUT4AB/FrameData[22] Tile_X1Y2_LUT4AB/FrameData[23]
+ Tile_X1Y2_LUT4AB/FrameData[24] Tile_X1Y2_LUT4AB/FrameData[25] Tile_X1Y2_LUT4AB/FrameData[26]
+ Tile_X1Y2_LUT4AB/FrameData[27] Tile_X1Y2_LUT4AB/FrameData[28] Tile_X1Y2_LUT4AB/FrameData[29]
+ Tile_X1Y2_LUT4AB/FrameData[2] Tile_X1Y2_LUT4AB/FrameData[30] Tile_X1Y2_LUT4AB/FrameData[31]
+ Tile_X1Y2_LUT4AB/FrameData[3] Tile_X1Y2_LUT4AB/FrameData[4] Tile_X1Y2_LUT4AB/FrameData[5]
+ Tile_X1Y2_LUT4AB/FrameData[6] Tile_X1Y2_LUT4AB/FrameData[7] Tile_X1Y2_LUT4AB/FrameData[8]
+ Tile_X1Y2_LUT4AB/FrameData[9] Tile_X0Y2_W_IO/FrameStrobe[0] Tile_X0Y2_W_IO/FrameStrobe[10]
+ Tile_X0Y2_W_IO/FrameStrobe[11] Tile_X0Y2_W_IO/FrameStrobe[12] Tile_X0Y2_W_IO/FrameStrobe[13]
+ Tile_X0Y2_W_IO/FrameStrobe[14] Tile_X0Y2_W_IO/FrameStrobe[15] Tile_X0Y2_W_IO/FrameStrobe[16]
+ Tile_X0Y2_W_IO/FrameStrobe[17] Tile_X0Y2_W_IO/FrameStrobe[18] Tile_X0Y2_W_IO/FrameStrobe[19]
+ Tile_X0Y2_W_IO/FrameStrobe[1] Tile_X0Y2_W_IO/FrameStrobe[2] Tile_X0Y2_W_IO/FrameStrobe[3]
+ Tile_X0Y2_W_IO/FrameStrobe[4] Tile_X0Y2_W_IO/FrameStrobe[5] Tile_X0Y2_W_IO/FrameStrobe[6]
+ Tile_X0Y2_W_IO/FrameStrobe[7] Tile_X0Y2_W_IO/FrameStrobe[8] Tile_X0Y2_W_IO/FrameStrobe[9]
+ Tile_X0Y1_W_IO/FrameStrobe[0] Tile_X0Y1_W_IO/FrameStrobe[10] Tile_X0Y1_W_IO/FrameStrobe[11]
+ Tile_X0Y1_W_IO/FrameStrobe[12] Tile_X0Y1_W_IO/FrameStrobe[13] Tile_X0Y1_W_IO/FrameStrobe[14]
+ Tile_X0Y1_W_IO/FrameStrobe[15] Tile_X0Y1_W_IO/FrameStrobe[16] Tile_X0Y1_W_IO/FrameStrobe[17]
+ Tile_X0Y1_W_IO/FrameStrobe[18] Tile_X0Y1_W_IO/FrameStrobe[19] Tile_X0Y1_W_IO/FrameStrobe[1]
+ Tile_X0Y1_W_IO/FrameStrobe[2] Tile_X0Y1_W_IO/FrameStrobe[3] Tile_X0Y1_W_IO/FrameStrobe[4]
+ Tile_X0Y1_W_IO/FrameStrobe[5] Tile_X0Y1_W_IO/FrameStrobe[6] Tile_X0Y1_W_IO/FrameStrobe[7]
+ Tile_X0Y1_W_IO/FrameStrobe[8] Tile_X0Y1_W_IO/FrameStrobe[9] Tile_X0Y2_W_IO/UserCLK
+ Tile_X0Y1_W_IO/UserCLK VGND VPWR Tile_X0Y2_W_IO/W1END[0] Tile_X0Y2_W_IO/W1END[1]
+ Tile_X0Y2_W_IO/W1END[2] Tile_X0Y2_W_IO/W1END[3] Tile_X0Y2_W_IO/W2END[0] Tile_X0Y2_W_IO/W2END[1]
+ Tile_X0Y2_W_IO/W2END[2] Tile_X0Y2_W_IO/W2END[3] Tile_X0Y2_W_IO/W2END[4] Tile_X0Y2_W_IO/W2END[5]
+ Tile_X0Y2_W_IO/W2END[6] Tile_X0Y2_W_IO/W2END[7] Tile_X0Y2_W_IO/W2MID[0] Tile_X0Y2_W_IO/W2MID[1]
+ Tile_X0Y2_W_IO/W2MID[2] Tile_X0Y2_W_IO/W2MID[3] Tile_X0Y2_W_IO/W2MID[4] Tile_X0Y2_W_IO/W2MID[5]
+ Tile_X0Y2_W_IO/W2MID[6] Tile_X0Y2_W_IO/W2MID[7] Tile_X0Y2_W_IO/W6END[0] Tile_X0Y2_W_IO/W6END[10]
+ Tile_X0Y2_W_IO/W6END[11] Tile_X0Y2_W_IO/W6END[1] Tile_X0Y2_W_IO/W6END[2] Tile_X0Y2_W_IO/W6END[3]
+ Tile_X0Y2_W_IO/W6END[4] Tile_X0Y2_W_IO/W6END[5] Tile_X0Y2_W_IO/W6END[6] Tile_X0Y2_W_IO/W6END[7]
+ Tile_X0Y2_W_IO/W6END[8] Tile_X0Y2_W_IO/W6END[9] Tile_X0Y2_W_IO/WW4END[0] Tile_X0Y2_W_IO/WW4END[10]
+ Tile_X0Y2_W_IO/WW4END[11] Tile_X0Y2_W_IO/WW4END[12] Tile_X0Y2_W_IO/WW4END[13] Tile_X0Y2_W_IO/WW4END[14]
+ Tile_X0Y2_W_IO/WW4END[15] Tile_X0Y2_W_IO/WW4END[1] Tile_X0Y2_W_IO/WW4END[2] Tile_X0Y2_W_IO/WW4END[3]
+ Tile_X0Y2_W_IO/WW4END[4] Tile_X0Y2_W_IO/WW4END[5] Tile_X0Y2_W_IO/WW4END[6] Tile_X0Y2_W_IO/WW4END[7]
+ Tile_X0Y2_W_IO/WW4END[8] Tile_X0Y2_W_IO/WW4END[9] W_IO
XTile_X4Y2_RegFile Tile_X5Y2_LUT4AB/E1END[0] Tile_X5Y2_LUT4AB/E1END[1] Tile_X5Y2_LUT4AB/E1END[2]
+ Tile_X5Y2_LUT4AB/E1END[3] Tile_X3Y2_LUT4AB/E1BEG[0] Tile_X3Y2_LUT4AB/E1BEG[1] Tile_X3Y2_LUT4AB/E1BEG[2]
+ Tile_X3Y2_LUT4AB/E1BEG[3] Tile_X5Y2_LUT4AB/E2MID[0] Tile_X5Y2_LUT4AB/E2MID[1] Tile_X5Y2_LUT4AB/E2MID[2]
+ Tile_X5Y2_LUT4AB/E2MID[3] Tile_X5Y2_LUT4AB/E2MID[4] Tile_X5Y2_LUT4AB/E2MID[5] Tile_X5Y2_LUT4AB/E2MID[6]
+ Tile_X5Y2_LUT4AB/E2MID[7] Tile_X5Y2_LUT4AB/E2END[0] Tile_X5Y2_LUT4AB/E2END[1] Tile_X5Y2_LUT4AB/E2END[2]
+ Tile_X5Y2_LUT4AB/E2END[3] Tile_X5Y2_LUT4AB/E2END[4] Tile_X5Y2_LUT4AB/E2END[5] Tile_X5Y2_LUT4AB/E2END[6]
+ Tile_X5Y2_LUT4AB/E2END[7] Tile_X4Y2_RegFile/E2END[0] Tile_X4Y2_RegFile/E2END[1]
+ Tile_X4Y2_RegFile/E2END[2] Tile_X4Y2_RegFile/E2END[3] Tile_X4Y2_RegFile/E2END[4]
+ Tile_X4Y2_RegFile/E2END[5] Tile_X4Y2_RegFile/E2END[6] Tile_X4Y2_RegFile/E2END[7]
+ Tile_X3Y2_LUT4AB/E2BEG[0] Tile_X3Y2_LUT4AB/E2BEG[1] Tile_X3Y2_LUT4AB/E2BEG[2] Tile_X3Y2_LUT4AB/E2BEG[3]
+ Tile_X3Y2_LUT4AB/E2BEG[4] Tile_X3Y2_LUT4AB/E2BEG[5] Tile_X3Y2_LUT4AB/E2BEG[6] Tile_X3Y2_LUT4AB/E2BEG[7]
+ Tile_X5Y2_LUT4AB/E6END[0] Tile_X5Y2_LUT4AB/E6END[10] Tile_X5Y2_LUT4AB/E6END[11]
+ Tile_X5Y2_LUT4AB/E6END[1] Tile_X5Y2_LUT4AB/E6END[2] Tile_X5Y2_LUT4AB/E6END[3] Tile_X5Y2_LUT4AB/E6END[4]
+ Tile_X5Y2_LUT4AB/E6END[5] Tile_X5Y2_LUT4AB/E6END[6] Tile_X5Y2_LUT4AB/E6END[7] Tile_X5Y2_LUT4AB/E6END[8]
+ Tile_X5Y2_LUT4AB/E6END[9] Tile_X3Y2_LUT4AB/E6BEG[0] Tile_X3Y2_LUT4AB/E6BEG[10] Tile_X3Y2_LUT4AB/E6BEG[11]
+ Tile_X3Y2_LUT4AB/E6BEG[1] Tile_X3Y2_LUT4AB/E6BEG[2] Tile_X3Y2_LUT4AB/E6BEG[3] Tile_X3Y2_LUT4AB/E6BEG[4]
+ Tile_X3Y2_LUT4AB/E6BEG[5] Tile_X3Y2_LUT4AB/E6BEG[6] Tile_X3Y2_LUT4AB/E6BEG[7] Tile_X3Y2_LUT4AB/E6BEG[8]
+ Tile_X3Y2_LUT4AB/E6BEG[9] Tile_X5Y2_LUT4AB/EE4END[0] Tile_X5Y2_LUT4AB/EE4END[10]
+ Tile_X5Y2_LUT4AB/EE4END[11] Tile_X5Y2_LUT4AB/EE4END[12] Tile_X5Y2_LUT4AB/EE4END[13]
+ Tile_X5Y2_LUT4AB/EE4END[14] Tile_X5Y2_LUT4AB/EE4END[15] Tile_X5Y2_LUT4AB/EE4END[1]
+ Tile_X5Y2_LUT4AB/EE4END[2] Tile_X5Y2_LUT4AB/EE4END[3] Tile_X5Y2_LUT4AB/EE4END[4]
+ Tile_X5Y2_LUT4AB/EE4END[5] Tile_X5Y2_LUT4AB/EE4END[6] Tile_X5Y2_LUT4AB/EE4END[7]
+ Tile_X5Y2_LUT4AB/EE4END[8] Tile_X5Y2_LUT4AB/EE4END[9] Tile_X3Y2_LUT4AB/EE4BEG[0]
+ Tile_X3Y2_LUT4AB/EE4BEG[10] Tile_X3Y2_LUT4AB/EE4BEG[11] Tile_X3Y2_LUT4AB/EE4BEG[12]
+ Tile_X3Y2_LUT4AB/EE4BEG[13] Tile_X3Y2_LUT4AB/EE4BEG[14] Tile_X3Y2_LUT4AB/EE4BEG[15]
+ Tile_X3Y2_LUT4AB/EE4BEG[1] Tile_X3Y2_LUT4AB/EE4BEG[2] Tile_X3Y2_LUT4AB/EE4BEG[3]
+ Tile_X3Y2_LUT4AB/EE4BEG[4] Tile_X3Y2_LUT4AB/EE4BEG[5] Tile_X3Y2_LUT4AB/EE4BEG[6]
+ Tile_X3Y2_LUT4AB/EE4BEG[7] Tile_X3Y2_LUT4AB/EE4BEG[8] Tile_X3Y2_LUT4AB/EE4BEG[9]
+ Tile_X4Y2_RegFile/FrameData[0] Tile_X4Y2_RegFile/FrameData[10] Tile_X4Y2_RegFile/FrameData[11]
+ Tile_X4Y2_RegFile/FrameData[12] Tile_X4Y2_RegFile/FrameData[13] Tile_X4Y2_RegFile/FrameData[14]
+ Tile_X4Y2_RegFile/FrameData[15] Tile_X4Y2_RegFile/FrameData[16] Tile_X4Y2_RegFile/FrameData[17]
+ Tile_X4Y2_RegFile/FrameData[18] Tile_X4Y2_RegFile/FrameData[19] Tile_X4Y2_RegFile/FrameData[1]
+ Tile_X4Y2_RegFile/FrameData[20] Tile_X4Y2_RegFile/FrameData[21] Tile_X4Y2_RegFile/FrameData[22]
+ Tile_X4Y2_RegFile/FrameData[23] Tile_X4Y2_RegFile/FrameData[24] Tile_X4Y2_RegFile/FrameData[25]
+ Tile_X4Y2_RegFile/FrameData[26] Tile_X4Y2_RegFile/FrameData[27] Tile_X4Y2_RegFile/FrameData[28]
+ Tile_X4Y2_RegFile/FrameData[29] Tile_X4Y2_RegFile/FrameData[2] Tile_X4Y2_RegFile/FrameData[30]
+ Tile_X4Y2_RegFile/FrameData[31] Tile_X4Y2_RegFile/FrameData[3] Tile_X4Y2_RegFile/FrameData[4]
+ Tile_X4Y2_RegFile/FrameData[5] Tile_X4Y2_RegFile/FrameData[6] Tile_X4Y2_RegFile/FrameData[7]
+ Tile_X4Y2_RegFile/FrameData[8] Tile_X4Y2_RegFile/FrameData[9] Tile_X5Y2_LUT4AB/FrameData[0]
+ Tile_X5Y2_LUT4AB/FrameData[10] Tile_X5Y2_LUT4AB/FrameData[11] Tile_X5Y2_LUT4AB/FrameData[12]
+ Tile_X5Y2_LUT4AB/FrameData[13] Tile_X5Y2_LUT4AB/FrameData[14] Tile_X5Y2_LUT4AB/FrameData[15]
+ Tile_X5Y2_LUT4AB/FrameData[16] Tile_X5Y2_LUT4AB/FrameData[17] Tile_X5Y2_LUT4AB/FrameData[18]
+ Tile_X5Y2_LUT4AB/FrameData[19] Tile_X5Y2_LUT4AB/FrameData[1] Tile_X5Y2_LUT4AB/FrameData[20]
+ Tile_X5Y2_LUT4AB/FrameData[21] Tile_X5Y2_LUT4AB/FrameData[22] Tile_X5Y2_LUT4AB/FrameData[23]
+ Tile_X5Y2_LUT4AB/FrameData[24] Tile_X5Y2_LUT4AB/FrameData[25] Tile_X5Y2_LUT4AB/FrameData[26]
+ Tile_X5Y2_LUT4AB/FrameData[27] Tile_X5Y2_LUT4AB/FrameData[28] Tile_X5Y2_LUT4AB/FrameData[29]
+ Tile_X5Y2_LUT4AB/FrameData[2] Tile_X5Y2_LUT4AB/FrameData[30] Tile_X5Y2_LUT4AB/FrameData[31]
+ Tile_X5Y2_LUT4AB/FrameData[3] Tile_X5Y2_LUT4AB/FrameData[4] Tile_X5Y2_LUT4AB/FrameData[5]
+ Tile_X5Y2_LUT4AB/FrameData[6] Tile_X5Y2_LUT4AB/FrameData[7] Tile_X5Y2_LUT4AB/FrameData[8]
+ Tile_X5Y2_LUT4AB/FrameData[9] Tile_X4Y2_RegFile/FrameStrobe[0] Tile_X4Y2_RegFile/FrameStrobe[10]
+ Tile_X4Y2_RegFile/FrameStrobe[11] Tile_X4Y2_RegFile/FrameStrobe[12] Tile_X4Y2_RegFile/FrameStrobe[13]
+ Tile_X4Y2_RegFile/FrameStrobe[14] Tile_X4Y2_RegFile/FrameStrobe[15] Tile_X4Y2_RegFile/FrameStrobe[16]
+ Tile_X4Y2_RegFile/FrameStrobe[17] Tile_X4Y2_RegFile/FrameStrobe[18] Tile_X4Y2_RegFile/FrameStrobe[19]
+ Tile_X4Y2_RegFile/FrameStrobe[1] Tile_X4Y2_RegFile/FrameStrobe[2] Tile_X4Y2_RegFile/FrameStrobe[3]
+ Tile_X4Y2_RegFile/FrameStrobe[4] Tile_X4Y2_RegFile/FrameStrobe[5] Tile_X4Y2_RegFile/FrameStrobe[6]
+ Tile_X4Y2_RegFile/FrameStrobe[7] Tile_X4Y2_RegFile/FrameStrobe[8] Tile_X4Y2_RegFile/FrameStrobe[9]
+ Tile_X4Y1_RegFile/FrameStrobe[0] Tile_X4Y1_RegFile/FrameStrobe[10] Tile_X4Y1_RegFile/FrameStrobe[11]
+ Tile_X4Y1_RegFile/FrameStrobe[12] Tile_X4Y1_RegFile/FrameStrobe[13] Tile_X4Y1_RegFile/FrameStrobe[14]
+ Tile_X4Y1_RegFile/FrameStrobe[15] Tile_X4Y1_RegFile/FrameStrobe[16] Tile_X4Y1_RegFile/FrameStrobe[17]
+ Tile_X4Y1_RegFile/FrameStrobe[18] Tile_X4Y1_RegFile/FrameStrobe[19] Tile_X4Y1_RegFile/FrameStrobe[1]
+ Tile_X4Y1_RegFile/FrameStrobe[2] Tile_X4Y1_RegFile/FrameStrobe[3] Tile_X4Y1_RegFile/FrameStrobe[4]
+ Tile_X4Y1_RegFile/FrameStrobe[5] Tile_X4Y1_RegFile/FrameStrobe[6] Tile_X4Y1_RegFile/FrameStrobe[7]
+ Tile_X4Y1_RegFile/FrameStrobe[8] Tile_X4Y1_RegFile/FrameStrobe[9] Tile_X4Y2_RegFile/N1BEG[0]
+ Tile_X4Y2_RegFile/N1BEG[1] Tile_X4Y2_RegFile/N1BEG[2] Tile_X4Y2_RegFile/N1BEG[3]
+ Tile_X4Y3_RegFile/N1BEG[0] Tile_X4Y3_RegFile/N1BEG[1] Tile_X4Y3_RegFile/N1BEG[2]
+ Tile_X4Y3_RegFile/N1BEG[3] Tile_X4Y2_RegFile/N2BEG[0] Tile_X4Y2_RegFile/N2BEG[1]
+ Tile_X4Y2_RegFile/N2BEG[2] Tile_X4Y2_RegFile/N2BEG[3] Tile_X4Y2_RegFile/N2BEG[4]
+ Tile_X4Y2_RegFile/N2BEG[5] Tile_X4Y2_RegFile/N2BEG[6] Tile_X4Y2_RegFile/N2BEG[7]
+ Tile_X4Y1_RegFile/N2END[0] Tile_X4Y1_RegFile/N2END[1] Tile_X4Y1_RegFile/N2END[2]
+ Tile_X4Y1_RegFile/N2END[3] Tile_X4Y1_RegFile/N2END[4] Tile_X4Y1_RegFile/N2END[5]
+ Tile_X4Y1_RegFile/N2END[6] Tile_X4Y1_RegFile/N2END[7] Tile_X4Y2_RegFile/N2END[0]
+ Tile_X4Y2_RegFile/N2END[1] Tile_X4Y2_RegFile/N2END[2] Tile_X4Y2_RegFile/N2END[3]
+ Tile_X4Y2_RegFile/N2END[4] Tile_X4Y2_RegFile/N2END[5] Tile_X4Y2_RegFile/N2END[6]
+ Tile_X4Y2_RegFile/N2END[7] Tile_X4Y3_RegFile/N2BEG[0] Tile_X4Y3_RegFile/N2BEG[1]
+ Tile_X4Y3_RegFile/N2BEG[2] Tile_X4Y3_RegFile/N2BEG[3] Tile_X4Y3_RegFile/N2BEG[4]
+ Tile_X4Y3_RegFile/N2BEG[5] Tile_X4Y3_RegFile/N2BEG[6] Tile_X4Y3_RegFile/N2BEG[7]
+ Tile_X4Y2_RegFile/N4BEG[0] Tile_X4Y2_RegFile/N4BEG[10] Tile_X4Y2_RegFile/N4BEG[11]
+ Tile_X4Y2_RegFile/N4BEG[12] Tile_X4Y2_RegFile/N4BEG[13] Tile_X4Y2_RegFile/N4BEG[14]
+ Tile_X4Y2_RegFile/N4BEG[15] Tile_X4Y2_RegFile/N4BEG[1] Tile_X4Y2_RegFile/N4BEG[2]
+ Tile_X4Y2_RegFile/N4BEG[3] Tile_X4Y2_RegFile/N4BEG[4] Tile_X4Y2_RegFile/N4BEG[5]
+ Tile_X4Y2_RegFile/N4BEG[6] Tile_X4Y2_RegFile/N4BEG[7] Tile_X4Y2_RegFile/N4BEG[8]
+ Tile_X4Y2_RegFile/N4BEG[9] Tile_X4Y3_RegFile/N4BEG[0] Tile_X4Y3_RegFile/N4BEG[10]
+ Tile_X4Y3_RegFile/N4BEG[11] Tile_X4Y3_RegFile/N4BEG[12] Tile_X4Y3_RegFile/N4BEG[13]
+ Tile_X4Y3_RegFile/N4BEG[14] Tile_X4Y3_RegFile/N4BEG[15] Tile_X4Y3_RegFile/N4BEG[1]
+ Tile_X4Y3_RegFile/N4BEG[2] Tile_X4Y3_RegFile/N4BEG[3] Tile_X4Y3_RegFile/N4BEG[4]
+ Tile_X4Y3_RegFile/N4BEG[5] Tile_X4Y3_RegFile/N4BEG[6] Tile_X4Y3_RegFile/N4BEG[7]
+ Tile_X4Y3_RegFile/N4BEG[8] Tile_X4Y3_RegFile/N4BEG[9] Tile_X4Y2_RegFile/NN4BEG[0]
+ Tile_X4Y2_RegFile/NN4BEG[10] Tile_X4Y2_RegFile/NN4BEG[11] Tile_X4Y2_RegFile/NN4BEG[12]
+ Tile_X4Y2_RegFile/NN4BEG[13] Tile_X4Y2_RegFile/NN4BEG[14] Tile_X4Y2_RegFile/NN4BEG[15]
+ Tile_X4Y2_RegFile/NN4BEG[1] Tile_X4Y2_RegFile/NN4BEG[2] Tile_X4Y2_RegFile/NN4BEG[3]
+ Tile_X4Y2_RegFile/NN4BEG[4] Tile_X4Y2_RegFile/NN4BEG[5] Tile_X4Y2_RegFile/NN4BEG[6]
+ Tile_X4Y2_RegFile/NN4BEG[7] Tile_X4Y2_RegFile/NN4BEG[8] Tile_X4Y2_RegFile/NN4BEG[9]
+ Tile_X4Y3_RegFile/NN4BEG[0] Tile_X4Y3_RegFile/NN4BEG[10] Tile_X4Y3_RegFile/NN4BEG[11]
+ Tile_X4Y3_RegFile/NN4BEG[12] Tile_X4Y3_RegFile/NN4BEG[13] Tile_X4Y3_RegFile/NN4BEG[14]
+ Tile_X4Y3_RegFile/NN4BEG[15] Tile_X4Y3_RegFile/NN4BEG[1] Tile_X4Y3_RegFile/NN4BEG[2]
+ Tile_X4Y3_RegFile/NN4BEG[3] Tile_X4Y3_RegFile/NN4BEG[4] Tile_X4Y3_RegFile/NN4BEG[5]
+ Tile_X4Y3_RegFile/NN4BEG[6] Tile_X4Y3_RegFile/NN4BEG[7] Tile_X4Y3_RegFile/NN4BEG[8]
+ Tile_X4Y3_RegFile/NN4BEG[9] Tile_X4Y3_RegFile/S1END[0] Tile_X4Y3_RegFile/S1END[1]
+ Tile_X4Y3_RegFile/S1END[2] Tile_X4Y3_RegFile/S1END[3] Tile_X4Y2_RegFile/S1END[0]
+ Tile_X4Y2_RegFile/S1END[1] Tile_X4Y2_RegFile/S1END[2] Tile_X4Y2_RegFile/S1END[3]
+ Tile_X4Y3_RegFile/S2MID[0] Tile_X4Y3_RegFile/S2MID[1] Tile_X4Y3_RegFile/S2MID[2]
+ Tile_X4Y3_RegFile/S2MID[3] Tile_X4Y3_RegFile/S2MID[4] Tile_X4Y3_RegFile/S2MID[5]
+ Tile_X4Y3_RegFile/S2MID[6] Tile_X4Y3_RegFile/S2MID[7] Tile_X4Y3_RegFile/S2END[0]
+ Tile_X4Y3_RegFile/S2END[1] Tile_X4Y3_RegFile/S2END[2] Tile_X4Y3_RegFile/S2END[3]
+ Tile_X4Y3_RegFile/S2END[4] Tile_X4Y3_RegFile/S2END[5] Tile_X4Y3_RegFile/S2END[6]
+ Tile_X4Y3_RegFile/S2END[7] Tile_X4Y2_RegFile/S2END[0] Tile_X4Y2_RegFile/S2END[1]
+ Tile_X4Y2_RegFile/S2END[2] Tile_X4Y2_RegFile/S2END[3] Tile_X4Y2_RegFile/S2END[4]
+ Tile_X4Y2_RegFile/S2END[5] Tile_X4Y2_RegFile/S2END[6] Tile_X4Y2_RegFile/S2END[7]
+ Tile_X4Y2_RegFile/S2MID[0] Tile_X4Y2_RegFile/S2MID[1] Tile_X4Y2_RegFile/S2MID[2]
+ Tile_X4Y2_RegFile/S2MID[3] Tile_X4Y2_RegFile/S2MID[4] Tile_X4Y2_RegFile/S2MID[5]
+ Tile_X4Y2_RegFile/S2MID[6] Tile_X4Y2_RegFile/S2MID[7] Tile_X4Y3_RegFile/S4END[0]
+ Tile_X4Y3_RegFile/S4END[10] Tile_X4Y3_RegFile/S4END[11] Tile_X4Y3_RegFile/S4END[12]
+ Tile_X4Y3_RegFile/S4END[13] Tile_X4Y3_RegFile/S4END[14] Tile_X4Y3_RegFile/S4END[15]
+ Tile_X4Y3_RegFile/S4END[1] Tile_X4Y3_RegFile/S4END[2] Tile_X4Y3_RegFile/S4END[3]
+ Tile_X4Y3_RegFile/S4END[4] Tile_X4Y3_RegFile/S4END[5] Tile_X4Y3_RegFile/S4END[6]
+ Tile_X4Y3_RegFile/S4END[7] Tile_X4Y3_RegFile/S4END[8] Tile_X4Y3_RegFile/S4END[9]
+ Tile_X4Y2_RegFile/S4END[0] Tile_X4Y2_RegFile/S4END[10] Tile_X4Y2_RegFile/S4END[11]
+ Tile_X4Y2_RegFile/S4END[12] Tile_X4Y2_RegFile/S4END[13] Tile_X4Y2_RegFile/S4END[14]
+ Tile_X4Y2_RegFile/S4END[15] Tile_X4Y2_RegFile/S4END[1] Tile_X4Y2_RegFile/S4END[2]
+ Tile_X4Y2_RegFile/S4END[3] Tile_X4Y2_RegFile/S4END[4] Tile_X4Y2_RegFile/S4END[5]
+ Tile_X4Y2_RegFile/S4END[6] Tile_X4Y2_RegFile/S4END[7] Tile_X4Y2_RegFile/S4END[8]
+ Tile_X4Y2_RegFile/S4END[9] Tile_X4Y3_RegFile/SS4END[0] Tile_X4Y3_RegFile/SS4END[10]
+ Tile_X4Y3_RegFile/SS4END[11] Tile_X4Y3_RegFile/SS4END[12] Tile_X4Y3_RegFile/SS4END[13]
+ Tile_X4Y3_RegFile/SS4END[14] Tile_X4Y3_RegFile/SS4END[15] Tile_X4Y3_RegFile/SS4END[1]
+ Tile_X4Y3_RegFile/SS4END[2] Tile_X4Y3_RegFile/SS4END[3] Tile_X4Y3_RegFile/SS4END[4]
+ Tile_X4Y3_RegFile/SS4END[5] Tile_X4Y3_RegFile/SS4END[6] Tile_X4Y3_RegFile/SS4END[7]
+ Tile_X4Y3_RegFile/SS4END[8] Tile_X4Y3_RegFile/SS4END[9] Tile_X4Y2_RegFile/SS4END[0]
+ Tile_X4Y2_RegFile/SS4END[10] Tile_X4Y2_RegFile/SS4END[11] Tile_X4Y2_RegFile/SS4END[12]
+ Tile_X4Y2_RegFile/SS4END[13] Tile_X4Y2_RegFile/SS4END[14] Tile_X4Y2_RegFile/SS4END[15]
+ Tile_X4Y2_RegFile/SS4END[1] Tile_X4Y2_RegFile/SS4END[2] Tile_X4Y2_RegFile/SS4END[3]
+ Tile_X4Y2_RegFile/SS4END[4] Tile_X4Y2_RegFile/SS4END[5] Tile_X4Y2_RegFile/SS4END[6]
+ Tile_X4Y2_RegFile/SS4END[7] Tile_X4Y2_RegFile/SS4END[8] Tile_X4Y2_RegFile/SS4END[9]
+ Tile_X4Y2_RegFile/UserCLK Tile_X4Y1_RegFile/UserCLK VGND VPWR Tile_X3Y2_LUT4AB/W1END[0]
+ Tile_X3Y2_LUT4AB/W1END[1] Tile_X3Y2_LUT4AB/W1END[2] Tile_X3Y2_LUT4AB/W1END[3] Tile_X5Y2_LUT4AB/W1BEG[0]
+ Tile_X5Y2_LUT4AB/W1BEG[1] Tile_X5Y2_LUT4AB/W1BEG[2] Tile_X5Y2_LUT4AB/W1BEG[3] Tile_X3Y2_LUT4AB/W2MID[0]
+ Tile_X3Y2_LUT4AB/W2MID[1] Tile_X3Y2_LUT4AB/W2MID[2] Tile_X3Y2_LUT4AB/W2MID[3] Tile_X3Y2_LUT4AB/W2MID[4]
+ Tile_X3Y2_LUT4AB/W2MID[5] Tile_X3Y2_LUT4AB/W2MID[6] Tile_X3Y2_LUT4AB/W2MID[7] Tile_X3Y2_LUT4AB/W2END[0]
+ Tile_X3Y2_LUT4AB/W2END[1] Tile_X3Y2_LUT4AB/W2END[2] Tile_X3Y2_LUT4AB/W2END[3] Tile_X3Y2_LUT4AB/W2END[4]
+ Tile_X3Y2_LUT4AB/W2END[5] Tile_X3Y2_LUT4AB/W2END[6] Tile_X3Y2_LUT4AB/W2END[7] Tile_X5Y2_LUT4AB/W2BEGb[0]
+ Tile_X5Y2_LUT4AB/W2BEGb[1] Tile_X5Y2_LUT4AB/W2BEGb[2] Tile_X5Y2_LUT4AB/W2BEGb[3]
+ Tile_X5Y2_LUT4AB/W2BEGb[4] Tile_X5Y2_LUT4AB/W2BEGb[5] Tile_X5Y2_LUT4AB/W2BEGb[6]
+ Tile_X5Y2_LUT4AB/W2BEGb[7] Tile_X5Y2_LUT4AB/W2BEG[0] Tile_X5Y2_LUT4AB/W2BEG[1] Tile_X5Y2_LUT4AB/W2BEG[2]
+ Tile_X5Y2_LUT4AB/W2BEG[3] Tile_X5Y2_LUT4AB/W2BEG[4] Tile_X5Y2_LUT4AB/W2BEG[5] Tile_X5Y2_LUT4AB/W2BEG[6]
+ Tile_X5Y2_LUT4AB/W2BEG[7] Tile_X3Y2_LUT4AB/W6END[0] Tile_X3Y2_LUT4AB/W6END[10] Tile_X3Y2_LUT4AB/W6END[11]
+ Tile_X3Y2_LUT4AB/W6END[1] Tile_X3Y2_LUT4AB/W6END[2] Tile_X3Y2_LUT4AB/W6END[3] Tile_X3Y2_LUT4AB/W6END[4]
+ Tile_X3Y2_LUT4AB/W6END[5] Tile_X3Y2_LUT4AB/W6END[6] Tile_X3Y2_LUT4AB/W6END[7] Tile_X3Y2_LUT4AB/W6END[8]
+ Tile_X3Y2_LUT4AB/W6END[9] Tile_X5Y2_LUT4AB/W6BEG[0] Tile_X5Y2_LUT4AB/W6BEG[10] Tile_X5Y2_LUT4AB/W6BEG[11]
+ Tile_X5Y2_LUT4AB/W6BEG[1] Tile_X5Y2_LUT4AB/W6BEG[2] Tile_X5Y2_LUT4AB/W6BEG[3] Tile_X5Y2_LUT4AB/W6BEG[4]
+ Tile_X5Y2_LUT4AB/W6BEG[5] Tile_X5Y2_LUT4AB/W6BEG[6] Tile_X5Y2_LUT4AB/W6BEG[7] Tile_X5Y2_LUT4AB/W6BEG[8]
+ Tile_X5Y2_LUT4AB/W6BEG[9] Tile_X3Y2_LUT4AB/WW4END[0] Tile_X3Y2_LUT4AB/WW4END[10]
+ Tile_X3Y2_LUT4AB/WW4END[11] Tile_X3Y2_LUT4AB/WW4END[12] Tile_X3Y2_LUT4AB/WW4END[13]
+ Tile_X3Y2_LUT4AB/WW4END[14] Tile_X3Y2_LUT4AB/WW4END[15] Tile_X3Y2_LUT4AB/WW4END[1]
+ Tile_X3Y2_LUT4AB/WW4END[2] Tile_X3Y2_LUT4AB/WW4END[3] Tile_X3Y2_LUT4AB/WW4END[4]
+ Tile_X3Y2_LUT4AB/WW4END[5] Tile_X3Y2_LUT4AB/WW4END[6] Tile_X3Y2_LUT4AB/WW4END[7]
+ Tile_X3Y2_LUT4AB/WW4END[8] Tile_X3Y2_LUT4AB/WW4END[9] Tile_X5Y2_LUT4AB/WW4BEG[0]
+ Tile_X5Y2_LUT4AB/WW4BEG[10] Tile_X5Y2_LUT4AB/WW4BEG[11] Tile_X5Y2_LUT4AB/WW4BEG[12]
+ Tile_X5Y2_LUT4AB/WW4BEG[13] Tile_X5Y2_LUT4AB/WW4BEG[14] Tile_X5Y2_LUT4AB/WW4BEG[15]
+ Tile_X5Y2_LUT4AB/WW4BEG[1] Tile_X5Y2_LUT4AB/WW4BEG[2] Tile_X5Y2_LUT4AB/WW4BEG[3]
+ Tile_X5Y2_LUT4AB/WW4BEG[4] Tile_X5Y2_LUT4AB/WW4BEG[5] Tile_X5Y2_LUT4AB/WW4BEG[6]
+ Tile_X5Y2_LUT4AB/WW4BEG[7] Tile_X5Y2_LUT4AB/WW4BEG[8] Tile_X5Y2_LUT4AB/WW4BEG[9]
+ RegFile
XTile_X9Y9_LUT4AB Tile_X9Y9_LUT4AB/Ci Tile_X9Y9_LUT4AB/Co Tile_X9Y9_LUT4AB/E1BEG[0]
+ Tile_X9Y9_LUT4AB/E1BEG[1] Tile_X9Y9_LUT4AB/E1BEG[2] Tile_X9Y9_LUT4AB/E1BEG[3] Tile_X9Y9_LUT4AB/E1END[0]
+ Tile_X9Y9_LUT4AB/E1END[1] Tile_X9Y9_LUT4AB/E1END[2] Tile_X9Y9_LUT4AB/E1END[3] Tile_X9Y9_LUT4AB/E2BEG[0]
+ Tile_X9Y9_LUT4AB/E2BEG[1] Tile_X9Y9_LUT4AB/E2BEG[2] Tile_X9Y9_LUT4AB/E2BEG[3] Tile_X9Y9_LUT4AB/E2BEG[4]
+ Tile_X9Y9_LUT4AB/E2BEG[5] Tile_X9Y9_LUT4AB/E2BEG[6] Tile_X9Y9_LUT4AB/E2BEG[7] Tile_X9Y9_LUT4AB/E2BEGb[0]
+ Tile_X9Y9_LUT4AB/E2BEGb[1] Tile_X9Y9_LUT4AB/E2BEGb[2] Tile_X9Y9_LUT4AB/E2BEGb[3]
+ Tile_X9Y9_LUT4AB/E2BEGb[4] Tile_X9Y9_LUT4AB/E2BEGb[5] Tile_X9Y9_LUT4AB/E2BEGb[6]
+ Tile_X9Y9_LUT4AB/E2BEGb[7] Tile_X9Y9_LUT4AB/E2END[0] Tile_X9Y9_LUT4AB/E2END[1] Tile_X9Y9_LUT4AB/E2END[2]
+ Tile_X9Y9_LUT4AB/E2END[3] Tile_X9Y9_LUT4AB/E2END[4] Tile_X9Y9_LUT4AB/E2END[5] Tile_X9Y9_LUT4AB/E2END[6]
+ Tile_X9Y9_LUT4AB/E2END[7] Tile_X9Y9_LUT4AB/E2MID[0] Tile_X9Y9_LUT4AB/E2MID[1] Tile_X9Y9_LUT4AB/E2MID[2]
+ Tile_X9Y9_LUT4AB/E2MID[3] Tile_X9Y9_LUT4AB/E2MID[4] Tile_X9Y9_LUT4AB/E2MID[5] Tile_X9Y9_LUT4AB/E2MID[6]
+ Tile_X9Y9_LUT4AB/E2MID[7] Tile_X9Y9_LUT4AB/E6BEG[0] Tile_X9Y9_LUT4AB/E6BEG[10] Tile_X9Y9_LUT4AB/E6BEG[11]
+ Tile_X9Y9_LUT4AB/E6BEG[1] Tile_X9Y9_LUT4AB/E6BEG[2] Tile_X9Y9_LUT4AB/E6BEG[3] Tile_X9Y9_LUT4AB/E6BEG[4]
+ Tile_X9Y9_LUT4AB/E6BEG[5] Tile_X9Y9_LUT4AB/E6BEG[6] Tile_X9Y9_LUT4AB/E6BEG[7] Tile_X9Y9_LUT4AB/E6BEG[8]
+ Tile_X9Y9_LUT4AB/E6BEG[9] Tile_X9Y9_LUT4AB/E6END[0] Tile_X9Y9_LUT4AB/E6END[10] Tile_X9Y9_LUT4AB/E6END[11]
+ Tile_X9Y9_LUT4AB/E6END[1] Tile_X9Y9_LUT4AB/E6END[2] Tile_X9Y9_LUT4AB/E6END[3] Tile_X9Y9_LUT4AB/E6END[4]
+ Tile_X9Y9_LUT4AB/E6END[5] Tile_X9Y9_LUT4AB/E6END[6] Tile_X9Y9_LUT4AB/E6END[7] Tile_X9Y9_LUT4AB/E6END[8]
+ Tile_X9Y9_LUT4AB/E6END[9] Tile_X9Y9_LUT4AB/EE4BEG[0] Tile_X9Y9_LUT4AB/EE4BEG[10]
+ Tile_X9Y9_LUT4AB/EE4BEG[11] Tile_X9Y9_LUT4AB/EE4BEG[12] Tile_X9Y9_LUT4AB/EE4BEG[13]
+ Tile_X9Y9_LUT4AB/EE4BEG[14] Tile_X9Y9_LUT4AB/EE4BEG[15] Tile_X9Y9_LUT4AB/EE4BEG[1]
+ Tile_X9Y9_LUT4AB/EE4BEG[2] Tile_X9Y9_LUT4AB/EE4BEG[3] Tile_X9Y9_LUT4AB/EE4BEG[4]
+ Tile_X9Y9_LUT4AB/EE4BEG[5] Tile_X9Y9_LUT4AB/EE4BEG[6] Tile_X9Y9_LUT4AB/EE4BEG[7]
+ Tile_X9Y9_LUT4AB/EE4BEG[8] Tile_X9Y9_LUT4AB/EE4BEG[9] Tile_X9Y9_LUT4AB/EE4END[0]
+ Tile_X9Y9_LUT4AB/EE4END[10] Tile_X9Y9_LUT4AB/EE4END[11] Tile_X9Y9_LUT4AB/EE4END[12]
+ Tile_X9Y9_LUT4AB/EE4END[13] Tile_X9Y9_LUT4AB/EE4END[14] Tile_X9Y9_LUT4AB/EE4END[15]
+ Tile_X9Y9_LUT4AB/EE4END[1] Tile_X9Y9_LUT4AB/EE4END[2] Tile_X9Y9_LUT4AB/EE4END[3]
+ Tile_X9Y9_LUT4AB/EE4END[4] Tile_X9Y9_LUT4AB/EE4END[5] Tile_X9Y9_LUT4AB/EE4END[6]
+ Tile_X9Y9_LUT4AB/EE4END[7] Tile_X9Y9_LUT4AB/EE4END[8] Tile_X9Y9_LUT4AB/EE4END[9]
+ Tile_X9Y9_LUT4AB/FrameData[0] Tile_X9Y9_LUT4AB/FrameData[10] Tile_X9Y9_LUT4AB/FrameData[11]
+ Tile_X9Y9_LUT4AB/FrameData[12] Tile_X9Y9_LUT4AB/FrameData[13] Tile_X9Y9_LUT4AB/FrameData[14]
+ Tile_X9Y9_LUT4AB/FrameData[15] Tile_X9Y9_LUT4AB/FrameData[16] Tile_X9Y9_LUT4AB/FrameData[17]
+ Tile_X9Y9_LUT4AB/FrameData[18] Tile_X9Y9_LUT4AB/FrameData[19] Tile_X9Y9_LUT4AB/FrameData[1]
+ Tile_X9Y9_LUT4AB/FrameData[20] Tile_X9Y9_LUT4AB/FrameData[21] Tile_X9Y9_LUT4AB/FrameData[22]
+ Tile_X9Y9_LUT4AB/FrameData[23] Tile_X9Y9_LUT4AB/FrameData[24] Tile_X9Y9_LUT4AB/FrameData[25]
+ Tile_X9Y9_LUT4AB/FrameData[26] Tile_X9Y9_LUT4AB/FrameData[27] Tile_X9Y9_LUT4AB/FrameData[28]
+ Tile_X9Y9_LUT4AB/FrameData[29] Tile_X9Y9_LUT4AB/FrameData[2] Tile_X9Y9_LUT4AB/FrameData[30]
+ Tile_X9Y9_LUT4AB/FrameData[31] Tile_X9Y9_LUT4AB/FrameData[3] Tile_X9Y9_LUT4AB/FrameData[4]
+ Tile_X9Y9_LUT4AB/FrameData[5] Tile_X9Y9_LUT4AB/FrameData[6] Tile_X9Y9_LUT4AB/FrameData[7]
+ Tile_X9Y9_LUT4AB/FrameData[8] Tile_X9Y9_LUT4AB/FrameData[9] Tile_X9Y9_LUT4AB/FrameData_O[0]
+ Tile_X9Y9_LUT4AB/FrameData_O[10] Tile_X9Y9_LUT4AB/FrameData_O[11] Tile_X9Y9_LUT4AB/FrameData_O[12]
+ Tile_X9Y9_LUT4AB/FrameData_O[13] Tile_X9Y9_LUT4AB/FrameData_O[14] Tile_X9Y9_LUT4AB/FrameData_O[15]
+ Tile_X9Y9_LUT4AB/FrameData_O[16] Tile_X9Y9_LUT4AB/FrameData_O[17] Tile_X9Y9_LUT4AB/FrameData_O[18]
+ Tile_X9Y9_LUT4AB/FrameData_O[19] Tile_X9Y9_LUT4AB/FrameData_O[1] Tile_X9Y9_LUT4AB/FrameData_O[20]
+ Tile_X9Y9_LUT4AB/FrameData_O[21] Tile_X9Y9_LUT4AB/FrameData_O[22] Tile_X9Y9_LUT4AB/FrameData_O[23]
+ Tile_X9Y9_LUT4AB/FrameData_O[24] Tile_X9Y9_LUT4AB/FrameData_O[25] Tile_X9Y9_LUT4AB/FrameData_O[26]
+ Tile_X9Y9_LUT4AB/FrameData_O[27] Tile_X9Y9_LUT4AB/FrameData_O[28] Tile_X9Y9_LUT4AB/FrameData_O[29]
+ Tile_X9Y9_LUT4AB/FrameData_O[2] Tile_X9Y9_LUT4AB/FrameData_O[30] Tile_X9Y9_LUT4AB/FrameData_O[31]
+ Tile_X9Y9_LUT4AB/FrameData_O[3] Tile_X9Y9_LUT4AB/FrameData_O[4] Tile_X9Y9_LUT4AB/FrameData_O[5]
+ Tile_X9Y9_LUT4AB/FrameData_O[6] Tile_X9Y9_LUT4AB/FrameData_O[7] Tile_X9Y9_LUT4AB/FrameData_O[8]
+ Tile_X9Y9_LUT4AB/FrameData_O[9] Tile_X9Y9_LUT4AB/FrameStrobe[0] Tile_X9Y9_LUT4AB/FrameStrobe[10]
+ Tile_X9Y9_LUT4AB/FrameStrobe[11] Tile_X9Y9_LUT4AB/FrameStrobe[12] Tile_X9Y9_LUT4AB/FrameStrobe[13]
+ Tile_X9Y9_LUT4AB/FrameStrobe[14] Tile_X9Y9_LUT4AB/FrameStrobe[15] Tile_X9Y9_LUT4AB/FrameStrobe[16]
+ Tile_X9Y9_LUT4AB/FrameStrobe[17] Tile_X9Y9_LUT4AB/FrameStrobe[18] Tile_X9Y9_LUT4AB/FrameStrobe[19]
+ Tile_X9Y9_LUT4AB/FrameStrobe[1] Tile_X9Y9_LUT4AB/FrameStrobe[2] Tile_X9Y9_LUT4AB/FrameStrobe[3]
+ Tile_X9Y9_LUT4AB/FrameStrobe[4] Tile_X9Y9_LUT4AB/FrameStrobe[5] Tile_X9Y9_LUT4AB/FrameStrobe[6]
+ Tile_X9Y9_LUT4AB/FrameStrobe[7] Tile_X9Y9_LUT4AB/FrameStrobe[8] Tile_X9Y9_LUT4AB/FrameStrobe[9]
+ Tile_X9Y8_LUT4AB/FrameStrobe[0] Tile_X9Y8_LUT4AB/FrameStrobe[10] Tile_X9Y8_LUT4AB/FrameStrobe[11]
+ Tile_X9Y8_LUT4AB/FrameStrobe[12] Tile_X9Y8_LUT4AB/FrameStrobe[13] Tile_X9Y8_LUT4AB/FrameStrobe[14]
+ Tile_X9Y8_LUT4AB/FrameStrobe[15] Tile_X9Y8_LUT4AB/FrameStrobe[16] Tile_X9Y8_LUT4AB/FrameStrobe[17]
+ Tile_X9Y8_LUT4AB/FrameStrobe[18] Tile_X9Y8_LUT4AB/FrameStrobe[19] Tile_X9Y8_LUT4AB/FrameStrobe[1]
+ Tile_X9Y8_LUT4AB/FrameStrobe[2] Tile_X9Y8_LUT4AB/FrameStrobe[3] Tile_X9Y8_LUT4AB/FrameStrobe[4]
+ Tile_X9Y8_LUT4AB/FrameStrobe[5] Tile_X9Y8_LUT4AB/FrameStrobe[6] Tile_X9Y8_LUT4AB/FrameStrobe[7]
+ Tile_X9Y8_LUT4AB/FrameStrobe[8] Tile_X9Y8_LUT4AB/FrameStrobe[9] Tile_X9Y9_LUT4AB/N1BEG[0]
+ Tile_X9Y9_LUT4AB/N1BEG[1] Tile_X9Y9_LUT4AB/N1BEG[2] Tile_X9Y9_LUT4AB/N1BEG[3] Tile_X9Y9_LUT4AB/N1END[0]
+ Tile_X9Y9_LUT4AB/N1END[1] Tile_X9Y9_LUT4AB/N1END[2] Tile_X9Y9_LUT4AB/N1END[3] Tile_X9Y9_LUT4AB/N2BEG[0]
+ Tile_X9Y9_LUT4AB/N2BEG[1] Tile_X9Y9_LUT4AB/N2BEG[2] Tile_X9Y9_LUT4AB/N2BEG[3] Tile_X9Y9_LUT4AB/N2BEG[4]
+ Tile_X9Y9_LUT4AB/N2BEG[5] Tile_X9Y9_LUT4AB/N2BEG[6] Tile_X9Y9_LUT4AB/N2BEG[7] Tile_X9Y8_LUT4AB/N2END[0]
+ Tile_X9Y8_LUT4AB/N2END[1] Tile_X9Y8_LUT4AB/N2END[2] Tile_X9Y8_LUT4AB/N2END[3] Tile_X9Y8_LUT4AB/N2END[4]
+ Tile_X9Y8_LUT4AB/N2END[5] Tile_X9Y8_LUT4AB/N2END[6] Tile_X9Y8_LUT4AB/N2END[7] Tile_X9Y9_LUT4AB/N2END[0]
+ Tile_X9Y9_LUT4AB/N2END[1] Tile_X9Y9_LUT4AB/N2END[2] Tile_X9Y9_LUT4AB/N2END[3] Tile_X9Y9_LUT4AB/N2END[4]
+ Tile_X9Y9_LUT4AB/N2END[5] Tile_X9Y9_LUT4AB/N2END[6] Tile_X9Y9_LUT4AB/N2END[7] Tile_X9Y9_LUT4AB/N2MID[0]
+ Tile_X9Y9_LUT4AB/N2MID[1] Tile_X9Y9_LUT4AB/N2MID[2] Tile_X9Y9_LUT4AB/N2MID[3] Tile_X9Y9_LUT4AB/N2MID[4]
+ Tile_X9Y9_LUT4AB/N2MID[5] Tile_X9Y9_LUT4AB/N2MID[6] Tile_X9Y9_LUT4AB/N2MID[7] Tile_X9Y9_LUT4AB/N4BEG[0]
+ Tile_X9Y9_LUT4AB/N4BEG[10] Tile_X9Y9_LUT4AB/N4BEG[11] Tile_X9Y9_LUT4AB/N4BEG[12]
+ Tile_X9Y9_LUT4AB/N4BEG[13] Tile_X9Y9_LUT4AB/N4BEG[14] Tile_X9Y9_LUT4AB/N4BEG[15]
+ Tile_X9Y9_LUT4AB/N4BEG[1] Tile_X9Y9_LUT4AB/N4BEG[2] Tile_X9Y9_LUT4AB/N4BEG[3] Tile_X9Y9_LUT4AB/N4BEG[4]
+ Tile_X9Y9_LUT4AB/N4BEG[5] Tile_X9Y9_LUT4AB/N4BEG[6] Tile_X9Y9_LUT4AB/N4BEG[7] Tile_X9Y9_LUT4AB/N4BEG[8]
+ Tile_X9Y9_LUT4AB/N4BEG[9] Tile_X9Y9_LUT4AB/N4END[0] Tile_X9Y9_LUT4AB/N4END[10] Tile_X9Y9_LUT4AB/N4END[11]
+ Tile_X9Y9_LUT4AB/N4END[12] Tile_X9Y9_LUT4AB/N4END[13] Tile_X9Y9_LUT4AB/N4END[14]
+ Tile_X9Y9_LUT4AB/N4END[15] Tile_X9Y9_LUT4AB/N4END[1] Tile_X9Y9_LUT4AB/N4END[2] Tile_X9Y9_LUT4AB/N4END[3]
+ Tile_X9Y9_LUT4AB/N4END[4] Tile_X9Y9_LUT4AB/N4END[5] Tile_X9Y9_LUT4AB/N4END[6] Tile_X9Y9_LUT4AB/N4END[7]
+ Tile_X9Y9_LUT4AB/N4END[8] Tile_X9Y9_LUT4AB/N4END[9] Tile_X9Y9_LUT4AB/NN4BEG[0] Tile_X9Y9_LUT4AB/NN4BEG[10]
+ Tile_X9Y9_LUT4AB/NN4BEG[11] Tile_X9Y9_LUT4AB/NN4BEG[12] Tile_X9Y9_LUT4AB/NN4BEG[13]
+ Tile_X9Y9_LUT4AB/NN4BEG[14] Tile_X9Y9_LUT4AB/NN4BEG[15] Tile_X9Y9_LUT4AB/NN4BEG[1]
+ Tile_X9Y9_LUT4AB/NN4BEG[2] Tile_X9Y9_LUT4AB/NN4BEG[3] Tile_X9Y9_LUT4AB/NN4BEG[4]
+ Tile_X9Y9_LUT4AB/NN4BEG[5] Tile_X9Y9_LUT4AB/NN4BEG[6] Tile_X9Y9_LUT4AB/NN4BEG[7]
+ Tile_X9Y9_LUT4AB/NN4BEG[8] Tile_X9Y9_LUT4AB/NN4BEG[9] Tile_X9Y9_LUT4AB/NN4END[0]
+ Tile_X9Y9_LUT4AB/NN4END[10] Tile_X9Y9_LUT4AB/NN4END[11] Tile_X9Y9_LUT4AB/NN4END[12]
+ Tile_X9Y9_LUT4AB/NN4END[13] Tile_X9Y9_LUT4AB/NN4END[14] Tile_X9Y9_LUT4AB/NN4END[15]
+ Tile_X9Y9_LUT4AB/NN4END[1] Tile_X9Y9_LUT4AB/NN4END[2] Tile_X9Y9_LUT4AB/NN4END[3]
+ Tile_X9Y9_LUT4AB/NN4END[4] Tile_X9Y9_LUT4AB/NN4END[5] Tile_X9Y9_LUT4AB/NN4END[6]
+ Tile_X9Y9_LUT4AB/NN4END[7] Tile_X9Y9_LUT4AB/NN4END[8] Tile_X9Y9_LUT4AB/NN4END[9]
+ Tile_X9Y9_LUT4AB/S1BEG[0] Tile_X9Y9_LUT4AB/S1BEG[1] Tile_X9Y9_LUT4AB/S1BEG[2] Tile_X9Y9_LUT4AB/S1BEG[3]
+ Tile_X9Y9_LUT4AB/S1END[0] Tile_X9Y9_LUT4AB/S1END[1] Tile_X9Y9_LUT4AB/S1END[2] Tile_X9Y9_LUT4AB/S1END[3]
+ Tile_X9Y9_LUT4AB/S2BEG[0] Tile_X9Y9_LUT4AB/S2BEG[1] Tile_X9Y9_LUT4AB/S2BEG[2] Tile_X9Y9_LUT4AB/S2BEG[3]
+ Tile_X9Y9_LUT4AB/S2BEG[4] Tile_X9Y9_LUT4AB/S2BEG[5] Tile_X9Y9_LUT4AB/S2BEG[6] Tile_X9Y9_LUT4AB/S2BEG[7]
+ Tile_X9Y9_LUT4AB/S2BEGb[0] Tile_X9Y9_LUT4AB/S2BEGb[1] Tile_X9Y9_LUT4AB/S2BEGb[2]
+ Tile_X9Y9_LUT4AB/S2BEGb[3] Tile_X9Y9_LUT4AB/S2BEGb[4] Tile_X9Y9_LUT4AB/S2BEGb[5]
+ Tile_X9Y9_LUT4AB/S2BEGb[6] Tile_X9Y9_LUT4AB/S2BEGb[7] Tile_X9Y9_LUT4AB/S2END[0]
+ Tile_X9Y9_LUT4AB/S2END[1] Tile_X9Y9_LUT4AB/S2END[2] Tile_X9Y9_LUT4AB/S2END[3] Tile_X9Y9_LUT4AB/S2END[4]
+ Tile_X9Y9_LUT4AB/S2END[5] Tile_X9Y9_LUT4AB/S2END[6] Tile_X9Y9_LUT4AB/S2END[7] Tile_X9Y9_LUT4AB/S2MID[0]
+ Tile_X9Y9_LUT4AB/S2MID[1] Tile_X9Y9_LUT4AB/S2MID[2] Tile_X9Y9_LUT4AB/S2MID[3] Tile_X9Y9_LUT4AB/S2MID[4]
+ Tile_X9Y9_LUT4AB/S2MID[5] Tile_X9Y9_LUT4AB/S2MID[6] Tile_X9Y9_LUT4AB/S2MID[7] Tile_X9Y9_LUT4AB/S4BEG[0]
+ Tile_X9Y9_LUT4AB/S4BEG[10] Tile_X9Y9_LUT4AB/S4BEG[11] Tile_X9Y9_LUT4AB/S4BEG[12]
+ Tile_X9Y9_LUT4AB/S4BEG[13] Tile_X9Y9_LUT4AB/S4BEG[14] Tile_X9Y9_LUT4AB/S4BEG[15]
+ Tile_X9Y9_LUT4AB/S4BEG[1] Tile_X9Y9_LUT4AB/S4BEG[2] Tile_X9Y9_LUT4AB/S4BEG[3] Tile_X9Y9_LUT4AB/S4BEG[4]
+ Tile_X9Y9_LUT4AB/S4BEG[5] Tile_X9Y9_LUT4AB/S4BEG[6] Tile_X9Y9_LUT4AB/S4BEG[7] Tile_X9Y9_LUT4AB/S4BEG[8]
+ Tile_X9Y9_LUT4AB/S4BEG[9] Tile_X9Y9_LUT4AB/S4END[0] Tile_X9Y9_LUT4AB/S4END[10] Tile_X9Y9_LUT4AB/S4END[11]
+ Tile_X9Y9_LUT4AB/S4END[12] Tile_X9Y9_LUT4AB/S4END[13] Tile_X9Y9_LUT4AB/S4END[14]
+ Tile_X9Y9_LUT4AB/S4END[15] Tile_X9Y9_LUT4AB/S4END[1] Tile_X9Y9_LUT4AB/S4END[2] Tile_X9Y9_LUT4AB/S4END[3]
+ Tile_X9Y9_LUT4AB/S4END[4] Tile_X9Y9_LUT4AB/S4END[5] Tile_X9Y9_LUT4AB/S4END[6] Tile_X9Y9_LUT4AB/S4END[7]
+ Tile_X9Y9_LUT4AB/S4END[8] Tile_X9Y9_LUT4AB/S4END[9] Tile_X9Y9_LUT4AB/SS4BEG[0] Tile_X9Y9_LUT4AB/SS4BEG[10]
+ Tile_X9Y9_LUT4AB/SS4BEG[11] Tile_X9Y9_LUT4AB/SS4BEG[12] Tile_X9Y9_LUT4AB/SS4BEG[13]
+ Tile_X9Y9_LUT4AB/SS4BEG[14] Tile_X9Y9_LUT4AB/SS4BEG[15] Tile_X9Y9_LUT4AB/SS4BEG[1]
+ Tile_X9Y9_LUT4AB/SS4BEG[2] Tile_X9Y9_LUT4AB/SS4BEG[3] Tile_X9Y9_LUT4AB/SS4BEG[4]
+ Tile_X9Y9_LUT4AB/SS4BEG[5] Tile_X9Y9_LUT4AB/SS4BEG[6] Tile_X9Y9_LUT4AB/SS4BEG[7]
+ Tile_X9Y9_LUT4AB/SS4BEG[8] Tile_X9Y9_LUT4AB/SS4BEG[9] Tile_X9Y9_LUT4AB/SS4END[0]
+ Tile_X9Y9_LUT4AB/SS4END[10] Tile_X9Y9_LUT4AB/SS4END[11] Tile_X9Y9_LUT4AB/SS4END[12]
+ Tile_X9Y9_LUT4AB/SS4END[13] Tile_X9Y9_LUT4AB/SS4END[14] Tile_X9Y9_LUT4AB/SS4END[15]
+ Tile_X9Y9_LUT4AB/SS4END[1] Tile_X9Y9_LUT4AB/SS4END[2] Tile_X9Y9_LUT4AB/SS4END[3]
+ Tile_X9Y9_LUT4AB/SS4END[4] Tile_X9Y9_LUT4AB/SS4END[5] Tile_X9Y9_LUT4AB/SS4END[6]
+ Tile_X9Y9_LUT4AB/SS4END[7] Tile_X9Y9_LUT4AB/SS4END[8] Tile_X9Y9_LUT4AB/SS4END[9]
+ Tile_X9Y9_LUT4AB/UserCLK Tile_X9Y8_LUT4AB/UserCLK VGND VPWR Tile_X9Y9_LUT4AB/W1BEG[0]
+ Tile_X9Y9_LUT4AB/W1BEG[1] Tile_X9Y9_LUT4AB/W1BEG[2] Tile_X9Y9_LUT4AB/W1BEG[3] Tile_X9Y9_LUT4AB/W1END[0]
+ Tile_X9Y9_LUT4AB/W1END[1] Tile_X9Y9_LUT4AB/W1END[2] Tile_X9Y9_LUT4AB/W1END[3] Tile_X9Y9_LUT4AB/W2BEG[0]
+ Tile_X9Y9_LUT4AB/W2BEG[1] Tile_X9Y9_LUT4AB/W2BEG[2] Tile_X9Y9_LUT4AB/W2BEG[3] Tile_X9Y9_LUT4AB/W2BEG[4]
+ Tile_X9Y9_LUT4AB/W2BEG[5] Tile_X9Y9_LUT4AB/W2BEG[6] Tile_X9Y9_LUT4AB/W2BEG[7] Tile_X8Y9_LUT4AB/W2END[0]
+ Tile_X8Y9_LUT4AB/W2END[1] Tile_X8Y9_LUT4AB/W2END[2] Tile_X8Y9_LUT4AB/W2END[3] Tile_X8Y9_LUT4AB/W2END[4]
+ Tile_X8Y9_LUT4AB/W2END[5] Tile_X8Y9_LUT4AB/W2END[6] Tile_X8Y9_LUT4AB/W2END[7] Tile_X9Y9_LUT4AB/W2END[0]
+ Tile_X9Y9_LUT4AB/W2END[1] Tile_X9Y9_LUT4AB/W2END[2] Tile_X9Y9_LUT4AB/W2END[3] Tile_X9Y9_LUT4AB/W2END[4]
+ Tile_X9Y9_LUT4AB/W2END[5] Tile_X9Y9_LUT4AB/W2END[6] Tile_X9Y9_LUT4AB/W2END[7] Tile_X9Y9_LUT4AB/W2MID[0]
+ Tile_X9Y9_LUT4AB/W2MID[1] Tile_X9Y9_LUT4AB/W2MID[2] Tile_X9Y9_LUT4AB/W2MID[3] Tile_X9Y9_LUT4AB/W2MID[4]
+ Tile_X9Y9_LUT4AB/W2MID[5] Tile_X9Y9_LUT4AB/W2MID[6] Tile_X9Y9_LUT4AB/W2MID[7] Tile_X9Y9_LUT4AB/W6BEG[0]
+ Tile_X9Y9_LUT4AB/W6BEG[10] Tile_X9Y9_LUT4AB/W6BEG[11] Tile_X9Y9_LUT4AB/W6BEG[1]
+ Tile_X9Y9_LUT4AB/W6BEG[2] Tile_X9Y9_LUT4AB/W6BEG[3] Tile_X9Y9_LUT4AB/W6BEG[4] Tile_X9Y9_LUT4AB/W6BEG[5]
+ Tile_X9Y9_LUT4AB/W6BEG[6] Tile_X9Y9_LUT4AB/W6BEG[7] Tile_X9Y9_LUT4AB/W6BEG[8] Tile_X9Y9_LUT4AB/W6BEG[9]
+ Tile_X9Y9_LUT4AB/W6END[0] Tile_X9Y9_LUT4AB/W6END[10] Tile_X9Y9_LUT4AB/W6END[11]
+ Tile_X9Y9_LUT4AB/W6END[1] Tile_X9Y9_LUT4AB/W6END[2] Tile_X9Y9_LUT4AB/W6END[3] Tile_X9Y9_LUT4AB/W6END[4]
+ Tile_X9Y9_LUT4AB/W6END[5] Tile_X9Y9_LUT4AB/W6END[6] Tile_X9Y9_LUT4AB/W6END[7] Tile_X9Y9_LUT4AB/W6END[8]
+ Tile_X9Y9_LUT4AB/W6END[9] Tile_X9Y9_LUT4AB/WW4BEG[0] Tile_X9Y9_LUT4AB/WW4BEG[10]
+ Tile_X9Y9_LUT4AB/WW4BEG[11] Tile_X9Y9_LUT4AB/WW4BEG[12] Tile_X9Y9_LUT4AB/WW4BEG[13]
+ Tile_X9Y9_LUT4AB/WW4BEG[14] Tile_X9Y9_LUT4AB/WW4BEG[15] Tile_X9Y9_LUT4AB/WW4BEG[1]
+ Tile_X9Y9_LUT4AB/WW4BEG[2] Tile_X9Y9_LUT4AB/WW4BEG[3] Tile_X9Y9_LUT4AB/WW4BEG[4]
+ Tile_X9Y9_LUT4AB/WW4BEG[5] Tile_X9Y9_LUT4AB/WW4BEG[6] Tile_X9Y9_LUT4AB/WW4BEG[7]
+ Tile_X9Y9_LUT4AB/WW4BEG[8] Tile_X9Y9_LUT4AB/WW4BEG[9] Tile_X9Y9_LUT4AB/WW4END[0]
+ Tile_X9Y9_LUT4AB/WW4END[10] Tile_X9Y9_LUT4AB/WW4END[11] Tile_X9Y9_LUT4AB/WW4END[12]
+ Tile_X9Y9_LUT4AB/WW4END[13] Tile_X9Y9_LUT4AB/WW4END[14] Tile_X9Y9_LUT4AB/WW4END[15]
+ Tile_X9Y9_LUT4AB/WW4END[1] Tile_X9Y9_LUT4AB/WW4END[2] Tile_X9Y9_LUT4AB/WW4END[3]
+ Tile_X9Y9_LUT4AB/WW4END[4] Tile_X9Y9_LUT4AB/WW4END[5] Tile_X9Y9_LUT4AB/WW4END[6]
+ Tile_X9Y9_LUT4AB/WW4END[7] Tile_X9Y9_LUT4AB/WW4END[8] Tile_X9Y9_LUT4AB/WW4END[9]
+ LUT4AB
XTile_X6Y4_LUT4AB Tile_X6Y5_LUT4AB/Co Tile_X6Y4_LUT4AB/Co Tile_X6Y4_LUT4AB/E1BEG[0]
+ Tile_X6Y4_LUT4AB/E1BEG[1] Tile_X6Y4_LUT4AB/E1BEG[2] Tile_X6Y4_LUT4AB/E1BEG[3] Tile_X6Y4_LUT4AB/E1END[0]
+ Tile_X6Y4_LUT4AB/E1END[1] Tile_X6Y4_LUT4AB/E1END[2] Tile_X6Y4_LUT4AB/E1END[3] Tile_X6Y4_LUT4AB/E2BEG[0]
+ Tile_X6Y4_LUT4AB/E2BEG[1] Tile_X6Y4_LUT4AB/E2BEG[2] Tile_X6Y4_LUT4AB/E2BEG[3] Tile_X6Y4_LUT4AB/E2BEG[4]
+ Tile_X6Y4_LUT4AB/E2BEG[5] Tile_X6Y4_LUT4AB/E2BEG[6] Tile_X6Y4_LUT4AB/E2BEG[7] Tile_X6Y4_LUT4AB/E2BEGb[0]
+ Tile_X6Y4_LUT4AB/E2BEGb[1] Tile_X6Y4_LUT4AB/E2BEGb[2] Tile_X6Y4_LUT4AB/E2BEGb[3]
+ Tile_X6Y4_LUT4AB/E2BEGb[4] Tile_X6Y4_LUT4AB/E2BEGb[5] Tile_X6Y4_LUT4AB/E2BEGb[6]
+ Tile_X6Y4_LUT4AB/E2BEGb[7] Tile_X6Y4_LUT4AB/E2END[0] Tile_X6Y4_LUT4AB/E2END[1] Tile_X6Y4_LUT4AB/E2END[2]
+ Tile_X6Y4_LUT4AB/E2END[3] Tile_X6Y4_LUT4AB/E2END[4] Tile_X6Y4_LUT4AB/E2END[5] Tile_X6Y4_LUT4AB/E2END[6]
+ Tile_X6Y4_LUT4AB/E2END[7] Tile_X6Y4_LUT4AB/E2MID[0] Tile_X6Y4_LUT4AB/E2MID[1] Tile_X6Y4_LUT4AB/E2MID[2]
+ Tile_X6Y4_LUT4AB/E2MID[3] Tile_X6Y4_LUT4AB/E2MID[4] Tile_X6Y4_LUT4AB/E2MID[5] Tile_X6Y4_LUT4AB/E2MID[6]
+ Tile_X6Y4_LUT4AB/E2MID[7] Tile_X6Y4_LUT4AB/E6BEG[0] Tile_X6Y4_LUT4AB/E6BEG[10] Tile_X6Y4_LUT4AB/E6BEG[11]
+ Tile_X6Y4_LUT4AB/E6BEG[1] Tile_X6Y4_LUT4AB/E6BEG[2] Tile_X6Y4_LUT4AB/E6BEG[3] Tile_X6Y4_LUT4AB/E6BEG[4]
+ Tile_X6Y4_LUT4AB/E6BEG[5] Tile_X6Y4_LUT4AB/E6BEG[6] Tile_X6Y4_LUT4AB/E6BEG[7] Tile_X6Y4_LUT4AB/E6BEG[8]
+ Tile_X6Y4_LUT4AB/E6BEG[9] Tile_X6Y4_LUT4AB/E6END[0] Tile_X6Y4_LUT4AB/E6END[10] Tile_X6Y4_LUT4AB/E6END[11]
+ Tile_X6Y4_LUT4AB/E6END[1] Tile_X6Y4_LUT4AB/E6END[2] Tile_X6Y4_LUT4AB/E6END[3] Tile_X6Y4_LUT4AB/E6END[4]
+ Tile_X6Y4_LUT4AB/E6END[5] Tile_X6Y4_LUT4AB/E6END[6] Tile_X6Y4_LUT4AB/E6END[7] Tile_X6Y4_LUT4AB/E6END[8]
+ Tile_X6Y4_LUT4AB/E6END[9] Tile_X6Y4_LUT4AB/EE4BEG[0] Tile_X6Y4_LUT4AB/EE4BEG[10]
+ Tile_X6Y4_LUT4AB/EE4BEG[11] Tile_X6Y4_LUT4AB/EE4BEG[12] Tile_X6Y4_LUT4AB/EE4BEG[13]
+ Tile_X6Y4_LUT4AB/EE4BEG[14] Tile_X6Y4_LUT4AB/EE4BEG[15] Tile_X6Y4_LUT4AB/EE4BEG[1]
+ Tile_X6Y4_LUT4AB/EE4BEG[2] Tile_X6Y4_LUT4AB/EE4BEG[3] Tile_X6Y4_LUT4AB/EE4BEG[4]
+ Tile_X6Y4_LUT4AB/EE4BEG[5] Tile_X6Y4_LUT4AB/EE4BEG[6] Tile_X6Y4_LUT4AB/EE4BEG[7]
+ Tile_X6Y4_LUT4AB/EE4BEG[8] Tile_X6Y4_LUT4AB/EE4BEG[9] Tile_X6Y4_LUT4AB/EE4END[0]
+ Tile_X6Y4_LUT4AB/EE4END[10] Tile_X6Y4_LUT4AB/EE4END[11] Tile_X6Y4_LUT4AB/EE4END[12]
+ Tile_X6Y4_LUT4AB/EE4END[13] Tile_X6Y4_LUT4AB/EE4END[14] Tile_X6Y4_LUT4AB/EE4END[15]
+ Tile_X6Y4_LUT4AB/EE4END[1] Tile_X6Y4_LUT4AB/EE4END[2] Tile_X6Y4_LUT4AB/EE4END[3]
+ Tile_X6Y4_LUT4AB/EE4END[4] Tile_X6Y4_LUT4AB/EE4END[5] Tile_X6Y4_LUT4AB/EE4END[6]
+ Tile_X6Y4_LUT4AB/EE4END[7] Tile_X6Y4_LUT4AB/EE4END[8] Tile_X6Y4_LUT4AB/EE4END[9]
+ Tile_X6Y4_LUT4AB/FrameData[0] Tile_X6Y4_LUT4AB/FrameData[10] Tile_X6Y4_LUT4AB/FrameData[11]
+ Tile_X6Y4_LUT4AB/FrameData[12] Tile_X6Y4_LUT4AB/FrameData[13] Tile_X6Y4_LUT4AB/FrameData[14]
+ Tile_X6Y4_LUT4AB/FrameData[15] Tile_X6Y4_LUT4AB/FrameData[16] Tile_X6Y4_LUT4AB/FrameData[17]
+ Tile_X6Y4_LUT4AB/FrameData[18] Tile_X6Y4_LUT4AB/FrameData[19] Tile_X6Y4_LUT4AB/FrameData[1]
+ Tile_X6Y4_LUT4AB/FrameData[20] Tile_X6Y4_LUT4AB/FrameData[21] Tile_X6Y4_LUT4AB/FrameData[22]
+ Tile_X6Y4_LUT4AB/FrameData[23] Tile_X6Y4_LUT4AB/FrameData[24] Tile_X6Y4_LUT4AB/FrameData[25]
+ Tile_X6Y4_LUT4AB/FrameData[26] Tile_X6Y4_LUT4AB/FrameData[27] Tile_X6Y4_LUT4AB/FrameData[28]
+ Tile_X6Y4_LUT4AB/FrameData[29] Tile_X6Y4_LUT4AB/FrameData[2] Tile_X6Y4_LUT4AB/FrameData[30]
+ Tile_X6Y4_LUT4AB/FrameData[31] Tile_X6Y4_LUT4AB/FrameData[3] Tile_X6Y4_LUT4AB/FrameData[4]
+ Tile_X6Y4_LUT4AB/FrameData[5] Tile_X6Y4_LUT4AB/FrameData[6] Tile_X6Y4_LUT4AB/FrameData[7]
+ Tile_X6Y4_LUT4AB/FrameData[8] Tile_X6Y4_LUT4AB/FrameData[9] Tile_X6Y4_LUT4AB/FrameData_O[0]
+ Tile_X6Y4_LUT4AB/FrameData_O[10] Tile_X6Y4_LUT4AB/FrameData_O[11] Tile_X6Y4_LUT4AB/FrameData_O[12]
+ Tile_X6Y4_LUT4AB/FrameData_O[13] Tile_X6Y4_LUT4AB/FrameData_O[14] Tile_X6Y4_LUT4AB/FrameData_O[15]
+ Tile_X6Y4_LUT4AB/FrameData_O[16] Tile_X6Y4_LUT4AB/FrameData_O[17] Tile_X6Y4_LUT4AB/FrameData_O[18]
+ Tile_X6Y4_LUT4AB/FrameData_O[19] Tile_X6Y4_LUT4AB/FrameData_O[1] Tile_X6Y4_LUT4AB/FrameData_O[20]
+ Tile_X6Y4_LUT4AB/FrameData_O[21] Tile_X6Y4_LUT4AB/FrameData_O[22] Tile_X6Y4_LUT4AB/FrameData_O[23]
+ Tile_X6Y4_LUT4AB/FrameData_O[24] Tile_X6Y4_LUT4AB/FrameData_O[25] Tile_X6Y4_LUT4AB/FrameData_O[26]
+ Tile_X6Y4_LUT4AB/FrameData_O[27] Tile_X6Y4_LUT4AB/FrameData_O[28] Tile_X6Y4_LUT4AB/FrameData_O[29]
+ Tile_X6Y4_LUT4AB/FrameData_O[2] Tile_X6Y4_LUT4AB/FrameData_O[30] Tile_X6Y4_LUT4AB/FrameData_O[31]
+ Tile_X6Y4_LUT4AB/FrameData_O[3] Tile_X6Y4_LUT4AB/FrameData_O[4] Tile_X6Y4_LUT4AB/FrameData_O[5]
+ Tile_X6Y4_LUT4AB/FrameData_O[6] Tile_X6Y4_LUT4AB/FrameData_O[7] Tile_X6Y4_LUT4AB/FrameData_O[8]
+ Tile_X6Y4_LUT4AB/FrameData_O[9] Tile_X6Y4_LUT4AB/FrameStrobe[0] Tile_X6Y4_LUT4AB/FrameStrobe[10]
+ Tile_X6Y4_LUT4AB/FrameStrobe[11] Tile_X6Y4_LUT4AB/FrameStrobe[12] Tile_X6Y4_LUT4AB/FrameStrobe[13]
+ Tile_X6Y4_LUT4AB/FrameStrobe[14] Tile_X6Y4_LUT4AB/FrameStrobe[15] Tile_X6Y4_LUT4AB/FrameStrobe[16]
+ Tile_X6Y4_LUT4AB/FrameStrobe[17] Tile_X6Y4_LUT4AB/FrameStrobe[18] Tile_X6Y4_LUT4AB/FrameStrobe[19]
+ Tile_X6Y4_LUT4AB/FrameStrobe[1] Tile_X6Y4_LUT4AB/FrameStrobe[2] Tile_X6Y4_LUT4AB/FrameStrobe[3]
+ Tile_X6Y4_LUT4AB/FrameStrobe[4] Tile_X6Y4_LUT4AB/FrameStrobe[5] Tile_X6Y4_LUT4AB/FrameStrobe[6]
+ Tile_X6Y4_LUT4AB/FrameStrobe[7] Tile_X6Y4_LUT4AB/FrameStrobe[8] Tile_X6Y4_LUT4AB/FrameStrobe[9]
+ Tile_X6Y3_LUT4AB/FrameStrobe[0] Tile_X6Y3_LUT4AB/FrameStrobe[10] Tile_X6Y3_LUT4AB/FrameStrobe[11]
+ Tile_X6Y3_LUT4AB/FrameStrobe[12] Tile_X6Y3_LUT4AB/FrameStrobe[13] Tile_X6Y3_LUT4AB/FrameStrobe[14]
+ Tile_X6Y3_LUT4AB/FrameStrobe[15] Tile_X6Y3_LUT4AB/FrameStrobe[16] Tile_X6Y3_LUT4AB/FrameStrobe[17]
+ Tile_X6Y3_LUT4AB/FrameStrobe[18] Tile_X6Y3_LUT4AB/FrameStrobe[19] Tile_X6Y3_LUT4AB/FrameStrobe[1]
+ Tile_X6Y3_LUT4AB/FrameStrobe[2] Tile_X6Y3_LUT4AB/FrameStrobe[3] Tile_X6Y3_LUT4AB/FrameStrobe[4]
+ Tile_X6Y3_LUT4AB/FrameStrobe[5] Tile_X6Y3_LUT4AB/FrameStrobe[6] Tile_X6Y3_LUT4AB/FrameStrobe[7]
+ Tile_X6Y3_LUT4AB/FrameStrobe[8] Tile_X6Y3_LUT4AB/FrameStrobe[9] Tile_X6Y4_LUT4AB/N1BEG[0]
+ Tile_X6Y4_LUT4AB/N1BEG[1] Tile_X6Y4_LUT4AB/N1BEG[2] Tile_X6Y4_LUT4AB/N1BEG[3] Tile_X6Y5_LUT4AB/N1BEG[0]
+ Tile_X6Y5_LUT4AB/N1BEG[1] Tile_X6Y5_LUT4AB/N1BEG[2] Tile_X6Y5_LUT4AB/N1BEG[3] Tile_X6Y4_LUT4AB/N2BEG[0]
+ Tile_X6Y4_LUT4AB/N2BEG[1] Tile_X6Y4_LUT4AB/N2BEG[2] Tile_X6Y4_LUT4AB/N2BEG[3] Tile_X6Y4_LUT4AB/N2BEG[4]
+ Tile_X6Y4_LUT4AB/N2BEG[5] Tile_X6Y4_LUT4AB/N2BEG[6] Tile_X6Y4_LUT4AB/N2BEG[7] Tile_X6Y3_LUT4AB/N2END[0]
+ Tile_X6Y3_LUT4AB/N2END[1] Tile_X6Y3_LUT4AB/N2END[2] Tile_X6Y3_LUT4AB/N2END[3] Tile_X6Y3_LUT4AB/N2END[4]
+ Tile_X6Y3_LUT4AB/N2END[5] Tile_X6Y3_LUT4AB/N2END[6] Tile_X6Y3_LUT4AB/N2END[7] Tile_X6Y4_LUT4AB/N2END[0]
+ Tile_X6Y4_LUT4AB/N2END[1] Tile_X6Y4_LUT4AB/N2END[2] Tile_X6Y4_LUT4AB/N2END[3] Tile_X6Y4_LUT4AB/N2END[4]
+ Tile_X6Y4_LUT4AB/N2END[5] Tile_X6Y4_LUT4AB/N2END[6] Tile_X6Y4_LUT4AB/N2END[7] Tile_X6Y5_LUT4AB/N2BEG[0]
+ Tile_X6Y5_LUT4AB/N2BEG[1] Tile_X6Y5_LUT4AB/N2BEG[2] Tile_X6Y5_LUT4AB/N2BEG[3] Tile_X6Y5_LUT4AB/N2BEG[4]
+ Tile_X6Y5_LUT4AB/N2BEG[5] Tile_X6Y5_LUT4AB/N2BEG[6] Tile_X6Y5_LUT4AB/N2BEG[7] Tile_X6Y4_LUT4AB/N4BEG[0]
+ Tile_X6Y4_LUT4AB/N4BEG[10] Tile_X6Y4_LUT4AB/N4BEG[11] Tile_X6Y4_LUT4AB/N4BEG[12]
+ Tile_X6Y4_LUT4AB/N4BEG[13] Tile_X6Y4_LUT4AB/N4BEG[14] Tile_X6Y4_LUT4AB/N4BEG[15]
+ Tile_X6Y4_LUT4AB/N4BEG[1] Tile_X6Y4_LUT4AB/N4BEG[2] Tile_X6Y4_LUT4AB/N4BEG[3] Tile_X6Y4_LUT4AB/N4BEG[4]
+ Tile_X6Y4_LUT4AB/N4BEG[5] Tile_X6Y4_LUT4AB/N4BEG[6] Tile_X6Y4_LUT4AB/N4BEG[7] Tile_X6Y4_LUT4AB/N4BEG[8]
+ Tile_X6Y4_LUT4AB/N4BEG[9] Tile_X6Y5_LUT4AB/N4BEG[0] Tile_X6Y5_LUT4AB/N4BEG[10] Tile_X6Y5_LUT4AB/N4BEG[11]
+ Tile_X6Y5_LUT4AB/N4BEG[12] Tile_X6Y5_LUT4AB/N4BEG[13] Tile_X6Y5_LUT4AB/N4BEG[14]
+ Tile_X6Y5_LUT4AB/N4BEG[15] Tile_X6Y5_LUT4AB/N4BEG[1] Tile_X6Y5_LUT4AB/N4BEG[2] Tile_X6Y5_LUT4AB/N4BEG[3]
+ Tile_X6Y5_LUT4AB/N4BEG[4] Tile_X6Y5_LUT4AB/N4BEG[5] Tile_X6Y5_LUT4AB/N4BEG[6] Tile_X6Y5_LUT4AB/N4BEG[7]
+ Tile_X6Y5_LUT4AB/N4BEG[8] Tile_X6Y5_LUT4AB/N4BEG[9] Tile_X6Y4_LUT4AB/NN4BEG[0] Tile_X6Y4_LUT4AB/NN4BEG[10]
+ Tile_X6Y4_LUT4AB/NN4BEG[11] Tile_X6Y4_LUT4AB/NN4BEG[12] Tile_X6Y4_LUT4AB/NN4BEG[13]
+ Tile_X6Y4_LUT4AB/NN4BEG[14] Tile_X6Y4_LUT4AB/NN4BEG[15] Tile_X6Y4_LUT4AB/NN4BEG[1]
+ Tile_X6Y4_LUT4AB/NN4BEG[2] Tile_X6Y4_LUT4AB/NN4BEG[3] Tile_X6Y4_LUT4AB/NN4BEG[4]
+ Tile_X6Y4_LUT4AB/NN4BEG[5] Tile_X6Y4_LUT4AB/NN4BEG[6] Tile_X6Y4_LUT4AB/NN4BEG[7]
+ Tile_X6Y4_LUT4AB/NN4BEG[8] Tile_X6Y4_LUT4AB/NN4BEG[9] Tile_X6Y5_LUT4AB/NN4BEG[0]
+ Tile_X6Y5_LUT4AB/NN4BEG[10] Tile_X6Y5_LUT4AB/NN4BEG[11] Tile_X6Y5_LUT4AB/NN4BEG[12]
+ Tile_X6Y5_LUT4AB/NN4BEG[13] Tile_X6Y5_LUT4AB/NN4BEG[14] Tile_X6Y5_LUT4AB/NN4BEG[15]
+ Tile_X6Y5_LUT4AB/NN4BEG[1] Tile_X6Y5_LUT4AB/NN4BEG[2] Tile_X6Y5_LUT4AB/NN4BEG[3]
+ Tile_X6Y5_LUT4AB/NN4BEG[4] Tile_X6Y5_LUT4AB/NN4BEG[5] Tile_X6Y5_LUT4AB/NN4BEG[6]
+ Tile_X6Y5_LUT4AB/NN4BEG[7] Tile_X6Y5_LUT4AB/NN4BEG[8] Tile_X6Y5_LUT4AB/NN4BEG[9]
+ Tile_X6Y5_LUT4AB/S1END[0] Tile_X6Y5_LUT4AB/S1END[1] Tile_X6Y5_LUT4AB/S1END[2] Tile_X6Y5_LUT4AB/S1END[3]
+ Tile_X6Y4_LUT4AB/S1END[0] Tile_X6Y4_LUT4AB/S1END[1] Tile_X6Y4_LUT4AB/S1END[2] Tile_X6Y4_LUT4AB/S1END[3]
+ Tile_X6Y5_LUT4AB/S2MID[0] Tile_X6Y5_LUT4AB/S2MID[1] Tile_X6Y5_LUT4AB/S2MID[2] Tile_X6Y5_LUT4AB/S2MID[3]
+ Tile_X6Y5_LUT4AB/S2MID[4] Tile_X6Y5_LUT4AB/S2MID[5] Tile_X6Y5_LUT4AB/S2MID[6] Tile_X6Y5_LUT4AB/S2MID[7]
+ Tile_X6Y5_LUT4AB/S2END[0] Tile_X6Y5_LUT4AB/S2END[1] Tile_X6Y5_LUT4AB/S2END[2] Tile_X6Y5_LUT4AB/S2END[3]
+ Tile_X6Y5_LUT4AB/S2END[4] Tile_X6Y5_LUT4AB/S2END[5] Tile_X6Y5_LUT4AB/S2END[6] Tile_X6Y5_LUT4AB/S2END[7]
+ Tile_X6Y4_LUT4AB/S2END[0] Tile_X6Y4_LUT4AB/S2END[1] Tile_X6Y4_LUT4AB/S2END[2] Tile_X6Y4_LUT4AB/S2END[3]
+ Tile_X6Y4_LUT4AB/S2END[4] Tile_X6Y4_LUT4AB/S2END[5] Tile_X6Y4_LUT4AB/S2END[6] Tile_X6Y4_LUT4AB/S2END[7]
+ Tile_X6Y4_LUT4AB/S2MID[0] Tile_X6Y4_LUT4AB/S2MID[1] Tile_X6Y4_LUT4AB/S2MID[2] Tile_X6Y4_LUT4AB/S2MID[3]
+ Tile_X6Y4_LUT4AB/S2MID[4] Tile_X6Y4_LUT4AB/S2MID[5] Tile_X6Y4_LUT4AB/S2MID[6] Tile_X6Y4_LUT4AB/S2MID[7]
+ Tile_X6Y5_LUT4AB/S4END[0] Tile_X6Y5_LUT4AB/S4END[10] Tile_X6Y5_LUT4AB/S4END[11]
+ Tile_X6Y5_LUT4AB/S4END[12] Tile_X6Y5_LUT4AB/S4END[13] Tile_X6Y5_LUT4AB/S4END[14]
+ Tile_X6Y5_LUT4AB/S4END[15] Tile_X6Y5_LUT4AB/S4END[1] Tile_X6Y5_LUT4AB/S4END[2] Tile_X6Y5_LUT4AB/S4END[3]
+ Tile_X6Y5_LUT4AB/S4END[4] Tile_X6Y5_LUT4AB/S4END[5] Tile_X6Y5_LUT4AB/S4END[6] Tile_X6Y5_LUT4AB/S4END[7]
+ Tile_X6Y5_LUT4AB/S4END[8] Tile_X6Y5_LUT4AB/S4END[9] Tile_X6Y4_LUT4AB/S4END[0] Tile_X6Y4_LUT4AB/S4END[10]
+ Tile_X6Y4_LUT4AB/S4END[11] Tile_X6Y4_LUT4AB/S4END[12] Tile_X6Y4_LUT4AB/S4END[13]
+ Tile_X6Y4_LUT4AB/S4END[14] Tile_X6Y4_LUT4AB/S4END[15] Tile_X6Y4_LUT4AB/S4END[1]
+ Tile_X6Y4_LUT4AB/S4END[2] Tile_X6Y4_LUT4AB/S4END[3] Tile_X6Y4_LUT4AB/S4END[4] Tile_X6Y4_LUT4AB/S4END[5]
+ Tile_X6Y4_LUT4AB/S4END[6] Tile_X6Y4_LUT4AB/S4END[7] Tile_X6Y4_LUT4AB/S4END[8] Tile_X6Y4_LUT4AB/S4END[9]
+ Tile_X6Y5_LUT4AB/SS4END[0] Tile_X6Y5_LUT4AB/SS4END[10] Tile_X6Y5_LUT4AB/SS4END[11]
+ Tile_X6Y5_LUT4AB/SS4END[12] Tile_X6Y5_LUT4AB/SS4END[13] Tile_X6Y5_LUT4AB/SS4END[14]
+ Tile_X6Y5_LUT4AB/SS4END[15] Tile_X6Y5_LUT4AB/SS4END[1] Tile_X6Y5_LUT4AB/SS4END[2]
+ Tile_X6Y5_LUT4AB/SS4END[3] Tile_X6Y5_LUT4AB/SS4END[4] Tile_X6Y5_LUT4AB/SS4END[5]
+ Tile_X6Y5_LUT4AB/SS4END[6] Tile_X6Y5_LUT4AB/SS4END[7] Tile_X6Y5_LUT4AB/SS4END[8]
+ Tile_X6Y5_LUT4AB/SS4END[9] Tile_X6Y4_LUT4AB/SS4END[0] Tile_X6Y4_LUT4AB/SS4END[10]
+ Tile_X6Y4_LUT4AB/SS4END[11] Tile_X6Y4_LUT4AB/SS4END[12] Tile_X6Y4_LUT4AB/SS4END[13]
+ Tile_X6Y4_LUT4AB/SS4END[14] Tile_X6Y4_LUT4AB/SS4END[15] Tile_X6Y4_LUT4AB/SS4END[1]
+ Tile_X6Y4_LUT4AB/SS4END[2] Tile_X6Y4_LUT4AB/SS4END[3] Tile_X6Y4_LUT4AB/SS4END[4]
+ Tile_X6Y4_LUT4AB/SS4END[5] Tile_X6Y4_LUT4AB/SS4END[6] Tile_X6Y4_LUT4AB/SS4END[7]
+ Tile_X6Y4_LUT4AB/SS4END[8] Tile_X6Y4_LUT4AB/SS4END[9] Tile_X6Y4_LUT4AB/UserCLK Tile_X6Y3_LUT4AB/UserCLK
+ VGND VPWR Tile_X6Y4_LUT4AB/W1BEG[0] Tile_X6Y4_LUT4AB/W1BEG[1] Tile_X6Y4_LUT4AB/W1BEG[2]
+ Tile_X6Y4_LUT4AB/W1BEG[3] Tile_X6Y4_LUT4AB/W1END[0] Tile_X6Y4_LUT4AB/W1END[1] Tile_X6Y4_LUT4AB/W1END[2]
+ Tile_X6Y4_LUT4AB/W1END[3] Tile_X6Y4_LUT4AB/W2BEG[0] Tile_X6Y4_LUT4AB/W2BEG[1] Tile_X6Y4_LUT4AB/W2BEG[2]
+ Tile_X6Y4_LUT4AB/W2BEG[3] Tile_X6Y4_LUT4AB/W2BEG[4] Tile_X6Y4_LUT4AB/W2BEG[5] Tile_X6Y4_LUT4AB/W2BEG[6]
+ Tile_X6Y4_LUT4AB/W2BEG[7] Tile_X5Y4_LUT4AB/W2END[0] Tile_X5Y4_LUT4AB/W2END[1] Tile_X5Y4_LUT4AB/W2END[2]
+ Tile_X5Y4_LUT4AB/W2END[3] Tile_X5Y4_LUT4AB/W2END[4] Tile_X5Y4_LUT4AB/W2END[5] Tile_X5Y4_LUT4AB/W2END[6]
+ Tile_X5Y4_LUT4AB/W2END[7] Tile_X6Y4_LUT4AB/W2END[0] Tile_X6Y4_LUT4AB/W2END[1] Tile_X6Y4_LUT4AB/W2END[2]
+ Tile_X6Y4_LUT4AB/W2END[3] Tile_X6Y4_LUT4AB/W2END[4] Tile_X6Y4_LUT4AB/W2END[5] Tile_X6Y4_LUT4AB/W2END[6]
+ Tile_X6Y4_LUT4AB/W2END[7] Tile_X6Y4_LUT4AB/W2MID[0] Tile_X6Y4_LUT4AB/W2MID[1] Tile_X6Y4_LUT4AB/W2MID[2]
+ Tile_X6Y4_LUT4AB/W2MID[3] Tile_X6Y4_LUT4AB/W2MID[4] Tile_X6Y4_LUT4AB/W2MID[5] Tile_X6Y4_LUT4AB/W2MID[6]
+ Tile_X6Y4_LUT4AB/W2MID[7] Tile_X6Y4_LUT4AB/W6BEG[0] Tile_X6Y4_LUT4AB/W6BEG[10] Tile_X6Y4_LUT4AB/W6BEG[11]
+ Tile_X6Y4_LUT4AB/W6BEG[1] Tile_X6Y4_LUT4AB/W6BEG[2] Tile_X6Y4_LUT4AB/W6BEG[3] Tile_X6Y4_LUT4AB/W6BEG[4]
+ Tile_X6Y4_LUT4AB/W6BEG[5] Tile_X6Y4_LUT4AB/W6BEG[6] Tile_X6Y4_LUT4AB/W6BEG[7] Tile_X6Y4_LUT4AB/W6BEG[8]
+ Tile_X6Y4_LUT4AB/W6BEG[9] Tile_X6Y4_LUT4AB/W6END[0] Tile_X6Y4_LUT4AB/W6END[10] Tile_X6Y4_LUT4AB/W6END[11]
+ Tile_X6Y4_LUT4AB/W6END[1] Tile_X6Y4_LUT4AB/W6END[2] Tile_X6Y4_LUT4AB/W6END[3] Tile_X6Y4_LUT4AB/W6END[4]
+ Tile_X6Y4_LUT4AB/W6END[5] Tile_X6Y4_LUT4AB/W6END[6] Tile_X6Y4_LUT4AB/W6END[7] Tile_X6Y4_LUT4AB/W6END[8]
+ Tile_X6Y4_LUT4AB/W6END[9] Tile_X6Y4_LUT4AB/WW4BEG[0] Tile_X6Y4_LUT4AB/WW4BEG[10]
+ Tile_X6Y4_LUT4AB/WW4BEG[11] Tile_X6Y4_LUT4AB/WW4BEG[12] Tile_X6Y4_LUT4AB/WW4BEG[13]
+ Tile_X6Y4_LUT4AB/WW4BEG[14] Tile_X6Y4_LUT4AB/WW4BEG[15] Tile_X6Y4_LUT4AB/WW4BEG[1]
+ Tile_X6Y4_LUT4AB/WW4BEG[2] Tile_X6Y4_LUT4AB/WW4BEG[3] Tile_X6Y4_LUT4AB/WW4BEG[4]
+ Tile_X6Y4_LUT4AB/WW4BEG[5] Tile_X6Y4_LUT4AB/WW4BEG[6] Tile_X6Y4_LUT4AB/WW4BEG[7]
+ Tile_X6Y4_LUT4AB/WW4BEG[8] Tile_X6Y4_LUT4AB/WW4BEG[9] Tile_X6Y4_LUT4AB/WW4END[0]
+ Tile_X6Y4_LUT4AB/WW4END[10] Tile_X6Y4_LUT4AB/WW4END[11] Tile_X6Y4_LUT4AB/WW4END[12]
+ Tile_X6Y4_LUT4AB/WW4END[13] Tile_X6Y4_LUT4AB/WW4END[14] Tile_X6Y4_LUT4AB/WW4END[15]
+ Tile_X6Y4_LUT4AB/WW4END[1] Tile_X6Y4_LUT4AB/WW4END[2] Tile_X6Y4_LUT4AB/WW4END[3]
+ Tile_X6Y4_LUT4AB/WW4END[4] Tile_X6Y4_LUT4AB/WW4END[5] Tile_X6Y4_LUT4AB/WW4END[6]
+ Tile_X6Y4_LUT4AB/WW4END[7] Tile_X6Y4_LUT4AB/WW4END[8] Tile_X6Y4_LUT4AB/WW4END[9]
+ LUT4AB
XTile_X0Y13_W_IO Tile_X0Y13_A_I_top Tile_X0Y13_A_O_top Tile_X0Y13_A_T_top Tile_X0Y13_A_config_C_bit0
+ Tile_X0Y13_A_config_C_bit1 Tile_X0Y13_A_config_C_bit2 Tile_X0Y13_A_config_C_bit3
+ Tile_X0Y13_B_I_top Tile_X0Y13_B_O_top Tile_X0Y13_B_T_top Tile_X0Y13_B_config_C_bit0
+ Tile_X0Y13_B_config_C_bit1 Tile_X0Y13_B_config_C_bit2 Tile_X0Y13_B_config_C_bit3
+ Tile_X0Y13_W_IO/E1BEG[0] Tile_X0Y13_W_IO/E1BEG[1] Tile_X0Y13_W_IO/E1BEG[2] Tile_X0Y13_W_IO/E1BEG[3]
+ Tile_X0Y13_W_IO/E2BEG[0] Tile_X0Y13_W_IO/E2BEG[1] Tile_X0Y13_W_IO/E2BEG[2] Tile_X0Y13_W_IO/E2BEG[3]
+ Tile_X0Y13_W_IO/E2BEG[4] Tile_X0Y13_W_IO/E2BEG[5] Tile_X0Y13_W_IO/E2BEG[6] Tile_X0Y13_W_IO/E2BEG[7]
+ Tile_X0Y13_W_IO/E2BEGb[0] Tile_X0Y13_W_IO/E2BEGb[1] Tile_X0Y13_W_IO/E2BEGb[2] Tile_X0Y13_W_IO/E2BEGb[3]
+ Tile_X0Y13_W_IO/E2BEGb[4] Tile_X0Y13_W_IO/E2BEGb[5] Tile_X0Y13_W_IO/E2BEGb[6] Tile_X0Y13_W_IO/E2BEGb[7]
+ Tile_X0Y13_W_IO/E6BEG[0] Tile_X0Y13_W_IO/E6BEG[10] Tile_X0Y13_W_IO/E6BEG[11] Tile_X0Y13_W_IO/E6BEG[1]
+ Tile_X0Y13_W_IO/E6BEG[2] Tile_X0Y13_W_IO/E6BEG[3] Tile_X0Y13_W_IO/E6BEG[4] Tile_X0Y13_W_IO/E6BEG[5]
+ Tile_X0Y13_W_IO/E6BEG[6] Tile_X0Y13_W_IO/E6BEG[7] Tile_X0Y13_W_IO/E6BEG[8] Tile_X0Y13_W_IO/E6BEG[9]
+ Tile_X0Y13_W_IO/EE4BEG[0] Tile_X0Y13_W_IO/EE4BEG[10] Tile_X0Y13_W_IO/EE4BEG[11]
+ Tile_X0Y13_W_IO/EE4BEG[12] Tile_X0Y13_W_IO/EE4BEG[13] Tile_X0Y13_W_IO/EE4BEG[14]
+ Tile_X0Y13_W_IO/EE4BEG[15] Tile_X0Y13_W_IO/EE4BEG[1] Tile_X0Y13_W_IO/EE4BEG[2] Tile_X0Y13_W_IO/EE4BEG[3]
+ Tile_X0Y13_W_IO/EE4BEG[4] Tile_X0Y13_W_IO/EE4BEG[5] Tile_X0Y13_W_IO/EE4BEG[6] Tile_X0Y13_W_IO/EE4BEG[7]
+ Tile_X0Y13_W_IO/EE4BEG[8] Tile_X0Y13_W_IO/EE4BEG[9] FrameData[416] FrameData[426]
+ FrameData[427] FrameData[428] FrameData[429] FrameData[430] FrameData[431] FrameData[432]
+ FrameData[433] FrameData[434] FrameData[435] FrameData[417] FrameData[436] FrameData[437]
+ FrameData[438] FrameData[439] FrameData[440] FrameData[441] FrameData[442] FrameData[443]
+ FrameData[444] FrameData[445] FrameData[418] FrameData[446] FrameData[447] FrameData[419]
+ FrameData[420] FrameData[421] FrameData[422] FrameData[423] FrameData[424] FrameData[425]
+ Tile_X1Y13_LUT4AB/FrameData[0] Tile_X1Y13_LUT4AB/FrameData[10] Tile_X1Y13_LUT4AB/FrameData[11]
+ Tile_X1Y13_LUT4AB/FrameData[12] Tile_X1Y13_LUT4AB/FrameData[13] Tile_X1Y13_LUT4AB/FrameData[14]
+ Tile_X1Y13_LUT4AB/FrameData[15] Tile_X1Y13_LUT4AB/FrameData[16] Tile_X1Y13_LUT4AB/FrameData[17]
+ Tile_X1Y13_LUT4AB/FrameData[18] Tile_X1Y13_LUT4AB/FrameData[19] Tile_X1Y13_LUT4AB/FrameData[1]
+ Tile_X1Y13_LUT4AB/FrameData[20] Tile_X1Y13_LUT4AB/FrameData[21] Tile_X1Y13_LUT4AB/FrameData[22]
+ Tile_X1Y13_LUT4AB/FrameData[23] Tile_X1Y13_LUT4AB/FrameData[24] Tile_X1Y13_LUT4AB/FrameData[25]
+ Tile_X1Y13_LUT4AB/FrameData[26] Tile_X1Y13_LUT4AB/FrameData[27] Tile_X1Y13_LUT4AB/FrameData[28]
+ Tile_X1Y13_LUT4AB/FrameData[29] Tile_X1Y13_LUT4AB/FrameData[2] Tile_X1Y13_LUT4AB/FrameData[30]
+ Tile_X1Y13_LUT4AB/FrameData[31] Tile_X1Y13_LUT4AB/FrameData[3] Tile_X1Y13_LUT4AB/FrameData[4]
+ Tile_X1Y13_LUT4AB/FrameData[5] Tile_X1Y13_LUT4AB/FrameData[6] Tile_X1Y13_LUT4AB/FrameData[7]
+ Tile_X1Y13_LUT4AB/FrameData[8] Tile_X1Y13_LUT4AB/FrameData[9] Tile_X0Y13_W_IO/FrameStrobe[0]
+ Tile_X0Y13_W_IO/FrameStrobe[10] Tile_X0Y13_W_IO/FrameStrobe[11] Tile_X0Y13_W_IO/FrameStrobe[12]
+ Tile_X0Y13_W_IO/FrameStrobe[13] Tile_X0Y13_W_IO/FrameStrobe[14] Tile_X0Y13_W_IO/FrameStrobe[15]
+ Tile_X0Y13_W_IO/FrameStrobe[16] Tile_X0Y13_W_IO/FrameStrobe[17] Tile_X0Y13_W_IO/FrameStrobe[18]
+ Tile_X0Y13_W_IO/FrameStrobe[19] Tile_X0Y13_W_IO/FrameStrobe[1] Tile_X0Y13_W_IO/FrameStrobe[2]
+ Tile_X0Y13_W_IO/FrameStrobe[3] Tile_X0Y13_W_IO/FrameStrobe[4] Tile_X0Y13_W_IO/FrameStrobe[5]
+ Tile_X0Y13_W_IO/FrameStrobe[6] Tile_X0Y13_W_IO/FrameStrobe[7] Tile_X0Y13_W_IO/FrameStrobe[8]
+ Tile_X0Y13_W_IO/FrameStrobe[9] Tile_X0Y12_W_IO/FrameStrobe[0] Tile_X0Y12_W_IO/FrameStrobe[10]
+ Tile_X0Y12_W_IO/FrameStrobe[11] Tile_X0Y12_W_IO/FrameStrobe[12] Tile_X0Y12_W_IO/FrameStrobe[13]
+ Tile_X0Y12_W_IO/FrameStrobe[14] Tile_X0Y12_W_IO/FrameStrobe[15] Tile_X0Y12_W_IO/FrameStrobe[16]
+ Tile_X0Y12_W_IO/FrameStrobe[17] Tile_X0Y12_W_IO/FrameStrobe[18] Tile_X0Y12_W_IO/FrameStrobe[19]
+ Tile_X0Y12_W_IO/FrameStrobe[1] Tile_X0Y12_W_IO/FrameStrobe[2] Tile_X0Y12_W_IO/FrameStrobe[3]
+ Tile_X0Y12_W_IO/FrameStrobe[4] Tile_X0Y12_W_IO/FrameStrobe[5] Tile_X0Y12_W_IO/FrameStrobe[6]
+ Tile_X0Y12_W_IO/FrameStrobe[7] Tile_X0Y12_W_IO/FrameStrobe[8] Tile_X0Y12_W_IO/FrameStrobe[9]
+ Tile_X0Y13_W_IO/UserCLK Tile_X0Y12_W_IO/UserCLK VGND VPWR Tile_X0Y13_W_IO/W1END[0]
+ Tile_X0Y13_W_IO/W1END[1] Tile_X0Y13_W_IO/W1END[2] Tile_X0Y13_W_IO/W1END[3] Tile_X0Y13_W_IO/W2END[0]
+ Tile_X0Y13_W_IO/W2END[1] Tile_X0Y13_W_IO/W2END[2] Tile_X0Y13_W_IO/W2END[3] Tile_X0Y13_W_IO/W2END[4]
+ Tile_X0Y13_W_IO/W2END[5] Tile_X0Y13_W_IO/W2END[6] Tile_X0Y13_W_IO/W2END[7] Tile_X0Y13_W_IO/W2MID[0]
+ Tile_X0Y13_W_IO/W2MID[1] Tile_X0Y13_W_IO/W2MID[2] Tile_X0Y13_W_IO/W2MID[3] Tile_X0Y13_W_IO/W2MID[4]
+ Tile_X0Y13_W_IO/W2MID[5] Tile_X0Y13_W_IO/W2MID[6] Tile_X0Y13_W_IO/W2MID[7] Tile_X0Y13_W_IO/W6END[0]
+ Tile_X0Y13_W_IO/W6END[10] Tile_X0Y13_W_IO/W6END[11] Tile_X0Y13_W_IO/W6END[1] Tile_X0Y13_W_IO/W6END[2]
+ Tile_X0Y13_W_IO/W6END[3] Tile_X0Y13_W_IO/W6END[4] Tile_X0Y13_W_IO/W6END[5] Tile_X0Y13_W_IO/W6END[6]
+ Tile_X0Y13_W_IO/W6END[7] Tile_X0Y13_W_IO/W6END[8] Tile_X0Y13_W_IO/W6END[9] Tile_X0Y13_W_IO/WW4END[0]
+ Tile_X0Y13_W_IO/WW4END[10] Tile_X0Y13_W_IO/WW4END[11] Tile_X0Y13_W_IO/WW4END[12]
+ Tile_X0Y13_W_IO/WW4END[13] Tile_X0Y13_W_IO/WW4END[14] Tile_X0Y13_W_IO/WW4END[15]
+ Tile_X0Y13_W_IO/WW4END[1] Tile_X0Y13_W_IO/WW4END[2] Tile_X0Y13_W_IO/WW4END[3] Tile_X0Y13_W_IO/WW4END[4]
+ Tile_X0Y13_W_IO/WW4END[5] Tile_X0Y13_W_IO/WW4END[6] Tile_X0Y13_W_IO/WW4END[7] Tile_X0Y13_W_IO/WW4END[8]
+ Tile_X0Y13_W_IO/WW4END[9] W_IO
XTile_X8Y13_LUT4AB Tile_X8Y14_LUT4AB/Co Tile_X8Y13_LUT4AB/Co Tile_X9Y13_LUT4AB/E1END[0]
+ Tile_X9Y13_LUT4AB/E1END[1] Tile_X9Y13_LUT4AB/E1END[2] Tile_X9Y13_LUT4AB/E1END[3]
+ Tile_X8Y13_LUT4AB/E1END[0] Tile_X8Y13_LUT4AB/E1END[1] Tile_X8Y13_LUT4AB/E1END[2]
+ Tile_X8Y13_LUT4AB/E1END[3] Tile_X9Y13_LUT4AB/E2MID[0] Tile_X9Y13_LUT4AB/E2MID[1]
+ Tile_X9Y13_LUT4AB/E2MID[2] Tile_X9Y13_LUT4AB/E2MID[3] Tile_X9Y13_LUT4AB/E2MID[4]
+ Tile_X9Y13_LUT4AB/E2MID[5] Tile_X9Y13_LUT4AB/E2MID[6] Tile_X9Y13_LUT4AB/E2MID[7]
+ Tile_X9Y13_LUT4AB/E2END[0] Tile_X9Y13_LUT4AB/E2END[1] Tile_X9Y13_LUT4AB/E2END[2]
+ Tile_X9Y13_LUT4AB/E2END[3] Tile_X9Y13_LUT4AB/E2END[4] Tile_X9Y13_LUT4AB/E2END[5]
+ Tile_X9Y13_LUT4AB/E2END[6] Tile_X9Y13_LUT4AB/E2END[7] Tile_X8Y13_LUT4AB/E2END[0]
+ Tile_X8Y13_LUT4AB/E2END[1] Tile_X8Y13_LUT4AB/E2END[2] Tile_X8Y13_LUT4AB/E2END[3]
+ Tile_X8Y13_LUT4AB/E2END[4] Tile_X8Y13_LUT4AB/E2END[5] Tile_X8Y13_LUT4AB/E2END[6]
+ Tile_X8Y13_LUT4AB/E2END[7] Tile_X8Y13_LUT4AB/E2MID[0] Tile_X8Y13_LUT4AB/E2MID[1]
+ Tile_X8Y13_LUT4AB/E2MID[2] Tile_X8Y13_LUT4AB/E2MID[3] Tile_X8Y13_LUT4AB/E2MID[4]
+ Tile_X8Y13_LUT4AB/E2MID[5] Tile_X8Y13_LUT4AB/E2MID[6] Tile_X8Y13_LUT4AB/E2MID[7]
+ Tile_X9Y13_LUT4AB/E6END[0] Tile_X9Y13_LUT4AB/E6END[10] Tile_X9Y13_LUT4AB/E6END[11]
+ Tile_X9Y13_LUT4AB/E6END[1] Tile_X9Y13_LUT4AB/E6END[2] Tile_X9Y13_LUT4AB/E6END[3]
+ Tile_X9Y13_LUT4AB/E6END[4] Tile_X9Y13_LUT4AB/E6END[5] Tile_X9Y13_LUT4AB/E6END[6]
+ Tile_X9Y13_LUT4AB/E6END[7] Tile_X9Y13_LUT4AB/E6END[8] Tile_X9Y13_LUT4AB/E6END[9]
+ Tile_X8Y13_LUT4AB/E6END[0] Tile_X8Y13_LUT4AB/E6END[10] Tile_X8Y13_LUT4AB/E6END[11]
+ Tile_X8Y13_LUT4AB/E6END[1] Tile_X8Y13_LUT4AB/E6END[2] Tile_X8Y13_LUT4AB/E6END[3]
+ Tile_X8Y13_LUT4AB/E6END[4] Tile_X8Y13_LUT4AB/E6END[5] Tile_X8Y13_LUT4AB/E6END[6]
+ Tile_X8Y13_LUT4AB/E6END[7] Tile_X8Y13_LUT4AB/E6END[8] Tile_X8Y13_LUT4AB/E6END[9]
+ Tile_X9Y13_LUT4AB/EE4END[0] Tile_X9Y13_LUT4AB/EE4END[10] Tile_X9Y13_LUT4AB/EE4END[11]
+ Tile_X9Y13_LUT4AB/EE4END[12] Tile_X9Y13_LUT4AB/EE4END[13] Tile_X9Y13_LUT4AB/EE4END[14]
+ Tile_X9Y13_LUT4AB/EE4END[15] Tile_X9Y13_LUT4AB/EE4END[1] Tile_X9Y13_LUT4AB/EE4END[2]
+ Tile_X9Y13_LUT4AB/EE4END[3] Tile_X9Y13_LUT4AB/EE4END[4] Tile_X9Y13_LUT4AB/EE4END[5]
+ Tile_X9Y13_LUT4AB/EE4END[6] Tile_X9Y13_LUT4AB/EE4END[7] Tile_X9Y13_LUT4AB/EE4END[8]
+ Tile_X9Y13_LUT4AB/EE4END[9] Tile_X8Y13_LUT4AB/EE4END[0] Tile_X8Y13_LUT4AB/EE4END[10]
+ Tile_X8Y13_LUT4AB/EE4END[11] Tile_X8Y13_LUT4AB/EE4END[12] Tile_X8Y13_LUT4AB/EE4END[13]
+ Tile_X8Y13_LUT4AB/EE4END[14] Tile_X8Y13_LUT4AB/EE4END[15] Tile_X8Y13_LUT4AB/EE4END[1]
+ Tile_X8Y13_LUT4AB/EE4END[2] Tile_X8Y13_LUT4AB/EE4END[3] Tile_X8Y13_LUT4AB/EE4END[4]
+ Tile_X8Y13_LUT4AB/EE4END[5] Tile_X8Y13_LUT4AB/EE4END[6] Tile_X8Y13_LUT4AB/EE4END[7]
+ Tile_X8Y13_LUT4AB/EE4END[8] Tile_X8Y13_LUT4AB/EE4END[9] Tile_X8Y13_LUT4AB/FrameData[0]
+ Tile_X8Y13_LUT4AB/FrameData[10] Tile_X8Y13_LUT4AB/FrameData[11] Tile_X8Y13_LUT4AB/FrameData[12]
+ Tile_X8Y13_LUT4AB/FrameData[13] Tile_X8Y13_LUT4AB/FrameData[14] Tile_X8Y13_LUT4AB/FrameData[15]
+ Tile_X8Y13_LUT4AB/FrameData[16] Tile_X8Y13_LUT4AB/FrameData[17] Tile_X8Y13_LUT4AB/FrameData[18]
+ Tile_X8Y13_LUT4AB/FrameData[19] Tile_X8Y13_LUT4AB/FrameData[1] Tile_X8Y13_LUT4AB/FrameData[20]
+ Tile_X8Y13_LUT4AB/FrameData[21] Tile_X8Y13_LUT4AB/FrameData[22] Tile_X8Y13_LUT4AB/FrameData[23]
+ Tile_X8Y13_LUT4AB/FrameData[24] Tile_X8Y13_LUT4AB/FrameData[25] Tile_X8Y13_LUT4AB/FrameData[26]
+ Tile_X8Y13_LUT4AB/FrameData[27] Tile_X8Y13_LUT4AB/FrameData[28] Tile_X8Y13_LUT4AB/FrameData[29]
+ Tile_X8Y13_LUT4AB/FrameData[2] Tile_X8Y13_LUT4AB/FrameData[30] Tile_X8Y13_LUT4AB/FrameData[31]
+ Tile_X8Y13_LUT4AB/FrameData[3] Tile_X8Y13_LUT4AB/FrameData[4] Tile_X8Y13_LUT4AB/FrameData[5]
+ Tile_X8Y13_LUT4AB/FrameData[6] Tile_X8Y13_LUT4AB/FrameData[7] Tile_X8Y13_LUT4AB/FrameData[8]
+ Tile_X8Y13_LUT4AB/FrameData[9] Tile_X9Y13_LUT4AB/FrameData[0] Tile_X9Y13_LUT4AB/FrameData[10]
+ Tile_X9Y13_LUT4AB/FrameData[11] Tile_X9Y13_LUT4AB/FrameData[12] Tile_X9Y13_LUT4AB/FrameData[13]
+ Tile_X9Y13_LUT4AB/FrameData[14] Tile_X9Y13_LUT4AB/FrameData[15] Tile_X9Y13_LUT4AB/FrameData[16]
+ Tile_X9Y13_LUT4AB/FrameData[17] Tile_X9Y13_LUT4AB/FrameData[18] Tile_X9Y13_LUT4AB/FrameData[19]
+ Tile_X9Y13_LUT4AB/FrameData[1] Tile_X9Y13_LUT4AB/FrameData[20] Tile_X9Y13_LUT4AB/FrameData[21]
+ Tile_X9Y13_LUT4AB/FrameData[22] Tile_X9Y13_LUT4AB/FrameData[23] Tile_X9Y13_LUT4AB/FrameData[24]
+ Tile_X9Y13_LUT4AB/FrameData[25] Tile_X9Y13_LUT4AB/FrameData[26] Tile_X9Y13_LUT4AB/FrameData[27]
+ Tile_X9Y13_LUT4AB/FrameData[28] Tile_X9Y13_LUT4AB/FrameData[29] Tile_X9Y13_LUT4AB/FrameData[2]
+ Tile_X9Y13_LUT4AB/FrameData[30] Tile_X9Y13_LUT4AB/FrameData[31] Tile_X9Y13_LUT4AB/FrameData[3]
+ Tile_X9Y13_LUT4AB/FrameData[4] Tile_X9Y13_LUT4AB/FrameData[5] Tile_X9Y13_LUT4AB/FrameData[6]
+ Tile_X9Y13_LUT4AB/FrameData[7] Tile_X9Y13_LUT4AB/FrameData[8] Tile_X9Y13_LUT4AB/FrameData[9]
+ Tile_X8Y13_LUT4AB/FrameStrobe[0] Tile_X8Y13_LUT4AB/FrameStrobe[10] Tile_X8Y13_LUT4AB/FrameStrobe[11]
+ Tile_X8Y13_LUT4AB/FrameStrobe[12] Tile_X8Y13_LUT4AB/FrameStrobe[13] Tile_X8Y13_LUT4AB/FrameStrobe[14]
+ Tile_X8Y13_LUT4AB/FrameStrobe[15] Tile_X8Y13_LUT4AB/FrameStrobe[16] Tile_X8Y13_LUT4AB/FrameStrobe[17]
+ Tile_X8Y13_LUT4AB/FrameStrobe[18] Tile_X8Y13_LUT4AB/FrameStrobe[19] Tile_X8Y13_LUT4AB/FrameStrobe[1]
+ Tile_X8Y13_LUT4AB/FrameStrobe[2] Tile_X8Y13_LUT4AB/FrameStrobe[3] Tile_X8Y13_LUT4AB/FrameStrobe[4]
+ Tile_X8Y13_LUT4AB/FrameStrobe[5] Tile_X8Y13_LUT4AB/FrameStrobe[6] Tile_X8Y13_LUT4AB/FrameStrobe[7]
+ Tile_X8Y13_LUT4AB/FrameStrobe[8] Tile_X8Y13_LUT4AB/FrameStrobe[9] Tile_X8Y12_LUT4AB/FrameStrobe[0]
+ Tile_X8Y12_LUT4AB/FrameStrobe[10] Tile_X8Y12_LUT4AB/FrameStrobe[11] Tile_X8Y12_LUT4AB/FrameStrobe[12]
+ Tile_X8Y12_LUT4AB/FrameStrobe[13] Tile_X8Y12_LUT4AB/FrameStrobe[14] Tile_X8Y12_LUT4AB/FrameStrobe[15]
+ Tile_X8Y12_LUT4AB/FrameStrobe[16] Tile_X8Y12_LUT4AB/FrameStrobe[17] Tile_X8Y12_LUT4AB/FrameStrobe[18]
+ Tile_X8Y12_LUT4AB/FrameStrobe[19] Tile_X8Y12_LUT4AB/FrameStrobe[1] Tile_X8Y12_LUT4AB/FrameStrobe[2]
+ Tile_X8Y12_LUT4AB/FrameStrobe[3] Tile_X8Y12_LUT4AB/FrameStrobe[4] Tile_X8Y12_LUT4AB/FrameStrobe[5]
+ Tile_X8Y12_LUT4AB/FrameStrobe[6] Tile_X8Y12_LUT4AB/FrameStrobe[7] Tile_X8Y12_LUT4AB/FrameStrobe[8]
+ Tile_X8Y12_LUT4AB/FrameStrobe[9] Tile_X8Y13_LUT4AB/N1BEG[0] Tile_X8Y13_LUT4AB/N1BEG[1]
+ Tile_X8Y13_LUT4AB/N1BEG[2] Tile_X8Y13_LUT4AB/N1BEG[3] Tile_X8Y14_LUT4AB/N1BEG[0]
+ Tile_X8Y14_LUT4AB/N1BEG[1] Tile_X8Y14_LUT4AB/N1BEG[2] Tile_X8Y14_LUT4AB/N1BEG[3]
+ Tile_X8Y13_LUT4AB/N2BEG[0] Tile_X8Y13_LUT4AB/N2BEG[1] Tile_X8Y13_LUT4AB/N2BEG[2]
+ Tile_X8Y13_LUT4AB/N2BEG[3] Tile_X8Y13_LUT4AB/N2BEG[4] Tile_X8Y13_LUT4AB/N2BEG[5]
+ Tile_X8Y13_LUT4AB/N2BEG[6] Tile_X8Y13_LUT4AB/N2BEG[7] Tile_X8Y12_LUT4AB/N2END[0]
+ Tile_X8Y12_LUT4AB/N2END[1] Tile_X8Y12_LUT4AB/N2END[2] Tile_X8Y12_LUT4AB/N2END[3]
+ Tile_X8Y12_LUT4AB/N2END[4] Tile_X8Y12_LUT4AB/N2END[5] Tile_X8Y12_LUT4AB/N2END[6]
+ Tile_X8Y12_LUT4AB/N2END[7] Tile_X8Y13_LUT4AB/N2END[0] Tile_X8Y13_LUT4AB/N2END[1]
+ Tile_X8Y13_LUT4AB/N2END[2] Tile_X8Y13_LUT4AB/N2END[3] Tile_X8Y13_LUT4AB/N2END[4]
+ Tile_X8Y13_LUT4AB/N2END[5] Tile_X8Y13_LUT4AB/N2END[6] Tile_X8Y13_LUT4AB/N2END[7]
+ Tile_X8Y14_LUT4AB/N2BEG[0] Tile_X8Y14_LUT4AB/N2BEG[1] Tile_X8Y14_LUT4AB/N2BEG[2]
+ Tile_X8Y14_LUT4AB/N2BEG[3] Tile_X8Y14_LUT4AB/N2BEG[4] Tile_X8Y14_LUT4AB/N2BEG[5]
+ Tile_X8Y14_LUT4AB/N2BEG[6] Tile_X8Y14_LUT4AB/N2BEG[7] Tile_X8Y13_LUT4AB/N4BEG[0]
+ Tile_X8Y13_LUT4AB/N4BEG[10] Tile_X8Y13_LUT4AB/N4BEG[11] Tile_X8Y13_LUT4AB/N4BEG[12]
+ Tile_X8Y13_LUT4AB/N4BEG[13] Tile_X8Y13_LUT4AB/N4BEG[14] Tile_X8Y13_LUT4AB/N4BEG[15]
+ Tile_X8Y13_LUT4AB/N4BEG[1] Tile_X8Y13_LUT4AB/N4BEG[2] Tile_X8Y13_LUT4AB/N4BEG[3]
+ Tile_X8Y13_LUT4AB/N4BEG[4] Tile_X8Y13_LUT4AB/N4BEG[5] Tile_X8Y13_LUT4AB/N4BEG[6]
+ Tile_X8Y13_LUT4AB/N4BEG[7] Tile_X8Y13_LUT4AB/N4BEG[8] Tile_X8Y13_LUT4AB/N4BEG[9]
+ Tile_X8Y14_LUT4AB/N4BEG[0] Tile_X8Y14_LUT4AB/N4BEG[10] Tile_X8Y14_LUT4AB/N4BEG[11]
+ Tile_X8Y14_LUT4AB/N4BEG[12] Tile_X8Y14_LUT4AB/N4BEG[13] Tile_X8Y14_LUT4AB/N4BEG[14]
+ Tile_X8Y14_LUT4AB/N4BEG[15] Tile_X8Y14_LUT4AB/N4BEG[1] Tile_X8Y14_LUT4AB/N4BEG[2]
+ Tile_X8Y14_LUT4AB/N4BEG[3] Tile_X8Y14_LUT4AB/N4BEG[4] Tile_X8Y14_LUT4AB/N4BEG[5]
+ Tile_X8Y14_LUT4AB/N4BEG[6] Tile_X8Y14_LUT4AB/N4BEG[7] Tile_X8Y14_LUT4AB/N4BEG[8]
+ Tile_X8Y14_LUT4AB/N4BEG[9] Tile_X8Y13_LUT4AB/NN4BEG[0] Tile_X8Y13_LUT4AB/NN4BEG[10]
+ Tile_X8Y13_LUT4AB/NN4BEG[11] Tile_X8Y13_LUT4AB/NN4BEG[12] Tile_X8Y13_LUT4AB/NN4BEG[13]
+ Tile_X8Y13_LUT4AB/NN4BEG[14] Tile_X8Y13_LUT4AB/NN4BEG[15] Tile_X8Y13_LUT4AB/NN4BEG[1]
+ Tile_X8Y13_LUT4AB/NN4BEG[2] Tile_X8Y13_LUT4AB/NN4BEG[3] Tile_X8Y13_LUT4AB/NN4BEG[4]
+ Tile_X8Y13_LUT4AB/NN4BEG[5] Tile_X8Y13_LUT4AB/NN4BEG[6] Tile_X8Y13_LUT4AB/NN4BEG[7]
+ Tile_X8Y13_LUT4AB/NN4BEG[8] Tile_X8Y13_LUT4AB/NN4BEG[9] Tile_X8Y14_LUT4AB/NN4BEG[0]
+ Tile_X8Y14_LUT4AB/NN4BEG[10] Tile_X8Y14_LUT4AB/NN4BEG[11] Tile_X8Y14_LUT4AB/NN4BEG[12]
+ Tile_X8Y14_LUT4AB/NN4BEG[13] Tile_X8Y14_LUT4AB/NN4BEG[14] Tile_X8Y14_LUT4AB/NN4BEG[15]
+ Tile_X8Y14_LUT4AB/NN4BEG[1] Tile_X8Y14_LUT4AB/NN4BEG[2] Tile_X8Y14_LUT4AB/NN4BEG[3]
+ Tile_X8Y14_LUT4AB/NN4BEG[4] Tile_X8Y14_LUT4AB/NN4BEG[5] Tile_X8Y14_LUT4AB/NN4BEG[6]
+ Tile_X8Y14_LUT4AB/NN4BEG[7] Tile_X8Y14_LUT4AB/NN4BEG[8] Tile_X8Y14_LUT4AB/NN4BEG[9]
+ Tile_X8Y14_LUT4AB/S1END[0] Tile_X8Y14_LUT4AB/S1END[1] Tile_X8Y14_LUT4AB/S1END[2]
+ Tile_X8Y14_LUT4AB/S1END[3] Tile_X8Y13_LUT4AB/S1END[0] Tile_X8Y13_LUT4AB/S1END[1]
+ Tile_X8Y13_LUT4AB/S1END[2] Tile_X8Y13_LUT4AB/S1END[3] Tile_X8Y14_LUT4AB/S2MID[0]
+ Tile_X8Y14_LUT4AB/S2MID[1] Tile_X8Y14_LUT4AB/S2MID[2] Tile_X8Y14_LUT4AB/S2MID[3]
+ Tile_X8Y14_LUT4AB/S2MID[4] Tile_X8Y14_LUT4AB/S2MID[5] Tile_X8Y14_LUT4AB/S2MID[6]
+ Tile_X8Y14_LUT4AB/S2MID[7] Tile_X8Y14_LUT4AB/S2END[0] Tile_X8Y14_LUT4AB/S2END[1]
+ Tile_X8Y14_LUT4AB/S2END[2] Tile_X8Y14_LUT4AB/S2END[3] Tile_X8Y14_LUT4AB/S2END[4]
+ Tile_X8Y14_LUT4AB/S2END[5] Tile_X8Y14_LUT4AB/S2END[6] Tile_X8Y14_LUT4AB/S2END[7]
+ Tile_X8Y13_LUT4AB/S2END[0] Tile_X8Y13_LUT4AB/S2END[1] Tile_X8Y13_LUT4AB/S2END[2]
+ Tile_X8Y13_LUT4AB/S2END[3] Tile_X8Y13_LUT4AB/S2END[4] Tile_X8Y13_LUT4AB/S2END[5]
+ Tile_X8Y13_LUT4AB/S2END[6] Tile_X8Y13_LUT4AB/S2END[7] Tile_X8Y13_LUT4AB/S2MID[0]
+ Tile_X8Y13_LUT4AB/S2MID[1] Tile_X8Y13_LUT4AB/S2MID[2] Tile_X8Y13_LUT4AB/S2MID[3]
+ Tile_X8Y13_LUT4AB/S2MID[4] Tile_X8Y13_LUT4AB/S2MID[5] Tile_X8Y13_LUT4AB/S2MID[6]
+ Tile_X8Y13_LUT4AB/S2MID[7] Tile_X8Y14_LUT4AB/S4END[0] Tile_X8Y14_LUT4AB/S4END[10]
+ Tile_X8Y14_LUT4AB/S4END[11] Tile_X8Y14_LUT4AB/S4END[12] Tile_X8Y14_LUT4AB/S4END[13]
+ Tile_X8Y14_LUT4AB/S4END[14] Tile_X8Y14_LUT4AB/S4END[15] Tile_X8Y14_LUT4AB/S4END[1]
+ Tile_X8Y14_LUT4AB/S4END[2] Tile_X8Y14_LUT4AB/S4END[3] Tile_X8Y14_LUT4AB/S4END[4]
+ Tile_X8Y14_LUT4AB/S4END[5] Tile_X8Y14_LUT4AB/S4END[6] Tile_X8Y14_LUT4AB/S4END[7]
+ Tile_X8Y14_LUT4AB/S4END[8] Tile_X8Y14_LUT4AB/S4END[9] Tile_X8Y13_LUT4AB/S4END[0]
+ Tile_X8Y13_LUT4AB/S4END[10] Tile_X8Y13_LUT4AB/S4END[11] Tile_X8Y13_LUT4AB/S4END[12]
+ Tile_X8Y13_LUT4AB/S4END[13] Tile_X8Y13_LUT4AB/S4END[14] Tile_X8Y13_LUT4AB/S4END[15]
+ Tile_X8Y13_LUT4AB/S4END[1] Tile_X8Y13_LUT4AB/S4END[2] Tile_X8Y13_LUT4AB/S4END[3]
+ Tile_X8Y13_LUT4AB/S4END[4] Tile_X8Y13_LUT4AB/S4END[5] Tile_X8Y13_LUT4AB/S4END[6]
+ Tile_X8Y13_LUT4AB/S4END[7] Tile_X8Y13_LUT4AB/S4END[8] Tile_X8Y13_LUT4AB/S4END[9]
+ Tile_X8Y14_LUT4AB/SS4END[0] Tile_X8Y14_LUT4AB/SS4END[10] Tile_X8Y14_LUT4AB/SS4END[11]
+ Tile_X8Y14_LUT4AB/SS4END[12] Tile_X8Y14_LUT4AB/SS4END[13] Tile_X8Y14_LUT4AB/SS4END[14]
+ Tile_X8Y14_LUT4AB/SS4END[15] Tile_X8Y14_LUT4AB/SS4END[1] Tile_X8Y14_LUT4AB/SS4END[2]
+ Tile_X8Y14_LUT4AB/SS4END[3] Tile_X8Y14_LUT4AB/SS4END[4] Tile_X8Y14_LUT4AB/SS4END[5]
+ Tile_X8Y14_LUT4AB/SS4END[6] Tile_X8Y14_LUT4AB/SS4END[7] Tile_X8Y14_LUT4AB/SS4END[8]
+ Tile_X8Y14_LUT4AB/SS4END[9] Tile_X8Y13_LUT4AB/SS4END[0] Tile_X8Y13_LUT4AB/SS4END[10]
+ Tile_X8Y13_LUT4AB/SS4END[11] Tile_X8Y13_LUT4AB/SS4END[12] Tile_X8Y13_LUT4AB/SS4END[13]
+ Tile_X8Y13_LUT4AB/SS4END[14] Tile_X8Y13_LUT4AB/SS4END[15] Tile_X8Y13_LUT4AB/SS4END[1]
+ Tile_X8Y13_LUT4AB/SS4END[2] Tile_X8Y13_LUT4AB/SS4END[3] Tile_X8Y13_LUT4AB/SS4END[4]
+ Tile_X8Y13_LUT4AB/SS4END[5] Tile_X8Y13_LUT4AB/SS4END[6] Tile_X8Y13_LUT4AB/SS4END[7]
+ Tile_X8Y13_LUT4AB/SS4END[8] Tile_X8Y13_LUT4AB/SS4END[9] Tile_X8Y13_LUT4AB/UserCLK
+ Tile_X8Y12_LUT4AB/UserCLK VGND VPWR Tile_X8Y13_LUT4AB/W1BEG[0] Tile_X8Y13_LUT4AB/W1BEG[1]
+ Tile_X8Y13_LUT4AB/W1BEG[2] Tile_X8Y13_LUT4AB/W1BEG[3] Tile_X9Y13_LUT4AB/W1BEG[0]
+ Tile_X9Y13_LUT4AB/W1BEG[1] Tile_X9Y13_LUT4AB/W1BEG[2] Tile_X9Y13_LUT4AB/W1BEG[3]
+ Tile_X8Y13_LUT4AB/W2BEG[0] Tile_X8Y13_LUT4AB/W2BEG[1] Tile_X8Y13_LUT4AB/W2BEG[2]
+ Tile_X8Y13_LUT4AB/W2BEG[3] Tile_X8Y13_LUT4AB/W2BEG[4] Tile_X8Y13_LUT4AB/W2BEG[5]
+ Tile_X8Y13_LUT4AB/W2BEG[6] Tile_X8Y13_LUT4AB/W2BEG[7] Tile_X8Y13_LUT4AB/W2BEGb[0]
+ Tile_X8Y13_LUT4AB/W2BEGb[1] Tile_X8Y13_LUT4AB/W2BEGb[2] Tile_X8Y13_LUT4AB/W2BEGb[3]
+ Tile_X8Y13_LUT4AB/W2BEGb[4] Tile_X8Y13_LUT4AB/W2BEGb[5] Tile_X8Y13_LUT4AB/W2BEGb[6]
+ Tile_X8Y13_LUT4AB/W2BEGb[7] Tile_X8Y13_LUT4AB/W2END[0] Tile_X8Y13_LUT4AB/W2END[1]
+ Tile_X8Y13_LUT4AB/W2END[2] Tile_X8Y13_LUT4AB/W2END[3] Tile_X8Y13_LUT4AB/W2END[4]
+ Tile_X8Y13_LUT4AB/W2END[5] Tile_X8Y13_LUT4AB/W2END[6] Tile_X8Y13_LUT4AB/W2END[7]
+ Tile_X9Y13_LUT4AB/W2BEG[0] Tile_X9Y13_LUT4AB/W2BEG[1] Tile_X9Y13_LUT4AB/W2BEG[2]
+ Tile_X9Y13_LUT4AB/W2BEG[3] Tile_X9Y13_LUT4AB/W2BEG[4] Tile_X9Y13_LUT4AB/W2BEG[5]
+ Tile_X9Y13_LUT4AB/W2BEG[6] Tile_X9Y13_LUT4AB/W2BEG[7] Tile_X8Y13_LUT4AB/W6BEG[0]
+ Tile_X8Y13_LUT4AB/W6BEG[10] Tile_X8Y13_LUT4AB/W6BEG[11] Tile_X8Y13_LUT4AB/W6BEG[1]
+ Tile_X8Y13_LUT4AB/W6BEG[2] Tile_X8Y13_LUT4AB/W6BEG[3] Tile_X8Y13_LUT4AB/W6BEG[4]
+ Tile_X8Y13_LUT4AB/W6BEG[5] Tile_X8Y13_LUT4AB/W6BEG[6] Tile_X8Y13_LUT4AB/W6BEG[7]
+ Tile_X8Y13_LUT4AB/W6BEG[8] Tile_X8Y13_LUT4AB/W6BEG[9] Tile_X9Y13_LUT4AB/W6BEG[0]
+ Tile_X9Y13_LUT4AB/W6BEG[10] Tile_X9Y13_LUT4AB/W6BEG[11] Tile_X9Y13_LUT4AB/W6BEG[1]
+ Tile_X9Y13_LUT4AB/W6BEG[2] Tile_X9Y13_LUT4AB/W6BEG[3] Tile_X9Y13_LUT4AB/W6BEG[4]
+ Tile_X9Y13_LUT4AB/W6BEG[5] Tile_X9Y13_LUT4AB/W6BEG[6] Tile_X9Y13_LUT4AB/W6BEG[7]
+ Tile_X9Y13_LUT4AB/W6BEG[8] Tile_X9Y13_LUT4AB/W6BEG[9] Tile_X8Y13_LUT4AB/WW4BEG[0]
+ Tile_X8Y13_LUT4AB/WW4BEG[10] Tile_X8Y13_LUT4AB/WW4BEG[11] Tile_X8Y13_LUT4AB/WW4BEG[12]
+ Tile_X8Y13_LUT4AB/WW4BEG[13] Tile_X8Y13_LUT4AB/WW4BEG[14] Tile_X8Y13_LUT4AB/WW4BEG[15]
+ Tile_X8Y13_LUT4AB/WW4BEG[1] Tile_X8Y13_LUT4AB/WW4BEG[2] Tile_X8Y13_LUT4AB/WW4BEG[3]
+ Tile_X8Y13_LUT4AB/WW4BEG[4] Tile_X8Y13_LUT4AB/WW4BEG[5] Tile_X8Y13_LUT4AB/WW4BEG[6]
+ Tile_X8Y13_LUT4AB/WW4BEG[7] Tile_X8Y13_LUT4AB/WW4BEG[8] Tile_X8Y13_LUT4AB/WW4BEG[9]
+ Tile_X9Y13_LUT4AB/WW4BEG[0] Tile_X9Y13_LUT4AB/WW4BEG[10] Tile_X9Y13_LUT4AB/WW4BEG[11]
+ Tile_X9Y13_LUT4AB/WW4BEG[12] Tile_X9Y13_LUT4AB/WW4BEG[13] Tile_X9Y13_LUT4AB/WW4BEG[14]
+ Tile_X9Y13_LUT4AB/WW4BEG[15] Tile_X9Y13_LUT4AB/WW4BEG[1] Tile_X9Y13_LUT4AB/WW4BEG[2]
+ Tile_X9Y13_LUT4AB/WW4BEG[3] Tile_X9Y13_LUT4AB/WW4BEG[4] Tile_X9Y13_LUT4AB/WW4BEG[5]
+ Tile_X9Y13_LUT4AB/WW4BEG[6] Tile_X9Y13_LUT4AB/WW4BEG[7] Tile_X9Y13_LUT4AB/WW4BEG[8]
+ Tile_X9Y13_LUT4AB/WW4BEG[9] LUT4AB
XTile_X2Y3_LUT4AB Tile_X2Y4_LUT4AB/Co Tile_X2Y3_LUT4AB/Co Tile_X3Y3_LUT4AB/E1END[0]
+ Tile_X3Y3_LUT4AB/E1END[1] Tile_X3Y3_LUT4AB/E1END[2] Tile_X3Y3_LUT4AB/E1END[3] Tile_X2Y3_LUT4AB/E1END[0]
+ Tile_X2Y3_LUT4AB/E1END[1] Tile_X2Y3_LUT4AB/E1END[2] Tile_X2Y3_LUT4AB/E1END[3] Tile_X3Y3_LUT4AB/E2MID[0]
+ Tile_X3Y3_LUT4AB/E2MID[1] Tile_X3Y3_LUT4AB/E2MID[2] Tile_X3Y3_LUT4AB/E2MID[3] Tile_X3Y3_LUT4AB/E2MID[4]
+ Tile_X3Y3_LUT4AB/E2MID[5] Tile_X3Y3_LUT4AB/E2MID[6] Tile_X3Y3_LUT4AB/E2MID[7] Tile_X3Y3_LUT4AB/E2END[0]
+ Tile_X3Y3_LUT4AB/E2END[1] Tile_X3Y3_LUT4AB/E2END[2] Tile_X3Y3_LUT4AB/E2END[3] Tile_X3Y3_LUT4AB/E2END[4]
+ Tile_X3Y3_LUT4AB/E2END[5] Tile_X3Y3_LUT4AB/E2END[6] Tile_X3Y3_LUT4AB/E2END[7] Tile_X2Y3_LUT4AB/E2END[0]
+ Tile_X2Y3_LUT4AB/E2END[1] Tile_X2Y3_LUT4AB/E2END[2] Tile_X2Y3_LUT4AB/E2END[3] Tile_X2Y3_LUT4AB/E2END[4]
+ Tile_X2Y3_LUT4AB/E2END[5] Tile_X2Y3_LUT4AB/E2END[6] Tile_X2Y3_LUT4AB/E2END[7] Tile_X2Y3_LUT4AB/E2MID[0]
+ Tile_X2Y3_LUT4AB/E2MID[1] Tile_X2Y3_LUT4AB/E2MID[2] Tile_X2Y3_LUT4AB/E2MID[3] Tile_X2Y3_LUT4AB/E2MID[4]
+ Tile_X2Y3_LUT4AB/E2MID[5] Tile_X2Y3_LUT4AB/E2MID[6] Tile_X2Y3_LUT4AB/E2MID[7] Tile_X3Y3_LUT4AB/E6END[0]
+ Tile_X3Y3_LUT4AB/E6END[10] Tile_X3Y3_LUT4AB/E6END[11] Tile_X3Y3_LUT4AB/E6END[1]
+ Tile_X3Y3_LUT4AB/E6END[2] Tile_X3Y3_LUT4AB/E6END[3] Tile_X3Y3_LUT4AB/E6END[4] Tile_X3Y3_LUT4AB/E6END[5]
+ Tile_X3Y3_LUT4AB/E6END[6] Tile_X3Y3_LUT4AB/E6END[7] Tile_X3Y3_LUT4AB/E6END[8] Tile_X3Y3_LUT4AB/E6END[9]
+ Tile_X2Y3_LUT4AB/E6END[0] Tile_X2Y3_LUT4AB/E6END[10] Tile_X2Y3_LUT4AB/E6END[11]
+ Tile_X2Y3_LUT4AB/E6END[1] Tile_X2Y3_LUT4AB/E6END[2] Tile_X2Y3_LUT4AB/E6END[3] Tile_X2Y3_LUT4AB/E6END[4]
+ Tile_X2Y3_LUT4AB/E6END[5] Tile_X2Y3_LUT4AB/E6END[6] Tile_X2Y3_LUT4AB/E6END[7] Tile_X2Y3_LUT4AB/E6END[8]
+ Tile_X2Y3_LUT4AB/E6END[9] Tile_X3Y3_LUT4AB/EE4END[0] Tile_X3Y3_LUT4AB/EE4END[10]
+ Tile_X3Y3_LUT4AB/EE4END[11] Tile_X3Y3_LUT4AB/EE4END[12] Tile_X3Y3_LUT4AB/EE4END[13]
+ Tile_X3Y3_LUT4AB/EE4END[14] Tile_X3Y3_LUT4AB/EE4END[15] Tile_X3Y3_LUT4AB/EE4END[1]
+ Tile_X3Y3_LUT4AB/EE4END[2] Tile_X3Y3_LUT4AB/EE4END[3] Tile_X3Y3_LUT4AB/EE4END[4]
+ Tile_X3Y3_LUT4AB/EE4END[5] Tile_X3Y3_LUT4AB/EE4END[6] Tile_X3Y3_LUT4AB/EE4END[7]
+ Tile_X3Y3_LUT4AB/EE4END[8] Tile_X3Y3_LUT4AB/EE4END[9] Tile_X2Y3_LUT4AB/EE4END[0]
+ Tile_X2Y3_LUT4AB/EE4END[10] Tile_X2Y3_LUT4AB/EE4END[11] Tile_X2Y3_LUT4AB/EE4END[12]
+ Tile_X2Y3_LUT4AB/EE4END[13] Tile_X2Y3_LUT4AB/EE4END[14] Tile_X2Y3_LUT4AB/EE4END[15]
+ Tile_X2Y3_LUT4AB/EE4END[1] Tile_X2Y3_LUT4AB/EE4END[2] Tile_X2Y3_LUT4AB/EE4END[3]
+ Tile_X2Y3_LUT4AB/EE4END[4] Tile_X2Y3_LUT4AB/EE4END[5] Tile_X2Y3_LUT4AB/EE4END[6]
+ Tile_X2Y3_LUT4AB/EE4END[7] Tile_X2Y3_LUT4AB/EE4END[8] Tile_X2Y3_LUT4AB/EE4END[9]
+ Tile_X2Y3_LUT4AB/FrameData[0] Tile_X2Y3_LUT4AB/FrameData[10] Tile_X2Y3_LUT4AB/FrameData[11]
+ Tile_X2Y3_LUT4AB/FrameData[12] Tile_X2Y3_LUT4AB/FrameData[13] Tile_X2Y3_LUT4AB/FrameData[14]
+ Tile_X2Y3_LUT4AB/FrameData[15] Tile_X2Y3_LUT4AB/FrameData[16] Tile_X2Y3_LUT4AB/FrameData[17]
+ Tile_X2Y3_LUT4AB/FrameData[18] Tile_X2Y3_LUT4AB/FrameData[19] Tile_X2Y3_LUT4AB/FrameData[1]
+ Tile_X2Y3_LUT4AB/FrameData[20] Tile_X2Y3_LUT4AB/FrameData[21] Tile_X2Y3_LUT4AB/FrameData[22]
+ Tile_X2Y3_LUT4AB/FrameData[23] Tile_X2Y3_LUT4AB/FrameData[24] Tile_X2Y3_LUT4AB/FrameData[25]
+ Tile_X2Y3_LUT4AB/FrameData[26] Tile_X2Y3_LUT4AB/FrameData[27] Tile_X2Y3_LUT4AB/FrameData[28]
+ Tile_X2Y3_LUT4AB/FrameData[29] Tile_X2Y3_LUT4AB/FrameData[2] Tile_X2Y3_LUT4AB/FrameData[30]
+ Tile_X2Y3_LUT4AB/FrameData[31] Tile_X2Y3_LUT4AB/FrameData[3] Tile_X2Y3_LUT4AB/FrameData[4]
+ Tile_X2Y3_LUT4AB/FrameData[5] Tile_X2Y3_LUT4AB/FrameData[6] Tile_X2Y3_LUT4AB/FrameData[7]
+ Tile_X2Y3_LUT4AB/FrameData[8] Tile_X2Y3_LUT4AB/FrameData[9] Tile_X3Y3_LUT4AB/FrameData[0]
+ Tile_X3Y3_LUT4AB/FrameData[10] Tile_X3Y3_LUT4AB/FrameData[11] Tile_X3Y3_LUT4AB/FrameData[12]
+ Tile_X3Y3_LUT4AB/FrameData[13] Tile_X3Y3_LUT4AB/FrameData[14] Tile_X3Y3_LUT4AB/FrameData[15]
+ Tile_X3Y3_LUT4AB/FrameData[16] Tile_X3Y3_LUT4AB/FrameData[17] Tile_X3Y3_LUT4AB/FrameData[18]
+ Tile_X3Y3_LUT4AB/FrameData[19] Tile_X3Y3_LUT4AB/FrameData[1] Tile_X3Y3_LUT4AB/FrameData[20]
+ Tile_X3Y3_LUT4AB/FrameData[21] Tile_X3Y3_LUT4AB/FrameData[22] Tile_X3Y3_LUT4AB/FrameData[23]
+ Tile_X3Y3_LUT4AB/FrameData[24] Tile_X3Y3_LUT4AB/FrameData[25] Tile_X3Y3_LUT4AB/FrameData[26]
+ Tile_X3Y3_LUT4AB/FrameData[27] Tile_X3Y3_LUT4AB/FrameData[28] Tile_X3Y3_LUT4AB/FrameData[29]
+ Tile_X3Y3_LUT4AB/FrameData[2] Tile_X3Y3_LUT4AB/FrameData[30] Tile_X3Y3_LUT4AB/FrameData[31]
+ Tile_X3Y3_LUT4AB/FrameData[3] Tile_X3Y3_LUT4AB/FrameData[4] Tile_X3Y3_LUT4AB/FrameData[5]
+ Tile_X3Y3_LUT4AB/FrameData[6] Tile_X3Y3_LUT4AB/FrameData[7] Tile_X3Y3_LUT4AB/FrameData[8]
+ Tile_X3Y3_LUT4AB/FrameData[9] Tile_X2Y3_LUT4AB/FrameStrobe[0] Tile_X2Y3_LUT4AB/FrameStrobe[10]
+ Tile_X2Y3_LUT4AB/FrameStrobe[11] Tile_X2Y3_LUT4AB/FrameStrobe[12] Tile_X2Y3_LUT4AB/FrameStrobe[13]
+ Tile_X2Y3_LUT4AB/FrameStrobe[14] Tile_X2Y3_LUT4AB/FrameStrobe[15] Tile_X2Y3_LUT4AB/FrameStrobe[16]
+ Tile_X2Y3_LUT4AB/FrameStrobe[17] Tile_X2Y3_LUT4AB/FrameStrobe[18] Tile_X2Y3_LUT4AB/FrameStrobe[19]
+ Tile_X2Y3_LUT4AB/FrameStrobe[1] Tile_X2Y3_LUT4AB/FrameStrobe[2] Tile_X2Y3_LUT4AB/FrameStrobe[3]
+ Tile_X2Y3_LUT4AB/FrameStrobe[4] Tile_X2Y3_LUT4AB/FrameStrobe[5] Tile_X2Y3_LUT4AB/FrameStrobe[6]
+ Tile_X2Y3_LUT4AB/FrameStrobe[7] Tile_X2Y3_LUT4AB/FrameStrobe[8] Tile_X2Y3_LUT4AB/FrameStrobe[9]
+ Tile_X2Y2_LUT4AB/FrameStrobe[0] Tile_X2Y2_LUT4AB/FrameStrobe[10] Tile_X2Y2_LUT4AB/FrameStrobe[11]
+ Tile_X2Y2_LUT4AB/FrameStrobe[12] Tile_X2Y2_LUT4AB/FrameStrobe[13] Tile_X2Y2_LUT4AB/FrameStrobe[14]
+ Tile_X2Y2_LUT4AB/FrameStrobe[15] Tile_X2Y2_LUT4AB/FrameStrobe[16] Tile_X2Y2_LUT4AB/FrameStrobe[17]
+ Tile_X2Y2_LUT4AB/FrameStrobe[18] Tile_X2Y2_LUT4AB/FrameStrobe[19] Tile_X2Y2_LUT4AB/FrameStrobe[1]
+ Tile_X2Y2_LUT4AB/FrameStrobe[2] Tile_X2Y2_LUT4AB/FrameStrobe[3] Tile_X2Y2_LUT4AB/FrameStrobe[4]
+ Tile_X2Y2_LUT4AB/FrameStrobe[5] Tile_X2Y2_LUT4AB/FrameStrobe[6] Tile_X2Y2_LUT4AB/FrameStrobe[7]
+ Tile_X2Y2_LUT4AB/FrameStrobe[8] Tile_X2Y2_LUT4AB/FrameStrobe[9] Tile_X2Y3_LUT4AB/N1BEG[0]
+ Tile_X2Y3_LUT4AB/N1BEG[1] Tile_X2Y3_LUT4AB/N1BEG[2] Tile_X2Y3_LUT4AB/N1BEG[3] Tile_X2Y4_LUT4AB/N1BEG[0]
+ Tile_X2Y4_LUT4AB/N1BEG[1] Tile_X2Y4_LUT4AB/N1BEG[2] Tile_X2Y4_LUT4AB/N1BEG[3] Tile_X2Y3_LUT4AB/N2BEG[0]
+ Tile_X2Y3_LUT4AB/N2BEG[1] Tile_X2Y3_LUT4AB/N2BEG[2] Tile_X2Y3_LUT4AB/N2BEG[3] Tile_X2Y3_LUT4AB/N2BEG[4]
+ Tile_X2Y3_LUT4AB/N2BEG[5] Tile_X2Y3_LUT4AB/N2BEG[6] Tile_X2Y3_LUT4AB/N2BEG[7] Tile_X2Y2_LUT4AB/N2END[0]
+ Tile_X2Y2_LUT4AB/N2END[1] Tile_X2Y2_LUT4AB/N2END[2] Tile_X2Y2_LUT4AB/N2END[3] Tile_X2Y2_LUT4AB/N2END[4]
+ Tile_X2Y2_LUT4AB/N2END[5] Tile_X2Y2_LUT4AB/N2END[6] Tile_X2Y2_LUT4AB/N2END[7] Tile_X2Y3_LUT4AB/N2END[0]
+ Tile_X2Y3_LUT4AB/N2END[1] Tile_X2Y3_LUT4AB/N2END[2] Tile_X2Y3_LUT4AB/N2END[3] Tile_X2Y3_LUT4AB/N2END[4]
+ Tile_X2Y3_LUT4AB/N2END[5] Tile_X2Y3_LUT4AB/N2END[6] Tile_X2Y3_LUT4AB/N2END[7] Tile_X2Y4_LUT4AB/N2BEG[0]
+ Tile_X2Y4_LUT4AB/N2BEG[1] Tile_X2Y4_LUT4AB/N2BEG[2] Tile_X2Y4_LUT4AB/N2BEG[3] Tile_X2Y4_LUT4AB/N2BEG[4]
+ Tile_X2Y4_LUT4AB/N2BEG[5] Tile_X2Y4_LUT4AB/N2BEG[6] Tile_X2Y4_LUT4AB/N2BEG[7] Tile_X2Y3_LUT4AB/N4BEG[0]
+ Tile_X2Y3_LUT4AB/N4BEG[10] Tile_X2Y3_LUT4AB/N4BEG[11] Tile_X2Y3_LUT4AB/N4BEG[12]
+ Tile_X2Y3_LUT4AB/N4BEG[13] Tile_X2Y3_LUT4AB/N4BEG[14] Tile_X2Y3_LUT4AB/N4BEG[15]
+ Tile_X2Y3_LUT4AB/N4BEG[1] Tile_X2Y3_LUT4AB/N4BEG[2] Tile_X2Y3_LUT4AB/N4BEG[3] Tile_X2Y3_LUT4AB/N4BEG[4]
+ Tile_X2Y3_LUT4AB/N4BEG[5] Tile_X2Y3_LUT4AB/N4BEG[6] Tile_X2Y3_LUT4AB/N4BEG[7] Tile_X2Y3_LUT4AB/N4BEG[8]
+ Tile_X2Y3_LUT4AB/N4BEG[9] Tile_X2Y4_LUT4AB/N4BEG[0] Tile_X2Y4_LUT4AB/N4BEG[10] Tile_X2Y4_LUT4AB/N4BEG[11]
+ Tile_X2Y4_LUT4AB/N4BEG[12] Tile_X2Y4_LUT4AB/N4BEG[13] Tile_X2Y4_LUT4AB/N4BEG[14]
+ Tile_X2Y4_LUT4AB/N4BEG[15] Tile_X2Y4_LUT4AB/N4BEG[1] Tile_X2Y4_LUT4AB/N4BEG[2] Tile_X2Y4_LUT4AB/N4BEG[3]
+ Tile_X2Y4_LUT4AB/N4BEG[4] Tile_X2Y4_LUT4AB/N4BEG[5] Tile_X2Y4_LUT4AB/N4BEG[6] Tile_X2Y4_LUT4AB/N4BEG[7]
+ Tile_X2Y4_LUT4AB/N4BEG[8] Tile_X2Y4_LUT4AB/N4BEG[9] Tile_X2Y3_LUT4AB/NN4BEG[0] Tile_X2Y3_LUT4AB/NN4BEG[10]
+ Tile_X2Y3_LUT4AB/NN4BEG[11] Tile_X2Y3_LUT4AB/NN4BEG[12] Tile_X2Y3_LUT4AB/NN4BEG[13]
+ Tile_X2Y3_LUT4AB/NN4BEG[14] Tile_X2Y3_LUT4AB/NN4BEG[15] Tile_X2Y3_LUT4AB/NN4BEG[1]
+ Tile_X2Y3_LUT4AB/NN4BEG[2] Tile_X2Y3_LUT4AB/NN4BEG[3] Tile_X2Y3_LUT4AB/NN4BEG[4]
+ Tile_X2Y3_LUT4AB/NN4BEG[5] Tile_X2Y3_LUT4AB/NN4BEG[6] Tile_X2Y3_LUT4AB/NN4BEG[7]
+ Tile_X2Y3_LUT4AB/NN4BEG[8] Tile_X2Y3_LUT4AB/NN4BEG[9] Tile_X2Y4_LUT4AB/NN4BEG[0]
+ Tile_X2Y4_LUT4AB/NN4BEG[10] Tile_X2Y4_LUT4AB/NN4BEG[11] Tile_X2Y4_LUT4AB/NN4BEG[12]
+ Tile_X2Y4_LUT4AB/NN4BEG[13] Tile_X2Y4_LUT4AB/NN4BEG[14] Tile_X2Y4_LUT4AB/NN4BEG[15]
+ Tile_X2Y4_LUT4AB/NN4BEG[1] Tile_X2Y4_LUT4AB/NN4BEG[2] Tile_X2Y4_LUT4AB/NN4BEG[3]
+ Tile_X2Y4_LUT4AB/NN4BEG[4] Tile_X2Y4_LUT4AB/NN4BEG[5] Tile_X2Y4_LUT4AB/NN4BEG[6]
+ Tile_X2Y4_LUT4AB/NN4BEG[7] Tile_X2Y4_LUT4AB/NN4BEG[8] Tile_X2Y4_LUT4AB/NN4BEG[9]
+ Tile_X2Y4_LUT4AB/S1END[0] Tile_X2Y4_LUT4AB/S1END[1] Tile_X2Y4_LUT4AB/S1END[2] Tile_X2Y4_LUT4AB/S1END[3]
+ Tile_X2Y3_LUT4AB/S1END[0] Tile_X2Y3_LUT4AB/S1END[1] Tile_X2Y3_LUT4AB/S1END[2] Tile_X2Y3_LUT4AB/S1END[3]
+ Tile_X2Y4_LUT4AB/S2MID[0] Tile_X2Y4_LUT4AB/S2MID[1] Tile_X2Y4_LUT4AB/S2MID[2] Tile_X2Y4_LUT4AB/S2MID[3]
+ Tile_X2Y4_LUT4AB/S2MID[4] Tile_X2Y4_LUT4AB/S2MID[5] Tile_X2Y4_LUT4AB/S2MID[6] Tile_X2Y4_LUT4AB/S2MID[7]
+ Tile_X2Y4_LUT4AB/S2END[0] Tile_X2Y4_LUT4AB/S2END[1] Tile_X2Y4_LUT4AB/S2END[2] Tile_X2Y4_LUT4AB/S2END[3]
+ Tile_X2Y4_LUT4AB/S2END[4] Tile_X2Y4_LUT4AB/S2END[5] Tile_X2Y4_LUT4AB/S2END[6] Tile_X2Y4_LUT4AB/S2END[7]
+ Tile_X2Y3_LUT4AB/S2END[0] Tile_X2Y3_LUT4AB/S2END[1] Tile_X2Y3_LUT4AB/S2END[2] Tile_X2Y3_LUT4AB/S2END[3]
+ Tile_X2Y3_LUT4AB/S2END[4] Tile_X2Y3_LUT4AB/S2END[5] Tile_X2Y3_LUT4AB/S2END[6] Tile_X2Y3_LUT4AB/S2END[7]
+ Tile_X2Y3_LUT4AB/S2MID[0] Tile_X2Y3_LUT4AB/S2MID[1] Tile_X2Y3_LUT4AB/S2MID[2] Tile_X2Y3_LUT4AB/S2MID[3]
+ Tile_X2Y3_LUT4AB/S2MID[4] Tile_X2Y3_LUT4AB/S2MID[5] Tile_X2Y3_LUT4AB/S2MID[6] Tile_X2Y3_LUT4AB/S2MID[7]
+ Tile_X2Y4_LUT4AB/S4END[0] Tile_X2Y4_LUT4AB/S4END[10] Tile_X2Y4_LUT4AB/S4END[11]
+ Tile_X2Y4_LUT4AB/S4END[12] Tile_X2Y4_LUT4AB/S4END[13] Tile_X2Y4_LUT4AB/S4END[14]
+ Tile_X2Y4_LUT4AB/S4END[15] Tile_X2Y4_LUT4AB/S4END[1] Tile_X2Y4_LUT4AB/S4END[2] Tile_X2Y4_LUT4AB/S4END[3]
+ Tile_X2Y4_LUT4AB/S4END[4] Tile_X2Y4_LUT4AB/S4END[5] Tile_X2Y4_LUT4AB/S4END[6] Tile_X2Y4_LUT4AB/S4END[7]
+ Tile_X2Y4_LUT4AB/S4END[8] Tile_X2Y4_LUT4AB/S4END[9] Tile_X2Y3_LUT4AB/S4END[0] Tile_X2Y3_LUT4AB/S4END[10]
+ Tile_X2Y3_LUT4AB/S4END[11] Tile_X2Y3_LUT4AB/S4END[12] Tile_X2Y3_LUT4AB/S4END[13]
+ Tile_X2Y3_LUT4AB/S4END[14] Tile_X2Y3_LUT4AB/S4END[15] Tile_X2Y3_LUT4AB/S4END[1]
+ Tile_X2Y3_LUT4AB/S4END[2] Tile_X2Y3_LUT4AB/S4END[3] Tile_X2Y3_LUT4AB/S4END[4] Tile_X2Y3_LUT4AB/S4END[5]
+ Tile_X2Y3_LUT4AB/S4END[6] Tile_X2Y3_LUT4AB/S4END[7] Tile_X2Y3_LUT4AB/S4END[8] Tile_X2Y3_LUT4AB/S4END[9]
+ Tile_X2Y4_LUT4AB/SS4END[0] Tile_X2Y4_LUT4AB/SS4END[10] Tile_X2Y4_LUT4AB/SS4END[11]
+ Tile_X2Y4_LUT4AB/SS4END[12] Tile_X2Y4_LUT4AB/SS4END[13] Tile_X2Y4_LUT4AB/SS4END[14]
+ Tile_X2Y4_LUT4AB/SS4END[15] Tile_X2Y4_LUT4AB/SS4END[1] Tile_X2Y4_LUT4AB/SS4END[2]
+ Tile_X2Y4_LUT4AB/SS4END[3] Tile_X2Y4_LUT4AB/SS4END[4] Tile_X2Y4_LUT4AB/SS4END[5]
+ Tile_X2Y4_LUT4AB/SS4END[6] Tile_X2Y4_LUT4AB/SS4END[7] Tile_X2Y4_LUT4AB/SS4END[8]
+ Tile_X2Y4_LUT4AB/SS4END[9] Tile_X2Y3_LUT4AB/SS4END[0] Tile_X2Y3_LUT4AB/SS4END[10]
+ Tile_X2Y3_LUT4AB/SS4END[11] Tile_X2Y3_LUT4AB/SS4END[12] Tile_X2Y3_LUT4AB/SS4END[13]
+ Tile_X2Y3_LUT4AB/SS4END[14] Tile_X2Y3_LUT4AB/SS4END[15] Tile_X2Y3_LUT4AB/SS4END[1]
+ Tile_X2Y3_LUT4AB/SS4END[2] Tile_X2Y3_LUT4AB/SS4END[3] Tile_X2Y3_LUT4AB/SS4END[4]
+ Tile_X2Y3_LUT4AB/SS4END[5] Tile_X2Y3_LUT4AB/SS4END[6] Tile_X2Y3_LUT4AB/SS4END[7]
+ Tile_X2Y3_LUT4AB/SS4END[8] Tile_X2Y3_LUT4AB/SS4END[9] Tile_X2Y3_LUT4AB/UserCLK Tile_X2Y2_LUT4AB/UserCLK
+ VGND VPWR Tile_X2Y3_LUT4AB/W1BEG[0] Tile_X2Y3_LUT4AB/W1BEG[1] Tile_X2Y3_LUT4AB/W1BEG[2]
+ Tile_X2Y3_LUT4AB/W1BEG[3] Tile_X3Y3_LUT4AB/W1BEG[0] Tile_X3Y3_LUT4AB/W1BEG[1] Tile_X3Y3_LUT4AB/W1BEG[2]
+ Tile_X3Y3_LUT4AB/W1BEG[3] Tile_X2Y3_LUT4AB/W2BEG[0] Tile_X2Y3_LUT4AB/W2BEG[1] Tile_X2Y3_LUT4AB/W2BEG[2]
+ Tile_X2Y3_LUT4AB/W2BEG[3] Tile_X2Y3_LUT4AB/W2BEG[4] Tile_X2Y3_LUT4AB/W2BEG[5] Tile_X2Y3_LUT4AB/W2BEG[6]
+ Tile_X2Y3_LUT4AB/W2BEG[7] Tile_X1Y3_LUT4AB/W2END[0] Tile_X1Y3_LUT4AB/W2END[1] Tile_X1Y3_LUT4AB/W2END[2]
+ Tile_X1Y3_LUT4AB/W2END[3] Tile_X1Y3_LUT4AB/W2END[4] Tile_X1Y3_LUT4AB/W2END[5] Tile_X1Y3_LUT4AB/W2END[6]
+ Tile_X1Y3_LUT4AB/W2END[7] Tile_X2Y3_LUT4AB/W2END[0] Tile_X2Y3_LUT4AB/W2END[1] Tile_X2Y3_LUT4AB/W2END[2]
+ Tile_X2Y3_LUT4AB/W2END[3] Tile_X2Y3_LUT4AB/W2END[4] Tile_X2Y3_LUT4AB/W2END[5] Tile_X2Y3_LUT4AB/W2END[6]
+ Tile_X2Y3_LUT4AB/W2END[7] Tile_X3Y3_LUT4AB/W2BEG[0] Tile_X3Y3_LUT4AB/W2BEG[1] Tile_X3Y3_LUT4AB/W2BEG[2]
+ Tile_X3Y3_LUT4AB/W2BEG[3] Tile_X3Y3_LUT4AB/W2BEG[4] Tile_X3Y3_LUT4AB/W2BEG[5] Tile_X3Y3_LUT4AB/W2BEG[6]
+ Tile_X3Y3_LUT4AB/W2BEG[7] Tile_X2Y3_LUT4AB/W6BEG[0] Tile_X2Y3_LUT4AB/W6BEG[10] Tile_X2Y3_LUT4AB/W6BEG[11]
+ Tile_X2Y3_LUT4AB/W6BEG[1] Tile_X2Y3_LUT4AB/W6BEG[2] Tile_X2Y3_LUT4AB/W6BEG[3] Tile_X2Y3_LUT4AB/W6BEG[4]
+ Tile_X2Y3_LUT4AB/W6BEG[5] Tile_X2Y3_LUT4AB/W6BEG[6] Tile_X2Y3_LUT4AB/W6BEG[7] Tile_X2Y3_LUT4AB/W6BEG[8]
+ Tile_X2Y3_LUT4AB/W6BEG[9] Tile_X3Y3_LUT4AB/W6BEG[0] Tile_X3Y3_LUT4AB/W6BEG[10] Tile_X3Y3_LUT4AB/W6BEG[11]
+ Tile_X3Y3_LUT4AB/W6BEG[1] Tile_X3Y3_LUT4AB/W6BEG[2] Tile_X3Y3_LUT4AB/W6BEG[3] Tile_X3Y3_LUT4AB/W6BEG[4]
+ Tile_X3Y3_LUT4AB/W6BEG[5] Tile_X3Y3_LUT4AB/W6BEG[6] Tile_X3Y3_LUT4AB/W6BEG[7] Tile_X3Y3_LUT4AB/W6BEG[8]
+ Tile_X3Y3_LUT4AB/W6BEG[9] Tile_X2Y3_LUT4AB/WW4BEG[0] Tile_X2Y3_LUT4AB/WW4BEG[10]
+ Tile_X2Y3_LUT4AB/WW4BEG[11] Tile_X2Y3_LUT4AB/WW4BEG[12] Tile_X2Y3_LUT4AB/WW4BEG[13]
+ Tile_X2Y3_LUT4AB/WW4BEG[14] Tile_X2Y3_LUT4AB/WW4BEG[15] Tile_X2Y3_LUT4AB/WW4BEG[1]
+ Tile_X2Y3_LUT4AB/WW4BEG[2] Tile_X2Y3_LUT4AB/WW4BEG[3] Tile_X2Y3_LUT4AB/WW4BEG[4]
+ Tile_X2Y3_LUT4AB/WW4BEG[5] Tile_X2Y3_LUT4AB/WW4BEG[6] Tile_X2Y3_LUT4AB/WW4BEG[7]
+ Tile_X2Y3_LUT4AB/WW4BEG[8] Tile_X2Y3_LUT4AB/WW4BEG[9] Tile_X3Y3_LUT4AB/WW4BEG[0]
+ Tile_X3Y3_LUT4AB/WW4BEG[10] Tile_X3Y3_LUT4AB/WW4BEG[11] Tile_X3Y3_LUT4AB/WW4BEG[12]
+ Tile_X3Y3_LUT4AB/WW4BEG[13] Tile_X3Y3_LUT4AB/WW4BEG[14] Tile_X3Y3_LUT4AB/WW4BEG[15]
+ Tile_X3Y3_LUT4AB/WW4BEG[1] Tile_X3Y3_LUT4AB/WW4BEG[2] Tile_X3Y3_LUT4AB/WW4BEG[3]
+ Tile_X3Y3_LUT4AB/WW4BEG[4] Tile_X3Y3_LUT4AB/WW4BEG[5] Tile_X3Y3_LUT4AB/WW4BEG[6]
+ Tile_X3Y3_LUT4AB/WW4BEG[7] Tile_X3Y3_LUT4AB/WW4BEG[8] Tile_X3Y3_LUT4AB/WW4BEG[9]
+ LUT4AB
XTile_X5Y8_LUT4AB Tile_X5Y9_LUT4AB/Co Tile_X5Y8_LUT4AB/Co Tile_X6Y8_LUT4AB/E1END[0]
+ Tile_X6Y8_LUT4AB/E1END[1] Tile_X6Y8_LUT4AB/E1END[2] Tile_X6Y8_LUT4AB/E1END[3] Tile_X5Y8_LUT4AB/E1END[0]
+ Tile_X5Y8_LUT4AB/E1END[1] Tile_X5Y8_LUT4AB/E1END[2] Tile_X5Y8_LUT4AB/E1END[3] Tile_X6Y8_LUT4AB/E2MID[0]
+ Tile_X6Y8_LUT4AB/E2MID[1] Tile_X6Y8_LUT4AB/E2MID[2] Tile_X6Y8_LUT4AB/E2MID[3] Tile_X6Y8_LUT4AB/E2MID[4]
+ Tile_X6Y8_LUT4AB/E2MID[5] Tile_X6Y8_LUT4AB/E2MID[6] Tile_X6Y8_LUT4AB/E2MID[7] Tile_X6Y8_LUT4AB/E2END[0]
+ Tile_X6Y8_LUT4AB/E2END[1] Tile_X6Y8_LUT4AB/E2END[2] Tile_X6Y8_LUT4AB/E2END[3] Tile_X6Y8_LUT4AB/E2END[4]
+ Tile_X6Y8_LUT4AB/E2END[5] Tile_X6Y8_LUT4AB/E2END[6] Tile_X6Y8_LUT4AB/E2END[7] Tile_X5Y8_LUT4AB/E2END[0]
+ Tile_X5Y8_LUT4AB/E2END[1] Tile_X5Y8_LUT4AB/E2END[2] Tile_X5Y8_LUT4AB/E2END[3] Tile_X5Y8_LUT4AB/E2END[4]
+ Tile_X5Y8_LUT4AB/E2END[5] Tile_X5Y8_LUT4AB/E2END[6] Tile_X5Y8_LUT4AB/E2END[7] Tile_X5Y8_LUT4AB/E2MID[0]
+ Tile_X5Y8_LUT4AB/E2MID[1] Tile_X5Y8_LUT4AB/E2MID[2] Tile_X5Y8_LUT4AB/E2MID[3] Tile_X5Y8_LUT4AB/E2MID[4]
+ Tile_X5Y8_LUT4AB/E2MID[5] Tile_X5Y8_LUT4AB/E2MID[6] Tile_X5Y8_LUT4AB/E2MID[7] Tile_X6Y8_LUT4AB/E6END[0]
+ Tile_X6Y8_LUT4AB/E6END[10] Tile_X6Y8_LUT4AB/E6END[11] Tile_X6Y8_LUT4AB/E6END[1]
+ Tile_X6Y8_LUT4AB/E6END[2] Tile_X6Y8_LUT4AB/E6END[3] Tile_X6Y8_LUT4AB/E6END[4] Tile_X6Y8_LUT4AB/E6END[5]
+ Tile_X6Y8_LUT4AB/E6END[6] Tile_X6Y8_LUT4AB/E6END[7] Tile_X6Y8_LUT4AB/E6END[8] Tile_X6Y8_LUT4AB/E6END[9]
+ Tile_X5Y8_LUT4AB/E6END[0] Tile_X5Y8_LUT4AB/E6END[10] Tile_X5Y8_LUT4AB/E6END[11]
+ Tile_X5Y8_LUT4AB/E6END[1] Tile_X5Y8_LUT4AB/E6END[2] Tile_X5Y8_LUT4AB/E6END[3] Tile_X5Y8_LUT4AB/E6END[4]
+ Tile_X5Y8_LUT4AB/E6END[5] Tile_X5Y8_LUT4AB/E6END[6] Tile_X5Y8_LUT4AB/E6END[7] Tile_X5Y8_LUT4AB/E6END[8]
+ Tile_X5Y8_LUT4AB/E6END[9] Tile_X6Y8_LUT4AB/EE4END[0] Tile_X6Y8_LUT4AB/EE4END[10]
+ Tile_X6Y8_LUT4AB/EE4END[11] Tile_X6Y8_LUT4AB/EE4END[12] Tile_X6Y8_LUT4AB/EE4END[13]
+ Tile_X6Y8_LUT4AB/EE4END[14] Tile_X6Y8_LUT4AB/EE4END[15] Tile_X6Y8_LUT4AB/EE4END[1]
+ Tile_X6Y8_LUT4AB/EE4END[2] Tile_X6Y8_LUT4AB/EE4END[3] Tile_X6Y8_LUT4AB/EE4END[4]
+ Tile_X6Y8_LUT4AB/EE4END[5] Tile_X6Y8_LUT4AB/EE4END[6] Tile_X6Y8_LUT4AB/EE4END[7]
+ Tile_X6Y8_LUT4AB/EE4END[8] Tile_X6Y8_LUT4AB/EE4END[9] Tile_X5Y8_LUT4AB/EE4END[0]
+ Tile_X5Y8_LUT4AB/EE4END[10] Tile_X5Y8_LUT4AB/EE4END[11] Tile_X5Y8_LUT4AB/EE4END[12]
+ Tile_X5Y8_LUT4AB/EE4END[13] Tile_X5Y8_LUT4AB/EE4END[14] Tile_X5Y8_LUT4AB/EE4END[15]
+ Tile_X5Y8_LUT4AB/EE4END[1] Tile_X5Y8_LUT4AB/EE4END[2] Tile_X5Y8_LUT4AB/EE4END[3]
+ Tile_X5Y8_LUT4AB/EE4END[4] Tile_X5Y8_LUT4AB/EE4END[5] Tile_X5Y8_LUT4AB/EE4END[6]
+ Tile_X5Y8_LUT4AB/EE4END[7] Tile_X5Y8_LUT4AB/EE4END[8] Tile_X5Y8_LUT4AB/EE4END[9]
+ Tile_X5Y8_LUT4AB/FrameData[0] Tile_X5Y8_LUT4AB/FrameData[10] Tile_X5Y8_LUT4AB/FrameData[11]
+ Tile_X5Y8_LUT4AB/FrameData[12] Tile_X5Y8_LUT4AB/FrameData[13] Tile_X5Y8_LUT4AB/FrameData[14]
+ Tile_X5Y8_LUT4AB/FrameData[15] Tile_X5Y8_LUT4AB/FrameData[16] Tile_X5Y8_LUT4AB/FrameData[17]
+ Tile_X5Y8_LUT4AB/FrameData[18] Tile_X5Y8_LUT4AB/FrameData[19] Tile_X5Y8_LUT4AB/FrameData[1]
+ Tile_X5Y8_LUT4AB/FrameData[20] Tile_X5Y8_LUT4AB/FrameData[21] Tile_X5Y8_LUT4AB/FrameData[22]
+ Tile_X5Y8_LUT4AB/FrameData[23] Tile_X5Y8_LUT4AB/FrameData[24] Tile_X5Y8_LUT4AB/FrameData[25]
+ Tile_X5Y8_LUT4AB/FrameData[26] Tile_X5Y8_LUT4AB/FrameData[27] Tile_X5Y8_LUT4AB/FrameData[28]
+ Tile_X5Y8_LUT4AB/FrameData[29] Tile_X5Y8_LUT4AB/FrameData[2] Tile_X5Y8_LUT4AB/FrameData[30]
+ Tile_X5Y8_LUT4AB/FrameData[31] Tile_X5Y8_LUT4AB/FrameData[3] Tile_X5Y8_LUT4AB/FrameData[4]
+ Tile_X5Y8_LUT4AB/FrameData[5] Tile_X5Y8_LUT4AB/FrameData[6] Tile_X5Y8_LUT4AB/FrameData[7]
+ Tile_X5Y8_LUT4AB/FrameData[8] Tile_X5Y8_LUT4AB/FrameData[9] Tile_X6Y8_LUT4AB/FrameData[0]
+ Tile_X6Y8_LUT4AB/FrameData[10] Tile_X6Y8_LUT4AB/FrameData[11] Tile_X6Y8_LUT4AB/FrameData[12]
+ Tile_X6Y8_LUT4AB/FrameData[13] Tile_X6Y8_LUT4AB/FrameData[14] Tile_X6Y8_LUT4AB/FrameData[15]
+ Tile_X6Y8_LUT4AB/FrameData[16] Tile_X6Y8_LUT4AB/FrameData[17] Tile_X6Y8_LUT4AB/FrameData[18]
+ Tile_X6Y8_LUT4AB/FrameData[19] Tile_X6Y8_LUT4AB/FrameData[1] Tile_X6Y8_LUT4AB/FrameData[20]
+ Tile_X6Y8_LUT4AB/FrameData[21] Tile_X6Y8_LUT4AB/FrameData[22] Tile_X6Y8_LUT4AB/FrameData[23]
+ Tile_X6Y8_LUT4AB/FrameData[24] Tile_X6Y8_LUT4AB/FrameData[25] Tile_X6Y8_LUT4AB/FrameData[26]
+ Tile_X6Y8_LUT4AB/FrameData[27] Tile_X6Y8_LUT4AB/FrameData[28] Tile_X6Y8_LUT4AB/FrameData[29]
+ Tile_X6Y8_LUT4AB/FrameData[2] Tile_X6Y8_LUT4AB/FrameData[30] Tile_X6Y8_LUT4AB/FrameData[31]
+ Tile_X6Y8_LUT4AB/FrameData[3] Tile_X6Y8_LUT4AB/FrameData[4] Tile_X6Y8_LUT4AB/FrameData[5]
+ Tile_X6Y8_LUT4AB/FrameData[6] Tile_X6Y8_LUT4AB/FrameData[7] Tile_X6Y8_LUT4AB/FrameData[8]
+ Tile_X6Y8_LUT4AB/FrameData[9] Tile_X5Y8_LUT4AB/FrameStrobe[0] Tile_X5Y8_LUT4AB/FrameStrobe[10]
+ Tile_X5Y8_LUT4AB/FrameStrobe[11] Tile_X5Y8_LUT4AB/FrameStrobe[12] Tile_X5Y8_LUT4AB/FrameStrobe[13]
+ Tile_X5Y8_LUT4AB/FrameStrobe[14] Tile_X5Y8_LUT4AB/FrameStrobe[15] Tile_X5Y8_LUT4AB/FrameStrobe[16]
+ Tile_X5Y8_LUT4AB/FrameStrobe[17] Tile_X5Y8_LUT4AB/FrameStrobe[18] Tile_X5Y8_LUT4AB/FrameStrobe[19]
+ Tile_X5Y8_LUT4AB/FrameStrobe[1] Tile_X5Y8_LUT4AB/FrameStrobe[2] Tile_X5Y8_LUT4AB/FrameStrobe[3]
+ Tile_X5Y8_LUT4AB/FrameStrobe[4] Tile_X5Y8_LUT4AB/FrameStrobe[5] Tile_X5Y8_LUT4AB/FrameStrobe[6]
+ Tile_X5Y8_LUT4AB/FrameStrobe[7] Tile_X5Y8_LUT4AB/FrameStrobe[8] Tile_X5Y8_LUT4AB/FrameStrobe[9]
+ Tile_X5Y7_LUT4AB/FrameStrobe[0] Tile_X5Y7_LUT4AB/FrameStrobe[10] Tile_X5Y7_LUT4AB/FrameStrobe[11]
+ Tile_X5Y7_LUT4AB/FrameStrobe[12] Tile_X5Y7_LUT4AB/FrameStrobe[13] Tile_X5Y7_LUT4AB/FrameStrobe[14]
+ Tile_X5Y7_LUT4AB/FrameStrobe[15] Tile_X5Y7_LUT4AB/FrameStrobe[16] Tile_X5Y7_LUT4AB/FrameStrobe[17]
+ Tile_X5Y7_LUT4AB/FrameStrobe[18] Tile_X5Y7_LUT4AB/FrameStrobe[19] Tile_X5Y7_LUT4AB/FrameStrobe[1]
+ Tile_X5Y7_LUT4AB/FrameStrobe[2] Tile_X5Y7_LUT4AB/FrameStrobe[3] Tile_X5Y7_LUT4AB/FrameStrobe[4]
+ Tile_X5Y7_LUT4AB/FrameStrobe[5] Tile_X5Y7_LUT4AB/FrameStrobe[6] Tile_X5Y7_LUT4AB/FrameStrobe[7]
+ Tile_X5Y7_LUT4AB/FrameStrobe[8] Tile_X5Y7_LUT4AB/FrameStrobe[9] Tile_X5Y8_LUT4AB/N1BEG[0]
+ Tile_X5Y8_LUT4AB/N1BEG[1] Tile_X5Y8_LUT4AB/N1BEG[2] Tile_X5Y8_LUT4AB/N1BEG[3] Tile_X5Y9_LUT4AB/N1BEG[0]
+ Tile_X5Y9_LUT4AB/N1BEG[1] Tile_X5Y9_LUT4AB/N1BEG[2] Tile_X5Y9_LUT4AB/N1BEG[3] Tile_X5Y8_LUT4AB/N2BEG[0]
+ Tile_X5Y8_LUT4AB/N2BEG[1] Tile_X5Y8_LUT4AB/N2BEG[2] Tile_X5Y8_LUT4AB/N2BEG[3] Tile_X5Y8_LUT4AB/N2BEG[4]
+ Tile_X5Y8_LUT4AB/N2BEG[5] Tile_X5Y8_LUT4AB/N2BEG[6] Tile_X5Y8_LUT4AB/N2BEG[7] Tile_X5Y7_LUT4AB/N2END[0]
+ Tile_X5Y7_LUT4AB/N2END[1] Tile_X5Y7_LUT4AB/N2END[2] Tile_X5Y7_LUT4AB/N2END[3] Tile_X5Y7_LUT4AB/N2END[4]
+ Tile_X5Y7_LUT4AB/N2END[5] Tile_X5Y7_LUT4AB/N2END[6] Tile_X5Y7_LUT4AB/N2END[7] Tile_X5Y8_LUT4AB/N2END[0]
+ Tile_X5Y8_LUT4AB/N2END[1] Tile_X5Y8_LUT4AB/N2END[2] Tile_X5Y8_LUT4AB/N2END[3] Tile_X5Y8_LUT4AB/N2END[4]
+ Tile_X5Y8_LUT4AB/N2END[5] Tile_X5Y8_LUT4AB/N2END[6] Tile_X5Y8_LUT4AB/N2END[7] Tile_X5Y9_LUT4AB/N2BEG[0]
+ Tile_X5Y9_LUT4AB/N2BEG[1] Tile_X5Y9_LUT4AB/N2BEG[2] Tile_X5Y9_LUT4AB/N2BEG[3] Tile_X5Y9_LUT4AB/N2BEG[4]
+ Tile_X5Y9_LUT4AB/N2BEG[5] Tile_X5Y9_LUT4AB/N2BEG[6] Tile_X5Y9_LUT4AB/N2BEG[7] Tile_X5Y8_LUT4AB/N4BEG[0]
+ Tile_X5Y8_LUT4AB/N4BEG[10] Tile_X5Y8_LUT4AB/N4BEG[11] Tile_X5Y8_LUT4AB/N4BEG[12]
+ Tile_X5Y8_LUT4AB/N4BEG[13] Tile_X5Y8_LUT4AB/N4BEG[14] Tile_X5Y8_LUT4AB/N4BEG[15]
+ Tile_X5Y8_LUT4AB/N4BEG[1] Tile_X5Y8_LUT4AB/N4BEG[2] Tile_X5Y8_LUT4AB/N4BEG[3] Tile_X5Y8_LUT4AB/N4BEG[4]
+ Tile_X5Y8_LUT4AB/N4BEG[5] Tile_X5Y8_LUT4AB/N4BEG[6] Tile_X5Y8_LUT4AB/N4BEG[7] Tile_X5Y8_LUT4AB/N4BEG[8]
+ Tile_X5Y8_LUT4AB/N4BEG[9] Tile_X5Y9_LUT4AB/N4BEG[0] Tile_X5Y9_LUT4AB/N4BEG[10] Tile_X5Y9_LUT4AB/N4BEG[11]
+ Tile_X5Y9_LUT4AB/N4BEG[12] Tile_X5Y9_LUT4AB/N4BEG[13] Tile_X5Y9_LUT4AB/N4BEG[14]
+ Tile_X5Y9_LUT4AB/N4BEG[15] Tile_X5Y9_LUT4AB/N4BEG[1] Tile_X5Y9_LUT4AB/N4BEG[2] Tile_X5Y9_LUT4AB/N4BEG[3]
+ Tile_X5Y9_LUT4AB/N4BEG[4] Tile_X5Y9_LUT4AB/N4BEG[5] Tile_X5Y9_LUT4AB/N4BEG[6] Tile_X5Y9_LUT4AB/N4BEG[7]
+ Tile_X5Y9_LUT4AB/N4BEG[8] Tile_X5Y9_LUT4AB/N4BEG[9] Tile_X5Y8_LUT4AB/NN4BEG[0] Tile_X5Y8_LUT4AB/NN4BEG[10]
+ Tile_X5Y8_LUT4AB/NN4BEG[11] Tile_X5Y8_LUT4AB/NN4BEG[12] Tile_X5Y8_LUT4AB/NN4BEG[13]
+ Tile_X5Y8_LUT4AB/NN4BEG[14] Tile_X5Y8_LUT4AB/NN4BEG[15] Tile_X5Y8_LUT4AB/NN4BEG[1]
+ Tile_X5Y8_LUT4AB/NN4BEG[2] Tile_X5Y8_LUT4AB/NN4BEG[3] Tile_X5Y8_LUT4AB/NN4BEG[4]
+ Tile_X5Y8_LUT4AB/NN4BEG[5] Tile_X5Y8_LUT4AB/NN4BEG[6] Tile_X5Y8_LUT4AB/NN4BEG[7]
+ Tile_X5Y8_LUT4AB/NN4BEG[8] Tile_X5Y8_LUT4AB/NN4BEG[9] Tile_X5Y9_LUT4AB/NN4BEG[0]
+ Tile_X5Y9_LUT4AB/NN4BEG[10] Tile_X5Y9_LUT4AB/NN4BEG[11] Tile_X5Y9_LUT4AB/NN4BEG[12]
+ Tile_X5Y9_LUT4AB/NN4BEG[13] Tile_X5Y9_LUT4AB/NN4BEG[14] Tile_X5Y9_LUT4AB/NN4BEG[15]
+ Tile_X5Y9_LUT4AB/NN4BEG[1] Tile_X5Y9_LUT4AB/NN4BEG[2] Tile_X5Y9_LUT4AB/NN4BEG[3]
+ Tile_X5Y9_LUT4AB/NN4BEG[4] Tile_X5Y9_LUT4AB/NN4BEG[5] Tile_X5Y9_LUT4AB/NN4BEG[6]
+ Tile_X5Y9_LUT4AB/NN4BEG[7] Tile_X5Y9_LUT4AB/NN4BEG[8] Tile_X5Y9_LUT4AB/NN4BEG[9]
+ Tile_X5Y9_LUT4AB/S1END[0] Tile_X5Y9_LUT4AB/S1END[1] Tile_X5Y9_LUT4AB/S1END[2] Tile_X5Y9_LUT4AB/S1END[3]
+ Tile_X5Y8_LUT4AB/S1END[0] Tile_X5Y8_LUT4AB/S1END[1] Tile_X5Y8_LUT4AB/S1END[2] Tile_X5Y8_LUT4AB/S1END[3]
+ Tile_X5Y9_LUT4AB/S2MID[0] Tile_X5Y9_LUT4AB/S2MID[1] Tile_X5Y9_LUT4AB/S2MID[2] Tile_X5Y9_LUT4AB/S2MID[3]
+ Tile_X5Y9_LUT4AB/S2MID[4] Tile_X5Y9_LUT4AB/S2MID[5] Tile_X5Y9_LUT4AB/S2MID[6] Tile_X5Y9_LUT4AB/S2MID[7]
+ Tile_X5Y9_LUT4AB/S2END[0] Tile_X5Y9_LUT4AB/S2END[1] Tile_X5Y9_LUT4AB/S2END[2] Tile_X5Y9_LUT4AB/S2END[3]
+ Tile_X5Y9_LUT4AB/S2END[4] Tile_X5Y9_LUT4AB/S2END[5] Tile_X5Y9_LUT4AB/S2END[6] Tile_X5Y9_LUT4AB/S2END[7]
+ Tile_X5Y8_LUT4AB/S2END[0] Tile_X5Y8_LUT4AB/S2END[1] Tile_X5Y8_LUT4AB/S2END[2] Tile_X5Y8_LUT4AB/S2END[3]
+ Tile_X5Y8_LUT4AB/S2END[4] Tile_X5Y8_LUT4AB/S2END[5] Tile_X5Y8_LUT4AB/S2END[6] Tile_X5Y8_LUT4AB/S2END[7]
+ Tile_X5Y8_LUT4AB/S2MID[0] Tile_X5Y8_LUT4AB/S2MID[1] Tile_X5Y8_LUT4AB/S2MID[2] Tile_X5Y8_LUT4AB/S2MID[3]
+ Tile_X5Y8_LUT4AB/S2MID[4] Tile_X5Y8_LUT4AB/S2MID[5] Tile_X5Y8_LUT4AB/S2MID[6] Tile_X5Y8_LUT4AB/S2MID[7]
+ Tile_X5Y9_LUT4AB/S4END[0] Tile_X5Y9_LUT4AB/S4END[10] Tile_X5Y9_LUT4AB/S4END[11]
+ Tile_X5Y9_LUT4AB/S4END[12] Tile_X5Y9_LUT4AB/S4END[13] Tile_X5Y9_LUT4AB/S4END[14]
+ Tile_X5Y9_LUT4AB/S4END[15] Tile_X5Y9_LUT4AB/S4END[1] Tile_X5Y9_LUT4AB/S4END[2] Tile_X5Y9_LUT4AB/S4END[3]
+ Tile_X5Y9_LUT4AB/S4END[4] Tile_X5Y9_LUT4AB/S4END[5] Tile_X5Y9_LUT4AB/S4END[6] Tile_X5Y9_LUT4AB/S4END[7]
+ Tile_X5Y9_LUT4AB/S4END[8] Tile_X5Y9_LUT4AB/S4END[9] Tile_X5Y8_LUT4AB/S4END[0] Tile_X5Y8_LUT4AB/S4END[10]
+ Tile_X5Y8_LUT4AB/S4END[11] Tile_X5Y8_LUT4AB/S4END[12] Tile_X5Y8_LUT4AB/S4END[13]
+ Tile_X5Y8_LUT4AB/S4END[14] Tile_X5Y8_LUT4AB/S4END[15] Tile_X5Y8_LUT4AB/S4END[1]
+ Tile_X5Y8_LUT4AB/S4END[2] Tile_X5Y8_LUT4AB/S4END[3] Tile_X5Y8_LUT4AB/S4END[4] Tile_X5Y8_LUT4AB/S4END[5]
+ Tile_X5Y8_LUT4AB/S4END[6] Tile_X5Y8_LUT4AB/S4END[7] Tile_X5Y8_LUT4AB/S4END[8] Tile_X5Y8_LUT4AB/S4END[9]
+ Tile_X5Y9_LUT4AB/SS4END[0] Tile_X5Y9_LUT4AB/SS4END[10] Tile_X5Y9_LUT4AB/SS4END[11]
+ Tile_X5Y9_LUT4AB/SS4END[12] Tile_X5Y9_LUT4AB/SS4END[13] Tile_X5Y9_LUT4AB/SS4END[14]
+ Tile_X5Y9_LUT4AB/SS4END[15] Tile_X5Y9_LUT4AB/SS4END[1] Tile_X5Y9_LUT4AB/SS4END[2]
+ Tile_X5Y9_LUT4AB/SS4END[3] Tile_X5Y9_LUT4AB/SS4END[4] Tile_X5Y9_LUT4AB/SS4END[5]
+ Tile_X5Y9_LUT4AB/SS4END[6] Tile_X5Y9_LUT4AB/SS4END[7] Tile_X5Y9_LUT4AB/SS4END[8]
+ Tile_X5Y9_LUT4AB/SS4END[9] Tile_X5Y8_LUT4AB/SS4END[0] Tile_X5Y8_LUT4AB/SS4END[10]
+ Tile_X5Y8_LUT4AB/SS4END[11] Tile_X5Y8_LUT4AB/SS4END[12] Tile_X5Y8_LUT4AB/SS4END[13]
+ Tile_X5Y8_LUT4AB/SS4END[14] Tile_X5Y8_LUT4AB/SS4END[15] Tile_X5Y8_LUT4AB/SS4END[1]
+ Tile_X5Y8_LUT4AB/SS4END[2] Tile_X5Y8_LUT4AB/SS4END[3] Tile_X5Y8_LUT4AB/SS4END[4]
+ Tile_X5Y8_LUT4AB/SS4END[5] Tile_X5Y8_LUT4AB/SS4END[6] Tile_X5Y8_LUT4AB/SS4END[7]
+ Tile_X5Y8_LUT4AB/SS4END[8] Tile_X5Y8_LUT4AB/SS4END[9] Tile_X5Y8_LUT4AB/UserCLK Tile_X5Y7_LUT4AB/UserCLK
+ VGND VPWR Tile_X5Y8_LUT4AB/W1BEG[0] Tile_X5Y8_LUT4AB/W1BEG[1] Tile_X5Y8_LUT4AB/W1BEG[2]
+ Tile_X5Y8_LUT4AB/W1BEG[3] Tile_X6Y8_LUT4AB/W1BEG[0] Tile_X6Y8_LUT4AB/W1BEG[1] Tile_X6Y8_LUT4AB/W1BEG[2]
+ Tile_X6Y8_LUT4AB/W1BEG[3] Tile_X5Y8_LUT4AB/W2BEG[0] Tile_X5Y8_LUT4AB/W2BEG[1] Tile_X5Y8_LUT4AB/W2BEG[2]
+ Tile_X5Y8_LUT4AB/W2BEG[3] Tile_X5Y8_LUT4AB/W2BEG[4] Tile_X5Y8_LUT4AB/W2BEG[5] Tile_X5Y8_LUT4AB/W2BEG[6]
+ Tile_X5Y8_LUT4AB/W2BEG[7] Tile_X5Y8_LUT4AB/W2BEGb[0] Tile_X5Y8_LUT4AB/W2BEGb[1]
+ Tile_X5Y8_LUT4AB/W2BEGb[2] Tile_X5Y8_LUT4AB/W2BEGb[3] Tile_X5Y8_LUT4AB/W2BEGb[4]
+ Tile_X5Y8_LUT4AB/W2BEGb[5] Tile_X5Y8_LUT4AB/W2BEGb[6] Tile_X5Y8_LUT4AB/W2BEGb[7]
+ Tile_X5Y8_LUT4AB/W2END[0] Tile_X5Y8_LUT4AB/W2END[1] Tile_X5Y8_LUT4AB/W2END[2] Tile_X5Y8_LUT4AB/W2END[3]
+ Tile_X5Y8_LUT4AB/W2END[4] Tile_X5Y8_LUT4AB/W2END[5] Tile_X5Y8_LUT4AB/W2END[6] Tile_X5Y8_LUT4AB/W2END[7]
+ Tile_X6Y8_LUT4AB/W2BEG[0] Tile_X6Y8_LUT4AB/W2BEG[1] Tile_X6Y8_LUT4AB/W2BEG[2] Tile_X6Y8_LUT4AB/W2BEG[3]
+ Tile_X6Y8_LUT4AB/W2BEG[4] Tile_X6Y8_LUT4AB/W2BEG[5] Tile_X6Y8_LUT4AB/W2BEG[6] Tile_X6Y8_LUT4AB/W2BEG[7]
+ Tile_X5Y8_LUT4AB/W6BEG[0] Tile_X5Y8_LUT4AB/W6BEG[10] Tile_X5Y8_LUT4AB/W6BEG[11]
+ Tile_X5Y8_LUT4AB/W6BEG[1] Tile_X5Y8_LUT4AB/W6BEG[2] Tile_X5Y8_LUT4AB/W6BEG[3] Tile_X5Y8_LUT4AB/W6BEG[4]
+ Tile_X5Y8_LUT4AB/W6BEG[5] Tile_X5Y8_LUT4AB/W6BEG[6] Tile_X5Y8_LUT4AB/W6BEG[7] Tile_X5Y8_LUT4AB/W6BEG[8]
+ Tile_X5Y8_LUT4AB/W6BEG[9] Tile_X6Y8_LUT4AB/W6BEG[0] Tile_X6Y8_LUT4AB/W6BEG[10] Tile_X6Y8_LUT4AB/W6BEG[11]
+ Tile_X6Y8_LUT4AB/W6BEG[1] Tile_X6Y8_LUT4AB/W6BEG[2] Tile_X6Y8_LUT4AB/W6BEG[3] Tile_X6Y8_LUT4AB/W6BEG[4]
+ Tile_X6Y8_LUT4AB/W6BEG[5] Tile_X6Y8_LUT4AB/W6BEG[6] Tile_X6Y8_LUT4AB/W6BEG[7] Tile_X6Y8_LUT4AB/W6BEG[8]
+ Tile_X6Y8_LUT4AB/W6BEG[9] Tile_X5Y8_LUT4AB/WW4BEG[0] Tile_X5Y8_LUT4AB/WW4BEG[10]
+ Tile_X5Y8_LUT4AB/WW4BEG[11] Tile_X5Y8_LUT4AB/WW4BEG[12] Tile_X5Y8_LUT4AB/WW4BEG[13]
+ Tile_X5Y8_LUT4AB/WW4BEG[14] Tile_X5Y8_LUT4AB/WW4BEG[15] Tile_X5Y8_LUT4AB/WW4BEG[1]
+ Tile_X5Y8_LUT4AB/WW4BEG[2] Tile_X5Y8_LUT4AB/WW4BEG[3] Tile_X5Y8_LUT4AB/WW4BEG[4]
+ Tile_X5Y8_LUT4AB/WW4BEG[5] Tile_X5Y8_LUT4AB/WW4BEG[6] Tile_X5Y8_LUT4AB/WW4BEG[7]
+ Tile_X5Y8_LUT4AB/WW4BEG[8] Tile_X5Y8_LUT4AB/WW4BEG[9] Tile_X6Y8_LUT4AB/WW4BEG[0]
+ Tile_X6Y8_LUT4AB/WW4BEG[10] Tile_X6Y8_LUT4AB/WW4BEG[11] Tile_X6Y8_LUT4AB/WW4BEG[12]
+ Tile_X6Y8_LUT4AB/WW4BEG[13] Tile_X6Y8_LUT4AB/WW4BEG[14] Tile_X6Y8_LUT4AB/WW4BEG[15]
+ Tile_X6Y8_LUT4AB/WW4BEG[1] Tile_X6Y8_LUT4AB/WW4BEG[2] Tile_X6Y8_LUT4AB/WW4BEG[3]
+ Tile_X6Y8_LUT4AB/WW4BEG[4] Tile_X6Y8_LUT4AB/WW4BEG[5] Tile_X6Y8_LUT4AB/WW4BEG[6]
+ Tile_X6Y8_LUT4AB/WW4BEG[7] Tile_X6Y8_LUT4AB/WW4BEG[8] Tile_X6Y8_LUT4AB/WW4BEG[9]
+ LUT4AB
XTile_X1Y7_LUT4AB Tile_X1Y8_LUT4AB/Co Tile_X1Y7_LUT4AB/Co Tile_X2Y7_LUT4AB/E1END[0]
+ Tile_X2Y7_LUT4AB/E1END[1] Tile_X2Y7_LUT4AB/E1END[2] Tile_X2Y7_LUT4AB/E1END[3] Tile_X0Y7_W_IO/E1BEG[0]
+ Tile_X0Y7_W_IO/E1BEG[1] Tile_X0Y7_W_IO/E1BEG[2] Tile_X0Y7_W_IO/E1BEG[3] Tile_X2Y7_LUT4AB/E2MID[0]
+ Tile_X2Y7_LUT4AB/E2MID[1] Tile_X2Y7_LUT4AB/E2MID[2] Tile_X2Y7_LUT4AB/E2MID[3] Tile_X2Y7_LUT4AB/E2MID[4]
+ Tile_X2Y7_LUT4AB/E2MID[5] Tile_X2Y7_LUT4AB/E2MID[6] Tile_X2Y7_LUT4AB/E2MID[7] Tile_X2Y7_LUT4AB/E2END[0]
+ Tile_X2Y7_LUT4AB/E2END[1] Tile_X2Y7_LUT4AB/E2END[2] Tile_X2Y7_LUT4AB/E2END[3] Tile_X2Y7_LUT4AB/E2END[4]
+ Tile_X2Y7_LUT4AB/E2END[5] Tile_X2Y7_LUT4AB/E2END[6] Tile_X2Y7_LUT4AB/E2END[7] Tile_X0Y7_W_IO/E2BEGb[0]
+ Tile_X0Y7_W_IO/E2BEGb[1] Tile_X0Y7_W_IO/E2BEGb[2] Tile_X0Y7_W_IO/E2BEGb[3] Tile_X0Y7_W_IO/E2BEGb[4]
+ Tile_X0Y7_W_IO/E2BEGb[5] Tile_X0Y7_W_IO/E2BEGb[6] Tile_X0Y7_W_IO/E2BEGb[7] Tile_X0Y7_W_IO/E2BEG[0]
+ Tile_X0Y7_W_IO/E2BEG[1] Tile_X0Y7_W_IO/E2BEG[2] Tile_X0Y7_W_IO/E2BEG[3] Tile_X0Y7_W_IO/E2BEG[4]
+ Tile_X0Y7_W_IO/E2BEG[5] Tile_X0Y7_W_IO/E2BEG[6] Tile_X0Y7_W_IO/E2BEG[7] Tile_X2Y7_LUT4AB/E6END[0]
+ Tile_X2Y7_LUT4AB/E6END[10] Tile_X2Y7_LUT4AB/E6END[11] Tile_X2Y7_LUT4AB/E6END[1]
+ Tile_X2Y7_LUT4AB/E6END[2] Tile_X2Y7_LUT4AB/E6END[3] Tile_X2Y7_LUT4AB/E6END[4] Tile_X2Y7_LUT4AB/E6END[5]
+ Tile_X2Y7_LUT4AB/E6END[6] Tile_X2Y7_LUT4AB/E6END[7] Tile_X2Y7_LUT4AB/E6END[8] Tile_X2Y7_LUT4AB/E6END[9]
+ Tile_X0Y7_W_IO/E6BEG[0] Tile_X0Y7_W_IO/E6BEG[10] Tile_X0Y7_W_IO/E6BEG[11] Tile_X0Y7_W_IO/E6BEG[1]
+ Tile_X0Y7_W_IO/E6BEG[2] Tile_X0Y7_W_IO/E6BEG[3] Tile_X0Y7_W_IO/E6BEG[4] Tile_X0Y7_W_IO/E6BEG[5]
+ Tile_X0Y7_W_IO/E6BEG[6] Tile_X0Y7_W_IO/E6BEG[7] Tile_X0Y7_W_IO/E6BEG[8] Tile_X0Y7_W_IO/E6BEG[9]
+ Tile_X2Y7_LUT4AB/EE4END[0] Tile_X2Y7_LUT4AB/EE4END[10] Tile_X2Y7_LUT4AB/EE4END[11]
+ Tile_X2Y7_LUT4AB/EE4END[12] Tile_X2Y7_LUT4AB/EE4END[13] Tile_X2Y7_LUT4AB/EE4END[14]
+ Tile_X2Y7_LUT4AB/EE4END[15] Tile_X2Y7_LUT4AB/EE4END[1] Tile_X2Y7_LUT4AB/EE4END[2]
+ Tile_X2Y7_LUT4AB/EE4END[3] Tile_X2Y7_LUT4AB/EE4END[4] Tile_X2Y7_LUT4AB/EE4END[5]
+ Tile_X2Y7_LUT4AB/EE4END[6] Tile_X2Y7_LUT4AB/EE4END[7] Tile_X2Y7_LUT4AB/EE4END[8]
+ Tile_X2Y7_LUT4AB/EE4END[9] Tile_X0Y7_W_IO/EE4BEG[0] Tile_X0Y7_W_IO/EE4BEG[10] Tile_X0Y7_W_IO/EE4BEG[11]
+ Tile_X0Y7_W_IO/EE4BEG[12] Tile_X0Y7_W_IO/EE4BEG[13] Tile_X0Y7_W_IO/EE4BEG[14] Tile_X0Y7_W_IO/EE4BEG[15]
+ Tile_X0Y7_W_IO/EE4BEG[1] Tile_X0Y7_W_IO/EE4BEG[2] Tile_X0Y7_W_IO/EE4BEG[3] Tile_X0Y7_W_IO/EE4BEG[4]
+ Tile_X0Y7_W_IO/EE4BEG[5] Tile_X0Y7_W_IO/EE4BEG[6] Tile_X0Y7_W_IO/EE4BEG[7] Tile_X0Y7_W_IO/EE4BEG[8]
+ Tile_X0Y7_W_IO/EE4BEG[9] Tile_X1Y7_LUT4AB/FrameData[0] Tile_X1Y7_LUT4AB/FrameData[10]
+ Tile_X1Y7_LUT4AB/FrameData[11] Tile_X1Y7_LUT4AB/FrameData[12] Tile_X1Y7_LUT4AB/FrameData[13]
+ Tile_X1Y7_LUT4AB/FrameData[14] Tile_X1Y7_LUT4AB/FrameData[15] Tile_X1Y7_LUT4AB/FrameData[16]
+ Tile_X1Y7_LUT4AB/FrameData[17] Tile_X1Y7_LUT4AB/FrameData[18] Tile_X1Y7_LUT4AB/FrameData[19]
+ Tile_X1Y7_LUT4AB/FrameData[1] Tile_X1Y7_LUT4AB/FrameData[20] Tile_X1Y7_LUT4AB/FrameData[21]
+ Tile_X1Y7_LUT4AB/FrameData[22] Tile_X1Y7_LUT4AB/FrameData[23] Tile_X1Y7_LUT4AB/FrameData[24]
+ Tile_X1Y7_LUT4AB/FrameData[25] Tile_X1Y7_LUT4AB/FrameData[26] Tile_X1Y7_LUT4AB/FrameData[27]
+ Tile_X1Y7_LUT4AB/FrameData[28] Tile_X1Y7_LUT4AB/FrameData[29] Tile_X1Y7_LUT4AB/FrameData[2]
+ Tile_X1Y7_LUT4AB/FrameData[30] Tile_X1Y7_LUT4AB/FrameData[31] Tile_X1Y7_LUT4AB/FrameData[3]
+ Tile_X1Y7_LUT4AB/FrameData[4] Tile_X1Y7_LUT4AB/FrameData[5] Tile_X1Y7_LUT4AB/FrameData[6]
+ Tile_X1Y7_LUT4AB/FrameData[7] Tile_X1Y7_LUT4AB/FrameData[8] Tile_X1Y7_LUT4AB/FrameData[9]
+ Tile_X2Y7_LUT4AB/FrameData[0] Tile_X2Y7_LUT4AB/FrameData[10] Tile_X2Y7_LUT4AB/FrameData[11]
+ Tile_X2Y7_LUT4AB/FrameData[12] Tile_X2Y7_LUT4AB/FrameData[13] Tile_X2Y7_LUT4AB/FrameData[14]
+ Tile_X2Y7_LUT4AB/FrameData[15] Tile_X2Y7_LUT4AB/FrameData[16] Tile_X2Y7_LUT4AB/FrameData[17]
+ Tile_X2Y7_LUT4AB/FrameData[18] Tile_X2Y7_LUT4AB/FrameData[19] Tile_X2Y7_LUT4AB/FrameData[1]
+ Tile_X2Y7_LUT4AB/FrameData[20] Tile_X2Y7_LUT4AB/FrameData[21] Tile_X2Y7_LUT4AB/FrameData[22]
+ Tile_X2Y7_LUT4AB/FrameData[23] Tile_X2Y7_LUT4AB/FrameData[24] Tile_X2Y7_LUT4AB/FrameData[25]
+ Tile_X2Y7_LUT4AB/FrameData[26] Tile_X2Y7_LUT4AB/FrameData[27] Tile_X2Y7_LUT4AB/FrameData[28]
+ Tile_X2Y7_LUT4AB/FrameData[29] Tile_X2Y7_LUT4AB/FrameData[2] Tile_X2Y7_LUT4AB/FrameData[30]
+ Tile_X2Y7_LUT4AB/FrameData[31] Tile_X2Y7_LUT4AB/FrameData[3] Tile_X2Y7_LUT4AB/FrameData[4]
+ Tile_X2Y7_LUT4AB/FrameData[5] Tile_X2Y7_LUT4AB/FrameData[6] Tile_X2Y7_LUT4AB/FrameData[7]
+ Tile_X2Y7_LUT4AB/FrameData[8] Tile_X2Y7_LUT4AB/FrameData[9] Tile_X1Y7_LUT4AB/FrameStrobe[0]
+ Tile_X1Y7_LUT4AB/FrameStrobe[10] Tile_X1Y7_LUT4AB/FrameStrobe[11] Tile_X1Y7_LUT4AB/FrameStrobe[12]
+ Tile_X1Y7_LUT4AB/FrameStrobe[13] Tile_X1Y7_LUT4AB/FrameStrobe[14] Tile_X1Y7_LUT4AB/FrameStrobe[15]
+ Tile_X1Y7_LUT4AB/FrameStrobe[16] Tile_X1Y7_LUT4AB/FrameStrobe[17] Tile_X1Y7_LUT4AB/FrameStrobe[18]
+ Tile_X1Y7_LUT4AB/FrameStrobe[19] Tile_X1Y7_LUT4AB/FrameStrobe[1] Tile_X1Y7_LUT4AB/FrameStrobe[2]
+ Tile_X1Y7_LUT4AB/FrameStrobe[3] Tile_X1Y7_LUT4AB/FrameStrobe[4] Tile_X1Y7_LUT4AB/FrameStrobe[5]
+ Tile_X1Y7_LUT4AB/FrameStrobe[6] Tile_X1Y7_LUT4AB/FrameStrobe[7] Tile_X1Y7_LUT4AB/FrameStrobe[8]
+ Tile_X1Y7_LUT4AB/FrameStrobe[9] Tile_X1Y6_LUT4AB/FrameStrobe[0] Tile_X1Y6_LUT4AB/FrameStrobe[10]
+ Tile_X1Y6_LUT4AB/FrameStrobe[11] Tile_X1Y6_LUT4AB/FrameStrobe[12] Tile_X1Y6_LUT4AB/FrameStrobe[13]
+ Tile_X1Y6_LUT4AB/FrameStrobe[14] Tile_X1Y6_LUT4AB/FrameStrobe[15] Tile_X1Y6_LUT4AB/FrameStrobe[16]
+ Tile_X1Y6_LUT4AB/FrameStrobe[17] Tile_X1Y6_LUT4AB/FrameStrobe[18] Tile_X1Y6_LUT4AB/FrameStrobe[19]
+ Tile_X1Y6_LUT4AB/FrameStrobe[1] Tile_X1Y6_LUT4AB/FrameStrobe[2] Tile_X1Y6_LUT4AB/FrameStrobe[3]
+ Tile_X1Y6_LUT4AB/FrameStrobe[4] Tile_X1Y6_LUT4AB/FrameStrobe[5] Tile_X1Y6_LUT4AB/FrameStrobe[6]
+ Tile_X1Y6_LUT4AB/FrameStrobe[7] Tile_X1Y6_LUT4AB/FrameStrobe[8] Tile_X1Y6_LUT4AB/FrameStrobe[9]
+ Tile_X1Y7_LUT4AB/N1BEG[0] Tile_X1Y7_LUT4AB/N1BEG[1] Tile_X1Y7_LUT4AB/N1BEG[2] Tile_X1Y7_LUT4AB/N1BEG[3]
+ Tile_X1Y8_LUT4AB/N1BEG[0] Tile_X1Y8_LUT4AB/N1BEG[1] Tile_X1Y8_LUT4AB/N1BEG[2] Tile_X1Y8_LUT4AB/N1BEG[3]
+ Tile_X1Y7_LUT4AB/N2BEG[0] Tile_X1Y7_LUT4AB/N2BEG[1] Tile_X1Y7_LUT4AB/N2BEG[2] Tile_X1Y7_LUT4AB/N2BEG[3]
+ Tile_X1Y7_LUT4AB/N2BEG[4] Tile_X1Y7_LUT4AB/N2BEG[5] Tile_X1Y7_LUT4AB/N2BEG[6] Tile_X1Y7_LUT4AB/N2BEG[7]
+ Tile_X1Y6_LUT4AB/N2END[0] Tile_X1Y6_LUT4AB/N2END[1] Tile_X1Y6_LUT4AB/N2END[2] Tile_X1Y6_LUT4AB/N2END[3]
+ Tile_X1Y6_LUT4AB/N2END[4] Tile_X1Y6_LUT4AB/N2END[5] Tile_X1Y6_LUT4AB/N2END[6] Tile_X1Y6_LUT4AB/N2END[7]
+ Tile_X1Y7_LUT4AB/N2END[0] Tile_X1Y7_LUT4AB/N2END[1] Tile_X1Y7_LUT4AB/N2END[2] Tile_X1Y7_LUT4AB/N2END[3]
+ Tile_X1Y7_LUT4AB/N2END[4] Tile_X1Y7_LUT4AB/N2END[5] Tile_X1Y7_LUT4AB/N2END[6] Tile_X1Y7_LUT4AB/N2END[7]
+ Tile_X1Y8_LUT4AB/N2BEG[0] Tile_X1Y8_LUT4AB/N2BEG[1] Tile_X1Y8_LUT4AB/N2BEG[2] Tile_X1Y8_LUT4AB/N2BEG[3]
+ Tile_X1Y8_LUT4AB/N2BEG[4] Tile_X1Y8_LUT4AB/N2BEG[5] Tile_X1Y8_LUT4AB/N2BEG[6] Tile_X1Y8_LUT4AB/N2BEG[7]
+ Tile_X1Y7_LUT4AB/N4BEG[0] Tile_X1Y7_LUT4AB/N4BEG[10] Tile_X1Y7_LUT4AB/N4BEG[11]
+ Tile_X1Y7_LUT4AB/N4BEG[12] Tile_X1Y7_LUT4AB/N4BEG[13] Tile_X1Y7_LUT4AB/N4BEG[14]
+ Tile_X1Y7_LUT4AB/N4BEG[15] Tile_X1Y7_LUT4AB/N4BEG[1] Tile_X1Y7_LUT4AB/N4BEG[2] Tile_X1Y7_LUT4AB/N4BEG[3]
+ Tile_X1Y7_LUT4AB/N4BEG[4] Tile_X1Y7_LUT4AB/N4BEG[5] Tile_X1Y7_LUT4AB/N4BEG[6] Tile_X1Y7_LUT4AB/N4BEG[7]
+ Tile_X1Y7_LUT4AB/N4BEG[8] Tile_X1Y7_LUT4AB/N4BEG[9] Tile_X1Y8_LUT4AB/N4BEG[0] Tile_X1Y8_LUT4AB/N4BEG[10]
+ Tile_X1Y8_LUT4AB/N4BEG[11] Tile_X1Y8_LUT4AB/N4BEG[12] Tile_X1Y8_LUT4AB/N4BEG[13]
+ Tile_X1Y8_LUT4AB/N4BEG[14] Tile_X1Y8_LUT4AB/N4BEG[15] Tile_X1Y8_LUT4AB/N4BEG[1]
+ Tile_X1Y8_LUT4AB/N4BEG[2] Tile_X1Y8_LUT4AB/N4BEG[3] Tile_X1Y8_LUT4AB/N4BEG[4] Tile_X1Y8_LUT4AB/N4BEG[5]
+ Tile_X1Y8_LUT4AB/N4BEG[6] Tile_X1Y8_LUT4AB/N4BEG[7] Tile_X1Y8_LUT4AB/N4BEG[8] Tile_X1Y8_LUT4AB/N4BEG[9]
+ Tile_X1Y7_LUT4AB/NN4BEG[0] Tile_X1Y7_LUT4AB/NN4BEG[10] Tile_X1Y7_LUT4AB/NN4BEG[11]
+ Tile_X1Y7_LUT4AB/NN4BEG[12] Tile_X1Y7_LUT4AB/NN4BEG[13] Tile_X1Y7_LUT4AB/NN4BEG[14]
+ Tile_X1Y7_LUT4AB/NN4BEG[15] Tile_X1Y7_LUT4AB/NN4BEG[1] Tile_X1Y7_LUT4AB/NN4BEG[2]
+ Tile_X1Y7_LUT4AB/NN4BEG[3] Tile_X1Y7_LUT4AB/NN4BEG[4] Tile_X1Y7_LUT4AB/NN4BEG[5]
+ Tile_X1Y7_LUT4AB/NN4BEG[6] Tile_X1Y7_LUT4AB/NN4BEG[7] Tile_X1Y7_LUT4AB/NN4BEG[8]
+ Tile_X1Y7_LUT4AB/NN4BEG[9] Tile_X1Y8_LUT4AB/NN4BEG[0] Tile_X1Y8_LUT4AB/NN4BEG[10]
+ Tile_X1Y8_LUT4AB/NN4BEG[11] Tile_X1Y8_LUT4AB/NN4BEG[12] Tile_X1Y8_LUT4AB/NN4BEG[13]
+ Tile_X1Y8_LUT4AB/NN4BEG[14] Tile_X1Y8_LUT4AB/NN4BEG[15] Tile_X1Y8_LUT4AB/NN4BEG[1]
+ Tile_X1Y8_LUT4AB/NN4BEG[2] Tile_X1Y8_LUT4AB/NN4BEG[3] Tile_X1Y8_LUT4AB/NN4BEG[4]
+ Tile_X1Y8_LUT4AB/NN4BEG[5] Tile_X1Y8_LUT4AB/NN4BEG[6] Tile_X1Y8_LUT4AB/NN4BEG[7]
+ Tile_X1Y8_LUT4AB/NN4BEG[8] Tile_X1Y8_LUT4AB/NN4BEG[9] Tile_X1Y8_LUT4AB/S1END[0]
+ Tile_X1Y8_LUT4AB/S1END[1] Tile_X1Y8_LUT4AB/S1END[2] Tile_X1Y8_LUT4AB/S1END[3] Tile_X1Y7_LUT4AB/S1END[0]
+ Tile_X1Y7_LUT4AB/S1END[1] Tile_X1Y7_LUT4AB/S1END[2] Tile_X1Y7_LUT4AB/S1END[3] Tile_X1Y8_LUT4AB/S2MID[0]
+ Tile_X1Y8_LUT4AB/S2MID[1] Tile_X1Y8_LUT4AB/S2MID[2] Tile_X1Y8_LUT4AB/S2MID[3] Tile_X1Y8_LUT4AB/S2MID[4]
+ Tile_X1Y8_LUT4AB/S2MID[5] Tile_X1Y8_LUT4AB/S2MID[6] Tile_X1Y8_LUT4AB/S2MID[7] Tile_X1Y8_LUT4AB/S2END[0]
+ Tile_X1Y8_LUT4AB/S2END[1] Tile_X1Y8_LUT4AB/S2END[2] Tile_X1Y8_LUT4AB/S2END[3] Tile_X1Y8_LUT4AB/S2END[4]
+ Tile_X1Y8_LUT4AB/S2END[5] Tile_X1Y8_LUT4AB/S2END[6] Tile_X1Y8_LUT4AB/S2END[7] Tile_X1Y7_LUT4AB/S2END[0]
+ Tile_X1Y7_LUT4AB/S2END[1] Tile_X1Y7_LUT4AB/S2END[2] Tile_X1Y7_LUT4AB/S2END[3] Tile_X1Y7_LUT4AB/S2END[4]
+ Tile_X1Y7_LUT4AB/S2END[5] Tile_X1Y7_LUT4AB/S2END[6] Tile_X1Y7_LUT4AB/S2END[7] Tile_X1Y7_LUT4AB/S2MID[0]
+ Tile_X1Y7_LUT4AB/S2MID[1] Tile_X1Y7_LUT4AB/S2MID[2] Tile_X1Y7_LUT4AB/S2MID[3] Tile_X1Y7_LUT4AB/S2MID[4]
+ Tile_X1Y7_LUT4AB/S2MID[5] Tile_X1Y7_LUT4AB/S2MID[6] Tile_X1Y7_LUT4AB/S2MID[7] Tile_X1Y8_LUT4AB/S4END[0]
+ Tile_X1Y8_LUT4AB/S4END[10] Tile_X1Y8_LUT4AB/S4END[11] Tile_X1Y8_LUT4AB/S4END[12]
+ Tile_X1Y8_LUT4AB/S4END[13] Tile_X1Y8_LUT4AB/S4END[14] Tile_X1Y8_LUT4AB/S4END[15]
+ Tile_X1Y8_LUT4AB/S4END[1] Tile_X1Y8_LUT4AB/S4END[2] Tile_X1Y8_LUT4AB/S4END[3] Tile_X1Y8_LUT4AB/S4END[4]
+ Tile_X1Y8_LUT4AB/S4END[5] Tile_X1Y8_LUT4AB/S4END[6] Tile_X1Y8_LUT4AB/S4END[7] Tile_X1Y8_LUT4AB/S4END[8]
+ Tile_X1Y8_LUT4AB/S4END[9] Tile_X1Y7_LUT4AB/S4END[0] Tile_X1Y7_LUT4AB/S4END[10] Tile_X1Y7_LUT4AB/S4END[11]
+ Tile_X1Y7_LUT4AB/S4END[12] Tile_X1Y7_LUT4AB/S4END[13] Tile_X1Y7_LUT4AB/S4END[14]
+ Tile_X1Y7_LUT4AB/S4END[15] Tile_X1Y7_LUT4AB/S4END[1] Tile_X1Y7_LUT4AB/S4END[2] Tile_X1Y7_LUT4AB/S4END[3]
+ Tile_X1Y7_LUT4AB/S4END[4] Tile_X1Y7_LUT4AB/S4END[5] Tile_X1Y7_LUT4AB/S4END[6] Tile_X1Y7_LUT4AB/S4END[7]
+ Tile_X1Y7_LUT4AB/S4END[8] Tile_X1Y7_LUT4AB/S4END[9] Tile_X1Y8_LUT4AB/SS4END[0] Tile_X1Y8_LUT4AB/SS4END[10]
+ Tile_X1Y8_LUT4AB/SS4END[11] Tile_X1Y8_LUT4AB/SS4END[12] Tile_X1Y8_LUT4AB/SS4END[13]
+ Tile_X1Y8_LUT4AB/SS4END[14] Tile_X1Y8_LUT4AB/SS4END[15] Tile_X1Y8_LUT4AB/SS4END[1]
+ Tile_X1Y8_LUT4AB/SS4END[2] Tile_X1Y8_LUT4AB/SS4END[3] Tile_X1Y8_LUT4AB/SS4END[4]
+ Tile_X1Y8_LUT4AB/SS4END[5] Tile_X1Y8_LUT4AB/SS4END[6] Tile_X1Y8_LUT4AB/SS4END[7]
+ Tile_X1Y8_LUT4AB/SS4END[8] Tile_X1Y8_LUT4AB/SS4END[9] Tile_X1Y7_LUT4AB/SS4END[0]
+ Tile_X1Y7_LUT4AB/SS4END[10] Tile_X1Y7_LUT4AB/SS4END[11] Tile_X1Y7_LUT4AB/SS4END[12]
+ Tile_X1Y7_LUT4AB/SS4END[13] Tile_X1Y7_LUT4AB/SS4END[14] Tile_X1Y7_LUT4AB/SS4END[15]
+ Tile_X1Y7_LUT4AB/SS4END[1] Tile_X1Y7_LUT4AB/SS4END[2] Tile_X1Y7_LUT4AB/SS4END[3]
+ Tile_X1Y7_LUT4AB/SS4END[4] Tile_X1Y7_LUT4AB/SS4END[5] Tile_X1Y7_LUT4AB/SS4END[6]
+ Tile_X1Y7_LUT4AB/SS4END[7] Tile_X1Y7_LUT4AB/SS4END[8] Tile_X1Y7_LUT4AB/SS4END[9]
+ Tile_X1Y7_LUT4AB/UserCLK Tile_X1Y6_LUT4AB/UserCLK VGND VPWR Tile_X0Y7_W_IO/W1END[0]
+ Tile_X0Y7_W_IO/W1END[1] Tile_X0Y7_W_IO/W1END[2] Tile_X0Y7_W_IO/W1END[3] Tile_X2Y7_LUT4AB/W1BEG[0]
+ Tile_X2Y7_LUT4AB/W1BEG[1] Tile_X2Y7_LUT4AB/W1BEG[2] Tile_X2Y7_LUT4AB/W1BEG[3] Tile_X0Y7_W_IO/W2MID[0]
+ Tile_X0Y7_W_IO/W2MID[1] Tile_X0Y7_W_IO/W2MID[2] Tile_X0Y7_W_IO/W2MID[3] Tile_X0Y7_W_IO/W2MID[4]
+ Tile_X0Y7_W_IO/W2MID[5] Tile_X0Y7_W_IO/W2MID[6] Tile_X0Y7_W_IO/W2MID[7] Tile_X0Y7_W_IO/W2END[0]
+ Tile_X0Y7_W_IO/W2END[1] Tile_X0Y7_W_IO/W2END[2] Tile_X0Y7_W_IO/W2END[3] Tile_X0Y7_W_IO/W2END[4]
+ Tile_X0Y7_W_IO/W2END[5] Tile_X0Y7_W_IO/W2END[6] Tile_X0Y7_W_IO/W2END[7] Tile_X1Y7_LUT4AB/W2END[0]
+ Tile_X1Y7_LUT4AB/W2END[1] Tile_X1Y7_LUT4AB/W2END[2] Tile_X1Y7_LUT4AB/W2END[3] Tile_X1Y7_LUT4AB/W2END[4]
+ Tile_X1Y7_LUT4AB/W2END[5] Tile_X1Y7_LUT4AB/W2END[6] Tile_X1Y7_LUT4AB/W2END[7] Tile_X2Y7_LUT4AB/W2BEG[0]
+ Tile_X2Y7_LUT4AB/W2BEG[1] Tile_X2Y7_LUT4AB/W2BEG[2] Tile_X2Y7_LUT4AB/W2BEG[3] Tile_X2Y7_LUT4AB/W2BEG[4]
+ Tile_X2Y7_LUT4AB/W2BEG[5] Tile_X2Y7_LUT4AB/W2BEG[6] Tile_X2Y7_LUT4AB/W2BEG[7] Tile_X0Y7_W_IO/W6END[0]
+ Tile_X0Y7_W_IO/W6END[10] Tile_X0Y7_W_IO/W6END[11] Tile_X0Y7_W_IO/W6END[1] Tile_X0Y7_W_IO/W6END[2]
+ Tile_X0Y7_W_IO/W6END[3] Tile_X0Y7_W_IO/W6END[4] Tile_X0Y7_W_IO/W6END[5] Tile_X0Y7_W_IO/W6END[6]
+ Tile_X0Y7_W_IO/W6END[7] Tile_X0Y7_W_IO/W6END[8] Tile_X0Y7_W_IO/W6END[9] Tile_X2Y7_LUT4AB/W6BEG[0]
+ Tile_X2Y7_LUT4AB/W6BEG[10] Tile_X2Y7_LUT4AB/W6BEG[11] Tile_X2Y7_LUT4AB/W6BEG[1]
+ Tile_X2Y7_LUT4AB/W6BEG[2] Tile_X2Y7_LUT4AB/W6BEG[3] Tile_X2Y7_LUT4AB/W6BEG[4] Tile_X2Y7_LUT4AB/W6BEG[5]
+ Tile_X2Y7_LUT4AB/W6BEG[6] Tile_X2Y7_LUT4AB/W6BEG[7] Tile_X2Y7_LUT4AB/W6BEG[8] Tile_X2Y7_LUT4AB/W6BEG[9]
+ Tile_X0Y7_W_IO/WW4END[0] Tile_X0Y7_W_IO/WW4END[10] Tile_X0Y7_W_IO/WW4END[11] Tile_X0Y7_W_IO/WW4END[12]
+ Tile_X0Y7_W_IO/WW4END[13] Tile_X0Y7_W_IO/WW4END[14] Tile_X0Y7_W_IO/WW4END[15] Tile_X0Y7_W_IO/WW4END[1]
+ Tile_X0Y7_W_IO/WW4END[2] Tile_X0Y7_W_IO/WW4END[3] Tile_X0Y7_W_IO/WW4END[4] Tile_X0Y7_W_IO/WW4END[5]
+ Tile_X0Y7_W_IO/WW4END[6] Tile_X0Y7_W_IO/WW4END[7] Tile_X0Y7_W_IO/WW4END[8] Tile_X0Y7_W_IO/WW4END[9]
+ Tile_X2Y7_LUT4AB/WW4BEG[0] Tile_X2Y7_LUT4AB/WW4BEG[10] Tile_X2Y7_LUT4AB/WW4BEG[11]
+ Tile_X2Y7_LUT4AB/WW4BEG[12] Tile_X2Y7_LUT4AB/WW4BEG[13] Tile_X2Y7_LUT4AB/WW4BEG[14]
+ Tile_X2Y7_LUT4AB/WW4BEG[15] Tile_X2Y7_LUT4AB/WW4BEG[1] Tile_X2Y7_LUT4AB/WW4BEG[2]
+ Tile_X2Y7_LUT4AB/WW4BEG[3] Tile_X2Y7_LUT4AB/WW4BEG[4] Tile_X2Y7_LUT4AB/WW4BEG[5]
+ Tile_X2Y7_LUT4AB/WW4BEG[6] Tile_X2Y7_LUT4AB/WW4BEG[7] Tile_X2Y7_LUT4AB/WW4BEG[8]
+ Tile_X2Y7_LUT4AB/WW4BEG[9] LUT4AB
XTile_X4Y11_RegFile Tile_X5Y11_LUT4AB/E1END[0] Tile_X5Y11_LUT4AB/E1END[1] Tile_X5Y11_LUT4AB/E1END[2]
+ Tile_X5Y11_LUT4AB/E1END[3] Tile_X3Y11_LUT4AB/E1BEG[0] Tile_X3Y11_LUT4AB/E1BEG[1]
+ Tile_X3Y11_LUT4AB/E1BEG[2] Tile_X3Y11_LUT4AB/E1BEG[3] Tile_X5Y11_LUT4AB/E2MID[0]
+ Tile_X5Y11_LUT4AB/E2MID[1] Tile_X5Y11_LUT4AB/E2MID[2] Tile_X5Y11_LUT4AB/E2MID[3]
+ Tile_X5Y11_LUT4AB/E2MID[4] Tile_X5Y11_LUT4AB/E2MID[5] Tile_X5Y11_LUT4AB/E2MID[6]
+ Tile_X5Y11_LUT4AB/E2MID[7] Tile_X5Y11_LUT4AB/E2END[0] Tile_X5Y11_LUT4AB/E2END[1]
+ Tile_X5Y11_LUT4AB/E2END[2] Tile_X5Y11_LUT4AB/E2END[3] Tile_X5Y11_LUT4AB/E2END[4]
+ Tile_X5Y11_LUT4AB/E2END[5] Tile_X5Y11_LUT4AB/E2END[6] Tile_X5Y11_LUT4AB/E2END[7]
+ Tile_X4Y11_RegFile/E2END[0] Tile_X4Y11_RegFile/E2END[1] Tile_X4Y11_RegFile/E2END[2]
+ Tile_X4Y11_RegFile/E2END[3] Tile_X4Y11_RegFile/E2END[4] Tile_X4Y11_RegFile/E2END[5]
+ Tile_X4Y11_RegFile/E2END[6] Tile_X4Y11_RegFile/E2END[7] Tile_X3Y11_LUT4AB/E2BEG[0]
+ Tile_X3Y11_LUT4AB/E2BEG[1] Tile_X3Y11_LUT4AB/E2BEG[2] Tile_X3Y11_LUT4AB/E2BEG[3]
+ Tile_X3Y11_LUT4AB/E2BEG[4] Tile_X3Y11_LUT4AB/E2BEG[5] Tile_X3Y11_LUT4AB/E2BEG[6]
+ Tile_X3Y11_LUT4AB/E2BEG[7] Tile_X5Y11_LUT4AB/E6END[0] Tile_X5Y11_LUT4AB/E6END[10]
+ Tile_X5Y11_LUT4AB/E6END[11] Tile_X5Y11_LUT4AB/E6END[1] Tile_X5Y11_LUT4AB/E6END[2]
+ Tile_X5Y11_LUT4AB/E6END[3] Tile_X5Y11_LUT4AB/E6END[4] Tile_X5Y11_LUT4AB/E6END[5]
+ Tile_X5Y11_LUT4AB/E6END[6] Tile_X5Y11_LUT4AB/E6END[7] Tile_X5Y11_LUT4AB/E6END[8]
+ Tile_X5Y11_LUT4AB/E6END[9] Tile_X3Y11_LUT4AB/E6BEG[0] Tile_X3Y11_LUT4AB/E6BEG[10]
+ Tile_X3Y11_LUT4AB/E6BEG[11] Tile_X3Y11_LUT4AB/E6BEG[1] Tile_X3Y11_LUT4AB/E6BEG[2]
+ Tile_X3Y11_LUT4AB/E6BEG[3] Tile_X3Y11_LUT4AB/E6BEG[4] Tile_X3Y11_LUT4AB/E6BEG[5]
+ Tile_X3Y11_LUT4AB/E6BEG[6] Tile_X3Y11_LUT4AB/E6BEG[7] Tile_X3Y11_LUT4AB/E6BEG[8]
+ Tile_X3Y11_LUT4AB/E6BEG[9] Tile_X5Y11_LUT4AB/EE4END[0] Tile_X5Y11_LUT4AB/EE4END[10]
+ Tile_X5Y11_LUT4AB/EE4END[11] Tile_X5Y11_LUT4AB/EE4END[12] Tile_X5Y11_LUT4AB/EE4END[13]
+ Tile_X5Y11_LUT4AB/EE4END[14] Tile_X5Y11_LUT4AB/EE4END[15] Tile_X5Y11_LUT4AB/EE4END[1]
+ Tile_X5Y11_LUT4AB/EE4END[2] Tile_X5Y11_LUT4AB/EE4END[3] Tile_X5Y11_LUT4AB/EE4END[4]
+ Tile_X5Y11_LUT4AB/EE4END[5] Tile_X5Y11_LUT4AB/EE4END[6] Tile_X5Y11_LUT4AB/EE4END[7]
+ Tile_X5Y11_LUT4AB/EE4END[8] Tile_X5Y11_LUT4AB/EE4END[9] Tile_X3Y11_LUT4AB/EE4BEG[0]
+ Tile_X3Y11_LUT4AB/EE4BEG[10] Tile_X3Y11_LUT4AB/EE4BEG[11] Tile_X3Y11_LUT4AB/EE4BEG[12]
+ Tile_X3Y11_LUT4AB/EE4BEG[13] Tile_X3Y11_LUT4AB/EE4BEG[14] Tile_X3Y11_LUT4AB/EE4BEG[15]
+ Tile_X3Y11_LUT4AB/EE4BEG[1] Tile_X3Y11_LUT4AB/EE4BEG[2] Tile_X3Y11_LUT4AB/EE4BEG[3]
+ Tile_X3Y11_LUT4AB/EE4BEG[4] Tile_X3Y11_LUT4AB/EE4BEG[5] Tile_X3Y11_LUT4AB/EE4BEG[6]
+ Tile_X3Y11_LUT4AB/EE4BEG[7] Tile_X3Y11_LUT4AB/EE4BEG[8] Tile_X3Y11_LUT4AB/EE4BEG[9]
+ Tile_X4Y11_RegFile/FrameData[0] Tile_X4Y11_RegFile/FrameData[10] Tile_X4Y11_RegFile/FrameData[11]
+ Tile_X4Y11_RegFile/FrameData[12] Tile_X4Y11_RegFile/FrameData[13] Tile_X4Y11_RegFile/FrameData[14]
+ Tile_X4Y11_RegFile/FrameData[15] Tile_X4Y11_RegFile/FrameData[16] Tile_X4Y11_RegFile/FrameData[17]
+ Tile_X4Y11_RegFile/FrameData[18] Tile_X4Y11_RegFile/FrameData[19] Tile_X4Y11_RegFile/FrameData[1]
+ Tile_X4Y11_RegFile/FrameData[20] Tile_X4Y11_RegFile/FrameData[21] Tile_X4Y11_RegFile/FrameData[22]
+ Tile_X4Y11_RegFile/FrameData[23] Tile_X4Y11_RegFile/FrameData[24] Tile_X4Y11_RegFile/FrameData[25]
+ Tile_X4Y11_RegFile/FrameData[26] Tile_X4Y11_RegFile/FrameData[27] Tile_X4Y11_RegFile/FrameData[28]
+ Tile_X4Y11_RegFile/FrameData[29] Tile_X4Y11_RegFile/FrameData[2] Tile_X4Y11_RegFile/FrameData[30]
+ Tile_X4Y11_RegFile/FrameData[31] Tile_X4Y11_RegFile/FrameData[3] Tile_X4Y11_RegFile/FrameData[4]
+ Tile_X4Y11_RegFile/FrameData[5] Tile_X4Y11_RegFile/FrameData[6] Tile_X4Y11_RegFile/FrameData[7]
+ Tile_X4Y11_RegFile/FrameData[8] Tile_X4Y11_RegFile/FrameData[9] Tile_X5Y11_LUT4AB/FrameData[0]
+ Tile_X5Y11_LUT4AB/FrameData[10] Tile_X5Y11_LUT4AB/FrameData[11] Tile_X5Y11_LUT4AB/FrameData[12]
+ Tile_X5Y11_LUT4AB/FrameData[13] Tile_X5Y11_LUT4AB/FrameData[14] Tile_X5Y11_LUT4AB/FrameData[15]
+ Tile_X5Y11_LUT4AB/FrameData[16] Tile_X5Y11_LUT4AB/FrameData[17] Tile_X5Y11_LUT4AB/FrameData[18]
+ Tile_X5Y11_LUT4AB/FrameData[19] Tile_X5Y11_LUT4AB/FrameData[1] Tile_X5Y11_LUT4AB/FrameData[20]
+ Tile_X5Y11_LUT4AB/FrameData[21] Tile_X5Y11_LUT4AB/FrameData[22] Tile_X5Y11_LUT4AB/FrameData[23]
+ Tile_X5Y11_LUT4AB/FrameData[24] Tile_X5Y11_LUT4AB/FrameData[25] Tile_X5Y11_LUT4AB/FrameData[26]
+ Tile_X5Y11_LUT4AB/FrameData[27] Tile_X5Y11_LUT4AB/FrameData[28] Tile_X5Y11_LUT4AB/FrameData[29]
+ Tile_X5Y11_LUT4AB/FrameData[2] Tile_X5Y11_LUT4AB/FrameData[30] Tile_X5Y11_LUT4AB/FrameData[31]
+ Tile_X5Y11_LUT4AB/FrameData[3] Tile_X5Y11_LUT4AB/FrameData[4] Tile_X5Y11_LUT4AB/FrameData[5]
+ Tile_X5Y11_LUT4AB/FrameData[6] Tile_X5Y11_LUT4AB/FrameData[7] Tile_X5Y11_LUT4AB/FrameData[8]
+ Tile_X5Y11_LUT4AB/FrameData[9] Tile_X4Y11_RegFile/FrameStrobe[0] Tile_X4Y11_RegFile/FrameStrobe[10]
+ Tile_X4Y11_RegFile/FrameStrobe[11] Tile_X4Y11_RegFile/FrameStrobe[12] Tile_X4Y11_RegFile/FrameStrobe[13]
+ Tile_X4Y11_RegFile/FrameStrobe[14] Tile_X4Y11_RegFile/FrameStrobe[15] Tile_X4Y11_RegFile/FrameStrobe[16]
+ Tile_X4Y11_RegFile/FrameStrobe[17] Tile_X4Y11_RegFile/FrameStrobe[18] Tile_X4Y11_RegFile/FrameStrobe[19]
+ Tile_X4Y11_RegFile/FrameStrobe[1] Tile_X4Y11_RegFile/FrameStrobe[2] Tile_X4Y11_RegFile/FrameStrobe[3]
+ Tile_X4Y11_RegFile/FrameStrobe[4] Tile_X4Y11_RegFile/FrameStrobe[5] Tile_X4Y11_RegFile/FrameStrobe[6]
+ Tile_X4Y11_RegFile/FrameStrobe[7] Tile_X4Y11_RegFile/FrameStrobe[8] Tile_X4Y11_RegFile/FrameStrobe[9]
+ Tile_X4Y10_RegFile/FrameStrobe[0] Tile_X4Y10_RegFile/FrameStrobe[10] Tile_X4Y10_RegFile/FrameStrobe[11]
+ Tile_X4Y10_RegFile/FrameStrobe[12] Tile_X4Y10_RegFile/FrameStrobe[13] Tile_X4Y10_RegFile/FrameStrobe[14]
+ Tile_X4Y10_RegFile/FrameStrobe[15] Tile_X4Y10_RegFile/FrameStrobe[16] Tile_X4Y10_RegFile/FrameStrobe[17]
+ Tile_X4Y10_RegFile/FrameStrobe[18] Tile_X4Y10_RegFile/FrameStrobe[19] Tile_X4Y10_RegFile/FrameStrobe[1]
+ Tile_X4Y10_RegFile/FrameStrobe[2] Tile_X4Y10_RegFile/FrameStrobe[3] Tile_X4Y10_RegFile/FrameStrobe[4]
+ Tile_X4Y10_RegFile/FrameStrobe[5] Tile_X4Y10_RegFile/FrameStrobe[6] Tile_X4Y10_RegFile/FrameStrobe[7]
+ Tile_X4Y10_RegFile/FrameStrobe[8] Tile_X4Y10_RegFile/FrameStrobe[9] Tile_X4Y11_RegFile/N1BEG[0]
+ Tile_X4Y11_RegFile/N1BEG[1] Tile_X4Y11_RegFile/N1BEG[2] Tile_X4Y11_RegFile/N1BEG[3]
+ Tile_X4Y12_RegFile/N1BEG[0] Tile_X4Y12_RegFile/N1BEG[1] Tile_X4Y12_RegFile/N1BEG[2]
+ Tile_X4Y12_RegFile/N1BEG[3] Tile_X4Y11_RegFile/N2BEG[0] Tile_X4Y11_RegFile/N2BEG[1]
+ Tile_X4Y11_RegFile/N2BEG[2] Tile_X4Y11_RegFile/N2BEG[3] Tile_X4Y11_RegFile/N2BEG[4]
+ Tile_X4Y11_RegFile/N2BEG[5] Tile_X4Y11_RegFile/N2BEG[6] Tile_X4Y11_RegFile/N2BEG[7]
+ Tile_X4Y10_RegFile/N2END[0] Tile_X4Y10_RegFile/N2END[1] Tile_X4Y10_RegFile/N2END[2]
+ Tile_X4Y10_RegFile/N2END[3] Tile_X4Y10_RegFile/N2END[4] Tile_X4Y10_RegFile/N2END[5]
+ Tile_X4Y10_RegFile/N2END[6] Tile_X4Y10_RegFile/N2END[7] Tile_X4Y11_RegFile/N2END[0]
+ Tile_X4Y11_RegFile/N2END[1] Tile_X4Y11_RegFile/N2END[2] Tile_X4Y11_RegFile/N2END[3]
+ Tile_X4Y11_RegFile/N2END[4] Tile_X4Y11_RegFile/N2END[5] Tile_X4Y11_RegFile/N2END[6]
+ Tile_X4Y11_RegFile/N2END[7] Tile_X4Y12_RegFile/N2BEG[0] Tile_X4Y12_RegFile/N2BEG[1]
+ Tile_X4Y12_RegFile/N2BEG[2] Tile_X4Y12_RegFile/N2BEG[3] Tile_X4Y12_RegFile/N2BEG[4]
+ Tile_X4Y12_RegFile/N2BEG[5] Tile_X4Y12_RegFile/N2BEG[6] Tile_X4Y12_RegFile/N2BEG[7]
+ Tile_X4Y11_RegFile/N4BEG[0] Tile_X4Y11_RegFile/N4BEG[10] Tile_X4Y11_RegFile/N4BEG[11]
+ Tile_X4Y11_RegFile/N4BEG[12] Tile_X4Y11_RegFile/N4BEG[13] Tile_X4Y11_RegFile/N4BEG[14]
+ Tile_X4Y11_RegFile/N4BEG[15] Tile_X4Y11_RegFile/N4BEG[1] Tile_X4Y11_RegFile/N4BEG[2]
+ Tile_X4Y11_RegFile/N4BEG[3] Tile_X4Y11_RegFile/N4BEG[4] Tile_X4Y11_RegFile/N4BEG[5]
+ Tile_X4Y11_RegFile/N4BEG[6] Tile_X4Y11_RegFile/N4BEG[7] Tile_X4Y11_RegFile/N4BEG[8]
+ Tile_X4Y11_RegFile/N4BEG[9] Tile_X4Y12_RegFile/N4BEG[0] Tile_X4Y12_RegFile/N4BEG[10]
+ Tile_X4Y12_RegFile/N4BEG[11] Tile_X4Y12_RegFile/N4BEG[12] Tile_X4Y12_RegFile/N4BEG[13]
+ Tile_X4Y12_RegFile/N4BEG[14] Tile_X4Y12_RegFile/N4BEG[15] Tile_X4Y12_RegFile/N4BEG[1]
+ Tile_X4Y12_RegFile/N4BEG[2] Tile_X4Y12_RegFile/N4BEG[3] Tile_X4Y12_RegFile/N4BEG[4]
+ Tile_X4Y12_RegFile/N4BEG[5] Tile_X4Y12_RegFile/N4BEG[6] Tile_X4Y12_RegFile/N4BEG[7]
+ Tile_X4Y12_RegFile/N4BEG[8] Tile_X4Y12_RegFile/N4BEG[9] Tile_X4Y11_RegFile/NN4BEG[0]
+ Tile_X4Y11_RegFile/NN4BEG[10] Tile_X4Y11_RegFile/NN4BEG[11] Tile_X4Y11_RegFile/NN4BEG[12]
+ Tile_X4Y11_RegFile/NN4BEG[13] Tile_X4Y11_RegFile/NN4BEG[14] Tile_X4Y11_RegFile/NN4BEG[15]
+ Tile_X4Y11_RegFile/NN4BEG[1] Tile_X4Y11_RegFile/NN4BEG[2] Tile_X4Y11_RegFile/NN4BEG[3]
+ Tile_X4Y11_RegFile/NN4BEG[4] Tile_X4Y11_RegFile/NN4BEG[5] Tile_X4Y11_RegFile/NN4BEG[6]
+ Tile_X4Y11_RegFile/NN4BEG[7] Tile_X4Y11_RegFile/NN4BEG[8] Tile_X4Y11_RegFile/NN4BEG[9]
+ Tile_X4Y12_RegFile/NN4BEG[0] Tile_X4Y12_RegFile/NN4BEG[10] Tile_X4Y12_RegFile/NN4BEG[11]
+ Tile_X4Y12_RegFile/NN4BEG[12] Tile_X4Y12_RegFile/NN4BEG[13] Tile_X4Y12_RegFile/NN4BEG[14]
+ Tile_X4Y12_RegFile/NN4BEG[15] Tile_X4Y12_RegFile/NN4BEG[1] Tile_X4Y12_RegFile/NN4BEG[2]
+ Tile_X4Y12_RegFile/NN4BEG[3] Tile_X4Y12_RegFile/NN4BEG[4] Tile_X4Y12_RegFile/NN4BEG[5]
+ Tile_X4Y12_RegFile/NN4BEG[6] Tile_X4Y12_RegFile/NN4BEG[7] Tile_X4Y12_RegFile/NN4BEG[8]
+ Tile_X4Y12_RegFile/NN4BEG[9] Tile_X4Y12_RegFile/S1END[0] Tile_X4Y12_RegFile/S1END[1]
+ Tile_X4Y12_RegFile/S1END[2] Tile_X4Y12_RegFile/S1END[3] Tile_X4Y11_RegFile/S1END[0]
+ Tile_X4Y11_RegFile/S1END[1] Tile_X4Y11_RegFile/S1END[2] Tile_X4Y11_RegFile/S1END[3]
+ Tile_X4Y12_RegFile/S2MID[0] Tile_X4Y12_RegFile/S2MID[1] Tile_X4Y12_RegFile/S2MID[2]
+ Tile_X4Y12_RegFile/S2MID[3] Tile_X4Y12_RegFile/S2MID[4] Tile_X4Y12_RegFile/S2MID[5]
+ Tile_X4Y12_RegFile/S2MID[6] Tile_X4Y12_RegFile/S2MID[7] Tile_X4Y12_RegFile/S2END[0]
+ Tile_X4Y12_RegFile/S2END[1] Tile_X4Y12_RegFile/S2END[2] Tile_X4Y12_RegFile/S2END[3]
+ Tile_X4Y12_RegFile/S2END[4] Tile_X4Y12_RegFile/S2END[5] Tile_X4Y12_RegFile/S2END[6]
+ Tile_X4Y12_RegFile/S2END[7] Tile_X4Y11_RegFile/S2END[0] Tile_X4Y11_RegFile/S2END[1]
+ Tile_X4Y11_RegFile/S2END[2] Tile_X4Y11_RegFile/S2END[3] Tile_X4Y11_RegFile/S2END[4]
+ Tile_X4Y11_RegFile/S2END[5] Tile_X4Y11_RegFile/S2END[6] Tile_X4Y11_RegFile/S2END[7]
+ Tile_X4Y11_RegFile/S2MID[0] Tile_X4Y11_RegFile/S2MID[1] Tile_X4Y11_RegFile/S2MID[2]
+ Tile_X4Y11_RegFile/S2MID[3] Tile_X4Y11_RegFile/S2MID[4] Tile_X4Y11_RegFile/S2MID[5]
+ Tile_X4Y11_RegFile/S2MID[6] Tile_X4Y11_RegFile/S2MID[7] Tile_X4Y12_RegFile/S4END[0]
+ Tile_X4Y12_RegFile/S4END[10] Tile_X4Y12_RegFile/S4END[11] Tile_X4Y12_RegFile/S4END[12]
+ Tile_X4Y12_RegFile/S4END[13] Tile_X4Y12_RegFile/S4END[14] Tile_X4Y12_RegFile/S4END[15]
+ Tile_X4Y12_RegFile/S4END[1] Tile_X4Y12_RegFile/S4END[2] Tile_X4Y12_RegFile/S4END[3]
+ Tile_X4Y12_RegFile/S4END[4] Tile_X4Y12_RegFile/S4END[5] Tile_X4Y12_RegFile/S4END[6]
+ Tile_X4Y12_RegFile/S4END[7] Tile_X4Y12_RegFile/S4END[8] Tile_X4Y12_RegFile/S4END[9]
+ Tile_X4Y11_RegFile/S4END[0] Tile_X4Y11_RegFile/S4END[10] Tile_X4Y11_RegFile/S4END[11]
+ Tile_X4Y11_RegFile/S4END[12] Tile_X4Y11_RegFile/S4END[13] Tile_X4Y11_RegFile/S4END[14]
+ Tile_X4Y11_RegFile/S4END[15] Tile_X4Y11_RegFile/S4END[1] Tile_X4Y11_RegFile/S4END[2]
+ Tile_X4Y11_RegFile/S4END[3] Tile_X4Y11_RegFile/S4END[4] Tile_X4Y11_RegFile/S4END[5]
+ Tile_X4Y11_RegFile/S4END[6] Tile_X4Y11_RegFile/S4END[7] Tile_X4Y11_RegFile/S4END[8]
+ Tile_X4Y11_RegFile/S4END[9] Tile_X4Y12_RegFile/SS4END[0] Tile_X4Y12_RegFile/SS4END[10]
+ Tile_X4Y12_RegFile/SS4END[11] Tile_X4Y12_RegFile/SS4END[12] Tile_X4Y12_RegFile/SS4END[13]
+ Tile_X4Y12_RegFile/SS4END[14] Tile_X4Y12_RegFile/SS4END[15] Tile_X4Y12_RegFile/SS4END[1]
+ Tile_X4Y12_RegFile/SS4END[2] Tile_X4Y12_RegFile/SS4END[3] Tile_X4Y12_RegFile/SS4END[4]
+ Tile_X4Y12_RegFile/SS4END[5] Tile_X4Y12_RegFile/SS4END[6] Tile_X4Y12_RegFile/SS4END[7]
+ Tile_X4Y12_RegFile/SS4END[8] Tile_X4Y12_RegFile/SS4END[9] Tile_X4Y11_RegFile/SS4END[0]
+ Tile_X4Y11_RegFile/SS4END[10] Tile_X4Y11_RegFile/SS4END[11] Tile_X4Y11_RegFile/SS4END[12]
+ Tile_X4Y11_RegFile/SS4END[13] Tile_X4Y11_RegFile/SS4END[14] Tile_X4Y11_RegFile/SS4END[15]
+ Tile_X4Y11_RegFile/SS4END[1] Tile_X4Y11_RegFile/SS4END[2] Tile_X4Y11_RegFile/SS4END[3]
+ Tile_X4Y11_RegFile/SS4END[4] Tile_X4Y11_RegFile/SS4END[5] Tile_X4Y11_RegFile/SS4END[6]
+ Tile_X4Y11_RegFile/SS4END[7] Tile_X4Y11_RegFile/SS4END[8] Tile_X4Y11_RegFile/SS4END[9]
+ Tile_X4Y11_RegFile/UserCLK Tile_X4Y10_RegFile/UserCLK VGND VPWR Tile_X3Y11_LUT4AB/W1END[0]
+ Tile_X3Y11_LUT4AB/W1END[1] Tile_X3Y11_LUT4AB/W1END[2] Tile_X3Y11_LUT4AB/W1END[3]
+ Tile_X5Y11_LUT4AB/W1BEG[0] Tile_X5Y11_LUT4AB/W1BEG[1] Tile_X5Y11_LUT4AB/W1BEG[2]
+ Tile_X5Y11_LUT4AB/W1BEG[3] Tile_X3Y11_LUT4AB/W2MID[0] Tile_X3Y11_LUT4AB/W2MID[1]
+ Tile_X3Y11_LUT4AB/W2MID[2] Tile_X3Y11_LUT4AB/W2MID[3] Tile_X3Y11_LUT4AB/W2MID[4]
+ Tile_X3Y11_LUT4AB/W2MID[5] Tile_X3Y11_LUT4AB/W2MID[6] Tile_X3Y11_LUT4AB/W2MID[7]
+ Tile_X3Y11_LUT4AB/W2END[0] Tile_X3Y11_LUT4AB/W2END[1] Tile_X3Y11_LUT4AB/W2END[2]
+ Tile_X3Y11_LUT4AB/W2END[3] Tile_X3Y11_LUT4AB/W2END[4] Tile_X3Y11_LUT4AB/W2END[5]
+ Tile_X3Y11_LUT4AB/W2END[6] Tile_X3Y11_LUT4AB/W2END[7] Tile_X5Y11_LUT4AB/W2BEGb[0]
+ Tile_X5Y11_LUT4AB/W2BEGb[1] Tile_X5Y11_LUT4AB/W2BEGb[2] Tile_X5Y11_LUT4AB/W2BEGb[3]
+ Tile_X5Y11_LUT4AB/W2BEGb[4] Tile_X5Y11_LUT4AB/W2BEGb[5] Tile_X5Y11_LUT4AB/W2BEGb[6]
+ Tile_X5Y11_LUT4AB/W2BEGb[7] Tile_X5Y11_LUT4AB/W2BEG[0] Tile_X5Y11_LUT4AB/W2BEG[1]
+ Tile_X5Y11_LUT4AB/W2BEG[2] Tile_X5Y11_LUT4AB/W2BEG[3] Tile_X5Y11_LUT4AB/W2BEG[4]
+ Tile_X5Y11_LUT4AB/W2BEG[5] Tile_X5Y11_LUT4AB/W2BEG[6] Tile_X5Y11_LUT4AB/W2BEG[7]
+ Tile_X3Y11_LUT4AB/W6END[0] Tile_X3Y11_LUT4AB/W6END[10] Tile_X3Y11_LUT4AB/W6END[11]
+ Tile_X3Y11_LUT4AB/W6END[1] Tile_X3Y11_LUT4AB/W6END[2] Tile_X3Y11_LUT4AB/W6END[3]
+ Tile_X3Y11_LUT4AB/W6END[4] Tile_X3Y11_LUT4AB/W6END[5] Tile_X3Y11_LUT4AB/W6END[6]
+ Tile_X3Y11_LUT4AB/W6END[7] Tile_X3Y11_LUT4AB/W6END[8] Tile_X3Y11_LUT4AB/W6END[9]
+ Tile_X5Y11_LUT4AB/W6BEG[0] Tile_X5Y11_LUT4AB/W6BEG[10] Tile_X5Y11_LUT4AB/W6BEG[11]
+ Tile_X5Y11_LUT4AB/W6BEG[1] Tile_X5Y11_LUT4AB/W6BEG[2] Tile_X5Y11_LUT4AB/W6BEG[3]
+ Tile_X5Y11_LUT4AB/W6BEG[4] Tile_X5Y11_LUT4AB/W6BEG[5] Tile_X5Y11_LUT4AB/W6BEG[6]
+ Tile_X5Y11_LUT4AB/W6BEG[7] Tile_X5Y11_LUT4AB/W6BEG[8] Tile_X5Y11_LUT4AB/W6BEG[9]
+ Tile_X3Y11_LUT4AB/WW4END[0] Tile_X3Y11_LUT4AB/WW4END[10] Tile_X3Y11_LUT4AB/WW4END[11]
+ Tile_X3Y11_LUT4AB/WW4END[12] Tile_X3Y11_LUT4AB/WW4END[13] Tile_X3Y11_LUT4AB/WW4END[14]
+ Tile_X3Y11_LUT4AB/WW4END[15] Tile_X3Y11_LUT4AB/WW4END[1] Tile_X3Y11_LUT4AB/WW4END[2]
+ Tile_X3Y11_LUT4AB/WW4END[3] Tile_X3Y11_LUT4AB/WW4END[4] Tile_X3Y11_LUT4AB/WW4END[5]
+ Tile_X3Y11_LUT4AB/WW4END[6] Tile_X3Y11_LUT4AB/WW4END[7] Tile_X3Y11_LUT4AB/WW4END[8]
+ Tile_X3Y11_LUT4AB/WW4END[9] Tile_X5Y11_LUT4AB/WW4BEG[0] Tile_X5Y11_LUT4AB/WW4BEG[10]
+ Tile_X5Y11_LUT4AB/WW4BEG[11] Tile_X5Y11_LUT4AB/WW4BEG[12] Tile_X5Y11_LUT4AB/WW4BEG[13]
+ Tile_X5Y11_LUT4AB/WW4BEG[14] Tile_X5Y11_LUT4AB/WW4BEG[15] Tile_X5Y11_LUT4AB/WW4BEG[1]
+ Tile_X5Y11_LUT4AB/WW4BEG[2] Tile_X5Y11_LUT4AB/WW4BEG[3] Tile_X5Y11_LUT4AB/WW4BEG[4]
+ Tile_X5Y11_LUT4AB/WW4BEG[5] Tile_X5Y11_LUT4AB/WW4BEG[6] Tile_X5Y11_LUT4AB/WW4BEG[7]
+ Tile_X5Y11_LUT4AB/WW4BEG[8] Tile_X5Y11_LUT4AB/WW4BEG[9] RegFile
XTile_X8Y2_LUT4AB Tile_X8Y3_LUT4AB/Co Tile_X8Y2_LUT4AB/Co Tile_X9Y2_LUT4AB/E1END[0]
+ Tile_X9Y2_LUT4AB/E1END[1] Tile_X9Y2_LUT4AB/E1END[2] Tile_X9Y2_LUT4AB/E1END[3] Tile_X8Y2_LUT4AB/E1END[0]
+ Tile_X8Y2_LUT4AB/E1END[1] Tile_X8Y2_LUT4AB/E1END[2] Tile_X8Y2_LUT4AB/E1END[3] Tile_X9Y2_LUT4AB/E2MID[0]
+ Tile_X9Y2_LUT4AB/E2MID[1] Tile_X9Y2_LUT4AB/E2MID[2] Tile_X9Y2_LUT4AB/E2MID[3] Tile_X9Y2_LUT4AB/E2MID[4]
+ Tile_X9Y2_LUT4AB/E2MID[5] Tile_X9Y2_LUT4AB/E2MID[6] Tile_X9Y2_LUT4AB/E2MID[7] Tile_X9Y2_LUT4AB/E2END[0]
+ Tile_X9Y2_LUT4AB/E2END[1] Tile_X9Y2_LUT4AB/E2END[2] Tile_X9Y2_LUT4AB/E2END[3] Tile_X9Y2_LUT4AB/E2END[4]
+ Tile_X9Y2_LUT4AB/E2END[5] Tile_X9Y2_LUT4AB/E2END[6] Tile_X9Y2_LUT4AB/E2END[7] Tile_X8Y2_LUT4AB/E2END[0]
+ Tile_X8Y2_LUT4AB/E2END[1] Tile_X8Y2_LUT4AB/E2END[2] Tile_X8Y2_LUT4AB/E2END[3] Tile_X8Y2_LUT4AB/E2END[4]
+ Tile_X8Y2_LUT4AB/E2END[5] Tile_X8Y2_LUT4AB/E2END[6] Tile_X8Y2_LUT4AB/E2END[7] Tile_X8Y2_LUT4AB/E2MID[0]
+ Tile_X8Y2_LUT4AB/E2MID[1] Tile_X8Y2_LUT4AB/E2MID[2] Tile_X8Y2_LUT4AB/E2MID[3] Tile_X8Y2_LUT4AB/E2MID[4]
+ Tile_X8Y2_LUT4AB/E2MID[5] Tile_X8Y2_LUT4AB/E2MID[6] Tile_X8Y2_LUT4AB/E2MID[7] Tile_X9Y2_LUT4AB/E6END[0]
+ Tile_X9Y2_LUT4AB/E6END[10] Tile_X9Y2_LUT4AB/E6END[11] Tile_X9Y2_LUT4AB/E6END[1]
+ Tile_X9Y2_LUT4AB/E6END[2] Tile_X9Y2_LUT4AB/E6END[3] Tile_X9Y2_LUT4AB/E6END[4] Tile_X9Y2_LUT4AB/E6END[5]
+ Tile_X9Y2_LUT4AB/E6END[6] Tile_X9Y2_LUT4AB/E6END[7] Tile_X9Y2_LUT4AB/E6END[8] Tile_X9Y2_LUT4AB/E6END[9]
+ Tile_X8Y2_LUT4AB/E6END[0] Tile_X8Y2_LUT4AB/E6END[10] Tile_X8Y2_LUT4AB/E6END[11]
+ Tile_X8Y2_LUT4AB/E6END[1] Tile_X8Y2_LUT4AB/E6END[2] Tile_X8Y2_LUT4AB/E6END[3] Tile_X8Y2_LUT4AB/E6END[4]
+ Tile_X8Y2_LUT4AB/E6END[5] Tile_X8Y2_LUT4AB/E6END[6] Tile_X8Y2_LUT4AB/E6END[7] Tile_X8Y2_LUT4AB/E6END[8]
+ Tile_X8Y2_LUT4AB/E6END[9] Tile_X9Y2_LUT4AB/EE4END[0] Tile_X9Y2_LUT4AB/EE4END[10]
+ Tile_X9Y2_LUT4AB/EE4END[11] Tile_X9Y2_LUT4AB/EE4END[12] Tile_X9Y2_LUT4AB/EE4END[13]
+ Tile_X9Y2_LUT4AB/EE4END[14] Tile_X9Y2_LUT4AB/EE4END[15] Tile_X9Y2_LUT4AB/EE4END[1]
+ Tile_X9Y2_LUT4AB/EE4END[2] Tile_X9Y2_LUT4AB/EE4END[3] Tile_X9Y2_LUT4AB/EE4END[4]
+ Tile_X9Y2_LUT4AB/EE4END[5] Tile_X9Y2_LUT4AB/EE4END[6] Tile_X9Y2_LUT4AB/EE4END[7]
+ Tile_X9Y2_LUT4AB/EE4END[8] Tile_X9Y2_LUT4AB/EE4END[9] Tile_X8Y2_LUT4AB/EE4END[0]
+ Tile_X8Y2_LUT4AB/EE4END[10] Tile_X8Y2_LUT4AB/EE4END[11] Tile_X8Y2_LUT4AB/EE4END[12]
+ Tile_X8Y2_LUT4AB/EE4END[13] Tile_X8Y2_LUT4AB/EE4END[14] Tile_X8Y2_LUT4AB/EE4END[15]
+ Tile_X8Y2_LUT4AB/EE4END[1] Tile_X8Y2_LUT4AB/EE4END[2] Tile_X8Y2_LUT4AB/EE4END[3]
+ Tile_X8Y2_LUT4AB/EE4END[4] Tile_X8Y2_LUT4AB/EE4END[5] Tile_X8Y2_LUT4AB/EE4END[6]
+ Tile_X8Y2_LUT4AB/EE4END[7] Tile_X8Y2_LUT4AB/EE4END[8] Tile_X8Y2_LUT4AB/EE4END[9]
+ Tile_X8Y2_LUT4AB/FrameData[0] Tile_X8Y2_LUT4AB/FrameData[10] Tile_X8Y2_LUT4AB/FrameData[11]
+ Tile_X8Y2_LUT4AB/FrameData[12] Tile_X8Y2_LUT4AB/FrameData[13] Tile_X8Y2_LUT4AB/FrameData[14]
+ Tile_X8Y2_LUT4AB/FrameData[15] Tile_X8Y2_LUT4AB/FrameData[16] Tile_X8Y2_LUT4AB/FrameData[17]
+ Tile_X8Y2_LUT4AB/FrameData[18] Tile_X8Y2_LUT4AB/FrameData[19] Tile_X8Y2_LUT4AB/FrameData[1]
+ Tile_X8Y2_LUT4AB/FrameData[20] Tile_X8Y2_LUT4AB/FrameData[21] Tile_X8Y2_LUT4AB/FrameData[22]
+ Tile_X8Y2_LUT4AB/FrameData[23] Tile_X8Y2_LUT4AB/FrameData[24] Tile_X8Y2_LUT4AB/FrameData[25]
+ Tile_X8Y2_LUT4AB/FrameData[26] Tile_X8Y2_LUT4AB/FrameData[27] Tile_X8Y2_LUT4AB/FrameData[28]
+ Tile_X8Y2_LUT4AB/FrameData[29] Tile_X8Y2_LUT4AB/FrameData[2] Tile_X8Y2_LUT4AB/FrameData[30]
+ Tile_X8Y2_LUT4AB/FrameData[31] Tile_X8Y2_LUT4AB/FrameData[3] Tile_X8Y2_LUT4AB/FrameData[4]
+ Tile_X8Y2_LUT4AB/FrameData[5] Tile_X8Y2_LUT4AB/FrameData[6] Tile_X8Y2_LUT4AB/FrameData[7]
+ Tile_X8Y2_LUT4AB/FrameData[8] Tile_X8Y2_LUT4AB/FrameData[9] Tile_X9Y2_LUT4AB/FrameData[0]
+ Tile_X9Y2_LUT4AB/FrameData[10] Tile_X9Y2_LUT4AB/FrameData[11] Tile_X9Y2_LUT4AB/FrameData[12]
+ Tile_X9Y2_LUT4AB/FrameData[13] Tile_X9Y2_LUT4AB/FrameData[14] Tile_X9Y2_LUT4AB/FrameData[15]
+ Tile_X9Y2_LUT4AB/FrameData[16] Tile_X9Y2_LUT4AB/FrameData[17] Tile_X9Y2_LUT4AB/FrameData[18]
+ Tile_X9Y2_LUT4AB/FrameData[19] Tile_X9Y2_LUT4AB/FrameData[1] Tile_X9Y2_LUT4AB/FrameData[20]
+ Tile_X9Y2_LUT4AB/FrameData[21] Tile_X9Y2_LUT4AB/FrameData[22] Tile_X9Y2_LUT4AB/FrameData[23]
+ Tile_X9Y2_LUT4AB/FrameData[24] Tile_X9Y2_LUT4AB/FrameData[25] Tile_X9Y2_LUT4AB/FrameData[26]
+ Tile_X9Y2_LUT4AB/FrameData[27] Tile_X9Y2_LUT4AB/FrameData[28] Tile_X9Y2_LUT4AB/FrameData[29]
+ Tile_X9Y2_LUT4AB/FrameData[2] Tile_X9Y2_LUT4AB/FrameData[30] Tile_X9Y2_LUT4AB/FrameData[31]
+ Tile_X9Y2_LUT4AB/FrameData[3] Tile_X9Y2_LUT4AB/FrameData[4] Tile_X9Y2_LUT4AB/FrameData[5]
+ Tile_X9Y2_LUT4AB/FrameData[6] Tile_X9Y2_LUT4AB/FrameData[7] Tile_X9Y2_LUT4AB/FrameData[8]
+ Tile_X9Y2_LUT4AB/FrameData[9] Tile_X8Y2_LUT4AB/FrameStrobe[0] Tile_X8Y2_LUT4AB/FrameStrobe[10]
+ Tile_X8Y2_LUT4AB/FrameStrobe[11] Tile_X8Y2_LUT4AB/FrameStrobe[12] Tile_X8Y2_LUT4AB/FrameStrobe[13]
+ Tile_X8Y2_LUT4AB/FrameStrobe[14] Tile_X8Y2_LUT4AB/FrameStrobe[15] Tile_X8Y2_LUT4AB/FrameStrobe[16]
+ Tile_X8Y2_LUT4AB/FrameStrobe[17] Tile_X8Y2_LUT4AB/FrameStrobe[18] Tile_X8Y2_LUT4AB/FrameStrobe[19]
+ Tile_X8Y2_LUT4AB/FrameStrobe[1] Tile_X8Y2_LUT4AB/FrameStrobe[2] Tile_X8Y2_LUT4AB/FrameStrobe[3]
+ Tile_X8Y2_LUT4AB/FrameStrobe[4] Tile_X8Y2_LUT4AB/FrameStrobe[5] Tile_X8Y2_LUT4AB/FrameStrobe[6]
+ Tile_X8Y2_LUT4AB/FrameStrobe[7] Tile_X8Y2_LUT4AB/FrameStrobe[8] Tile_X8Y2_LUT4AB/FrameStrobe[9]
+ Tile_X8Y1_LUT4AB/FrameStrobe[0] Tile_X8Y1_LUT4AB/FrameStrobe[10] Tile_X8Y1_LUT4AB/FrameStrobe[11]
+ Tile_X8Y1_LUT4AB/FrameStrobe[12] Tile_X8Y1_LUT4AB/FrameStrobe[13] Tile_X8Y1_LUT4AB/FrameStrobe[14]
+ Tile_X8Y1_LUT4AB/FrameStrobe[15] Tile_X8Y1_LUT4AB/FrameStrobe[16] Tile_X8Y1_LUT4AB/FrameStrobe[17]
+ Tile_X8Y1_LUT4AB/FrameStrobe[18] Tile_X8Y1_LUT4AB/FrameStrobe[19] Tile_X8Y1_LUT4AB/FrameStrobe[1]
+ Tile_X8Y1_LUT4AB/FrameStrobe[2] Tile_X8Y1_LUT4AB/FrameStrobe[3] Tile_X8Y1_LUT4AB/FrameStrobe[4]
+ Tile_X8Y1_LUT4AB/FrameStrobe[5] Tile_X8Y1_LUT4AB/FrameStrobe[6] Tile_X8Y1_LUT4AB/FrameStrobe[7]
+ Tile_X8Y1_LUT4AB/FrameStrobe[8] Tile_X8Y1_LUT4AB/FrameStrobe[9] Tile_X8Y2_LUT4AB/N1BEG[0]
+ Tile_X8Y2_LUT4AB/N1BEG[1] Tile_X8Y2_LUT4AB/N1BEG[2] Tile_X8Y2_LUT4AB/N1BEG[3] Tile_X8Y3_LUT4AB/N1BEG[0]
+ Tile_X8Y3_LUT4AB/N1BEG[1] Tile_X8Y3_LUT4AB/N1BEG[2] Tile_X8Y3_LUT4AB/N1BEG[3] Tile_X8Y2_LUT4AB/N2BEG[0]
+ Tile_X8Y2_LUT4AB/N2BEG[1] Tile_X8Y2_LUT4AB/N2BEG[2] Tile_X8Y2_LUT4AB/N2BEG[3] Tile_X8Y2_LUT4AB/N2BEG[4]
+ Tile_X8Y2_LUT4AB/N2BEG[5] Tile_X8Y2_LUT4AB/N2BEG[6] Tile_X8Y2_LUT4AB/N2BEG[7] Tile_X8Y1_LUT4AB/N2END[0]
+ Tile_X8Y1_LUT4AB/N2END[1] Tile_X8Y1_LUT4AB/N2END[2] Tile_X8Y1_LUT4AB/N2END[3] Tile_X8Y1_LUT4AB/N2END[4]
+ Tile_X8Y1_LUT4AB/N2END[5] Tile_X8Y1_LUT4AB/N2END[6] Tile_X8Y1_LUT4AB/N2END[7] Tile_X8Y2_LUT4AB/N2END[0]
+ Tile_X8Y2_LUT4AB/N2END[1] Tile_X8Y2_LUT4AB/N2END[2] Tile_X8Y2_LUT4AB/N2END[3] Tile_X8Y2_LUT4AB/N2END[4]
+ Tile_X8Y2_LUT4AB/N2END[5] Tile_X8Y2_LUT4AB/N2END[6] Tile_X8Y2_LUT4AB/N2END[7] Tile_X8Y3_LUT4AB/N2BEG[0]
+ Tile_X8Y3_LUT4AB/N2BEG[1] Tile_X8Y3_LUT4AB/N2BEG[2] Tile_X8Y3_LUT4AB/N2BEG[3] Tile_X8Y3_LUT4AB/N2BEG[4]
+ Tile_X8Y3_LUT4AB/N2BEG[5] Tile_X8Y3_LUT4AB/N2BEG[6] Tile_X8Y3_LUT4AB/N2BEG[7] Tile_X8Y2_LUT4AB/N4BEG[0]
+ Tile_X8Y2_LUT4AB/N4BEG[10] Tile_X8Y2_LUT4AB/N4BEG[11] Tile_X8Y2_LUT4AB/N4BEG[12]
+ Tile_X8Y2_LUT4AB/N4BEG[13] Tile_X8Y2_LUT4AB/N4BEG[14] Tile_X8Y2_LUT4AB/N4BEG[15]
+ Tile_X8Y2_LUT4AB/N4BEG[1] Tile_X8Y2_LUT4AB/N4BEG[2] Tile_X8Y2_LUT4AB/N4BEG[3] Tile_X8Y2_LUT4AB/N4BEG[4]
+ Tile_X8Y2_LUT4AB/N4BEG[5] Tile_X8Y2_LUT4AB/N4BEG[6] Tile_X8Y2_LUT4AB/N4BEG[7] Tile_X8Y2_LUT4AB/N4BEG[8]
+ Tile_X8Y2_LUT4AB/N4BEG[9] Tile_X8Y3_LUT4AB/N4BEG[0] Tile_X8Y3_LUT4AB/N4BEG[10] Tile_X8Y3_LUT4AB/N4BEG[11]
+ Tile_X8Y3_LUT4AB/N4BEG[12] Tile_X8Y3_LUT4AB/N4BEG[13] Tile_X8Y3_LUT4AB/N4BEG[14]
+ Tile_X8Y3_LUT4AB/N4BEG[15] Tile_X8Y3_LUT4AB/N4BEG[1] Tile_X8Y3_LUT4AB/N4BEG[2] Tile_X8Y3_LUT4AB/N4BEG[3]
+ Tile_X8Y3_LUT4AB/N4BEG[4] Tile_X8Y3_LUT4AB/N4BEG[5] Tile_X8Y3_LUT4AB/N4BEG[6] Tile_X8Y3_LUT4AB/N4BEG[7]
+ Tile_X8Y3_LUT4AB/N4BEG[8] Tile_X8Y3_LUT4AB/N4BEG[9] Tile_X8Y2_LUT4AB/NN4BEG[0] Tile_X8Y2_LUT4AB/NN4BEG[10]
+ Tile_X8Y2_LUT4AB/NN4BEG[11] Tile_X8Y2_LUT4AB/NN4BEG[12] Tile_X8Y2_LUT4AB/NN4BEG[13]
+ Tile_X8Y2_LUT4AB/NN4BEG[14] Tile_X8Y2_LUT4AB/NN4BEG[15] Tile_X8Y2_LUT4AB/NN4BEG[1]
+ Tile_X8Y2_LUT4AB/NN4BEG[2] Tile_X8Y2_LUT4AB/NN4BEG[3] Tile_X8Y2_LUT4AB/NN4BEG[4]
+ Tile_X8Y2_LUT4AB/NN4BEG[5] Tile_X8Y2_LUT4AB/NN4BEG[6] Tile_X8Y2_LUT4AB/NN4BEG[7]
+ Tile_X8Y2_LUT4AB/NN4BEG[8] Tile_X8Y2_LUT4AB/NN4BEG[9] Tile_X8Y3_LUT4AB/NN4BEG[0]
+ Tile_X8Y3_LUT4AB/NN4BEG[10] Tile_X8Y3_LUT4AB/NN4BEG[11] Tile_X8Y3_LUT4AB/NN4BEG[12]
+ Tile_X8Y3_LUT4AB/NN4BEG[13] Tile_X8Y3_LUT4AB/NN4BEG[14] Tile_X8Y3_LUT4AB/NN4BEG[15]
+ Tile_X8Y3_LUT4AB/NN4BEG[1] Tile_X8Y3_LUT4AB/NN4BEG[2] Tile_X8Y3_LUT4AB/NN4BEG[3]
+ Tile_X8Y3_LUT4AB/NN4BEG[4] Tile_X8Y3_LUT4AB/NN4BEG[5] Tile_X8Y3_LUT4AB/NN4BEG[6]
+ Tile_X8Y3_LUT4AB/NN4BEG[7] Tile_X8Y3_LUT4AB/NN4BEG[8] Tile_X8Y3_LUT4AB/NN4BEG[9]
+ Tile_X8Y3_LUT4AB/S1END[0] Tile_X8Y3_LUT4AB/S1END[1] Tile_X8Y3_LUT4AB/S1END[2] Tile_X8Y3_LUT4AB/S1END[3]
+ Tile_X8Y2_LUT4AB/S1END[0] Tile_X8Y2_LUT4AB/S1END[1] Tile_X8Y2_LUT4AB/S1END[2] Tile_X8Y2_LUT4AB/S1END[3]
+ Tile_X8Y3_LUT4AB/S2MID[0] Tile_X8Y3_LUT4AB/S2MID[1] Tile_X8Y3_LUT4AB/S2MID[2] Tile_X8Y3_LUT4AB/S2MID[3]
+ Tile_X8Y3_LUT4AB/S2MID[4] Tile_X8Y3_LUT4AB/S2MID[5] Tile_X8Y3_LUT4AB/S2MID[6] Tile_X8Y3_LUT4AB/S2MID[7]
+ Tile_X8Y3_LUT4AB/S2END[0] Tile_X8Y3_LUT4AB/S2END[1] Tile_X8Y3_LUT4AB/S2END[2] Tile_X8Y3_LUT4AB/S2END[3]
+ Tile_X8Y3_LUT4AB/S2END[4] Tile_X8Y3_LUT4AB/S2END[5] Tile_X8Y3_LUT4AB/S2END[6] Tile_X8Y3_LUT4AB/S2END[7]
+ Tile_X8Y2_LUT4AB/S2END[0] Tile_X8Y2_LUT4AB/S2END[1] Tile_X8Y2_LUT4AB/S2END[2] Tile_X8Y2_LUT4AB/S2END[3]
+ Tile_X8Y2_LUT4AB/S2END[4] Tile_X8Y2_LUT4AB/S2END[5] Tile_X8Y2_LUT4AB/S2END[6] Tile_X8Y2_LUT4AB/S2END[7]
+ Tile_X8Y2_LUT4AB/S2MID[0] Tile_X8Y2_LUT4AB/S2MID[1] Tile_X8Y2_LUT4AB/S2MID[2] Tile_X8Y2_LUT4AB/S2MID[3]
+ Tile_X8Y2_LUT4AB/S2MID[4] Tile_X8Y2_LUT4AB/S2MID[5] Tile_X8Y2_LUT4AB/S2MID[6] Tile_X8Y2_LUT4AB/S2MID[7]
+ Tile_X8Y3_LUT4AB/S4END[0] Tile_X8Y3_LUT4AB/S4END[10] Tile_X8Y3_LUT4AB/S4END[11]
+ Tile_X8Y3_LUT4AB/S4END[12] Tile_X8Y3_LUT4AB/S4END[13] Tile_X8Y3_LUT4AB/S4END[14]
+ Tile_X8Y3_LUT4AB/S4END[15] Tile_X8Y3_LUT4AB/S4END[1] Tile_X8Y3_LUT4AB/S4END[2] Tile_X8Y3_LUT4AB/S4END[3]
+ Tile_X8Y3_LUT4AB/S4END[4] Tile_X8Y3_LUT4AB/S4END[5] Tile_X8Y3_LUT4AB/S4END[6] Tile_X8Y3_LUT4AB/S4END[7]
+ Tile_X8Y3_LUT4AB/S4END[8] Tile_X8Y3_LUT4AB/S4END[9] Tile_X8Y2_LUT4AB/S4END[0] Tile_X8Y2_LUT4AB/S4END[10]
+ Tile_X8Y2_LUT4AB/S4END[11] Tile_X8Y2_LUT4AB/S4END[12] Tile_X8Y2_LUT4AB/S4END[13]
+ Tile_X8Y2_LUT4AB/S4END[14] Tile_X8Y2_LUT4AB/S4END[15] Tile_X8Y2_LUT4AB/S4END[1]
+ Tile_X8Y2_LUT4AB/S4END[2] Tile_X8Y2_LUT4AB/S4END[3] Tile_X8Y2_LUT4AB/S4END[4] Tile_X8Y2_LUT4AB/S4END[5]
+ Tile_X8Y2_LUT4AB/S4END[6] Tile_X8Y2_LUT4AB/S4END[7] Tile_X8Y2_LUT4AB/S4END[8] Tile_X8Y2_LUT4AB/S4END[9]
+ Tile_X8Y3_LUT4AB/SS4END[0] Tile_X8Y3_LUT4AB/SS4END[10] Tile_X8Y3_LUT4AB/SS4END[11]
+ Tile_X8Y3_LUT4AB/SS4END[12] Tile_X8Y3_LUT4AB/SS4END[13] Tile_X8Y3_LUT4AB/SS4END[14]
+ Tile_X8Y3_LUT4AB/SS4END[15] Tile_X8Y3_LUT4AB/SS4END[1] Tile_X8Y3_LUT4AB/SS4END[2]
+ Tile_X8Y3_LUT4AB/SS4END[3] Tile_X8Y3_LUT4AB/SS4END[4] Tile_X8Y3_LUT4AB/SS4END[5]
+ Tile_X8Y3_LUT4AB/SS4END[6] Tile_X8Y3_LUT4AB/SS4END[7] Tile_X8Y3_LUT4AB/SS4END[8]
+ Tile_X8Y3_LUT4AB/SS4END[9] Tile_X8Y2_LUT4AB/SS4END[0] Tile_X8Y2_LUT4AB/SS4END[10]
+ Tile_X8Y2_LUT4AB/SS4END[11] Tile_X8Y2_LUT4AB/SS4END[12] Tile_X8Y2_LUT4AB/SS4END[13]
+ Tile_X8Y2_LUT4AB/SS4END[14] Tile_X8Y2_LUT4AB/SS4END[15] Tile_X8Y2_LUT4AB/SS4END[1]
+ Tile_X8Y2_LUT4AB/SS4END[2] Tile_X8Y2_LUT4AB/SS4END[3] Tile_X8Y2_LUT4AB/SS4END[4]
+ Tile_X8Y2_LUT4AB/SS4END[5] Tile_X8Y2_LUT4AB/SS4END[6] Tile_X8Y2_LUT4AB/SS4END[7]
+ Tile_X8Y2_LUT4AB/SS4END[8] Tile_X8Y2_LUT4AB/SS4END[9] Tile_X8Y2_LUT4AB/UserCLK Tile_X8Y1_LUT4AB/UserCLK
+ VGND VPWR Tile_X8Y2_LUT4AB/W1BEG[0] Tile_X8Y2_LUT4AB/W1BEG[1] Tile_X8Y2_LUT4AB/W1BEG[2]
+ Tile_X8Y2_LUT4AB/W1BEG[3] Tile_X9Y2_LUT4AB/W1BEG[0] Tile_X9Y2_LUT4AB/W1BEG[1] Tile_X9Y2_LUT4AB/W1BEG[2]
+ Tile_X9Y2_LUT4AB/W1BEG[3] Tile_X8Y2_LUT4AB/W2BEG[0] Tile_X8Y2_LUT4AB/W2BEG[1] Tile_X8Y2_LUT4AB/W2BEG[2]
+ Tile_X8Y2_LUT4AB/W2BEG[3] Tile_X8Y2_LUT4AB/W2BEG[4] Tile_X8Y2_LUT4AB/W2BEG[5] Tile_X8Y2_LUT4AB/W2BEG[6]
+ Tile_X8Y2_LUT4AB/W2BEG[7] Tile_X8Y2_LUT4AB/W2BEGb[0] Tile_X8Y2_LUT4AB/W2BEGb[1]
+ Tile_X8Y2_LUT4AB/W2BEGb[2] Tile_X8Y2_LUT4AB/W2BEGb[3] Tile_X8Y2_LUT4AB/W2BEGb[4]
+ Tile_X8Y2_LUT4AB/W2BEGb[5] Tile_X8Y2_LUT4AB/W2BEGb[6] Tile_X8Y2_LUT4AB/W2BEGb[7]
+ Tile_X8Y2_LUT4AB/W2END[0] Tile_X8Y2_LUT4AB/W2END[1] Tile_X8Y2_LUT4AB/W2END[2] Tile_X8Y2_LUT4AB/W2END[3]
+ Tile_X8Y2_LUT4AB/W2END[4] Tile_X8Y2_LUT4AB/W2END[5] Tile_X8Y2_LUT4AB/W2END[6] Tile_X8Y2_LUT4AB/W2END[7]
+ Tile_X9Y2_LUT4AB/W2BEG[0] Tile_X9Y2_LUT4AB/W2BEG[1] Tile_X9Y2_LUT4AB/W2BEG[2] Tile_X9Y2_LUT4AB/W2BEG[3]
+ Tile_X9Y2_LUT4AB/W2BEG[4] Tile_X9Y2_LUT4AB/W2BEG[5] Tile_X9Y2_LUT4AB/W2BEG[6] Tile_X9Y2_LUT4AB/W2BEG[7]
+ Tile_X8Y2_LUT4AB/W6BEG[0] Tile_X8Y2_LUT4AB/W6BEG[10] Tile_X8Y2_LUT4AB/W6BEG[11]
+ Tile_X8Y2_LUT4AB/W6BEG[1] Tile_X8Y2_LUT4AB/W6BEG[2] Tile_X8Y2_LUT4AB/W6BEG[3] Tile_X8Y2_LUT4AB/W6BEG[4]
+ Tile_X8Y2_LUT4AB/W6BEG[5] Tile_X8Y2_LUT4AB/W6BEG[6] Tile_X8Y2_LUT4AB/W6BEG[7] Tile_X8Y2_LUT4AB/W6BEG[8]
+ Tile_X8Y2_LUT4AB/W6BEG[9] Tile_X9Y2_LUT4AB/W6BEG[0] Tile_X9Y2_LUT4AB/W6BEG[10] Tile_X9Y2_LUT4AB/W6BEG[11]
+ Tile_X9Y2_LUT4AB/W6BEG[1] Tile_X9Y2_LUT4AB/W6BEG[2] Tile_X9Y2_LUT4AB/W6BEG[3] Tile_X9Y2_LUT4AB/W6BEG[4]
+ Tile_X9Y2_LUT4AB/W6BEG[5] Tile_X9Y2_LUT4AB/W6BEG[6] Tile_X9Y2_LUT4AB/W6BEG[7] Tile_X9Y2_LUT4AB/W6BEG[8]
+ Tile_X9Y2_LUT4AB/W6BEG[9] Tile_X8Y2_LUT4AB/WW4BEG[0] Tile_X8Y2_LUT4AB/WW4BEG[10]
+ Tile_X8Y2_LUT4AB/WW4BEG[11] Tile_X8Y2_LUT4AB/WW4BEG[12] Tile_X8Y2_LUT4AB/WW4BEG[13]
+ Tile_X8Y2_LUT4AB/WW4BEG[14] Tile_X8Y2_LUT4AB/WW4BEG[15] Tile_X8Y2_LUT4AB/WW4BEG[1]
+ Tile_X8Y2_LUT4AB/WW4BEG[2] Tile_X8Y2_LUT4AB/WW4BEG[3] Tile_X8Y2_LUT4AB/WW4BEG[4]
+ Tile_X8Y2_LUT4AB/WW4BEG[5] Tile_X8Y2_LUT4AB/WW4BEG[6] Tile_X8Y2_LUT4AB/WW4BEG[7]
+ Tile_X8Y2_LUT4AB/WW4BEG[8] Tile_X8Y2_LUT4AB/WW4BEG[9] Tile_X9Y2_LUT4AB/WW4BEG[0]
+ Tile_X9Y2_LUT4AB/WW4BEG[10] Tile_X9Y2_LUT4AB/WW4BEG[11] Tile_X9Y2_LUT4AB/WW4BEG[12]
+ Tile_X9Y2_LUT4AB/WW4BEG[13] Tile_X9Y2_LUT4AB/WW4BEG[14] Tile_X9Y2_LUT4AB/WW4BEG[15]
+ Tile_X9Y2_LUT4AB/WW4BEG[1] Tile_X9Y2_LUT4AB/WW4BEG[2] Tile_X9Y2_LUT4AB/WW4BEG[3]
+ Tile_X9Y2_LUT4AB/WW4BEG[4] Tile_X9Y2_LUT4AB/WW4BEG[5] Tile_X9Y2_LUT4AB/WW4BEG[6]
+ Tile_X9Y2_LUT4AB/WW4BEG[7] Tile_X9Y2_LUT4AB/WW4BEG[8] Tile_X9Y2_LUT4AB/WW4BEG[9]
+ LUT4AB
XTile_X3Y12_LUT4AB Tile_X3Y13_LUT4AB/Co Tile_X3Y12_LUT4AB/Co Tile_X3Y12_LUT4AB/E1BEG[0]
+ Tile_X3Y12_LUT4AB/E1BEG[1] Tile_X3Y12_LUT4AB/E1BEG[2] Tile_X3Y12_LUT4AB/E1BEG[3]
+ Tile_X3Y12_LUT4AB/E1END[0] Tile_X3Y12_LUT4AB/E1END[1] Tile_X3Y12_LUT4AB/E1END[2]
+ Tile_X3Y12_LUT4AB/E1END[3] Tile_X3Y12_LUT4AB/E2BEG[0] Tile_X3Y12_LUT4AB/E2BEG[1]
+ Tile_X3Y12_LUT4AB/E2BEG[2] Tile_X3Y12_LUT4AB/E2BEG[3] Tile_X3Y12_LUT4AB/E2BEG[4]
+ Tile_X3Y12_LUT4AB/E2BEG[5] Tile_X3Y12_LUT4AB/E2BEG[6] Tile_X3Y12_LUT4AB/E2BEG[7]
+ Tile_X4Y12_RegFile/E2END[0] Tile_X4Y12_RegFile/E2END[1] Tile_X4Y12_RegFile/E2END[2]
+ Tile_X4Y12_RegFile/E2END[3] Tile_X4Y12_RegFile/E2END[4] Tile_X4Y12_RegFile/E2END[5]
+ Tile_X4Y12_RegFile/E2END[6] Tile_X4Y12_RegFile/E2END[7] Tile_X3Y12_LUT4AB/E2END[0]
+ Tile_X3Y12_LUT4AB/E2END[1] Tile_X3Y12_LUT4AB/E2END[2] Tile_X3Y12_LUT4AB/E2END[3]
+ Tile_X3Y12_LUT4AB/E2END[4] Tile_X3Y12_LUT4AB/E2END[5] Tile_X3Y12_LUT4AB/E2END[6]
+ Tile_X3Y12_LUT4AB/E2END[7] Tile_X3Y12_LUT4AB/E2MID[0] Tile_X3Y12_LUT4AB/E2MID[1]
+ Tile_X3Y12_LUT4AB/E2MID[2] Tile_X3Y12_LUT4AB/E2MID[3] Tile_X3Y12_LUT4AB/E2MID[4]
+ Tile_X3Y12_LUT4AB/E2MID[5] Tile_X3Y12_LUT4AB/E2MID[6] Tile_X3Y12_LUT4AB/E2MID[7]
+ Tile_X3Y12_LUT4AB/E6BEG[0] Tile_X3Y12_LUT4AB/E6BEG[10] Tile_X3Y12_LUT4AB/E6BEG[11]
+ Tile_X3Y12_LUT4AB/E6BEG[1] Tile_X3Y12_LUT4AB/E6BEG[2] Tile_X3Y12_LUT4AB/E6BEG[3]
+ Tile_X3Y12_LUT4AB/E6BEG[4] Tile_X3Y12_LUT4AB/E6BEG[5] Tile_X3Y12_LUT4AB/E6BEG[6]
+ Tile_X3Y12_LUT4AB/E6BEG[7] Tile_X3Y12_LUT4AB/E6BEG[8] Tile_X3Y12_LUT4AB/E6BEG[9]
+ Tile_X3Y12_LUT4AB/E6END[0] Tile_X3Y12_LUT4AB/E6END[10] Tile_X3Y12_LUT4AB/E6END[11]
+ Tile_X3Y12_LUT4AB/E6END[1] Tile_X3Y12_LUT4AB/E6END[2] Tile_X3Y12_LUT4AB/E6END[3]
+ Tile_X3Y12_LUT4AB/E6END[4] Tile_X3Y12_LUT4AB/E6END[5] Tile_X3Y12_LUT4AB/E6END[6]
+ Tile_X3Y12_LUT4AB/E6END[7] Tile_X3Y12_LUT4AB/E6END[8] Tile_X3Y12_LUT4AB/E6END[9]
+ Tile_X3Y12_LUT4AB/EE4BEG[0] Tile_X3Y12_LUT4AB/EE4BEG[10] Tile_X3Y12_LUT4AB/EE4BEG[11]
+ Tile_X3Y12_LUT4AB/EE4BEG[12] Tile_X3Y12_LUT4AB/EE4BEG[13] Tile_X3Y12_LUT4AB/EE4BEG[14]
+ Tile_X3Y12_LUT4AB/EE4BEG[15] Tile_X3Y12_LUT4AB/EE4BEG[1] Tile_X3Y12_LUT4AB/EE4BEG[2]
+ Tile_X3Y12_LUT4AB/EE4BEG[3] Tile_X3Y12_LUT4AB/EE4BEG[4] Tile_X3Y12_LUT4AB/EE4BEG[5]
+ Tile_X3Y12_LUT4AB/EE4BEG[6] Tile_X3Y12_LUT4AB/EE4BEG[7] Tile_X3Y12_LUT4AB/EE4BEG[8]
+ Tile_X3Y12_LUT4AB/EE4BEG[9] Tile_X3Y12_LUT4AB/EE4END[0] Tile_X3Y12_LUT4AB/EE4END[10]
+ Tile_X3Y12_LUT4AB/EE4END[11] Tile_X3Y12_LUT4AB/EE4END[12] Tile_X3Y12_LUT4AB/EE4END[13]
+ Tile_X3Y12_LUT4AB/EE4END[14] Tile_X3Y12_LUT4AB/EE4END[15] Tile_X3Y12_LUT4AB/EE4END[1]
+ Tile_X3Y12_LUT4AB/EE4END[2] Tile_X3Y12_LUT4AB/EE4END[3] Tile_X3Y12_LUT4AB/EE4END[4]
+ Tile_X3Y12_LUT4AB/EE4END[5] Tile_X3Y12_LUT4AB/EE4END[6] Tile_X3Y12_LUT4AB/EE4END[7]
+ Tile_X3Y12_LUT4AB/EE4END[8] Tile_X3Y12_LUT4AB/EE4END[9] Tile_X3Y12_LUT4AB/FrameData[0]
+ Tile_X3Y12_LUT4AB/FrameData[10] Tile_X3Y12_LUT4AB/FrameData[11] Tile_X3Y12_LUT4AB/FrameData[12]
+ Tile_X3Y12_LUT4AB/FrameData[13] Tile_X3Y12_LUT4AB/FrameData[14] Tile_X3Y12_LUT4AB/FrameData[15]
+ Tile_X3Y12_LUT4AB/FrameData[16] Tile_X3Y12_LUT4AB/FrameData[17] Tile_X3Y12_LUT4AB/FrameData[18]
+ Tile_X3Y12_LUT4AB/FrameData[19] Tile_X3Y12_LUT4AB/FrameData[1] Tile_X3Y12_LUT4AB/FrameData[20]
+ Tile_X3Y12_LUT4AB/FrameData[21] Tile_X3Y12_LUT4AB/FrameData[22] Tile_X3Y12_LUT4AB/FrameData[23]
+ Tile_X3Y12_LUT4AB/FrameData[24] Tile_X3Y12_LUT4AB/FrameData[25] Tile_X3Y12_LUT4AB/FrameData[26]
+ Tile_X3Y12_LUT4AB/FrameData[27] Tile_X3Y12_LUT4AB/FrameData[28] Tile_X3Y12_LUT4AB/FrameData[29]
+ Tile_X3Y12_LUT4AB/FrameData[2] Tile_X3Y12_LUT4AB/FrameData[30] Tile_X3Y12_LUT4AB/FrameData[31]
+ Tile_X3Y12_LUT4AB/FrameData[3] Tile_X3Y12_LUT4AB/FrameData[4] Tile_X3Y12_LUT4AB/FrameData[5]
+ Tile_X3Y12_LUT4AB/FrameData[6] Tile_X3Y12_LUT4AB/FrameData[7] Tile_X3Y12_LUT4AB/FrameData[8]
+ Tile_X3Y12_LUT4AB/FrameData[9] Tile_X4Y12_RegFile/FrameData[0] Tile_X4Y12_RegFile/FrameData[10]
+ Tile_X4Y12_RegFile/FrameData[11] Tile_X4Y12_RegFile/FrameData[12] Tile_X4Y12_RegFile/FrameData[13]
+ Tile_X4Y12_RegFile/FrameData[14] Tile_X4Y12_RegFile/FrameData[15] Tile_X4Y12_RegFile/FrameData[16]
+ Tile_X4Y12_RegFile/FrameData[17] Tile_X4Y12_RegFile/FrameData[18] Tile_X4Y12_RegFile/FrameData[19]
+ Tile_X4Y12_RegFile/FrameData[1] Tile_X4Y12_RegFile/FrameData[20] Tile_X4Y12_RegFile/FrameData[21]
+ Tile_X4Y12_RegFile/FrameData[22] Tile_X4Y12_RegFile/FrameData[23] Tile_X4Y12_RegFile/FrameData[24]
+ Tile_X4Y12_RegFile/FrameData[25] Tile_X4Y12_RegFile/FrameData[26] Tile_X4Y12_RegFile/FrameData[27]
+ Tile_X4Y12_RegFile/FrameData[28] Tile_X4Y12_RegFile/FrameData[29] Tile_X4Y12_RegFile/FrameData[2]
+ Tile_X4Y12_RegFile/FrameData[30] Tile_X4Y12_RegFile/FrameData[31] Tile_X4Y12_RegFile/FrameData[3]
+ Tile_X4Y12_RegFile/FrameData[4] Tile_X4Y12_RegFile/FrameData[5] Tile_X4Y12_RegFile/FrameData[6]
+ Tile_X4Y12_RegFile/FrameData[7] Tile_X4Y12_RegFile/FrameData[8] Tile_X4Y12_RegFile/FrameData[9]
+ Tile_X3Y12_LUT4AB/FrameStrobe[0] Tile_X3Y12_LUT4AB/FrameStrobe[10] Tile_X3Y12_LUT4AB/FrameStrobe[11]
+ Tile_X3Y12_LUT4AB/FrameStrobe[12] Tile_X3Y12_LUT4AB/FrameStrobe[13] Tile_X3Y12_LUT4AB/FrameStrobe[14]
+ Tile_X3Y12_LUT4AB/FrameStrobe[15] Tile_X3Y12_LUT4AB/FrameStrobe[16] Tile_X3Y12_LUT4AB/FrameStrobe[17]
+ Tile_X3Y12_LUT4AB/FrameStrobe[18] Tile_X3Y12_LUT4AB/FrameStrobe[19] Tile_X3Y12_LUT4AB/FrameStrobe[1]
+ Tile_X3Y12_LUT4AB/FrameStrobe[2] Tile_X3Y12_LUT4AB/FrameStrobe[3] Tile_X3Y12_LUT4AB/FrameStrobe[4]
+ Tile_X3Y12_LUT4AB/FrameStrobe[5] Tile_X3Y12_LUT4AB/FrameStrobe[6] Tile_X3Y12_LUT4AB/FrameStrobe[7]
+ Tile_X3Y12_LUT4AB/FrameStrobe[8] Tile_X3Y12_LUT4AB/FrameStrobe[9] Tile_X3Y11_LUT4AB/FrameStrobe[0]
+ Tile_X3Y11_LUT4AB/FrameStrobe[10] Tile_X3Y11_LUT4AB/FrameStrobe[11] Tile_X3Y11_LUT4AB/FrameStrobe[12]
+ Tile_X3Y11_LUT4AB/FrameStrobe[13] Tile_X3Y11_LUT4AB/FrameStrobe[14] Tile_X3Y11_LUT4AB/FrameStrobe[15]
+ Tile_X3Y11_LUT4AB/FrameStrobe[16] Tile_X3Y11_LUT4AB/FrameStrobe[17] Tile_X3Y11_LUT4AB/FrameStrobe[18]
+ Tile_X3Y11_LUT4AB/FrameStrobe[19] Tile_X3Y11_LUT4AB/FrameStrobe[1] Tile_X3Y11_LUT4AB/FrameStrobe[2]
+ Tile_X3Y11_LUT4AB/FrameStrobe[3] Tile_X3Y11_LUT4AB/FrameStrobe[4] Tile_X3Y11_LUT4AB/FrameStrobe[5]
+ Tile_X3Y11_LUT4AB/FrameStrobe[6] Tile_X3Y11_LUT4AB/FrameStrobe[7] Tile_X3Y11_LUT4AB/FrameStrobe[8]
+ Tile_X3Y11_LUT4AB/FrameStrobe[9] Tile_X3Y12_LUT4AB/N1BEG[0] Tile_X3Y12_LUT4AB/N1BEG[1]
+ Tile_X3Y12_LUT4AB/N1BEG[2] Tile_X3Y12_LUT4AB/N1BEG[3] Tile_X3Y13_LUT4AB/N1BEG[0]
+ Tile_X3Y13_LUT4AB/N1BEG[1] Tile_X3Y13_LUT4AB/N1BEG[2] Tile_X3Y13_LUT4AB/N1BEG[3]
+ Tile_X3Y12_LUT4AB/N2BEG[0] Tile_X3Y12_LUT4AB/N2BEG[1] Tile_X3Y12_LUT4AB/N2BEG[2]
+ Tile_X3Y12_LUT4AB/N2BEG[3] Tile_X3Y12_LUT4AB/N2BEG[4] Tile_X3Y12_LUT4AB/N2BEG[5]
+ Tile_X3Y12_LUT4AB/N2BEG[6] Tile_X3Y12_LUT4AB/N2BEG[7] Tile_X3Y11_LUT4AB/N2END[0]
+ Tile_X3Y11_LUT4AB/N2END[1] Tile_X3Y11_LUT4AB/N2END[2] Tile_X3Y11_LUT4AB/N2END[3]
+ Tile_X3Y11_LUT4AB/N2END[4] Tile_X3Y11_LUT4AB/N2END[5] Tile_X3Y11_LUT4AB/N2END[6]
+ Tile_X3Y11_LUT4AB/N2END[7] Tile_X3Y12_LUT4AB/N2END[0] Tile_X3Y12_LUT4AB/N2END[1]
+ Tile_X3Y12_LUT4AB/N2END[2] Tile_X3Y12_LUT4AB/N2END[3] Tile_X3Y12_LUT4AB/N2END[4]
+ Tile_X3Y12_LUT4AB/N2END[5] Tile_X3Y12_LUT4AB/N2END[6] Tile_X3Y12_LUT4AB/N2END[7]
+ Tile_X3Y13_LUT4AB/N2BEG[0] Tile_X3Y13_LUT4AB/N2BEG[1] Tile_X3Y13_LUT4AB/N2BEG[2]
+ Tile_X3Y13_LUT4AB/N2BEG[3] Tile_X3Y13_LUT4AB/N2BEG[4] Tile_X3Y13_LUT4AB/N2BEG[5]
+ Tile_X3Y13_LUT4AB/N2BEG[6] Tile_X3Y13_LUT4AB/N2BEG[7] Tile_X3Y12_LUT4AB/N4BEG[0]
+ Tile_X3Y12_LUT4AB/N4BEG[10] Tile_X3Y12_LUT4AB/N4BEG[11] Tile_X3Y12_LUT4AB/N4BEG[12]
+ Tile_X3Y12_LUT4AB/N4BEG[13] Tile_X3Y12_LUT4AB/N4BEG[14] Tile_X3Y12_LUT4AB/N4BEG[15]
+ Tile_X3Y12_LUT4AB/N4BEG[1] Tile_X3Y12_LUT4AB/N4BEG[2] Tile_X3Y12_LUT4AB/N4BEG[3]
+ Tile_X3Y12_LUT4AB/N4BEG[4] Tile_X3Y12_LUT4AB/N4BEG[5] Tile_X3Y12_LUT4AB/N4BEG[6]
+ Tile_X3Y12_LUT4AB/N4BEG[7] Tile_X3Y12_LUT4AB/N4BEG[8] Tile_X3Y12_LUT4AB/N4BEG[9]
+ Tile_X3Y13_LUT4AB/N4BEG[0] Tile_X3Y13_LUT4AB/N4BEG[10] Tile_X3Y13_LUT4AB/N4BEG[11]
+ Tile_X3Y13_LUT4AB/N4BEG[12] Tile_X3Y13_LUT4AB/N4BEG[13] Tile_X3Y13_LUT4AB/N4BEG[14]
+ Tile_X3Y13_LUT4AB/N4BEG[15] Tile_X3Y13_LUT4AB/N4BEG[1] Tile_X3Y13_LUT4AB/N4BEG[2]
+ Tile_X3Y13_LUT4AB/N4BEG[3] Tile_X3Y13_LUT4AB/N4BEG[4] Tile_X3Y13_LUT4AB/N4BEG[5]
+ Tile_X3Y13_LUT4AB/N4BEG[6] Tile_X3Y13_LUT4AB/N4BEG[7] Tile_X3Y13_LUT4AB/N4BEG[8]
+ Tile_X3Y13_LUT4AB/N4BEG[9] Tile_X3Y12_LUT4AB/NN4BEG[0] Tile_X3Y12_LUT4AB/NN4BEG[10]
+ Tile_X3Y12_LUT4AB/NN4BEG[11] Tile_X3Y12_LUT4AB/NN4BEG[12] Tile_X3Y12_LUT4AB/NN4BEG[13]
+ Tile_X3Y12_LUT4AB/NN4BEG[14] Tile_X3Y12_LUT4AB/NN4BEG[15] Tile_X3Y12_LUT4AB/NN4BEG[1]
+ Tile_X3Y12_LUT4AB/NN4BEG[2] Tile_X3Y12_LUT4AB/NN4BEG[3] Tile_X3Y12_LUT4AB/NN4BEG[4]
+ Tile_X3Y12_LUT4AB/NN4BEG[5] Tile_X3Y12_LUT4AB/NN4BEG[6] Tile_X3Y12_LUT4AB/NN4BEG[7]
+ Tile_X3Y12_LUT4AB/NN4BEG[8] Tile_X3Y12_LUT4AB/NN4BEG[9] Tile_X3Y13_LUT4AB/NN4BEG[0]
+ Tile_X3Y13_LUT4AB/NN4BEG[10] Tile_X3Y13_LUT4AB/NN4BEG[11] Tile_X3Y13_LUT4AB/NN4BEG[12]
+ Tile_X3Y13_LUT4AB/NN4BEG[13] Tile_X3Y13_LUT4AB/NN4BEG[14] Tile_X3Y13_LUT4AB/NN4BEG[15]
+ Tile_X3Y13_LUT4AB/NN4BEG[1] Tile_X3Y13_LUT4AB/NN4BEG[2] Tile_X3Y13_LUT4AB/NN4BEG[3]
+ Tile_X3Y13_LUT4AB/NN4BEG[4] Tile_X3Y13_LUT4AB/NN4BEG[5] Tile_X3Y13_LUT4AB/NN4BEG[6]
+ Tile_X3Y13_LUT4AB/NN4BEG[7] Tile_X3Y13_LUT4AB/NN4BEG[8] Tile_X3Y13_LUT4AB/NN4BEG[9]
+ Tile_X3Y13_LUT4AB/S1END[0] Tile_X3Y13_LUT4AB/S1END[1] Tile_X3Y13_LUT4AB/S1END[2]
+ Tile_X3Y13_LUT4AB/S1END[3] Tile_X3Y12_LUT4AB/S1END[0] Tile_X3Y12_LUT4AB/S1END[1]
+ Tile_X3Y12_LUT4AB/S1END[2] Tile_X3Y12_LUT4AB/S1END[3] Tile_X3Y13_LUT4AB/S2MID[0]
+ Tile_X3Y13_LUT4AB/S2MID[1] Tile_X3Y13_LUT4AB/S2MID[2] Tile_X3Y13_LUT4AB/S2MID[3]
+ Tile_X3Y13_LUT4AB/S2MID[4] Tile_X3Y13_LUT4AB/S2MID[5] Tile_X3Y13_LUT4AB/S2MID[6]
+ Tile_X3Y13_LUT4AB/S2MID[7] Tile_X3Y13_LUT4AB/S2END[0] Tile_X3Y13_LUT4AB/S2END[1]
+ Tile_X3Y13_LUT4AB/S2END[2] Tile_X3Y13_LUT4AB/S2END[3] Tile_X3Y13_LUT4AB/S2END[4]
+ Tile_X3Y13_LUT4AB/S2END[5] Tile_X3Y13_LUT4AB/S2END[6] Tile_X3Y13_LUT4AB/S2END[7]
+ Tile_X3Y12_LUT4AB/S2END[0] Tile_X3Y12_LUT4AB/S2END[1] Tile_X3Y12_LUT4AB/S2END[2]
+ Tile_X3Y12_LUT4AB/S2END[3] Tile_X3Y12_LUT4AB/S2END[4] Tile_X3Y12_LUT4AB/S2END[5]
+ Tile_X3Y12_LUT4AB/S2END[6] Tile_X3Y12_LUT4AB/S2END[7] Tile_X3Y12_LUT4AB/S2MID[0]
+ Tile_X3Y12_LUT4AB/S2MID[1] Tile_X3Y12_LUT4AB/S2MID[2] Tile_X3Y12_LUT4AB/S2MID[3]
+ Tile_X3Y12_LUT4AB/S2MID[4] Tile_X3Y12_LUT4AB/S2MID[5] Tile_X3Y12_LUT4AB/S2MID[6]
+ Tile_X3Y12_LUT4AB/S2MID[7] Tile_X3Y13_LUT4AB/S4END[0] Tile_X3Y13_LUT4AB/S4END[10]
+ Tile_X3Y13_LUT4AB/S4END[11] Tile_X3Y13_LUT4AB/S4END[12] Tile_X3Y13_LUT4AB/S4END[13]
+ Tile_X3Y13_LUT4AB/S4END[14] Tile_X3Y13_LUT4AB/S4END[15] Tile_X3Y13_LUT4AB/S4END[1]
+ Tile_X3Y13_LUT4AB/S4END[2] Tile_X3Y13_LUT4AB/S4END[3] Tile_X3Y13_LUT4AB/S4END[4]
+ Tile_X3Y13_LUT4AB/S4END[5] Tile_X3Y13_LUT4AB/S4END[6] Tile_X3Y13_LUT4AB/S4END[7]
+ Tile_X3Y13_LUT4AB/S4END[8] Tile_X3Y13_LUT4AB/S4END[9] Tile_X3Y12_LUT4AB/S4END[0]
+ Tile_X3Y12_LUT4AB/S4END[10] Tile_X3Y12_LUT4AB/S4END[11] Tile_X3Y12_LUT4AB/S4END[12]
+ Tile_X3Y12_LUT4AB/S4END[13] Tile_X3Y12_LUT4AB/S4END[14] Tile_X3Y12_LUT4AB/S4END[15]
+ Tile_X3Y12_LUT4AB/S4END[1] Tile_X3Y12_LUT4AB/S4END[2] Tile_X3Y12_LUT4AB/S4END[3]
+ Tile_X3Y12_LUT4AB/S4END[4] Tile_X3Y12_LUT4AB/S4END[5] Tile_X3Y12_LUT4AB/S4END[6]
+ Tile_X3Y12_LUT4AB/S4END[7] Tile_X3Y12_LUT4AB/S4END[8] Tile_X3Y12_LUT4AB/S4END[9]
+ Tile_X3Y13_LUT4AB/SS4END[0] Tile_X3Y13_LUT4AB/SS4END[10] Tile_X3Y13_LUT4AB/SS4END[11]
+ Tile_X3Y13_LUT4AB/SS4END[12] Tile_X3Y13_LUT4AB/SS4END[13] Tile_X3Y13_LUT4AB/SS4END[14]
+ Tile_X3Y13_LUT4AB/SS4END[15] Tile_X3Y13_LUT4AB/SS4END[1] Tile_X3Y13_LUT4AB/SS4END[2]
+ Tile_X3Y13_LUT4AB/SS4END[3] Tile_X3Y13_LUT4AB/SS4END[4] Tile_X3Y13_LUT4AB/SS4END[5]
+ Tile_X3Y13_LUT4AB/SS4END[6] Tile_X3Y13_LUT4AB/SS4END[7] Tile_X3Y13_LUT4AB/SS4END[8]
+ Tile_X3Y13_LUT4AB/SS4END[9] Tile_X3Y12_LUT4AB/SS4END[0] Tile_X3Y12_LUT4AB/SS4END[10]
+ Tile_X3Y12_LUT4AB/SS4END[11] Tile_X3Y12_LUT4AB/SS4END[12] Tile_X3Y12_LUT4AB/SS4END[13]
+ Tile_X3Y12_LUT4AB/SS4END[14] Tile_X3Y12_LUT4AB/SS4END[15] Tile_X3Y12_LUT4AB/SS4END[1]
+ Tile_X3Y12_LUT4AB/SS4END[2] Tile_X3Y12_LUT4AB/SS4END[3] Tile_X3Y12_LUT4AB/SS4END[4]
+ Tile_X3Y12_LUT4AB/SS4END[5] Tile_X3Y12_LUT4AB/SS4END[6] Tile_X3Y12_LUT4AB/SS4END[7]
+ Tile_X3Y12_LUT4AB/SS4END[8] Tile_X3Y12_LUT4AB/SS4END[9] Tile_X3Y12_LUT4AB/UserCLK
+ Tile_X3Y11_LUT4AB/UserCLK VGND VPWR Tile_X3Y12_LUT4AB/W1BEG[0] Tile_X3Y12_LUT4AB/W1BEG[1]
+ Tile_X3Y12_LUT4AB/W1BEG[2] Tile_X3Y12_LUT4AB/W1BEG[3] Tile_X3Y12_LUT4AB/W1END[0]
+ Tile_X3Y12_LUT4AB/W1END[1] Tile_X3Y12_LUT4AB/W1END[2] Tile_X3Y12_LUT4AB/W1END[3]
+ Tile_X3Y12_LUT4AB/W2BEG[0] Tile_X3Y12_LUT4AB/W2BEG[1] Tile_X3Y12_LUT4AB/W2BEG[2]
+ Tile_X3Y12_LUT4AB/W2BEG[3] Tile_X3Y12_LUT4AB/W2BEG[4] Tile_X3Y12_LUT4AB/W2BEG[5]
+ Tile_X3Y12_LUT4AB/W2BEG[6] Tile_X3Y12_LUT4AB/W2BEG[7] Tile_X2Y12_LUT4AB/W2END[0]
+ Tile_X2Y12_LUT4AB/W2END[1] Tile_X2Y12_LUT4AB/W2END[2] Tile_X2Y12_LUT4AB/W2END[3]
+ Tile_X2Y12_LUT4AB/W2END[4] Tile_X2Y12_LUT4AB/W2END[5] Tile_X2Y12_LUT4AB/W2END[6]
+ Tile_X2Y12_LUT4AB/W2END[7] Tile_X3Y12_LUT4AB/W2END[0] Tile_X3Y12_LUT4AB/W2END[1]
+ Tile_X3Y12_LUT4AB/W2END[2] Tile_X3Y12_LUT4AB/W2END[3] Tile_X3Y12_LUT4AB/W2END[4]
+ Tile_X3Y12_LUT4AB/W2END[5] Tile_X3Y12_LUT4AB/W2END[6] Tile_X3Y12_LUT4AB/W2END[7]
+ Tile_X3Y12_LUT4AB/W2MID[0] Tile_X3Y12_LUT4AB/W2MID[1] Tile_X3Y12_LUT4AB/W2MID[2]
+ Tile_X3Y12_LUT4AB/W2MID[3] Tile_X3Y12_LUT4AB/W2MID[4] Tile_X3Y12_LUT4AB/W2MID[5]
+ Tile_X3Y12_LUT4AB/W2MID[6] Tile_X3Y12_LUT4AB/W2MID[7] Tile_X3Y12_LUT4AB/W6BEG[0]
+ Tile_X3Y12_LUT4AB/W6BEG[10] Tile_X3Y12_LUT4AB/W6BEG[11] Tile_X3Y12_LUT4AB/W6BEG[1]
+ Tile_X3Y12_LUT4AB/W6BEG[2] Tile_X3Y12_LUT4AB/W6BEG[3] Tile_X3Y12_LUT4AB/W6BEG[4]
+ Tile_X3Y12_LUT4AB/W6BEG[5] Tile_X3Y12_LUT4AB/W6BEG[6] Tile_X3Y12_LUT4AB/W6BEG[7]
+ Tile_X3Y12_LUT4AB/W6BEG[8] Tile_X3Y12_LUT4AB/W6BEG[9] Tile_X3Y12_LUT4AB/W6END[0]
+ Tile_X3Y12_LUT4AB/W6END[10] Tile_X3Y12_LUT4AB/W6END[11] Tile_X3Y12_LUT4AB/W6END[1]
+ Tile_X3Y12_LUT4AB/W6END[2] Tile_X3Y12_LUT4AB/W6END[3] Tile_X3Y12_LUT4AB/W6END[4]
+ Tile_X3Y12_LUT4AB/W6END[5] Tile_X3Y12_LUT4AB/W6END[6] Tile_X3Y12_LUT4AB/W6END[7]
+ Tile_X3Y12_LUT4AB/W6END[8] Tile_X3Y12_LUT4AB/W6END[9] Tile_X3Y12_LUT4AB/WW4BEG[0]
+ Tile_X3Y12_LUT4AB/WW4BEG[10] Tile_X3Y12_LUT4AB/WW4BEG[11] Tile_X3Y12_LUT4AB/WW4BEG[12]
+ Tile_X3Y12_LUT4AB/WW4BEG[13] Tile_X3Y12_LUT4AB/WW4BEG[14] Tile_X3Y12_LUT4AB/WW4BEG[15]
+ Tile_X3Y12_LUT4AB/WW4BEG[1] Tile_X3Y12_LUT4AB/WW4BEG[2] Tile_X3Y12_LUT4AB/WW4BEG[3]
+ Tile_X3Y12_LUT4AB/WW4BEG[4] Tile_X3Y12_LUT4AB/WW4BEG[5] Tile_X3Y12_LUT4AB/WW4BEG[6]
+ Tile_X3Y12_LUT4AB/WW4BEG[7] Tile_X3Y12_LUT4AB/WW4BEG[8] Tile_X3Y12_LUT4AB/WW4BEG[9]
+ Tile_X3Y12_LUT4AB/WW4END[0] Tile_X3Y12_LUT4AB/WW4END[10] Tile_X3Y12_LUT4AB/WW4END[11]
+ Tile_X3Y12_LUT4AB/WW4END[12] Tile_X3Y12_LUT4AB/WW4END[13] Tile_X3Y12_LUT4AB/WW4END[14]
+ Tile_X3Y12_LUT4AB/WW4END[15] Tile_X3Y12_LUT4AB/WW4END[1] Tile_X3Y12_LUT4AB/WW4END[2]
+ Tile_X3Y12_LUT4AB/WW4END[3] Tile_X3Y12_LUT4AB/WW4END[4] Tile_X3Y12_LUT4AB/WW4END[5]
+ Tile_X3Y12_LUT4AB/WW4END[6] Tile_X3Y12_LUT4AB/WW4END[7] Tile_X3Y12_LUT4AB/WW4END[8]
+ Tile_X3Y12_LUT4AB/WW4END[9] LUT4AB
XTile_X0Y5_W_IO Tile_X0Y5_A_I_top Tile_X0Y5_A_O_top Tile_X0Y5_A_T_top Tile_X0Y5_A_config_C_bit0
+ Tile_X0Y5_A_config_C_bit1 Tile_X0Y5_A_config_C_bit2 Tile_X0Y5_A_config_C_bit3 Tile_X0Y5_B_I_top
+ Tile_X0Y5_B_O_top Tile_X0Y5_B_T_top Tile_X0Y5_B_config_C_bit0 Tile_X0Y5_B_config_C_bit1
+ Tile_X0Y5_B_config_C_bit2 Tile_X0Y5_B_config_C_bit3 Tile_X0Y5_W_IO/E1BEG[0] Tile_X0Y5_W_IO/E1BEG[1]
+ Tile_X0Y5_W_IO/E1BEG[2] Tile_X0Y5_W_IO/E1BEG[3] Tile_X0Y5_W_IO/E2BEG[0] Tile_X0Y5_W_IO/E2BEG[1]
+ Tile_X0Y5_W_IO/E2BEG[2] Tile_X0Y5_W_IO/E2BEG[3] Tile_X0Y5_W_IO/E2BEG[4] Tile_X0Y5_W_IO/E2BEG[5]
+ Tile_X0Y5_W_IO/E2BEG[6] Tile_X0Y5_W_IO/E2BEG[7] Tile_X0Y5_W_IO/E2BEGb[0] Tile_X0Y5_W_IO/E2BEGb[1]
+ Tile_X0Y5_W_IO/E2BEGb[2] Tile_X0Y5_W_IO/E2BEGb[3] Tile_X0Y5_W_IO/E2BEGb[4] Tile_X0Y5_W_IO/E2BEGb[5]
+ Tile_X0Y5_W_IO/E2BEGb[6] Tile_X0Y5_W_IO/E2BEGb[7] Tile_X0Y5_W_IO/E6BEG[0] Tile_X0Y5_W_IO/E6BEG[10]
+ Tile_X0Y5_W_IO/E6BEG[11] Tile_X0Y5_W_IO/E6BEG[1] Tile_X0Y5_W_IO/E6BEG[2] Tile_X0Y5_W_IO/E6BEG[3]
+ Tile_X0Y5_W_IO/E6BEG[4] Tile_X0Y5_W_IO/E6BEG[5] Tile_X0Y5_W_IO/E6BEG[6] Tile_X0Y5_W_IO/E6BEG[7]
+ Tile_X0Y5_W_IO/E6BEG[8] Tile_X0Y5_W_IO/E6BEG[9] Tile_X0Y5_W_IO/EE4BEG[0] Tile_X0Y5_W_IO/EE4BEG[10]
+ Tile_X0Y5_W_IO/EE4BEG[11] Tile_X0Y5_W_IO/EE4BEG[12] Tile_X0Y5_W_IO/EE4BEG[13] Tile_X0Y5_W_IO/EE4BEG[14]
+ Tile_X0Y5_W_IO/EE4BEG[15] Tile_X0Y5_W_IO/EE4BEG[1] Tile_X0Y5_W_IO/EE4BEG[2] Tile_X0Y5_W_IO/EE4BEG[3]
+ Tile_X0Y5_W_IO/EE4BEG[4] Tile_X0Y5_W_IO/EE4BEG[5] Tile_X0Y5_W_IO/EE4BEG[6] Tile_X0Y5_W_IO/EE4BEG[7]
+ Tile_X0Y5_W_IO/EE4BEG[8] Tile_X0Y5_W_IO/EE4BEG[9] FrameData[160] FrameData[170]
+ FrameData[171] FrameData[172] FrameData[173] FrameData[174] FrameData[175] FrameData[176]
+ FrameData[177] FrameData[178] FrameData[179] FrameData[161] FrameData[180] FrameData[181]
+ FrameData[182] FrameData[183] FrameData[184] FrameData[185] FrameData[186] FrameData[187]
+ FrameData[188] FrameData[189] FrameData[162] FrameData[190] FrameData[191] FrameData[163]
+ FrameData[164] FrameData[165] FrameData[166] FrameData[167] FrameData[168] FrameData[169]
+ Tile_X1Y5_LUT4AB/FrameData[0] Tile_X1Y5_LUT4AB/FrameData[10] Tile_X1Y5_LUT4AB/FrameData[11]
+ Tile_X1Y5_LUT4AB/FrameData[12] Tile_X1Y5_LUT4AB/FrameData[13] Tile_X1Y5_LUT4AB/FrameData[14]
+ Tile_X1Y5_LUT4AB/FrameData[15] Tile_X1Y5_LUT4AB/FrameData[16] Tile_X1Y5_LUT4AB/FrameData[17]
+ Tile_X1Y5_LUT4AB/FrameData[18] Tile_X1Y5_LUT4AB/FrameData[19] Tile_X1Y5_LUT4AB/FrameData[1]
+ Tile_X1Y5_LUT4AB/FrameData[20] Tile_X1Y5_LUT4AB/FrameData[21] Tile_X1Y5_LUT4AB/FrameData[22]
+ Tile_X1Y5_LUT4AB/FrameData[23] Tile_X1Y5_LUT4AB/FrameData[24] Tile_X1Y5_LUT4AB/FrameData[25]
+ Tile_X1Y5_LUT4AB/FrameData[26] Tile_X1Y5_LUT4AB/FrameData[27] Tile_X1Y5_LUT4AB/FrameData[28]
+ Tile_X1Y5_LUT4AB/FrameData[29] Tile_X1Y5_LUT4AB/FrameData[2] Tile_X1Y5_LUT4AB/FrameData[30]
+ Tile_X1Y5_LUT4AB/FrameData[31] Tile_X1Y5_LUT4AB/FrameData[3] Tile_X1Y5_LUT4AB/FrameData[4]
+ Tile_X1Y5_LUT4AB/FrameData[5] Tile_X1Y5_LUT4AB/FrameData[6] Tile_X1Y5_LUT4AB/FrameData[7]
+ Tile_X1Y5_LUT4AB/FrameData[8] Tile_X1Y5_LUT4AB/FrameData[9] Tile_X0Y5_W_IO/FrameStrobe[0]
+ Tile_X0Y5_W_IO/FrameStrobe[10] Tile_X0Y5_W_IO/FrameStrobe[11] Tile_X0Y5_W_IO/FrameStrobe[12]
+ Tile_X0Y5_W_IO/FrameStrobe[13] Tile_X0Y5_W_IO/FrameStrobe[14] Tile_X0Y5_W_IO/FrameStrobe[15]
+ Tile_X0Y5_W_IO/FrameStrobe[16] Tile_X0Y5_W_IO/FrameStrobe[17] Tile_X0Y5_W_IO/FrameStrobe[18]
+ Tile_X0Y5_W_IO/FrameStrobe[19] Tile_X0Y5_W_IO/FrameStrobe[1] Tile_X0Y5_W_IO/FrameStrobe[2]
+ Tile_X0Y5_W_IO/FrameStrobe[3] Tile_X0Y5_W_IO/FrameStrobe[4] Tile_X0Y5_W_IO/FrameStrobe[5]
+ Tile_X0Y5_W_IO/FrameStrobe[6] Tile_X0Y5_W_IO/FrameStrobe[7] Tile_X0Y5_W_IO/FrameStrobe[8]
+ Tile_X0Y5_W_IO/FrameStrobe[9] Tile_X0Y4_W_IO/FrameStrobe[0] Tile_X0Y4_W_IO/FrameStrobe[10]
+ Tile_X0Y4_W_IO/FrameStrobe[11] Tile_X0Y4_W_IO/FrameStrobe[12] Tile_X0Y4_W_IO/FrameStrobe[13]
+ Tile_X0Y4_W_IO/FrameStrobe[14] Tile_X0Y4_W_IO/FrameStrobe[15] Tile_X0Y4_W_IO/FrameStrobe[16]
+ Tile_X0Y4_W_IO/FrameStrobe[17] Tile_X0Y4_W_IO/FrameStrobe[18] Tile_X0Y4_W_IO/FrameStrobe[19]
+ Tile_X0Y4_W_IO/FrameStrobe[1] Tile_X0Y4_W_IO/FrameStrobe[2] Tile_X0Y4_W_IO/FrameStrobe[3]
+ Tile_X0Y4_W_IO/FrameStrobe[4] Tile_X0Y4_W_IO/FrameStrobe[5] Tile_X0Y4_W_IO/FrameStrobe[6]
+ Tile_X0Y4_W_IO/FrameStrobe[7] Tile_X0Y4_W_IO/FrameStrobe[8] Tile_X0Y4_W_IO/FrameStrobe[9]
+ Tile_X0Y5_W_IO/UserCLK Tile_X0Y4_W_IO/UserCLK VGND VPWR Tile_X0Y5_W_IO/W1END[0]
+ Tile_X0Y5_W_IO/W1END[1] Tile_X0Y5_W_IO/W1END[2] Tile_X0Y5_W_IO/W1END[3] Tile_X0Y5_W_IO/W2END[0]
+ Tile_X0Y5_W_IO/W2END[1] Tile_X0Y5_W_IO/W2END[2] Tile_X0Y5_W_IO/W2END[3] Tile_X0Y5_W_IO/W2END[4]
+ Tile_X0Y5_W_IO/W2END[5] Tile_X0Y5_W_IO/W2END[6] Tile_X0Y5_W_IO/W2END[7] Tile_X0Y5_W_IO/W2MID[0]
+ Tile_X0Y5_W_IO/W2MID[1] Tile_X0Y5_W_IO/W2MID[2] Tile_X0Y5_W_IO/W2MID[3] Tile_X0Y5_W_IO/W2MID[4]
+ Tile_X0Y5_W_IO/W2MID[5] Tile_X0Y5_W_IO/W2MID[6] Tile_X0Y5_W_IO/W2MID[7] Tile_X0Y5_W_IO/W6END[0]
+ Tile_X0Y5_W_IO/W6END[10] Tile_X0Y5_W_IO/W6END[11] Tile_X0Y5_W_IO/W6END[1] Tile_X0Y5_W_IO/W6END[2]
+ Tile_X0Y5_W_IO/W6END[3] Tile_X0Y5_W_IO/W6END[4] Tile_X0Y5_W_IO/W6END[5] Tile_X0Y5_W_IO/W6END[6]
+ Tile_X0Y5_W_IO/W6END[7] Tile_X0Y5_W_IO/W6END[8] Tile_X0Y5_W_IO/W6END[9] Tile_X0Y5_W_IO/WW4END[0]
+ Tile_X0Y5_W_IO/WW4END[10] Tile_X0Y5_W_IO/WW4END[11] Tile_X0Y5_W_IO/WW4END[12] Tile_X0Y5_W_IO/WW4END[13]
+ Tile_X0Y5_W_IO/WW4END[14] Tile_X0Y5_W_IO/WW4END[15] Tile_X0Y5_W_IO/WW4END[1] Tile_X0Y5_W_IO/WW4END[2]
+ Tile_X0Y5_W_IO/WW4END[3] Tile_X0Y5_W_IO/WW4END[4] Tile_X0Y5_W_IO/WW4END[5] Tile_X0Y5_W_IO/WW4END[6]
+ Tile_X0Y5_W_IO/WW4END[7] Tile_X0Y5_W_IO/WW4END[8] Tile_X0Y5_W_IO/WW4END[9] W_IO
XTile_X8Y0_N_term_single Tile_X8Y1_LUT4AB/Co Tile_X7Y0_N_term_DSP/FrameData_O[0] Tile_X7Y0_N_term_DSP/FrameData_O[10]
+ Tile_X7Y0_N_term_DSP/FrameData_O[11] Tile_X7Y0_N_term_DSP/FrameData_O[12] Tile_X7Y0_N_term_DSP/FrameData_O[13]
+ Tile_X7Y0_N_term_DSP/FrameData_O[14] Tile_X7Y0_N_term_DSP/FrameData_O[15] Tile_X7Y0_N_term_DSP/FrameData_O[16]
+ Tile_X7Y0_N_term_DSP/FrameData_O[17] Tile_X7Y0_N_term_DSP/FrameData_O[18] Tile_X7Y0_N_term_DSP/FrameData_O[19]
+ Tile_X7Y0_N_term_DSP/FrameData_O[1] Tile_X7Y0_N_term_DSP/FrameData_O[20] Tile_X7Y0_N_term_DSP/FrameData_O[21]
+ Tile_X7Y0_N_term_DSP/FrameData_O[22] Tile_X7Y0_N_term_DSP/FrameData_O[23] Tile_X7Y0_N_term_DSP/FrameData_O[24]
+ Tile_X7Y0_N_term_DSP/FrameData_O[25] Tile_X7Y0_N_term_DSP/FrameData_O[26] Tile_X7Y0_N_term_DSP/FrameData_O[27]
+ Tile_X7Y0_N_term_DSP/FrameData_O[28] Tile_X7Y0_N_term_DSP/FrameData_O[29] Tile_X7Y0_N_term_DSP/FrameData_O[2]
+ Tile_X7Y0_N_term_DSP/FrameData_O[30] Tile_X7Y0_N_term_DSP/FrameData_O[31] Tile_X7Y0_N_term_DSP/FrameData_O[3]
+ Tile_X7Y0_N_term_DSP/FrameData_O[4] Tile_X7Y0_N_term_DSP/FrameData_O[5] Tile_X7Y0_N_term_DSP/FrameData_O[6]
+ Tile_X7Y0_N_term_DSP/FrameData_O[7] Tile_X7Y0_N_term_DSP/FrameData_O[8] Tile_X7Y0_N_term_DSP/FrameData_O[9]
+ Tile_X9Y0_N_term_single/FrameData[0] Tile_X9Y0_N_term_single/FrameData[10] Tile_X9Y0_N_term_single/FrameData[11]
+ Tile_X9Y0_N_term_single/FrameData[12] Tile_X9Y0_N_term_single/FrameData[13] Tile_X9Y0_N_term_single/FrameData[14]
+ Tile_X9Y0_N_term_single/FrameData[15] Tile_X9Y0_N_term_single/FrameData[16] Tile_X9Y0_N_term_single/FrameData[17]
+ Tile_X9Y0_N_term_single/FrameData[18] Tile_X9Y0_N_term_single/FrameData[19] Tile_X9Y0_N_term_single/FrameData[1]
+ Tile_X9Y0_N_term_single/FrameData[20] Tile_X9Y0_N_term_single/FrameData[21] Tile_X9Y0_N_term_single/FrameData[22]
+ Tile_X9Y0_N_term_single/FrameData[23] Tile_X9Y0_N_term_single/FrameData[24] Tile_X9Y0_N_term_single/FrameData[25]
+ Tile_X9Y0_N_term_single/FrameData[26] Tile_X9Y0_N_term_single/FrameData[27] Tile_X9Y0_N_term_single/FrameData[28]
+ Tile_X9Y0_N_term_single/FrameData[29] Tile_X9Y0_N_term_single/FrameData[2] Tile_X9Y0_N_term_single/FrameData[30]
+ Tile_X9Y0_N_term_single/FrameData[31] Tile_X9Y0_N_term_single/FrameData[3] Tile_X9Y0_N_term_single/FrameData[4]
+ Tile_X9Y0_N_term_single/FrameData[5] Tile_X9Y0_N_term_single/FrameData[6] Tile_X9Y0_N_term_single/FrameData[7]
+ Tile_X9Y0_N_term_single/FrameData[8] Tile_X9Y0_N_term_single/FrameData[9] Tile_X8Y1_LUT4AB/FrameStrobe_O[0]
+ Tile_X8Y1_LUT4AB/FrameStrobe_O[10] Tile_X8Y1_LUT4AB/FrameStrobe_O[11] Tile_X8Y1_LUT4AB/FrameStrobe_O[12]
+ Tile_X8Y1_LUT4AB/FrameStrobe_O[13] Tile_X8Y1_LUT4AB/FrameStrobe_O[14] Tile_X8Y1_LUT4AB/FrameStrobe_O[15]
+ Tile_X8Y1_LUT4AB/FrameStrobe_O[16] Tile_X8Y1_LUT4AB/FrameStrobe_O[17] Tile_X8Y1_LUT4AB/FrameStrobe_O[18]
+ Tile_X8Y1_LUT4AB/FrameStrobe_O[19] Tile_X8Y1_LUT4AB/FrameStrobe_O[1] Tile_X8Y1_LUT4AB/FrameStrobe_O[2]
+ Tile_X8Y1_LUT4AB/FrameStrobe_O[3] Tile_X8Y1_LUT4AB/FrameStrobe_O[4] Tile_X8Y1_LUT4AB/FrameStrobe_O[5]
+ Tile_X8Y1_LUT4AB/FrameStrobe_O[6] Tile_X8Y1_LUT4AB/FrameStrobe_O[7] Tile_X8Y1_LUT4AB/FrameStrobe_O[8]
+ Tile_X8Y1_LUT4AB/FrameStrobe_O[9] Tile_X8Y0_N_term_single/FrameStrobe_O[0] Tile_X8Y0_N_term_single/FrameStrobe_O[10]
+ Tile_X8Y0_N_term_single/FrameStrobe_O[11] Tile_X8Y0_N_term_single/FrameStrobe_O[12]
+ Tile_X8Y0_N_term_single/FrameStrobe_O[13] Tile_X8Y0_N_term_single/FrameStrobe_O[14]
+ Tile_X8Y0_N_term_single/FrameStrobe_O[15] Tile_X8Y0_N_term_single/FrameStrobe_O[16]
+ Tile_X8Y0_N_term_single/FrameStrobe_O[17] Tile_X8Y0_N_term_single/FrameStrobe_O[18]
+ Tile_X8Y0_N_term_single/FrameStrobe_O[19] Tile_X8Y0_N_term_single/FrameStrobe_O[1]
+ Tile_X8Y0_N_term_single/FrameStrobe_O[2] Tile_X8Y0_N_term_single/FrameStrobe_O[3]
+ Tile_X8Y0_N_term_single/FrameStrobe_O[4] Tile_X8Y0_N_term_single/FrameStrobe_O[5]
+ Tile_X8Y0_N_term_single/FrameStrobe_O[6] Tile_X8Y0_N_term_single/FrameStrobe_O[7]
+ Tile_X8Y0_N_term_single/FrameStrobe_O[8] Tile_X8Y0_N_term_single/FrameStrobe_O[9]
+ Tile_X8Y1_LUT4AB/N1BEG[0] Tile_X8Y1_LUT4AB/N1BEG[1] Tile_X8Y1_LUT4AB/N1BEG[2] Tile_X8Y1_LUT4AB/N1BEG[3]
+ Tile_X8Y1_LUT4AB/N2BEGb[0] Tile_X8Y1_LUT4AB/N2BEGb[1] Tile_X8Y1_LUT4AB/N2BEGb[2]
+ Tile_X8Y1_LUT4AB/N2BEGb[3] Tile_X8Y1_LUT4AB/N2BEGb[4] Tile_X8Y1_LUT4AB/N2BEGb[5]
+ Tile_X8Y1_LUT4AB/N2BEGb[6] Tile_X8Y1_LUT4AB/N2BEGb[7] Tile_X8Y1_LUT4AB/N2BEG[0]
+ Tile_X8Y1_LUT4AB/N2BEG[1] Tile_X8Y1_LUT4AB/N2BEG[2] Tile_X8Y1_LUT4AB/N2BEG[3] Tile_X8Y1_LUT4AB/N2BEG[4]
+ Tile_X8Y1_LUT4AB/N2BEG[5] Tile_X8Y1_LUT4AB/N2BEG[6] Tile_X8Y1_LUT4AB/N2BEG[7] Tile_X8Y1_LUT4AB/N4BEG[0]
+ Tile_X8Y1_LUT4AB/N4BEG[10] Tile_X8Y1_LUT4AB/N4BEG[11] Tile_X8Y1_LUT4AB/N4BEG[12]
+ Tile_X8Y1_LUT4AB/N4BEG[13] Tile_X8Y1_LUT4AB/N4BEG[14] Tile_X8Y1_LUT4AB/N4BEG[15]
+ Tile_X8Y1_LUT4AB/N4BEG[1] Tile_X8Y1_LUT4AB/N4BEG[2] Tile_X8Y1_LUT4AB/N4BEG[3] Tile_X8Y1_LUT4AB/N4BEG[4]
+ Tile_X8Y1_LUT4AB/N4BEG[5] Tile_X8Y1_LUT4AB/N4BEG[6] Tile_X8Y1_LUT4AB/N4BEG[7] Tile_X8Y1_LUT4AB/N4BEG[8]
+ Tile_X8Y1_LUT4AB/N4BEG[9] Tile_X8Y1_LUT4AB/NN4BEG[0] Tile_X8Y1_LUT4AB/NN4BEG[10]
+ Tile_X8Y1_LUT4AB/NN4BEG[11] Tile_X8Y1_LUT4AB/NN4BEG[12] Tile_X8Y1_LUT4AB/NN4BEG[13]
+ Tile_X8Y1_LUT4AB/NN4BEG[14] Tile_X8Y1_LUT4AB/NN4BEG[15] Tile_X8Y1_LUT4AB/NN4BEG[1]
+ Tile_X8Y1_LUT4AB/NN4BEG[2] Tile_X8Y1_LUT4AB/NN4BEG[3] Tile_X8Y1_LUT4AB/NN4BEG[4]
+ Tile_X8Y1_LUT4AB/NN4BEG[5] Tile_X8Y1_LUT4AB/NN4BEG[6] Tile_X8Y1_LUT4AB/NN4BEG[7]
+ Tile_X8Y1_LUT4AB/NN4BEG[8] Tile_X8Y1_LUT4AB/NN4BEG[9] Tile_X8Y1_LUT4AB/S1END[0]
+ Tile_X8Y1_LUT4AB/S1END[1] Tile_X8Y1_LUT4AB/S1END[2] Tile_X8Y1_LUT4AB/S1END[3] Tile_X8Y1_LUT4AB/S2MID[0]
+ Tile_X8Y1_LUT4AB/S2MID[1] Tile_X8Y1_LUT4AB/S2MID[2] Tile_X8Y1_LUT4AB/S2MID[3] Tile_X8Y1_LUT4AB/S2MID[4]
+ Tile_X8Y1_LUT4AB/S2MID[5] Tile_X8Y1_LUT4AB/S2MID[6] Tile_X8Y1_LUT4AB/S2MID[7] Tile_X8Y1_LUT4AB/S2END[0]
+ Tile_X8Y1_LUT4AB/S2END[1] Tile_X8Y1_LUT4AB/S2END[2] Tile_X8Y1_LUT4AB/S2END[3] Tile_X8Y1_LUT4AB/S2END[4]
+ Tile_X8Y1_LUT4AB/S2END[5] Tile_X8Y1_LUT4AB/S2END[6] Tile_X8Y1_LUT4AB/S2END[7] Tile_X8Y1_LUT4AB/S4END[0]
+ Tile_X8Y1_LUT4AB/S4END[10] Tile_X8Y1_LUT4AB/S4END[11] Tile_X8Y1_LUT4AB/S4END[12]
+ Tile_X8Y1_LUT4AB/S4END[13] Tile_X8Y1_LUT4AB/S4END[14] Tile_X8Y1_LUT4AB/S4END[15]
+ Tile_X8Y1_LUT4AB/S4END[1] Tile_X8Y1_LUT4AB/S4END[2] Tile_X8Y1_LUT4AB/S4END[3] Tile_X8Y1_LUT4AB/S4END[4]
+ Tile_X8Y1_LUT4AB/S4END[5] Tile_X8Y1_LUT4AB/S4END[6] Tile_X8Y1_LUT4AB/S4END[7] Tile_X8Y1_LUT4AB/S4END[8]
+ Tile_X8Y1_LUT4AB/S4END[9] Tile_X8Y1_LUT4AB/SS4END[0] Tile_X8Y1_LUT4AB/SS4END[10]
+ Tile_X8Y1_LUT4AB/SS4END[11] Tile_X8Y1_LUT4AB/SS4END[12] Tile_X8Y1_LUT4AB/SS4END[13]
+ Tile_X8Y1_LUT4AB/SS4END[14] Tile_X8Y1_LUT4AB/SS4END[15] Tile_X8Y1_LUT4AB/SS4END[1]
+ Tile_X8Y1_LUT4AB/SS4END[2] Tile_X8Y1_LUT4AB/SS4END[3] Tile_X8Y1_LUT4AB/SS4END[4]
+ Tile_X8Y1_LUT4AB/SS4END[5] Tile_X8Y1_LUT4AB/SS4END[6] Tile_X8Y1_LUT4AB/SS4END[7]
+ Tile_X8Y1_LUT4AB/SS4END[8] Tile_X8Y1_LUT4AB/SS4END[9] Tile_X8Y1_LUT4AB/UserCLKo
+ Tile_X8Y0_N_term_single/UserCLKo VGND VPWR N_term_single
XTile_X10Y1_IHP_SRAM Tile_X10Y2_ADDR_SRAM0 Tile_X10Y2_ADDR_SRAM1 Tile_X10Y2_ADDR_SRAM2
+ Tile_X10Y2_ADDR_SRAM3 Tile_X10Y2_ADDR_SRAM4 Tile_X10Y2_ADDR_SRAM5 Tile_X10Y2_ADDR_SRAM6
+ Tile_X10Y2_ADDR_SRAM7 Tile_X10Y2_ADDR_SRAM8 Tile_X10Y2_ADDR_SRAM9 Tile_X10Y2_BM_SRAM0
+ Tile_X10Y2_BM_SRAM1 Tile_X10Y2_BM_SRAM10 Tile_X10Y2_BM_SRAM11 Tile_X10Y2_BM_SRAM12
+ Tile_X10Y2_BM_SRAM13 Tile_X10Y2_BM_SRAM14 Tile_X10Y2_BM_SRAM15 Tile_X10Y2_BM_SRAM16
+ Tile_X10Y2_BM_SRAM17 Tile_X10Y2_BM_SRAM18 Tile_X10Y2_BM_SRAM19 Tile_X10Y2_BM_SRAM2
+ Tile_X10Y2_BM_SRAM20 Tile_X10Y2_BM_SRAM21 Tile_X10Y2_BM_SRAM22 Tile_X10Y2_BM_SRAM23
+ Tile_X10Y2_BM_SRAM24 Tile_X10Y2_BM_SRAM25 Tile_X10Y2_BM_SRAM26 Tile_X10Y2_BM_SRAM27
+ Tile_X10Y2_BM_SRAM28 Tile_X10Y2_BM_SRAM29 Tile_X10Y2_BM_SRAM3 Tile_X10Y2_BM_SRAM30
+ Tile_X10Y2_BM_SRAM31 Tile_X10Y2_BM_SRAM4 Tile_X10Y2_BM_SRAM5 Tile_X10Y2_BM_SRAM6
+ Tile_X10Y2_BM_SRAM7 Tile_X10Y2_BM_SRAM8 Tile_X10Y2_BM_SRAM9 Tile_X10Y2_CLK_SRAM
+ Tile_X10Y2_CONFIGURED_top Tile_X10Y2_DIN_SRAM0 Tile_X10Y2_DIN_SRAM1 Tile_X10Y2_DIN_SRAM10
+ Tile_X10Y2_DIN_SRAM11 Tile_X10Y2_DIN_SRAM12 Tile_X10Y2_DIN_SRAM13 Tile_X10Y2_DIN_SRAM14
+ Tile_X10Y2_DIN_SRAM15 Tile_X10Y2_DIN_SRAM16 Tile_X10Y2_DIN_SRAM17 Tile_X10Y2_DIN_SRAM18
+ Tile_X10Y2_DIN_SRAM19 Tile_X10Y2_DIN_SRAM2 Tile_X10Y2_DIN_SRAM20 Tile_X10Y2_DIN_SRAM21
+ Tile_X10Y2_DIN_SRAM22 Tile_X10Y2_DIN_SRAM23 Tile_X10Y2_DIN_SRAM24 Tile_X10Y2_DIN_SRAM25
+ Tile_X10Y2_DIN_SRAM26 Tile_X10Y2_DIN_SRAM27 Tile_X10Y2_DIN_SRAM28 Tile_X10Y2_DIN_SRAM29
+ Tile_X10Y2_DIN_SRAM3 Tile_X10Y2_DIN_SRAM30 Tile_X10Y2_DIN_SRAM31 Tile_X10Y2_DIN_SRAM4
+ Tile_X10Y2_DIN_SRAM5 Tile_X10Y2_DIN_SRAM6 Tile_X10Y2_DIN_SRAM7 Tile_X10Y2_DIN_SRAM8
+ Tile_X10Y2_DIN_SRAM9 Tile_X10Y2_DOUT_SRAM0 Tile_X10Y2_DOUT_SRAM1 Tile_X10Y2_DOUT_SRAM10
+ Tile_X10Y2_DOUT_SRAM11 Tile_X10Y2_DOUT_SRAM12 Tile_X10Y2_DOUT_SRAM13 Tile_X10Y2_DOUT_SRAM14
+ Tile_X10Y2_DOUT_SRAM15 Tile_X10Y2_DOUT_SRAM16 Tile_X10Y2_DOUT_SRAM17 Tile_X10Y2_DOUT_SRAM18
+ Tile_X10Y2_DOUT_SRAM19 Tile_X10Y2_DOUT_SRAM2 Tile_X10Y2_DOUT_SRAM20 Tile_X10Y2_DOUT_SRAM21
+ Tile_X10Y2_DOUT_SRAM22 Tile_X10Y2_DOUT_SRAM23 Tile_X10Y2_DOUT_SRAM24 Tile_X10Y2_DOUT_SRAM25
+ Tile_X10Y2_DOUT_SRAM26 Tile_X10Y2_DOUT_SRAM27 Tile_X10Y2_DOUT_SRAM28 Tile_X10Y2_DOUT_SRAM29
+ Tile_X10Y2_DOUT_SRAM3 Tile_X10Y2_DOUT_SRAM30 Tile_X10Y2_DOUT_SRAM31 Tile_X10Y2_DOUT_SRAM4
+ Tile_X10Y2_DOUT_SRAM5 Tile_X10Y2_DOUT_SRAM6 Tile_X10Y2_DOUT_SRAM7 Tile_X10Y2_DOUT_SRAM8
+ Tile_X10Y2_DOUT_SRAM9 Tile_X10Y2_MEN_SRAM Tile_X10Y2_REN_SRAM Tile_X10Y2_TIE_HIGH_SRAM
+ Tile_X10Y2_TIE_LOW_SRAM Tile_X9Y1_LUT4AB/E1BEG[0] Tile_X9Y1_LUT4AB/E1BEG[1] Tile_X9Y1_LUT4AB/E1BEG[2]
+ Tile_X9Y1_LUT4AB/E1BEG[3] Tile_X9Y1_LUT4AB/E2BEGb[0] Tile_X9Y1_LUT4AB/E2BEGb[1]
+ Tile_X9Y1_LUT4AB/E2BEGb[2] Tile_X9Y1_LUT4AB/E2BEGb[3] Tile_X9Y1_LUT4AB/E2BEGb[4]
+ Tile_X9Y1_LUT4AB/E2BEGb[5] Tile_X9Y1_LUT4AB/E2BEGb[6] Tile_X9Y1_LUT4AB/E2BEGb[7]
+ Tile_X9Y1_LUT4AB/E2BEG[0] Tile_X9Y1_LUT4AB/E2BEG[1] Tile_X9Y1_LUT4AB/E2BEG[2] Tile_X9Y1_LUT4AB/E2BEG[3]
+ Tile_X9Y1_LUT4AB/E2BEG[4] Tile_X9Y1_LUT4AB/E2BEG[5] Tile_X9Y1_LUT4AB/E2BEG[6] Tile_X9Y1_LUT4AB/E2BEG[7]
+ Tile_X9Y1_LUT4AB/E6BEG[0] Tile_X9Y1_LUT4AB/E6BEG[10] Tile_X9Y1_LUT4AB/E6BEG[11]
+ Tile_X9Y1_LUT4AB/E6BEG[1] Tile_X9Y1_LUT4AB/E6BEG[2] Tile_X9Y1_LUT4AB/E6BEG[3] Tile_X9Y1_LUT4AB/E6BEG[4]
+ Tile_X9Y1_LUT4AB/E6BEG[5] Tile_X9Y1_LUT4AB/E6BEG[6] Tile_X9Y1_LUT4AB/E6BEG[7] Tile_X9Y1_LUT4AB/E6BEG[8]
+ Tile_X9Y1_LUT4AB/E6BEG[9] Tile_X9Y1_LUT4AB/EE4BEG[0] Tile_X9Y1_LUT4AB/EE4BEG[10]
+ Tile_X9Y1_LUT4AB/EE4BEG[11] Tile_X9Y1_LUT4AB/EE4BEG[12] Tile_X9Y1_LUT4AB/EE4BEG[13]
+ Tile_X9Y1_LUT4AB/EE4BEG[14] Tile_X9Y1_LUT4AB/EE4BEG[15] Tile_X9Y1_LUT4AB/EE4BEG[1]
+ Tile_X9Y1_LUT4AB/EE4BEG[2] Tile_X9Y1_LUT4AB/EE4BEG[3] Tile_X9Y1_LUT4AB/EE4BEG[4]
+ Tile_X9Y1_LUT4AB/EE4BEG[5] Tile_X9Y1_LUT4AB/EE4BEG[6] Tile_X9Y1_LUT4AB/EE4BEG[7]
+ Tile_X9Y1_LUT4AB/EE4BEG[8] Tile_X9Y1_LUT4AB/EE4BEG[9] Tile_X9Y1_LUT4AB/FrameData_O[0]
+ Tile_X9Y1_LUT4AB/FrameData_O[10] Tile_X9Y1_LUT4AB/FrameData_O[11] Tile_X9Y1_LUT4AB/FrameData_O[12]
+ Tile_X9Y1_LUT4AB/FrameData_O[13] Tile_X9Y1_LUT4AB/FrameData_O[14] Tile_X9Y1_LUT4AB/FrameData_O[15]
+ Tile_X9Y1_LUT4AB/FrameData_O[16] Tile_X9Y1_LUT4AB/FrameData_O[17] Tile_X9Y1_LUT4AB/FrameData_O[18]
+ Tile_X9Y1_LUT4AB/FrameData_O[19] Tile_X9Y1_LUT4AB/FrameData_O[1] Tile_X9Y1_LUT4AB/FrameData_O[20]
+ Tile_X9Y1_LUT4AB/FrameData_O[21] Tile_X9Y1_LUT4AB/FrameData_O[22] Tile_X9Y1_LUT4AB/FrameData_O[23]
+ Tile_X9Y1_LUT4AB/FrameData_O[24] Tile_X9Y1_LUT4AB/FrameData_O[25] Tile_X9Y1_LUT4AB/FrameData_O[26]
+ Tile_X9Y1_LUT4AB/FrameData_O[27] Tile_X9Y1_LUT4AB/FrameData_O[28] Tile_X9Y1_LUT4AB/FrameData_O[29]
+ Tile_X9Y1_LUT4AB/FrameData_O[2] Tile_X9Y1_LUT4AB/FrameData_O[30] Tile_X9Y1_LUT4AB/FrameData_O[31]
+ Tile_X9Y1_LUT4AB/FrameData_O[3] Tile_X9Y1_LUT4AB/FrameData_O[4] Tile_X9Y1_LUT4AB/FrameData_O[5]
+ Tile_X9Y1_LUT4AB/FrameData_O[6] Tile_X9Y1_LUT4AB/FrameData_O[7] Tile_X9Y1_LUT4AB/FrameData_O[8]
+ Tile_X9Y1_LUT4AB/FrameData_O[9] Tile_X10Y1_IHP_SRAM/Tile_X0Y0_FrameData_O[0] Tile_X10Y1_IHP_SRAM/Tile_X0Y0_FrameData_O[10]
+ Tile_X10Y1_IHP_SRAM/Tile_X0Y0_FrameData_O[11] Tile_X10Y1_IHP_SRAM/Tile_X0Y0_FrameData_O[12]
+ Tile_X10Y1_IHP_SRAM/Tile_X0Y0_FrameData_O[13] Tile_X10Y1_IHP_SRAM/Tile_X0Y0_FrameData_O[14]
+ Tile_X10Y1_IHP_SRAM/Tile_X0Y0_FrameData_O[15] Tile_X10Y1_IHP_SRAM/Tile_X0Y0_FrameData_O[16]
+ Tile_X10Y1_IHP_SRAM/Tile_X0Y0_FrameData_O[17] Tile_X10Y1_IHP_SRAM/Tile_X0Y0_FrameData_O[18]
+ Tile_X10Y1_IHP_SRAM/Tile_X0Y0_FrameData_O[19] Tile_X10Y1_IHP_SRAM/Tile_X0Y0_FrameData_O[1]
+ Tile_X10Y1_IHP_SRAM/Tile_X0Y0_FrameData_O[20] Tile_X10Y1_IHP_SRAM/Tile_X0Y0_FrameData_O[21]
+ Tile_X10Y1_IHP_SRAM/Tile_X0Y0_FrameData_O[22] Tile_X10Y1_IHP_SRAM/Tile_X0Y0_FrameData_O[23]
+ Tile_X10Y1_IHP_SRAM/Tile_X0Y0_FrameData_O[24] Tile_X10Y1_IHP_SRAM/Tile_X0Y0_FrameData_O[25]
+ Tile_X10Y1_IHP_SRAM/Tile_X0Y0_FrameData_O[26] Tile_X10Y1_IHP_SRAM/Tile_X0Y0_FrameData_O[27]
+ Tile_X10Y1_IHP_SRAM/Tile_X0Y0_FrameData_O[28] Tile_X10Y1_IHP_SRAM/Tile_X0Y0_FrameData_O[29]
+ Tile_X10Y1_IHP_SRAM/Tile_X0Y0_FrameData_O[2] Tile_X10Y1_IHP_SRAM/Tile_X0Y0_FrameData_O[30]
+ Tile_X10Y1_IHP_SRAM/Tile_X0Y0_FrameData_O[31] Tile_X10Y1_IHP_SRAM/Tile_X0Y0_FrameData_O[3]
+ Tile_X10Y1_IHP_SRAM/Tile_X0Y0_FrameData_O[4] Tile_X10Y1_IHP_SRAM/Tile_X0Y0_FrameData_O[5]
+ Tile_X10Y1_IHP_SRAM/Tile_X0Y0_FrameData_O[6] Tile_X10Y1_IHP_SRAM/Tile_X0Y0_FrameData_O[7]
+ Tile_X10Y1_IHP_SRAM/Tile_X0Y0_FrameData_O[8] Tile_X10Y1_IHP_SRAM/Tile_X0Y0_FrameData_O[9]
+ Tile_X10Y0_N_term_IHP_SRAM/FrameStrobe[0] Tile_X10Y0_N_term_IHP_SRAM/FrameStrobe[10]
+ Tile_X10Y0_N_term_IHP_SRAM/FrameStrobe[11] Tile_X10Y0_N_term_IHP_SRAM/FrameStrobe[12]
+ Tile_X10Y0_N_term_IHP_SRAM/FrameStrobe[13] Tile_X10Y0_N_term_IHP_SRAM/FrameStrobe[14]
+ Tile_X10Y0_N_term_IHP_SRAM/FrameStrobe[15] Tile_X10Y0_N_term_IHP_SRAM/FrameStrobe[16]
+ Tile_X10Y0_N_term_IHP_SRAM/FrameStrobe[17] Tile_X10Y0_N_term_IHP_SRAM/FrameStrobe[18]
+ Tile_X10Y0_N_term_IHP_SRAM/FrameStrobe[19] Tile_X10Y0_N_term_IHP_SRAM/FrameStrobe[1]
+ Tile_X10Y0_N_term_IHP_SRAM/FrameStrobe[2] Tile_X10Y0_N_term_IHP_SRAM/FrameStrobe[3]
+ Tile_X10Y0_N_term_IHP_SRAM/FrameStrobe[4] Tile_X10Y0_N_term_IHP_SRAM/FrameStrobe[5]
+ Tile_X10Y0_N_term_IHP_SRAM/FrameStrobe[6] Tile_X10Y0_N_term_IHP_SRAM/FrameStrobe[7]
+ Tile_X10Y0_N_term_IHP_SRAM/FrameStrobe[8] Tile_X10Y0_N_term_IHP_SRAM/FrameStrobe[9]
+ Tile_X10Y0_N_term_IHP_SRAM/N1END[0] Tile_X10Y0_N_term_IHP_SRAM/N1END[1] Tile_X10Y0_N_term_IHP_SRAM/N1END[2]
+ Tile_X10Y0_N_term_IHP_SRAM/N1END[3] Tile_X10Y0_N_term_IHP_SRAM/N2MID[0] Tile_X10Y0_N_term_IHP_SRAM/N2MID[1]
+ Tile_X10Y0_N_term_IHP_SRAM/N2MID[2] Tile_X10Y0_N_term_IHP_SRAM/N2MID[3] Tile_X10Y0_N_term_IHP_SRAM/N2MID[4]
+ Tile_X10Y0_N_term_IHP_SRAM/N2MID[5] Tile_X10Y0_N_term_IHP_SRAM/N2MID[6] Tile_X10Y0_N_term_IHP_SRAM/N2MID[7]
+ Tile_X10Y0_N_term_IHP_SRAM/N2END[0] Tile_X10Y0_N_term_IHP_SRAM/N2END[1] Tile_X10Y0_N_term_IHP_SRAM/N2END[2]
+ Tile_X10Y0_N_term_IHP_SRAM/N2END[3] Tile_X10Y0_N_term_IHP_SRAM/N2END[4] Tile_X10Y0_N_term_IHP_SRAM/N2END[5]
+ Tile_X10Y0_N_term_IHP_SRAM/N2END[6] Tile_X10Y0_N_term_IHP_SRAM/N2END[7] Tile_X10Y0_N_term_IHP_SRAM/N4END[0]
+ Tile_X10Y0_N_term_IHP_SRAM/N4END[10] Tile_X10Y0_N_term_IHP_SRAM/N4END[11] Tile_X10Y0_N_term_IHP_SRAM/N4END[12]
+ Tile_X10Y0_N_term_IHP_SRAM/N4END[13] Tile_X10Y0_N_term_IHP_SRAM/N4END[14] Tile_X10Y0_N_term_IHP_SRAM/N4END[15]
+ Tile_X10Y0_N_term_IHP_SRAM/N4END[1] Tile_X10Y0_N_term_IHP_SRAM/N4END[2] Tile_X10Y0_N_term_IHP_SRAM/N4END[3]
+ Tile_X10Y0_N_term_IHP_SRAM/N4END[4] Tile_X10Y0_N_term_IHP_SRAM/N4END[5] Tile_X10Y0_N_term_IHP_SRAM/N4END[6]
+ Tile_X10Y0_N_term_IHP_SRAM/N4END[7] Tile_X10Y0_N_term_IHP_SRAM/N4END[8] Tile_X10Y0_N_term_IHP_SRAM/N4END[9]
+ Tile_X10Y0_N_term_IHP_SRAM/S1BEG[0] Tile_X10Y0_N_term_IHP_SRAM/S1BEG[1] Tile_X10Y0_N_term_IHP_SRAM/S1BEG[2]
+ Tile_X10Y0_N_term_IHP_SRAM/S1BEG[3] Tile_X10Y0_N_term_IHP_SRAM/S2BEGb[0] Tile_X10Y0_N_term_IHP_SRAM/S2BEGb[1]
+ Tile_X10Y0_N_term_IHP_SRAM/S2BEGb[2] Tile_X10Y0_N_term_IHP_SRAM/S2BEGb[3] Tile_X10Y0_N_term_IHP_SRAM/S2BEGb[4]
+ Tile_X10Y0_N_term_IHP_SRAM/S2BEGb[5] Tile_X10Y0_N_term_IHP_SRAM/S2BEGb[6] Tile_X10Y0_N_term_IHP_SRAM/S2BEGb[7]
+ Tile_X10Y0_N_term_IHP_SRAM/S2BEG[0] Tile_X10Y0_N_term_IHP_SRAM/S2BEG[1] Tile_X10Y0_N_term_IHP_SRAM/S2BEG[2]
+ Tile_X10Y0_N_term_IHP_SRAM/S2BEG[3] Tile_X10Y0_N_term_IHP_SRAM/S2BEG[4] Tile_X10Y0_N_term_IHP_SRAM/S2BEG[5]
+ Tile_X10Y0_N_term_IHP_SRAM/S2BEG[6] Tile_X10Y0_N_term_IHP_SRAM/S2BEG[7] Tile_X10Y0_N_term_IHP_SRAM/S4BEG[0]
+ Tile_X10Y0_N_term_IHP_SRAM/S4BEG[10] Tile_X10Y0_N_term_IHP_SRAM/S4BEG[11] Tile_X10Y0_N_term_IHP_SRAM/S4BEG[12]
+ Tile_X10Y0_N_term_IHP_SRAM/S4BEG[13] Tile_X10Y0_N_term_IHP_SRAM/S4BEG[14] Tile_X10Y0_N_term_IHP_SRAM/S4BEG[15]
+ Tile_X10Y0_N_term_IHP_SRAM/S4BEG[1] Tile_X10Y0_N_term_IHP_SRAM/S4BEG[2] Tile_X10Y0_N_term_IHP_SRAM/S4BEG[3]
+ Tile_X10Y0_N_term_IHP_SRAM/S4BEG[4] Tile_X10Y0_N_term_IHP_SRAM/S4BEG[5] Tile_X10Y0_N_term_IHP_SRAM/S4BEG[6]
+ Tile_X10Y0_N_term_IHP_SRAM/S4BEG[7] Tile_X10Y0_N_term_IHP_SRAM/S4BEG[8] Tile_X10Y0_N_term_IHP_SRAM/S4BEG[9]
+ Tile_X10Y0_N_term_IHP_SRAM/UserCLK Tile_X9Y1_LUT4AB/W1END[0] Tile_X9Y1_LUT4AB/W1END[1]
+ Tile_X9Y1_LUT4AB/W1END[2] Tile_X9Y1_LUT4AB/W1END[3] Tile_X9Y1_LUT4AB/W2MID[0] Tile_X9Y1_LUT4AB/W2MID[1]
+ Tile_X9Y1_LUT4AB/W2MID[2] Tile_X9Y1_LUT4AB/W2MID[3] Tile_X9Y1_LUT4AB/W2MID[4] Tile_X9Y1_LUT4AB/W2MID[5]
+ Tile_X9Y1_LUT4AB/W2MID[6] Tile_X9Y1_LUT4AB/W2MID[7] Tile_X9Y1_LUT4AB/W2END[0] Tile_X9Y1_LUT4AB/W2END[1]
+ Tile_X9Y1_LUT4AB/W2END[2] Tile_X9Y1_LUT4AB/W2END[3] Tile_X9Y1_LUT4AB/W2END[4] Tile_X9Y1_LUT4AB/W2END[5]
+ Tile_X9Y1_LUT4AB/W2END[6] Tile_X9Y1_LUT4AB/W2END[7] Tile_X9Y1_LUT4AB/W6END[0] Tile_X9Y1_LUT4AB/W6END[10]
+ Tile_X9Y1_LUT4AB/W6END[11] Tile_X9Y1_LUT4AB/W6END[1] Tile_X9Y1_LUT4AB/W6END[2] Tile_X9Y1_LUT4AB/W6END[3]
+ Tile_X9Y1_LUT4AB/W6END[4] Tile_X9Y1_LUT4AB/W6END[5] Tile_X9Y1_LUT4AB/W6END[6] Tile_X9Y1_LUT4AB/W6END[7]
+ Tile_X9Y1_LUT4AB/W6END[8] Tile_X9Y1_LUT4AB/W6END[9] Tile_X9Y1_LUT4AB/WW4END[0] Tile_X9Y1_LUT4AB/WW4END[10]
+ Tile_X9Y1_LUT4AB/WW4END[11] Tile_X9Y1_LUT4AB/WW4END[12] Tile_X9Y1_LUT4AB/WW4END[13]
+ Tile_X9Y1_LUT4AB/WW4END[14] Tile_X9Y1_LUT4AB/WW4END[15] Tile_X9Y1_LUT4AB/WW4END[1]
+ Tile_X9Y1_LUT4AB/WW4END[2] Tile_X9Y1_LUT4AB/WW4END[3] Tile_X9Y1_LUT4AB/WW4END[4]
+ Tile_X9Y1_LUT4AB/WW4END[5] Tile_X9Y1_LUT4AB/WW4END[6] Tile_X9Y1_LUT4AB/WW4END[7]
+ Tile_X9Y1_LUT4AB/WW4END[8] Tile_X9Y1_LUT4AB/WW4END[9] Tile_X9Y2_LUT4AB/E1BEG[0]
+ Tile_X9Y2_LUT4AB/E1BEG[1] Tile_X9Y2_LUT4AB/E1BEG[2] Tile_X9Y2_LUT4AB/E1BEG[3] Tile_X9Y2_LUT4AB/E2BEGb[0]
+ Tile_X9Y2_LUT4AB/E2BEGb[1] Tile_X9Y2_LUT4AB/E2BEGb[2] Tile_X9Y2_LUT4AB/E2BEGb[3]
+ Tile_X9Y2_LUT4AB/E2BEGb[4] Tile_X9Y2_LUT4AB/E2BEGb[5] Tile_X9Y2_LUT4AB/E2BEGb[6]
+ Tile_X9Y2_LUT4AB/E2BEGb[7] Tile_X9Y2_LUT4AB/E2BEG[0] Tile_X9Y2_LUT4AB/E2BEG[1] Tile_X9Y2_LUT4AB/E2BEG[2]
+ Tile_X9Y2_LUT4AB/E2BEG[3] Tile_X9Y2_LUT4AB/E2BEG[4] Tile_X9Y2_LUT4AB/E2BEG[5] Tile_X9Y2_LUT4AB/E2BEG[6]
+ Tile_X9Y2_LUT4AB/E2BEG[7] Tile_X9Y2_LUT4AB/E6BEG[0] Tile_X9Y2_LUT4AB/E6BEG[10] Tile_X9Y2_LUT4AB/E6BEG[11]
+ Tile_X9Y2_LUT4AB/E6BEG[1] Tile_X9Y2_LUT4AB/E6BEG[2] Tile_X9Y2_LUT4AB/E6BEG[3] Tile_X9Y2_LUT4AB/E6BEG[4]
+ Tile_X9Y2_LUT4AB/E6BEG[5] Tile_X9Y2_LUT4AB/E6BEG[6] Tile_X9Y2_LUT4AB/E6BEG[7] Tile_X9Y2_LUT4AB/E6BEG[8]
+ Tile_X9Y2_LUT4AB/E6BEG[9] Tile_X9Y2_LUT4AB/EE4BEG[0] Tile_X9Y2_LUT4AB/EE4BEG[10]
+ Tile_X9Y2_LUT4AB/EE4BEG[11] Tile_X9Y2_LUT4AB/EE4BEG[12] Tile_X9Y2_LUT4AB/EE4BEG[13]
+ Tile_X9Y2_LUT4AB/EE4BEG[14] Tile_X9Y2_LUT4AB/EE4BEG[15] Tile_X9Y2_LUT4AB/EE4BEG[1]
+ Tile_X9Y2_LUT4AB/EE4BEG[2] Tile_X9Y2_LUT4AB/EE4BEG[3] Tile_X9Y2_LUT4AB/EE4BEG[4]
+ Tile_X9Y2_LUT4AB/EE4BEG[5] Tile_X9Y2_LUT4AB/EE4BEG[6] Tile_X9Y2_LUT4AB/EE4BEG[7]
+ Tile_X9Y2_LUT4AB/EE4BEG[8] Tile_X9Y2_LUT4AB/EE4BEG[9] Tile_X9Y2_LUT4AB/FrameData_O[0]
+ Tile_X9Y2_LUT4AB/FrameData_O[10] Tile_X9Y2_LUT4AB/FrameData_O[11] Tile_X9Y2_LUT4AB/FrameData_O[12]
+ Tile_X9Y2_LUT4AB/FrameData_O[13] Tile_X9Y2_LUT4AB/FrameData_O[14] Tile_X9Y2_LUT4AB/FrameData_O[15]
+ Tile_X9Y2_LUT4AB/FrameData_O[16] Tile_X9Y2_LUT4AB/FrameData_O[17] Tile_X9Y2_LUT4AB/FrameData_O[18]
+ Tile_X9Y2_LUT4AB/FrameData_O[19] Tile_X9Y2_LUT4AB/FrameData_O[1] Tile_X9Y2_LUT4AB/FrameData_O[20]
+ Tile_X9Y2_LUT4AB/FrameData_O[21] Tile_X9Y2_LUT4AB/FrameData_O[22] Tile_X9Y2_LUT4AB/FrameData_O[23]
+ Tile_X9Y2_LUT4AB/FrameData_O[24] Tile_X9Y2_LUT4AB/FrameData_O[25] Tile_X9Y2_LUT4AB/FrameData_O[26]
+ Tile_X9Y2_LUT4AB/FrameData_O[27] Tile_X9Y2_LUT4AB/FrameData_O[28] Tile_X9Y2_LUT4AB/FrameData_O[29]
+ Tile_X9Y2_LUT4AB/FrameData_O[2] Tile_X9Y2_LUT4AB/FrameData_O[30] Tile_X9Y2_LUT4AB/FrameData_O[31]
+ Tile_X9Y2_LUT4AB/FrameData_O[3] Tile_X9Y2_LUT4AB/FrameData_O[4] Tile_X9Y2_LUT4AB/FrameData_O[5]
+ Tile_X9Y2_LUT4AB/FrameData_O[6] Tile_X9Y2_LUT4AB/FrameData_O[7] Tile_X9Y2_LUT4AB/FrameData_O[8]
+ Tile_X9Y2_LUT4AB/FrameData_O[9] Tile_X10Y1_IHP_SRAM/Tile_X0Y1_FrameData_O[0] Tile_X10Y1_IHP_SRAM/Tile_X0Y1_FrameData_O[10]
+ Tile_X10Y1_IHP_SRAM/Tile_X0Y1_FrameData_O[11] Tile_X10Y1_IHP_SRAM/Tile_X0Y1_FrameData_O[12]
+ Tile_X10Y1_IHP_SRAM/Tile_X0Y1_FrameData_O[13] Tile_X10Y1_IHP_SRAM/Tile_X0Y1_FrameData_O[14]
+ Tile_X10Y1_IHP_SRAM/Tile_X0Y1_FrameData_O[15] Tile_X10Y1_IHP_SRAM/Tile_X0Y1_FrameData_O[16]
+ Tile_X10Y1_IHP_SRAM/Tile_X0Y1_FrameData_O[17] Tile_X10Y1_IHP_SRAM/Tile_X0Y1_FrameData_O[18]
+ Tile_X10Y1_IHP_SRAM/Tile_X0Y1_FrameData_O[19] Tile_X10Y1_IHP_SRAM/Tile_X0Y1_FrameData_O[1]
+ Tile_X10Y1_IHP_SRAM/Tile_X0Y1_FrameData_O[20] Tile_X10Y1_IHP_SRAM/Tile_X0Y1_FrameData_O[21]
+ Tile_X10Y1_IHP_SRAM/Tile_X0Y1_FrameData_O[22] Tile_X10Y1_IHP_SRAM/Tile_X0Y1_FrameData_O[23]
+ Tile_X10Y1_IHP_SRAM/Tile_X0Y1_FrameData_O[24] Tile_X10Y1_IHP_SRAM/Tile_X0Y1_FrameData_O[25]
+ Tile_X10Y1_IHP_SRAM/Tile_X0Y1_FrameData_O[26] Tile_X10Y1_IHP_SRAM/Tile_X0Y1_FrameData_O[27]
+ Tile_X10Y1_IHP_SRAM/Tile_X0Y1_FrameData_O[28] Tile_X10Y1_IHP_SRAM/Tile_X0Y1_FrameData_O[29]
+ Tile_X10Y1_IHP_SRAM/Tile_X0Y1_FrameData_O[2] Tile_X10Y1_IHP_SRAM/Tile_X0Y1_FrameData_O[30]
+ Tile_X10Y1_IHP_SRAM/Tile_X0Y1_FrameData_O[31] Tile_X10Y1_IHP_SRAM/Tile_X0Y1_FrameData_O[3]
+ Tile_X10Y1_IHP_SRAM/Tile_X0Y1_FrameData_O[4] Tile_X10Y1_IHP_SRAM/Tile_X0Y1_FrameData_O[5]
+ Tile_X10Y1_IHP_SRAM/Tile_X0Y1_FrameData_O[6] Tile_X10Y1_IHP_SRAM/Tile_X0Y1_FrameData_O[7]
+ Tile_X10Y1_IHP_SRAM/Tile_X0Y1_FrameData_O[8] Tile_X10Y1_IHP_SRAM/Tile_X0Y1_FrameData_O[9]
+ Tile_X10Y1_IHP_SRAM/Tile_X0Y1_FrameStrobe[0] Tile_X10Y1_IHP_SRAM/Tile_X0Y1_FrameStrobe[10]
+ Tile_X10Y1_IHP_SRAM/Tile_X0Y1_FrameStrobe[11] Tile_X10Y1_IHP_SRAM/Tile_X0Y1_FrameStrobe[12]
+ Tile_X10Y1_IHP_SRAM/Tile_X0Y1_FrameStrobe[13] Tile_X10Y1_IHP_SRAM/Tile_X0Y1_FrameStrobe[14]
+ Tile_X10Y1_IHP_SRAM/Tile_X0Y1_FrameStrobe[15] Tile_X10Y1_IHP_SRAM/Tile_X0Y1_FrameStrobe[16]
+ Tile_X10Y1_IHP_SRAM/Tile_X0Y1_FrameStrobe[17] Tile_X10Y1_IHP_SRAM/Tile_X0Y1_FrameStrobe[18]
+ Tile_X10Y1_IHP_SRAM/Tile_X0Y1_FrameStrobe[19] Tile_X10Y1_IHP_SRAM/Tile_X0Y1_FrameStrobe[1]
+ Tile_X10Y1_IHP_SRAM/Tile_X0Y1_FrameStrobe[2] Tile_X10Y1_IHP_SRAM/Tile_X0Y1_FrameStrobe[3]
+ Tile_X10Y1_IHP_SRAM/Tile_X0Y1_FrameStrobe[4] Tile_X10Y1_IHP_SRAM/Tile_X0Y1_FrameStrobe[5]
+ Tile_X10Y1_IHP_SRAM/Tile_X0Y1_FrameStrobe[6] Tile_X10Y1_IHP_SRAM/Tile_X0Y1_FrameStrobe[7]
+ Tile_X10Y1_IHP_SRAM/Tile_X0Y1_FrameStrobe[8] Tile_X10Y1_IHP_SRAM/Tile_X0Y1_FrameStrobe[9]
+ Tile_X10Y3_IHP_SRAM/Tile_X0Y0_N1BEG[0] Tile_X10Y3_IHP_SRAM/Tile_X0Y0_N1BEG[1] Tile_X10Y3_IHP_SRAM/Tile_X0Y0_N1BEG[2]
+ Tile_X10Y3_IHP_SRAM/Tile_X0Y0_N1BEG[3] Tile_X10Y1_IHP_SRAM/Tile_X0Y1_N2END[0] Tile_X10Y1_IHP_SRAM/Tile_X0Y1_N2END[1]
+ Tile_X10Y1_IHP_SRAM/Tile_X0Y1_N2END[2] Tile_X10Y1_IHP_SRAM/Tile_X0Y1_N2END[3] Tile_X10Y1_IHP_SRAM/Tile_X0Y1_N2END[4]
+ Tile_X10Y1_IHP_SRAM/Tile_X0Y1_N2END[5] Tile_X10Y1_IHP_SRAM/Tile_X0Y1_N2END[6] Tile_X10Y1_IHP_SRAM/Tile_X0Y1_N2END[7]
+ Tile_X10Y3_IHP_SRAM/Tile_X0Y0_N2BEG[0] Tile_X10Y3_IHP_SRAM/Tile_X0Y0_N2BEG[1] Tile_X10Y3_IHP_SRAM/Tile_X0Y0_N2BEG[2]
+ Tile_X10Y3_IHP_SRAM/Tile_X0Y0_N2BEG[3] Tile_X10Y3_IHP_SRAM/Tile_X0Y0_N2BEG[4] Tile_X10Y3_IHP_SRAM/Tile_X0Y0_N2BEG[5]
+ Tile_X10Y3_IHP_SRAM/Tile_X0Y0_N2BEG[6] Tile_X10Y3_IHP_SRAM/Tile_X0Y0_N2BEG[7] Tile_X10Y3_IHP_SRAM/Tile_X0Y0_N4BEG[0]
+ Tile_X10Y3_IHP_SRAM/Tile_X0Y0_N4BEG[10] Tile_X10Y3_IHP_SRAM/Tile_X0Y0_N4BEG[11]
+ Tile_X10Y3_IHP_SRAM/Tile_X0Y0_N4BEG[12] Tile_X10Y3_IHP_SRAM/Tile_X0Y0_N4BEG[13]
+ Tile_X10Y3_IHP_SRAM/Tile_X0Y0_N4BEG[14] Tile_X10Y3_IHP_SRAM/Tile_X0Y0_N4BEG[15]
+ Tile_X10Y3_IHP_SRAM/Tile_X0Y0_N4BEG[1] Tile_X10Y3_IHP_SRAM/Tile_X0Y0_N4BEG[2] Tile_X10Y3_IHP_SRAM/Tile_X0Y0_N4BEG[3]
+ Tile_X10Y3_IHP_SRAM/Tile_X0Y0_N4BEG[4] Tile_X10Y3_IHP_SRAM/Tile_X0Y0_N4BEG[5] Tile_X10Y3_IHP_SRAM/Tile_X0Y0_N4BEG[6]
+ Tile_X10Y3_IHP_SRAM/Tile_X0Y0_N4BEG[7] Tile_X10Y3_IHP_SRAM/Tile_X0Y0_N4BEG[8] Tile_X10Y3_IHP_SRAM/Tile_X0Y0_N4BEG[9]
+ Tile_X10Y3_IHP_SRAM/Tile_X0Y0_S1END[0] Tile_X10Y3_IHP_SRAM/Tile_X0Y0_S1END[1] Tile_X10Y3_IHP_SRAM/Tile_X0Y0_S1END[2]
+ Tile_X10Y3_IHP_SRAM/Tile_X0Y0_S1END[3] Tile_X10Y3_IHP_SRAM/Tile_X0Y0_S2MID[0] Tile_X10Y3_IHP_SRAM/Tile_X0Y0_S2MID[1]
+ Tile_X10Y3_IHP_SRAM/Tile_X0Y0_S2MID[2] Tile_X10Y3_IHP_SRAM/Tile_X0Y0_S2MID[3] Tile_X10Y3_IHP_SRAM/Tile_X0Y0_S2MID[4]
+ Tile_X10Y3_IHP_SRAM/Tile_X0Y0_S2MID[5] Tile_X10Y3_IHP_SRAM/Tile_X0Y0_S2MID[6] Tile_X10Y3_IHP_SRAM/Tile_X0Y0_S2MID[7]
+ Tile_X10Y3_IHP_SRAM/Tile_X0Y0_S2END[0] Tile_X10Y3_IHP_SRAM/Tile_X0Y0_S2END[1] Tile_X10Y3_IHP_SRAM/Tile_X0Y0_S2END[2]
+ Tile_X10Y3_IHP_SRAM/Tile_X0Y0_S2END[3] Tile_X10Y3_IHP_SRAM/Tile_X0Y0_S2END[4] Tile_X10Y3_IHP_SRAM/Tile_X0Y0_S2END[5]
+ Tile_X10Y3_IHP_SRAM/Tile_X0Y0_S2END[6] Tile_X10Y3_IHP_SRAM/Tile_X0Y0_S2END[7] Tile_X10Y3_IHP_SRAM/Tile_X0Y0_S4END[0]
+ Tile_X10Y3_IHP_SRAM/Tile_X0Y0_S4END[10] Tile_X10Y3_IHP_SRAM/Tile_X0Y0_S4END[11]
+ Tile_X10Y3_IHP_SRAM/Tile_X0Y0_S4END[12] Tile_X10Y3_IHP_SRAM/Tile_X0Y0_S4END[13]
+ Tile_X10Y3_IHP_SRAM/Tile_X0Y0_S4END[14] Tile_X10Y3_IHP_SRAM/Tile_X0Y0_S4END[15]
+ Tile_X10Y3_IHP_SRAM/Tile_X0Y0_S4END[1] Tile_X10Y3_IHP_SRAM/Tile_X0Y0_S4END[2] Tile_X10Y3_IHP_SRAM/Tile_X0Y0_S4END[3]
+ Tile_X10Y3_IHP_SRAM/Tile_X0Y0_S4END[4] Tile_X10Y3_IHP_SRAM/Tile_X0Y0_S4END[5] Tile_X10Y3_IHP_SRAM/Tile_X0Y0_S4END[6]
+ Tile_X10Y3_IHP_SRAM/Tile_X0Y0_S4END[7] Tile_X10Y3_IHP_SRAM/Tile_X0Y0_S4END[8] Tile_X10Y3_IHP_SRAM/Tile_X0Y0_S4END[9]
+ Tile_X10Y1_IHP_SRAM/Tile_X0Y1_UserCLK Tile_X9Y2_LUT4AB/W1END[0] Tile_X9Y2_LUT4AB/W1END[1]
+ Tile_X9Y2_LUT4AB/W1END[2] Tile_X9Y2_LUT4AB/W1END[3] Tile_X9Y2_LUT4AB/W2MID[0] Tile_X9Y2_LUT4AB/W2MID[1]
+ Tile_X9Y2_LUT4AB/W2MID[2] Tile_X9Y2_LUT4AB/W2MID[3] Tile_X9Y2_LUT4AB/W2MID[4] Tile_X9Y2_LUT4AB/W2MID[5]
+ Tile_X9Y2_LUT4AB/W2MID[6] Tile_X9Y2_LUT4AB/W2MID[7] Tile_X9Y2_LUT4AB/W2END[0] Tile_X9Y2_LUT4AB/W2END[1]
+ Tile_X9Y2_LUT4AB/W2END[2] Tile_X9Y2_LUT4AB/W2END[3] Tile_X9Y2_LUT4AB/W2END[4] Tile_X9Y2_LUT4AB/W2END[5]
+ Tile_X9Y2_LUT4AB/W2END[6] Tile_X9Y2_LUT4AB/W2END[7] Tile_X9Y2_LUT4AB/W6END[0] Tile_X9Y2_LUT4AB/W6END[10]
+ Tile_X9Y2_LUT4AB/W6END[11] Tile_X9Y2_LUT4AB/W6END[1] Tile_X9Y2_LUT4AB/W6END[2] Tile_X9Y2_LUT4AB/W6END[3]
+ Tile_X9Y2_LUT4AB/W6END[4] Tile_X9Y2_LUT4AB/W6END[5] Tile_X9Y2_LUT4AB/W6END[6] Tile_X9Y2_LUT4AB/W6END[7]
+ Tile_X9Y2_LUT4AB/W6END[8] Tile_X9Y2_LUT4AB/W6END[9] Tile_X9Y2_LUT4AB/WW4END[0] Tile_X9Y2_LUT4AB/WW4END[10]
+ Tile_X9Y2_LUT4AB/WW4END[11] Tile_X9Y2_LUT4AB/WW4END[12] Tile_X9Y2_LUT4AB/WW4END[13]
+ Tile_X9Y2_LUT4AB/WW4END[14] Tile_X9Y2_LUT4AB/WW4END[15] Tile_X9Y2_LUT4AB/WW4END[1]
+ Tile_X9Y2_LUT4AB/WW4END[2] Tile_X9Y2_LUT4AB/WW4END[3] Tile_X9Y2_LUT4AB/WW4END[4]
+ Tile_X9Y2_LUT4AB/WW4END[5] Tile_X9Y2_LUT4AB/WW4END[6] Tile_X9Y2_LUT4AB/WW4END[7]
+ Tile_X9Y2_LUT4AB/WW4END[8] Tile_X9Y2_LUT4AB/WW4END[9] VGND VPWR Tile_X10Y2_WEN_SRAM
+ IHP_SRAM
XTile_X3Y5_LUT4AB Tile_X3Y6_LUT4AB/Co Tile_X3Y5_LUT4AB/Co Tile_X3Y5_LUT4AB/E1BEG[0]
+ Tile_X3Y5_LUT4AB/E1BEG[1] Tile_X3Y5_LUT4AB/E1BEG[2] Tile_X3Y5_LUT4AB/E1BEG[3] Tile_X3Y5_LUT4AB/E1END[0]
+ Tile_X3Y5_LUT4AB/E1END[1] Tile_X3Y5_LUT4AB/E1END[2] Tile_X3Y5_LUT4AB/E1END[3] Tile_X3Y5_LUT4AB/E2BEG[0]
+ Tile_X3Y5_LUT4AB/E2BEG[1] Tile_X3Y5_LUT4AB/E2BEG[2] Tile_X3Y5_LUT4AB/E2BEG[3] Tile_X3Y5_LUT4AB/E2BEG[4]
+ Tile_X3Y5_LUT4AB/E2BEG[5] Tile_X3Y5_LUT4AB/E2BEG[6] Tile_X3Y5_LUT4AB/E2BEG[7] Tile_X4Y5_RegFile/E2END[0]
+ Tile_X4Y5_RegFile/E2END[1] Tile_X4Y5_RegFile/E2END[2] Tile_X4Y5_RegFile/E2END[3]
+ Tile_X4Y5_RegFile/E2END[4] Tile_X4Y5_RegFile/E2END[5] Tile_X4Y5_RegFile/E2END[6]
+ Tile_X4Y5_RegFile/E2END[7] Tile_X3Y5_LUT4AB/E2END[0] Tile_X3Y5_LUT4AB/E2END[1] Tile_X3Y5_LUT4AB/E2END[2]
+ Tile_X3Y5_LUT4AB/E2END[3] Tile_X3Y5_LUT4AB/E2END[4] Tile_X3Y5_LUT4AB/E2END[5] Tile_X3Y5_LUT4AB/E2END[6]
+ Tile_X3Y5_LUT4AB/E2END[7] Tile_X3Y5_LUT4AB/E2MID[0] Tile_X3Y5_LUT4AB/E2MID[1] Tile_X3Y5_LUT4AB/E2MID[2]
+ Tile_X3Y5_LUT4AB/E2MID[3] Tile_X3Y5_LUT4AB/E2MID[4] Tile_X3Y5_LUT4AB/E2MID[5] Tile_X3Y5_LUT4AB/E2MID[6]
+ Tile_X3Y5_LUT4AB/E2MID[7] Tile_X3Y5_LUT4AB/E6BEG[0] Tile_X3Y5_LUT4AB/E6BEG[10] Tile_X3Y5_LUT4AB/E6BEG[11]
+ Tile_X3Y5_LUT4AB/E6BEG[1] Tile_X3Y5_LUT4AB/E6BEG[2] Tile_X3Y5_LUT4AB/E6BEG[3] Tile_X3Y5_LUT4AB/E6BEG[4]
+ Tile_X3Y5_LUT4AB/E6BEG[5] Tile_X3Y5_LUT4AB/E6BEG[6] Tile_X3Y5_LUT4AB/E6BEG[7] Tile_X3Y5_LUT4AB/E6BEG[8]
+ Tile_X3Y5_LUT4AB/E6BEG[9] Tile_X3Y5_LUT4AB/E6END[0] Tile_X3Y5_LUT4AB/E6END[10] Tile_X3Y5_LUT4AB/E6END[11]
+ Tile_X3Y5_LUT4AB/E6END[1] Tile_X3Y5_LUT4AB/E6END[2] Tile_X3Y5_LUT4AB/E6END[3] Tile_X3Y5_LUT4AB/E6END[4]
+ Tile_X3Y5_LUT4AB/E6END[5] Tile_X3Y5_LUT4AB/E6END[6] Tile_X3Y5_LUT4AB/E6END[7] Tile_X3Y5_LUT4AB/E6END[8]
+ Tile_X3Y5_LUT4AB/E6END[9] Tile_X3Y5_LUT4AB/EE4BEG[0] Tile_X3Y5_LUT4AB/EE4BEG[10]
+ Tile_X3Y5_LUT4AB/EE4BEG[11] Tile_X3Y5_LUT4AB/EE4BEG[12] Tile_X3Y5_LUT4AB/EE4BEG[13]
+ Tile_X3Y5_LUT4AB/EE4BEG[14] Tile_X3Y5_LUT4AB/EE4BEG[15] Tile_X3Y5_LUT4AB/EE4BEG[1]
+ Tile_X3Y5_LUT4AB/EE4BEG[2] Tile_X3Y5_LUT4AB/EE4BEG[3] Tile_X3Y5_LUT4AB/EE4BEG[4]
+ Tile_X3Y5_LUT4AB/EE4BEG[5] Tile_X3Y5_LUT4AB/EE4BEG[6] Tile_X3Y5_LUT4AB/EE4BEG[7]
+ Tile_X3Y5_LUT4AB/EE4BEG[8] Tile_X3Y5_LUT4AB/EE4BEG[9] Tile_X3Y5_LUT4AB/EE4END[0]
+ Tile_X3Y5_LUT4AB/EE4END[10] Tile_X3Y5_LUT4AB/EE4END[11] Tile_X3Y5_LUT4AB/EE4END[12]
+ Tile_X3Y5_LUT4AB/EE4END[13] Tile_X3Y5_LUT4AB/EE4END[14] Tile_X3Y5_LUT4AB/EE4END[15]
+ Tile_X3Y5_LUT4AB/EE4END[1] Tile_X3Y5_LUT4AB/EE4END[2] Tile_X3Y5_LUT4AB/EE4END[3]
+ Tile_X3Y5_LUT4AB/EE4END[4] Tile_X3Y5_LUT4AB/EE4END[5] Tile_X3Y5_LUT4AB/EE4END[6]
+ Tile_X3Y5_LUT4AB/EE4END[7] Tile_X3Y5_LUT4AB/EE4END[8] Tile_X3Y5_LUT4AB/EE4END[9]
+ Tile_X3Y5_LUT4AB/FrameData[0] Tile_X3Y5_LUT4AB/FrameData[10] Tile_X3Y5_LUT4AB/FrameData[11]
+ Tile_X3Y5_LUT4AB/FrameData[12] Tile_X3Y5_LUT4AB/FrameData[13] Tile_X3Y5_LUT4AB/FrameData[14]
+ Tile_X3Y5_LUT4AB/FrameData[15] Tile_X3Y5_LUT4AB/FrameData[16] Tile_X3Y5_LUT4AB/FrameData[17]
+ Tile_X3Y5_LUT4AB/FrameData[18] Tile_X3Y5_LUT4AB/FrameData[19] Tile_X3Y5_LUT4AB/FrameData[1]
+ Tile_X3Y5_LUT4AB/FrameData[20] Tile_X3Y5_LUT4AB/FrameData[21] Tile_X3Y5_LUT4AB/FrameData[22]
+ Tile_X3Y5_LUT4AB/FrameData[23] Tile_X3Y5_LUT4AB/FrameData[24] Tile_X3Y5_LUT4AB/FrameData[25]
+ Tile_X3Y5_LUT4AB/FrameData[26] Tile_X3Y5_LUT4AB/FrameData[27] Tile_X3Y5_LUT4AB/FrameData[28]
+ Tile_X3Y5_LUT4AB/FrameData[29] Tile_X3Y5_LUT4AB/FrameData[2] Tile_X3Y5_LUT4AB/FrameData[30]
+ Tile_X3Y5_LUT4AB/FrameData[31] Tile_X3Y5_LUT4AB/FrameData[3] Tile_X3Y5_LUT4AB/FrameData[4]
+ Tile_X3Y5_LUT4AB/FrameData[5] Tile_X3Y5_LUT4AB/FrameData[6] Tile_X3Y5_LUT4AB/FrameData[7]
+ Tile_X3Y5_LUT4AB/FrameData[8] Tile_X3Y5_LUT4AB/FrameData[9] Tile_X4Y5_RegFile/FrameData[0]
+ Tile_X4Y5_RegFile/FrameData[10] Tile_X4Y5_RegFile/FrameData[11] Tile_X4Y5_RegFile/FrameData[12]
+ Tile_X4Y5_RegFile/FrameData[13] Tile_X4Y5_RegFile/FrameData[14] Tile_X4Y5_RegFile/FrameData[15]
+ Tile_X4Y5_RegFile/FrameData[16] Tile_X4Y5_RegFile/FrameData[17] Tile_X4Y5_RegFile/FrameData[18]
+ Tile_X4Y5_RegFile/FrameData[19] Tile_X4Y5_RegFile/FrameData[1] Tile_X4Y5_RegFile/FrameData[20]
+ Tile_X4Y5_RegFile/FrameData[21] Tile_X4Y5_RegFile/FrameData[22] Tile_X4Y5_RegFile/FrameData[23]
+ Tile_X4Y5_RegFile/FrameData[24] Tile_X4Y5_RegFile/FrameData[25] Tile_X4Y5_RegFile/FrameData[26]
+ Tile_X4Y5_RegFile/FrameData[27] Tile_X4Y5_RegFile/FrameData[28] Tile_X4Y5_RegFile/FrameData[29]
+ Tile_X4Y5_RegFile/FrameData[2] Tile_X4Y5_RegFile/FrameData[30] Tile_X4Y5_RegFile/FrameData[31]
+ Tile_X4Y5_RegFile/FrameData[3] Tile_X4Y5_RegFile/FrameData[4] Tile_X4Y5_RegFile/FrameData[5]
+ Tile_X4Y5_RegFile/FrameData[6] Tile_X4Y5_RegFile/FrameData[7] Tile_X4Y5_RegFile/FrameData[8]
+ Tile_X4Y5_RegFile/FrameData[9] Tile_X3Y5_LUT4AB/FrameStrobe[0] Tile_X3Y5_LUT4AB/FrameStrobe[10]
+ Tile_X3Y5_LUT4AB/FrameStrobe[11] Tile_X3Y5_LUT4AB/FrameStrobe[12] Tile_X3Y5_LUT4AB/FrameStrobe[13]
+ Tile_X3Y5_LUT4AB/FrameStrobe[14] Tile_X3Y5_LUT4AB/FrameStrobe[15] Tile_X3Y5_LUT4AB/FrameStrobe[16]
+ Tile_X3Y5_LUT4AB/FrameStrobe[17] Tile_X3Y5_LUT4AB/FrameStrobe[18] Tile_X3Y5_LUT4AB/FrameStrobe[19]
+ Tile_X3Y5_LUT4AB/FrameStrobe[1] Tile_X3Y5_LUT4AB/FrameStrobe[2] Tile_X3Y5_LUT4AB/FrameStrobe[3]
+ Tile_X3Y5_LUT4AB/FrameStrobe[4] Tile_X3Y5_LUT4AB/FrameStrobe[5] Tile_X3Y5_LUT4AB/FrameStrobe[6]
+ Tile_X3Y5_LUT4AB/FrameStrobe[7] Tile_X3Y5_LUT4AB/FrameStrobe[8] Tile_X3Y5_LUT4AB/FrameStrobe[9]
+ Tile_X3Y4_LUT4AB/FrameStrobe[0] Tile_X3Y4_LUT4AB/FrameStrobe[10] Tile_X3Y4_LUT4AB/FrameStrobe[11]
+ Tile_X3Y4_LUT4AB/FrameStrobe[12] Tile_X3Y4_LUT4AB/FrameStrobe[13] Tile_X3Y4_LUT4AB/FrameStrobe[14]
+ Tile_X3Y4_LUT4AB/FrameStrobe[15] Tile_X3Y4_LUT4AB/FrameStrobe[16] Tile_X3Y4_LUT4AB/FrameStrobe[17]
+ Tile_X3Y4_LUT4AB/FrameStrobe[18] Tile_X3Y4_LUT4AB/FrameStrobe[19] Tile_X3Y4_LUT4AB/FrameStrobe[1]
+ Tile_X3Y4_LUT4AB/FrameStrobe[2] Tile_X3Y4_LUT4AB/FrameStrobe[3] Tile_X3Y4_LUT4AB/FrameStrobe[4]
+ Tile_X3Y4_LUT4AB/FrameStrobe[5] Tile_X3Y4_LUT4AB/FrameStrobe[6] Tile_X3Y4_LUT4AB/FrameStrobe[7]
+ Tile_X3Y4_LUT4AB/FrameStrobe[8] Tile_X3Y4_LUT4AB/FrameStrobe[9] Tile_X3Y5_LUT4AB/N1BEG[0]
+ Tile_X3Y5_LUT4AB/N1BEG[1] Tile_X3Y5_LUT4AB/N1BEG[2] Tile_X3Y5_LUT4AB/N1BEG[3] Tile_X3Y6_LUT4AB/N1BEG[0]
+ Tile_X3Y6_LUT4AB/N1BEG[1] Tile_X3Y6_LUT4AB/N1BEG[2] Tile_X3Y6_LUT4AB/N1BEG[3] Tile_X3Y5_LUT4AB/N2BEG[0]
+ Tile_X3Y5_LUT4AB/N2BEG[1] Tile_X3Y5_LUT4AB/N2BEG[2] Tile_X3Y5_LUT4AB/N2BEG[3] Tile_X3Y5_LUT4AB/N2BEG[4]
+ Tile_X3Y5_LUT4AB/N2BEG[5] Tile_X3Y5_LUT4AB/N2BEG[6] Tile_X3Y5_LUT4AB/N2BEG[7] Tile_X3Y4_LUT4AB/N2END[0]
+ Tile_X3Y4_LUT4AB/N2END[1] Tile_X3Y4_LUT4AB/N2END[2] Tile_X3Y4_LUT4AB/N2END[3] Tile_X3Y4_LUT4AB/N2END[4]
+ Tile_X3Y4_LUT4AB/N2END[5] Tile_X3Y4_LUT4AB/N2END[6] Tile_X3Y4_LUT4AB/N2END[7] Tile_X3Y5_LUT4AB/N2END[0]
+ Tile_X3Y5_LUT4AB/N2END[1] Tile_X3Y5_LUT4AB/N2END[2] Tile_X3Y5_LUT4AB/N2END[3] Tile_X3Y5_LUT4AB/N2END[4]
+ Tile_X3Y5_LUT4AB/N2END[5] Tile_X3Y5_LUT4AB/N2END[6] Tile_X3Y5_LUT4AB/N2END[7] Tile_X3Y6_LUT4AB/N2BEG[0]
+ Tile_X3Y6_LUT4AB/N2BEG[1] Tile_X3Y6_LUT4AB/N2BEG[2] Tile_X3Y6_LUT4AB/N2BEG[3] Tile_X3Y6_LUT4AB/N2BEG[4]
+ Tile_X3Y6_LUT4AB/N2BEG[5] Tile_X3Y6_LUT4AB/N2BEG[6] Tile_X3Y6_LUT4AB/N2BEG[7] Tile_X3Y5_LUT4AB/N4BEG[0]
+ Tile_X3Y5_LUT4AB/N4BEG[10] Tile_X3Y5_LUT4AB/N4BEG[11] Tile_X3Y5_LUT4AB/N4BEG[12]
+ Tile_X3Y5_LUT4AB/N4BEG[13] Tile_X3Y5_LUT4AB/N4BEG[14] Tile_X3Y5_LUT4AB/N4BEG[15]
+ Tile_X3Y5_LUT4AB/N4BEG[1] Tile_X3Y5_LUT4AB/N4BEG[2] Tile_X3Y5_LUT4AB/N4BEG[3] Tile_X3Y5_LUT4AB/N4BEG[4]
+ Tile_X3Y5_LUT4AB/N4BEG[5] Tile_X3Y5_LUT4AB/N4BEG[6] Tile_X3Y5_LUT4AB/N4BEG[7] Tile_X3Y5_LUT4AB/N4BEG[8]
+ Tile_X3Y5_LUT4AB/N4BEG[9] Tile_X3Y6_LUT4AB/N4BEG[0] Tile_X3Y6_LUT4AB/N4BEG[10] Tile_X3Y6_LUT4AB/N4BEG[11]
+ Tile_X3Y6_LUT4AB/N4BEG[12] Tile_X3Y6_LUT4AB/N4BEG[13] Tile_X3Y6_LUT4AB/N4BEG[14]
+ Tile_X3Y6_LUT4AB/N4BEG[15] Tile_X3Y6_LUT4AB/N4BEG[1] Tile_X3Y6_LUT4AB/N4BEG[2] Tile_X3Y6_LUT4AB/N4BEG[3]
+ Tile_X3Y6_LUT4AB/N4BEG[4] Tile_X3Y6_LUT4AB/N4BEG[5] Tile_X3Y6_LUT4AB/N4BEG[6] Tile_X3Y6_LUT4AB/N4BEG[7]
+ Tile_X3Y6_LUT4AB/N4BEG[8] Tile_X3Y6_LUT4AB/N4BEG[9] Tile_X3Y5_LUT4AB/NN4BEG[0] Tile_X3Y5_LUT4AB/NN4BEG[10]
+ Tile_X3Y5_LUT4AB/NN4BEG[11] Tile_X3Y5_LUT4AB/NN4BEG[12] Tile_X3Y5_LUT4AB/NN4BEG[13]
+ Tile_X3Y5_LUT4AB/NN4BEG[14] Tile_X3Y5_LUT4AB/NN4BEG[15] Tile_X3Y5_LUT4AB/NN4BEG[1]
+ Tile_X3Y5_LUT4AB/NN4BEG[2] Tile_X3Y5_LUT4AB/NN4BEG[3] Tile_X3Y5_LUT4AB/NN4BEG[4]
+ Tile_X3Y5_LUT4AB/NN4BEG[5] Tile_X3Y5_LUT4AB/NN4BEG[6] Tile_X3Y5_LUT4AB/NN4BEG[7]
+ Tile_X3Y5_LUT4AB/NN4BEG[8] Tile_X3Y5_LUT4AB/NN4BEG[9] Tile_X3Y6_LUT4AB/NN4BEG[0]
+ Tile_X3Y6_LUT4AB/NN4BEG[10] Tile_X3Y6_LUT4AB/NN4BEG[11] Tile_X3Y6_LUT4AB/NN4BEG[12]
+ Tile_X3Y6_LUT4AB/NN4BEG[13] Tile_X3Y6_LUT4AB/NN4BEG[14] Tile_X3Y6_LUT4AB/NN4BEG[15]
+ Tile_X3Y6_LUT4AB/NN4BEG[1] Tile_X3Y6_LUT4AB/NN4BEG[2] Tile_X3Y6_LUT4AB/NN4BEG[3]
+ Tile_X3Y6_LUT4AB/NN4BEG[4] Tile_X3Y6_LUT4AB/NN4BEG[5] Tile_X3Y6_LUT4AB/NN4BEG[6]
+ Tile_X3Y6_LUT4AB/NN4BEG[7] Tile_X3Y6_LUT4AB/NN4BEG[8] Tile_X3Y6_LUT4AB/NN4BEG[9]
+ Tile_X3Y6_LUT4AB/S1END[0] Tile_X3Y6_LUT4AB/S1END[1] Tile_X3Y6_LUT4AB/S1END[2] Tile_X3Y6_LUT4AB/S1END[3]
+ Tile_X3Y5_LUT4AB/S1END[0] Tile_X3Y5_LUT4AB/S1END[1] Tile_X3Y5_LUT4AB/S1END[2] Tile_X3Y5_LUT4AB/S1END[3]
+ Tile_X3Y6_LUT4AB/S2MID[0] Tile_X3Y6_LUT4AB/S2MID[1] Tile_X3Y6_LUT4AB/S2MID[2] Tile_X3Y6_LUT4AB/S2MID[3]
+ Tile_X3Y6_LUT4AB/S2MID[4] Tile_X3Y6_LUT4AB/S2MID[5] Tile_X3Y6_LUT4AB/S2MID[6] Tile_X3Y6_LUT4AB/S2MID[7]
+ Tile_X3Y6_LUT4AB/S2END[0] Tile_X3Y6_LUT4AB/S2END[1] Tile_X3Y6_LUT4AB/S2END[2] Tile_X3Y6_LUT4AB/S2END[3]
+ Tile_X3Y6_LUT4AB/S2END[4] Tile_X3Y6_LUT4AB/S2END[5] Tile_X3Y6_LUT4AB/S2END[6] Tile_X3Y6_LUT4AB/S2END[7]
+ Tile_X3Y5_LUT4AB/S2END[0] Tile_X3Y5_LUT4AB/S2END[1] Tile_X3Y5_LUT4AB/S2END[2] Tile_X3Y5_LUT4AB/S2END[3]
+ Tile_X3Y5_LUT4AB/S2END[4] Tile_X3Y5_LUT4AB/S2END[5] Tile_X3Y5_LUT4AB/S2END[6] Tile_X3Y5_LUT4AB/S2END[7]
+ Tile_X3Y5_LUT4AB/S2MID[0] Tile_X3Y5_LUT4AB/S2MID[1] Tile_X3Y5_LUT4AB/S2MID[2] Tile_X3Y5_LUT4AB/S2MID[3]
+ Tile_X3Y5_LUT4AB/S2MID[4] Tile_X3Y5_LUT4AB/S2MID[5] Tile_X3Y5_LUT4AB/S2MID[6] Tile_X3Y5_LUT4AB/S2MID[7]
+ Tile_X3Y6_LUT4AB/S4END[0] Tile_X3Y6_LUT4AB/S4END[10] Tile_X3Y6_LUT4AB/S4END[11]
+ Tile_X3Y6_LUT4AB/S4END[12] Tile_X3Y6_LUT4AB/S4END[13] Tile_X3Y6_LUT4AB/S4END[14]
+ Tile_X3Y6_LUT4AB/S4END[15] Tile_X3Y6_LUT4AB/S4END[1] Tile_X3Y6_LUT4AB/S4END[2] Tile_X3Y6_LUT4AB/S4END[3]
+ Tile_X3Y6_LUT4AB/S4END[4] Tile_X3Y6_LUT4AB/S4END[5] Tile_X3Y6_LUT4AB/S4END[6] Tile_X3Y6_LUT4AB/S4END[7]
+ Tile_X3Y6_LUT4AB/S4END[8] Tile_X3Y6_LUT4AB/S4END[9] Tile_X3Y5_LUT4AB/S4END[0] Tile_X3Y5_LUT4AB/S4END[10]
+ Tile_X3Y5_LUT4AB/S4END[11] Tile_X3Y5_LUT4AB/S4END[12] Tile_X3Y5_LUT4AB/S4END[13]
+ Tile_X3Y5_LUT4AB/S4END[14] Tile_X3Y5_LUT4AB/S4END[15] Tile_X3Y5_LUT4AB/S4END[1]
+ Tile_X3Y5_LUT4AB/S4END[2] Tile_X3Y5_LUT4AB/S4END[3] Tile_X3Y5_LUT4AB/S4END[4] Tile_X3Y5_LUT4AB/S4END[5]
+ Tile_X3Y5_LUT4AB/S4END[6] Tile_X3Y5_LUT4AB/S4END[7] Tile_X3Y5_LUT4AB/S4END[8] Tile_X3Y5_LUT4AB/S4END[9]
+ Tile_X3Y6_LUT4AB/SS4END[0] Tile_X3Y6_LUT4AB/SS4END[10] Tile_X3Y6_LUT4AB/SS4END[11]
+ Tile_X3Y6_LUT4AB/SS4END[12] Tile_X3Y6_LUT4AB/SS4END[13] Tile_X3Y6_LUT4AB/SS4END[14]
+ Tile_X3Y6_LUT4AB/SS4END[15] Tile_X3Y6_LUT4AB/SS4END[1] Tile_X3Y6_LUT4AB/SS4END[2]
+ Tile_X3Y6_LUT4AB/SS4END[3] Tile_X3Y6_LUT4AB/SS4END[4] Tile_X3Y6_LUT4AB/SS4END[5]
+ Tile_X3Y6_LUT4AB/SS4END[6] Tile_X3Y6_LUT4AB/SS4END[7] Tile_X3Y6_LUT4AB/SS4END[8]
+ Tile_X3Y6_LUT4AB/SS4END[9] Tile_X3Y5_LUT4AB/SS4END[0] Tile_X3Y5_LUT4AB/SS4END[10]
+ Tile_X3Y5_LUT4AB/SS4END[11] Tile_X3Y5_LUT4AB/SS4END[12] Tile_X3Y5_LUT4AB/SS4END[13]
+ Tile_X3Y5_LUT4AB/SS4END[14] Tile_X3Y5_LUT4AB/SS4END[15] Tile_X3Y5_LUT4AB/SS4END[1]
+ Tile_X3Y5_LUT4AB/SS4END[2] Tile_X3Y5_LUT4AB/SS4END[3] Tile_X3Y5_LUT4AB/SS4END[4]
+ Tile_X3Y5_LUT4AB/SS4END[5] Tile_X3Y5_LUT4AB/SS4END[6] Tile_X3Y5_LUT4AB/SS4END[7]
+ Tile_X3Y5_LUT4AB/SS4END[8] Tile_X3Y5_LUT4AB/SS4END[9] Tile_X3Y5_LUT4AB/UserCLK Tile_X3Y4_LUT4AB/UserCLK
+ VGND VPWR Tile_X3Y5_LUT4AB/W1BEG[0] Tile_X3Y5_LUT4AB/W1BEG[1] Tile_X3Y5_LUT4AB/W1BEG[2]
+ Tile_X3Y5_LUT4AB/W1BEG[3] Tile_X3Y5_LUT4AB/W1END[0] Tile_X3Y5_LUT4AB/W1END[1] Tile_X3Y5_LUT4AB/W1END[2]
+ Tile_X3Y5_LUT4AB/W1END[3] Tile_X3Y5_LUT4AB/W2BEG[0] Tile_X3Y5_LUT4AB/W2BEG[1] Tile_X3Y5_LUT4AB/W2BEG[2]
+ Tile_X3Y5_LUT4AB/W2BEG[3] Tile_X3Y5_LUT4AB/W2BEG[4] Tile_X3Y5_LUT4AB/W2BEG[5] Tile_X3Y5_LUT4AB/W2BEG[6]
+ Tile_X3Y5_LUT4AB/W2BEG[7] Tile_X2Y5_LUT4AB/W2END[0] Tile_X2Y5_LUT4AB/W2END[1] Tile_X2Y5_LUT4AB/W2END[2]
+ Tile_X2Y5_LUT4AB/W2END[3] Tile_X2Y5_LUT4AB/W2END[4] Tile_X2Y5_LUT4AB/W2END[5] Tile_X2Y5_LUT4AB/W2END[6]
+ Tile_X2Y5_LUT4AB/W2END[7] Tile_X3Y5_LUT4AB/W2END[0] Tile_X3Y5_LUT4AB/W2END[1] Tile_X3Y5_LUT4AB/W2END[2]
+ Tile_X3Y5_LUT4AB/W2END[3] Tile_X3Y5_LUT4AB/W2END[4] Tile_X3Y5_LUT4AB/W2END[5] Tile_X3Y5_LUT4AB/W2END[6]
+ Tile_X3Y5_LUT4AB/W2END[7] Tile_X3Y5_LUT4AB/W2MID[0] Tile_X3Y5_LUT4AB/W2MID[1] Tile_X3Y5_LUT4AB/W2MID[2]
+ Tile_X3Y5_LUT4AB/W2MID[3] Tile_X3Y5_LUT4AB/W2MID[4] Tile_X3Y5_LUT4AB/W2MID[5] Tile_X3Y5_LUT4AB/W2MID[6]
+ Tile_X3Y5_LUT4AB/W2MID[7] Tile_X3Y5_LUT4AB/W6BEG[0] Tile_X3Y5_LUT4AB/W6BEG[10] Tile_X3Y5_LUT4AB/W6BEG[11]
+ Tile_X3Y5_LUT4AB/W6BEG[1] Tile_X3Y5_LUT4AB/W6BEG[2] Tile_X3Y5_LUT4AB/W6BEG[3] Tile_X3Y5_LUT4AB/W6BEG[4]
+ Tile_X3Y5_LUT4AB/W6BEG[5] Tile_X3Y5_LUT4AB/W6BEG[6] Tile_X3Y5_LUT4AB/W6BEG[7] Tile_X3Y5_LUT4AB/W6BEG[8]
+ Tile_X3Y5_LUT4AB/W6BEG[9] Tile_X3Y5_LUT4AB/W6END[0] Tile_X3Y5_LUT4AB/W6END[10] Tile_X3Y5_LUT4AB/W6END[11]
+ Tile_X3Y5_LUT4AB/W6END[1] Tile_X3Y5_LUT4AB/W6END[2] Tile_X3Y5_LUT4AB/W6END[3] Tile_X3Y5_LUT4AB/W6END[4]
+ Tile_X3Y5_LUT4AB/W6END[5] Tile_X3Y5_LUT4AB/W6END[6] Tile_X3Y5_LUT4AB/W6END[7] Tile_X3Y5_LUT4AB/W6END[8]
+ Tile_X3Y5_LUT4AB/W6END[9] Tile_X3Y5_LUT4AB/WW4BEG[0] Tile_X3Y5_LUT4AB/WW4BEG[10]
+ Tile_X3Y5_LUT4AB/WW4BEG[11] Tile_X3Y5_LUT4AB/WW4BEG[12] Tile_X3Y5_LUT4AB/WW4BEG[13]
+ Tile_X3Y5_LUT4AB/WW4BEG[14] Tile_X3Y5_LUT4AB/WW4BEG[15] Tile_X3Y5_LUT4AB/WW4BEG[1]
+ Tile_X3Y5_LUT4AB/WW4BEG[2] Tile_X3Y5_LUT4AB/WW4BEG[3] Tile_X3Y5_LUT4AB/WW4BEG[4]
+ Tile_X3Y5_LUT4AB/WW4BEG[5] Tile_X3Y5_LUT4AB/WW4BEG[6] Tile_X3Y5_LUT4AB/WW4BEG[7]
+ Tile_X3Y5_LUT4AB/WW4BEG[8] Tile_X3Y5_LUT4AB/WW4BEG[9] Tile_X3Y5_LUT4AB/WW4END[0]
+ Tile_X3Y5_LUT4AB/WW4END[10] Tile_X3Y5_LUT4AB/WW4END[11] Tile_X3Y5_LUT4AB/WW4END[12]
+ Tile_X3Y5_LUT4AB/WW4END[13] Tile_X3Y5_LUT4AB/WW4END[14] Tile_X3Y5_LUT4AB/WW4END[15]
+ Tile_X3Y5_LUT4AB/WW4END[1] Tile_X3Y5_LUT4AB/WW4END[2] Tile_X3Y5_LUT4AB/WW4END[3]
+ Tile_X3Y5_LUT4AB/WW4END[4] Tile_X3Y5_LUT4AB/WW4END[5] Tile_X3Y5_LUT4AB/WW4END[6]
+ Tile_X3Y5_LUT4AB/WW4END[7] Tile_X3Y5_LUT4AB/WW4END[8] Tile_X3Y5_LUT4AB/WW4END[9]
+ LUT4AB
XTile_X2Y9_LUT4AB Tile_X2Y9_LUT4AB/Ci Tile_X2Y9_LUT4AB/Co Tile_X3Y9_LUT4AB/E1END[0]
+ Tile_X3Y9_LUT4AB/E1END[1] Tile_X3Y9_LUT4AB/E1END[2] Tile_X3Y9_LUT4AB/E1END[3] Tile_X2Y9_LUT4AB/E1END[0]
+ Tile_X2Y9_LUT4AB/E1END[1] Tile_X2Y9_LUT4AB/E1END[2] Tile_X2Y9_LUT4AB/E1END[3] Tile_X3Y9_LUT4AB/E2MID[0]
+ Tile_X3Y9_LUT4AB/E2MID[1] Tile_X3Y9_LUT4AB/E2MID[2] Tile_X3Y9_LUT4AB/E2MID[3] Tile_X3Y9_LUT4AB/E2MID[4]
+ Tile_X3Y9_LUT4AB/E2MID[5] Tile_X3Y9_LUT4AB/E2MID[6] Tile_X3Y9_LUT4AB/E2MID[7] Tile_X3Y9_LUT4AB/E2END[0]
+ Tile_X3Y9_LUT4AB/E2END[1] Tile_X3Y9_LUT4AB/E2END[2] Tile_X3Y9_LUT4AB/E2END[3] Tile_X3Y9_LUT4AB/E2END[4]
+ Tile_X3Y9_LUT4AB/E2END[5] Tile_X3Y9_LUT4AB/E2END[6] Tile_X3Y9_LUT4AB/E2END[7] Tile_X2Y9_LUT4AB/E2END[0]
+ Tile_X2Y9_LUT4AB/E2END[1] Tile_X2Y9_LUT4AB/E2END[2] Tile_X2Y9_LUT4AB/E2END[3] Tile_X2Y9_LUT4AB/E2END[4]
+ Tile_X2Y9_LUT4AB/E2END[5] Tile_X2Y9_LUT4AB/E2END[6] Tile_X2Y9_LUT4AB/E2END[7] Tile_X2Y9_LUT4AB/E2MID[0]
+ Tile_X2Y9_LUT4AB/E2MID[1] Tile_X2Y9_LUT4AB/E2MID[2] Tile_X2Y9_LUT4AB/E2MID[3] Tile_X2Y9_LUT4AB/E2MID[4]
+ Tile_X2Y9_LUT4AB/E2MID[5] Tile_X2Y9_LUT4AB/E2MID[6] Tile_X2Y9_LUT4AB/E2MID[7] Tile_X3Y9_LUT4AB/E6END[0]
+ Tile_X3Y9_LUT4AB/E6END[10] Tile_X3Y9_LUT4AB/E6END[11] Tile_X3Y9_LUT4AB/E6END[1]
+ Tile_X3Y9_LUT4AB/E6END[2] Tile_X3Y9_LUT4AB/E6END[3] Tile_X3Y9_LUT4AB/E6END[4] Tile_X3Y9_LUT4AB/E6END[5]
+ Tile_X3Y9_LUT4AB/E6END[6] Tile_X3Y9_LUT4AB/E6END[7] Tile_X3Y9_LUT4AB/E6END[8] Tile_X3Y9_LUT4AB/E6END[9]
+ Tile_X2Y9_LUT4AB/E6END[0] Tile_X2Y9_LUT4AB/E6END[10] Tile_X2Y9_LUT4AB/E6END[11]
+ Tile_X2Y9_LUT4AB/E6END[1] Tile_X2Y9_LUT4AB/E6END[2] Tile_X2Y9_LUT4AB/E6END[3] Tile_X2Y9_LUT4AB/E6END[4]
+ Tile_X2Y9_LUT4AB/E6END[5] Tile_X2Y9_LUT4AB/E6END[6] Tile_X2Y9_LUT4AB/E6END[7] Tile_X2Y9_LUT4AB/E6END[8]
+ Tile_X2Y9_LUT4AB/E6END[9] Tile_X3Y9_LUT4AB/EE4END[0] Tile_X3Y9_LUT4AB/EE4END[10]
+ Tile_X3Y9_LUT4AB/EE4END[11] Tile_X3Y9_LUT4AB/EE4END[12] Tile_X3Y9_LUT4AB/EE4END[13]
+ Tile_X3Y9_LUT4AB/EE4END[14] Tile_X3Y9_LUT4AB/EE4END[15] Tile_X3Y9_LUT4AB/EE4END[1]
+ Tile_X3Y9_LUT4AB/EE4END[2] Tile_X3Y9_LUT4AB/EE4END[3] Tile_X3Y9_LUT4AB/EE4END[4]
+ Tile_X3Y9_LUT4AB/EE4END[5] Tile_X3Y9_LUT4AB/EE4END[6] Tile_X3Y9_LUT4AB/EE4END[7]
+ Tile_X3Y9_LUT4AB/EE4END[8] Tile_X3Y9_LUT4AB/EE4END[9] Tile_X2Y9_LUT4AB/EE4END[0]
+ Tile_X2Y9_LUT4AB/EE4END[10] Tile_X2Y9_LUT4AB/EE4END[11] Tile_X2Y9_LUT4AB/EE4END[12]
+ Tile_X2Y9_LUT4AB/EE4END[13] Tile_X2Y9_LUT4AB/EE4END[14] Tile_X2Y9_LUT4AB/EE4END[15]
+ Tile_X2Y9_LUT4AB/EE4END[1] Tile_X2Y9_LUT4AB/EE4END[2] Tile_X2Y9_LUT4AB/EE4END[3]
+ Tile_X2Y9_LUT4AB/EE4END[4] Tile_X2Y9_LUT4AB/EE4END[5] Tile_X2Y9_LUT4AB/EE4END[6]
+ Tile_X2Y9_LUT4AB/EE4END[7] Tile_X2Y9_LUT4AB/EE4END[8] Tile_X2Y9_LUT4AB/EE4END[9]
+ Tile_X2Y9_LUT4AB/FrameData[0] Tile_X2Y9_LUT4AB/FrameData[10] Tile_X2Y9_LUT4AB/FrameData[11]
+ Tile_X2Y9_LUT4AB/FrameData[12] Tile_X2Y9_LUT4AB/FrameData[13] Tile_X2Y9_LUT4AB/FrameData[14]
+ Tile_X2Y9_LUT4AB/FrameData[15] Tile_X2Y9_LUT4AB/FrameData[16] Tile_X2Y9_LUT4AB/FrameData[17]
+ Tile_X2Y9_LUT4AB/FrameData[18] Tile_X2Y9_LUT4AB/FrameData[19] Tile_X2Y9_LUT4AB/FrameData[1]
+ Tile_X2Y9_LUT4AB/FrameData[20] Tile_X2Y9_LUT4AB/FrameData[21] Tile_X2Y9_LUT4AB/FrameData[22]
+ Tile_X2Y9_LUT4AB/FrameData[23] Tile_X2Y9_LUT4AB/FrameData[24] Tile_X2Y9_LUT4AB/FrameData[25]
+ Tile_X2Y9_LUT4AB/FrameData[26] Tile_X2Y9_LUT4AB/FrameData[27] Tile_X2Y9_LUT4AB/FrameData[28]
+ Tile_X2Y9_LUT4AB/FrameData[29] Tile_X2Y9_LUT4AB/FrameData[2] Tile_X2Y9_LUT4AB/FrameData[30]
+ Tile_X2Y9_LUT4AB/FrameData[31] Tile_X2Y9_LUT4AB/FrameData[3] Tile_X2Y9_LUT4AB/FrameData[4]
+ Tile_X2Y9_LUT4AB/FrameData[5] Tile_X2Y9_LUT4AB/FrameData[6] Tile_X2Y9_LUT4AB/FrameData[7]
+ Tile_X2Y9_LUT4AB/FrameData[8] Tile_X2Y9_LUT4AB/FrameData[9] Tile_X3Y9_LUT4AB/FrameData[0]
+ Tile_X3Y9_LUT4AB/FrameData[10] Tile_X3Y9_LUT4AB/FrameData[11] Tile_X3Y9_LUT4AB/FrameData[12]
+ Tile_X3Y9_LUT4AB/FrameData[13] Tile_X3Y9_LUT4AB/FrameData[14] Tile_X3Y9_LUT4AB/FrameData[15]
+ Tile_X3Y9_LUT4AB/FrameData[16] Tile_X3Y9_LUT4AB/FrameData[17] Tile_X3Y9_LUT4AB/FrameData[18]
+ Tile_X3Y9_LUT4AB/FrameData[19] Tile_X3Y9_LUT4AB/FrameData[1] Tile_X3Y9_LUT4AB/FrameData[20]
+ Tile_X3Y9_LUT4AB/FrameData[21] Tile_X3Y9_LUT4AB/FrameData[22] Tile_X3Y9_LUT4AB/FrameData[23]
+ Tile_X3Y9_LUT4AB/FrameData[24] Tile_X3Y9_LUT4AB/FrameData[25] Tile_X3Y9_LUT4AB/FrameData[26]
+ Tile_X3Y9_LUT4AB/FrameData[27] Tile_X3Y9_LUT4AB/FrameData[28] Tile_X3Y9_LUT4AB/FrameData[29]
+ Tile_X3Y9_LUT4AB/FrameData[2] Tile_X3Y9_LUT4AB/FrameData[30] Tile_X3Y9_LUT4AB/FrameData[31]
+ Tile_X3Y9_LUT4AB/FrameData[3] Tile_X3Y9_LUT4AB/FrameData[4] Tile_X3Y9_LUT4AB/FrameData[5]
+ Tile_X3Y9_LUT4AB/FrameData[6] Tile_X3Y9_LUT4AB/FrameData[7] Tile_X3Y9_LUT4AB/FrameData[8]
+ Tile_X3Y9_LUT4AB/FrameData[9] Tile_X2Y9_LUT4AB/FrameStrobe[0] Tile_X2Y9_LUT4AB/FrameStrobe[10]
+ Tile_X2Y9_LUT4AB/FrameStrobe[11] Tile_X2Y9_LUT4AB/FrameStrobe[12] Tile_X2Y9_LUT4AB/FrameStrobe[13]
+ Tile_X2Y9_LUT4AB/FrameStrobe[14] Tile_X2Y9_LUT4AB/FrameStrobe[15] Tile_X2Y9_LUT4AB/FrameStrobe[16]
+ Tile_X2Y9_LUT4AB/FrameStrobe[17] Tile_X2Y9_LUT4AB/FrameStrobe[18] Tile_X2Y9_LUT4AB/FrameStrobe[19]
+ Tile_X2Y9_LUT4AB/FrameStrobe[1] Tile_X2Y9_LUT4AB/FrameStrobe[2] Tile_X2Y9_LUT4AB/FrameStrobe[3]
+ Tile_X2Y9_LUT4AB/FrameStrobe[4] Tile_X2Y9_LUT4AB/FrameStrobe[5] Tile_X2Y9_LUT4AB/FrameStrobe[6]
+ Tile_X2Y9_LUT4AB/FrameStrobe[7] Tile_X2Y9_LUT4AB/FrameStrobe[8] Tile_X2Y9_LUT4AB/FrameStrobe[9]
+ Tile_X2Y8_LUT4AB/FrameStrobe[0] Tile_X2Y8_LUT4AB/FrameStrobe[10] Tile_X2Y8_LUT4AB/FrameStrobe[11]
+ Tile_X2Y8_LUT4AB/FrameStrobe[12] Tile_X2Y8_LUT4AB/FrameStrobe[13] Tile_X2Y8_LUT4AB/FrameStrobe[14]
+ Tile_X2Y8_LUT4AB/FrameStrobe[15] Tile_X2Y8_LUT4AB/FrameStrobe[16] Tile_X2Y8_LUT4AB/FrameStrobe[17]
+ Tile_X2Y8_LUT4AB/FrameStrobe[18] Tile_X2Y8_LUT4AB/FrameStrobe[19] Tile_X2Y8_LUT4AB/FrameStrobe[1]
+ Tile_X2Y8_LUT4AB/FrameStrobe[2] Tile_X2Y8_LUT4AB/FrameStrobe[3] Tile_X2Y8_LUT4AB/FrameStrobe[4]
+ Tile_X2Y8_LUT4AB/FrameStrobe[5] Tile_X2Y8_LUT4AB/FrameStrobe[6] Tile_X2Y8_LUT4AB/FrameStrobe[7]
+ Tile_X2Y8_LUT4AB/FrameStrobe[8] Tile_X2Y8_LUT4AB/FrameStrobe[9] Tile_X2Y9_LUT4AB/N1BEG[0]
+ Tile_X2Y9_LUT4AB/N1BEG[1] Tile_X2Y9_LUT4AB/N1BEG[2] Tile_X2Y9_LUT4AB/N1BEG[3] Tile_X2Y9_LUT4AB/N1END[0]
+ Tile_X2Y9_LUT4AB/N1END[1] Tile_X2Y9_LUT4AB/N1END[2] Tile_X2Y9_LUT4AB/N1END[3] Tile_X2Y9_LUT4AB/N2BEG[0]
+ Tile_X2Y9_LUT4AB/N2BEG[1] Tile_X2Y9_LUT4AB/N2BEG[2] Tile_X2Y9_LUT4AB/N2BEG[3] Tile_X2Y9_LUT4AB/N2BEG[4]
+ Tile_X2Y9_LUT4AB/N2BEG[5] Tile_X2Y9_LUT4AB/N2BEG[6] Tile_X2Y9_LUT4AB/N2BEG[7] Tile_X2Y8_LUT4AB/N2END[0]
+ Tile_X2Y8_LUT4AB/N2END[1] Tile_X2Y8_LUT4AB/N2END[2] Tile_X2Y8_LUT4AB/N2END[3] Tile_X2Y8_LUT4AB/N2END[4]
+ Tile_X2Y8_LUT4AB/N2END[5] Tile_X2Y8_LUT4AB/N2END[6] Tile_X2Y8_LUT4AB/N2END[7] Tile_X2Y9_LUT4AB/N2END[0]
+ Tile_X2Y9_LUT4AB/N2END[1] Tile_X2Y9_LUT4AB/N2END[2] Tile_X2Y9_LUT4AB/N2END[3] Tile_X2Y9_LUT4AB/N2END[4]
+ Tile_X2Y9_LUT4AB/N2END[5] Tile_X2Y9_LUT4AB/N2END[6] Tile_X2Y9_LUT4AB/N2END[7] Tile_X2Y9_LUT4AB/N2MID[0]
+ Tile_X2Y9_LUT4AB/N2MID[1] Tile_X2Y9_LUT4AB/N2MID[2] Tile_X2Y9_LUT4AB/N2MID[3] Tile_X2Y9_LUT4AB/N2MID[4]
+ Tile_X2Y9_LUT4AB/N2MID[5] Tile_X2Y9_LUT4AB/N2MID[6] Tile_X2Y9_LUT4AB/N2MID[7] Tile_X2Y9_LUT4AB/N4BEG[0]
+ Tile_X2Y9_LUT4AB/N4BEG[10] Tile_X2Y9_LUT4AB/N4BEG[11] Tile_X2Y9_LUT4AB/N4BEG[12]
+ Tile_X2Y9_LUT4AB/N4BEG[13] Tile_X2Y9_LUT4AB/N4BEG[14] Tile_X2Y9_LUT4AB/N4BEG[15]
+ Tile_X2Y9_LUT4AB/N4BEG[1] Tile_X2Y9_LUT4AB/N4BEG[2] Tile_X2Y9_LUT4AB/N4BEG[3] Tile_X2Y9_LUT4AB/N4BEG[4]
+ Tile_X2Y9_LUT4AB/N4BEG[5] Tile_X2Y9_LUT4AB/N4BEG[6] Tile_X2Y9_LUT4AB/N4BEG[7] Tile_X2Y9_LUT4AB/N4BEG[8]
+ Tile_X2Y9_LUT4AB/N4BEG[9] Tile_X2Y9_LUT4AB/N4END[0] Tile_X2Y9_LUT4AB/N4END[10] Tile_X2Y9_LUT4AB/N4END[11]
+ Tile_X2Y9_LUT4AB/N4END[12] Tile_X2Y9_LUT4AB/N4END[13] Tile_X2Y9_LUT4AB/N4END[14]
+ Tile_X2Y9_LUT4AB/N4END[15] Tile_X2Y9_LUT4AB/N4END[1] Tile_X2Y9_LUT4AB/N4END[2] Tile_X2Y9_LUT4AB/N4END[3]
+ Tile_X2Y9_LUT4AB/N4END[4] Tile_X2Y9_LUT4AB/N4END[5] Tile_X2Y9_LUT4AB/N4END[6] Tile_X2Y9_LUT4AB/N4END[7]
+ Tile_X2Y9_LUT4AB/N4END[8] Tile_X2Y9_LUT4AB/N4END[9] Tile_X2Y9_LUT4AB/NN4BEG[0] Tile_X2Y9_LUT4AB/NN4BEG[10]
+ Tile_X2Y9_LUT4AB/NN4BEG[11] Tile_X2Y9_LUT4AB/NN4BEG[12] Tile_X2Y9_LUT4AB/NN4BEG[13]
+ Tile_X2Y9_LUT4AB/NN4BEG[14] Tile_X2Y9_LUT4AB/NN4BEG[15] Tile_X2Y9_LUT4AB/NN4BEG[1]
+ Tile_X2Y9_LUT4AB/NN4BEG[2] Tile_X2Y9_LUT4AB/NN4BEG[3] Tile_X2Y9_LUT4AB/NN4BEG[4]
+ Tile_X2Y9_LUT4AB/NN4BEG[5] Tile_X2Y9_LUT4AB/NN4BEG[6] Tile_X2Y9_LUT4AB/NN4BEG[7]
+ Tile_X2Y9_LUT4AB/NN4BEG[8] Tile_X2Y9_LUT4AB/NN4BEG[9] Tile_X2Y9_LUT4AB/NN4END[0]
+ Tile_X2Y9_LUT4AB/NN4END[10] Tile_X2Y9_LUT4AB/NN4END[11] Tile_X2Y9_LUT4AB/NN4END[12]
+ Tile_X2Y9_LUT4AB/NN4END[13] Tile_X2Y9_LUT4AB/NN4END[14] Tile_X2Y9_LUT4AB/NN4END[15]
+ Tile_X2Y9_LUT4AB/NN4END[1] Tile_X2Y9_LUT4AB/NN4END[2] Tile_X2Y9_LUT4AB/NN4END[3]
+ Tile_X2Y9_LUT4AB/NN4END[4] Tile_X2Y9_LUT4AB/NN4END[5] Tile_X2Y9_LUT4AB/NN4END[6]
+ Tile_X2Y9_LUT4AB/NN4END[7] Tile_X2Y9_LUT4AB/NN4END[8] Tile_X2Y9_LUT4AB/NN4END[9]
+ Tile_X2Y9_LUT4AB/S1BEG[0] Tile_X2Y9_LUT4AB/S1BEG[1] Tile_X2Y9_LUT4AB/S1BEG[2] Tile_X2Y9_LUT4AB/S1BEG[3]
+ Tile_X2Y9_LUT4AB/S1END[0] Tile_X2Y9_LUT4AB/S1END[1] Tile_X2Y9_LUT4AB/S1END[2] Tile_X2Y9_LUT4AB/S1END[3]
+ Tile_X2Y9_LUT4AB/S2BEG[0] Tile_X2Y9_LUT4AB/S2BEG[1] Tile_X2Y9_LUT4AB/S2BEG[2] Tile_X2Y9_LUT4AB/S2BEG[3]
+ Tile_X2Y9_LUT4AB/S2BEG[4] Tile_X2Y9_LUT4AB/S2BEG[5] Tile_X2Y9_LUT4AB/S2BEG[6] Tile_X2Y9_LUT4AB/S2BEG[7]
+ Tile_X2Y9_LUT4AB/S2BEGb[0] Tile_X2Y9_LUT4AB/S2BEGb[1] Tile_X2Y9_LUT4AB/S2BEGb[2]
+ Tile_X2Y9_LUT4AB/S2BEGb[3] Tile_X2Y9_LUT4AB/S2BEGb[4] Tile_X2Y9_LUT4AB/S2BEGb[5]
+ Tile_X2Y9_LUT4AB/S2BEGb[6] Tile_X2Y9_LUT4AB/S2BEGb[7] Tile_X2Y9_LUT4AB/S2END[0]
+ Tile_X2Y9_LUT4AB/S2END[1] Tile_X2Y9_LUT4AB/S2END[2] Tile_X2Y9_LUT4AB/S2END[3] Tile_X2Y9_LUT4AB/S2END[4]
+ Tile_X2Y9_LUT4AB/S2END[5] Tile_X2Y9_LUT4AB/S2END[6] Tile_X2Y9_LUT4AB/S2END[7] Tile_X2Y9_LUT4AB/S2MID[0]
+ Tile_X2Y9_LUT4AB/S2MID[1] Tile_X2Y9_LUT4AB/S2MID[2] Tile_X2Y9_LUT4AB/S2MID[3] Tile_X2Y9_LUT4AB/S2MID[4]
+ Tile_X2Y9_LUT4AB/S2MID[5] Tile_X2Y9_LUT4AB/S2MID[6] Tile_X2Y9_LUT4AB/S2MID[7] Tile_X2Y9_LUT4AB/S4BEG[0]
+ Tile_X2Y9_LUT4AB/S4BEG[10] Tile_X2Y9_LUT4AB/S4BEG[11] Tile_X2Y9_LUT4AB/S4BEG[12]
+ Tile_X2Y9_LUT4AB/S4BEG[13] Tile_X2Y9_LUT4AB/S4BEG[14] Tile_X2Y9_LUT4AB/S4BEG[15]
+ Tile_X2Y9_LUT4AB/S4BEG[1] Tile_X2Y9_LUT4AB/S4BEG[2] Tile_X2Y9_LUT4AB/S4BEG[3] Tile_X2Y9_LUT4AB/S4BEG[4]
+ Tile_X2Y9_LUT4AB/S4BEG[5] Tile_X2Y9_LUT4AB/S4BEG[6] Tile_X2Y9_LUT4AB/S4BEG[7] Tile_X2Y9_LUT4AB/S4BEG[8]
+ Tile_X2Y9_LUT4AB/S4BEG[9] Tile_X2Y9_LUT4AB/S4END[0] Tile_X2Y9_LUT4AB/S4END[10] Tile_X2Y9_LUT4AB/S4END[11]
+ Tile_X2Y9_LUT4AB/S4END[12] Tile_X2Y9_LUT4AB/S4END[13] Tile_X2Y9_LUT4AB/S4END[14]
+ Tile_X2Y9_LUT4AB/S4END[15] Tile_X2Y9_LUT4AB/S4END[1] Tile_X2Y9_LUT4AB/S4END[2] Tile_X2Y9_LUT4AB/S4END[3]
+ Tile_X2Y9_LUT4AB/S4END[4] Tile_X2Y9_LUT4AB/S4END[5] Tile_X2Y9_LUT4AB/S4END[6] Tile_X2Y9_LUT4AB/S4END[7]
+ Tile_X2Y9_LUT4AB/S4END[8] Tile_X2Y9_LUT4AB/S4END[9] Tile_X2Y9_LUT4AB/SS4BEG[0] Tile_X2Y9_LUT4AB/SS4BEG[10]
+ Tile_X2Y9_LUT4AB/SS4BEG[11] Tile_X2Y9_LUT4AB/SS4BEG[12] Tile_X2Y9_LUT4AB/SS4BEG[13]
+ Tile_X2Y9_LUT4AB/SS4BEG[14] Tile_X2Y9_LUT4AB/SS4BEG[15] Tile_X2Y9_LUT4AB/SS4BEG[1]
+ Tile_X2Y9_LUT4AB/SS4BEG[2] Tile_X2Y9_LUT4AB/SS4BEG[3] Tile_X2Y9_LUT4AB/SS4BEG[4]
+ Tile_X2Y9_LUT4AB/SS4BEG[5] Tile_X2Y9_LUT4AB/SS4BEG[6] Tile_X2Y9_LUT4AB/SS4BEG[7]
+ Tile_X2Y9_LUT4AB/SS4BEG[8] Tile_X2Y9_LUT4AB/SS4BEG[9] Tile_X2Y9_LUT4AB/SS4END[0]
+ Tile_X2Y9_LUT4AB/SS4END[10] Tile_X2Y9_LUT4AB/SS4END[11] Tile_X2Y9_LUT4AB/SS4END[12]
+ Tile_X2Y9_LUT4AB/SS4END[13] Tile_X2Y9_LUT4AB/SS4END[14] Tile_X2Y9_LUT4AB/SS4END[15]
+ Tile_X2Y9_LUT4AB/SS4END[1] Tile_X2Y9_LUT4AB/SS4END[2] Tile_X2Y9_LUT4AB/SS4END[3]
+ Tile_X2Y9_LUT4AB/SS4END[4] Tile_X2Y9_LUT4AB/SS4END[5] Tile_X2Y9_LUT4AB/SS4END[6]
+ Tile_X2Y9_LUT4AB/SS4END[7] Tile_X2Y9_LUT4AB/SS4END[8] Tile_X2Y9_LUT4AB/SS4END[9]
+ Tile_X2Y9_LUT4AB/UserCLK Tile_X2Y8_LUT4AB/UserCLK VGND VPWR Tile_X2Y9_LUT4AB/W1BEG[0]
+ Tile_X2Y9_LUT4AB/W1BEG[1] Tile_X2Y9_LUT4AB/W1BEG[2] Tile_X2Y9_LUT4AB/W1BEG[3] Tile_X3Y9_LUT4AB/W1BEG[0]
+ Tile_X3Y9_LUT4AB/W1BEG[1] Tile_X3Y9_LUT4AB/W1BEG[2] Tile_X3Y9_LUT4AB/W1BEG[3] Tile_X2Y9_LUT4AB/W2BEG[0]
+ Tile_X2Y9_LUT4AB/W2BEG[1] Tile_X2Y9_LUT4AB/W2BEG[2] Tile_X2Y9_LUT4AB/W2BEG[3] Tile_X2Y9_LUT4AB/W2BEG[4]
+ Tile_X2Y9_LUT4AB/W2BEG[5] Tile_X2Y9_LUT4AB/W2BEG[6] Tile_X2Y9_LUT4AB/W2BEG[7] Tile_X1Y9_LUT4AB/W2END[0]
+ Tile_X1Y9_LUT4AB/W2END[1] Tile_X1Y9_LUT4AB/W2END[2] Tile_X1Y9_LUT4AB/W2END[3] Tile_X1Y9_LUT4AB/W2END[4]
+ Tile_X1Y9_LUT4AB/W2END[5] Tile_X1Y9_LUT4AB/W2END[6] Tile_X1Y9_LUT4AB/W2END[7] Tile_X2Y9_LUT4AB/W2END[0]
+ Tile_X2Y9_LUT4AB/W2END[1] Tile_X2Y9_LUT4AB/W2END[2] Tile_X2Y9_LUT4AB/W2END[3] Tile_X2Y9_LUT4AB/W2END[4]
+ Tile_X2Y9_LUT4AB/W2END[5] Tile_X2Y9_LUT4AB/W2END[6] Tile_X2Y9_LUT4AB/W2END[7] Tile_X3Y9_LUT4AB/W2BEG[0]
+ Tile_X3Y9_LUT4AB/W2BEG[1] Tile_X3Y9_LUT4AB/W2BEG[2] Tile_X3Y9_LUT4AB/W2BEG[3] Tile_X3Y9_LUT4AB/W2BEG[4]
+ Tile_X3Y9_LUT4AB/W2BEG[5] Tile_X3Y9_LUT4AB/W2BEG[6] Tile_X3Y9_LUT4AB/W2BEG[7] Tile_X2Y9_LUT4AB/W6BEG[0]
+ Tile_X2Y9_LUT4AB/W6BEG[10] Tile_X2Y9_LUT4AB/W6BEG[11] Tile_X2Y9_LUT4AB/W6BEG[1]
+ Tile_X2Y9_LUT4AB/W6BEG[2] Tile_X2Y9_LUT4AB/W6BEG[3] Tile_X2Y9_LUT4AB/W6BEG[4] Tile_X2Y9_LUT4AB/W6BEG[5]
+ Tile_X2Y9_LUT4AB/W6BEG[6] Tile_X2Y9_LUT4AB/W6BEG[7] Tile_X2Y9_LUT4AB/W6BEG[8] Tile_X2Y9_LUT4AB/W6BEG[9]
+ Tile_X3Y9_LUT4AB/W6BEG[0] Tile_X3Y9_LUT4AB/W6BEG[10] Tile_X3Y9_LUT4AB/W6BEG[11]
+ Tile_X3Y9_LUT4AB/W6BEG[1] Tile_X3Y9_LUT4AB/W6BEG[2] Tile_X3Y9_LUT4AB/W6BEG[3] Tile_X3Y9_LUT4AB/W6BEG[4]
+ Tile_X3Y9_LUT4AB/W6BEG[5] Tile_X3Y9_LUT4AB/W6BEG[6] Tile_X3Y9_LUT4AB/W6BEG[7] Tile_X3Y9_LUT4AB/W6BEG[8]
+ Tile_X3Y9_LUT4AB/W6BEG[9] Tile_X2Y9_LUT4AB/WW4BEG[0] Tile_X2Y9_LUT4AB/WW4BEG[10]
+ Tile_X2Y9_LUT4AB/WW4BEG[11] Tile_X2Y9_LUT4AB/WW4BEG[12] Tile_X2Y9_LUT4AB/WW4BEG[13]
+ Tile_X2Y9_LUT4AB/WW4BEG[14] Tile_X2Y9_LUT4AB/WW4BEG[15] Tile_X2Y9_LUT4AB/WW4BEG[1]
+ Tile_X2Y9_LUT4AB/WW4BEG[2] Tile_X2Y9_LUT4AB/WW4BEG[3] Tile_X2Y9_LUT4AB/WW4BEG[4]
+ Tile_X2Y9_LUT4AB/WW4BEG[5] Tile_X2Y9_LUT4AB/WW4BEG[6] Tile_X2Y9_LUT4AB/WW4BEG[7]
+ Tile_X2Y9_LUT4AB/WW4BEG[8] Tile_X2Y9_LUT4AB/WW4BEG[9] Tile_X3Y9_LUT4AB/WW4BEG[0]
+ Tile_X3Y9_LUT4AB/WW4BEG[10] Tile_X3Y9_LUT4AB/WW4BEG[11] Tile_X3Y9_LUT4AB/WW4BEG[12]
+ Tile_X3Y9_LUT4AB/WW4BEG[13] Tile_X3Y9_LUT4AB/WW4BEG[14] Tile_X3Y9_LUT4AB/WW4BEG[15]
+ Tile_X3Y9_LUT4AB/WW4BEG[1] Tile_X3Y9_LUT4AB/WW4BEG[2] Tile_X3Y9_LUT4AB/WW4BEG[3]
+ Tile_X3Y9_LUT4AB/WW4BEG[4] Tile_X3Y9_LUT4AB/WW4BEG[5] Tile_X3Y9_LUT4AB/WW4BEG[6]
+ Tile_X3Y9_LUT4AB/WW4BEG[7] Tile_X3Y9_LUT4AB/WW4BEG[8] Tile_X3Y9_LUT4AB/WW4BEG[9]
+ LUT4AB
XTile_X7Y7_DSP Tile_X8Y7_LUT4AB/E1END[0] Tile_X8Y7_LUT4AB/E1END[1] Tile_X8Y7_LUT4AB/E1END[2]
+ Tile_X8Y7_LUT4AB/E1END[3] Tile_X6Y7_LUT4AB/E1BEG[0] Tile_X6Y7_LUT4AB/E1BEG[1] Tile_X6Y7_LUT4AB/E1BEG[2]
+ Tile_X6Y7_LUT4AB/E1BEG[3] Tile_X8Y7_LUT4AB/E2MID[0] Tile_X8Y7_LUT4AB/E2MID[1] Tile_X8Y7_LUT4AB/E2MID[2]
+ Tile_X8Y7_LUT4AB/E2MID[3] Tile_X8Y7_LUT4AB/E2MID[4] Tile_X8Y7_LUT4AB/E2MID[5] Tile_X8Y7_LUT4AB/E2MID[6]
+ Tile_X8Y7_LUT4AB/E2MID[7] Tile_X8Y7_LUT4AB/E2END[0] Tile_X8Y7_LUT4AB/E2END[1] Tile_X8Y7_LUT4AB/E2END[2]
+ Tile_X8Y7_LUT4AB/E2END[3] Tile_X8Y7_LUT4AB/E2END[4] Tile_X8Y7_LUT4AB/E2END[5] Tile_X8Y7_LUT4AB/E2END[6]
+ Tile_X8Y7_LUT4AB/E2END[7] Tile_X6Y7_LUT4AB/E2BEGb[0] Tile_X6Y7_LUT4AB/E2BEGb[1]
+ Tile_X6Y7_LUT4AB/E2BEGb[2] Tile_X6Y7_LUT4AB/E2BEGb[3] Tile_X6Y7_LUT4AB/E2BEGb[4]
+ Tile_X6Y7_LUT4AB/E2BEGb[5] Tile_X6Y7_LUT4AB/E2BEGb[6] Tile_X6Y7_LUT4AB/E2BEGb[7]
+ Tile_X6Y7_LUT4AB/E2BEG[0] Tile_X6Y7_LUT4AB/E2BEG[1] Tile_X6Y7_LUT4AB/E2BEG[2] Tile_X6Y7_LUT4AB/E2BEG[3]
+ Tile_X6Y7_LUT4AB/E2BEG[4] Tile_X6Y7_LUT4AB/E2BEG[5] Tile_X6Y7_LUT4AB/E2BEG[6] Tile_X6Y7_LUT4AB/E2BEG[7]
+ Tile_X8Y7_LUT4AB/E6END[0] Tile_X8Y7_LUT4AB/E6END[10] Tile_X8Y7_LUT4AB/E6END[11]
+ Tile_X8Y7_LUT4AB/E6END[1] Tile_X8Y7_LUT4AB/E6END[2] Tile_X8Y7_LUT4AB/E6END[3] Tile_X8Y7_LUT4AB/E6END[4]
+ Tile_X8Y7_LUT4AB/E6END[5] Tile_X8Y7_LUT4AB/E6END[6] Tile_X8Y7_LUT4AB/E6END[7] Tile_X8Y7_LUT4AB/E6END[8]
+ Tile_X8Y7_LUT4AB/E6END[9] Tile_X6Y7_LUT4AB/E6BEG[0] Tile_X6Y7_LUT4AB/E6BEG[10] Tile_X6Y7_LUT4AB/E6BEG[11]
+ Tile_X6Y7_LUT4AB/E6BEG[1] Tile_X6Y7_LUT4AB/E6BEG[2] Tile_X6Y7_LUT4AB/E6BEG[3] Tile_X6Y7_LUT4AB/E6BEG[4]
+ Tile_X6Y7_LUT4AB/E6BEG[5] Tile_X6Y7_LUT4AB/E6BEG[6] Tile_X6Y7_LUT4AB/E6BEG[7] Tile_X6Y7_LUT4AB/E6BEG[8]
+ Tile_X6Y7_LUT4AB/E6BEG[9] Tile_X8Y7_LUT4AB/EE4END[0] Tile_X8Y7_LUT4AB/EE4END[10]
+ Tile_X8Y7_LUT4AB/EE4END[11] Tile_X8Y7_LUT4AB/EE4END[12] Tile_X8Y7_LUT4AB/EE4END[13]
+ Tile_X8Y7_LUT4AB/EE4END[14] Tile_X8Y7_LUT4AB/EE4END[15] Tile_X8Y7_LUT4AB/EE4END[1]
+ Tile_X8Y7_LUT4AB/EE4END[2] Tile_X8Y7_LUT4AB/EE4END[3] Tile_X8Y7_LUT4AB/EE4END[4]
+ Tile_X8Y7_LUT4AB/EE4END[5] Tile_X8Y7_LUT4AB/EE4END[6] Tile_X8Y7_LUT4AB/EE4END[7]
+ Tile_X8Y7_LUT4AB/EE4END[8] Tile_X8Y7_LUT4AB/EE4END[9] Tile_X6Y7_LUT4AB/EE4BEG[0]
+ Tile_X6Y7_LUT4AB/EE4BEG[10] Tile_X6Y7_LUT4AB/EE4BEG[11] Tile_X6Y7_LUT4AB/EE4BEG[12]
+ Tile_X6Y7_LUT4AB/EE4BEG[13] Tile_X6Y7_LUT4AB/EE4BEG[14] Tile_X6Y7_LUT4AB/EE4BEG[15]
+ Tile_X6Y7_LUT4AB/EE4BEG[1] Tile_X6Y7_LUT4AB/EE4BEG[2] Tile_X6Y7_LUT4AB/EE4BEG[3]
+ Tile_X6Y7_LUT4AB/EE4BEG[4] Tile_X6Y7_LUT4AB/EE4BEG[5] Tile_X6Y7_LUT4AB/EE4BEG[6]
+ Tile_X6Y7_LUT4AB/EE4BEG[7] Tile_X6Y7_LUT4AB/EE4BEG[8] Tile_X6Y7_LUT4AB/EE4BEG[9]
+ Tile_X6Y7_LUT4AB/FrameData_O[0] Tile_X6Y7_LUT4AB/FrameData_O[10] Tile_X6Y7_LUT4AB/FrameData_O[11]
+ Tile_X6Y7_LUT4AB/FrameData_O[12] Tile_X6Y7_LUT4AB/FrameData_O[13] Tile_X6Y7_LUT4AB/FrameData_O[14]
+ Tile_X6Y7_LUT4AB/FrameData_O[15] Tile_X6Y7_LUT4AB/FrameData_O[16] Tile_X6Y7_LUT4AB/FrameData_O[17]
+ Tile_X6Y7_LUT4AB/FrameData_O[18] Tile_X6Y7_LUT4AB/FrameData_O[19] Tile_X6Y7_LUT4AB/FrameData_O[1]
+ Tile_X6Y7_LUT4AB/FrameData_O[20] Tile_X6Y7_LUT4AB/FrameData_O[21] Tile_X6Y7_LUT4AB/FrameData_O[22]
+ Tile_X6Y7_LUT4AB/FrameData_O[23] Tile_X6Y7_LUT4AB/FrameData_O[24] Tile_X6Y7_LUT4AB/FrameData_O[25]
+ Tile_X6Y7_LUT4AB/FrameData_O[26] Tile_X6Y7_LUT4AB/FrameData_O[27] Tile_X6Y7_LUT4AB/FrameData_O[28]
+ Tile_X6Y7_LUT4AB/FrameData_O[29] Tile_X6Y7_LUT4AB/FrameData_O[2] Tile_X6Y7_LUT4AB/FrameData_O[30]
+ Tile_X6Y7_LUT4AB/FrameData_O[31] Tile_X6Y7_LUT4AB/FrameData_O[3] Tile_X6Y7_LUT4AB/FrameData_O[4]
+ Tile_X6Y7_LUT4AB/FrameData_O[5] Tile_X6Y7_LUT4AB/FrameData_O[6] Tile_X6Y7_LUT4AB/FrameData_O[7]
+ Tile_X6Y7_LUT4AB/FrameData_O[8] Tile_X6Y7_LUT4AB/FrameData_O[9] Tile_X8Y7_LUT4AB/FrameData[0]
+ Tile_X8Y7_LUT4AB/FrameData[10] Tile_X8Y7_LUT4AB/FrameData[11] Tile_X8Y7_LUT4AB/FrameData[12]
+ Tile_X8Y7_LUT4AB/FrameData[13] Tile_X8Y7_LUT4AB/FrameData[14] Tile_X8Y7_LUT4AB/FrameData[15]
+ Tile_X8Y7_LUT4AB/FrameData[16] Tile_X8Y7_LUT4AB/FrameData[17] Tile_X8Y7_LUT4AB/FrameData[18]
+ Tile_X8Y7_LUT4AB/FrameData[19] Tile_X8Y7_LUT4AB/FrameData[1] Tile_X8Y7_LUT4AB/FrameData[20]
+ Tile_X8Y7_LUT4AB/FrameData[21] Tile_X8Y7_LUT4AB/FrameData[22] Tile_X8Y7_LUT4AB/FrameData[23]
+ Tile_X8Y7_LUT4AB/FrameData[24] Tile_X8Y7_LUT4AB/FrameData[25] Tile_X8Y7_LUT4AB/FrameData[26]
+ Tile_X8Y7_LUT4AB/FrameData[27] Tile_X8Y7_LUT4AB/FrameData[28] Tile_X8Y7_LUT4AB/FrameData[29]
+ Tile_X8Y7_LUT4AB/FrameData[2] Tile_X8Y7_LUT4AB/FrameData[30] Tile_X8Y7_LUT4AB/FrameData[31]
+ Tile_X8Y7_LUT4AB/FrameData[3] Tile_X8Y7_LUT4AB/FrameData[4] Tile_X8Y7_LUT4AB/FrameData[5]
+ Tile_X8Y7_LUT4AB/FrameData[6] Tile_X8Y7_LUT4AB/FrameData[7] Tile_X8Y7_LUT4AB/FrameData[8]
+ Tile_X8Y7_LUT4AB/FrameData[9] Tile_X7Y5_DSP/Tile_X0Y1_FrameStrobe[0] Tile_X7Y5_DSP/Tile_X0Y1_FrameStrobe[10]
+ Tile_X7Y5_DSP/Tile_X0Y1_FrameStrobe[11] Tile_X7Y5_DSP/Tile_X0Y1_FrameStrobe[12]
+ Tile_X7Y5_DSP/Tile_X0Y1_FrameStrobe[13] Tile_X7Y5_DSP/Tile_X0Y1_FrameStrobe[14]
+ Tile_X7Y5_DSP/Tile_X0Y1_FrameStrobe[15] Tile_X7Y5_DSP/Tile_X0Y1_FrameStrobe[16]
+ Tile_X7Y5_DSP/Tile_X0Y1_FrameStrobe[17] Tile_X7Y5_DSP/Tile_X0Y1_FrameStrobe[18]
+ Tile_X7Y5_DSP/Tile_X0Y1_FrameStrobe[19] Tile_X7Y5_DSP/Tile_X0Y1_FrameStrobe[1] Tile_X7Y5_DSP/Tile_X0Y1_FrameStrobe[2]
+ Tile_X7Y5_DSP/Tile_X0Y1_FrameStrobe[3] Tile_X7Y5_DSP/Tile_X0Y1_FrameStrobe[4] Tile_X7Y5_DSP/Tile_X0Y1_FrameStrobe[5]
+ Tile_X7Y5_DSP/Tile_X0Y1_FrameStrobe[6] Tile_X7Y5_DSP/Tile_X0Y1_FrameStrobe[7] Tile_X7Y5_DSP/Tile_X0Y1_FrameStrobe[8]
+ Tile_X7Y5_DSP/Tile_X0Y1_FrameStrobe[9] Tile_X7Y7_DSP/Tile_X0Y0_N1BEG[0] Tile_X7Y7_DSP/Tile_X0Y0_N1BEG[1]
+ Tile_X7Y7_DSP/Tile_X0Y0_N1BEG[2] Tile_X7Y7_DSP/Tile_X0Y0_N1BEG[3] Tile_X7Y7_DSP/Tile_X0Y0_N2BEG[0]
+ Tile_X7Y7_DSP/Tile_X0Y0_N2BEG[1] Tile_X7Y7_DSP/Tile_X0Y0_N2BEG[2] Tile_X7Y7_DSP/Tile_X0Y0_N2BEG[3]
+ Tile_X7Y7_DSP/Tile_X0Y0_N2BEG[4] Tile_X7Y7_DSP/Tile_X0Y0_N2BEG[5] Tile_X7Y7_DSP/Tile_X0Y0_N2BEG[6]
+ Tile_X7Y7_DSP/Tile_X0Y0_N2BEG[7] Tile_X7Y5_DSP/Tile_X0Y1_N2END[0] Tile_X7Y5_DSP/Tile_X0Y1_N2END[1]
+ Tile_X7Y5_DSP/Tile_X0Y1_N2END[2] Tile_X7Y5_DSP/Tile_X0Y1_N2END[3] Tile_X7Y5_DSP/Tile_X0Y1_N2END[4]
+ Tile_X7Y5_DSP/Tile_X0Y1_N2END[5] Tile_X7Y5_DSP/Tile_X0Y1_N2END[6] Tile_X7Y5_DSP/Tile_X0Y1_N2END[7]
+ Tile_X7Y7_DSP/Tile_X0Y0_N4BEG[0] Tile_X7Y7_DSP/Tile_X0Y0_N4BEG[10] Tile_X7Y7_DSP/Tile_X0Y0_N4BEG[11]
+ Tile_X7Y7_DSP/Tile_X0Y0_N4BEG[12] Tile_X7Y7_DSP/Tile_X0Y0_N4BEG[13] Tile_X7Y7_DSP/Tile_X0Y0_N4BEG[14]
+ Tile_X7Y7_DSP/Tile_X0Y0_N4BEG[15] Tile_X7Y7_DSP/Tile_X0Y0_N4BEG[1] Tile_X7Y7_DSP/Tile_X0Y0_N4BEG[2]
+ Tile_X7Y7_DSP/Tile_X0Y0_N4BEG[3] Tile_X7Y7_DSP/Tile_X0Y0_N4BEG[4] Tile_X7Y7_DSP/Tile_X0Y0_N4BEG[5]
+ Tile_X7Y7_DSP/Tile_X0Y0_N4BEG[6] Tile_X7Y7_DSP/Tile_X0Y0_N4BEG[7] Tile_X7Y7_DSP/Tile_X0Y0_N4BEG[8]
+ Tile_X7Y7_DSP/Tile_X0Y0_N4BEG[9] Tile_X7Y7_DSP/Tile_X0Y0_NN4BEG[0] Tile_X7Y7_DSP/Tile_X0Y0_NN4BEG[10]
+ Tile_X7Y7_DSP/Tile_X0Y0_NN4BEG[11] Tile_X7Y7_DSP/Tile_X0Y0_NN4BEG[12] Tile_X7Y7_DSP/Tile_X0Y0_NN4BEG[13]
+ Tile_X7Y7_DSP/Tile_X0Y0_NN4BEG[14] Tile_X7Y7_DSP/Tile_X0Y0_NN4BEG[15] Tile_X7Y7_DSP/Tile_X0Y0_NN4BEG[1]
+ Tile_X7Y7_DSP/Tile_X0Y0_NN4BEG[2] Tile_X7Y7_DSP/Tile_X0Y0_NN4BEG[3] Tile_X7Y7_DSP/Tile_X0Y0_NN4BEG[4]
+ Tile_X7Y7_DSP/Tile_X0Y0_NN4BEG[5] Tile_X7Y7_DSP/Tile_X0Y0_NN4BEG[6] Tile_X7Y7_DSP/Tile_X0Y0_NN4BEG[7]
+ Tile_X7Y7_DSP/Tile_X0Y0_NN4BEG[8] Tile_X7Y7_DSP/Tile_X0Y0_NN4BEG[9] Tile_X7Y7_DSP/Tile_X0Y0_S1END[0]
+ Tile_X7Y7_DSP/Tile_X0Y0_S1END[1] Tile_X7Y7_DSP/Tile_X0Y0_S1END[2] Tile_X7Y7_DSP/Tile_X0Y0_S1END[3]
+ Tile_X7Y7_DSP/Tile_X0Y0_S2END[0] Tile_X7Y7_DSP/Tile_X0Y0_S2END[1] Tile_X7Y7_DSP/Tile_X0Y0_S2END[2]
+ Tile_X7Y7_DSP/Tile_X0Y0_S2END[3] Tile_X7Y7_DSP/Tile_X0Y0_S2END[4] Tile_X7Y7_DSP/Tile_X0Y0_S2END[5]
+ Tile_X7Y7_DSP/Tile_X0Y0_S2END[6] Tile_X7Y7_DSP/Tile_X0Y0_S2END[7] Tile_X7Y7_DSP/Tile_X0Y0_S2MID[0]
+ Tile_X7Y7_DSP/Tile_X0Y0_S2MID[1] Tile_X7Y7_DSP/Tile_X0Y0_S2MID[2] Tile_X7Y7_DSP/Tile_X0Y0_S2MID[3]
+ Tile_X7Y7_DSP/Tile_X0Y0_S2MID[4] Tile_X7Y7_DSP/Tile_X0Y0_S2MID[5] Tile_X7Y7_DSP/Tile_X0Y0_S2MID[6]
+ Tile_X7Y7_DSP/Tile_X0Y0_S2MID[7] Tile_X7Y7_DSP/Tile_X0Y0_S4END[0] Tile_X7Y7_DSP/Tile_X0Y0_S4END[10]
+ Tile_X7Y7_DSP/Tile_X0Y0_S4END[11] Tile_X7Y7_DSP/Tile_X0Y0_S4END[12] Tile_X7Y7_DSP/Tile_X0Y0_S4END[13]
+ Tile_X7Y7_DSP/Tile_X0Y0_S4END[14] Tile_X7Y7_DSP/Tile_X0Y0_S4END[15] Tile_X7Y7_DSP/Tile_X0Y0_S4END[1]
+ Tile_X7Y7_DSP/Tile_X0Y0_S4END[2] Tile_X7Y7_DSP/Tile_X0Y0_S4END[3] Tile_X7Y7_DSP/Tile_X0Y0_S4END[4]
+ Tile_X7Y7_DSP/Tile_X0Y0_S4END[5] Tile_X7Y7_DSP/Tile_X0Y0_S4END[6] Tile_X7Y7_DSP/Tile_X0Y0_S4END[7]
+ Tile_X7Y7_DSP/Tile_X0Y0_S4END[8] Tile_X7Y7_DSP/Tile_X0Y0_S4END[9] Tile_X7Y7_DSP/Tile_X0Y0_SS4END[0]
+ Tile_X7Y7_DSP/Tile_X0Y0_SS4END[10] Tile_X7Y7_DSP/Tile_X0Y0_SS4END[11] Tile_X7Y7_DSP/Tile_X0Y0_SS4END[12]
+ Tile_X7Y7_DSP/Tile_X0Y0_SS4END[13] Tile_X7Y7_DSP/Tile_X0Y0_SS4END[14] Tile_X7Y7_DSP/Tile_X0Y0_SS4END[15]
+ Tile_X7Y7_DSP/Tile_X0Y0_SS4END[1] Tile_X7Y7_DSP/Tile_X0Y0_SS4END[2] Tile_X7Y7_DSP/Tile_X0Y0_SS4END[3]
+ Tile_X7Y7_DSP/Tile_X0Y0_SS4END[4] Tile_X7Y7_DSP/Tile_X0Y0_SS4END[5] Tile_X7Y7_DSP/Tile_X0Y0_SS4END[6]
+ Tile_X7Y7_DSP/Tile_X0Y0_SS4END[7] Tile_X7Y7_DSP/Tile_X0Y0_SS4END[8] Tile_X7Y7_DSP/Tile_X0Y0_SS4END[9]
+ Tile_X7Y5_DSP/Tile_X0Y1_UserCLK Tile_X6Y7_LUT4AB/W1END[0] Tile_X6Y7_LUT4AB/W1END[1]
+ Tile_X6Y7_LUT4AB/W1END[2] Tile_X6Y7_LUT4AB/W1END[3] Tile_X8Y7_LUT4AB/W1BEG[0] Tile_X8Y7_LUT4AB/W1BEG[1]
+ Tile_X8Y7_LUT4AB/W1BEG[2] Tile_X8Y7_LUT4AB/W1BEG[3] Tile_X6Y7_LUT4AB/W2MID[0] Tile_X6Y7_LUT4AB/W2MID[1]
+ Tile_X6Y7_LUT4AB/W2MID[2] Tile_X6Y7_LUT4AB/W2MID[3] Tile_X6Y7_LUT4AB/W2MID[4] Tile_X6Y7_LUT4AB/W2MID[5]
+ Tile_X6Y7_LUT4AB/W2MID[6] Tile_X6Y7_LUT4AB/W2MID[7] Tile_X6Y7_LUT4AB/W2END[0] Tile_X6Y7_LUT4AB/W2END[1]
+ Tile_X6Y7_LUT4AB/W2END[2] Tile_X6Y7_LUT4AB/W2END[3] Tile_X6Y7_LUT4AB/W2END[4] Tile_X6Y7_LUT4AB/W2END[5]
+ Tile_X6Y7_LUT4AB/W2END[6] Tile_X6Y7_LUT4AB/W2END[7] Tile_X8Y7_LUT4AB/W2BEGb[0] Tile_X8Y7_LUT4AB/W2BEGb[1]
+ Tile_X8Y7_LUT4AB/W2BEGb[2] Tile_X8Y7_LUT4AB/W2BEGb[3] Tile_X8Y7_LUT4AB/W2BEGb[4]
+ Tile_X8Y7_LUT4AB/W2BEGb[5] Tile_X8Y7_LUT4AB/W2BEGb[6] Tile_X8Y7_LUT4AB/W2BEGb[7]
+ Tile_X8Y7_LUT4AB/W2BEG[0] Tile_X8Y7_LUT4AB/W2BEG[1] Tile_X8Y7_LUT4AB/W2BEG[2] Tile_X8Y7_LUT4AB/W2BEG[3]
+ Tile_X8Y7_LUT4AB/W2BEG[4] Tile_X8Y7_LUT4AB/W2BEG[5] Tile_X8Y7_LUT4AB/W2BEG[6] Tile_X8Y7_LUT4AB/W2BEG[7]
+ Tile_X6Y7_LUT4AB/W6END[0] Tile_X6Y7_LUT4AB/W6END[10] Tile_X6Y7_LUT4AB/W6END[11]
+ Tile_X6Y7_LUT4AB/W6END[1] Tile_X6Y7_LUT4AB/W6END[2] Tile_X6Y7_LUT4AB/W6END[3] Tile_X6Y7_LUT4AB/W6END[4]
+ Tile_X6Y7_LUT4AB/W6END[5] Tile_X6Y7_LUT4AB/W6END[6] Tile_X6Y7_LUT4AB/W6END[7] Tile_X6Y7_LUT4AB/W6END[8]
+ Tile_X6Y7_LUT4AB/W6END[9] Tile_X8Y7_LUT4AB/W6BEG[0] Tile_X8Y7_LUT4AB/W6BEG[10] Tile_X8Y7_LUT4AB/W6BEG[11]
+ Tile_X8Y7_LUT4AB/W6BEG[1] Tile_X8Y7_LUT4AB/W6BEG[2] Tile_X8Y7_LUT4AB/W6BEG[3] Tile_X8Y7_LUT4AB/W6BEG[4]
+ Tile_X8Y7_LUT4AB/W6BEG[5] Tile_X8Y7_LUT4AB/W6BEG[6] Tile_X8Y7_LUT4AB/W6BEG[7] Tile_X8Y7_LUT4AB/W6BEG[8]
+ Tile_X8Y7_LUT4AB/W6BEG[9] Tile_X6Y7_LUT4AB/WW4END[0] Tile_X6Y7_LUT4AB/WW4END[10]
+ Tile_X6Y7_LUT4AB/WW4END[11] Tile_X6Y7_LUT4AB/WW4END[12] Tile_X6Y7_LUT4AB/WW4END[13]
+ Tile_X6Y7_LUT4AB/WW4END[14] Tile_X6Y7_LUT4AB/WW4END[15] Tile_X6Y7_LUT4AB/WW4END[1]
+ Tile_X6Y7_LUT4AB/WW4END[2] Tile_X6Y7_LUT4AB/WW4END[3] Tile_X6Y7_LUT4AB/WW4END[4]
+ Tile_X6Y7_LUT4AB/WW4END[5] Tile_X6Y7_LUT4AB/WW4END[6] Tile_X6Y7_LUT4AB/WW4END[7]
+ Tile_X6Y7_LUT4AB/WW4END[8] Tile_X6Y7_LUT4AB/WW4END[9] Tile_X8Y7_LUT4AB/WW4BEG[0]
+ Tile_X8Y7_LUT4AB/WW4BEG[10] Tile_X8Y7_LUT4AB/WW4BEG[11] Tile_X8Y7_LUT4AB/WW4BEG[12]
+ Tile_X8Y7_LUT4AB/WW4BEG[13] Tile_X8Y7_LUT4AB/WW4BEG[14] Tile_X8Y7_LUT4AB/WW4BEG[15]
+ Tile_X8Y7_LUT4AB/WW4BEG[1] Tile_X8Y7_LUT4AB/WW4BEG[2] Tile_X8Y7_LUT4AB/WW4BEG[3]
+ Tile_X8Y7_LUT4AB/WW4BEG[4] Tile_X8Y7_LUT4AB/WW4BEG[5] Tile_X8Y7_LUT4AB/WW4BEG[6]
+ Tile_X8Y7_LUT4AB/WW4BEG[7] Tile_X8Y7_LUT4AB/WW4BEG[8] Tile_X8Y7_LUT4AB/WW4BEG[9]
+ Tile_X8Y8_LUT4AB/E1END[0] Tile_X8Y8_LUT4AB/E1END[1] Tile_X8Y8_LUT4AB/E1END[2] Tile_X8Y8_LUT4AB/E1END[3]
+ Tile_X6Y8_LUT4AB/E1BEG[0] Tile_X6Y8_LUT4AB/E1BEG[1] Tile_X6Y8_LUT4AB/E1BEG[2] Tile_X6Y8_LUT4AB/E1BEG[3]
+ Tile_X8Y8_LUT4AB/E2MID[0] Tile_X8Y8_LUT4AB/E2MID[1] Tile_X8Y8_LUT4AB/E2MID[2] Tile_X8Y8_LUT4AB/E2MID[3]
+ Tile_X8Y8_LUT4AB/E2MID[4] Tile_X8Y8_LUT4AB/E2MID[5] Tile_X8Y8_LUT4AB/E2MID[6] Tile_X8Y8_LUT4AB/E2MID[7]
+ Tile_X8Y8_LUT4AB/E2END[0] Tile_X8Y8_LUT4AB/E2END[1] Tile_X8Y8_LUT4AB/E2END[2] Tile_X8Y8_LUT4AB/E2END[3]
+ Tile_X8Y8_LUT4AB/E2END[4] Tile_X8Y8_LUT4AB/E2END[5] Tile_X8Y8_LUT4AB/E2END[6] Tile_X8Y8_LUT4AB/E2END[7]
+ Tile_X6Y8_LUT4AB/E2BEGb[0] Tile_X6Y8_LUT4AB/E2BEGb[1] Tile_X6Y8_LUT4AB/E2BEGb[2]
+ Tile_X6Y8_LUT4AB/E2BEGb[3] Tile_X6Y8_LUT4AB/E2BEGb[4] Tile_X6Y8_LUT4AB/E2BEGb[5]
+ Tile_X6Y8_LUT4AB/E2BEGb[6] Tile_X6Y8_LUT4AB/E2BEGb[7] Tile_X6Y8_LUT4AB/E2BEG[0]
+ Tile_X6Y8_LUT4AB/E2BEG[1] Tile_X6Y8_LUT4AB/E2BEG[2] Tile_X6Y8_LUT4AB/E2BEG[3] Tile_X6Y8_LUT4AB/E2BEG[4]
+ Tile_X6Y8_LUT4AB/E2BEG[5] Tile_X6Y8_LUT4AB/E2BEG[6] Tile_X6Y8_LUT4AB/E2BEG[7] Tile_X8Y8_LUT4AB/E6END[0]
+ Tile_X8Y8_LUT4AB/E6END[10] Tile_X8Y8_LUT4AB/E6END[11] Tile_X8Y8_LUT4AB/E6END[1]
+ Tile_X8Y8_LUT4AB/E6END[2] Tile_X8Y8_LUT4AB/E6END[3] Tile_X8Y8_LUT4AB/E6END[4] Tile_X8Y8_LUT4AB/E6END[5]
+ Tile_X8Y8_LUT4AB/E6END[6] Tile_X8Y8_LUT4AB/E6END[7] Tile_X8Y8_LUT4AB/E6END[8] Tile_X8Y8_LUT4AB/E6END[9]
+ Tile_X6Y8_LUT4AB/E6BEG[0] Tile_X6Y8_LUT4AB/E6BEG[10] Tile_X6Y8_LUT4AB/E6BEG[11]
+ Tile_X6Y8_LUT4AB/E6BEG[1] Tile_X6Y8_LUT4AB/E6BEG[2] Tile_X6Y8_LUT4AB/E6BEG[3] Tile_X6Y8_LUT4AB/E6BEG[4]
+ Tile_X6Y8_LUT4AB/E6BEG[5] Tile_X6Y8_LUT4AB/E6BEG[6] Tile_X6Y8_LUT4AB/E6BEG[7] Tile_X6Y8_LUT4AB/E6BEG[8]
+ Tile_X6Y8_LUT4AB/E6BEG[9] Tile_X8Y8_LUT4AB/EE4END[0] Tile_X8Y8_LUT4AB/EE4END[10]
+ Tile_X8Y8_LUT4AB/EE4END[11] Tile_X8Y8_LUT4AB/EE4END[12] Tile_X8Y8_LUT4AB/EE4END[13]
+ Tile_X8Y8_LUT4AB/EE4END[14] Tile_X8Y8_LUT4AB/EE4END[15] Tile_X8Y8_LUT4AB/EE4END[1]
+ Tile_X8Y8_LUT4AB/EE4END[2] Tile_X8Y8_LUT4AB/EE4END[3] Tile_X8Y8_LUT4AB/EE4END[4]
+ Tile_X8Y8_LUT4AB/EE4END[5] Tile_X8Y8_LUT4AB/EE4END[6] Tile_X8Y8_LUT4AB/EE4END[7]
+ Tile_X8Y8_LUT4AB/EE4END[8] Tile_X8Y8_LUT4AB/EE4END[9] Tile_X6Y8_LUT4AB/EE4BEG[0]
+ Tile_X6Y8_LUT4AB/EE4BEG[10] Tile_X6Y8_LUT4AB/EE4BEG[11] Tile_X6Y8_LUT4AB/EE4BEG[12]
+ Tile_X6Y8_LUT4AB/EE4BEG[13] Tile_X6Y8_LUT4AB/EE4BEG[14] Tile_X6Y8_LUT4AB/EE4BEG[15]
+ Tile_X6Y8_LUT4AB/EE4BEG[1] Tile_X6Y8_LUT4AB/EE4BEG[2] Tile_X6Y8_LUT4AB/EE4BEG[3]
+ Tile_X6Y8_LUT4AB/EE4BEG[4] Tile_X6Y8_LUT4AB/EE4BEG[5] Tile_X6Y8_LUT4AB/EE4BEG[6]
+ Tile_X6Y8_LUT4AB/EE4BEG[7] Tile_X6Y8_LUT4AB/EE4BEG[8] Tile_X6Y8_LUT4AB/EE4BEG[9]
+ Tile_X6Y8_LUT4AB/FrameData_O[0] Tile_X6Y8_LUT4AB/FrameData_O[10] Tile_X6Y8_LUT4AB/FrameData_O[11]
+ Tile_X6Y8_LUT4AB/FrameData_O[12] Tile_X6Y8_LUT4AB/FrameData_O[13] Tile_X6Y8_LUT4AB/FrameData_O[14]
+ Tile_X6Y8_LUT4AB/FrameData_O[15] Tile_X6Y8_LUT4AB/FrameData_O[16] Tile_X6Y8_LUT4AB/FrameData_O[17]
+ Tile_X6Y8_LUT4AB/FrameData_O[18] Tile_X6Y8_LUT4AB/FrameData_O[19] Tile_X6Y8_LUT4AB/FrameData_O[1]
+ Tile_X6Y8_LUT4AB/FrameData_O[20] Tile_X6Y8_LUT4AB/FrameData_O[21] Tile_X6Y8_LUT4AB/FrameData_O[22]
+ Tile_X6Y8_LUT4AB/FrameData_O[23] Tile_X6Y8_LUT4AB/FrameData_O[24] Tile_X6Y8_LUT4AB/FrameData_O[25]
+ Tile_X6Y8_LUT4AB/FrameData_O[26] Tile_X6Y8_LUT4AB/FrameData_O[27] Tile_X6Y8_LUT4AB/FrameData_O[28]
+ Tile_X6Y8_LUT4AB/FrameData_O[29] Tile_X6Y8_LUT4AB/FrameData_O[2] Tile_X6Y8_LUT4AB/FrameData_O[30]
+ Tile_X6Y8_LUT4AB/FrameData_O[31] Tile_X6Y8_LUT4AB/FrameData_O[3] Tile_X6Y8_LUT4AB/FrameData_O[4]
+ Tile_X6Y8_LUT4AB/FrameData_O[5] Tile_X6Y8_LUT4AB/FrameData_O[6] Tile_X6Y8_LUT4AB/FrameData_O[7]
+ Tile_X6Y8_LUT4AB/FrameData_O[8] Tile_X6Y8_LUT4AB/FrameData_O[9] Tile_X8Y8_LUT4AB/FrameData[0]
+ Tile_X8Y8_LUT4AB/FrameData[10] Tile_X8Y8_LUT4AB/FrameData[11] Tile_X8Y8_LUT4AB/FrameData[12]
+ Tile_X8Y8_LUT4AB/FrameData[13] Tile_X8Y8_LUT4AB/FrameData[14] Tile_X8Y8_LUT4AB/FrameData[15]
+ Tile_X8Y8_LUT4AB/FrameData[16] Tile_X8Y8_LUT4AB/FrameData[17] Tile_X8Y8_LUT4AB/FrameData[18]
+ Tile_X8Y8_LUT4AB/FrameData[19] Tile_X8Y8_LUT4AB/FrameData[1] Tile_X8Y8_LUT4AB/FrameData[20]
+ Tile_X8Y8_LUT4AB/FrameData[21] Tile_X8Y8_LUT4AB/FrameData[22] Tile_X8Y8_LUT4AB/FrameData[23]
+ Tile_X8Y8_LUT4AB/FrameData[24] Tile_X8Y8_LUT4AB/FrameData[25] Tile_X8Y8_LUT4AB/FrameData[26]
+ Tile_X8Y8_LUT4AB/FrameData[27] Tile_X8Y8_LUT4AB/FrameData[28] Tile_X8Y8_LUT4AB/FrameData[29]
+ Tile_X8Y8_LUT4AB/FrameData[2] Tile_X8Y8_LUT4AB/FrameData[30] Tile_X8Y8_LUT4AB/FrameData[31]
+ Tile_X8Y8_LUT4AB/FrameData[3] Tile_X8Y8_LUT4AB/FrameData[4] Tile_X8Y8_LUT4AB/FrameData[5]
+ Tile_X8Y8_LUT4AB/FrameData[6] Tile_X8Y8_LUT4AB/FrameData[7] Tile_X8Y8_LUT4AB/FrameData[8]
+ Tile_X8Y8_LUT4AB/FrameData[9] Tile_X7Y7_DSP/Tile_X0Y1_FrameStrobe[0] Tile_X7Y7_DSP/Tile_X0Y1_FrameStrobe[10]
+ Tile_X7Y7_DSP/Tile_X0Y1_FrameStrobe[11] Tile_X7Y7_DSP/Tile_X0Y1_FrameStrobe[12]
+ Tile_X7Y7_DSP/Tile_X0Y1_FrameStrobe[13] Tile_X7Y7_DSP/Tile_X0Y1_FrameStrobe[14]
+ Tile_X7Y7_DSP/Tile_X0Y1_FrameStrobe[15] Tile_X7Y7_DSP/Tile_X0Y1_FrameStrobe[16]
+ Tile_X7Y7_DSP/Tile_X0Y1_FrameStrobe[17] Tile_X7Y7_DSP/Tile_X0Y1_FrameStrobe[18]
+ Tile_X7Y7_DSP/Tile_X0Y1_FrameStrobe[19] Tile_X7Y7_DSP/Tile_X0Y1_FrameStrobe[1] Tile_X7Y7_DSP/Tile_X0Y1_FrameStrobe[2]
+ Tile_X7Y7_DSP/Tile_X0Y1_FrameStrobe[3] Tile_X7Y7_DSP/Tile_X0Y1_FrameStrobe[4] Tile_X7Y7_DSP/Tile_X0Y1_FrameStrobe[5]
+ Tile_X7Y7_DSP/Tile_X0Y1_FrameStrobe[6] Tile_X7Y7_DSP/Tile_X0Y1_FrameStrobe[7] Tile_X7Y7_DSP/Tile_X0Y1_FrameStrobe[8]
+ Tile_X7Y7_DSP/Tile_X0Y1_FrameStrobe[9] Tile_X7Y9_DSP/Tile_X0Y0_N1BEG[0] Tile_X7Y9_DSP/Tile_X0Y0_N1BEG[1]
+ Tile_X7Y9_DSP/Tile_X0Y0_N1BEG[2] Tile_X7Y9_DSP/Tile_X0Y0_N1BEG[3] Tile_X7Y7_DSP/Tile_X0Y1_N2END[0]
+ Tile_X7Y7_DSP/Tile_X0Y1_N2END[1] Tile_X7Y7_DSP/Tile_X0Y1_N2END[2] Tile_X7Y7_DSP/Tile_X0Y1_N2END[3]
+ Tile_X7Y7_DSP/Tile_X0Y1_N2END[4] Tile_X7Y7_DSP/Tile_X0Y1_N2END[5] Tile_X7Y7_DSP/Tile_X0Y1_N2END[6]
+ Tile_X7Y7_DSP/Tile_X0Y1_N2END[7] Tile_X7Y9_DSP/Tile_X0Y0_N2BEG[0] Tile_X7Y9_DSP/Tile_X0Y0_N2BEG[1]
+ Tile_X7Y9_DSP/Tile_X0Y0_N2BEG[2] Tile_X7Y9_DSP/Tile_X0Y0_N2BEG[3] Tile_X7Y9_DSP/Tile_X0Y0_N2BEG[4]
+ Tile_X7Y9_DSP/Tile_X0Y0_N2BEG[5] Tile_X7Y9_DSP/Tile_X0Y0_N2BEG[6] Tile_X7Y9_DSP/Tile_X0Y0_N2BEG[7]
+ Tile_X7Y9_DSP/Tile_X0Y0_N4BEG[0] Tile_X7Y9_DSP/Tile_X0Y0_N4BEG[10] Tile_X7Y9_DSP/Tile_X0Y0_N4BEG[11]
+ Tile_X7Y9_DSP/Tile_X0Y0_N4BEG[12] Tile_X7Y9_DSP/Tile_X0Y0_N4BEG[13] Tile_X7Y9_DSP/Tile_X0Y0_N4BEG[14]
+ Tile_X7Y9_DSP/Tile_X0Y0_N4BEG[15] Tile_X7Y9_DSP/Tile_X0Y0_N4BEG[1] Tile_X7Y9_DSP/Tile_X0Y0_N4BEG[2]
+ Tile_X7Y9_DSP/Tile_X0Y0_N4BEG[3] Tile_X7Y9_DSP/Tile_X0Y0_N4BEG[4] Tile_X7Y9_DSP/Tile_X0Y0_N4BEG[5]
+ Tile_X7Y9_DSP/Tile_X0Y0_N4BEG[6] Tile_X7Y9_DSP/Tile_X0Y0_N4BEG[7] Tile_X7Y9_DSP/Tile_X0Y0_N4BEG[8]
+ Tile_X7Y9_DSP/Tile_X0Y0_N4BEG[9] Tile_X7Y9_DSP/Tile_X0Y0_NN4BEG[0] Tile_X7Y9_DSP/Tile_X0Y0_NN4BEG[10]
+ Tile_X7Y9_DSP/Tile_X0Y0_NN4BEG[11] Tile_X7Y9_DSP/Tile_X0Y0_NN4BEG[12] Tile_X7Y9_DSP/Tile_X0Y0_NN4BEG[13]
+ Tile_X7Y9_DSP/Tile_X0Y0_NN4BEG[14] Tile_X7Y9_DSP/Tile_X0Y0_NN4BEG[15] Tile_X7Y9_DSP/Tile_X0Y0_NN4BEG[1]
+ Tile_X7Y9_DSP/Tile_X0Y0_NN4BEG[2] Tile_X7Y9_DSP/Tile_X0Y0_NN4BEG[3] Tile_X7Y9_DSP/Tile_X0Y0_NN4BEG[4]
+ Tile_X7Y9_DSP/Tile_X0Y0_NN4BEG[5] Tile_X7Y9_DSP/Tile_X0Y0_NN4BEG[6] Tile_X7Y9_DSP/Tile_X0Y0_NN4BEG[7]
+ Tile_X7Y9_DSP/Tile_X0Y0_NN4BEG[8] Tile_X7Y9_DSP/Tile_X0Y0_NN4BEG[9] Tile_X7Y9_DSP/Tile_X0Y0_S1END[0]
+ Tile_X7Y9_DSP/Tile_X0Y0_S1END[1] Tile_X7Y9_DSP/Tile_X0Y0_S1END[2] Tile_X7Y9_DSP/Tile_X0Y0_S1END[3]
+ Tile_X7Y9_DSP/Tile_X0Y0_S2MID[0] Tile_X7Y9_DSP/Tile_X0Y0_S2MID[1] Tile_X7Y9_DSP/Tile_X0Y0_S2MID[2]
+ Tile_X7Y9_DSP/Tile_X0Y0_S2MID[3] Tile_X7Y9_DSP/Tile_X0Y0_S2MID[4] Tile_X7Y9_DSP/Tile_X0Y0_S2MID[5]
+ Tile_X7Y9_DSP/Tile_X0Y0_S2MID[6] Tile_X7Y9_DSP/Tile_X0Y0_S2MID[7] Tile_X7Y9_DSP/Tile_X0Y0_S2END[0]
+ Tile_X7Y9_DSP/Tile_X0Y0_S2END[1] Tile_X7Y9_DSP/Tile_X0Y0_S2END[2] Tile_X7Y9_DSP/Tile_X0Y0_S2END[3]
+ Tile_X7Y9_DSP/Tile_X0Y0_S2END[4] Tile_X7Y9_DSP/Tile_X0Y0_S2END[5] Tile_X7Y9_DSP/Tile_X0Y0_S2END[6]
+ Tile_X7Y9_DSP/Tile_X0Y0_S2END[7] Tile_X7Y9_DSP/Tile_X0Y0_S4END[0] Tile_X7Y9_DSP/Tile_X0Y0_S4END[10]
+ Tile_X7Y9_DSP/Tile_X0Y0_S4END[11] Tile_X7Y9_DSP/Tile_X0Y0_S4END[12] Tile_X7Y9_DSP/Tile_X0Y0_S4END[13]
+ Tile_X7Y9_DSP/Tile_X0Y0_S4END[14] Tile_X7Y9_DSP/Tile_X0Y0_S4END[15] Tile_X7Y9_DSP/Tile_X0Y0_S4END[1]
+ Tile_X7Y9_DSP/Tile_X0Y0_S4END[2] Tile_X7Y9_DSP/Tile_X0Y0_S4END[3] Tile_X7Y9_DSP/Tile_X0Y0_S4END[4]
+ Tile_X7Y9_DSP/Tile_X0Y0_S4END[5] Tile_X7Y9_DSP/Tile_X0Y0_S4END[6] Tile_X7Y9_DSP/Tile_X0Y0_S4END[7]
+ Tile_X7Y9_DSP/Tile_X0Y0_S4END[8] Tile_X7Y9_DSP/Tile_X0Y0_S4END[9] Tile_X7Y9_DSP/Tile_X0Y0_SS4END[0]
+ Tile_X7Y9_DSP/Tile_X0Y0_SS4END[10] Tile_X7Y9_DSP/Tile_X0Y0_SS4END[11] Tile_X7Y9_DSP/Tile_X0Y0_SS4END[12]
+ Tile_X7Y9_DSP/Tile_X0Y0_SS4END[13] Tile_X7Y9_DSP/Tile_X0Y0_SS4END[14] Tile_X7Y9_DSP/Tile_X0Y0_SS4END[15]
+ Tile_X7Y9_DSP/Tile_X0Y0_SS4END[1] Tile_X7Y9_DSP/Tile_X0Y0_SS4END[2] Tile_X7Y9_DSP/Tile_X0Y0_SS4END[3]
+ Tile_X7Y9_DSP/Tile_X0Y0_SS4END[4] Tile_X7Y9_DSP/Tile_X0Y0_SS4END[5] Tile_X7Y9_DSP/Tile_X0Y0_SS4END[6]
+ Tile_X7Y9_DSP/Tile_X0Y0_SS4END[7] Tile_X7Y9_DSP/Tile_X0Y0_SS4END[8] Tile_X7Y9_DSP/Tile_X0Y0_SS4END[9]
+ Tile_X7Y7_DSP/Tile_X0Y1_UserCLK Tile_X6Y8_LUT4AB/W1END[0] Tile_X6Y8_LUT4AB/W1END[1]
+ Tile_X6Y8_LUT4AB/W1END[2] Tile_X6Y8_LUT4AB/W1END[3] Tile_X8Y8_LUT4AB/W1BEG[0] Tile_X8Y8_LUT4AB/W1BEG[1]
+ Tile_X8Y8_LUT4AB/W1BEG[2] Tile_X8Y8_LUT4AB/W1BEG[3] Tile_X6Y8_LUT4AB/W2MID[0] Tile_X6Y8_LUT4AB/W2MID[1]
+ Tile_X6Y8_LUT4AB/W2MID[2] Tile_X6Y8_LUT4AB/W2MID[3] Tile_X6Y8_LUT4AB/W2MID[4] Tile_X6Y8_LUT4AB/W2MID[5]
+ Tile_X6Y8_LUT4AB/W2MID[6] Tile_X6Y8_LUT4AB/W2MID[7] Tile_X6Y8_LUT4AB/W2END[0] Tile_X6Y8_LUT4AB/W2END[1]
+ Tile_X6Y8_LUT4AB/W2END[2] Tile_X6Y8_LUT4AB/W2END[3] Tile_X6Y8_LUT4AB/W2END[4] Tile_X6Y8_LUT4AB/W2END[5]
+ Tile_X6Y8_LUT4AB/W2END[6] Tile_X6Y8_LUT4AB/W2END[7] Tile_X8Y8_LUT4AB/W2BEGb[0] Tile_X8Y8_LUT4AB/W2BEGb[1]
+ Tile_X8Y8_LUT4AB/W2BEGb[2] Tile_X8Y8_LUT4AB/W2BEGb[3] Tile_X8Y8_LUT4AB/W2BEGb[4]
+ Tile_X8Y8_LUT4AB/W2BEGb[5] Tile_X8Y8_LUT4AB/W2BEGb[6] Tile_X8Y8_LUT4AB/W2BEGb[7]
+ Tile_X8Y8_LUT4AB/W2BEG[0] Tile_X8Y8_LUT4AB/W2BEG[1] Tile_X8Y8_LUT4AB/W2BEG[2] Tile_X8Y8_LUT4AB/W2BEG[3]
+ Tile_X8Y8_LUT4AB/W2BEG[4] Tile_X8Y8_LUT4AB/W2BEG[5] Tile_X8Y8_LUT4AB/W2BEG[6] Tile_X8Y8_LUT4AB/W2BEG[7]
+ Tile_X6Y8_LUT4AB/W6END[0] Tile_X6Y8_LUT4AB/W6END[10] Tile_X6Y8_LUT4AB/W6END[11]
+ Tile_X6Y8_LUT4AB/W6END[1] Tile_X6Y8_LUT4AB/W6END[2] Tile_X6Y8_LUT4AB/W6END[3] Tile_X6Y8_LUT4AB/W6END[4]
+ Tile_X6Y8_LUT4AB/W6END[5] Tile_X6Y8_LUT4AB/W6END[6] Tile_X6Y8_LUT4AB/W6END[7] Tile_X6Y8_LUT4AB/W6END[8]
+ Tile_X6Y8_LUT4AB/W6END[9] Tile_X8Y8_LUT4AB/W6BEG[0] Tile_X8Y8_LUT4AB/W6BEG[10] Tile_X8Y8_LUT4AB/W6BEG[11]
+ Tile_X8Y8_LUT4AB/W6BEG[1] Tile_X8Y8_LUT4AB/W6BEG[2] Tile_X8Y8_LUT4AB/W6BEG[3] Tile_X8Y8_LUT4AB/W6BEG[4]
+ Tile_X8Y8_LUT4AB/W6BEG[5] Tile_X8Y8_LUT4AB/W6BEG[6] Tile_X8Y8_LUT4AB/W6BEG[7] Tile_X8Y8_LUT4AB/W6BEG[8]
+ Tile_X8Y8_LUT4AB/W6BEG[9] Tile_X6Y8_LUT4AB/WW4END[0] Tile_X6Y8_LUT4AB/WW4END[10]
+ Tile_X6Y8_LUT4AB/WW4END[11] Tile_X6Y8_LUT4AB/WW4END[12] Tile_X6Y8_LUT4AB/WW4END[13]
+ Tile_X6Y8_LUT4AB/WW4END[14] Tile_X6Y8_LUT4AB/WW4END[15] Tile_X6Y8_LUT4AB/WW4END[1]
+ Tile_X6Y8_LUT4AB/WW4END[2] Tile_X6Y8_LUT4AB/WW4END[3] Tile_X6Y8_LUT4AB/WW4END[4]
+ Tile_X6Y8_LUT4AB/WW4END[5] Tile_X6Y8_LUT4AB/WW4END[6] Tile_X6Y8_LUT4AB/WW4END[7]
+ Tile_X6Y8_LUT4AB/WW4END[8] Tile_X6Y8_LUT4AB/WW4END[9] Tile_X8Y8_LUT4AB/WW4BEG[0]
+ Tile_X8Y8_LUT4AB/WW4BEG[10] Tile_X8Y8_LUT4AB/WW4BEG[11] Tile_X8Y8_LUT4AB/WW4BEG[12]
+ Tile_X8Y8_LUT4AB/WW4BEG[13] Tile_X8Y8_LUT4AB/WW4BEG[14] Tile_X8Y8_LUT4AB/WW4BEG[15]
+ Tile_X8Y8_LUT4AB/WW4BEG[1] Tile_X8Y8_LUT4AB/WW4BEG[2] Tile_X8Y8_LUT4AB/WW4BEG[3]
+ Tile_X8Y8_LUT4AB/WW4BEG[4] Tile_X8Y8_LUT4AB/WW4BEG[5] Tile_X8Y8_LUT4AB/WW4BEG[6]
+ Tile_X8Y8_LUT4AB/WW4BEG[7] Tile_X8Y8_LUT4AB/WW4BEG[8] Tile_X8Y8_LUT4AB/WW4BEG[9]
+ VGND VPWR DSP
XTile_X4Y15_S_term_single2 Tile_X3Y15_S_CPU_IRQ/FrameData_O[0] Tile_X3Y15_S_CPU_IRQ/FrameData_O[10]
+ Tile_X3Y15_S_CPU_IRQ/FrameData_O[11] Tile_X3Y15_S_CPU_IRQ/FrameData_O[12] Tile_X3Y15_S_CPU_IRQ/FrameData_O[13]
+ Tile_X3Y15_S_CPU_IRQ/FrameData_O[14] Tile_X3Y15_S_CPU_IRQ/FrameData_O[15] Tile_X3Y15_S_CPU_IRQ/FrameData_O[16]
+ Tile_X3Y15_S_CPU_IRQ/FrameData_O[17] Tile_X3Y15_S_CPU_IRQ/FrameData_O[18] Tile_X3Y15_S_CPU_IRQ/FrameData_O[19]
+ Tile_X3Y15_S_CPU_IRQ/FrameData_O[1] Tile_X3Y15_S_CPU_IRQ/FrameData_O[20] Tile_X3Y15_S_CPU_IRQ/FrameData_O[21]
+ Tile_X3Y15_S_CPU_IRQ/FrameData_O[22] Tile_X3Y15_S_CPU_IRQ/FrameData_O[23] Tile_X3Y15_S_CPU_IRQ/FrameData_O[24]
+ Tile_X3Y15_S_CPU_IRQ/FrameData_O[25] Tile_X3Y15_S_CPU_IRQ/FrameData_O[26] Tile_X3Y15_S_CPU_IRQ/FrameData_O[27]
+ Tile_X3Y15_S_CPU_IRQ/FrameData_O[28] Tile_X3Y15_S_CPU_IRQ/FrameData_O[29] Tile_X3Y15_S_CPU_IRQ/FrameData_O[2]
+ Tile_X3Y15_S_CPU_IRQ/FrameData_O[30] Tile_X3Y15_S_CPU_IRQ/FrameData_O[31] Tile_X3Y15_S_CPU_IRQ/FrameData_O[3]
+ Tile_X3Y15_S_CPU_IRQ/FrameData_O[4] Tile_X3Y15_S_CPU_IRQ/FrameData_O[5] Tile_X3Y15_S_CPU_IRQ/FrameData_O[6]
+ Tile_X3Y15_S_CPU_IRQ/FrameData_O[7] Tile_X3Y15_S_CPU_IRQ/FrameData_O[8] Tile_X3Y15_S_CPU_IRQ/FrameData_O[9]
+ Tile_X5Y15_S_CPU_IF/FrameData[0] Tile_X5Y15_S_CPU_IF/FrameData[10] Tile_X5Y15_S_CPU_IF/FrameData[11]
+ Tile_X5Y15_S_CPU_IF/FrameData[12] Tile_X5Y15_S_CPU_IF/FrameData[13] Tile_X5Y15_S_CPU_IF/FrameData[14]
+ Tile_X5Y15_S_CPU_IF/FrameData[15] Tile_X5Y15_S_CPU_IF/FrameData[16] Tile_X5Y15_S_CPU_IF/FrameData[17]
+ Tile_X5Y15_S_CPU_IF/FrameData[18] Tile_X5Y15_S_CPU_IF/FrameData[19] Tile_X5Y15_S_CPU_IF/FrameData[1]
+ Tile_X5Y15_S_CPU_IF/FrameData[20] Tile_X5Y15_S_CPU_IF/FrameData[21] Tile_X5Y15_S_CPU_IF/FrameData[22]
+ Tile_X5Y15_S_CPU_IF/FrameData[23] Tile_X5Y15_S_CPU_IF/FrameData[24] Tile_X5Y15_S_CPU_IF/FrameData[25]
+ Tile_X5Y15_S_CPU_IF/FrameData[26] Tile_X5Y15_S_CPU_IF/FrameData[27] Tile_X5Y15_S_CPU_IF/FrameData[28]
+ Tile_X5Y15_S_CPU_IF/FrameData[29] Tile_X5Y15_S_CPU_IF/FrameData[2] Tile_X5Y15_S_CPU_IF/FrameData[30]
+ Tile_X5Y15_S_CPU_IF/FrameData[31] Tile_X5Y15_S_CPU_IF/FrameData[3] Tile_X5Y15_S_CPU_IF/FrameData[4]
+ Tile_X5Y15_S_CPU_IF/FrameData[5] Tile_X5Y15_S_CPU_IF/FrameData[6] Tile_X5Y15_S_CPU_IF/FrameData[7]
+ Tile_X5Y15_S_CPU_IF/FrameData[8] Tile_X5Y15_S_CPU_IF/FrameData[9] FrameStrobe[80]
+ FrameStrobe[90] FrameStrobe[91] FrameStrobe[92] FrameStrobe[93] FrameStrobe[94]
+ FrameStrobe[95] FrameStrobe[96] FrameStrobe[97] FrameStrobe[98] FrameStrobe[99]
+ FrameStrobe[81] FrameStrobe[82] FrameStrobe[83] FrameStrobe[84] FrameStrobe[85]
+ FrameStrobe[86] FrameStrobe[87] FrameStrobe[88] FrameStrobe[89] Tile_X4Y14_RegFile/FrameStrobe[0]
+ Tile_X4Y14_RegFile/FrameStrobe[10] Tile_X4Y14_RegFile/FrameStrobe[11] Tile_X4Y14_RegFile/FrameStrobe[12]
+ Tile_X4Y14_RegFile/FrameStrobe[13] Tile_X4Y14_RegFile/FrameStrobe[14] Tile_X4Y14_RegFile/FrameStrobe[15]
+ Tile_X4Y14_RegFile/FrameStrobe[16] Tile_X4Y14_RegFile/FrameStrobe[17] Tile_X4Y14_RegFile/FrameStrobe[18]
+ Tile_X4Y14_RegFile/FrameStrobe[19] Tile_X4Y14_RegFile/FrameStrobe[1] Tile_X4Y14_RegFile/FrameStrobe[2]
+ Tile_X4Y14_RegFile/FrameStrobe[3] Tile_X4Y14_RegFile/FrameStrobe[4] Tile_X4Y14_RegFile/FrameStrobe[5]
+ Tile_X4Y14_RegFile/FrameStrobe[6] Tile_X4Y14_RegFile/FrameStrobe[7] Tile_X4Y14_RegFile/FrameStrobe[8]
+ Tile_X4Y14_RegFile/FrameStrobe[9] Tile_X4Y14_RegFile/N1END[0] Tile_X4Y14_RegFile/N1END[1]
+ Tile_X4Y14_RegFile/N1END[2] Tile_X4Y14_RegFile/N1END[3] Tile_X4Y14_RegFile/N2MID[0]
+ Tile_X4Y14_RegFile/N2MID[1] Tile_X4Y14_RegFile/N2MID[2] Tile_X4Y14_RegFile/N2MID[3]
+ Tile_X4Y14_RegFile/N2MID[4] Tile_X4Y14_RegFile/N2MID[5] Tile_X4Y14_RegFile/N2MID[6]
+ Tile_X4Y14_RegFile/N2MID[7] Tile_X4Y14_RegFile/N2END[0] Tile_X4Y14_RegFile/N2END[1]
+ Tile_X4Y14_RegFile/N2END[2] Tile_X4Y14_RegFile/N2END[3] Tile_X4Y14_RegFile/N2END[4]
+ Tile_X4Y14_RegFile/N2END[5] Tile_X4Y14_RegFile/N2END[6] Tile_X4Y14_RegFile/N2END[7]
+ Tile_X4Y14_RegFile/N4END[0] Tile_X4Y14_RegFile/N4END[10] Tile_X4Y14_RegFile/N4END[11]
+ Tile_X4Y14_RegFile/N4END[12] Tile_X4Y14_RegFile/N4END[13] Tile_X4Y14_RegFile/N4END[14]
+ Tile_X4Y14_RegFile/N4END[15] Tile_X4Y14_RegFile/N4END[1] Tile_X4Y14_RegFile/N4END[2]
+ Tile_X4Y14_RegFile/N4END[3] Tile_X4Y14_RegFile/N4END[4] Tile_X4Y14_RegFile/N4END[5]
+ Tile_X4Y14_RegFile/N4END[6] Tile_X4Y14_RegFile/N4END[7] Tile_X4Y14_RegFile/N4END[8]
+ Tile_X4Y14_RegFile/N4END[9] Tile_X4Y14_RegFile/NN4END[0] Tile_X4Y14_RegFile/NN4END[10]
+ Tile_X4Y14_RegFile/NN4END[11] Tile_X4Y14_RegFile/NN4END[12] Tile_X4Y14_RegFile/NN4END[13]
+ Tile_X4Y14_RegFile/NN4END[14] Tile_X4Y14_RegFile/NN4END[15] Tile_X4Y14_RegFile/NN4END[1]
+ Tile_X4Y14_RegFile/NN4END[2] Tile_X4Y14_RegFile/NN4END[3] Tile_X4Y14_RegFile/NN4END[4]
+ Tile_X4Y14_RegFile/NN4END[5] Tile_X4Y14_RegFile/NN4END[6] Tile_X4Y14_RegFile/NN4END[7]
+ Tile_X4Y14_RegFile/NN4END[8] Tile_X4Y14_RegFile/NN4END[9] Tile_X4Y14_RegFile/S1BEG[0]
+ Tile_X4Y14_RegFile/S1BEG[1] Tile_X4Y14_RegFile/S1BEG[2] Tile_X4Y14_RegFile/S1BEG[3]
+ Tile_X4Y14_RegFile/S2BEGb[0] Tile_X4Y14_RegFile/S2BEGb[1] Tile_X4Y14_RegFile/S2BEGb[2]
+ Tile_X4Y14_RegFile/S2BEGb[3] Tile_X4Y14_RegFile/S2BEGb[4] Tile_X4Y14_RegFile/S2BEGb[5]
+ Tile_X4Y14_RegFile/S2BEGb[6] Tile_X4Y14_RegFile/S2BEGb[7] Tile_X4Y14_RegFile/S2BEG[0]
+ Tile_X4Y14_RegFile/S2BEG[1] Tile_X4Y14_RegFile/S2BEG[2] Tile_X4Y14_RegFile/S2BEG[3]
+ Tile_X4Y14_RegFile/S2BEG[4] Tile_X4Y14_RegFile/S2BEG[5] Tile_X4Y14_RegFile/S2BEG[6]
+ Tile_X4Y14_RegFile/S2BEG[7] Tile_X4Y14_RegFile/S4BEG[0] Tile_X4Y14_RegFile/S4BEG[10]
+ Tile_X4Y14_RegFile/S4BEG[11] Tile_X4Y14_RegFile/S4BEG[12] Tile_X4Y14_RegFile/S4BEG[13]
+ Tile_X4Y14_RegFile/S4BEG[14] Tile_X4Y14_RegFile/S4BEG[15] Tile_X4Y14_RegFile/S4BEG[1]
+ Tile_X4Y14_RegFile/S4BEG[2] Tile_X4Y14_RegFile/S4BEG[3] Tile_X4Y14_RegFile/S4BEG[4]
+ Tile_X4Y14_RegFile/S4BEG[5] Tile_X4Y14_RegFile/S4BEG[6] Tile_X4Y14_RegFile/S4BEG[7]
+ Tile_X4Y14_RegFile/S4BEG[8] Tile_X4Y14_RegFile/S4BEG[9] Tile_X4Y14_RegFile/SS4BEG[0]
+ Tile_X4Y14_RegFile/SS4BEG[10] Tile_X4Y14_RegFile/SS4BEG[11] Tile_X4Y14_RegFile/SS4BEG[12]
+ Tile_X4Y14_RegFile/SS4BEG[13] Tile_X4Y14_RegFile/SS4BEG[14] Tile_X4Y14_RegFile/SS4BEG[15]
+ Tile_X4Y14_RegFile/SS4BEG[1] Tile_X4Y14_RegFile/SS4BEG[2] Tile_X4Y14_RegFile/SS4BEG[3]
+ Tile_X4Y14_RegFile/SS4BEG[4] Tile_X4Y14_RegFile/SS4BEG[5] Tile_X4Y14_RegFile/SS4BEG[6]
+ Tile_X4Y14_RegFile/SS4BEG[7] Tile_X4Y14_RegFile/SS4BEG[8] Tile_X4Y14_RegFile/SS4BEG[9]
+ UserCLK Tile_X4Y14_RegFile/UserCLK VGND VPWR S_term_single2
XTile_X9Y4_LUT4AB Tile_X9Y5_LUT4AB/Co Tile_X9Y4_LUT4AB/Co Tile_X9Y4_LUT4AB/E1BEG[0]
+ Tile_X9Y4_LUT4AB/E1BEG[1] Tile_X9Y4_LUT4AB/E1BEG[2] Tile_X9Y4_LUT4AB/E1BEG[3] Tile_X9Y4_LUT4AB/E1END[0]
+ Tile_X9Y4_LUT4AB/E1END[1] Tile_X9Y4_LUT4AB/E1END[2] Tile_X9Y4_LUT4AB/E1END[3] Tile_X9Y4_LUT4AB/E2BEG[0]
+ Tile_X9Y4_LUT4AB/E2BEG[1] Tile_X9Y4_LUT4AB/E2BEG[2] Tile_X9Y4_LUT4AB/E2BEG[3] Tile_X9Y4_LUT4AB/E2BEG[4]
+ Tile_X9Y4_LUT4AB/E2BEG[5] Tile_X9Y4_LUT4AB/E2BEG[6] Tile_X9Y4_LUT4AB/E2BEG[7] Tile_X9Y4_LUT4AB/E2BEGb[0]
+ Tile_X9Y4_LUT4AB/E2BEGb[1] Tile_X9Y4_LUT4AB/E2BEGb[2] Tile_X9Y4_LUT4AB/E2BEGb[3]
+ Tile_X9Y4_LUT4AB/E2BEGb[4] Tile_X9Y4_LUT4AB/E2BEGb[5] Tile_X9Y4_LUT4AB/E2BEGb[6]
+ Tile_X9Y4_LUT4AB/E2BEGb[7] Tile_X9Y4_LUT4AB/E2END[0] Tile_X9Y4_LUT4AB/E2END[1] Tile_X9Y4_LUT4AB/E2END[2]
+ Tile_X9Y4_LUT4AB/E2END[3] Tile_X9Y4_LUT4AB/E2END[4] Tile_X9Y4_LUT4AB/E2END[5] Tile_X9Y4_LUT4AB/E2END[6]
+ Tile_X9Y4_LUT4AB/E2END[7] Tile_X9Y4_LUT4AB/E2MID[0] Tile_X9Y4_LUT4AB/E2MID[1] Tile_X9Y4_LUT4AB/E2MID[2]
+ Tile_X9Y4_LUT4AB/E2MID[3] Tile_X9Y4_LUT4AB/E2MID[4] Tile_X9Y4_LUT4AB/E2MID[5] Tile_X9Y4_LUT4AB/E2MID[6]
+ Tile_X9Y4_LUT4AB/E2MID[7] Tile_X9Y4_LUT4AB/E6BEG[0] Tile_X9Y4_LUT4AB/E6BEG[10] Tile_X9Y4_LUT4AB/E6BEG[11]
+ Tile_X9Y4_LUT4AB/E6BEG[1] Tile_X9Y4_LUT4AB/E6BEG[2] Tile_X9Y4_LUT4AB/E6BEG[3] Tile_X9Y4_LUT4AB/E6BEG[4]
+ Tile_X9Y4_LUT4AB/E6BEG[5] Tile_X9Y4_LUT4AB/E6BEG[6] Tile_X9Y4_LUT4AB/E6BEG[7] Tile_X9Y4_LUT4AB/E6BEG[8]
+ Tile_X9Y4_LUT4AB/E6BEG[9] Tile_X9Y4_LUT4AB/E6END[0] Tile_X9Y4_LUT4AB/E6END[10] Tile_X9Y4_LUT4AB/E6END[11]
+ Tile_X9Y4_LUT4AB/E6END[1] Tile_X9Y4_LUT4AB/E6END[2] Tile_X9Y4_LUT4AB/E6END[3] Tile_X9Y4_LUT4AB/E6END[4]
+ Tile_X9Y4_LUT4AB/E6END[5] Tile_X9Y4_LUT4AB/E6END[6] Tile_X9Y4_LUT4AB/E6END[7] Tile_X9Y4_LUT4AB/E6END[8]
+ Tile_X9Y4_LUT4AB/E6END[9] Tile_X9Y4_LUT4AB/EE4BEG[0] Tile_X9Y4_LUT4AB/EE4BEG[10]
+ Tile_X9Y4_LUT4AB/EE4BEG[11] Tile_X9Y4_LUT4AB/EE4BEG[12] Tile_X9Y4_LUT4AB/EE4BEG[13]
+ Tile_X9Y4_LUT4AB/EE4BEG[14] Tile_X9Y4_LUT4AB/EE4BEG[15] Tile_X9Y4_LUT4AB/EE4BEG[1]
+ Tile_X9Y4_LUT4AB/EE4BEG[2] Tile_X9Y4_LUT4AB/EE4BEG[3] Tile_X9Y4_LUT4AB/EE4BEG[4]
+ Tile_X9Y4_LUT4AB/EE4BEG[5] Tile_X9Y4_LUT4AB/EE4BEG[6] Tile_X9Y4_LUT4AB/EE4BEG[7]
+ Tile_X9Y4_LUT4AB/EE4BEG[8] Tile_X9Y4_LUT4AB/EE4BEG[9] Tile_X9Y4_LUT4AB/EE4END[0]
+ Tile_X9Y4_LUT4AB/EE4END[10] Tile_X9Y4_LUT4AB/EE4END[11] Tile_X9Y4_LUT4AB/EE4END[12]
+ Tile_X9Y4_LUT4AB/EE4END[13] Tile_X9Y4_LUT4AB/EE4END[14] Tile_X9Y4_LUT4AB/EE4END[15]
+ Tile_X9Y4_LUT4AB/EE4END[1] Tile_X9Y4_LUT4AB/EE4END[2] Tile_X9Y4_LUT4AB/EE4END[3]
+ Tile_X9Y4_LUT4AB/EE4END[4] Tile_X9Y4_LUT4AB/EE4END[5] Tile_X9Y4_LUT4AB/EE4END[6]
+ Tile_X9Y4_LUT4AB/EE4END[7] Tile_X9Y4_LUT4AB/EE4END[8] Tile_X9Y4_LUT4AB/EE4END[9]
+ Tile_X9Y4_LUT4AB/FrameData[0] Tile_X9Y4_LUT4AB/FrameData[10] Tile_X9Y4_LUT4AB/FrameData[11]
+ Tile_X9Y4_LUT4AB/FrameData[12] Tile_X9Y4_LUT4AB/FrameData[13] Tile_X9Y4_LUT4AB/FrameData[14]
+ Tile_X9Y4_LUT4AB/FrameData[15] Tile_X9Y4_LUT4AB/FrameData[16] Tile_X9Y4_LUT4AB/FrameData[17]
+ Tile_X9Y4_LUT4AB/FrameData[18] Tile_X9Y4_LUT4AB/FrameData[19] Tile_X9Y4_LUT4AB/FrameData[1]
+ Tile_X9Y4_LUT4AB/FrameData[20] Tile_X9Y4_LUT4AB/FrameData[21] Tile_X9Y4_LUT4AB/FrameData[22]
+ Tile_X9Y4_LUT4AB/FrameData[23] Tile_X9Y4_LUT4AB/FrameData[24] Tile_X9Y4_LUT4AB/FrameData[25]
+ Tile_X9Y4_LUT4AB/FrameData[26] Tile_X9Y4_LUT4AB/FrameData[27] Tile_X9Y4_LUT4AB/FrameData[28]
+ Tile_X9Y4_LUT4AB/FrameData[29] Tile_X9Y4_LUT4AB/FrameData[2] Tile_X9Y4_LUT4AB/FrameData[30]
+ Tile_X9Y4_LUT4AB/FrameData[31] Tile_X9Y4_LUT4AB/FrameData[3] Tile_X9Y4_LUT4AB/FrameData[4]
+ Tile_X9Y4_LUT4AB/FrameData[5] Tile_X9Y4_LUT4AB/FrameData[6] Tile_X9Y4_LUT4AB/FrameData[7]
+ Tile_X9Y4_LUT4AB/FrameData[8] Tile_X9Y4_LUT4AB/FrameData[9] Tile_X9Y4_LUT4AB/FrameData_O[0]
+ Tile_X9Y4_LUT4AB/FrameData_O[10] Tile_X9Y4_LUT4AB/FrameData_O[11] Tile_X9Y4_LUT4AB/FrameData_O[12]
+ Tile_X9Y4_LUT4AB/FrameData_O[13] Tile_X9Y4_LUT4AB/FrameData_O[14] Tile_X9Y4_LUT4AB/FrameData_O[15]
+ Tile_X9Y4_LUT4AB/FrameData_O[16] Tile_X9Y4_LUT4AB/FrameData_O[17] Tile_X9Y4_LUT4AB/FrameData_O[18]
+ Tile_X9Y4_LUT4AB/FrameData_O[19] Tile_X9Y4_LUT4AB/FrameData_O[1] Tile_X9Y4_LUT4AB/FrameData_O[20]
+ Tile_X9Y4_LUT4AB/FrameData_O[21] Tile_X9Y4_LUT4AB/FrameData_O[22] Tile_X9Y4_LUT4AB/FrameData_O[23]
+ Tile_X9Y4_LUT4AB/FrameData_O[24] Tile_X9Y4_LUT4AB/FrameData_O[25] Tile_X9Y4_LUT4AB/FrameData_O[26]
+ Tile_X9Y4_LUT4AB/FrameData_O[27] Tile_X9Y4_LUT4AB/FrameData_O[28] Tile_X9Y4_LUT4AB/FrameData_O[29]
+ Tile_X9Y4_LUT4AB/FrameData_O[2] Tile_X9Y4_LUT4AB/FrameData_O[30] Tile_X9Y4_LUT4AB/FrameData_O[31]
+ Tile_X9Y4_LUT4AB/FrameData_O[3] Tile_X9Y4_LUT4AB/FrameData_O[4] Tile_X9Y4_LUT4AB/FrameData_O[5]
+ Tile_X9Y4_LUT4AB/FrameData_O[6] Tile_X9Y4_LUT4AB/FrameData_O[7] Tile_X9Y4_LUT4AB/FrameData_O[8]
+ Tile_X9Y4_LUT4AB/FrameData_O[9] Tile_X9Y4_LUT4AB/FrameStrobe[0] Tile_X9Y4_LUT4AB/FrameStrobe[10]
+ Tile_X9Y4_LUT4AB/FrameStrobe[11] Tile_X9Y4_LUT4AB/FrameStrobe[12] Tile_X9Y4_LUT4AB/FrameStrobe[13]
+ Tile_X9Y4_LUT4AB/FrameStrobe[14] Tile_X9Y4_LUT4AB/FrameStrobe[15] Tile_X9Y4_LUT4AB/FrameStrobe[16]
+ Tile_X9Y4_LUT4AB/FrameStrobe[17] Tile_X9Y4_LUT4AB/FrameStrobe[18] Tile_X9Y4_LUT4AB/FrameStrobe[19]
+ Tile_X9Y4_LUT4AB/FrameStrobe[1] Tile_X9Y4_LUT4AB/FrameStrobe[2] Tile_X9Y4_LUT4AB/FrameStrobe[3]
+ Tile_X9Y4_LUT4AB/FrameStrobe[4] Tile_X9Y4_LUT4AB/FrameStrobe[5] Tile_X9Y4_LUT4AB/FrameStrobe[6]
+ Tile_X9Y4_LUT4AB/FrameStrobe[7] Tile_X9Y4_LUT4AB/FrameStrobe[8] Tile_X9Y4_LUT4AB/FrameStrobe[9]
+ Tile_X9Y3_LUT4AB/FrameStrobe[0] Tile_X9Y3_LUT4AB/FrameStrobe[10] Tile_X9Y3_LUT4AB/FrameStrobe[11]
+ Tile_X9Y3_LUT4AB/FrameStrobe[12] Tile_X9Y3_LUT4AB/FrameStrobe[13] Tile_X9Y3_LUT4AB/FrameStrobe[14]
+ Tile_X9Y3_LUT4AB/FrameStrobe[15] Tile_X9Y3_LUT4AB/FrameStrobe[16] Tile_X9Y3_LUT4AB/FrameStrobe[17]
+ Tile_X9Y3_LUT4AB/FrameStrobe[18] Tile_X9Y3_LUT4AB/FrameStrobe[19] Tile_X9Y3_LUT4AB/FrameStrobe[1]
+ Tile_X9Y3_LUT4AB/FrameStrobe[2] Tile_X9Y3_LUT4AB/FrameStrobe[3] Tile_X9Y3_LUT4AB/FrameStrobe[4]
+ Tile_X9Y3_LUT4AB/FrameStrobe[5] Tile_X9Y3_LUT4AB/FrameStrobe[6] Tile_X9Y3_LUT4AB/FrameStrobe[7]
+ Tile_X9Y3_LUT4AB/FrameStrobe[8] Tile_X9Y3_LUT4AB/FrameStrobe[9] Tile_X9Y4_LUT4AB/N1BEG[0]
+ Tile_X9Y4_LUT4AB/N1BEG[1] Tile_X9Y4_LUT4AB/N1BEG[2] Tile_X9Y4_LUT4AB/N1BEG[3] Tile_X9Y5_LUT4AB/N1BEG[0]
+ Tile_X9Y5_LUT4AB/N1BEG[1] Tile_X9Y5_LUT4AB/N1BEG[2] Tile_X9Y5_LUT4AB/N1BEG[3] Tile_X9Y4_LUT4AB/N2BEG[0]
+ Tile_X9Y4_LUT4AB/N2BEG[1] Tile_X9Y4_LUT4AB/N2BEG[2] Tile_X9Y4_LUT4AB/N2BEG[3] Tile_X9Y4_LUT4AB/N2BEG[4]
+ Tile_X9Y4_LUT4AB/N2BEG[5] Tile_X9Y4_LUT4AB/N2BEG[6] Tile_X9Y4_LUT4AB/N2BEG[7] Tile_X9Y3_LUT4AB/N2END[0]
+ Tile_X9Y3_LUT4AB/N2END[1] Tile_X9Y3_LUT4AB/N2END[2] Tile_X9Y3_LUT4AB/N2END[3] Tile_X9Y3_LUT4AB/N2END[4]
+ Tile_X9Y3_LUT4AB/N2END[5] Tile_X9Y3_LUT4AB/N2END[6] Tile_X9Y3_LUT4AB/N2END[7] Tile_X9Y4_LUT4AB/N2END[0]
+ Tile_X9Y4_LUT4AB/N2END[1] Tile_X9Y4_LUT4AB/N2END[2] Tile_X9Y4_LUT4AB/N2END[3] Tile_X9Y4_LUT4AB/N2END[4]
+ Tile_X9Y4_LUT4AB/N2END[5] Tile_X9Y4_LUT4AB/N2END[6] Tile_X9Y4_LUT4AB/N2END[7] Tile_X9Y5_LUT4AB/N2BEG[0]
+ Tile_X9Y5_LUT4AB/N2BEG[1] Tile_X9Y5_LUT4AB/N2BEG[2] Tile_X9Y5_LUT4AB/N2BEG[3] Tile_X9Y5_LUT4AB/N2BEG[4]
+ Tile_X9Y5_LUT4AB/N2BEG[5] Tile_X9Y5_LUT4AB/N2BEG[6] Tile_X9Y5_LUT4AB/N2BEG[7] Tile_X9Y4_LUT4AB/N4BEG[0]
+ Tile_X9Y4_LUT4AB/N4BEG[10] Tile_X9Y4_LUT4AB/N4BEG[11] Tile_X9Y4_LUT4AB/N4BEG[12]
+ Tile_X9Y4_LUT4AB/N4BEG[13] Tile_X9Y4_LUT4AB/N4BEG[14] Tile_X9Y4_LUT4AB/N4BEG[15]
+ Tile_X9Y4_LUT4AB/N4BEG[1] Tile_X9Y4_LUT4AB/N4BEG[2] Tile_X9Y4_LUT4AB/N4BEG[3] Tile_X9Y4_LUT4AB/N4BEG[4]
+ Tile_X9Y4_LUT4AB/N4BEG[5] Tile_X9Y4_LUT4AB/N4BEG[6] Tile_X9Y4_LUT4AB/N4BEG[7] Tile_X9Y4_LUT4AB/N4BEG[8]
+ Tile_X9Y4_LUT4AB/N4BEG[9] Tile_X9Y5_LUT4AB/N4BEG[0] Tile_X9Y5_LUT4AB/N4BEG[10] Tile_X9Y5_LUT4AB/N4BEG[11]
+ Tile_X9Y5_LUT4AB/N4BEG[12] Tile_X9Y5_LUT4AB/N4BEG[13] Tile_X9Y5_LUT4AB/N4BEG[14]
+ Tile_X9Y5_LUT4AB/N4BEG[15] Tile_X9Y5_LUT4AB/N4BEG[1] Tile_X9Y5_LUT4AB/N4BEG[2] Tile_X9Y5_LUT4AB/N4BEG[3]
+ Tile_X9Y5_LUT4AB/N4BEG[4] Tile_X9Y5_LUT4AB/N4BEG[5] Tile_X9Y5_LUT4AB/N4BEG[6] Tile_X9Y5_LUT4AB/N4BEG[7]
+ Tile_X9Y5_LUT4AB/N4BEG[8] Tile_X9Y5_LUT4AB/N4BEG[9] Tile_X9Y4_LUT4AB/NN4BEG[0] Tile_X9Y4_LUT4AB/NN4BEG[10]
+ Tile_X9Y4_LUT4AB/NN4BEG[11] Tile_X9Y4_LUT4AB/NN4BEG[12] Tile_X9Y4_LUT4AB/NN4BEG[13]
+ Tile_X9Y4_LUT4AB/NN4BEG[14] Tile_X9Y4_LUT4AB/NN4BEG[15] Tile_X9Y4_LUT4AB/NN4BEG[1]
+ Tile_X9Y4_LUT4AB/NN4BEG[2] Tile_X9Y4_LUT4AB/NN4BEG[3] Tile_X9Y4_LUT4AB/NN4BEG[4]
+ Tile_X9Y4_LUT4AB/NN4BEG[5] Tile_X9Y4_LUT4AB/NN4BEG[6] Tile_X9Y4_LUT4AB/NN4BEG[7]
+ Tile_X9Y4_LUT4AB/NN4BEG[8] Tile_X9Y4_LUT4AB/NN4BEG[9] Tile_X9Y5_LUT4AB/NN4BEG[0]
+ Tile_X9Y5_LUT4AB/NN4BEG[10] Tile_X9Y5_LUT4AB/NN4BEG[11] Tile_X9Y5_LUT4AB/NN4BEG[12]
+ Tile_X9Y5_LUT4AB/NN4BEG[13] Tile_X9Y5_LUT4AB/NN4BEG[14] Tile_X9Y5_LUT4AB/NN4BEG[15]
+ Tile_X9Y5_LUT4AB/NN4BEG[1] Tile_X9Y5_LUT4AB/NN4BEG[2] Tile_X9Y5_LUT4AB/NN4BEG[3]
+ Tile_X9Y5_LUT4AB/NN4BEG[4] Tile_X9Y5_LUT4AB/NN4BEG[5] Tile_X9Y5_LUT4AB/NN4BEG[6]
+ Tile_X9Y5_LUT4AB/NN4BEG[7] Tile_X9Y5_LUT4AB/NN4BEG[8] Tile_X9Y5_LUT4AB/NN4BEG[9]
+ Tile_X9Y5_LUT4AB/S1END[0] Tile_X9Y5_LUT4AB/S1END[1] Tile_X9Y5_LUT4AB/S1END[2] Tile_X9Y5_LUT4AB/S1END[3]
+ Tile_X9Y4_LUT4AB/S1END[0] Tile_X9Y4_LUT4AB/S1END[1] Tile_X9Y4_LUT4AB/S1END[2] Tile_X9Y4_LUT4AB/S1END[3]
+ Tile_X9Y5_LUT4AB/S2MID[0] Tile_X9Y5_LUT4AB/S2MID[1] Tile_X9Y5_LUT4AB/S2MID[2] Tile_X9Y5_LUT4AB/S2MID[3]
+ Tile_X9Y5_LUT4AB/S2MID[4] Tile_X9Y5_LUT4AB/S2MID[5] Tile_X9Y5_LUT4AB/S2MID[6] Tile_X9Y5_LUT4AB/S2MID[7]
+ Tile_X9Y5_LUT4AB/S2END[0] Tile_X9Y5_LUT4AB/S2END[1] Tile_X9Y5_LUT4AB/S2END[2] Tile_X9Y5_LUT4AB/S2END[3]
+ Tile_X9Y5_LUT4AB/S2END[4] Tile_X9Y5_LUT4AB/S2END[5] Tile_X9Y5_LUT4AB/S2END[6] Tile_X9Y5_LUT4AB/S2END[7]
+ Tile_X9Y4_LUT4AB/S2END[0] Tile_X9Y4_LUT4AB/S2END[1] Tile_X9Y4_LUT4AB/S2END[2] Tile_X9Y4_LUT4AB/S2END[3]
+ Tile_X9Y4_LUT4AB/S2END[4] Tile_X9Y4_LUT4AB/S2END[5] Tile_X9Y4_LUT4AB/S2END[6] Tile_X9Y4_LUT4AB/S2END[7]
+ Tile_X9Y4_LUT4AB/S2MID[0] Tile_X9Y4_LUT4AB/S2MID[1] Tile_X9Y4_LUT4AB/S2MID[2] Tile_X9Y4_LUT4AB/S2MID[3]
+ Tile_X9Y4_LUT4AB/S2MID[4] Tile_X9Y4_LUT4AB/S2MID[5] Tile_X9Y4_LUT4AB/S2MID[6] Tile_X9Y4_LUT4AB/S2MID[7]
+ Tile_X9Y5_LUT4AB/S4END[0] Tile_X9Y5_LUT4AB/S4END[10] Tile_X9Y5_LUT4AB/S4END[11]
+ Tile_X9Y5_LUT4AB/S4END[12] Tile_X9Y5_LUT4AB/S4END[13] Tile_X9Y5_LUT4AB/S4END[14]
+ Tile_X9Y5_LUT4AB/S4END[15] Tile_X9Y5_LUT4AB/S4END[1] Tile_X9Y5_LUT4AB/S4END[2] Tile_X9Y5_LUT4AB/S4END[3]
+ Tile_X9Y5_LUT4AB/S4END[4] Tile_X9Y5_LUT4AB/S4END[5] Tile_X9Y5_LUT4AB/S4END[6] Tile_X9Y5_LUT4AB/S4END[7]
+ Tile_X9Y5_LUT4AB/S4END[8] Tile_X9Y5_LUT4AB/S4END[9] Tile_X9Y4_LUT4AB/S4END[0] Tile_X9Y4_LUT4AB/S4END[10]
+ Tile_X9Y4_LUT4AB/S4END[11] Tile_X9Y4_LUT4AB/S4END[12] Tile_X9Y4_LUT4AB/S4END[13]
+ Tile_X9Y4_LUT4AB/S4END[14] Tile_X9Y4_LUT4AB/S4END[15] Tile_X9Y4_LUT4AB/S4END[1]
+ Tile_X9Y4_LUT4AB/S4END[2] Tile_X9Y4_LUT4AB/S4END[3] Tile_X9Y4_LUT4AB/S4END[4] Tile_X9Y4_LUT4AB/S4END[5]
+ Tile_X9Y4_LUT4AB/S4END[6] Tile_X9Y4_LUT4AB/S4END[7] Tile_X9Y4_LUT4AB/S4END[8] Tile_X9Y4_LUT4AB/S4END[9]
+ Tile_X9Y5_LUT4AB/SS4END[0] Tile_X9Y5_LUT4AB/SS4END[10] Tile_X9Y5_LUT4AB/SS4END[11]
+ Tile_X9Y5_LUT4AB/SS4END[12] Tile_X9Y5_LUT4AB/SS4END[13] Tile_X9Y5_LUT4AB/SS4END[14]
+ Tile_X9Y5_LUT4AB/SS4END[15] Tile_X9Y5_LUT4AB/SS4END[1] Tile_X9Y5_LUT4AB/SS4END[2]
+ Tile_X9Y5_LUT4AB/SS4END[3] Tile_X9Y5_LUT4AB/SS4END[4] Tile_X9Y5_LUT4AB/SS4END[5]
+ Tile_X9Y5_LUT4AB/SS4END[6] Tile_X9Y5_LUT4AB/SS4END[7] Tile_X9Y5_LUT4AB/SS4END[8]
+ Tile_X9Y5_LUT4AB/SS4END[9] Tile_X9Y4_LUT4AB/SS4END[0] Tile_X9Y4_LUT4AB/SS4END[10]
+ Tile_X9Y4_LUT4AB/SS4END[11] Tile_X9Y4_LUT4AB/SS4END[12] Tile_X9Y4_LUT4AB/SS4END[13]
+ Tile_X9Y4_LUT4AB/SS4END[14] Tile_X9Y4_LUT4AB/SS4END[15] Tile_X9Y4_LUT4AB/SS4END[1]
+ Tile_X9Y4_LUT4AB/SS4END[2] Tile_X9Y4_LUT4AB/SS4END[3] Tile_X9Y4_LUT4AB/SS4END[4]
+ Tile_X9Y4_LUT4AB/SS4END[5] Tile_X9Y4_LUT4AB/SS4END[6] Tile_X9Y4_LUT4AB/SS4END[7]
+ Tile_X9Y4_LUT4AB/SS4END[8] Tile_X9Y4_LUT4AB/SS4END[9] Tile_X9Y4_LUT4AB/UserCLK Tile_X9Y3_LUT4AB/UserCLK
+ VGND VPWR Tile_X9Y4_LUT4AB/W1BEG[0] Tile_X9Y4_LUT4AB/W1BEG[1] Tile_X9Y4_LUT4AB/W1BEG[2]
+ Tile_X9Y4_LUT4AB/W1BEG[3] Tile_X9Y4_LUT4AB/W1END[0] Tile_X9Y4_LUT4AB/W1END[1] Tile_X9Y4_LUT4AB/W1END[2]
+ Tile_X9Y4_LUT4AB/W1END[3] Tile_X9Y4_LUT4AB/W2BEG[0] Tile_X9Y4_LUT4AB/W2BEG[1] Tile_X9Y4_LUT4AB/W2BEG[2]
+ Tile_X9Y4_LUT4AB/W2BEG[3] Tile_X9Y4_LUT4AB/W2BEG[4] Tile_X9Y4_LUT4AB/W2BEG[5] Tile_X9Y4_LUT4AB/W2BEG[6]
+ Tile_X9Y4_LUT4AB/W2BEG[7] Tile_X8Y4_LUT4AB/W2END[0] Tile_X8Y4_LUT4AB/W2END[1] Tile_X8Y4_LUT4AB/W2END[2]
+ Tile_X8Y4_LUT4AB/W2END[3] Tile_X8Y4_LUT4AB/W2END[4] Tile_X8Y4_LUT4AB/W2END[5] Tile_X8Y4_LUT4AB/W2END[6]
+ Tile_X8Y4_LUT4AB/W2END[7] Tile_X9Y4_LUT4AB/W2END[0] Tile_X9Y4_LUT4AB/W2END[1] Tile_X9Y4_LUT4AB/W2END[2]
+ Tile_X9Y4_LUT4AB/W2END[3] Tile_X9Y4_LUT4AB/W2END[4] Tile_X9Y4_LUT4AB/W2END[5] Tile_X9Y4_LUT4AB/W2END[6]
+ Tile_X9Y4_LUT4AB/W2END[7] Tile_X9Y4_LUT4AB/W2MID[0] Tile_X9Y4_LUT4AB/W2MID[1] Tile_X9Y4_LUT4AB/W2MID[2]
+ Tile_X9Y4_LUT4AB/W2MID[3] Tile_X9Y4_LUT4AB/W2MID[4] Tile_X9Y4_LUT4AB/W2MID[5] Tile_X9Y4_LUT4AB/W2MID[6]
+ Tile_X9Y4_LUT4AB/W2MID[7] Tile_X9Y4_LUT4AB/W6BEG[0] Tile_X9Y4_LUT4AB/W6BEG[10] Tile_X9Y4_LUT4AB/W6BEG[11]
+ Tile_X9Y4_LUT4AB/W6BEG[1] Tile_X9Y4_LUT4AB/W6BEG[2] Tile_X9Y4_LUT4AB/W6BEG[3] Tile_X9Y4_LUT4AB/W6BEG[4]
+ Tile_X9Y4_LUT4AB/W6BEG[5] Tile_X9Y4_LUT4AB/W6BEG[6] Tile_X9Y4_LUT4AB/W6BEG[7] Tile_X9Y4_LUT4AB/W6BEG[8]
+ Tile_X9Y4_LUT4AB/W6BEG[9] Tile_X9Y4_LUT4AB/W6END[0] Tile_X9Y4_LUT4AB/W6END[10] Tile_X9Y4_LUT4AB/W6END[11]
+ Tile_X9Y4_LUT4AB/W6END[1] Tile_X9Y4_LUT4AB/W6END[2] Tile_X9Y4_LUT4AB/W6END[3] Tile_X9Y4_LUT4AB/W6END[4]
+ Tile_X9Y4_LUT4AB/W6END[5] Tile_X9Y4_LUT4AB/W6END[6] Tile_X9Y4_LUT4AB/W6END[7] Tile_X9Y4_LUT4AB/W6END[8]
+ Tile_X9Y4_LUT4AB/W6END[9] Tile_X9Y4_LUT4AB/WW4BEG[0] Tile_X9Y4_LUT4AB/WW4BEG[10]
+ Tile_X9Y4_LUT4AB/WW4BEG[11] Tile_X9Y4_LUT4AB/WW4BEG[12] Tile_X9Y4_LUT4AB/WW4BEG[13]
+ Tile_X9Y4_LUT4AB/WW4BEG[14] Tile_X9Y4_LUT4AB/WW4BEG[15] Tile_X9Y4_LUT4AB/WW4BEG[1]
+ Tile_X9Y4_LUT4AB/WW4BEG[2] Tile_X9Y4_LUT4AB/WW4BEG[3] Tile_X9Y4_LUT4AB/WW4BEG[4]
+ Tile_X9Y4_LUT4AB/WW4BEG[5] Tile_X9Y4_LUT4AB/WW4BEG[6] Tile_X9Y4_LUT4AB/WW4BEG[7]
+ Tile_X9Y4_LUT4AB/WW4BEG[8] Tile_X9Y4_LUT4AB/WW4BEG[9] Tile_X9Y4_LUT4AB/WW4END[0]
+ Tile_X9Y4_LUT4AB/WW4END[10] Tile_X9Y4_LUT4AB/WW4END[11] Tile_X9Y4_LUT4AB/WW4END[12]
+ Tile_X9Y4_LUT4AB/WW4END[13] Tile_X9Y4_LUT4AB/WW4END[14] Tile_X9Y4_LUT4AB/WW4END[15]
+ Tile_X9Y4_LUT4AB/WW4END[1] Tile_X9Y4_LUT4AB/WW4END[2] Tile_X9Y4_LUT4AB/WW4END[3]
+ Tile_X9Y4_LUT4AB/WW4END[4] Tile_X9Y4_LUT4AB/WW4END[5] Tile_X9Y4_LUT4AB/WW4END[6]
+ Tile_X9Y4_LUT4AB/WW4END[7] Tile_X9Y4_LUT4AB/WW4END[8] Tile_X9Y4_LUT4AB/WW4END[9]
+ LUT4AB
XTile_X2Y11_LUT4AB Tile_X2Y12_LUT4AB/Co Tile_X2Y11_LUT4AB/Co Tile_X3Y11_LUT4AB/E1END[0]
+ Tile_X3Y11_LUT4AB/E1END[1] Tile_X3Y11_LUT4AB/E1END[2] Tile_X3Y11_LUT4AB/E1END[3]
+ Tile_X2Y11_LUT4AB/E1END[0] Tile_X2Y11_LUT4AB/E1END[1] Tile_X2Y11_LUT4AB/E1END[2]
+ Tile_X2Y11_LUT4AB/E1END[3] Tile_X3Y11_LUT4AB/E2MID[0] Tile_X3Y11_LUT4AB/E2MID[1]
+ Tile_X3Y11_LUT4AB/E2MID[2] Tile_X3Y11_LUT4AB/E2MID[3] Tile_X3Y11_LUT4AB/E2MID[4]
+ Tile_X3Y11_LUT4AB/E2MID[5] Tile_X3Y11_LUT4AB/E2MID[6] Tile_X3Y11_LUT4AB/E2MID[7]
+ Tile_X3Y11_LUT4AB/E2END[0] Tile_X3Y11_LUT4AB/E2END[1] Tile_X3Y11_LUT4AB/E2END[2]
+ Tile_X3Y11_LUT4AB/E2END[3] Tile_X3Y11_LUT4AB/E2END[4] Tile_X3Y11_LUT4AB/E2END[5]
+ Tile_X3Y11_LUT4AB/E2END[6] Tile_X3Y11_LUT4AB/E2END[7] Tile_X2Y11_LUT4AB/E2END[0]
+ Tile_X2Y11_LUT4AB/E2END[1] Tile_X2Y11_LUT4AB/E2END[2] Tile_X2Y11_LUT4AB/E2END[3]
+ Tile_X2Y11_LUT4AB/E2END[4] Tile_X2Y11_LUT4AB/E2END[5] Tile_X2Y11_LUT4AB/E2END[6]
+ Tile_X2Y11_LUT4AB/E2END[7] Tile_X2Y11_LUT4AB/E2MID[0] Tile_X2Y11_LUT4AB/E2MID[1]
+ Tile_X2Y11_LUT4AB/E2MID[2] Tile_X2Y11_LUT4AB/E2MID[3] Tile_X2Y11_LUT4AB/E2MID[4]
+ Tile_X2Y11_LUT4AB/E2MID[5] Tile_X2Y11_LUT4AB/E2MID[6] Tile_X2Y11_LUT4AB/E2MID[7]
+ Tile_X3Y11_LUT4AB/E6END[0] Tile_X3Y11_LUT4AB/E6END[10] Tile_X3Y11_LUT4AB/E6END[11]
+ Tile_X3Y11_LUT4AB/E6END[1] Tile_X3Y11_LUT4AB/E6END[2] Tile_X3Y11_LUT4AB/E6END[3]
+ Tile_X3Y11_LUT4AB/E6END[4] Tile_X3Y11_LUT4AB/E6END[5] Tile_X3Y11_LUT4AB/E6END[6]
+ Tile_X3Y11_LUT4AB/E6END[7] Tile_X3Y11_LUT4AB/E6END[8] Tile_X3Y11_LUT4AB/E6END[9]
+ Tile_X2Y11_LUT4AB/E6END[0] Tile_X2Y11_LUT4AB/E6END[10] Tile_X2Y11_LUT4AB/E6END[11]
+ Tile_X2Y11_LUT4AB/E6END[1] Tile_X2Y11_LUT4AB/E6END[2] Tile_X2Y11_LUT4AB/E6END[3]
+ Tile_X2Y11_LUT4AB/E6END[4] Tile_X2Y11_LUT4AB/E6END[5] Tile_X2Y11_LUT4AB/E6END[6]
+ Tile_X2Y11_LUT4AB/E6END[7] Tile_X2Y11_LUT4AB/E6END[8] Tile_X2Y11_LUT4AB/E6END[9]
+ Tile_X3Y11_LUT4AB/EE4END[0] Tile_X3Y11_LUT4AB/EE4END[10] Tile_X3Y11_LUT4AB/EE4END[11]
+ Tile_X3Y11_LUT4AB/EE4END[12] Tile_X3Y11_LUT4AB/EE4END[13] Tile_X3Y11_LUT4AB/EE4END[14]
+ Tile_X3Y11_LUT4AB/EE4END[15] Tile_X3Y11_LUT4AB/EE4END[1] Tile_X3Y11_LUT4AB/EE4END[2]
+ Tile_X3Y11_LUT4AB/EE4END[3] Tile_X3Y11_LUT4AB/EE4END[4] Tile_X3Y11_LUT4AB/EE4END[5]
+ Tile_X3Y11_LUT4AB/EE4END[6] Tile_X3Y11_LUT4AB/EE4END[7] Tile_X3Y11_LUT4AB/EE4END[8]
+ Tile_X3Y11_LUT4AB/EE4END[9] Tile_X2Y11_LUT4AB/EE4END[0] Tile_X2Y11_LUT4AB/EE4END[10]
+ Tile_X2Y11_LUT4AB/EE4END[11] Tile_X2Y11_LUT4AB/EE4END[12] Tile_X2Y11_LUT4AB/EE4END[13]
+ Tile_X2Y11_LUT4AB/EE4END[14] Tile_X2Y11_LUT4AB/EE4END[15] Tile_X2Y11_LUT4AB/EE4END[1]
+ Tile_X2Y11_LUT4AB/EE4END[2] Tile_X2Y11_LUT4AB/EE4END[3] Tile_X2Y11_LUT4AB/EE4END[4]
+ Tile_X2Y11_LUT4AB/EE4END[5] Tile_X2Y11_LUT4AB/EE4END[6] Tile_X2Y11_LUT4AB/EE4END[7]
+ Tile_X2Y11_LUT4AB/EE4END[8] Tile_X2Y11_LUT4AB/EE4END[9] Tile_X2Y11_LUT4AB/FrameData[0]
+ Tile_X2Y11_LUT4AB/FrameData[10] Tile_X2Y11_LUT4AB/FrameData[11] Tile_X2Y11_LUT4AB/FrameData[12]
+ Tile_X2Y11_LUT4AB/FrameData[13] Tile_X2Y11_LUT4AB/FrameData[14] Tile_X2Y11_LUT4AB/FrameData[15]
+ Tile_X2Y11_LUT4AB/FrameData[16] Tile_X2Y11_LUT4AB/FrameData[17] Tile_X2Y11_LUT4AB/FrameData[18]
+ Tile_X2Y11_LUT4AB/FrameData[19] Tile_X2Y11_LUT4AB/FrameData[1] Tile_X2Y11_LUT4AB/FrameData[20]
+ Tile_X2Y11_LUT4AB/FrameData[21] Tile_X2Y11_LUT4AB/FrameData[22] Tile_X2Y11_LUT4AB/FrameData[23]
+ Tile_X2Y11_LUT4AB/FrameData[24] Tile_X2Y11_LUT4AB/FrameData[25] Tile_X2Y11_LUT4AB/FrameData[26]
+ Tile_X2Y11_LUT4AB/FrameData[27] Tile_X2Y11_LUT4AB/FrameData[28] Tile_X2Y11_LUT4AB/FrameData[29]
+ Tile_X2Y11_LUT4AB/FrameData[2] Tile_X2Y11_LUT4AB/FrameData[30] Tile_X2Y11_LUT4AB/FrameData[31]
+ Tile_X2Y11_LUT4AB/FrameData[3] Tile_X2Y11_LUT4AB/FrameData[4] Tile_X2Y11_LUT4AB/FrameData[5]
+ Tile_X2Y11_LUT4AB/FrameData[6] Tile_X2Y11_LUT4AB/FrameData[7] Tile_X2Y11_LUT4AB/FrameData[8]
+ Tile_X2Y11_LUT4AB/FrameData[9] Tile_X3Y11_LUT4AB/FrameData[0] Tile_X3Y11_LUT4AB/FrameData[10]
+ Tile_X3Y11_LUT4AB/FrameData[11] Tile_X3Y11_LUT4AB/FrameData[12] Tile_X3Y11_LUT4AB/FrameData[13]
+ Tile_X3Y11_LUT4AB/FrameData[14] Tile_X3Y11_LUT4AB/FrameData[15] Tile_X3Y11_LUT4AB/FrameData[16]
+ Tile_X3Y11_LUT4AB/FrameData[17] Tile_X3Y11_LUT4AB/FrameData[18] Tile_X3Y11_LUT4AB/FrameData[19]
+ Tile_X3Y11_LUT4AB/FrameData[1] Tile_X3Y11_LUT4AB/FrameData[20] Tile_X3Y11_LUT4AB/FrameData[21]
+ Tile_X3Y11_LUT4AB/FrameData[22] Tile_X3Y11_LUT4AB/FrameData[23] Tile_X3Y11_LUT4AB/FrameData[24]
+ Tile_X3Y11_LUT4AB/FrameData[25] Tile_X3Y11_LUT4AB/FrameData[26] Tile_X3Y11_LUT4AB/FrameData[27]
+ Tile_X3Y11_LUT4AB/FrameData[28] Tile_X3Y11_LUT4AB/FrameData[29] Tile_X3Y11_LUT4AB/FrameData[2]
+ Tile_X3Y11_LUT4AB/FrameData[30] Tile_X3Y11_LUT4AB/FrameData[31] Tile_X3Y11_LUT4AB/FrameData[3]
+ Tile_X3Y11_LUT4AB/FrameData[4] Tile_X3Y11_LUT4AB/FrameData[5] Tile_X3Y11_LUT4AB/FrameData[6]
+ Tile_X3Y11_LUT4AB/FrameData[7] Tile_X3Y11_LUT4AB/FrameData[8] Tile_X3Y11_LUT4AB/FrameData[9]
+ Tile_X2Y11_LUT4AB/FrameStrobe[0] Tile_X2Y11_LUT4AB/FrameStrobe[10] Tile_X2Y11_LUT4AB/FrameStrobe[11]
+ Tile_X2Y11_LUT4AB/FrameStrobe[12] Tile_X2Y11_LUT4AB/FrameStrobe[13] Tile_X2Y11_LUT4AB/FrameStrobe[14]
+ Tile_X2Y11_LUT4AB/FrameStrobe[15] Tile_X2Y11_LUT4AB/FrameStrobe[16] Tile_X2Y11_LUT4AB/FrameStrobe[17]
+ Tile_X2Y11_LUT4AB/FrameStrobe[18] Tile_X2Y11_LUT4AB/FrameStrobe[19] Tile_X2Y11_LUT4AB/FrameStrobe[1]
+ Tile_X2Y11_LUT4AB/FrameStrobe[2] Tile_X2Y11_LUT4AB/FrameStrobe[3] Tile_X2Y11_LUT4AB/FrameStrobe[4]
+ Tile_X2Y11_LUT4AB/FrameStrobe[5] Tile_X2Y11_LUT4AB/FrameStrobe[6] Tile_X2Y11_LUT4AB/FrameStrobe[7]
+ Tile_X2Y11_LUT4AB/FrameStrobe[8] Tile_X2Y11_LUT4AB/FrameStrobe[9] Tile_X2Y10_LUT4AB/FrameStrobe[0]
+ Tile_X2Y10_LUT4AB/FrameStrobe[10] Tile_X2Y10_LUT4AB/FrameStrobe[11] Tile_X2Y10_LUT4AB/FrameStrobe[12]
+ Tile_X2Y10_LUT4AB/FrameStrobe[13] Tile_X2Y10_LUT4AB/FrameStrobe[14] Tile_X2Y10_LUT4AB/FrameStrobe[15]
+ Tile_X2Y10_LUT4AB/FrameStrobe[16] Tile_X2Y10_LUT4AB/FrameStrobe[17] Tile_X2Y10_LUT4AB/FrameStrobe[18]
+ Tile_X2Y10_LUT4AB/FrameStrobe[19] Tile_X2Y10_LUT4AB/FrameStrobe[1] Tile_X2Y10_LUT4AB/FrameStrobe[2]
+ Tile_X2Y10_LUT4AB/FrameStrobe[3] Tile_X2Y10_LUT4AB/FrameStrobe[4] Tile_X2Y10_LUT4AB/FrameStrobe[5]
+ Tile_X2Y10_LUT4AB/FrameStrobe[6] Tile_X2Y10_LUT4AB/FrameStrobe[7] Tile_X2Y10_LUT4AB/FrameStrobe[8]
+ Tile_X2Y10_LUT4AB/FrameStrobe[9] Tile_X2Y11_LUT4AB/N1BEG[0] Tile_X2Y11_LUT4AB/N1BEG[1]
+ Tile_X2Y11_LUT4AB/N1BEG[2] Tile_X2Y11_LUT4AB/N1BEG[3] Tile_X2Y12_LUT4AB/N1BEG[0]
+ Tile_X2Y12_LUT4AB/N1BEG[1] Tile_X2Y12_LUT4AB/N1BEG[2] Tile_X2Y12_LUT4AB/N1BEG[3]
+ Tile_X2Y11_LUT4AB/N2BEG[0] Tile_X2Y11_LUT4AB/N2BEG[1] Tile_X2Y11_LUT4AB/N2BEG[2]
+ Tile_X2Y11_LUT4AB/N2BEG[3] Tile_X2Y11_LUT4AB/N2BEG[4] Tile_X2Y11_LUT4AB/N2BEG[5]
+ Tile_X2Y11_LUT4AB/N2BEG[6] Tile_X2Y11_LUT4AB/N2BEG[7] Tile_X2Y10_LUT4AB/N2END[0]
+ Tile_X2Y10_LUT4AB/N2END[1] Tile_X2Y10_LUT4AB/N2END[2] Tile_X2Y10_LUT4AB/N2END[3]
+ Tile_X2Y10_LUT4AB/N2END[4] Tile_X2Y10_LUT4AB/N2END[5] Tile_X2Y10_LUT4AB/N2END[6]
+ Tile_X2Y10_LUT4AB/N2END[7] Tile_X2Y11_LUT4AB/N2END[0] Tile_X2Y11_LUT4AB/N2END[1]
+ Tile_X2Y11_LUT4AB/N2END[2] Tile_X2Y11_LUT4AB/N2END[3] Tile_X2Y11_LUT4AB/N2END[4]
+ Tile_X2Y11_LUT4AB/N2END[5] Tile_X2Y11_LUT4AB/N2END[6] Tile_X2Y11_LUT4AB/N2END[7]
+ Tile_X2Y12_LUT4AB/N2BEG[0] Tile_X2Y12_LUT4AB/N2BEG[1] Tile_X2Y12_LUT4AB/N2BEG[2]
+ Tile_X2Y12_LUT4AB/N2BEG[3] Tile_X2Y12_LUT4AB/N2BEG[4] Tile_X2Y12_LUT4AB/N2BEG[5]
+ Tile_X2Y12_LUT4AB/N2BEG[6] Tile_X2Y12_LUT4AB/N2BEG[7] Tile_X2Y11_LUT4AB/N4BEG[0]
+ Tile_X2Y11_LUT4AB/N4BEG[10] Tile_X2Y11_LUT4AB/N4BEG[11] Tile_X2Y11_LUT4AB/N4BEG[12]
+ Tile_X2Y11_LUT4AB/N4BEG[13] Tile_X2Y11_LUT4AB/N4BEG[14] Tile_X2Y11_LUT4AB/N4BEG[15]
+ Tile_X2Y11_LUT4AB/N4BEG[1] Tile_X2Y11_LUT4AB/N4BEG[2] Tile_X2Y11_LUT4AB/N4BEG[3]
+ Tile_X2Y11_LUT4AB/N4BEG[4] Tile_X2Y11_LUT4AB/N4BEG[5] Tile_X2Y11_LUT4AB/N4BEG[6]
+ Tile_X2Y11_LUT4AB/N4BEG[7] Tile_X2Y11_LUT4AB/N4BEG[8] Tile_X2Y11_LUT4AB/N4BEG[9]
+ Tile_X2Y12_LUT4AB/N4BEG[0] Tile_X2Y12_LUT4AB/N4BEG[10] Tile_X2Y12_LUT4AB/N4BEG[11]
+ Tile_X2Y12_LUT4AB/N4BEG[12] Tile_X2Y12_LUT4AB/N4BEG[13] Tile_X2Y12_LUT4AB/N4BEG[14]
+ Tile_X2Y12_LUT4AB/N4BEG[15] Tile_X2Y12_LUT4AB/N4BEG[1] Tile_X2Y12_LUT4AB/N4BEG[2]
+ Tile_X2Y12_LUT4AB/N4BEG[3] Tile_X2Y12_LUT4AB/N4BEG[4] Tile_X2Y12_LUT4AB/N4BEG[5]
+ Tile_X2Y12_LUT4AB/N4BEG[6] Tile_X2Y12_LUT4AB/N4BEG[7] Tile_X2Y12_LUT4AB/N4BEG[8]
+ Tile_X2Y12_LUT4AB/N4BEG[9] Tile_X2Y11_LUT4AB/NN4BEG[0] Tile_X2Y11_LUT4AB/NN4BEG[10]
+ Tile_X2Y11_LUT4AB/NN4BEG[11] Tile_X2Y11_LUT4AB/NN4BEG[12] Tile_X2Y11_LUT4AB/NN4BEG[13]
+ Tile_X2Y11_LUT4AB/NN4BEG[14] Tile_X2Y11_LUT4AB/NN4BEG[15] Tile_X2Y11_LUT4AB/NN4BEG[1]
+ Tile_X2Y11_LUT4AB/NN4BEG[2] Tile_X2Y11_LUT4AB/NN4BEG[3] Tile_X2Y11_LUT4AB/NN4BEG[4]
+ Tile_X2Y11_LUT4AB/NN4BEG[5] Tile_X2Y11_LUT4AB/NN4BEG[6] Tile_X2Y11_LUT4AB/NN4BEG[7]
+ Tile_X2Y11_LUT4AB/NN4BEG[8] Tile_X2Y11_LUT4AB/NN4BEG[9] Tile_X2Y12_LUT4AB/NN4BEG[0]
+ Tile_X2Y12_LUT4AB/NN4BEG[10] Tile_X2Y12_LUT4AB/NN4BEG[11] Tile_X2Y12_LUT4AB/NN4BEG[12]
+ Tile_X2Y12_LUT4AB/NN4BEG[13] Tile_X2Y12_LUT4AB/NN4BEG[14] Tile_X2Y12_LUT4AB/NN4BEG[15]
+ Tile_X2Y12_LUT4AB/NN4BEG[1] Tile_X2Y12_LUT4AB/NN4BEG[2] Tile_X2Y12_LUT4AB/NN4BEG[3]
+ Tile_X2Y12_LUT4AB/NN4BEG[4] Tile_X2Y12_LUT4AB/NN4BEG[5] Tile_X2Y12_LUT4AB/NN4BEG[6]
+ Tile_X2Y12_LUT4AB/NN4BEG[7] Tile_X2Y12_LUT4AB/NN4BEG[8] Tile_X2Y12_LUT4AB/NN4BEG[9]
+ Tile_X2Y12_LUT4AB/S1END[0] Tile_X2Y12_LUT4AB/S1END[1] Tile_X2Y12_LUT4AB/S1END[2]
+ Tile_X2Y12_LUT4AB/S1END[3] Tile_X2Y11_LUT4AB/S1END[0] Tile_X2Y11_LUT4AB/S1END[1]
+ Tile_X2Y11_LUT4AB/S1END[2] Tile_X2Y11_LUT4AB/S1END[3] Tile_X2Y12_LUT4AB/S2MID[0]
+ Tile_X2Y12_LUT4AB/S2MID[1] Tile_X2Y12_LUT4AB/S2MID[2] Tile_X2Y12_LUT4AB/S2MID[3]
+ Tile_X2Y12_LUT4AB/S2MID[4] Tile_X2Y12_LUT4AB/S2MID[5] Tile_X2Y12_LUT4AB/S2MID[6]
+ Tile_X2Y12_LUT4AB/S2MID[7] Tile_X2Y12_LUT4AB/S2END[0] Tile_X2Y12_LUT4AB/S2END[1]
+ Tile_X2Y12_LUT4AB/S2END[2] Tile_X2Y12_LUT4AB/S2END[3] Tile_X2Y12_LUT4AB/S2END[4]
+ Tile_X2Y12_LUT4AB/S2END[5] Tile_X2Y12_LUT4AB/S2END[6] Tile_X2Y12_LUT4AB/S2END[7]
+ Tile_X2Y11_LUT4AB/S2END[0] Tile_X2Y11_LUT4AB/S2END[1] Tile_X2Y11_LUT4AB/S2END[2]
+ Tile_X2Y11_LUT4AB/S2END[3] Tile_X2Y11_LUT4AB/S2END[4] Tile_X2Y11_LUT4AB/S2END[5]
+ Tile_X2Y11_LUT4AB/S2END[6] Tile_X2Y11_LUT4AB/S2END[7] Tile_X2Y11_LUT4AB/S2MID[0]
+ Tile_X2Y11_LUT4AB/S2MID[1] Tile_X2Y11_LUT4AB/S2MID[2] Tile_X2Y11_LUT4AB/S2MID[3]
+ Tile_X2Y11_LUT4AB/S2MID[4] Tile_X2Y11_LUT4AB/S2MID[5] Tile_X2Y11_LUT4AB/S2MID[6]
+ Tile_X2Y11_LUT4AB/S2MID[7] Tile_X2Y12_LUT4AB/S4END[0] Tile_X2Y12_LUT4AB/S4END[10]
+ Tile_X2Y12_LUT4AB/S4END[11] Tile_X2Y12_LUT4AB/S4END[12] Tile_X2Y12_LUT4AB/S4END[13]
+ Tile_X2Y12_LUT4AB/S4END[14] Tile_X2Y12_LUT4AB/S4END[15] Tile_X2Y12_LUT4AB/S4END[1]
+ Tile_X2Y12_LUT4AB/S4END[2] Tile_X2Y12_LUT4AB/S4END[3] Tile_X2Y12_LUT4AB/S4END[4]
+ Tile_X2Y12_LUT4AB/S4END[5] Tile_X2Y12_LUT4AB/S4END[6] Tile_X2Y12_LUT4AB/S4END[7]
+ Tile_X2Y12_LUT4AB/S4END[8] Tile_X2Y12_LUT4AB/S4END[9] Tile_X2Y11_LUT4AB/S4END[0]
+ Tile_X2Y11_LUT4AB/S4END[10] Tile_X2Y11_LUT4AB/S4END[11] Tile_X2Y11_LUT4AB/S4END[12]
+ Tile_X2Y11_LUT4AB/S4END[13] Tile_X2Y11_LUT4AB/S4END[14] Tile_X2Y11_LUT4AB/S4END[15]
+ Tile_X2Y11_LUT4AB/S4END[1] Tile_X2Y11_LUT4AB/S4END[2] Tile_X2Y11_LUT4AB/S4END[3]
+ Tile_X2Y11_LUT4AB/S4END[4] Tile_X2Y11_LUT4AB/S4END[5] Tile_X2Y11_LUT4AB/S4END[6]
+ Tile_X2Y11_LUT4AB/S4END[7] Tile_X2Y11_LUT4AB/S4END[8] Tile_X2Y11_LUT4AB/S4END[9]
+ Tile_X2Y12_LUT4AB/SS4END[0] Tile_X2Y12_LUT4AB/SS4END[10] Tile_X2Y12_LUT4AB/SS4END[11]
+ Tile_X2Y12_LUT4AB/SS4END[12] Tile_X2Y12_LUT4AB/SS4END[13] Tile_X2Y12_LUT4AB/SS4END[14]
+ Tile_X2Y12_LUT4AB/SS4END[15] Tile_X2Y12_LUT4AB/SS4END[1] Tile_X2Y12_LUT4AB/SS4END[2]
+ Tile_X2Y12_LUT4AB/SS4END[3] Tile_X2Y12_LUT4AB/SS4END[4] Tile_X2Y12_LUT4AB/SS4END[5]
+ Tile_X2Y12_LUT4AB/SS4END[6] Tile_X2Y12_LUT4AB/SS4END[7] Tile_X2Y12_LUT4AB/SS4END[8]
+ Tile_X2Y12_LUT4AB/SS4END[9] Tile_X2Y11_LUT4AB/SS4END[0] Tile_X2Y11_LUT4AB/SS4END[10]
+ Tile_X2Y11_LUT4AB/SS4END[11] Tile_X2Y11_LUT4AB/SS4END[12] Tile_X2Y11_LUT4AB/SS4END[13]
+ Tile_X2Y11_LUT4AB/SS4END[14] Tile_X2Y11_LUT4AB/SS4END[15] Tile_X2Y11_LUT4AB/SS4END[1]
+ Tile_X2Y11_LUT4AB/SS4END[2] Tile_X2Y11_LUT4AB/SS4END[3] Tile_X2Y11_LUT4AB/SS4END[4]
+ Tile_X2Y11_LUT4AB/SS4END[5] Tile_X2Y11_LUT4AB/SS4END[6] Tile_X2Y11_LUT4AB/SS4END[7]
+ Tile_X2Y11_LUT4AB/SS4END[8] Tile_X2Y11_LUT4AB/SS4END[9] Tile_X2Y11_LUT4AB/UserCLK
+ Tile_X2Y10_LUT4AB/UserCLK VGND VPWR Tile_X2Y11_LUT4AB/W1BEG[0] Tile_X2Y11_LUT4AB/W1BEG[1]
+ Tile_X2Y11_LUT4AB/W1BEG[2] Tile_X2Y11_LUT4AB/W1BEG[3] Tile_X3Y11_LUT4AB/W1BEG[0]
+ Tile_X3Y11_LUT4AB/W1BEG[1] Tile_X3Y11_LUT4AB/W1BEG[2] Tile_X3Y11_LUT4AB/W1BEG[3]
+ Tile_X2Y11_LUT4AB/W2BEG[0] Tile_X2Y11_LUT4AB/W2BEG[1] Tile_X2Y11_LUT4AB/W2BEG[2]
+ Tile_X2Y11_LUT4AB/W2BEG[3] Tile_X2Y11_LUT4AB/W2BEG[4] Tile_X2Y11_LUT4AB/W2BEG[5]
+ Tile_X2Y11_LUT4AB/W2BEG[6] Tile_X2Y11_LUT4AB/W2BEG[7] Tile_X1Y11_LUT4AB/W2END[0]
+ Tile_X1Y11_LUT4AB/W2END[1] Tile_X1Y11_LUT4AB/W2END[2] Tile_X1Y11_LUT4AB/W2END[3]
+ Tile_X1Y11_LUT4AB/W2END[4] Tile_X1Y11_LUT4AB/W2END[5] Tile_X1Y11_LUT4AB/W2END[6]
+ Tile_X1Y11_LUT4AB/W2END[7] Tile_X2Y11_LUT4AB/W2END[0] Tile_X2Y11_LUT4AB/W2END[1]
+ Tile_X2Y11_LUT4AB/W2END[2] Tile_X2Y11_LUT4AB/W2END[3] Tile_X2Y11_LUT4AB/W2END[4]
+ Tile_X2Y11_LUT4AB/W2END[5] Tile_X2Y11_LUT4AB/W2END[6] Tile_X2Y11_LUT4AB/W2END[7]
+ Tile_X3Y11_LUT4AB/W2BEG[0] Tile_X3Y11_LUT4AB/W2BEG[1] Tile_X3Y11_LUT4AB/W2BEG[2]
+ Tile_X3Y11_LUT4AB/W2BEG[3] Tile_X3Y11_LUT4AB/W2BEG[4] Tile_X3Y11_LUT4AB/W2BEG[5]
+ Tile_X3Y11_LUT4AB/W2BEG[6] Tile_X3Y11_LUT4AB/W2BEG[7] Tile_X2Y11_LUT4AB/W6BEG[0]
+ Tile_X2Y11_LUT4AB/W6BEG[10] Tile_X2Y11_LUT4AB/W6BEG[11] Tile_X2Y11_LUT4AB/W6BEG[1]
+ Tile_X2Y11_LUT4AB/W6BEG[2] Tile_X2Y11_LUT4AB/W6BEG[3] Tile_X2Y11_LUT4AB/W6BEG[4]
+ Tile_X2Y11_LUT4AB/W6BEG[5] Tile_X2Y11_LUT4AB/W6BEG[6] Tile_X2Y11_LUT4AB/W6BEG[7]
+ Tile_X2Y11_LUT4AB/W6BEG[8] Tile_X2Y11_LUT4AB/W6BEG[9] Tile_X3Y11_LUT4AB/W6BEG[0]
+ Tile_X3Y11_LUT4AB/W6BEG[10] Tile_X3Y11_LUT4AB/W6BEG[11] Tile_X3Y11_LUT4AB/W6BEG[1]
+ Tile_X3Y11_LUT4AB/W6BEG[2] Tile_X3Y11_LUT4AB/W6BEG[3] Tile_X3Y11_LUT4AB/W6BEG[4]
+ Tile_X3Y11_LUT4AB/W6BEG[5] Tile_X3Y11_LUT4AB/W6BEG[6] Tile_X3Y11_LUT4AB/W6BEG[7]
+ Tile_X3Y11_LUT4AB/W6BEG[8] Tile_X3Y11_LUT4AB/W6BEG[9] Tile_X2Y11_LUT4AB/WW4BEG[0]
+ Tile_X2Y11_LUT4AB/WW4BEG[10] Tile_X2Y11_LUT4AB/WW4BEG[11] Tile_X2Y11_LUT4AB/WW4BEG[12]
+ Tile_X2Y11_LUT4AB/WW4BEG[13] Tile_X2Y11_LUT4AB/WW4BEG[14] Tile_X2Y11_LUT4AB/WW4BEG[15]
+ Tile_X2Y11_LUT4AB/WW4BEG[1] Tile_X2Y11_LUT4AB/WW4BEG[2] Tile_X2Y11_LUT4AB/WW4BEG[3]
+ Tile_X2Y11_LUT4AB/WW4BEG[4] Tile_X2Y11_LUT4AB/WW4BEG[5] Tile_X2Y11_LUT4AB/WW4BEG[6]
+ Tile_X2Y11_LUT4AB/WW4BEG[7] Tile_X2Y11_LUT4AB/WW4BEG[8] Tile_X2Y11_LUT4AB/WW4BEG[9]
+ Tile_X3Y11_LUT4AB/WW4BEG[0] Tile_X3Y11_LUT4AB/WW4BEG[10] Tile_X3Y11_LUT4AB/WW4BEG[11]
+ Tile_X3Y11_LUT4AB/WW4BEG[12] Tile_X3Y11_LUT4AB/WW4BEG[13] Tile_X3Y11_LUT4AB/WW4BEG[14]
+ Tile_X3Y11_LUT4AB/WW4BEG[15] Tile_X3Y11_LUT4AB/WW4BEG[1] Tile_X3Y11_LUT4AB/WW4BEG[2]
+ Tile_X3Y11_LUT4AB/WW4BEG[3] Tile_X3Y11_LUT4AB/WW4BEG[4] Tile_X3Y11_LUT4AB/WW4BEG[5]
+ Tile_X3Y11_LUT4AB/WW4BEG[6] Tile_X3Y11_LUT4AB/WW4BEG[7] Tile_X3Y11_LUT4AB/WW4BEG[8]
+ Tile_X3Y11_LUT4AB/WW4BEG[9] LUT4AB
XTile_X3Y0_N_term_single Tile_X3Y1_LUT4AB/Co Tile_X2Y0_N_IO/FrameData_O[0] Tile_X2Y0_N_IO/FrameData_O[10]
+ Tile_X2Y0_N_IO/FrameData_O[11] Tile_X2Y0_N_IO/FrameData_O[12] Tile_X2Y0_N_IO/FrameData_O[13]
+ Tile_X2Y0_N_IO/FrameData_O[14] Tile_X2Y0_N_IO/FrameData_O[15] Tile_X2Y0_N_IO/FrameData_O[16]
+ Tile_X2Y0_N_IO/FrameData_O[17] Tile_X2Y0_N_IO/FrameData_O[18] Tile_X2Y0_N_IO/FrameData_O[19]
+ Tile_X2Y0_N_IO/FrameData_O[1] Tile_X2Y0_N_IO/FrameData_O[20] Tile_X2Y0_N_IO/FrameData_O[21]
+ Tile_X2Y0_N_IO/FrameData_O[22] Tile_X2Y0_N_IO/FrameData_O[23] Tile_X2Y0_N_IO/FrameData_O[24]
+ Tile_X2Y0_N_IO/FrameData_O[25] Tile_X2Y0_N_IO/FrameData_O[26] Tile_X2Y0_N_IO/FrameData_O[27]
+ Tile_X2Y0_N_IO/FrameData_O[28] Tile_X2Y0_N_IO/FrameData_O[29] Tile_X2Y0_N_IO/FrameData_O[2]
+ Tile_X2Y0_N_IO/FrameData_O[30] Tile_X2Y0_N_IO/FrameData_O[31] Tile_X2Y0_N_IO/FrameData_O[3]
+ Tile_X2Y0_N_IO/FrameData_O[4] Tile_X2Y0_N_IO/FrameData_O[5] Tile_X2Y0_N_IO/FrameData_O[6]
+ Tile_X2Y0_N_IO/FrameData_O[7] Tile_X2Y0_N_IO/FrameData_O[8] Tile_X2Y0_N_IO/FrameData_O[9]
+ Tile_X4Y0_N_term_single2/FrameData[0] Tile_X4Y0_N_term_single2/FrameData[10] Tile_X4Y0_N_term_single2/FrameData[11]
+ Tile_X4Y0_N_term_single2/FrameData[12] Tile_X4Y0_N_term_single2/FrameData[13] Tile_X4Y0_N_term_single2/FrameData[14]
+ Tile_X4Y0_N_term_single2/FrameData[15] Tile_X4Y0_N_term_single2/FrameData[16] Tile_X4Y0_N_term_single2/FrameData[17]
+ Tile_X4Y0_N_term_single2/FrameData[18] Tile_X4Y0_N_term_single2/FrameData[19] Tile_X4Y0_N_term_single2/FrameData[1]
+ Tile_X4Y0_N_term_single2/FrameData[20] Tile_X4Y0_N_term_single2/FrameData[21] Tile_X4Y0_N_term_single2/FrameData[22]
+ Tile_X4Y0_N_term_single2/FrameData[23] Tile_X4Y0_N_term_single2/FrameData[24] Tile_X4Y0_N_term_single2/FrameData[25]
+ Tile_X4Y0_N_term_single2/FrameData[26] Tile_X4Y0_N_term_single2/FrameData[27] Tile_X4Y0_N_term_single2/FrameData[28]
+ Tile_X4Y0_N_term_single2/FrameData[29] Tile_X4Y0_N_term_single2/FrameData[2] Tile_X4Y0_N_term_single2/FrameData[30]
+ Tile_X4Y0_N_term_single2/FrameData[31] Tile_X4Y0_N_term_single2/FrameData[3] Tile_X4Y0_N_term_single2/FrameData[4]
+ Tile_X4Y0_N_term_single2/FrameData[5] Tile_X4Y0_N_term_single2/FrameData[6] Tile_X4Y0_N_term_single2/FrameData[7]
+ Tile_X4Y0_N_term_single2/FrameData[8] Tile_X4Y0_N_term_single2/FrameData[9] Tile_X3Y1_LUT4AB/FrameStrobe_O[0]
+ Tile_X3Y1_LUT4AB/FrameStrobe_O[10] Tile_X3Y1_LUT4AB/FrameStrobe_O[11] Tile_X3Y1_LUT4AB/FrameStrobe_O[12]
+ Tile_X3Y1_LUT4AB/FrameStrobe_O[13] Tile_X3Y1_LUT4AB/FrameStrobe_O[14] Tile_X3Y1_LUT4AB/FrameStrobe_O[15]
+ Tile_X3Y1_LUT4AB/FrameStrobe_O[16] Tile_X3Y1_LUT4AB/FrameStrobe_O[17] Tile_X3Y1_LUT4AB/FrameStrobe_O[18]
+ Tile_X3Y1_LUT4AB/FrameStrobe_O[19] Tile_X3Y1_LUT4AB/FrameStrobe_O[1] Tile_X3Y1_LUT4AB/FrameStrobe_O[2]
+ Tile_X3Y1_LUT4AB/FrameStrobe_O[3] Tile_X3Y1_LUT4AB/FrameStrobe_O[4] Tile_X3Y1_LUT4AB/FrameStrobe_O[5]
+ Tile_X3Y1_LUT4AB/FrameStrobe_O[6] Tile_X3Y1_LUT4AB/FrameStrobe_O[7] Tile_X3Y1_LUT4AB/FrameStrobe_O[8]
+ Tile_X3Y1_LUT4AB/FrameStrobe_O[9] Tile_X3Y0_N_term_single/FrameStrobe_O[0] Tile_X3Y0_N_term_single/FrameStrobe_O[10]
+ Tile_X3Y0_N_term_single/FrameStrobe_O[11] Tile_X3Y0_N_term_single/FrameStrobe_O[12]
+ Tile_X3Y0_N_term_single/FrameStrobe_O[13] Tile_X3Y0_N_term_single/FrameStrobe_O[14]
+ Tile_X3Y0_N_term_single/FrameStrobe_O[15] Tile_X3Y0_N_term_single/FrameStrobe_O[16]
+ Tile_X3Y0_N_term_single/FrameStrobe_O[17] Tile_X3Y0_N_term_single/FrameStrobe_O[18]
+ Tile_X3Y0_N_term_single/FrameStrobe_O[19] Tile_X3Y0_N_term_single/FrameStrobe_O[1]
+ Tile_X3Y0_N_term_single/FrameStrobe_O[2] Tile_X3Y0_N_term_single/FrameStrobe_O[3]
+ Tile_X3Y0_N_term_single/FrameStrobe_O[4] Tile_X3Y0_N_term_single/FrameStrobe_O[5]
+ Tile_X3Y0_N_term_single/FrameStrobe_O[6] Tile_X3Y0_N_term_single/FrameStrobe_O[7]
+ Tile_X3Y0_N_term_single/FrameStrobe_O[8] Tile_X3Y0_N_term_single/FrameStrobe_O[9]
+ Tile_X3Y1_LUT4AB/N1BEG[0] Tile_X3Y1_LUT4AB/N1BEG[1] Tile_X3Y1_LUT4AB/N1BEG[2] Tile_X3Y1_LUT4AB/N1BEG[3]
+ Tile_X3Y1_LUT4AB/N2BEGb[0] Tile_X3Y1_LUT4AB/N2BEGb[1] Tile_X3Y1_LUT4AB/N2BEGb[2]
+ Tile_X3Y1_LUT4AB/N2BEGb[3] Tile_X3Y1_LUT4AB/N2BEGb[4] Tile_X3Y1_LUT4AB/N2BEGb[5]
+ Tile_X3Y1_LUT4AB/N2BEGb[6] Tile_X3Y1_LUT4AB/N2BEGb[7] Tile_X3Y1_LUT4AB/N2BEG[0]
+ Tile_X3Y1_LUT4AB/N2BEG[1] Tile_X3Y1_LUT4AB/N2BEG[2] Tile_X3Y1_LUT4AB/N2BEG[3] Tile_X3Y1_LUT4AB/N2BEG[4]
+ Tile_X3Y1_LUT4AB/N2BEG[5] Tile_X3Y1_LUT4AB/N2BEG[6] Tile_X3Y1_LUT4AB/N2BEG[7] Tile_X3Y1_LUT4AB/N4BEG[0]
+ Tile_X3Y1_LUT4AB/N4BEG[10] Tile_X3Y1_LUT4AB/N4BEG[11] Tile_X3Y1_LUT4AB/N4BEG[12]
+ Tile_X3Y1_LUT4AB/N4BEG[13] Tile_X3Y1_LUT4AB/N4BEG[14] Tile_X3Y1_LUT4AB/N4BEG[15]
+ Tile_X3Y1_LUT4AB/N4BEG[1] Tile_X3Y1_LUT4AB/N4BEG[2] Tile_X3Y1_LUT4AB/N4BEG[3] Tile_X3Y1_LUT4AB/N4BEG[4]
+ Tile_X3Y1_LUT4AB/N4BEG[5] Tile_X3Y1_LUT4AB/N4BEG[6] Tile_X3Y1_LUT4AB/N4BEG[7] Tile_X3Y1_LUT4AB/N4BEG[8]
+ Tile_X3Y1_LUT4AB/N4BEG[9] Tile_X3Y1_LUT4AB/NN4BEG[0] Tile_X3Y1_LUT4AB/NN4BEG[10]
+ Tile_X3Y1_LUT4AB/NN4BEG[11] Tile_X3Y1_LUT4AB/NN4BEG[12] Tile_X3Y1_LUT4AB/NN4BEG[13]
+ Tile_X3Y1_LUT4AB/NN4BEG[14] Tile_X3Y1_LUT4AB/NN4BEG[15] Tile_X3Y1_LUT4AB/NN4BEG[1]
+ Tile_X3Y1_LUT4AB/NN4BEG[2] Tile_X3Y1_LUT4AB/NN4BEG[3] Tile_X3Y1_LUT4AB/NN4BEG[4]
+ Tile_X3Y1_LUT4AB/NN4BEG[5] Tile_X3Y1_LUT4AB/NN4BEG[6] Tile_X3Y1_LUT4AB/NN4BEG[7]
+ Tile_X3Y1_LUT4AB/NN4BEG[8] Tile_X3Y1_LUT4AB/NN4BEG[9] Tile_X3Y1_LUT4AB/S1END[0]
+ Tile_X3Y1_LUT4AB/S1END[1] Tile_X3Y1_LUT4AB/S1END[2] Tile_X3Y1_LUT4AB/S1END[3] Tile_X3Y1_LUT4AB/S2MID[0]
+ Tile_X3Y1_LUT4AB/S2MID[1] Tile_X3Y1_LUT4AB/S2MID[2] Tile_X3Y1_LUT4AB/S2MID[3] Tile_X3Y1_LUT4AB/S2MID[4]
+ Tile_X3Y1_LUT4AB/S2MID[5] Tile_X3Y1_LUT4AB/S2MID[6] Tile_X3Y1_LUT4AB/S2MID[7] Tile_X3Y1_LUT4AB/S2END[0]
+ Tile_X3Y1_LUT4AB/S2END[1] Tile_X3Y1_LUT4AB/S2END[2] Tile_X3Y1_LUT4AB/S2END[3] Tile_X3Y1_LUT4AB/S2END[4]
+ Tile_X3Y1_LUT4AB/S2END[5] Tile_X3Y1_LUT4AB/S2END[6] Tile_X3Y1_LUT4AB/S2END[7] Tile_X3Y1_LUT4AB/S4END[0]
+ Tile_X3Y1_LUT4AB/S4END[10] Tile_X3Y1_LUT4AB/S4END[11] Tile_X3Y1_LUT4AB/S4END[12]
+ Tile_X3Y1_LUT4AB/S4END[13] Tile_X3Y1_LUT4AB/S4END[14] Tile_X3Y1_LUT4AB/S4END[15]
+ Tile_X3Y1_LUT4AB/S4END[1] Tile_X3Y1_LUT4AB/S4END[2] Tile_X3Y1_LUT4AB/S4END[3] Tile_X3Y1_LUT4AB/S4END[4]
+ Tile_X3Y1_LUT4AB/S4END[5] Tile_X3Y1_LUT4AB/S4END[6] Tile_X3Y1_LUT4AB/S4END[7] Tile_X3Y1_LUT4AB/S4END[8]
+ Tile_X3Y1_LUT4AB/S4END[9] Tile_X3Y1_LUT4AB/SS4END[0] Tile_X3Y1_LUT4AB/SS4END[10]
+ Tile_X3Y1_LUT4AB/SS4END[11] Tile_X3Y1_LUT4AB/SS4END[12] Tile_X3Y1_LUT4AB/SS4END[13]
+ Tile_X3Y1_LUT4AB/SS4END[14] Tile_X3Y1_LUT4AB/SS4END[15] Tile_X3Y1_LUT4AB/SS4END[1]
+ Tile_X3Y1_LUT4AB/SS4END[2] Tile_X3Y1_LUT4AB/SS4END[3] Tile_X3Y1_LUT4AB/SS4END[4]
+ Tile_X3Y1_LUT4AB/SS4END[5] Tile_X3Y1_LUT4AB/SS4END[6] Tile_X3Y1_LUT4AB/SS4END[7]
+ Tile_X3Y1_LUT4AB/SS4END[8] Tile_X3Y1_LUT4AB/SS4END[9] Tile_X3Y1_LUT4AB/UserCLKo
+ Tile_X3Y0_N_term_single/UserCLKo VGND VPWR N_term_single
XTile_X5Y3_LUT4AB Tile_X5Y4_LUT4AB/Co Tile_X5Y3_LUT4AB/Co Tile_X6Y3_LUT4AB/E1END[0]
+ Tile_X6Y3_LUT4AB/E1END[1] Tile_X6Y3_LUT4AB/E1END[2] Tile_X6Y3_LUT4AB/E1END[3] Tile_X5Y3_LUT4AB/E1END[0]
+ Tile_X5Y3_LUT4AB/E1END[1] Tile_X5Y3_LUT4AB/E1END[2] Tile_X5Y3_LUT4AB/E1END[3] Tile_X6Y3_LUT4AB/E2MID[0]
+ Tile_X6Y3_LUT4AB/E2MID[1] Tile_X6Y3_LUT4AB/E2MID[2] Tile_X6Y3_LUT4AB/E2MID[3] Tile_X6Y3_LUT4AB/E2MID[4]
+ Tile_X6Y3_LUT4AB/E2MID[5] Tile_X6Y3_LUT4AB/E2MID[6] Tile_X6Y3_LUT4AB/E2MID[7] Tile_X6Y3_LUT4AB/E2END[0]
+ Tile_X6Y3_LUT4AB/E2END[1] Tile_X6Y3_LUT4AB/E2END[2] Tile_X6Y3_LUT4AB/E2END[3] Tile_X6Y3_LUT4AB/E2END[4]
+ Tile_X6Y3_LUT4AB/E2END[5] Tile_X6Y3_LUT4AB/E2END[6] Tile_X6Y3_LUT4AB/E2END[7] Tile_X5Y3_LUT4AB/E2END[0]
+ Tile_X5Y3_LUT4AB/E2END[1] Tile_X5Y3_LUT4AB/E2END[2] Tile_X5Y3_LUT4AB/E2END[3] Tile_X5Y3_LUT4AB/E2END[4]
+ Tile_X5Y3_LUT4AB/E2END[5] Tile_X5Y3_LUT4AB/E2END[6] Tile_X5Y3_LUT4AB/E2END[7] Tile_X5Y3_LUT4AB/E2MID[0]
+ Tile_X5Y3_LUT4AB/E2MID[1] Tile_X5Y3_LUT4AB/E2MID[2] Tile_X5Y3_LUT4AB/E2MID[3] Tile_X5Y3_LUT4AB/E2MID[4]
+ Tile_X5Y3_LUT4AB/E2MID[5] Tile_X5Y3_LUT4AB/E2MID[6] Tile_X5Y3_LUT4AB/E2MID[7] Tile_X6Y3_LUT4AB/E6END[0]
+ Tile_X6Y3_LUT4AB/E6END[10] Tile_X6Y3_LUT4AB/E6END[11] Tile_X6Y3_LUT4AB/E6END[1]
+ Tile_X6Y3_LUT4AB/E6END[2] Tile_X6Y3_LUT4AB/E6END[3] Tile_X6Y3_LUT4AB/E6END[4] Tile_X6Y3_LUT4AB/E6END[5]
+ Tile_X6Y3_LUT4AB/E6END[6] Tile_X6Y3_LUT4AB/E6END[7] Tile_X6Y3_LUT4AB/E6END[8] Tile_X6Y3_LUT4AB/E6END[9]
+ Tile_X5Y3_LUT4AB/E6END[0] Tile_X5Y3_LUT4AB/E6END[10] Tile_X5Y3_LUT4AB/E6END[11]
+ Tile_X5Y3_LUT4AB/E6END[1] Tile_X5Y3_LUT4AB/E6END[2] Tile_X5Y3_LUT4AB/E6END[3] Tile_X5Y3_LUT4AB/E6END[4]
+ Tile_X5Y3_LUT4AB/E6END[5] Tile_X5Y3_LUT4AB/E6END[6] Tile_X5Y3_LUT4AB/E6END[7] Tile_X5Y3_LUT4AB/E6END[8]
+ Tile_X5Y3_LUT4AB/E6END[9] Tile_X6Y3_LUT4AB/EE4END[0] Tile_X6Y3_LUT4AB/EE4END[10]
+ Tile_X6Y3_LUT4AB/EE4END[11] Tile_X6Y3_LUT4AB/EE4END[12] Tile_X6Y3_LUT4AB/EE4END[13]
+ Tile_X6Y3_LUT4AB/EE4END[14] Tile_X6Y3_LUT4AB/EE4END[15] Tile_X6Y3_LUT4AB/EE4END[1]
+ Tile_X6Y3_LUT4AB/EE4END[2] Tile_X6Y3_LUT4AB/EE4END[3] Tile_X6Y3_LUT4AB/EE4END[4]
+ Tile_X6Y3_LUT4AB/EE4END[5] Tile_X6Y3_LUT4AB/EE4END[6] Tile_X6Y3_LUT4AB/EE4END[7]
+ Tile_X6Y3_LUT4AB/EE4END[8] Tile_X6Y3_LUT4AB/EE4END[9] Tile_X5Y3_LUT4AB/EE4END[0]
+ Tile_X5Y3_LUT4AB/EE4END[10] Tile_X5Y3_LUT4AB/EE4END[11] Tile_X5Y3_LUT4AB/EE4END[12]
+ Tile_X5Y3_LUT4AB/EE4END[13] Tile_X5Y3_LUT4AB/EE4END[14] Tile_X5Y3_LUT4AB/EE4END[15]
+ Tile_X5Y3_LUT4AB/EE4END[1] Tile_X5Y3_LUT4AB/EE4END[2] Tile_X5Y3_LUT4AB/EE4END[3]
+ Tile_X5Y3_LUT4AB/EE4END[4] Tile_X5Y3_LUT4AB/EE4END[5] Tile_X5Y3_LUT4AB/EE4END[6]
+ Tile_X5Y3_LUT4AB/EE4END[7] Tile_X5Y3_LUT4AB/EE4END[8] Tile_X5Y3_LUT4AB/EE4END[9]
+ Tile_X5Y3_LUT4AB/FrameData[0] Tile_X5Y3_LUT4AB/FrameData[10] Tile_X5Y3_LUT4AB/FrameData[11]
+ Tile_X5Y3_LUT4AB/FrameData[12] Tile_X5Y3_LUT4AB/FrameData[13] Tile_X5Y3_LUT4AB/FrameData[14]
+ Tile_X5Y3_LUT4AB/FrameData[15] Tile_X5Y3_LUT4AB/FrameData[16] Tile_X5Y3_LUT4AB/FrameData[17]
+ Tile_X5Y3_LUT4AB/FrameData[18] Tile_X5Y3_LUT4AB/FrameData[19] Tile_X5Y3_LUT4AB/FrameData[1]
+ Tile_X5Y3_LUT4AB/FrameData[20] Tile_X5Y3_LUT4AB/FrameData[21] Tile_X5Y3_LUT4AB/FrameData[22]
+ Tile_X5Y3_LUT4AB/FrameData[23] Tile_X5Y3_LUT4AB/FrameData[24] Tile_X5Y3_LUT4AB/FrameData[25]
+ Tile_X5Y3_LUT4AB/FrameData[26] Tile_X5Y3_LUT4AB/FrameData[27] Tile_X5Y3_LUT4AB/FrameData[28]
+ Tile_X5Y3_LUT4AB/FrameData[29] Tile_X5Y3_LUT4AB/FrameData[2] Tile_X5Y3_LUT4AB/FrameData[30]
+ Tile_X5Y3_LUT4AB/FrameData[31] Tile_X5Y3_LUT4AB/FrameData[3] Tile_X5Y3_LUT4AB/FrameData[4]
+ Tile_X5Y3_LUT4AB/FrameData[5] Tile_X5Y3_LUT4AB/FrameData[6] Tile_X5Y3_LUT4AB/FrameData[7]
+ Tile_X5Y3_LUT4AB/FrameData[8] Tile_X5Y3_LUT4AB/FrameData[9] Tile_X6Y3_LUT4AB/FrameData[0]
+ Tile_X6Y3_LUT4AB/FrameData[10] Tile_X6Y3_LUT4AB/FrameData[11] Tile_X6Y3_LUT4AB/FrameData[12]
+ Tile_X6Y3_LUT4AB/FrameData[13] Tile_X6Y3_LUT4AB/FrameData[14] Tile_X6Y3_LUT4AB/FrameData[15]
+ Tile_X6Y3_LUT4AB/FrameData[16] Tile_X6Y3_LUT4AB/FrameData[17] Tile_X6Y3_LUT4AB/FrameData[18]
+ Tile_X6Y3_LUT4AB/FrameData[19] Tile_X6Y3_LUT4AB/FrameData[1] Tile_X6Y3_LUT4AB/FrameData[20]
+ Tile_X6Y3_LUT4AB/FrameData[21] Tile_X6Y3_LUT4AB/FrameData[22] Tile_X6Y3_LUT4AB/FrameData[23]
+ Tile_X6Y3_LUT4AB/FrameData[24] Tile_X6Y3_LUT4AB/FrameData[25] Tile_X6Y3_LUT4AB/FrameData[26]
+ Tile_X6Y3_LUT4AB/FrameData[27] Tile_X6Y3_LUT4AB/FrameData[28] Tile_X6Y3_LUT4AB/FrameData[29]
+ Tile_X6Y3_LUT4AB/FrameData[2] Tile_X6Y3_LUT4AB/FrameData[30] Tile_X6Y3_LUT4AB/FrameData[31]
+ Tile_X6Y3_LUT4AB/FrameData[3] Tile_X6Y3_LUT4AB/FrameData[4] Tile_X6Y3_LUT4AB/FrameData[5]
+ Tile_X6Y3_LUT4AB/FrameData[6] Tile_X6Y3_LUT4AB/FrameData[7] Tile_X6Y3_LUT4AB/FrameData[8]
+ Tile_X6Y3_LUT4AB/FrameData[9] Tile_X5Y3_LUT4AB/FrameStrobe[0] Tile_X5Y3_LUT4AB/FrameStrobe[10]
+ Tile_X5Y3_LUT4AB/FrameStrobe[11] Tile_X5Y3_LUT4AB/FrameStrobe[12] Tile_X5Y3_LUT4AB/FrameStrobe[13]
+ Tile_X5Y3_LUT4AB/FrameStrobe[14] Tile_X5Y3_LUT4AB/FrameStrobe[15] Tile_X5Y3_LUT4AB/FrameStrobe[16]
+ Tile_X5Y3_LUT4AB/FrameStrobe[17] Tile_X5Y3_LUT4AB/FrameStrobe[18] Tile_X5Y3_LUT4AB/FrameStrobe[19]
+ Tile_X5Y3_LUT4AB/FrameStrobe[1] Tile_X5Y3_LUT4AB/FrameStrobe[2] Tile_X5Y3_LUT4AB/FrameStrobe[3]
+ Tile_X5Y3_LUT4AB/FrameStrobe[4] Tile_X5Y3_LUT4AB/FrameStrobe[5] Tile_X5Y3_LUT4AB/FrameStrobe[6]
+ Tile_X5Y3_LUT4AB/FrameStrobe[7] Tile_X5Y3_LUT4AB/FrameStrobe[8] Tile_X5Y3_LUT4AB/FrameStrobe[9]
+ Tile_X5Y2_LUT4AB/FrameStrobe[0] Tile_X5Y2_LUT4AB/FrameStrobe[10] Tile_X5Y2_LUT4AB/FrameStrobe[11]
+ Tile_X5Y2_LUT4AB/FrameStrobe[12] Tile_X5Y2_LUT4AB/FrameStrobe[13] Tile_X5Y2_LUT4AB/FrameStrobe[14]
+ Tile_X5Y2_LUT4AB/FrameStrobe[15] Tile_X5Y2_LUT4AB/FrameStrobe[16] Tile_X5Y2_LUT4AB/FrameStrobe[17]
+ Tile_X5Y2_LUT4AB/FrameStrobe[18] Tile_X5Y2_LUT4AB/FrameStrobe[19] Tile_X5Y2_LUT4AB/FrameStrobe[1]
+ Tile_X5Y2_LUT4AB/FrameStrobe[2] Tile_X5Y2_LUT4AB/FrameStrobe[3] Tile_X5Y2_LUT4AB/FrameStrobe[4]
+ Tile_X5Y2_LUT4AB/FrameStrobe[5] Tile_X5Y2_LUT4AB/FrameStrobe[6] Tile_X5Y2_LUT4AB/FrameStrobe[7]
+ Tile_X5Y2_LUT4AB/FrameStrobe[8] Tile_X5Y2_LUT4AB/FrameStrobe[9] Tile_X5Y3_LUT4AB/N1BEG[0]
+ Tile_X5Y3_LUT4AB/N1BEG[1] Tile_X5Y3_LUT4AB/N1BEG[2] Tile_X5Y3_LUT4AB/N1BEG[3] Tile_X5Y4_LUT4AB/N1BEG[0]
+ Tile_X5Y4_LUT4AB/N1BEG[1] Tile_X5Y4_LUT4AB/N1BEG[2] Tile_X5Y4_LUT4AB/N1BEG[3] Tile_X5Y3_LUT4AB/N2BEG[0]
+ Tile_X5Y3_LUT4AB/N2BEG[1] Tile_X5Y3_LUT4AB/N2BEG[2] Tile_X5Y3_LUT4AB/N2BEG[3] Tile_X5Y3_LUT4AB/N2BEG[4]
+ Tile_X5Y3_LUT4AB/N2BEG[5] Tile_X5Y3_LUT4AB/N2BEG[6] Tile_X5Y3_LUT4AB/N2BEG[7] Tile_X5Y2_LUT4AB/N2END[0]
+ Tile_X5Y2_LUT4AB/N2END[1] Tile_X5Y2_LUT4AB/N2END[2] Tile_X5Y2_LUT4AB/N2END[3] Tile_X5Y2_LUT4AB/N2END[4]
+ Tile_X5Y2_LUT4AB/N2END[5] Tile_X5Y2_LUT4AB/N2END[6] Tile_X5Y2_LUT4AB/N2END[7] Tile_X5Y3_LUT4AB/N2END[0]
+ Tile_X5Y3_LUT4AB/N2END[1] Tile_X5Y3_LUT4AB/N2END[2] Tile_X5Y3_LUT4AB/N2END[3] Tile_X5Y3_LUT4AB/N2END[4]
+ Tile_X5Y3_LUT4AB/N2END[5] Tile_X5Y3_LUT4AB/N2END[6] Tile_X5Y3_LUT4AB/N2END[7] Tile_X5Y4_LUT4AB/N2BEG[0]
+ Tile_X5Y4_LUT4AB/N2BEG[1] Tile_X5Y4_LUT4AB/N2BEG[2] Tile_X5Y4_LUT4AB/N2BEG[3] Tile_X5Y4_LUT4AB/N2BEG[4]
+ Tile_X5Y4_LUT4AB/N2BEG[5] Tile_X5Y4_LUT4AB/N2BEG[6] Tile_X5Y4_LUT4AB/N2BEG[7] Tile_X5Y3_LUT4AB/N4BEG[0]
+ Tile_X5Y3_LUT4AB/N4BEG[10] Tile_X5Y3_LUT4AB/N4BEG[11] Tile_X5Y3_LUT4AB/N4BEG[12]
+ Tile_X5Y3_LUT4AB/N4BEG[13] Tile_X5Y3_LUT4AB/N4BEG[14] Tile_X5Y3_LUT4AB/N4BEG[15]
+ Tile_X5Y3_LUT4AB/N4BEG[1] Tile_X5Y3_LUT4AB/N4BEG[2] Tile_X5Y3_LUT4AB/N4BEG[3] Tile_X5Y3_LUT4AB/N4BEG[4]
+ Tile_X5Y3_LUT4AB/N4BEG[5] Tile_X5Y3_LUT4AB/N4BEG[6] Tile_X5Y3_LUT4AB/N4BEG[7] Tile_X5Y3_LUT4AB/N4BEG[8]
+ Tile_X5Y3_LUT4AB/N4BEG[9] Tile_X5Y4_LUT4AB/N4BEG[0] Tile_X5Y4_LUT4AB/N4BEG[10] Tile_X5Y4_LUT4AB/N4BEG[11]
+ Tile_X5Y4_LUT4AB/N4BEG[12] Tile_X5Y4_LUT4AB/N4BEG[13] Tile_X5Y4_LUT4AB/N4BEG[14]
+ Tile_X5Y4_LUT4AB/N4BEG[15] Tile_X5Y4_LUT4AB/N4BEG[1] Tile_X5Y4_LUT4AB/N4BEG[2] Tile_X5Y4_LUT4AB/N4BEG[3]
+ Tile_X5Y4_LUT4AB/N4BEG[4] Tile_X5Y4_LUT4AB/N4BEG[5] Tile_X5Y4_LUT4AB/N4BEG[6] Tile_X5Y4_LUT4AB/N4BEG[7]
+ Tile_X5Y4_LUT4AB/N4BEG[8] Tile_X5Y4_LUT4AB/N4BEG[9] Tile_X5Y3_LUT4AB/NN4BEG[0] Tile_X5Y3_LUT4AB/NN4BEG[10]
+ Tile_X5Y3_LUT4AB/NN4BEG[11] Tile_X5Y3_LUT4AB/NN4BEG[12] Tile_X5Y3_LUT4AB/NN4BEG[13]
+ Tile_X5Y3_LUT4AB/NN4BEG[14] Tile_X5Y3_LUT4AB/NN4BEG[15] Tile_X5Y3_LUT4AB/NN4BEG[1]
+ Tile_X5Y3_LUT4AB/NN4BEG[2] Tile_X5Y3_LUT4AB/NN4BEG[3] Tile_X5Y3_LUT4AB/NN4BEG[4]
+ Tile_X5Y3_LUT4AB/NN4BEG[5] Tile_X5Y3_LUT4AB/NN4BEG[6] Tile_X5Y3_LUT4AB/NN4BEG[7]
+ Tile_X5Y3_LUT4AB/NN4BEG[8] Tile_X5Y3_LUT4AB/NN4BEG[9] Tile_X5Y4_LUT4AB/NN4BEG[0]
+ Tile_X5Y4_LUT4AB/NN4BEG[10] Tile_X5Y4_LUT4AB/NN4BEG[11] Tile_X5Y4_LUT4AB/NN4BEG[12]
+ Tile_X5Y4_LUT4AB/NN4BEG[13] Tile_X5Y4_LUT4AB/NN4BEG[14] Tile_X5Y4_LUT4AB/NN4BEG[15]
+ Tile_X5Y4_LUT4AB/NN4BEG[1] Tile_X5Y4_LUT4AB/NN4BEG[2] Tile_X5Y4_LUT4AB/NN4BEG[3]
+ Tile_X5Y4_LUT4AB/NN4BEG[4] Tile_X5Y4_LUT4AB/NN4BEG[5] Tile_X5Y4_LUT4AB/NN4BEG[6]
+ Tile_X5Y4_LUT4AB/NN4BEG[7] Tile_X5Y4_LUT4AB/NN4BEG[8] Tile_X5Y4_LUT4AB/NN4BEG[9]
+ Tile_X5Y4_LUT4AB/S1END[0] Tile_X5Y4_LUT4AB/S1END[1] Tile_X5Y4_LUT4AB/S1END[2] Tile_X5Y4_LUT4AB/S1END[3]
+ Tile_X5Y3_LUT4AB/S1END[0] Tile_X5Y3_LUT4AB/S1END[1] Tile_X5Y3_LUT4AB/S1END[2] Tile_X5Y3_LUT4AB/S1END[3]
+ Tile_X5Y4_LUT4AB/S2MID[0] Tile_X5Y4_LUT4AB/S2MID[1] Tile_X5Y4_LUT4AB/S2MID[2] Tile_X5Y4_LUT4AB/S2MID[3]
+ Tile_X5Y4_LUT4AB/S2MID[4] Tile_X5Y4_LUT4AB/S2MID[5] Tile_X5Y4_LUT4AB/S2MID[6] Tile_X5Y4_LUT4AB/S2MID[7]
+ Tile_X5Y4_LUT4AB/S2END[0] Tile_X5Y4_LUT4AB/S2END[1] Tile_X5Y4_LUT4AB/S2END[2] Tile_X5Y4_LUT4AB/S2END[3]
+ Tile_X5Y4_LUT4AB/S2END[4] Tile_X5Y4_LUT4AB/S2END[5] Tile_X5Y4_LUT4AB/S2END[6] Tile_X5Y4_LUT4AB/S2END[7]
+ Tile_X5Y3_LUT4AB/S2END[0] Tile_X5Y3_LUT4AB/S2END[1] Tile_X5Y3_LUT4AB/S2END[2] Tile_X5Y3_LUT4AB/S2END[3]
+ Tile_X5Y3_LUT4AB/S2END[4] Tile_X5Y3_LUT4AB/S2END[5] Tile_X5Y3_LUT4AB/S2END[6] Tile_X5Y3_LUT4AB/S2END[7]
+ Tile_X5Y3_LUT4AB/S2MID[0] Tile_X5Y3_LUT4AB/S2MID[1] Tile_X5Y3_LUT4AB/S2MID[2] Tile_X5Y3_LUT4AB/S2MID[3]
+ Tile_X5Y3_LUT4AB/S2MID[4] Tile_X5Y3_LUT4AB/S2MID[5] Tile_X5Y3_LUT4AB/S2MID[6] Tile_X5Y3_LUT4AB/S2MID[7]
+ Tile_X5Y4_LUT4AB/S4END[0] Tile_X5Y4_LUT4AB/S4END[10] Tile_X5Y4_LUT4AB/S4END[11]
+ Tile_X5Y4_LUT4AB/S4END[12] Tile_X5Y4_LUT4AB/S4END[13] Tile_X5Y4_LUT4AB/S4END[14]
+ Tile_X5Y4_LUT4AB/S4END[15] Tile_X5Y4_LUT4AB/S4END[1] Tile_X5Y4_LUT4AB/S4END[2] Tile_X5Y4_LUT4AB/S4END[3]
+ Tile_X5Y4_LUT4AB/S4END[4] Tile_X5Y4_LUT4AB/S4END[5] Tile_X5Y4_LUT4AB/S4END[6] Tile_X5Y4_LUT4AB/S4END[7]
+ Tile_X5Y4_LUT4AB/S4END[8] Tile_X5Y4_LUT4AB/S4END[9] Tile_X5Y3_LUT4AB/S4END[0] Tile_X5Y3_LUT4AB/S4END[10]
+ Tile_X5Y3_LUT4AB/S4END[11] Tile_X5Y3_LUT4AB/S4END[12] Tile_X5Y3_LUT4AB/S4END[13]
+ Tile_X5Y3_LUT4AB/S4END[14] Tile_X5Y3_LUT4AB/S4END[15] Tile_X5Y3_LUT4AB/S4END[1]
+ Tile_X5Y3_LUT4AB/S4END[2] Tile_X5Y3_LUT4AB/S4END[3] Tile_X5Y3_LUT4AB/S4END[4] Tile_X5Y3_LUT4AB/S4END[5]
+ Tile_X5Y3_LUT4AB/S4END[6] Tile_X5Y3_LUT4AB/S4END[7] Tile_X5Y3_LUT4AB/S4END[8] Tile_X5Y3_LUT4AB/S4END[9]
+ Tile_X5Y4_LUT4AB/SS4END[0] Tile_X5Y4_LUT4AB/SS4END[10] Tile_X5Y4_LUT4AB/SS4END[11]
+ Tile_X5Y4_LUT4AB/SS4END[12] Tile_X5Y4_LUT4AB/SS4END[13] Tile_X5Y4_LUT4AB/SS4END[14]
+ Tile_X5Y4_LUT4AB/SS4END[15] Tile_X5Y4_LUT4AB/SS4END[1] Tile_X5Y4_LUT4AB/SS4END[2]
+ Tile_X5Y4_LUT4AB/SS4END[3] Tile_X5Y4_LUT4AB/SS4END[4] Tile_X5Y4_LUT4AB/SS4END[5]
+ Tile_X5Y4_LUT4AB/SS4END[6] Tile_X5Y4_LUT4AB/SS4END[7] Tile_X5Y4_LUT4AB/SS4END[8]
+ Tile_X5Y4_LUT4AB/SS4END[9] Tile_X5Y3_LUT4AB/SS4END[0] Tile_X5Y3_LUT4AB/SS4END[10]
+ Tile_X5Y3_LUT4AB/SS4END[11] Tile_X5Y3_LUT4AB/SS4END[12] Tile_X5Y3_LUT4AB/SS4END[13]
+ Tile_X5Y3_LUT4AB/SS4END[14] Tile_X5Y3_LUT4AB/SS4END[15] Tile_X5Y3_LUT4AB/SS4END[1]
+ Tile_X5Y3_LUT4AB/SS4END[2] Tile_X5Y3_LUT4AB/SS4END[3] Tile_X5Y3_LUT4AB/SS4END[4]
+ Tile_X5Y3_LUT4AB/SS4END[5] Tile_X5Y3_LUT4AB/SS4END[6] Tile_X5Y3_LUT4AB/SS4END[7]
+ Tile_X5Y3_LUT4AB/SS4END[8] Tile_X5Y3_LUT4AB/SS4END[9] Tile_X5Y3_LUT4AB/UserCLK Tile_X5Y2_LUT4AB/UserCLK
+ VGND VPWR Tile_X5Y3_LUT4AB/W1BEG[0] Tile_X5Y3_LUT4AB/W1BEG[1] Tile_X5Y3_LUT4AB/W1BEG[2]
+ Tile_X5Y3_LUT4AB/W1BEG[3] Tile_X6Y3_LUT4AB/W1BEG[0] Tile_X6Y3_LUT4AB/W1BEG[1] Tile_X6Y3_LUT4AB/W1BEG[2]
+ Tile_X6Y3_LUT4AB/W1BEG[3] Tile_X5Y3_LUT4AB/W2BEG[0] Tile_X5Y3_LUT4AB/W2BEG[1] Tile_X5Y3_LUT4AB/W2BEG[2]
+ Tile_X5Y3_LUT4AB/W2BEG[3] Tile_X5Y3_LUT4AB/W2BEG[4] Tile_X5Y3_LUT4AB/W2BEG[5] Tile_X5Y3_LUT4AB/W2BEG[6]
+ Tile_X5Y3_LUT4AB/W2BEG[7] Tile_X5Y3_LUT4AB/W2BEGb[0] Tile_X5Y3_LUT4AB/W2BEGb[1]
+ Tile_X5Y3_LUT4AB/W2BEGb[2] Tile_X5Y3_LUT4AB/W2BEGb[3] Tile_X5Y3_LUT4AB/W2BEGb[4]
+ Tile_X5Y3_LUT4AB/W2BEGb[5] Tile_X5Y3_LUT4AB/W2BEGb[6] Tile_X5Y3_LUT4AB/W2BEGb[7]
+ Tile_X5Y3_LUT4AB/W2END[0] Tile_X5Y3_LUT4AB/W2END[1] Tile_X5Y3_LUT4AB/W2END[2] Tile_X5Y3_LUT4AB/W2END[3]
+ Tile_X5Y3_LUT4AB/W2END[4] Tile_X5Y3_LUT4AB/W2END[5] Tile_X5Y3_LUT4AB/W2END[6] Tile_X5Y3_LUT4AB/W2END[7]
+ Tile_X6Y3_LUT4AB/W2BEG[0] Tile_X6Y3_LUT4AB/W2BEG[1] Tile_X6Y3_LUT4AB/W2BEG[2] Tile_X6Y3_LUT4AB/W2BEG[3]
+ Tile_X6Y3_LUT4AB/W2BEG[4] Tile_X6Y3_LUT4AB/W2BEG[5] Tile_X6Y3_LUT4AB/W2BEG[6] Tile_X6Y3_LUT4AB/W2BEG[7]
+ Tile_X5Y3_LUT4AB/W6BEG[0] Tile_X5Y3_LUT4AB/W6BEG[10] Tile_X5Y3_LUT4AB/W6BEG[11]
+ Tile_X5Y3_LUT4AB/W6BEG[1] Tile_X5Y3_LUT4AB/W6BEG[2] Tile_X5Y3_LUT4AB/W6BEG[3] Tile_X5Y3_LUT4AB/W6BEG[4]
+ Tile_X5Y3_LUT4AB/W6BEG[5] Tile_X5Y3_LUT4AB/W6BEG[6] Tile_X5Y3_LUT4AB/W6BEG[7] Tile_X5Y3_LUT4AB/W6BEG[8]
+ Tile_X5Y3_LUT4AB/W6BEG[9] Tile_X6Y3_LUT4AB/W6BEG[0] Tile_X6Y3_LUT4AB/W6BEG[10] Tile_X6Y3_LUT4AB/W6BEG[11]
+ Tile_X6Y3_LUT4AB/W6BEG[1] Tile_X6Y3_LUT4AB/W6BEG[2] Tile_X6Y3_LUT4AB/W6BEG[3] Tile_X6Y3_LUT4AB/W6BEG[4]
+ Tile_X6Y3_LUT4AB/W6BEG[5] Tile_X6Y3_LUT4AB/W6BEG[6] Tile_X6Y3_LUT4AB/W6BEG[7] Tile_X6Y3_LUT4AB/W6BEG[8]
+ Tile_X6Y3_LUT4AB/W6BEG[9] Tile_X5Y3_LUT4AB/WW4BEG[0] Tile_X5Y3_LUT4AB/WW4BEG[10]
+ Tile_X5Y3_LUT4AB/WW4BEG[11] Tile_X5Y3_LUT4AB/WW4BEG[12] Tile_X5Y3_LUT4AB/WW4BEG[13]
+ Tile_X5Y3_LUT4AB/WW4BEG[14] Tile_X5Y3_LUT4AB/WW4BEG[15] Tile_X5Y3_LUT4AB/WW4BEG[1]
+ Tile_X5Y3_LUT4AB/WW4BEG[2] Tile_X5Y3_LUT4AB/WW4BEG[3] Tile_X5Y3_LUT4AB/WW4BEG[4]
+ Tile_X5Y3_LUT4AB/WW4BEG[5] Tile_X5Y3_LUT4AB/WW4BEG[6] Tile_X5Y3_LUT4AB/WW4BEG[7]
+ Tile_X5Y3_LUT4AB/WW4BEG[8] Tile_X5Y3_LUT4AB/WW4BEG[9] Tile_X6Y3_LUT4AB/WW4BEG[0]
+ Tile_X6Y3_LUT4AB/WW4BEG[10] Tile_X6Y3_LUT4AB/WW4BEG[11] Tile_X6Y3_LUT4AB/WW4BEG[12]
+ Tile_X6Y3_LUT4AB/WW4BEG[13] Tile_X6Y3_LUT4AB/WW4BEG[14] Tile_X6Y3_LUT4AB/WW4BEG[15]
+ Tile_X6Y3_LUT4AB/WW4BEG[1] Tile_X6Y3_LUT4AB/WW4BEG[2] Tile_X6Y3_LUT4AB/WW4BEG[3]
+ Tile_X6Y3_LUT4AB/WW4BEG[4] Tile_X6Y3_LUT4AB/WW4BEG[5] Tile_X6Y3_LUT4AB/WW4BEG[6]
+ Tile_X6Y3_LUT4AB/WW4BEG[7] Tile_X6Y3_LUT4AB/WW4BEG[8] Tile_X6Y3_LUT4AB/WW4BEG[9]
+ LUT4AB
XTile_X8Y8_LUT4AB Tile_X8Y9_LUT4AB/Co Tile_X8Y8_LUT4AB/Co Tile_X9Y8_LUT4AB/E1END[0]
+ Tile_X9Y8_LUT4AB/E1END[1] Tile_X9Y8_LUT4AB/E1END[2] Tile_X9Y8_LUT4AB/E1END[3] Tile_X8Y8_LUT4AB/E1END[0]
+ Tile_X8Y8_LUT4AB/E1END[1] Tile_X8Y8_LUT4AB/E1END[2] Tile_X8Y8_LUT4AB/E1END[3] Tile_X9Y8_LUT4AB/E2MID[0]
+ Tile_X9Y8_LUT4AB/E2MID[1] Tile_X9Y8_LUT4AB/E2MID[2] Tile_X9Y8_LUT4AB/E2MID[3] Tile_X9Y8_LUT4AB/E2MID[4]
+ Tile_X9Y8_LUT4AB/E2MID[5] Tile_X9Y8_LUT4AB/E2MID[6] Tile_X9Y8_LUT4AB/E2MID[7] Tile_X9Y8_LUT4AB/E2END[0]
+ Tile_X9Y8_LUT4AB/E2END[1] Tile_X9Y8_LUT4AB/E2END[2] Tile_X9Y8_LUT4AB/E2END[3] Tile_X9Y8_LUT4AB/E2END[4]
+ Tile_X9Y8_LUT4AB/E2END[5] Tile_X9Y8_LUT4AB/E2END[6] Tile_X9Y8_LUT4AB/E2END[7] Tile_X8Y8_LUT4AB/E2END[0]
+ Tile_X8Y8_LUT4AB/E2END[1] Tile_X8Y8_LUT4AB/E2END[2] Tile_X8Y8_LUT4AB/E2END[3] Tile_X8Y8_LUT4AB/E2END[4]
+ Tile_X8Y8_LUT4AB/E2END[5] Tile_X8Y8_LUT4AB/E2END[6] Tile_X8Y8_LUT4AB/E2END[7] Tile_X8Y8_LUT4AB/E2MID[0]
+ Tile_X8Y8_LUT4AB/E2MID[1] Tile_X8Y8_LUT4AB/E2MID[2] Tile_X8Y8_LUT4AB/E2MID[3] Tile_X8Y8_LUT4AB/E2MID[4]
+ Tile_X8Y8_LUT4AB/E2MID[5] Tile_X8Y8_LUT4AB/E2MID[6] Tile_X8Y8_LUT4AB/E2MID[7] Tile_X9Y8_LUT4AB/E6END[0]
+ Tile_X9Y8_LUT4AB/E6END[10] Tile_X9Y8_LUT4AB/E6END[11] Tile_X9Y8_LUT4AB/E6END[1]
+ Tile_X9Y8_LUT4AB/E6END[2] Tile_X9Y8_LUT4AB/E6END[3] Tile_X9Y8_LUT4AB/E6END[4] Tile_X9Y8_LUT4AB/E6END[5]
+ Tile_X9Y8_LUT4AB/E6END[6] Tile_X9Y8_LUT4AB/E6END[7] Tile_X9Y8_LUT4AB/E6END[8] Tile_X9Y8_LUT4AB/E6END[9]
+ Tile_X8Y8_LUT4AB/E6END[0] Tile_X8Y8_LUT4AB/E6END[10] Tile_X8Y8_LUT4AB/E6END[11]
+ Tile_X8Y8_LUT4AB/E6END[1] Tile_X8Y8_LUT4AB/E6END[2] Tile_X8Y8_LUT4AB/E6END[3] Tile_X8Y8_LUT4AB/E6END[4]
+ Tile_X8Y8_LUT4AB/E6END[5] Tile_X8Y8_LUT4AB/E6END[6] Tile_X8Y8_LUT4AB/E6END[7] Tile_X8Y8_LUT4AB/E6END[8]
+ Tile_X8Y8_LUT4AB/E6END[9] Tile_X9Y8_LUT4AB/EE4END[0] Tile_X9Y8_LUT4AB/EE4END[10]
+ Tile_X9Y8_LUT4AB/EE4END[11] Tile_X9Y8_LUT4AB/EE4END[12] Tile_X9Y8_LUT4AB/EE4END[13]
+ Tile_X9Y8_LUT4AB/EE4END[14] Tile_X9Y8_LUT4AB/EE4END[15] Tile_X9Y8_LUT4AB/EE4END[1]
+ Tile_X9Y8_LUT4AB/EE4END[2] Tile_X9Y8_LUT4AB/EE4END[3] Tile_X9Y8_LUT4AB/EE4END[4]
+ Tile_X9Y8_LUT4AB/EE4END[5] Tile_X9Y8_LUT4AB/EE4END[6] Tile_X9Y8_LUT4AB/EE4END[7]
+ Tile_X9Y8_LUT4AB/EE4END[8] Tile_X9Y8_LUT4AB/EE4END[9] Tile_X8Y8_LUT4AB/EE4END[0]
+ Tile_X8Y8_LUT4AB/EE4END[10] Tile_X8Y8_LUT4AB/EE4END[11] Tile_X8Y8_LUT4AB/EE4END[12]
+ Tile_X8Y8_LUT4AB/EE4END[13] Tile_X8Y8_LUT4AB/EE4END[14] Tile_X8Y8_LUT4AB/EE4END[15]
+ Tile_X8Y8_LUT4AB/EE4END[1] Tile_X8Y8_LUT4AB/EE4END[2] Tile_X8Y8_LUT4AB/EE4END[3]
+ Tile_X8Y8_LUT4AB/EE4END[4] Tile_X8Y8_LUT4AB/EE4END[5] Tile_X8Y8_LUT4AB/EE4END[6]
+ Tile_X8Y8_LUT4AB/EE4END[7] Tile_X8Y8_LUT4AB/EE4END[8] Tile_X8Y8_LUT4AB/EE4END[9]
+ Tile_X8Y8_LUT4AB/FrameData[0] Tile_X8Y8_LUT4AB/FrameData[10] Tile_X8Y8_LUT4AB/FrameData[11]
+ Tile_X8Y8_LUT4AB/FrameData[12] Tile_X8Y8_LUT4AB/FrameData[13] Tile_X8Y8_LUT4AB/FrameData[14]
+ Tile_X8Y8_LUT4AB/FrameData[15] Tile_X8Y8_LUT4AB/FrameData[16] Tile_X8Y8_LUT4AB/FrameData[17]
+ Tile_X8Y8_LUT4AB/FrameData[18] Tile_X8Y8_LUT4AB/FrameData[19] Tile_X8Y8_LUT4AB/FrameData[1]
+ Tile_X8Y8_LUT4AB/FrameData[20] Tile_X8Y8_LUT4AB/FrameData[21] Tile_X8Y8_LUT4AB/FrameData[22]
+ Tile_X8Y8_LUT4AB/FrameData[23] Tile_X8Y8_LUT4AB/FrameData[24] Tile_X8Y8_LUT4AB/FrameData[25]
+ Tile_X8Y8_LUT4AB/FrameData[26] Tile_X8Y8_LUT4AB/FrameData[27] Tile_X8Y8_LUT4AB/FrameData[28]
+ Tile_X8Y8_LUT4AB/FrameData[29] Tile_X8Y8_LUT4AB/FrameData[2] Tile_X8Y8_LUT4AB/FrameData[30]
+ Tile_X8Y8_LUT4AB/FrameData[31] Tile_X8Y8_LUT4AB/FrameData[3] Tile_X8Y8_LUT4AB/FrameData[4]
+ Tile_X8Y8_LUT4AB/FrameData[5] Tile_X8Y8_LUT4AB/FrameData[6] Tile_X8Y8_LUT4AB/FrameData[7]
+ Tile_X8Y8_LUT4AB/FrameData[8] Tile_X8Y8_LUT4AB/FrameData[9] Tile_X9Y8_LUT4AB/FrameData[0]
+ Tile_X9Y8_LUT4AB/FrameData[10] Tile_X9Y8_LUT4AB/FrameData[11] Tile_X9Y8_LUT4AB/FrameData[12]
+ Tile_X9Y8_LUT4AB/FrameData[13] Tile_X9Y8_LUT4AB/FrameData[14] Tile_X9Y8_LUT4AB/FrameData[15]
+ Tile_X9Y8_LUT4AB/FrameData[16] Tile_X9Y8_LUT4AB/FrameData[17] Tile_X9Y8_LUT4AB/FrameData[18]
+ Tile_X9Y8_LUT4AB/FrameData[19] Tile_X9Y8_LUT4AB/FrameData[1] Tile_X9Y8_LUT4AB/FrameData[20]
+ Tile_X9Y8_LUT4AB/FrameData[21] Tile_X9Y8_LUT4AB/FrameData[22] Tile_X9Y8_LUT4AB/FrameData[23]
+ Tile_X9Y8_LUT4AB/FrameData[24] Tile_X9Y8_LUT4AB/FrameData[25] Tile_X9Y8_LUT4AB/FrameData[26]
+ Tile_X9Y8_LUT4AB/FrameData[27] Tile_X9Y8_LUT4AB/FrameData[28] Tile_X9Y8_LUT4AB/FrameData[29]
+ Tile_X9Y8_LUT4AB/FrameData[2] Tile_X9Y8_LUT4AB/FrameData[30] Tile_X9Y8_LUT4AB/FrameData[31]
+ Tile_X9Y8_LUT4AB/FrameData[3] Tile_X9Y8_LUT4AB/FrameData[4] Tile_X9Y8_LUT4AB/FrameData[5]
+ Tile_X9Y8_LUT4AB/FrameData[6] Tile_X9Y8_LUT4AB/FrameData[7] Tile_X9Y8_LUT4AB/FrameData[8]
+ Tile_X9Y8_LUT4AB/FrameData[9] Tile_X8Y8_LUT4AB/FrameStrobe[0] Tile_X8Y8_LUT4AB/FrameStrobe[10]
+ Tile_X8Y8_LUT4AB/FrameStrobe[11] Tile_X8Y8_LUT4AB/FrameStrobe[12] Tile_X8Y8_LUT4AB/FrameStrobe[13]
+ Tile_X8Y8_LUT4AB/FrameStrobe[14] Tile_X8Y8_LUT4AB/FrameStrobe[15] Tile_X8Y8_LUT4AB/FrameStrobe[16]
+ Tile_X8Y8_LUT4AB/FrameStrobe[17] Tile_X8Y8_LUT4AB/FrameStrobe[18] Tile_X8Y8_LUT4AB/FrameStrobe[19]
+ Tile_X8Y8_LUT4AB/FrameStrobe[1] Tile_X8Y8_LUT4AB/FrameStrobe[2] Tile_X8Y8_LUT4AB/FrameStrobe[3]
+ Tile_X8Y8_LUT4AB/FrameStrobe[4] Tile_X8Y8_LUT4AB/FrameStrobe[5] Tile_X8Y8_LUT4AB/FrameStrobe[6]
+ Tile_X8Y8_LUT4AB/FrameStrobe[7] Tile_X8Y8_LUT4AB/FrameStrobe[8] Tile_X8Y8_LUT4AB/FrameStrobe[9]
+ Tile_X8Y7_LUT4AB/FrameStrobe[0] Tile_X8Y7_LUT4AB/FrameStrobe[10] Tile_X8Y7_LUT4AB/FrameStrobe[11]
+ Tile_X8Y7_LUT4AB/FrameStrobe[12] Tile_X8Y7_LUT4AB/FrameStrobe[13] Tile_X8Y7_LUT4AB/FrameStrobe[14]
+ Tile_X8Y7_LUT4AB/FrameStrobe[15] Tile_X8Y7_LUT4AB/FrameStrobe[16] Tile_X8Y7_LUT4AB/FrameStrobe[17]
+ Tile_X8Y7_LUT4AB/FrameStrobe[18] Tile_X8Y7_LUT4AB/FrameStrobe[19] Tile_X8Y7_LUT4AB/FrameStrobe[1]
+ Tile_X8Y7_LUT4AB/FrameStrobe[2] Tile_X8Y7_LUT4AB/FrameStrobe[3] Tile_X8Y7_LUT4AB/FrameStrobe[4]
+ Tile_X8Y7_LUT4AB/FrameStrobe[5] Tile_X8Y7_LUT4AB/FrameStrobe[6] Tile_X8Y7_LUT4AB/FrameStrobe[7]
+ Tile_X8Y7_LUT4AB/FrameStrobe[8] Tile_X8Y7_LUT4AB/FrameStrobe[9] Tile_X8Y8_LUT4AB/N1BEG[0]
+ Tile_X8Y8_LUT4AB/N1BEG[1] Tile_X8Y8_LUT4AB/N1BEG[2] Tile_X8Y8_LUT4AB/N1BEG[3] Tile_X8Y9_LUT4AB/N1BEG[0]
+ Tile_X8Y9_LUT4AB/N1BEG[1] Tile_X8Y9_LUT4AB/N1BEG[2] Tile_X8Y9_LUT4AB/N1BEG[3] Tile_X8Y8_LUT4AB/N2BEG[0]
+ Tile_X8Y8_LUT4AB/N2BEG[1] Tile_X8Y8_LUT4AB/N2BEG[2] Tile_X8Y8_LUT4AB/N2BEG[3] Tile_X8Y8_LUT4AB/N2BEG[4]
+ Tile_X8Y8_LUT4AB/N2BEG[5] Tile_X8Y8_LUT4AB/N2BEG[6] Tile_X8Y8_LUT4AB/N2BEG[7] Tile_X8Y7_LUT4AB/N2END[0]
+ Tile_X8Y7_LUT4AB/N2END[1] Tile_X8Y7_LUT4AB/N2END[2] Tile_X8Y7_LUT4AB/N2END[3] Tile_X8Y7_LUT4AB/N2END[4]
+ Tile_X8Y7_LUT4AB/N2END[5] Tile_X8Y7_LUT4AB/N2END[6] Tile_X8Y7_LUT4AB/N2END[7] Tile_X8Y8_LUT4AB/N2END[0]
+ Tile_X8Y8_LUT4AB/N2END[1] Tile_X8Y8_LUT4AB/N2END[2] Tile_X8Y8_LUT4AB/N2END[3] Tile_X8Y8_LUT4AB/N2END[4]
+ Tile_X8Y8_LUT4AB/N2END[5] Tile_X8Y8_LUT4AB/N2END[6] Tile_X8Y8_LUT4AB/N2END[7] Tile_X8Y9_LUT4AB/N2BEG[0]
+ Tile_X8Y9_LUT4AB/N2BEG[1] Tile_X8Y9_LUT4AB/N2BEG[2] Tile_X8Y9_LUT4AB/N2BEG[3] Tile_X8Y9_LUT4AB/N2BEG[4]
+ Tile_X8Y9_LUT4AB/N2BEG[5] Tile_X8Y9_LUT4AB/N2BEG[6] Tile_X8Y9_LUT4AB/N2BEG[7] Tile_X8Y8_LUT4AB/N4BEG[0]
+ Tile_X8Y8_LUT4AB/N4BEG[10] Tile_X8Y8_LUT4AB/N4BEG[11] Tile_X8Y8_LUT4AB/N4BEG[12]
+ Tile_X8Y8_LUT4AB/N4BEG[13] Tile_X8Y8_LUT4AB/N4BEG[14] Tile_X8Y8_LUT4AB/N4BEG[15]
+ Tile_X8Y8_LUT4AB/N4BEG[1] Tile_X8Y8_LUT4AB/N4BEG[2] Tile_X8Y8_LUT4AB/N4BEG[3] Tile_X8Y8_LUT4AB/N4BEG[4]
+ Tile_X8Y8_LUT4AB/N4BEG[5] Tile_X8Y8_LUT4AB/N4BEG[6] Tile_X8Y8_LUT4AB/N4BEG[7] Tile_X8Y8_LUT4AB/N4BEG[8]
+ Tile_X8Y8_LUT4AB/N4BEG[9] Tile_X8Y9_LUT4AB/N4BEG[0] Tile_X8Y9_LUT4AB/N4BEG[10] Tile_X8Y9_LUT4AB/N4BEG[11]
+ Tile_X8Y9_LUT4AB/N4BEG[12] Tile_X8Y9_LUT4AB/N4BEG[13] Tile_X8Y9_LUT4AB/N4BEG[14]
+ Tile_X8Y9_LUT4AB/N4BEG[15] Tile_X8Y9_LUT4AB/N4BEG[1] Tile_X8Y9_LUT4AB/N4BEG[2] Tile_X8Y9_LUT4AB/N4BEG[3]
+ Tile_X8Y9_LUT4AB/N4BEG[4] Tile_X8Y9_LUT4AB/N4BEG[5] Tile_X8Y9_LUT4AB/N4BEG[6] Tile_X8Y9_LUT4AB/N4BEG[7]
+ Tile_X8Y9_LUT4AB/N4BEG[8] Tile_X8Y9_LUT4AB/N4BEG[9] Tile_X8Y8_LUT4AB/NN4BEG[0] Tile_X8Y8_LUT4AB/NN4BEG[10]
+ Tile_X8Y8_LUT4AB/NN4BEG[11] Tile_X8Y8_LUT4AB/NN4BEG[12] Tile_X8Y8_LUT4AB/NN4BEG[13]
+ Tile_X8Y8_LUT4AB/NN4BEG[14] Tile_X8Y8_LUT4AB/NN4BEG[15] Tile_X8Y8_LUT4AB/NN4BEG[1]
+ Tile_X8Y8_LUT4AB/NN4BEG[2] Tile_X8Y8_LUT4AB/NN4BEG[3] Tile_X8Y8_LUT4AB/NN4BEG[4]
+ Tile_X8Y8_LUT4AB/NN4BEG[5] Tile_X8Y8_LUT4AB/NN4BEG[6] Tile_X8Y8_LUT4AB/NN4BEG[7]
+ Tile_X8Y8_LUT4AB/NN4BEG[8] Tile_X8Y8_LUT4AB/NN4BEG[9] Tile_X8Y9_LUT4AB/NN4BEG[0]
+ Tile_X8Y9_LUT4AB/NN4BEG[10] Tile_X8Y9_LUT4AB/NN4BEG[11] Tile_X8Y9_LUT4AB/NN4BEG[12]
+ Tile_X8Y9_LUT4AB/NN4BEG[13] Tile_X8Y9_LUT4AB/NN4BEG[14] Tile_X8Y9_LUT4AB/NN4BEG[15]
+ Tile_X8Y9_LUT4AB/NN4BEG[1] Tile_X8Y9_LUT4AB/NN4BEG[2] Tile_X8Y9_LUT4AB/NN4BEG[3]
+ Tile_X8Y9_LUT4AB/NN4BEG[4] Tile_X8Y9_LUT4AB/NN4BEG[5] Tile_X8Y9_LUT4AB/NN4BEG[6]
+ Tile_X8Y9_LUT4AB/NN4BEG[7] Tile_X8Y9_LUT4AB/NN4BEG[8] Tile_X8Y9_LUT4AB/NN4BEG[9]
+ Tile_X8Y9_LUT4AB/S1END[0] Tile_X8Y9_LUT4AB/S1END[1] Tile_X8Y9_LUT4AB/S1END[2] Tile_X8Y9_LUT4AB/S1END[3]
+ Tile_X8Y8_LUT4AB/S1END[0] Tile_X8Y8_LUT4AB/S1END[1] Tile_X8Y8_LUT4AB/S1END[2] Tile_X8Y8_LUT4AB/S1END[3]
+ Tile_X8Y9_LUT4AB/S2MID[0] Tile_X8Y9_LUT4AB/S2MID[1] Tile_X8Y9_LUT4AB/S2MID[2] Tile_X8Y9_LUT4AB/S2MID[3]
+ Tile_X8Y9_LUT4AB/S2MID[4] Tile_X8Y9_LUT4AB/S2MID[5] Tile_X8Y9_LUT4AB/S2MID[6] Tile_X8Y9_LUT4AB/S2MID[7]
+ Tile_X8Y9_LUT4AB/S2END[0] Tile_X8Y9_LUT4AB/S2END[1] Tile_X8Y9_LUT4AB/S2END[2] Tile_X8Y9_LUT4AB/S2END[3]
+ Tile_X8Y9_LUT4AB/S2END[4] Tile_X8Y9_LUT4AB/S2END[5] Tile_X8Y9_LUT4AB/S2END[6] Tile_X8Y9_LUT4AB/S2END[7]
+ Tile_X8Y8_LUT4AB/S2END[0] Tile_X8Y8_LUT4AB/S2END[1] Tile_X8Y8_LUT4AB/S2END[2] Tile_X8Y8_LUT4AB/S2END[3]
+ Tile_X8Y8_LUT4AB/S2END[4] Tile_X8Y8_LUT4AB/S2END[5] Tile_X8Y8_LUT4AB/S2END[6] Tile_X8Y8_LUT4AB/S2END[7]
+ Tile_X8Y8_LUT4AB/S2MID[0] Tile_X8Y8_LUT4AB/S2MID[1] Tile_X8Y8_LUT4AB/S2MID[2] Tile_X8Y8_LUT4AB/S2MID[3]
+ Tile_X8Y8_LUT4AB/S2MID[4] Tile_X8Y8_LUT4AB/S2MID[5] Tile_X8Y8_LUT4AB/S2MID[6] Tile_X8Y8_LUT4AB/S2MID[7]
+ Tile_X8Y9_LUT4AB/S4END[0] Tile_X8Y9_LUT4AB/S4END[10] Tile_X8Y9_LUT4AB/S4END[11]
+ Tile_X8Y9_LUT4AB/S4END[12] Tile_X8Y9_LUT4AB/S4END[13] Tile_X8Y9_LUT4AB/S4END[14]
+ Tile_X8Y9_LUT4AB/S4END[15] Tile_X8Y9_LUT4AB/S4END[1] Tile_X8Y9_LUT4AB/S4END[2] Tile_X8Y9_LUT4AB/S4END[3]
+ Tile_X8Y9_LUT4AB/S4END[4] Tile_X8Y9_LUT4AB/S4END[5] Tile_X8Y9_LUT4AB/S4END[6] Tile_X8Y9_LUT4AB/S4END[7]
+ Tile_X8Y9_LUT4AB/S4END[8] Tile_X8Y9_LUT4AB/S4END[9] Tile_X8Y8_LUT4AB/S4END[0] Tile_X8Y8_LUT4AB/S4END[10]
+ Tile_X8Y8_LUT4AB/S4END[11] Tile_X8Y8_LUT4AB/S4END[12] Tile_X8Y8_LUT4AB/S4END[13]
+ Tile_X8Y8_LUT4AB/S4END[14] Tile_X8Y8_LUT4AB/S4END[15] Tile_X8Y8_LUT4AB/S4END[1]
+ Tile_X8Y8_LUT4AB/S4END[2] Tile_X8Y8_LUT4AB/S4END[3] Tile_X8Y8_LUT4AB/S4END[4] Tile_X8Y8_LUT4AB/S4END[5]
+ Tile_X8Y8_LUT4AB/S4END[6] Tile_X8Y8_LUT4AB/S4END[7] Tile_X8Y8_LUT4AB/S4END[8] Tile_X8Y8_LUT4AB/S4END[9]
+ Tile_X8Y9_LUT4AB/SS4END[0] Tile_X8Y9_LUT4AB/SS4END[10] Tile_X8Y9_LUT4AB/SS4END[11]
+ Tile_X8Y9_LUT4AB/SS4END[12] Tile_X8Y9_LUT4AB/SS4END[13] Tile_X8Y9_LUT4AB/SS4END[14]
+ Tile_X8Y9_LUT4AB/SS4END[15] Tile_X8Y9_LUT4AB/SS4END[1] Tile_X8Y9_LUT4AB/SS4END[2]
+ Tile_X8Y9_LUT4AB/SS4END[3] Tile_X8Y9_LUT4AB/SS4END[4] Tile_X8Y9_LUT4AB/SS4END[5]
+ Tile_X8Y9_LUT4AB/SS4END[6] Tile_X8Y9_LUT4AB/SS4END[7] Tile_X8Y9_LUT4AB/SS4END[8]
+ Tile_X8Y9_LUT4AB/SS4END[9] Tile_X8Y8_LUT4AB/SS4END[0] Tile_X8Y8_LUT4AB/SS4END[10]
+ Tile_X8Y8_LUT4AB/SS4END[11] Tile_X8Y8_LUT4AB/SS4END[12] Tile_X8Y8_LUT4AB/SS4END[13]
+ Tile_X8Y8_LUT4AB/SS4END[14] Tile_X8Y8_LUT4AB/SS4END[15] Tile_X8Y8_LUT4AB/SS4END[1]
+ Tile_X8Y8_LUT4AB/SS4END[2] Tile_X8Y8_LUT4AB/SS4END[3] Tile_X8Y8_LUT4AB/SS4END[4]
+ Tile_X8Y8_LUT4AB/SS4END[5] Tile_X8Y8_LUT4AB/SS4END[6] Tile_X8Y8_LUT4AB/SS4END[7]
+ Tile_X8Y8_LUT4AB/SS4END[8] Tile_X8Y8_LUT4AB/SS4END[9] Tile_X8Y8_LUT4AB/UserCLK Tile_X8Y7_LUT4AB/UserCLK
+ VGND VPWR Tile_X8Y8_LUT4AB/W1BEG[0] Tile_X8Y8_LUT4AB/W1BEG[1] Tile_X8Y8_LUT4AB/W1BEG[2]
+ Tile_X8Y8_LUT4AB/W1BEG[3] Tile_X9Y8_LUT4AB/W1BEG[0] Tile_X9Y8_LUT4AB/W1BEG[1] Tile_X9Y8_LUT4AB/W1BEG[2]
+ Tile_X9Y8_LUT4AB/W1BEG[3] Tile_X8Y8_LUT4AB/W2BEG[0] Tile_X8Y8_LUT4AB/W2BEG[1] Tile_X8Y8_LUT4AB/W2BEG[2]
+ Tile_X8Y8_LUT4AB/W2BEG[3] Tile_X8Y8_LUT4AB/W2BEG[4] Tile_X8Y8_LUT4AB/W2BEG[5] Tile_X8Y8_LUT4AB/W2BEG[6]
+ Tile_X8Y8_LUT4AB/W2BEG[7] Tile_X8Y8_LUT4AB/W2BEGb[0] Tile_X8Y8_LUT4AB/W2BEGb[1]
+ Tile_X8Y8_LUT4AB/W2BEGb[2] Tile_X8Y8_LUT4AB/W2BEGb[3] Tile_X8Y8_LUT4AB/W2BEGb[4]
+ Tile_X8Y8_LUT4AB/W2BEGb[5] Tile_X8Y8_LUT4AB/W2BEGb[6] Tile_X8Y8_LUT4AB/W2BEGb[7]
+ Tile_X8Y8_LUT4AB/W2END[0] Tile_X8Y8_LUT4AB/W2END[1] Tile_X8Y8_LUT4AB/W2END[2] Tile_X8Y8_LUT4AB/W2END[3]
+ Tile_X8Y8_LUT4AB/W2END[4] Tile_X8Y8_LUT4AB/W2END[5] Tile_X8Y8_LUT4AB/W2END[6] Tile_X8Y8_LUT4AB/W2END[7]
+ Tile_X9Y8_LUT4AB/W2BEG[0] Tile_X9Y8_LUT4AB/W2BEG[1] Tile_X9Y8_LUT4AB/W2BEG[2] Tile_X9Y8_LUT4AB/W2BEG[3]
+ Tile_X9Y8_LUT4AB/W2BEG[4] Tile_X9Y8_LUT4AB/W2BEG[5] Tile_X9Y8_LUT4AB/W2BEG[6] Tile_X9Y8_LUT4AB/W2BEG[7]
+ Tile_X8Y8_LUT4AB/W6BEG[0] Tile_X8Y8_LUT4AB/W6BEG[10] Tile_X8Y8_LUT4AB/W6BEG[11]
+ Tile_X8Y8_LUT4AB/W6BEG[1] Tile_X8Y8_LUT4AB/W6BEG[2] Tile_X8Y8_LUT4AB/W6BEG[3] Tile_X8Y8_LUT4AB/W6BEG[4]
+ Tile_X8Y8_LUT4AB/W6BEG[5] Tile_X8Y8_LUT4AB/W6BEG[6] Tile_X8Y8_LUT4AB/W6BEG[7] Tile_X8Y8_LUT4AB/W6BEG[8]
+ Tile_X8Y8_LUT4AB/W6BEG[9] Tile_X9Y8_LUT4AB/W6BEG[0] Tile_X9Y8_LUT4AB/W6BEG[10] Tile_X9Y8_LUT4AB/W6BEG[11]
+ Tile_X9Y8_LUT4AB/W6BEG[1] Tile_X9Y8_LUT4AB/W6BEG[2] Tile_X9Y8_LUT4AB/W6BEG[3] Tile_X9Y8_LUT4AB/W6BEG[4]
+ Tile_X9Y8_LUT4AB/W6BEG[5] Tile_X9Y8_LUT4AB/W6BEG[6] Tile_X9Y8_LUT4AB/W6BEG[7] Tile_X9Y8_LUT4AB/W6BEG[8]
+ Tile_X9Y8_LUT4AB/W6BEG[9] Tile_X8Y8_LUT4AB/WW4BEG[0] Tile_X8Y8_LUT4AB/WW4BEG[10]
+ Tile_X8Y8_LUT4AB/WW4BEG[11] Tile_X8Y8_LUT4AB/WW4BEG[12] Tile_X8Y8_LUT4AB/WW4BEG[13]
+ Tile_X8Y8_LUT4AB/WW4BEG[14] Tile_X8Y8_LUT4AB/WW4BEG[15] Tile_X8Y8_LUT4AB/WW4BEG[1]
+ Tile_X8Y8_LUT4AB/WW4BEG[2] Tile_X8Y8_LUT4AB/WW4BEG[3] Tile_X8Y8_LUT4AB/WW4BEG[4]
+ Tile_X8Y8_LUT4AB/WW4BEG[5] Tile_X8Y8_LUT4AB/WW4BEG[6] Tile_X8Y8_LUT4AB/WW4BEG[7]
+ Tile_X8Y8_LUT4AB/WW4BEG[8] Tile_X8Y8_LUT4AB/WW4BEG[9] Tile_X9Y8_LUT4AB/WW4BEG[0]
+ Tile_X9Y8_LUT4AB/WW4BEG[10] Tile_X9Y8_LUT4AB/WW4BEG[11] Tile_X9Y8_LUT4AB/WW4BEG[12]
+ Tile_X9Y8_LUT4AB/WW4BEG[13] Tile_X9Y8_LUT4AB/WW4BEG[14] Tile_X9Y8_LUT4AB/WW4BEG[15]
+ Tile_X9Y8_LUT4AB/WW4BEG[1] Tile_X9Y8_LUT4AB/WW4BEG[2] Tile_X9Y8_LUT4AB/WW4BEG[3]
+ Tile_X9Y8_LUT4AB/WW4BEG[4] Tile_X9Y8_LUT4AB/WW4BEG[5] Tile_X9Y8_LUT4AB/WW4BEG[6]
+ Tile_X9Y8_LUT4AB/WW4BEG[7] Tile_X9Y8_LUT4AB/WW4BEG[8] Tile_X9Y8_LUT4AB/WW4BEG[9]
+ LUT4AB
XTile_X0Y8_W_IO Tile_X0Y8_A_I_top Tile_X0Y8_A_O_top Tile_X0Y8_A_T_top Tile_X0Y8_A_config_C_bit0
+ Tile_X0Y8_A_config_C_bit1 Tile_X0Y8_A_config_C_bit2 Tile_X0Y8_A_config_C_bit3 Tile_X0Y8_B_I_top
+ Tile_X0Y8_B_O_top Tile_X0Y8_B_T_top Tile_X0Y8_B_config_C_bit0 Tile_X0Y8_B_config_C_bit1
+ Tile_X0Y8_B_config_C_bit2 Tile_X0Y8_B_config_C_bit3 Tile_X0Y8_W_IO/E1BEG[0] Tile_X0Y8_W_IO/E1BEG[1]
+ Tile_X0Y8_W_IO/E1BEG[2] Tile_X0Y8_W_IO/E1BEG[3] Tile_X0Y8_W_IO/E2BEG[0] Tile_X0Y8_W_IO/E2BEG[1]
+ Tile_X0Y8_W_IO/E2BEG[2] Tile_X0Y8_W_IO/E2BEG[3] Tile_X0Y8_W_IO/E2BEG[4] Tile_X0Y8_W_IO/E2BEG[5]
+ Tile_X0Y8_W_IO/E2BEG[6] Tile_X0Y8_W_IO/E2BEG[7] Tile_X0Y8_W_IO/E2BEGb[0] Tile_X0Y8_W_IO/E2BEGb[1]
+ Tile_X0Y8_W_IO/E2BEGb[2] Tile_X0Y8_W_IO/E2BEGb[3] Tile_X0Y8_W_IO/E2BEGb[4] Tile_X0Y8_W_IO/E2BEGb[5]
+ Tile_X0Y8_W_IO/E2BEGb[6] Tile_X0Y8_W_IO/E2BEGb[7] Tile_X0Y8_W_IO/E6BEG[0] Tile_X0Y8_W_IO/E6BEG[10]
+ Tile_X0Y8_W_IO/E6BEG[11] Tile_X0Y8_W_IO/E6BEG[1] Tile_X0Y8_W_IO/E6BEG[2] Tile_X0Y8_W_IO/E6BEG[3]
+ Tile_X0Y8_W_IO/E6BEG[4] Tile_X0Y8_W_IO/E6BEG[5] Tile_X0Y8_W_IO/E6BEG[6] Tile_X0Y8_W_IO/E6BEG[7]
+ Tile_X0Y8_W_IO/E6BEG[8] Tile_X0Y8_W_IO/E6BEG[9] Tile_X0Y8_W_IO/EE4BEG[0] Tile_X0Y8_W_IO/EE4BEG[10]
+ Tile_X0Y8_W_IO/EE4BEG[11] Tile_X0Y8_W_IO/EE4BEG[12] Tile_X0Y8_W_IO/EE4BEG[13] Tile_X0Y8_W_IO/EE4BEG[14]
+ Tile_X0Y8_W_IO/EE4BEG[15] Tile_X0Y8_W_IO/EE4BEG[1] Tile_X0Y8_W_IO/EE4BEG[2] Tile_X0Y8_W_IO/EE4BEG[3]
+ Tile_X0Y8_W_IO/EE4BEG[4] Tile_X0Y8_W_IO/EE4BEG[5] Tile_X0Y8_W_IO/EE4BEG[6] Tile_X0Y8_W_IO/EE4BEG[7]
+ Tile_X0Y8_W_IO/EE4BEG[8] Tile_X0Y8_W_IO/EE4BEG[9] FrameData[256] FrameData[266]
+ FrameData[267] FrameData[268] FrameData[269] FrameData[270] FrameData[271] FrameData[272]
+ FrameData[273] FrameData[274] FrameData[275] FrameData[257] FrameData[276] FrameData[277]
+ FrameData[278] FrameData[279] FrameData[280] FrameData[281] FrameData[282] FrameData[283]
+ FrameData[284] FrameData[285] FrameData[258] FrameData[286] FrameData[287] FrameData[259]
+ FrameData[260] FrameData[261] FrameData[262] FrameData[263] FrameData[264] FrameData[265]
+ Tile_X1Y8_LUT4AB/FrameData[0] Tile_X1Y8_LUT4AB/FrameData[10] Tile_X1Y8_LUT4AB/FrameData[11]
+ Tile_X1Y8_LUT4AB/FrameData[12] Tile_X1Y8_LUT4AB/FrameData[13] Tile_X1Y8_LUT4AB/FrameData[14]
+ Tile_X1Y8_LUT4AB/FrameData[15] Tile_X1Y8_LUT4AB/FrameData[16] Tile_X1Y8_LUT4AB/FrameData[17]
+ Tile_X1Y8_LUT4AB/FrameData[18] Tile_X1Y8_LUT4AB/FrameData[19] Tile_X1Y8_LUT4AB/FrameData[1]
+ Tile_X1Y8_LUT4AB/FrameData[20] Tile_X1Y8_LUT4AB/FrameData[21] Tile_X1Y8_LUT4AB/FrameData[22]
+ Tile_X1Y8_LUT4AB/FrameData[23] Tile_X1Y8_LUT4AB/FrameData[24] Tile_X1Y8_LUT4AB/FrameData[25]
+ Tile_X1Y8_LUT4AB/FrameData[26] Tile_X1Y8_LUT4AB/FrameData[27] Tile_X1Y8_LUT4AB/FrameData[28]
+ Tile_X1Y8_LUT4AB/FrameData[29] Tile_X1Y8_LUT4AB/FrameData[2] Tile_X1Y8_LUT4AB/FrameData[30]
+ Tile_X1Y8_LUT4AB/FrameData[31] Tile_X1Y8_LUT4AB/FrameData[3] Tile_X1Y8_LUT4AB/FrameData[4]
+ Tile_X1Y8_LUT4AB/FrameData[5] Tile_X1Y8_LUT4AB/FrameData[6] Tile_X1Y8_LUT4AB/FrameData[7]
+ Tile_X1Y8_LUT4AB/FrameData[8] Tile_X1Y8_LUT4AB/FrameData[9] Tile_X0Y8_W_IO/FrameStrobe[0]
+ Tile_X0Y8_W_IO/FrameStrobe[10] Tile_X0Y8_W_IO/FrameStrobe[11] Tile_X0Y8_W_IO/FrameStrobe[12]
+ Tile_X0Y8_W_IO/FrameStrobe[13] Tile_X0Y8_W_IO/FrameStrobe[14] Tile_X0Y8_W_IO/FrameStrobe[15]
+ Tile_X0Y8_W_IO/FrameStrobe[16] Tile_X0Y8_W_IO/FrameStrobe[17] Tile_X0Y8_W_IO/FrameStrobe[18]
+ Tile_X0Y8_W_IO/FrameStrobe[19] Tile_X0Y8_W_IO/FrameStrobe[1] Tile_X0Y8_W_IO/FrameStrobe[2]
+ Tile_X0Y8_W_IO/FrameStrobe[3] Tile_X0Y8_W_IO/FrameStrobe[4] Tile_X0Y8_W_IO/FrameStrobe[5]
+ Tile_X0Y8_W_IO/FrameStrobe[6] Tile_X0Y8_W_IO/FrameStrobe[7] Tile_X0Y8_W_IO/FrameStrobe[8]
+ Tile_X0Y8_W_IO/FrameStrobe[9] Tile_X0Y7_W_IO/FrameStrobe[0] Tile_X0Y7_W_IO/FrameStrobe[10]
+ Tile_X0Y7_W_IO/FrameStrobe[11] Tile_X0Y7_W_IO/FrameStrobe[12] Tile_X0Y7_W_IO/FrameStrobe[13]
+ Tile_X0Y7_W_IO/FrameStrobe[14] Tile_X0Y7_W_IO/FrameStrobe[15] Tile_X0Y7_W_IO/FrameStrobe[16]
+ Tile_X0Y7_W_IO/FrameStrobe[17] Tile_X0Y7_W_IO/FrameStrobe[18] Tile_X0Y7_W_IO/FrameStrobe[19]
+ Tile_X0Y7_W_IO/FrameStrobe[1] Tile_X0Y7_W_IO/FrameStrobe[2] Tile_X0Y7_W_IO/FrameStrobe[3]
+ Tile_X0Y7_W_IO/FrameStrobe[4] Tile_X0Y7_W_IO/FrameStrobe[5] Tile_X0Y7_W_IO/FrameStrobe[6]
+ Tile_X0Y7_W_IO/FrameStrobe[7] Tile_X0Y7_W_IO/FrameStrobe[8] Tile_X0Y7_W_IO/FrameStrobe[9]
+ Tile_X0Y8_W_IO/UserCLK Tile_X0Y7_W_IO/UserCLK VGND VPWR Tile_X0Y8_W_IO/W1END[0]
+ Tile_X0Y8_W_IO/W1END[1] Tile_X0Y8_W_IO/W1END[2] Tile_X0Y8_W_IO/W1END[3] Tile_X0Y8_W_IO/W2END[0]
+ Tile_X0Y8_W_IO/W2END[1] Tile_X0Y8_W_IO/W2END[2] Tile_X0Y8_W_IO/W2END[3] Tile_X0Y8_W_IO/W2END[4]
+ Tile_X0Y8_W_IO/W2END[5] Tile_X0Y8_W_IO/W2END[6] Tile_X0Y8_W_IO/W2END[7] Tile_X0Y8_W_IO/W2MID[0]
+ Tile_X0Y8_W_IO/W2MID[1] Tile_X0Y8_W_IO/W2MID[2] Tile_X0Y8_W_IO/W2MID[3] Tile_X0Y8_W_IO/W2MID[4]
+ Tile_X0Y8_W_IO/W2MID[5] Tile_X0Y8_W_IO/W2MID[6] Tile_X0Y8_W_IO/W2MID[7] Tile_X0Y8_W_IO/W6END[0]
+ Tile_X0Y8_W_IO/W6END[10] Tile_X0Y8_W_IO/W6END[11] Tile_X0Y8_W_IO/W6END[1] Tile_X0Y8_W_IO/W6END[2]
+ Tile_X0Y8_W_IO/W6END[3] Tile_X0Y8_W_IO/W6END[4] Tile_X0Y8_W_IO/W6END[5] Tile_X0Y8_W_IO/W6END[6]
+ Tile_X0Y8_W_IO/W6END[7] Tile_X0Y8_W_IO/W6END[8] Tile_X0Y8_W_IO/W6END[9] Tile_X0Y8_W_IO/WW4END[0]
+ Tile_X0Y8_W_IO/WW4END[10] Tile_X0Y8_W_IO/WW4END[11] Tile_X0Y8_W_IO/WW4END[12] Tile_X0Y8_W_IO/WW4END[13]
+ Tile_X0Y8_W_IO/WW4END[14] Tile_X0Y8_W_IO/WW4END[15] Tile_X0Y8_W_IO/WW4END[1] Tile_X0Y8_W_IO/WW4END[2]
+ Tile_X0Y8_W_IO/WW4END[3] Tile_X0Y8_W_IO/WW4END[4] Tile_X0Y8_W_IO/WW4END[5] Tile_X0Y8_W_IO/WW4END[6]
+ Tile_X0Y8_W_IO/WW4END[7] Tile_X0Y8_W_IO/WW4END[8] Tile_X0Y8_W_IO/WW4END[9] W_IO
XTile_X1Y2_LUT4AB Tile_X1Y3_LUT4AB/Co Tile_X1Y2_LUT4AB/Co Tile_X2Y2_LUT4AB/E1END[0]
+ Tile_X2Y2_LUT4AB/E1END[1] Tile_X2Y2_LUT4AB/E1END[2] Tile_X2Y2_LUT4AB/E1END[3] Tile_X0Y2_W_IO/E1BEG[0]
+ Tile_X0Y2_W_IO/E1BEG[1] Tile_X0Y2_W_IO/E1BEG[2] Tile_X0Y2_W_IO/E1BEG[3] Tile_X2Y2_LUT4AB/E2MID[0]
+ Tile_X2Y2_LUT4AB/E2MID[1] Tile_X2Y2_LUT4AB/E2MID[2] Tile_X2Y2_LUT4AB/E2MID[3] Tile_X2Y2_LUT4AB/E2MID[4]
+ Tile_X2Y2_LUT4AB/E2MID[5] Tile_X2Y2_LUT4AB/E2MID[6] Tile_X2Y2_LUT4AB/E2MID[7] Tile_X2Y2_LUT4AB/E2END[0]
+ Tile_X2Y2_LUT4AB/E2END[1] Tile_X2Y2_LUT4AB/E2END[2] Tile_X2Y2_LUT4AB/E2END[3] Tile_X2Y2_LUT4AB/E2END[4]
+ Tile_X2Y2_LUT4AB/E2END[5] Tile_X2Y2_LUT4AB/E2END[6] Tile_X2Y2_LUT4AB/E2END[7] Tile_X0Y2_W_IO/E2BEGb[0]
+ Tile_X0Y2_W_IO/E2BEGb[1] Tile_X0Y2_W_IO/E2BEGb[2] Tile_X0Y2_W_IO/E2BEGb[3] Tile_X0Y2_W_IO/E2BEGb[4]
+ Tile_X0Y2_W_IO/E2BEGb[5] Tile_X0Y2_W_IO/E2BEGb[6] Tile_X0Y2_W_IO/E2BEGb[7] Tile_X0Y2_W_IO/E2BEG[0]
+ Tile_X0Y2_W_IO/E2BEG[1] Tile_X0Y2_W_IO/E2BEG[2] Tile_X0Y2_W_IO/E2BEG[3] Tile_X0Y2_W_IO/E2BEG[4]
+ Tile_X0Y2_W_IO/E2BEG[5] Tile_X0Y2_W_IO/E2BEG[6] Tile_X0Y2_W_IO/E2BEG[7] Tile_X2Y2_LUT4AB/E6END[0]
+ Tile_X2Y2_LUT4AB/E6END[10] Tile_X2Y2_LUT4AB/E6END[11] Tile_X2Y2_LUT4AB/E6END[1]
+ Tile_X2Y2_LUT4AB/E6END[2] Tile_X2Y2_LUT4AB/E6END[3] Tile_X2Y2_LUT4AB/E6END[4] Tile_X2Y2_LUT4AB/E6END[5]
+ Tile_X2Y2_LUT4AB/E6END[6] Tile_X2Y2_LUT4AB/E6END[7] Tile_X2Y2_LUT4AB/E6END[8] Tile_X2Y2_LUT4AB/E6END[9]
+ Tile_X0Y2_W_IO/E6BEG[0] Tile_X0Y2_W_IO/E6BEG[10] Tile_X0Y2_W_IO/E6BEG[11] Tile_X0Y2_W_IO/E6BEG[1]
+ Tile_X0Y2_W_IO/E6BEG[2] Tile_X0Y2_W_IO/E6BEG[3] Tile_X0Y2_W_IO/E6BEG[4] Tile_X0Y2_W_IO/E6BEG[5]
+ Tile_X0Y2_W_IO/E6BEG[6] Tile_X0Y2_W_IO/E6BEG[7] Tile_X0Y2_W_IO/E6BEG[8] Tile_X0Y2_W_IO/E6BEG[9]
+ Tile_X2Y2_LUT4AB/EE4END[0] Tile_X2Y2_LUT4AB/EE4END[10] Tile_X2Y2_LUT4AB/EE4END[11]
+ Tile_X2Y2_LUT4AB/EE4END[12] Tile_X2Y2_LUT4AB/EE4END[13] Tile_X2Y2_LUT4AB/EE4END[14]
+ Tile_X2Y2_LUT4AB/EE4END[15] Tile_X2Y2_LUT4AB/EE4END[1] Tile_X2Y2_LUT4AB/EE4END[2]
+ Tile_X2Y2_LUT4AB/EE4END[3] Tile_X2Y2_LUT4AB/EE4END[4] Tile_X2Y2_LUT4AB/EE4END[5]
+ Tile_X2Y2_LUT4AB/EE4END[6] Tile_X2Y2_LUT4AB/EE4END[7] Tile_X2Y2_LUT4AB/EE4END[8]
+ Tile_X2Y2_LUT4AB/EE4END[9] Tile_X0Y2_W_IO/EE4BEG[0] Tile_X0Y2_W_IO/EE4BEG[10] Tile_X0Y2_W_IO/EE4BEG[11]
+ Tile_X0Y2_W_IO/EE4BEG[12] Tile_X0Y2_W_IO/EE4BEG[13] Tile_X0Y2_W_IO/EE4BEG[14] Tile_X0Y2_W_IO/EE4BEG[15]
+ Tile_X0Y2_W_IO/EE4BEG[1] Tile_X0Y2_W_IO/EE4BEG[2] Tile_X0Y2_W_IO/EE4BEG[3] Tile_X0Y2_W_IO/EE4BEG[4]
+ Tile_X0Y2_W_IO/EE4BEG[5] Tile_X0Y2_W_IO/EE4BEG[6] Tile_X0Y2_W_IO/EE4BEG[7] Tile_X0Y2_W_IO/EE4BEG[8]
+ Tile_X0Y2_W_IO/EE4BEG[9] Tile_X1Y2_LUT4AB/FrameData[0] Tile_X1Y2_LUT4AB/FrameData[10]
+ Tile_X1Y2_LUT4AB/FrameData[11] Tile_X1Y2_LUT4AB/FrameData[12] Tile_X1Y2_LUT4AB/FrameData[13]
+ Tile_X1Y2_LUT4AB/FrameData[14] Tile_X1Y2_LUT4AB/FrameData[15] Tile_X1Y2_LUT4AB/FrameData[16]
+ Tile_X1Y2_LUT4AB/FrameData[17] Tile_X1Y2_LUT4AB/FrameData[18] Tile_X1Y2_LUT4AB/FrameData[19]
+ Tile_X1Y2_LUT4AB/FrameData[1] Tile_X1Y2_LUT4AB/FrameData[20] Tile_X1Y2_LUT4AB/FrameData[21]
+ Tile_X1Y2_LUT4AB/FrameData[22] Tile_X1Y2_LUT4AB/FrameData[23] Tile_X1Y2_LUT4AB/FrameData[24]
+ Tile_X1Y2_LUT4AB/FrameData[25] Tile_X1Y2_LUT4AB/FrameData[26] Tile_X1Y2_LUT4AB/FrameData[27]
+ Tile_X1Y2_LUT4AB/FrameData[28] Tile_X1Y2_LUT4AB/FrameData[29] Tile_X1Y2_LUT4AB/FrameData[2]
+ Tile_X1Y2_LUT4AB/FrameData[30] Tile_X1Y2_LUT4AB/FrameData[31] Tile_X1Y2_LUT4AB/FrameData[3]
+ Tile_X1Y2_LUT4AB/FrameData[4] Tile_X1Y2_LUT4AB/FrameData[5] Tile_X1Y2_LUT4AB/FrameData[6]
+ Tile_X1Y2_LUT4AB/FrameData[7] Tile_X1Y2_LUT4AB/FrameData[8] Tile_X1Y2_LUT4AB/FrameData[9]
+ Tile_X2Y2_LUT4AB/FrameData[0] Tile_X2Y2_LUT4AB/FrameData[10] Tile_X2Y2_LUT4AB/FrameData[11]
+ Tile_X2Y2_LUT4AB/FrameData[12] Tile_X2Y2_LUT4AB/FrameData[13] Tile_X2Y2_LUT4AB/FrameData[14]
+ Tile_X2Y2_LUT4AB/FrameData[15] Tile_X2Y2_LUT4AB/FrameData[16] Tile_X2Y2_LUT4AB/FrameData[17]
+ Tile_X2Y2_LUT4AB/FrameData[18] Tile_X2Y2_LUT4AB/FrameData[19] Tile_X2Y2_LUT4AB/FrameData[1]
+ Tile_X2Y2_LUT4AB/FrameData[20] Tile_X2Y2_LUT4AB/FrameData[21] Tile_X2Y2_LUT4AB/FrameData[22]
+ Tile_X2Y2_LUT4AB/FrameData[23] Tile_X2Y2_LUT4AB/FrameData[24] Tile_X2Y2_LUT4AB/FrameData[25]
+ Tile_X2Y2_LUT4AB/FrameData[26] Tile_X2Y2_LUT4AB/FrameData[27] Tile_X2Y2_LUT4AB/FrameData[28]
+ Tile_X2Y2_LUT4AB/FrameData[29] Tile_X2Y2_LUT4AB/FrameData[2] Tile_X2Y2_LUT4AB/FrameData[30]
+ Tile_X2Y2_LUT4AB/FrameData[31] Tile_X2Y2_LUT4AB/FrameData[3] Tile_X2Y2_LUT4AB/FrameData[4]
+ Tile_X2Y2_LUT4AB/FrameData[5] Tile_X2Y2_LUT4AB/FrameData[6] Tile_X2Y2_LUT4AB/FrameData[7]
+ Tile_X2Y2_LUT4AB/FrameData[8] Tile_X2Y2_LUT4AB/FrameData[9] Tile_X1Y2_LUT4AB/FrameStrobe[0]
+ Tile_X1Y2_LUT4AB/FrameStrobe[10] Tile_X1Y2_LUT4AB/FrameStrobe[11] Tile_X1Y2_LUT4AB/FrameStrobe[12]
+ Tile_X1Y2_LUT4AB/FrameStrobe[13] Tile_X1Y2_LUT4AB/FrameStrobe[14] Tile_X1Y2_LUT4AB/FrameStrobe[15]
+ Tile_X1Y2_LUT4AB/FrameStrobe[16] Tile_X1Y2_LUT4AB/FrameStrobe[17] Tile_X1Y2_LUT4AB/FrameStrobe[18]
+ Tile_X1Y2_LUT4AB/FrameStrobe[19] Tile_X1Y2_LUT4AB/FrameStrobe[1] Tile_X1Y2_LUT4AB/FrameStrobe[2]
+ Tile_X1Y2_LUT4AB/FrameStrobe[3] Tile_X1Y2_LUT4AB/FrameStrobe[4] Tile_X1Y2_LUT4AB/FrameStrobe[5]
+ Tile_X1Y2_LUT4AB/FrameStrobe[6] Tile_X1Y2_LUT4AB/FrameStrobe[7] Tile_X1Y2_LUT4AB/FrameStrobe[8]
+ Tile_X1Y2_LUT4AB/FrameStrobe[9] Tile_X1Y1_LUT4AB/FrameStrobe[0] Tile_X1Y1_LUT4AB/FrameStrobe[10]
+ Tile_X1Y1_LUT4AB/FrameStrobe[11] Tile_X1Y1_LUT4AB/FrameStrobe[12] Tile_X1Y1_LUT4AB/FrameStrobe[13]
+ Tile_X1Y1_LUT4AB/FrameStrobe[14] Tile_X1Y1_LUT4AB/FrameStrobe[15] Tile_X1Y1_LUT4AB/FrameStrobe[16]
+ Tile_X1Y1_LUT4AB/FrameStrobe[17] Tile_X1Y1_LUT4AB/FrameStrobe[18] Tile_X1Y1_LUT4AB/FrameStrobe[19]
+ Tile_X1Y1_LUT4AB/FrameStrobe[1] Tile_X1Y1_LUT4AB/FrameStrobe[2] Tile_X1Y1_LUT4AB/FrameStrobe[3]
+ Tile_X1Y1_LUT4AB/FrameStrobe[4] Tile_X1Y1_LUT4AB/FrameStrobe[5] Tile_X1Y1_LUT4AB/FrameStrobe[6]
+ Tile_X1Y1_LUT4AB/FrameStrobe[7] Tile_X1Y1_LUT4AB/FrameStrobe[8] Tile_X1Y1_LUT4AB/FrameStrobe[9]
+ Tile_X1Y2_LUT4AB/N1BEG[0] Tile_X1Y2_LUT4AB/N1BEG[1] Tile_X1Y2_LUT4AB/N1BEG[2] Tile_X1Y2_LUT4AB/N1BEG[3]
+ Tile_X1Y3_LUT4AB/N1BEG[0] Tile_X1Y3_LUT4AB/N1BEG[1] Tile_X1Y3_LUT4AB/N1BEG[2] Tile_X1Y3_LUT4AB/N1BEG[3]
+ Tile_X1Y2_LUT4AB/N2BEG[0] Tile_X1Y2_LUT4AB/N2BEG[1] Tile_X1Y2_LUT4AB/N2BEG[2] Tile_X1Y2_LUT4AB/N2BEG[3]
+ Tile_X1Y2_LUT4AB/N2BEG[4] Tile_X1Y2_LUT4AB/N2BEG[5] Tile_X1Y2_LUT4AB/N2BEG[6] Tile_X1Y2_LUT4AB/N2BEG[7]
+ Tile_X1Y1_LUT4AB/N2END[0] Tile_X1Y1_LUT4AB/N2END[1] Tile_X1Y1_LUT4AB/N2END[2] Tile_X1Y1_LUT4AB/N2END[3]
+ Tile_X1Y1_LUT4AB/N2END[4] Tile_X1Y1_LUT4AB/N2END[5] Tile_X1Y1_LUT4AB/N2END[6] Tile_X1Y1_LUT4AB/N2END[7]
+ Tile_X1Y2_LUT4AB/N2END[0] Tile_X1Y2_LUT4AB/N2END[1] Tile_X1Y2_LUT4AB/N2END[2] Tile_X1Y2_LUT4AB/N2END[3]
+ Tile_X1Y2_LUT4AB/N2END[4] Tile_X1Y2_LUT4AB/N2END[5] Tile_X1Y2_LUT4AB/N2END[6] Tile_X1Y2_LUT4AB/N2END[7]
+ Tile_X1Y3_LUT4AB/N2BEG[0] Tile_X1Y3_LUT4AB/N2BEG[1] Tile_X1Y3_LUT4AB/N2BEG[2] Tile_X1Y3_LUT4AB/N2BEG[3]
+ Tile_X1Y3_LUT4AB/N2BEG[4] Tile_X1Y3_LUT4AB/N2BEG[5] Tile_X1Y3_LUT4AB/N2BEG[6] Tile_X1Y3_LUT4AB/N2BEG[7]
+ Tile_X1Y2_LUT4AB/N4BEG[0] Tile_X1Y2_LUT4AB/N4BEG[10] Tile_X1Y2_LUT4AB/N4BEG[11]
+ Tile_X1Y2_LUT4AB/N4BEG[12] Tile_X1Y2_LUT4AB/N4BEG[13] Tile_X1Y2_LUT4AB/N4BEG[14]
+ Tile_X1Y2_LUT4AB/N4BEG[15] Tile_X1Y2_LUT4AB/N4BEG[1] Tile_X1Y2_LUT4AB/N4BEG[2] Tile_X1Y2_LUT4AB/N4BEG[3]
+ Tile_X1Y2_LUT4AB/N4BEG[4] Tile_X1Y2_LUT4AB/N4BEG[5] Tile_X1Y2_LUT4AB/N4BEG[6] Tile_X1Y2_LUT4AB/N4BEG[7]
+ Tile_X1Y2_LUT4AB/N4BEG[8] Tile_X1Y2_LUT4AB/N4BEG[9] Tile_X1Y3_LUT4AB/N4BEG[0] Tile_X1Y3_LUT4AB/N4BEG[10]
+ Tile_X1Y3_LUT4AB/N4BEG[11] Tile_X1Y3_LUT4AB/N4BEG[12] Tile_X1Y3_LUT4AB/N4BEG[13]
+ Tile_X1Y3_LUT4AB/N4BEG[14] Tile_X1Y3_LUT4AB/N4BEG[15] Tile_X1Y3_LUT4AB/N4BEG[1]
+ Tile_X1Y3_LUT4AB/N4BEG[2] Tile_X1Y3_LUT4AB/N4BEG[3] Tile_X1Y3_LUT4AB/N4BEG[4] Tile_X1Y3_LUT4AB/N4BEG[5]
+ Tile_X1Y3_LUT4AB/N4BEG[6] Tile_X1Y3_LUT4AB/N4BEG[7] Tile_X1Y3_LUT4AB/N4BEG[8] Tile_X1Y3_LUT4AB/N4BEG[9]
+ Tile_X1Y2_LUT4AB/NN4BEG[0] Tile_X1Y2_LUT4AB/NN4BEG[10] Tile_X1Y2_LUT4AB/NN4BEG[11]
+ Tile_X1Y2_LUT4AB/NN4BEG[12] Tile_X1Y2_LUT4AB/NN4BEG[13] Tile_X1Y2_LUT4AB/NN4BEG[14]
+ Tile_X1Y2_LUT4AB/NN4BEG[15] Tile_X1Y2_LUT4AB/NN4BEG[1] Tile_X1Y2_LUT4AB/NN4BEG[2]
+ Tile_X1Y2_LUT4AB/NN4BEG[3] Tile_X1Y2_LUT4AB/NN4BEG[4] Tile_X1Y2_LUT4AB/NN4BEG[5]
+ Tile_X1Y2_LUT4AB/NN4BEG[6] Tile_X1Y2_LUT4AB/NN4BEG[7] Tile_X1Y2_LUT4AB/NN4BEG[8]
+ Tile_X1Y2_LUT4AB/NN4BEG[9] Tile_X1Y3_LUT4AB/NN4BEG[0] Tile_X1Y3_LUT4AB/NN4BEG[10]
+ Tile_X1Y3_LUT4AB/NN4BEG[11] Tile_X1Y3_LUT4AB/NN4BEG[12] Tile_X1Y3_LUT4AB/NN4BEG[13]
+ Tile_X1Y3_LUT4AB/NN4BEG[14] Tile_X1Y3_LUT4AB/NN4BEG[15] Tile_X1Y3_LUT4AB/NN4BEG[1]
+ Tile_X1Y3_LUT4AB/NN4BEG[2] Tile_X1Y3_LUT4AB/NN4BEG[3] Tile_X1Y3_LUT4AB/NN4BEG[4]
+ Tile_X1Y3_LUT4AB/NN4BEG[5] Tile_X1Y3_LUT4AB/NN4BEG[6] Tile_X1Y3_LUT4AB/NN4BEG[7]
+ Tile_X1Y3_LUT4AB/NN4BEG[8] Tile_X1Y3_LUT4AB/NN4BEG[9] Tile_X1Y3_LUT4AB/S1END[0]
+ Tile_X1Y3_LUT4AB/S1END[1] Tile_X1Y3_LUT4AB/S1END[2] Tile_X1Y3_LUT4AB/S1END[3] Tile_X1Y2_LUT4AB/S1END[0]
+ Tile_X1Y2_LUT4AB/S1END[1] Tile_X1Y2_LUT4AB/S1END[2] Tile_X1Y2_LUT4AB/S1END[3] Tile_X1Y3_LUT4AB/S2MID[0]
+ Tile_X1Y3_LUT4AB/S2MID[1] Tile_X1Y3_LUT4AB/S2MID[2] Tile_X1Y3_LUT4AB/S2MID[3] Tile_X1Y3_LUT4AB/S2MID[4]
+ Tile_X1Y3_LUT4AB/S2MID[5] Tile_X1Y3_LUT4AB/S2MID[6] Tile_X1Y3_LUT4AB/S2MID[7] Tile_X1Y3_LUT4AB/S2END[0]
+ Tile_X1Y3_LUT4AB/S2END[1] Tile_X1Y3_LUT4AB/S2END[2] Tile_X1Y3_LUT4AB/S2END[3] Tile_X1Y3_LUT4AB/S2END[4]
+ Tile_X1Y3_LUT4AB/S2END[5] Tile_X1Y3_LUT4AB/S2END[6] Tile_X1Y3_LUT4AB/S2END[7] Tile_X1Y2_LUT4AB/S2END[0]
+ Tile_X1Y2_LUT4AB/S2END[1] Tile_X1Y2_LUT4AB/S2END[2] Tile_X1Y2_LUT4AB/S2END[3] Tile_X1Y2_LUT4AB/S2END[4]
+ Tile_X1Y2_LUT4AB/S2END[5] Tile_X1Y2_LUT4AB/S2END[6] Tile_X1Y2_LUT4AB/S2END[7] Tile_X1Y2_LUT4AB/S2MID[0]
+ Tile_X1Y2_LUT4AB/S2MID[1] Tile_X1Y2_LUT4AB/S2MID[2] Tile_X1Y2_LUT4AB/S2MID[3] Tile_X1Y2_LUT4AB/S2MID[4]
+ Tile_X1Y2_LUT4AB/S2MID[5] Tile_X1Y2_LUT4AB/S2MID[6] Tile_X1Y2_LUT4AB/S2MID[7] Tile_X1Y3_LUT4AB/S4END[0]
+ Tile_X1Y3_LUT4AB/S4END[10] Tile_X1Y3_LUT4AB/S4END[11] Tile_X1Y3_LUT4AB/S4END[12]
+ Tile_X1Y3_LUT4AB/S4END[13] Tile_X1Y3_LUT4AB/S4END[14] Tile_X1Y3_LUT4AB/S4END[15]
+ Tile_X1Y3_LUT4AB/S4END[1] Tile_X1Y3_LUT4AB/S4END[2] Tile_X1Y3_LUT4AB/S4END[3] Tile_X1Y3_LUT4AB/S4END[4]
+ Tile_X1Y3_LUT4AB/S4END[5] Tile_X1Y3_LUT4AB/S4END[6] Tile_X1Y3_LUT4AB/S4END[7] Tile_X1Y3_LUT4AB/S4END[8]
+ Tile_X1Y3_LUT4AB/S4END[9] Tile_X1Y2_LUT4AB/S4END[0] Tile_X1Y2_LUT4AB/S4END[10] Tile_X1Y2_LUT4AB/S4END[11]
+ Tile_X1Y2_LUT4AB/S4END[12] Tile_X1Y2_LUT4AB/S4END[13] Tile_X1Y2_LUT4AB/S4END[14]
+ Tile_X1Y2_LUT4AB/S4END[15] Tile_X1Y2_LUT4AB/S4END[1] Tile_X1Y2_LUT4AB/S4END[2] Tile_X1Y2_LUT4AB/S4END[3]
+ Tile_X1Y2_LUT4AB/S4END[4] Tile_X1Y2_LUT4AB/S4END[5] Tile_X1Y2_LUT4AB/S4END[6] Tile_X1Y2_LUT4AB/S4END[7]
+ Tile_X1Y2_LUT4AB/S4END[8] Tile_X1Y2_LUT4AB/S4END[9] Tile_X1Y3_LUT4AB/SS4END[0] Tile_X1Y3_LUT4AB/SS4END[10]
+ Tile_X1Y3_LUT4AB/SS4END[11] Tile_X1Y3_LUT4AB/SS4END[12] Tile_X1Y3_LUT4AB/SS4END[13]
+ Tile_X1Y3_LUT4AB/SS4END[14] Tile_X1Y3_LUT4AB/SS4END[15] Tile_X1Y3_LUT4AB/SS4END[1]
+ Tile_X1Y3_LUT4AB/SS4END[2] Tile_X1Y3_LUT4AB/SS4END[3] Tile_X1Y3_LUT4AB/SS4END[4]
+ Tile_X1Y3_LUT4AB/SS4END[5] Tile_X1Y3_LUT4AB/SS4END[6] Tile_X1Y3_LUT4AB/SS4END[7]
+ Tile_X1Y3_LUT4AB/SS4END[8] Tile_X1Y3_LUT4AB/SS4END[9] Tile_X1Y2_LUT4AB/SS4END[0]
+ Tile_X1Y2_LUT4AB/SS4END[10] Tile_X1Y2_LUT4AB/SS4END[11] Tile_X1Y2_LUT4AB/SS4END[12]
+ Tile_X1Y2_LUT4AB/SS4END[13] Tile_X1Y2_LUT4AB/SS4END[14] Tile_X1Y2_LUT4AB/SS4END[15]
+ Tile_X1Y2_LUT4AB/SS4END[1] Tile_X1Y2_LUT4AB/SS4END[2] Tile_X1Y2_LUT4AB/SS4END[3]
+ Tile_X1Y2_LUT4AB/SS4END[4] Tile_X1Y2_LUT4AB/SS4END[5] Tile_X1Y2_LUT4AB/SS4END[6]
+ Tile_X1Y2_LUT4AB/SS4END[7] Tile_X1Y2_LUT4AB/SS4END[8] Tile_X1Y2_LUT4AB/SS4END[9]
+ Tile_X1Y2_LUT4AB/UserCLK Tile_X1Y1_LUT4AB/UserCLK VGND VPWR Tile_X0Y2_W_IO/W1END[0]
+ Tile_X0Y2_W_IO/W1END[1] Tile_X0Y2_W_IO/W1END[2] Tile_X0Y2_W_IO/W1END[3] Tile_X2Y2_LUT4AB/W1BEG[0]
+ Tile_X2Y2_LUT4AB/W1BEG[1] Tile_X2Y2_LUT4AB/W1BEG[2] Tile_X2Y2_LUT4AB/W1BEG[3] Tile_X0Y2_W_IO/W2MID[0]
+ Tile_X0Y2_W_IO/W2MID[1] Tile_X0Y2_W_IO/W2MID[2] Tile_X0Y2_W_IO/W2MID[3] Tile_X0Y2_W_IO/W2MID[4]
+ Tile_X0Y2_W_IO/W2MID[5] Tile_X0Y2_W_IO/W2MID[6] Tile_X0Y2_W_IO/W2MID[7] Tile_X0Y2_W_IO/W2END[0]
+ Tile_X0Y2_W_IO/W2END[1] Tile_X0Y2_W_IO/W2END[2] Tile_X0Y2_W_IO/W2END[3] Tile_X0Y2_W_IO/W2END[4]
+ Tile_X0Y2_W_IO/W2END[5] Tile_X0Y2_W_IO/W2END[6] Tile_X0Y2_W_IO/W2END[7] Tile_X1Y2_LUT4AB/W2END[0]
+ Tile_X1Y2_LUT4AB/W2END[1] Tile_X1Y2_LUT4AB/W2END[2] Tile_X1Y2_LUT4AB/W2END[3] Tile_X1Y2_LUT4AB/W2END[4]
+ Tile_X1Y2_LUT4AB/W2END[5] Tile_X1Y2_LUT4AB/W2END[6] Tile_X1Y2_LUT4AB/W2END[7] Tile_X2Y2_LUT4AB/W2BEG[0]
+ Tile_X2Y2_LUT4AB/W2BEG[1] Tile_X2Y2_LUT4AB/W2BEG[2] Tile_X2Y2_LUT4AB/W2BEG[3] Tile_X2Y2_LUT4AB/W2BEG[4]
+ Tile_X2Y2_LUT4AB/W2BEG[5] Tile_X2Y2_LUT4AB/W2BEG[6] Tile_X2Y2_LUT4AB/W2BEG[7] Tile_X0Y2_W_IO/W6END[0]
+ Tile_X0Y2_W_IO/W6END[10] Tile_X0Y2_W_IO/W6END[11] Tile_X0Y2_W_IO/W6END[1] Tile_X0Y2_W_IO/W6END[2]
+ Tile_X0Y2_W_IO/W6END[3] Tile_X0Y2_W_IO/W6END[4] Tile_X0Y2_W_IO/W6END[5] Tile_X0Y2_W_IO/W6END[6]
+ Tile_X0Y2_W_IO/W6END[7] Tile_X0Y2_W_IO/W6END[8] Tile_X0Y2_W_IO/W6END[9] Tile_X2Y2_LUT4AB/W6BEG[0]
+ Tile_X2Y2_LUT4AB/W6BEG[10] Tile_X2Y2_LUT4AB/W6BEG[11] Tile_X2Y2_LUT4AB/W6BEG[1]
+ Tile_X2Y2_LUT4AB/W6BEG[2] Tile_X2Y2_LUT4AB/W6BEG[3] Tile_X2Y2_LUT4AB/W6BEG[4] Tile_X2Y2_LUT4AB/W6BEG[5]
+ Tile_X2Y2_LUT4AB/W6BEG[6] Tile_X2Y2_LUT4AB/W6BEG[7] Tile_X2Y2_LUT4AB/W6BEG[8] Tile_X2Y2_LUT4AB/W6BEG[9]
+ Tile_X0Y2_W_IO/WW4END[0] Tile_X0Y2_W_IO/WW4END[10] Tile_X0Y2_W_IO/WW4END[11] Tile_X0Y2_W_IO/WW4END[12]
+ Tile_X0Y2_W_IO/WW4END[13] Tile_X0Y2_W_IO/WW4END[14] Tile_X0Y2_W_IO/WW4END[15] Tile_X0Y2_W_IO/WW4END[1]
+ Tile_X0Y2_W_IO/WW4END[2] Tile_X0Y2_W_IO/WW4END[3] Tile_X0Y2_W_IO/WW4END[4] Tile_X0Y2_W_IO/WW4END[5]
+ Tile_X0Y2_W_IO/WW4END[6] Tile_X0Y2_W_IO/WW4END[7] Tile_X0Y2_W_IO/WW4END[8] Tile_X0Y2_W_IO/WW4END[9]
+ Tile_X2Y2_LUT4AB/WW4BEG[0] Tile_X2Y2_LUT4AB/WW4BEG[10] Tile_X2Y2_LUT4AB/WW4BEG[11]
+ Tile_X2Y2_LUT4AB/WW4BEG[12] Tile_X2Y2_LUT4AB/WW4BEG[13] Tile_X2Y2_LUT4AB/WW4BEG[14]
+ Tile_X2Y2_LUT4AB/WW4BEG[15] Tile_X2Y2_LUT4AB/WW4BEG[1] Tile_X2Y2_LUT4AB/WW4BEG[2]
+ Tile_X2Y2_LUT4AB/WW4BEG[3] Tile_X2Y2_LUT4AB/WW4BEG[4] Tile_X2Y2_LUT4AB/WW4BEG[5]
+ Tile_X2Y2_LUT4AB/WW4BEG[6] Tile_X2Y2_LUT4AB/WW4BEG[7] Tile_X2Y2_LUT4AB/WW4BEG[8]
+ Tile_X2Y2_LUT4AB/WW4BEG[9] LUT4AB
XTile_X6Y11_LUT4AB Tile_X6Y12_LUT4AB/Co Tile_X6Y11_LUT4AB/Co Tile_X6Y11_LUT4AB/E1BEG[0]
+ Tile_X6Y11_LUT4AB/E1BEG[1] Tile_X6Y11_LUT4AB/E1BEG[2] Tile_X6Y11_LUT4AB/E1BEG[3]
+ Tile_X6Y11_LUT4AB/E1END[0] Tile_X6Y11_LUT4AB/E1END[1] Tile_X6Y11_LUT4AB/E1END[2]
+ Tile_X6Y11_LUT4AB/E1END[3] Tile_X6Y11_LUT4AB/E2BEG[0] Tile_X6Y11_LUT4AB/E2BEG[1]
+ Tile_X6Y11_LUT4AB/E2BEG[2] Tile_X6Y11_LUT4AB/E2BEG[3] Tile_X6Y11_LUT4AB/E2BEG[4]
+ Tile_X6Y11_LUT4AB/E2BEG[5] Tile_X6Y11_LUT4AB/E2BEG[6] Tile_X6Y11_LUT4AB/E2BEG[7]
+ Tile_X6Y11_LUT4AB/E2BEGb[0] Tile_X6Y11_LUT4AB/E2BEGb[1] Tile_X6Y11_LUT4AB/E2BEGb[2]
+ Tile_X6Y11_LUT4AB/E2BEGb[3] Tile_X6Y11_LUT4AB/E2BEGb[4] Tile_X6Y11_LUT4AB/E2BEGb[5]
+ Tile_X6Y11_LUT4AB/E2BEGb[6] Tile_X6Y11_LUT4AB/E2BEGb[7] Tile_X6Y11_LUT4AB/E2END[0]
+ Tile_X6Y11_LUT4AB/E2END[1] Tile_X6Y11_LUT4AB/E2END[2] Tile_X6Y11_LUT4AB/E2END[3]
+ Tile_X6Y11_LUT4AB/E2END[4] Tile_X6Y11_LUT4AB/E2END[5] Tile_X6Y11_LUT4AB/E2END[6]
+ Tile_X6Y11_LUT4AB/E2END[7] Tile_X6Y11_LUT4AB/E2MID[0] Tile_X6Y11_LUT4AB/E2MID[1]
+ Tile_X6Y11_LUT4AB/E2MID[2] Tile_X6Y11_LUT4AB/E2MID[3] Tile_X6Y11_LUT4AB/E2MID[4]
+ Tile_X6Y11_LUT4AB/E2MID[5] Tile_X6Y11_LUT4AB/E2MID[6] Tile_X6Y11_LUT4AB/E2MID[7]
+ Tile_X6Y11_LUT4AB/E6BEG[0] Tile_X6Y11_LUT4AB/E6BEG[10] Tile_X6Y11_LUT4AB/E6BEG[11]
+ Tile_X6Y11_LUT4AB/E6BEG[1] Tile_X6Y11_LUT4AB/E6BEG[2] Tile_X6Y11_LUT4AB/E6BEG[3]
+ Tile_X6Y11_LUT4AB/E6BEG[4] Tile_X6Y11_LUT4AB/E6BEG[5] Tile_X6Y11_LUT4AB/E6BEG[6]
+ Tile_X6Y11_LUT4AB/E6BEG[7] Tile_X6Y11_LUT4AB/E6BEG[8] Tile_X6Y11_LUT4AB/E6BEG[9]
+ Tile_X6Y11_LUT4AB/E6END[0] Tile_X6Y11_LUT4AB/E6END[10] Tile_X6Y11_LUT4AB/E6END[11]
+ Tile_X6Y11_LUT4AB/E6END[1] Tile_X6Y11_LUT4AB/E6END[2] Tile_X6Y11_LUT4AB/E6END[3]
+ Tile_X6Y11_LUT4AB/E6END[4] Tile_X6Y11_LUT4AB/E6END[5] Tile_X6Y11_LUT4AB/E6END[6]
+ Tile_X6Y11_LUT4AB/E6END[7] Tile_X6Y11_LUT4AB/E6END[8] Tile_X6Y11_LUT4AB/E6END[9]
+ Tile_X6Y11_LUT4AB/EE4BEG[0] Tile_X6Y11_LUT4AB/EE4BEG[10] Tile_X6Y11_LUT4AB/EE4BEG[11]
+ Tile_X6Y11_LUT4AB/EE4BEG[12] Tile_X6Y11_LUT4AB/EE4BEG[13] Tile_X6Y11_LUT4AB/EE4BEG[14]
+ Tile_X6Y11_LUT4AB/EE4BEG[15] Tile_X6Y11_LUT4AB/EE4BEG[1] Tile_X6Y11_LUT4AB/EE4BEG[2]
+ Tile_X6Y11_LUT4AB/EE4BEG[3] Tile_X6Y11_LUT4AB/EE4BEG[4] Tile_X6Y11_LUT4AB/EE4BEG[5]
+ Tile_X6Y11_LUT4AB/EE4BEG[6] Tile_X6Y11_LUT4AB/EE4BEG[7] Tile_X6Y11_LUT4AB/EE4BEG[8]
+ Tile_X6Y11_LUT4AB/EE4BEG[9] Tile_X6Y11_LUT4AB/EE4END[0] Tile_X6Y11_LUT4AB/EE4END[10]
+ Tile_X6Y11_LUT4AB/EE4END[11] Tile_X6Y11_LUT4AB/EE4END[12] Tile_X6Y11_LUT4AB/EE4END[13]
+ Tile_X6Y11_LUT4AB/EE4END[14] Tile_X6Y11_LUT4AB/EE4END[15] Tile_X6Y11_LUT4AB/EE4END[1]
+ Tile_X6Y11_LUT4AB/EE4END[2] Tile_X6Y11_LUT4AB/EE4END[3] Tile_X6Y11_LUT4AB/EE4END[4]
+ Tile_X6Y11_LUT4AB/EE4END[5] Tile_X6Y11_LUT4AB/EE4END[6] Tile_X6Y11_LUT4AB/EE4END[7]
+ Tile_X6Y11_LUT4AB/EE4END[8] Tile_X6Y11_LUT4AB/EE4END[9] Tile_X6Y11_LUT4AB/FrameData[0]
+ Tile_X6Y11_LUT4AB/FrameData[10] Tile_X6Y11_LUT4AB/FrameData[11] Tile_X6Y11_LUT4AB/FrameData[12]
+ Tile_X6Y11_LUT4AB/FrameData[13] Tile_X6Y11_LUT4AB/FrameData[14] Tile_X6Y11_LUT4AB/FrameData[15]
+ Tile_X6Y11_LUT4AB/FrameData[16] Tile_X6Y11_LUT4AB/FrameData[17] Tile_X6Y11_LUT4AB/FrameData[18]
+ Tile_X6Y11_LUT4AB/FrameData[19] Tile_X6Y11_LUT4AB/FrameData[1] Tile_X6Y11_LUT4AB/FrameData[20]
+ Tile_X6Y11_LUT4AB/FrameData[21] Tile_X6Y11_LUT4AB/FrameData[22] Tile_X6Y11_LUT4AB/FrameData[23]
+ Tile_X6Y11_LUT4AB/FrameData[24] Tile_X6Y11_LUT4AB/FrameData[25] Tile_X6Y11_LUT4AB/FrameData[26]
+ Tile_X6Y11_LUT4AB/FrameData[27] Tile_X6Y11_LUT4AB/FrameData[28] Tile_X6Y11_LUT4AB/FrameData[29]
+ Tile_X6Y11_LUT4AB/FrameData[2] Tile_X6Y11_LUT4AB/FrameData[30] Tile_X6Y11_LUT4AB/FrameData[31]
+ Tile_X6Y11_LUT4AB/FrameData[3] Tile_X6Y11_LUT4AB/FrameData[4] Tile_X6Y11_LUT4AB/FrameData[5]
+ Tile_X6Y11_LUT4AB/FrameData[6] Tile_X6Y11_LUT4AB/FrameData[7] Tile_X6Y11_LUT4AB/FrameData[8]
+ Tile_X6Y11_LUT4AB/FrameData[9] Tile_X6Y11_LUT4AB/FrameData_O[0] Tile_X6Y11_LUT4AB/FrameData_O[10]
+ Tile_X6Y11_LUT4AB/FrameData_O[11] Tile_X6Y11_LUT4AB/FrameData_O[12] Tile_X6Y11_LUT4AB/FrameData_O[13]
+ Tile_X6Y11_LUT4AB/FrameData_O[14] Tile_X6Y11_LUT4AB/FrameData_O[15] Tile_X6Y11_LUT4AB/FrameData_O[16]
+ Tile_X6Y11_LUT4AB/FrameData_O[17] Tile_X6Y11_LUT4AB/FrameData_O[18] Tile_X6Y11_LUT4AB/FrameData_O[19]
+ Tile_X6Y11_LUT4AB/FrameData_O[1] Tile_X6Y11_LUT4AB/FrameData_O[20] Tile_X6Y11_LUT4AB/FrameData_O[21]
+ Tile_X6Y11_LUT4AB/FrameData_O[22] Tile_X6Y11_LUT4AB/FrameData_O[23] Tile_X6Y11_LUT4AB/FrameData_O[24]
+ Tile_X6Y11_LUT4AB/FrameData_O[25] Tile_X6Y11_LUT4AB/FrameData_O[26] Tile_X6Y11_LUT4AB/FrameData_O[27]
+ Tile_X6Y11_LUT4AB/FrameData_O[28] Tile_X6Y11_LUT4AB/FrameData_O[29] Tile_X6Y11_LUT4AB/FrameData_O[2]
+ Tile_X6Y11_LUT4AB/FrameData_O[30] Tile_X6Y11_LUT4AB/FrameData_O[31] Tile_X6Y11_LUT4AB/FrameData_O[3]
+ Tile_X6Y11_LUT4AB/FrameData_O[4] Tile_X6Y11_LUT4AB/FrameData_O[5] Tile_X6Y11_LUT4AB/FrameData_O[6]
+ Tile_X6Y11_LUT4AB/FrameData_O[7] Tile_X6Y11_LUT4AB/FrameData_O[8] Tile_X6Y11_LUT4AB/FrameData_O[9]
+ Tile_X6Y11_LUT4AB/FrameStrobe[0] Tile_X6Y11_LUT4AB/FrameStrobe[10] Tile_X6Y11_LUT4AB/FrameStrobe[11]
+ Tile_X6Y11_LUT4AB/FrameStrobe[12] Tile_X6Y11_LUT4AB/FrameStrobe[13] Tile_X6Y11_LUT4AB/FrameStrobe[14]
+ Tile_X6Y11_LUT4AB/FrameStrobe[15] Tile_X6Y11_LUT4AB/FrameStrobe[16] Tile_X6Y11_LUT4AB/FrameStrobe[17]
+ Tile_X6Y11_LUT4AB/FrameStrobe[18] Tile_X6Y11_LUT4AB/FrameStrobe[19] Tile_X6Y11_LUT4AB/FrameStrobe[1]
+ Tile_X6Y11_LUT4AB/FrameStrobe[2] Tile_X6Y11_LUT4AB/FrameStrobe[3] Tile_X6Y11_LUT4AB/FrameStrobe[4]
+ Tile_X6Y11_LUT4AB/FrameStrobe[5] Tile_X6Y11_LUT4AB/FrameStrobe[6] Tile_X6Y11_LUT4AB/FrameStrobe[7]
+ Tile_X6Y11_LUT4AB/FrameStrobe[8] Tile_X6Y11_LUT4AB/FrameStrobe[9] Tile_X6Y10_LUT4AB/FrameStrobe[0]
+ Tile_X6Y10_LUT4AB/FrameStrobe[10] Tile_X6Y10_LUT4AB/FrameStrobe[11] Tile_X6Y10_LUT4AB/FrameStrobe[12]
+ Tile_X6Y10_LUT4AB/FrameStrobe[13] Tile_X6Y10_LUT4AB/FrameStrobe[14] Tile_X6Y10_LUT4AB/FrameStrobe[15]
+ Tile_X6Y10_LUT4AB/FrameStrobe[16] Tile_X6Y10_LUT4AB/FrameStrobe[17] Tile_X6Y10_LUT4AB/FrameStrobe[18]
+ Tile_X6Y10_LUT4AB/FrameStrobe[19] Tile_X6Y10_LUT4AB/FrameStrobe[1] Tile_X6Y10_LUT4AB/FrameStrobe[2]
+ Tile_X6Y10_LUT4AB/FrameStrobe[3] Tile_X6Y10_LUT4AB/FrameStrobe[4] Tile_X6Y10_LUT4AB/FrameStrobe[5]
+ Tile_X6Y10_LUT4AB/FrameStrobe[6] Tile_X6Y10_LUT4AB/FrameStrobe[7] Tile_X6Y10_LUT4AB/FrameStrobe[8]
+ Tile_X6Y10_LUT4AB/FrameStrobe[9] Tile_X6Y11_LUT4AB/N1BEG[0] Tile_X6Y11_LUT4AB/N1BEG[1]
+ Tile_X6Y11_LUT4AB/N1BEG[2] Tile_X6Y11_LUT4AB/N1BEG[3] Tile_X6Y12_LUT4AB/N1BEG[0]
+ Tile_X6Y12_LUT4AB/N1BEG[1] Tile_X6Y12_LUT4AB/N1BEG[2] Tile_X6Y12_LUT4AB/N1BEG[3]
+ Tile_X6Y11_LUT4AB/N2BEG[0] Tile_X6Y11_LUT4AB/N2BEG[1] Tile_X6Y11_LUT4AB/N2BEG[2]
+ Tile_X6Y11_LUT4AB/N2BEG[3] Tile_X6Y11_LUT4AB/N2BEG[4] Tile_X6Y11_LUT4AB/N2BEG[5]
+ Tile_X6Y11_LUT4AB/N2BEG[6] Tile_X6Y11_LUT4AB/N2BEG[7] Tile_X6Y10_LUT4AB/N2END[0]
+ Tile_X6Y10_LUT4AB/N2END[1] Tile_X6Y10_LUT4AB/N2END[2] Tile_X6Y10_LUT4AB/N2END[3]
+ Tile_X6Y10_LUT4AB/N2END[4] Tile_X6Y10_LUT4AB/N2END[5] Tile_X6Y10_LUT4AB/N2END[6]
+ Tile_X6Y10_LUT4AB/N2END[7] Tile_X6Y11_LUT4AB/N2END[0] Tile_X6Y11_LUT4AB/N2END[1]
+ Tile_X6Y11_LUT4AB/N2END[2] Tile_X6Y11_LUT4AB/N2END[3] Tile_X6Y11_LUT4AB/N2END[4]
+ Tile_X6Y11_LUT4AB/N2END[5] Tile_X6Y11_LUT4AB/N2END[6] Tile_X6Y11_LUT4AB/N2END[7]
+ Tile_X6Y12_LUT4AB/N2BEG[0] Tile_X6Y12_LUT4AB/N2BEG[1] Tile_X6Y12_LUT4AB/N2BEG[2]
+ Tile_X6Y12_LUT4AB/N2BEG[3] Tile_X6Y12_LUT4AB/N2BEG[4] Tile_X6Y12_LUT4AB/N2BEG[5]
+ Tile_X6Y12_LUT4AB/N2BEG[6] Tile_X6Y12_LUT4AB/N2BEG[7] Tile_X6Y11_LUT4AB/N4BEG[0]
+ Tile_X6Y11_LUT4AB/N4BEG[10] Tile_X6Y11_LUT4AB/N4BEG[11] Tile_X6Y11_LUT4AB/N4BEG[12]
+ Tile_X6Y11_LUT4AB/N4BEG[13] Tile_X6Y11_LUT4AB/N4BEG[14] Tile_X6Y11_LUT4AB/N4BEG[15]
+ Tile_X6Y11_LUT4AB/N4BEG[1] Tile_X6Y11_LUT4AB/N4BEG[2] Tile_X6Y11_LUT4AB/N4BEG[3]
+ Tile_X6Y11_LUT4AB/N4BEG[4] Tile_X6Y11_LUT4AB/N4BEG[5] Tile_X6Y11_LUT4AB/N4BEG[6]
+ Tile_X6Y11_LUT4AB/N4BEG[7] Tile_X6Y11_LUT4AB/N4BEG[8] Tile_X6Y11_LUT4AB/N4BEG[9]
+ Tile_X6Y12_LUT4AB/N4BEG[0] Tile_X6Y12_LUT4AB/N4BEG[10] Tile_X6Y12_LUT4AB/N4BEG[11]
+ Tile_X6Y12_LUT4AB/N4BEG[12] Tile_X6Y12_LUT4AB/N4BEG[13] Tile_X6Y12_LUT4AB/N4BEG[14]
+ Tile_X6Y12_LUT4AB/N4BEG[15] Tile_X6Y12_LUT4AB/N4BEG[1] Tile_X6Y12_LUT4AB/N4BEG[2]
+ Tile_X6Y12_LUT4AB/N4BEG[3] Tile_X6Y12_LUT4AB/N4BEG[4] Tile_X6Y12_LUT4AB/N4BEG[5]
+ Tile_X6Y12_LUT4AB/N4BEG[6] Tile_X6Y12_LUT4AB/N4BEG[7] Tile_X6Y12_LUT4AB/N4BEG[8]
+ Tile_X6Y12_LUT4AB/N4BEG[9] Tile_X6Y11_LUT4AB/NN4BEG[0] Tile_X6Y11_LUT4AB/NN4BEG[10]
+ Tile_X6Y11_LUT4AB/NN4BEG[11] Tile_X6Y11_LUT4AB/NN4BEG[12] Tile_X6Y11_LUT4AB/NN4BEG[13]
+ Tile_X6Y11_LUT4AB/NN4BEG[14] Tile_X6Y11_LUT4AB/NN4BEG[15] Tile_X6Y11_LUT4AB/NN4BEG[1]
+ Tile_X6Y11_LUT4AB/NN4BEG[2] Tile_X6Y11_LUT4AB/NN4BEG[3] Tile_X6Y11_LUT4AB/NN4BEG[4]
+ Tile_X6Y11_LUT4AB/NN4BEG[5] Tile_X6Y11_LUT4AB/NN4BEG[6] Tile_X6Y11_LUT4AB/NN4BEG[7]
+ Tile_X6Y11_LUT4AB/NN4BEG[8] Tile_X6Y11_LUT4AB/NN4BEG[9] Tile_X6Y12_LUT4AB/NN4BEG[0]
+ Tile_X6Y12_LUT4AB/NN4BEG[10] Tile_X6Y12_LUT4AB/NN4BEG[11] Tile_X6Y12_LUT4AB/NN4BEG[12]
+ Tile_X6Y12_LUT4AB/NN4BEG[13] Tile_X6Y12_LUT4AB/NN4BEG[14] Tile_X6Y12_LUT4AB/NN4BEG[15]
+ Tile_X6Y12_LUT4AB/NN4BEG[1] Tile_X6Y12_LUT4AB/NN4BEG[2] Tile_X6Y12_LUT4AB/NN4BEG[3]
+ Tile_X6Y12_LUT4AB/NN4BEG[4] Tile_X6Y12_LUT4AB/NN4BEG[5] Tile_X6Y12_LUT4AB/NN4BEG[6]
+ Tile_X6Y12_LUT4AB/NN4BEG[7] Tile_X6Y12_LUT4AB/NN4BEG[8] Tile_X6Y12_LUT4AB/NN4BEG[9]
+ Tile_X6Y12_LUT4AB/S1END[0] Tile_X6Y12_LUT4AB/S1END[1] Tile_X6Y12_LUT4AB/S1END[2]
+ Tile_X6Y12_LUT4AB/S1END[3] Tile_X6Y11_LUT4AB/S1END[0] Tile_X6Y11_LUT4AB/S1END[1]
+ Tile_X6Y11_LUT4AB/S1END[2] Tile_X6Y11_LUT4AB/S1END[3] Tile_X6Y12_LUT4AB/S2MID[0]
+ Tile_X6Y12_LUT4AB/S2MID[1] Tile_X6Y12_LUT4AB/S2MID[2] Tile_X6Y12_LUT4AB/S2MID[3]
+ Tile_X6Y12_LUT4AB/S2MID[4] Tile_X6Y12_LUT4AB/S2MID[5] Tile_X6Y12_LUT4AB/S2MID[6]
+ Tile_X6Y12_LUT4AB/S2MID[7] Tile_X6Y12_LUT4AB/S2END[0] Tile_X6Y12_LUT4AB/S2END[1]
+ Tile_X6Y12_LUT4AB/S2END[2] Tile_X6Y12_LUT4AB/S2END[3] Tile_X6Y12_LUT4AB/S2END[4]
+ Tile_X6Y12_LUT4AB/S2END[5] Tile_X6Y12_LUT4AB/S2END[6] Tile_X6Y12_LUT4AB/S2END[7]
+ Tile_X6Y11_LUT4AB/S2END[0] Tile_X6Y11_LUT4AB/S2END[1] Tile_X6Y11_LUT4AB/S2END[2]
+ Tile_X6Y11_LUT4AB/S2END[3] Tile_X6Y11_LUT4AB/S2END[4] Tile_X6Y11_LUT4AB/S2END[5]
+ Tile_X6Y11_LUT4AB/S2END[6] Tile_X6Y11_LUT4AB/S2END[7] Tile_X6Y11_LUT4AB/S2MID[0]
+ Tile_X6Y11_LUT4AB/S2MID[1] Tile_X6Y11_LUT4AB/S2MID[2] Tile_X6Y11_LUT4AB/S2MID[3]
+ Tile_X6Y11_LUT4AB/S2MID[4] Tile_X6Y11_LUT4AB/S2MID[5] Tile_X6Y11_LUT4AB/S2MID[6]
+ Tile_X6Y11_LUT4AB/S2MID[7] Tile_X6Y12_LUT4AB/S4END[0] Tile_X6Y12_LUT4AB/S4END[10]
+ Tile_X6Y12_LUT4AB/S4END[11] Tile_X6Y12_LUT4AB/S4END[12] Tile_X6Y12_LUT4AB/S4END[13]
+ Tile_X6Y12_LUT4AB/S4END[14] Tile_X6Y12_LUT4AB/S4END[15] Tile_X6Y12_LUT4AB/S4END[1]
+ Tile_X6Y12_LUT4AB/S4END[2] Tile_X6Y12_LUT4AB/S4END[3] Tile_X6Y12_LUT4AB/S4END[4]
+ Tile_X6Y12_LUT4AB/S4END[5] Tile_X6Y12_LUT4AB/S4END[6] Tile_X6Y12_LUT4AB/S4END[7]
+ Tile_X6Y12_LUT4AB/S4END[8] Tile_X6Y12_LUT4AB/S4END[9] Tile_X6Y11_LUT4AB/S4END[0]
+ Tile_X6Y11_LUT4AB/S4END[10] Tile_X6Y11_LUT4AB/S4END[11] Tile_X6Y11_LUT4AB/S4END[12]
+ Tile_X6Y11_LUT4AB/S4END[13] Tile_X6Y11_LUT4AB/S4END[14] Tile_X6Y11_LUT4AB/S4END[15]
+ Tile_X6Y11_LUT4AB/S4END[1] Tile_X6Y11_LUT4AB/S4END[2] Tile_X6Y11_LUT4AB/S4END[3]
+ Tile_X6Y11_LUT4AB/S4END[4] Tile_X6Y11_LUT4AB/S4END[5] Tile_X6Y11_LUT4AB/S4END[6]
+ Tile_X6Y11_LUT4AB/S4END[7] Tile_X6Y11_LUT4AB/S4END[8] Tile_X6Y11_LUT4AB/S4END[9]
+ Tile_X6Y12_LUT4AB/SS4END[0] Tile_X6Y12_LUT4AB/SS4END[10] Tile_X6Y12_LUT4AB/SS4END[11]
+ Tile_X6Y12_LUT4AB/SS4END[12] Tile_X6Y12_LUT4AB/SS4END[13] Tile_X6Y12_LUT4AB/SS4END[14]
+ Tile_X6Y12_LUT4AB/SS4END[15] Tile_X6Y12_LUT4AB/SS4END[1] Tile_X6Y12_LUT4AB/SS4END[2]
+ Tile_X6Y12_LUT4AB/SS4END[3] Tile_X6Y12_LUT4AB/SS4END[4] Tile_X6Y12_LUT4AB/SS4END[5]
+ Tile_X6Y12_LUT4AB/SS4END[6] Tile_X6Y12_LUT4AB/SS4END[7] Tile_X6Y12_LUT4AB/SS4END[8]
+ Tile_X6Y12_LUT4AB/SS4END[9] Tile_X6Y11_LUT4AB/SS4END[0] Tile_X6Y11_LUT4AB/SS4END[10]
+ Tile_X6Y11_LUT4AB/SS4END[11] Tile_X6Y11_LUT4AB/SS4END[12] Tile_X6Y11_LUT4AB/SS4END[13]
+ Tile_X6Y11_LUT4AB/SS4END[14] Tile_X6Y11_LUT4AB/SS4END[15] Tile_X6Y11_LUT4AB/SS4END[1]
+ Tile_X6Y11_LUT4AB/SS4END[2] Tile_X6Y11_LUT4AB/SS4END[3] Tile_X6Y11_LUT4AB/SS4END[4]
+ Tile_X6Y11_LUT4AB/SS4END[5] Tile_X6Y11_LUT4AB/SS4END[6] Tile_X6Y11_LUT4AB/SS4END[7]
+ Tile_X6Y11_LUT4AB/SS4END[8] Tile_X6Y11_LUT4AB/SS4END[9] Tile_X6Y11_LUT4AB/UserCLK
+ Tile_X6Y10_LUT4AB/UserCLK VGND VPWR Tile_X6Y11_LUT4AB/W1BEG[0] Tile_X6Y11_LUT4AB/W1BEG[1]
+ Tile_X6Y11_LUT4AB/W1BEG[2] Tile_X6Y11_LUT4AB/W1BEG[3] Tile_X6Y11_LUT4AB/W1END[0]
+ Tile_X6Y11_LUT4AB/W1END[1] Tile_X6Y11_LUT4AB/W1END[2] Tile_X6Y11_LUT4AB/W1END[3]
+ Tile_X6Y11_LUT4AB/W2BEG[0] Tile_X6Y11_LUT4AB/W2BEG[1] Tile_X6Y11_LUT4AB/W2BEG[2]
+ Tile_X6Y11_LUT4AB/W2BEG[3] Tile_X6Y11_LUT4AB/W2BEG[4] Tile_X6Y11_LUT4AB/W2BEG[5]
+ Tile_X6Y11_LUT4AB/W2BEG[6] Tile_X6Y11_LUT4AB/W2BEG[7] Tile_X5Y11_LUT4AB/W2END[0]
+ Tile_X5Y11_LUT4AB/W2END[1] Tile_X5Y11_LUT4AB/W2END[2] Tile_X5Y11_LUT4AB/W2END[3]
+ Tile_X5Y11_LUT4AB/W2END[4] Tile_X5Y11_LUT4AB/W2END[5] Tile_X5Y11_LUT4AB/W2END[6]
+ Tile_X5Y11_LUT4AB/W2END[7] Tile_X6Y11_LUT4AB/W2END[0] Tile_X6Y11_LUT4AB/W2END[1]
+ Tile_X6Y11_LUT4AB/W2END[2] Tile_X6Y11_LUT4AB/W2END[3] Tile_X6Y11_LUT4AB/W2END[4]
+ Tile_X6Y11_LUT4AB/W2END[5] Tile_X6Y11_LUT4AB/W2END[6] Tile_X6Y11_LUT4AB/W2END[7]
+ Tile_X6Y11_LUT4AB/W2MID[0] Tile_X6Y11_LUT4AB/W2MID[1] Tile_X6Y11_LUT4AB/W2MID[2]
+ Tile_X6Y11_LUT4AB/W2MID[3] Tile_X6Y11_LUT4AB/W2MID[4] Tile_X6Y11_LUT4AB/W2MID[5]
+ Tile_X6Y11_LUT4AB/W2MID[6] Tile_X6Y11_LUT4AB/W2MID[7] Tile_X6Y11_LUT4AB/W6BEG[0]
+ Tile_X6Y11_LUT4AB/W6BEG[10] Tile_X6Y11_LUT4AB/W6BEG[11] Tile_X6Y11_LUT4AB/W6BEG[1]
+ Tile_X6Y11_LUT4AB/W6BEG[2] Tile_X6Y11_LUT4AB/W6BEG[3] Tile_X6Y11_LUT4AB/W6BEG[4]
+ Tile_X6Y11_LUT4AB/W6BEG[5] Tile_X6Y11_LUT4AB/W6BEG[6] Tile_X6Y11_LUT4AB/W6BEG[7]
+ Tile_X6Y11_LUT4AB/W6BEG[8] Tile_X6Y11_LUT4AB/W6BEG[9] Tile_X6Y11_LUT4AB/W6END[0]
+ Tile_X6Y11_LUT4AB/W6END[10] Tile_X6Y11_LUT4AB/W6END[11] Tile_X6Y11_LUT4AB/W6END[1]
+ Tile_X6Y11_LUT4AB/W6END[2] Tile_X6Y11_LUT4AB/W6END[3] Tile_X6Y11_LUT4AB/W6END[4]
+ Tile_X6Y11_LUT4AB/W6END[5] Tile_X6Y11_LUT4AB/W6END[6] Tile_X6Y11_LUT4AB/W6END[7]
+ Tile_X6Y11_LUT4AB/W6END[8] Tile_X6Y11_LUT4AB/W6END[9] Tile_X6Y11_LUT4AB/WW4BEG[0]
+ Tile_X6Y11_LUT4AB/WW4BEG[10] Tile_X6Y11_LUT4AB/WW4BEG[11] Tile_X6Y11_LUT4AB/WW4BEG[12]
+ Tile_X6Y11_LUT4AB/WW4BEG[13] Tile_X6Y11_LUT4AB/WW4BEG[14] Tile_X6Y11_LUT4AB/WW4BEG[15]
+ Tile_X6Y11_LUT4AB/WW4BEG[1] Tile_X6Y11_LUT4AB/WW4BEG[2] Tile_X6Y11_LUT4AB/WW4BEG[3]
+ Tile_X6Y11_LUT4AB/WW4BEG[4] Tile_X6Y11_LUT4AB/WW4BEG[5] Tile_X6Y11_LUT4AB/WW4BEG[6]
+ Tile_X6Y11_LUT4AB/WW4BEG[7] Tile_X6Y11_LUT4AB/WW4BEG[8] Tile_X6Y11_LUT4AB/WW4BEG[9]
+ Tile_X6Y11_LUT4AB/WW4END[0] Tile_X6Y11_LUT4AB/WW4END[10] Tile_X6Y11_LUT4AB/WW4END[11]
+ Tile_X6Y11_LUT4AB/WW4END[12] Tile_X6Y11_LUT4AB/WW4END[13] Tile_X6Y11_LUT4AB/WW4END[14]
+ Tile_X6Y11_LUT4AB/WW4END[15] Tile_X6Y11_LUT4AB/WW4END[1] Tile_X6Y11_LUT4AB/WW4END[2]
+ Tile_X6Y11_LUT4AB/WW4END[3] Tile_X6Y11_LUT4AB/WW4END[4] Tile_X6Y11_LUT4AB/WW4END[5]
+ Tile_X6Y11_LUT4AB/WW4END[6] Tile_X6Y11_LUT4AB/WW4END[7] Tile_X6Y11_LUT4AB/WW4END[8]
+ Tile_X6Y11_LUT4AB/WW4END[9] LUT4AB
XTile_X1Y10_LUT4AB Tile_X1Y11_LUT4AB/Co Tile_X1Y9_LUT4AB/Ci Tile_X2Y10_LUT4AB/E1END[0]
+ Tile_X2Y10_LUT4AB/E1END[1] Tile_X2Y10_LUT4AB/E1END[2] Tile_X2Y10_LUT4AB/E1END[3]
+ Tile_X0Y10_W_IO/E1BEG[0] Tile_X0Y10_W_IO/E1BEG[1] Tile_X0Y10_W_IO/E1BEG[2] Tile_X0Y10_W_IO/E1BEG[3]
+ Tile_X2Y10_LUT4AB/E2MID[0] Tile_X2Y10_LUT4AB/E2MID[1] Tile_X2Y10_LUT4AB/E2MID[2]
+ Tile_X2Y10_LUT4AB/E2MID[3] Tile_X2Y10_LUT4AB/E2MID[4] Tile_X2Y10_LUT4AB/E2MID[5]
+ Tile_X2Y10_LUT4AB/E2MID[6] Tile_X2Y10_LUT4AB/E2MID[7] Tile_X2Y10_LUT4AB/E2END[0]
+ Tile_X2Y10_LUT4AB/E2END[1] Tile_X2Y10_LUT4AB/E2END[2] Tile_X2Y10_LUT4AB/E2END[3]
+ Tile_X2Y10_LUT4AB/E2END[4] Tile_X2Y10_LUT4AB/E2END[5] Tile_X2Y10_LUT4AB/E2END[6]
+ Tile_X2Y10_LUT4AB/E2END[7] Tile_X0Y10_W_IO/E2BEGb[0] Tile_X0Y10_W_IO/E2BEGb[1] Tile_X0Y10_W_IO/E2BEGb[2]
+ Tile_X0Y10_W_IO/E2BEGb[3] Tile_X0Y10_W_IO/E2BEGb[4] Tile_X0Y10_W_IO/E2BEGb[5] Tile_X0Y10_W_IO/E2BEGb[6]
+ Tile_X0Y10_W_IO/E2BEGb[7] Tile_X0Y10_W_IO/E2BEG[0] Tile_X0Y10_W_IO/E2BEG[1] Tile_X0Y10_W_IO/E2BEG[2]
+ Tile_X0Y10_W_IO/E2BEG[3] Tile_X0Y10_W_IO/E2BEG[4] Tile_X0Y10_W_IO/E2BEG[5] Tile_X0Y10_W_IO/E2BEG[6]
+ Tile_X0Y10_W_IO/E2BEG[7] Tile_X2Y10_LUT4AB/E6END[0] Tile_X2Y10_LUT4AB/E6END[10]
+ Tile_X2Y10_LUT4AB/E6END[11] Tile_X2Y10_LUT4AB/E6END[1] Tile_X2Y10_LUT4AB/E6END[2]
+ Tile_X2Y10_LUT4AB/E6END[3] Tile_X2Y10_LUT4AB/E6END[4] Tile_X2Y10_LUT4AB/E6END[5]
+ Tile_X2Y10_LUT4AB/E6END[6] Tile_X2Y10_LUT4AB/E6END[7] Tile_X2Y10_LUT4AB/E6END[8]
+ Tile_X2Y10_LUT4AB/E6END[9] Tile_X0Y10_W_IO/E6BEG[0] Tile_X0Y10_W_IO/E6BEG[10] Tile_X0Y10_W_IO/E6BEG[11]
+ Tile_X0Y10_W_IO/E6BEG[1] Tile_X0Y10_W_IO/E6BEG[2] Tile_X0Y10_W_IO/E6BEG[3] Tile_X0Y10_W_IO/E6BEG[4]
+ Tile_X0Y10_W_IO/E6BEG[5] Tile_X0Y10_W_IO/E6BEG[6] Tile_X0Y10_W_IO/E6BEG[7] Tile_X0Y10_W_IO/E6BEG[8]
+ Tile_X0Y10_W_IO/E6BEG[9] Tile_X2Y10_LUT4AB/EE4END[0] Tile_X2Y10_LUT4AB/EE4END[10]
+ Tile_X2Y10_LUT4AB/EE4END[11] Tile_X2Y10_LUT4AB/EE4END[12] Tile_X2Y10_LUT4AB/EE4END[13]
+ Tile_X2Y10_LUT4AB/EE4END[14] Tile_X2Y10_LUT4AB/EE4END[15] Tile_X2Y10_LUT4AB/EE4END[1]
+ Tile_X2Y10_LUT4AB/EE4END[2] Tile_X2Y10_LUT4AB/EE4END[3] Tile_X2Y10_LUT4AB/EE4END[4]
+ Tile_X2Y10_LUT4AB/EE4END[5] Tile_X2Y10_LUT4AB/EE4END[6] Tile_X2Y10_LUT4AB/EE4END[7]
+ Tile_X2Y10_LUT4AB/EE4END[8] Tile_X2Y10_LUT4AB/EE4END[9] Tile_X0Y10_W_IO/EE4BEG[0]
+ Tile_X0Y10_W_IO/EE4BEG[10] Tile_X0Y10_W_IO/EE4BEG[11] Tile_X0Y10_W_IO/EE4BEG[12]
+ Tile_X0Y10_W_IO/EE4BEG[13] Tile_X0Y10_W_IO/EE4BEG[14] Tile_X0Y10_W_IO/EE4BEG[15]
+ Tile_X0Y10_W_IO/EE4BEG[1] Tile_X0Y10_W_IO/EE4BEG[2] Tile_X0Y10_W_IO/EE4BEG[3] Tile_X0Y10_W_IO/EE4BEG[4]
+ Tile_X0Y10_W_IO/EE4BEG[5] Tile_X0Y10_W_IO/EE4BEG[6] Tile_X0Y10_W_IO/EE4BEG[7] Tile_X0Y10_W_IO/EE4BEG[8]
+ Tile_X0Y10_W_IO/EE4BEG[9] Tile_X1Y10_LUT4AB/FrameData[0] Tile_X1Y10_LUT4AB/FrameData[10]
+ Tile_X1Y10_LUT4AB/FrameData[11] Tile_X1Y10_LUT4AB/FrameData[12] Tile_X1Y10_LUT4AB/FrameData[13]
+ Tile_X1Y10_LUT4AB/FrameData[14] Tile_X1Y10_LUT4AB/FrameData[15] Tile_X1Y10_LUT4AB/FrameData[16]
+ Tile_X1Y10_LUT4AB/FrameData[17] Tile_X1Y10_LUT4AB/FrameData[18] Tile_X1Y10_LUT4AB/FrameData[19]
+ Tile_X1Y10_LUT4AB/FrameData[1] Tile_X1Y10_LUT4AB/FrameData[20] Tile_X1Y10_LUT4AB/FrameData[21]
+ Tile_X1Y10_LUT4AB/FrameData[22] Tile_X1Y10_LUT4AB/FrameData[23] Tile_X1Y10_LUT4AB/FrameData[24]
+ Tile_X1Y10_LUT4AB/FrameData[25] Tile_X1Y10_LUT4AB/FrameData[26] Tile_X1Y10_LUT4AB/FrameData[27]
+ Tile_X1Y10_LUT4AB/FrameData[28] Tile_X1Y10_LUT4AB/FrameData[29] Tile_X1Y10_LUT4AB/FrameData[2]
+ Tile_X1Y10_LUT4AB/FrameData[30] Tile_X1Y10_LUT4AB/FrameData[31] Tile_X1Y10_LUT4AB/FrameData[3]
+ Tile_X1Y10_LUT4AB/FrameData[4] Tile_X1Y10_LUT4AB/FrameData[5] Tile_X1Y10_LUT4AB/FrameData[6]
+ Tile_X1Y10_LUT4AB/FrameData[7] Tile_X1Y10_LUT4AB/FrameData[8] Tile_X1Y10_LUT4AB/FrameData[9]
+ Tile_X2Y10_LUT4AB/FrameData[0] Tile_X2Y10_LUT4AB/FrameData[10] Tile_X2Y10_LUT4AB/FrameData[11]
+ Tile_X2Y10_LUT4AB/FrameData[12] Tile_X2Y10_LUT4AB/FrameData[13] Tile_X2Y10_LUT4AB/FrameData[14]
+ Tile_X2Y10_LUT4AB/FrameData[15] Tile_X2Y10_LUT4AB/FrameData[16] Tile_X2Y10_LUT4AB/FrameData[17]
+ Tile_X2Y10_LUT4AB/FrameData[18] Tile_X2Y10_LUT4AB/FrameData[19] Tile_X2Y10_LUT4AB/FrameData[1]
+ Tile_X2Y10_LUT4AB/FrameData[20] Tile_X2Y10_LUT4AB/FrameData[21] Tile_X2Y10_LUT4AB/FrameData[22]
+ Tile_X2Y10_LUT4AB/FrameData[23] Tile_X2Y10_LUT4AB/FrameData[24] Tile_X2Y10_LUT4AB/FrameData[25]
+ Tile_X2Y10_LUT4AB/FrameData[26] Tile_X2Y10_LUT4AB/FrameData[27] Tile_X2Y10_LUT4AB/FrameData[28]
+ Tile_X2Y10_LUT4AB/FrameData[29] Tile_X2Y10_LUT4AB/FrameData[2] Tile_X2Y10_LUT4AB/FrameData[30]
+ Tile_X2Y10_LUT4AB/FrameData[31] Tile_X2Y10_LUT4AB/FrameData[3] Tile_X2Y10_LUT4AB/FrameData[4]
+ Tile_X2Y10_LUT4AB/FrameData[5] Tile_X2Y10_LUT4AB/FrameData[6] Tile_X2Y10_LUT4AB/FrameData[7]
+ Tile_X2Y10_LUT4AB/FrameData[8] Tile_X2Y10_LUT4AB/FrameData[9] Tile_X1Y10_LUT4AB/FrameStrobe[0]
+ Tile_X1Y10_LUT4AB/FrameStrobe[10] Tile_X1Y10_LUT4AB/FrameStrobe[11] Tile_X1Y10_LUT4AB/FrameStrobe[12]
+ Tile_X1Y10_LUT4AB/FrameStrobe[13] Tile_X1Y10_LUT4AB/FrameStrobe[14] Tile_X1Y10_LUT4AB/FrameStrobe[15]
+ Tile_X1Y10_LUT4AB/FrameStrobe[16] Tile_X1Y10_LUT4AB/FrameStrobe[17] Tile_X1Y10_LUT4AB/FrameStrobe[18]
+ Tile_X1Y10_LUT4AB/FrameStrobe[19] Tile_X1Y10_LUT4AB/FrameStrobe[1] Tile_X1Y10_LUT4AB/FrameStrobe[2]
+ Tile_X1Y10_LUT4AB/FrameStrobe[3] Tile_X1Y10_LUT4AB/FrameStrobe[4] Tile_X1Y10_LUT4AB/FrameStrobe[5]
+ Tile_X1Y10_LUT4AB/FrameStrobe[6] Tile_X1Y10_LUT4AB/FrameStrobe[7] Tile_X1Y10_LUT4AB/FrameStrobe[8]
+ Tile_X1Y10_LUT4AB/FrameStrobe[9] Tile_X1Y9_LUT4AB/FrameStrobe[0] Tile_X1Y9_LUT4AB/FrameStrobe[10]
+ Tile_X1Y9_LUT4AB/FrameStrobe[11] Tile_X1Y9_LUT4AB/FrameStrobe[12] Tile_X1Y9_LUT4AB/FrameStrobe[13]
+ Tile_X1Y9_LUT4AB/FrameStrobe[14] Tile_X1Y9_LUT4AB/FrameStrobe[15] Tile_X1Y9_LUT4AB/FrameStrobe[16]
+ Tile_X1Y9_LUT4AB/FrameStrobe[17] Tile_X1Y9_LUT4AB/FrameStrobe[18] Tile_X1Y9_LUT4AB/FrameStrobe[19]
+ Tile_X1Y9_LUT4AB/FrameStrobe[1] Tile_X1Y9_LUT4AB/FrameStrobe[2] Tile_X1Y9_LUT4AB/FrameStrobe[3]
+ Tile_X1Y9_LUT4AB/FrameStrobe[4] Tile_X1Y9_LUT4AB/FrameStrobe[5] Tile_X1Y9_LUT4AB/FrameStrobe[6]
+ Tile_X1Y9_LUT4AB/FrameStrobe[7] Tile_X1Y9_LUT4AB/FrameStrobe[8] Tile_X1Y9_LUT4AB/FrameStrobe[9]
+ Tile_X1Y9_LUT4AB/N1END[0] Tile_X1Y9_LUT4AB/N1END[1] Tile_X1Y9_LUT4AB/N1END[2] Tile_X1Y9_LUT4AB/N1END[3]
+ Tile_X1Y11_LUT4AB/N1BEG[0] Tile_X1Y11_LUT4AB/N1BEG[1] Tile_X1Y11_LUT4AB/N1BEG[2]
+ Tile_X1Y11_LUT4AB/N1BEG[3] Tile_X1Y9_LUT4AB/N2MID[0] Tile_X1Y9_LUT4AB/N2MID[1] Tile_X1Y9_LUT4AB/N2MID[2]
+ Tile_X1Y9_LUT4AB/N2MID[3] Tile_X1Y9_LUT4AB/N2MID[4] Tile_X1Y9_LUT4AB/N2MID[5] Tile_X1Y9_LUT4AB/N2MID[6]
+ Tile_X1Y9_LUT4AB/N2MID[7] Tile_X1Y9_LUT4AB/N2END[0] Tile_X1Y9_LUT4AB/N2END[1] Tile_X1Y9_LUT4AB/N2END[2]
+ Tile_X1Y9_LUT4AB/N2END[3] Tile_X1Y9_LUT4AB/N2END[4] Tile_X1Y9_LUT4AB/N2END[5] Tile_X1Y9_LUT4AB/N2END[6]
+ Tile_X1Y9_LUT4AB/N2END[7] Tile_X1Y10_LUT4AB/N2END[0] Tile_X1Y10_LUT4AB/N2END[1]
+ Tile_X1Y10_LUT4AB/N2END[2] Tile_X1Y10_LUT4AB/N2END[3] Tile_X1Y10_LUT4AB/N2END[4]
+ Tile_X1Y10_LUT4AB/N2END[5] Tile_X1Y10_LUT4AB/N2END[6] Tile_X1Y10_LUT4AB/N2END[7]
+ Tile_X1Y11_LUT4AB/N2BEG[0] Tile_X1Y11_LUT4AB/N2BEG[1] Tile_X1Y11_LUT4AB/N2BEG[2]
+ Tile_X1Y11_LUT4AB/N2BEG[3] Tile_X1Y11_LUT4AB/N2BEG[4] Tile_X1Y11_LUT4AB/N2BEG[5]
+ Tile_X1Y11_LUT4AB/N2BEG[6] Tile_X1Y11_LUT4AB/N2BEG[7] Tile_X1Y9_LUT4AB/N4END[0]
+ Tile_X1Y9_LUT4AB/N4END[10] Tile_X1Y9_LUT4AB/N4END[11] Tile_X1Y9_LUT4AB/N4END[12]
+ Tile_X1Y9_LUT4AB/N4END[13] Tile_X1Y9_LUT4AB/N4END[14] Tile_X1Y9_LUT4AB/N4END[15]
+ Tile_X1Y9_LUT4AB/N4END[1] Tile_X1Y9_LUT4AB/N4END[2] Tile_X1Y9_LUT4AB/N4END[3] Tile_X1Y9_LUT4AB/N4END[4]
+ Tile_X1Y9_LUT4AB/N4END[5] Tile_X1Y9_LUT4AB/N4END[6] Tile_X1Y9_LUT4AB/N4END[7] Tile_X1Y9_LUT4AB/N4END[8]
+ Tile_X1Y9_LUT4AB/N4END[9] Tile_X1Y11_LUT4AB/N4BEG[0] Tile_X1Y11_LUT4AB/N4BEG[10]
+ Tile_X1Y11_LUT4AB/N4BEG[11] Tile_X1Y11_LUT4AB/N4BEG[12] Tile_X1Y11_LUT4AB/N4BEG[13]
+ Tile_X1Y11_LUT4AB/N4BEG[14] Tile_X1Y11_LUT4AB/N4BEG[15] Tile_X1Y11_LUT4AB/N4BEG[1]
+ Tile_X1Y11_LUT4AB/N4BEG[2] Tile_X1Y11_LUT4AB/N4BEG[3] Tile_X1Y11_LUT4AB/N4BEG[4]
+ Tile_X1Y11_LUT4AB/N4BEG[5] Tile_X1Y11_LUT4AB/N4BEG[6] Tile_X1Y11_LUT4AB/N4BEG[7]
+ Tile_X1Y11_LUT4AB/N4BEG[8] Tile_X1Y11_LUT4AB/N4BEG[9] Tile_X1Y9_LUT4AB/NN4END[0]
+ Tile_X1Y9_LUT4AB/NN4END[10] Tile_X1Y9_LUT4AB/NN4END[11] Tile_X1Y9_LUT4AB/NN4END[12]
+ Tile_X1Y9_LUT4AB/NN4END[13] Tile_X1Y9_LUT4AB/NN4END[14] Tile_X1Y9_LUT4AB/NN4END[15]
+ Tile_X1Y9_LUT4AB/NN4END[1] Tile_X1Y9_LUT4AB/NN4END[2] Tile_X1Y9_LUT4AB/NN4END[3]
+ Tile_X1Y9_LUT4AB/NN4END[4] Tile_X1Y9_LUT4AB/NN4END[5] Tile_X1Y9_LUT4AB/NN4END[6]
+ Tile_X1Y9_LUT4AB/NN4END[7] Tile_X1Y9_LUT4AB/NN4END[8] Tile_X1Y9_LUT4AB/NN4END[9]
+ Tile_X1Y11_LUT4AB/NN4BEG[0] Tile_X1Y11_LUT4AB/NN4BEG[10] Tile_X1Y11_LUT4AB/NN4BEG[11]
+ Tile_X1Y11_LUT4AB/NN4BEG[12] Tile_X1Y11_LUT4AB/NN4BEG[13] Tile_X1Y11_LUT4AB/NN4BEG[14]
+ Tile_X1Y11_LUT4AB/NN4BEG[15] Tile_X1Y11_LUT4AB/NN4BEG[1] Tile_X1Y11_LUT4AB/NN4BEG[2]
+ Tile_X1Y11_LUT4AB/NN4BEG[3] Tile_X1Y11_LUT4AB/NN4BEG[4] Tile_X1Y11_LUT4AB/NN4BEG[5]
+ Tile_X1Y11_LUT4AB/NN4BEG[6] Tile_X1Y11_LUT4AB/NN4BEG[7] Tile_X1Y11_LUT4AB/NN4BEG[8]
+ Tile_X1Y11_LUT4AB/NN4BEG[9] Tile_X1Y11_LUT4AB/S1END[0] Tile_X1Y11_LUT4AB/S1END[1]
+ Tile_X1Y11_LUT4AB/S1END[2] Tile_X1Y11_LUT4AB/S1END[3] Tile_X1Y9_LUT4AB/S1BEG[0]
+ Tile_X1Y9_LUT4AB/S1BEG[1] Tile_X1Y9_LUT4AB/S1BEG[2] Tile_X1Y9_LUT4AB/S1BEG[3] Tile_X1Y11_LUT4AB/S2MID[0]
+ Tile_X1Y11_LUT4AB/S2MID[1] Tile_X1Y11_LUT4AB/S2MID[2] Tile_X1Y11_LUT4AB/S2MID[3]
+ Tile_X1Y11_LUT4AB/S2MID[4] Tile_X1Y11_LUT4AB/S2MID[5] Tile_X1Y11_LUT4AB/S2MID[6]
+ Tile_X1Y11_LUT4AB/S2MID[7] Tile_X1Y11_LUT4AB/S2END[0] Tile_X1Y11_LUT4AB/S2END[1]
+ Tile_X1Y11_LUT4AB/S2END[2] Tile_X1Y11_LUT4AB/S2END[3] Tile_X1Y11_LUT4AB/S2END[4]
+ Tile_X1Y11_LUT4AB/S2END[5] Tile_X1Y11_LUT4AB/S2END[6] Tile_X1Y11_LUT4AB/S2END[7]
+ Tile_X1Y9_LUT4AB/S2BEGb[0] Tile_X1Y9_LUT4AB/S2BEGb[1] Tile_X1Y9_LUT4AB/S2BEGb[2]
+ Tile_X1Y9_LUT4AB/S2BEGb[3] Tile_X1Y9_LUT4AB/S2BEGb[4] Tile_X1Y9_LUT4AB/S2BEGb[5]
+ Tile_X1Y9_LUT4AB/S2BEGb[6] Tile_X1Y9_LUT4AB/S2BEGb[7] Tile_X1Y9_LUT4AB/S2BEG[0]
+ Tile_X1Y9_LUT4AB/S2BEG[1] Tile_X1Y9_LUT4AB/S2BEG[2] Tile_X1Y9_LUT4AB/S2BEG[3] Tile_X1Y9_LUT4AB/S2BEG[4]
+ Tile_X1Y9_LUT4AB/S2BEG[5] Tile_X1Y9_LUT4AB/S2BEG[6] Tile_X1Y9_LUT4AB/S2BEG[7] Tile_X1Y11_LUT4AB/S4END[0]
+ Tile_X1Y11_LUT4AB/S4END[10] Tile_X1Y11_LUT4AB/S4END[11] Tile_X1Y11_LUT4AB/S4END[12]
+ Tile_X1Y11_LUT4AB/S4END[13] Tile_X1Y11_LUT4AB/S4END[14] Tile_X1Y11_LUT4AB/S4END[15]
+ Tile_X1Y11_LUT4AB/S4END[1] Tile_X1Y11_LUT4AB/S4END[2] Tile_X1Y11_LUT4AB/S4END[3]
+ Tile_X1Y11_LUT4AB/S4END[4] Tile_X1Y11_LUT4AB/S4END[5] Tile_X1Y11_LUT4AB/S4END[6]
+ Tile_X1Y11_LUT4AB/S4END[7] Tile_X1Y11_LUT4AB/S4END[8] Tile_X1Y11_LUT4AB/S4END[9]
+ Tile_X1Y9_LUT4AB/S4BEG[0] Tile_X1Y9_LUT4AB/S4BEG[10] Tile_X1Y9_LUT4AB/S4BEG[11]
+ Tile_X1Y9_LUT4AB/S4BEG[12] Tile_X1Y9_LUT4AB/S4BEG[13] Tile_X1Y9_LUT4AB/S4BEG[14]
+ Tile_X1Y9_LUT4AB/S4BEG[15] Tile_X1Y9_LUT4AB/S4BEG[1] Tile_X1Y9_LUT4AB/S4BEG[2] Tile_X1Y9_LUT4AB/S4BEG[3]
+ Tile_X1Y9_LUT4AB/S4BEG[4] Tile_X1Y9_LUT4AB/S4BEG[5] Tile_X1Y9_LUT4AB/S4BEG[6] Tile_X1Y9_LUT4AB/S4BEG[7]
+ Tile_X1Y9_LUT4AB/S4BEG[8] Tile_X1Y9_LUT4AB/S4BEG[9] Tile_X1Y11_LUT4AB/SS4END[0]
+ Tile_X1Y11_LUT4AB/SS4END[10] Tile_X1Y11_LUT4AB/SS4END[11] Tile_X1Y11_LUT4AB/SS4END[12]
+ Tile_X1Y11_LUT4AB/SS4END[13] Tile_X1Y11_LUT4AB/SS4END[14] Tile_X1Y11_LUT4AB/SS4END[15]
+ Tile_X1Y11_LUT4AB/SS4END[1] Tile_X1Y11_LUT4AB/SS4END[2] Tile_X1Y11_LUT4AB/SS4END[3]
+ Tile_X1Y11_LUT4AB/SS4END[4] Tile_X1Y11_LUT4AB/SS4END[5] Tile_X1Y11_LUT4AB/SS4END[6]
+ Tile_X1Y11_LUT4AB/SS4END[7] Tile_X1Y11_LUT4AB/SS4END[8] Tile_X1Y11_LUT4AB/SS4END[9]
+ Tile_X1Y9_LUT4AB/SS4BEG[0] Tile_X1Y9_LUT4AB/SS4BEG[10] Tile_X1Y9_LUT4AB/SS4BEG[11]
+ Tile_X1Y9_LUT4AB/SS4BEG[12] Tile_X1Y9_LUT4AB/SS4BEG[13] Tile_X1Y9_LUT4AB/SS4BEG[14]
+ Tile_X1Y9_LUT4AB/SS4BEG[15] Tile_X1Y9_LUT4AB/SS4BEG[1] Tile_X1Y9_LUT4AB/SS4BEG[2]
+ Tile_X1Y9_LUT4AB/SS4BEG[3] Tile_X1Y9_LUT4AB/SS4BEG[4] Tile_X1Y9_LUT4AB/SS4BEG[5]
+ Tile_X1Y9_LUT4AB/SS4BEG[6] Tile_X1Y9_LUT4AB/SS4BEG[7] Tile_X1Y9_LUT4AB/SS4BEG[8]
+ Tile_X1Y9_LUT4AB/SS4BEG[9] Tile_X1Y10_LUT4AB/UserCLK Tile_X1Y9_LUT4AB/UserCLK VGND
+ VPWR Tile_X0Y10_W_IO/W1END[0] Tile_X0Y10_W_IO/W1END[1] Tile_X0Y10_W_IO/W1END[2]
+ Tile_X0Y10_W_IO/W1END[3] Tile_X2Y10_LUT4AB/W1BEG[0] Tile_X2Y10_LUT4AB/W1BEG[1] Tile_X2Y10_LUT4AB/W1BEG[2]
+ Tile_X2Y10_LUT4AB/W1BEG[3] Tile_X0Y10_W_IO/W2MID[0] Tile_X0Y10_W_IO/W2MID[1] Tile_X0Y10_W_IO/W2MID[2]
+ Tile_X0Y10_W_IO/W2MID[3] Tile_X0Y10_W_IO/W2MID[4] Tile_X0Y10_W_IO/W2MID[5] Tile_X0Y10_W_IO/W2MID[6]
+ Tile_X0Y10_W_IO/W2MID[7] Tile_X0Y10_W_IO/W2END[0] Tile_X0Y10_W_IO/W2END[1] Tile_X0Y10_W_IO/W2END[2]
+ Tile_X0Y10_W_IO/W2END[3] Tile_X0Y10_W_IO/W2END[4] Tile_X0Y10_W_IO/W2END[5] Tile_X0Y10_W_IO/W2END[6]
+ Tile_X0Y10_W_IO/W2END[7] Tile_X1Y10_LUT4AB/W2END[0] Tile_X1Y10_LUT4AB/W2END[1] Tile_X1Y10_LUT4AB/W2END[2]
+ Tile_X1Y10_LUT4AB/W2END[3] Tile_X1Y10_LUT4AB/W2END[4] Tile_X1Y10_LUT4AB/W2END[5]
+ Tile_X1Y10_LUT4AB/W2END[6] Tile_X1Y10_LUT4AB/W2END[7] Tile_X2Y10_LUT4AB/W2BEG[0]
+ Tile_X2Y10_LUT4AB/W2BEG[1] Tile_X2Y10_LUT4AB/W2BEG[2] Tile_X2Y10_LUT4AB/W2BEG[3]
+ Tile_X2Y10_LUT4AB/W2BEG[4] Tile_X2Y10_LUT4AB/W2BEG[5] Tile_X2Y10_LUT4AB/W2BEG[6]
+ Tile_X2Y10_LUT4AB/W2BEG[7] Tile_X0Y10_W_IO/W6END[0] Tile_X0Y10_W_IO/W6END[10] Tile_X0Y10_W_IO/W6END[11]
+ Tile_X0Y10_W_IO/W6END[1] Tile_X0Y10_W_IO/W6END[2] Tile_X0Y10_W_IO/W6END[3] Tile_X0Y10_W_IO/W6END[4]
+ Tile_X0Y10_W_IO/W6END[5] Tile_X0Y10_W_IO/W6END[6] Tile_X0Y10_W_IO/W6END[7] Tile_X0Y10_W_IO/W6END[8]
+ Tile_X0Y10_W_IO/W6END[9] Tile_X2Y10_LUT4AB/W6BEG[0] Tile_X2Y10_LUT4AB/W6BEG[10]
+ Tile_X2Y10_LUT4AB/W6BEG[11] Tile_X2Y10_LUT4AB/W6BEG[1] Tile_X2Y10_LUT4AB/W6BEG[2]
+ Tile_X2Y10_LUT4AB/W6BEG[3] Tile_X2Y10_LUT4AB/W6BEG[4] Tile_X2Y10_LUT4AB/W6BEG[5]
+ Tile_X2Y10_LUT4AB/W6BEG[6] Tile_X2Y10_LUT4AB/W6BEG[7] Tile_X2Y10_LUT4AB/W6BEG[8]
+ Tile_X2Y10_LUT4AB/W6BEG[9] Tile_X0Y10_W_IO/WW4END[0] Tile_X0Y10_W_IO/WW4END[10]
+ Tile_X0Y10_W_IO/WW4END[11] Tile_X0Y10_W_IO/WW4END[12] Tile_X0Y10_W_IO/WW4END[13]
+ Tile_X0Y10_W_IO/WW4END[14] Tile_X0Y10_W_IO/WW4END[15] Tile_X0Y10_W_IO/WW4END[1]
+ Tile_X0Y10_W_IO/WW4END[2] Tile_X0Y10_W_IO/WW4END[3] Tile_X0Y10_W_IO/WW4END[4] Tile_X0Y10_W_IO/WW4END[5]
+ Tile_X0Y10_W_IO/WW4END[6] Tile_X0Y10_W_IO/WW4END[7] Tile_X0Y10_W_IO/WW4END[8] Tile_X0Y10_W_IO/WW4END[9]
+ Tile_X2Y10_LUT4AB/WW4BEG[0] Tile_X2Y10_LUT4AB/WW4BEG[10] Tile_X2Y10_LUT4AB/WW4BEG[11]
+ Tile_X2Y10_LUT4AB/WW4BEG[12] Tile_X2Y10_LUT4AB/WW4BEG[13] Tile_X2Y10_LUT4AB/WW4BEG[14]
+ Tile_X2Y10_LUT4AB/WW4BEG[15] Tile_X2Y10_LUT4AB/WW4BEG[1] Tile_X2Y10_LUT4AB/WW4BEG[2]
+ Tile_X2Y10_LUT4AB/WW4BEG[3] Tile_X2Y10_LUT4AB/WW4BEG[4] Tile_X2Y10_LUT4AB/WW4BEG[5]
+ Tile_X2Y10_LUT4AB/WW4BEG[6] Tile_X2Y10_LUT4AB/WW4BEG[7] Tile_X2Y10_LUT4AB/WW4BEG[8]
+ Tile_X2Y10_LUT4AB/WW4BEG[9] LUT4AB
XTile_X6Y5_LUT4AB Tile_X6Y6_LUT4AB/Co Tile_X6Y5_LUT4AB/Co Tile_X6Y5_LUT4AB/E1BEG[0]
+ Tile_X6Y5_LUT4AB/E1BEG[1] Tile_X6Y5_LUT4AB/E1BEG[2] Tile_X6Y5_LUT4AB/E1BEG[3] Tile_X6Y5_LUT4AB/E1END[0]
+ Tile_X6Y5_LUT4AB/E1END[1] Tile_X6Y5_LUT4AB/E1END[2] Tile_X6Y5_LUT4AB/E1END[3] Tile_X6Y5_LUT4AB/E2BEG[0]
+ Tile_X6Y5_LUT4AB/E2BEG[1] Tile_X6Y5_LUT4AB/E2BEG[2] Tile_X6Y5_LUT4AB/E2BEG[3] Tile_X6Y5_LUT4AB/E2BEG[4]
+ Tile_X6Y5_LUT4AB/E2BEG[5] Tile_X6Y5_LUT4AB/E2BEG[6] Tile_X6Y5_LUT4AB/E2BEG[7] Tile_X6Y5_LUT4AB/E2BEGb[0]
+ Tile_X6Y5_LUT4AB/E2BEGb[1] Tile_X6Y5_LUT4AB/E2BEGb[2] Tile_X6Y5_LUT4AB/E2BEGb[3]
+ Tile_X6Y5_LUT4AB/E2BEGb[4] Tile_X6Y5_LUT4AB/E2BEGb[5] Tile_X6Y5_LUT4AB/E2BEGb[6]
+ Tile_X6Y5_LUT4AB/E2BEGb[7] Tile_X6Y5_LUT4AB/E2END[0] Tile_X6Y5_LUT4AB/E2END[1] Tile_X6Y5_LUT4AB/E2END[2]
+ Tile_X6Y5_LUT4AB/E2END[3] Tile_X6Y5_LUT4AB/E2END[4] Tile_X6Y5_LUT4AB/E2END[5] Tile_X6Y5_LUT4AB/E2END[6]
+ Tile_X6Y5_LUT4AB/E2END[7] Tile_X6Y5_LUT4AB/E2MID[0] Tile_X6Y5_LUT4AB/E2MID[1] Tile_X6Y5_LUT4AB/E2MID[2]
+ Tile_X6Y5_LUT4AB/E2MID[3] Tile_X6Y5_LUT4AB/E2MID[4] Tile_X6Y5_LUT4AB/E2MID[5] Tile_X6Y5_LUT4AB/E2MID[6]
+ Tile_X6Y5_LUT4AB/E2MID[7] Tile_X6Y5_LUT4AB/E6BEG[0] Tile_X6Y5_LUT4AB/E6BEG[10] Tile_X6Y5_LUT4AB/E6BEG[11]
+ Tile_X6Y5_LUT4AB/E6BEG[1] Tile_X6Y5_LUT4AB/E6BEG[2] Tile_X6Y5_LUT4AB/E6BEG[3] Tile_X6Y5_LUT4AB/E6BEG[4]
+ Tile_X6Y5_LUT4AB/E6BEG[5] Tile_X6Y5_LUT4AB/E6BEG[6] Tile_X6Y5_LUT4AB/E6BEG[7] Tile_X6Y5_LUT4AB/E6BEG[8]
+ Tile_X6Y5_LUT4AB/E6BEG[9] Tile_X6Y5_LUT4AB/E6END[0] Tile_X6Y5_LUT4AB/E6END[10] Tile_X6Y5_LUT4AB/E6END[11]
+ Tile_X6Y5_LUT4AB/E6END[1] Tile_X6Y5_LUT4AB/E6END[2] Tile_X6Y5_LUT4AB/E6END[3] Tile_X6Y5_LUT4AB/E6END[4]
+ Tile_X6Y5_LUT4AB/E6END[5] Tile_X6Y5_LUT4AB/E6END[6] Tile_X6Y5_LUT4AB/E6END[7] Tile_X6Y5_LUT4AB/E6END[8]
+ Tile_X6Y5_LUT4AB/E6END[9] Tile_X6Y5_LUT4AB/EE4BEG[0] Tile_X6Y5_LUT4AB/EE4BEG[10]
+ Tile_X6Y5_LUT4AB/EE4BEG[11] Tile_X6Y5_LUT4AB/EE4BEG[12] Tile_X6Y5_LUT4AB/EE4BEG[13]
+ Tile_X6Y5_LUT4AB/EE4BEG[14] Tile_X6Y5_LUT4AB/EE4BEG[15] Tile_X6Y5_LUT4AB/EE4BEG[1]
+ Tile_X6Y5_LUT4AB/EE4BEG[2] Tile_X6Y5_LUT4AB/EE4BEG[3] Tile_X6Y5_LUT4AB/EE4BEG[4]
+ Tile_X6Y5_LUT4AB/EE4BEG[5] Tile_X6Y5_LUT4AB/EE4BEG[6] Tile_X6Y5_LUT4AB/EE4BEG[7]
+ Tile_X6Y5_LUT4AB/EE4BEG[8] Tile_X6Y5_LUT4AB/EE4BEG[9] Tile_X6Y5_LUT4AB/EE4END[0]
+ Tile_X6Y5_LUT4AB/EE4END[10] Tile_X6Y5_LUT4AB/EE4END[11] Tile_X6Y5_LUT4AB/EE4END[12]
+ Tile_X6Y5_LUT4AB/EE4END[13] Tile_X6Y5_LUT4AB/EE4END[14] Tile_X6Y5_LUT4AB/EE4END[15]
+ Tile_X6Y5_LUT4AB/EE4END[1] Tile_X6Y5_LUT4AB/EE4END[2] Tile_X6Y5_LUT4AB/EE4END[3]
+ Tile_X6Y5_LUT4AB/EE4END[4] Tile_X6Y5_LUT4AB/EE4END[5] Tile_X6Y5_LUT4AB/EE4END[6]
+ Tile_X6Y5_LUT4AB/EE4END[7] Tile_X6Y5_LUT4AB/EE4END[8] Tile_X6Y5_LUT4AB/EE4END[9]
+ Tile_X6Y5_LUT4AB/FrameData[0] Tile_X6Y5_LUT4AB/FrameData[10] Tile_X6Y5_LUT4AB/FrameData[11]
+ Tile_X6Y5_LUT4AB/FrameData[12] Tile_X6Y5_LUT4AB/FrameData[13] Tile_X6Y5_LUT4AB/FrameData[14]
+ Tile_X6Y5_LUT4AB/FrameData[15] Tile_X6Y5_LUT4AB/FrameData[16] Tile_X6Y5_LUT4AB/FrameData[17]
+ Tile_X6Y5_LUT4AB/FrameData[18] Tile_X6Y5_LUT4AB/FrameData[19] Tile_X6Y5_LUT4AB/FrameData[1]
+ Tile_X6Y5_LUT4AB/FrameData[20] Tile_X6Y5_LUT4AB/FrameData[21] Tile_X6Y5_LUT4AB/FrameData[22]
+ Tile_X6Y5_LUT4AB/FrameData[23] Tile_X6Y5_LUT4AB/FrameData[24] Tile_X6Y5_LUT4AB/FrameData[25]
+ Tile_X6Y5_LUT4AB/FrameData[26] Tile_X6Y5_LUT4AB/FrameData[27] Tile_X6Y5_LUT4AB/FrameData[28]
+ Tile_X6Y5_LUT4AB/FrameData[29] Tile_X6Y5_LUT4AB/FrameData[2] Tile_X6Y5_LUT4AB/FrameData[30]
+ Tile_X6Y5_LUT4AB/FrameData[31] Tile_X6Y5_LUT4AB/FrameData[3] Tile_X6Y5_LUT4AB/FrameData[4]
+ Tile_X6Y5_LUT4AB/FrameData[5] Tile_X6Y5_LUT4AB/FrameData[6] Tile_X6Y5_LUT4AB/FrameData[7]
+ Tile_X6Y5_LUT4AB/FrameData[8] Tile_X6Y5_LUT4AB/FrameData[9] Tile_X6Y5_LUT4AB/FrameData_O[0]
+ Tile_X6Y5_LUT4AB/FrameData_O[10] Tile_X6Y5_LUT4AB/FrameData_O[11] Tile_X6Y5_LUT4AB/FrameData_O[12]
+ Tile_X6Y5_LUT4AB/FrameData_O[13] Tile_X6Y5_LUT4AB/FrameData_O[14] Tile_X6Y5_LUT4AB/FrameData_O[15]
+ Tile_X6Y5_LUT4AB/FrameData_O[16] Tile_X6Y5_LUT4AB/FrameData_O[17] Tile_X6Y5_LUT4AB/FrameData_O[18]
+ Tile_X6Y5_LUT4AB/FrameData_O[19] Tile_X6Y5_LUT4AB/FrameData_O[1] Tile_X6Y5_LUT4AB/FrameData_O[20]
+ Tile_X6Y5_LUT4AB/FrameData_O[21] Tile_X6Y5_LUT4AB/FrameData_O[22] Tile_X6Y5_LUT4AB/FrameData_O[23]
+ Tile_X6Y5_LUT4AB/FrameData_O[24] Tile_X6Y5_LUT4AB/FrameData_O[25] Tile_X6Y5_LUT4AB/FrameData_O[26]
+ Tile_X6Y5_LUT4AB/FrameData_O[27] Tile_X6Y5_LUT4AB/FrameData_O[28] Tile_X6Y5_LUT4AB/FrameData_O[29]
+ Tile_X6Y5_LUT4AB/FrameData_O[2] Tile_X6Y5_LUT4AB/FrameData_O[30] Tile_X6Y5_LUT4AB/FrameData_O[31]
+ Tile_X6Y5_LUT4AB/FrameData_O[3] Tile_X6Y5_LUT4AB/FrameData_O[4] Tile_X6Y5_LUT4AB/FrameData_O[5]
+ Tile_X6Y5_LUT4AB/FrameData_O[6] Tile_X6Y5_LUT4AB/FrameData_O[7] Tile_X6Y5_LUT4AB/FrameData_O[8]
+ Tile_X6Y5_LUT4AB/FrameData_O[9] Tile_X6Y5_LUT4AB/FrameStrobe[0] Tile_X6Y5_LUT4AB/FrameStrobe[10]
+ Tile_X6Y5_LUT4AB/FrameStrobe[11] Tile_X6Y5_LUT4AB/FrameStrobe[12] Tile_X6Y5_LUT4AB/FrameStrobe[13]
+ Tile_X6Y5_LUT4AB/FrameStrobe[14] Tile_X6Y5_LUT4AB/FrameStrobe[15] Tile_X6Y5_LUT4AB/FrameStrobe[16]
+ Tile_X6Y5_LUT4AB/FrameStrobe[17] Tile_X6Y5_LUT4AB/FrameStrobe[18] Tile_X6Y5_LUT4AB/FrameStrobe[19]
+ Tile_X6Y5_LUT4AB/FrameStrobe[1] Tile_X6Y5_LUT4AB/FrameStrobe[2] Tile_X6Y5_LUT4AB/FrameStrobe[3]
+ Tile_X6Y5_LUT4AB/FrameStrobe[4] Tile_X6Y5_LUT4AB/FrameStrobe[5] Tile_X6Y5_LUT4AB/FrameStrobe[6]
+ Tile_X6Y5_LUT4AB/FrameStrobe[7] Tile_X6Y5_LUT4AB/FrameStrobe[8] Tile_X6Y5_LUT4AB/FrameStrobe[9]
+ Tile_X6Y4_LUT4AB/FrameStrobe[0] Tile_X6Y4_LUT4AB/FrameStrobe[10] Tile_X6Y4_LUT4AB/FrameStrobe[11]
+ Tile_X6Y4_LUT4AB/FrameStrobe[12] Tile_X6Y4_LUT4AB/FrameStrobe[13] Tile_X6Y4_LUT4AB/FrameStrobe[14]
+ Tile_X6Y4_LUT4AB/FrameStrobe[15] Tile_X6Y4_LUT4AB/FrameStrobe[16] Tile_X6Y4_LUT4AB/FrameStrobe[17]
+ Tile_X6Y4_LUT4AB/FrameStrobe[18] Tile_X6Y4_LUT4AB/FrameStrobe[19] Tile_X6Y4_LUT4AB/FrameStrobe[1]
+ Tile_X6Y4_LUT4AB/FrameStrobe[2] Tile_X6Y4_LUT4AB/FrameStrobe[3] Tile_X6Y4_LUT4AB/FrameStrobe[4]
+ Tile_X6Y4_LUT4AB/FrameStrobe[5] Tile_X6Y4_LUT4AB/FrameStrobe[6] Tile_X6Y4_LUT4AB/FrameStrobe[7]
+ Tile_X6Y4_LUT4AB/FrameStrobe[8] Tile_X6Y4_LUT4AB/FrameStrobe[9] Tile_X6Y5_LUT4AB/N1BEG[0]
+ Tile_X6Y5_LUT4AB/N1BEG[1] Tile_X6Y5_LUT4AB/N1BEG[2] Tile_X6Y5_LUT4AB/N1BEG[3] Tile_X6Y6_LUT4AB/N1BEG[0]
+ Tile_X6Y6_LUT4AB/N1BEG[1] Tile_X6Y6_LUT4AB/N1BEG[2] Tile_X6Y6_LUT4AB/N1BEG[3] Tile_X6Y5_LUT4AB/N2BEG[0]
+ Tile_X6Y5_LUT4AB/N2BEG[1] Tile_X6Y5_LUT4AB/N2BEG[2] Tile_X6Y5_LUT4AB/N2BEG[3] Tile_X6Y5_LUT4AB/N2BEG[4]
+ Tile_X6Y5_LUT4AB/N2BEG[5] Tile_X6Y5_LUT4AB/N2BEG[6] Tile_X6Y5_LUT4AB/N2BEG[7] Tile_X6Y4_LUT4AB/N2END[0]
+ Tile_X6Y4_LUT4AB/N2END[1] Tile_X6Y4_LUT4AB/N2END[2] Tile_X6Y4_LUT4AB/N2END[3] Tile_X6Y4_LUT4AB/N2END[4]
+ Tile_X6Y4_LUT4AB/N2END[5] Tile_X6Y4_LUT4AB/N2END[6] Tile_X6Y4_LUT4AB/N2END[7] Tile_X6Y5_LUT4AB/N2END[0]
+ Tile_X6Y5_LUT4AB/N2END[1] Tile_X6Y5_LUT4AB/N2END[2] Tile_X6Y5_LUT4AB/N2END[3] Tile_X6Y5_LUT4AB/N2END[4]
+ Tile_X6Y5_LUT4AB/N2END[5] Tile_X6Y5_LUT4AB/N2END[6] Tile_X6Y5_LUT4AB/N2END[7] Tile_X6Y6_LUT4AB/N2BEG[0]
+ Tile_X6Y6_LUT4AB/N2BEG[1] Tile_X6Y6_LUT4AB/N2BEG[2] Tile_X6Y6_LUT4AB/N2BEG[3] Tile_X6Y6_LUT4AB/N2BEG[4]
+ Tile_X6Y6_LUT4AB/N2BEG[5] Tile_X6Y6_LUT4AB/N2BEG[6] Tile_X6Y6_LUT4AB/N2BEG[7] Tile_X6Y5_LUT4AB/N4BEG[0]
+ Tile_X6Y5_LUT4AB/N4BEG[10] Tile_X6Y5_LUT4AB/N4BEG[11] Tile_X6Y5_LUT4AB/N4BEG[12]
+ Tile_X6Y5_LUT4AB/N4BEG[13] Tile_X6Y5_LUT4AB/N4BEG[14] Tile_X6Y5_LUT4AB/N4BEG[15]
+ Tile_X6Y5_LUT4AB/N4BEG[1] Tile_X6Y5_LUT4AB/N4BEG[2] Tile_X6Y5_LUT4AB/N4BEG[3] Tile_X6Y5_LUT4AB/N4BEG[4]
+ Tile_X6Y5_LUT4AB/N4BEG[5] Tile_X6Y5_LUT4AB/N4BEG[6] Tile_X6Y5_LUT4AB/N4BEG[7] Tile_X6Y5_LUT4AB/N4BEG[8]
+ Tile_X6Y5_LUT4AB/N4BEG[9] Tile_X6Y6_LUT4AB/N4BEG[0] Tile_X6Y6_LUT4AB/N4BEG[10] Tile_X6Y6_LUT4AB/N4BEG[11]
+ Tile_X6Y6_LUT4AB/N4BEG[12] Tile_X6Y6_LUT4AB/N4BEG[13] Tile_X6Y6_LUT4AB/N4BEG[14]
+ Tile_X6Y6_LUT4AB/N4BEG[15] Tile_X6Y6_LUT4AB/N4BEG[1] Tile_X6Y6_LUT4AB/N4BEG[2] Tile_X6Y6_LUT4AB/N4BEG[3]
+ Tile_X6Y6_LUT4AB/N4BEG[4] Tile_X6Y6_LUT4AB/N4BEG[5] Tile_X6Y6_LUT4AB/N4BEG[6] Tile_X6Y6_LUT4AB/N4BEG[7]
+ Tile_X6Y6_LUT4AB/N4BEG[8] Tile_X6Y6_LUT4AB/N4BEG[9] Tile_X6Y5_LUT4AB/NN4BEG[0] Tile_X6Y5_LUT4AB/NN4BEG[10]
+ Tile_X6Y5_LUT4AB/NN4BEG[11] Tile_X6Y5_LUT4AB/NN4BEG[12] Tile_X6Y5_LUT4AB/NN4BEG[13]
+ Tile_X6Y5_LUT4AB/NN4BEG[14] Tile_X6Y5_LUT4AB/NN4BEG[15] Tile_X6Y5_LUT4AB/NN4BEG[1]
+ Tile_X6Y5_LUT4AB/NN4BEG[2] Tile_X6Y5_LUT4AB/NN4BEG[3] Tile_X6Y5_LUT4AB/NN4BEG[4]
+ Tile_X6Y5_LUT4AB/NN4BEG[5] Tile_X6Y5_LUT4AB/NN4BEG[6] Tile_X6Y5_LUT4AB/NN4BEG[7]
+ Tile_X6Y5_LUT4AB/NN4BEG[8] Tile_X6Y5_LUT4AB/NN4BEG[9] Tile_X6Y6_LUT4AB/NN4BEG[0]
+ Tile_X6Y6_LUT4AB/NN4BEG[10] Tile_X6Y6_LUT4AB/NN4BEG[11] Tile_X6Y6_LUT4AB/NN4BEG[12]
+ Tile_X6Y6_LUT4AB/NN4BEG[13] Tile_X6Y6_LUT4AB/NN4BEG[14] Tile_X6Y6_LUT4AB/NN4BEG[15]
+ Tile_X6Y6_LUT4AB/NN4BEG[1] Tile_X6Y6_LUT4AB/NN4BEG[2] Tile_X6Y6_LUT4AB/NN4BEG[3]
+ Tile_X6Y6_LUT4AB/NN4BEG[4] Tile_X6Y6_LUT4AB/NN4BEG[5] Tile_X6Y6_LUT4AB/NN4BEG[6]
+ Tile_X6Y6_LUT4AB/NN4BEG[7] Tile_X6Y6_LUT4AB/NN4BEG[8] Tile_X6Y6_LUT4AB/NN4BEG[9]
+ Tile_X6Y6_LUT4AB/S1END[0] Tile_X6Y6_LUT4AB/S1END[1] Tile_X6Y6_LUT4AB/S1END[2] Tile_X6Y6_LUT4AB/S1END[3]
+ Tile_X6Y5_LUT4AB/S1END[0] Tile_X6Y5_LUT4AB/S1END[1] Tile_X6Y5_LUT4AB/S1END[2] Tile_X6Y5_LUT4AB/S1END[3]
+ Tile_X6Y6_LUT4AB/S2MID[0] Tile_X6Y6_LUT4AB/S2MID[1] Tile_X6Y6_LUT4AB/S2MID[2] Tile_X6Y6_LUT4AB/S2MID[3]
+ Tile_X6Y6_LUT4AB/S2MID[4] Tile_X6Y6_LUT4AB/S2MID[5] Tile_X6Y6_LUT4AB/S2MID[6] Tile_X6Y6_LUT4AB/S2MID[7]
+ Tile_X6Y6_LUT4AB/S2END[0] Tile_X6Y6_LUT4AB/S2END[1] Tile_X6Y6_LUT4AB/S2END[2] Tile_X6Y6_LUT4AB/S2END[3]
+ Tile_X6Y6_LUT4AB/S2END[4] Tile_X6Y6_LUT4AB/S2END[5] Tile_X6Y6_LUT4AB/S2END[6] Tile_X6Y6_LUT4AB/S2END[7]
+ Tile_X6Y5_LUT4AB/S2END[0] Tile_X6Y5_LUT4AB/S2END[1] Tile_X6Y5_LUT4AB/S2END[2] Tile_X6Y5_LUT4AB/S2END[3]
+ Tile_X6Y5_LUT4AB/S2END[4] Tile_X6Y5_LUT4AB/S2END[5] Tile_X6Y5_LUT4AB/S2END[6] Tile_X6Y5_LUT4AB/S2END[7]
+ Tile_X6Y5_LUT4AB/S2MID[0] Tile_X6Y5_LUT4AB/S2MID[1] Tile_X6Y5_LUT4AB/S2MID[2] Tile_X6Y5_LUT4AB/S2MID[3]
+ Tile_X6Y5_LUT4AB/S2MID[4] Tile_X6Y5_LUT4AB/S2MID[5] Tile_X6Y5_LUT4AB/S2MID[6] Tile_X6Y5_LUT4AB/S2MID[7]
+ Tile_X6Y6_LUT4AB/S4END[0] Tile_X6Y6_LUT4AB/S4END[10] Tile_X6Y6_LUT4AB/S4END[11]
+ Tile_X6Y6_LUT4AB/S4END[12] Tile_X6Y6_LUT4AB/S4END[13] Tile_X6Y6_LUT4AB/S4END[14]
+ Tile_X6Y6_LUT4AB/S4END[15] Tile_X6Y6_LUT4AB/S4END[1] Tile_X6Y6_LUT4AB/S4END[2] Tile_X6Y6_LUT4AB/S4END[3]
+ Tile_X6Y6_LUT4AB/S4END[4] Tile_X6Y6_LUT4AB/S4END[5] Tile_X6Y6_LUT4AB/S4END[6] Tile_X6Y6_LUT4AB/S4END[7]
+ Tile_X6Y6_LUT4AB/S4END[8] Tile_X6Y6_LUT4AB/S4END[9] Tile_X6Y5_LUT4AB/S4END[0] Tile_X6Y5_LUT4AB/S4END[10]
+ Tile_X6Y5_LUT4AB/S4END[11] Tile_X6Y5_LUT4AB/S4END[12] Tile_X6Y5_LUT4AB/S4END[13]
+ Tile_X6Y5_LUT4AB/S4END[14] Tile_X6Y5_LUT4AB/S4END[15] Tile_X6Y5_LUT4AB/S4END[1]
+ Tile_X6Y5_LUT4AB/S4END[2] Tile_X6Y5_LUT4AB/S4END[3] Tile_X6Y5_LUT4AB/S4END[4] Tile_X6Y5_LUT4AB/S4END[5]
+ Tile_X6Y5_LUT4AB/S4END[6] Tile_X6Y5_LUT4AB/S4END[7] Tile_X6Y5_LUT4AB/S4END[8] Tile_X6Y5_LUT4AB/S4END[9]
+ Tile_X6Y6_LUT4AB/SS4END[0] Tile_X6Y6_LUT4AB/SS4END[10] Tile_X6Y6_LUT4AB/SS4END[11]
+ Tile_X6Y6_LUT4AB/SS4END[12] Tile_X6Y6_LUT4AB/SS4END[13] Tile_X6Y6_LUT4AB/SS4END[14]
+ Tile_X6Y6_LUT4AB/SS4END[15] Tile_X6Y6_LUT4AB/SS4END[1] Tile_X6Y6_LUT4AB/SS4END[2]
+ Tile_X6Y6_LUT4AB/SS4END[3] Tile_X6Y6_LUT4AB/SS4END[4] Tile_X6Y6_LUT4AB/SS4END[5]
+ Tile_X6Y6_LUT4AB/SS4END[6] Tile_X6Y6_LUT4AB/SS4END[7] Tile_X6Y6_LUT4AB/SS4END[8]
+ Tile_X6Y6_LUT4AB/SS4END[9] Tile_X6Y5_LUT4AB/SS4END[0] Tile_X6Y5_LUT4AB/SS4END[10]
+ Tile_X6Y5_LUT4AB/SS4END[11] Tile_X6Y5_LUT4AB/SS4END[12] Tile_X6Y5_LUT4AB/SS4END[13]
+ Tile_X6Y5_LUT4AB/SS4END[14] Tile_X6Y5_LUT4AB/SS4END[15] Tile_X6Y5_LUT4AB/SS4END[1]
+ Tile_X6Y5_LUT4AB/SS4END[2] Tile_X6Y5_LUT4AB/SS4END[3] Tile_X6Y5_LUT4AB/SS4END[4]
+ Tile_X6Y5_LUT4AB/SS4END[5] Tile_X6Y5_LUT4AB/SS4END[6] Tile_X6Y5_LUT4AB/SS4END[7]
+ Tile_X6Y5_LUT4AB/SS4END[8] Tile_X6Y5_LUT4AB/SS4END[9] Tile_X6Y5_LUT4AB/UserCLK Tile_X6Y4_LUT4AB/UserCLK
+ VGND VPWR Tile_X6Y5_LUT4AB/W1BEG[0] Tile_X6Y5_LUT4AB/W1BEG[1] Tile_X6Y5_LUT4AB/W1BEG[2]
+ Tile_X6Y5_LUT4AB/W1BEG[3] Tile_X6Y5_LUT4AB/W1END[0] Tile_X6Y5_LUT4AB/W1END[1] Tile_X6Y5_LUT4AB/W1END[2]
+ Tile_X6Y5_LUT4AB/W1END[3] Tile_X6Y5_LUT4AB/W2BEG[0] Tile_X6Y5_LUT4AB/W2BEG[1] Tile_X6Y5_LUT4AB/W2BEG[2]
+ Tile_X6Y5_LUT4AB/W2BEG[3] Tile_X6Y5_LUT4AB/W2BEG[4] Tile_X6Y5_LUT4AB/W2BEG[5] Tile_X6Y5_LUT4AB/W2BEG[6]
+ Tile_X6Y5_LUT4AB/W2BEG[7] Tile_X5Y5_LUT4AB/W2END[0] Tile_X5Y5_LUT4AB/W2END[1] Tile_X5Y5_LUT4AB/W2END[2]
+ Tile_X5Y5_LUT4AB/W2END[3] Tile_X5Y5_LUT4AB/W2END[4] Tile_X5Y5_LUT4AB/W2END[5] Tile_X5Y5_LUT4AB/W2END[6]
+ Tile_X5Y5_LUT4AB/W2END[7] Tile_X6Y5_LUT4AB/W2END[0] Tile_X6Y5_LUT4AB/W2END[1] Tile_X6Y5_LUT4AB/W2END[2]
+ Tile_X6Y5_LUT4AB/W2END[3] Tile_X6Y5_LUT4AB/W2END[4] Tile_X6Y5_LUT4AB/W2END[5] Tile_X6Y5_LUT4AB/W2END[6]
+ Tile_X6Y5_LUT4AB/W2END[7] Tile_X6Y5_LUT4AB/W2MID[0] Tile_X6Y5_LUT4AB/W2MID[1] Tile_X6Y5_LUT4AB/W2MID[2]
+ Tile_X6Y5_LUT4AB/W2MID[3] Tile_X6Y5_LUT4AB/W2MID[4] Tile_X6Y5_LUT4AB/W2MID[5] Tile_X6Y5_LUT4AB/W2MID[6]
+ Tile_X6Y5_LUT4AB/W2MID[7] Tile_X6Y5_LUT4AB/W6BEG[0] Tile_X6Y5_LUT4AB/W6BEG[10] Tile_X6Y5_LUT4AB/W6BEG[11]
+ Tile_X6Y5_LUT4AB/W6BEG[1] Tile_X6Y5_LUT4AB/W6BEG[2] Tile_X6Y5_LUT4AB/W6BEG[3] Tile_X6Y5_LUT4AB/W6BEG[4]
+ Tile_X6Y5_LUT4AB/W6BEG[5] Tile_X6Y5_LUT4AB/W6BEG[6] Tile_X6Y5_LUT4AB/W6BEG[7] Tile_X6Y5_LUT4AB/W6BEG[8]
+ Tile_X6Y5_LUT4AB/W6BEG[9] Tile_X6Y5_LUT4AB/W6END[0] Tile_X6Y5_LUT4AB/W6END[10] Tile_X6Y5_LUT4AB/W6END[11]
+ Tile_X6Y5_LUT4AB/W6END[1] Tile_X6Y5_LUT4AB/W6END[2] Tile_X6Y5_LUT4AB/W6END[3] Tile_X6Y5_LUT4AB/W6END[4]
+ Tile_X6Y5_LUT4AB/W6END[5] Tile_X6Y5_LUT4AB/W6END[6] Tile_X6Y5_LUT4AB/W6END[7] Tile_X6Y5_LUT4AB/W6END[8]
+ Tile_X6Y5_LUT4AB/W6END[9] Tile_X6Y5_LUT4AB/WW4BEG[0] Tile_X6Y5_LUT4AB/WW4BEG[10]
+ Tile_X6Y5_LUT4AB/WW4BEG[11] Tile_X6Y5_LUT4AB/WW4BEG[12] Tile_X6Y5_LUT4AB/WW4BEG[13]
+ Tile_X6Y5_LUT4AB/WW4BEG[14] Tile_X6Y5_LUT4AB/WW4BEG[15] Tile_X6Y5_LUT4AB/WW4BEG[1]
+ Tile_X6Y5_LUT4AB/WW4BEG[2] Tile_X6Y5_LUT4AB/WW4BEG[3] Tile_X6Y5_LUT4AB/WW4BEG[4]
+ Tile_X6Y5_LUT4AB/WW4BEG[5] Tile_X6Y5_LUT4AB/WW4BEG[6] Tile_X6Y5_LUT4AB/WW4BEG[7]
+ Tile_X6Y5_LUT4AB/WW4BEG[8] Tile_X6Y5_LUT4AB/WW4BEG[9] Tile_X6Y5_LUT4AB/WW4END[0]
+ Tile_X6Y5_LUT4AB/WW4END[10] Tile_X6Y5_LUT4AB/WW4END[11] Tile_X6Y5_LUT4AB/WW4END[12]
+ Tile_X6Y5_LUT4AB/WW4END[13] Tile_X6Y5_LUT4AB/WW4END[14] Tile_X6Y5_LUT4AB/WW4END[15]
+ Tile_X6Y5_LUT4AB/WW4END[1] Tile_X6Y5_LUT4AB/WW4END[2] Tile_X6Y5_LUT4AB/WW4END[3]
+ Tile_X6Y5_LUT4AB/WW4END[4] Tile_X6Y5_LUT4AB/WW4END[5] Tile_X6Y5_LUT4AB/WW4END[6]
+ Tile_X6Y5_LUT4AB/WW4END[7] Tile_X6Y5_LUT4AB/WW4END[8] Tile_X6Y5_LUT4AB/WW4END[9]
+ LUT4AB
XTile_X8Y14_LUT4AB Tile_X8Y14_LUT4AB/Ci Tile_X8Y14_LUT4AB/Co Tile_X9Y14_LUT4AB/E1END[0]
+ Tile_X9Y14_LUT4AB/E1END[1] Tile_X9Y14_LUT4AB/E1END[2] Tile_X9Y14_LUT4AB/E1END[3]
+ Tile_X8Y14_LUT4AB/E1END[0] Tile_X8Y14_LUT4AB/E1END[1] Tile_X8Y14_LUT4AB/E1END[2]
+ Tile_X8Y14_LUT4AB/E1END[3] Tile_X9Y14_LUT4AB/E2MID[0] Tile_X9Y14_LUT4AB/E2MID[1]
+ Tile_X9Y14_LUT4AB/E2MID[2] Tile_X9Y14_LUT4AB/E2MID[3] Tile_X9Y14_LUT4AB/E2MID[4]
+ Tile_X9Y14_LUT4AB/E2MID[5] Tile_X9Y14_LUT4AB/E2MID[6] Tile_X9Y14_LUT4AB/E2MID[7]
+ Tile_X9Y14_LUT4AB/E2END[0] Tile_X9Y14_LUT4AB/E2END[1] Tile_X9Y14_LUT4AB/E2END[2]
+ Tile_X9Y14_LUT4AB/E2END[3] Tile_X9Y14_LUT4AB/E2END[4] Tile_X9Y14_LUT4AB/E2END[5]
+ Tile_X9Y14_LUT4AB/E2END[6] Tile_X9Y14_LUT4AB/E2END[7] Tile_X8Y14_LUT4AB/E2END[0]
+ Tile_X8Y14_LUT4AB/E2END[1] Tile_X8Y14_LUT4AB/E2END[2] Tile_X8Y14_LUT4AB/E2END[3]
+ Tile_X8Y14_LUT4AB/E2END[4] Tile_X8Y14_LUT4AB/E2END[5] Tile_X8Y14_LUT4AB/E2END[6]
+ Tile_X8Y14_LUT4AB/E2END[7] Tile_X8Y14_LUT4AB/E2MID[0] Tile_X8Y14_LUT4AB/E2MID[1]
+ Tile_X8Y14_LUT4AB/E2MID[2] Tile_X8Y14_LUT4AB/E2MID[3] Tile_X8Y14_LUT4AB/E2MID[4]
+ Tile_X8Y14_LUT4AB/E2MID[5] Tile_X8Y14_LUT4AB/E2MID[6] Tile_X8Y14_LUT4AB/E2MID[7]
+ Tile_X9Y14_LUT4AB/E6END[0] Tile_X9Y14_LUT4AB/E6END[10] Tile_X9Y14_LUT4AB/E6END[11]
+ Tile_X9Y14_LUT4AB/E6END[1] Tile_X9Y14_LUT4AB/E6END[2] Tile_X9Y14_LUT4AB/E6END[3]
+ Tile_X9Y14_LUT4AB/E6END[4] Tile_X9Y14_LUT4AB/E6END[5] Tile_X9Y14_LUT4AB/E6END[6]
+ Tile_X9Y14_LUT4AB/E6END[7] Tile_X9Y14_LUT4AB/E6END[8] Tile_X9Y14_LUT4AB/E6END[9]
+ Tile_X8Y14_LUT4AB/E6END[0] Tile_X8Y14_LUT4AB/E6END[10] Tile_X8Y14_LUT4AB/E6END[11]
+ Tile_X8Y14_LUT4AB/E6END[1] Tile_X8Y14_LUT4AB/E6END[2] Tile_X8Y14_LUT4AB/E6END[3]
+ Tile_X8Y14_LUT4AB/E6END[4] Tile_X8Y14_LUT4AB/E6END[5] Tile_X8Y14_LUT4AB/E6END[6]
+ Tile_X8Y14_LUT4AB/E6END[7] Tile_X8Y14_LUT4AB/E6END[8] Tile_X8Y14_LUT4AB/E6END[9]
+ Tile_X9Y14_LUT4AB/EE4END[0] Tile_X9Y14_LUT4AB/EE4END[10] Tile_X9Y14_LUT4AB/EE4END[11]
+ Tile_X9Y14_LUT4AB/EE4END[12] Tile_X9Y14_LUT4AB/EE4END[13] Tile_X9Y14_LUT4AB/EE4END[14]
+ Tile_X9Y14_LUT4AB/EE4END[15] Tile_X9Y14_LUT4AB/EE4END[1] Tile_X9Y14_LUT4AB/EE4END[2]
+ Tile_X9Y14_LUT4AB/EE4END[3] Tile_X9Y14_LUT4AB/EE4END[4] Tile_X9Y14_LUT4AB/EE4END[5]
+ Tile_X9Y14_LUT4AB/EE4END[6] Tile_X9Y14_LUT4AB/EE4END[7] Tile_X9Y14_LUT4AB/EE4END[8]
+ Tile_X9Y14_LUT4AB/EE4END[9] Tile_X8Y14_LUT4AB/EE4END[0] Tile_X8Y14_LUT4AB/EE4END[10]
+ Tile_X8Y14_LUT4AB/EE4END[11] Tile_X8Y14_LUT4AB/EE4END[12] Tile_X8Y14_LUT4AB/EE4END[13]
+ Tile_X8Y14_LUT4AB/EE4END[14] Tile_X8Y14_LUT4AB/EE4END[15] Tile_X8Y14_LUT4AB/EE4END[1]
+ Tile_X8Y14_LUT4AB/EE4END[2] Tile_X8Y14_LUT4AB/EE4END[3] Tile_X8Y14_LUT4AB/EE4END[4]
+ Tile_X8Y14_LUT4AB/EE4END[5] Tile_X8Y14_LUT4AB/EE4END[6] Tile_X8Y14_LUT4AB/EE4END[7]
+ Tile_X8Y14_LUT4AB/EE4END[8] Tile_X8Y14_LUT4AB/EE4END[9] Tile_X8Y14_LUT4AB/FrameData[0]
+ Tile_X8Y14_LUT4AB/FrameData[10] Tile_X8Y14_LUT4AB/FrameData[11] Tile_X8Y14_LUT4AB/FrameData[12]
+ Tile_X8Y14_LUT4AB/FrameData[13] Tile_X8Y14_LUT4AB/FrameData[14] Tile_X8Y14_LUT4AB/FrameData[15]
+ Tile_X8Y14_LUT4AB/FrameData[16] Tile_X8Y14_LUT4AB/FrameData[17] Tile_X8Y14_LUT4AB/FrameData[18]
+ Tile_X8Y14_LUT4AB/FrameData[19] Tile_X8Y14_LUT4AB/FrameData[1] Tile_X8Y14_LUT4AB/FrameData[20]
+ Tile_X8Y14_LUT4AB/FrameData[21] Tile_X8Y14_LUT4AB/FrameData[22] Tile_X8Y14_LUT4AB/FrameData[23]
+ Tile_X8Y14_LUT4AB/FrameData[24] Tile_X8Y14_LUT4AB/FrameData[25] Tile_X8Y14_LUT4AB/FrameData[26]
+ Tile_X8Y14_LUT4AB/FrameData[27] Tile_X8Y14_LUT4AB/FrameData[28] Tile_X8Y14_LUT4AB/FrameData[29]
+ Tile_X8Y14_LUT4AB/FrameData[2] Tile_X8Y14_LUT4AB/FrameData[30] Tile_X8Y14_LUT4AB/FrameData[31]
+ Tile_X8Y14_LUT4AB/FrameData[3] Tile_X8Y14_LUT4AB/FrameData[4] Tile_X8Y14_LUT4AB/FrameData[5]
+ Tile_X8Y14_LUT4AB/FrameData[6] Tile_X8Y14_LUT4AB/FrameData[7] Tile_X8Y14_LUT4AB/FrameData[8]
+ Tile_X8Y14_LUT4AB/FrameData[9] Tile_X9Y14_LUT4AB/FrameData[0] Tile_X9Y14_LUT4AB/FrameData[10]
+ Tile_X9Y14_LUT4AB/FrameData[11] Tile_X9Y14_LUT4AB/FrameData[12] Tile_X9Y14_LUT4AB/FrameData[13]
+ Tile_X9Y14_LUT4AB/FrameData[14] Tile_X9Y14_LUT4AB/FrameData[15] Tile_X9Y14_LUT4AB/FrameData[16]
+ Tile_X9Y14_LUT4AB/FrameData[17] Tile_X9Y14_LUT4AB/FrameData[18] Tile_X9Y14_LUT4AB/FrameData[19]
+ Tile_X9Y14_LUT4AB/FrameData[1] Tile_X9Y14_LUT4AB/FrameData[20] Tile_X9Y14_LUT4AB/FrameData[21]
+ Tile_X9Y14_LUT4AB/FrameData[22] Tile_X9Y14_LUT4AB/FrameData[23] Tile_X9Y14_LUT4AB/FrameData[24]
+ Tile_X9Y14_LUT4AB/FrameData[25] Tile_X9Y14_LUT4AB/FrameData[26] Tile_X9Y14_LUT4AB/FrameData[27]
+ Tile_X9Y14_LUT4AB/FrameData[28] Tile_X9Y14_LUT4AB/FrameData[29] Tile_X9Y14_LUT4AB/FrameData[2]
+ Tile_X9Y14_LUT4AB/FrameData[30] Tile_X9Y14_LUT4AB/FrameData[31] Tile_X9Y14_LUT4AB/FrameData[3]
+ Tile_X9Y14_LUT4AB/FrameData[4] Tile_X9Y14_LUT4AB/FrameData[5] Tile_X9Y14_LUT4AB/FrameData[6]
+ Tile_X9Y14_LUT4AB/FrameData[7] Tile_X9Y14_LUT4AB/FrameData[8] Tile_X9Y14_LUT4AB/FrameData[9]
+ Tile_X8Y14_LUT4AB/FrameStrobe[0] Tile_X8Y14_LUT4AB/FrameStrobe[10] Tile_X8Y14_LUT4AB/FrameStrobe[11]
+ Tile_X8Y14_LUT4AB/FrameStrobe[12] Tile_X8Y14_LUT4AB/FrameStrobe[13] Tile_X8Y14_LUT4AB/FrameStrobe[14]
+ Tile_X8Y14_LUT4AB/FrameStrobe[15] Tile_X8Y14_LUT4AB/FrameStrobe[16] Tile_X8Y14_LUT4AB/FrameStrobe[17]
+ Tile_X8Y14_LUT4AB/FrameStrobe[18] Tile_X8Y14_LUT4AB/FrameStrobe[19] Tile_X8Y14_LUT4AB/FrameStrobe[1]
+ Tile_X8Y14_LUT4AB/FrameStrobe[2] Tile_X8Y14_LUT4AB/FrameStrobe[3] Tile_X8Y14_LUT4AB/FrameStrobe[4]
+ Tile_X8Y14_LUT4AB/FrameStrobe[5] Tile_X8Y14_LUT4AB/FrameStrobe[6] Tile_X8Y14_LUT4AB/FrameStrobe[7]
+ Tile_X8Y14_LUT4AB/FrameStrobe[8] Tile_X8Y14_LUT4AB/FrameStrobe[9] Tile_X8Y13_LUT4AB/FrameStrobe[0]
+ Tile_X8Y13_LUT4AB/FrameStrobe[10] Tile_X8Y13_LUT4AB/FrameStrobe[11] Tile_X8Y13_LUT4AB/FrameStrobe[12]
+ Tile_X8Y13_LUT4AB/FrameStrobe[13] Tile_X8Y13_LUT4AB/FrameStrobe[14] Tile_X8Y13_LUT4AB/FrameStrobe[15]
+ Tile_X8Y13_LUT4AB/FrameStrobe[16] Tile_X8Y13_LUT4AB/FrameStrobe[17] Tile_X8Y13_LUT4AB/FrameStrobe[18]
+ Tile_X8Y13_LUT4AB/FrameStrobe[19] Tile_X8Y13_LUT4AB/FrameStrobe[1] Tile_X8Y13_LUT4AB/FrameStrobe[2]
+ Tile_X8Y13_LUT4AB/FrameStrobe[3] Tile_X8Y13_LUT4AB/FrameStrobe[4] Tile_X8Y13_LUT4AB/FrameStrobe[5]
+ Tile_X8Y13_LUT4AB/FrameStrobe[6] Tile_X8Y13_LUT4AB/FrameStrobe[7] Tile_X8Y13_LUT4AB/FrameStrobe[8]
+ Tile_X8Y13_LUT4AB/FrameStrobe[9] Tile_X8Y14_LUT4AB/N1BEG[0] Tile_X8Y14_LUT4AB/N1BEG[1]
+ Tile_X8Y14_LUT4AB/N1BEG[2] Tile_X8Y14_LUT4AB/N1BEG[3] Tile_X8Y14_LUT4AB/N1END[0]
+ Tile_X8Y14_LUT4AB/N1END[1] Tile_X8Y14_LUT4AB/N1END[2] Tile_X8Y14_LUT4AB/N1END[3]
+ Tile_X8Y14_LUT4AB/N2BEG[0] Tile_X8Y14_LUT4AB/N2BEG[1] Tile_X8Y14_LUT4AB/N2BEG[2]
+ Tile_X8Y14_LUT4AB/N2BEG[3] Tile_X8Y14_LUT4AB/N2BEG[4] Tile_X8Y14_LUT4AB/N2BEG[5]
+ Tile_X8Y14_LUT4AB/N2BEG[6] Tile_X8Y14_LUT4AB/N2BEG[7] Tile_X8Y13_LUT4AB/N2END[0]
+ Tile_X8Y13_LUT4AB/N2END[1] Tile_X8Y13_LUT4AB/N2END[2] Tile_X8Y13_LUT4AB/N2END[3]
+ Tile_X8Y13_LUT4AB/N2END[4] Tile_X8Y13_LUT4AB/N2END[5] Tile_X8Y13_LUT4AB/N2END[6]
+ Tile_X8Y13_LUT4AB/N2END[7] Tile_X8Y14_LUT4AB/N2END[0] Tile_X8Y14_LUT4AB/N2END[1]
+ Tile_X8Y14_LUT4AB/N2END[2] Tile_X8Y14_LUT4AB/N2END[3] Tile_X8Y14_LUT4AB/N2END[4]
+ Tile_X8Y14_LUT4AB/N2END[5] Tile_X8Y14_LUT4AB/N2END[6] Tile_X8Y14_LUT4AB/N2END[7]
+ Tile_X8Y14_LUT4AB/N2MID[0] Tile_X8Y14_LUT4AB/N2MID[1] Tile_X8Y14_LUT4AB/N2MID[2]
+ Tile_X8Y14_LUT4AB/N2MID[3] Tile_X8Y14_LUT4AB/N2MID[4] Tile_X8Y14_LUT4AB/N2MID[5]
+ Tile_X8Y14_LUT4AB/N2MID[6] Tile_X8Y14_LUT4AB/N2MID[7] Tile_X8Y14_LUT4AB/N4BEG[0]
+ Tile_X8Y14_LUT4AB/N4BEG[10] Tile_X8Y14_LUT4AB/N4BEG[11] Tile_X8Y14_LUT4AB/N4BEG[12]
+ Tile_X8Y14_LUT4AB/N4BEG[13] Tile_X8Y14_LUT4AB/N4BEG[14] Tile_X8Y14_LUT4AB/N4BEG[15]
+ Tile_X8Y14_LUT4AB/N4BEG[1] Tile_X8Y14_LUT4AB/N4BEG[2] Tile_X8Y14_LUT4AB/N4BEG[3]
+ Tile_X8Y14_LUT4AB/N4BEG[4] Tile_X8Y14_LUT4AB/N4BEG[5] Tile_X8Y14_LUT4AB/N4BEG[6]
+ Tile_X8Y14_LUT4AB/N4BEG[7] Tile_X8Y14_LUT4AB/N4BEG[8] Tile_X8Y14_LUT4AB/N4BEG[9]
+ Tile_X8Y14_LUT4AB/N4END[0] Tile_X8Y14_LUT4AB/N4END[10] Tile_X8Y14_LUT4AB/N4END[11]
+ Tile_X8Y14_LUT4AB/N4END[12] Tile_X8Y14_LUT4AB/N4END[13] Tile_X8Y14_LUT4AB/N4END[14]
+ Tile_X8Y14_LUT4AB/N4END[15] Tile_X8Y14_LUT4AB/N4END[1] Tile_X8Y14_LUT4AB/N4END[2]
+ Tile_X8Y14_LUT4AB/N4END[3] Tile_X8Y14_LUT4AB/N4END[4] Tile_X8Y14_LUT4AB/N4END[5]
+ Tile_X8Y14_LUT4AB/N4END[6] Tile_X8Y14_LUT4AB/N4END[7] Tile_X8Y14_LUT4AB/N4END[8]
+ Tile_X8Y14_LUT4AB/N4END[9] Tile_X8Y14_LUT4AB/NN4BEG[0] Tile_X8Y14_LUT4AB/NN4BEG[10]
+ Tile_X8Y14_LUT4AB/NN4BEG[11] Tile_X8Y14_LUT4AB/NN4BEG[12] Tile_X8Y14_LUT4AB/NN4BEG[13]
+ Tile_X8Y14_LUT4AB/NN4BEG[14] Tile_X8Y14_LUT4AB/NN4BEG[15] Tile_X8Y14_LUT4AB/NN4BEG[1]
+ Tile_X8Y14_LUT4AB/NN4BEG[2] Tile_X8Y14_LUT4AB/NN4BEG[3] Tile_X8Y14_LUT4AB/NN4BEG[4]
+ Tile_X8Y14_LUT4AB/NN4BEG[5] Tile_X8Y14_LUT4AB/NN4BEG[6] Tile_X8Y14_LUT4AB/NN4BEG[7]
+ Tile_X8Y14_LUT4AB/NN4BEG[8] Tile_X8Y14_LUT4AB/NN4BEG[9] Tile_X8Y14_LUT4AB/NN4END[0]
+ Tile_X8Y14_LUT4AB/NN4END[10] Tile_X8Y14_LUT4AB/NN4END[11] Tile_X8Y14_LUT4AB/NN4END[12]
+ Tile_X8Y14_LUT4AB/NN4END[13] Tile_X8Y14_LUT4AB/NN4END[14] Tile_X8Y14_LUT4AB/NN4END[15]
+ Tile_X8Y14_LUT4AB/NN4END[1] Tile_X8Y14_LUT4AB/NN4END[2] Tile_X8Y14_LUT4AB/NN4END[3]
+ Tile_X8Y14_LUT4AB/NN4END[4] Tile_X8Y14_LUT4AB/NN4END[5] Tile_X8Y14_LUT4AB/NN4END[6]
+ Tile_X8Y14_LUT4AB/NN4END[7] Tile_X8Y14_LUT4AB/NN4END[8] Tile_X8Y14_LUT4AB/NN4END[9]
+ Tile_X8Y14_LUT4AB/S1BEG[0] Tile_X8Y14_LUT4AB/S1BEG[1] Tile_X8Y14_LUT4AB/S1BEG[2]
+ Tile_X8Y14_LUT4AB/S1BEG[3] Tile_X8Y14_LUT4AB/S1END[0] Tile_X8Y14_LUT4AB/S1END[1]
+ Tile_X8Y14_LUT4AB/S1END[2] Tile_X8Y14_LUT4AB/S1END[3] Tile_X8Y14_LUT4AB/S2BEG[0]
+ Tile_X8Y14_LUT4AB/S2BEG[1] Tile_X8Y14_LUT4AB/S2BEG[2] Tile_X8Y14_LUT4AB/S2BEG[3]
+ Tile_X8Y14_LUT4AB/S2BEG[4] Tile_X8Y14_LUT4AB/S2BEG[5] Tile_X8Y14_LUT4AB/S2BEG[6]
+ Tile_X8Y14_LUT4AB/S2BEG[7] Tile_X8Y14_LUT4AB/S2BEGb[0] Tile_X8Y14_LUT4AB/S2BEGb[1]
+ Tile_X8Y14_LUT4AB/S2BEGb[2] Tile_X8Y14_LUT4AB/S2BEGb[3] Tile_X8Y14_LUT4AB/S2BEGb[4]
+ Tile_X8Y14_LUT4AB/S2BEGb[5] Tile_X8Y14_LUT4AB/S2BEGb[6] Tile_X8Y14_LUT4AB/S2BEGb[7]
+ Tile_X8Y14_LUT4AB/S2END[0] Tile_X8Y14_LUT4AB/S2END[1] Tile_X8Y14_LUT4AB/S2END[2]
+ Tile_X8Y14_LUT4AB/S2END[3] Tile_X8Y14_LUT4AB/S2END[4] Tile_X8Y14_LUT4AB/S2END[5]
+ Tile_X8Y14_LUT4AB/S2END[6] Tile_X8Y14_LUT4AB/S2END[7] Tile_X8Y14_LUT4AB/S2MID[0]
+ Tile_X8Y14_LUT4AB/S2MID[1] Tile_X8Y14_LUT4AB/S2MID[2] Tile_X8Y14_LUT4AB/S2MID[3]
+ Tile_X8Y14_LUT4AB/S2MID[4] Tile_X8Y14_LUT4AB/S2MID[5] Tile_X8Y14_LUT4AB/S2MID[6]
+ Tile_X8Y14_LUT4AB/S2MID[7] Tile_X8Y14_LUT4AB/S4BEG[0] Tile_X8Y14_LUT4AB/S4BEG[10]
+ Tile_X8Y14_LUT4AB/S4BEG[11] Tile_X8Y14_LUT4AB/S4BEG[12] Tile_X8Y14_LUT4AB/S4BEG[13]
+ Tile_X8Y14_LUT4AB/S4BEG[14] Tile_X8Y14_LUT4AB/S4BEG[15] Tile_X8Y14_LUT4AB/S4BEG[1]
+ Tile_X8Y14_LUT4AB/S4BEG[2] Tile_X8Y14_LUT4AB/S4BEG[3] Tile_X8Y14_LUT4AB/S4BEG[4]
+ Tile_X8Y14_LUT4AB/S4BEG[5] Tile_X8Y14_LUT4AB/S4BEG[6] Tile_X8Y14_LUT4AB/S4BEG[7]
+ Tile_X8Y14_LUT4AB/S4BEG[8] Tile_X8Y14_LUT4AB/S4BEG[9] Tile_X8Y14_LUT4AB/S4END[0]
+ Tile_X8Y14_LUT4AB/S4END[10] Tile_X8Y14_LUT4AB/S4END[11] Tile_X8Y14_LUT4AB/S4END[12]
+ Tile_X8Y14_LUT4AB/S4END[13] Tile_X8Y14_LUT4AB/S4END[14] Tile_X8Y14_LUT4AB/S4END[15]
+ Tile_X8Y14_LUT4AB/S4END[1] Tile_X8Y14_LUT4AB/S4END[2] Tile_X8Y14_LUT4AB/S4END[3]
+ Tile_X8Y14_LUT4AB/S4END[4] Tile_X8Y14_LUT4AB/S4END[5] Tile_X8Y14_LUT4AB/S4END[6]
+ Tile_X8Y14_LUT4AB/S4END[7] Tile_X8Y14_LUT4AB/S4END[8] Tile_X8Y14_LUT4AB/S4END[9]
+ Tile_X8Y14_LUT4AB/SS4BEG[0] Tile_X8Y14_LUT4AB/SS4BEG[10] Tile_X8Y14_LUT4AB/SS4BEG[11]
+ Tile_X8Y14_LUT4AB/SS4BEG[12] Tile_X8Y14_LUT4AB/SS4BEG[13] Tile_X8Y14_LUT4AB/SS4BEG[14]
+ Tile_X8Y14_LUT4AB/SS4BEG[15] Tile_X8Y14_LUT4AB/SS4BEG[1] Tile_X8Y14_LUT4AB/SS4BEG[2]
+ Tile_X8Y14_LUT4AB/SS4BEG[3] Tile_X8Y14_LUT4AB/SS4BEG[4] Tile_X8Y14_LUT4AB/SS4BEG[5]
+ Tile_X8Y14_LUT4AB/SS4BEG[6] Tile_X8Y14_LUT4AB/SS4BEG[7] Tile_X8Y14_LUT4AB/SS4BEG[8]
+ Tile_X8Y14_LUT4AB/SS4BEG[9] Tile_X8Y14_LUT4AB/SS4END[0] Tile_X8Y14_LUT4AB/SS4END[10]
+ Tile_X8Y14_LUT4AB/SS4END[11] Tile_X8Y14_LUT4AB/SS4END[12] Tile_X8Y14_LUT4AB/SS4END[13]
+ Tile_X8Y14_LUT4AB/SS4END[14] Tile_X8Y14_LUT4AB/SS4END[15] Tile_X8Y14_LUT4AB/SS4END[1]
+ Tile_X8Y14_LUT4AB/SS4END[2] Tile_X8Y14_LUT4AB/SS4END[3] Tile_X8Y14_LUT4AB/SS4END[4]
+ Tile_X8Y14_LUT4AB/SS4END[5] Tile_X8Y14_LUT4AB/SS4END[6] Tile_X8Y14_LUT4AB/SS4END[7]
+ Tile_X8Y14_LUT4AB/SS4END[8] Tile_X8Y14_LUT4AB/SS4END[9] Tile_X8Y14_LUT4AB/UserCLK
+ Tile_X8Y13_LUT4AB/UserCLK VGND VPWR Tile_X8Y14_LUT4AB/W1BEG[0] Tile_X8Y14_LUT4AB/W1BEG[1]
+ Tile_X8Y14_LUT4AB/W1BEG[2] Tile_X8Y14_LUT4AB/W1BEG[3] Tile_X9Y14_LUT4AB/W1BEG[0]
+ Tile_X9Y14_LUT4AB/W1BEG[1] Tile_X9Y14_LUT4AB/W1BEG[2] Tile_X9Y14_LUT4AB/W1BEG[3]
+ Tile_X8Y14_LUT4AB/W2BEG[0] Tile_X8Y14_LUT4AB/W2BEG[1] Tile_X8Y14_LUT4AB/W2BEG[2]
+ Tile_X8Y14_LUT4AB/W2BEG[3] Tile_X8Y14_LUT4AB/W2BEG[4] Tile_X8Y14_LUT4AB/W2BEG[5]
+ Tile_X8Y14_LUT4AB/W2BEG[6] Tile_X8Y14_LUT4AB/W2BEG[7] Tile_X8Y14_LUT4AB/W2BEGb[0]
+ Tile_X8Y14_LUT4AB/W2BEGb[1] Tile_X8Y14_LUT4AB/W2BEGb[2] Tile_X8Y14_LUT4AB/W2BEGb[3]
+ Tile_X8Y14_LUT4AB/W2BEGb[4] Tile_X8Y14_LUT4AB/W2BEGb[5] Tile_X8Y14_LUT4AB/W2BEGb[6]
+ Tile_X8Y14_LUT4AB/W2BEGb[7] Tile_X8Y14_LUT4AB/W2END[0] Tile_X8Y14_LUT4AB/W2END[1]
+ Tile_X8Y14_LUT4AB/W2END[2] Tile_X8Y14_LUT4AB/W2END[3] Tile_X8Y14_LUT4AB/W2END[4]
+ Tile_X8Y14_LUT4AB/W2END[5] Tile_X8Y14_LUT4AB/W2END[6] Tile_X8Y14_LUT4AB/W2END[7]
+ Tile_X9Y14_LUT4AB/W2BEG[0] Tile_X9Y14_LUT4AB/W2BEG[1] Tile_X9Y14_LUT4AB/W2BEG[2]
+ Tile_X9Y14_LUT4AB/W2BEG[3] Tile_X9Y14_LUT4AB/W2BEG[4] Tile_X9Y14_LUT4AB/W2BEG[5]
+ Tile_X9Y14_LUT4AB/W2BEG[6] Tile_X9Y14_LUT4AB/W2BEG[7] Tile_X8Y14_LUT4AB/W6BEG[0]
+ Tile_X8Y14_LUT4AB/W6BEG[10] Tile_X8Y14_LUT4AB/W6BEG[11] Tile_X8Y14_LUT4AB/W6BEG[1]
+ Tile_X8Y14_LUT4AB/W6BEG[2] Tile_X8Y14_LUT4AB/W6BEG[3] Tile_X8Y14_LUT4AB/W6BEG[4]
+ Tile_X8Y14_LUT4AB/W6BEG[5] Tile_X8Y14_LUT4AB/W6BEG[6] Tile_X8Y14_LUT4AB/W6BEG[7]
+ Tile_X8Y14_LUT4AB/W6BEG[8] Tile_X8Y14_LUT4AB/W6BEG[9] Tile_X9Y14_LUT4AB/W6BEG[0]
+ Tile_X9Y14_LUT4AB/W6BEG[10] Tile_X9Y14_LUT4AB/W6BEG[11] Tile_X9Y14_LUT4AB/W6BEG[1]
+ Tile_X9Y14_LUT4AB/W6BEG[2] Tile_X9Y14_LUT4AB/W6BEG[3] Tile_X9Y14_LUT4AB/W6BEG[4]
+ Tile_X9Y14_LUT4AB/W6BEG[5] Tile_X9Y14_LUT4AB/W6BEG[6] Tile_X9Y14_LUT4AB/W6BEG[7]
+ Tile_X9Y14_LUT4AB/W6BEG[8] Tile_X9Y14_LUT4AB/W6BEG[9] Tile_X8Y14_LUT4AB/WW4BEG[0]
+ Tile_X8Y14_LUT4AB/WW4BEG[10] Tile_X8Y14_LUT4AB/WW4BEG[11] Tile_X8Y14_LUT4AB/WW4BEG[12]
+ Tile_X8Y14_LUT4AB/WW4BEG[13] Tile_X8Y14_LUT4AB/WW4BEG[14] Tile_X8Y14_LUT4AB/WW4BEG[15]
+ Tile_X8Y14_LUT4AB/WW4BEG[1] Tile_X8Y14_LUT4AB/WW4BEG[2] Tile_X8Y14_LUT4AB/WW4BEG[3]
+ Tile_X8Y14_LUT4AB/WW4BEG[4] Tile_X8Y14_LUT4AB/WW4BEG[5] Tile_X8Y14_LUT4AB/WW4BEG[6]
+ Tile_X8Y14_LUT4AB/WW4BEG[7] Tile_X8Y14_LUT4AB/WW4BEG[8] Tile_X8Y14_LUT4AB/WW4BEG[9]
+ Tile_X9Y14_LUT4AB/WW4BEG[0] Tile_X9Y14_LUT4AB/WW4BEG[10] Tile_X9Y14_LUT4AB/WW4BEG[11]
+ Tile_X9Y14_LUT4AB/WW4BEG[12] Tile_X9Y14_LUT4AB/WW4BEG[13] Tile_X9Y14_LUT4AB/WW4BEG[14]
+ Tile_X9Y14_LUT4AB/WW4BEG[15] Tile_X9Y14_LUT4AB/WW4BEG[1] Tile_X9Y14_LUT4AB/WW4BEG[2]
+ Tile_X9Y14_LUT4AB/WW4BEG[3] Tile_X9Y14_LUT4AB/WW4BEG[4] Tile_X9Y14_LUT4AB/WW4BEG[5]
+ Tile_X9Y14_LUT4AB/WW4BEG[6] Tile_X9Y14_LUT4AB/WW4BEG[7] Tile_X9Y14_LUT4AB/WW4BEG[8]
+ Tile_X9Y14_LUT4AB/WW4BEG[9] LUT4AB
XTile_X5Y9_LUT4AB Tile_X5Y9_LUT4AB/Ci Tile_X5Y9_LUT4AB/Co Tile_X6Y9_LUT4AB/E1END[0]
+ Tile_X6Y9_LUT4AB/E1END[1] Tile_X6Y9_LUT4AB/E1END[2] Tile_X6Y9_LUT4AB/E1END[3] Tile_X5Y9_LUT4AB/E1END[0]
+ Tile_X5Y9_LUT4AB/E1END[1] Tile_X5Y9_LUT4AB/E1END[2] Tile_X5Y9_LUT4AB/E1END[3] Tile_X6Y9_LUT4AB/E2MID[0]
+ Tile_X6Y9_LUT4AB/E2MID[1] Tile_X6Y9_LUT4AB/E2MID[2] Tile_X6Y9_LUT4AB/E2MID[3] Tile_X6Y9_LUT4AB/E2MID[4]
+ Tile_X6Y9_LUT4AB/E2MID[5] Tile_X6Y9_LUT4AB/E2MID[6] Tile_X6Y9_LUT4AB/E2MID[7] Tile_X6Y9_LUT4AB/E2END[0]
+ Tile_X6Y9_LUT4AB/E2END[1] Tile_X6Y9_LUT4AB/E2END[2] Tile_X6Y9_LUT4AB/E2END[3] Tile_X6Y9_LUT4AB/E2END[4]
+ Tile_X6Y9_LUT4AB/E2END[5] Tile_X6Y9_LUT4AB/E2END[6] Tile_X6Y9_LUT4AB/E2END[7] Tile_X5Y9_LUT4AB/E2END[0]
+ Tile_X5Y9_LUT4AB/E2END[1] Tile_X5Y9_LUT4AB/E2END[2] Tile_X5Y9_LUT4AB/E2END[3] Tile_X5Y9_LUT4AB/E2END[4]
+ Tile_X5Y9_LUT4AB/E2END[5] Tile_X5Y9_LUT4AB/E2END[6] Tile_X5Y9_LUT4AB/E2END[7] Tile_X5Y9_LUT4AB/E2MID[0]
+ Tile_X5Y9_LUT4AB/E2MID[1] Tile_X5Y9_LUT4AB/E2MID[2] Tile_X5Y9_LUT4AB/E2MID[3] Tile_X5Y9_LUT4AB/E2MID[4]
+ Tile_X5Y9_LUT4AB/E2MID[5] Tile_X5Y9_LUT4AB/E2MID[6] Tile_X5Y9_LUT4AB/E2MID[7] Tile_X6Y9_LUT4AB/E6END[0]
+ Tile_X6Y9_LUT4AB/E6END[10] Tile_X6Y9_LUT4AB/E6END[11] Tile_X6Y9_LUT4AB/E6END[1]
+ Tile_X6Y9_LUT4AB/E6END[2] Tile_X6Y9_LUT4AB/E6END[3] Tile_X6Y9_LUT4AB/E6END[4] Tile_X6Y9_LUT4AB/E6END[5]
+ Tile_X6Y9_LUT4AB/E6END[6] Tile_X6Y9_LUT4AB/E6END[7] Tile_X6Y9_LUT4AB/E6END[8] Tile_X6Y9_LUT4AB/E6END[9]
+ Tile_X5Y9_LUT4AB/E6END[0] Tile_X5Y9_LUT4AB/E6END[10] Tile_X5Y9_LUT4AB/E6END[11]
+ Tile_X5Y9_LUT4AB/E6END[1] Tile_X5Y9_LUT4AB/E6END[2] Tile_X5Y9_LUT4AB/E6END[3] Tile_X5Y9_LUT4AB/E6END[4]
+ Tile_X5Y9_LUT4AB/E6END[5] Tile_X5Y9_LUT4AB/E6END[6] Tile_X5Y9_LUT4AB/E6END[7] Tile_X5Y9_LUT4AB/E6END[8]
+ Tile_X5Y9_LUT4AB/E6END[9] Tile_X6Y9_LUT4AB/EE4END[0] Tile_X6Y9_LUT4AB/EE4END[10]
+ Tile_X6Y9_LUT4AB/EE4END[11] Tile_X6Y9_LUT4AB/EE4END[12] Tile_X6Y9_LUT4AB/EE4END[13]
+ Tile_X6Y9_LUT4AB/EE4END[14] Tile_X6Y9_LUT4AB/EE4END[15] Tile_X6Y9_LUT4AB/EE4END[1]
+ Tile_X6Y9_LUT4AB/EE4END[2] Tile_X6Y9_LUT4AB/EE4END[3] Tile_X6Y9_LUT4AB/EE4END[4]
+ Tile_X6Y9_LUT4AB/EE4END[5] Tile_X6Y9_LUT4AB/EE4END[6] Tile_X6Y9_LUT4AB/EE4END[7]
+ Tile_X6Y9_LUT4AB/EE4END[8] Tile_X6Y9_LUT4AB/EE4END[9] Tile_X5Y9_LUT4AB/EE4END[0]
+ Tile_X5Y9_LUT4AB/EE4END[10] Tile_X5Y9_LUT4AB/EE4END[11] Tile_X5Y9_LUT4AB/EE4END[12]
+ Tile_X5Y9_LUT4AB/EE4END[13] Tile_X5Y9_LUT4AB/EE4END[14] Tile_X5Y9_LUT4AB/EE4END[15]
+ Tile_X5Y9_LUT4AB/EE4END[1] Tile_X5Y9_LUT4AB/EE4END[2] Tile_X5Y9_LUT4AB/EE4END[3]
+ Tile_X5Y9_LUT4AB/EE4END[4] Tile_X5Y9_LUT4AB/EE4END[5] Tile_X5Y9_LUT4AB/EE4END[6]
+ Tile_X5Y9_LUT4AB/EE4END[7] Tile_X5Y9_LUT4AB/EE4END[8] Tile_X5Y9_LUT4AB/EE4END[9]
+ Tile_X5Y9_LUT4AB/FrameData[0] Tile_X5Y9_LUT4AB/FrameData[10] Tile_X5Y9_LUT4AB/FrameData[11]
+ Tile_X5Y9_LUT4AB/FrameData[12] Tile_X5Y9_LUT4AB/FrameData[13] Tile_X5Y9_LUT4AB/FrameData[14]
+ Tile_X5Y9_LUT4AB/FrameData[15] Tile_X5Y9_LUT4AB/FrameData[16] Tile_X5Y9_LUT4AB/FrameData[17]
+ Tile_X5Y9_LUT4AB/FrameData[18] Tile_X5Y9_LUT4AB/FrameData[19] Tile_X5Y9_LUT4AB/FrameData[1]
+ Tile_X5Y9_LUT4AB/FrameData[20] Tile_X5Y9_LUT4AB/FrameData[21] Tile_X5Y9_LUT4AB/FrameData[22]
+ Tile_X5Y9_LUT4AB/FrameData[23] Tile_X5Y9_LUT4AB/FrameData[24] Tile_X5Y9_LUT4AB/FrameData[25]
+ Tile_X5Y9_LUT4AB/FrameData[26] Tile_X5Y9_LUT4AB/FrameData[27] Tile_X5Y9_LUT4AB/FrameData[28]
+ Tile_X5Y9_LUT4AB/FrameData[29] Tile_X5Y9_LUT4AB/FrameData[2] Tile_X5Y9_LUT4AB/FrameData[30]
+ Tile_X5Y9_LUT4AB/FrameData[31] Tile_X5Y9_LUT4AB/FrameData[3] Tile_X5Y9_LUT4AB/FrameData[4]
+ Tile_X5Y9_LUT4AB/FrameData[5] Tile_X5Y9_LUT4AB/FrameData[6] Tile_X5Y9_LUT4AB/FrameData[7]
+ Tile_X5Y9_LUT4AB/FrameData[8] Tile_X5Y9_LUT4AB/FrameData[9] Tile_X6Y9_LUT4AB/FrameData[0]
+ Tile_X6Y9_LUT4AB/FrameData[10] Tile_X6Y9_LUT4AB/FrameData[11] Tile_X6Y9_LUT4AB/FrameData[12]
+ Tile_X6Y9_LUT4AB/FrameData[13] Tile_X6Y9_LUT4AB/FrameData[14] Tile_X6Y9_LUT4AB/FrameData[15]
+ Tile_X6Y9_LUT4AB/FrameData[16] Tile_X6Y9_LUT4AB/FrameData[17] Tile_X6Y9_LUT4AB/FrameData[18]
+ Tile_X6Y9_LUT4AB/FrameData[19] Tile_X6Y9_LUT4AB/FrameData[1] Tile_X6Y9_LUT4AB/FrameData[20]
+ Tile_X6Y9_LUT4AB/FrameData[21] Tile_X6Y9_LUT4AB/FrameData[22] Tile_X6Y9_LUT4AB/FrameData[23]
+ Tile_X6Y9_LUT4AB/FrameData[24] Tile_X6Y9_LUT4AB/FrameData[25] Tile_X6Y9_LUT4AB/FrameData[26]
+ Tile_X6Y9_LUT4AB/FrameData[27] Tile_X6Y9_LUT4AB/FrameData[28] Tile_X6Y9_LUT4AB/FrameData[29]
+ Tile_X6Y9_LUT4AB/FrameData[2] Tile_X6Y9_LUT4AB/FrameData[30] Tile_X6Y9_LUT4AB/FrameData[31]
+ Tile_X6Y9_LUT4AB/FrameData[3] Tile_X6Y9_LUT4AB/FrameData[4] Tile_X6Y9_LUT4AB/FrameData[5]
+ Tile_X6Y9_LUT4AB/FrameData[6] Tile_X6Y9_LUT4AB/FrameData[7] Tile_X6Y9_LUT4AB/FrameData[8]
+ Tile_X6Y9_LUT4AB/FrameData[9] Tile_X5Y9_LUT4AB/FrameStrobe[0] Tile_X5Y9_LUT4AB/FrameStrobe[10]
+ Tile_X5Y9_LUT4AB/FrameStrobe[11] Tile_X5Y9_LUT4AB/FrameStrobe[12] Tile_X5Y9_LUT4AB/FrameStrobe[13]
+ Tile_X5Y9_LUT4AB/FrameStrobe[14] Tile_X5Y9_LUT4AB/FrameStrobe[15] Tile_X5Y9_LUT4AB/FrameStrobe[16]
+ Tile_X5Y9_LUT4AB/FrameStrobe[17] Tile_X5Y9_LUT4AB/FrameStrobe[18] Tile_X5Y9_LUT4AB/FrameStrobe[19]
+ Tile_X5Y9_LUT4AB/FrameStrobe[1] Tile_X5Y9_LUT4AB/FrameStrobe[2] Tile_X5Y9_LUT4AB/FrameStrobe[3]
+ Tile_X5Y9_LUT4AB/FrameStrobe[4] Tile_X5Y9_LUT4AB/FrameStrobe[5] Tile_X5Y9_LUT4AB/FrameStrobe[6]
+ Tile_X5Y9_LUT4AB/FrameStrobe[7] Tile_X5Y9_LUT4AB/FrameStrobe[8] Tile_X5Y9_LUT4AB/FrameStrobe[9]
+ Tile_X5Y8_LUT4AB/FrameStrobe[0] Tile_X5Y8_LUT4AB/FrameStrobe[10] Tile_X5Y8_LUT4AB/FrameStrobe[11]
+ Tile_X5Y8_LUT4AB/FrameStrobe[12] Tile_X5Y8_LUT4AB/FrameStrobe[13] Tile_X5Y8_LUT4AB/FrameStrobe[14]
+ Tile_X5Y8_LUT4AB/FrameStrobe[15] Tile_X5Y8_LUT4AB/FrameStrobe[16] Tile_X5Y8_LUT4AB/FrameStrobe[17]
+ Tile_X5Y8_LUT4AB/FrameStrobe[18] Tile_X5Y8_LUT4AB/FrameStrobe[19] Tile_X5Y8_LUT4AB/FrameStrobe[1]
+ Tile_X5Y8_LUT4AB/FrameStrobe[2] Tile_X5Y8_LUT4AB/FrameStrobe[3] Tile_X5Y8_LUT4AB/FrameStrobe[4]
+ Tile_X5Y8_LUT4AB/FrameStrobe[5] Tile_X5Y8_LUT4AB/FrameStrobe[6] Tile_X5Y8_LUT4AB/FrameStrobe[7]
+ Tile_X5Y8_LUT4AB/FrameStrobe[8] Tile_X5Y8_LUT4AB/FrameStrobe[9] Tile_X5Y9_LUT4AB/N1BEG[0]
+ Tile_X5Y9_LUT4AB/N1BEG[1] Tile_X5Y9_LUT4AB/N1BEG[2] Tile_X5Y9_LUT4AB/N1BEG[3] Tile_X5Y9_LUT4AB/N1END[0]
+ Tile_X5Y9_LUT4AB/N1END[1] Tile_X5Y9_LUT4AB/N1END[2] Tile_X5Y9_LUT4AB/N1END[3] Tile_X5Y9_LUT4AB/N2BEG[0]
+ Tile_X5Y9_LUT4AB/N2BEG[1] Tile_X5Y9_LUT4AB/N2BEG[2] Tile_X5Y9_LUT4AB/N2BEG[3] Tile_X5Y9_LUT4AB/N2BEG[4]
+ Tile_X5Y9_LUT4AB/N2BEG[5] Tile_X5Y9_LUT4AB/N2BEG[6] Tile_X5Y9_LUT4AB/N2BEG[7] Tile_X5Y8_LUT4AB/N2END[0]
+ Tile_X5Y8_LUT4AB/N2END[1] Tile_X5Y8_LUT4AB/N2END[2] Tile_X5Y8_LUT4AB/N2END[3] Tile_X5Y8_LUT4AB/N2END[4]
+ Tile_X5Y8_LUT4AB/N2END[5] Tile_X5Y8_LUT4AB/N2END[6] Tile_X5Y8_LUT4AB/N2END[7] Tile_X5Y9_LUT4AB/N2END[0]
+ Tile_X5Y9_LUT4AB/N2END[1] Tile_X5Y9_LUT4AB/N2END[2] Tile_X5Y9_LUT4AB/N2END[3] Tile_X5Y9_LUT4AB/N2END[4]
+ Tile_X5Y9_LUT4AB/N2END[5] Tile_X5Y9_LUT4AB/N2END[6] Tile_X5Y9_LUT4AB/N2END[7] Tile_X5Y9_LUT4AB/N2MID[0]
+ Tile_X5Y9_LUT4AB/N2MID[1] Tile_X5Y9_LUT4AB/N2MID[2] Tile_X5Y9_LUT4AB/N2MID[3] Tile_X5Y9_LUT4AB/N2MID[4]
+ Tile_X5Y9_LUT4AB/N2MID[5] Tile_X5Y9_LUT4AB/N2MID[6] Tile_X5Y9_LUT4AB/N2MID[7] Tile_X5Y9_LUT4AB/N4BEG[0]
+ Tile_X5Y9_LUT4AB/N4BEG[10] Tile_X5Y9_LUT4AB/N4BEG[11] Tile_X5Y9_LUT4AB/N4BEG[12]
+ Tile_X5Y9_LUT4AB/N4BEG[13] Tile_X5Y9_LUT4AB/N4BEG[14] Tile_X5Y9_LUT4AB/N4BEG[15]
+ Tile_X5Y9_LUT4AB/N4BEG[1] Tile_X5Y9_LUT4AB/N4BEG[2] Tile_X5Y9_LUT4AB/N4BEG[3] Tile_X5Y9_LUT4AB/N4BEG[4]
+ Tile_X5Y9_LUT4AB/N4BEG[5] Tile_X5Y9_LUT4AB/N4BEG[6] Tile_X5Y9_LUT4AB/N4BEG[7] Tile_X5Y9_LUT4AB/N4BEG[8]
+ Tile_X5Y9_LUT4AB/N4BEG[9] Tile_X5Y9_LUT4AB/N4END[0] Tile_X5Y9_LUT4AB/N4END[10] Tile_X5Y9_LUT4AB/N4END[11]
+ Tile_X5Y9_LUT4AB/N4END[12] Tile_X5Y9_LUT4AB/N4END[13] Tile_X5Y9_LUT4AB/N4END[14]
+ Tile_X5Y9_LUT4AB/N4END[15] Tile_X5Y9_LUT4AB/N4END[1] Tile_X5Y9_LUT4AB/N4END[2] Tile_X5Y9_LUT4AB/N4END[3]
+ Tile_X5Y9_LUT4AB/N4END[4] Tile_X5Y9_LUT4AB/N4END[5] Tile_X5Y9_LUT4AB/N4END[6] Tile_X5Y9_LUT4AB/N4END[7]
+ Tile_X5Y9_LUT4AB/N4END[8] Tile_X5Y9_LUT4AB/N4END[9] Tile_X5Y9_LUT4AB/NN4BEG[0] Tile_X5Y9_LUT4AB/NN4BEG[10]
+ Tile_X5Y9_LUT4AB/NN4BEG[11] Tile_X5Y9_LUT4AB/NN4BEG[12] Tile_X5Y9_LUT4AB/NN4BEG[13]
+ Tile_X5Y9_LUT4AB/NN4BEG[14] Tile_X5Y9_LUT4AB/NN4BEG[15] Tile_X5Y9_LUT4AB/NN4BEG[1]
+ Tile_X5Y9_LUT4AB/NN4BEG[2] Tile_X5Y9_LUT4AB/NN4BEG[3] Tile_X5Y9_LUT4AB/NN4BEG[4]
+ Tile_X5Y9_LUT4AB/NN4BEG[5] Tile_X5Y9_LUT4AB/NN4BEG[6] Tile_X5Y9_LUT4AB/NN4BEG[7]
+ Tile_X5Y9_LUT4AB/NN4BEG[8] Tile_X5Y9_LUT4AB/NN4BEG[9] Tile_X5Y9_LUT4AB/NN4END[0]
+ Tile_X5Y9_LUT4AB/NN4END[10] Tile_X5Y9_LUT4AB/NN4END[11] Tile_X5Y9_LUT4AB/NN4END[12]
+ Tile_X5Y9_LUT4AB/NN4END[13] Tile_X5Y9_LUT4AB/NN4END[14] Tile_X5Y9_LUT4AB/NN4END[15]
+ Tile_X5Y9_LUT4AB/NN4END[1] Tile_X5Y9_LUT4AB/NN4END[2] Tile_X5Y9_LUT4AB/NN4END[3]
+ Tile_X5Y9_LUT4AB/NN4END[4] Tile_X5Y9_LUT4AB/NN4END[5] Tile_X5Y9_LUT4AB/NN4END[6]
+ Tile_X5Y9_LUT4AB/NN4END[7] Tile_X5Y9_LUT4AB/NN4END[8] Tile_X5Y9_LUT4AB/NN4END[9]
+ Tile_X5Y9_LUT4AB/S1BEG[0] Tile_X5Y9_LUT4AB/S1BEG[1] Tile_X5Y9_LUT4AB/S1BEG[2] Tile_X5Y9_LUT4AB/S1BEG[3]
+ Tile_X5Y9_LUT4AB/S1END[0] Tile_X5Y9_LUT4AB/S1END[1] Tile_X5Y9_LUT4AB/S1END[2] Tile_X5Y9_LUT4AB/S1END[3]
+ Tile_X5Y9_LUT4AB/S2BEG[0] Tile_X5Y9_LUT4AB/S2BEG[1] Tile_X5Y9_LUT4AB/S2BEG[2] Tile_X5Y9_LUT4AB/S2BEG[3]
+ Tile_X5Y9_LUT4AB/S2BEG[4] Tile_X5Y9_LUT4AB/S2BEG[5] Tile_X5Y9_LUT4AB/S2BEG[6] Tile_X5Y9_LUT4AB/S2BEG[7]
+ Tile_X5Y9_LUT4AB/S2BEGb[0] Tile_X5Y9_LUT4AB/S2BEGb[1] Tile_X5Y9_LUT4AB/S2BEGb[2]
+ Tile_X5Y9_LUT4AB/S2BEGb[3] Tile_X5Y9_LUT4AB/S2BEGb[4] Tile_X5Y9_LUT4AB/S2BEGb[5]
+ Tile_X5Y9_LUT4AB/S2BEGb[6] Tile_X5Y9_LUT4AB/S2BEGb[7] Tile_X5Y9_LUT4AB/S2END[0]
+ Tile_X5Y9_LUT4AB/S2END[1] Tile_X5Y9_LUT4AB/S2END[2] Tile_X5Y9_LUT4AB/S2END[3] Tile_X5Y9_LUT4AB/S2END[4]
+ Tile_X5Y9_LUT4AB/S2END[5] Tile_X5Y9_LUT4AB/S2END[6] Tile_X5Y9_LUT4AB/S2END[7] Tile_X5Y9_LUT4AB/S2MID[0]
+ Tile_X5Y9_LUT4AB/S2MID[1] Tile_X5Y9_LUT4AB/S2MID[2] Tile_X5Y9_LUT4AB/S2MID[3] Tile_X5Y9_LUT4AB/S2MID[4]
+ Tile_X5Y9_LUT4AB/S2MID[5] Tile_X5Y9_LUT4AB/S2MID[6] Tile_X5Y9_LUT4AB/S2MID[7] Tile_X5Y9_LUT4AB/S4BEG[0]
+ Tile_X5Y9_LUT4AB/S4BEG[10] Tile_X5Y9_LUT4AB/S4BEG[11] Tile_X5Y9_LUT4AB/S4BEG[12]
+ Tile_X5Y9_LUT4AB/S4BEG[13] Tile_X5Y9_LUT4AB/S4BEG[14] Tile_X5Y9_LUT4AB/S4BEG[15]
+ Tile_X5Y9_LUT4AB/S4BEG[1] Tile_X5Y9_LUT4AB/S4BEG[2] Tile_X5Y9_LUT4AB/S4BEG[3] Tile_X5Y9_LUT4AB/S4BEG[4]
+ Tile_X5Y9_LUT4AB/S4BEG[5] Tile_X5Y9_LUT4AB/S4BEG[6] Tile_X5Y9_LUT4AB/S4BEG[7] Tile_X5Y9_LUT4AB/S4BEG[8]
+ Tile_X5Y9_LUT4AB/S4BEG[9] Tile_X5Y9_LUT4AB/S4END[0] Tile_X5Y9_LUT4AB/S4END[10] Tile_X5Y9_LUT4AB/S4END[11]
+ Tile_X5Y9_LUT4AB/S4END[12] Tile_X5Y9_LUT4AB/S4END[13] Tile_X5Y9_LUT4AB/S4END[14]
+ Tile_X5Y9_LUT4AB/S4END[15] Tile_X5Y9_LUT4AB/S4END[1] Tile_X5Y9_LUT4AB/S4END[2] Tile_X5Y9_LUT4AB/S4END[3]
+ Tile_X5Y9_LUT4AB/S4END[4] Tile_X5Y9_LUT4AB/S4END[5] Tile_X5Y9_LUT4AB/S4END[6] Tile_X5Y9_LUT4AB/S4END[7]
+ Tile_X5Y9_LUT4AB/S4END[8] Tile_X5Y9_LUT4AB/S4END[9] Tile_X5Y9_LUT4AB/SS4BEG[0] Tile_X5Y9_LUT4AB/SS4BEG[10]
+ Tile_X5Y9_LUT4AB/SS4BEG[11] Tile_X5Y9_LUT4AB/SS4BEG[12] Tile_X5Y9_LUT4AB/SS4BEG[13]
+ Tile_X5Y9_LUT4AB/SS4BEG[14] Tile_X5Y9_LUT4AB/SS4BEG[15] Tile_X5Y9_LUT4AB/SS4BEG[1]
+ Tile_X5Y9_LUT4AB/SS4BEG[2] Tile_X5Y9_LUT4AB/SS4BEG[3] Tile_X5Y9_LUT4AB/SS4BEG[4]
+ Tile_X5Y9_LUT4AB/SS4BEG[5] Tile_X5Y9_LUT4AB/SS4BEG[6] Tile_X5Y9_LUT4AB/SS4BEG[7]
+ Tile_X5Y9_LUT4AB/SS4BEG[8] Tile_X5Y9_LUT4AB/SS4BEG[9] Tile_X5Y9_LUT4AB/SS4END[0]
+ Tile_X5Y9_LUT4AB/SS4END[10] Tile_X5Y9_LUT4AB/SS4END[11] Tile_X5Y9_LUT4AB/SS4END[12]
+ Tile_X5Y9_LUT4AB/SS4END[13] Tile_X5Y9_LUT4AB/SS4END[14] Tile_X5Y9_LUT4AB/SS4END[15]
+ Tile_X5Y9_LUT4AB/SS4END[1] Tile_X5Y9_LUT4AB/SS4END[2] Tile_X5Y9_LUT4AB/SS4END[3]
+ Tile_X5Y9_LUT4AB/SS4END[4] Tile_X5Y9_LUT4AB/SS4END[5] Tile_X5Y9_LUT4AB/SS4END[6]
+ Tile_X5Y9_LUT4AB/SS4END[7] Tile_X5Y9_LUT4AB/SS4END[8] Tile_X5Y9_LUT4AB/SS4END[9]
+ Tile_X5Y9_LUT4AB/UserCLK Tile_X5Y8_LUT4AB/UserCLK VGND VPWR Tile_X5Y9_LUT4AB/W1BEG[0]
+ Tile_X5Y9_LUT4AB/W1BEG[1] Tile_X5Y9_LUT4AB/W1BEG[2] Tile_X5Y9_LUT4AB/W1BEG[3] Tile_X6Y9_LUT4AB/W1BEG[0]
+ Tile_X6Y9_LUT4AB/W1BEG[1] Tile_X6Y9_LUT4AB/W1BEG[2] Tile_X6Y9_LUT4AB/W1BEG[3] Tile_X5Y9_LUT4AB/W2BEG[0]
+ Tile_X5Y9_LUT4AB/W2BEG[1] Tile_X5Y9_LUT4AB/W2BEG[2] Tile_X5Y9_LUT4AB/W2BEG[3] Tile_X5Y9_LUT4AB/W2BEG[4]
+ Tile_X5Y9_LUT4AB/W2BEG[5] Tile_X5Y9_LUT4AB/W2BEG[6] Tile_X5Y9_LUT4AB/W2BEG[7] Tile_X5Y9_LUT4AB/W2BEGb[0]
+ Tile_X5Y9_LUT4AB/W2BEGb[1] Tile_X5Y9_LUT4AB/W2BEGb[2] Tile_X5Y9_LUT4AB/W2BEGb[3]
+ Tile_X5Y9_LUT4AB/W2BEGb[4] Tile_X5Y9_LUT4AB/W2BEGb[5] Tile_X5Y9_LUT4AB/W2BEGb[6]
+ Tile_X5Y9_LUT4AB/W2BEGb[7] Tile_X5Y9_LUT4AB/W2END[0] Tile_X5Y9_LUT4AB/W2END[1] Tile_X5Y9_LUT4AB/W2END[2]
+ Tile_X5Y9_LUT4AB/W2END[3] Tile_X5Y9_LUT4AB/W2END[4] Tile_X5Y9_LUT4AB/W2END[5] Tile_X5Y9_LUT4AB/W2END[6]
+ Tile_X5Y9_LUT4AB/W2END[7] Tile_X6Y9_LUT4AB/W2BEG[0] Tile_X6Y9_LUT4AB/W2BEG[1] Tile_X6Y9_LUT4AB/W2BEG[2]
+ Tile_X6Y9_LUT4AB/W2BEG[3] Tile_X6Y9_LUT4AB/W2BEG[4] Tile_X6Y9_LUT4AB/W2BEG[5] Tile_X6Y9_LUT4AB/W2BEG[6]
+ Tile_X6Y9_LUT4AB/W2BEG[7] Tile_X5Y9_LUT4AB/W6BEG[0] Tile_X5Y9_LUT4AB/W6BEG[10] Tile_X5Y9_LUT4AB/W6BEG[11]
+ Tile_X5Y9_LUT4AB/W6BEG[1] Tile_X5Y9_LUT4AB/W6BEG[2] Tile_X5Y9_LUT4AB/W6BEG[3] Tile_X5Y9_LUT4AB/W6BEG[4]
+ Tile_X5Y9_LUT4AB/W6BEG[5] Tile_X5Y9_LUT4AB/W6BEG[6] Tile_X5Y9_LUT4AB/W6BEG[7] Tile_X5Y9_LUT4AB/W6BEG[8]
+ Tile_X5Y9_LUT4AB/W6BEG[9] Tile_X6Y9_LUT4AB/W6BEG[0] Tile_X6Y9_LUT4AB/W6BEG[10] Tile_X6Y9_LUT4AB/W6BEG[11]
+ Tile_X6Y9_LUT4AB/W6BEG[1] Tile_X6Y9_LUT4AB/W6BEG[2] Tile_X6Y9_LUT4AB/W6BEG[3] Tile_X6Y9_LUT4AB/W6BEG[4]
+ Tile_X6Y9_LUT4AB/W6BEG[5] Tile_X6Y9_LUT4AB/W6BEG[6] Tile_X6Y9_LUT4AB/W6BEG[7] Tile_X6Y9_LUT4AB/W6BEG[8]
+ Tile_X6Y9_LUT4AB/W6BEG[9] Tile_X5Y9_LUT4AB/WW4BEG[0] Tile_X5Y9_LUT4AB/WW4BEG[10]
+ Tile_X5Y9_LUT4AB/WW4BEG[11] Tile_X5Y9_LUT4AB/WW4BEG[12] Tile_X5Y9_LUT4AB/WW4BEG[13]
+ Tile_X5Y9_LUT4AB/WW4BEG[14] Tile_X5Y9_LUT4AB/WW4BEG[15] Tile_X5Y9_LUT4AB/WW4BEG[1]
+ Tile_X5Y9_LUT4AB/WW4BEG[2] Tile_X5Y9_LUT4AB/WW4BEG[3] Tile_X5Y9_LUT4AB/WW4BEG[4]
+ Tile_X5Y9_LUT4AB/WW4BEG[5] Tile_X5Y9_LUT4AB/WW4BEG[6] Tile_X5Y9_LUT4AB/WW4BEG[7]
+ Tile_X5Y9_LUT4AB/WW4BEG[8] Tile_X5Y9_LUT4AB/WW4BEG[9] Tile_X6Y9_LUT4AB/WW4BEG[0]
+ Tile_X6Y9_LUT4AB/WW4BEG[10] Tile_X6Y9_LUT4AB/WW4BEG[11] Tile_X6Y9_LUT4AB/WW4BEG[12]
+ Tile_X6Y9_LUT4AB/WW4BEG[13] Tile_X6Y9_LUT4AB/WW4BEG[14] Tile_X6Y9_LUT4AB/WW4BEG[15]
+ Tile_X6Y9_LUT4AB/WW4BEG[1] Tile_X6Y9_LUT4AB/WW4BEG[2] Tile_X6Y9_LUT4AB/WW4BEG[3]
+ Tile_X6Y9_LUT4AB/WW4BEG[4] Tile_X6Y9_LUT4AB/WW4BEG[5] Tile_X6Y9_LUT4AB/WW4BEG[6]
+ Tile_X6Y9_LUT4AB/WW4BEG[7] Tile_X6Y9_LUT4AB/WW4BEG[8] Tile_X6Y9_LUT4AB/WW4BEG[9]
+ LUT4AB
XTile_X2Y4_LUT4AB Tile_X2Y5_LUT4AB/Co Tile_X2Y4_LUT4AB/Co Tile_X3Y4_LUT4AB/E1END[0]
+ Tile_X3Y4_LUT4AB/E1END[1] Tile_X3Y4_LUT4AB/E1END[2] Tile_X3Y4_LUT4AB/E1END[3] Tile_X2Y4_LUT4AB/E1END[0]
+ Tile_X2Y4_LUT4AB/E1END[1] Tile_X2Y4_LUT4AB/E1END[2] Tile_X2Y4_LUT4AB/E1END[3] Tile_X3Y4_LUT4AB/E2MID[0]
+ Tile_X3Y4_LUT4AB/E2MID[1] Tile_X3Y4_LUT4AB/E2MID[2] Tile_X3Y4_LUT4AB/E2MID[3] Tile_X3Y4_LUT4AB/E2MID[4]
+ Tile_X3Y4_LUT4AB/E2MID[5] Tile_X3Y4_LUT4AB/E2MID[6] Tile_X3Y4_LUT4AB/E2MID[7] Tile_X3Y4_LUT4AB/E2END[0]
+ Tile_X3Y4_LUT4AB/E2END[1] Tile_X3Y4_LUT4AB/E2END[2] Tile_X3Y4_LUT4AB/E2END[3] Tile_X3Y4_LUT4AB/E2END[4]
+ Tile_X3Y4_LUT4AB/E2END[5] Tile_X3Y4_LUT4AB/E2END[6] Tile_X3Y4_LUT4AB/E2END[7] Tile_X2Y4_LUT4AB/E2END[0]
+ Tile_X2Y4_LUT4AB/E2END[1] Tile_X2Y4_LUT4AB/E2END[2] Tile_X2Y4_LUT4AB/E2END[3] Tile_X2Y4_LUT4AB/E2END[4]
+ Tile_X2Y4_LUT4AB/E2END[5] Tile_X2Y4_LUT4AB/E2END[6] Tile_X2Y4_LUT4AB/E2END[7] Tile_X2Y4_LUT4AB/E2MID[0]
+ Tile_X2Y4_LUT4AB/E2MID[1] Tile_X2Y4_LUT4AB/E2MID[2] Tile_X2Y4_LUT4AB/E2MID[3] Tile_X2Y4_LUT4AB/E2MID[4]
+ Tile_X2Y4_LUT4AB/E2MID[5] Tile_X2Y4_LUT4AB/E2MID[6] Tile_X2Y4_LUT4AB/E2MID[7] Tile_X3Y4_LUT4AB/E6END[0]
+ Tile_X3Y4_LUT4AB/E6END[10] Tile_X3Y4_LUT4AB/E6END[11] Tile_X3Y4_LUT4AB/E6END[1]
+ Tile_X3Y4_LUT4AB/E6END[2] Tile_X3Y4_LUT4AB/E6END[3] Tile_X3Y4_LUT4AB/E6END[4] Tile_X3Y4_LUT4AB/E6END[5]
+ Tile_X3Y4_LUT4AB/E6END[6] Tile_X3Y4_LUT4AB/E6END[7] Tile_X3Y4_LUT4AB/E6END[8] Tile_X3Y4_LUT4AB/E6END[9]
+ Tile_X2Y4_LUT4AB/E6END[0] Tile_X2Y4_LUT4AB/E6END[10] Tile_X2Y4_LUT4AB/E6END[11]
+ Tile_X2Y4_LUT4AB/E6END[1] Tile_X2Y4_LUT4AB/E6END[2] Tile_X2Y4_LUT4AB/E6END[3] Tile_X2Y4_LUT4AB/E6END[4]
+ Tile_X2Y4_LUT4AB/E6END[5] Tile_X2Y4_LUT4AB/E6END[6] Tile_X2Y4_LUT4AB/E6END[7] Tile_X2Y4_LUT4AB/E6END[8]
+ Tile_X2Y4_LUT4AB/E6END[9] Tile_X3Y4_LUT4AB/EE4END[0] Tile_X3Y4_LUT4AB/EE4END[10]
+ Tile_X3Y4_LUT4AB/EE4END[11] Tile_X3Y4_LUT4AB/EE4END[12] Tile_X3Y4_LUT4AB/EE4END[13]
+ Tile_X3Y4_LUT4AB/EE4END[14] Tile_X3Y4_LUT4AB/EE4END[15] Tile_X3Y4_LUT4AB/EE4END[1]
+ Tile_X3Y4_LUT4AB/EE4END[2] Tile_X3Y4_LUT4AB/EE4END[3] Tile_X3Y4_LUT4AB/EE4END[4]
+ Tile_X3Y4_LUT4AB/EE4END[5] Tile_X3Y4_LUT4AB/EE4END[6] Tile_X3Y4_LUT4AB/EE4END[7]
+ Tile_X3Y4_LUT4AB/EE4END[8] Tile_X3Y4_LUT4AB/EE4END[9] Tile_X2Y4_LUT4AB/EE4END[0]
+ Tile_X2Y4_LUT4AB/EE4END[10] Tile_X2Y4_LUT4AB/EE4END[11] Tile_X2Y4_LUT4AB/EE4END[12]
+ Tile_X2Y4_LUT4AB/EE4END[13] Tile_X2Y4_LUT4AB/EE4END[14] Tile_X2Y4_LUT4AB/EE4END[15]
+ Tile_X2Y4_LUT4AB/EE4END[1] Tile_X2Y4_LUT4AB/EE4END[2] Tile_X2Y4_LUT4AB/EE4END[3]
+ Tile_X2Y4_LUT4AB/EE4END[4] Tile_X2Y4_LUT4AB/EE4END[5] Tile_X2Y4_LUT4AB/EE4END[6]
+ Tile_X2Y4_LUT4AB/EE4END[7] Tile_X2Y4_LUT4AB/EE4END[8] Tile_X2Y4_LUT4AB/EE4END[9]
+ Tile_X2Y4_LUT4AB/FrameData[0] Tile_X2Y4_LUT4AB/FrameData[10] Tile_X2Y4_LUT4AB/FrameData[11]
+ Tile_X2Y4_LUT4AB/FrameData[12] Tile_X2Y4_LUT4AB/FrameData[13] Tile_X2Y4_LUT4AB/FrameData[14]
+ Tile_X2Y4_LUT4AB/FrameData[15] Tile_X2Y4_LUT4AB/FrameData[16] Tile_X2Y4_LUT4AB/FrameData[17]
+ Tile_X2Y4_LUT4AB/FrameData[18] Tile_X2Y4_LUT4AB/FrameData[19] Tile_X2Y4_LUT4AB/FrameData[1]
+ Tile_X2Y4_LUT4AB/FrameData[20] Tile_X2Y4_LUT4AB/FrameData[21] Tile_X2Y4_LUT4AB/FrameData[22]
+ Tile_X2Y4_LUT4AB/FrameData[23] Tile_X2Y4_LUT4AB/FrameData[24] Tile_X2Y4_LUT4AB/FrameData[25]
+ Tile_X2Y4_LUT4AB/FrameData[26] Tile_X2Y4_LUT4AB/FrameData[27] Tile_X2Y4_LUT4AB/FrameData[28]
+ Tile_X2Y4_LUT4AB/FrameData[29] Tile_X2Y4_LUT4AB/FrameData[2] Tile_X2Y4_LUT4AB/FrameData[30]
+ Tile_X2Y4_LUT4AB/FrameData[31] Tile_X2Y4_LUT4AB/FrameData[3] Tile_X2Y4_LUT4AB/FrameData[4]
+ Tile_X2Y4_LUT4AB/FrameData[5] Tile_X2Y4_LUT4AB/FrameData[6] Tile_X2Y4_LUT4AB/FrameData[7]
+ Tile_X2Y4_LUT4AB/FrameData[8] Tile_X2Y4_LUT4AB/FrameData[9] Tile_X3Y4_LUT4AB/FrameData[0]
+ Tile_X3Y4_LUT4AB/FrameData[10] Tile_X3Y4_LUT4AB/FrameData[11] Tile_X3Y4_LUT4AB/FrameData[12]
+ Tile_X3Y4_LUT4AB/FrameData[13] Tile_X3Y4_LUT4AB/FrameData[14] Tile_X3Y4_LUT4AB/FrameData[15]
+ Tile_X3Y4_LUT4AB/FrameData[16] Tile_X3Y4_LUT4AB/FrameData[17] Tile_X3Y4_LUT4AB/FrameData[18]
+ Tile_X3Y4_LUT4AB/FrameData[19] Tile_X3Y4_LUT4AB/FrameData[1] Tile_X3Y4_LUT4AB/FrameData[20]
+ Tile_X3Y4_LUT4AB/FrameData[21] Tile_X3Y4_LUT4AB/FrameData[22] Tile_X3Y4_LUT4AB/FrameData[23]
+ Tile_X3Y4_LUT4AB/FrameData[24] Tile_X3Y4_LUT4AB/FrameData[25] Tile_X3Y4_LUT4AB/FrameData[26]
+ Tile_X3Y4_LUT4AB/FrameData[27] Tile_X3Y4_LUT4AB/FrameData[28] Tile_X3Y4_LUT4AB/FrameData[29]
+ Tile_X3Y4_LUT4AB/FrameData[2] Tile_X3Y4_LUT4AB/FrameData[30] Tile_X3Y4_LUT4AB/FrameData[31]
+ Tile_X3Y4_LUT4AB/FrameData[3] Tile_X3Y4_LUT4AB/FrameData[4] Tile_X3Y4_LUT4AB/FrameData[5]
+ Tile_X3Y4_LUT4AB/FrameData[6] Tile_X3Y4_LUT4AB/FrameData[7] Tile_X3Y4_LUT4AB/FrameData[8]
+ Tile_X3Y4_LUT4AB/FrameData[9] Tile_X2Y4_LUT4AB/FrameStrobe[0] Tile_X2Y4_LUT4AB/FrameStrobe[10]
+ Tile_X2Y4_LUT4AB/FrameStrobe[11] Tile_X2Y4_LUT4AB/FrameStrobe[12] Tile_X2Y4_LUT4AB/FrameStrobe[13]
+ Tile_X2Y4_LUT4AB/FrameStrobe[14] Tile_X2Y4_LUT4AB/FrameStrobe[15] Tile_X2Y4_LUT4AB/FrameStrobe[16]
+ Tile_X2Y4_LUT4AB/FrameStrobe[17] Tile_X2Y4_LUT4AB/FrameStrobe[18] Tile_X2Y4_LUT4AB/FrameStrobe[19]
+ Tile_X2Y4_LUT4AB/FrameStrobe[1] Tile_X2Y4_LUT4AB/FrameStrobe[2] Tile_X2Y4_LUT4AB/FrameStrobe[3]
+ Tile_X2Y4_LUT4AB/FrameStrobe[4] Tile_X2Y4_LUT4AB/FrameStrobe[5] Tile_X2Y4_LUT4AB/FrameStrobe[6]
+ Tile_X2Y4_LUT4AB/FrameStrobe[7] Tile_X2Y4_LUT4AB/FrameStrobe[8] Tile_X2Y4_LUT4AB/FrameStrobe[9]
+ Tile_X2Y3_LUT4AB/FrameStrobe[0] Tile_X2Y3_LUT4AB/FrameStrobe[10] Tile_X2Y3_LUT4AB/FrameStrobe[11]
+ Tile_X2Y3_LUT4AB/FrameStrobe[12] Tile_X2Y3_LUT4AB/FrameStrobe[13] Tile_X2Y3_LUT4AB/FrameStrobe[14]
+ Tile_X2Y3_LUT4AB/FrameStrobe[15] Tile_X2Y3_LUT4AB/FrameStrobe[16] Tile_X2Y3_LUT4AB/FrameStrobe[17]
+ Tile_X2Y3_LUT4AB/FrameStrobe[18] Tile_X2Y3_LUT4AB/FrameStrobe[19] Tile_X2Y3_LUT4AB/FrameStrobe[1]
+ Tile_X2Y3_LUT4AB/FrameStrobe[2] Tile_X2Y3_LUT4AB/FrameStrobe[3] Tile_X2Y3_LUT4AB/FrameStrobe[4]
+ Tile_X2Y3_LUT4AB/FrameStrobe[5] Tile_X2Y3_LUT4AB/FrameStrobe[6] Tile_X2Y3_LUT4AB/FrameStrobe[7]
+ Tile_X2Y3_LUT4AB/FrameStrobe[8] Tile_X2Y3_LUT4AB/FrameStrobe[9] Tile_X2Y4_LUT4AB/N1BEG[0]
+ Tile_X2Y4_LUT4AB/N1BEG[1] Tile_X2Y4_LUT4AB/N1BEG[2] Tile_X2Y4_LUT4AB/N1BEG[3] Tile_X2Y5_LUT4AB/N1BEG[0]
+ Tile_X2Y5_LUT4AB/N1BEG[1] Tile_X2Y5_LUT4AB/N1BEG[2] Tile_X2Y5_LUT4AB/N1BEG[3] Tile_X2Y4_LUT4AB/N2BEG[0]
+ Tile_X2Y4_LUT4AB/N2BEG[1] Tile_X2Y4_LUT4AB/N2BEG[2] Tile_X2Y4_LUT4AB/N2BEG[3] Tile_X2Y4_LUT4AB/N2BEG[4]
+ Tile_X2Y4_LUT4AB/N2BEG[5] Tile_X2Y4_LUT4AB/N2BEG[6] Tile_X2Y4_LUT4AB/N2BEG[7] Tile_X2Y3_LUT4AB/N2END[0]
+ Tile_X2Y3_LUT4AB/N2END[1] Tile_X2Y3_LUT4AB/N2END[2] Tile_X2Y3_LUT4AB/N2END[3] Tile_X2Y3_LUT4AB/N2END[4]
+ Tile_X2Y3_LUT4AB/N2END[5] Tile_X2Y3_LUT4AB/N2END[6] Tile_X2Y3_LUT4AB/N2END[7] Tile_X2Y4_LUT4AB/N2END[0]
+ Tile_X2Y4_LUT4AB/N2END[1] Tile_X2Y4_LUT4AB/N2END[2] Tile_X2Y4_LUT4AB/N2END[3] Tile_X2Y4_LUT4AB/N2END[4]
+ Tile_X2Y4_LUT4AB/N2END[5] Tile_X2Y4_LUT4AB/N2END[6] Tile_X2Y4_LUT4AB/N2END[7] Tile_X2Y5_LUT4AB/N2BEG[0]
+ Tile_X2Y5_LUT4AB/N2BEG[1] Tile_X2Y5_LUT4AB/N2BEG[2] Tile_X2Y5_LUT4AB/N2BEG[3] Tile_X2Y5_LUT4AB/N2BEG[4]
+ Tile_X2Y5_LUT4AB/N2BEG[5] Tile_X2Y5_LUT4AB/N2BEG[6] Tile_X2Y5_LUT4AB/N2BEG[7] Tile_X2Y4_LUT4AB/N4BEG[0]
+ Tile_X2Y4_LUT4AB/N4BEG[10] Tile_X2Y4_LUT4AB/N4BEG[11] Tile_X2Y4_LUT4AB/N4BEG[12]
+ Tile_X2Y4_LUT4AB/N4BEG[13] Tile_X2Y4_LUT4AB/N4BEG[14] Tile_X2Y4_LUT4AB/N4BEG[15]
+ Tile_X2Y4_LUT4AB/N4BEG[1] Tile_X2Y4_LUT4AB/N4BEG[2] Tile_X2Y4_LUT4AB/N4BEG[3] Tile_X2Y4_LUT4AB/N4BEG[4]
+ Tile_X2Y4_LUT4AB/N4BEG[5] Tile_X2Y4_LUT4AB/N4BEG[6] Tile_X2Y4_LUT4AB/N4BEG[7] Tile_X2Y4_LUT4AB/N4BEG[8]
+ Tile_X2Y4_LUT4AB/N4BEG[9] Tile_X2Y5_LUT4AB/N4BEG[0] Tile_X2Y5_LUT4AB/N4BEG[10] Tile_X2Y5_LUT4AB/N4BEG[11]
+ Tile_X2Y5_LUT4AB/N4BEG[12] Tile_X2Y5_LUT4AB/N4BEG[13] Tile_X2Y5_LUT4AB/N4BEG[14]
+ Tile_X2Y5_LUT4AB/N4BEG[15] Tile_X2Y5_LUT4AB/N4BEG[1] Tile_X2Y5_LUT4AB/N4BEG[2] Tile_X2Y5_LUT4AB/N4BEG[3]
+ Tile_X2Y5_LUT4AB/N4BEG[4] Tile_X2Y5_LUT4AB/N4BEG[5] Tile_X2Y5_LUT4AB/N4BEG[6] Tile_X2Y5_LUT4AB/N4BEG[7]
+ Tile_X2Y5_LUT4AB/N4BEG[8] Tile_X2Y5_LUT4AB/N4BEG[9] Tile_X2Y4_LUT4AB/NN4BEG[0] Tile_X2Y4_LUT4AB/NN4BEG[10]
+ Tile_X2Y4_LUT4AB/NN4BEG[11] Tile_X2Y4_LUT4AB/NN4BEG[12] Tile_X2Y4_LUT4AB/NN4BEG[13]
+ Tile_X2Y4_LUT4AB/NN4BEG[14] Tile_X2Y4_LUT4AB/NN4BEG[15] Tile_X2Y4_LUT4AB/NN4BEG[1]
+ Tile_X2Y4_LUT4AB/NN4BEG[2] Tile_X2Y4_LUT4AB/NN4BEG[3] Tile_X2Y4_LUT4AB/NN4BEG[4]
+ Tile_X2Y4_LUT4AB/NN4BEG[5] Tile_X2Y4_LUT4AB/NN4BEG[6] Tile_X2Y4_LUT4AB/NN4BEG[7]
+ Tile_X2Y4_LUT4AB/NN4BEG[8] Tile_X2Y4_LUT4AB/NN4BEG[9] Tile_X2Y5_LUT4AB/NN4BEG[0]
+ Tile_X2Y5_LUT4AB/NN4BEG[10] Tile_X2Y5_LUT4AB/NN4BEG[11] Tile_X2Y5_LUT4AB/NN4BEG[12]
+ Tile_X2Y5_LUT4AB/NN4BEG[13] Tile_X2Y5_LUT4AB/NN4BEG[14] Tile_X2Y5_LUT4AB/NN4BEG[15]
+ Tile_X2Y5_LUT4AB/NN4BEG[1] Tile_X2Y5_LUT4AB/NN4BEG[2] Tile_X2Y5_LUT4AB/NN4BEG[3]
+ Tile_X2Y5_LUT4AB/NN4BEG[4] Tile_X2Y5_LUT4AB/NN4BEG[5] Tile_X2Y5_LUT4AB/NN4BEG[6]
+ Tile_X2Y5_LUT4AB/NN4BEG[7] Tile_X2Y5_LUT4AB/NN4BEG[8] Tile_X2Y5_LUT4AB/NN4BEG[9]
+ Tile_X2Y5_LUT4AB/S1END[0] Tile_X2Y5_LUT4AB/S1END[1] Tile_X2Y5_LUT4AB/S1END[2] Tile_X2Y5_LUT4AB/S1END[3]
+ Tile_X2Y4_LUT4AB/S1END[0] Tile_X2Y4_LUT4AB/S1END[1] Tile_X2Y4_LUT4AB/S1END[2] Tile_X2Y4_LUT4AB/S1END[3]
+ Tile_X2Y5_LUT4AB/S2MID[0] Tile_X2Y5_LUT4AB/S2MID[1] Tile_X2Y5_LUT4AB/S2MID[2] Tile_X2Y5_LUT4AB/S2MID[3]
+ Tile_X2Y5_LUT4AB/S2MID[4] Tile_X2Y5_LUT4AB/S2MID[5] Tile_X2Y5_LUT4AB/S2MID[6] Tile_X2Y5_LUT4AB/S2MID[7]
+ Tile_X2Y5_LUT4AB/S2END[0] Tile_X2Y5_LUT4AB/S2END[1] Tile_X2Y5_LUT4AB/S2END[2] Tile_X2Y5_LUT4AB/S2END[3]
+ Tile_X2Y5_LUT4AB/S2END[4] Tile_X2Y5_LUT4AB/S2END[5] Tile_X2Y5_LUT4AB/S2END[6] Tile_X2Y5_LUT4AB/S2END[7]
+ Tile_X2Y4_LUT4AB/S2END[0] Tile_X2Y4_LUT4AB/S2END[1] Tile_X2Y4_LUT4AB/S2END[2] Tile_X2Y4_LUT4AB/S2END[3]
+ Tile_X2Y4_LUT4AB/S2END[4] Tile_X2Y4_LUT4AB/S2END[5] Tile_X2Y4_LUT4AB/S2END[6] Tile_X2Y4_LUT4AB/S2END[7]
+ Tile_X2Y4_LUT4AB/S2MID[0] Tile_X2Y4_LUT4AB/S2MID[1] Tile_X2Y4_LUT4AB/S2MID[2] Tile_X2Y4_LUT4AB/S2MID[3]
+ Tile_X2Y4_LUT4AB/S2MID[4] Tile_X2Y4_LUT4AB/S2MID[5] Tile_X2Y4_LUT4AB/S2MID[6] Tile_X2Y4_LUT4AB/S2MID[7]
+ Tile_X2Y5_LUT4AB/S4END[0] Tile_X2Y5_LUT4AB/S4END[10] Tile_X2Y5_LUT4AB/S4END[11]
+ Tile_X2Y5_LUT4AB/S4END[12] Tile_X2Y5_LUT4AB/S4END[13] Tile_X2Y5_LUT4AB/S4END[14]
+ Tile_X2Y5_LUT4AB/S4END[15] Tile_X2Y5_LUT4AB/S4END[1] Tile_X2Y5_LUT4AB/S4END[2] Tile_X2Y5_LUT4AB/S4END[3]
+ Tile_X2Y5_LUT4AB/S4END[4] Tile_X2Y5_LUT4AB/S4END[5] Tile_X2Y5_LUT4AB/S4END[6] Tile_X2Y5_LUT4AB/S4END[7]
+ Tile_X2Y5_LUT4AB/S4END[8] Tile_X2Y5_LUT4AB/S4END[9] Tile_X2Y4_LUT4AB/S4END[0] Tile_X2Y4_LUT4AB/S4END[10]
+ Tile_X2Y4_LUT4AB/S4END[11] Tile_X2Y4_LUT4AB/S4END[12] Tile_X2Y4_LUT4AB/S4END[13]
+ Tile_X2Y4_LUT4AB/S4END[14] Tile_X2Y4_LUT4AB/S4END[15] Tile_X2Y4_LUT4AB/S4END[1]
+ Tile_X2Y4_LUT4AB/S4END[2] Tile_X2Y4_LUT4AB/S4END[3] Tile_X2Y4_LUT4AB/S4END[4] Tile_X2Y4_LUT4AB/S4END[5]
+ Tile_X2Y4_LUT4AB/S4END[6] Tile_X2Y4_LUT4AB/S4END[7] Tile_X2Y4_LUT4AB/S4END[8] Tile_X2Y4_LUT4AB/S4END[9]
+ Tile_X2Y5_LUT4AB/SS4END[0] Tile_X2Y5_LUT4AB/SS4END[10] Tile_X2Y5_LUT4AB/SS4END[11]
+ Tile_X2Y5_LUT4AB/SS4END[12] Tile_X2Y5_LUT4AB/SS4END[13] Tile_X2Y5_LUT4AB/SS4END[14]
+ Tile_X2Y5_LUT4AB/SS4END[15] Tile_X2Y5_LUT4AB/SS4END[1] Tile_X2Y5_LUT4AB/SS4END[2]
+ Tile_X2Y5_LUT4AB/SS4END[3] Tile_X2Y5_LUT4AB/SS4END[4] Tile_X2Y5_LUT4AB/SS4END[5]
+ Tile_X2Y5_LUT4AB/SS4END[6] Tile_X2Y5_LUT4AB/SS4END[7] Tile_X2Y5_LUT4AB/SS4END[8]
+ Tile_X2Y5_LUT4AB/SS4END[9] Tile_X2Y4_LUT4AB/SS4END[0] Tile_X2Y4_LUT4AB/SS4END[10]
+ Tile_X2Y4_LUT4AB/SS4END[11] Tile_X2Y4_LUT4AB/SS4END[12] Tile_X2Y4_LUT4AB/SS4END[13]
+ Tile_X2Y4_LUT4AB/SS4END[14] Tile_X2Y4_LUT4AB/SS4END[15] Tile_X2Y4_LUT4AB/SS4END[1]
+ Tile_X2Y4_LUT4AB/SS4END[2] Tile_X2Y4_LUT4AB/SS4END[3] Tile_X2Y4_LUT4AB/SS4END[4]
+ Tile_X2Y4_LUT4AB/SS4END[5] Tile_X2Y4_LUT4AB/SS4END[6] Tile_X2Y4_LUT4AB/SS4END[7]
+ Tile_X2Y4_LUT4AB/SS4END[8] Tile_X2Y4_LUT4AB/SS4END[9] Tile_X2Y4_LUT4AB/UserCLK Tile_X2Y3_LUT4AB/UserCLK
+ VGND VPWR Tile_X2Y4_LUT4AB/W1BEG[0] Tile_X2Y4_LUT4AB/W1BEG[1] Tile_X2Y4_LUT4AB/W1BEG[2]
+ Tile_X2Y4_LUT4AB/W1BEG[3] Tile_X3Y4_LUT4AB/W1BEG[0] Tile_X3Y4_LUT4AB/W1BEG[1] Tile_X3Y4_LUT4AB/W1BEG[2]
+ Tile_X3Y4_LUT4AB/W1BEG[3] Tile_X2Y4_LUT4AB/W2BEG[0] Tile_X2Y4_LUT4AB/W2BEG[1] Tile_X2Y4_LUT4AB/W2BEG[2]
+ Tile_X2Y4_LUT4AB/W2BEG[3] Tile_X2Y4_LUT4AB/W2BEG[4] Tile_X2Y4_LUT4AB/W2BEG[5] Tile_X2Y4_LUT4AB/W2BEG[6]
+ Tile_X2Y4_LUT4AB/W2BEG[7] Tile_X1Y4_LUT4AB/W2END[0] Tile_X1Y4_LUT4AB/W2END[1] Tile_X1Y4_LUT4AB/W2END[2]
+ Tile_X1Y4_LUT4AB/W2END[3] Tile_X1Y4_LUT4AB/W2END[4] Tile_X1Y4_LUT4AB/W2END[5] Tile_X1Y4_LUT4AB/W2END[6]
+ Tile_X1Y4_LUT4AB/W2END[7] Tile_X2Y4_LUT4AB/W2END[0] Tile_X2Y4_LUT4AB/W2END[1] Tile_X2Y4_LUT4AB/W2END[2]
+ Tile_X2Y4_LUT4AB/W2END[3] Tile_X2Y4_LUT4AB/W2END[4] Tile_X2Y4_LUT4AB/W2END[5] Tile_X2Y4_LUT4AB/W2END[6]
+ Tile_X2Y4_LUT4AB/W2END[7] Tile_X3Y4_LUT4AB/W2BEG[0] Tile_X3Y4_LUT4AB/W2BEG[1] Tile_X3Y4_LUT4AB/W2BEG[2]
+ Tile_X3Y4_LUT4AB/W2BEG[3] Tile_X3Y4_LUT4AB/W2BEG[4] Tile_X3Y4_LUT4AB/W2BEG[5] Tile_X3Y4_LUT4AB/W2BEG[6]
+ Tile_X3Y4_LUT4AB/W2BEG[7] Tile_X2Y4_LUT4AB/W6BEG[0] Tile_X2Y4_LUT4AB/W6BEG[10] Tile_X2Y4_LUT4AB/W6BEG[11]
+ Tile_X2Y4_LUT4AB/W6BEG[1] Tile_X2Y4_LUT4AB/W6BEG[2] Tile_X2Y4_LUT4AB/W6BEG[3] Tile_X2Y4_LUT4AB/W6BEG[4]
+ Tile_X2Y4_LUT4AB/W6BEG[5] Tile_X2Y4_LUT4AB/W6BEG[6] Tile_X2Y4_LUT4AB/W6BEG[7] Tile_X2Y4_LUT4AB/W6BEG[8]
+ Tile_X2Y4_LUT4AB/W6BEG[9] Tile_X3Y4_LUT4AB/W6BEG[0] Tile_X3Y4_LUT4AB/W6BEG[10] Tile_X3Y4_LUT4AB/W6BEG[11]
+ Tile_X3Y4_LUT4AB/W6BEG[1] Tile_X3Y4_LUT4AB/W6BEG[2] Tile_X3Y4_LUT4AB/W6BEG[3] Tile_X3Y4_LUT4AB/W6BEG[4]
+ Tile_X3Y4_LUT4AB/W6BEG[5] Tile_X3Y4_LUT4AB/W6BEG[6] Tile_X3Y4_LUT4AB/W6BEG[7] Tile_X3Y4_LUT4AB/W6BEG[8]
+ Tile_X3Y4_LUT4AB/W6BEG[9] Tile_X2Y4_LUT4AB/WW4BEG[0] Tile_X2Y4_LUT4AB/WW4BEG[10]
+ Tile_X2Y4_LUT4AB/WW4BEG[11] Tile_X2Y4_LUT4AB/WW4BEG[12] Tile_X2Y4_LUT4AB/WW4BEG[13]
+ Tile_X2Y4_LUT4AB/WW4BEG[14] Tile_X2Y4_LUT4AB/WW4BEG[15] Tile_X2Y4_LUT4AB/WW4BEG[1]
+ Tile_X2Y4_LUT4AB/WW4BEG[2] Tile_X2Y4_LUT4AB/WW4BEG[3] Tile_X2Y4_LUT4AB/WW4BEG[4]
+ Tile_X2Y4_LUT4AB/WW4BEG[5] Tile_X2Y4_LUT4AB/WW4BEG[6] Tile_X2Y4_LUT4AB/WW4BEG[7]
+ Tile_X2Y4_LUT4AB/WW4BEG[8] Tile_X2Y4_LUT4AB/WW4BEG[9] Tile_X3Y4_LUT4AB/WW4BEG[0]
+ Tile_X3Y4_LUT4AB/WW4BEG[10] Tile_X3Y4_LUT4AB/WW4BEG[11] Tile_X3Y4_LUT4AB/WW4BEG[12]
+ Tile_X3Y4_LUT4AB/WW4BEG[13] Tile_X3Y4_LUT4AB/WW4BEG[14] Tile_X3Y4_LUT4AB/WW4BEG[15]
+ Tile_X3Y4_LUT4AB/WW4BEG[1] Tile_X3Y4_LUT4AB/WW4BEG[2] Tile_X3Y4_LUT4AB/WW4BEG[3]
+ Tile_X3Y4_LUT4AB/WW4BEG[4] Tile_X3Y4_LUT4AB/WW4BEG[5] Tile_X3Y4_LUT4AB/WW4BEG[6]
+ Tile_X3Y4_LUT4AB/WW4BEG[7] Tile_X3Y4_LUT4AB/WW4BEG[8] Tile_X3Y4_LUT4AB/WW4BEG[9]
+ LUT4AB
XTile_X7Y13_DSP Tile_X8Y13_LUT4AB/E1END[0] Tile_X8Y13_LUT4AB/E1END[1] Tile_X8Y13_LUT4AB/E1END[2]
+ Tile_X8Y13_LUT4AB/E1END[3] Tile_X6Y13_LUT4AB/E1BEG[0] Tile_X6Y13_LUT4AB/E1BEG[1]
+ Tile_X6Y13_LUT4AB/E1BEG[2] Tile_X6Y13_LUT4AB/E1BEG[3] Tile_X8Y13_LUT4AB/E2MID[0]
+ Tile_X8Y13_LUT4AB/E2MID[1] Tile_X8Y13_LUT4AB/E2MID[2] Tile_X8Y13_LUT4AB/E2MID[3]
+ Tile_X8Y13_LUT4AB/E2MID[4] Tile_X8Y13_LUT4AB/E2MID[5] Tile_X8Y13_LUT4AB/E2MID[6]
+ Tile_X8Y13_LUT4AB/E2MID[7] Tile_X8Y13_LUT4AB/E2END[0] Tile_X8Y13_LUT4AB/E2END[1]
+ Tile_X8Y13_LUT4AB/E2END[2] Tile_X8Y13_LUT4AB/E2END[3] Tile_X8Y13_LUT4AB/E2END[4]
+ Tile_X8Y13_LUT4AB/E2END[5] Tile_X8Y13_LUT4AB/E2END[6] Tile_X8Y13_LUT4AB/E2END[7]
+ Tile_X6Y13_LUT4AB/E2BEGb[0] Tile_X6Y13_LUT4AB/E2BEGb[1] Tile_X6Y13_LUT4AB/E2BEGb[2]
+ Tile_X6Y13_LUT4AB/E2BEGb[3] Tile_X6Y13_LUT4AB/E2BEGb[4] Tile_X6Y13_LUT4AB/E2BEGb[5]
+ Tile_X6Y13_LUT4AB/E2BEGb[6] Tile_X6Y13_LUT4AB/E2BEGb[7] Tile_X6Y13_LUT4AB/E2BEG[0]
+ Tile_X6Y13_LUT4AB/E2BEG[1] Tile_X6Y13_LUT4AB/E2BEG[2] Tile_X6Y13_LUT4AB/E2BEG[3]
+ Tile_X6Y13_LUT4AB/E2BEG[4] Tile_X6Y13_LUT4AB/E2BEG[5] Tile_X6Y13_LUT4AB/E2BEG[6]
+ Tile_X6Y13_LUT4AB/E2BEG[7] Tile_X8Y13_LUT4AB/E6END[0] Tile_X8Y13_LUT4AB/E6END[10]
+ Tile_X8Y13_LUT4AB/E6END[11] Tile_X8Y13_LUT4AB/E6END[1] Tile_X8Y13_LUT4AB/E6END[2]
+ Tile_X8Y13_LUT4AB/E6END[3] Tile_X8Y13_LUT4AB/E6END[4] Tile_X8Y13_LUT4AB/E6END[5]
+ Tile_X8Y13_LUT4AB/E6END[6] Tile_X8Y13_LUT4AB/E6END[7] Tile_X8Y13_LUT4AB/E6END[8]
+ Tile_X8Y13_LUT4AB/E6END[9] Tile_X6Y13_LUT4AB/E6BEG[0] Tile_X6Y13_LUT4AB/E6BEG[10]
+ Tile_X6Y13_LUT4AB/E6BEG[11] Tile_X6Y13_LUT4AB/E6BEG[1] Tile_X6Y13_LUT4AB/E6BEG[2]
+ Tile_X6Y13_LUT4AB/E6BEG[3] Tile_X6Y13_LUT4AB/E6BEG[4] Tile_X6Y13_LUT4AB/E6BEG[5]
+ Tile_X6Y13_LUT4AB/E6BEG[6] Tile_X6Y13_LUT4AB/E6BEG[7] Tile_X6Y13_LUT4AB/E6BEG[8]
+ Tile_X6Y13_LUT4AB/E6BEG[9] Tile_X8Y13_LUT4AB/EE4END[0] Tile_X8Y13_LUT4AB/EE4END[10]
+ Tile_X8Y13_LUT4AB/EE4END[11] Tile_X8Y13_LUT4AB/EE4END[12] Tile_X8Y13_LUT4AB/EE4END[13]
+ Tile_X8Y13_LUT4AB/EE4END[14] Tile_X8Y13_LUT4AB/EE4END[15] Tile_X8Y13_LUT4AB/EE4END[1]
+ Tile_X8Y13_LUT4AB/EE4END[2] Tile_X8Y13_LUT4AB/EE4END[3] Tile_X8Y13_LUT4AB/EE4END[4]
+ Tile_X8Y13_LUT4AB/EE4END[5] Tile_X8Y13_LUT4AB/EE4END[6] Tile_X8Y13_LUT4AB/EE4END[7]
+ Tile_X8Y13_LUT4AB/EE4END[8] Tile_X8Y13_LUT4AB/EE4END[9] Tile_X6Y13_LUT4AB/EE4BEG[0]
+ Tile_X6Y13_LUT4AB/EE4BEG[10] Tile_X6Y13_LUT4AB/EE4BEG[11] Tile_X6Y13_LUT4AB/EE4BEG[12]
+ Tile_X6Y13_LUT4AB/EE4BEG[13] Tile_X6Y13_LUT4AB/EE4BEG[14] Tile_X6Y13_LUT4AB/EE4BEG[15]
+ Tile_X6Y13_LUT4AB/EE4BEG[1] Tile_X6Y13_LUT4AB/EE4BEG[2] Tile_X6Y13_LUT4AB/EE4BEG[3]
+ Tile_X6Y13_LUT4AB/EE4BEG[4] Tile_X6Y13_LUT4AB/EE4BEG[5] Tile_X6Y13_LUT4AB/EE4BEG[6]
+ Tile_X6Y13_LUT4AB/EE4BEG[7] Tile_X6Y13_LUT4AB/EE4BEG[8] Tile_X6Y13_LUT4AB/EE4BEG[9]
+ Tile_X6Y13_LUT4AB/FrameData_O[0] Tile_X6Y13_LUT4AB/FrameData_O[10] Tile_X6Y13_LUT4AB/FrameData_O[11]
+ Tile_X6Y13_LUT4AB/FrameData_O[12] Tile_X6Y13_LUT4AB/FrameData_O[13] Tile_X6Y13_LUT4AB/FrameData_O[14]
+ Tile_X6Y13_LUT4AB/FrameData_O[15] Tile_X6Y13_LUT4AB/FrameData_O[16] Tile_X6Y13_LUT4AB/FrameData_O[17]
+ Tile_X6Y13_LUT4AB/FrameData_O[18] Tile_X6Y13_LUT4AB/FrameData_O[19] Tile_X6Y13_LUT4AB/FrameData_O[1]
+ Tile_X6Y13_LUT4AB/FrameData_O[20] Tile_X6Y13_LUT4AB/FrameData_O[21] Tile_X6Y13_LUT4AB/FrameData_O[22]
+ Tile_X6Y13_LUT4AB/FrameData_O[23] Tile_X6Y13_LUT4AB/FrameData_O[24] Tile_X6Y13_LUT4AB/FrameData_O[25]
+ Tile_X6Y13_LUT4AB/FrameData_O[26] Tile_X6Y13_LUT4AB/FrameData_O[27] Tile_X6Y13_LUT4AB/FrameData_O[28]
+ Tile_X6Y13_LUT4AB/FrameData_O[29] Tile_X6Y13_LUT4AB/FrameData_O[2] Tile_X6Y13_LUT4AB/FrameData_O[30]
+ Tile_X6Y13_LUT4AB/FrameData_O[31] Tile_X6Y13_LUT4AB/FrameData_O[3] Tile_X6Y13_LUT4AB/FrameData_O[4]
+ Tile_X6Y13_LUT4AB/FrameData_O[5] Tile_X6Y13_LUT4AB/FrameData_O[6] Tile_X6Y13_LUT4AB/FrameData_O[7]
+ Tile_X6Y13_LUT4AB/FrameData_O[8] Tile_X6Y13_LUT4AB/FrameData_O[9] Tile_X8Y13_LUT4AB/FrameData[0]
+ Tile_X8Y13_LUT4AB/FrameData[10] Tile_X8Y13_LUT4AB/FrameData[11] Tile_X8Y13_LUT4AB/FrameData[12]
+ Tile_X8Y13_LUT4AB/FrameData[13] Tile_X8Y13_LUT4AB/FrameData[14] Tile_X8Y13_LUT4AB/FrameData[15]
+ Tile_X8Y13_LUT4AB/FrameData[16] Tile_X8Y13_LUT4AB/FrameData[17] Tile_X8Y13_LUT4AB/FrameData[18]
+ Tile_X8Y13_LUT4AB/FrameData[19] Tile_X8Y13_LUT4AB/FrameData[1] Tile_X8Y13_LUT4AB/FrameData[20]
+ Tile_X8Y13_LUT4AB/FrameData[21] Tile_X8Y13_LUT4AB/FrameData[22] Tile_X8Y13_LUT4AB/FrameData[23]
+ Tile_X8Y13_LUT4AB/FrameData[24] Tile_X8Y13_LUT4AB/FrameData[25] Tile_X8Y13_LUT4AB/FrameData[26]
+ Tile_X8Y13_LUT4AB/FrameData[27] Tile_X8Y13_LUT4AB/FrameData[28] Tile_X8Y13_LUT4AB/FrameData[29]
+ Tile_X8Y13_LUT4AB/FrameData[2] Tile_X8Y13_LUT4AB/FrameData[30] Tile_X8Y13_LUT4AB/FrameData[31]
+ Tile_X8Y13_LUT4AB/FrameData[3] Tile_X8Y13_LUT4AB/FrameData[4] Tile_X8Y13_LUT4AB/FrameData[5]
+ Tile_X8Y13_LUT4AB/FrameData[6] Tile_X8Y13_LUT4AB/FrameData[7] Tile_X8Y13_LUT4AB/FrameData[8]
+ Tile_X8Y13_LUT4AB/FrameData[9] Tile_X7Y11_DSP/Tile_X0Y1_FrameStrobe[0] Tile_X7Y11_DSP/Tile_X0Y1_FrameStrobe[10]
+ Tile_X7Y11_DSP/Tile_X0Y1_FrameStrobe[11] Tile_X7Y11_DSP/Tile_X0Y1_FrameStrobe[12]
+ Tile_X7Y11_DSP/Tile_X0Y1_FrameStrobe[13] Tile_X7Y11_DSP/Tile_X0Y1_FrameStrobe[14]
+ Tile_X7Y11_DSP/Tile_X0Y1_FrameStrobe[15] Tile_X7Y11_DSP/Tile_X0Y1_FrameStrobe[16]
+ Tile_X7Y11_DSP/Tile_X0Y1_FrameStrobe[17] Tile_X7Y11_DSP/Tile_X0Y1_FrameStrobe[18]
+ Tile_X7Y11_DSP/Tile_X0Y1_FrameStrobe[19] Tile_X7Y11_DSP/Tile_X0Y1_FrameStrobe[1]
+ Tile_X7Y11_DSP/Tile_X0Y1_FrameStrobe[2] Tile_X7Y11_DSP/Tile_X0Y1_FrameStrobe[3]
+ Tile_X7Y11_DSP/Tile_X0Y1_FrameStrobe[4] Tile_X7Y11_DSP/Tile_X0Y1_FrameStrobe[5]
+ Tile_X7Y11_DSP/Tile_X0Y1_FrameStrobe[6] Tile_X7Y11_DSP/Tile_X0Y1_FrameStrobe[7]
+ Tile_X7Y11_DSP/Tile_X0Y1_FrameStrobe[8] Tile_X7Y11_DSP/Tile_X0Y1_FrameStrobe[9]
+ Tile_X7Y13_DSP/Tile_X0Y0_N1BEG[0] Tile_X7Y13_DSP/Tile_X0Y0_N1BEG[1] Tile_X7Y13_DSP/Tile_X0Y0_N1BEG[2]
+ Tile_X7Y13_DSP/Tile_X0Y0_N1BEG[3] Tile_X7Y13_DSP/Tile_X0Y0_N2BEG[0] Tile_X7Y13_DSP/Tile_X0Y0_N2BEG[1]
+ Tile_X7Y13_DSP/Tile_X0Y0_N2BEG[2] Tile_X7Y13_DSP/Tile_X0Y0_N2BEG[3] Tile_X7Y13_DSP/Tile_X0Y0_N2BEG[4]
+ Tile_X7Y13_DSP/Tile_X0Y0_N2BEG[5] Tile_X7Y13_DSP/Tile_X0Y0_N2BEG[6] Tile_X7Y13_DSP/Tile_X0Y0_N2BEG[7]
+ Tile_X7Y11_DSP/Tile_X0Y1_N2END[0] Tile_X7Y11_DSP/Tile_X0Y1_N2END[1] Tile_X7Y11_DSP/Tile_X0Y1_N2END[2]
+ Tile_X7Y11_DSP/Tile_X0Y1_N2END[3] Tile_X7Y11_DSP/Tile_X0Y1_N2END[4] Tile_X7Y11_DSP/Tile_X0Y1_N2END[5]
+ Tile_X7Y11_DSP/Tile_X0Y1_N2END[6] Tile_X7Y11_DSP/Tile_X0Y1_N2END[7] Tile_X7Y13_DSP/Tile_X0Y0_N4BEG[0]
+ Tile_X7Y13_DSP/Tile_X0Y0_N4BEG[10] Tile_X7Y13_DSP/Tile_X0Y0_N4BEG[11] Tile_X7Y13_DSP/Tile_X0Y0_N4BEG[12]
+ Tile_X7Y13_DSP/Tile_X0Y0_N4BEG[13] Tile_X7Y13_DSP/Tile_X0Y0_N4BEG[14] Tile_X7Y13_DSP/Tile_X0Y0_N4BEG[15]
+ Tile_X7Y13_DSP/Tile_X0Y0_N4BEG[1] Tile_X7Y13_DSP/Tile_X0Y0_N4BEG[2] Tile_X7Y13_DSP/Tile_X0Y0_N4BEG[3]
+ Tile_X7Y13_DSP/Tile_X0Y0_N4BEG[4] Tile_X7Y13_DSP/Tile_X0Y0_N4BEG[5] Tile_X7Y13_DSP/Tile_X0Y0_N4BEG[6]
+ Tile_X7Y13_DSP/Tile_X0Y0_N4BEG[7] Tile_X7Y13_DSP/Tile_X0Y0_N4BEG[8] Tile_X7Y13_DSP/Tile_X0Y0_N4BEG[9]
+ Tile_X7Y13_DSP/Tile_X0Y0_NN4BEG[0] Tile_X7Y13_DSP/Tile_X0Y0_NN4BEG[10] Tile_X7Y13_DSP/Tile_X0Y0_NN4BEG[11]
+ Tile_X7Y13_DSP/Tile_X0Y0_NN4BEG[12] Tile_X7Y13_DSP/Tile_X0Y0_NN4BEG[13] Tile_X7Y13_DSP/Tile_X0Y0_NN4BEG[14]
+ Tile_X7Y13_DSP/Tile_X0Y0_NN4BEG[15] Tile_X7Y13_DSP/Tile_X0Y0_NN4BEG[1] Tile_X7Y13_DSP/Tile_X0Y0_NN4BEG[2]
+ Tile_X7Y13_DSP/Tile_X0Y0_NN4BEG[3] Tile_X7Y13_DSP/Tile_X0Y0_NN4BEG[4] Tile_X7Y13_DSP/Tile_X0Y0_NN4BEG[5]
+ Tile_X7Y13_DSP/Tile_X0Y0_NN4BEG[6] Tile_X7Y13_DSP/Tile_X0Y0_NN4BEG[7] Tile_X7Y13_DSP/Tile_X0Y0_NN4BEG[8]
+ Tile_X7Y13_DSP/Tile_X0Y0_NN4BEG[9] Tile_X7Y13_DSP/Tile_X0Y0_S1END[0] Tile_X7Y13_DSP/Tile_X0Y0_S1END[1]
+ Tile_X7Y13_DSP/Tile_X0Y0_S1END[2] Tile_X7Y13_DSP/Tile_X0Y0_S1END[3] Tile_X7Y13_DSP/Tile_X0Y0_S2END[0]
+ Tile_X7Y13_DSP/Tile_X0Y0_S2END[1] Tile_X7Y13_DSP/Tile_X0Y0_S2END[2] Tile_X7Y13_DSP/Tile_X0Y0_S2END[3]
+ Tile_X7Y13_DSP/Tile_X0Y0_S2END[4] Tile_X7Y13_DSP/Tile_X0Y0_S2END[5] Tile_X7Y13_DSP/Tile_X0Y0_S2END[6]
+ Tile_X7Y13_DSP/Tile_X0Y0_S2END[7] Tile_X7Y13_DSP/Tile_X0Y0_S2MID[0] Tile_X7Y13_DSP/Tile_X0Y0_S2MID[1]
+ Tile_X7Y13_DSP/Tile_X0Y0_S2MID[2] Tile_X7Y13_DSP/Tile_X0Y0_S2MID[3] Tile_X7Y13_DSP/Tile_X0Y0_S2MID[4]
+ Tile_X7Y13_DSP/Tile_X0Y0_S2MID[5] Tile_X7Y13_DSP/Tile_X0Y0_S2MID[6] Tile_X7Y13_DSP/Tile_X0Y0_S2MID[7]
+ Tile_X7Y13_DSP/Tile_X0Y0_S4END[0] Tile_X7Y13_DSP/Tile_X0Y0_S4END[10] Tile_X7Y13_DSP/Tile_X0Y0_S4END[11]
+ Tile_X7Y13_DSP/Tile_X0Y0_S4END[12] Tile_X7Y13_DSP/Tile_X0Y0_S4END[13] Tile_X7Y13_DSP/Tile_X0Y0_S4END[14]
+ Tile_X7Y13_DSP/Tile_X0Y0_S4END[15] Tile_X7Y13_DSP/Tile_X0Y0_S4END[1] Tile_X7Y13_DSP/Tile_X0Y0_S4END[2]
+ Tile_X7Y13_DSP/Tile_X0Y0_S4END[3] Tile_X7Y13_DSP/Tile_X0Y0_S4END[4] Tile_X7Y13_DSP/Tile_X0Y0_S4END[5]
+ Tile_X7Y13_DSP/Tile_X0Y0_S4END[6] Tile_X7Y13_DSP/Tile_X0Y0_S4END[7] Tile_X7Y13_DSP/Tile_X0Y0_S4END[8]
+ Tile_X7Y13_DSP/Tile_X0Y0_S4END[9] Tile_X7Y13_DSP/Tile_X0Y0_SS4END[0] Tile_X7Y13_DSP/Tile_X0Y0_SS4END[10]
+ Tile_X7Y13_DSP/Tile_X0Y0_SS4END[11] Tile_X7Y13_DSP/Tile_X0Y0_SS4END[12] Tile_X7Y13_DSP/Tile_X0Y0_SS4END[13]
+ Tile_X7Y13_DSP/Tile_X0Y0_SS4END[14] Tile_X7Y13_DSP/Tile_X0Y0_SS4END[15] Tile_X7Y13_DSP/Tile_X0Y0_SS4END[1]
+ Tile_X7Y13_DSP/Tile_X0Y0_SS4END[2] Tile_X7Y13_DSP/Tile_X0Y0_SS4END[3] Tile_X7Y13_DSP/Tile_X0Y0_SS4END[4]
+ Tile_X7Y13_DSP/Tile_X0Y0_SS4END[5] Tile_X7Y13_DSP/Tile_X0Y0_SS4END[6] Tile_X7Y13_DSP/Tile_X0Y0_SS4END[7]
+ Tile_X7Y13_DSP/Tile_X0Y0_SS4END[8] Tile_X7Y13_DSP/Tile_X0Y0_SS4END[9] Tile_X7Y11_DSP/Tile_X0Y1_UserCLK
+ Tile_X6Y13_LUT4AB/W1END[0] Tile_X6Y13_LUT4AB/W1END[1] Tile_X6Y13_LUT4AB/W1END[2]
+ Tile_X6Y13_LUT4AB/W1END[3] Tile_X8Y13_LUT4AB/W1BEG[0] Tile_X8Y13_LUT4AB/W1BEG[1]
+ Tile_X8Y13_LUT4AB/W1BEG[2] Tile_X8Y13_LUT4AB/W1BEG[3] Tile_X6Y13_LUT4AB/W2MID[0]
+ Tile_X6Y13_LUT4AB/W2MID[1] Tile_X6Y13_LUT4AB/W2MID[2] Tile_X6Y13_LUT4AB/W2MID[3]
+ Tile_X6Y13_LUT4AB/W2MID[4] Tile_X6Y13_LUT4AB/W2MID[5] Tile_X6Y13_LUT4AB/W2MID[6]
+ Tile_X6Y13_LUT4AB/W2MID[7] Tile_X6Y13_LUT4AB/W2END[0] Tile_X6Y13_LUT4AB/W2END[1]
+ Tile_X6Y13_LUT4AB/W2END[2] Tile_X6Y13_LUT4AB/W2END[3] Tile_X6Y13_LUT4AB/W2END[4]
+ Tile_X6Y13_LUT4AB/W2END[5] Tile_X6Y13_LUT4AB/W2END[6] Tile_X6Y13_LUT4AB/W2END[7]
+ Tile_X8Y13_LUT4AB/W2BEGb[0] Tile_X8Y13_LUT4AB/W2BEGb[1] Tile_X8Y13_LUT4AB/W2BEGb[2]
+ Tile_X8Y13_LUT4AB/W2BEGb[3] Tile_X8Y13_LUT4AB/W2BEGb[4] Tile_X8Y13_LUT4AB/W2BEGb[5]
+ Tile_X8Y13_LUT4AB/W2BEGb[6] Tile_X8Y13_LUT4AB/W2BEGb[7] Tile_X8Y13_LUT4AB/W2BEG[0]
+ Tile_X8Y13_LUT4AB/W2BEG[1] Tile_X8Y13_LUT4AB/W2BEG[2] Tile_X8Y13_LUT4AB/W2BEG[3]
+ Tile_X8Y13_LUT4AB/W2BEG[4] Tile_X8Y13_LUT4AB/W2BEG[5] Tile_X8Y13_LUT4AB/W2BEG[6]
+ Tile_X8Y13_LUT4AB/W2BEG[7] Tile_X6Y13_LUT4AB/W6END[0] Tile_X6Y13_LUT4AB/W6END[10]
+ Tile_X6Y13_LUT4AB/W6END[11] Tile_X6Y13_LUT4AB/W6END[1] Tile_X6Y13_LUT4AB/W6END[2]
+ Tile_X6Y13_LUT4AB/W6END[3] Tile_X6Y13_LUT4AB/W6END[4] Tile_X6Y13_LUT4AB/W6END[5]
+ Tile_X6Y13_LUT4AB/W6END[6] Tile_X6Y13_LUT4AB/W6END[7] Tile_X6Y13_LUT4AB/W6END[8]
+ Tile_X6Y13_LUT4AB/W6END[9] Tile_X8Y13_LUT4AB/W6BEG[0] Tile_X8Y13_LUT4AB/W6BEG[10]
+ Tile_X8Y13_LUT4AB/W6BEG[11] Tile_X8Y13_LUT4AB/W6BEG[1] Tile_X8Y13_LUT4AB/W6BEG[2]
+ Tile_X8Y13_LUT4AB/W6BEG[3] Tile_X8Y13_LUT4AB/W6BEG[4] Tile_X8Y13_LUT4AB/W6BEG[5]
+ Tile_X8Y13_LUT4AB/W6BEG[6] Tile_X8Y13_LUT4AB/W6BEG[7] Tile_X8Y13_LUT4AB/W6BEG[8]
+ Tile_X8Y13_LUT4AB/W6BEG[9] Tile_X6Y13_LUT4AB/WW4END[0] Tile_X6Y13_LUT4AB/WW4END[10]
+ Tile_X6Y13_LUT4AB/WW4END[11] Tile_X6Y13_LUT4AB/WW4END[12] Tile_X6Y13_LUT4AB/WW4END[13]
+ Tile_X6Y13_LUT4AB/WW4END[14] Tile_X6Y13_LUT4AB/WW4END[15] Tile_X6Y13_LUT4AB/WW4END[1]
+ Tile_X6Y13_LUT4AB/WW4END[2] Tile_X6Y13_LUT4AB/WW4END[3] Tile_X6Y13_LUT4AB/WW4END[4]
+ Tile_X6Y13_LUT4AB/WW4END[5] Tile_X6Y13_LUT4AB/WW4END[6] Tile_X6Y13_LUT4AB/WW4END[7]
+ Tile_X6Y13_LUT4AB/WW4END[8] Tile_X6Y13_LUT4AB/WW4END[9] Tile_X8Y13_LUT4AB/WW4BEG[0]
+ Tile_X8Y13_LUT4AB/WW4BEG[10] Tile_X8Y13_LUT4AB/WW4BEG[11] Tile_X8Y13_LUT4AB/WW4BEG[12]
+ Tile_X8Y13_LUT4AB/WW4BEG[13] Tile_X8Y13_LUT4AB/WW4BEG[14] Tile_X8Y13_LUT4AB/WW4BEG[15]
+ Tile_X8Y13_LUT4AB/WW4BEG[1] Tile_X8Y13_LUT4AB/WW4BEG[2] Tile_X8Y13_LUT4AB/WW4BEG[3]
+ Tile_X8Y13_LUT4AB/WW4BEG[4] Tile_X8Y13_LUT4AB/WW4BEG[5] Tile_X8Y13_LUT4AB/WW4BEG[6]
+ Tile_X8Y13_LUT4AB/WW4BEG[7] Tile_X8Y13_LUT4AB/WW4BEG[8] Tile_X8Y13_LUT4AB/WW4BEG[9]
+ Tile_X8Y14_LUT4AB/E1END[0] Tile_X8Y14_LUT4AB/E1END[1] Tile_X8Y14_LUT4AB/E1END[2]
+ Tile_X8Y14_LUT4AB/E1END[3] Tile_X6Y14_LUT4AB/E1BEG[0] Tile_X6Y14_LUT4AB/E1BEG[1]
+ Tile_X6Y14_LUT4AB/E1BEG[2] Tile_X6Y14_LUT4AB/E1BEG[3] Tile_X8Y14_LUT4AB/E2MID[0]
+ Tile_X8Y14_LUT4AB/E2MID[1] Tile_X8Y14_LUT4AB/E2MID[2] Tile_X8Y14_LUT4AB/E2MID[3]
+ Tile_X8Y14_LUT4AB/E2MID[4] Tile_X8Y14_LUT4AB/E2MID[5] Tile_X8Y14_LUT4AB/E2MID[6]
+ Tile_X8Y14_LUT4AB/E2MID[7] Tile_X8Y14_LUT4AB/E2END[0] Tile_X8Y14_LUT4AB/E2END[1]
+ Tile_X8Y14_LUT4AB/E2END[2] Tile_X8Y14_LUT4AB/E2END[3] Tile_X8Y14_LUT4AB/E2END[4]
+ Tile_X8Y14_LUT4AB/E2END[5] Tile_X8Y14_LUT4AB/E2END[6] Tile_X8Y14_LUT4AB/E2END[7]
+ Tile_X6Y14_LUT4AB/E2BEGb[0] Tile_X6Y14_LUT4AB/E2BEGb[1] Tile_X6Y14_LUT4AB/E2BEGb[2]
+ Tile_X6Y14_LUT4AB/E2BEGb[3] Tile_X6Y14_LUT4AB/E2BEGb[4] Tile_X6Y14_LUT4AB/E2BEGb[5]
+ Tile_X6Y14_LUT4AB/E2BEGb[6] Tile_X6Y14_LUT4AB/E2BEGb[7] Tile_X6Y14_LUT4AB/E2BEG[0]
+ Tile_X6Y14_LUT4AB/E2BEG[1] Tile_X6Y14_LUT4AB/E2BEG[2] Tile_X6Y14_LUT4AB/E2BEG[3]
+ Tile_X6Y14_LUT4AB/E2BEG[4] Tile_X6Y14_LUT4AB/E2BEG[5] Tile_X6Y14_LUT4AB/E2BEG[6]
+ Tile_X6Y14_LUT4AB/E2BEG[7] Tile_X8Y14_LUT4AB/E6END[0] Tile_X8Y14_LUT4AB/E6END[10]
+ Tile_X8Y14_LUT4AB/E6END[11] Tile_X8Y14_LUT4AB/E6END[1] Tile_X8Y14_LUT4AB/E6END[2]
+ Tile_X8Y14_LUT4AB/E6END[3] Tile_X8Y14_LUT4AB/E6END[4] Tile_X8Y14_LUT4AB/E6END[5]
+ Tile_X8Y14_LUT4AB/E6END[6] Tile_X8Y14_LUT4AB/E6END[7] Tile_X8Y14_LUT4AB/E6END[8]
+ Tile_X8Y14_LUT4AB/E6END[9] Tile_X6Y14_LUT4AB/E6BEG[0] Tile_X6Y14_LUT4AB/E6BEG[10]
+ Tile_X6Y14_LUT4AB/E6BEG[11] Tile_X6Y14_LUT4AB/E6BEG[1] Tile_X6Y14_LUT4AB/E6BEG[2]
+ Tile_X6Y14_LUT4AB/E6BEG[3] Tile_X6Y14_LUT4AB/E6BEG[4] Tile_X6Y14_LUT4AB/E6BEG[5]
+ Tile_X6Y14_LUT4AB/E6BEG[6] Tile_X6Y14_LUT4AB/E6BEG[7] Tile_X6Y14_LUT4AB/E6BEG[8]
+ Tile_X6Y14_LUT4AB/E6BEG[9] Tile_X8Y14_LUT4AB/EE4END[0] Tile_X8Y14_LUT4AB/EE4END[10]
+ Tile_X8Y14_LUT4AB/EE4END[11] Tile_X8Y14_LUT4AB/EE4END[12] Tile_X8Y14_LUT4AB/EE4END[13]
+ Tile_X8Y14_LUT4AB/EE4END[14] Tile_X8Y14_LUT4AB/EE4END[15] Tile_X8Y14_LUT4AB/EE4END[1]
+ Tile_X8Y14_LUT4AB/EE4END[2] Tile_X8Y14_LUT4AB/EE4END[3] Tile_X8Y14_LUT4AB/EE4END[4]
+ Tile_X8Y14_LUT4AB/EE4END[5] Tile_X8Y14_LUT4AB/EE4END[6] Tile_X8Y14_LUT4AB/EE4END[7]
+ Tile_X8Y14_LUT4AB/EE4END[8] Tile_X8Y14_LUT4AB/EE4END[9] Tile_X6Y14_LUT4AB/EE4BEG[0]
+ Tile_X6Y14_LUT4AB/EE4BEG[10] Tile_X6Y14_LUT4AB/EE4BEG[11] Tile_X6Y14_LUT4AB/EE4BEG[12]
+ Tile_X6Y14_LUT4AB/EE4BEG[13] Tile_X6Y14_LUT4AB/EE4BEG[14] Tile_X6Y14_LUT4AB/EE4BEG[15]
+ Tile_X6Y14_LUT4AB/EE4BEG[1] Tile_X6Y14_LUT4AB/EE4BEG[2] Tile_X6Y14_LUT4AB/EE4BEG[3]
+ Tile_X6Y14_LUT4AB/EE4BEG[4] Tile_X6Y14_LUT4AB/EE4BEG[5] Tile_X6Y14_LUT4AB/EE4BEG[6]
+ Tile_X6Y14_LUT4AB/EE4BEG[7] Tile_X6Y14_LUT4AB/EE4BEG[8] Tile_X6Y14_LUT4AB/EE4BEG[9]
+ Tile_X6Y14_LUT4AB/FrameData_O[0] Tile_X6Y14_LUT4AB/FrameData_O[10] Tile_X6Y14_LUT4AB/FrameData_O[11]
+ Tile_X6Y14_LUT4AB/FrameData_O[12] Tile_X6Y14_LUT4AB/FrameData_O[13] Tile_X6Y14_LUT4AB/FrameData_O[14]
+ Tile_X6Y14_LUT4AB/FrameData_O[15] Tile_X6Y14_LUT4AB/FrameData_O[16] Tile_X6Y14_LUT4AB/FrameData_O[17]
+ Tile_X6Y14_LUT4AB/FrameData_O[18] Tile_X6Y14_LUT4AB/FrameData_O[19] Tile_X6Y14_LUT4AB/FrameData_O[1]
+ Tile_X6Y14_LUT4AB/FrameData_O[20] Tile_X6Y14_LUT4AB/FrameData_O[21] Tile_X6Y14_LUT4AB/FrameData_O[22]
+ Tile_X6Y14_LUT4AB/FrameData_O[23] Tile_X6Y14_LUT4AB/FrameData_O[24] Tile_X6Y14_LUT4AB/FrameData_O[25]
+ Tile_X6Y14_LUT4AB/FrameData_O[26] Tile_X6Y14_LUT4AB/FrameData_O[27] Tile_X6Y14_LUT4AB/FrameData_O[28]
+ Tile_X6Y14_LUT4AB/FrameData_O[29] Tile_X6Y14_LUT4AB/FrameData_O[2] Tile_X6Y14_LUT4AB/FrameData_O[30]
+ Tile_X6Y14_LUT4AB/FrameData_O[31] Tile_X6Y14_LUT4AB/FrameData_O[3] Tile_X6Y14_LUT4AB/FrameData_O[4]
+ Tile_X6Y14_LUT4AB/FrameData_O[5] Tile_X6Y14_LUT4AB/FrameData_O[6] Tile_X6Y14_LUT4AB/FrameData_O[7]
+ Tile_X6Y14_LUT4AB/FrameData_O[8] Tile_X6Y14_LUT4AB/FrameData_O[9] Tile_X8Y14_LUT4AB/FrameData[0]
+ Tile_X8Y14_LUT4AB/FrameData[10] Tile_X8Y14_LUT4AB/FrameData[11] Tile_X8Y14_LUT4AB/FrameData[12]
+ Tile_X8Y14_LUT4AB/FrameData[13] Tile_X8Y14_LUT4AB/FrameData[14] Tile_X8Y14_LUT4AB/FrameData[15]
+ Tile_X8Y14_LUT4AB/FrameData[16] Tile_X8Y14_LUT4AB/FrameData[17] Tile_X8Y14_LUT4AB/FrameData[18]
+ Tile_X8Y14_LUT4AB/FrameData[19] Tile_X8Y14_LUT4AB/FrameData[1] Tile_X8Y14_LUT4AB/FrameData[20]
+ Tile_X8Y14_LUT4AB/FrameData[21] Tile_X8Y14_LUT4AB/FrameData[22] Tile_X8Y14_LUT4AB/FrameData[23]
+ Tile_X8Y14_LUT4AB/FrameData[24] Tile_X8Y14_LUT4AB/FrameData[25] Tile_X8Y14_LUT4AB/FrameData[26]
+ Tile_X8Y14_LUT4AB/FrameData[27] Tile_X8Y14_LUT4AB/FrameData[28] Tile_X8Y14_LUT4AB/FrameData[29]
+ Tile_X8Y14_LUT4AB/FrameData[2] Tile_X8Y14_LUT4AB/FrameData[30] Tile_X8Y14_LUT4AB/FrameData[31]
+ Tile_X8Y14_LUT4AB/FrameData[3] Tile_X8Y14_LUT4AB/FrameData[4] Tile_X8Y14_LUT4AB/FrameData[5]
+ Tile_X8Y14_LUT4AB/FrameData[6] Tile_X8Y14_LUT4AB/FrameData[7] Tile_X8Y14_LUT4AB/FrameData[8]
+ Tile_X8Y14_LUT4AB/FrameData[9] Tile_X7Y15_S_term_DSP/FrameStrobe_O[0] Tile_X7Y15_S_term_DSP/FrameStrobe_O[10]
+ Tile_X7Y15_S_term_DSP/FrameStrobe_O[11] Tile_X7Y15_S_term_DSP/FrameStrobe_O[12]
+ Tile_X7Y15_S_term_DSP/FrameStrobe_O[13] Tile_X7Y15_S_term_DSP/FrameStrobe_O[14]
+ Tile_X7Y15_S_term_DSP/FrameStrobe_O[15] Tile_X7Y15_S_term_DSP/FrameStrobe_O[16]
+ Tile_X7Y15_S_term_DSP/FrameStrobe_O[17] Tile_X7Y15_S_term_DSP/FrameStrobe_O[18]
+ Tile_X7Y15_S_term_DSP/FrameStrobe_O[19] Tile_X7Y15_S_term_DSP/FrameStrobe_O[1] Tile_X7Y15_S_term_DSP/FrameStrobe_O[2]
+ Tile_X7Y15_S_term_DSP/FrameStrobe_O[3] Tile_X7Y15_S_term_DSP/FrameStrobe_O[4] Tile_X7Y15_S_term_DSP/FrameStrobe_O[5]
+ Tile_X7Y15_S_term_DSP/FrameStrobe_O[6] Tile_X7Y15_S_term_DSP/FrameStrobe_O[7] Tile_X7Y15_S_term_DSP/FrameStrobe_O[8]
+ Tile_X7Y15_S_term_DSP/FrameStrobe_O[9] Tile_X7Y15_S_term_DSP/N1BEG[0] Tile_X7Y15_S_term_DSP/N1BEG[1]
+ Tile_X7Y15_S_term_DSP/N1BEG[2] Tile_X7Y15_S_term_DSP/N1BEG[3] Tile_X7Y15_S_term_DSP/N2BEGb[0]
+ Tile_X7Y15_S_term_DSP/N2BEGb[1] Tile_X7Y15_S_term_DSP/N2BEGb[2] Tile_X7Y15_S_term_DSP/N2BEGb[3]
+ Tile_X7Y15_S_term_DSP/N2BEGb[4] Tile_X7Y15_S_term_DSP/N2BEGb[5] Tile_X7Y15_S_term_DSP/N2BEGb[6]
+ Tile_X7Y15_S_term_DSP/N2BEGb[7] Tile_X7Y15_S_term_DSP/N2BEG[0] Tile_X7Y15_S_term_DSP/N2BEG[1]
+ Tile_X7Y15_S_term_DSP/N2BEG[2] Tile_X7Y15_S_term_DSP/N2BEG[3] Tile_X7Y15_S_term_DSP/N2BEG[4]
+ Tile_X7Y15_S_term_DSP/N2BEG[5] Tile_X7Y15_S_term_DSP/N2BEG[6] Tile_X7Y15_S_term_DSP/N2BEG[7]
+ Tile_X7Y15_S_term_DSP/N4BEG[0] Tile_X7Y15_S_term_DSP/N4BEG[10] Tile_X7Y15_S_term_DSP/N4BEG[11]
+ Tile_X7Y15_S_term_DSP/N4BEG[12] Tile_X7Y15_S_term_DSP/N4BEG[13] Tile_X7Y15_S_term_DSP/N4BEG[14]
+ Tile_X7Y15_S_term_DSP/N4BEG[15] Tile_X7Y15_S_term_DSP/N4BEG[1] Tile_X7Y15_S_term_DSP/N4BEG[2]
+ Tile_X7Y15_S_term_DSP/N4BEG[3] Tile_X7Y15_S_term_DSP/N4BEG[4] Tile_X7Y15_S_term_DSP/N4BEG[5]
+ Tile_X7Y15_S_term_DSP/N4BEG[6] Tile_X7Y15_S_term_DSP/N4BEG[7] Tile_X7Y15_S_term_DSP/N4BEG[8]
+ Tile_X7Y15_S_term_DSP/N4BEG[9] Tile_X7Y15_S_term_DSP/NN4BEG[0] Tile_X7Y15_S_term_DSP/NN4BEG[10]
+ Tile_X7Y15_S_term_DSP/NN4BEG[11] Tile_X7Y15_S_term_DSP/NN4BEG[12] Tile_X7Y15_S_term_DSP/NN4BEG[13]
+ Tile_X7Y15_S_term_DSP/NN4BEG[14] Tile_X7Y15_S_term_DSP/NN4BEG[15] Tile_X7Y15_S_term_DSP/NN4BEG[1]
+ Tile_X7Y15_S_term_DSP/NN4BEG[2] Tile_X7Y15_S_term_DSP/NN4BEG[3] Tile_X7Y15_S_term_DSP/NN4BEG[4]
+ Tile_X7Y15_S_term_DSP/NN4BEG[5] Tile_X7Y15_S_term_DSP/NN4BEG[6] Tile_X7Y15_S_term_DSP/NN4BEG[7]
+ Tile_X7Y15_S_term_DSP/NN4BEG[8] Tile_X7Y15_S_term_DSP/NN4BEG[9] Tile_X7Y15_S_term_DSP/S1END[0]
+ Tile_X7Y15_S_term_DSP/S1END[1] Tile_X7Y15_S_term_DSP/S1END[2] Tile_X7Y15_S_term_DSP/S1END[3]
+ Tile_X7Y15_S_term_DSP/S2MID[0] Tile_X7Y15_S_term_DSP/S2MID[1] Tile_X7Y15_S_term_DSP/S2MID[2]
+ Tile_X7Y15_S_term_DSP/S2MID[3] Tile_X7Y15_S_term_DSP/S2MID[4] Tile_X7Y15_S_term_DSP/S2MID[5]
+ Tile_X7Y15_S_term_DSP/S2MID[6] Tile_X7Y15_S_term_DSP/S2MID[7] Tile_X7Y15_S_term_DSP/S2END[0]
+ Tile_X7Y15_S_term_DSP/S2END[1] Tile_X7Y15_S_term_DSP/S2END[2] Tile_X7Y15_S_term_DSP/S2END[3]
+ Tile_X7Y15_S_term_DSP/S2END[4] Tile_X7Y15_S_term_DSP/S2END[5] Tile_X7Y15_S_term_DSP/S2END[6]
+ Tile_X7Y15_S_term_DSP/S2END[7] Tile_X7Y15_S_term_DSP/S4END[0] Tile_X7Y15_S_term_DSP/S4END[10]
+ Tile_X7Y15_S_term_DSP/S4END[11] Tile_X7Y15_S_term_DSP/S4END[12] Tile_X7Y15_S_term_DSP/S4END[13]
+ Tile_X7Y15_S_term_DSP/S4END[14] Tile_X7Y15_S_term_DSP/S4END[15] Tile_X7Y15_S_term_DSP/S4END[1]
+ Tile_X7Y15_S_term_DSP/S4END[2] Tile_X7Y15_S_term_DSP/S4END[3] Tile_X7Y15_S_term_DSP/S4END[4]
+ Tile_X7Y15_S_term_DSP/S4END[5] Tile_X7Y15_S_term_DSP/S4END[6] Tile_X7Y15_S_term_DSP/S4END[7]
+ Tile_X7Y15_S_term_DSP/S4END[8] Tile_X7Y15_S_term_DSP/S4END[9] Tile_X7Y15_S_term_DSP/SS4END[0]
+ Tile_X7Y15_S_term_DSP/SS4END[10] Tile_X7Y15_S_term_DSP/SS4END[11] Tile_X7Y15_S_term_DSP/SS4END[12]
+ Tile_X7Y15_S_term_DSP/SS4END[13] Tile_X7Y15_S_term_DSP/SS4END[14] Tile_X7Y15_S_term_DSP/SS4END[15]
+ Tile_X7Y15_S_term_DSP/SS4END[1] Tile_X7Y15_S_term_DSP/SS4END[2] Tile_X7Y15_S_term_DSP/SS4END[3]
+ Tile_X7Y15_S_term_DSP/SS4END[4] Tile_X7Y15_S_term_DSP/SS4END[5] Tile_X7Y15_S_term_DSP/SS4END[6]
+ Tile_X7Y15_S_term_DSP/SS4END[7] Tile_X7Y15_S_term_DSP/SS4END[8] Tile_X7Y15_S_term_DSP/SS4END[9]
+ Tile_X7Y15_S_term_DSP/UserCLKo Tile_X6Y14_LUT4AB/W1END[0] Tile_X6Y14_LUT4AB/W1END[1]
+ Tile_X6Y14_LUT4AB/W1END[2] Tile_X6Y14_LUT4AB/W1END[3] Tile_X8Y14_LUT4AB/W1BEG[0]
+ Tile_X8Y14_LUT4AB/W1BEG[1] Tile_X8Y14_LUT4AB/W1BEG[2] Tile_X8Y14_LUT4AB/W1BEG[3]
+ Tile_X6Y14_LUT4AB/W2MID[0] Tile_X6Y14_LUT4AB/W2MID[1] Tile_X6Y14_LUT4AB/W2MID[2]
+ Tile_X6Y14_LUT4AB/W2MID[3] Tile_X6Y14_LUT4AB/W2MID[4] Tile_X6Y14_LUT4AB/W2MID[5]
+ Tile_X6Y14_LUT4AB/W2MID[6] Tile_X6Y14_LUT4AB/W2MID[7] Tile_X6Y14_LUT4AB/W2END[0]
+ Tile_X6Y14_LUT4AB/W2END[1] Tile_X6Y14_LUT4AB/W2END[2] Tile_X6Y14_LUT4AB/W2END[3]
+ Tile_X6Y14_LUT4AB/W2END[4] Tile_X6Y14_LUT4AB/W2END[5] Tile_X6Y14_LUT4AB/W2END[6]
+ Tile_X6Y14_LUT4AB/W2END[7] Tile_X8Y14_LUT4AB/W2BEGb[0] Tile_X8Y14_LUT4AB/W2BEGb[1]
+ Tile_X8Y14_LUT4AB/W2BEGb[2] Tile_X8Y14_LUT4AB/W2BEGb[3] Tile_X8Y14_LUT4AB/W2BEGb[4]
+ Tile_X8Y14_LUT4AB/W2BEGb[5] Tile_X8Y14_LUT4AB/W2BEGb[6] Tile_X8Y14_LUT4AB/W2BEGb[7]
+ Tile_X8Y14_LUT4AB/W2BEG[0] Tile_X8Y14_LUT4AB/W2BEG[1] Tile_X8Y14_LUT4AB/W2BEG[2]
+ Tile_X8Y14_LUT4AB/W2BEG[3] Tile_X8Y14_LUT4AB/W2BEG[4] Tile_X8Y14_LUT4AB/W2BEG[5]
+ Tile_X8Y14_LUT4AB/W2BEG[6] Tile_X8Y14_LUT4AB/W2BEG[7] Tile_X6Y14_LUT4AB/W6END[0]
+ Tile_X6Y14_LUT4AB/W6END[10] Tile_X6Y14_LUT4AB/W6END[11] Tile_X6Y14_LUT4AB/W6END[1]
+ Tile_X6Y14_LUT4AB/W6END[2] Tile_X6Y14_LUT4AB/W6END[3] Tile_X6Y14_LUT4AB/W6END[4]
+ Tile_X6Y14_LUT4AB/W6END[5] Tile_X6Y14_LUT4AB/W6END[6] Tile_X6Y14_LUT4AB/W6END[7]
+ Tile_X6Y14_LUT4AB/W6END[8] Tile_X6Y14_LUT4AB/W6END[9] Tile_X8Y14_LUT4AB/W6BEG[0]
+ Tile_X8Y14_LUT4AB/W6BEG[10] Tile_X8Y14_LUT4AB/W6BEG[11] Tile_X8Y14_LUT4AB/W6BEG[1]
+ Tile_X8Y14_LUT4AB/W6BEG[2] Tile_X8Y14_LUT4AB/W6BEG[3] Tile_X8Y14_LUT4AB/W6BEG[4]
+ Tile_X8Y14_LUT4AB/W6BEG[5] Tile_X8Y14_LUT4AB/W6BEG[6] Tile_X8Y14_LUT4AB/W6BEG[7]
+ Tile_X8Y14_LUT4AB/W6BEG[8] Tile_X8Y14_LUT4AB/W6BEG[9] Tile_X6Y14_LUT4AB/WW4END[0]
+ Tile_X6Y14_LUT4AB/WW4END[10] Tile_X6Y14_LUT4AB/WW4END[11] Tile_X6Y14_LUT4AB/WW4END[12]
+ Tile_X6Y14_LUT4AB/WW4END[13] Tile_X6Y14_LUT4AB/WW4END[14] Tile_X6Y14_LUT4AB/WW4END[15]
+ Tile_X6Y14_LUT4AB/WW4END[1] Tile_X6Y14_LUT4AB/WW4END[2] Tile_X6Y14_LUT4AB/WW4END[3]
+ Tile_X6Y14_LUT4AB/WW4END[4] Tile_X6Y14_LUT4AB/WW4END[5] Tile_X6Y14_LUT4AB/WW4END[6]
+ Tile_X6Y14_LUT4AB/WW4END[7] Tile_X6Y14_LUT4AB/WW4END[8] Tile_X6Y14_LUT4AB/WW4END[9]
+ Tile_X8Y14_LUT4AB/WW4BEG[0] Tile_X8Y14_LUT4AB/WW4BEG[10] Tile_X8Y14_LUT4AB/WW4BEG[11]
+ Tile_X8Y14_LUT4AB/WW4BEG[12] Tile_X8Y14_LUT4AB/WW4BEG[13] Tile_X8Y14_LUT4AB/WW4BEG[14]
+ Tile_X8Y14_LUT4AB/WW4BEG[15] Tile_X8Y14_LUT4AB/WW4BEG[1] Tile_X8Y14_LUT4AB/WW4BEG[2]
+ Tile_X8Y14_LUT4AB/WW4BEG[3] Tile_X8Y14_LUT4AB/WW4BEG[4] Tile_X8Y14_LUT4AB/WW4BEG[5]
+ Tile_X8Y14_LUT4AB/WW4BEG[6] Tile_X8Y14_LUT4AB/WW4BEG[7] Tile_X8Y14_LUT4AB/WW4BEG[8]
+ Tile_X8Y14_LUT4AB/WW4BEG[9] VGND VPWR DSP
XTile_X4Y9_RegFile Tile_X5Y9_LUT4AB/E1END[0] Tile_X5Y9_LUT4AB/E1END[1] Tile_X5Y9_LUT4AB/E1END[2]
+ Tile_X5Y9_LUT4AB/E1END[3] Tile_X3Y9_LUT4AB/E1BEG[0] Tile_X3Y9_LUT4AB/E1BEG[1] Tile_X3Y9_LUT4AB/E1BEG[2]
+ Tile_X3Y9_LUT4AB/E1BEG[3] Tile_X5Y9_LUT4AB/E2MID[0] Tile_X5Y9_LUT4AB/E2MID[1] Tile_X5Y9_LUT4AB/E2MID[2]
+ Tile_X5Y9_LUT4AB/E2MID[3] Tile_X5Y9_LUT4AB/E2MID[4] Tile_X5Y9_LUT4AB/E2MID[5] Tile_X5Y9_LUT4AB/E2MID[6]
+ Tile_X5Y9_LUT4AB/E2MID[7] Tile_X5Y9_LUT4AB/E2END[0] Tile_X5Y9_LUT4AB/E2END[1] Tile_X5Y9_LUT4AB/E2END[2]
+ Tile_X5Y9_LUT4AB/E2END[3] Tile_X5Y9_LUT4AB/E2END[4] Tile_X5Y9_LUT4AB/E2END[5] Tile_X5Y9_LUT4AB/E2END[6]
+ Tile_X5Y9_LUT4AB/E2END[7] Tile_X4Y9_RegFile/E2END[0] Tile_X4Y9_RegFile/E2END[1]
+ Tile_X4Y9_RegFile/E2END[2] Tile_X4Y9_RegFile/E2END[3] Tile_X4Y9_RegFile/E2END[4]
+ Tile_X4Y9_RegFile/E2END[5] Tile_X4Y9_RegFile/E2END[6] Tile_X4Y9_RegFile/E2END[7]
+ Tile_X3Y9_LUT4AB/E2BEG[0] Tile_X3Y9_LUT4AB/E2BEG[1] Tile_X3Y9_LUT4AB/E2BEG[2] Tile_X3Y9_LUT4AB/E2BEG[3]
+ Tile_X3Y9_LUT4AB/E2BEG[4] Tile_X3Y9_LUT4AB/E2BEG[5] Tile_X3Y9_LUT4AB/E2BEG[6] Tile_X3Y9_LUT4AB/E2BEG[7]
+ Tile_X5Y9_LUT4AB/E6END[0] Tile_X5Y9_LUT4AB/E6END[10] Tile_X5Y9_LUT4AB/E6END[11]
+ Tile_X5Y9_LUT4AB/E6END[1] Tile_X5Y9_LUT4AB/E6END[2] Tile_X5Y9_LUT4AB/E6END[3] Tile_X5Y9_LUT4AB/E6END[4]
+ Tile_X5Y9_LUT4AB/E6END[5] Tile_X5Y9_LUT4AB/E6END[6] Tile_X5Y9_LUT4AB/E6END[7] Tile_X5Y9_LUT4AB/E6END[8]
+ Tile_X5Y9_LUT4AB/E6END[9] Tile_X3Y9_LUT4AB/E6BEG[0] Tile_X3Y9_LUT4AB/E6BEG[10] Tile_X3Y9_LUT4AB/E6BEG[11]
+ Tile_X3Y9_LUT4AB/E6BEG[1] Tile_X3Y9_LUT4AB/E6BEG[2] Tile_X3Y9_LUT4AB/E6BEG[3] Tile_X3Y9_LUT4AB/E6BEG[4]
+ Tile_X3Y9_LUT4AB/E6BEG[5] Tile_X3Y9_LUT4AB/E6BEG[6] Tile_X3Y9_LUT4AB/E6BEG[7] Tile_X3Y9_LUT4AB/E6BEG[8]
+ Tile_X3Y9_LUT4AB/E6BEG[9] Tile_X5Y9_LUT4AB/EE4END[0] Tile_X5Y9_LUT4AB/EE4END[10]
+ Tile_X5Y9_LUT4AB/EE4END[11] Tile_X5Y9_LUT4AB/EE4END[12] Tile_X5Y9_LUT4AB/EE4END[13]
+ Tile_X5Y9_LUT4AB/EE4END[14] Tile_X5Y9_LUT4AB/EE4END[15] Tile_X5Y9_LUT4AB/EE4END[1]
+ Tile_X5Y9_LUT4AB/EE4END[2] Tile_X5Y9_LUT4AB/EE4END[3] Tile_X5Y9_LUT4AB/EE4END[4]
+ Tile_X5Y9_LUT4AB/EE4END[5] Tile_X5Y9_LUT4AB/EE4END[6] Tile_X5Y9_LUT4AB/EE4END[7]
+ Tile_X5Y9_LUT4AB/EE4END[8] Tile_X5Y9_LUT4AB/EE4END[9] Tile_X3Y9_LUT4AB/EE4BEG[0]
+ Tile_X3Y9_LUT4AB/EE4BEG[10] Tile_X3Y9_LUT4AB/EE4BEG[11] Tile_X3Y9_LUT4AB/EE4BEG[12]
+ Tile_X3Y9_LUT4AB/EE4BEG[13] Tile_X3Y9_LUT4AB/EE4BEG[14] Tile_X3Y9_LUT4AB/EE4BEG[15]
+ Tile_X3Y9_LUT4AB/EE4BEG[1] Tile_X3Y9_LUT4AB/EE4BEG[2] Tile_X3Y9_LUT4AB/EE4BEG[3]
+ Tile_X3Y9_LUT4AB/EE4BEG[4] Tile_X3Y9_LUT4AB/EE4BEG[5] Tile_X3Y9_LUT4AB/EE4BEG[6]
+ Tile_X3Y9_LUT4AB/EE4BEG[7] Tile_X3Y9_LUT4AB/EE4BEG[8] Tile_X3Y9_LUT4AB/EE4BEG[9]
+ Tile_X4Y9_RegFile/FrameData[0] Tile_X4Y9_RegFile/FrameData[10] Tile_X4Y9_RegFile/FrameData[11]
+ Tile_X4Y9_RegFile/FrameData[12] Tile_X4Y9_RegFile/FrameData[13] Tile_X4Y9_RegFile/FrameData[14]
+ Tile_X4Y9_RegFile/FrameData[15] Tile_X4Y9_RegFile/FrameData[16] Tile_X4Y9_RegFile/FrameData[17]
+ Tile_X4Y9_RegFile/FrameData[18] Tile_X4Y9_RegFile/FrameData[19] Tile_X4Y9_RegFile/FrameData[1]
+ Tile_X4Y9_RegFile/FrameData[20] Tile_X4Y9_RegFile/FrameData[21] Tile_X4Y9_RegFile/FrameData[22]
+ Tile_X4Y9_RegFile/FrameData[23] Tile_X4Y9_RegFile/FrameData[24] Tile_X4Y9_RegFile/FrameData[25]
+ Tile_X4Y9_RegFile/FrameData[26] Tile_X4Y9_RegFile/FrameData[27] Tile_X4Y9_RegFile/FrameData[28]
+ Tile_X4Y9_RegFile/FrameData[29] Tile_X4Y9_RegFile/FrameData[2] Tile_X4Y9_RegFile/FrameData[30]
+ Tile_X4Y9_RegFile/FrameData[31] Tile_X4Y9_RegFile/FrameData[3] Tile_X4Y9_RegFile/FrameData[4]
+ Tile_X4Y9_RegFile/FrameData[5] Tile_X4Y9_RegFile/FrameData[6] Tile_X4Y9_RegFile/FrameData[7]
+ Tile_X4Y9_RegFile/FrameData[8] Tile_X4Y9_RegFile/FrameData[9] Tile_X5Y9_LUT4AB/FrameData[0]
+ Tile_X5Y9_LUT4AB/FrameData[10] Tile_X5Y9_LUT4AB/FrameData[11] Tile_X5Y9_LUT4AB/FrameData[12]
+ Tile_X5Y9_LUT4AB/FrameData[13] Tile_X5Y9_LUT4AB/FrameData[14] Tile_X5Y9_LUT4AB/FrameData[15]
+ Tile_X5Y9_LUT4AB/FrameData[16] Tile_X5Y9_LUT4AB/FrameData[17] Tile_X5Y9_LUT4AB/FrameData[18]
+ Tile_X5Y9_LUT4AB/FrameData[19] Tile_X5Y9_LUT4AB/FrameData[1] Tile_X5Y9_LUT4AB/FrameData[20]
+ Tile_X5Y9_LUT4AB/FrameData[21] Tile_X5Y9_LUT4AB/FrameData[22] Tile_X5Y9_LUT4AB/FrameData[23]
+ Tile_X5Y9_LUT4AB/FrameData[24] Tile_X5Y9_LUT4AB/FrameData[25] Tile_X5Y9_LUT4AB/FrameData[26]
+ Tile_X5Y9_LUT4AB/FrameData[27] Tile_X5Y9_LUT4AB/FrameData[28] Tile_X5Y9_LUT4AB/FrameData[29]
+ Tile_X5Y9_LUT4AB/FrameData[2] Tile_X5Y9_LUT4AB/FrameData[30] Tile_X5Y9_LUT4AB/FrameData[31]
+ Tile_X5Y9_LUT4AB/FrameData[3] Tile_X5Y9_LUT4AB/FrameData[4] Tile_X5Y9_LUT4AB/FrameData[5]
+ Tile_X5Y9_LUT4AB/FrameData[6] Tile_X5Y9_LUT4AB/FrameData[7] Tile_X5Y9_LUT4AB/FrameData[8]
+ Tile_X5Y9_LUT4AB/FrameData[9] Tile_X4Y9_RegFile/FrameStrobe[0] Tile_X4Y9_RegFile/FrameStrobe[10]
+ Tile_X4Y9_RegFile/FrameStrobe[11] Tile_X4Y9_RegFile/FrameStrobe[12] Tile_X4Y9_RegFile/FrameStrobe[13]
+ Tile_X4Y9_RegFile/FrameStrobe[14] Tile_X4Y9_RegFile/FrameStrobe[15] Tile_X4Y9_RegFile/FrameStrobe[16]
+ Tile_X4Y9_RegFile/FrameStrobe[17] Tile_X4Y9_RegFile/FrameStrobe[18] Tile_X4Y9_RegFile/FrameStrobe[19]
+ Tile_X4Y9_RegFile/FrameStrobe[1] Tile_X4Y9_RegFile/FrameStrobe[2] Tile_X4Y9_RegFile/FrameStrobe[3]
+ Tile_X4Y9_RegFile/FrameStrobe[4] Tile_X4Y9_RegFile/FrameStrobe[5] Tile_X4Y9_RegFile/FrameStrobe[6]
+ Tile_X4Y9_RegFile/FrameStrobe[7] Tile_X4Y9_RegFile/FrameStrobe[8] Tile_X4Y9_RegFile/FrameStrobe[9]
+ Tile_X4Y8_RegFile/FrameStrobe[0] Tile_X4Y8_RegFile/FrameStrobe[10] Tile_X4Y8_RegFile/FrameStrobe[11]
+ Tile_X4Y8_RegFile/FrameStrobe[12] Tile_X4Y8_RegFile/FrameStrobe[13] Tile_X4Y8_RegFile/FrameStrobe[14]
+ Tile_X4Y8_RegFile/FrameStrobe[15] Tile_X4Y8_RegFile/FrameStrobe[16] Tile_X4Y8_RegFile/FrameStrobe[17]
+ Tile_X4Y8_RegFile/FrameStrobe[18] Tile_X4Y8_RegFile/FrameStrobe[19] Tile_X4Y8_RegFile/FrameStrobe[1]
+ Tile_X4Y8_RegFile/FrameStrobe[2] Tile_X4Y8_RegFile/FrameStrobe[3] Tile_X4Y8_RegFile/FrameStrobe[4]
+ Tile_X4Y8_RegFile/FrameStrobe[5] Tile_X4Y8_RegFile/FrameStrobe[6] Tile_X4Y8_RegFile/FrameStrobe[7]
+ Tile_X4Y8_RegFile/FrameStrobe[8] Tile_X4Y8_RegFile/FrameStrobe[9] Tile_X4Y9_RegFile/N1BEG[0]
+ Tile_X4Y9_RegFile/N1BEG[1] Tile_X4Y9_RegFile/N1BEG[2] Tile_X4Y9_RegFile/N1BEG[3]
+ Tile_X4Y9_RegFile/N1END[0] Tile_X4Y9_RegFile/N1END[1] Tile_X4Y9_RegFile/N1END[2]
+ Tile_X4Y9_RegFile/N1END[3] Tile_X4Y9_RegFile/N2BEG[0] Tile_X4Y9_RegFile/N2BEG[1]
+ Tile_X4Y9_RegFile/N2BEG[2] Tile_X4Y9_RegFile/N2BEG[3] Tile_X4Y9_RegFile/N2BEG[4]
+ Tile_X4Y9_RegFile/N2BEG[5] Tile_X4Y9_RegFile/N2BEG[6] Tile_X4Y9_RegFile/N2BEG[7]
+ Tile_X4Y8_RegFile/N2END[0] Tile_X4Y8_RegFile/N2END[1] Tile_X4Y8_RegFile/N2END[2]
+ Tile_X4Y8_RegFile/N2END[3] Tile_X4Y8_RegFile/N2END[4] Tile_X4Y8_RegFile/N2END[5]
+ Tile_X4Y8_RegFile/N2END[6] Tile_X4Y8_RegFile/N2END[7] Tile_X4Y9_RegFile/N2END[0]
+ Tile_X4Y9_RegFile/N2END[1] Tile_X4Y9_RegFile/N2END[2] Tile_X4Y9_RegFile/N2END[3]
+ Tile_X4Y9_RegFile/N2END[4] Tile_X4Y9_RegFile/N2END[5] Tile_X4Y9_RegFile/N2END[6]
+ Tile_X4Y9_RegFile/N2END[7] Tile_X4Y9_RegFile/N2MID[0] Tile_X4Y9_RegFile/N2MID[1]
+ Tile_X4Y9_RegFile/N2MID[2] Tile_X4Y9_RegFile/N2MID[3] Tile_X4Y9_RegFile/N2MID[4]
+ Tile_X4Y9_RegFile/N2MID[5] Tile_X4Y9_RegFile/N2MID[6] Tile_X4Y9_RegFile/N2MID[7]
+ Tile_X4Y9_RegFile/N4BEG[0] Tile_X4Y9_RegFile/N4BEG[10] Tile_X4Y9_RegFile/N4BEG[11]
+ Tile_X4Y9_RegFile/N4BEG[12] Tile_X4Y9_RegFile/N4BEG[13] Tile_X4Y9_RegFile/N4BEG[14]
+ Tile_X4Y9_RegFile/N4BEG[15] Tile_X4Y9_RegFile/N4BEG[1] Tile_X4Y9_RegFile/N4BEG[2]
+ Tile_X4Y9_RegFile/N4BEG[3] Tile_X4Y9_RegFile/N4BEG[4] Tile_X4Y9_RegFile/N4BEG[5]
+ Tile_X4Y9_RegFile/N4BEG[6] Tile_X4Y9_RegFile/N4BEG[7] Tile_X4Y9_RegFile/N4BEG[8]
+ Tile_X4Y9_RegFile/N4BEG[9] Tile_X4Y9_RegFile/N4END[0] Tile_X4Y9_RegFile/N4END[10]
+ Tile_X4Y9_RegFile/N4END[11] Tile_X4Y9_RegFile/N4END[12] Tile_X4Y9_RegFile/N4END[13]
+ Tile_X4Y9_RegFile/N4END[14] Tile_X4Y9_RegFile/N4END[15] Tile_X4Y9_RegFile/N4END[1]
+ Tile_X4Y9_RegFile/N4END[2] Tile_X4Y9_RegFile/N4END[3] Tile_X4Y9_RegFile/N4END[4]
+ Tile_X4Y9_RegFile/N4END[5] Tile_X4Y9_RegFile/N4END[6] Tile_X4Y9_RegFile/N4END[7]
+ Tile_X4Y9_RegFile/N4END[8] Tile_X4Y9_RegFile/N4END[9] Tile_X4Y9_RegFile/NN4BEG[0]
+ Tile_X4Y9_RegFile/NN4BEG[10] Tile_X4Y9_RegFile/NN4BEG[11] Tile_X4Y9_RegFile/NN4BEG[12]
+ Tile_X4Y9_RegFile/NN4BEG[13] Tile_X4Y9_RegFile/NN4BEG[14] Tile_X4Y9_RegFile/NN4BEG[15]
+ Tile_X4Y9_RegFile/NN4BEG[1] Tile_X4Y9_RegFile/NN4BEG[2] Tile_X4Y9_RegFile/NN4BEG[3]
+ Tile_X4Y9_RegFile/NN4BEG[4] Tile_X4Y9_RegFile/NN4BEG[5] Tile_X4Y9_RegFile/NN4BEG[6]
+ Tile_X4Y9_RegFile/NN4BEG[7] Tile_X4Y9_RegFile/NN4BEG[8] Tile_X4Y9_RegFile/NN4BEG[9]
+ Tile_X4Y9_RegFile/NN4END[0] Tile_X4Y9_RegFile/NN4END[10] Tile_X4Y9_RegFile/NN4END[11]
+ Tile_X4Y9_RegFile/NN4END[12] Tile_X4Y9_RegFile/NN4END[13] Tile_X4Y9_RegFile/NN4END[14]
+ Tile_X4Y9_RegFile/NN4END[15] Tile_X4Y9_RegFile/NN4END[1] Tile_X4Y9_RegFile/NN4END[2]
+ Tile_X4Y9_RegFile/NN4END[3] Tile_X4Y9_RegFile/NN4END[4] Tile_X4Y9_RegFile/NN4END[5]
+ Tile_X4Y9_RegFile/NN4END[6] Tile_X4Y9_RegFile/NN4END[7] Tile_X4Y9_RegFile/NN4END[8]
+ Tile_X4Y9_RegFile/NN4END[9] Tile_X4Y9_RegFile/S1BEG[0] Tile_X4Y9_RegFile/S1BEG[1]
+ Tile_X4Y9_RegFile/S1BEG[2] Tile_X4Y9_RegFile/S1BEG[3] Tile_X4Y9_RegFile/S1END[0]
+ Tile_X4Y9_RegFile/S1END[1] Tile_X4Y9_RegFile/S1END[2] Tile_X4Y9_RegFile/S1END[3]
+ Tile_X4Y9_RegFile/S2BEG[0] Tile_X4Y9_RegFile/S2BEG[1] Tile_X4Y9_RegFile/S2BEG[2]
+ Tile_X4Y9_RegFile/S2BEG[3] Tile_X4Y9_RegFile/S2BEG[4] Tile_X4Y9_RegFile/S2BEG[5]
+ Tile_X4Y9_RegFile/S2BEG[6] Tile_X4Y9_RegFile/S2BEG[7] Tile_X4Y9_RegFile/S2BEGb[0]
+ Tile_X4Y9_RegFile/S2BEGb[1] Tile_X4Y9_RegFile/S2BEGb[2] Tile_X4Y9_RegFile/S2BEGb[3]
+ Tile_X4Y9_RegFile/S2BEGb[4] Tile_X4Y9_RegFile/S2BEGb[5] Tile_X4Y9_RegFile/S2BEGb[6]
+ Tile_X4Y9_RegFile/S2BEGb[7] Tile_X4Y9_RegFile/S2END[0] Tile_X4Y9_RegFile/S2END[1]
+ Tile_X4Y9_RegFile/S2END[2] Tile_X4Y9_RegFile/S2END[3] Tile_X4Y9_RegFile/S2END[4]
+ Tile_X4Y9_RegFile/S2END[5] Tile_X4Y9_RegFile/S2END[6] Tile_X4Y9_RegFile/S2END[7]
+ Tile_X4Y9_RegFile/S2MID[0] Tile_X4Y9_RegFile/S2MID[1] Tile_X4Y9_RegFile/S2MID[2]
+ Tile_X4Y9_RegFile/S2MID[3] Tile_X4Y9_RegFile/S2MID[4] Tile_X4Y9_RegFile/S2MID[5]
+ Tile_X4Y9_RegFile/S2MID[6] Tile_X4Y9_RegFile/S2MID[7] Tile_X4Y9_RegFile/S4BEG[0]
+ Tile_X4Y9_RegFile/S4BEG[10] Tile_X4Y9_RegFile/S4BEG[11] Tile_X4Y9_RegFile/S4BEG[12]
+ Tile_X4Y9_RegFile/S4BEG[13] Tile_X4Y9_RegFile/S4BEG[14] Tile_X4Y9_RegFile/S4BEG[15]
+ Tile_X4Y9_RegFile/S4BEG[1] Tile_X4Y9_RegFile/S4BEG[2] Tile_X4Y9_RegFile/S4BEG[3]
+ Tile_X4Y9_RegFile/S4BEG[4] Tile_X4Y9_RegFile/S4BEG[5] Tile_X4Y9_RegFile/S4BEG[6]
+ Tile_X4Y9_RegFile/S4BEG[7] Tile_X4Y9_RegFile/S4BEG[8] Tile_X4Y9_RegFile/S4BEG[9]
+ Tile_X4Y9_RegFile/S4END[0] Tile_X4Y9_RegFile/S4END[10] Tile_X4Y9_RegFile/S4END[11]
+ Tile_X4Y9_RegFile/S4END[12] Tile_X4Y9_RegFile/S4END[13] Tile_X4Y9_RegFile/S4END[14]
+ Tile_X4Y9_RegFile/S4END[15] Tile_X4Y9_RegFile/S4END[1] Tile_X4Y9_RegFile/S4END[2]
+ Tile_X4Y9_RegFile/S4END[3] Tile_X4Y9_RegFile/S4END[4] Tile_X4Y9_RegFile/S4END[5]
+ Tile_X4Y9_RegFile/S4END[6] Tile_X4Y9_RegFile/S4END[7] Tile_X4Y9_RegFile/S4END[8]
+ Tile_X4Y9_RegFile/S4END[9] Tile_X4Y9_RegFile/SS4BEG[0] Tile_X4Y9_RegFile/SS4BEG[10]
+ Tile_X4Y9_RegFile/SS4BEG[11] Tile_X4Y9_RegFile/SS4BEG[12] Tile_X4Y9_RegFile/SS4BEG[13]
+ Tile_X4Y9_RegFile/SS4BEG[14] Tile_X4Y9_RegFile/SS4BEG[15] Tile_X4Y9_RegFile/SS4BEG[1]
+ Tile_X4Y9_RegFile/SS4BEG[2] Tile_X4Y9_RegFile/SS4BEG[3] Tile_X4Y9_RegFile/SS4BEG[4]
+ Tile_X4Y9_RegFile/SS4BEG[5] Tile_X4Y9_RegFile/SS4BEG[6] Tile_X4Y9_RegFile/SS4BEG[7]
+ Tile_X4Y9_RegFile/SS4BEG[8] Tile_X4Y9_RegFile/SS4BEG[9] Tile_X4Y9_RegFile/SS4END[0]
+ Tile_X4Y9_RegFile/SS4END[10] Tile_X4Y9_RegFile/SS4END[11] Tile_X4Y9_RegFile/SS4END[12]
+ Tile_X4Y9_RegFile/SS4END[13] Tile_X4Y9_RegFile/SS4END[14] Tile_X4Y9_RegFile/SS4END[15]
+ Tile_X4Y9_RegFile/SS4END[1] Tile_X4Y9_RegFile/SS4END[2] Tile_X4Y9_RegFile/SS4END[3]
+ Tile_X4Y9_RegFile/SS4END[4] Tile_X4Y9_RegFile/SS4END[5] Tile_X4Y9_RegFile/SS4END[6]
+ Tile_X4Y9_RegFile/SS4END[7] Tile_X4Y9_RegFile/SS4END[8] Tile_X4Y9_RegFile/SS4END[9]
+ Tile_X4Y9_RegFile/UserCLK Tile_X4Y8_RegFile/UserCLK VGND VPWR Tile_X3Y9_LUT4AB/W1END[0]
+ Tile_X3Y9_LUT4AB/W1END[1] Tile_X3Y9_LUT4AB/W1END[2] Tile_X3Y9_LUT4AB/W1END[3] Tile_X5Y9_LUT4AB/W1BEG[0]
+ Tile_X5Y9_LUT4AB/W1BEG[1] Tile_X5Y9_LUT4AB/W1BEG[2] Tile_X5Y9_LUT4AB/W1BEG[3] Tile_X3Y9_LUT4AB/W2MID[0]
+ Tile_X3Y9_LUT4AB/W2MID[1] Tile_X3Y9_LUT4AB/W2MID[2] Tile_X3Y9_LUT4AB/W2MID[3] Tile_X3Y9_LUT4AB/W2MID[4]
+ Tile_X3Y9_LUT4AB/W2MID[5] Tile_X3Y9_LUT4AB/W2MID[6] Tile_X3Y9_LUT4AB/W2MID[7] Tile_X3Y9_LUT4AB/W2END[0]
+ Tile_X3Y9_LUT4AB/W2END[1] Tile_X3Y9_LUT4AB/W2END[2] Tile_X3Y9_LUT4AB/W2END[3] Tile_X3Y9_LUT4AB/W2END[4]
+ Tile_X3Y9_LUT4AB/W2END[5] Tile_X3Y9_LUT4AB/W2END[6] Tile_X3Y9_LUT4AB/W2END[7] Tile_X5Y9_LUT4AB/W2BEGb[0]
+ Tile_X5Y9_LUT4AB/W2BEGb[1] Tile_X5Y9_LUT4AB/W2BEGb[2] Tile_X5Y9_LUT4AB/W2BEGb[3]
+ Tile_X5Y9_LUT4AB/W2BEGb[4] Tile_X5Y9_LUT4AB/W2BEGb[5] Tile_X5Y9_LUT4AB/W2BEGb[6]
+ Tile_X5Y9_LUT4AB/W2BEGb[7] Tile_X5Y9_LUT4AB/W2BEG[0] Tile_X5Y9_LUT4AB/W2BEG[1] Tile_X5Y9_LUT4AB/W2BEG[2]
+ Tile_X5Y9_LUT4AB/W2BEG[3] Tile_X5Y9_LUT4AB/W2BEG[4] Tile_X5Y9_LUT4AB/W2BEG[5] Tile_X5Y9_LUT4AB/W2BEG[6]
+ Tile_X5Y9_LUT4AB/W2BEG[7] Tile_X3Y9_LUT4AB/W6END[0] Tile_X3Y9_LUT4AB/W6END[10] Tile_X3Y9_LUT4AB/W6END[11]
+ Tile_X3Y9_LUT4AB/W6END[1] Tile_X3Y9_LUT4AB/W6END[2] Tile_X3Y9_LUT4AB/W6END[3] Tile_X3Y9_LUT4AB/W6END[4]
+ Tile_X3Y9_LUT4AB/W6END[5] Tile_X3Y9_LUT4AB/W6END[6] Tile_X3Y9_LUT4AB/W6END[7] Tile_X3Y9_LUT4AB/W6END[8]
+ Tile_X3Y9_LUT4AB/W6END[9] Tile_X5Y9_LUT4AB/W6BEG[0] Tile_X5Y9_LUT4AB/W6BEG[10] Tile_X5Y9_LUT4AB/W6BEG[11]
+ Tile_X5Y9_LUT4AB/W6BEG[1] Tile_X5Y9_LUT4AB/W6BEG[2] Tile_X5Y9_LUT4AB/W6BEG[3] Tile_X5Y9_LUT4AB/W6BEG[4]
+ Tile_X5Y9_LUT4AB/W6BEG[5] Tile_X5Y9_LUT4AB/W6BEG[6] Tile_X5Y9_LUT4AB/W6BEG[7] Tile_X5Y9_LUT4AB/W6BEG[8]
+ Tile_X5Y9_LUT4AB/W6BEG[9] Tile_X3Y9_LUT4AB/WW4END[0] Tile_X3Y9_LUT4AB/WW4END[10]
+ Tile_X3Y9_LUT4AB/WW4END[11] Tile_X3Y9_LUT4AB/WW4END[12] Tile_X3Y9_LUT4AB/WW4END[13]
+ Tile_X3Y9_LUT4AB/WW4END[14] Tile_X3Y9_LUT4AB/WW4END[15] Tile_X3Y9_LUT4AB/WW4END[1]
+ Tile_X3Y9_LUT4AB/WW4END[2] Tile_X3Y9_LUT4AB/WW4END[3] Tile_X3Y9_LUT4AB/WW4END[4]
+ Tile_X3Y9_LUT4AB/WW4END[5] Tile_X3Y9_LUT4AB/WW4END[6] Tile_X3Y9_LUT4AB/WW4END[7]
+ Tile_X3Y9_LUT4AB/WW4END[8] Tile_X3Y9_LUT4AB/WW4END[9] Tile_X5Y9_LUT4AB/WW4BEG[0]
+ Tile_X5Y9_LUT4AB/WW4BEG[10] Tile_X5Y9_LUT4AB/WW4BEG[11] Tile_X5Y9_LUT4AB/WW4BEG[12]
+ Tile_X5Y9_LUT4AB/WW4BEG[13] Tile_X5Y9_LUT4AB/WW4BEG[14] Tile_X5Y9_LUT4AB/WW4BEG[15]
+ Tile_X5Y9_LUT4AB/WW4BEG[1] Tile_X5Y9_LUT4AB/WW4BEG[2] Tile_X5Y9_LUT4AB/WW4BEG[3]
+ Tile_X5Y9_LUT4AB/WW4BEG[4] Tile_X5Y9_LUT4AB/WW4BEG[5] Tile_X5Y9_LUT4AB/WW4BEG[6]
+ Tile_X5Y9_LUT4AB/WW4BEG[7] Tile_X5Y9_LUT4AB/WW4BEG[8] Tile_X5Y9_LUT4AB/WW4BEG[9]
+ RegFile
XTile_X5Y10_LUT4AB Tile_X5Y11_LUT4AB/Co Tile_X5Y9_LUT4AB/Ci Tile_X6Y10_LUT4AB/E1END[0]
+ Tile_X6Y10_LUT4AB/E1END[1] Tile_X6Y10_LUT4AB/E1END[2] Tile_X6Y10_LUT4AB/E1END[3]
+ Tile_X5Y10_LUT4AB/E1END[0] Tile_X5Y10_LUT4AB/E1END[1] Tile_X5Y10_LUT4AB/E1END[2]
+ Tile_X5Y10_LUT4AB/E1END[3] Tile_X6Y10_LUT4AB/E2MID[0] Tile_X6Y10_LUT4AB/E2MID[1]
+ Tile_X6Y10_LUT4AB/E2MID[2] Tile_X6Y10_LUT4AB/E2MID[3] Tile_X6Y10_LUT4AB/E2MID[4]
+ Tile_X6Y10_LUT4AB/E2MID[5] Tile_X6Y10_LUT4AB/E2MID[6] Tile_X6Y10_LUT4AB/E2MID[7]
+ Tile_X6Y10_LUT4AB/E2END[0] Tile_X6Y10_LUT4AB/E2END[1] Tile_X6Y10_LUT4AB/E2END[2]
+ Tile_X6Y10_LUT4AB/E2END[3] Tile_X6Y10_LUT4AB/E2END[4] Tile_X6Y10_LUT4AB/E2END[5]
+ Tile_X6Y10_LUT4AB/E2END[6] Tile_X6Y10_LUT4AB/E2END[7] Tile_X5Y10_LUT4AB/E2END[0]
+ Tile_X5Y10_LUT4AB/E2END[1] Tile_X5Y10_LUT4AB/E2END[2] Tile_X5Y10_LUT4AB/E2END[3]
+ Tile_X5Y10_LUT4AB/E2END[4] Tile_X5Y10_LUT4AB/E2END[5] Tile_X5Y10_LUT4AB/E2END[6]
+ Tile_X5Y10_LUT4AB/E2END[7] Tile_X5Y10_LUT4AB/E2MID[0] Tile_X5Y10_LUT4AB/E2MID[1]
+ Tile_X5Y10_LUT4AB/E2MID[2] Tile_X5Y10_LUT4AB/E2MID[3] Tile_X5Y10_LUT4AB/E2MID[4]
+ Tile_X5Y10_LUT4AB/E2MID[5] Tile_X5Y10_LUT4AB/E2MID[6] Tile_X5Y10_LUT4AB/E2MID[7]
+ Tile_X6Y10_LUT4AB/E6END[0] Tile_X6Y10_LUT4AB/E6END[10] Tile_X6Y10_LUT4AB/E6END[11]
+ Tile_X6Y10_LUT4AB/E6END[1] Tile_X6Y10_LUT4AB/E6END[2] Tile_X6Y10_LUT4AB/E6END[3]
+ Tile_X6Y10_LUT4AB/E6END[4] Tile_X6Y10_LUT4AB/E6END[5] Tile_X6Y10_LUT4AB/E6END[6]
+ Tile_X6Y10_LUT4AB/E6END[7] Tile_X6Y10_LUT4AB/E6END[8] Tile_X6Y10_LUT4AB/E6END[9]
+ Tile_X5Y10_LUT4AB/E6END[0] Tile_X5Y10_LUT4AB/E6END[10] Tile_X5Y10_LUT4AB/E6END[11]
+ Tile_X5Y10_LUT4AB/E6END[1] Tile_X5Y10_LUT4AB/E6END[2] Tile_X5Y10_LUT4AB/E6END[3]
+ Tile_X5Y10_LUT4AB/E6END[4] Tile_X5Y10_LUT4AB/E6END[5] Tile_X5Y10_LUT4AB/E6END[6]
+ Tile_X5Y10_LUT4AB/E6END[7] Tile_X5Y10_LUT4AB/E6END[8] Tile_X5Y10_LUT4AB/E6END[9]
+ Tile_X6Y10_LUT4AB/EE4END[0] Tile_X6Y10_LUT4AB/EE4END[10] Tile_X6Y10_LUT4AB/EE4END[11]
+ Tile_X6Y10_LUT4AB/EE4END[12] Tile_X6Y10_LUT4AB/EE4END[13] Tile_X6Y10_LUT4AB/EE4END[14]
+ Tile_X6Y10_LUT4AB/EE4END[15] Tile_X6Y10_LUT4AB/EE4END[1] Tile_X6Y10_LUT4AB/EE4END[2]
+ Tile_X6Y10_LUT4AB/EE4END[3] Tile_X6Y10_LUT4AB/EE4END[4] Tile_X6Y10_LUT4AB/EE4END[5]
+ Tile_X6Y10_LUT4AB/EE4END[6] Tile_X6Y10_LUT4AB/EE4END[7] Tile_X6Y10_LUT4AB/EE4END[8]
+ Tile_X6Y10_LUT4AB/EE4END[9] Tile_X5Y10_LUT4AB/EE4END[0] Tile_X5Y10_LUT4AB/EE4END[10]
+ Tile_X5Y10_LUT4AB/EE4END[11] Tile_X5Y10_LUT4AB/EE4END[12] Tile_X5Y10_LUT4AB/EE4END[13]
+ Tile_X5Y10_LUT4AB/EE4END[14] Tile_X5Y10_LUT4AB/EE4END[15] Tile_X5Y10_LUT4AB/EE4END[1]
+ Tile_X5Y10_LUT4AB/EE4END[2] Tile_X5Y10_LUT4AB/EE4END[3] Tile_X5Y10_LUT4AB/EE4END[4]
+ Tile_X5Y10_LUT4AB/EE4END[5] Tile_X5Y10_LUT4AB/EE4END[6] Tile_X5Y10_LUT4AB/EE4END[7]
+ Tile_X5Y10_LUT4AB/EE4END[8] Tile_X5Y10_LUT4AB/EE4END[9] Tile_X5Y10_LUT4AB/FrameData[0]
+ Tile_X5Y10_LUT4AB/FrameData[10] Tile_X5Y10_LUT4AB/FrameData[11] Tile_X5Y10_LUT4AB/FrameData[12]
+ Tile_X5Y10_LUT4AB/FrameData[13] Tile_X5Y10_LUT4AB/FrameData[14] Tile_X5Y10_LUT4AB/FrameData[15]
+ Tile_X5Y10_LUT4AB/FrameData[16] Tile_X5Y10_LUT4AB/FrameData[17] Tile_X5Y10_LUT4AB/FrameData[18]
+ Tile_X5Y10_LUT4AB/FrameData[19] Tile_X5Y10_LUT4AB/FrameData[1] Tile_X5Y10_LUT4AB/FrameData[20]
+ Tile_X5Y10_LUT4AB/FrameData[21] Tile_X5Y10_LUT4AB/FrameData[22] Tile_X5Y10_LUT4AB/FrameData[23]
+ Tile_X5Y10_LUT4AB/FrameData[24] Tile_X5Y10_LUT4AB/FrameData[25] Tile_X5Y10_LUT4AB/FrameData[26]
+ Tile_X5Y10_LUT4AB/FrameData[27] Tile_X5Y10_LUT4AB/FrameData[28] Tile_X5Y10_LUT4AB/FrameData[29]
+ Tile_X5Y10_LUT4AB/FrameData[2] Tile_X5Y10_LUT4AB/FrameData[30] Tile_X5Y10_LUT4AB/FrameData[31]
+ Tile_X5Y10_LUT4AB/FrameData[3] Tile_X5Y10_LUT4AB/FrameData[4] Tile_X5Y10_LUT4AB/FrameData[5]
+ Tile_X5Y10_LUT4AB/FrameData[6] Tile_X5Y10_LUT4AB/FrameData[7] Tile_X5Y10_LUT4AB/FrameData[8]
+ Tile_X5Y10_LUT4AB/FrameData[9] Tile_X6Y10_LUT4AB/FrameData[0] Tile_X6Y10_LUT4AB/FrameData[10]
+ Tile_X6Y10_LUT4AB/FrameData[11] Tile_X6Y10_LUT4AB/FrameData[12] Tile_X6Y10_LUT4AB/FrameData[13]
+ Tile_X6Y10_LUT4AB/FrameData[14] Tile_X6Y10_LUT4AB/FrameData[15] Tile_X6Y10_LUT4AB/FrameData[16]
+ Tile_X6Y10_LUT4AB/FrameData[17] Tile_X6Y10_LUT4AB/FrameData[18] Tile_X6Y10_LUT4AB/FrameData[19]
+ Tile_X6Y10_LUT4AB/FrameData[1] Tile_X6Y10_LUT4AB/FrameData[20] Tile_X6Y10_LUT4AB/FrameData[21]
+ Tile_X6Y10_LUT4AB/FrameData[22] Tile_X6Y10_LUT4AB/FrameData[23] Tile_X6Y10_LUT4AB/FrameData[24]
+ Tile_X6Y10_LUT4AB/FrameData[25] Tile_X6Y10_LUT4AB/FrameData[26] Tile_X6Y10_LUT4AB/FrameData[27]
+ Tile_X6Y10_LUT4AB/FrameData[28] Tile_X6Y10_LUT4AB/FrameData[29] Tile_X6Y10_LUT4AB/FrameData[2]
+ Tile_X6Y10_LUT4AB/FrameData[30] Tile_X6Y10_LUT4AB/FrameData[31] Tile_X6Y10_LUT4AB/FrameData[3]
+ Tile_X6Y10_LUT4AB/FrameData[4] Tile_X6Y10_LUT4AB/FrameData[5] Tile_X6Y10_LUT4AB/FrameData[6]
+ Tile_X6Y10_LUT4AB/FrameData[7] Tile_X6Y10_LUT4AB/FrameData[8] Tile_X6Y10_LUT4AB/FrameData[9]
+ Tile_X5Y10_LUT4AB/FrameStrobe[0] Tile_X5Y10_LUT4AB/FrameStrobe[10] Tile_X5Y10_LUT4AB/FrameStrobe[11]
+ Tile_X5Y10_LUT4AB/FrameStrobe[12] Tile_X5Y10_LUT4AB/FrameStrobe[13] Tile_X5Y10_LUT4AB/FrameStrobe[14]
+ Tile_X5Y10_LUT4AB/FrameStrobe[15] Tile_X5Y10_LUT4AB/FrameStrobe[16] Tile_X5Y10_LUT4AB/FrameStrobe[17]
+ Tile_X5Y10_LUT4AB/FrameStrobe[18] Tile_X5Y10_LUT4AB/FrameStrobe[19] Tile_X5Y10_LUT4AB/FrameStrobe[1]
+ Tile_X5Y10_LUT4AB/FrameStrobe[2] Tile_X5Y10_LUT4AB/FrameStrobe[3] Tile_X5Y10_LUT4AB/FrameStrobe[4]
+ Tile_X5Y10_LUT4AB/FrameStrobe[5] Tile_X5Y10_LUT4AB/FrameStrobe[6] Tile_X5Y10_LUT4AB/FrameStrobe[7]
+ Tile_X5Y10_LUT4AB/FrameStrobe[8] Tile_X5Y10_LUT4AB/FrameStrobe[9] Tile_X5Y9_LUT4AB/FrameStrobe[0]
+ Tile_X5Y9_LUT4AB/FrameStrobe[10] Tile_X5Y9_LUT4AB/FrameStrobe[11] Tile_X5Y9_LUT4AB/FrameStrobe[12]
+ Tile_X5Y9_LUT4AB/FrameStrobe[13] Tile_X5Y9_LUT4AB/FrameStrobe[14] Tile_X5Y9_LUT4AB/FrameStrobe[15]
+ Tile_X5Y9_LUT4AB/FrameStrobe[16] Tile_X5Y9_LUT4AB/FrameStrobe[17] Tile_X5Y9_LUT4AB/FrameStrobe[18]
+ Tile_X5Y9_LUT4AB/FrameStrobe[19] Tile_X5Y9_LUT4AB/FrameStrobe[1] Tile_X5Y9_LUT4AB/FrameStrobe[2]
+ Tile_X5Y9_LUT4AB/FrameStrobe[3] Tile_X5Y9_LUT4AB/FrameStrobe[4] Tile_X5Y9_LUT4AB/FrameStrobe[5]
+ Tile_X5Y9_LUT4AB/FrameStrobe[6] Tile_X5Y9_LUT4AB/FrameStrobe[7] Tile_X5Y9_LUT4AB/FrameStrobe[8]
+ Tile_X5Y9_LUT4AB/FrameStrobe[9] Tile_X5Y9_LUT4AB/N1END[0] Tile_X5Y9_LUT4AB/N1END[1]
+ Tile_X5Y9_LUT4AB/N1END[2] Tile_X5Y9_LUT4AB/N1END[3] Tile_X5Y11_LUT4AB/N1BEG[0] Tile_X5Y11_LUT4AB/N1BEG[1]
+ Tile_X5Y11_LUT4AB/N1BEG[2] Tile_X5Y11_LUT4AB/N1BEG[3] Tile_X5Y9_LUT4AB/N2MID[0]
+ Tile_X5Y9_LUT4AB/N2MID[1] Tile_X5Y9_LUT4AB/N2MID[2] Tile_X5Y9_LUT4AB/N2MID[3] Tile_X5Y9_LUT4AB/N2MID[4]
+ Tile_X5Y9_LUT4AB/N2MID[5] Tile_X5Y9_LUT4AB/N2MID[6] Tile_X5Y9_LUT4AB/N2MID[7] Tile_X5Y9_LUT4AB/N2END[0]
+ Tile_X5Y9_LUT4AB/N2END[1] Tile_X5Y9_LUT4AB/N2END[2] Tile_X5Y9_LUT4AB/N2END[3] Tile_X5Y9_LUT4AB/N2END[4]
+ Tile_X5Y9_LUT4AB/N2END[5] Tile_X5Y9_LUT4AB/N2END[6] Tile_X5Y9_LUT4AB/N2END[7] Tile_X5Y10_LUT4AB/N2END[0]
+ Tile_X5Y10_LUT4AB/N2END[1] Tile_X5Y10_LUT4AB/N2END[2] Tile_X5Y10_LUT4AB/N2END[3]
+ Tile_X5Y10_LUT4AB/N2END[4] Tile_X5Y10_LUT4AB/N2END[5] Tile_X5Y10_LUT4AB/N2END[6]
+ Tile_X5Y10_LUT4AB/N2END[7] Tile_X5Y11_LUT4AB/N2BEG[0] Tile_X5Y11_LUT4AB/N2BEG[1]
+ Tile_X5Y11_LUT4AB/N2BEG[2] Tile_X5Y11_LUT4AB/N2BEG[3] Tile_X5Y11_LUT4AB/N2BEG[4]
+ Tile_X5Y11_LUT4AB/N2BEG[5] Tile_X5Y11_LUT4AB/N2BEG[6] Tile_X5Y11_LUT4AB/N2BEG[7]
+ Tile_X5Y9_LUT4AB/N4END[0] Tile_X5Y9_LUT4AB/N4END[10] Tile_X5Y9_LUT4AB/N4END[11]
+ Tile_X5Y9_LUT4AB/N4END[12] Tile_X5Y9_LUT4AB/N4END[13] Tile_X5Y9_LUT4AB/N4END[14]
+ Tile_X5Y9_LUT4AB/N4END[15] Tile_X5Y9_LUT4AB/N4END[1] Tile_X5Y9_LUT4AB/N4END[2] Tile_X5Y9_LUT4AB/N4END[3]
+ Tile_X5Y9_LUT4AB/N4END[4] Tile_X5Y9_LUT4AB/N4END[5] Tile_X5Y9_LUT4AB/N4END[6] Tile_X5Y9_LUT4AB/N4END[7]
+ Tile_X5Y9_LUT4AB/N4END[8] Tile_X5Y9_LUT4AB/N4END[9] Tile_X5Y11_LUT4AB/N4BEG[0] Tile_X5Y11_LUT4AB/N4BEG[10]
+ Tile_X5Y11_LUT4AB/N4BEG[11] Tile_X5Y11_LUT4AB/N4BEG[12] Tile_X5Y11_LUT4AB/N4BEG[13]
+ Tile_X5Y11_LUT4AB/N4BEG[14] Tile_X5Y11_LUT4AB/N4BEG[15] Tile_X5Y11_LUT4AB/N4BEG[1]
+ Tile_X5Y11_LUT4AB/N4BEG[2] Tile_X5Y11_LUT4AB/N4BEG[3] Tile_X5Y11_LUT4AB/N4BEG[4]
+ Tile_X5Y11_LUT4AB/N4BEG[5] Tile_X5Y11_LUT4AB/N4BEG[6] Tile_X5Y11_LUT4AB/N4BEG[7]
+ Tile_X5Y11_LUT4AB/N4BEG[8] Tile_X5Y11_LUT4AB/N4BEG[9] Tile_X5Y9_LUT4AB/NN4END[0]
+ Tile_X5Y9_LUT4AB/NN4END[10] Tile_X5Y9_LUT4AB/NN4END[11] Tile_X5Y9_LUT4AB/NN4END[12]
+ Tile_X5Y9_LUT4AB/NN4END[13] Tile_X5Y9_LUT4AB/NN4END[14] Tile_X5Y9_LUT4AB/NN4END[15]
+ Tile_X5Y9_LUT4AB/NN4END[1] Tile_X5Y9_LUT4AB/NN4END[2] Tile_X5Y9_LUT4AB/NN4END[3]
+ Tile_X5Y9_LUT4AB/NN4END[4] Tile_X5Y9_LUT4AB/NN4END[5] Tile_X5Y9_LUT4AB/NN4END[6]
+ Tile_X5Y9_LUT4AB/NN4END[7] Tile_X5Y9_LUT4AB/NN4END[8] Tile_X5Y9_LUT4AB/NN4END[9]
+ Tile_X5Y11_LUT4AB/NN4BEG[0] Tile_X5Y11_LUT4AB/NN4BEG[10] Tile_X5Y11_LUT4AB/NN4BEG[11]
+ Tile_X5Y11_LUT4AB/NN4BEG[12] Tile_X5Y11_LUT4AB/NN4BEG[13] Tile_X5Y11_LUT4AB/NN4BEG[14]
+ Tile_X5Y11_LUT4AB/NN4BEG[15] Tile_X5Y11_LUT4AB/NN4BEG[1] Tile_X5Y11_LUT4AB/NN4BEG[2]
+ Tile_X5Y11_LUT4AB/NN4BEG[3] Tile_X5Y11_LUT4AB/NN4BEG[4] Tile_X5Y11_LUT4AB/NN4BEG[5]
+ Tile_X5Y11_LUT4AB/NN4BEG[6] Tile_X5Y11_LUT4AB/NN4BEG[7] Tile_X5Y11_LUT4AB/NN4BEG[8]
+ Tile_X5Y11_LUT4AB/NN4BEG[9] Tile_X5Y11_LUT4AB/S1END[0] Tile_X5Y11_LUT4AB/S1END[1]
+ Tile_X5Y11_LUT4AB/S1END[2] Tile_X5Y11_LUT4AB/S1END[3] Tile_X5Y9_LUT4AB/S1BEG[0]
+ Tile_X5Y9_LUT4AB/S1BEG[1] Tile_X5Y9_LUT4AB/S1BEG[2] Tile_X5Y9_LUT4AB/S1BEG[3] Tile_X5Y11_LUT4AB/S2MID[0]
+ Tile_X5Y11_LUT4AB/S2MID[1] Tile_X5Y11_LUT4AB/S2MID[2] Tile_X5Y11_LUT4AB/S2MID[3]
+ Tile_X5Y11_LUT4AB/S2MID[4] Tile_X5Y11_LUT4AB/S2MID[5] Tile_X5Y11_LUT4AB/S2MID[6]
+ Tile_X5Y11_LUT4AB/S2MID[7] Tile_X5Y11_LUT4AB/S2END[0] Tile_X5Y11_LUT4AB/S2END[1]
+ Tile_X5Y11_LUT4AB/S2END[2] Tile_X5Y11_LUT4AB/S2END[3] Tile_X5Y11_LUT4AB/S2END[4]
+ Tile_X5Y11_LUT4AB/S2END[5] Tile_X5Y11_LUT4AB/S2END[6] Tile_X5Y11_LUT4AB/S2END[7]
+ Tile_X5Y9_LUT4AB/S2BEGb[0] Tile_X5Y9_LUT4AB/S2BEGb[1] Tile_X5Y9_LUT4AB/S2BEGb[2]
+ Tile_X5Y9_LUT4AB/S2BEGb[3] Tile_X5Y9_LUT4AB/S2BEGb[4] Tile_X5Y9_LUT4AB/S2BEGb[5]
+ Tile_X5Y9_LUT4AB/S2BEGb[6] Tile_X5Y9_LUT4AB/S2BEGb[7] Tile_X5Y9_LUT4AB/S2BEG[0]
+ Tile_X5Y9_LUT4AB/S2BEG[1] Tile_X5Y9_LUT4AB/S2BEG[2] Tile_X5Y9_LUT4AB/S2BEG[3] Tile_X5Y9_LUT4AB/S2BEG[4]
+ Tile_X5Y9_LUT4AB/S2BEG[5] Tile_X5Y9_LUT4AB/S2BEG[6] Tile_X5Y9_LUT4AB/S2BEG[7] Tile_X5Y11_LUT4AB/S4END[0]
+ Tile_X5Y11_LUT4AB/S4END[10] Tile_X5Y11_LUT4AB/S4END[11] Tile_X5Y11_LUT4AB/S4END[12]
+ Tile_X5Y11_LUT4AB/S4END[13] Tile_X5Y11_LUT4AB/S4END[14] Tile_X5Y11_LUT4AB/S4END[15]
+ Tile_X5Y11_LUT4AB/S4END[1] Tile_X5Y11_LUT4AB/S4END[2] Tile_X5Y11_LUT4AB/S4END[3]
+ Tile_X5Y11_LUT4AB/S4END[4] Tile_X5Y11_LUT4AB/S4END[5] Tile_X5Y11_LUT4AB/S4END[6]
+ Tile_X5Y11_LUT4AB/S4END[7] Tile_X5Y11_LUT4AB/S4END[8] Tile_X5Y11_LUT4AB/S4END[9]
+ Tile_X5Y9_LUT4AB/S4BEG[0] Tile_X5Y9_LUT4AB/S4BEG[10] Tile_X5Y9_LUT4AB/S4BEG[11]
+ Tile_X5Y9_LUT4AB/S4BEG[12] Tile_X5Y9_LUT4AB/S4BEG[13] Tile_X5Y9_LUT4AB/S4BEG[14]
+ Tile_X5Y9_LUT4AB/S4BEG[15] Tile_X5Y9_LUT4AB/S4BEG[1] Tile_X5Y9_LUT4AB/S4BEG[2] Tile_X5Y9_LUT4AB/S4BEG[3]
+ Tile_X5Y9_LUT4AB/S4BEG[4] Tile_X5Y9_LUT4AB/S4BEG[5] Tile_X5Y9_LUT4AB/S4BEG[6] Tile_X5Y9_LUT4AB/S4BEG[7]
+ Tile_X5Y9_LUT4AB/S4BEG[8] Tile_X5Y9_LUT4AB/S4BEG[9] Tile_X5Y11_LUT4AB/SS4END[0]
+ Tile_X5Y11_LUT4AB/SS4END[10] Tile_X5Y11_LUT4AB/SS4END[11] Tile_X5Y11_LUT4AB/SS4END[12]
+ Tile_X5Y11_LUT4AB/SS4END[13] Tile_X5Y11_LUT4AB/SS4END[14] Tile_X5Y11_LUT4AB/SS4END[15]
+ Tile_X5Y11_LUT4AB/SS4END[1] Tile_X5Y11_LUT4AB/SS4END[2] Tile_X5Y11_LUT4AB/SS4END[3]
+ Tile_X5Y11_LUT4AB/SS4END[4] Tile_X5Y11_LUT4AB/SS4END[5] Tile_X5Y11_LUT4AB/SS4END[6]
+ Tile_X5Y11_LUT4AB/SS4END[7] Tile_X5Y11_LUT4AB/SS4END[8] Tile_X5Y11_LUT4AB/SS4END[9]
+ Tile_X5Y9_LUT4AB/SS4BEG[0] Tile_X5Y9_LUT4AB/SS4BEG[10] Tile_X5Y9_LUT4AB/SS4BEG[11]
+ Tile_X5Y9_LUT4AB/SS4BEG[12] Tile_X5Y9_LUT4AB/SS4BEG[13] Tile_X5Y9_LUT4AB/SS4BEG[14]
+ Tile_X5Y9_LUT4AB/SS4BEG[15] Tile_X5Y9_LUT4AB/SS4BEG[1] Tile_X5Y9_LUT4AB/SS4BEG[2]
+ Tile_X5Y9_LUT4AB/SS4BEG[3] Tile_X5Y9_LUT4AB/SS4BEG[4] Tile_X5Y9_LUT4AB/SS4BEG[5]
+ Tile_X5Y9_LUT4AB/SS4BEG[6] Tile_X5Y9_LUT4AB/SS4BEG[7] Tile_X5Y9_LUT4AB/SS4BEG[8]
+ Tile_X5Y9_LUT4AB/SS4BEG[9] Tile_X5Y10_LUT4AB/UserCLK Tile_X5Y9_LUT4AB/UserCLK VGND
+ VPWR Tile_X5Y10_LUT4AB/W1BEG[0] Tile_X5Y10_LUT4AB/W1BEG[1] Tile_X5Y10_LUT4AB/W1BEG[2]
+ Tile_X5Y10_LUT4AB/W1BEG[3] Tile_X6Y10_LUT4AB/W1BEG[0] Tile_X6Y10_LUT4AB/W1BEG[1]
+ Tile_X6Y10_LUT4AB/W1BEG[2] Tile_X6Y10_LUT4AB/W1BEG[3] Tile_X5Y10_LUT4AB/W2BEG[0]
+ Tile_X5Y10_LUT4AB/W2BEG[1] Tile_X5Y10_LUT4AB/W2BEG[2] Tile_X5Y10_LUT4AB/W2BEG[3]
+ Tile_X5Y10_LUT4AB/W2BEG[4] Tile_X5Y10_LUT4AB/W2BEG[5] Tile_X5Y10_LUT4AB/W2BEG[6]
+ Tile_X5Y10_LUT4AB/W2BEG[7] Tile_X5Y10_LUT4AB/W2BEGb[0] Tile_X5Y10_LUT4AB/W2BEGb[1]
+ Tile_X5Y10_LUT4AB/W2BEGb[2] Tile_X5Y10_LUT4AB/W2BEGb[3] Tile_X5Y10_LUT4AB/W2BEGb[4]
+ Tile_X5Y10_LUT4AB/W2BEGb[5] Tile_X5Y10_LUT4AB/W2BEGb[6] Tile_X5Y10_LUT4AB/W2BEGb[7]
+ Tile_X5Y10_LUT4AB/W2END[0] Tile_X5Y10_LUT4AB/W2END[1] Tile_X5Y10_LUT4AB/W2END[2]
+ Tile_X5Y10_LUT4AB/W2END[3] Tile_X5Y10_LUT4AB/W2END[4] Tile_X5Y10_LUT4AB/W2END[5]
+ Tile_X5Y10_LUT4AB/W2END[6] Tile_X5Y10_LUT4AB/W2END[7] Tile_X6Y10_LUT4AB/W2BEG[0]
+ Tile_X6Y10_LUT4AB/W2BEG[1] Tile_X6Y10_LUT4AB/W2BEG[2] Tile_X6Y10_LUT4AB/W2BEG[3]
+ Tile_X6Y10_LUT4AB/W2BEG[4] Tile_X6Y10_LUT4AB/W2BEG[5] Tile_X6Y10_LUT4AB/W2BEG[6]
+ Tile_X6Y10_LUT4AB/W2BEG[7] Tile_X5Y10_LUT4AB/W6BEG[0] Tile_X5Y10_LUT4AB/W6BEG[10]
+ Tile_X5Y10_LUT4AB/W6BEG[11] Tile_X5Y10_LUT4AB/W6BEG[1] Tile_X5Y10_LUT4AB/W6BEG[2]
+ Tile_X5Y10_LUT4AB/W6BEG[3] Tile_X5Y10_LUT4AB/W6BEG[4] Tile_X5Y10_LUT4AB/W6BEG[5]
+ Tile_X5Y10_LUT4AB/W6BEG[6] Tile_X5Y10_LUT4AB/W6BEG[7] Tile_X5Y10_LUT4AB/W6BEG[8]
+ Tile_X5Y10_LUT4AB/W6BEG[9] Tile_X6Y10_LUT4AB/W6BEG[0] Tile_X6Y10_LUT4AB/W6BEG[10]
+ Tile_X6Y10_LUT4AB/W6BEG[11] Tile_X6Y10_LUT4AB/W6BEG[1] Tile_X6Y10_LUT4AB/W6BEG[2]
+ Tile_X6Y10_LUT4AB/W6BEG[3] Tile_X6Y10_LUT4AB/W6BEG[4] Tile_X6Y10_LUT4AB/W6BEG[5]
+ Tile_X6Y10_LUT4AB/W6BEG[6] Tile_X6Y10_LUT4AB/W6BEG[7] Tile_X6Y10_LUT4AB/W6BEG[8]
+ Tile_X6Y10_LUT4AB/W6BEG[9] Tile_X5Y10_LUT4AB/WW4BEG[0] Tile_X5Y10_LUT4AB/WW4BEG[10]
+ Tile_X5Y10_LUT4AB/WW4BEG[11] Tile_X5Y10_LUT4AB/WW4BEG[12] Tile_X5Y10_LUT4AB/WW4BEG[13]
+ Tile_X5Y10_LUT4AB/WW4BEG[14] Tile_X5Y10_LUT4AB/WW4BEG[15] Tile_X5Y10_LUT4AB/WW4BEG[1]
+ Tile_X5Y10_LUT4AB/WW4BEG[2] Tile_X5Y10_LUT4AB/WW4BEG[3] Tile_X5Y10_LUT4AB/WW4BEG[4]
+ Tile_X5Y10_LUT4AB/WW4BEG[5] Tile_X5Y10_LUT4AB/WW4BEG[6] Tile_X5Y10_LUT4AB/WW4BEG[7]
+ Tile_X5Y10_LUT4AB/WW4BEG[8] Tile_X5Y10_LUT4AB/WW4BEG[9] Tile_X6Y10_LUT4AB/WW4BEG[0]
+ Tile_X6Y10_LUT4AB/WW4BEG[10] Tile_X6Y10_LUT4AB/WW4BEG[11] Tile_X6Y10_LUT4AB/WW4BEG[12]
+ Tile_X6Y10_LUT4AB/WW4BEG[13] Tile_X6Y10_LUT4AB/WW4BEG[14] Tile_X6Y10_LUT4AB/WW4BEG[15]
+ Tile_X6Y10_LUT4AB/WW4BEG[1] Tile_X6Y10_LUT4AB/WW4BEG[2] Tile_X6Y10_LUT4AB/WW4BEG[3]
+ Tile_X6Y10_LUT4AB/WW4BEG[4] Tile_X6Y10_LUT4AB/WW4BEG[5] Tile_X6Y10_LUT4AB/WW4BEG[6]
+ Tile_X6Y10_LUT4AB/WW4BEG[7] Tile_X6Y10_LUT4AB/WW4BEG[8] Tile_X6Y10_LUT4AB/WW4BEG[9]
+ LUT4AB
XTile_X1Y8_LUT4AB Tile_X1Y9_LUT4AB/Co Tile_X1Y8_LUT4AB/Co Tile_X2Y8_LUT4AB/E1END[0]
+ Tile_X2Y8_LUT4AB/E1END[1] Tile_X2Y8_LUT4AB/E1END[2] Tile_X2Y8_LUT4AB/E1END[3] Tile_X0Y8_W_IO/E1BEG[0]
+ Tile_X0Y8_W_IO/E1BEG[1] Tile_X0Y8_W_IO/E1BEG[2] Tile_X0Y8_W_IO/E1BEG[3] Tile_X2Y8_LUT4AB/E2MID[0]
+ Tile_X2Y8_LUT4AB/E2MID[1] Tile_X2Y8_LUT4AB/E2MID[2] Tile_X2Y8_LUT4AB/E2MID[3] Tile_X2Y8_LUT4AB/E2MID[4]
+ Tile_X2Y8_LUT4AB/E2MID[5] Tile_X2Y8_LUT4AB/E2MID[6] Tile_X2Y8_LUT4AB/E2MID[7] Tile_X2Y8_LUT4AB/E2END[0]
+ Tile_X2Y8_LUT4AB/E2END[1] Tile_X2Y8_LUT4AB/E2END[2] Tile_X2Y8_LUT4AB/E2END[3] Tile_X2Y8_LUT4AB/E2END[4]
+ Tile_X2Y8_LUT4AB/E2END[5] Tile_X2Y8_LUT4AB/E2END[6] Tile_X2Y8_LUT4AB/E2END[7] Tile_X0Y8_W_IO/E2BEGb[0]
+ Tile_X0Y8_W_IO/E2BEGb[1] Tile_X0Y8_W_IO/E2BEGb[2] Tile_X0Y8_W_IO/E2BEGb[3] Tile_X0Y8_W_IO/E2BEGb[4]
+ Tile_X0Y8_W_IO/E2BEGb[5] Tile_X0Y8_W_IO/E2BEGb[6] Tile_X0Y8_W_IO/E2BEGb[7] Tile_X0Y8_W_IO/E2BEG[0]
+ Tile_X0Y8_W_IO/E2BEG[1] Tile_X0Y8_W_IO/E2BEG[2] Tile_X0Y8_W_IO/E2BEG[3] Tile_X0Y8_W_IO/E2BEG[4]
+ Tile_X0Y8_W_IO/E2BEG[5] Tile_X0Y8_W_IO/E2BEG[6] Tile_X0Y8_W_IO/E2BEG[7] Tile_X2Y8_LUT4AB/E6END[0]
+ Tile_X2Y8_LUT4AB/E6END[10] Tile_X2Y8_LUT4AB/E6END[11] Tile_X2Y8_LUT4AB/E6END[1]
+ Tile_X2Y8_LUT4AB/E6END[2] Tile_X2Y8_LUT4AB/E6END[3] Tile_X2Y8_LUT4AB/E6END[4] Tile_X2Y8_LUT4AB/E6END[5]
+ Tile_X2Y8_LUT4AB/E6END[6] Tile_X2Y8_LUT4AB/E6END[7] Tile_X2Y8_LUT4AB/E6END[8] Tile_X2Y8_LUT4AB/E6END[9]
+ Tile_X0Y8_W_IO/E6BEG[0] Tile_X0Y8_W_IO/E6BEG[10] Tile_X0Y8_W_IO/E6BEG[11] Tile_X0Y8_W_IO/E6BEG[1]
+ Tile_X0Y8_W_IO/E6BEG[2] Tile_X0Y8_W_IO/E6BEG[3] Tile_X0Y8_W_IO/E6BEG[4] Tile_X0Y8_W_IO/E6BEG[5]
+ Tile_X0Y8_W_IO/E6BEG[6] Tile_X0Y8_W_IO/E6BEG[7] Tile_X0Y8_W_IO/E6BEG[8] Tile_X0Y8_W_IO/E6BEG[9]
+ Tile_X2Y8_LUT4AB/EE4END[0] Tile_X2Y8_LUT4AB/EE4END[10] Tile_X2Y8_LUT4AB/EE4END[11]
+ Tile_X2Y8_LUT4AB/EE4END[12] Tile_X2Y8_LUT4AB/EE4END[13] Tile_X2Y8_LUT4AB/EE4END[14]
+ Tile_X2Y8_LUT4AB/EE4END[15] Tile_X2Y8_LUT4AB/EE4END[1] Tile_X2Y8_LUT4AB/EE4END[2]
+ Tile_X2Y8_LUT4AB/EE4END[3] Tile_X2Y8_LUT4AB/EE4END[4] Tile_X2Y8_LUT4AB/EE4END[5]
+ Tile_X2Y8_LUT4AB/EE4END[6] Tile_X2Y8_LUT4AB/EE4END[7] Tile_X2Y8_LUT4AB/EE4END[8]
+ Tile_X2Y8_LUT4AB/EE4END[9] Tile_X0Y8_W_IO/EE4BEG[0] Tile_X0Y8_W_IO/EE4BEG[10] Tile_X0Y8_W_IO/EE4BEG[11]
+ Tile_X0Y8_W_IO/EE4BEG[12] Tile_X0Y8_W_IO/EE4BEG[13] Tile_X0Y8_W_IO/EE4BEG[14] Tile_X0Y8_W_IO/EE4BEG[15]
+ Tile_X0Y8_W_IO/EE4BEG[1] Tile_X0Y8_W_IO/EE4BEG[2] Tile_X0Y8_W_IO/EE4BEG[3] Tile_X0Y8_W_IO/EE4BEG[4]
+ Tile_X0Y8_W_IO/EE4BEG[5] Tile_X0Y8_W_IO/EE4BEG[6] Tile_X0Y8_W_IO/EE4BEG[7] Tile_X0Y8_W_IO/EE4BEG[8]
+ Tile_X0Y8_W_IO/EE4BEG[9] Tile_X1Y8_LUT4AB/FrameData[0] Tile_X1Y8_LUT4AB/FrameData[10]
+ Tile_X1Y8_LUT4AB/FrameData[11] Tile_X1Y8_LUT4AB/FrameData[12] Tile_X1Y8_LUT4AB/FrameData[13]
+ Tile_X1Y8_LUT4AB/FrameData[14] Tile_X1Y8_LUT4AB/FrameData[15] Tile_X1Y8_LUT4AB/FrameData[16]
+ Tile_X1Y8_LUT4AB/FrameData[17] Tile_X1Y8_LUT4AB/FrameData[18] Tile_X1Y8_LUT4AB/FrameData[19]
+ Tile_X1Y8_LUT4AB/FrameData[1] Tile_X1Y8_LUT4AB/FrameData[20] Tile_X1Y8_LUT4AB/FrameData[21]
+ Tile_X1Y8_LUT4AB/FrameData[22] Tile_X1Y8_LUT4AB/FrameData[23] Tile_X1Y8_LUT4AB/FrameData[24]
+ Tile_X1Y8_LUT4AB/FrameData[25] Tile_X1Y8_LUT4AB/FrameData[26] Tile_X1Y8_LUT4AB/FrameData[27]
+ Tile_X1Y8_LUT4AB/FrameData[28] Tile_X1Y8_LUT4AB/FrameData[29] Tile_X1Y8_LUT4AB/FrameData[2]
+ Tile_X1Y8_LUT4AB/FrameData[30] Tile_X1Y8_LUT4AB/FrameData[31] Tile_X1Y8_LUT4AB/FrameData[3]
+ Tile_X1Y8_LUT4AB/FrameData[4] Tile_X1Y8_LUT4AB/FrameData[5] Tile_X1Y8_LUT4AB/FrameData[6]
+ Tile_X1Y8_LUT4AB/FrameData[7] Tile_X1Y8_LUT4AB/FrameData[8] Tile_X1Y8_LUT4AB/FrameData[9]
+ Tile_X2Y8_LUT4AB/FrameData[0] Tile_X2Y8_LUT4AB/FrameData[10] Tile_X2Y8_LUT4AB/FrameData[11]
+ Tile_X2Y8_LUT4AB/FrameData[12] Tile_X2Y8_LUT4AB/FrameData[13] Tile_X2Y8_LUT4AB/FrameData[14]
+ Tile_X2Y8_LUT4AB/FrameData[15] Tile_X2Y8_LUT4AB/FrameData[16] Tile_X2Y8_LUT4AB/FrameData[17]
+ Tile_X2Y8_LUT4AB/FrameData[18] Tile_X2Y8_LUT4AB/FrameData[19] Tile_X2Y8_LUT4AB/FrameData[1]
+ Tile_X2Y8_LUT4AB/FrameData[20] Tile_X2Y8_LUT4AB/FrameData[21] Tile_X2Y8_LUT4AB/FrameData[22]
+ Tile_X2Y8_LUT4AB/FrameData[23] Tile_X2Y8_LUT4AB/FrameData[24] Tile_X2Y8_LUT4AB/FrameData[25]
+ Tile_X2Y8_LUT4AB/FrameData[26] Tile_X2Y8_LUT4AB/FrameData[27] Tile_X2Y8_LUT4AB/FrameData[28]
+ Tile_X2Y8_LUT4AB/FrameData[29] Tile_X2Y8_LUT4AB/FrameData[2] Tile_X2Y8_LUT4AB/FrameData[30]
+ Tile_X2Y8_LUT4AB/FrameData[31] Tile_X2Y8_LUT4AB/FrameData[3] Tile_X2Y8_LUT4AB/FrameData[4]
+ Tile_X2Y8_LUT4AB/FrameData[5] Tile_X2Y8_LUT4AB/FrameData[6] Tile_X2Y8_LUT4AB/FrameData[7]
+ Tile_X2Y8_LUT4AB/FrameData[8] Tile_X2Y8_LUT4AB/FrameData[9] Tile_X1Y8_LUT4AB/FrameStrobe[0]
+ Tile_X1Y8_LUT4AB/FrameStrobe[10] Tile_X1Y8_LUT4AB/FrameStrobe[11] Tile_X1Y8_LUT4AB/FrameStrobe[12]
+ Tile_X1Y8_LUT4AB/FrameStrobe[13] Tile_X1Y8_LUT4AB/FrameStrobe[14] Tile_X1Y8_LUT4AB/FrameStrobe[15]
+ Tile_X1Y8_LUT4AB/FrameStrobe[16] Tile_X1Y8_LUT4AB/FrameStrobe[17] Tile_X1Y8_LUT4AB/FrameStrobe[18]
+ Tile_X1Y8_LUT4AB/FrameStrobe[19] Tile_X1Y8_LUT4AB/FrameStrobe[1] Tile_X1Y8_LUT4AB/FrameStrobe[2]
+ Tile_X1Y8_LUT4AB/FrameStrobe[3] Tile_X1Y8_LUT4AB/FrameStrobe[4] Tile_X1Y8_LUT4AB/FrameStrobe[5]
+ Tile_X1Y8_LUT4AB/FrameStrobe[6] Tile_X1Y8_LUT4AB/FrameStrobe[7] Tile_X1Y8_LUT4AB/FrameStrobe[8]
+ Tile_X1Y8_LUT4AB/FrameStrobe[9] Tile_X1Y7_LUT4AB/FrameStrobe[0] Tile_X1Y7_LUT4AB/FrameStrobe[10]
+ Tile_X1Y7_LUT4AB/FrameStrobe[11] Tile_X1Y7_LUT4AB/FrameStrobe[12] Tile_X1Y7_LUT4AB/FrameStrobe[13]
+ Tile_X1Y7_LUT4AB/FrameStrobe[14] Tile_X1Y7_LUT4AB/FrameStrobe[15] Tile_X1Y7_LUT4AB/FrameStrobe[16]
+ Tile_X1Y7_LUT4AB/FrameStrobe[17] Tile_X1Y7_LUT4AB/FrameStrobe[18] Tile_X1Y7_LUT4AB/FrameStrobe[19]
+ Tile_X1Y7_LUT4AB/FrameStrobe[1] Tile_X1Y7_LUT4AB/FrameStrobe[2] Tile_X1Y7_LUT4AB/FrameStrobe[3]
+ Tile_X1Y7_LUT4AB/FrameStrobe[4] Tile_X1Y7_LUT4AB/FrameStrobe[5] Tile_X1Y7_LUT4AB/FrameStrobe[6]
+ Tile_X1Y7_LUT4AB/FrameStrobe[7] Tile_X1Y7_LUT4AB/FrameStrobe[8] Tile_X1Y7_LUT4AB/FrameStrobe[9]
+ Tile_X1Y8_LUT4AB/N1BEG[0] Tile_X1Y8_LUT4AB/N1BEG[1] Tile_X1Y8_LUT4AB/N1BEG[2] Tile_X1Y8_LUT4AB/N1BEG[3]
+ Tile_X1Y9_LUT4AB/N1BEG[0] Tile_X1Y9_LUT4AB/N1BEG[1] Tile_X1Y9_LUT4AB/N1BEG[2] Tile_X1Y9_LUT4AB/N1BEG[3]
+ Tile_X1Y8_LUT4AB/N2BEG[0] Tile_X1Y8_LUT4AB/N2BEG[1] Tile_X1Y8_LUT4AB/N2BEG[2] Tile_X1Y8_LUT4AB/N2BEG[3]
+ Tile_X1Y8_LUT4AB/N2BEG[4] Tile_X1Y8_LUT4AB/N2BEG[5] Tile_X1Y8_LUT4AB/N2BEG[6] Tile_X1Y8_LUT4AB/N2BEG[7]
+ Tile_X1Y7_LUT4AB/N2END[0] Tile_X1Y7_LUT4AB/N2END[1] Tile_X1Y7_LUT4AB/N2END[2] Tile_X1Y7_LUT4AB/N2END[3]
+ Tile_X1Y7_LUT4AB/N2END[4] Tile_X1Y7_LUT4AB/N2END[5] Tile_X1Y7_LUT4AB/N2END[6] Tile_X1Y7_LUT4AB/N2END[7]
+ Tile_X1Y8_LUT4AB/N2END[0] Tile_X1Y8_LUT4AB/N2END[1] Tile_X1Y8_LUT4AB/N2END[2] Tile_X1Y8_LUT4AB/N2END[3]
+ Tile_X1Y8_LUT4AB/N2END[4] Tile_X1Y8_LUT4AB/N2END[5] Tile_X1Y8_LUT4AB/N2END[6] Tile_X1Y8_LUT4AB/N2END[7]
+ Tile_X1Y9_LUT4AB/N2BEG[0] Tile_X1Y9_LUT4AB/N2BEG[1] Tile_X1Y9_LUT4AB/N2BEG[2] Tile_X1Y9_LUT4AB/N2BEG[3]
+ Tile_X1Y9_LUT4AB/N2BEG[4] Tile_X1Y9_LUT4AB/N2BEG[5] Tile_X1Y9_LUT4AB/N2BEG[6] Tile_X1Y9_LUT4AB/N2BEG[7]
+ Tile_X1Y8_LUT4AB/N4BEG[0] Tile_X1Y8_LUT4AB/N4BEG[10] Tile_X1Y8_LUT4AB/N4BEG[11]
+ Tile_X1Y8_LUT4AB/N4BEG[12] Tile_X1Y8_LUT4AB/N4BEG[13] Tile_X1Y8_LUT4AB/N4BEG[14]
+ Tile_X1Y8_LUT4AB/N4BEG[15] Tile_X1Y8_LUT4AB/N4BEG[1] Tile_X1Y8_LUT4AB/N4BEG[2] Tile_X1Y8_LUT4AB/N4BEG[3]
+ Tile_X1Y8_LUT4AB/N4BEG[4] Tile_X1Y8_LUT4AB/N4BEG[5] Tile_X1Y8_LUT4AB/N4BEG[6] Tile_X1Y8_LUT4AB/N4BEG[7]
+ Tile_X1Y8_LUT4AB/N4BEG[8] Tile_X1Y8_LUT4AB/N4BEG[9] Tile_X1Y9_LUT4AB/N4BEG[0] Tile_X1Y9_LUT4AB/N4BEG[10]
+ Tile_X1Y9_LUT4AB/N4BEG[11] Tile_X1Y9_LUT4AB/N4BEG[12] Tile_X1Y9_LUT4AB/N4BEG[13]
+ Tile_X1Y9_LUT4AB/N4BEG[14] Tile_X1Y9_LUT4AB/N4BEG[15] Tile_X1Y9_LUT4AB/N4BEG[1]
+ Tile_X1Y9_LUT4AB/N4BEG[2] Tile_X1Y9_LUT4AB/N4BEG[3] Tile_X1Y9_LUT4AB/N4BEG[4] Tile_X1Y9_LUT4AB/N4BEG[5]
+ Tile_X1Y9_LUT4AB/N4BEG[6] Tile_X1Y9_LUT4AB/N4BEG[7] Tile_X1Y9_LUT4AB/N4BEG[8] Tile_X1Y9_LUT4AB/N4BEG[9]
+ Tile_X1Y8_LUT4AB/NN4BEG[0] Tile_X1Y8_LUT4AB/NN4BEG[10] Tile_X1Y8_LUT4AB/NN4BEG[11]
+ Tile_X1Y8_LUT4AB/NN4BEG[12] Tile_X1Y8_LUT4AB/NN4BEG[13] Tile_X1Y8_LUT4AB/NN4BEG[14]
+ Tile_X1Y8_LUT4AB/NN4BEG[15] Tile_X1Y8_LUT4AB/NN4BEG[1] Tile_X1Y8_LUT4AB/NN4BEG[2]
+ Tile_X1Y8_LUT4AB/NN4BEG[3] Tile_X1Y8_LUT4AB/NN4BEG[4] Tile_X1Y8_LUT4AB/NN4BEG[5]
+ Tile_X1Y8_LUT4AB/NN4BEG[6] Tile_X1Y8_LUT4AB/NN4BEG[7] Tile_X1Y8_LUT4AB/NN4BEG[8]
+ Tile_X1Y8_LUT4AB/NN4BEG[9] Tile_X1Y9_LUT4AB/NN4BEG[0] Tile_X1Y9_LUT4AB/NN4BEG[10]
+ Tile_X1Y9_LUT4AB/NN4BEG[11] Tile_X1Y9_LUT4AB/NN4BEG[12] Tile_X1Y9_LUT4AB/NN4BEG[13]
+ Tile_X1Y9_LUT4AB/NN4BEG[14] Tile_X1Y9_LUT4AB/NN4BEG[15] Tile_X1Y9_LUT4AB/NN4BEG[1]
+ Tile_X1Y9_LUT4AB/NN4BEG[2] Tile_X1Y9_LUT4AB/NN4BEG[3] Tile_X1Y9_LUT4AB/NN4BEG[4]
+ Tile_X1Y9_LUT4AB/NN4BEG[5] Tile_X1Y9_LUT4AB/NN4BEG[6] Tile_X1Y9_LUT4AB/NN4BEG[7]
+ Tile_X1Y9_LUT4AB/NN4BEG[8] Tile_X1Y9_LUT4AB/NN4BEG[9] Tile_X1Y9_LUT4AB/S1END[0]
+ Tile_X1Y9_LUT4AB/S1END[1] Tile_X1Y9_LUT4AB/S1END[2] Tile_X1Y9_LUT4AB/S1END[3] Tile_X1Y8_LUT4AB/S1END[0]
+ Tile_X1Y8_LUT4AB/S1END[1] Tile_X1Y8_LUT4AB/S1END[2] Tile_X1Y8_LUT4AB/S1END[3] Tile_X1Y9_LUT4AB/S2MID[0]
+ Tile_X1Y9_LUT4AB/S2MID[1] Tile_X1Y9_LUT4AB/S2MID[2] Tile_X1Y9_LUT4AB/S2MID[3] Tile_X1Y9_LUT4AB/S2MID[4]
+ Tile_X1Y9_LUT4AB/S2MID[5] Tile_X1Y9_LUT4AB/S2MID[6] Tile_X1Y9_LUT4AB/S2MID[7] Tile_X1Y9_LUT4AB/S2END[0]
+ Tile_X1Y9_LUT4AB/S2END[1] Tile_X1Y9_LUT4AB/S2END[2] Tile_X1Y9_LUT4AB/S2END[3] Tile_X1Y9_LUT4AB/S2END[4]
+ Tile_X1Y9_LUT4AB/S2END[5] Tile_X1Y9_LUT4AB/S2END[6] Tile_X1Y9_LUT4AB/S2END[7] Tile_X1Y8_LUT4AB/S2END[0]
+ Tile_X1Y8_LUT4AB/S2END[1] Tile_X1Y8_LUT4AB/S2END[2] Tile_X1Y8_LUT4AB/S2END[3] Tile_X1Y8_LUT4AB/S2END[4]
+ Tile_X1Y8_LUT4AB/S2END[5] Tile_X1Y8_LUT4AB/S2END[6] Tile_X1Y8_LUT4AB/S2END[7] Tile_X1Y8_LUT4AB/S2MID[0]
+ Tile_X1Y8_LUT4AB/S2MID[1] Tile_X1Y8_LUT4AB/S2MID[2] Tile_X1Y8_LUT4AB/S2MID[3] Tile_X1Y8_LUT4AB/S2MID[4]
+ Tile_X1Y8_LUT4AB/S2MID[5] Tile_X1Y8_LUT4AB/S2MID[6] Tile_X1Y8_LUT4AB/S2MID[7] Tile_X1Y9_LUT4AB/S4END[0]
+ Tile_X1Y9_LUT4AB/S4END[10] Tile_X1Y9_LUT4AB/S4END[11] Tile_X1Y9_LUT4AB/S4END[12]
+ Tile_X1Y9_LUT4AB/S4END[13] Tile_X1Y9_LUT4AB/S4END[14] Tile_X1Y9_LUT4AB/S4END[15]
+ Tile_X1Y9_LUT4AB/S4END[1] Tile_X1Y9_LUT4AB/S4END[2] Tile_X1Y9_LUT4AB/S4END[3] Tile_X1Y9_LUT4AB/S4END[4]
+ Tile_X1Y9_LUT4AB/S4END[5] Tile_X1Y9_LUT4AB/S4END[6] Tile_X1Y9_LUT4AB/S4END[7] Tile_X1Y9_LUT4AB/S4END[8]
+ Tile_X1Y9_LUT4AB/S4END[9] Tile_X1Y8_LUT4AB/S4END[0] Tile_X1Y8_LUT4AB/S4END[10] Tile_X1Y8_LUT4AB/S4END[11]
+ Tile_X1Y8_LUT4AB/S4END[12] Tile_X1Y8_LUT4AB/S4END[13] Tile_X1Y8_LUT4AB/S4END[14]
+ Tile_X1Y8_LUT4AB/S4END[15] Tile_X1Y8_LUT4AB/S4END[1] Tile_X1Y8_LUT4AB/S4END[2] Tile_X1Y8_LUT4AB/S4END[3]
+ Tile_X1Y8_LUT4AB/S4END[4] Tile_X1Y8_LUT4AB/S4END[5] Tile_X1Y8_LUT4AB/S4END[6] Tile_X1Y8_LUT4AB/S4END[7]
+ Tile_X1Y8_LUT4AB/S4END[8] Tile_X1Y8_LUT4AB/S4END[9] Tile_X1Y9_LUT4AB/SS4END[0] Tile_X1Y9_LUT4AB/SS4END[10]
+ Tile_X1Y9_LUT4AB/SS4END[11] Tile_X1Y9_LUT4AB/SS4END[12] Tile_X1Y9_LUT4AB/SS4END[13]
+ Tile_X1Y9_LUT4AB/SS4END[14] Tile_X1Y9_LUT4AB/SS4END[15] Tile_X1Y9_LUT4AB/SS4END[1]
+ Tile_X1Y9_LUT4AB/SS4END[2] Tile_X1Y9_LUT4AB/SS4END[3] Tile_X1Y9_LUT4AB/SS4END[4]
+ Tile_X1Y9_LUT4AB/SS4END[5] Tile_X1Y9_LUT4AB/SS4END[6] Tile_X1Y9_LUT4AB/SS4END[7]
+ Tile_X1Y9_LUT4AB/SS4END[8] Tile_X1Y9_LUT4AB/SS4END[9] Tile_X1Y8_LUT4AB/SS4END[0]
+ Tile_X1Y8_LUT4AB/SS4END[10] Tile_X1Y8_LUT4AB/SS4END[11] Tile_X1Y8_LUT4AB/SS4END[12]
+ Tile_X1Y8_LUT4AB/SS4END[13] Tile_X1Y8_LUT4AB/SS4END[14] Tile_X1Y8_LUT4AB/SS4END[15]
+ Tile_X1Y8_LUT4AB/SS4END[1] Tile_X1Y8_LUT4AB/SS4END[2] Tile_X1Y8_LUT4AB/SS4END[3]
+ Tile_X1Y8_LUT4AB/SS4END[4] Tile_X1Y8_LUT4AB/SS4END[5] Tile_X1Y8_LUT4AB/SS4END[6]
+ Tile_X1Y8_LUT4AB/SS4END[7] Tile_X1Y8_LUT4AB/SS4END[8] Tile_X1Y8_LUT4AB/SS4END[9]
+ Tile_X1Y8_LUT4AB/UserCLK Tile_X1Y7_LUT4AB/UserCLK VGND VPWR Tile_X0Y8_W_IO/W1END[0]
+ Tile_X0Y8_W_IO/W1END[1] Tile_X0Y8_W_IO/W1END[2] Tile_X0Y8_W_IO/W1END[3] Tile_X2Y8_LUT4AB/W1BEG[0]
+ Tile_X2Y8_LUT4AB/W1BEG[1] Tile_X2Y8_LUT4AB/W1BEG[2] Tile_X2Y8_LUT4AB/W1BEG[3] Tile_X0Y8_W_IO/W2MID[0]
+ Tile_X0Y8_W_IO/W2MID[1] Tile_X0Y8_W_IO/W2MID[2] Tile_X0Y8_W_IO/W2MID[3] Tile_X0Y8_W_IO/W2MID[4]
+ Tile_X0Y8_W_IO/W2MID[5] Tile_X0Y8_W_IO/W2MID[6] Tile_X0Y8_W_IO/W2MID[7] Tile_X0Y8_W_IO/W2END[0]
+ Tile_X0Y8_W_IO/W2END[1] Tile_X0Y8_W_IO/W2END[2] Tile_X0Y8_W_IO/W2END[3] Tile_X0Y8_W_IO/W2END[4]
+ Tile_X0Y8_W_IO/W2END[5] Tile_X0Y8_W_IO/W2END[6] Tile_X0Y8_W_IO/W2END[7] Tile_X1Y8_LUT4AB/W2END[0]
+ Tile_X1Y8_LUT4AB/W2END[1] Tile_X1Y8_LUT4AB/W2END[2] Tile_X1Y8_LUT4AB/W2END[3] Tile_X1Y8_LUT4AB/W2END[4]
+ Tile_X1Y8_LUT4AB/W2END[5] Tile_X1Y8_LUT4AB/W2END[6] Tile_X1Y8_LUT4AB/W2END[7] Tile_X2Y8_LUT4AB/W2BEG[0]
+ Tile_X2Y8_LUT4AB/W2BEG[1] Tile_X2Y8_LUT4AB/W2BEG[2] Tile_X2Y8_LUT4AB/W2BEG[3] Tile_X2Y8_LUT4AB/W2BEG[4]
+ Tile_X2Y8_LUT4AB/W2BEG[5] Tile_X2Y8_LUT4AB/W2BEG[6] Tile_X2Y8_LUT4AB/W2BEG[7] Tile_X0Y8_W_IO/W6END[0]
+ Tile_X0Y8_W_IO/W6END[10] Tile_X0Y8_W_IO/W6END[11] Tile_X0Y8_W_IO/W6END[1] Tile_X0Y8_W_IO/W6END[2]
+ Tile_X0Y8_W_IO/W6END[3] Tile_X0Y8_W_IO/W6END[4] Tile_X0Y8_W_IO/W6END[5] Tile_X0Y8_W_IO/W6END[6]
+ Tile_X0Y8_W_IO/W6END[7] Tile_X0Y8_W_IO/W6END[8] Tile_X0Y8_W_IO/W6END[9] Tile_X2Y8_LUT4AB/W6BEG[0]
+ Tile_X2Y8_LUT4AB/W6BEG[10] Tile_X2Y8_LUT4AB/W6BEG[11] Tile_X2Y8_LUT4AB/W6BEG[1]
+ Tile_X2Y8_LUT4AB/W6BEG[2] Tile_X2Y8_LUT4AB/W6BEG[3] Tile_X2Y8_LUT4AB/W6BEG[4] Tile_X2Y8_LUT4AB/W6BEG[5]
+ Tile_X2Y8_LUT4AB/W6BEG[6] Tile_X2Y8_LUT4AB/W6BEG[7] Tile_X2Y8_LUT4AB/W6BEG[8] Tile_X2Y8_LUT4AB/W6BEG[9]
+ Tile_X0Y8_W_IO/WW4END[0] Tile_X0Y8_W_IO/WW4END[10] Tile_X0Y8_W_IO/WW4END[11] Tile_X0Y8_W_IO/WW4END[12]
+ Tile_X0Y8_W_IO/WW4END[13] Tile_X0Y8_W_IO/WW4END[14] Tile_X0Y8_W_IO/WW4END[15] Tile_X0Y8_W_IO/WW4END[1]
+ Tile_X0Y8_W_IO/WW4END[2] Tile_X0Y8_W_IO/WW4END[3] Tile_X0Y8_W_IO/WW4END[4] Tile_X0Y8_W_IO/WW4END[5]
+ Tile_X0Y8_W_IO/WW4END[6] Tile_X0Y8_W_IO/WW4END[7] Tile_X0Y8_W_IO/WW4END[8] Tile_X0Y8_W_IO/WW4END[9]
+ Tile_X2Y8_LUT4AB/WW4BEG[0] Tile_X2Y8_LUT4AB/WW4BEG[10] Tile_X2Y8_LUT4AB/WW4BEG[11]
+ Tile_X2Y8_LUT4AB/WW4BEG[12] Tile_X2Y8_LUT4AB/WW4BEG[13] Tile_X2Y8_LUT4AB/WW4BEG[14]
+ Tile_X2Y8_LUT4AB/WW4BEG[15] Tile_X2Y8_LUT4AB/WW4BEG[1] Tile_X2Y8_LUT4AB/WW4BEG[2]
+ Tile_X2Y8_LUT4AB/WW4BEG[3] Tile_X2Y8_LUT4AB/WW4BEG[4] Tile_X2Y8_LUT4AB/WW4BEG[5]
+ Tile_X2Y8_LUT4AB/WW4BEG[6] Tile_X2Y8_LUT4AB/WW4BEG[7] Tile_X2Y8_LUT4AB/WW4BEG[8]
+ Tile_X2Y8_LUT4AB/WW4BEG[9] LUT4AB
XTile_X4Y5_RegFile Tile_X5Y5_LUT4AB/E1END[0] Tile_X5Y5_LUT4AB/E1END[1] Tile_X5Y5_LUT4AB/E1END[2]
+ Tile_X5Y5_LUT4AB/E1END[3] Tile_X3Y5_LUT4AB/E1BEG[0] Tile_X3Y5_LUT4AB/E1BEG[1] Tile_X3Y5_LUT4AB/E1BEG[2]
+ Tile_X3Y5_LUT4AB/E1BEG[3] Tile_X5Y5_LUT4AB/E2MID[0] Tile_X5Y5_LUT4AB/E2MID[1] Tile_X5Y5_LUT4AB/E2MID[2]
+ Tile_X5Y5_LUT4AB/E2MID[3] Tile_X5Y5_LUT4AB/E2MID[4] Tile_X5Y5_LUT4AB/E2MID[5] Tile_X5Y5_LUT4AB/E2MID[6]
+ Tile_X5Y5_LUT4AB/E2MID[7] Tile_X5Y5_LUT4AB/E2END[0] Tile_X5Y5_LUT4AB/E2END[1] Tile_X5Y5_LUT4AB/E2END[2]
+ Tile_X5Y5_LUT4AB/E2END[3] Tile_X5Y5_LUT4AB/E2END[4] Tile_X5Y5_LUT4AB/E2END[5] Tile_X5Y5_LUT4AB/E2END[6]
+ Tile_X5Y5_LUT4AB/E2END[7] Tile_X4Y5_RegFile/E2END[0] Tile_X4Y5_RegFile/E2END[1]
+ Tile_X4Y5_RegFile/E2END[2] Tile_X4Y5_RegFile/E2END[3] Tile_X4Y5_RegFile/E2END[4]
+ Tile_X4Y5_RegFile/E2END[5] Tile_X4Y5_RegFile/E2END[6] Tile_X4Y5_RegFile/E2END[7]
+ Tile_X3Y5_LUT4AB/E2BEG[0] Tile_X3Y5_LUT4AB/E2BEG[1] Tile_X3Y5_LUT4AB/E2BEG[2] Tile_X3Y5_LUT4AB/E2BEG[3]
+ Tile_X3Y5_LUT4AB/E2BEG[4] Tile_X3Y5_LUT4AB/E2BEG[5] Tile_X3Y5_LUT4AB/E2BEG[6] Tile_X3Y5_LUT4AB/E2BEG[7]
+ Tile_X5Y5_LUT4AB/E6END[0] Tile_X5Y5_LUT4AB/E6END[10] Tile_X5Y5_LUT4AB/E6END[11]
+ Tile_X5Y5_LUT4AB/E6END[1] Tile_X5Y5_LUT4AB/E6END[2] Tile_X5Y5_LUT4AB/E6END[3] Tile_X5Y5_LUT4AB/E6END[4]
+ Tile_X5Y5_LUT4AB/E6END[5] Tile_X5Y5_LUT4AB/E6END[6] Tile_X5Y5_LUT4AB/E6END[7] Tile_X5Y5_LUT4AB/E6END[8]
+ Tile_X5Y5_LUT4AB/E6END[9] Tile_X3Y5_LUT4AB/E6BEG[0] Tile_X3Y5_LUT4AB/E6BEG[10] Tile_X3Y5_LUT4AB/E6BEG[11]
+ Tile_X3Y5_LUT4AB/E6BEG[1] Tile_X3Y5_LUT4AB/E6BEG[2] Tile_X3Y5_LUT4AB/E6BEG[3] Tile_X3Y5_LUT4AB/E6BEG[4]
+ Tile_X3Y5_LUT4AB/E6BEG[5] Tile_X3Y5_LUT4AB/E6BEG[6] Tile_X3Y5_LUT4AB/E6BEG[7] Tile_X3Y5_LUT4AB/E6BEG[8]
+ Tile_X3Y5_LUT4AB/E6BEG[9] Tile_X5Y5_LUT4AB/EE4END[0] Tile_X5Y5_LUT4AB/EE4END[10]
+ Tile_X5Y5_LUT4AB/EE4END[11] Tile_X5Y5_LUT4AB/EE4END[12] Tile_X5Y5_LUT4AB/EE4END[13]
+ Tile_X5Y5_LUT4AB/EE4END[14] Tile_X5Y5_LUT4AB/EE4END[15] Tile_X5Y5_LUT4AB/EE4END[1]
+ Tile_X5Y5_LUT4AB/EE4END[2] Tile_X5Y5_LUT4AB/EE4END[3] Tile_X5Y5_LUT4AB/EE4END[4]
+ Tile_X5Y5_LUT4AB/EE4END[5] Tile_X5Y5_LUT4AB/EE4END[6] Tile_X5Y5_LUT4AB/EE4END[7]
+ Tile_X5Y5_LUT4AB/EE4END[8] Tile_X5Y5_LUT4AB/EE4END[9] Tile_X3Y5_LUT4AB/EE4BEG[0]
+ Tile_X3Y5_LUT4AB/EE4BEG[10] Tile_X3Y5_LUT4AB/EE4BEG[11] Tile_X3Y5_LUT4AB/EE4BEG[12]
+ Tile_X3Y5_LUT4AB/EE4BEG[13] Tile_X3Y5_LUT4AB/EE4BEG[14] Tile_X3Y5_LUT4AB/EE4BEG[15]
+ Tile_X3Y5_LUT4AB/EE4BEG[1] Tile_X3Y5_LUT4AB/EE4BEG[2] Tile_X3Y5_LUT4AB/EE4BEG[3]
+ Tile_X3Y5_LUT4AB/EE4BEG[4] Tile_X3Y5_LUT4AB/EE4BEG[5] Tile_X3Y5_LUT4AB/EE4BEG[6]
+ Tile_X3Y5_LUT4AB/EE4BEG[7] Tile_X3Y5_LUT4AB/EE4BEG[8] Tile_X3Y5_LUT4AB/EE4BEG[9]
+ Tile_X4Y5_RegFile/FrameData[0] Tile_X4Y5_RegFile/FrameData[10] Tile_X4Y5_RegFile/FrameData[11]
+ Tile_X4Y5_RegFile/FrameData[12] Tile_X4Y5_RegFile/FrameData[13] Tile_X4Y5_RegFile/FrameData[14]
+ Tile_X4Y5_RegFile/FrameData[15] Tile_X4Y5_RegFile/FrameData[16] Tile_X4Y5_RegFile/FrameData[17]
+ Tile_X4Y5_RegFile/FrameData[18] Tile_X4Y5_RegFile/FrameData[19] Tile_X4Y5_RegFile/FrameData[1]
+ Tile_X4Y5_RegFile/FrameData[20] Tile_X4Y5_RegFile/FrameData[21] Tile_X4Y5_RegFile/FrameData[22]
+ Tile_X4Y5_RegFile/FrameData[23] Tile_X4Y5_RegFile/FrameData[24] Tile_X4Y5_RegFile/FrameData[25]
+ Tile_X4Y5_RegFile/FrameData[26] Tile_X4Y5_RegFile/FrameData[27] Tile_X4Y5_RegFile/FrameData[28]
+ Tile_X4Y5_RegFile/FrameData[29] Tile_X4Y5_RegFile/FrameData[2] Tile_X4Y5_RegFile/FrameData[30]
+ Tile_X4Y5_RegFile/FrameData[31] Tile_X4Y5_RegFile/FrameData[3] Tile_X4Y5_RegFile/FrameData[4]
+ Tile_X4Y5_RegFile/FrameData[5] Tile_X4Y5_RegFile/FrameData[6] Tile_X4Y5_RegFile/FrameData[7]
+ Tile_X4Y5_RegFile/FrameData[8] Tile_X4Y5_RegFile/FrameData[9] Tile_X5Y5_LUT4AB/FrameData[0]
+ Tile_X5Y5_LUT4AB/FrameData[10] Tile_X5Y5_LUT4AB/FrameData[11] Tile_X5Y5_LUT4AB/FrameData[12]
+ Tile_X5Y5_LUT4AB/FrameData[13] Tile_X5Y5_LUT4AB/FrameData[14] Tile_X5Y5_LUT4AB/FrameData[15]
+ Tile_X5Y5_LUT4AB/FrameData[16] Tile_X5Y5_LUT4AB/FrameData[17] Tile_X5Y5_LUT4AB/FrameData[18]
+ Tile_X5Y5_LUT4AB/FrameData[19] Tile_X5Y5_LUT4AB/FrameData[1] Tile_X5Y5_LUT4AB/FrameData[20]
+ Tile_X5Y5_LUT4AB/FrameData[21] Tile_X5Y5_LUT4AB/FrameData[22] Tile_X5Y5_LUT4AB/FrameData[23]
+ Tile_X5Y5_LUT4AB/FrameData[24] Tile_X5Y5_LUT4AB/FrameData[25] Tile_X5Y5_LUT4AB/FrameData[26]
+ Tile_X5Y5_LUT4AB/FrameData[27] Tile_X5Y5_LUT4AB/FrameData[28] Tile_X5Y5_LUT4AB/FrameData[29]
+ Tile_X5Y5_LUT4AB/FrameData[2] Tile_X5Y5_LUT4AB/FrameData[30] Tile_X5Y5_LUT4AB/FrameData[31]
+ Tile_X5Y5_LUT4AB/FrameData[3] Tile_X5Y5_LUT4AB/FrameData[4] Tile_X5Y5_LUT4AB/FrameData[5]
+ Tile_X5Y5_LUT4AB/FrameData[6] Tile_X5Y5_LUT4AB/FrameData[7] Tile_X5Y5_LUT4AB/FrameData[8]
+ Tile_X5Y5_LUT4AB/FrameData[9] Tile_X4Y5_RegFile/FrameStrobe[0] Tile_X4Y5_RegFile/FrameStrobe[10]
+ Tile_X4Y5_RegFile/FrameStrobe[11] Tile_X4Y5_RegFile/FrameStrobe[12] Tile_X4Y5_RegFile/FrameStrobe[13]
+ Tile_X4Y5_RegFile/FrameStrobe[14] Tile_X4Y5_RegFile/FrameStrobe[15] Tile_X4Y5_RegFile/FrameStrobe[16]
+ Tile_X4Y5_RegFile/FrameStrobe[17] Tile_X4Y5_RegFile/FrameStrobe[18] Tile_X4Y5_RegFile/FrameStrobe[19]
+ Tile_X4Y5_RegFile/FrameStrobe[1] Tile_X4Y5_RegFile/FrameStrobe[2] Tile_X4Y5_RegFile/FrameStrobe[3]
+ Tile_X4Y5_RegFile/FrameStrobe[4] Tile_X4Y5_RegFile/FrameStrobe[5] Tile_X4Y5_RegFile/FrameStrobe[6]
+ Tile_X4Y5_RegFile/FrameStrobe[7] Tile_X4Y5_RegFile/FrameStrobe[8] Tile_X4Y5_RegFile/FrameStrobe[9]
+ Tile_X4Y4_RegFile/FrameStrobe[0] Tile_X4Y4_RegFile/FrameStrobe[10] Tile_X4Y4_RegFile/FrameStrobe[11]
+ Tile_X4Y4_RegFile/FrameStrobe[12] Tile_X4Y4_RegFile/FrameStrobe[13] Tile_X4Y4_RegFile/FrameStrobe[14]
+ Tile_X4Y4_RegFile/FrameStrobe[15] Tile_X4Y4_RegFile/FrameStrobe[16] Tile_X4Y4_RegFile/FrameStrobe[17]
+ Tile_X4Y4_RegFile/FrameStrobe[18] Tile_X4Y4_RegFile/FrameStrobe[19] Tile_X4Y4_RegFile/FrameStrobe[1]
+ Tile_X4Y4_RegFile/FrameStrobe[2] Tile_X4Y4_RegFile/FrameStrobe[3] Tile_X4Y4_RegFile/FrameStrobe[4]
+ Tile_X4Y4_RegFile/FrameStrobe[5] Tile_X4Y4_RegFile/FrameStrobe[6] Tile_X4Y4_RegFile/FrameStrobe[7]
+ Tile_X4Y4_RegFile/FrameStrobe[8] Tile_X4Y4_RegFile/FrameStrobe[9] Tile_X4Y5_RegFile/N1BEG[0]
+ Tile_X4Y5_RegFile/N1BEG[1] Tile_X4Y5_RegFile/N1BEG[2] Tile_X4Y5_RegFile/N1BEG[3]
+ Tile_X4Y6_RegFile/N1BEG[0] Tile_X4Y6_RegFile/N1BEG[1] Tile_X4Y6_RegFile/N1BEG[2]
+ Tile_X4Y6_RegFile/N1BEG[3] Tile_X4Y5_RegFile/N2BEG[0] Tile_X4Y5_RegFile/N2BEG[1]
+ Tile_X4Y5_RegFile/N2BEG[2] Tile_X4Y5_RegFile/N2BEG[3] Tile_X4Y5_RegFile/N2BEG[4]
+ Tile_X4Y5_RegFile/N2BEG[5] Tile_X4Y5_RegFile/N2BEG[6] Tile_X4Y5_RegFile/N2BEG[7]
+ Tile_X4Y4_RegFile/N2END[0] Tile_X4Y4_RegFile/N2END[1] Tile_X4Y4_RegFile/N2END[2]
+ Tile_X4Y4_RegFile/N2END[3] Tile_X4Y4_RegFile/N2END[4] Tile_X4Y4_RegFile/N2END[5]
+ Tile_X4Y4_RegFile/N2END[6] Tile_X4Y4_RegFile/N2END[7] Tile_X4Y5_RegFile/N2END[0]
+ Tile_X4Y5_RegFile/N2END[1] Tile_X4Y5_RegFile/N2END[2] Tile_X4Y5_RegFile/N2END[3]
+ Tile_X4Y5_RegFile/N2END[4] Tile_X4Y5_RegFile/N2END[5] Tile_X4Y5_RegFile/N2END[6]
+ Tile_X4Y5_RegFile/N2END[7] Tile_X4Y6_RegFile/N2BEG[0] Tile_X4Y6_RegFile/N2BEG[1]
+ Tile_X4Y6_RegFile/N2BEG[2] Tile_X4Y6_RegFile/N2BEG[3] Tile_X4Y6_RegFile/N2BEG[4]
+ Tile_X4Y6_RegFile/N2BEG[5] Tile_X4Y6_RegFile/N2BEG[6] Tile_X4Y6_RegFile/N2BEG[7]
+ Tile_X4Y5_RegFile/N4BEG[0] Tile_X4Y5_RegFile/N4BEG[10] Tile_X4Y5_RegFile/N4BEG[11]
+ Tile_X4Y5_RegFile/N4BEG[12] Tile_X4Y5_RegFile/N4BEG[13] Tile_X4Y5_RegFile/N4BEG[14]
+ Tile_X4Y5_RegFile/N4BEG[15] Tile_X4Y5_RegFile/N4BEG[1] Tile_X4Y5_RegFile/N4BEG[2]
+ Tile_X4Y5_RegFile/N4BEG[3] Tile_X4Y5_RegFile/N4BEG[4] Tile_X4Y5_RegFile/N4BEG[5]
+ Tile_X4Y5_RegFile/N4BEG[6] Tile_X4Y5_RegFile/N4BEG[7] Tile_X4Y5_RegFile/N4BEG[8]
+ Tile_X4Y5_RegFile/N4BEG[9] Tile_X4Y6_RegFile/N4BEG[0] Tile_X4Y6_RegFile/N4BEG[10]
+ Tile_X4Y6_RegFile/N4BEG[11] Tile_X4Y6_RegFile/N4BEG[12] Tile_X4Y6_RegFile/N4BEG[13]
+ Tile_X4Y6_RegFile/N4BEG[14] Tile_X4Y6_RegFile/N4BEG[15] Tile_X4Y6_RegFile/N4BEG[1]
+ Tile_X4Y6_RegFile/N4BEG[2] Tile_X4Y6_RegFile/N4BEG[3] Tile_X4Y6_RegFile/N4BEG[4]
+ Tile_X4Y6_RegFile/N4BEG[5] Tile_X4Y6_RegFile/N4BEG[6] Tile_X4Y6_RegFile/N4BEG[7]
+ Tile_X4Y6_RegFile/N4BEG[8] Tile_X4Y6_RegFile/N4BEG[9] Tile_X4Y5_RegFile/NN4BEG[0]
+ Tile_X4Y5_RegFile/NN4BEG[10] Tile_X4Y5_RegFile/NN4BEG[11] Tile_X4Y5_RegFile/NN4BEG[12]
+ Tile_X4Y5_RegFile/NN4BEG[13] Tile_X4Y5_RegFile/NN4BEG[14] Tile_X4Y5_RegFile/NN4BEG[15]
+ Tile_X4Y5_RegFile/NN4BEG[1] Tile_X4Y5_RegFile/NN4BEG[2] Tile_X4Y5_RegFile/NN4BEG[3]
+ Tile_X4Y5_RegFile/NN4BEG[4] Tile_X4Y5_RegFile/NN4BEG[5] Tile_X4Y5_RegFile/NN4BEG[6]
+ Tile_X4Y5_RegFile/NN4BEG[7] Tile_X4Y5_RegFile/NN4BEG[8] Tile_X4Y5_RegFile/NN4BEG[9]
+ Tile_X4Y6_RegFile/NN4BEG[0] Tile_X4Y6_RegFile/NN4BEG[10] Tile_X4Y6_RegFile/NN4BEG[11]
+ Tile_X4Y6_RegFile/NN4BEG[12] Tile_X4Y6_RegFile/NN4BEG[13] Tile_X4Y6_RegFile/NN4BEG[14]
+ Tile_X4Y6_RegFile/NN4BEG[15] Tile_X4Y6_RegFile/NN4BEG[1] Tile_X4Y6_RegFile/NN4BEG[2]
+ Tile_X4Y6_RegFile/NN4BEG[3] Tile_X4Y6_RegFile/NN4BEG[4] Tile_X4Y6_RegFile/NN4BEG[5]
+ Tile_X4Y6_RegFile/NN4BEG[6] Tile_X4Y6_RegFile/NN4BEG[7] Tile_X4Y6_RegFile/NN4BEG[8]
+ Tile_X4Y6_RegFile/NN4BEG[9] Tile_X4Y6_RegFile/S1END[0] Tile_X4Y6_RegFile/S1END[1]
+ Tile_X4Y6_RegFile/S1END[2] Tile_X4Y6_RegFile/S1END[3] Tile_X4Y5_RegFile/S1END[0]
+ Tile_X4Y5_RegFile/S1END[1] Tile_X4Y5_RegFile/S1END[2] Tile_X4Y5_RegFile/S1END[3]
+ Tile_X4Y6_RegFile/S2MID[0] Tile_X4Y6_RegFile/S2MID[1] Tile_X4Y6_RegFile/S2MID[2]
+ Tile_X4Y6_RegFile/S2MID[3] Tile_X4Y6_RegFile/S2MID[4] Tile_X4Y6_RegFile/S2MID[5]
+ Tile_X4Y6_RegFile/S2MID[6] Tile_X4Y6_RegFile/S2MID[7] Tile_X4Y6_RegFile/S2END[0]
+ Tile_X4Y6_RegFile/S2END[1] Tile_X4Y6_RegFile/S2END[2] Tile_X4Y6_RegFile/S2END[3]
+ Tile_X4Y6_RegFile/S2END[4] Tile_X4Y6_RegFile/S2END[5] Tile_X4Y6_RegFile/S2END[6]
+ Tile_X4Y6_RegFile/S2END[7] Tile_X4Y5_RegFile/S2END[0] Tile_X4Y5_RegFile/S2END[1]
+ Tile_X4Y5_RegFile/S2END[2] Tile_X4Y5_RegFile/S2END[3] Tile_X4Y5_RegFile/S2END[4]
+ Tile_X4Y5_RegFile/S2END[5] Tile_X4Y5_RegFile/S2END[6] Tile_X4Y5_RegFile/S2END[7]
+ Tile_X4Y5_RegFile/S2MID[0] Tile_X4Y5_RegFile/S2MID[1] Tile_X4Y5_RegFile/S2MID[2]
+ Tile_X4Y5_RegFile/S2MID[3] Tile_X4Y5_RegFile/S2MID[4] Tile_X4Y5_RegFile/S2MID[5]
+ Tile_X4Y5_RegFile/S2MID[6] Tile_X4Y5_RegFile/S2MID[7] Tile_X4Y6_RegFile/S4END[0]
+ Tile_X4Y6_RegFile/S4END[10] Tile_X4Y6_RegFile/S4END[11] Tile_X4Y6_RegFile/S4END[12]
+ Tile_X4Y6_RegFile/S4END[13] Tile_X4Y6_RegFile/S4END[14] Tile_X4Y6_RegFile/S4END[15]
+ Tile_X4Y6_RegFile/S4END[1] Tile_X4Y6_RegFile/S4END[2] Tile_X4Y6_RegFile/S4END[3]
+ Tile_X4Y6_RegFile/S4END[4] Tile_X4Y6_RegFile/S4END[5] Tile_X4Y6_RegFile/S4END[6]
+ Tile_X4Y6_RegFile/S4END[7] Tile_X4Y6_RegFile/S4END[8] Tile_X4Y6_RegFile/S4END[9]
+ Tile_X4Y5_RegFile/S4END[0] Tile_X4Y5_RegFile/S4END[10] Tile_X4Y5_RegFile/S4END[11]
+ Tile_X4Y5_RegFile/S4END[12] Tile_X4Y5_RegFile/S4END[13] Tile_X4Y5_RegFile/S4END[14]
+ Tile_X4Y5_RegFile/S4END[15] Tile_X4Y5_RegFile/S4END[1] Tile_X4Y5_RegFile/S4END[2]
+ Tile_X4Y5_RegFile/S4END[3] Tile_X4Y5_RegFile/S4END[4] Tile_X4Y5_RegFile/S4END[5]
+ Tile_X4Y5_RegFile/S4END[6] Tile_X4Y5_RegFile/S4END[7] Tile_X4Y5_RegFile/S4END[8]
+ Tile_X4Y5_RegFile/S4END[9] Tile_X4Y6_RegFile/SS4END[0] Tile_X4Y6_RegFile/SS4END[10]
+ Tile_X4Y6_RegFile/SS4END[11] Tile_X4Y6_RegFile/SS4END[12] Tile_X4Y6_RegFile/SS4END[13]
+ Tile_X4Y6_RegFile/SS4END[14] Tile_X4Y6_RegFile/SS4END[15] Tile_X4Y6_RegFile/SS4END[1]
+ Tile_X4Y6_RegFile/SS4END[2] Tile_X4Y6_RegFile/SS4END[3] Tile_X4Y6_RegFile/SS4END[4]
+ Tile_X4Y6_RegFile/SS4END[5] Tile_X4Y6_RegFile/SS4END[6] Tile_X4Y6_RegFile/SS4END[7]
+ Tile_X4Y6_RegFile/SS4END[8] Tile_X4Y6_RegFile/SS4END[9] Tile_X4Y5_RegFile/SS4END[0]
+ Tile_X4Y5_RegFile/SS4END[10] Tile_X4Y5_RegFile/SS4END[11] Tile_X4Y5_RegFile/SS4END[12]
+ Tile_X4Y5_RegFile/SS4END[13] Tile_X4Y5_RegFile/SS4END[14] Tile_X4Y5_RegFile/SS4END[15]
+ Tile_X4Y5_RegFile/SS4END[1] Tile_X4Y5_RegFile/SS4END[2] Tile_X4Y5_RegFile/SS4END[3]
+ Tile_X4Y5_RegFile/SS4END[4] Tile_X4Y5_RegFile/SS4END[5] Tile_X4Y5_RegFile/SS4END[6]
+ Tile_X4Y5_RegFile/SS4END[7] Tile_X4Y5_RegFile/SS4END[8] Tile_X4Y5_RegFile/SS4END[9]
+ Tile_X4Y5_RegFile/UserCLK Tile_X4Y4_RegFile/UserCLK VGND VPWR Tile_X3Y5_LUT4AB/W1END[0]
+ Tile_X3Y5_LUT4AB/W1END[1] Tile_X3Y5_LUT4AB/W1END[2] Tile_X3Y5_LUT4AB/W1END[3] Tile_X5Y5_LUT4AB/W1BEG[0]
+ Tile_X5Y5_LUT4AB/W1BEG[1] Tile_X5Y5_LUT4AB/W1BEG[2] Tile_X5Y5_LUT4AB/W1BEG[3] Tile_X3Y5_LUT4AB/W2MID[0]
+ Tile_X3Y5_LUT4AB/W2MID[1] Tile_X3Y5_LUT4AB/W2MID[2] Tile_X3Y5_LUT4AB/W2MID[3] Tile_X3Y5_LUT4AB/W2MID[4]
+ Tile_X3Y5_LUT4AB/W2MID[5] Tile_X3Y5_LUT4AB/W2MID[6] Tile_X3Y5_LUT4AB/W2MID[7] Tile_X3Y5_LUT4AB/W2END[0]
+ Tile_X3Y5_LUT4AB/W2END[1] Tile_X3Y5_LUT4AB/W2END[2] Tile_X3Y5_LUT4AB/W2END[3] Tile_X3Y5_LUT4AB/W2END[4]
+ Tile_X3Y5_LUT4AB/W2END[5] Tile_X3Y5_LUT4AB/W2END[6] Tile_X3Y5_LUT4AB/W2END[7] Tile_X5Y5_LUT4AB/W2BEGb[0]
+ Tile_X5Y5_LUT4AB/W2BEGb[1] Tile_X5Y5_LUT4AB/W2BEGb[2] Tile_X5Y5_LUT4AB/W2BEGb[3]
+ Tile_X5Y5_LUT4AB/W2BEGb[4] Tile_X5Y5_LUT4AB/W2BEGb[5] Tile_X5Y5_LUT4AB/W2BEGb[6]
+ Tile_X5Y5_LUT4AB/W2BEGb[7] Tile_X5Y5_LUT4AB/W2BEG[0] Tile_X5Y5_LUT4AB/W2BEG[1] Tile_X5Y5_LUT4AB/W2BEG[2]
+ Tile_X5Y5_LUT4AB/W2BEG[3] Tile_X5Y5_LUT4AB/W2BEG[4] Tile_X5Y5_LUT4AB/W2BEG[5] Tile_X5Y5_LUT4AB/W2BEG[6]
+ Tile_X5Y5_LUT4AB/W2BEG[7] Tile_X3Y5_LUT4AB/W6END[0] Tile_X3Y5_LUT4AB/W6END[10] Tile_X3Y5_LUT4AB/W6END[11]
+ Tile_X3Y5_LUT4AB/W6END[1] Tile_X3Y5_LUT4AB/W6END[2] Tile_X3Y5_LUT4AB/W6END[3] Tile_X3Y5_LUT4AB/W6END[4]
+ Tile_X3Y5_LUT4AB/W6END[5] Tile_X3Y5_LUT4AB/W6END[6] Tile_X3Y5_LUT4AB/W6END[7] Tile_X3Y5_LUT4AB/W6END[8]
+ Tile_X3Y5_LUT4AB/W6END[9] Tile_X5Y5_LUT4AB/W6BEG[0] Tile_X5Y5_LUT4AB/W6BEG[10] Tile_X5Y5_LUT4AB/W6BEG[11]
+ Tile_X5Y5_LUT4AB/W6BEG[1] Tile_X5Y5_LUT4AB/W6BEG[2] Tile_X5Y5_LUT4AB/W6BEG[3] Tile_X5Y5_LUT4AB/W6BEG[4]
+ Tile_X5Y5_LUT4AB/W6BEG[5] Tile_X5Y5_LUT4AB/W6BEG[6] Tile_X5Y5_LUT4AB/W6BEG[7] Tile_X5Y5_LUT4AB/W6BEG[8]
+ Tile_X5Y5_LUT4AB/W6BEG[9] Tile_X3Y5_LUT4AB/WW4END[0] Tile_X3Y5_LUT4AB/WW4END[10]
+ Tile_X3Y5_LUT4AB/WW4END[11] Tile_X3Y5_LUT4AB/WW4END[12] Tile_X3Y5_LUT4AB/WW4END[13]
+ Tile_X3Y5_LUT4AB/WW4END[14] Tile_X3Y5_LUT4AB/WW4END[15] Tile_X3Y5_LUT4AB/WW4END[1]
+ Tile_X3Y5_LUT4AB/WW4END[2] Tile_X3Y5_LUT4AB/WW4END[3] Tile_X3Y5_LUT4AB/WW4END[4]
+ Tile_X3Y5_LUT4AB/WW4END[5] Tile_X3Y5_LUT4AB/WW4END[6] Tile_X3Y5_LUT4AB/WW4END[7]
+ Tile_X3Y5_LUT4AB/WW4END[8] Tile_X3Y5_LUT4AB/WW4END[9] Tile_X5Y5_LUT4AB/WW4BEG[0]
+ Tile_X5Y5_LUT4AB/WW4BEG[10] Tile_X5Y5_LUT4AB/WW4BEG[11] Tile_X5Y5_LUT4AB/WW4BEG[12]
+ Tile_X5Y5_LUT4AB/WW4BEG[13] Tile_X5Y5_LUT4AB/WW4BEG[14] Tile_X5Y5_LUT4AB/WW4BEG[15]
+ Tile_X5Y5_LUT4AB/WW4BEG[1] Tile_X5Y5_LUT4AB/WW4BEG[2] Tile_X5Y5_LUT4AB/WW4BEG[3]
+ Tile_X5Y5_LUT4AB/WW4BEG[4] Tile_X5Y5_LUT4AB/WW4BEG[5] Tile_X5Y5_LUT4AB/WW4BEG[6]
+ Tile_X5Y5_LUT4AB/WW4BEG[7] Tile_X5Y5_LUT4AB/WW4BEG[8] Tile_X5Y5_LUT4AB/WW4BEG[9]
+ RegFile
XTile_X8Y3_LUT4AB Tile_X8Y4_LUT4AB/Co Tile_X8Y3_LUT4AB/Co Tile_X9Y3_LUT4AB/E1END[0]
+ Tile_X9Y3_LUT4AB/E1END[1] Tile_X9Y3_LUT4AB/E1END[2] Tile_X9Y3_LUT4AB/E1END[3] Tile_X8Y3_LUT4AB/E1END[0]
+ Tile_X8Y3_LUT4AB/E1END[1] Tile_X8Y3_LUT4AB/E1END[2] Tile_X8Y3_LUT4AB/E1END[3] Tile_X9Y3_LUT4AB/E2MID[0]
+ Tile_X9Y3_LUT4AB/E2MID[1] Tile_X9Y3_LUT4AB/E2MID[2] Tile_X9Y3_LUT4AB/E2MID[3] Tile_X9Y3_LUT4AB/E2MID[4]
+ Tile_X9Y3_LUT4AB/E2MID[5] Tile_X9Y3_LUT4AB/E2MID[6] Tile_X9Y3_LUT4AB/E2MID[7] Tile_X9Y3_LUT4AB/E2END[0]
+ Tile_X9Y3_LUT4AB/E2END[1] Tile_X9Y3_LUT4AB/E2END[2] Tile_X9Y3_LUT4AB/E2END[3] Tile_X9Y3_LUT4AB/E2END[4]
+ Tile_X9Y3_LUT4AB/E2END[5] Tile_X9Y3_LUT4AB/E2END[6] Tile_X9Y3_LUT4AB/E2END[7] Tile_X8Y3_LUT4AB/E2END[0]
+ Tile_X8Y3_LUT4AB/E2END[1] Tile_X8Y3_LUT4AB/E2END[2] Tile_X8Y3_LUT4AB/E2END[3] Tile_X8Y3_LUT4AB/E2END[4]
+ Tile_X8Y3_LUT4AB/E2END[5] Tile_X8Y3_LUT4AB/E2END[6] Tile_X8Y3_LUT4AB/E2END[7] Tile_X8Y3_LUT4AB/E2MID[0]
+ Tile_X8Y3_LUT4AB/E2MID[1] Tile_X8Y3_LUT4AB/E2MID[2] Tile_X8Y3_LUT4AB/E2MID[3] Tile_X8Y3_LUT4AB/E2MID[4]
+ Tile_X8Y3_LUT4AB/E2MID[5] Tile_X8Y3_LUT4AB/E2MID[6] Tile_X8Y3_LUT4AB/E2MID[7] Tile_X9Y3_LUT4AB/E6END[0]
+ Tile_X9Y3_LUT4AB/E6END[10] Tile_X9Y3_LUT4AB/E6END[11] Tile_X9Y3_LUT4AB/E6END[1]
+ Tile_X9Y3_LUT4AB/E6END[2] Tile_X9Y3_LUT4AB/E6END[3] Tile_X9Y3_LUT4AB/E6END[4] Tile_X9Y3_LUT4AB/E6END[5]
+ Tile_X9Y3_LUT4AB/E6END[6] Tile_X9Y3_LUT4AB/E6END[7] Tile_X9Y3_LUT4AB/E6END[8] Tile_X9Y3_LUT4AB/E6END[9]
+ Tile_X8Y3_LUT4AB/E6END[0] Tile_X8Y3_LUT4AB/E6END[10] Tile_X8Y3_LUT4AB/E6END[11]
+ Tile_X8Y3_LUT4AB/E6END[1] Tile_X8Y3_LUT4AB/E6END[2] Tile_X8Y3_LUT4AB/E6END[3] Tile_X8Y3_LUT4AB/E6END[4]
+ Tile_X8Y3_LUT4AB/E6END[5] Tile_X8Y3_LUT4AB/E6END[6] Tile_X8Y3_LUT4AB/E6END[7] Tile_X8Y3_LUT4AB/E6END[8]
+ Tile_X8Y3_LUT4AB/E6END[9] Tile_X9Y3_LUT4AB/EE4END[0] Tile_X9Y3_LUT4AB/EE4END[10]
+ Tile_X9Y3_LUT4AB/EE4END[11] Tile_X9Y3_LUT4AB/EE4END[12] Tile_X9Y3_LUT4AB/EE4END[13]
+ Tile_X9Y3_LUT4AB/EE4END[14] Tile_X9Y3_LUT4AB/EE4END[15] Tile_X9Y3_LUT4AB/EE4END[1]
+ Tile_X9Y3_LUT4AB/EE4END[2] Tile_X9Y3_LUT4AB/EE4END[3] Tile_X9Y3_LUT4AB/EE4END[4]
+ Tile_X9Y3_LUT4AB/EE4END[5] Tile_X9Y3_LUT4AB/EE4END[6] Tile_X9Y3_LUT4AB/EE4END[7]
+ Tile_X9Y3_LUT4AB/EE4END[8] Tile_X9Y3_LUT4AB/EE4END[9] Tile_X8Y3_LUT4AB/EE4END[0]
+ Tile_X8Y3_LUT4AB/EE4END[10] Tile_X8Y3_LUT4AB/EE4END[11] Tile_X8Y3_LUT4AB/EE4END[12]
+ Tile_X8Y3_LUT4AB/EE4END[13] Tile_X8Y3_LUT4AB/EE4END[14] Tile_X8Y3_LUT4AB/EE4END[15]
+ Tile_X8Y3_LUT4AB/EE4END[1] Tile_X8Y3_LUT4AB/EE4END[2] Tile_X8Y3_LUT4AB/EE4END[3]
+ Tile_X8Y3_LUT4AB/EE4END[4] Tile_X8Y3_LUT4AB/EE4END[5] Tile_X8Y3_LUT4AB/EE4END[6]
+ Tile_X8Y3_LUT4AB/EE4END[7] Tile_X8Y3_LUT4AB/EE4END[8] Tile_X8Y3_LUT4AB/EE4END[9]
+ Tile_X8Y3_LUT4AB/FrameData[0] Tile_X8Y3_LUT4AB/FrameData[10] Tile_X8Y3_LUT4AB/FrameData[11]
+ Tile_X8Y3_LUT4AB/FrameData[12] Tile_X8Y3_LUT4AB/FrameData[13] Tile_X8Y3_LUT4AB/FrameData[14]
+ Tile_X8Y3_LUT4AB/FrameData[15] Tile_X8Y3_LUT4AB/FrameData[16] Tile_X8Y3_LUT4AB/FrameData[17]
+ Tile_X8Y3_LUT4AB/FrameData[18] Tile_X8Y3_LUT4AB/FrameData[19] Tile_X8Y3_LUT4AB/FrameData[1]
+ Tile_X8Y3_LUT4AB/FrameData[20] Tile_X8Y3_LUT4AB/FrameData[21] Tile_X8Y3_LUT4AB/FrameData[22]
+ Tile_X8Y3_LUT4AB/FrameData[23] Tile_X8Y3_LUT4AB/FrameData[24] Tile_X8Y3_LUT4AB/FrameData[25]
+ Tile_X8Y3_LUT4AB/FrameData[26] Tile_X8Y3_LUT4AB/FrameData[27] Tile_X8Y3_LUT4AB/FrameData[28]
+ Tile_X8Y3_LUT4AB/FrameData[29] Tile_X8Y3_LUT4AB/FrameData[2] Tile_X8Y3_LUT4AB/FrameData[30]
+ Tile_X8Y3_LUT4AB/FrameData[31] Tile_X8Y3_LUT4AB/FrameData[3] Tile_X8Y3_LUT4AB/FrameData[4]
+ Tile_X8Y3_LUT4AB/FrameData[5] Tile_X8Y3_LUT4AB/FrameData[6] Tile_X8Y3_LUT4AB/FrameData[7]
+ Tile_X8Y3_LUT4AB/FrameData[8] Tile_X8Y3_LUT4AB/FrameData[9] Tile_X9Y3_LUT4AB/FrameData[0]
+ Tile_X9Y3_LUT4AB/FrameData[10] Tile_X9Y3_LUT4AB/FrameData[11] Tile_X9Y3_LUT4AB/FrameData[12]
+ Tile_X9Y3_LUT4AB/FrameData[13] Tile_X9Y3_LUT4AB/FrameData[14] Tile_X9Y3_LUT4AB/FrameData[15]
+ Tile_X9Y3_LUT4AB/FrameData[16] Tile_X9Y3_LUT4AB/FrameData[17] Tile_X9Y3_LUT4AB/FrameData[18]
+ Tile_X9Y3_LUT4AB/FrameData[19] Tile_X9Y3_LUT4AB/FrameData[1] Tile_X9Y3_LUT4AB/FrameData[20]
+ Tile_X9Y3_LUT4AB/FrameData[21] Tile_X9Y3_LUT4AB/FrameData[22] Tile_X9Y3_LUT4AB/FrameData[23]
+ Tile_X9Y3_LUT4AB/FrameData[24] Tile_X9Y3_LUT4AB/FrameData[25] Tile_X9Y3_LUT4AB/FrameData[26]
+ Tile_X9Y3_LUT4AB/FrameData[27] Tile_X9Y3_LUT4AB/FrameData[28] Tile_X9Y3_LUT4AB/FrameData[29]
+ Tile_X9Y3_LUT4AB/FrameData[2] Tile_X9Y3_LUT4AB/FrameData[30] Tile_X9Y3_LUT4AB/FrameData[31]
+ Tile_X9Y3_LUT4AB/FrameData[3] Tile_X9Y3_LUT4AB/FrameData[4] Tile_X9Y3_LUT4AB/FrameData[5]
+ Tile_X9Y3_LUT4AB/FrameData[6] Tile_X9Y3_LUT4AB/FrameData[7] Tile_X9Y3_LUT4AB/FrameData[8]
+ Tile_X9Y3_LUT4AB/FrameData[9] Tile_X8Y3_LUT4AB/FrameStrobe[0] Tile_X8Y3_LUT4AB/FrameStrobe[10]
+ Tile_X8Y3_LUT4AB/FrameStrobe[11] Tile_X8Y3_LUT4AB/FrameStrobe[12] Tile_X8Y3_LUT4AB/FrameStrobe[13]
+ Tile_X8Y3_LUT4AB/FrameStrobe[14] Tile_X8Y3_LUT4AB/FrameStrobe[15] Tile_X8Y3_LUT4AB/FrameStrobe[16]
+ Tile_X8Y3_LUT4AB/FrameStrobe[17] Tile_X8Y3_LUT4AB/FrameStrobe[18] Tile_X8Y3_LUT4AB/FrameStrobe[19]
+ Tile_X8Y3_LUT4AB/FrameStrobe[1] Tile_X8Y3_LUT4AB/FrameStrobe[2] Tile_X8Y3_LUT4AB/FrameStrobe[3]
+ Tile_X8Y3_LUT4AB/FrameStrobe[4] Tile_X8Y3_LUT4AB/FrameStrobe[5] Tile_X8Y3_LUT4AB/FrameStrobe[6]
+ Tile_X8Y3_LUT4AB/FrameStrobe[7] Tile_X8Y3_LUT4AB/FrameStrobe[8] Tile_X8Y3_LUT4AB/FrameStrobe[9]
+ Tile_X8Y2_LUT4AB/FrameStrobe[0] Tile_X8Y2_LUT4AB/FrameStrobe[10] Tile_X8Y2_LUT4AB/FrameStrobe[11]
+ Tile_X8Y2_LUT4AB/FrameStrobe[12] Tile_X8Y2_LUT4AB/FrameStrobe[13] Tile_X8Y2_LUT4AB/FrameStrobe[14]
+ Tile_X8Y2_LUT4AB/FrameStrobe[15] Tile_X8Y2_LUT4AB/FrameStrobe[16] Tile_X8Y2_LUT4AB/FrameStrobe[17]
+ Tile_X8Y2_LUT4AB/FrameStrobe[18] Tile_X8Y2_LUT4AB/FrameStrobe[19] Tile_X8Y2_LUT4AB/FrameStrobe[1]
+ Tile_X8Y2_LUT4AB/FrameStrobe[2] Tile_X8Y2_LUT4AB/FrameStrobe[3] Tile_X8Y2_LUT4AB/FrameStrobe[4]
+ Tile_X8Y2_LUT4AB/FrameStrobe[5] Tile_X8Y2_LUT4AB/FrameStrobe[6] Tile_X8Y2_LUT4AB/FrameStrobe[7]
+ Tile_X8Y2_LUT4AB/FrameStrobe[8] Tile_X8Y2_LUT4AB/FrameStrobe[9] Tile_X8Y3_LUT4AB/N1BEG[0]
+ Tile_X8Y3_LUT4AB/N1BEG[1] Tile_X8Y3_LUT4AB/N1BEG[2] Tile_X8Y3_LUT4AB/N1BEG[3] Tile_X8Y4_LUT4AB/N1BEG[0]
+ Tile_X8Y4_LUT4AB/N1BEG[1] Tile_X8Y4_LUT4AB/N1BEG[2] Tile_X8Y4_LUT4AB/N1BEG[3] Tile_X8Y3_LUT4AB/N2BEG[0]
+ Tile_X8Y3_LUT4AB/N2BEG[1] Tile_X8Y3_LUT4AB/N2BEG[2] Tile_X8Y3_LUT4AB/N2BEG[3] Tile_X8Y3_LUT4AB/N2BEG[4]
+ Tile_X8Y3_LUT4AB/N2BEG[5] Tile_X8Y3_LUT4AB/N2BEG[6] Tile_X8Y3_LUT4AB/N2BEG[7] Tile_X8Y2_LUT4AB/N2END[0]
+ Tile_X8Y2_LUT4AB/N2END[1] Tile_X8Y2_LUT4AB/N2END[2] Tile_X8Y2_LUT4AB/N2END[3] Tile_X8Y2_LUT4AB/N2END[4]
+ Tile_X8Y2_LUT4AB/N2END[5] Tile_X8Y2_LUT4AB/N2END[6] Tile_X8Y2_LUT4AB/N2END[7] Tile_X8Y3_LUT4AB/N2END[0]
+ Tile_X8Y3_LUT4AB/N2END[1] Tile_X8Y3_LUT4AB/N2END[2] Tile_X8Y3_LUT4AB/N2END[3] Tile_X8Y3_LUT4AB/N2END[4]
+ Tile_X8Y3_LUT4AB/N2END[5] Tile_X8Y3_LUT4AB/N2END[6] Tile_X8Y3_LUT4AB/N2END[7] Tile_X8Y4_LUT4AB/N2BEG[0]
+ Tile_X8Y4_LUT4AB/N2BEG[1] Tile_X8Y4_LUT4AB/N2BEG[2] Tile_X8Y4_LUT4AB/N2BEG[3] Tile_X8Y4_LUT4AB/N2BEG[4]
+ Tile_X8Y4_LUT4AB/N2BEG[5] Tile_X8Y4_LUT4AB/N2BEG[6] Tile_X8Y4_LUT4AB/N2BEG[7] Tile_X8Y3_LUT4AB/N4BEG[0]
+ Tile_X8Y3_LUT4AB/N4BEG[10] Tile_X8Y3_LUT4AB/N4BEG[11] Tile_X8Y3_LUT4AB/N4BEG[12]
+ Tile_X8Y3_LUT4AB/N4BEG[13] Tile_X8Y3_LUT4AB/N4BEG[14] Tile_X8Y3_LUT4AB/N4BEG[15]
+ Tile_X8Y3_LUT4AB/N4BEG[1] Tile_X8Y3_LUT4AB/N4BEG[2] Tile_X8Y3_LUT4AB/N4BEG[3] Tile_X8Y3_LUT4AB/N4BEG[4]
+ Tile_X8Y3_LUT4AB/N4BEG[5] Tile_X8Y3_LUT4AB/N4BEG[6] Tile_X8Y3_LUT4AB/N4BEG[7] Tile_X8Y3_LUT4AB/N4BEG[8]
+ Tile_X8Y3_LUT4AB/N4BEG[9] Tile_X8Y4_LUT4AB/N4BEG[0] Tile_X8Y4_LUT4AB/N4BEG[10] Tile_X8Y4_LUT4AB/N4BEG[11]
+ Tile_X8Y4_LUT4AB/N4BEG[12] Tile_X8Y4_LUT4AB/N4BEG[13] Tile_X8Y4_LUT4AB/N4BEG[14]
+ Tile_X8Y4_LUT4AB/N4BEG[15] Tile_X8Y4_LUT4AB/N4BEG[1] Tile_X8Y4_LUT4AB/N4BEG[2] Tile_X8Y4_LUT4AB/N4BEG[3]
+ Tile_X8Y4_LUT4AB/N4BEG[4] Tile_X8Y4_LUT4AB/N4BEG[5] Tile_X8Y4_LUT4AB/N4BEG[6] Tile_X8Y4_LUT4AB/N4BEG[7]
+ Tile_X8Y4_LUT4AB/N4BEG[8] Tile_X8Y4_LUT4AB/N4BEG[9] Tile_X8Y3_LUT4AB/NN4BEG[0] Tile_X8Y3_LUT4AB/NN4BEG[10]
+ Tile_X8Y3_LUT4AB/NN4BEG[11] Tile_X8Y3_LUT4AB/NN4BEG[12] Tile_X8Y3_LUT4AB/NN4BEG[13]
+ Tile_X8Y3_LUT4AB/NN4BEG[14] Tile_X8Y3_LUT4AB/NN4BEG[15] Tile_X8Y3_LUT4AB/NN4BEG[1]
+ Tile_X8Y3_LUT4AB/NN4BEG[2] Tile_X8Y3_LUT4AB/NN4BEG[3] Tile_X8Y3_LUT4AB/NN4BEG[4]
+ Tile_X8Y3_LUT4AB/NN4BEG[5] Tile_X8Y3_LUT4AB/NN4BEG[6] Tile_X8Y3_LUT4AB/NN4BEG[7]
+ Tile_X8Y3_LUT4AB/NN4BEG[8] Tile_X8Y3_LUT4AB/NN4BEG[9] Tile_X8Y4_LUT4AB/NN4BEG[0]
+ Tile_X8Y4_LUT4AB/NN4BEG[10] Tile_X8Y4_LUT4AB/NN4BEG[11] Tile_X8Y4_LUT4AB/NN4BEG[12]
+ Tile_X8Y4_LUT4AB/NN4BEG[13] Tile_X8Y4_LUT4AB/NN4BEG[14] Tile_X8Y4_LUT4AB/NN4BEG[15]
+ Tile_X8Y4_LUT4AB/NN4BEG[1] Tile_X8Y4_LUT4AB/NN4BEG[2] Tile_X8Y4_LUT4AB/NN4BEG[3]
+ Tile_X8Y4_LUT4AB/NN4BEG[4] Tile_X8Y4_LUT4AB/NN4BEG[5] Tile_X8Y4_LUT4AB/NN4BEG[6]
+ Tile_X8Y4_LUT4AB/NN4BEG[7] Tile_X8Y4_LUT4AB/NN4BEG[8] Tile_X8Y4_LUT4AB/NN4BEG[9]
+ Tile_X8Y4_LUT4AB/S1END[0] Tile_X8Y4_LUT4AB/S1END[1] Tile_X8Y4_LUT4AB/S1END[2] Tile_X8Y4_LUT4AB/S1END[3]
+ Tile_X8Y3_LUT4AB/S1END[0] Tile_X8Y3_LUT4AB/S1END[1] Tile_X8Y3_LUT4AB/S1END[2] Tile_X8Y3_LUT4AB/S1END[3]
+ Tile_X8Y4_LUT4AB/S2MID[0] Tile_X8Y4_LUT4AB/S2MID[1] Tile_X8Y4_LUT4AB/S2MID[2] Tile_X8Y4_LUT4AB/S2MID[3]
+ Tile_X8Y4_LUT4AB/S2MID[4] Tile_X8Y4_LUT4AB/S2MID[5] Tile_X8Y4_LUT4AB/S2MID[6] Tile_X8Y4_LUT4AB/S2MID[7]
+ Tile_X8Y4_LUT4AB/S2END[0] Tile_X8Y4_LUT4AB/S2END[1] Tile_X8Y4_LUT4AB/S2END[2] Tile_X8Y4_LUT4AB/S2END[3]
+ Tile_X8Y4_LUT4AB/S2END[4] Tile_X8Y4_LUT4AB/S2END[5] Tile_X8Y4_LUT4AB/S2END[6] Tile_X8Y4_LUT4AB/S2END[7]
+ Tile_X8Y3_LUT4AB/S2END[0] Tile_X8Y3_LUT4AB/S2END[1] Tile_X8Y3_LUT4AB/S2END[2] Tile_X8Y3_LUT4AB/S2END[3]
+ Tile_X8Y3_LUT4AB/S2END[4] Tile_X8Y3_LUT4AB/S2END[5] Tile_X8Y3_LUT4AB/S2END[6] Tile_X8Y3_LUT4AB/S2END[7]
+ Tile_X8Y3_LUT4AB/S2MID[0] Tile_X8Y3_LUT4AB/S2MID[1] Tile_X8Y3_LUT4AB/S2MID[2] Tile_X8Y3_LUT4AB/S2MID[3]
+ Tile_X8Y3_LUT4AB/S2MID[4] Tile_X8Y3_LUT4AB/S2MID[5] Tile_X8Y3_LUT4AB/S2MID[6] Tile_X8Y3_LUT4AB/S2MID[7]
+ Tile_X8Y4_LUT4AB/S4END[0] Tile_X8Y4_LUT4AB/S4END[10] Tile_X8Y4_LUT4AB/S4END[11]
+ Tile_X8Y4_LUT4AB/S4END[12] Tile_X8Y4_LUT4AB/S4END[13] Tile_X8Y4_LUT4AB/S4END[14]
+ Tile_X8Y4_LUT4AB/S4END[15] Tile_X8Y4_LUT4AB/S4END[1] Tile_X8Y4_LUT4AB/S4END[2] Tile_X8Y4_LUT4AB/S4END[3]
+ Tile_X8Y4_LUT4AB/S4END[4] Tile_X8Y4_LUT4AB/S4END[5] Tile_X8Y4_LUT4AB/S4END[6] Tile_X8Y4_LUT4AB/S4END[7]
+ Tile_X8Y4_LUT4AB/S4END[8] Tile_X8Y4_LUT4AB/S4END[9] Tile_X8Y3_LUT4AB/S4END[0] Tile_X8Y3_LUT4AB/S4END[10]
+ Tile_X8Y3_LUT4AB/S4END[11] Tile_X8Y3_LUT4AB/S4END[12] Tile_X8Y3_LUT4AB/S4END[13]
+ Tile_X8Y3_LUT4AB/S4END[14] Tile_X8Y3_LUT4AB/S4END[15] Tile_X8Y3_LUT4AB/S4END[1]
+ Tile_X8Y3_LUT4AB/S4END[2] Tile_X8Y3_LUT4AB/S4END[3] Tile_X8Y3_LUT4AB/S4END[4] Tile_X8Y3_LUT4AB/S4END[5]
+ Tile_X8Y3_LUT4AB/S4END[6] Tile_X8Y3_LUT4AB/S4END[7] Tile_X8Y3_LUT4AB/S4END[8] Tile_X8Y3_LUT4AB/S4END[9]
+ Tile_X8Y4_LUT4AB/SS4END[0] Tile_X8Y4_LUT4AB/SS4END[10] Tile_X8Y4_LUT4AB/SS4END[11]
+ Tile_X8Y4_LUT4AB/SS4END[12] Tile_X8Y4_LUT4AB/SS4END[13] Tile_X8Y4_LUT4AB/SS4END[14]
+ Tile_X8Y4_LUT4AB/SS4END[15] Tile_X8Y4_LUT4AB/SS4END[1] Tile_X8Y4_LUT4AB/SS4END[2]
+ Tile_X8Y4_LUT4AB/SS4END[3] Tile_X8Y4_LUT4AB/SS4END[4] Tile_X8Y4_LUT4AB/SS4END[5]
+ Tile_X8Y4_LUT4AB/SS4END[6] Tile_X8Y4_LUT4AB/SS4END[7] Tile_X8Y4_LUT4AB/SS4END[8]
+ Tile_X8Y4_LUT4AB/SS4END[9] Tile_X8Y3_LUT4AB/SS4END[0] Tile_X8Y3_LUT4AB/SS4END[10]
+ Tile_X8Y3_LUT4AB/SS4END[11] Tile_X8Y3_LUT4AB/SS4END[12] Tile_X8Y3_LUT4AB/SS4END[13]
+ Tile_X8Y3_LUT4AB/SS4END[14] Tile_X8Y3_LUT4AB/SS4END[15] Tile_X8Y3_LUT4AB/SS4END[1]
+ Tile_X8Y3_LUT4AB/SS4END[2] Tile_X8Y3_LUT4AB/SS4END[3] Tile_X8Y3_LUT4AB/SS4END[4]
+ Tile_X8Y3_LUT4AB/SS4END[5] Tile_X8Y3_LUT4AB/SS4END[6] Tile_X8Y3_LUT4AB/SS4END[7]
+ Tile_X8Y3_LUT4AB/SS4END[8] Tile_X8Y3_LUT4AB/SS4END[9] Tile_X8Y3_LUT4AB/UserCLK Tile_X8Y2_LUT4AB/UserCLK
+ VGND VPWR Tile_X8Y3_LUT4AB/W1BEG[0] Tile_X8Y3_LUT4AB/W1BEG[1] Tile_X8Y3_LUT4AB/W1BEG[2]
+ Tile_X8Y3_LUT4AB/W1BEG[3] Tile_X9Y3_LUT4AB/W1BEG[0] Tile_X9Y3_LUT4AB/W1BEG[1] Tile_X9Y3_LUT4AB/W1BEG[2]
+ Tile_X9Y3_LUT4AB/W1BEG[3] Tile_X8Y3_LUT4AB/W2BEG[0] Tile_X8Y3_LUT4AB/W2BEG[1] Tile_X8Y3_LUT4AB/W2BEG[2]
+ Tile_X8Y3_LUT4AB/W2BEG[3] Tile_X8Y3_LUT4AB/W2BEG[4] Tile_X8Y3_LUT4AB/W2BEG[5] Tile_X8Y3_LUT4AB/W2BEG[6]
+ Tile_X8Y3_LUT4AB/W2BEG[7] Tile_X8Y3_LUT4AB/W2BEGb[0] Tile_X8Y3_LUT4AB/W2BEGb[1]
+ Tile_X8Y3_LUT4AB/W2BEGb[2] Tile_X8Y3_LUT4AB/W2BEGb[3] Tile_X8Y3_LUT4AB/W2BEGb[4]
+ Tile_X8Y3_LUT4AB/W2BEGb[5] Tile_X8Y3_LUT4AB/W2BEGb[6] Tile_X8Y3_LUT4AB/W2BEGb[7]
+ Tile_X8Y3_LUT4AB/W2END[0] Tile_X8Y3_LUT4AB/W2END[1] Tile_X8Y3_LUT4AB/W2END[2] Tile_X8Y3_LUT4AB/W2END[3]
+ Tile_X8Y3_LUT4AB/W2END[4] Tile_X8Y3_LUT4AB/W2END[5] Tile_X8Y3_LUT4AB/W2END[6] Tile_X8Y3_LUT4AB/W2END[7]
+ Tile_X9Y3_LUT4AB/W2BEG[0] Tile_X9Y3_LUT4AB/W2BEG[1] Tile_X9Y3_LUT4AB/W2BEG[2] Tile_X9Y3_LUT4AB/W2BEG[3]
+ Tile_X9Y3_LUT4AB/W2BEG[4] Tile_X9Y3_LUT4AB/W2BEG[5] Tile_X9Y3_LUT4AB/W2BEG[6] Tile_X9Y3_LUT4AB/W2BEG[7]
+ Tile_X8Y3_LUT4AB/W6BEG[0] Tile_X8Y3_LUT4AB/W6BEG[10] Tile_X8Y3_LUT4AB/W6BEG[11]
+ Tile_X8Y3_LUT4AB/W6BEG[1] Tile_X8Y3_LUT4AB/W6BEG[2] Tile_X8Y3_LUT4AB/W6BEG[3] Tile_X8Y3_LUT4AB/W6BEG[4]
+ Tile_X8Y3_LUT4AB/W6BEG[5] Tile_X8Y3_LUT4AB/W6BEG[6] Tile_X8Y3_LUT4AB/W6BEG[7] Tile_X8Y3_LUT4AB/W6BEG[8]
+ Tile_X8Y3_LUT4AB/W6BEG[9] Tile_X9Y3_LUT4AB/W6BEG[0] Tile_X9Y3_LUT4AB/W6BEG[10] Tile_X9Y3_LUT4AB/W6BEG[11]
+ Tile_X9Y3_LUT4AB/W6BEG[1] Tile_X9Y3_LUT4AB/W6BEG[2] Tile_X9Y3_LUT4AB/W6BEG[3] Tile_X9Y3_LUT4AB/W6BEG[4]
+ Tile_X9Y3_LUT4AB/W6BEG[5] Tile_X9Y3_LUT4AB/W6BEG[6] Tile_X9Y3_LUT4AB/W6BEG[7] Tile_X9Y3_LUT4AB/W6BEG[8]
+ Tile_X9Y3_LUT4AB/W6BEG[9] Tile_X8Y3_LUT4AB/WW4BEG[0] Tile_X8Y3_LUT4AB/WW4BEG[10]
+ Tile_X8Y3_LUT4AB/WW4BEG[11] Tile_X8Y3_LUT4AB/WW4BEG[12] Tile_X8Y3_LUT4AB/WW4BEG[13]
+ Tile_X8Y3_LUT4AB/WW4BEG[14] Tile_X8Y3_LUT4AB/WW4BEG[15] Tile_X8Y3_LUT4AB/WW4BEG[1]
+ Tile_X8Y3_LUT4AB/WW4BEG[2] Tile_X8Y3_LUT4AB/WW4BEG[3] Tile_X8Y3_LUT4AB/WW4BEG[4]
+ Tile_X8Y3_LUT4AB/WW4BEG[5] Tile_X8Y3_LUT4AB/WW4BEG[6] Tile_X8Y3_LUT4AB/WW4BEG[7]
+ Tile_X8Y3_LUT4AB/WW4BEG[8] Tile_X8Y3_LUT4AB/WW4BEG[9] Tile_X9Y3_LUT4AB/WW4BEG[0]
+ Tile_X9Y3_LUT4AB/WW4BEG[10] Tile_X9Y3_LUT4AB/WW4BEG[11] Tile_X9Y3_LUT4AB/WW4BEG[12]
+ Tile_X9Y3_LUT4AB/WW4BEG[13] Tile_X9Y3_LUT4AB/WW4BEG[14] Tile_X9Y3_LUT4AB/WW4BEG[15]
+ Tile_X9Y3_LUT4AB/WW4BEG[1] Tile_X9Y3_LUT4AB/WW4BEG[2] Tile_X9Y3_LUT4AB/WW4BEG[3]
+ Tile_X9Y3_LUT4AB/WW4BEG[4] Tile_X9Y3_LUT4AB/WW4BEG[5] Tile_X9Y3_LUT4AB/WW4BEG[6]
+ Tile_X9Y3_LUT4AB/WW4BEG[7] Tile_X9Y3_LUT4AB/WW4BEG[8] Tile_X9Y3_LUT4AB/WW4BEG[9]
+ LUT4AB
XTile_X3Y13_LUT4AB Tile_X3Y14_LUT4AB/Co Tile_X3Y13_LUT4AB/Co Tile_X3Y13_LUT4AB/E1BEG[0]
+ Tile_X3Y13_LUT4AB/E1BEG[1] Tile_X3Y13_LUT4AB/E1BEG[2] Tile_X3Y13_LUT4AB/E1BEG[3]
+ Tile_X3Y13_LUT4AB/E1END[0] Tile_X3Y13_LUT4AB/E1END[1] Tile_X3Y13_LUT4AB/E1END[2]
+ Tile_X3Y13_LUT4AB/E1END[3] Tile_X3Y13_LUT4AB/E2BEG[0] Tile_X3Y13_LUT4AB/E2BEG[1]
+ Tile_X3Y13_LUT4AB/E2BEG[2] Tile_X3Y13_LUT4AB/E2BEG[3] Tile_X3Y13_LUT4AB/E2BEG[4]
+ Tile_X3Y13_LUT4AB/E2BEG[5] Tile_X3Y13_LUT4AB/E2BEG[6] Tile_X3Y13_LUT4AB/E2BEG[7]
+ Tile_X4Y13_RegFile/E2END[0] Tile_X4Y13_RegFile/E2END[1] Tile_X4Y13_RegFile/E2END[2]
+ Tile_X4Y13_RegFile/E2END[3] Tile_X4Y13_RegFile/E2END[4] Tile_X4Y13_RegFile/E2END[5]
+ Tile_X4Y13_RegFile/E2END[6] Tile_X4Y13_RegFile/E2END[7] Tile_X3Y13_LUT4AB/E2END[0]
+ Tile_X3Y13_LUT4AB/E2END[1] Tile_X3Y13_LUT4AB/E2END[2] Tile_X3Y13_LUT4AB/E2END[3]
+ Tile_X3Y13_LUT4AB/E2END[4] Tile_X3Y13_LUT4AB/E2END[5] Tile_X3Y13_LUT4AB/E2END[6]
+ Tile_X3Y13_LUT4AB/E2END[7] Tile_X3Y13_LUT4AB/E2MID[0] Tile_X3Y13_LUT4AB/E2MID[1]
+ Tile_X3Y13_LUT4AB/E2MID[2] Tile_X3Y13_LUT4AB/E2MID[3] Tile_X3Y13_LUT4AB/E2MID[4]
+ Tile_X3Y13_LUT4AB/E2MID[5] Tile_X3Y13_LUT4AB/E2MID[6] Tile_X3Y13_LUT4AB/E2MID[7]
+ Tile_X3Y13_LUT4AB/E6BEG[0] Tile_X3Y13_LUT4AB/E6BEG[10] Tile_X3Y13_LUT4AB/E6BEG[11]
+ Tile_X3Y13_LUT4AB/E6BEG[1] Tile_X3Y13_LUT4AB/E6BEG[2] Tile_X3Y13_LUT4AB/E6BEG[3]
+ Tile_X3Y13_LUT4AB/E6BEG[4] Tile_X3Y13_LUT4AB/E6BEG[5] Tile_X3Y13_LUT4AB/E6BEG[6]
+ Tile_X3Y13_LUT4AB/E6BEG[7] Tile_X3Y13_LUT4AB/E6BEG[8] Tile_X3Y13_LUT4AB/E6BEG[9]
+ Tile_X3Y13_LUT4AB/E6END[0] Tile_X3Y13_LUT4AB/E6END[10] Tile_X3Y13_LUT4AB/E6END[11]
+ Tile_X3Y13_LUT4AB/E6END[1] Tile_X3Y13_LUT4AB/E6END[2] Tile_X3Y13_LUT4AB/E6END[3]
+ Tile_X3Y13_LUT4AB/E6END[4] Tile_X3Y13_LUT4AB/E6END[5] Tile_X3Y13_LUT4AB/E6END[6]
+ Tile_X3Y13_LUT4AB/E6END[7] Tile_X3Y13_LUT4AB/E6END[8] Tile_X3Y13_LUT4AB/E6END[9]
+ Tile_X3Y13_LUT4AB/EE4BEG[0] Tile_X3Y13_LUT4AB/EE4BEG[10] Tile_X3Y13_LUT4AB/EE4BEG[11]
+ Tile_X3Y13_LUT4AB/EE4BEG[12] Tile_X3Y13_LUT4AB/EE4BEG[13] Tile_X3Y13_LUT4AB/EE4BEG[14]
+ Tile_X3Y13_LUT4AB/EE4BEG[15] Tile_X3Y13_LUT4AB/EE4BEG[1] Tile_X3Y13_LUT4AB/EE4BEG[2]
+ Tile_X3Y13_LUT4AB/EE4BEG[3] Tile_X3Y13_LUT4AB/EE4BEG[4] Tile_X3Y13_LUT4AB/EE4BEG[5]
+ Tile_X3Y13_LUT4AB/EE4BEG[6] Tile_X3Y13_LUT4AB/EE4BEG[7] Tile_X3Y13_LUT4AB/EE4BEG[8]
+ Tile_X3Y13_LUT4AB/EE4BEG[9] Tile_X3Y13_LUT4AB/EE4END[0] Tile_X3Y13_LUT4AB/EE4END[10]
+ Tile_X3Y13_LUT4AB/EE4END[11] Tile_X3Y13_LUT4AB/EE4END[12] Tile_X3Y13_LUT4AB/EE4END[13]
+ Tile_X3Y13_LUT4AB/EE4END[14] Tile_X3Y13_LUT4AB/EE4END[15] Tile_X3Y13_LUT4AB/EE4END[1]
+ Tile_X3Y13_LUT4AB/EE4END[2] Tile_X3Y13_LUT4AB/EE4END[3] Tile_X3Y13_LUT4AB/EE4END[4]
+ Tile_X3Y13_LUT4AB/EE4END[5] Tile_X3Y13_LUT4AB/EE4END[6] Tile_X3Y13_LUT4AB/EE4END[7]
+ Tile_X3Y13_LUT4AB/EE4END[8] Tile_X3Y13_LUT4AB/EE4END[9] Tile_X3Y13_LUT4AB/FrameData[0]
+ Tile_X3Y13_LUT4AB/FrameData[10] Tile_X3Y13_LUT4AB/FrameData[11] Tile_X3Y13_LUT4AB/FrameData[12]
+ Tile_X3Y13_LUT4AB/FrameData[13] Tile_X3Y13_LUT4AB/FrameData[14] Tile_X3Y13_LUT4AB/FrameData[15]
+ Tile_X3Y13_LUT4AB/FrameData[16] Tile_X3Y13_LUT4AB/FrameData[17] Tile_X3Y13_LUT4AB/FrameData[18]
+ Tile_X3Y13_LUT4AB/FrameData[19] Tile_X3Y13_LUT4AB/FrameData[1] Tile_X3Y13_LUT4AB/FrameData[20]
+ Tile_X3Y13_LUT4AB/FrameData[21] Tile_X3Y13_LUT4AB/FrameData[22] Tile_X3Y13_LUT4AB/FrameData[23]
+ Tile_X3Y13_LUT4AB/FrameData[24] Tile_X3Y13_LUT4AB/FrameData[25] Tile_X3Y13_LUT4AB/FrameData[26]
+ Tile_X3Y13_LUT4AB/FrameData[27] Tile_X3Y13_LUT4AB/FrameData[28] Tile_X3Y13_LUT4AB/FrameData[29]
+ Tile_X3Y13_LUT4AB/FrameData[2] Tile_X3Y13_LUT4AB/FrameData[30] Tile_X3Y13_LUT4AB/FrameData[31]
+ Tile_X3Y13_LUT4AB/FrameData[3] Tile_X3Y13_LUT4AB/FrameData[4] Tile_X3Y13_LUT4AB/FrameData[5]
+ Tile_X3Y13_LUT4AB/FrameData[6] Tile_X3Y13_LUT4AB/FrameData[7] Tile_X3Y13_LUT4AB/FrameData[8]
+ Tile_X3Y13_LUT4AB/FrameData[9] Tile_X4Y13_RegFile/FrameData[0] Tile_X4Y13_RegFile/FrameData[10]
+ Tile_X4Y13_RegFile/FrameData[11] Tile_X4Y13_RegFile/FrameData[12] Tile_X4Y13_RegFile/FrameData[13]
+ Tile_X4Y13_RegFile/FrameData[14] Tile_X4Y13_RegFile/FrameData[15] Tile_X4Y13_RegFile/FrameData[16]
+ Tile_X4Y13_RegFile/FrameData[17] Tile_X4Y13_RegFile/FrameData[18] Tile_X4Y13_RegFile/FrameData[19]
+ Tile_X4Y13_RegFile/FrameData[1] Tile_X4Y13_RegFile/FrameData[20] Tile_X4Y13_RegFile/FrameData[21]
+ Tile_X4Y13_RegFile/FrameData[22] Tile_X4Y13_RegFile/FrameData[23] Tile_X4Y13_RegFile/FrameData[24]
+ Tile_X4Y13_RegFile/FrameData[25] Tile_X4Y13_RegFile/FrameData[26] Tile_X4Y13_RegFile/FrameData[27]
+ Tile_X4Y13_RegFile/FrameData[28] Tile_X4Y13_RegFile/FrameData[29] Tile_X4Y13_RegFile/FrameData[2]
+ Tile_X4Y13_RegFile/FrameData[30] Tile_X4Y13_RegFile/FrameData[31] Tile_X4Y13_RegFile/FrameData[3]
+ Tile_X4Y13_RegFile/FrameData[4] Tile_X4Y13_RegFile/FrameData[5] Tile_X4Y13_RegFile/FrameData[6]
+ Tile_X4Y13_RegFile/FrameData[7] Tile_X4Y13_RegFile/FrameData[8] Tile_X4Y13_RegFile/FrameData[9]
+ Tile_X3Y13_LUT4AB/FrameStrobe[0] Tile_X3Y13_LUT4AB/FrameStrobe[10] Tile_X3Y13_LUT4AB/FrameStrobe[11]
+ Tile_X3Y13_LUT4AB/FrameStrobe[12] Tile_X3Y13_LUT4AB/FrameStrobe[13] Tile_X3Y13_LUT4AB/FrameStrobe[14]
+ Tile_X3Y13_LUT4AB/FrameStrobe[15] Tile_X3Y13_LUT4AB/FrameStrobe[16] Tile_X3Y13_LUT4AB/FrameStrobe[17]
+ Tile_X3Y13_LUT4AB/FrameStrobe[18] Tile_X3Y13_LUT4AB/FrameStrobe[19] Tile_X3Y13_LUT4AB/FrameStrobe[1]
+ Tile_X3Y13_LUT4AB/FrameStrobe[2] Tile_X3Y13_LUT4AB/FrameStrobe[3] Tile_X3Y13_LUT4AB/FrameStrobe[4]
+ Tile_X3Y13_LUT4AB/FrameStrobe[5] Tile_X3Y13_LUT4AB/FrameStrobe[6] Tile_X3Y13_LUT4AB/FrameStrobe[7]
+ Tile_X3Y13_LUT4AB/FrameStrobe[8] Tile_X3Y13_LUT4AB/FrameStrobe[9] Tile_X3Y12_LUT4AB/FrameStrobe[0]
+ Tile_X3Y12_LUT4AB/FrameStrobe[10] Tile_X3Y12_LUT4AB/FrameStrobe[11] Tile_X3Y12_LUT4AB/FrameStrobe[12]
+ Tile_X3Y12_LUT4AB/FrameStrobe[13] Tile_X3Y12_LUT4AB/FrameStrobe[14] Tile_X3Y12_LUT4AB/FrameStrobe[15]
+ Tile_X3Y12_LUT4AB/FrameStrobe[16] Tile_X3Y12_LUT4AB/FrameStrobe[17] Tile_X3Y12_LUT4AB/FrameStrobe[18]
+ Tile_X3Y12_LUT4AB/FrameStrobe[19] Tile_X3Y12_LUT4AB/FrameStrobe[1] Tile_X3Y12_LUT4AB/FrameStrobe[2]
+ Tile_X3Y12_LUT4AB/FrameStrobe[3] Tile_X3Y12_LUT4AB/FrameStrobe[4] Tile_X3Y12_LUT4AB/FrameStrobe[5]
+ Tile_X3Y12_LUT4AB/FrameStrobe[6] Tile_X3Y12_LUT4AB/FrameStrobe[7] Tile_X3Y12_LUT4AB/FrameStrobe[8]
+ Tile_X3Y12_LUT4AB/FrameStrobe[9] Tile_X3Y13_LUT4AB/N1BEG[0] Tile_X3Y13_LUT4AB/N1BEG[1]
+ Tile_X3Y13_LUT4AB/N1BEG[2] Tile_X3Y13_LUT4AB/N1BEG[3] Tile_X3Y14_LUT4AB/N1BEG[0]
+ Tile_X3Y14_LUT4AB/N1BEG[1] Tile_X3Y14_LUT4AB/N1BEG[2] Tile_X3Y14_LUT4AB/N1BEG[3]
+ Tile_X3Y13_LUT4AB/N2BEG[0] Tile_X3Y13_LUT4AB/N2BEG[1] Tile_X3Y13_LUT4AB/N2BEG[2]
+ Tile_X3Y13_LUT4AB/N2BEG[3] Tile_X3Y13_LUT4AB/N2BEG[4] Tile_X3Y13_LUT4AB/N2BEG[5]
+ Tile_X3Y13_LUT4AB/N2BEG[6] Tile_X3Y13_LUT4AB/N2BEG[7] Tile_X3Y12_LUT4AB/N2END[0]
+ Tile_X3Y12_LUT4AB/N2END[1] Tile_X3Y12_LUT4AB/N2END[2] Tile_X3Y12_LUT4AB/N2END[3]
+ Tile_X3Y12_LUT4AB/N2END[4] Tile_X3Y12_LUT4AB/N2END[5] Tile_X3Y12_LUT4AB/N2END[6]
+ Tile_X3Y12_LUT4AB/N2END[7] Tile_X3Y13_LUT4AB/N2END[0] Tile_X3Y13_LUT4AB/N2END[1]
+ Tile_X3Y13_LUT4AB/N2END[2] Tile_X3Y13_LUT4AB/N2END[3] Tile_X3Y13_LUT4AB/N2END[4]
+ Tile_X3Y13_LUT4AB/N2END[5] Tile_X3Y13_LUT4AB/N2END[6] Tile_X3Y13_LUT4AB/N2END[7]
+ Tile_X3Y14_LUT4AB/N2BEG[0] Tile_X3Y14_LUT4AB/N2BEG[1] Tile_X3Y14_LUT4AB/N2BEG[2]
+ Tile_X3Y14_LUT4AB/N2BEG[3] Tile_X3Y14_LUT4AB/N2BEG[4] Tile_X3Y14_LUT4AB/N2BEG[5]
+ Tile_X3Y14_LUT4AB/N2BEG[6] Tile_X3Y14_LUT4AB/N2BEG[7] Tile_X3Y13_LUT4AB/N4BEG[0]
+ Tile_X3Y13_LUT4AB/N4BEG[10] Tile_X3Y13_LUT4AB/N4BEG[11] Tile_X3Y13_LUT4AB/N4BEG[12]
+ Tile_X3Y13_LUT4AB/N4BEG[13] Tile_X3Y13_LUT4AB/N4BEG[14] Tile_X3Y13_LUT4AB/N4BEG[15]
+ Tile_X3Y13_LUT4AB/N4BEG[1] Tile_X3Y13_LUT4AB/N4BEG[2] Tile_X3Y13_LUT4AB/N4BEG[3]
+ Tile_X3Y13_LUT4AB/N4BEG[4] Tile_X3Y13_LUT4AB/N4BEG[5] Tile_X3Y13_LUT4AB/N4BEG[6]
+ Tile_X3Y13_LUT4AB/N4BEG[7] Tile_X3Y13_LUT4AB/N4BEG[8] Tile_X3Y13_LUT4AB/N4BEG[9]
+ Tile_X3Y14_LUT4AB/N4BEG[0] Tile_X3Y14_LUT4AB/N4BEG[10] Tile_X3Y14_LUT4AB/N4BEG[11]
+ Tile_X3Y14_LUT4AB/N4BEG[12] Tile_X3Y14_LUT4AB/N4BEG[13] Tile_X3Y14_LUT4AB/N4BEG[14]
+ Tile_X3Y14_LUT4AB/N4BEG[15] Tile_X3Y14_LUT4AB/N4BEG[1] Tile_X3Y14_LUT4AB/N4BEG[2]
+ Tile_X3Y14_LUT4AB/N4BEG[3] Tile_X3Y14_LUT4AB/N4BEG[4] Tile_X3Y14_LUT4AB/N4BEG[5]
+ Tile_X3Y14_LUT4AB/N4BEG[6] Tile_X3Y14_LUT4AB/N4BEG[7] Tile_X3Y14_LUT4AB/N4BEG[8]
+ Tile_X3Y14_LUT4AB/N4BEG[9] Tile_X3Y13_LUT4AB/NN4BEG[0] Tile_X3Y13_LUT4AB/NN4BEG[10]
+ Tile_X3Y13_LUT4AB/NN4BEG[11] Tile_X3Y13_LUT4AB/NN4BEG[12] Tile_X3Y13_LUT4AB/NN4BEG[13]
+ Tile_X3Y13_LUT4AB/NN4BEG[14] Tile_X3Y13_LUT4AB/NN4BEG[15] Tile_X3Y13_LUT4AB/NN4BEG[1]
+ Tile_X3Y13_LUT4AB/NN4BEG[2] Tile_X3Y13_LUT4AB/NN4BEG[3] Tile_X3Y13_LUT4AB/NN4BEG[4]
+ Tile_X3Y13_LUT4AB/NN4BEG[5] Tile_X3Y13_LUT4AB/NN4BEG[6] Tile_X3Y13_LUT4AB/NN4BEG[7]
+ Tile_X3Y13_LUT4AB/NN4BEG[8] Tile_X3Y13_LUT4AB/NN4BEG[9] Tile_X3Y14_LUT4AB/NN4BEG[0]
+ Tile_X3Y14_LUT4AB/NN4BEG[10] Tile_X3Y14_LUT4AB/NN4BEG[11] Tile_X3Y14_LUT4AB/NN4BEG[12]
+ Tile_X3Y14_LUT4AB/NN4BEG[13] Tile_X3Y14_LUT4AB/NN4BEG[14] Tile_X3Y14_LUT4AB/NN4BEG[15]
+ Tile_X3Y14_LUT4AB/NN4BEG[1] Tile_X3Y14_LUT4AB/NN4BEG[2] Tile_X3Y14_LUT4AB/NN4BEG[3]
+ Tile_X3Y14_LUT4AB/NN4BEG[4] Tile_X3Y14_LUT4AB/NN4BEG[5] Tile_X3Y14_LUT4AB/NN4BEG[6]
+ Tile_X3Y14_LUT4AB/NN4BEG[7] Tile_X3Y14_LUT4AB/NN4BEG[8] Tile_X3Y14_LUT4AB/NN4BEG[9]
+ Tile_X3Y14_LUT4AB/S1END[0] Tile_X3Y14_LUT4AB/S1END[1] Tile_X3Y14_LUT4AB/S1END[2]
+ Tile_X3Y14_LUT4AB/S1END[3] Tile_X3Y13_LUT4AB/S1END[0] Tile_X3Y13_LUT4AB/S1END[1]
+ Tile_X3Y13_LUT4AB/S1END[2] Tile_X3Y13_LUT4AB/S1END[3] Tile_X3Y14_LUT4AB/S2MID[0]
+ Tile_X3Y14_LUT4AB/S2MID[1] Tile_X3Y14_LUT4AB/S2MID[2] Tile_X3Y14_LUT4AB/S2MID[3]
+ Tile_X3Y14_LUT4AB/S2MID[4] Tile_X3Y14_LUT4AB/S2MID[5] Tile_X3Y14_LUT4AB/S2MID[6]
+ Tile_X3Y14_LUT4AB/S2MID[7] Tile_X3Y14_LUT4AB/S2END[0] Tile_X3Y14_LUT4AB/S2END[1]
+ Tile_X3Y14_LUT4AB/S2END[2] Tile_X3Y14_LUT4AB/S2END[3] Tile_X3Y14_LUT4AB/S2END[4]
+ Tile_X3Y14_LUT4AB/S2END[5] Tile_X3Y14_LUT4AB/S2END[6] Tile_X3Y14_LUT4AB/S2END[7]
+ Tile_X3Y13_LUT4AB/S2END[0] Tile_X3Y13_LUT4AB/S2END[1] Tile_X3Y13_LUT4AB/S2END[2]
+ Tile_X3Y13_LUT4AB/S2END[3] Tile_X3Y13_LUT4AB/S2END[4] Tile_X3Y13_LUT4AB/S2END[5]
+ Tile_X3Y13_LUT4AB/S2END[6] Tile_X3Y13_LUT4AB/S2END[7] Tile_X3Y13_LUT4AB/S2MID[0]
+ Tile_X3Y13_LUT4AB/S2MID[1] Tile_X3Y13_LUT4AB/S2MID[2] Tile_X3Y13_LUT4AB/S2MID[3]
+ Tile_X3Y13_LUT4AB/S2MID[4] Tile_X3Y13_LUT4AB/S2MID[5] Tile_X3Y13_LUT4AB/S2MID[6]
+ Tile_X3Y13_LUT4AB/S2MID[7] Tile_X3Y14_LUT4AB/S4END[0] Tile_X3Y14_LUT4AB/S4END[10]
+ Tile_X3Y14_LUT4AB/S4END[11] Tile_X3Y14_LUT4AB/S4END[12] Tile_X3Y14_LUT4AB/S4END[13]
+ Tile_X3Y14_LUT4AB/S4END[14] Tile_X3Y14_LUT4AB/S4END[15] Tile_X3Y14_LUT4AB/S4END[1]
+ Tile_X3Y14_LUT4AB/S4END[2] Tile_X3Y14_LUT4AB/S4END[3] Tile_X3Y14_LUT4AB/S4END[4]
+ Tile_X3Y14_LUT4AB/S4END[5] Tile_X3Y14_LUT4AB/S4END[6] Tile_X3Y14_LUT4AB/S4END[7]
+ Tile_X3Y14_LUT4AB/S4END[8] Tile_X3Y14_LUT4AB/S4END[9] Tile_X3Y13_LUT4AB/S4END[0]
+ Tile_X3Y13_LUT4AB/S4END[10] Tile_X3Y13_LUT4AB/S4END[11] Tile_X3Y13_LUT4AB/S4END[12]
+ Tile_X3Y13_LUT4AB/S4END[13] Tile_X3Y13_LUT4AB/S4END[14] Tile_X3Y13_LUT4AB/S4END[15]
+ Tile_X3Y13_LUT4AB/S4END[1] Tile_X3Y13_LUT4AB/S4END[2] Tile_X3Y13_LUT4AB/S4END[3]
+ Tile_X3Y13_LUT4AB/S4END[4] Tile_X3Y13_LUT4AB/S4END[5] Tile_X3Y13_LUT4AB/S4END[6]
+ Tile_X3Y13_LUT4AB/S4END[7] Tile_X3Y13_LUT4AB/S4END[8] Tile_X3Y13_LUT4AB/S4END[9]
+ Tile_X3Y14_LUT4AB/SS4END[0] Tile_X3Y14_LUT4AB/SS4END[10] Tile_X3Y14_LUT4AB/SS4END[11]
+ Tile_X3Y14_LUT4AB/SS4END[12] Tile_X3Y14_LUT4AB/SS4END[13] Tile_X3Y14_LUT4AB/SS4END[14]
+ Tile_X3Y14_LUT4AB/SS4END[15] Tile_X3Y14_LUT4AB/SS4END[1] Tile_X3Y14_LUT4AB/SS4END[2]
+ Tile_X3Y14_LUT4AB/SS4END[3] Tile_X3Y14_LUT4AB/SS4END[4] Tile_X3Y14_LUT4AB/SS4END[5]
+ Tile_X3Y14_LUT4AB/SS4END[6] Tile_X3Y14_LUT4AB/SS4END[7] Tile_X3Y14_LUT4AB/SS4END[8]
+ Tile_X3Y14_LUT4AB/SS4END[9] Tile_X3Y13_LUT4AB/SS4END[0] Tile_X3Y13_LUT4AB/SS4END[10]
+ Tile_X3Y13_LUT4AB/SS4END[11] Tile_X3Y13_LUT4AB/SS4END[12] Tile_X3Y13_LUT4AB/SS4END[13]
+ Tile_X3Y13_LUT4AB/SS4END[14] Tile_X3Y13_LUT4AB/SS4END[15] Tile_X3Y13_LUT4AB/SS4END[1]
+ Tile_X3Y13_LUT4AB/SS4END[2] Tile_X3Y13_LUT4AB/SS4END[3] Tile_X3Y13_LUT4AB/SS4END[4]
+ Tile_X3Y13_LUT4AB/SS4END[5] Tile_X3Y13_LUT4AB/SS4END[6] Tile_X3Y13_LUT4AB/SS4END[7]
+ Tile_X3Y13_LUT4AB/SS4END[8] Tile_X3Y13_LUT4AB/SS4END[9] Tile_X3Y13_LUT4AB/UserCLK
+ Tile_X3Y12_LUT4AB/UserCLK VGND VPWR Tile_X3Y13_LUT4AB/W1BEG[0] Tile_X3Y13_LUT4AB/W1BEG[1]
+ Tile_X3Y13_LUT4AB/W1BEG[2] Tile_X3Y13_LUT4AB/W1BEG[3] Tile_X3Y13_LUT4AB/W1END[0]
+ Tile_X3Y13_LUT4AB/W1END[1] Tile_X3Y13_LUT4AB/W1END[2] Tile_X3Y13_LUT4AB/W1END[3]
+ Tile_X3Y13_LUT4AB/W2BEG[0] Tile_X3Y13_LUT4AB/W2BEG[1] Tile_X3Y13_LUT4AB/W2BEG[2]
+ Tile_X3Y13_LUT4AB/W2BEG[3] Tile_X3Y13_LUT4AB/W2BEG[4] Tile_X3Y13_LUT4AB/W2BEG[5]
+ Tile_X3Y13_LUT4AB/W2BEG[6] Tile_X3Y13_LUT4AB/W2BEG[7] Tile_X2Y13_LUT4AB/W2END[0]
+ Tile_X2Y13_LUT4AB/W2END[1] Tile_X2Y13_LUT4AB/W2END[2] Tile_X2Y13_LUT4AB/W2END[3]
+ Tile_X2Y13_LUT4AB/W2END[4] Tile_X2Y13_LUT4AB/W2END[5] Tile_X2Y13_LUT4AB/W2END[6]
+ Tile_X2Y13_LUT4AB/W2END[7] Tile_X3Y13_LUT4AB/W2END[0] Tile_X3Y13_LUT4AB/W2END[1]
+ Tile_X3Y13_LUT4AB/W2END[2] Tile_X3Y13_LUT4AB/W2END[3] Tile_X3Y13_LUT4AB/W2END[4]
+ Tile_X3Y13_LUT4AB/W2END[5] Tile_X3Y13_LUT4AB/W2END[6] Tile_X3Y13_LUT4AB/W2END[7]
+ Tile_X3Y13_LUT4AB/W2MID[0] Tile_X3Y13_LUT4AB/W2MID[1] Tile_X3Y13_LUT4AB/W2MID[2]
+ Tile_X3Y13_LUT4AB/W2MID[3] Tile_X3Y13_LUT4AB/W2MID[4] Tile_X3Y13_LUT4AB/W2MID[5]
+ Tile_X3Y13_LUT4AB/W2MID[6] Tile_X3Y13_LUT4AB/W2MID[7] Tile_X3Y13_LUT4AB/W6BEG[0]
+ Tile_X3Y13_LUT4AB/W6BEG[10] Tile_X3Y13_LUT4AB/W6BEG[11] Tile_X3Y13_LUT4AB/W6BEG[1]
+ Tile_X3Y13_LUT4AB/W6BEG[2] Tile_X3Y13_LUT4AB/W6BEG[3] Tile_X3Y13_LUT4AB/W6BEG[4]
+ Tile_X3Y13_LUT4AB/W6BEG[5] Tile_X3Y13_LUT4AB/W6BEG[6] Tile_X3Y13_LUT4AB/W6BEG[7]
+ Tile_X3Y13_LUT4AB/W6BEG[8] Tile_X3Y13_LUT4AB/W6BEG[9] Tile_X3Y13_LUT4AB/W6END[0]
+ Tile_X3Y13_LUT4AB/W6END[10] Tile_X3Y13_LUT4AB/W6END[11] Tile_X3Y13_LUT4AB/W6END[1]
+ Tile_X3Y13_LUT4AB/W6END[2] Tile_X3Y13_LUT4AB/W6END[3] Tile_X3Y13_LUT4AB/W6END[4]
+ Tile_X3Y13_LUT4AB/W6END[5] Tile_X3Y13_LUT4AB/W6END[6] Tile_X3Y13_LUT4AB/W6END[7]
+ Tile_X3Y13_LUT4AB/W6END[8] Tile_X3Y13_LUT4AB/W6END[9] Tile_X3Y13_LUT4AB/WW4BEG[0]
+ Tile_X3Y13_LUT4AB/WW4BEG[10] Tile_X3Y13_LUT4AB/WW4BEG[11] Tile_X3Y13_LUT4AB/WW4BEG[12]
+ Tile_X3Y13_LUT4AB/WW4BEG[13] Tile_X3Y13_LUT4AB/WW4BEG[14] Tile_X3Y13_LUT4AB/WW4BEG[15]
+ Tile_X3Y13_LUT4AB/WW4BEG[1] Tile_X3Y13_LUT4AB/WW4BEG[2] Tile_X3Y13_LUT4AB/WW4BEG[3]
+ Tile_X3Y13_LUT4AB/WW4BEG[4] Tile_X3Y13_LUT4AB/WW4BEG[5] Tile_X3Y13_LUT4AB/WW4BEG[6]
+ Tile_X3Y13_LUT4AB/WW4BEG[7] Tile_X3Y13_LUT4AB/WW4BEG[8] Tile_X3Y13_LUT4AB/WW4BEG[9]
+ Tile_X3Y13_LUT4AB/WW4END[0] Tile_X3Y13_LUT4AB/WW4END[10] Tile_X3Y13_LUT4AB/WW4END[11]
+ Tile_X3Y13_LUT4AB/WW4END[12] Tile_X3Y13_LUT4AB/WW4END[13] Tile_X3Y13_LUT4AB/WW4END[14]
+ Tile_X3Y13_LUT4AB/WW4END[15] Tile_X3Y13_LUT4AB/WW4END[1] Tile_X3Y13_LUT4AB/WW4END[2]
+ Tile_X3Y13_LUT4AB/WW4END[3] Tile_X3Y13_LUT4AB/WW4END[4] Tile_X3Y13_LUT4AB/WW4END[5]
+ Tile_X3Y13_LUT4AB/WW4END[6] Tile_X3Y13_LUT4AB/WW4END[7] Tile_X3Y13_LUT4AB/WW4END[8]
+ Tile_X3Y13_LUT4AB/WW4END[9] LUT4AB
XTile_X9Y10_LUT4AB Tile_X9Y11_LUT4AB/Co Tile_X9Y9_LUT4AB/Ci Tile_X9Y10_LUT4AB/E1BEG[0]
+ Tile_X9Y10_LUT4AB/E1BEG[1] Tile_X9Y10_LUT4AB/E1BEG[2] Tile_X9Y10_LUT4AB/E1BEG[3]
+ Tile_X9Y10_LUT4AB/E1END[0] Tile_X9Y10_LUT4AB/E1END[1] Tile_X9Y10_LUT4AB/E1END[2]
+ Tile_X9Y10_LUT4AB/E1END[3] Tile_X9Y10_LUT4AB/E2BEG[0] Tile_X9Y10_LUT4AB/E2BEG[1]
+ Tile_X9Y10_LUT4AB/E2BEG[2] Tile_X9Y10_LUT4AB/E2BEG[3] Tile_X9Y10_LUT4AB/E2BEG[4]
+ Tile_X9Y10_LUT4AB/E2BEG[5] Tile_X9Y10_LUT4AB/E2BEG[6] Tile_X9Y10_LUT4AB/E2BEG[7]
+ Tile_X9Y10_LUT4AB/E2BEGb[0] Tile_X9Y10_LUT4AB/E2BEGb[1] Tile_X9Y10_LUT4AB/E2BEGb[2]
+ Tile_X9Y10_LUT4AB/E2BEGb[3] Tile_X9Y10_LUT4AB/E2BEGb[4] Tile_X9Y10_LUT4AB/E2BEGb[5]
+ Tile_X9Y10_LUT4AB/E2BEGb[6] Tile_X9Y10_LUT4AB/E2BEGb[7] Tile_X9Y10_LUT4AB/E2END[0]
+ Tile_X9Y10_LUT4AB/E2END[1] Tile_X9Y10_LUT4AB/E2END[2] Tile_X9Y10_LUT4AB/E2END[3]
+ Tile_X9Y10_LUT4AB/E2END[4] Tile_X9Y10_LUT4AB/E2END[5] Tile_X9Y10_LUT4AB/E2END[6]
+ Tile_X9Y10_LUT4AB/E2END[7] Tile_X9Y10_LUT4AB/E2MID[0] Tile_X9Y10_LUT4AB/E2MID[1]
+ Tile_X9Y10_LUT4AB/E2MID[2] Tile_X9Y10_LUT4AB/E2MID[3] Tile_X9Y10_LUT4AB/E2MID[4]
+ Tile_X9Y10_LUT4AB/E2MID[5] Tile_X9Y10_LUT4AB/E2MID[6] Tile_X9Y10_LUT4AB/E2MID[7]
+ Tile_X9Y10_LUT4AB/E6BEG[0] Tile_X9Y10_LUT4AB/E6BEG[10] Tile_X9Y10_LUT4AB/E6BEG[11]
+ Tile_X9Y10_LUT4AB/E6BEG[1] Tile_X9Y10_LUT4AB/E6BEG[2] Tile_X9Y10_LUT4AB/E6BEG[3]
+ Tile_X9Y10_LUT4AB/E6BEG[4] Tile_X9Y10_LUT4AB/E6BEG[5] Tile_X9Y10_LUT4AB/E6BEG[6]
+ Tile_X9Y10_LUT4AB/E6BEG[7] Tile_X9Y10_LUT4AB/E6BEG[8] Tile_X9Y10_LUT4AB/E6BEG[9]
+ Tile_X9Y10_LUT4AB/E6END[0] Tile_X9Y10_LUT4AB/E6END[10] Tile_X9Y10_LUT4AB/E6END[11]
+ Tile_X9Y10_LUT4AB/E6END[1] Tile_X9Y10_LUT4AB/E6END[2] Tile_X9Y10_LUT4AB/E6END[3]
+ Tile_X9Y10_LUT4AB/E6END[4] Tile_X9Y10_LUT4AB/E6END[5] Tile_X9Y10_LUT4AB/E6END[6]
+ Tile_X9Y10_LUT4AB/E6END[7] Tile_X9Y10_LUT4AB/E6END[8] Tile_X9Y10_LUT4AB/E6END[9]
+ Tile_X9Y10_LUT4AB/EE4BEG[0] Tile_X9Y10_LUT4AB/EE4BEG[10] Tile_X9Y10_LUT4AB/EE4BEG[11]
+ Tile_X9Y10_LUT4AB/EE4BEG[12] Tile_X9Y10_LUT4AB/EE4BEG[13] Tile_X9Y10_LUT4AB/EE4BEG[14]
+ Tile_X9Y10_LUT4AB/EE4BEG[15] Tile_X9Y10_LUT4AB/EE4BEG[1] Tile_X9Y10_LUT4AB/EE4BEG[2]
+ Tile_X9Y10_LUT4AB/EE4BEG[3] Tile_X9Y10_LUT4AB/EE4BEG[4] Tile_X9Y10_LUT4AB/EE4BEG[5]
+ Tile_X9Y10_LUT4AB/EE4BEG[6] Tile_X9Y10_LUT4AB/EE4BEG[7] Tile_X9Y10_LUT4AB/EE4BEG[8]
+ Tile_X9Y10_LUT4AB/EE4BEG[9] Tile_X9Y10_LUT4AB/EE4END[0] Tile_X9Y10_LUT4AB/EE4END[10]
+ Tile_X9Y10_LUT4AB/EE4END[11] Tile_X9Y10_LUT4AB/EE4END[12] Tile_X9Y10_LUT4AB/EE4END[13]
+ Tile_X9Y10_LUT4AB/EE4END[14] Tile_X9Y10_LUT4AB/EE4END[15] Tile_X9Y10_LUT4AB/EE4END[1]
+ Tile_X9Y10_LUT4AB/EE4END[2] Tile_X9Y10_LUT4AB/EE4END[3] Tile_X9Y10_LUT4AB/EE4END[4]
+ Tile_X9Y10_LUT4AB/EE4END[5] Tile_X9Y10_LUT4AB/EE4END[6] Tile_X9Y10_LUT4AB/EE4END[7]
+ Tile_X9Y10_LUT4AB/EE4END[8] Tile_X9Y10_LUT4AB/EE4END[9] Tile_X9Y10_LUT4AB/FrameData[0]
+ Tile_X9Y10_LUT4AB/FrameData[10] Tile_X9Y10_LUT4AB/FrameData[11] Tile_X9Y10_LUT4AB/FrameData[12]
+ Tile_X9Y10_LUT4AB/FrameData[13] Tile_X9Y10_LUT4AB/FrameData[14] Tile_X9Y10_LUT4AB/FrameData[15]
+ Tile_X9Y10_LUT4AB/FrameData[16] Tile_X9Y10_LUT4AB/FrameData[17] Tile_X9Y10_LUT4AB/FrameData[18]
+ Tile_X9Y10_LUT4AB/FrameData[19] Tile_X9Y10_LUT4AB/FrameData[1] Tile_X9Y10_LUT4AB/FrameData[20]
+ Tile_X9Y10_LUT4AB/FrameData[21] Tile_X9Y10_LUT4AB/FrameData[22] Tile_X9Y10_LUT4AB/FrameData[23]
+ Tile_X9Y10_LUT4AB/FrameData[24] Tile_X9Y10_LUT4AB/FrameData[25] Tile_X9Y10_LUT4AB/FrameData[26]
+ Tile_X9Y10_LUT4AB/FrameData[27] Tile_X9Y10_LUT4AB/FrameData[28] Tile_X9Y10_LUT4AB/FrameData[29]
+ Tile_X9Y10_LUT4AB/FrameData[2] Tile_X9Y10_LUT4AB/FrameData[30] Tile_X9Y10_LUT4AB/FrameData[31]
+ Tile_X9Y10_LUT4AB/FrameData[3] Tile_X9Y10_LUT4AB/FrameData[4] Tile_X9Y10_LUT4AB/FrameData[5]
+ Tile_X9Y10_LUT4AB/FrameData[6] Tile_X9Y10_LUT4AB/FrameData[7] Tile_X9Y10_LUT4AB/FrameData[8]
+ Tile_X9Y10_LUT4AB/FrameData[9] Tile_X9Y10_LUT4AB/FrameData_O[0] Tile_X9Y10_LUT4AB/FrameData_O[10]
+ Tile_X9Y10_LUT4AB/FrameData_O[11] Tile_X9Y10_LUT4AB/FrameData_O[12] Tile_X9Y10_LUT4AB/FrameData_O[13]
+ Tile_X9Y10_LUT4AB/FrameData_O[14] Tile_X9Y10_LUT4AB/FrameData_O[15] Tile_X9Y10_LUT4AB/FrameData_O[16]
+ Tile_X9Y10_LUT4AB/FrameData_O[17] Tile_X9Y10_LUT4AB/FrameData_O[18] Tile_X9Y10_LUT4AB/FrameData_O[19]
+ Tile_X9Y10_LUT4AB/FrameData_O[1] Tile_X9Y10_LUT4AB/FrameData_O[20] Tile_X9Y10_LUT4AB/FrameData_O[21]
+ Tile_X9Y10_LUT4AB/FrameData_O[22] Tile_X9Y10_LUT4AB/FrameData_O[23] Tile_X9Y10_LUT4AB/FrameData_O[24]
+ Tile_X9Y10_LUT4AB/FrameData_O[25] Tile_X9Y10_LUT4AB/FrameData_O[26] Tile_X9Y10_LUT4AB/FrameData_O[27]
+ Tile_X9Y10_LUT4AB/FrameData_O[28] Tile_X9Y10_LUT4AB/FrameData_O[29] Tile_X9Y10_LUT4AB/FrameData_O[2]
+ Tile_X9Y10_LUT4AB/FrameData_O[30] Tile_X9Y10_LUT4AB/FrameData_O[31] Tile_X9Y10_LUT4AB/FrameData_O[3]
+ Tile_X9Y10_LUT4AB/FrameData_O[4] Tile_X9Y10_LUT4AB/FrameData_O[5] Tile_X9Y10_LUT4AB/FrameData_O[6]
+ Tile_X9Y10_LUT4AB/FrameData_O[7] Tile_X9Y10_LUT4AB/FrameData_O[8] Tile_X9Y10_LUT4AB/FrameData_O[9]
+ Tile_X9Y10_LUT4AB/FrameStrobe[0] Tile_X9Y10_LUT4AB/FrameStrobe[10] Tile_X9Y10_LUT4AB/FrameStrobe[11]
+ Tile_X9Y10_LUT4AB/FrameStrobe[12] Tile_X9Y10_LUT4AB/FrameStrobe[13] Tile_X9Y10_LUT4AB/FrameStrobe[14]
+ Tile_X9Y10_LUT4AB/FrameStrobe[15] Tile_X9Y10_LUT4AB/FrameStrobe[16] Tile_X9Y10_LUT4AB/FrameStrobe[17]
+ Tile_X9Y10_LUT4AB/FrameStrobe[18] Tile_X9Y10_LUT4AB/FrameStrobe[19] Tile_X9Y10_LUT4AB/FrameStrobe[1]
+ Tile_X9Y10_LUT4AB/FrameStrobe[2] Tile_X9Y10_LUT4AB/FrameStrobe[3] Tile_X9Y10_LUT4AB/FrameStrobe[4]
+ Tile_X9Y10_LUT4AB/FrameStrobe[5] Tile_X9Y10_LUT4AB/FrameStrobe[6] Tile_X9Y10_LUT4AB/FrameStrobe[7]
+ Tile_X9Y10_LUT4AB/FrameStrobe[8] Tile_X9Y10_LUT4AB/FrameStrobe[9] Tile_X9Y9_LUT4AB/FrameStrobe[0]
+ Tile_X9Y9_LUT4AB/FrameStrobe[10] Tile_X9Y9_LUT4AB/FrameStrobe[11] Tile_X9Y9_LUT4AB/FrameStrobe[12]
+ Tile_X9Y9_LUT4AB/FrameStrobe[13] Tile_X9Y9_LUT4AB/FrameStrobe[14] Tile_X9Y9_LUT4AB/FrameStrobe[15]
+ Tile_X9Y9_LUT4AB/FrameStrobe[16] Tile_X9Y9_LUT4AB/FrameStrobe[17] Tile_X9Y9_LUT4AB/FrameStrobe[18]
+ Tile_X9Y9_LUT4AB/FrameStrobe[19] Tile_X9Y9_LUT4AB/FrameStrobe[1] Tile_X9Y9_LUT4AB/FrameStrobe[2]
+ Tile_X9Y9_LUT4AB/FrameStrobe[3] Tile_X9Y9_LUT4AB/FrameStrobe[4] Tile_X9Y9_LUT4AB/FrameStrobe[5]
+ Tile_X9Y9_LUT4AB/FrameStrobe[6] Tile_X9Y9_LUT4AB/FrameStrobe[7] Tile_X9Y9_LUT4AB/FrameStrobe[8]
+ Tile_X9Y9_LUT4AB/FrameStrobe[9] Tile_X9Y9_LUT4AB/N1END[0] Tile_X9Y9_LUT4AB/N1END[1]
+ Tile_X9Y9_LUT4AB/N1END[2] Tile_X9Y9_LUT4AB/N1END[3] Tile_X9Y11_LUT4AB/N1BEG[0] Tile_X9Y11_LUT4AB/N1BEG[1]
+ Tile_X9Y11_LUT4AB/N1BEG[2] Tile_X9Y11_LUT4AB/N1BEG[3] Tile_X9Y9_LUT4AB/N2MID[0]
+ Tile_X9Y9_LUT4AB/N2MID[1] Tile_X9Y9_LUT4AB/N2MID[2] Tile_X9Y9_LUT4AB/N2MID[3] Tile_X9Y9_LUT4AB/N2MID[4]
+ Tile_X9Y9_LUT4AB/N2MID[5] Tile_X9Y9_LUT4AB/N2MID[6] Tile_X9Y9_LUT4AB/N2MID[7] Tile_X9Y9_LUT4AB/N2END[0]
+ Tile_X9Y9_LUT4AB/N2END[1] Tile_X9Y9_LUT4AB/N2END[2] Tile_X9Y9_LUT4AB/N2END[3] Tile_X9Y9_LUT4AB/N2END[4]
+ Tile_X9Y9_LUT4AB/N2END[5] Tile_X9Y9_LUT4AB/N2END[6] Tile_X9Y9_LUT4AB/N2END[7] Tile_X9Y10_LUT4AB/N2END[0]
+ Tile_X9Y10_LUT4AB/N2END[1] Tile_X9Y10_LUT4AB/N2END[2] Tile_X9Y10_LUT4AB/N2END[3]
+ Tile_X9Y10_LUT4AB/N2END[4] Tile_X9Y10_LUT4AB/N2END[5] Tile_X9Y10_LUT4AB/N2END[6]
+ Tile_X9Y10_LUT4AB/N2END[7] Tile_X9Y11_LUT4AB/N2BEG[0] Tile_X9Y11_LUT4AB/N2BEG[1]
+ Tile_X9Y11_LUT4AB/N2BEG[2] Tile_X9Y11_LUT4AB/N2BEG[3] Tile_X9Y11_LUT4AB/N2BEG[4]
+ Tile_X9Y11_LUT4AB/N2BEG[5] Tile_X9Y11_LUT4AB/N2BEG[6] Tile_X9Y11_LUT4AB/N2BEG[7]
+ Tile_X9Y9_LUT4AB/N4END[0] Tile_X9Y9_LUT4AB/N4END[10] Tile_X9Y9_LUT4AB/N4END[11]
+ Tile_X9Y9_LUT4AB/N4END[12] Tile_X9Y9_LUT4AB/N4END[13] Tile_X9Y9_LUT4AB/N4END[14]
+ Tile_X9Y9_LUT4AB/N4END[15] Tile_X9Y9_LUT4AB/N4END[1] Tile_X9Y9_LUT4AB/N4END[2] Tile_X9Y9_LUT4AB/N4END[3]
+ Tile_X9Y9_LUT4AB/N4END[4] Tile_X9Y9_LUT4AB/N4END[5] Tile_X9Y9_LUT4AB/N4END[6] Tile_X9Y9_LUT4AB/N4END[7]
+ Tile_X9Y9_LUT4AB/N4END[8] Tile_X9Y9_LUT4AB/N4END[9] Tile_X9Y11_LUT4AB/N4BEG[0] Tile_X9Y11_LUT4AB/N4BEG[10]
+ Tile_X9Y11_LUT4AB/N4BEG[11] Tile_X9Y11_LUT4AB/N4BEG[12] Tile_X9Y11_LUT4AB/N4BEG[13]
+ Tile_X9Y11_LUT4AB/N4BEG[14] Tile_X9Y11_LUT4AB/N4BEG[15] Tile_X9Y11_LUT4AB/N4BEG[1]
+ Tile_X9Y11_LUT4AB/N4BEG[2] Tile_X9Y11_LUT4AB/N4BEG[3] Tile_X9Y11_LUT4AB/N4BEG[4]
+ Tile_X9Y11_LUT4AB/N4BEG[5] Tile_X9Y11_LUT4AB/N4BEG[6] Tile_X9Y11_LUT4AB/N4BEG[7]
+ Tile_X9Y11_LUT4AB/N4BEG[8] Tile_X9Y11_LUT4AB/N4BEG[9] Tile_X9Y9_LUT4AB/NN4END[0]
+ Tile_X9Y9_LUT4AB/NN4END[10] Tile_X9Y9_LUT4AB/NN4END[11] Tile_X9Y9_LUT4AB/NN4END[12]
+ Tile_X9Y9_LUT4AB/NN4END[13] Tile_X9Y9_LUT4AB/NN4END[14] Tile_X9Y9_LUT4AB/NN4END[15]
+ Tile_X9Y9_LUT4AB/NN4END[1] Tile_X9Y9_LUT4AB/NN4END[2] Tile_X9Y9_LUT4AB/NN4END[3]
+ Tile_X9Y9_LUT4AB/NN4END[4] Tile_X9Y9_LUT4AB/NN4END[5] Tile_X9Y9_LUT4AB/NN4END[6]
+ Tile_X9Y9_LUT4AB/NN4END[7] Tile_X9Y9_LUT4AB/NN4END[8] Tile_X9Y9_LUT4AB/NN4END[9]
+ Tile_X9Y11_LUT4AB/NN4BEG[0] Tile_X9Y11_LUT4AB/NN4BEG[10] Tile_X9Y11_LUT4AB/NN4BEG[11]
+ Tile_X9Y11_LUT4AB/NN4BEG[12] Tile_X9Y11_LUT4AB/NN4BEG[13] Tile_X9Y11_LUT4AB/NN4BEG[14]
+ Tile_X9Y11_LUT4AB/NN4BEG[15] Tile_X9Y11_LUT4AB/NN4BEG[1] Tile_X9Y11_LUT4AB/NN4BEG[2]
+ Tile_X9Y11_LUT4AB/NN4BEG[3] Tile_X9Y11_LUT4AB/NN4BEG[4] Tile_X9Y11_LUT4AB/NN4BEG[5]
+ Tile_X9Y11_LUT4AB/NN4BEG[6] Tile_X9Y11_LUT4AB/NN4BEG[7] Tile_X9Y11_LUT4AB/NN4BEG[8]
+ Tile_X9Y11_LUT4AB/NN4BEG[9] Tile_X9Y11_LUT4AB/S1END[0] Tile_X9Y11_LUT4AB/S1END[1]
+ Tile_X9Y11_LUT4AB/S1END[2] Tile_X9Y11_LUT4AB/S1END[3] Tile_X9Y9_LUT4AB/S1BEG[0]
+ Tile_X9Y9_LUT4AB/S1BEG[1] Tile_X9Y9_LUT4AB/S1BEG[2] Tile_X9Y9_LUT4AB/S1BEG[3] Tile_X9Y11_LUT4AB/S2MID[0]
+ Tile_X9Y11_LUT4AB/S2MID[1] Tile_X9Y11_LUT4AB/S2MID[2] Tile_X9Y11_LUT4AB/S2MID[3]
+ Tile_X9Y11_LUT4AB/S2MID[4] Tile_X9Y11_LUT4AB/S2MID[5] Tile_X9Y11_LUT4AB/S2MID[6]
+ Tile_X9Y11_LUT4AB/S2MID[7] Tile_X9Y11_LUT4AB/S2END[0] Tile_X9Y11_LUT4AB/S2END[1]
+ Tile_X9Y11_LUT4AB/S2END[2] Tile_X9Y11_LUT4AB/S2END[3] Tile_X9Y11_LUT4AB/S2END[4]
+ Tile_X9Y11_LUT4AB/S2END[5] Tile_X9Y11_LUT4AB/S2END[6] Tile_X9Y11_LUT4AB/S2END[7]
+ Tile_X9Y9_LUT4AB/S2BEGb[0] Tile_X9Y9_LUT4AB/S2BEGb[1] Tile_X9Y9_LUT4AB/S2BEGb[2]
+ Tile_X9Y9_LUT4AB/S2BEGb[3] Tile_X9Y9_LUT4AB/S2BEGb[4] Tile_X9Y9_LUT4AB/S2BEGb[5]
+ Tile_X9Y9_LUT4AB/S2BEGb[6] Tile_X9Y9_LUT4AB/S2BEGb[7] Tile_X9Y9_LUT4AB/S2BEG[0]
+ Tile_X9Y9_LUT4AB/S2BEG[1] Tile_X9Y9_LUT4AB/S2BEG[2] Tile_X9Y9_LUT4AB/S2BEG[3] Tile_X9Y9_LUT4AB/S2BEG[4]
+ Tile_X9Y9_LUT4AB/S2BEG[5] Tile_X9Y9_LUT4AB/S2BEG[6] Tile_X9Y9_LUT4AB/S2BEG[7] Tile_X9Y11_LUT4AB/S4END[0]
+ Tile_X9Y11_LUT4AB/S4END[10] Tile_X9Y11_LUT4AB/S4END[11] Tile_X9Y11_LUT4AB/S4END[12]
+ Tile_X9Y11_LUT4AB/S4END[13] Tile_X9Y11_LUT4AB/S4END[14] Tile_X9Y11_LUT4AB/S4END[15]
+ Tile_X9Y11_LUT4AB/S4END[1] Tile_X9Y11_LUT4AB/S4END[2] Tile_X9Y11_LUT4AB/S4END[3]
+ Tile_X9Y11_LUT4AB/S4END[4] Tile_X9Y11_LUT4AB/S4END[5] Tile_X9Y11_LUT4AB/S4END[6]
+ Tile_X9Y11_LUT4AB/S4END[7] Tile_X9Y11_LUT4AB/S4END[8] Tile_X9Y11_LUT4AB/S4END[9]
+ Tile_X9Y9_LUT4AB/S4BEG[0] Tile_X9Y9_LUT4AB/S4BEG[10] Tile_X9Y9_LUT4AB/S4BEG[11]
+ Tile_X9Y9_LUT4AB/S4BEG[12] Tile_X9Y9_LUT4AB/S4BEG[13] Tile_X9Y9_LUT4AB/S4BEG[14]
+ Tile_X9Y9_LUT4AB/S4BEG[15] Tile_X9Y9_LUT4AB/S4BEG[1] Tile_X9Y9_LUT4AB/S4BEG[2] Tile_X9Y9_LUT4AB/S4BEG[3]
+ Tile_X9Y9_LUT4AB/S4BEG[4] Tile_X9Y9_LUT4AB/S4BEG[5] Tile_X9Y9_LUT4AB/S4BEG[6] Tile_X9Y9_LUT4AB/S4BEG[7]
+ Tile_X9Y9_LUT4AB/S4BEG[8] Tile_X9Y9_LUT4AB/S4BEG[9] Tile_X9Y11_LUT4AB/SS4END[0]
+ Tile_X9Y11_LUT4AB/SS4END[10] Tile_X9Y11_LUT4AB/SS4END[11] Tile_X9Y11_LUT4AB/SS4END[12]
+ Tile_X9Y11_LUT4AB/SS4END[13] Tile_X9Y11_LUT4AB/SS4END[14] Tile_X9Y11_LUT4AB/SS4END[15]
+ Tile_X9Y11_LUT4AB/SS4END[1] Tile_X9Y11_LUT4AB/SS4END[2] Tile_X9Y11_LUT4AB/SS4END[3]
+ Tile_X9Y11_LUT4AB/SS4END[4] Tile_X9Y11_LUT4AB/SS4END[5] Tile_X9Y11_LUT4AB/SS4END[6]
+ Tile_X9Y11_LUT4AB/SS4END[7] Tile_X9Y11_LUT4AB/SS4END[8] Tile_X9Y11_LUT4AB/SS4END[9]
+ Tile_X9Y9_LUT4AB/SS4BEG[0] Tile_X9Y9_LUT4AB/SS4BEG[10] Tile_X9Y9_LUT4AB/SS4BEG[11]
+ Tile_X9Y9_LUT4AB/SS4BEG[12] Tile_X9Y9_LUT4AB/SS4BEG[13] Tile_X9Y9_LUT4AB/SS4BEG[14]
+ Tile_X9Y9_LUT4AB/SS4BEG[15] Tile_X9Y9_LUT4AB/SS4BEG[1] Tile_X9Y9_LUT4AB/SS4BEG[2]
+ Tile_X9Y9_LUT4AB/SS4BEG[3] Tile_X9Y9_LUT4AB/SS4BEG[4] Tile_X9Y9_LUT4AB/SS4BEG[5]
+ Tile_X9Y9_LUT4AB/SS4BEG[6] Tile_X9Y9_LUT4AB/SS4BEG[7] Tile_X9Y9_LUT4AB/SS4BEG[8]
+ Tile_X9Y9_LUT4AB/SS4BEG[9] Tile_X9Y10_LUT4AB/UserCLK Tile_X9Y9_LUT4AB/UserCLK VGND
+ VPWR Tile_X9Y10_LUT4AB/W1BEG[0] Tile_X9Y10_LUT4AB/W1BEG[1] Tile_X9Y10_LUT4AB/W1BEG[2]
+ Tile_X9Y10_LUT4AB/W1BEG[3] Tile_X9Y10_LUT4AB/W1END[0] Tile_X9Y10_LUT4AB/W1END[1]
+ Tile_X9Y10_LUT4AB/W1END[2] Tile_X9Y10_LUT4AB/W1END[3] Tile_X9Y10_LUT4AB/W2BEG[0]
+ Tile_X9Y10_LUT4AB/W2BEG[1] Tile_X9Y10_LUT4AB/W2BEG[2] Tile_X9Y10_LUT4AB/W2BEG[3]
+ Tile_X9Y10_LUT4AB/W2BEG[4] Tile_X9Y10_LUT4AB/W2BEG[5] Tile_X9Y10_LUT4AB/W2BEG[6]
+ Tile_X9Y10_LUT4AB/W2BEG[7] Tile_X8Y10_LUT4AB/W2END[0] Tile_X8Y10_LUT4AB/W2END[1]
+ Tile_X8Y10_LUT4AB/W2END[2] Tile_X8Y10_LUT4AB/W2END[3] Tile_X8Y10_LUT4AB/W2END[4]
+ Tile_X8Y10_LUT4AB/W2END[5] Tile_X8Y10_LUT4AB/W2END[6] Tile_X8Y10_LUT4AB/W2END[7]
+ Tile_X9Y10_LUT4AB/W2END[0] Tile_X9Y10_LUT4AB/W2END[1] Tile_X9Y10_LUT4AB/W2END[2]
+ Tile_X9Y10_LUT4AB/W2END[3] Tile_X9Y10_LUT4AB/W2END[4] Tile_X9Y10_LUT4AB/W2END[5]
+ Tile_X9Y10_LUT4AB/W2END[6] Tile_X9Y10_LUT4AB/W2END[7] Tile_X9Y10_LUT4AB/W2MID[0]
+ Tile_X9Y10_LUT4AB/W2MID[1] Tile_X9Y10_LUT4AB/W2MID[2] Tile_X9Y10_LUT4AB/W2MID[3]
+ Tile_X9Y10_LUT4AB/W2MID[4] Tile_X9Y10_LUT4AB/W2MID[5] Tile_X9Y10_LUT4AB/W2MID[6]
+ Tile_X9Y10_LUT4AB/W2MID[7] Tile_X9Y10_LUT4AB/W6BEG[0] Tile_X9Y10_LUT4AB/W6BEG[10]
+ Tile_X9Y10_LUT4AB/W6BEG[11] Tile_X9Y10_LUT4AB/W6BEG[1] Tile_X9Y10_LUT4AB/W6BEG[2]
+ Tile_X9Y10_LUT4AB/W6BEG[3] Tile_X9Y10_LUT4AB/W6BEG[4] Tile_X9Y10_LUT4AB/W6BEG[5]
+ Tile_X9Y10_LUT4AB/W6BEG[6] Tile_X9Y10_LUT4AB/W6BEG[7] Tile_X9Y10_LUT4AB/W6BEG[8]
+ Tile_X9Y10_LUT4AB/W6BEG[9] Tile_X9Y10_LUT4AB/W6END[0] Tile_X9Y10_LUT4AB/W6END[10]
+ Tile_X9Y10_LUT4AB/W6END[11] Tile_X9Y10_LUT4AB/W6END[1] Tile_X9Y10_LUT4AB/W6END[2]
+ Tile_X9Y10_LUT4AB/W6END[3] Tile_X9Y10_LUT4AB/W6END[4] Tile_X9Y10_LUT4AB/W6END[5]
+ Tile_X9Y10_LUT4AB/W6END[6] Tile_X9Y10_LUT4AB/W6END[7] Tile_X9Y10_LUT4AB/W6END[8]
+ Tile_X9Y10_LUT4AB/W6END[9] Tile_X9Y10_LUT4AB/WW4BEG[0] Tile_X9Y10_LUT4AB/WW4BEG[10]
+ Tile_X9Y10_LUT4AB/WW4BEG[11] Tile_X9Y10_LUT4AB/WW4BEG[12] Tile_X9Y10_LUT4AB/WW4BEG[13]
+ Tile_X9Y10_LUT4AB/WW4BEG[14] Tile_X9Y10_LUT4AB/WW4BEG[15] Tile_X9Y10_LUT4AB/WW4BEG[1]
+ Tile_X9Y10_LUT4AB/WW4BEG[2] Tile_X9Y10_LUT4AB/WW4BEG[3] Tile_X9Y10_LUT4AB/WW4BEG[4]
+ Tile_X9Y10_LUT4AB/WW4BEG[5] Tile_X9Y10_LUT4AB/WW4BEG[6] Tile_X9Y10_LUT4AB/WW4BEG[7]
+ Tile_X9Y10_LUT4AB/WW4BEG[8] Tile_X9Y10_LUT4AB/WW4BEG[9] Tile_X9Y10_LUT4AB/WW4END[0]
+ Tile_X9Y10_LUT4AB/WW4END[10] Tile_X9Y10_LUT4AB/WW4END[11] Tile_X9Y10_LUT4AB/WW4END[12]
+ Tile_X9Y10_LUT4AB/WW4END[13] Tile_X9Y10_LUT4AB/WW4END[14] Tile_X9Y10_LUT4AB/WW4END[15]
+ Tile_X9Y10_LUT4AB/WW4END[1] Tile_X9Y10_LUT4AB/WW4END[2] Tile_X9Y10_LUT4AB/WW4END[3]
+ Tile_X9Y10_LUT4AB/WW4END[4] Tile_X9Y10_LUT4AB/WW4END[5] Tile_X9Y10_LUT4AB/WW4END[6]
+ Tile_X9Y10_LUT4AB/WW4END[7] Tile_X9Y10_LUT4AB/WW4END[8] Tile_X9Y10_LUT4AB/WW4END[9]
+ LUT4AB
XTile_X4Y1_RegFile Tile_X5Y1_LUT4AB/E1END[0] Tile_X5Y1_LUT4AB/E1END[1] Tile_X5Y1_LUT4AB/E1END[2]
+ Tile_X5Y1_LUT4AB/E1END[3] Tile_X3Y1_LUT4AB/E1BEG[0] Tile_X3Y1_LUT4AB/E1BEG[1] Tile_X3Y1_LUT4AB/E1BEG[2]
+ Tile_X3Y1_LUT4AB/E1BEG[3] Tile_X5Y1_LUT4AB/E2MID[0] Tile_X5Y1_LUT4AB/E2MID[1] Tile_X5Y1_LUT4AB/E2MID[2]
+ Tile_X5Y1_LUT4AB/E2MID[3] Tile_X5Y1_LUT4AB/E2MID[4] Tile_X5Y1_LUT4AB/E2MID[5] Tile_X5Y1_LUT4AB/E2MID[6]
+ Tile_X5Y1_LUT4AB/E2MID[7] Tile_X5Y1_LUT4AB/E2END[0] Tile_X5Y1_LUT4AB/E2END[1] Tile_X5Y1_LUT4AB/E2END[2]
+ Tile_X5Y1_LUT4AB/E2END[3] Tile_X5Y1_LUT4AB/E2END[4] Tile_X5Y1_LUT4AB/E2END[5] Tile_X5Y1_LUT4AB/E2END[6]
+ Tile_X5Y1_LUT4AB/E2END[7] Tile_X4Y1_RegFile/E2END[0] Tile_X4Y1_RegFile/E2END[1]
+ Tile_X4Y1_RegFile/E2END[2] Tile_X4Y1_RegFile/E2END[3] Tile_X4Y1_RegFile/E2END[4]
+ Tile_X4Y1_RegFile/E2END[5] Tile_X4Y1_RegFile/E2END[6] Tile_X4Y1_RegFile/E2END[7]
+ Tile_X3Y1_LUT4AB/E2BEG[0] Tile_X3Y1_LUT4AB/E2BEG[1] Tile_X3Y1_LUT4AB/E2BEG[2] Tile_X3Y1_LUT4AB/E2BEG[3]
+ Tile_X3Y1_LUT4AB/E2BEG[4] Tile_X3Y1_LUT4AB/E2BEG[5] Tile_X3Y1_LUT4AB/E2BEG[6] Tile_X3Y1_LUT4AB/E2BEG[7]
+ Tile_X5Y1_LUT4AB/E6END[0] Tile_X5Y1_LUT4AB/E6END[10] Tile_X5Y1_LUT4AB/E6END[11]
+ Tile_X5Y1_LUT4AB/E6END[1] Tile_X5Y1_LUT4AB/E6END[2] Tile_X5Y1_LUT4AB/E6END[3] Tile_X5Y1_LUT4AB/E6END[4]
+ Tile_X5Y1_LUT4AB/E6END[5] Tile_X5Y1_LUT4AB/E6END[6] Tile_X5Y1_LUT4AB/E6END[7] Tile_X5Y1_LUT4AB/E6END[8]
+ Tile_X5Y1_LUT4AB/E6END[9] Tile_X3Y1_LUT4AB/E6BEG[0] Tile_X3Y1_LUT4AB/E6BEG[10] Tile_X3Y1_LUT4AB/E6BEG[11]
+ Tile_X3Y1_LUT4AB/E6BEG[1] Tile_X3Y1_LUT4AB/E6BEG[2] Tile_X3Y1_LUT4AB/E6BEG[3] Tile_X3Y1_LUT4AB/E6BEG[4]
+ Tile_X3Y1_LUT4AB/E6BEG[5] Tile_X3Y1_LUT4AB/E6BEG[6] Tile_X3Y1_LUT4AB/E6BEG[7] Tile_X3Y1_LUT4AB/E6BEG[8]
+ Tile_X3Y1_LUT4AB/E6BEG[9] Tile_X5Y1_LUT4AB/EE4END[0] Tile_X5Y1_LUT4AB/EE4END[10]
+ Tile_X5Y1_LUT4AB/EE4END[11] Tile_X5Y1_LUT4AB/EE4END[12] Tile_X5Y1_LUT4AB/EE4END[13]
+ Tile_X5Y1_LUT4AB/EE4END[14] Tile_X5Y1_LUT4AB/EE4END[15] Tile_X5Y1_LUT4AB/EE4END[1]
+ Tile_X5Y1_LUT4AB/EE4END[2] Tile_X5Y1_LUT4AB/EE4END[3] Tile_X5Y1_LUT4AB/EE4END[4]
+ Tile_X5Y1_LUT4AB/EE4END[5] Tile_X5Y1_LUT4AB/EE4END[6] Tile_X5Y1_LUT4AB/EE4END[7]
+ Tile_X5Y1_LUT4AB/EE4END[8] Tile_X5Y1_LUT4AB/EE4END[9] Tile_X3Y1_LUT4AB/EE4BEG[0]
+ Tile_X3Y1_LUT4AB/EE4BEG[10] Tile_X3Y1_LUT4AB/EE4BEG[11] Tile_X3Y1_LUT4AB/EE4BEG[12]
+ Tile_X3Y1_LUT4AB/EE4BEG[13] Tile_X3Y1_LUT4AB/EE4BEG[14] Tile_X3Y1_LUT4AB/EE4BEG[15]
+ Tile_X3Y1_LUT4AB/EE4BEG[1] Tile_X3Y1_LUT4AB/EE4BEG[2] Tile_X3Y1_LUT4AB/EE4BEG[3]
+ Tile_X3Y1_LUT4AB/EE4BEG[4] Tile_X3Y1_LUT4AB/EE4BEG[5] Tile_X3Y1_LUT4AB/EE4BEG[6]
+ Tile_X3Y1_LUT4AB/EE4BEG[7] Tile_X3Y1_LUT4AB/EE4BEG[8] Tile_X3Y1_LUT4AB/EE4BEG[9]
+ Tile_X4Y1_RegFile/FrameData[0] Tile_X4Y1_RegFile/FrameData[10] Tile_X4Y1_RegFile/FrameData[11]
+ Tile_X4Y1_RegFile/FrameData[12] Tile_X4Y1_RegFile/FrameData[13] Tile_X4Y1_RegFile/FrameData[14]
+ Tile_X4Y1_RegFile/FrameData[15] Tile_X4Y1_RegFile/FrameData[16] Tile_X4Y1_RegFile/FrameData[17]
+ Tile_X4Y1_RegFile/FrameData[18] Tile_X4Y1_RegFile/FrameData[19] Tile_X4Y1_RegFile/FrameData[1]
+ Tile_X4Y1_RegFile/FrameData[20] Tile_X4Y1_RegFile/FrameData[21] Tile_X4Y1_RegFile/FrameData[22]
+ Tile_X4Y1_RegFile/FrameData[23] Tile_X4Y1_RegFile/FrameData[24] Tile_X4Y1_RegFile/FrameData[25]
+ Tile_X4Y1_RegFile/FrameData[26] Tile_X4Y1_RegFile/FrameData[27] Tile_X4Y1_RegFile/FrameData[28]
+ Tile_X4Y1_RegFile/FrameData[29] Tile_X4Y1_RegFile/FrameData[2] Tile_X4Y1_RegFile/FrameData[30]
+ Tile_X4Y1_RegFile/FrameData[31] Tile_X4Y1_RegFile/FrameData[3] Tile_X4Y1_RegFile/FrameData[4]
+ Tile_X4Y1_RegFile/FrameData[5] Tile_X4Y1_RegFile/FrameData[6] Tile_X4Y1_RegFile/FrameData[7]
+ Tile_X4Y1_RegFile/FrameData[8] Tile_X4Y1_RegFile/FrameData[9] Tile_X5Y1_LUT4AB/FrameData[0]
+ Tile_X5Y1_LUT4AB/FrameData[10] Tile_X5Y1_LUT4AB/FrameData[11] Tile_X5Y1_LUT4AB/FrameData[12]
+ Tile_X5Y1_LUT4AB/FrameData[13] Tile_X5Y1_LUT4AB/FrameData[14] Tile_X5Y1_LUT4AB/FrameData[15]
+ Tile_X5Y1_LUT4AB/FrameData[16] Tile_X5Y1_LUT4AB/FrameData[17] Tile_X5Y1_LUT4AB/FrameData[18]
+ Tile_X5Y1_LUT4AB/FrameData[19] Tile_X5Y1_LUT4AB/FrameData[1] Tile_X5Y1_LUT4AB/FrameData[20]
+ Tile_X5Y1_LUT4AB/FrameData[21] Tile_X5Y1_LUT4AB/FrameData[22] Tile_X5Y1_LUT4AB/FrameData[23]
+ Tile_X5Y1_LUT4AB/FrameData[24] Tile_X5Y1_LUT4AB/FrameData[25] Tile_X5Y1_LUT4AB/FrameData[26]
+ Tile_X5Y1_LUT4AB/FrameData[27] Tile_X5Y1_LUT4AB/FrameData[28] Tile_X5Y1_LUT4AB/FrameData[29]
+ Tile_X5Y1_LUT4AB/FrameData[2] Tile_X5Y1_LUT4AB/FrameData[30] Tile_X5Y1_LUT4AB/FrameData[31]
+ Tile_X5Y1_LUT4AB/FrameData[3] Tile_X5Y1_LUT4AB/FrameData[4] Tile_X5Y1_LUT4AB/FrameData[5]
+ Tile_X5Y1_LUT4AB/FrameData[6] Tile_X5Y1_LUT4AB/FrameData[7] Tile_X5Y1_LUT4AB/FrameData[8]
+ Tile_X5Y1_LUT4AB/FrameData[9] Tile_X4Y1_RegFile/FrameStrobe[0] Tile_X4Y1_RegFile/FrameStrobe[10]
+ Tile_X4Y1_RegFile/FrameStrobe[11] Tile_X4Y1_RegFile/FrameStrobe[12] Tile_X4Y1_RegFile/FrameStrobe[13]
+ Tile_X4Y1_RegFile/FrameStrobe[14] Tile_X4Y1_RegFile/FrameStrobe[15] Tile_X4Y1_RegFile/FrameStrobe[16]
+ Tile_X4Y1_RegFile/FrameStrobe[17] Tile_X4Y1_RegFile/FrameStrobe[18] Tile_X4Y1_RegFile/FrameStrobe[19]
+ Tile_X4Y1_RegFile/FrameStrobe[1] Tile_X4Y1_RegFile/FrameStrobe[2] Tile_X4Y1_RegFile/FrameStrobe[3]
+ Tile_X4Y1_RegFile/FrameStrobe[4] Tile_X4Y1_RegFile/FrameStrobe[5] Tile_X4Y1_RegFile/FrameStrobe[6]
+ Tile_X4Y1_RegFile/FrameStrobe[7] Tile_X4Y1_RegFile/FrameStrobe[8] Tile_X4Y1_RegFile/FrameStrobe[9]
+ Tile_X4Y1_RegFile/FrameStrobe_O[0] Tile_X4Y1_RegFile/FrameStrobe_O[10] Tile_X4Y1_RegFile/FrameStrobe_O[11]
+ Tile_X4Y1_RegFile/FrameStrobe_O[12] Tile_X4Y1_RegFile/FrameStrobe_O[13] Tile_X4Y1_RegFile/FrameStrobe_O[14]
+ Tile_X4Y1_RegFile/FrameStrobe_O[15] Tile_X4Y1_RegFile/FrameStrobe_O[16] Tile_X4Y1_RegFile/FrameStrobe_O[17]
+ Tile_X4Y1_RegFile/FrameStrobe_O[18] Tile_X4Y1_RegFile/FrameStrobe_O[19] Tile_X4Y1_RegFile/FrameStrobe_O[1]
+ Tile_X4Y1_RegFile/FrameStrobe_O[2] Tile_X4Y1_RegFile/FrameStrobe_O[3] Tile_X4Y1_RegFile/FrameStrobe_O[4]
+ Tile_X4Y1_RegFile/FrameStrobe_O[5] Tile_X4Y1_RegFile/FrameStrobe_O[6] Tile_X4Y1_RegFile/FrameStrobe_O[7]
+ Tile_X4Y1_RegFile/FrameStrobe_O[8] Tile_X4Y1_RegFile/FrameStrobe_O[9] Tile_X4Y1_RegFile/N1BEG[0]
+ Tile_X4Y1_RegFile/N1BEG[1] Tile_X4Y1_RegFile/N1BEG[2] Tile_X4Y1_RegFile/N1BEG[3]
+ Tile_X4Y2_RegFile/N1BEG[0] Tile_X4Y2_RegFile/N1BEG[1] Tile_X4Y2_RegFile/N1BEG[2]
+ Tile_X4Y2_RegFile/N1BEG[3] Tile_X4Y1_RegFile/N2BEG[0] Tile_X4Y1_RegFile/N2BEG[1]
+ Tile_X4Y1_RegFile/N2BEG[2] Tile_X4Y1_RegFile/N2BEG[3] Tile_X4Y1_RegFile/N2BEG[4]
+ Tile_X4Y1_RegFile/N2BEG[5] Tile_X4Y1_RegFile/N2BEG[6] Tile_X4Y1_RegFile/N2BEG[7]
+ Tile_X4Y1_RegFile/N2BEGb[0] Tile_X4Y1_RegFile/N2BEGb[1] Tile_X4Y1_RegFile/N2BEGb[2]
+ Tile_X4Y1_RegFile/N2BEGb[3] Tile_X4Y1_RegFile/N2BEGb[4] Tile_X4Y1_RegFile/N2BEGb[5]
+ Tile_X4Y1_RegFile/N2BEGb[6] Tile_X4Y1_RegFile/N2BEGb[7] Tile_X4Y1_RegFile/N2END[0]
+ Tile_X4Y1_RegFile/N2END[1] Tile_X4Y1_RegFile/N2END[2] Tile_X4Y1_RegFile/N2END[3]
+ Tile_X4Y1_RegFile/N2END[4] Tile_X4Y1_RegFile/N2END[5] Tile_X4Y1_RegFile/N2END[6]
+ Tile_X4Y1_RegFile/N2END[7] Tile_X4Y2_RegFile/N2BEG[0] Tile_X4Y2_RegFile/N2BEG[1]
+ Tile_X4Y2_RegFile/N2BEG[2] Tile_X4Y2_RegFile/N2BEG[3] Tile_X4Y2_RegFile/N2BEG[4]
+ Tile_X4Y2_RegFile/N2BEG[5] Tile_X4Y2_RegFile/N2BEG[6] Tile_X4Y2_RegFile/N2BEG[7]
+ Tile_X4Y1_RegFile/N4BEG[0] Tile_X4Y1_RegFile/N4BEG[10] Tile_X4Y1_RegFile/N4BEG[11]
+ Tile_X4Y1_RegFile/N4BEG[12] Tile_X4Y1_RegFile/N4BEG[13] Tile_X4Y1_RegFile/N4BEG[14]
+ Tile_X4Y1_RegFile/N4BEG[15] Tile_X4Y1_RegFile/N4BEG[1] Tile_X4Y1_RegFile/N4BEG[2]
+ Tile_X4Y1_RegFile/N4BEG[3] Tile_X4Y1_RegFile/N4BEG[4] Tile_X4Y1_RegFile/N4BEG[5]
+ Tile_X4Y1_RegFile/N4BEG[6] Tile_X4Y1_RegFile/N4BEG[7] Tile_X4Y1_RegFile/N4BEG[8]
+ Tile_X4Y1_RegFile/N4BEG[9] Tile_X4Y2_RegFile/N4BEG[0] Tile_X4Y2_RegFile/N4BEG[10]
+ Tile_X4Y2_RegFile/N4BEG[11] Tile_X4Y2_RegFile/N4BEG[12] Tile_X4Y2_RegFile/N4BEG[13]
+ Tile_X4Y2_RegFile/N4BEG[14] Tile_X4Y2_RegFile/N4BEG[15] Tile_X4Y2_RegFile/N4BEG[1]
+ Tile_X4Y2_RegFile/N4BEG[2] Tile_X4Y2_RegFile/N4BEG[3] Tile_X4Y2_RegFile/N4BEG[4]
+ Tile_X4Y2_RegFile/N4BEG[5] Tile_X4Y2_RegFile/N4BEG[6] Tile_X4Y2_RegFile/N4BEG[7]
+ Tile_X4Y2_RegFile/N4BEG[8] Tile_X4Y2_RegFile/N4BEG[9] Tile_X4Y1_RegFile/NN4BEG[0]
+ Tile_X4Y1_RegFile/NN4BEG[10] Tile_X4Y1_RegFile/NN4BEG[11] Tile_X4Y1_RegFile/NN4BEG[12]
+ Tile_X4Y1_RegFile/NN4BEG[13] Tile_X4Y1_RegFile/NN4BEG[14] Tile_X4Y1_RegFile/NN4BEG[15]
+ Tile_X4Y1_RegFile/NN4BEG[1] Tile_X4Y1_RegFile/NN4BEG[2] Tile_X4Y1_RegFile/NN4BEG[3]
+ Tile_X4Y1_RegFile/NN4BEG[4] Tile_X4Y1_RegFile/NN4BEG[5] Tile_X4Y1_RegFile/NN4BEG[6]
+ Tile_X4Y1_RegFile/NN4BEG[7] Tile_X4Y1_RegFile/NN4BEG[8] Tile_X4Y1_RegFile/NN4BEG[9]
+ Tile_X4Y2_RegFile/NN4BEG[0] Tile_X4Y2_RegFile/NN4BEG[10] Tile_X4Y2_RegFile/NN4BEG[11]
+ Tile_X4Y2_RegFile/NN4BEG[12] Tile_X4Y2_RegFile/NN4BEG[13] Tile_X4Y2_RegFile/NN4BEG[14]
+ Tile_X4Y2_RegFile/NN4BEG[15] Tile_X4Y2_RegFile/NN4BEG[1] Tile_X4Y2_RegFile/NN4BEG[2]
+ Tile_X4Y2_RegFile/NN4BEG[3] Tile_X4Y2_RegFile/NN4BEG[4] Tile_X4Y2_RegFile/NN4BEG[5]
+ Tile_X4Y2_RegFile/NN4BEG[6] Tile_X4Y2_RegFile/NN4BEG[7] Tile_X4Y2_RegFile/NN4BEG[8]
+ Tile_X4Y2_RegFile/NN4BEG[9] Tile_X4Y2_RegFile/S1END[0] Tile_X4Y2_RegFile/S1END[1]
+ Tile_X4Y2_RegFile/S1END[2] Tile_X4Y2_RegFile/S1END[3] Tile_X4Y1_RegFile/S1END[0]
+ Tile_X4Y1_RegFile/S1END[1] Tile_X4Y1_RegFile/S1END[2] Tile_X4Y1_RegFile/S1END[3]
+ Tile_X4Y2_RegFile/S2MID[0] Tile_X4Y2_RegFile/S2MID[1] Tile_X4Y2_RegFile/S2MID[2]
+ Tile_X4Y2_RegFile/S2MID[3] Tile_X4Y2_RegFile/S2MID[4] Tile_X4Y2_RegFile/S2MID[5]
+ Tile_X4Y2_RegFile/S2MID[6] Tile_X4Y2_RegFile/S2MID[7] Tile_X4Y2_RegFile/S2END[0]
+ Tile_X4Y2_RegFile/S2END[1] Tile_X4Y2_RegFile/S2END[2] Tile_X4Y2_RegFile/S2END[3]
+ Tile_X4Y2_RegFile/S2END[4] Tile_X4Y2_RegFile/S2END[5] Tile_X4Y2_RegFile/S2END[6]
+ Tile_X4Y2_RegFile/S2END[7] Tile_X4Y1_RegFile/S2END[0] Tile_X4Y1_RegFile/S2END[1]
+ Tile_X4Y1_RegFile/S2END[2] Tile_X4Y1_RegFile/S2END[3] Tile_X4Y1_RegFile/S2END[4]
+ Tile_X4Y1_RegFile/S2END[5] Tile_X4Y1_RegFile/S2END[6] Tile_X4Y1_RegFile/S2END[7]
+ Tile_X4Y1_RegFile/S2MID[0] Tile_X4Y1_RegFile/S2MID[1] Tile_X4Y1_RegFile/S2MID[2]
+ Tile_X4Y1_RegFile/S2MID[3] Tile_X4Y1_RegFile/S2MID[4] Tile_X4Y1_RegFile/S2MID[5]
+ Tile_X4Y1_RegFile/S2MID[6] Tile_X4Y1_RegFile/S2MID[7] Tile_X4Y2_RegFile/S4END[0]
+ Tile_X4Y2_RegFile/S4END[10] Tile_X4Y2_RegFile/S4END[11] Tile_X4Y2_RegFile/S4END[12]
+ Tile_X4Y2_RegFile/S4END[13] Tile_X4Y2_RegFile/S4END[14] Tile_X4Y2_RegFile/S4END[15]
+ Tile_X4Y2_RegFile/S4END[1] Tile_X4Y2_RegFile/S4END[2] Tile_X4Y2_RegFile/S4END[3]
+ Tile_X4Y2_RegFile/S4END[4] Tile_X4Y2_RegFile/S4END[5] Tile_X4Y2_RegFile/S4END[6]
+ Tile_X4Y2_RegFile/S4END[7] Tile_X4Y2_RegFile/S4END[8] Tile_X4Y2_RegFile/S4END[9]
+ Tile_X4Y1_RegFile/S4END[0] Tile_X4Y1_RegFile/S4END[10] Tile_X4Y1_RegFile/S4END[11]
+ Tile_X4Y1_RegFile/S4END[12] Tile_X4Y1_RegFile/S4END[13] Tile_X4Y1_RegFile/S4END[14]
+ Tile_X4Y1_RegFile/S4END[15] Tile_X4Y1_RegFile/S4END[1] Tile_X4Y1_RegFile/S4END[2]
+ Tile_X4Y1_RegFile/S4END[3] Tile_X4Y1_RegFile/S4END[4] Tile_X4Y1_RegFile/S4END[5]
+ Tile_X4Y1_RegFile/S4END[6] Tile_X4Y1_RegFile/S4END[7] Tile_X4Y1_RegFile/S4END[8]
+ Tile_X4Y1_RegFile/S4END[9] Tile_X4Y2_RegFile/SS4END[0] Tile_X4Y2_RegFile/SS4END[10]
+ Tile_X4Y2_RegFile/SS4END[11] Tile_X4Y2_RegFile/SS4END[12] Tile_X4Y2_RegFile/SS4END[13]
+ Tile_X4Y2_RegFile/SS4END[14] Tile_X4Y2_RegFile/SS4END[15] Tile_X4Y2_RegFile/SS4END[1]
+ Tile_X4Y2_RegFile/SS4END[2] Tile_X4Y2_RegFile/SS4END[3] Tile_X4Y2_RegFile/SS4END[4]
+ Tile_X4Y2_RegFile/SS4END[5] Tile_X4Y2_RegFile/SS4END[6] Tile_X4Y2_RegFile/SS4END[7]
+ Tile_X4Y2_RegFile/SS4END[8] Tile_X4Y2_RegFile/SS4END[9] Tile_X4Y1_RegFile/SS4END[0]
+ Tile_X4Y1_RegFile/SS4END[10] Tile_X4Y1_RegFile/SS4END[11] Tile_X4Y1_RegFile/SS4END[12]
+ Tile_X4Y1_RegFile/SS4END[13] Tile_X4Y1_RegFile/SS4END[14] Tile_X4Y1_RegFile/SS4END[15]
+ Tile_X4Y1_RegFile/SS4END[1] Tile_X4Y1_RegFile/SS4END[2] Tile_X4Y1_RegFile/SS4END[3]
+ Tile_X4Y1_RegFile/SS4END[4] Tile_X4Y1_RegFile/SS4END[5] Tile_X4Y1_RegFile/SS4END[6]
+ Tile_X4Y1_RegFile/SS4END[7] Tile_X4Y1_RegFile/SS4END[8] Tile_X4Y1_RegFile/SS4END[9]
+ Tile_X4Y1_RegFile/UserCLK Tile_X4Y1_RegFile/UserCLKo VGND VPWR Tile_X3Y1_LUT4AB/W1END[0]
+ Tile_X3Y1_LUT4AB/W1END[1] Tile_X3Y1_LUT4AB/W1END[2] Tile_X3Y1_LUT4AB/W1END[3] Tile_X5Y1_LUT4AB/W1BEG[0]
+ Tile_X5Y1_LUT4AB/W1BEG[1] Tile_X5Y1_LUT4AB/W1BEG[2] Tile_X5Y1_LUT4AB/W1BEG[3] Tile_X3Y1_LUT4AB/W2MID[0]
+ Tile_X3Y1_LUT4AB/W2MID[1] Tile_X3Y1_LUT4AB/W2MID[2] Tile_X3Y1_LUT4AB/W2MID[3] Tile_X3Y1_LUT4AB/W2MID[4]
+ Tile_X3Y1_LUT4AB/W2MID[5] Tile_X3Y1_LUT4AB/W2MID[6] Tile_X3Y1_LUT4AB/W2MID[7] Tile_X3Y1_LUT4AB/W2END[0]
+ Tile_X3Y1_LUT4AB/W2END[1] Tile_X3Y1_LUT4AB/W2END[2] Tile_X3Y1_LUT4AB/W2END[3] Tile_X3Y1_LUT4AB/W2END[4]
+ Tile_X3Y1_LUT4AB/W2END[5] Tile_X3Y1_LUT4AB/W2END[6] Tile_X3Y1_LUT4AB/W2END[7] Tile_X5Y1_LUT4AB/W2BEGb[0]
+ Tile_X5Y1_LUT4AB/W2BEGb[1] Tile_X5Y1_LUT4AB/W2BEGb[2] Tile_X5Y1_LUT4AB/W2BEGb[3]
+ Tile_X5Y1_LUT4AB/W2BEGb[4] Tile_X5Y1_LUT4AB/W2BEGb[5] Tile_X5Y1_LUT4AB/W2BEGb[6]
+ Tile_X5Y1_LUT4AB/W2BEGb[7] Tile_X5Y1_LUT4AB/W2BEG[0] Tile_X5Y1_LUT4AB/W2BEG[1] Tile_X5Y1_LUT4AB/W2BEG[2]
+ Tile_X5Y1_LUT4AB/W2BEG[3] Tile_X5Y1_LUT4AB/W2BEG[4] Tile_X5Y1_LUT4AB/W2BEG[5] Tile_X5Y1_LUT4AB/W2BEG[6]
+ Tile_X5Y1_LUT4AB/W2BEG[7] Tile_X3Y1_LUT4AB/W6END[0] Tile_X3Y1_LUT4AB/W6END[10] Tile_X3Y1_LUT4AB/W6END[11]
+ Tile_X3Y1_LUT4AB/W6END[1] Tile_X3Y1_LUT4AB/W6END[2] Tile_X3Y1_LUT4AB/W6END[3] Tile_X3Y1_LUT4AB/W6END[4]
+ Tile_X3Y1_LUT4AB/W6END[5] Tile_X3Y1_LUT4AB/W6END[6] Tile_X3Y1_LUT4AB/W6END[7] Tile_X3Y1_LUT4AB/W6END[8]
+ Tile_X3Y1_LUT4AB/W6END[9] Tile_X5Y1_LUT4AB/W6BEG[0] Tile_X5Y1_LUT4AB/W6BEG[10] Tile_X5Y1_LUT4AB/W6BEG[11]
+ Tile_X5Y1_LUT4AB/W6BEG[1] Tile_X5Y1_LUT4AB/W6BEG[2] Tile_X5Y1_LUT4AB/W6BEG[3] Tile_X5Y1_LUT4AB/W6BEG[4]
+ Tile_X5Y1_LUT4AB/W6BEG[5] Tile_X5Y1_LUT4AB/W6BEG[6] Tile_X5Y1_LUT4AB/W6BEG[7] Tile_X5Y1_LUT4AB/W6BEG[8]
+ Tile_X5Y1_LUT4AB/W6BEG[9] Tile_X3Y1_LUT4AB/WW4END[0] Tile_X3Y1_LUT4AB/WW4END[10]
+ Tile_X3Y1_LUT4AB/WW4END[11] Tile_X3Y1_LUT4AB/WW4END[12] Tile_X3Y1_LUT4AB/WW4END[13]
+ Tile_X3Y1_LUT4AB/WW4END[14] Tile_X3Y1_LUT4AB/WW4END[15] Tile_X3Y1_LUT4AB/WW4END[1]
+ Tile_X3Y1_LUT4AB/WW4END[2] Tile_X3Y1_LUT4AB/WW4END[3] Tile_X3Y1_LUT4AB/WW4END[4]
+ Tile_X3Y1_LUT4AB/WW4END[5] Tile_X3Y1_LUT4AB/WW4END[6] Tile_X3Y1_LUT4AB/WW4END[7]
+ Tile_X3Y1_LUT4AB/WW4END[8] Tile_X3Y1_LUT4AB/WW4END[9] Tile_X5Y1_LUT4AB/WW4BEG[0]
+ Tile_X5Y1_LUT4AB/WW4BEG[10] Tile_X5Y1_LUT4AB/WW4BEG[11] Tile_X5Y1_LUT4AB/WW4BEG[12]
+ Tile_X5Y1_LUT4AB/WW4BEG[13] Tile_X5Y1_LUT4AB/WW4BEG[14] Tile_X5Y1_LUT4AB/WW4BEG[15]
+ Tile_X5Y1_LUT4AB/WW4BEG[1] Tile_X5Y1_LUT4AB/WW4BEG[2] Tile_X5Y1_LUT4AB/WW4BEG[3]
+ Tile_X5Y1_LUT4AB/WW4BEG[4] Tile_X5Y1_LUT4AB/WW4BEG[5] Tile_X5Y1_LUT4AB/WW4BEG[6]
+ Tile_X5Y1_LUT4AB/WW4BEG[7] Tile_X5Y1_LUT4AB/WW4BEG[8] Tile_X5Y1_LUT4AB/WW4BEG[9]
+ RegFile
XTile_X1Y15_S_term_single Tile_X1Y14_LUT4AB/Ci FrameData[480] FrameData[490] FrameData[491]
+ FrameData[492] FrameData[493] FrameData[494] FrameData[495] FrameData[496] FrameData[497]
+ FrameData[498] FrameData[499] FrameData[481] FrameData[500] FrameData[501] FrameData[502]
+ FrameData[503] FrameData[504] FrameData[505] FrameData[506] FrameData[507] FrameData[508]
+ FrameData[509] FrameData[482] FrameData[510] FrameData[511] FrameData[483] FrameData[484]
+ FrameData[485] FrameData[486] FrameData[487] FrameData[488] FrameData[489] Tile_X2Y15_S_WARMBOOT/FrameData[0]
+ Tile_X2Y15_S_WARMBOOT/FrameData[10] Tile_X2Y15_S_WARMBOOT/FrameData[11] Tile_X2Y15_S_WARMBOOT/FrameData[12]
+ Tile_X2Y15_S_WARMBOOT/FrameData[13] Tile_X2Y15_S_WARMBOOT/FrameData[14] Tile_X2Y15_S_WARMBOOT/FrameData[15]
+ Tile_X2Y15_S_WARMBOOT/FrameData[16] Tile_X2Y15_S_WARMBOOT/FrameData[17] Tile_X2Y15_S_WARMBOOT/FrameData[18]
+ Tile_X2Y15_S_WARMBOOT/FrameData[19] Tile_X2Y15_S_WARMBOOT/FrameData[1] Tile_X2Y15_S_WARMBOOT/FrameData[20]
+ Tile_X2Y15_S_WARMBOOT/FrameData[21] Tile_X2Y15_S_WARMBOOT/FrameData[22] Tile_X2Y15_S_WARMBOOT/FrameData[23]
+ Tile_X2Y15_S_WARMBOOT/FrameData[24] Tile_X2Y15_S_WARMBOOT/FrameData[25] Tile_X2Y15_S_WARMBOOT/FrameData[26]
+ Tile_X2Y15_S_WARMBOOT/FrameData[27] Tile_X2Y15_S_WARMBOOT/FrameData[28] Tile_X2Y15_S_WARMBOOT/FrameData[29]
+ Tile_X2Y15_S_WARMBOOT/FrameData[2] Tile_X2Y15_S_WARMBOOT/FrameData[30] Tile_X2Y15_S_WARMBOOT/FrameData[31]
+ Tile_X2Y15_S_WARMBOOT/FrameData[3] Tile_X2Y15_S_WARMBOOT/FrameData[4] Tile_X2Y15_S_WARMBOOT/FrameData[5]
+ Tile_X2Y15_S_WARMBOOT/FrameData[6] Tile_X2Y15_S_WARMBOOT/FrameData[7] Tile_X2Y15_S_WARMBOOT/FrameData[8]
+ Tile_X2Y15_S_WARMBOOT/FrameData[9] FrameStrobe[20] FrameStrobe[30] FrameStrobe[31]
+ FrameStrobe[32] FrameStrobe[33] FrameStrobe[34] FrameStrobe[35] FrameStrobe[36]
+ FrameStrobe[37] FrameStrobe[38] FrameStrobe[39] FrameStrobe[21] FrameStrobe[22]
+ FrameStrobe[23] FrameStrobe[24] FrameStrobe[25] FrameStrobe[26] FrameStrobe[27]
+ FrameStrobe[28] FrameStrobe[29] Tile_X1Y14_LUT4AB/FrameStrobe[0] Tile_X1Y14_LUT4AB/FrameStrobe[10]
+ Tile_X1Y14_LUT4AB/FrameStrobe[11] Tile_X1Y14_LUT4AB/FrameStrobe[12] Tile_X1Y14_LUT4AB/FrameStrobe[13]
+ Tile_X1Y14_LUT4AB/FrameStrobe[14] Tile_X1Y14_LUT4AB/FrameStrobe[15] Tile_X1Y14_LUT4AB/FrameStrobe[16]
+ Tile_X1Y14_LUT4AB/FrameStrobe[17] Tile_X1Y14_LUT4AB/FrameStrobe[18] Tile_X1Y14_LUT4AB/FrameStrobe[19]
+ Tile_X1Y14_LUT4AB/FrameStrobe[1] Tile_X1Y14_LUT4AB/FrameStrobe[2] Tile_X1Y14_LUT4AB/FrameStrobe[3]
+ Tile_X1Y14_LUT4AB/FrameStrobe[4] Tile_X1Y14_LUT4AB/FrameStrobe[5] Tile_X1Y14_LUT4AB/FrameStrobe[6]
+ Tile_X1Y14_LUT4AB/FrameStrobe[7] Tile_X1Y14_LUT4AB/FrameStrobe[8] Tile_X1Y14_LUT4AB/FrameStrobe[9]
+ Tile_X1Y14_LUT4AB/N1END[0] Tile_X1Y14_LUT4AB/N1END[1] Tile_X1Y14_LUT4AB/N1END[2]
+ Tile_X1Y14_LUT4AB/N1END[3] Tile_X1Y14_LUT4AB/N2MID[0] Tile_X1Y14_LUT4AB/N2MID[1]
+ Tile_X1Y14_LUT4AB/N2MID[2] Tile_X1Y14_LUT4AB/N2MID[3] Tile_X1Y14_LUT4AB/N2MID[4]
+ Tile_X1Y14_LUT4AB/N2MID[5] Tile_X1Y14_LUT4AB/N2MID[6] Tile_X1Y14_LUT4AB/N2MID[7]
+ Tile_X1Y14_LUT4AB/N2END[0] Tile_X1Y14_LUT4AB/N2END[1] Tile_X1Y14_LUT4AB/N2END[2]
+ Tile_X1Y14_LUT4AB/N2END[3] Tile_X1Y14_LUT4AB/N2END[4] Tile_X1Y14_LUT4AB/N2END[5]
+ Tile_X1Y14_LUT4AB/N2END[6] Tile_X1Y14_LUT4AB/N2END[7] Tile_X1Y14_LUT4AB/N4END[0]
+ Tile_X1Y14_LUT4AB/N4END[10] Tile_X1Y14_LUT4AB/N4END[11] Tile_X1Y14_LUT4AB/N4END[12]
+ Tile_X1Y14_LUT4AB/N4END[13] Tile_X1Y14_LUT4AB/N4END[14] Tile_X1Y14_LUT4AB/N4END[15]
+ Tile_X1Y14_LUT4AB/N4END[1] Tile_X1Y14_LUT4AB/N4END[2] Tile_X1Y14_LUT4AB/N4END[3]
+ Tile_X1Y14_LUT4AB/N4END[4] Tile_X1Y14_LUT4AB/N4END[5] Tile_X1Y14_LUT4AB/N4END[6]
+ Tile_X1Y14_LUT4AB/N4END[7] Tile_X1Y14_LUT4AB/N4END[8] Tile_X1Y14_LUT4AB/N4END[9]
+ Tile_X1Y14_LUT4AB/NN4END[0] Tile_X1Y14_LUT4AB/NN4END[10] Tile_X1Y14_LUT4AB/NN4END[11]
+ Tile_X1Y14_LUT4AB/NN4END[12] Tile_X1Y14_LUT4AB/NN4END[13] Tile_X1Y14_LUT4AB/NN4END[14]
+ Tile_X1Y14_LUT4AB/NN4END[15] Tile_X1Y14_LUT4AB/NN4END[1] Tile_X1Y14_LUT4AB/NN4END[2]
+ Tile_X1Y14_LUT4AB/NN4END[3] Tile_X1Y14_LUT4AB/NN4END[4] Tile_X1Y14_LUT4AB/NN4END[5]
+ Tile_X1Y14_LUT4AB/NN4END[6] Tile_X1Y14_LUT4AB/NN4END[7] Tile_X1Y14_LUT4AB/NN4END[8]
+ Tile_X1Y14_LUT4AB/NN4END[9] Tile_X1Y14_LUT4AB/S1BEG[0] Tile_X1Y14_LUT4AB/S1BEG[1]
+ Tile_X1Y14_LUT4AB/S1BEG[2] Tile_X1Y14_LUT4AB/S1BEG[3] Tile_X1Y14_LUT4AB/S2BEGb[0]
+ Tile_X1Y14_LUT4AB/S2BEGb[1] Tile_X1Y14_LUT4AB/S2BEGb[2] Tile_X1Y14_LUT4AB/S2BEGb[3]
+ Tile_X1Y14_LUT4AB/S2BEGb[4] Tile_X1Y14_LUT4AB/S2BEGb[5] Tile_X1Y14_LUT4AB/S2BEGb[6]
+ Tile_X1Y14_LUT4AB/S2BEGb[7] Tile_X1Y14_LUT4AB/S2BEG[0] Tile_X1Y14_LUT4AB/S2BEG[1]
+ Tile_X1Y14_LUT4AB/S2BEG[2] Tile_X1Y14_LUT4AB/S2BEG[3] Tile_X1Y14_LUT4AB/S2BEG[4]
+ Tile_X1Y14_LUT4AB/S2BEG[5] Tile_X1Y14_LUT4AB/S2BEG[6] Tile_X1Y14_LUT4AB/S2BEG[7]
+ Tile_X1Y14_LUT4AB/S4BEG[0] Tile_X1Y14_LUT4AB/S4BEG[10] Tile_X1Y14_LUT4AB/S4BEG[11]
+ Tile_X1Y14_LUT4AB/S4BEG[12] Tile_X1Y14_LUT4AB/S4BEG[13] Tile_X1Y14_LUT4AB/S4BEG[14]
+ Tile_X1Y14_LUT4AB/S4BEG[15] Tile_X1Y14_LUT4AB/S4BEG[1] Tile_X1Y14_LUT4AB/S4BEG[2]
+ Tile_X1Y14_LUT4AB/S4BEG[3] Tile_X1Y14_LUT4AB/S4BEG[4] Tile_X1Y14_LUT4AB/S4BEG[5]
+ Tile_X1Y14_LUT4AB/S4BEG[6] Tile_X1Y14_LUT4AB/S4BEG[7] Tile_X1Y14_LUT4AB/S4BEG[8]
+ Tile_X1Y14_LUT4AB/S4BEG[9] Tile_X1Y14_LUT4AB/SS4BEG[0] Tile_X1Y14_LUT4AB/SS4BEG[10]
+ Tile_X1Y14_LUT4AB/SS4BEG[11] Tile_X1Y14_LUT4AB/SS4BEG[12] Tile_X1Y14_LUT4AB/SS4BEG[13]
+ Tile_X1Y14_LUT4AB/SS4BEG[14] Tile_X1Y14_LUT4AB/SS4BEG[15] Tile_X1Y14_LUT4AB/SS4BEG[1]
+ Tile_X1Y14_LUT4AB/SS4BEG[2] Tile_X1Y14_LUT4AB/SS4BEG[3] Tile_X1Y14_LUT4AB/SS4BEG[4]
+ Tile_X1Y14_LUT4AB/SS4BEG[5] Tile_X1Y14_LUT4AB/SS4BEG[6] Tile_X1Y14_LUT4AB/SS4BEG[7]
+ Tile_X1Y14_LUT4AB/SS4BEG[8] Tile_X1Y14_LUT4AB/SS4BEG[9] UserCLK Tile_X1Y14_LUT4AB/UserCLK
+ VGND VPWR S_term_single
XTile_X9Y0_N_term_single Tile_X9Y1_LUT4AB/Co Tile_X9Y0_N_term_single/FrameData[0]
+ Tile_X9Y0_N_term_single/FrameData[10] Tile_X9Y0_N_term_single/FrameData[11] Tile_X9Y0_N_term_single/FrameData[12]
+ Tile_X9Y0_N_term_single/FrameData[13] Tile_X9Y0_N_term_single/FrameData[14] Tile_X9Y0_N_term_single/FrameData[15]
+ Tile_X9Y0_N_term_single/FrameData[16] Tile_X9Y0_N_term_single/FrameData[17] Tile_X9Y0_N_term_single/FrameData[18]
+ Tile_X9Y0_N_term_single/FrameData[19] Tile_X9Y0_N_term_single/FrameData[1] Tile_X9Y0_N_term_single/FrameData[20]
+ Tile_X9Y0_N_term_single/FrameData[21] Tile_X9Y0_N_term_single/FrameData[22] Tile_X9Y0_N_term_single/FrameData[23]
+ Tile_X9Y0_N_term_single/FrameData[24] Tile_X9Y0_N_term_single/FrameData[25] Tile_X9Y0_N_term_single/FrameData[26]
+ Tile_X9Y0_N_term_single/FrameData[27] Tile_X9Y0_N_term_single/FrameData[28] Tile_X9Y0_N_term_single/FrameData[29]
+ Tile_X9Y0_N_term_single/FrameData[2] Tile_X9Y0_N_term_single/FrameData[30] Tile_X9Y0_N_term_single/FrameData[31]
+ Tile_X9Y0_N_term_single/FrameData[3] Tile_X9Y0_N_term_single/FrameData[4] Tile_X9Y0_N_term_single/FrameData[5]
+ Tile_X9Y0_N_term_single/FrameData[6] Tile_X9Y0_N_term_single/FrameData[7] Tile_X9Y0_N_term_single/FrameData[8]
+ Tile_X9Y0_N_term_single/FrameData[9] Tile_X9Y0_N_term_single/FrameData_O[0] Tile_X9Y0_N_term_single/FrameData_O[10]
+ Tile_X9Y0_N_term_single/FrameData_O[11] Tile_X9Y0_N_term_single/FrameData_O[12]
+ Tile_X9Y0_N_term_single/FrameData_O[13] Tile_X9Y0_N_term_single/FrameData_O[14]
+ Tile_X9Y0_N_term_single/FrameData_O[15] Tile_X9Y0_N_term_single/FrameData_O[16]
+ Tile_X9Y0_N_term_single/FrameData_O[17] Tile_X9Y0_N_term_single/FrameData_O[18]
+ Tile_X9Y0_N_term_single/FrameData_O[19] Tile_X9Y0_N_term_single/FrameData_O[1] Tile_X9Y0_N_term_single/FrameData_O[20]
+ Tile_X9Y0_N_term_single/FrameData_O[21] Tile_X9Y0_N_term_single/FrameData_O[22]
+ Tile_X9Y0_N_term_single/FrameData_O[23] Tile_X9Y0_N_term_single/FrameData_O[24]
+ Tile_X9Y0_N_term_single/FrameData_O[25] Tile_X9Y0_N_term_single/FrameData_O[26]
+ Tile_X9Y0_N_term_single/FrameData_O[27] Tile_X9Y0_N_term_single/FrameData_O[28]
+ Tile_X9Y0_N_term_single/FrameData_O[29] Tile_X9Y0_N_term_single/FrameData_O[2] Tile_X9Y0_N_term_single/FrameData_O[30]
+ Tile_X9Y0_N_term_single/FrameData_O[31] Tile_X9Y0_N_term_single/FrameData_O[3] Tile_X9Y0_N_term_single/FrameData_O[4]
+ Tile_X9Y0_N_term_single/FrameData_O[5] Tile_X9Y0_N_term_single/FrameData_O[6] Tile_X9Y0_N_term_single/FrameData_O[7]
+ Tile_X9Y0_N_term_single/FrameData_O[8] Tile_X9Y0_N_term_single/FrameData_O[9] Tile_X9Y1_LUT4AB/FrameStrobe_O[0]
+ Tile_X9Y1_LUT4AB/FrameStrobe_O[10] Tile_X9Y1_LUT4AB/FrameStrobe_O[11] Tile_X9Y1_LUT4AB/FrameStrobe_O[12]
+ Tile_X9Y1_LUT4AB/FrameStrobe_O[13] Tile_X9Y1_LUT4AB/FrameStrobe_O[14] Tile_X9Y1_LUT4AB/FrameStrobe_O[15]
+ Tile_X9Y1_LUT4AB/FrameStrobe_O[16] Tile_X9Y1_LUT4AB/FrameStrobe_O[17] Tile_X9Y1_LUT4AB/FrameStrobe_O[18]
+ Tile_X9Y1_LUT4AB/FrameStrobe_O[19] Tile_X9Y1_LUT4AB/FrameStrobe_O[1] Tile_X9Y1_LUT4AB/FrameStrobe_O[2]
+ Tile_X9Y1_LUT4AB/FrameStrobe_O[3] Tile_X9Y1_LUT4AB/FrameStrobe_O[4] Tile_X9Y1_LUT4AB/FrameStrobe_O[5]
+ Tile_X9Y1_LUT4AB/FrameStrobe_O[6] Tile_X9Y1_LUT4AB/FrameStrobe_O[7] Tile_X9Y1_LUT4AB/FrameStrobe_O[8]
+ Tile_X9Y1_LUT4AB/FrameStrobe_O[9] Tile_X9Y0_N_term_single/FrameStrobe_O[0] Tile_X9Y0_N_term_single/FrameStrobe_O[10]
+ Tile_X9Y0_N_term_single/FrameStrobe_O[11] Tile_X9Y0_N_term_single/FrameStrobe_O[12]
+ Tile_X9Y0_N_term_single/FrameStrobe_O[13] Tile_X9Y0_N_term_single/FrameStrobe_O[14]
+ Tile_X9Y0_N_term_single/FrameStrobe_O[15] Tile_X9Y0_N_term_single/FrameStrobe_O[16]
+ Tile_X9Y0_N_term_single/FrameStrobe_O[17] Tile_X9Y0_N_term_single/FrameStrobe_O[18]
+ Tile_X9Y0_N_term_single/FrameStrobe_O[19] Tile_X9Y0_N_term_single/FrameStrobe_O[1]
+ Tile_X9Y0_N_term_single/FrameStrobe_O[2] Tile_X9Y0_N_term_single/FrameStrobe_O[3]
+ Tile_X9Y0_N_term_single/FrameStrobe_O[4] Tile_X9Y0_N_term_single/FrameStrobe_O[5]
+ Tile_X9Y0_N_term_single/FrameStrobe_O[6] Tile_X9Y0_N_term_single/FrameStrobe_O[7]
+ Tile_X9Y0_N_term_single/FrameStrobe_O[8] Tile_X9Y0_N_term_single/FrameStrobe_O[9]
+ Tile_X9Y1_LUT4AB/N1BEG[0] Tile_X9Y1_LUT4AB/N1BEG[1] Tile_X9Y1_LUT4AB/N1BEG[2] Tile_X9Y1_LUT4AB/N1BEG[3]
+ Tile_X9Y1_LUT4AB/N2BEGb[0] Tile_X9Y1_LUT4AB/N2BEGb[1] Tile_X9Y1_LUT4AB/N2BEGb[2]
+ Tile_X9Y1_LUT4AB/N2BEGb[3] Tile_X9Y1_LUT4AB/N2BEGb[4] Tile_X9Y1_LUT4AB/N2BEGb[5]
+ Tile_X9Y1_LUT4AB/N2BEGb[6] Tile_X9Y1_LUT4AB/N2BEGb[7] Tile_X9Y1_LUT4AB/N2BEG[0]
+ Tile_X9Y1_LUT4AB/N2BEG[1] Tile_X9Y1_LUT4AB/N2BEG[2] Tile_X9Y1_LUT4AB/N2BEG[3] Tile_X9Y1_LUT4AB/N2BEG[4]
+ Tile_X9Y1_LUT4AB/N2BEG[5] Tile_X9Y1_LUT4AB/N2BEG[6] Tile_X9Y1_LUT4AB/N2BEG[7] Tile_X9Y1_LUT4AB/N4BEG[0]
+ Tile_X9Y1_LUT4AB/N4BEG[10] Tile_X9Y1_LUT4AB/N4BEG[11] Tile_X9Y1_LUT4AB/N4BEG[12]
+ Tile_X9Y1_LUT4AB/N4BEG[13] Tile_X9Y1_LUT4AB/N4BEG[14] Tile_X9Y1_LUT4AB/N4BEG[15]
+ Tile_X9Y1_LUT4AB/N4BEG[1] Tile_X9Y1_LUT4AB/N4BEG[2] Tile_X9Y1_LUT4AB/N4BEG[3] Tile_X9Y1_LUT4AB/N4BEG[4]
+ Tile_X9Y1_LUT4AB/N4BEG[5] Tile_X9Y1_LUT4AB/N4BEG[6] Tile_X9Y1_LUT4AB/N4BEG[7] Tile_X9Y1_LUT4AB/N4BEG[8]
+ Tile_X9Y1_LUT4AB/N4BEG[9] Tile_X9Y1_LUT4AB/NN4BEG[0] Tile_X9Y1_LUT4AB/NN4BEG[10]
+ Tile_X9Y1_LUT4AB/NN4BEG[11] Tile_X9Y1_LUT4AB/NN4BEG[12] Tile_X9Y1_LUT4AB/NN4BEG[13]
+ Tile_X9Y1_LUT4AB/NN4BEG[14] Tile_X9Y1_LUT4AB/NN4BEG[15] Tile_X9Y1_LUT4AB/NN4BEG[1]
+ Tile_X9Y1_LUT4AB/NN4BEG[2] Tile_X9Y1_LUT4AB/NN4BEG[3] Tile_X9Y1_LUT4AB/NN4BEG[4]
+ Tile_X9Y1_LUT4AB/NN4BEG[5] Tile_X9Y1_LUT4AB/NN4BEG[6] Tile_X9Y1_LUT4AB/NN4BEG[7]
+ Tile_X9Y1_LUT4AB/NN4BEG[8] Tile_X9Y1_LUT4AB/NN4BEG[9] Tile_X9Y1_LUT4AB/S1END[0]
+ Tile_X9Y1_LUT4AB/S1END[1] Tile_X9Y1_LUT4AB/S1END[2] Tile_X9Y1_LUT4AB/S1END[3] Tile_X9Y1_LUT4AB/S2MID[0]
+ Tile_X9Y1_LUT4AB/S2MID[1] Tile_X9Y1_LUT4AB/S2MID[2] Tile_X9Y1_LUT4AB/S2MID[3] Tile_X9Y1_LUT4AB/S2MID[4]
+ Tile_X9Y1_LUT4AB/S2MID[5] Tile_X9Y1_LUT4AB/S2MID[6] Tile_X9Y1_LUT4AB/S2MID[7] Tile_X9Y1_LUT4AB/S2END[0]
+ Tile_X9Y1_LUT4AB/S2END[1] Tile_X9Y1_LUT4AB/S2END[2] Tile_X9Y1_LUT4AB/S2END[3] Tile_X9Y1_LUT4AB/S2END[4]
+ Tile_X9Y1_LUT4AB/S2END[5] Tile_X9Y1_LUT4AB/S2END[6] Tile_X9Y1_LUT4AB/S2END[7] Tile_X9Y1_LUT4AB/S4END[0]
+ Tile_X9Y1_LUT4AB/S4END[10] Tile_X9Y1_LUT4AB/S4END[11] Tile_X9Y1_LUT4AB/S4END[12]
+ Tile_X9Y1_LUT4AB/S4END[13] Tile_X9Y1_LUT4AB/S4END[14] Tile_X9Y1_LUT4AB/S4END[15]
+ Tile_X9Y1_LUT4AB/S4END[1] Tile_X9Y1_LUT4AB/S4END[2] Tile_X9Y1_LUT4AB/S4END[3] Tile_X9Y1_LUT4AB/S4END[4]
+ Tile_X9Y1_LUT4AB/S4END[5] Tile_X9Y1_LUT4AB/S4END[6] Tile_X9Y1_LUT4AB/S4END[7] Tile_X9Y1_LUT4AB/S4END[8]
+ Tile_X9Y1_LUT4AB/S4END[9] Tile_X9Y1_LUT4AB/SS4END[0] Tile_X9Y1_LUT4AB/SS4END[10]
+ Tile_X9Y1_LUT4AB/SS4END[11] Tile_X9Y1_LUT4AB/SS4END[12] Tile_X9Y1_LUT4AB/SS4END[13]
+ Tile_X9Y1_LUT4AB/SS4END[14] Tile_X9Y1_LUT4AB/SS4END[15] Tile_X9Y1_LUT4AB/SS4END[1]
+ Tile_X9Y1_LUT4AB/SS4END[2] Tile_X9Y1_LUT4AB/SS4END[3] Tile_X9Y1_LUT4AB/SS4END[4]
+ Tile_X9Y1_LUT4AB/SS4END[5] Tile_X9Y1_LUT4AB/SS4END[6] Tile_X9Y1_LUT4AB/SS4END[7]
+ Tile_X9Y1_LUT4AB/SS4END[8] Tile_X9Y1_LUT4AB/SS4END[9] Tile_X9Y1_LUT4AB/UserCLKo
+ Tile_X9Y0_N_term_single/UserCLKo VGND VPWR N_term_single
XTile_X3Y6_LUT4AB Tile_X3Y7_LUT4AB/Co Tile_X3Y6_LUT4AB/Co Tile_X3Y6_LUT4AB/E1BEG[0]
+ Tile_X3Y6_LUT4AB/E1BEG[1] Tile_X3Y6_LUT4AB/E1BEG[2] Tile_X3Y6_LUT4AB/E1BEG[3] Tile_X3Y6_LUT4AB/E1END[0]
+ Tile_X3Y6_LUT4AB/E1END[1] Tile_X3Y6_LUT4AB/E1END[2] Tile_X3Y6_LUT4AB/E1END[3] Tile_X3Y6_LUT4AB/E2BEG[0]
+ Tile_X3Y6_LUT4AB/E2BEG[1] Tile_X3Y6_LUT4AB/E2BEG[2] Tile_X3Y6_LUT4AB/E2BEG[3] Tile_X3Y6_LUT4AB/E2BEG[4]
+ Tile_X3Y6_LUT4AB/E2BEG[5] Tile_X3Y6_LUT4AB/E2BEG[6] Tile_X3Y6_LUT4AB/E2BEG[7] Tile_X4Y6_RegFile/E2END[0]
+ Tile_X4Y6_RegFile/E2END[1] Tile_X4Y6_RegFile/E2END[2] Tile_X4Y6_RegFile/E2END[3]
+ Tile_X4Y6_RegFile/E2END[4] Tile_X4Y6_RegFile/E2END[5] Tile_X4Y6_RegFile/E2END[6]
+ Tile_X4Y6_RegFile/E2END[7] Tile_X3Y6_LUT4AB/E2END[0] Tile_X3Y6_LUT4AB/E2END[1] Tile_X3Y6_LUT4AB/E2END[2]
+ Tile_X3Y6_LUT4AB/E2END[3] Tile_X3Y6_LUT4AB/E2END[4] Tile_X3Y6_LUT4AB/E2END[5] Tile_X3Y6_LUT4AB/E2END[6]
+ Tile_X3Y6_LUT4AB/E2END[7] Tile_X3Y6_LUT4AB/E2MID[0] Tile_X3Y6_LUT4AB/E2MID[1] Tile_X3Y6_LUT4AB/E2MID[2]
+ Tile_X3Y6_LUT4AB/E2MID[3] Tile_X3Y6_LUT4AB/E2MID[4] Tile_X3Y6_LUT4AB/E2MID[5] Tile_X3Y6_LUT4AB/E2MID[6]
+ Tile_X3Y6_LUT4AB/E2MID[7] Tile_X3Y6_LUT4AB/E6BEG[0] Tile_X3Y6_LUT4AB/E6BEG[10] Tile_X3Y6_LUT4AB/E6BEG[11]
+ Tile_X3Y6_LUT4AB/E6BEG[1] Tile_X3Y6_LUT4AB/E6BEG[2] Tile_X3Y6_LUT4AB/E6BEG[3] Tile_X3Y6_LUT4AB/E6BEG[4]
+ Tile_X3Y6_LUT4AB/E6BEG[5] Tile_X3Y6_LUT4AB/E6BEG[6] Tile_X3Y6_LUT4AB/E6BEG[7] Tile_X3Y6_LUT4AB/E6BEG[8]
+ Tile_X3Y6_LUT4AB/E6BEG[9] Tile_X3Y6_LUT4AB/E6END[0] Tile_X3Y6_LUT4AB/E6END[10] Tile_X3Y6_LUT4AB/E6END[11]
+ Tile_X3Y6_LUT4AB/E6END[1] Tile_X3Y6_LUT4AB/E6END[2] Tile_X3Y6_LUT4AB/E6END[3] Tile_X3Y6_LUT4AB/E6END[4]
+ Tile_X3Y6_LUT4AB/E6END[5] Tile_X3Y6_LUT4AB/E6END[6] Tile_X3Y6_LUT4AB/E6END[7] Tile_X3Y6_LUT4AB/E6END[8]
+ Tile_X3Y6_LUT4AB/E6END[9] Tile_X3Y6_LUT4AB/EE4BEG[0] Tile_X3Y6_LUT4AB/EE4BEG[10]
+ Tile_X3Y6_LUT4AB/EE4BEG[11] Tile_X3Y6_LUT4AB/EE4BEG[12] Tile_X3Y6_LUT4AB/EE4BEG[13]
+ Tile_X3Y6_LUT4AB/EE4BEG[14] Tile_X3Y6_LUT4AB/EE4BEG[15] Tile_X3Y6_LUT4AB/EE4BEG[1]
+ Tile_X3Y6_LUT4AB/EE4BEG[2] Tile_X3Y6_LUT4AB/EE4BEG[3] Tile_X3Y6_LUT4AB/EE4BEG[4]
+ Tile_X3Y6_LUT4AB/EE4BEG[5] Tile_X3Y6_LUT4AB/EE4BEG[6] Tile_X3Y6_LUT4AB/EE4BEG[7]
+ Tile_X3Y6_LUT4AB/EE4BEG[8] Tile_X3Y6_LUT4AB/EE4BEG[9] Tile_X3Y6_LUT4AB/EE4END[0]
+ Tile_X3Y6_LUT4AB/EE4END[10] Tile_X3Y6_LUT4AB/EE4END[11] Tile_X3Y6_LUT4AB/EE4END[12]
+ Tile_X3Y6_LUT4AB/EE4END[13] Tile_X3Y6_LUT4AB/EE4END[14] Tile_X3Y6_LUT4AB/EE4END[15]
+ Tile_X3Y6_LUT4AB/EE4END[1] Tile_X3Y6_LUT4AB/EE4END[2] Tile_X3Y6_LUT4AB/EE4END[3]
+ Tile_X3Y6_LUT4AB/EE4END[4] Tile_X3Y6_LUT4AB/EE4END[5] Tile_X3Y6_LUT4AB/EE4END[6]
+ Tile_X3Y6_LUT4AB/EE4END[7] Tile_X3Y6_LUT4AB/EE4END[8] Tile_X3Y6_LUT4AB/EE4END[9]
+ Tile_X3Y6_LUT4AB/FrameData[0] Tile_X3Y6_LUT4AB/FrameData[10] Tile_X3Y6_LUT4AB/FrameData[11]
+ Tile_X3Y6_LUT4AB/FrameData[12] Tile_X3Y6_LUT4AB/FrameData[13] Tile_X3Y6_LUT4AB/FrameData[14]
+ Tile_X3Y6_LUT4AB/FrameData[15] Tile_X3Y6_LUT4AB/FrameData[16] Tile_X3Y6_LUT4AB/FrameData[17]
+ Tile_X3Y6_LUT4AB/FrameData[18] Tile_X3Y6_LUT4AB/FrameData[19] Tile_X3Y6_LUT4AB/FrameData[1]
+ Tile_X3Y6_LUT4AB/FrameData[20] Tile_X3Y6_LUT4AB/FrameData[21] Tile_X3Y6_LUT4AB/FrameData[22]
+ Tile_X3Y6_LUT4AB/FrameData[23] Tile_X3Y6_LUT4AB/FrameData[24] Tile_X3Y6_LUT4AB/FrameData[25]
+ Tile_X3Y6_LUT4AB/FrameData[26] Tile_X3Y6_LUT4AB/FrameData[27] Tile_X3Y6_LUT4AB/FrameData[28]
+ Tile_X3Y6_LUT4AB/FrameData[29] Tile_X3Y6_LUT4AB/FrameData[2] Tile_X3Y6_LUT4AB/FrameData[30]
+ Tile_X3Y6_LUT4AB/FrameData[31] Tile_X3Y6_LUT4AB/FrameData[3] Tile_X3Y6_LUT4AB/FrameData[4]
+ Tile_X3Y6_LUT4AB/FrameData[5] Tile_X3Y6_LUT4AB/FrameData[6] Tile_X3Y6_LUT4AB/FrameData[7]
+ Tile_X3Y6_LUT4AB/FrameData[8] Tile_X3Y6_LUT4AB/FrameData[9] Tile_X4Y6_RegFile/FrameData[0]
+ Tile_X4Y6_RegFile/FrameData[10] Tile_X4Y6_RegFile/FrameData[11] Tile_X4Y6_RegFile/FrameData[12]
+ Tile_X4Y6_RegFile/FrameData[13] Tile_X4Y6_RegFile/FrameData[14] Tile_X4Y6_RegFile/FrameData[15]
+ Tile_X4Y6_RegFile/FrameData[16] Tile_X4Y6_RegFile/FrameData[17] Tile_X4Y6_RegFile/FrameData[18]
+ Tile_X4Y6_RegFile/FrameData[19] Tile_X4Y6_RegFile/FrameData[1] Tile_X4Y6_RegFile/FrameData[20]
+ Tile_X4Y6_RegFile/FrameData[21] Tile_X4Y6_RegFile/FrameData[22] Tile_X4Y6_RegFile/FrameData[23]
+ Tile_X4Y6_RegFile/FrameData[24] Tile_X4Y6_RegFile/FrameData[25] Tile_X4Y6_RegFile/FrameData[26]
+ Tile_X4Y6_RegFile/FrameData[27] Tile_X4Y6_RegFile/FrameData[28] Tile_X4Y6_RegFile/FrameData[29]
+ Tile_X4Y6_RegFile/FrameData[2] Tile_X4Y6_RegFile/FrameData[30] Tile_X4Y6_RegFile/FrameData[31]
+ Tile_X4Y6_RegFile/FrameData[3] Tile_X4Y6_RegFile/FrameData[4] Tile_X4Y6_RegFile/FrameData[5]
+ Tile_X4Y6_RegFile/FrameData[6] Tile_X4Y6_RegFile/FrameData[7] Tile_X4Y6_RegFile/FrameData[8]
+ Tile_X4Y6_RegFile/FrameData[9] Tile_X3Y6_LUT4AB/FrameStrobe[0] Tile_X3Y6_LUT4AB/FrameStrobe[10]
+ Tile_X3Y6_LUT4AB/FrameStrobe[11] Tile_X3Y6_LUT4AB/FrameStrobe[12] Tile_X3Y6_LUT4AB/FrameStrobe[13]
+ Tile_X3Y6_LUT4AB/FrameStrobe[14] Tile_X3Y6_LUT4AB/FrameStrobe[15] Tile_X3Y6_LUT4AB/FrameStrobe[16]
+ Tile_X3Y6_LUT4AB/FrameStrobe[17] Tile_X3Y6_LUT4AB/FrameStrobe[18] Tile_X3Y6_LUT4AB/FrameStrobe[19]
+ Tile_X3Y6_LUT4AB/FrameStrobe[1] Tile_X3Y6_LUT4AB/FrameStrobe[2] Tile_X3Y6_LUT4AB/FrameStrobe[3]
+ Tile_X3Y6_LUT4AB/FrameStrobe[4] Tile_X3Y6_LUT4AB/FrameStrobe[5] Tile_X3Y6_LUT4AB/FrameStrobe[6]
+ Tile_X3Y6_LUT4AB/FrameStrobe[7] Tile_X3Y6_LUT4AB/FrameStrobe[8] Tile_X3Y6_LUT4AB/FrameStrobe[9]
+ Tile_X3Y5_LUT4AB/FrameStrobe[0] Tile_X3Y5_LUT4AB/FrameStrobe[10] Tile_X3Y5_LUT4AB/FrameStrobe[11]
+ Tile_X3Y5_LUT4AB/FrameStrobe[12] Tile_X3Y5_LUT4AB/FrameStrobe[13] Tile_X3Y5_LUT4AB/FrameStrobe[14]
+ Tile_X3Y5_LUT4AB/FrameStrobe[15] Tile_X3Y5_LUT4AB/FrameStrobe[16] Tile_X3Y5_LUT4AB/FrameStrobe[17]
+ Tile_X3Y5_LUT4AB/FrameStrobe[18] Tile_X3Y5_LUT4AB/FrameStrobe[19] Tile_X3Y5_LUT4AB/FrameStrobe[1]
+ Tile_X3Y5_LUT4AB/FrameStrobe[2] Tile_X3Y5_LUT4AB/FrameStrobe[3] Tile_X3Y5_LUT4AB/FrameStrobe[4]
+ Tile_X3Y5_LUT4AB/FrameStrobe[5] Tile_X3Y5_LUT4AB/FrameStrobe[6] Tile_X3Y5_LUT4AB/FrameStrobe[7]
+ Tile_X3Y5_LUT4AB/FrameStrobe[8] Tile_X3Y5_LUT4AB/FrameStrobe[9] Tile_X3Y6_LUT4AB/N1BEG[0]
+ Tile_X3Y6_LUT4AB/N1BEG[1] Tile_X3Y6_LUT4AB/N1BEG[2] Tile_X3Y6_LUT4AB/N1BEG[3] Tile_X3Y7_LUT4AB/N1BEG[0]
+ Tile_X3Y7_LUT4AB/N1BEG[1] Tile_X3Y7_LUT4AB/N1BEG[2] Tile_X3Y7_LUT4AB/N1BEG[3] Tile_X3Y6_LUT4AB/N2BEG[0]
+ Tile_X3Y6_LUT4AB/N2BEG[1] Tile_X3Y6_LUT4AB/N2BEG[2] Tile_X3Y6_LUT4AB/N2BEG[3] Tile_X3Y6_LUT4AB/N2BEG[4]
+ Tile_X3Y6_LUT4AB/N2BEG[5] Tile_X3Y6_LUT4AB/N2BEG[6] Tile_X3Y6_LUT4AB/N2BEG[7] Tile_X3Y5_LUT4AB/N2END[0]
+ Tile_X3Y5_LUT4AB/N2END[1] Tile_X3Y5_LUT4AB/N2END[2] Tile_X3Y5_LUT4AB/N2END[3] Tile_X3Y5_LUT4AB/N2END[4]
+ Tile_X3Y5_LUT4AB/N2END[5] Tile_X3Y5_LUT4AB/N2END[6] Tile_X3Y5_LUT4AB/N2END[7] Tile_X3Y6_LUT4AB/N2END[0]
+ Tile_X3Y6_LUT4AB/N2END[1] Tile_X3Y6_LUT4AB/N2END[2] Tile_X3Y6_LUT4AB/N2END[3] Tile_X3Y6_LUT4AB/N2END[4]
+ Tile_X3Y6_LUT4AB/N2END[5] Tile_X3Y6_LUT4AB/N2END[6] Tile_X3Y6_LUT4AB/N2END[7] Tile_X3Y7_LUT4AB/N2BEG[0]
+ Tile_X3Y7_LUT4AB/N2BEG[1] Tile_X3Y7_LUT4AB/N2BEG[2] Tile_X3Y7_LUT4AB/N2BEG[3] Tile_X3Y7_LUT4AB/N2BEG[4]
+ Tile_X3Y7_LUT4AB/N2BEG[5] Tile_X3Y7_LUT4AB/N2BEG[6] Tile_X3Y7_LUT4AB/N2BEG[7] Tile_X3Y6_LUT4AB/N4BEG[0]
+ Tile_X3Y6_LUT4AB/N4BEG[10] Tile_X3Y6_LUT4AB/N4BEG[11] Tile_X3Y6_LUT4AB/N4BEG[12]
+ Tile_X3Y6_LUT4AB/N4BEG[13] Tile_X3Y6_LUT4AB/N4BEG[14] Tile_X3Y6_LUT4AB/N4BEG[15]
+ Tile_X3Y6_LUT4AB/N4BEG[1] Tile_X3Y6_LUT4AB/N4BEG[2] Tile_X3Y6_LUT4AB/N4BEG[3] Tile_X3Y6_LUT4AB/N4BEG[4]
+ Tile_X3Y6_LUT4AB/N4BEG[5] Tile_X3Y6_LUT4AB/N4BEG[6] Tile_X3Y6_LUT4AB/N4BEG[7] Tile_X3Y6_LUT4AB/N4BEG[8]
+ Tile_X3Y6_LUT4AB/N4BEG[9] Tile_X3Y7_LUT4AB/N4BEG[0] Tile_X3Y7_LUT4AB/N4BEG[10] Tile_X3Y7_LUT4AB/N4BEG[11]
+ Tile_X3Y7_LUT4AB/N4BEG[12] Tile_X3Y7_LUT4AB/N4BEG[13] Tile_X3Y7_LUT4AB/N4BEG[14]
+ Tile_X3Y7_LUT4AB/N4BEG[15] Tile_X3Y7_LUT4AB/N4BEG[1] Tile_X3Y7_LUT4AB/N4BEG[2] Tile_X3Y7_LUT4AB/N4BEG[3]
+ Tile_X3Y7_LUT4AB/N4BEG[4] Tile_X3Y7_LUT4AB/N4BEG[5] Tile_X3Y7_LUT4AB/N4BEG[6] Tile_X3Y7_LUT4AB/N4BEG[7]
+ Tile_X3Y7_LUT4AB/N4BEG[8] Tile_X3Y7_LUT4AB/N4BEG[9] Tile_X3Y6_LUT4AB/NN4BEG[0] Tile_X3Y6_LUT4AB/NN4BEG[10]
+ Tile_X3Y6_LUT4AB/NN4BEG[11] Tile_X3Y6_LUT4AB/NN4BEG[12] Tile_X3Y6_LUT4AB/NN4BEG[13]
+ Tile_X3Y6_LUT4AB/NN4BEG[14] Tile_X3Y6_LUT4AB/NN4BEG[15] Tile_X3Y6_LUT4AB/NN4BEG[1]
+ Tile_X3Y6_LUT4AB/NN4BEG[2] Tile_X3Y6_LUT4AB/NN4BEG[3] Tile_X3Y6_LUT4AB/NN4BEG[4]
+ Tile_X3Y6_LUT4AB/NN4BEG[5] Tile_X3Y6_LUT4AB/NN4BEG[6] Tile_X3Y6_LUT4AB/NN4BEG[7]
+ Tile_X3Y6_LUT4AB/NN4BEG[8] Tile_X3Y6_LUT4AB/NN4BEG[9] Tile_X3Y7_LUT4AB/NN4BEG[0]
+ Tile_X3Y7_LUT4AB/NN4BEG[10] Tile_X3Y7_LUT4AB/NN4BEG[11] Tile_X3Y7_LUT4AB/NN4BEG[12]
+ Tile_X3Y7_LUT4AB/NN4BEG[13] Tile_X3Y7_LUT4AB/NN4BEG[14] Tile_X3Y7_LUT4AB/NN4BEG[15]
+ Tile_X3Y7_LUT4AB/NN4BEG[1] Tile_X3Y7_LUT4AB/NN4BEG[2] Tile_X3Y7_LUT4AB/NN4BEG[3]
+ Tile_X3Y7_LUT4AB/NN4BEG[4] Tile_X3Y7_LUT4AB/NN4BEG[5] Tile_X3Y7_LUT4AB/NN4BEG[6]
+ Tile_X3Y7_LUT4AB/NN4BEG[7] Tile_X3Y7_LUT4AB/NN4BEG[8] Tile_X3Y7_LUT4AB/NN4BEG[9]
+ Tile_X3Y7_LUT4AB/S1END[0] Tile_X3Y7_LUT4AB/S1END[1] Tile_X3Y7_LUT4AB/S1END[2] Tile_X3Y7_LUT4AB/S1END[3]
+ Tile_X3Y6_LUT4AB/S1END[0] Tile_X3Y6_LUT4AB/S1END[1] Tile_X3Y6_LUT4AB/S1END[2] Tile_X3Y6_LUT4AB/S1END[3]
+ Tile_X3Y7_LUT4AB/S2MID[0] Tile_X3Y7_LUT4AB/S2MID[1] Tile_X3Y7_LUT4AB/S2MID[2] Tile_X3Y7_LUT4AB/S2MID[3]
+ Tile_X3Y7_LUT4AB/S2MID[4] Tile_X3Y7_LUT4AB/S2MID[5] Tile_X3Y7_LUT4AB/S2MID[6] Tile_X3Y7_LUT4AB/S2MID[7]
+ Tile_X3Y7_LUT4AB/S2END[0] Tile_X3Y7_LUT4AB/S2END[1] Tile_X3Y7_LUT4AB/S2END[2] Tile_X3Y7_LUT4AB/S2END[3]
+ Tile_X3Y7_LUT4AB/S2END[4] Tile_X3Y7_LUT4AB/S2END[5] Tile_X3Y7_LUT4AB/S2END[6] Tile_X3Y7_LUT4AB/S2END[7]
+ Tile_X3Y6_LUT4AB/S2END[0] Tile_X3Y6_LUT4AB/S2END[1] Tile_X3Y6_LUT4AB/S2END[2] Tile_X3Y6_LUT4AB/S2END[3]
+ Tile_X3Y6_LUT4AB/S2END[4] Tile_X3Y6_LUT4AB/S2END[5] Tile_X3Y6_LUT4AB/S2END[6] Tile_X3Y6_LUT4AB/S2END[7]
+ Tile_X3Y6_LUT4AB/S2MID[0] Tile_X3Y6_LUT4AB/S2MID[1] Tile_X3Y6_LUT4AB/S2MID[2] Tile_X3Y6_LUT4AB/S2MID[3]
+ Tile_X3Y6_LUT4AB/S2MID[4] Tile_X3Y6_LUT4AB/S2MID[5] Tile_X3Y6_LUT4AB/S2MID[6] Tile_X3Y6_LUT4AB/S2MID[7]
+ Tile_X3Y7_LUT4AB/S4END[0] Tile_X3Y7_LUT4AB/S4END[10] Tile_X3Y7_LUT4AB/S4END[11]
+ Tile_X3Y7_LUT4AB/S4END[12] Tile_X3Y7_LUT4AB/S4END[13] Tile_X3Y7_LUT4AB/S4END[14]
+ Tile_X3Y7_LUT4AB/S4END[15] Tile_X3Y7_LUT4AB/S4END[1] Tile_X3Y7_LUT4AB/S4END[2] Tile_X3Y7_LUT4AB/S4END[3]
+ Tile_X3Y7_LUT4AB/S4END[4] Tile_X3Y7_LUT4AB/S4END[5] Tile_X3Y7_LUT4AB/S4END[6] Tile_X3Y7_LUT4AB/S4END[7]
+ Tile_X3Y7_LUT4AB/S4END[8] Tile_X3Y7_LUT4AB/S4END[9] Tile_X3Y6_LUT4AB/S4END[0] Tile_X3Y6_LUT4AB/S4END[10]
+ Tile_X3Y6_LUT4AB/S4END[11] Tile_X3Y6_LUT4AB/S4END[12] Tile_X3Y6_LUT4AB/S4END[13]
+ Tile_X3Y6_LUT4AB/S4END[14] Tile_X3Y6_LUT4AB/S4END[15] Tile_X3Y6_LUT4AB/S4END[1]
+ Tile_X3Y6_LUT4AB/S4END[2] Tile_X3Y6_LUT4AB/S4END[3] Tile_X3Y6_LUT4AB/S4END[4] Tile_X3Y6_LUT4AB/S4END[5]
+ Tile_X3Y6_LUT4AB/S4END[6] Tile_X3Y6_LUT4AB/S4END[7] Tile_X3Y6_LUT4AB/S4END[8] Tile_X3Y6_LUT4AB/S4END[9]
+ Tile_X3Y7_LUT4AB/SS4END[0] Tile_X3Y7_LUT4AB/SS4END[10] Tile_X3Y7_LUT4AB/SS4END[11]
+ Tile_X3Y7_LUT4AB/SS4END[12] Tile_X3Y7_LUT4AB/SS4END[13] Tile_X3Y7_LUT4AB/SS4END[14]
+ Tile_X3Y7_LUT4AB/SS4END[15] Tile_X3Y7_LUT4AB/SS4END[1] Tile_X3Y7_LUT4AB/SS4END[2]
+ Tile_X3Y7_LUT4AB/SS4END[3] Tile_X3Y7_LUT4AB/SS4END[4] Tile_X3Y7_LUT4AB/SS4END[5]
+ Tile_X3Y7_LUT4AB/SS4END[6] Tile_X3Y7_LUT4AB/SS4END[7] Tile_X3Y7_LUT4AB/SS4END[8]
+ Tile_X3Y7_LUT4AB/SS4END[9] Tile_X3Y6_LUT4AB/SS4END[0] Tile_X3Y6_LUT4AB/SS4END[10]
+ Tile_X3Y6_LUT4AB/SS4END[11] Tile_X3Y6_LUT4AB/SS4END[12] Tile_X3Y6_LUT4AB/SS4END[13]
+ Tile_X3Y6_LUT4AB/SS4END[14] Tile_X3Y6_LUT4AB/SS4END[15] Tile_X3Y6_LUT4AB/SS4END[1]
+ Tile_X3Y6_LUT4AB/SS4END[2] Tile_X3Y6_LUT4AB/SS4END[3] Tile_X3Y6_LUT4AB/SS4END[4]
+ Tile_X3Y6_LUT4AB/SS4END[5] Tile_X3Y6_LUT4AB/SS4END[6] Tile_X3Y6_LUT4AB/SS4END[7]
+ Tile_X3Y6_LUT4AB/SS4END[8] Tile_X3Y6_LUT4AB/SS4END[9] Tile_X3Y6_LUT4AB/UserCLK Tile_X3Y5_LUT4AB/UserCLK
+ VGND VPWR Tile_X3Y6_LUT4AB/W1BEG[0] Tile_X3Y6_LUT4AB/W1BEG[1] Tile_X3Y6_LUT4AB/W1BEG[2]
+ Tile_X3Y6_LUT4AB/W1BEG[3] Tile_X3Y6_LUT4AB/W1END[0] Tile_X3Y6_LUT4AB/W1END[1] Tile_X3Y6_LUT4AB/W1END[2]
+ Tile_X3Y6_LUT4AB/W1END[3] Tile_X3Y6_LUT4AB/W2BEG[0] Tile_X3Y6_LUT4AB/W2BEG[1] Tile_X3Y6_LUT4AB/W2BEG[2]
+ Tile_X3Y6_LUT4AB/W2BEG[3] Tile_X3Y6_LUT4AB/W2BEG[4] Tile_X3Y6_LUT4AB/W2BEG[5] Tile_X3Y6_LUT4AB/W2BEG[6]
+ Tile_X3Y6_LUT4AB/W2BEG[7] Tile_X2Y6_LUT4AB/W2END[0] Tile_X2Y6_LUT4AB/W2END[1] Tile_X2Y6_LUT4AB/W2END[2]
+ Tile_X2Y6_LUT4AB/W2END[3] Tile_X2Y6_LUT4AB/W2END[4] Tile_X2Y6_LUT4AB/W2END[5] Tile_X2Y6_LUT4AB/W2END[6]
+ Tile_X2Y6_LUT4AB/W2END[7] Tile_X3Y6_LUT4AB/W2END[0] Tile_X3Y6_LUT4AB/W2END[1] Tile_X3Y6_LUT4AB/W2END[2]
+ Tile_X3Y6_LUT4AB/W2END[3] Tile_X3Y6_LUT4AB/W2END[4] Tile_X3Y6_LUT4AB/W2END[5] Tile_X3Y6_LUT4AB/W2END[6]
+ Tile_X3Y6_LUT4AB/W2END[7] Tile_X3Y6_LUT4AB/W2MID[0] Tile_X3Y6_LUT4AB/W2MID[1] Tile_X3Y6_LUT4AB/W2MID[2]
+ Tile_X3Y6_LUT4AB/W2MID[3] Tile_X3Y6_LUT4AB/W2MID[4] Tile_X3Y6_LUT4AB/W2MID[5] Tile_X3Y6_LUT4AB/W2MID[6]
+ Tile_X3Y6_LUT4AB/W2MID[7] Tile_X3Y6_LUT4AB/W6BEG[0] Tile_X3Y6_LUT4AB/W6BEG[10] Tile_X3Y6_LUT4AB/W6BEG[11]
+ Tile_X3Y6_LUT4AB/W6BEG[1] Tile_X3Y6_LUT4AB/W6BEG[2] Tile_X3Y6_LUT4AB/W6BEG[3] Tile_X3Y6_LUT4AB/W6BEG[4]
+ Tile_X3Y6_LUT4AB/W6BEG[5] Tile_X3Y6_LUT4AB/W6BEG[6] Tile_X3Y6_LUT4AB/W6BEG[7] Tile_X3Y6_LUT4AB/W6BEG[8]
+ Tile_X3Y6_LUT4AB/W6BEG[9] Tile_X3Y6_LUT4AB/W6END[0] Tile_X3Y6_LUT4AB/W6END[10] Tile_X3Y6_LUT4AB/W6END[11]
+ Tile_X3Y6_LUT4AB/W6END[1] Tile_X3Y6_LUT4AB/W6END[2] Tile_X3Y6_LUT4AB/W6END[3] Tile_X3Y6_LUT4AB/W6END[4]
+ Tile_X3Y6_LUT4AB/W6END[5] Tile_X3Y6_LUT4AB/W6END[6] Tile_X3Y6_LUT4AB/W6END[7] Tile_X3Y6_LUT4AB/W6END[8]
+ Tile_X3Y6_LUT4AB/W6END[9] Tile_X3Y6_LUT4AB/WW4BEG[0] Tile_X3Y6_LUT4AB/WW4BEG[10]
+ Tile_X3Y6_LUT4AB/WW4BEG[11] Tile_X3Y6_LUT4AB/WW4BEG[12] Tile_X3Y6_LUT4AB/WW4BEG[13]
+ Tile_X3Y6_LUT4AB/WW4BEG[14] Tile_X3Y6_LUT4AB/WW4BEG[15] Tile_X3Y6_LUT4AB/WW4BEG[1]
+ Tile_X3Y6_LUT4AB/WW4BEG[2] Tile_X3Y6_LUT4AB/WW4BEG[3] Tile_X3Y6_LUT4AB/WW4BEG[4]
+ Tile_X3Y6_LUT4AB/WW4BEG[5] Tile_X3Y6_LUT4AB/WW4BEG[6] Tile_X3Y6_LUT4AB/WW4BEG[7]
+ Tile_X3Y6_LUT4AB/WW4BEG[8] Tile_X3Y6_LUT4AB/WW4BEG[9] Tile_X3Y6_LUT4AB/WW4END[0]
+ Tile_X3Y6_LUT4AB/WW4END[10] Tile_X3Y6_LUT4AB/WW4END[11] Tile_X3Y6_LUT4AB/WW4END[12]
+ Tile_X3Y6_LUT4AB/WW4END[13] Tile_X3Y6_LUT4AB/WW4END[14] Tile_X3Y6_LUT4AB/WW4END[15]
+ Tile_X3Y6_LUT4AB/WW4END[1] Tile_X3Y6_LUT4AB/WW4END[2] Tile_X3Y6_LUT4AB/WW4END[3]
+ Tile_X3Y6_LUT4AB/WW4END[4] Tile_X3Y6_LUT4AB/WW4END[5] Tile_X3Y6_LUT4AB/WW4END[6]
+ Tile_X3Y6_LUT4AB/WW4END[7] Tile_X3Y6_LUT4AB/WW4END[8] Tile_X3Y6_LUT4AB/WW4END[9]
+ LUT4AB
XTile_X4Y14_RegFile Tile_X5Y14_LUT4AB/E1END[0] Tile_X5Y14_LUT4AB/E1END[1] Tile_X5Y14_LUT4AB/E1END[2]
+ Tile_X5Y14_LUT4AB/E1END[3] Tile_X3Y14_LUT4AB/E1BEG[0] Tile_X3Y14_LUT4AB/E1BEG[1]
+ Tile_X3Y14_LUT4AB/E1BEG[2] Tile_X3Y14_LUT4AB/E1BEG[3] Tile_X5Y14_LUT4AB/E2MID[0]
+ Tile_X5Y14_LUT4AB/E2MID[1] Tile_X5Y14_LUT4AB/E2MID[2] Tile_X5Y14_LUT4AB/E2MID[3]
+ Tile_X5Y14_LUT4AB/E2MID[4] Tile_X5Y14_LUT4AB/E2MID[5] Tile_X5Y14_LUT4AB/E2MID[6]
+ Tile_X5Y14_LUT4AB/E2MID[7] Tile_X5Y14_LUT4AB/E2END[0] Tile_X5Y14_LUT4AB/E2END[1]
+ Tile_X5Y14_LUT4AB/E2END[2] Tile_X5Y14_LUT4AB/E2END[3] Tile_X5Y14_LUT4AB/E2END[4]
+ Tile_X5Y14_LUT4AB/E2END[5] Tile_X5Y14_LUT4AB/E2END[6] Tile_X5Y14_LUT4AB/E2END[7]
+ Tile_X4Y14_RegFile/E2END[0] Tile_X4Y14_RegFile/E2END[1] Tile_X4Y14_RegFile/E2END[2]
+ Tile_X4Y14_RegFile/E2END[3] Tile_X4Y14_RegFile/E2END[4] Tile_X4Y14_RegFile/E2END[5]
+ Tile_X4Y14_RegFile/E2END[6] Tile_X4Y14_RegFile/E2END[7] Tile_X3Y14_LUT4AB/E2BEG[0]
+ Tile_X3Y14_LUT4AB/E2BEG[1] Tile_X3Y14_LUT4AB/E2BEG[2] Tile_X3Y14_LUT4AB/E2BEG[3]
+ Tile_X3Y14_LUT4AB/E2BEG[4] Tile_X3Y14_LUT4AB/E2BEG[5] Tile_X3Y14_LUT4AB/E2BEG[6]
+ Tile_X3Y14_LUT4AB/E2BEG[7] Tile_X5Y14_LUT4AB/E6END[0] Tile_X5Y14_LUT4AB/E6END[10]
+ Tile_X5Y14_LUT4AB/E6END[11] Tile_X5Y14_LUT4AB/E6END[1] Tile_X5Y14_LUT4AB/E6END[2]
+ Tile_X5Y14_LUT4AB/E6END[3] Tile_X5Y14_LUT4AB/E6END[4] Tile_X5Y14_LUT4AB/E6END[5]
+ Tile_X5Y14_LUT4AB/E6END[6] Tile_X5Y14_LUT4AB/E6END[7] Tile_X5Y14_LUT4AB/E6END[8]
+ Tile_X5Y14_LUT4AB/E6END[9] Tile_X3Y14_LUT4AB/E6BEG[0] Tile_X3Y14_LUT4AB/E6BEG[10]
+ Tile_X3Y14_LUT4AB/E6BEG[11] Tile_X3Y14_LUT4AB/E6BEG[1] Tile_X3Y14_LUT4AB/E6BEG[2]
+ Tile_X3Y14_LUT4AB/E6BEG[3] Tile_X3Y14_LUT4AB/E6BEG[4] Tile_X3Y14_LUT4AB/E6BEG[5]
+ Tile_X3Y14_LUT4AB/E6BEG[6] Tile_X3Y14_LUT4AB/E6BEG[7] Tile_X3Y14_LUT4AB/E6BEG[8]
+ Tile_X3Y14_LUT4AB/E6BEG[9] Tile_X5Y14_LUT4AB/EE4END[0] Tile_X5Y14_LUT4AB/EE4END[10]
+ Tile_X5Y14_LUT4AB/EE4END[11] Tile_X5Y14_LUT4AB/EE4END[12] Tile_X5Y14_LUT4AB/EE4END[13]
+ Tile_X5Y14_LUT4AB/EE4END[14] Tile_X5Y14_LUT4AB/EE4END[15] Tile_X5Y14_LUT4AB/EE4END[1]
+ Tile_X5Y14_LUT4AB/EE4END[2] Tile_X5Y14_LUT4AB/EE4END[3] Tile_X5Y14_LUT4AB/EE4END[4]
+ Tile_X5Y14_LUT4AB/EE4END[5] Tile_X5Y14_LUT4AB/EE4END[6] Tile_X5Y14_LUT4AB/EE4END[7]
+ Tile_X5Y14_LUT4AB/EE4END[8] Tile_X5Y14_LUT4AB/EE4END[9] Tile_X3Y14_LUT4AB/EE4BEG[0]
+ Tile_X3Y14_LUT4AB/EE4BEG[10] Tile_X3Y14_LUT4AB/EE4BEG[11] Tile_X3Y14_LUT4AB/EE4BEG[12]
+ Tile_X3Y14_LUT4AB/EE4BEG[13] Tile_X3Y14_LUT4AB/EE4BEG[14] Tile_X3Y14_LUT4AB/EE4BEG[15]
+ Tile_X3Y14_LUT4AB/EE4BEG[1] Tile_X3Y14_LUT4AB/EE4BEG[2] Tile_X3Y14_LUT4AB/EE4BEG[3]
+ Tile_X3Y14_LUT4AB/EE4BEG[4] Tile_X3Y14_LUT4AB/EE4BEG[5] Tile_X3Y14_LUT4AB/EE4BEG[6]
+ Tile_X3Y14_LUT4AB/EE4BEG[7] Tile_X3Y14_LUT4AB/EE4BEG[8] Tile_X3Y14_LUT4AB/EE4BEG[9]
+ Tile_X4Y14_RegFile/FrameData[0] Tile_X4Y14_RegFile/FrameData[10] Tile_X4Y14_RegFile/FrameData[11]
+ Tile_X4Y14_RegFile/FrameData[12] Tile_X4Y14_RegFile/FrameData[13] Tile_X4Y14_RegFile/FrameData[14]
+ Tile_X4Y14_RegFile/FrameData[15] Tile_X4Y14_RegFile/FrameData[16] Tile_X4Y14_RegFile/FrameData[17]
+ Tile_X4Y14_RegFile/FrameData[18] Tile_X4Y14_RegFile/FrameData[19] Tile_X4Y14_RegFile/FrameData[1]
+ Tile_X4Y14_RegFile/FrameData[20] Tile_X4Y14_RegFile/FrameData[21] Tile_X4Y14_RegFile/FrameData[22]
+ Tile_X4Y14_RegFile/FrameData[23] Tile_X4Y14_RegFile/FrameData[24] Tile_X4Y14_RegFile/FrameData[25]
+ Tile_X4Y14_RegFile/FrameData[26] Tile_X4Y14_RegFile/FrameData[27] Tile_X4Y14_RegFile/FrameData[28]
+ Tile_X4Y14_RegFile/FrameData[29] Tile_X4Y14_RegFile/FrameData[2] Tile_X4Y14_RegFile/FrameData[30]
+ Tile_X4Y14_RegFile/FrameData[31] Tile_X4Y14_RegFile/FrameData[3] Tile_X4Y14_RegFile/FrameData[4]
+ Tile_X4Y14_RegFile/FrameData[5] Tile_X4Y14_RegFile/FrameData[6] Tile_X4Y14_RegFile/FrameData[7]
+ Tile_X4Y14_RegFile/FrameData[8] Tile_X4Y14_RegFile/FrameData[9] Tile_X5Y14_LUT4AB/FrameData[0]
+ Tile_X5Y14_LUT4AB/FrameData[10] Tile_X5Y14_LUT4AB/FrameData[11] Tile_X5Y14_LUT4AB/FrameData[12]
+ Tile_X5Y14_LUT4AB/FrameData[13] Tile_X5Y14_LUT4AB/FrameData[14] Tile_X5Y14_LUT4AB/FrameData[15]
+ Tile_X5Y14_LUT4AB/FrameData[16] Tile_X5Y14_LUT4AB/FrameData[17] Tile_X5Y14_LUT4AB/FrameData[18]
+ Tile_X5Y14_LUT4AB/FrameData[19] Tile_X5Y14_LUT4AB/FrameData[1] Tile_X5Y14_LUT4AB/FrameData[20]
+ Tile_X5Y14_LUT4AB/FrameData[21] Tile_X5Y14_LUT4AB/FrameData[22] Tile_X5Y14_LUT4AB/FrameData[23]
+ Tile_X5Y14_LUT4AB/FrameData[24] Tile_X5Y14_LUT4AB/FrameData[25] Tile_X5Y14_LUT4AB/FrameData[26]
+ Tile_X5Y14_LUT4AB/FrameData[27] Tile_X5Y14_LUT4AB/FrameData[28] Tile_X5Y14_LUT4AB/FrameData[29]
+ Tile_X5Y14_LUT4AB/FrameData[2] Tile_X5Y14_LUT4AB/FrameData[30] Tile_X5Y14_LUT4AB/FrameData[31]
+ Tile_X5Y14_LUT4AB/FrameData[3] Tile_X5Y14_LUT4AB/FrameData[4] Tile_X5Y14_LUT4AB/FrameData[5]
+ Tile_X5Y14_LUT4AB/FrameData[6] Tile_X5Y14_LUT4AB/FrameData[7] Tile_X5Y14_LUT4AB/FrameData[8]
+ Tile_X5Y14_LUT4AB/FrameData[9] Tile_X4Y14_RegFile/FrameStrobe[0] Tile_X4Y14_RegFile/FrameStrobe[10]
+ Tile_X4Y14_RegFile/FrameStrobe[11] Tile_X4Y14_RegFile/FrameStrobe[12] Tile_X4Y14_RegFile/FrameStrobe[13]
+ Tile_X4Y14_RegFile/FrameStrobe[14] Tile_X4Y14_RegFile/FrameStrobe[15] Tile_X4Y14_RegFile/FrameStrobe[16]
+ Tile_X4Y14_RegFile/FrameStrobe[17] Tile_X4Y14_RegFile/FrameStrobe[18] Tile_X4Y14_RegFile/FrameStrobe[19]
+ Tile_X4Y14_RegFile/FrameStrobe[1] Tile_X4Y14_RegFile/FrameStrobe[2] Tile_X4Y14_RegFile/FrameStrobe[3]
+ Tile_X4Y14_RegFile/FrameStrobe[4] Tile_X4Y14_RegFile/FrameStrobe[5] Tile_X4Y14_RegFile/FrameStrobe[6]
+ Tile_X4Y14_RegFile/FrameStrobe[7] Tile_X4Y14_RegFile/FrameStrobe[8] Tile_X4Y14_RegFile/FrameStrobe[9]
+ Tile_X4Y13_RegFile/FrameStrobe[0] Tile_X4Y13_RegFile/FrameStrobe[10] Tile_X4Y13_RegFile/FrameStrobe[11]
+ Tile_X4Y13_RegFile/FrameStrobe[12] Tile_X4Y13_RegFile/FrameStrobe[13] Tile_X4Y13_RegFile/FrameStrobe[14]
+ Tile_X4Y13_RegFile/FrameStrobe[15] Tile_X4Y13_RegFile/FrameStrobe[16] Tile_X4Y13_RegFile/FrameStrobe[17]
+ Tile_X4Y13_RegFile/FrameStrobe[18] Tile_X4Y13_RegFile/FrameStrobe[19] Tile_X4Y13_RegFile/FrameStrobe[1]
+ Tile_X4Y13_RegFile/FrameStrobe[2] Tile_X4Y13_RegFile/FrameStrobe[3] Tile_X4Y13_RegFile/FrameStrobe[4]
+ Tile_X4Y13_RegFile/FrameStrobe[5] Tile_X4Y13_RegFile/FrameStrobe[6] Tile_X4Y13_RegFile/FrameStrobe[7]
+ Tile_X4Y13_RegFile/FrameStrobe[8] Tile_X4Y13_RegFile/FrameStrobe[9] Tile_X4Y14_RegFile/N1BEG[0]
+ Tile_X4Y14_RegFile/N1BEG[1] Tile_X4Y14_RegFile/N1BEG[2] Tile_X4Y14_RegFile/N1BEG[3]
+ Tile_X4Y14_RegFile/N1END[0] Tile_X4Y14_RegFile/N1END[1] Tile_X4Y14_RegFile/N1END[2]
+ Tile_X4Y14_RegFile/N1END[3] Tile_X4Y14_RegFile/N2BEG[0] Tile_X4Y14_RegFile/N2BEG[1]
+ Tile_X4Y14_RegFile/N2BEG[2] Tile_X4Y14_RegFile/N2BEG[3] Tile_X4Y14_RegFile/N2BEG[4]
+ Tile_X4Y14_RegFile/N2BEG[5] Tile_X4Y14_RegFile/N2BEG[6] Tile_X4Y14_RegFile/N2BEG[7]
+ Tile_X4Y13_RegFile/N2END[0] Tile_X4Y13_RegFile/N2END[1] Tile_X4Y13_RegFile/N2END[2]
+ Tile_X4Y13_RegFile/N2END[3] Tile_X4Y13_RegFile/N2END[4] Tile_X4Y13_RegFile/N2END[5]
+ Tile_X4Y13_RegFile/N2END[6] Tile_X4Y13_RegFile/N2END[7] Tile_X4Y14_RegFile/N2END[0]
+ Tile_X4Y14_RegFile/N2END[1] Tile_X4Y14_RegFile/N2END[2] Tile_X4Y14_RegFile/N2END[3]
+ Tile_X4Y14_RegFile/N2END[4] Tile_X4Y14_RegFile/N2END[5] Tile_X4Y14_RegFile/N2END[6]
+ Tile_X4Y14_RegFile/N2END[7] Tile_X4Y14_RegFile/N2MID[0] Tile_X4Y14_RegFile/N2MID[1]
+ Tile_X4Y14_RegFile/N2MID[2] Tile_X4Y14_RegFile/N2MID[3] Tile_X4Y14_RegFile/N2MID[4]
+ Tile_X4Y14_RegFile/N2MID[5] Tile_X4Y14_RegFile/N2MID[6] Tile_X4Y14_RegFile/N2MID[7]
+ Tile_X4Y14_RegFile/N4BEG[0] Tile_X4Y14_RegFile/N4BEG[10] Tile_X4Y14_RegFile/N4BEG[11]
+ Tile_X4Y14_RegFile/N4BEG[12] Tile_X4Y14_RegFile/N4BEG[13] Tile_X4Y14_RegFile/N4BEG[14]
+ Tile_X4Y14_RegFile/N4BEG[15] Tile_X4Y14_RegFile/N4BEG[1] Tile_X4Y14_RegFile/N4BEG[2]
+ Tile_X4Y14_RegFile/N4BEG[3] Tile_X4Y14_RegFile/N4BEG[4] Tile_X4Y14_RegFile/N4BEG[5]
+ Tile_X4Y14_RegFile/N4BEG[6] Tile_X4Y14_RegFile/N4BEG[7] Tile_X4Y14_RegFile/N4BEG[8]
+ Tile_X4Y14_RegFile/N4BEG[9] Tile_X4Y14_RegFile/N4END[0] Tile_X4Y14_RegFile/N4END[10]
+ Tile_X4Y14_RegFile/N4END[11] Tile_X4Y14_RegFile/N4END[12] Tile_X4Y14_RegFile/N4END[13]
+ Tile_X4Y14_RegFile/N4END[14] Tile_X4Y14_RegFile/N4END[15] Tile_X4Y14_RegFile/N4END[1]
+ Tile_X4Y14_RegFile/N4END[2] Tile_X4Y14_RegFile/N4END[3] Tile_X4Y14_RegFile/N4END[4]
+ Tile_X4Y14_RegFile/N4END[5] Tile_X4Y14_RegFile/N4END[6] Tile_X4Y14_RegFile/N4END[7]
+ Tile_X4Y14_RegFile/N4END[8] Tile_X4Y14_RegFile/N4END[9] Tile_X4Y14_RegFile/NN4BEG[0]
+ Tile_X4Y14_RegFile/NN4BEG[10] Tile_X4Y14_RegFile/NN4BEG[11] Tile_X4Y14_RegFile/NN4BEG[12]
+ Tile_X4Y14_RegFile/NN4BEG[13] Tile_X4Y14_RegFile/NN4BEG[14] Tile_X4Y14_RegFile/NN4BEG[15]
+ Tile_X4Y14_RegFile/NN4BEG[1] Tile_X4Y14_RegFile/NN4BEG[2] Tile_X4Y14_RegFile/NN4BEG[3]
+ Tile_X4Y14_RegFile/NN4BEG[4] Tile_X4Y14_RegFile/NN4BEG[5] Tile_X4Y14_RegFile/NN4BEG[6]
+ Tile_X4Y14_RegFile/NN4BEG[7] Tile_X4Y14_RegFile/NN4BEG[8] Tile_X4Y14_RegFile/NN4BEG[9]
+ Tile_X4Y14_RegFile/NN4END[0] Tile_X4Y14_RegFile/NN4END[10] Tile_X4Y14_RegFile/NN4END[11]
+ Tile_X4Y14_RegFile/NN4END[12] Tile_X4Y14_RegFile/NN4END[13] Tile_X4Y14_RegFile/NN4END[14]
+ Tile_X4Y14_RegFile/NN4END[15] Tile_X4Y14_RegFile/NN4END[1] Tile_X4Y14_RegFile/NN4END[2]
+ Tile_X4Y14_RegFile/NN4END[3] Tile_X4Y14_RegFile/NN4END[4] Tile_X4Y14_RegFile/NN4END[5]
+ Tile_X4Y14_RegFile/NN4END[6] Tile_X4Y14_RegFile/NN4END[7] Tile_X4Y14_RegFile/NN4END[8]
+ Tile_X4Y14_RegFile/NN4END[9] Tile_X4Y14_RegFile/S1BEG[0] Tile_X4Y14_RegFile/S1BEG[1]
+ Tile_X4Y14_RegFile/S1BEG[2] Tile_X4Y14_RegFile/S1BEG[3] Tile_X4Y14_RegFile/S1END[0]
+ Tile_X4Y14_RegFile/S1END[1] Tile_X4Y14_RegFile/S1END[2] Tile_X4Y14_RegFile/S1END[3]
+ Tile_X4Y14_RegFile/S2BEG[0] Tile_X4Y14_RegFile/S2BEG[1] Tile_X4Y14_RegFile/S2BEG[2]
+ Tile_X4Y14_RegFile/S2BEG[3] Tile_X4Y14_RegFile/S2BEG[4] Tile_X4Y14_RegFile/S2BEG[5]
+ Tile_X4Y14_RegFile/S2BEG[6] Tile_X4Y14_RegFile/S2BEG[7] Tile_X4Y14_RegFile/S2BEGb[0]
+ Tile_X4Y14_RegFile/S2BEGb[1] Tile_X4Y14_RegFile/S2BEGb[2] Tile_X4Y14_RegFile/S2BEGb[3]
+ Tile_X4Y14_RegFile/S2BEGb[4] Tile_X4Y14_RegFile/S2BEGb[5] Tile_X4Y14_RegFile/S2BEGb[6]
+ Tile_X4Y14_RegFile/S2BEGb[7] Tile_X4Y14_RegFile/S2END[0] Tile_X4Y14_RegFile/S2END[1]
+ Tile_X4Y14_RegFile/S2END[2] Tile_X4Y14_RegFile/S2END[3] Tile_X4Y14_RegFile/S2END[4]
+ Tile_X4Y14_RegFile/S2END[5] Tile_X4Y14_RegFile/S2END[6] Tile_X4Y14_RegFile/S2END[7]
+ Tile_X4Y14_RegFile/S2MID[0] Tile_X4Y14_RegFile/S2MID[1] Tile_X4Y14_RegFile/S2MID[2]
+ Tile_X4Y14_RegFile/S2MID[3] Tile_X4Y14_RegFile/S2MID[4] Tile_X4Y14_RegFile/S2MID[5]
+ Tile_X4Y14_RegFile/S2MID[6] Tile_X4Y14_RegFile/S2MID[7] Tile_X4Y14_RegFile/S4BEG[0]
+ Tile_X4Y14_RegFile/S4BEG[10] Tile_X4Y14_RegFile/S4BEG[11] Tile_X4Y14_RegFile/S4BEG[12]
+ Tile_X4Y14_RegFile/S4BEG[13] Tile_X4Y14_RegFile/S4BEG[14] Tile_X4Y14_RegFile/S4BEG[15]
+ Tile_X4Y14_RegFile/S4BEG[1] Tile_X4Y14_RegFile/S4BEG[2] Tile_X4Y14_RegFile/S4BEG[3]
+ Tile_X4Y14_RegFile/S4BEG[4] Tile_X4Y14_RegFile/S4BEG[5] Tile_X4Y14_RegFile/S4BEG[6]
+ Tile_X4Y14_RegFile/S4BEG[7] Tile_X4Y14_RegFile/S4BEG[8] Tile_X4Y14_RegFile/S4BEG[9]
+ Tile_X4Y14_RegFile/S4END[0] Tile_X4Y14_RegFile/S4END[10] Tile_X4Y14_RegFile/S4END[11]
+ Tile_X4Y14_RegFile/S4END[12] Tile_X4Y14_RegFile/S4END[13] Tile_X4Y14_RegFile/S4END[14]
+ Tile_X4Y14_RegFile/S4END[15] Tile_X4Y14_RegFile/S4END[1] Tile_X4Y14_RegFile/S4END[2]
+ Tile_X4Y14_RegFile/S4END[3] Tile_X4Y14_RegFile/S4END[4] Tile_X4Y14_RegFile/S4END[5]
+ Tile_X4Y14_RegFile/S4END[6] Tile_X4Y14_RegFile/S4END[7] Tile_X4Y14_RegFile/S4END[8]
+ Tile_X4Y14_RegFile/S4END[9] Tile_X4Y14_RegFile/SS4BEG[0] Tile_X4Y14_RegFile/SS4BEG[10]
+ Tile_X4Y14_RegFile/SS4BEG[11] Tile_X4Y14_RegFile/SS4BEG[12] Tile_X4Y14_RegFile/SS4BEG[13]
+ Tile_X4Y14_RegFile/SS4BEG[14] Tile_X4Y14_RegFile/SS4BEG[15] Tile_X4Y14_RegFile/SS4BEG[1]
+ Tile_X4Y14_RegFile/SS4BEG[2] Tile_X4Y14_RegFile/SS4BEG[3] Tile_X4Y14_RegFile/SS4BEG[4]
+ Tile_X4Y14_RegFile/SS4BEG[5] Tile_X4Y14_RegFile/SS4BEG[6] Tile_X4Y14_RegFile/SS4BEG[7]
+ Tile_X4Y14_RegFile/SS4BEG[8] Tile_X4Y14_RegFile/SS4BEG[9] Tile_X4Y14_RegFile/SS4END[0]
+ Tile_X4Y14_RegFile/SS4END[10] Tile_X4Y14_RegFile/SS4END[11] Tile_X4Y14_RegFile/SS4END[12]
+ Tile_X4Y14_RegFile/SS4END[13] Tile_X4Y14_RegFile/SS4END[14] Tile_X4Y14_RegFile/SS4END[15]
+ Tile_X4Y14_RegFile/SS4END[1] Tile_X4Y14_RegFile/SS4END[2] Tile_X4Y14_RegFile/SS4END[3]
+ Tile_X4Y14_RegFile/SS4END[4] Tile_X4Y14_RegFile/SS4END[5] Tile_X4Y14_RegFile/SS4END[6]
+ Tile_X4Y14_RegFile/SS4END[7] Tile_X4Y14_RegFile/SS4END[8] Tile_X4Y14_RegFile/SS4END[9]
+ Tile_X4Y14_RegFile/UserCLK Tile_X4Y13_RegFile/UserCLK VGND VPWR Tile_X3Y14_LUT4AB/W1END[0]
+ Tile_X3Y14_LUT4AB/W1END[1] Tile_X3Y14_LUT4AB/W1END[2] Tile_X3Y14_LUT4AB/W1END[3]
+ Tile_X5Y14_LUT4AB/W1BEG[0] Tile_X5Y14_LUT4AB/W1BEG[1] Tile_X5Y14_LUT4AB/W1BEG[2]
+ Tile_X5Y14_LUT4AB/W1BEG[3] Tile_X3Y14_LUT4AB/W2MID[0] Tile_X3Y14_LUT4AB/W2MID[1]
+ Tile_X3Y14_LUT4AB/W2MID[2] Tile_X3Y14_LUT4AB/W2MID[3] Tile_X3Y14_LUT4AB/W2MID[4]
+ Tile_X3Y14_LUT4AB/W2MID[5] Tile_X3Y14_LUT4AB/W2MID[6] Tile_X3Y14_LUT4AB/W2MID[7]
+ Tile_X3Y14_LUT4AB/W2END[0] Tile_X3Y14_LUT4AB/W2END[1] Tile_X3Y14_LUT4AB/W2END[2]
+ Tile_X3Y14_LUT4AB/W2END[3] Tile_X3Y14_LUT4AB/W2END[4] Tile_X3Y14_LUT4AB/W2END[5]
+ Tile_X3Y14_LUT4AB/W2END[6] Tile_X3Y14_LUT4AB/W2END[7] Tile_X5Y14_LUT4AB/W2BEGb[0]
+ Tile_X5Y14_LUT4AB/W2BEGb[1] Tile_X5Y14_LUT4AB/W2BEGb[2] Tile_X5Y14_LUT4AB/W2BEGb[3]
+ Tile_X5Y14_LUT4AB/W2BEGb[4] Tile_X5Y14_LUT4AB/W2BEGb[5] Tile_X5Y14_LUT4AB/W2BEGb[6]
+ Tile_X5Y14_LUT4AB/W2BEGb[7] Tile_X5Y14_LUT4AB/W2BEG[0] Tile_X5Y14_LUT4AB/W2BEG[1]
+ Tile_X5Y14_LUT4AB/W2BEG[2] Tile_X5Y14_LUT4AB/W2BEG[3] Tile_X5Y14_LUT4AB/W2BEG[4]
+ Tile_X5Y14_LUT4AB/W2BEG[5] Tile_X5Y14_LUT4AB/W2BEG[6] Tile_X5Y14_LUT4AB/W2BEG[7]
+ Tile_X3Y14_LUT4AB/W6END[0] Tile_X3Y14_LUT4AB/W6END[10] Tile_X3Y14_LUT4AB/W6END[11]
+ Tile_X3Y14_LUT4AB/W6END[1] Tile_X3Y14_LUT4AB/W6END[2] Tile_X3Y14_LUT4AB/W6END[3]
+ Tile_X3Y14_LUT4AB/W6END[4] Tile_X3Y14_LUT4AB/W6END[5] Tile_X3Y14_LUT4AB/W6END[6]
+ Tile_X3Y14_LUT4AB/W6END[7] Tile_X3Y14_LUT4AB/W6END[8] Tile_X3Y14_LUT4AB/W6END[9]
+ Tile_X5Y14_LUT4AB/W6BEG[0] Tile_X5Y14_LUT4AB/W6BEG[10] Tile_X5Y14_LUT4AB/W6BEG[11]
+ Tile_X5Y14_LUT4AB/W6BEG[1] Tile_X5Y14_LUT4AB/W6BEG[2] Tile_X5Y14_LUT4AB/W6BEG[3]
+ Tile_X5Y14_LUT4AB/W6BEG[4] Tile_X5Y14_LUT4AB/W6BEG[5] Tile_X5Y14_LUT4AB/W6BEG[6]
+ Tile_X5Y14_LUT4AB/W6BEG[7] Tile_X5Y14_LUT4AB/W6BEG[8] Tile_X5Y14_LUT4AB/W6BEG[9]
+ Tile_X3Y14_LUT4AB/WW4END[0] Tile_X3Y14_LUT4AB/WW4END[10] Tile_X3Y14_LUT4AB/WW4END[11]
+ Tile_X3Y14_LUT4AB/WW4END[12] Tile_X3Y14_LUT4AB/WW4END[13] Tile_X3Y14_LUT4AB/WW4END[14]
+ Tile_X3Y14_LUT4AB/WW4END[15] Tile_X3Y14_LUT4AB/WW4END[1] Tile_X3Y14_LUT4AB/WW4END[2]
+ Tile_X3Y14_LUT4AB/WW4END[3] Tile_X3Y14_LUT4AB/WW4END[4] Tile_X3Y14_LUT4AB/WW4END[5]
+ Tile_X3Y14_LUT4AB/WW4END[6] Tile_X3Y14_LUT4AB/WW4END[7] Tile_X3Y14_LUT4AB/WW4END[8]
+ Tile_X3Y14_LUT4AB/WW4END[9] Tile_X5Y14_LUT4AB/WW4BEG[0] Tile_X5Y14_LUT4AB/WW4BEG[10]
+ Tile_X5Y14_LUT4AB/WW4BEG[11] Tile_X5Y14_LUT4AB/WW4BEG[12] Tile_X5Y14_LUT4AB/WW4BEG[13]
+ Tile_X5Y14_LUT4AB/WW4BEG[14] Tile_X5Y14_LUT4AB/WW4BEG[15] Tile_X5Y14_LUT4AB/WW4BEG[1]
+ Tile_X5Y14_LUT4AB/WW4BEG[2] Tile_X5Y14_LUT4AB/WW4BEG[3] Tile_X5Y14_LUT4AB/WW4BEG[4]
+ Tile_X5Y14_LUT4AB/WW4BEG[5] Tile_X5Y14_LUT4AB/WW4BEG[6] Tile_X5Y14_LUT4AB/WW4BEG[7]
+ Tile_X5Y14_LUT4AB/WW4BEG[8] Tile_X5Y14_LUT4AB/WW4BEG[9] RegFile
XTile_X10Y7_IHP_SRAM Tile_X10Y8_ADDR_SRAM0 Tile_X10Y8_ADDR_SRAM1 Tile_X10Y8_ADDR_SRAM2
+ Tile_X10Y8_ADDR_SRAM3 Tile_X10Y8_ADDR_SRAM4 Tile_X10Y8_ADDR_SRAM5 Tile_X10Y8_ADDR_SRAM6
+ Tile_X10Y8_ADDR_SRAM7 Tile_X10Y8_ADDR_SRAM8 Tile_X10Y8_ADDR_SRAM9 Tile_X10Y8_BM_SRAM0
+ Tile_X10Y8_BM_SRAM1 Tile_X10Y8_BM_SRAM10 Tile_X10Y8_BM_SRAM11 Tile_X10Y8_BM_SRAM12
+ Tile_X10Y8_BM_SRAM13 Tile_X10Y8_BM_SRAM14 Tile_X10Y8_BM_SRAM15 Tile_X10Y8_BM_SRAM16
+ Tile_X10Y8_BM_SRAM17 Tile_X10Y8_BM_SRAM18 Tile_X10Y8_BM_SRAM19 Tile_X10Y8_BM_SRAM2
+ Tile_X10Y8_BM_SRAM20 Tile_X10Y8_BM_SRAM21 Tile_X10Y8_BM_SRAM22 Tile_X10Y8_BM_SRAM23
+ Tile_X10Y8_BM_SRAM24 Tile_X10Y8_BM_SRAM25 Tile_X10Y8_BM_SRAM26 Tile_X10Y8_BM_SRAM27
+ Tile_X10Y8_BM_SRAM28 Tile_X10Y8_BM_SRAM29 Tile_X10Y8_BM_SRAM3 Tile_X10Y8_BM_SRAM30
+ Tile_X10Y8_BM_SRAM31 Tile_X10Y8_BM_SRAM4 Tile_X10Y8_BM_SRAM5 Tile_X10Y8_BM_SRAM6
+ Tile_X10Y8_BM_SRAM7 Tile_X10Y8_BM_SRAM8 Tile_X10Y8_BM_SRAM9 Tile_X10Y8_CLK_SRAM
+ Tile_X10Y8_CONFIGURED_top Tile_X10Y8_DIN_SRAM0 Tile_X10Y8_DIN_SRAM1 Tile_X10Y8_DIN_SRAM10
+ Tile_X10Y8_DIN_SRAM11 Tile_X10Y8_DIN_SRAM12 Tile_X10Y8_DIN_SRAM13 Tile_X10Y8_DIN_SRAM14
+ Tile_X10Y8_DIN_SRAM15 Tile_X10Y8_DIN_SRAM16 Tile_X10Y8_DIN_SRAM17 Tile_X10Y8_DIN_SRAM18
+ Tile_X10Y8_DIN_SRAM19 Tile_X10Y8_DIN_SRAM2 Tile_X10Y8_DIN_SRAM20 Tile_X10Y8_DIN_SRAM21
+ Tile_X10Y8_DIN_SRAM22 Tile_X10Y8_DIN_SRAM23 Tile_X10Y8_DIN_SRAM24 Tile_X10Y8_DIN_SRAM25
+ Tile_X10Y8_DIN_SRAM26 Tile_X10Y8_DIN_SRAM27 Tile_X10Y8_DIN_SRAM28 Tile_X10Y8_DIN_SRAM29
+ Tile_X10Y8_DIN_SRAM3 Tile_X10Y8_DIN_SRAM30 Tile_X10Y8_DIN_SRAM31 Tile_X10Y8_DIN_SRAM4
+ Tile_X10Y8_DIN_SRAM5 Tile_X10Y8_DIN_SRAM6 Tile_X10Y8_DIN_SRAM7 Tile_X10Y8_DIN_SRAM8
+ Tile_X10Y8_DIN_SRAM9 Tile_X10Y8_DOUT_SRAM0 Tile_X10Y8_DOUT_SRAM1 Tile_X10Y8_DOUT_SRAM10
+ Tile_X10Y8_DOUT_SRAM11 Tile_X10Y8_DOUT_SRAM12 Tile_X10Y8_DOUT_SRAM13 Tile_X10Y8_DOUT_SRAM14
+ Tile_X10Y8_DOUT_SRAM15 Tile_X10Y8_DOUT_SRAM16 Tile_X10Y8_DOUT_SRAM17 Tile_X10Y8_DOUT_SRAM18
+ Tile_X10Y8_DOUT_SRAM19 Tile_X10Y8_DOUT_SRAM2 Tile_X10Y8_DOUT_SRAM20 Tile_X10Y8_DOUT_SRAM21
+ Tile_X10Y8_DOUT_SRAM22 Tile_X10Y8_DOUT_SRAM23 Tile_X10Y8_DOUT_SRAM24 Tile_X10Y8_DOUT_SRAM25
+ Tile_X10Y8_DOUT_SRAM26 Tile_X10Y8_DOUT_SRAM27 Tile_X10Y8_DOUT_SRAM28 Tile_X10Y8_DOUT_SRAM29
+ Tile_X10Y8_DOUT_SRAM3 Tile_X10Y8_DOUT_SRAM30 Tile_X10Y8_DOUT_SRAM31 Tile_X10Y8_DOUT_SRAM4
+ Tile_X10Y8_DOUT_SRAM5 Tile_X10Y8_DOUT_SRAM6 Tile_X10Y8_DOUT_SRAM7 Tile_X10Y8_DOUT_SRAM8
+ Tile_X10Y8_DOUT_SRAM9 Tile_X10Y8_MEN_SRAM Tile_X10Y8_REN_SRAM Tile_X10Y8_TIE_HIGH_SRAM
+ Tile_X10Y8_TIE_LOW_SRAM Tile_X9Y7_LUT4AB/E1BEG[0] Tile_X9Y7_LUT4AB/E1BEG[1] Tile_X9Y7_LUT4AB/E1BEG[2]
+ Tile_X9Y7_LUT4AB/E1BEG[3] Tile_X9Y7_LUT4AB/E2BEGb[0] Tile_X9Y7_LUT4AB/E2BEGb[1]
+ Tile_X9Y7_LUT4AB/E2BEGb[2] Tile_X9Y7_LUT4AB/E2BEGb[3] Tile_X9Y7_LUT4AB/E2BEGb[4]
+ Tile_X9Y7_LUT4AB/E2BEGb[5] Tile_X9Y7_LUT4AB/E2BEGb[6] Tile_X9Y7_LUT4AB/E2BEGb[7]
+ Tile_X9Y7_LUT4AB/E2BEG[0] Tile_X9Y7_LUT4AB/E2BEG[1] Tile_X9Y7_LUT4AB/E2BEG[2] Tile_X9Y7_LUT4AB/E2BEG[3]
+ Tile_X9Y7_LUT4AB/E2BEG[4] Tile_X9Y7_LUT4AB/E2BEG[5] Tile_X9Y7_LUT4AB/E2BEG[6] Tile_X9Y7_LUT4AB/E2BEG[7]
+ Tile_X9Y7_LUT4AB/E6BEG[0] Tile_X9Y7_LUT4AB/E6BEG[10] Tile_X9Y7_LUT4AB/E6BEG[11]
+ Tile_X9Y7_LUT4AB/E6BEG[1] Tile_X9Y7_LUT4AB/E6BEG[2] Tile_X9Y7_LUT4AB/E6BEG[3] Tile_X9Y7_LUT4AB/E6BEG[4]
+ Tile_X9Y7_LUT4AB/E6BEG[5] Tile_X9Y7_LUT4AB/E6BEG[6] Tile_X9Y7_LUT4AB/E6BEG[7] Tile_X9Y7_LUT4AB/E6BEG[8]
+ Tile_X9Y7_LUT4AB/E6BEG[9] Tile_X9Y7_LUT4AB/EE4BEG[0] Tile_X9Y7_LUT4AB/EE4BEG[10]
+ Tile_X9Y7_LUT4AB/EE4BEG[11] Tile_X9Y7_LUT4AB/EE4BEG[12] Tile_X9Y7_LUT4AB/EE4BEG[13]
+ Tile_X9Y7_LUT4AB/EE4BEG[14] Tile_X9Y7_LUT4AB/EE4BEG[15] Tile_X9Y7_LUT4AB/EE4BEG[1]
+ Tile_X9Y7_LUT4AB/EE4BEG[2] Tile_X9Y7_LUT4AB/EE4BEG[3] Tile_X9Y7_LUT4AB/EE4BEG[4]
+ Tile_X9Y7_LUT4AB/EE4BEG[5] Tile_X9Y7_LUT4AB/EE4BEG[6] Tile_X9Y7_LUT4AB/EE4BEG[7]
+ Tile_X9Y7_LUT4AB/EE4BEG[8] Tile_X9Y7_LUT4AB/EE4BEG[9] Tile_X9Y7_LUT4AB/FrameData_O[0]
+ Tile_X9Y7_LUT4AB/FrameData_O[10] Tile_X9Y7_LUT4AB/FrameData_O[11] Tile_X9Y7_LUT4AB/FrameData_O[12]
+ Tile_X9Y7_LUT4AB/FrameData_O[13] Tile_X9Y7_LUT4AB/FrameData_O[14] Tile_X9Y7_LUT4AB/FrameData_O[15]
+ Tile_X9Y7_LUT4AB/FrameData_O[16] Tile_X9Y7_LUT4AB/FrameData_O[17] Tile_X9Y7_LUT4AB/FrameData_O[18]
+ Tile_X9Y7_LUT4AB/FrameData_O[19] Tile_X9Y7_LUT4AB/FrameData_O[1] Tile_X9Y7_LUT4AB/FrameData_O[20]
+ Tile_X9Y7_LUT4AB/FrameData_O[21] Tile_X9Y7_LUT4AB/FrameData_O[22] Tile_X9Y7_LUT4AB/FrameData_O[23]
+ Tile_X9Y7_LUT4AB/FrameData_O[24] Tile_X9Y7_LUT4AB/FrameData_O[25] Tile_X9Y7_LUT4AB/FrameData_O[26]
+ Tile_X9Y7_LUT4AB/FrameData_O[27] Tile_X9Y7_LUT4AB/FrameData_O[28] Tile_X9Y7_LUT4AB/FrameData_O[29]
+ Tile_X9Y7_LUT4AB/FrameData_O[2] Tile_X9Y7_LUT4AB/FrameData_O[30] Tile_X9Y7_LUT4AB/FrameData_O[31]
+ Tile_X9Y7_LUT4AB/FrameData_O[3] Tile_X9Y7_LUT4AB/FrameData_O[4] Tile_X9Y7_LUT4AB/FrameData_O[5]
+ Tile_X9Y7_LUT4AB/FrameData_O[6] Tile_X9Y7_LUT4AB/FrameData_O[7] Tile_X9Y7_LUT4AB/FrameData_O[8]
+ Tile_X9Y7_LUT4AB/FrameData_O[9] Tile_X10Y7_IHP_SRAM/Tile_X0Y0_FrameData_O[0] Tile_X10Y7_IHP_SRAM/Tile_X0Y0_FrameData_O[10]
+ Tile_X10Y7_IHP_SRAM/Tile_X0Y0_FrameData_O[11] Tile_X10Y7_IHP_SRAM/Tile_X0Y0_FrameData_O[12]
+ Tile_X10Y7_IHP_SRAM/Tile_X0Y0_FrameData_O[13] Tile_X10Y7_IHP_SRAM/Tile_X0Y0_FrameData_O[14]
+ Tile_X10Y7_IHP_SRAM/Tile_X0Y0_FrameData_O[15] Tile_X10Y7_IHP_SRAM/Tile_X0Y0_FrameData_O[16]
+ Tile_X10Y7_IHP_SRAM/Tile_X0Y0_FrameData_O[17] Tile_X10Y7_IHP_SRAM/Tile_X0Y0_FrameData_O[18]
+ Tile_X10Y7_IHP_SRAM/Tile_X0Y0_FrameData_O[19] Tile_X10Y7_IHP_SRAM/Tile_X0Y0_FrameData_O[1]
+ Tile_X10Y7_IHP_SRAM/Tile_X0Y0_FrameData_O[20] Tile_X10Y7_IHP_SRAM/Tile_X0Y0_FrameData_O[21]
+ Tile_X10Y7_IHP_SRAM/Tile_X0Y0_FrameData_O[22] Tile_X10Y7_IHP_SRAM/Tile_X0Y0_FrameData_O[23]
+ Tile_X10Y7_IHP_SRAM/Tile_X0Y0_FrameData_O[24] Tile_X10Y7_IHP_SRAM/Tile_X0Y0_FrameData_O[25]
+ Tile_X10Y7_IHP_SRAM/Tile_X0Y0_FrameData_O[26] Tile_X10Y7_IHP_SRAM/Tile_X0Y0_FrameData_O[27]
+ Tile_X10Y7_IHP_SRAM/Tile_X0Y0_FrameData_O[28] Tile_X10Y7_IHP_SRAM/Tile_X0Y0_FrameData_O[29]
+ Tile_X10Y7_IHP_SRAM/Tile_X0Y0_FrameData_O[2] Tile_X10Y7_IHP_SRAM/Tile_X0Y0_FrameData_O[30]
+ Tile_X10Y7_IHP_SRAM/Tile_X0Y0_FrameData_O[31] Tile_X10Y7_IHP_SRAM/Tile_X0Y0_FrameData_O[3]
+ Tile_X10Y7_IHP_SRAM/Tile_X0Y0_FrameData_O[4] Tile_X10Y7_IHP_SRAM/Tile_X0Y0_FrameData_O[5]
+ Tile_X10Y7_IHP_SRAM/Tile_X0Y0_FrameData_O[6] Tile_X10Y7_IHP_SRAM/Tile_X0Y0_FrameData_O[7]
+ Tile_X10Y7_IHP_SRAM/Tile_X0Y0_FrameData_O[8] Tile_X10Y7_IHP_SRAM/Tile_X0Y0_FrameData_O[9]
+ Tile_X10Y5_IHP_SRAM/Tile_X0Y1_FrameStrobe[0] Tile_X10Y5_IHP_SRAM/Tile_X0Y1_FrameStrobe[10]
+ Tile_X10Y5_IHP_SRAM/Tile_X0Y1_FrameStrobe[11] Tile_X10Y5_IHP_SRAM/Tile_X0Y1_FrameStrobe[12]
+ Tile_X10Y5_IHP_SRAM/Tile_X0Y1_FrameStrobe[13] Tile_X10Y5_IHP_SRAM/Tile_X0Y1_FrameStrobe[14]
+ Tile_X10Y5_IHP_SRAM/Tile_X0Y1_FrameStrobe[15] Tile_X10Y5_IHP_SRAM/Tile_X0Y1_FrameStrobe[16]
+ Tile_X10Y5_IHP_SRAM/Tile_X0Y1_FrameStrobe[17] Tile_X10Y5_IHP_SRAM/Tile_X0Y1_FrameStrobe[18]
+ Tile_X10Y5_IHP_SRAM/Tile_X0Y1_FrameStrobe[19] Tile_X10Y5_IHP_SRAM/Tile_X0Y1_FrameStrobe[1]
+ Tile_X10Y5_IHP_SRAM/Tile_X0Y1_FrameStrobe[2] Tile_X10Y5_IHP_SRAM/Tile_X0Y1_FrameStrobe[3]
+ Tile_X10Y5_IHP_SRAM/Tile_X0Y1_FrameStrobe[4] Tile_X10Y5_IHP_SRAM/Tile_X0Y1_FrameStrobe[5]
+ Tile_X10Y5_IHP_SRAM/Tile_X0Y1_FrameStrobe[6] Tile_X10Y5_IHP_SRAM/Tile_X0Y1_FrameStrobe[7]
+ Tile_X10Y5_IHP_SRAM/Tile_X0Y1_FrameStrobe[8] Tile_X10Y5_IHP_SRAM/Tile_X0Y1_FrameStrobe[9]
+ Tile_X10Y7_IHP_SRAM/Tile_X0Y0_N1BEG[0] Tile_X10Y7_IHP_SRAM/Tile_X0Y0_N1BEG[1] Tile_X10Y7_IHP_SRAM/Tile_X0Y0_N1BEG[2]
+ Tile_X10Y7_IHP_SRAM/Tile_X0Y0_N1BEG[3] Tile_X10Y7_IHP_SRAM/Tile_X0Y0_N2BEG[0] Tile_X10Y7_IHP_SRAM/Tile_X0Y0_N2BEG[1]
+ Tile_X10Y7_IHP_SRAM/Tile_X0Y0_N2BEG[2] Tile_X10Y7_IHP_SRAM/Tile_X0Y0_N2BEG[3] Tile_X10Y7_IHP_SRAM/Tile_X0Y0_N2BEG[4]
+ Tile_X10Y7_IHP_SRAM/Tile_X0Y0_N2BEG[5] Tile_X10Y7_IHP_SRAM/Tile_X0Y0_N2BEG[6] Tile_X10Y7_IHP_SRAM/Tile_X0Y0_N2BEG[7]
+ Tile_X10Y5_IHP_SRAM/Tile_X0Y1_N2END[0] Tile_X10Y5_IHP_SRAM/Tile_X0Y1_N2END[1] Tile_X10Y5_IHP_SRAM/Tile_X0Y1_N2END[2]
+ Tile_X10Y5_IHP_SRAM/Tile_X0Y1_N2END[3] Tile_X10Y5_IHP_SRAM/Tile_X0Y1_N2END[4] Tile_X10Y5_IHP_SRAM/Tile_X0Y1_N2END[5]
+ Tile_X10Y5_IHP_SRAM/Tile_X0Y1_N2END[6] Tile_X10Y5_IHP_SRAM/Tile_X0Y1_N2END[7] Tile_X10Y7_IHP_SRAM/Tile_X0Y0_N4BEG[0]
+ Tile_X10Y7_IHP_SRAM/Tile_X0Y0_N4BEG[10] Tile_X10Y7_IHP_SRAM/Tile_X0Y0_N4BEG[11]
+ Tile_X10Y7_IHP_SRAM/Tile_X0Y0_N4BEG[12] Tile_X10Y7_IHP_SRAM/Tile_X0Y0_N4BEG[13]
+ Tile_X10Y7_IHP_SRAM/Tile_X0Y0_N4BEG[14] Tile_X10Y7_IHP_SRAM/Tile_X0Y0_N4BEG[15]
+ Tile_X10Y7_IHP_SRAM/Tile_X0Y0_N4BEG[1] Tile_X10Y7_IHP_SRAM/Tile_X0Y0_N4BEG[2] Tile_X10Y7_IHP_SRAM/Tile_X0Y0_N4BEG[3]
+ Tile_X10Y7_IHP_SRAM/Tile_X0Y0_N4BEG[4] Tile_X10Y7_IHP_SRAM/Tile_X0Y0_N4BEG[5] Tile_X10Y7_IHP_SRAM/Tile_X0Y0_N4BEG[6]
+ Tile_X10Y7_IHP_SRAM/Tile_X0Y0_N4BEG[7] Tile_X10Y7_IHP_SRAM/Tile_X0Y0_N4BEG[8] Tile_X10Y7_IHP_SRAM/Tile_X0Y0_N4BEG[9]
+ Tile_X10Y7_IHP_SRAM/Tile_X0Y0_S1END[0] Tile_X10Y7_IHP_SRAM/Tile_X0Y0_S1END[1] Tile_X10Y7_IHP_SRAM/Tile_X0Y0_S1END[2]
+ Tile_X10Y7_IHP_SRAM/Tile_X0Y0_S1END[3] Tile_X10Y7_IHP_SRAM/Tile_X0Y0_S2END[0] Tile_X10Y7_IHP_SRAM/Tile_X0Y0_S2END[1]
+ Tile_X10Y7_IHP_SRAM/Tile_X0Y0_S2END[2] Tile_X10Y7_IHP_SRAM/Tile_X0Y0_S2END[3] Tile_X10Y7_IHP_SRAM/Tile_X0Y0_S2END[4]
+ Tile_X10Y7_IHP_SRAM/Tile_X0Y0_S2END[5] Tile_X10Y7_IHP_SRAM/Tile_X0Y0_S2END[6] Tile_X10Y7_IHP_SRAM/Tile_X0Y0_S2END[7]
+ Tile_X10Y7_IHP_SRAM/Tile_X0Y0_S2MID[0] Tile_X10Y7_IHP_SRAM/Tile_X0Y0_S2MID[1] Tile_X10Y7_IHP_SRAM/Tile_X0Y0_S2MID[2]
+ Tile_X10Y7_IHP_SRAM/Tile_X0Y0_S2MID[3] Tile_X10Y7_IHP_SRAM/Tile_X0Y0_S2MID[4] Tile_X10Y7_IHP_SRAM/Tile_X0Y0_S2MID[5]
+ Tile_X10Y7_IHP_SRAM/Tile_X0Y0_S2MID[6] Tile_X10Y7_IHP_SRAM/Tile_X0Y0_S2MID[7] Tile_X10Y7_IHP_SRAM/Tile_X0Y0_S4END[0]
+ Tile_X10Y7_IHP_SRAM/Tile_X0Y0_S4END[10] Tile_X10Y7_IHP_SRAM/Tile_X0Y0_S4END[11]
+ Tile_X10Y7_IHP_SRAM/Tile_X0Y0_S4END[12] Tile_X10Y7_IHP_SRAM/Tile_X0Y0_S4END[13]
+ Tile_X10Y7_IHP_SRAM/Tile_X0Y0_S4END[14] Tile_X10Y7_IHP_SRAM/Tile_X0Y0_S4END[15]
+ Tile_X10Y7_IHP_SRAM/Tile_X0Y0_S4END[1] Tile_X10Y7_IHP_SRAM/Tile_X0Y0_S4END[2] Tile_X10Y7_IHP_SRAM/Tile_X0Y0_S4END[3]
+ Tile_X10Y7_IHP_SRAM/Tile_X0Y0_S4END[4] Tile_X10Y7_IHP_SRAM/Tile_X0Y0_S4END[5] Tile_X10Y7_IHP_SRAM/Tile_X0Y0_S4END[6]
+ Tile_X10Y7_IHP_SRAM/Tile_X0Y0_S4END[7] Tile_X10Y7_IHP_SRAM/Tile_X0Y0_S4END[8] Tile_X10Y7_IHP_SRAM/Tile_X0Y0_S4END[9]
+ Tile_X10Y5_IHP_SRAM/Tile_X0Y1_UserCLK Tile_X9Y7_LUT4AB/W1END[0] Tile_X9Y7_LUT4AB/W1END[1]
+ Tile_X9Y7_LUT4AB/W1END[2] Tile_X9Y7_LUT4AB/W1END[3] Tile_X9Y7_LUT4AB/W2MID[0] Tile_X9Y7_LUT4AB/W2MID[1]
+ Tile_X9Y7_LUT4AB/W2MID[2] Tile_X9Y7_LUT4AB/W2MID[3] Tile_X9Y7_LUT4AB/W2MID[4] Tile_X9Y7_LUT4AB/W2MID[5]
+ Tile_X9Y7_LUT4AB/W2MID[6] Tile_X9Y7_LUT4AB/W2MID[7] Tile_X9Y7_LUT4AB/W2END[0] Tile_X9Y7_LUT4AB/W2END[1]
+ Tile_X9Y7_LUT4AB/W2END[2] Tile_X9Y7_LUT4AB/W2END[3] Tile_X9Y7_LUT4AB/W2END[4] Tile_X9Y7_LUT4AB/W2END[5]
+ Tile_X9Y7_LUT4AB/W2END[6] Tile_X9Y7_LUT4AB/W2END[7] Tile_X9Y7_LUT4AB/W6END[0] Tile_X9Y7_LUT4AB/W6END[10]
+ Tile_X9Y7_LUT4AB/W6END[11] Tile_X9Y7_LUT4AB/W6END[1] Tile_X9Y7_LUT4AB/W6END[2] Tile_X9Y7_LUT4AB/W6END[3]
+ Tile_X9Y7_LUT4AB/W6END[4] Tile_X9Y7_LUT4AB/W6END[5] Tile_X9Y7_LUT4AB/W6END[6] Tile_X9Y7_LUT4AB/W6END[7]
+ Tile_X9Y7_LUT4AB/W6END[8] Tile_X9Y7_LUT4AB/W6END[9] Tile_X9Y7_LUT4AB/WW4END[0] Tile_X9Y7_LUT4AB/WW4END[10]
+ Tile_X9Y7_LUT4AB/WW4END[11] Tile_X9Y7_LUT4AB/WW4END[12] Tile_X9Y7_LUT4AB/WW4END[13]
+ Tile_X9Y7_LUT4AB/WW4END[14] Tile_X9Y7_LUT4AB/WW4END[15] Tile_X9Y7_LUT4AB/WW4END[1]
+ Tile_X9Y7_LUT4AB/WW4END[2] Tile_X9Y7_LUT4AB/WW4END[3] Tile_X9Y7_LUT4AB/WW4END[4]
+ Tile_X9Y7_LUT4AB/WW4END[5] Tile_X9Y7_LUT4AB/WW4END[6] Tile_X9Y7_LUT4AB/WW4END[7]
+ Tile_X9Y7_LUT4AB/WW4END[8] Tile_X9Y7_LUT4AB/WW4END[9] Tile_X9Y8_LUT4AB/E1BEG[0]
+ Tile_X9Y8_LUT4AB/E1BEG[1] Tile_X9Y8_LUT4AB/E1BEG[2] Tile_X9Y8_LUT4AB/E1BEG[3] Tile_X9Y8_LUT4AB/E2BEGb[0]
+ Tile_X9Y8_LUT4AB/E2BEGb[1] Tile_X9Y8_LUT4AB/E2BEGb[2] Tile_X9Y8_LUT4AB/E2BEGb[3]
+ Tile_X9Y8_LUT4AB/E2BEGb[4] Tile_X9Y8_LUT4AB/E2BEGb[5] Tile_X9Y8_LUT4AB/E2BEGb[6]
+ Tile_X9Y8_LUT4AB/E2BEGb[7] Tile_X9Y8_LUT4AB/E2BEG[0] Tile_X9Y8_LUT4AB/E2BEG[1] Tile_X9Y8_LUT4AB/E2BEG[2]
+ Tile_X9Y8_LUT4AB/E2BEG[3] Tile_X9Y8_LUT4AB/E2BEG[4] Tile_X9Y8_LUT4AB/E2BEG[5] Tile_X9Y8_LUT4AB/E2BEG[6]
+ Tile_X9Y8_LUT4AB/E2BEG[7] Tile_X9Y8_LUT4AB/E6BEG[0] Tile_X9Y8_LUT4AB/E6BEG[10] Tile_X9Y8_LUT4AB/E6BEG[11]
+ Tile_X9Y8_LUT4AB/E6BEG[1] Tile_X9Y8_LUT4AB/E6BEG[2] Tile_X9Y8_LUT4AB/E6BEG[3] Tile_X9Y8_LUT4AB/E6BEG[4]
+ Tile_X9Y8_LUT4AB/E6BEG[5] Tile_X9Y8_LUT4AB/E6BEG[6] Tile_X9Y8_LUT4AB/E6BEG[7] Tile_X9Y8_LUT4AB/E6BEG[8]
+ Tile_X9Y8_LUT4AB/E6BEG[9] Tile_X9Y8_LUT4AB/EE4BEG[0] Tile_X9Y8_LUT4AB/EE4BEG[10]
+ Tile_X9Y8_LUT4AB/EE4BEG[11] Tile_X9Y8_LUT4AB/EE4BEG[12] Tile_X9Y8_LUT4AB/EE4BEG[13]
+ Tile_X9Y8_LUT4AB/EE4BEG[14] Tile_X9Y8_LUT4AB/EE4BEG[15] Tile_X9Y8_LUT4AB/EE4BEG[1]
+ Tile_X9Y8_LUT4AB/EE4BEG[2] Tile_X9Y8_LUT4AB/EE4BEG[3] Tile_X9Y8_LUT4AB/EE4BEG[4]
+ Tile_X9Y8_LUT4AB/EE4BEG[5] Tile_X9Y8_LUT4AB/EE4BEG[6] Tile_X9Y8_LUT4AB/EE4BEG[7]
+ Tile_X9Y8_LUT4AB/EE4BEG[8] Tile_X9Y8_LUT4AB/EE4BEG[9] Tile_X9Y8_LUT4AB/FrameData_O[0]
+ Tile_X9Y8_LUT4AB/FrameData_O[10] Tile_X9Y8_LUT4AB/FrameData_O[11] Tile_X9Y8_LUT4AB/FrameData_O[12]
+ Tile_X9Y8_LUT4AB/FrameData_O[13] Tile_X9Y8_LUT4AB/FrameData_O[14] Tile_X9Y8_LUT4AB/FrameData_O[15]
+ Tile_X9Y8_LUT4AB/FrameData_O[16] Tile_X9Y8_LUT4AB/FrameData_O[17] Tile_X9Y8_LUT4AB/FrameData_O[18]
+ Tile_X9Y8_LUT4AB/FrameData_O[19] Tile_X9Y8_LUT4AB/FrameData_O[1] Tile_X9Y8_LUT4AB/FrameData_O[20]
+ Tile_X9Y8_LUT4AB/FrameData_O[21] Tile_X9Y8_LUT4AB/FrameData_O[22] Tile_X9Y8_LUT4AB/FrameData_O[23]
+ Tile_X9Y8_LUT4AB/FrameData_O[24] Tile_X9Y8_LUT4AB/FrameData_O[25] Tile_X9Y8_LUT4AB/FrameData_O[26]
+ Tile_X9Y8_LUT4AB/FrameData_O[27] Tile_X9Y8_LUT4AB/FrameData_O[28] Tile_X9Y8_LUT4AB/FrameData_O[29]
+ Tile_X9Y8_LUT4AB/FrameData_O[2] Tile_X9Y8_LUT4AB/FrameData_O[30] Tile_X9Y8_LUT4AB/FrameData_O[31]
+ Tile_X9Y8_LUT4AB/FrameData_O[3] Tile_X9Y8_LUT4AB/FrameData_O[4] Tile_X9Y8_LUT4AB/FrameData_O[5]
+ Tile_X9Y8_LUT4AB/FrameData_O[6] Tile_X9Y8_LUT4AB/FrameData_O[7] Tile_X9Y8_LUT4AB/FrameData_O[8]
+ Tile_X9Y8_LUT4AB/FrameData_O[9] Tile_X10Y7_IHP_SRAM/Tile_X0Y1_FrameData_O[0] Tile_X10Y7_IHP_SRAM/Tile_X0Y1_FrameData_O[10]
+ Tile_X10Y7_IHP_SRAM/Tile_X0Y1_FrameData_O[11] Tile_X10Y7_IHP_SRAM/Tile_X0Y1_FrameData_O[12]
+ Tile_X10Y7_IHP_SRAM/Tile_X0Y1_FrameData_O[13] Tile_X10Y7_IHP_SRAM/Tile_X0Y1_FrameData_O[14]
+ Tile_X10Y7_IHP_SRAM/Tile_X0Y1_FrameData_O[15] Tile_X10Y7_IHP_SRAM/Tile_X0Y1_FrameData_O[16]
+ Tile_X10Y7_IHP_SRAM/Tile_X0Y1_FrameData_O[17] Tile_X10Y7_IHP_SRAM/Tile_X0Y1_FrameData_O[18]
+ Tile_X10Y7_IHP_SRAM/Tile_X0Y1_FrameData_O[19] Tile_X10Y7_IHP_SRAM/Tile_X0Y1_FrameData_O[1]
+ Tile_X10Y7_IHP_SRAM/Tile_X0Y1_FrameData_O[20] Tile_X10Y7_IHP_SRAM/Tile_X0Y1_FrameData_O[21]
+ Tile_X10Y7_IHP_SRAM/Tile_X0Y1_FrameData_O[22] Tile_X10Y7_IHP_SRAM/Tile_X0Y1_FrameData_O[23]
+ Tile_X10Y7_IHP_SRAM/Tile_X0Y1_FrameData_O[24] Tile_X10Y7_IHP_SRAM/Tile_X0Y1_FrameData_O[25]
+ Tile_X10Y7_IHP_SRAM/Tile_X0Y1_FrameData_O[26] Tile_X10Y7_IHP_SRAM/Tile_X0Y1_FrameData_O[27]
+ Tile_X10Y7_IHP_SRAM/Tile_X0Y1_FrameData_O[28] Tile_X10Y7_IHP_SRAM/Tile_X0Y1_FrameData_O[29]
+ Tile_X10Y7_IHP_SRAM/Tile_X0Y1_FrameData_O[2] Tile_X10Y7_IHP_SRAM/Tile_X0Y1_FrameData_O[30]
+ Tile_X10Y7_IHP_SRAM/Tile_X0Y1_FrameData_O[31] Tile_X10Y7_IHP_SRAM/Tile_X0Y1_FrameData_O[3]
+ Tile_X10Y7_IHP_SRAM/Tile_X0Y1_FrameData_O[4] Tile_X10Y7_IHP_SRAM/Tile_X0Y1_FrameData_O[5]
+ Tile_X10Y7_IHP_SRAM/Tile_X0Y1_FrameData_O[6] Tile_X10Y7_IHP_SRAM/Tile_X0Y1_FrameData_O[7]
+ Tile_X10Y7_IHP_SRAM/Tile_X0Y1_FrameData_O[8] Tile_X10Y7_IHP_SRAM/Tile_X0Y1_FrameData_O[9]
+ Tile_X10Y7_IHP_SRAM/Tile_X0Y1_FrameStrobe[0] Tile_X10Y7_IHP_SRAM/Tile_X0Y1_FrameStrobe[10]
+ Tile_X10Y7_IHP_SRAM/Tile_X0Y1_FrameStrobe[11] Tile_X10Y7_IHP_SRAM/Tile_X0Y1_FrameStrobe[12]
+ Tile_X10Y7_IHP_SRAM/Tile_X0Y1_FrameStrobe[13] Tile_X10Y7_IHP_SRAM/Tile_X0Y1_FrameStrobe[14]
+ Tile_X10Y7_IHP_SRAM/Tile_X0Y1_FrameStrobe[15] Tile_X10Y7_IHP_SRAM/Tile_X0Y1_FrameStrobe[16]
+ Tile_X10Y7_IHP_SRAM/Tile_X0Y1_FrameStrobe[17] Tile_X10Y7_IHP_SRAM/Tile_X0Y1_FrameStrobe[18]
+ Tile_X10Y7_IHP_SRAM/Tile_X0Y1_FrameStrobe[19] Tile_X10Y7_IHP_SRAM/Tile_X0Y1_FrameStrobe[1]
+ Tile_X10Y7_IHP_SRAM/Tile_X0Y1_FrameStrobe[2] Tile_X10Y7_IHP_SRAM/Tile_X0Y1_FrameStrobe[3]
+ Tile_X10Y7_IHP_SRAM/Tile_X0Y1_FrameStrobe[4] Tile_X10Y7_IHP_SRAM/Tile_X0Y1_FrameStrobe[5]
+ Tile_X10Y7_IHP_SRAM/Tile_X0Y1_FrameStrobe[6] Tile_X10Y7_IHP_SRAM/Tile_X0Y1_FrameStrobe[7]
+ Tile_X10Y7_IHP_SRAM/Tile_X0Y1_FrameStrobe[8] Tile_X10Y7_IHP_SRAM/Tile_X0Y1_FrameStrobe[9]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y0_N1BEG[0] Tile_X10Y9_IHP_SRAM/Tile_X0Y0_N1BEG[1] Tile_X10Y9_IHP_SRAM/Tile_X0Y0_N1BEG[2]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y0_N1BEG[3] Tile_X10Y7_IHP_SRAM/Tile_X0Y1_N2END[0] Tile_X10Y7_IHP_SRAM/Tile_X0Y1_N2END[1]
+ Tile_X10Y7_IHP_SRAM/Tile_X0Y1_N2END[2] Tile_X10Y7_IHP_SRAM/Tile_X0Y1_N2END[3] Tile_X10Y7_IHP_SRAM/Tile_X0Y1_N2END[4]
+ Tile_X10Y7_IHP_SRAM/Tile_X0Y1_N2END[5] Tile_X10Y7_IHP_SRAM/Tile_X0Y1_N2END[6] Tile_X10Y7_IHP_SRAM/Tile_X0Y1_N2END[7]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y0_N2BEG[0] Tile_X10Y9_IHP_SRAM/Tile_X0Y0_N2BEG[1] Tile_X10Y9_IHP_SRAM/Tile_X0Y0_N2BEG[2]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y0_N2BEG[3] Tile_X10Y9_IHP_SRAM/Tile_X0Y0_N2BEG[4] Tile_X10Y9_IHP_SRAM/Tile_X0Y0_N2BEG[5]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y0_N2BEG[6] Tile_X10Y9_IHP_SRAM/Tile_X0Y0_N2BEG[7] Tile_X10Y9_IHP_SRAM/Tile_X0Y0_N4BEG[0]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y0_N4BEG[10] Tile_X10Y9_IHP_SRAM/Tile_X0Y0_N4BEG[11]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y0_N4BEG[12] Tile_X10Y9_IHP_SRAM/Tile_X0Y0_N4BEG[13]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y0_N4BEG[14] Tile_X10Y9_IHP_SRAM/Tile_X0Y0_N4BEG[15]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y0_N4BEG[1] Tile_X10Y9_IHP_SRAM/Tile_X0Y0_N4BEG[2] Tile_X10Y9_IHP_SRAM/Tile_X0Y0_N4BEG[3]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y0_N4BEG[4] Tile_X10Y9_IHP_SRAM/Tile_X0Y0_N4BEG[5] Tile_X10Y9_IHP_SRAM/Tile_X0Y0_N4BEG[6]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y0_N4BEG[7] Tile_X10Y9_IHP_SRAM/Tile_X0Y0_N4BEG[8] Tile_X10Y9_IHP_SRAM/Tile_X0Y0_N4BEG[9]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y0_S1END[0] Tile_X10Y9_IHP_SRAM/Tile_X0Y0_S1END[1] Tile_X10Y9_IHP_SRAM/Tile_X0Y0_S1END[2]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y0_S1END[3] Tile_X10Y9_IHP_SRAM/Tile_X0Y0_S2MID[0] Tile_X10Y9_IHP_SRAM/Tile_X0Y0_S2MID[1]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y0_S2MID[2] Tile_X10Y9_IHP_SRAM/Tile_X0Y0_S2MID[3] Tile_X10Y9_IHP_SRAM/Tile_X0Y0_S2MID[4]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y0_S2MID[5] Tile_X10Y9_IHP_SRAM/Tile_X0Y0_S2MID[6] Tile_X10Y9_IHP_SRAM/Tile_X0Y0_S2MID[7]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y0_S2END[0] Tile_X10Y9_IHP_SRAM/Tile_X0Y0_S2END[1] Tile_X10Y9_IHP_SRAM/Tile_X0Y0_S2END[2]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y0_S2END[3] Tile_X10Y9_IHP_SRAM/Tile_X0Y0_S2END[4] Tile_X10Y9_IHP_SRAM/Tile_X0Y0_S2END[5]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y0_S2END[6] Tile_X10Y9_IHP_SRAM/Tile_X0Y0_S2END[7] Tile_X10Y9_IHP_SRAM/Tile_X0Y0_S4END[0]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y0_S4END[10] Tile_X10Y9_IHP_SRAM/Tile_X0Y0_S4END[11]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y0_S4END[12] Tile_X10Y9_IHP_SRAM/Tile_X0Y0_S4END[13]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y0_S4END[14] Tile_X10Y9_IHP_SRAM/Tile_X0Y0_S4END[15]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y0_S4END[1] Tile_X10Y9_IHP_SRAM/Tile_X0Y0_S4END[2] Tile_X10Y9_IHP_SRAM/Tile_X0Y0_S4END[3]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y0_S4END[4] Tile_X10Y9_IHP_SRAM/Tile_X0Y0_S4END[5] Tile_X10Y9_IHP_SRAM/Tile_X0Y0_S4END[6]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y0_S4END[7] Tile_X10Y9_IHP_SRAM/Tile_X0Y0_S4END[8] Tile_X10Y9_IHP_SRAM/Tile_X0Y0_S4END[9]
+ Tile_X10Y7_IHP_SRAM/Tile_X0Y1_UserCLK Tile_X9Y8_LUT4AB/W1END[0] Tile_X9Y8_LUT4AB/W1END[1]
+ Tile_X9Y8_LUT4AB/W1END[2] Tile_X9Y8_LUT4AB/W1END[3] Tile_X9Y8_LUT4AB/W2MID[0] Tile_X9Y8_LUT4AB/W2MID[1]
+ Tile_X9Y8_LUT4AB/W2MID[2] Tile_X9Y8_LUT4AB/W2MID[3] Tile_X9Y8_LUT4AB/W2MID[4] Tile_X9Y8_LUT4AB/W2MID[5]
+ Tile_X9Y8_LUT4AB/W2MID[6] Tile_X9Y8_LUT4AB/W2MID[7] Tile_X9Y8_LUT4AB/W2END[0] Tile_X9Y8_LUT4AB/W2END[1]
+ Tile_X9Y8_LUT4AB/W2END[2] Tile_X9Y8_LUT4AB/W2END[3] Tile_X9Y8_LUT4AB/W2END[4] Tile_X9Y8_LUT4AB/W2END[5]
+ Tile_X9Y8_LUT4AB/W2END[6] Tile_X9Y8_LUT4AB/W2END[7] Tile_X9Y8_LUT4AB/W6END[0] Tile_X9Y8_LUT4AB/W6END[10]
+ Tile_X9Y8_LUT4AB/W6END[11] Tile_X9Y8_LUT4AB/W6END[1] Tile_X9Y8_LUT4AB/W6END[2] Tile_X9Y8_LUT4AB/W6END[3]
+ Tile_X9Y8_LUT4AB/W6END[4] Tile_X9Y8_LUT4AB/W6END[5] Tile_X9Y8_LUT4AB/W6END[6] Tile_X9Y8_LUT4AB/W6END[7]
+ Tile_X9Y8_LUT4AB/W6END[8] Tile_X9Y8_LUT4AB/W6END[9] Tile_X9Y8_LUT4AB/WW4END[0] Tile_X9Y8_LUT4AB/WW4END[10]
+ Tile_X9Y8_LUT4AB/WW4END[11] Tile_X9Y8_LUT4AB/WW4END[12] Tile_X9Y8_LUT4AB/WW4END[13]
+ Tile_X9Y8_LUT4AB/WW4END[14] Tile_X9Y8_LUT4AB/WW4END[15] Tile_X9Y8_LUT4AB/WW4END[1]
+ Tile_X9Y8_LUT4AB/WW4END[2] Tile_X9Y8_LUT4AB/WW4END[3] Tile_X9Y8_LUT4AB/WW4END[4]
+ Tile_X9Y8_LUT4AB/WW4END[5] Tile_X9Y8_LUT4AB/WW4END[6] Tile_X9Y8_LUT4AB/WW4END[7]
+ Tile_X9Y8_LUT4AB/WW4END[8] Tile_X9Y8_LUT4AB/WW4END[9] VGND VPWR Tile_X10Y8_WEN_SRAM
+ IHP_SRAM
XTile_X9Y5_LUT4AB Tile_X9Y6_LUT4AB/Co Tile_X9Y5_LUT4AB/Co Tile_X9Y5_LUT4AB/E1BEG[0]
+ Tile_X9Y5_LUT4AB/E1BEG[1] Tile_X9Y5_LUT4AB/E1BEG[2] Tile_X9Y5_LUT4AB/E1BEG[3] Tile_X9Y5_LUT4AB/E1END[0]
+ Tile_X9Y5_LUT4AB/E1END[1] Tile_X9Y5_LUT4AB/E1END[2] Tile_X9Y5_LUT4AB/E1END[3] Tile_X9Y5_LUT4AB/E2BEG[0]
+ Tile_X9Y5_LUT4AB/E2BEG[1] Tile_X9Y5_LUT4AB/E2BEG[2] Tile_X9Y5_LUT4AB/E2BEG[3] Tile_X9Y5_LUT4AB/E2BEG[4]
+ Tile_X9Y5_LUT4AB/E2BEG[5] Tile_X9Y5_LUT4AB/E2BEG[6] Tile_X9Y5_LUT4AB/E2BEG[7] Tile_X9Y5_LUT4AB/E2BEGb[0]
+ Tile_X9Y5_LUT4AB/E2BEGb[1] Tile_X9Y5_LUT4AB/E2BEGb[2] Tile_X9Y5_LUT4AB/E2BEGb[3]
+ Tile_X9Y5_LUT4AB/E2BEGb[4] Tile_X9Y5_LUT4AB/E2BEGb[5] Tile_X9Y5_LUT4AB/E2BEGb[6]
+ Tile_X9Y5_LUT4AB/E2BEGb[7] Tile_X9Y5_LUT4AB/E2END[0] Tile_X9Y5_LUT4AB/E2END[1] Tile_X9Y5_LUT4AB/E2END[2]
+ Tile_X9Y5_LUT4AB/E2END[3] Tile_X9Y5_LUT4AB/E2END[4] Tile_X9Y5_LUT4AB/E2END[5] Tile_X9Y5_LUT4AB/E2END[6]
+ Tile_X9Y5_LUT4AB/E2END[7] Tile_X9Y5_LUT4AB/E2MID[0] Tile_X9Y5_LUT4AB/E2MID[1] Tile_X9Y5_LUT4AB/E2MID[2]
+ Tile_X9Y5_LUT4AB/E2MID[3] Tile_X9Y5_LUT4AB/E2MID[4] Tile_X9Y5_LUT4AB/E2MID[5] Tile_X9Y5_LUT4AB/E2MID[6]
+ Tile_X9Y5_LUT4AB/E2MID[7] Tile_X9Y5_LUT4AB/E6BEG[0] Tile_X9Y5_LUT4AB/E6BEG[10] Tile_X9Y5_LUT4AB/E6BEG[11]
+ Tile_X9Y5_LUT4AB/E6BEG[1] Tile_X9Y5_LUT4AB/E6BEG[2] Tile_X9Y5_LUT4AB/E6BEG[3] Tile_X9Y5_LUT4AB/E6BEG[4]
+ Tile_X9Y5_LUT4AB/E6BEG[5] Tile_X9Y5_LUT4AB/E6BEG[6] Tile_X9Y5_LUT4AB/E6BEG[7] Tile_X9Y5_LUT4AB/E6BEG[8]
+ Tile_X9Y5_LUT4AB/E6BEG[9] Tile_X9Y5_LUT4AB/E6END[0] Tile_X9Y5_LUT4AB/E6END[10] Tile_X9Y5_LUT4AB/E6END[11]
+ Tile_X9Y5_LUT4AB/E6END[1] Tile_X9Y5_LUT4AB/E6END[2] Tile_X9Y5_LUT4AB/E6END[3] Tile_X9Y5_LUT4AB/E6END[4]
+ Tile_X9Y5_LUT4AB/E6END[5] Tile_X9Y5_LUT4AB/E6END[6] Tile_X9Y5_LUT4AB/E6END[7] Tile_X9Y5_LUT4AB/E6END[8]
+ Tile_X9Y5_LUT4AB/E6END[9] Tile_X9Y5_LUT4AB/EE4BEG[0] Tile_X9Y5_LUT4AB/EE4BEG[10]
+ Tile_X9Y5_LUT4AB/EE4BEG[11] Tile_X9Y5_LUT4AB/EE4BEG[12] Tile_X9Y5_LUT4AB/EE4BEG[13]
+ Tile_X9Y5_LUT4AB/EE4BEG[14] Tile_X9Y5_LUT4AB/EE4BEG[15] Tile_X9Y5_LUT4AB/EE4BEG[1]
+ Tile_X9Y5_LUT4AB/EE4BEG[2] Tile_X9Y5_LUT4AB/EE4BEG[3] Tile_X9Y5_LUT4AB/EE4BEG[4]
+ Tile_X9Y5_LUT4AB/EE4BEG[5] Tile_X9Y5_LUT4AB/EE4BEG[6] Tile_X9Y5_LUT4AB/EE4BEG[7]
+ Tile_X9Y5_LUT4AB/EE4BEG[8] Tile_X9Y5_LUT4AB/EE4BEG[9] Tile_X9Y5_LUT4AB/EE4END[0]
+ Tile_X9Y5_LUT4AB/EE4END[10] Tile_X9Y5_LUT4AB/EE4END[11] Tile_X9Y5_LUT4AB/EE4END[12]
+ Tile_X9Y5_LUT4AB/EE4END[13] Tile_X9Y5_LUT4AB/EE4END[14] Tile_X9Y5_LUT4AB/EE4END[15]
+ Tile_X9Y5_LUT4AB/EE4END[1] Tile_X9Y5_LUT4AB/EE4END[2] Tile_X9Y5_LUT4AB/EE4END[3]
+ Tile_X9Y5_LUT4AB/EE4END[4] Tile_X9Y5_LUT4AB/EE4END[5] Tile_X9Y5_LUT4AB/EE4END[6]
+ Tile_X9Y5_LUT4AB/EE4END[7] Tile_X9Y5_LUT4AB/EE4END[8] Tile_X9Y5_LUT4AB/EE4END[9]
+ Tile_X9Y5_LUT4AB/FrameData[0] Tile_X9Y5_LUT4AB/FrameData[10] Tile_X9Y5_LUT4AB/FrameData[11]
+ Tile_X9Y5_LUT4AB/FrameData[12] Tile_X9Y5_LUT4AB/FrameData[13] Tile_X9Y5_LUT4AB/FrameData[14]
+ Tile_X9Y5_LUT4AB/FrameData[15] Tile_X9Y5_LUT4AB/FrameData[16] Tile_X9Y5_LUT4AB/FrameData[17]
+ Tile_X9Y5_LUT4AB/FrameData[18] Tile_X9Y5_LUT4AB/FrameData[19] Tile_X9Y5_LUT4AB/FrameData[1]
+ Tile_X9Y5_LUT4AB/FrameData[20] Tile_X9Y5_LUT4AB/FrameData[21] Tile_X9Y5_LUT4AB/FrameData[22]
+ Tile_X9Y5_LUT4AB/FrameData[23] Tile_X9Y5_LUT4AB/FrameData[24] Tile_X9Y5_LUT4AB/FrameData[25]
+ Tile_X9Y5_LUT4AB/FrameData[26] Tile_X9Y5_LUT4AB/FrameData[27] Tile_X9Y5_LUT4AB/FrameData[28]
+ Tile_X9Y5_LUT4AB/FrameData[29] Tile_X9Y5_LUT4AB/FrameData[2] Tile_X9Y5_LUT4AB/FrameData[30]
+ Tile_X9Y5_LUT4AB/FrameData[31] Tile_X9Y5_LUT4AB/FrameData[3] Tile_X9Y5_LUT4AB/FrameData[4]
+ Tile_X9Y5_LUT4AB/FrameData[5] Tile_X9Y5_LUT4AB/FrameData[6] Tile_X9Y5_LUT4AB/FrameData[7]
+ Tile_X9Y5_LUT4AB/FrameData[8] Tile_X9Y5_LUT4AB/FrameData[9] Tile_X9Y5_LUT4AB/FrameData_O[0]
+ Tile_X9Y5_LUT4AB/FrameData_O[10] Tile_X9Y5_LUT4AB/FrameData_O[11] Tile_X9Y5_LUT4AB/FrameData_O[12]
+ Tile_X9Y5_LUT4AB/FrameData_O[13] Tile_X9Y5_LUT4AB/FrameData_O[14] Tile_X9Y5_LUT4AB/FrameData_O[15]
+ Tile_X9Y5_LUT4AB/FrameData_O[16] Tile_X9Y5_LUT4AB/FrameData_O[17] Tile_X9Y5_LUT4AB/FrameData_O[18]
+ Tile_X9Y5_LUT4AB/FrameData_O[19] Tile_X9Y5_LUT4AB/FrameData_O[1] Tile_X9Y5_LUT4AB/FrameData_O[20]
+ Tile_X9Y5_LUT4AB/FrameData_O[21] Tile_X9Y5_LUT4AB/FrameData_O[22] Tile_X9Y5_LUT4AB/FrameData_O[23]
+ Tile_X9Y5_LUT4AB/FrameData_O[24] Tile_X9Y5_LUT4AB/FrameData_O[25] Tile_X9Y5_LUT4AB/FrameData_O[26]
+ Tile_X9Y5_LUT4AB/FrameData_O[27] Tile_X9Y5_LUT4AB/FrameData_O[28] Tile_X9Y5_LUT4AB/FrameData_O[29]
+ Tile_X9Y5_LUT4AB/FrameData_O[2] Tile_X9Y5_LUT4AB/FrameData_O[30] Tile_X9Y5_LUT4AB/FrameData_O[31]
+ Tile_X9Y5_LUT4AB/FrameData_O[3] Tile_X9Y5_LUT4AB/FrameData_O[4] Tile_X9Y5_LUT4AB/FrameData_O[5]
+ Tile_X9Y5_LUT4AB/FrameData_O[6] Tile_X9Y5_LUT4AB/FrameData_O[7] Tile_X9Y5_LUT4AB/FrameData_O[8]
+ Tile_X9Y5_LUT4AB/FrameData_O[9] Tile_X9Y5_LUT4AB/FrameStrobe[0] Tile_X9Y5_LUT4AB/FrameStrobe[10]
+ Tile_X9Y5_LUT4AB/FrameStrobe[11] Tile_X9Y5_LUT4AB/FrameStrobe[12] Tile_X9Y5_LUT4AB/FrameStrobe[13]
+ Tile_X9Y5_LUT4AB/FrameStrobe[14] Tile_X9Y5_LUT4AB/FrameStrobe[15] Tile_X9Y5_LUT4AB/FrameStrobe[16]
+ Tile_X9Y5_LUT4AB/FrameStrobe[17] Tile_X9Y5_LUT4AB/FrameStrobe[18] Tile_X9Y5_LUT4AB/FrameStrobe[19]
+ Tile_X9Y5_LUT4AB/FrameStrobe[1] Tile_X9Y5_LUT4AB/FrameStrobe[2] Tile_X9Y5_LUT4AB/FrameStrobe[3]
+ Tile_X9Y5_LUT4AB/FrameStrobe[4] Tile_X9Y5_LUT4AB/FrameStrobe[5] Tile_X9Y5_LUT4AB/FrameStrobe[6]
+ Tile_X9Y5_LUT4AB/FrameStrobe[7] Tile_X9Y5_LUT4AB/FrameStrobe[8] Tile_X9Y5_LUT4AB/FrameStrobe[9]
+ Tile_X9Y4_LUT4AB/FrameStrobe[0] Tile_X9Y4_LUT4AB/FrameStrobe[10] Tile_X9Y4_LUT4AB/FrameStrobe[11]
+ Tile_X9Y4_LUT4AB/FrameStrobe[12] Tile_X9Y4_LUT4AB/FrameStrobe[13] Tile_X9Y4_LUT4AB/FrameStrobe[14]
+ Tile_X9Y4_LUT4AB/FrameStrobe[15] Tile_X9Y4_LUT4AB/FrameStrobe[16] Tile_X9Y4_LUT4AB/FrameStrobe[17]
+ Tile_X9Y4_LUT4AB/FrameStrobe[18] Tile_X9Y4_LUT4AB/FrameStrobe[19] Tile_X9Y4_LUT4AB/FrameStrobe[1]
+ Tile_X9Y4_LUT4AB/FrameStrobe[2] Tile_X9Y4_LUT4AB/FrameStrobe[3] Tile_X9Y4_LUT4AB/FrameStrobe[4]
+ Tile_X9Y4_LUT4AB/FrameStrobe[5] Tile_X9Y4_LUT4AB/FrameStrobe[6] Tile_X9Y4_LUT4AB/FrameStrobe[7]
+ Tile_X9Y4_LUT4AB/FrameStrobe[8] Tile_X9Y4_LUT4AB/FrameStrobe[9] Tile_X9Y5_LUT4AB/N1BEG[0]
+ Tile_X9Y5_LUT4AB/N1BEG[1] Tile_X9Y5_LUT4AB/N1BEG[2] Tile_X9Y5_LUT4AB/N1BEG[3] Tile_X9Y6_LUT4AB/N1BEG[0]
+ Tile_X9Y6_LUT4AB/N1BEG[1] Tile_X9Y6_LUT4AB/N1BEG[2] Tile_X9Y6_LUT4AB/N1BEG[3] Tile_X9Y5_LUT4AB/N2BEG[0]
+ Tile_X9Y5_LUT4AB/N2BEG[1] Tile_X9Y5_LUT4AB/N2BEG[2] Tile_X9Y5_LUT4AB/N2BEG[3] Tile_X9Y5_LUT4AB/N2BEG[4]
+ Tile_X9Y5_LUT4AB/N2BEG[5] Tile_X9Y5_LUT4AB/N2BEG[6] Tile_X9Y5_LUT4AB/N2BEG[7] Tile_X9Y4_LUT4AB/N2END[0]
+ Tile_X9Y4_LUT4AB/N2END[1] Tile_X9Y4_LUT4AB/N2END[2] Tile_X9Y4_LUT4AB/N2END[3] Tile_X9Y4_LUT4AB/N2END[4]
+ Tile_X9Y4_LUT4AB/N2END[5] Tile_X9Y4_LUT4AB/N2END[6] Tile_X9Y4_LUT4AB/N2END[7] Tile_X9Y5_LUT4AB/N2END[0]
+ Tile_X9Y5_LUT4AB/N2END[1] Tile_X9Y5_LUT4AB/N2END[2] Tile_X9Y5_LUT4AB/N2END[3] Tile_X9Y5_LUT4AB/N2END[4]
+ Tile_X9Y5_LUT4AB/N2END[5] Tile_X9Y5_LUT4AB/N2END[6] Tile_X9Y5_LUT4AB/N2END[7] Tile_X9Y6_LUT4AB/N2BEG[0]
+ Tile_X9Y6_LUT4AB/N2BEG[1] Tile_X9Y6_LUT4AB/N2BEG[2] Tile_X9Y6_LUT4AB/N2BEG[3] Tile_X9Y6_LUT4AB/N2BEG[4]
+ Tile_X9Y6_LUT4AB/N2BEG[5] Tile_X9Y6_LUT4AB/N2BEG[6] Tile_X9Y6_LUT4AB/N2BEG[7] Tile_X9Y5_LUT4AB/N4BEG[0]
+ Tile_X9Y5_LUT4AB/N4BEG[10] Tile_X9Y5_LUT4AB/N4BEG[11] Tile_X9Y5_LUT4AB/N4BEG[12]
+ Tile_X9Y5_LUT4AB/N4BEG[13] Tile_X9Y5_LUT4AB/N4BEG[14] Tile_X9Y5_LUT4AB/N4BEG[15]
+ Tile_X9Y5_LUT4AB/N4BEG[1] Tile_X9Y5_LUT4AB/N4BEG[2] Tile_X9Y5_LUT4AB/N4BEG[3] Tile_X9Y5_LUT4AB/N4BEG[4]
+ Tile_X9Y5_LUT4AB/N4BEG[5] Tile_X9Y5_LUT4AB/N4BEG[6] Tile_X9Y5_LUT4AB/N4BEG[7] Tile_X9Y5_LUT4AB/N4BEG[8]
+ Tile_X9Y5_LUT4AB/N4BEG[9] Tile_X9Y6_LUT4AB/N4BEG[0] Tile_X9Y6_LUT4AB/N4BEG[10] Tile_X9Y6_LUT4AB/N4BEG[11]
+ Tile_X9Y6_LUT4AB/N4BEG[12] Tile_X9Y6_LUT4AB/N4BEG[13] Tile_X9Y6_LUT4AB/N4BEG[14]
+ Tile_X9Y6_LUT4AB/N4BEG[15] Tile_X9Y6_LUT4AB/N4BEG[1] Tile_X9Y6_LUT4AB/N4BEG[2] Tile_X9Y6_LUT4AB/N4BEG[3]
+ Tile_X9Y6_LUT4AB/N4BEG[4] Tile_X9Y6_LUT4AB/N4BEG[5] Tile_X9Y6_LUT4AB/N4BEG[6] Tile_X9Y6_LUT4AB/N4BEG[7]
+ Tile_X9Y6_LUT4AB/N4BEG[8] Tile_X9Y6_LUT4AB/N4BEG[9] Tile_X9Y5_LUT4AB/NN4BEG[0] Tile_X9Y5_LUT4AB/NN4BEG[10]
+ Tile_X9Y5_LUT4AB/NN4BEG[11] Tile_X9Y5_LUT4AB/NN4BEG[12] Tile_X9Y5_LUT4AB/NN4BEG[13]
+ Tile_X9Y5_LUT4AB/NN4BEG[14] Tile_X9Y5_LUT4AB/NN4BEG[15] Tile_X9Y5_LUT4AB/NN4BEG[1]
+ Tile_X9Y5_LUT4AB/NN4BEG[2] Tile_X9Y5_LUT4AB/NN4BEG[3] Tile_X9Y5_LUT4AB/NN4BEG[4]
+ Tile_X9Y5_LUT4AB/NN4BEG[5] Tile_X9Y5_LUT4AB/NN4BEG[6] Tile_X9Y5_LUT4AB/NN4BEG[7]
+ Tile_X9Y5_LUT4AB/NN4BEG[8] Tile_X9Y5_LUT4AB/NN4BEG[9] Tile_X9Y6_LUT4AB/NN4BEG[0]
+ Tile_X9Y6_LUT4AB/NN4BEG[10] Tile_X9Y6_LUT4AB/NN4BEG[11] Tile_X9Y6_LUT4AB/NN4BEG[12]
+ Tile_X9Y6_LUT4AB/NN4BEG[13] Tile_X9Y6_LUT4AB/NN4BEG[14] Tile_X9Y6_LUT4AB/NN4BEG[15]
+ Tile_X9Y6_LUT4AB/NN4BEG[1] Tile_X9Y6_LUT4AB/NN4BEG[2] Tile_X9Y6_LUT4AB/NN4BEG[3]
+ Tile_X9Y6_LUT4AB/NN4BEG[4] Tile_X9Y6_LUT4AB/NN4BEG[5] Tile_X9Y6_LUT4AB/NN4BEG[6]
+ Tile_X9Y6_LUT4AB/NN4BEG[7] Tile_X9Y6_LUT4AB/NN4BEG[8] Tile_X9Y6_LUT4AB/NN4BEG[9]
+ Tile_X9Y6_LUT4AB/S1END[0] Tile_X9Y6_LUT4AB/S1END[1] Tile_X9Y6_LUT4AB/S1END[2] Tile_X9Y6_LUT4AB/S1END[3]
+ Tile_X9Y5_LUT4AB/S1END[0] Tile_X9Y5_LUT4AB/S1END[1] Tile_X9Y5_LUT4AB/S1END[2] Tile_X9Y5_LUT4AB/S1END[3]
+ Tile_X9Y6_LUT4AB/S2MID[0] Tile_X9Y6_LUT4AB/S2MID[1] Tile_X9Y6_LUT4AB/S2MID[2] Tile_X9Y6_LUT4AB/S2MID[3]
+ Tile_X9Y6_LUT4AB/S2MID[4] Tile_X9Y6_LUT4AB/S2MID[5] Tile_X9Y6_LUT4AB/S2MID[6] Tile_X9Y6_LUT4AB/S2MID[7]
+ Tile_X9Y6_LUT4AB/S2END[0] Tile_X9Y6_LUT4AB/S2END[1] Tile_X9Y6_LUT4AB/S2END[2] Tile_X9Y6_LUT4AB/S2END[3]
+ Tile_X9Y6_LUT4AB/S2END[4] Tile_X9Y6_LUT4AB/S2END[5] Tile_X9Y6_LUT4AB/S2END[6] Tile_X9Y6_LUT4AB/S2END[7]
+ Tile_X9Y5_LUT4AB/S2END[0] Tile_X9Y5_LUT4AB/S2END[1] Tile_X9Y5_LUT4AB/S2END[2] Tile_X9Y5_LUT4AB/S2END[3]
+ Tile_X9Y5_LUT4AB/S2END[4] Tile_X9Y5_LUT4AB/S2END[5] Tile_X9Y5_LUT4AB/S2END[6] Tile_X9Y5_LUT4AB/S2END[7]
+ Tile_X9Y5_LUT4AB/S2MID[0] Tile_X9Y5_LUT4AB/S2MID[1] Tile_X9Y5_LUT4AB/S2MID[2] Tile_X9Y5_LUT4AB/S2MID[3]
+ Tile_X9Y5_LUT4AB/S2MID[4] Tile_X9Y5_LUT4AB/S2MID[5] Tile_X9Y5_LUT4AB/S2MID[6] Tile_X9Y5_LUT4AB/S2MID[7]
+ Tile_X9Y6_LUT4AB/S4END[0] Tile_X9Y6_LUT4AB/S4END[10] Tile_X9Y6_LUT4AB/S4END[11]
+ Tile_X9Y6_LUT4AB/S4END[12] Tile_X9Y6_LUT4AB/S4END[13] Tile_X9Y6_LUT4AB/S4END[14]
+ Tile_X9Y6_LUT4AB/S4END[15] Tile_X9Y6_LUT4AB/S4END[1] Tile_X9Y6_LUT4AB/S4END[2] Tile_X9Y6_LUT4AB/S4END[3]
+ Tile_X9Y6_LUT4AB/S4END[4] Tile_X9Y6_LUT4AB/S4END[5] Tile_X9Y6_LUT4AB/S4END[6] Tile_X9Y6_LUT4AB/S4END[7]
+ Tile_X9Y6_LUT4AB/S4END[8] Tile_X9Y6_LUT4AB/S4END[9] Tile_X9Y5_LUT4AB/S4END[0] Tile_X9Y5_LUT4AB/S4END[10]
+ Tile_X9Y5_LUT4AB/S4END[11] Tile_X9Y5_LUT4AB/S4END[12] Tile_X9Y5_LUT4AB/S4END[13]
+ Tile_X9Y5_LUT4AB/S4END[14] Tile_X9Y5_LUT4AB/S4END[15] Tile_X9Y5_LUT4AB/S4END[1]
+ Tile_X9Y5_LUT4AB/S4END[2] Tile_X9Y5_LUT4AB/S4END[3] Tile_X9Y5_LUT4AB/S4END[4] Tile_X9Y5_LUT4AB/S4END[5]
+ Tile_X9Y5_LUT4AB/S4END[6] Tile_X9Y5_LUT4AB/S4END[7] Tile_X9Y5_LUT4AB/S4END[8] Tile_X9Y5_LUT4AB/S4END[9]
+ Tile_X9Y6_LUT4AB/SS4END[0] Tile_X9Y6_LUT4AB/SS4END[10] Tile_X9Y6_LUT4AB/SS4END[11]
+ Tile_X9Y6_LUT4AB/SS4END[12] Tile_X9Y6_LUT4AB/SS4END[13] Tile_X9Y6_LUT4AB/SS4END[14]
+ Tile_X9Y6_LUT4AB/SS4END[15] Tile_X9Y6_LUT4AB/SS4END[1] Tile_X9Y6_LUT4AB/SS4END[2]
+ Tile_X9Y6_LUT4AB/SS4END[3] Tile_X9Y6_LUT4AB/SS4END[4] Tile_X9Y6_LUT4AB/SS4END[5]
+ Tile_X9Y6_LUT4AB/SS4END[6] Tile_X9Y6_LUT4AB/SS4END[7] Tile_X9Y6_LUT4AB/SS4END[8]
+ Tile_X9Y6_LUT4AB/SS4END[9] Tile_X9Y5_LUT4AB/SS4END[0] Tile_X9Y5_LUT4AB/SS4END[10]
+ Tile_X9Y5_LUT4AB/SS4END[11] Tile_X9Y5_LUT4AB/SS4END[12] Tile_X9Y5_LUT4AB/SS4END[13]
+ Tile_X9Y5_LUT4AB/SS4END[14] Tile_X9Y5_LUT4AB/SS4END[15] Tile_X9Y5_LUT4AB/SS4END[1]
+ Tile_X9Y5_LUT4AB/SS4END[2] Tile_X9Y5_LUT4AB/SS4END[3] Tile_X9Y5_LUT4AB/SS4END[4]
+ Tile_X9Y5_LUT4AB/SS4END[5] Tile_X9Y5_LUT4AB/SS4END[6] Tile_X9Y5_LUT4AB/SS4END[7]
+ Tile_X9Y5_LUT4AB/SS4END[8] Tile_X9Y5_LUT4AB/SS4END[9] Tile_X9Y5_LUT4AB/UserCLK Tile_X9Y4_LUT4AB/UserCLK
+ VGND VPWR Tile_X9Y5_LUT4AB/W1BEG[0] Tile_X9Y5_LUT4AB/W1BEG[1] Tile_X9Y5_LUT4AB/W1BEG[2]
+ Tile_X9Y5_LUT4AB/W1BEG[3] Tile_X9Y5_LUT4AB/W1END[0] Tile_X9Y5_LUT4AB/W1END[1] Tile_X9Y5_LUT4AB/W1END[2]
+ Tile_X9Y5_LUT4AB/W1END[3] Tile_X9Y5_LUT4AB/W2BEG[0] Tile_X9Y5_LUT4AB/W2BEG[1] Tile_X9Y5_LUT4AB/W2BEG[2]
+ Tile_X9Y5_LUT4AB/W2BEG[3] Tile_X9Y5_LUT4AB/W2BEG[4] Tile_X9Y5_LUT4AB/W2BEG[5] Tile_X9Y5_LUT4AB/W2BEG[6]
+ Tile_X9Y5_LUT4AB/W2BEG[7] Tile_X8Y5_LUT4AB/W2END[0] Tile_X8Y5_LUT4AB/W2END[1] Tile_X8Y5_LUT4AB/W2END[2]
+ Tile_X8Y5_LUT4AB/W2END[3] Tile_X8Y5_LUT4AB/W2END[4] Tile_X8Y5_LUT4AB/W2END[5] Tile_X8Y5_LUT4AB/W2END[6]
+ Tile_X8Y5_LUT4AB/W2END[7] Tile_X9Y5_LUT4AB/W2END[0] Tile_X9Y5_LUT4AB/W2END[1] Tile_X9Y5_LUT4AB/W2END[2]
+ Tile_X9Y5_LUT4AB/W2END[3] Tile_X9Y5_LUT4AB/W2END[4] Tile_X9Y5_LUT4AB/W2END[5] Tile_X9Y5_LUT4AB/W2END[6]
+ Tile_X9Y5_LUT4AB/W2END[7] Tile_X9Y5_LUT4AB/W2MID[0] Tile_X9Y5_LUT4AB/W2MID[1] Tile_X9Y5_LUT4AB/W2MID[2]
+ Tile_X9Y5_LUT4AB/W2MID[3] Tile_X9Y5_LUT4AB/W2MID[4] Tile_X9Y5_LUT4AB/W2MID[5] Tile_X9Y5_LUT4AB/W2MID[6]
+ Tile_X9Y5_LUT4AB/W2MID[7] Tile_X9Y5_LUT4AB/W6BEG[0] Tile_X9Y5_LUT4AB/W6BEG[10] Tile_X9Y5_LUT4AB/W6BEG[11]
+ Tile_X9Y5_LUT4AB/W6BEG[1] Tile_X9Y5_LUT4AB/W6BEG[2] Tile_X9Y5_LUT4AB/W6BEG[3] Tile_X9Y5_LUT4AB/W6BEG[4]
+ Tile_X9Y5_LUT4AB/W6BEG[5] Tile_X9Y5_LUT4AB/W6BEG[6] Tile_X9Y5_LUT4AB/W6BEG[7] Tile_X9Y5_LUT4AB/W6BEG[8]
+ Tile_X9Y5_LUT4AB/W6BEG[9] Tile_X9Y5_LUT4AB/W6END[0] Tile_X9Y5_LUT4AB/W6END[10] Tile_X9Y5_LUT4AB/W6END[11]
+ Tile_X9Y5_LUT4AB/W6END[1] Tile_X9Y5_LUT4AB/W6END[2] Tile_X9Y5_LUT4AB/W6END[3] Tile_X9Y5_LUT4AB/W6END[4]
+ Tile_X9Y5_LUT4AB/W6END[5] Tile_X9Y5_LUT4AB/W6END[6] Tile_X9Y5_LUT4AB/W6END[7] Tile_X9Y5_LUT4AB/W6END[8]
+ Tile_X9Y5_LUT4AB/W6END[9] Tile_X9Y5_LUT4AB/WW4BEG[0] Tile_X9Y5_LUT4AB/WW4BEG[10]
+ Tile_X9Y5_LUT4AB/WW4BEG[11] Tile_X9Y5_LUT4AB/WW4BEG[12] Tile_X9Y5_LUT4AB/WW4BEG[13]
+ Tile_X9Y5_LUT4AB/WW4BEG[14] Tile_X9Y5_LUT4AB/WW4BEG[15] Tile_X9Y5_LUT4AB/WW4BEG[1]
+ Tile_X9Y5_LUT4AB/WW4BEG[2] Tile_X9Y5_LUT4AB/WW4BEG[3] Tile_X9Y5_LUT4AB/WW4BEG[4]
+ Tile_X9Y5_LUT4AB/WW4BEG[5] Tile_X9Y5_LUT4AB/WW4BEG[6] Tile_X9Y5_LUT4AB/WW4BEG[7]
+ Tile_X9Y5_LUT4AB/WW4BEG[8] Tile_X9Y5_LUT4AB/WW4BEG[9] Tile_X9Y5_LUT4AB/WW4END[0]
+ Tile_X9Y5_LUT4AB/WW4END[10] Tile_X9Y5_LUT4AB/WW4END[11] Tile_X9Y5_LUT4AB/WW4END[12]
+ Tile_X9Y5_LUT4AB/WW4END[13] Tile_X9Y5_LUT4AB/WW4END[14] Tile_X9Y5_LUT4AB/WW4END[15]
+ Tile_X9Y5_LUT4AB/WW4END[1] Tile_X9Y5_LUT4AB/WW4END[2] Tile_X9Y5_LUT4AB/WW4END[3]
+ Tile_X9Y5_LUT4AB/WW4END[4] Tile_X9Y5_LUT4AB/WW4END[5] Tile_X9Y5_LUT4AB/WW4END[6]
+ Tile_X9Y5_LUT4AB/WW4END[7] Tile_X9Y5_LUT4AB/WW4END[8] Tile_X9Y5_LUT4AB/WW4END[9]
+ LUT4AB
XTile_X0Y1_W_IO Tile_X0Y1_A_I_top Tile_X0Y1_A_O_top Tile_X0Y1_A_T_top Tile_X0Y1_A_config_C_bit0
+ Tile_X0Y1_A_config_C_bit1 Tile_X0Y1_A_config_C_bit2 Tile_X0Y1_A_config_C_bit3 Tile_X0Y1_B_I_top
+ Tile_X0Y1_B_O_top Tile_X0Y1_B_T_top Tile_X0Y1_B_config_C_bit0 Tile_X0Y1_B_config_C_bit1
+ Tile_X0Y1_B_config_C_bit2 Tile_X0Y1_B_config_C_bit3 Tile_X0Y1_W_IO/E1BEG[0] Tile_X0Y1_W_IO/E1BEG[1]
+ Tile_X0Y1_W_IO/E1BEG[2] Tile_X0Y1_W_IO/E1BEG[3] Tile_X0Y1_W_IO/E2BEG[0] Tile_X0Y1_W_IO/E2BEG[1]
+ Tile_X0Y1_W_IO/E2BEG[2] Tile_X0Y1_W_IO/E2BEG[3] Tile_X0Y1_W_IO/E2BEG[4] Tile_X0Y1_W_IO/E2BEG[5]
+ Tile_X0Y1_W_IO/E2BEG[6] Tile_X0Y1_W_IO/E2BEG[7] Tile_X0Y1_W_IO/E2BEGb[0] Tile_X0Y1_W_IO/E2BEGb[1]
+ Tile_X0Y1_W_IO/E2BEGb[2] Tile_X0Y1_W_IO/E2BEGb[3] Tile_X0Y1_W_IO/E2BEGb[4] Tile_X0Y1_W_IO/E2BEGb[5]
+ Tile_X0Y1_W_IO/E2BEGb[6] Tile_X0Y1_W_IO/E2BEGb[7] Tile_X0Y1_W_IO/E6BEG[0] Tile_X0Y1_W_IO/E6BEG[10]
+ Tile_X0Y1_W_IO/E6BEG[11] Tile_X0Y1_W_IO/E6BEG[1] Tile_X0Y1_W_IO/E6BEG[2] Tile_X0Y1_W_IO/E6BEG[3]
+ Tile_X0Y1_W_IO/E6BEG[4] Tile_X0Y1_W_IO/E6BEG[5] Tile_X0Y1_W_IO/E6BEG[6] Tile_X0Y1_W_IO/E6BEG[7]
+ Tile_X0Y1_W_IO/E6BEG[8] Tile_X0Y1_W_IO/E6BEG[9] Tile_X0Y1_W_IO/EE4BEG[0] Tile_X0Y1_W_IO/EE4BEG[10]
+ Tile_X0Y1_W_IO/EE4BEG[11] Tile_X0Y1_W_IO/EE4BEG[12] Tile_X0Y1_W_IO/EE4BEG[13] Tile_X0Y1_W_IO/EE4BEG[14]
+ Tile_X0Y1_W_IO/EE4BEG[15] Tile_X0Y1_W_IO/EE4BEG[1] Tile_X0Y1_W_IO/EE4BEG[2] Tile_X0Y1_W_IO/EE4BEG[3]
+ Tile_X0Y1_W_IO/EE4BEG[4] Tile_X0Y1_W_IO/EE4BEG[5] Tile_X0Y1_W_IO/EE4BEG[6] Tile_X0Y1_W_IO/EE4BEG[7]
+ Tile_X0Y1_W_IO/EE4BEG[8] Tile_X0Y1_W_IO/EE4BEG[9] FrameData[32] FrameData[42] FrameData[43]
+ FrameData[44] FrameData[45] FrameData[46] FrameData[47] FrameData[48] FrameData[49]
+ FrameData[50] FrameData[51] FrameData[33] FrameData[52] FrameData[53] FrameData[54]
+ FrameData[55] FrameData[56] FrameData[57] FrameData[58] FrameData[59] FrameData[60]
+ FrameData[61] FrameData[34] FrameData[62] FrameData[63] FrameData[35] FrameData[36]
+ FrameData[37] FrameData[38] FrameData[39] FrameData[40] FrameData[41] Tile_X1Y1_LUT4AB/FrameData[0]
+ Tile_X1Y1_LUT4AB/FrameData[10] Tile_X1Y1_LUT4AB/FrameData[11] Tile_X1Y1_LUT4AB/FrameData[12]
+ Tile_X1Y1_LUT4AB/FrameData[13] Tile_X1Y1_LUT4AB/FrameData[14] Tile_X1Y1_LUT4AB/FrameData[15]
+ Tile_X1Y1_LUT4AB/FrameData[16] Tile_X1Y1_LUT4AB/FrameData[17] Tile_X1Y1_LUT4AB/FrameData[18]
+ Tile_X1Y1_LUT4AB/FrameData[19] Tile_X1Y1_LUT4AB/FrameData[1] Tile_X1Y1_LUT4AB/FrameData[20]
+ Tile_X1Y1_LUT4AB/FrameData[21] Tile_X1Y1_LUT4AB/FrameData[22] Tile_X1Y1_LUT4AB/FrameData[23]
+ Tile_X1Y1_LUT4AB/FrameData[24] Tile_X1Y1_LUT4AB/FrameData[25] Tile_X1Y1_LUT4AB/FrameData[26]
+ Tile_X1Y1_LUT4AB/FrameData[27] Tile_X1Y1_LUT4AB/FrameData[28] Tile_X1Y1_LUT4AB/FrameData[29]
+ Tile_X1Y1_LUT4AB/FrameData[2] Tile_X1Y1_LUT4AB/FrameData[30] Tile_X1Y1_LUT4AB/FrameData[31]
+ Tile_X1Y1_LUT4AB/FrameData[3] Tile_X1Y1_LUT4AB/FrameData[4] Tile_X1Y1_LUT4AB/FrameData[5]
+ Tile_X1Y1_LUT4AB/FrameData[6] Tile_X1Y1_LUT4AB/FrameData[7] Tile_X1Y1_LUT4AB/FrameData[8]
+ Tile_X1Y1_LUT4AB/FrameData[9] Tile_X0Y1_W_IO/FrameStrobe[0] Tile_X0Y1_W_IO/FrameStrobe[10]
+ Tile_X0Y1_W_IO/FrameStrobe[11] Tile_X0Y1_W_IO/FrameStrobe[12] Tile_X0Y1_W_IO/FrameStrobe[13]
+ Tile_X0Y1_W_IO/FrameStrobe[14] Tile_X0Y1_W_IO/FrameStrobe[15] Tile_X0Y1_W_IO/FrameStrobe[16]
+ Tile_X0Y1_W_IO/FrameStrobe[17] Tile_X0Y1_W_IO/FrameStrobe[18] Tile_X0Y1_W_IO/FrameStrobe[19]
+ Tile_X0Y1_W_IO/FrameStrobe[1] Tile_X0Y1_W_IO/FrameStrobe[2] Tile_X0Y1_W_IO/FrameStrobe[3]
+ Tile_X0Y1_W_IO/FrameStrobe[4] Tile_X0Y1_W_IO/FrameStrobe[5] Tile_X0Y1_W_IO/FrameStrobe[6]
+ Tile_X0Y1_W_IO/FrameStrobe[7] Tile_X0Y1_W_IO/FrameStrobe[8] Tile_X0Y1_W_IO/FrameStrobe[9]
+ Tile_X0Y1_W_IO/FrameStrobe_O[0] Tile_X0Y1_W_IO/FrameStrobe_O[10] Tile_X0Y1_W_IO/FrameStrobe_O[11]
+ Tile_X0Y1_W_IO/FrameStrobe_O[12] Tile_X0Y1_W_IO/FrameStrobe_O[13] Tile_X0Y1_W_IO/FrameStrobe_O[14]
+ Tile_X0Y1_W_IO/FrameStrobe_O[15] Tile_X0Y1_W_IO/FrameStrobe_O[16] Tile_X0Y1_W_IO/FrameStrobe_O[17]
+ Tile_X0Y1_W_IO/FrameStrobe_O[18] Tile_X0Y1_W_IO/FrameStrobe_O[19] Tile_X0Y1_W_IO/FrameStrobe_O[1]
+ Tile_X0Y1_W_IO/FrameStrobe_O[2] Tile_X0Y1_W_IO/FrameStrobe_O[3] Tile_X0Y1_W_IO/FrameStrobe_O[4]
+ Tile_X0Y1_W_IO/FrameStrobe_O[5] Tile_X0Y1_W_IO/FrameStrobe_O[6] Tile_X0Y1_W_IO/FrameStrobe_O[7]
+ Tile_X0Y1_W_IO/FrameStrobe_O[8] Tile_X0Y1_W_IO/FrameStrobe_O[9] Tile_X0Y1_W_IO/UserCLK
+ Tile_X0Y1_W_IO/UserCLKo VGND VPWR Tile_X0Y1_W_IO/W1END[0] Tile_X0Y1_W_IO/W1END[1]
+ Tile_X0Y1_W_IO/W1END[2] Tile_X0Y1_W_IO/W1END[3] Tile_X0Y1_W_IO/W2END[0] Tile_X0Y1_W_IO/W2END[1]
+ Tile_X0Y1_W_IO/W2END[2] Tile_X0Y1_W_IO/W2END[3] Tile_X0Y1_W_IO/W2END[4] Tile_X0Y1_W_IO/W2END[5]
+ Tile_X0Y1_W_IO/W2END[6] Tile_X0Y1_W_IO/W2END[7] Tile_X0Y1_W_IO/W2MID[0] Tile_X0Y1_W_IO/W2MID[1]
+ Tile_X0Y1_W_IO/W2MID[2] Tile_X0Y1_W_IO/W2MID[3] Tile_X0Y1_W_IO/W2MID[4] Tile_X0Y1_W_IO/W2MID[5]
+ Tile_X0Y1_W_IO/W2MID[6] Tile_X0Y1_W_IO/W2MID[7] Tile_X0Y1_W_IO/W6END[0] Tile_X0Y1_W_IO/W6END[10]
+ Tile_X0Y1_W_IO/W6END[11] Tile_X0Y1_W_IO/W6END[1] Tile_X0Y1_W_IO/W6END[2] Tile_X0Y1_W_IO/W6END[3]
+ Tile_X0Y1_W_IO/W6END[4] Tile_X0Y1_W_IO/W6END[5] Tile_X0Y1_W_IO/W6END[6] Tile_X0Y1_W_IO/W6END[7]
+ Tile_X0Y1_W_IO/W6END[8] Tile_X0Y1_W_IO/W6END[9] Tile_X0Y1_W_IO/WW4END[0] Tile_X0Y1_W_IO/WW4END[10]
+ Tile_X0Y1_W_IO/WW4END[11] Tile_X0Y1_W_IO/WW4END[12] Tile_X0Y1_W_IO/WW4END[13] Tile_X0Y1_W_IO/WW4END[14]
+ Tile_X0Y1_W_IO/WW4END[15] Tile_X0Y1_W_IO/WW4END[1] Tile_X0Y1_W_IO/WW4END[2] Tile_X0Y1_W_IO/WW4END[3]
+ Tile_X0Y1_W_IO/WW4END[4] Tile_X0Y1_W_IO/WW4END[5] Tile_X0Y1_W_IO/WW4END[6] Tile_X0Y1_W_IO/WW4END[7]
+ Tile_X0Y1_W_IO/WW4END[8] Tile_X0Y1_W_IO/WW4END[9] W_IO
XTile_X2Y12_LUT4AB Tile_X2Y13_LUT4AB/Co Tile_X2Y12_LUT4AB/Co Tile_X3Y12_LUT4AB/E1END[0]
+ Tile_X3Y12_LUT4AB/E1END[1] Tile_X3Y12_LUT4AB/E1END[2] Tile_X3Y12_LUT4AB/E1END[3]
+ Tile_X2Y12_LUT4AB/E1END[0] Tile_X2Y12_LUT4AB/E1END[1] Tile_X2Y12_LUT4AB/E1END[2]
+ Tile_X2Y12_LUT4AB/E1END[3] Tile_X3Y12_LUT4AB/E2MID[0] Tile_X3Y12_LUT4AB/E2MID[1]
+ Tile_X3Y12_LUT4AB/E2MID[2] Tile_X3Y12_LUT4AB/E2MID[3] Tile_X3Y12_LUT4AB/E2MID[4]
+ Tile_X3Y12_LUT4AB/E2MID[5] Tile_X3Y12_LUT4AB/E2MID[6] Tile_X3Y12_LUT4AB/E2MID[7]
+ Tile_X3Y12_LUT4AB/E2END[0] Tile_X3Y12_LUT4AB/E2END[1] Tile_X3Y12_LUT4AB/E2END[2]
+ Tile_X3Y12_LUT4AB/E2END[3] Tile_X3Y12_LUT4AB/E2END[4] Tile_X3Y12_LUT4AB/E2END[5]
+ Tile_X3Y12_LUT4AB/E2END[6] Tile_X3Y12_LUT4AB/E2END[7] Tile_X2Y12_LUT4AB/E2END[0]
+ Tile_X2Y12_LUT4AB/E2END[1] Tile_X2Y12_LUT4AB/E2END[2] Tile_X2Y12_LUT4AB/E2END[3]
+ Tile_X2Y12_LUT4AB/E2END[4] Tile_X2Y12_LUT4AB/E2END[5] Tile_X2Y12_LUT4AB/E2END[6]
+ Tile_X2Y12_LUT4AB/E2END[7] Tile_X2Y12_LUT4AB/E2MID[0] Tile_X2Y12_LUT4AB/E2MID[1]
+ Tile_X2Y12_LUT4AB/E2MID[2] Tile_X2Y12_LUT4AB/E2MID[3] Tile_X2Y12_LUT4AB/E2MID[4]
+ Tile_X2Y12_LUT4AB/E2MID[5] Tile_X2Y12_LUT4AB/E2MID[6] Tile_X2Y12_LUT4AB/E2MID[7]
+ Tile_X3Y12_LUT4AB/E6END[0] Tile_X3Y12_LUT4AB/E6END[10] Tile_X3Y12_LUT4AB/E6END[11]
+ Tile_X3Y12_LUT4AB/E6END[1] Tile_X3Y12_LUT4AB/E6END[2] Tile_X3Y12_LUT4AB/E6END[3]
+ Tile_X3Y12_LUT4AB/E6END[4] Tile_X3Y12_LUT4AB/E6END[5] Tile_X3Y12_LUT4AB/E6END[6]
+ Tile_X3Y12_LUT4AB/E6END[7] Tile_X3Y12_LUT4AB/E6END[8] Tile_X3Y12_LUT4AB/E6END[9]
+ Tile_X2Y12_LUT4AB/E6END[0] Tile_X2Y12_LUT4AB/E6END[10] Tile_X2Y12_LUT4AB/E6END[11]
+ Tile_X2Y12_LUT4AB/E6END[1] Tile_X2Y12_LUT4AB/E6END[2] Tile_X2Y12_LUT4AB/E6END[3]
+ Tile_X2Y12_LUT4AB/E6END[4] Tile_X2Y12_LUT4AB/E6END[5] Tile_X2Y12_LUT4AB/E6END[6]
+ Tile_X2Y12_LUT4AB/E6END[7] Tile_X2Y12_LUT4AB/E6END[8] Tile_X2Y12_LUT4AB/E6END[9]
+ Tile_X3Y12_LUT4AB/EE4END[0] Tile_X3Y12_LUT4AB/EE4END[10] Tile_X3Y12_LUT4AB/EE4END[11]
+ Tile_X3Y12_LUT4AB/EE4END[12] Tile_X3Y12_LUT4AB/EE4END[13] Tile_X3Y12_LUT4AB/EE4END[14]
+ Tile_X3Y12_LUT4AB/EE4END[15] Tile_X3Y12_LUT4AB/EE4END[1] Tile_X3Y12_LUT4AB/EE4END[2]
+ Tile_X3Y12_LUT4AB/EE4END[3] Tile_X3Y12_LUT4AB/EE4END[4] Tile_X3Y12_LUT4AB/EE4END[5]
+ Tile_X3Y12_LUT4AB/EE4END[6] Tile_X3Y12_LUT4AB/EE4END[7] Tile_X3Y12_LUT4AB/EE4END[8]
+ Tile_X3Y12_LUT4AB/EE4END[9] Tile_X2Y12_LUT4AB/EE4END[0] Tile_X2Y12_LUT4AB/EE4END[10]
+ Tile_X2Y12_LUT4AB/EE4END[11] Tile_X2Y12_LUT4AB/EE4END[12] Tile_X2Y12_LUT4AB/EE4END[13]
+ Tile_X2Y12_LUT4AB/EE4END[14] Tile_X2Y12_LUT4AB/EE4END[15] Tile_X2Y12_LUT4AB/EE4END[1]
+ Tile_X2Y12_LUT4AB/EE4END[2] Tile_X2Y12_LUT4AB/EE4END[3] Tile_X2Y12_LUT4AB/EE4END[4]
+ Tile_X2Y12_LUT4AB/EE4END[5] Tile_X2Y12_LUT4AB/EE4END[6] Tile_X2Y12_LUT4AB/EE4END[7]
+ Tile_X2Y12_LUT4AB/EE4END[8] Tile_X2Y12_LUT4AB/EE4END[9] Tile_X2Y12_LUT4AB/FrameData[0]
+ Tile_X2Y12_LUT4AB/FrameData[10] Tile_X2Y12_LUT4AB/FrameData[11] Tile_X2Y12_LUT4AB/FrameData[12]
+ Tile_X2Y12_LUT4AB/FrameData[13] Tile_X2Y12_LUT4AB/FrameData[14] Tile_X2Y12_LUT4AB/FrameData[15]
+ Tile_X2Y12_LUT4AB/FrameData[16] Tile_X2Y12_LUT4AB/FrameData[17] Tile_X2Y12_LUT4AB/FrameData[18]
+ Tile_X2Y12_LUT4AB/FrameData[19] Tile_X2Y12_LUT4AB/FrameData[1] Tile_X2Y12_LUT4AB/FrameData[20]
+ Tile_X2Y12_LUT4AB/FrameData[21] Tile_X2Y12_LUT4AB/FrameData[22] Tile_X2Y12_LUT4AB/FrameData[23]
+ Tile_X2Y12_LUT4AB/FrameData[24] Tile_X2Y12_LUT4AB/FrameData[25] Tile_X2Y12_LUT4AB/FrameData[26]
+ Tile_X2Y12_LUT4AB/FrameData[27] Tile_X2Y12_LUT4AB/FrameData[28] Tile_X2Y12_LUT4AB/FrameData[29]
+ Tile_X2Y12_LUT4AB/FrameData[2] Tile_X2Y12_LUT4AB/FrameData[30] Tile_X2Y12_LUT4AB/FrameData[31]
+ Tile_X2Y12_LUT4AB/FrameData[3] Tile_X2Y12_LUT4AB/FrameData[4] Tile_X2Y12_LUT4AB/FrameData[5]
+ Tile_X2Y12_LUT4AB/FrameData[6] Tile_X2Y12_LUT4AB/FrameData[7] Tile_X2Y12_LUT4AB/FrameData[8]
+ Tile_X2Y12_LUT4AB/FrameData[9] Tile_X3Y12_LUT4AB/FrameData[0] Tile_X3Y12_LUT4AB/FrameData[10]
+ Tile_X3Y12_LUT4AB/FrameData[11] Tile_X3Y12_LUT4AB/FrameData[12] Tile_X3Y12_LUT4AB/FrameData[13]
+ Tile_X3Y12_LUT4AB/FrameData[14] Tile_X3Y12_LUT4AB/FrameData[15] Tile_X3Y12_LUT4AB/FrameData[16]
+ Tile_X3Y12_LUT4AB/FrameData[17] Tile_X3Y12_LUT4AB/FrameData[18] Tile_X3Y12_LUT4AB/FrameData[19]
+ Tile_X3Y12_LUT4AB/FrameData[1] Tile_X3Y12_LUT4AB/FrameData[20] Tile_X3Y12_LUT4AB/FrameData[21]
+ Tile_X3Y12_LUT4AB/FrameData[22] Tile_X3Y12_LUT4AB/FrameData[23] Tile_X3Y12_LUT4AB/FrameData[24]
+ Tile_X3Y12_LUT4AB/FrameData[25] Tile_X3Y12_LUT4AB/FrameData[26] Tile_X3Y12_LUT4AB/FrameData[27]
+ Tile_X3Y12_LUT4AB/FrameData[28] Tile_X3Y12_LUT4AB/FrameData[29] Tile_X3Y12_LUT4AB/FrameData[2]
+ Tile_X3Y12_LUT4AB/FrameData[30] Tile_X3Y12_LUT4AB/FrameData[31] Tile_X3Y12_LUT4AB/FrameData[3]
+ Tile_X3Y12_LUT4AB/FrameData[4] Tile_X3Y12_LUT4AB/FrameData[5] Tile_X3Y12_LUT4AB/FrameData[6]
+ Tile_X3Y12_LUT4AB/FrameData[7] Tile_X3Y12_LUT4AB/FrameData[8] Tile_X3Y12_LUT4AB/FrameData[9]
+ Tile_X2Y12_LUT4AB/FrameStrobe[0] Tile_X2Y12_LUT4AB/FrameStrobe[10] Tile_X2Y12_LUT4AB/FrameStrobe[11]
+ Tile_X2Y12_LUT4AB/FrameStrobe[12] Tile_X2Y12_LUT4AB/FrameStrobe[13] Tile_X2Y12_LUT4AB/FrameStrobe[14]
+ Tile_X2Y12_LUT4AB/FrameStrobe[15] Tile_X2Y12_LUT4AB/FrameStrobe[16] Tile_X2Y12_LUT4AB/FrameStrobe[17]
+ Tile_X2Y12_LUT4AB/FrameStrobe[18] Tile_X2Y12_LUT4AB/FrameStrobe[19] Tile_X2Y12_LUT4AB/FrameStrobe[1]
+ Tile_X2Y12_LUT4AB/FrameStrobe[2] Tile_X2Y12_LUT4AB/FrameStrobe[3] Tile_X2Y12_LUT4AB/FrameStrobe[4]
+ Tile_X2Y12_LUT4AB/FrameStrobe[5] Tile_X2Y12_LUT4AB/FrameStrobe[6] Tile_X2Y12_LUT4AB/FrameStrobe[7]
+ Tile_X2Y12_LUT4AB/FrameStrobe[8] Tile_X2Y12_LUT4AB/FrameStrobe[9] Tile_X2Y11_LUT4AB/FrameStrobe[0]
+ Tile_X2Y11_LUT4AB/FrameStrobe[10] Tile_X2Y11_LUT4AB/FrameStrobe[11] Tile_X2Y11_LUT4AB/FrameStrobe[12]
+ Tile_X2Y11_LUT4AB/FrameStrobe[13] Tile_X2Y11_LUT4AB/FrameStrobe[14] Tile_X2Y11_LUT4AB/FrameStrobe[15]
+ Tile_X2Y11_LUT4AB/FrameStrobe[16] Tile_X2Y11_LUT4AB/FrameStrobe[17] Tile_X2Y11_LUT4AB/FrameStrobe[18]
+ Tile_X2Y11_LUT4AB/FrameStrobe[19] Tile_X2Y11_LUT4AB/FrameStrobe[1] Tile_X2Y11_LUT4AB/FrameStrobe[2]
+ Tile_X2Y11_LUT4AB/FrameStrobe[3] Tile_X2Y11_LUT4AB/FrameStrobe[4] Tile_X2Y11_LUT4AB/FrameStrobe[5]
+ Tile_X2Y11_LUT4AB/FrameStrobe[6] Tile_X2Y11_LUT4AB/FrameStrobe[7] Tile_X2Y11_LUT4AB/FrameStrobe[8]
+ Tile_X2Y11_LUT4AB/FrameStrobe[9] Tile_X2Y12_LUT4AB/N1BEG[0] Tile_X2Y12_LUT4AB/N1BEG[1]
+ Tile_X2Y12_LUT4AB/N1BEG[2] Tile_X2Y12_LUT4AB/N1BEG[3] Tile_X2Y13_LUT4AB/N1BEG[0]
+ Tile_X2Y13_LUT4AB/N1BEG[1] Tile_X2Y13_LUT4AB/N1BEG[2] Tile_X2Y13_LUT4AB/N1BEG[3]
+ Tile_X2Y12_LUT4AB/N2BEG[0] Tile_X2Y12_LUT4AB/N2BEG[1] Tile_X2Y12_LUT4AB/N2BEG[2]
+ Tile_X2Y12_LUT4AB/N2BEG[3] Tile_X2Y12_LUT4AB/N2BEG[4] Tile_X2Y12_LUT4AB/N2BEG[5]
+ Tile_X2Y12_LUT4AB/N2BEG[6] Tile_X2Y12_LUT4AB/N2BEG[7] Tile_X2Y11_LUT4AB/N2END[0]
+ Tile_X2Y11_LUT4AB/N2END[1] Tile_X2Y11_LUT4AB/N2END[2] Tile_X2Y11_LUT4AB/N2END[3]
+ Tile_X2Y11_LUT4AB/N2END[4] Tile_X2Y11_LUT4AB/N2END[5] Tile_X2Y11_LUT4AB/N2END[6]
+ Tile_X2Y11_LUT4AB/N2END[7] Tile_X2Y12_LUT4AB/N2END[0] Tile_X2Y12_LUT4AB/N2END[1]
+ Tile_X2Y12_LUT4AB/N2END[2] Tile_X2Y12_LUT4AB/N2END[3] Tile_X2Y12_LUT4AB/N2END[4]
+ Tile_X2Y12_LUT4AB/N2END[5] Tile_X2Y12_LUT4AB/N2END[6] Tile_X2Y12_LUT4AB/N2END[7]
+ Tile_X2Y13_LUT4AB/N2BEG[0] Tile_X2Y13_LUT4AB/N2BEG[1] Tile_X2Y13_LUT4AB/N2BEG[2]
+ Tile_X2Y13_LUT4AB/N2BEG[3] Tile_X2Y13_LUT4AB/N2BEG[4] Tile_X2Y13_LUT4AB/N2BEG[5]
+ Tile_X2Y13_LUT4AB/N2BEG[6] Tile_X2Y13_LUT4AB/N2BEG[7] Tile_X2Y12_LUT4AB/N4BEG[0]
+ Tile_X2Y12_LUT4AB/N4BEG[10] Tile_X2Y12_LUT4AB/N4BEG[11] Tile_X2Y12_LUT4AB/N4BEG[12]
+ Tile_X2Y12_LUT4AB/N4BEG[13] Tile_X2Y12_LUT4AB/N4BEG[14] Tile_X2Y12_LUT4AB/N4BEG[15]
+ Tile_X2Y12_LUT4AB/N4BEG[1] Tile_X2Y12_LUT4AB/N4BEG[2] Tile_X2Y12_LUT4AB/N4BEG[3]
+ Tile_X2Y12_LUT4AB/N4BEG[4] Tile_X2Y12_LUT4AB/N4BEG[5] Tile_X2Y12_LUT4AB/N4BEG[6]
+ Tile_X2Y12_LUT4AB/N4BEG[7] Tile_X2Y12_LUT4AB/N4BEG[8] Tile_X2Y12_LUT4AB/N4BEG[9]
+ Tile_X2Y13_LUT4AB/N4BEG[0] Tile_X2Y13_LUT4AB/N4BEG[10] Tile_X2Y13_LUT4AB/N4BEG[11]
+ Tile_X2Y13_LUT4AB/N4BEG[12] Tile_X2Y13_LUT4AB/N4BEG[13] Tile_X2Y13_LUT4AB/N4BEG[14]
+ Tile_X2Y13_LUT4AB/N4BEG[15] Tile_X2Y13_LUT4AB/N4BEG[1] Tile_X2Y13_LUT4AB/N4BEG[2]
+ Tile_X2Y13_LUT4AB/N4BEG[3] Tile_X2Y13_LUT4AB/N4BEG[4] Tile_X2Y13_LUT4AB/N4BEG[5]
+ Tile_X2Y13_LUT4AB/N4BEG[6] Tile_X2Y13_LUT4AB/N4BEG[7] Tile_X2Y13_LUT4AB/N4BEG[8]
+ Tile_X2Y13_LUT4AB/N4BEG[9] Tile_X2Y12_LUT4AB/NN4BEG[0] Tile_X2Y12_LUT4AB/NN4BEG[10]
+ Tile_X2Y12_LUT4AB/NN4BEG[11] Tile_X2Y12_LUT4AB/NN4BEG[12] Tile_X2Y12_LUT4AB/NN4BEG[13]
+ Tile_X2Y12_LUT4AB/NN4BEG[14] Tile_X2Y12_LUT4AB/NN4BEG[15] Tile_X2Y12_LUT4AB/NN4BEG[1]
+ Tile_X2Y12_LUT4AB/NN4BEG[2] Tile_X2Y12_LUT4AB/NN4BEG[3] Tile_X2Y12_LUT4AB/NN4BEG[4]
+ Tile_X2Y12_LUT4AB/NN4BEG[5] Tile_X2Y12_LUT4AB/NN4BEG[6] Tile_X2Y12_LUT4AB/NN4BEG[7]
+ Tile_X2Y12_LUT4AB/NN4BEG[8] Tile_X2Y12_LUT4AB/NN4BEG[9] Tile_X2Y13_LUT4AB/NN4BEG[0]
+ Tile_X2Y13_LUT4AB/NN4BEG[10] Tile_X2Y13_LUT4AB/NN4BEG[11] Tile_X2Y13_LUT4AB/NN4BEG[12]
+ Tile_X2Y13_LUT4AB/NN4BEG[13] Tile_X2Y13_LUT4AB/NN4BEG[14] Tile_X2Y13_LUT4AB/NN4BEG[15]
+ Tile_X2Y13_LUT4AB/NN4BEG[1] Tile_X2Y13_LUT4AB/NN4BEG[2] Tile_X2Y13_LUT4AB/NN4BEG[3]
+ Tile_X2Y13_LUT4AB/NN4BEG[4] Tile_X2Y13_LUT4AB/NN4BEG[5] Tile_X2Y13_LUT4AB/NN4BEG[6]
+ Tile_X2Y13_LUT4AB/NN4BEG[7] Tile_X2Y13_LUT4AB/NN4BEG[8] Tile_X2Y13_LUT4AB/NN4BEG[9]
+ Tile_X2Y13_LUT4AB/S1END[0] Tile_X2Y13_LUT4AB/S1END[1] Tile_X2Y13_LUT4AB/S1END[2]
+ Tile_X2Y13_LUT4AB/S1END[3] Tile_X2Y12_LUT4AB/S1END[0] Tile_X2Y12_LUT4AB/S1END[1]
+ Tile_X2Y12_LUT4AB/S1END[2] Tile_X2Y12_LUT4AB/S1END[3] Tile_X2Y13_LUT4AB/S2MID[0]
+ Tile_X2Y13_LUT4AB/S2MID[1] Tile_X2Y13_LUT4AB/S2MID[2] Tile_X2Y13_LUT4AB/S2MID[3]
+ Tile_X2Y13_LUT4AB/S2MID[4] Tile_X2Y13_LUT4AB/S2MID[5] Tile_X2Y13_LUT4AB/S2MID[6]
+ Tile_X2Y13_LUT4AB/S2MID[7] Tile_X2Y13_LUT4AB/S2END[0] Tile_X2Y13_LUT4AB/S2END[1]
+ Tile_X2Y13_LUT4AB/S2END[2] Tile_X2Y13_LUT4AB/S2END[3] Tile_X2Y13_LUT4AB/S2END[4]
+ Tile_X2Y13_LUT4AB/S2END[5] Tile_X2Y13_LUT4AB/S2END[6] Tile_X2Y13_LUT4AB/S2END[7]
+ Tile_X2Y12_LUT4AB/S2END[0] Tile_X2Y12_LUT4AB/S2END[1] Tile_X2Y12_LUT4AB/S2END[2]
+ Tile_X2Y12_LUT4AB/S2END[3] Tile_X2Y12_LUT4AB/S2END[4] Tile_X2Y12_LUT4AB/S2END[5]
+ Tile_X2Y12_LUT4AB/S2END[6] Tile_X2Y12_LUT4AB/S2END[7] Tile_X2Y12_LUT4AB/S2MID[0]
+ Tile_X2Y12_LUT4AB/S2MID[1] Tile_X2Y12_LUT4AB/S2MID[2] Tile_X2Y12_LUT4AB/S2MID[3]
+ Tile_X2Y12_LUT4AB/S2MID[4] Tile_X2Y12_LUT4AB/S2MID[5] Tile_X2Y12_LUT4AB/S2MID[6]
+ Tile_X2Y12_LUT4AB/S2MID[7] Tile_X2Y13_LUT4AB/S4END[0] Tile_X2Y13_LUT4AB/S4END[10]
+ Tile_X2Y13_LUT4AB/S4END[11] Tile_X2Y13_LUT4AB/S4END[12] Tile_X2Y13_LUT4AB/S4END[13]
+ Tile_X2Y13_LUT4AB/S4END[14] Tile_X2Y13_LUT4AB/S4END[15] Tile_X2Y13_LUT4AB/S4END[1]
+ Tile_X2Y13_LUT4AB/S4END[2] Tile_X2Y13_LUT4AB/S4END[3] Tile_X2Y13_LUT4AB/S4END[4]
+ Tile_X2Y13_LUT4AB/S4END[5] Tile_X2Y13_LUT4AB/S4END[6] Tile_X2Y13_LUT4AB/S4END[7]
+ Tile_X2Y13_LUT4AB/S4END[8] Tile_X2Y13_LUT4AB/S4END[9] Tile_X2Y12_LUT4AB/S4END[0]
+ Tile_X2Y12_LUT4AB/S4END[10] Tile_X2Y12_LUT4AB/S4END[11] Tile_X2Y12_LUT4AB/S4END[12]
+ Tile_X2Y12_LUT4AB/S4END[13] Tile_X2Y12_LUT4AB/S4END[14] Tile_X2Y12_LUT4AB/S4END[15]
+ Tile_X2Y12_LUT4AB/S4END[1] Tile_X2Y12_LUT4AB/S4END[2] Tile_X2Y12_LUT4AB/S4END[3]
+ Tile_X2Y12_LUT4AB/S4END[4] Tile_X2Y12_LUT4AB/S4END[5] Tile_X2Y12_LUT4AB/S4END[6]
+ Tile_X2Y12_LUT4AB/S4END[7] Tile_X2Y12_LUT4AB/S4END[8] Tile_X2Y12_LUT4AB/S4END[9]
+ Tile_X2Y13_LUT4AB/SS4END[0] Tile_X2Y13_LUT4AB/SS4END[10] Tile_X2Y13_LUT4AB/SS4END[11]
+ Tile_X2Y13_LUT4AB/SS4END[12] Tile_X2Y13_LUT4AB/SS4END[13] Tile_X2Y13_LUT4AB/SS4END[14]
+ Tile_X2Y13_LUT4AB/SS4END[15] Tile_X2Y13_LUT4AB/SS4END[1] Tile_X2Y13_LUT4AB/SS4END[2]
+ Tile_X2Y13_LUT4AB/SS4END[3] Tile_X2Y13_LUT4AB/SS4END[4] Tile_X2Y13_LUT4AB/SS4END[5]
+ Tile_X2Y13_LUT4AB/SS4END[6] Tile_X2Y13_LUT4AB/SS4END[7] Tile_X2Y13_LUT4AB/SS4END[8]
+ Tile_X2Y13_LUT4AB/SS4END[9] Tile_X2Y12_LUT4AB/SS4END[0] Tile_X2Y12_LUT4AB/SS4END[10]
+ Tile_X2Y12_LUT4AB/SS4END[11] Tile_X2Y12_LUT4AB/SS4END[12] Tile_X2Y12_LUT4AB/SS4END[13]
+ Tile_X2Y12_LUT4AB/SS4END[14] Tile_X2Y12_LUT4AB/SS4END[15] Tile_X2Y12_LUT4AB/SS4END[1]
+ Tile_X2Y12_LUT4AB/SS4END[2] Tile_X2Y12_LUT4AB/SS4END[3] Tile_X2Y12_LUT4AB/SS4END[4]
+ Tile_X2Y12_LUT4AB/SS4END[5] Tile_X2Y12_LUT4AB/SS4END[6] Tile_X2Y12_LUT4AB/SS4END[7]
+ Tile_X2Y12_LUT4AB/SS4END[8] Tile_X2Y12_LUT4AB/SS4END[9] Tile_X2Y12_LUT4AB/UserCLK
+ Tile_X2Y11_LUT4AB/UserCLK VGND VPWR Tile_X2Y12_LUT4AB/W1BEG[0] Tile_X2Y12_LUT4AB/W1BEG[1]
+ Tile_X2Y12_LUT4AB/W1BEG[2] Tile_X2Y12_LUT4AB/W1BEG[3] Tile_X3Y12_LUT4AB/W1BEG[0]
+ Tile_X3Y12_LUT4AB/W1BEG[1] Tile_X3Y12_LUT4AB/W1BEG[2] Tile_X3Y12_LUT4AB/W1BEG[3]
+ Tile_X2Y12_LUT4AB/W2BEG[0] Tile_X2Y12_LUT4AB/W2BEG[1] Tile_X2Y12_LUT4AB/W2BEG[2]
+ Tile_X2Y12_LUT4AB/W2BEG[3] Tile_X2Y12_LUT4AB/W2BEG[4] Tile_X2Y12_LUT4AB/W2BEG[5]
+ Tile_X2Y12_LUT4AB/W2BEG[6] Tile_X2Y12_LUT4AB/W2BEG[7] Tile_X1Y12_LUT4AB/W2END[0]
+ Tile_X1Y12_LUT4AB/W2END[1] Tile_X1Y12_LUT4AB/W2END[2] Tile_X1Y12_LUT4AB/W2END[3]
+ Tile_X1Y12_LUT4AB/W2END[4] Tile_X1Y12_LUT4AB/W2END[5] Tile_X1Y12_LUT4AB/W2END[6]
+ Tile_X1Y12_LUT4AB/W2END[7] Tile_X2Y12_LUT4AB/W2END[0] Tile_X2Y12_LUT4AB/W2END[1]
+ Tile_X2Y12_LUT4AB/W2END[2] Tile_X2Y12_LUT4AB/W2END[3] Tile_X2Y12_LUT4AB/W2END[4]
+ Tile_X2Y12_LUT4AB/W2END[5] Tile_X2Y12_LUT4AB/W2END[6] Tile_X2Y12_LUT4AB/W2END[7]
+ Tile_X3Y12_LUT4AB/W2BEG[0] Tile_X3Y12_LUT4AB/W2BEG[1] Tile_X3Y12_LUT4AB/W2BEG[2]
+ Tile_X3Y12_LUT4AB/W2BEG[3] Tile_X3Y12_LUT4AB/W2BEG[4] Tile_X3Y12_LUT4AB/W2BEG[5]
+ Tile_X3Y12_LUT4AB/W2BEG[6] Tile_X3Y12_LUT4AB/W2BEG[7] Tile_X2Y12_LUT4AB/W6BEG[0]
+ Tile_X2Y12_LUT4AB/W6BEG[10] Tile_X2Y12_LUT4AB/W6BEG[11] Tile_X2Y12_LUT4AB/W6BEG[1]
+ Tile_X2Y12_LUT4AB/W6BEG[2] Tile_X2Y12_LUT4AB/W6BEG[3] Tile_X2Y12_LUT4AB/W6BEG[4]
+ Tile_X2Y12_LUT4AB/W6BEG[5] Tile_X2Y12_LUT4AB/W6BEG[6] Tile_X2Y12_LUT4AB/W6BEG[7]
+ Tile_X2Y12_LUT4AB/W6BEG[8] Tile_X2Y12_LUT4AB/W6BEG[9] Tile_X3Y12_LUT4AB/W6BEG[0]
+ Tile_X3Y12_LUT4AB/W6BEG[10] Tile_X3Y12_LUT4AB/W6BEG[11] Tile_X3Y12_LUT4AB/W6BEG[1]
+ Tile_X3Y12_LUT4AB/W6BEG[2] Tile_X3Y12_LUT4AB/W6BEG[3] Tile_X3Y12_LUT4AB/W6BEG[4]
+ Tile_X3Y12_LUT4AB/W6BEG[5] Tile_X3Y12_LUT4AB/W6BEG[6] Tile_X3Y12_LUT4AB/W6BEG[7]
+ Tile_X3Y12_LUT4AB/W6BEG[8] Tile_X3Y12_LUT4AB/W6BEG[9] Tile_X2Y12_LUT4AB/WW4BEG[0]
+ Tile_X2Y12_LUT4AB/WW4BEG[10] Tile_X2Y12_LUT4AB/WW4BEG[11] Tile_X2Y12_LUT4AB/WW4BEG[12]
+ Tile_X2Y12_LUT4AB/WW4BEG[13] Tile_X2Y12_LUT4AB/WW4BEG[14] Tile_X2Y12_LUT4AB/WW4BEG[15]
+ Tile_X2Y12_LUT4AB/WW4BEG[1] Tile_X2Y12_LUT4AB/WW4BEG[2] Tile_X2Y12_LUT4AB/WW4BEG[3]
+ Tile_X2Y12_LUT4AB/WW4BEG[4] Tile_X2Y12_LUT4AB/WW4BEG[5] Tile_X2Y12_LUT4AB/WW4BEG[6]
+ Tile_X2Y12_LUT4AB/WW4BEG[7] Tile_X2Y12_LUT4AB/WW4BEG[8] Tile_X2Y12_LUT4AB/WW4BEG[9]
+ Tile_X3Y12_LUT4AB/WW4BEG[0] Tile_X3Y12_LUT4AB/WW4BEG[10] Tile_X3Y12_LUT4AB/WW4BEG[11]
+ Tile_X3Y12_LUT4AB/WW4BEG[12] Tile_X3Y12_LUT4AB/WW4BEG[13] Tile_X3Y12_LUT4AB/WW4BEG[14]
+ Tile_X3Y12_LUT4AB/WW4BEG[15] Tile_X3Y12_LUT4AB/WW4BEG[1] Tile_X3Y12_LUT4AB/WW4BEG[2]
+ Tile_X3Y12_LUT4AB/WW4BEG[3] Tile_X3Y12_LUT4AB/WW4BEG[4] Tile_X3Y12_LUT4AB/WW4BEG[5]
+ Tile_X3Y12_LUT4AB/WW4BEG[6] Tile_X3Y12_LUT4AB/WW4BEG[7] Tile_X3Y12_LUT4AB/WW4BEG[8]
+ Tile_X3Y12_LUT4AB/WW4BEG[9] LUT4AB
XTile_X5Y4_LUT4AB Tile_X5Y5_LUT4AB/Co Tile_X5Y4_LUT4AB/Co Tile_X6Y4_LUT4AB/E1END[0]
+ Tile_X6Y4_LUT4AB/E1END[1] Tile_X6Y4_LUT4AB/E1END[2] Tile_X6Y4_LUT4AB/E1END[3] Tile_X5Y4_LUT4AB/E1END[0]
+ Tile_X5Y4_LUT4AB/E1END[1] Tile_X5Y4_LUT4AB/E1END[2] Tile_X5Y4_LUT4AB/E1END[3] Tile_X6Y4_LUT4AB/E2MID[0]
+ Tile_X6Y4_LUT4AB/E2MID[1] Tile_X6Y4_LUT4AB/E2MID[2] Tile_X6Y4_LUT4AB/E2MID[3] Tile_X6Y4_LUT4AB/E2MID[4]
+ Tile_X6Y4_LUT4AB/E2MID[5] Tile_X6Y4_LUT4AB/E2MID[6] Tile_X6Y4_LUT4AB/E2MID[7] Tile_X6Y4_LUT4AB/E2END[0]
+ Tile_X6Y4_LUT4AB/E2END[1] Tile_X6Y4_LUT4AB/E2END[2] Tile_X6Y4_LUT4AB/E2END[3] Tile_X6Y4_LUT4AB/E2END[4]
+ Tile_X6Y4_LUT4AB/E2END[5] Tile_X6Y4_LUT4AB/E2END[6] Tile_X6Y4_LUT4AB/E2END[7] Tile_X5Y4_LUT4AB/E2END[0]
+ Tile_X5Y4_LUT4AB/E2END[1] Tile_X5Y4_LUT4AB/E2END[2] Tile_X5Y4_LUT4AB/E2END[3] Tile_X5Y4_LUT4AB/E2END[4]
+ Tile_X5Y4_LUT4AB/E2END[5] Tile_X5Y4_LUT4AB/E2END[6] Tile_X5Y4_LUT4AB/E2END[7] Tile_X5Y4_LUT4AB/E2MID[0]
+ Tile_X5Y4_LUT4AB/E2MID[1] Tile_X5Y4_LUT4AB/E2MID[2] Tile_X5Y4_LUT4AB/E2MID[3] Tile_X5Y4_LUT4AB/E2MID[4]
+ Tile_X5Y4_LUT4AB/E2MID[5] Tile_X5Y4_LUT4AB/E2MID[6] Tile_X5Y4_LUT4AB/E2MID[7] Tile_X6Y4_LUT4AB/E6END[0]
+ Tile_X6Y4_LUT4AB/E6END[10] Tile_X6Y4_LUT4AB/E6END[11] Tile_X6Y4_LUT4AB/E6END[1]
+ Tile_X6Y4_LUT4AB/E6END[2] Tile_X6Y4_LUT4AB/E6END[3] Tile_X6Y4_LUT4AB/E6END[4] Tile_X6Y4_LUT4AB/E6END[5]
+ Tile_X6Y4_LUT4AB/E6END[6] Tile_X6Y4_LUT4AB/E6END[7] Tile_X6Y4_LUT4AB/E6END[8] Tile_X6Y4_LUT4AB/E6END[9]
+ Tile_X5Y4_LUT4AB/E6END[0] Tile_X5Y4_LUT4AB/E6END[10] Tile_X5Y4_LUT4AB/E6END[11]
+ Tile_X5Y4_LUT4AB/E6END[1] Tile_X5Y4_LUT4AB/E6END[2] Tile_X5Y4_LUT4AB/E6END[3] Tile_X5Y4_LUT4AB/E6END[4]
+ Tile_X5Y4_LUT4AB/E6END[5] Tile_X5Y4_LUT4AB/E6END[6] Tile_X5Y4_LUT4AB/E6END[7] Tile_X5Y4_LUT4AB/E6END[8]
+ Tile_X5Y4_LUT4AB/E6END[9] Tile_X6Y4_LUT4AB/EE4END[0] Tile_X6Y4_LUT4AB/EE4END[10]
+ Tile_X6Y4_LUT4AB/EE4END[11] Tile_X6Y4_LUT4AB/EE4END[12] Tile_X6Y4_LUT4AB/EE4END[13]
+ Tile_X6Y4_LUT4AB/EE4END[14] Tile_X6Y4_LUT4AB/EE4END[15] Tile_X6Y4_LUT4AB/EE4END[1]
+ Tile_X6Y4_LUT4AB/EE4END[2] Tile_X6Y4_LUT4AB/EE4END[3] Tile_X6Y4_LUT4AB/EE4END[4]
+ Tile_X6Y4_LUT4AB/EE4END[5] Tile_X6Y4_LUT4AB/EE4END[6] Tile_X6Y4_LUT4AB/EE4END[7]
+ Tile_X6Y4_LUT4AB/EE4END[8] Tile_X6Y4_LUT4AB/EE4END[9] Tile_X5Y4_LUT4AB/EE4END[0]
+ Tile_X5Y4_LUT4AB/EE4END[10] Tile_X5Y4_LUT4AB/EE4END[11] Tile_X5Y4_LUT4AB/EE4END[12]
+ Tile_X5Y4_LUT4AB/EE4END[13] Tile_X5Y4_LUT4AB/EE4END[14] Tile_X5Y4_LUT4AB/EE4END[15]
+ Tile_X5Y4_LUT4AB/EE4END[1] Tile_X5Y4_LUT4AB/EE4END[2] Tile_X5Y4_LUT4AB/EE4END[3]
+ Tile_X5Y4_LUT4AB/EE4END[4] Tile_X5Y4_LUT4AB/EE4END[5] Tile_X5Y4_LUT4AB/EE4END[6]
+ Tile_X5Y4_LUT4AB/EE4END[7] Tile_X5Y4_LUT4AB/EE4END[8] Tile_X5Y4_LUT4AB/EE4END[9]
+ Tile_X5Y4_LUT4AB/FrameData[0] Tile_X5Y4_LUT4AB/FrameData[10] Tile_X5Y4_LUT4AB/FrameData[11]
+ Tile_X5Y4_LUT4AB/FrameData[12] Tile_X5Y4_LUT4AB/FrameData[13] Tile_X5Y4_LUT4AB/FrameData[14]
+ Tile_X5Y4_LUT4AB/FrameData[15] Tile_X5Y4_LUT4AB/FrameData[16] Tile_X5Y4_LUT4AB/FrameData[17]
+ Tile_X5Y4_LUT4AB/FrameData[18] Tile_X5Y4_LUT4AB/FrameData[19] Tile_X5Y4_LUT4AB/FrameData[1]
+ Tile_X5Y4_LUT4AB/FrameData[20] Tile_X5Y4_LUT4AB/FrameData[21] Tile_X5Y4_LUT4AB/FrameData[22]
+ Tile_X5Y4_LUT4AB/FrameData[23] Tile_X5Y4_LUT4AB/FrameData[24] Tile_X5Y4_LUT4AB/FrameData[25]
+ Tile_X5Y4_LUT4AB/FrameData[26] Tile_X5Y4_LUT4AB/FrameData[27] Tile_X5Y4_LUT4AB/FrameData[28]
+ Tile_X5Y4_LUT4AB/FrameData[29] Tile_X5Y4_LUT4AB/FrameData[2] Tile_X5Y4_LUT4AB/FrameData[30]
+ Tile_X5Y4_LUT4AB/FrameData[31] Tile_X5Y4_LUT4AB/FrameData[3] Tile_X5Y4_LUT4AB/FrameData[4]
+ Tile_X5Y4_LUT4AB/FrameData[5] Tile_X5Y4_LUT4AB/FrameData[6] Tile_X5Y4_LUT4AB/FrameData[7]
+ Tile_X5Y4_LUT4AB/FrameData[8] Tile_X5Y4_LUT4AB/FrameData[9] Tile_X6Y4_LUT4AB/FrameData[0]
+ Tile_X6Y4_LUT4AB/FrameData[10] Tile_X6Y4_LUT4AB/FrameData[11] Tile_X6Y4_LUT4AB/FrameData[12]
+ Tile_X6Y4_LUT4AB/FrameData[13] Tile_X6Y4_LUT4AB/FrameData[14] Tile_X6Y4_LUT4AB/FrameData[15]
+ Tile_X6Y4_LUT4AB/FrameData[16] Tile_X6Y4_LUT4AB/FrameData[17] Tile_X6Y4_LUT4AB/FrameData[18]
+ Tile_X6Y4_LUT4AB/FrameData[19] Tile_X6Y4_LUT4AB/FrameData[1] Tile_X6Y4_LUT4AB/FrameData[20]
+ Tile_X6Y4_LUT4AB/FrameData[21] Tile_X6Y4_LUT4AB/FrameData[22] Tile_X6Y4_LUT4AB/FrameData[23]
+ Tile_X6Y4_LUT4AB/FrameData[24] Tile_X6Y4_LUT4AB/FrameData[25] Tile_X6Y4_LUT4AB/FrameData[26]
+ Tile_X6Y4_LUT4AB/FrameData[27] Tile_X6Y4_LUT4AB/FrameData[28] Tile_X6Y4_LUT4AB/FrameData[29]
+ Tile_X6Y4_LUT4AB/FrameData[2] Tile_X6Y4_LUT4AB/FrameData[30] Tile_X6Y4_LUT4AB/FrameData[31]
+ Tile_X6Y4_LUT4AB/FrameData[3] Tile_X6Y4_LUT4AB/FrameData[4] Tile_X6Y4_LUT4AB/FrameData[5]
+ Tile_X6Y4_LUT4AB/FrameData[6] Tile_X6Y4_LUT4AB/FrameData[7] Tile_X6Y4_LUT4AB/FrameData[8]
+ Tile_X6Y4_LUT4AB/FrameData[9] Tile_X5Y4_LUT4AB/FrameStrobe[0] Tile_X5Y4_LUT4AB/FrameStrobe[10]
+ Tile_X5Y4_LUT4AB/FrameStrobe[11] Tile_X5Y4_LUT4AB/FrameStrobe[12] Tile_X5Y4_LUT4AB/FrameStrobe[13]
+ Tile_X5Y4_LUT4AB/FrameStrobe[14] Tile_X5Y4_LUT4AB/FrameStrobe[15] Tile_X5Y4_LUT4AB/FrameStrobe[16]
+ Tile_X5Y4_LUT4AB/FrameStrobe[17] Tile_X5Y4_LUT4AB/FrameStrobe[18] Tile_X5Y4_LUT4AB/FrameStrobe[19]
+ Tile_X5Y4_LUT4AB/FrameStrobe[1] Tile_X5Y4_LUT4AB/FrameStrobe[2] Tile_X5Y4_LUT4AB/FrameStrobe[3]
+ Tile_X5Y4_LUT4AB/FrameStrobe[4] Tile_X5Y4_LUT4AB/FrameStrobe[5] Tile_X5Y4_LUT4AB/FrameStrobe[6]
+ Tile_X5Y4_LUT4AB/FrameStrobe[7] Tile_X5Y4_LUT4AB/FrameStrobe[8] Tile_X5Y4_LUT4AB/FrameStrobe[9]
+ Tile_X5Y3_LUT4AB/FrameStrobe[0] Tile_X5Y3_LUT4AB/FrameStrobe[10] Tile_X5Y3_LUT4AB/FrameStrobe[11]
+ Tile_X5Y3_LUT4AB/FrameStrobe[12] Tile_X5Y3_LUT4AB/FrameStrobe[13] Tile_X5Y3_LUT4AB/FrameStrobe[14]
+ Tile_X5Y3_LUT4AB/FrameStrobe[15] Tile_X5Y3_LUT4AB/FrameStrobe[16] Tile_X5Y3_LUT4AB/FrameStrobe[17]
+ Tile_X5Y3_LUT4AB/FrameStrobe[18] Tile_X5Y3_LUT4AB/FrameStrobe[19] Tile_X5Y3_LUT4AB/FrameStrobe[1]
+ Tile_X5Y3_LUT4AB/FrameStrobe[2] Tile_X5Y3_LUT4AB/FrameStrobe[3] Tile_X5Y3_LUT4AB/FrameStrobe[4]
+ Tile_X5Y3_LUT4AB/FrameStrobe[5] Tile_X5Y3_LUT4AB/FrameStrobe[6] Tile_X5Y3_LUT4AB/FrameStrobe[7]
+ Tile_X5Y3_LUT4AB/FrameStrobe[8] Tile_X5Y3_LUT4AB/FrameStrobe[9] Tile_X5Y4_LUT4AB/N1BEG[0]
+ Tile_X5Y4_LUT4AB/N1BEG[1] Tile_X5Y4_LUT4AB/N1BEG[2] Tile_X5Y4_LUT4AB/N1BEG[3] Tile_X5Y5_LUT4AB/N1BEG[0]
+ Tile_X5Y5_LUT4AB/N1BEG[1] Tile_X5Y5_LUT4AB/N1BEG[2] Tile_X5Y5_LUT4AB/N1BEG[3] Tile_X5Y4_LUT4AB/N2BEG[0]
+ Tile_X5Y4_LUT4AB/N2BEG[1] Tile_X5Y4_LUT4AB/N2BEG[2] Tile_X5Y4_LUT4AB/N2BEG[3] Tile_X5Y4_LUT4AB/N2BEG[4]
+ Tile_X5Y4_LUT4AB/N2BEG[5] Tile_X5Y4_LUT4AB/N2BEG[6] Tile_X5Y4_LUT4AB/N2BEG[7] Tile_X5Y3_LUT4AB/N2END[0]
+ Tile_X5Y3_LUT4AB/N2END[1] Tile_X5Y3_LUT4AB/N2END[2] Tile_X5Y3_LUT4AB/N2END[3] Tile_X5Y3_LUT4AB/N2END[4]
+ Tile_X5Y3_LUT4AB/N2END[5] Tile_X5Y3_LUT4AB/N2END[6] Tile_X5Y3_LUT4AB/N2END[7] Tile_X5Y4_LUT4AB/N2END[0]
+ Tile_X5Y4_LUT4AB/N2END[1] Tile_X5Y4_LUT4AB/N2END[2] Tile_X5Y4_LUT4AB/N2END[3] Tile_X5Y4_LUT4AB/N2END[4]
+ Tile_X5Y4_LUT4AB/N2END[5] Tile_X5Y4_LUT4AB/N2END[6] Tile_X5Y4_LUT4AB/N2END[7] Tile_X5Y5_LUT4AB/N2BEG[0]
+ Tile_X5Y5_LUT4AB/N2BEG[1] Tile_X5Y5_LUT4AB/N2BEG[2] Tile_X5Y5_LUT4AB/N2BEG[3] Tile_X5Y5_LUT4AB/N2BEG[4]
+ Tile_X5Y5_LUT4AB/N2BEG[5] Tile_X5Y5_LUT4AB/N2BEG[6] Tile_X5Y5_LUT4AB/N2BEG[7] Tile_X5Y4_LUT4AB/N4BEG[0]
+ Tile_X5Y4_LUT4AB/N4BEG[10] Tile_X5Y4_LUT4AB/N4BEG[11] Tile_X5Y4_LUT4AB/N4BEG[12]
+ Tile_X5Y4_LUT4AB/N4BEG[13] Tile_X5Y4_LUT4AB/N4BEG[14] Tile_X5Y4_LUT4AB/N4BEG[15]
+ Tile_X5Y4_LUT4AB/N4BEG[1] Tile_X5Y4_LUT4AB/N4BEG[2] Tile_X5Y4_LUT4AB/N4BEG[3] Tile_X5Y4_LUT4AB/N4BEG[4]
+ Tile_X5Y4_LUT4AB/N4BEG[5] Tile_X5Y4_LUT4AB/N4BEG[6] Tile_X5Y4_LUT4AB/N4BEG[7] Tile_X5Y4_LUT4AB/N4BEG[8]
+ Tile_X5Y4_LUT4AB/N4BEG[9] Tile_X5Y5_LUT4AB/N4BEG[0] Tile_X5Y5_LUT4AB/N4BEG[10] Tile_X5Y5_LUT4AB/N4BEG[11]
+ Tile_X5Y5_LUT4AB/N4BEG[12] Tile_X5Y5_LUT4AB/N4BEG[13] Tile_X5Y5_LUT4AB/N4BEG[14]
+ Tile_X5Y5_LUT4AB/N4BEG[15] Tile_X5Y5_LUT4AB/N4BEG[1] Tile_X5Y5_LUT4AB/N4BEG[2] Tile_X5Y5_LUT4AB/N4BEG[3]
+ Tile_X5Y5_LUT4AB/N4BEG[4] Tile_X5Y5_LUT4AB/N4BEG[5] Tile_X5Y5_LUT4AB/N4BEG[6] Tile_X5Y5_LUT4AB/N4BEG[7]
+ Tile_X5Y5_LUT4AB/N4BEG[8] Tile_X5Y5_LUT4AB/N4BEG[9] Tile_X5Y4_LUT4AB/NN4BEG[0] Tile_X5Y4_LUT4AB/NN4BEG[10]
+ Tile_X5Y4_LUT4AB/NN4BEG[11] Tile_X5Y4_LUT4AB/NN4BEG[12] Tile_X5Y4_LUT4AB/NN4BEG[13]
+ Tile_X5Y4_LUT4AB/NN4BEG[14] Tile_X5Y4_LUT4AB/NN4BEG[15] Tile_X5Y4_LUT4AB/NN4BEG[1]
+ Tile_X5Y4_LUT4AB/NN4BEG[2] Tile_X5Y4_LUT4AB/NN4BEG[3] Tile_X5Y4_LUT4AB/NN4BEG[4]
+ Tile_X5Y4_LUT4AB/NN4BEG[5] Tile_X5Y4_LUT4AB/NN4BEG[6] Tile_X5Y4_LUT4AB/NN4BEG[7]
+ Tile_X5Y4_LUT4AB/NN4BEG[8] Tile_X5Y4_LUT4AB/NN4BEG[9] Tile_X5Y5_LUT4AB/NN4BEG[0]
+ Tile_X5Y5_LUT4AB/NN4BEG[10] Tile_X5Y5_LUT4AB/NN4BEG[11] Tile_X5Y5_LUT4AB/NN4BEG[12]
+ Tile_X5Y5_LUT4AB/NN4BEG[13] Tile_X5Y5_LUT4AB/NN4BEG[14] Tile_X5Y5_LUT4AB/NN4BEG[15]
+ Tile_X5Y5_LUT4AB/NN4BEG[1] Tile_X5Y5_LUT4AB/NN4BEG[2] Tile_X5Y5_LUT4AB/NN4BEG[3]
+ Tile_X5Y5_LUT4AB/NN4BEG[4] Tile_X5Y5_LUT4AB/NN4BEG[5] Tile_X5Y5_LUT4AB/NN4BEG[6]
+ Tile_X5Y5_LUT4AB/NN4BEG[7] Tile_X5Y5_LUT4AB/NN4BEG[8] Tile_X5Y5_LUT4AB/NN4BEG[9]
+ Tile_X5Y5_LUT4AB/S1END[0] Tile_X5Y5_LUT4AB/S1END[1] Tile_X5Y5_LUT4AB/S1END[2] Tile_X5Y5_LUT4AB/S1END[3]
+ Tile_X5Y4_LUT4AB/S1END[0] Tile_X5Y4_LUT4AB/S1END[1] Tile_X5Y4_LUT4AB/S1END[2] Tile_X5Y4_LUT4AB/S1END[3]
+ Tile_X5Y5_LUT4AB/S2MID[0] Tile_X5Y5_LUT4AB/S2MID[1] Tile_X5Y5_LUT4AB/S2MID[2] Tile_X5Y5_LUT4AB/S2MID[3]
+ Tile_X5Y5_LUT4AB/S2MID[4] Tile_X5Y5_LUT4AB/S2MID[5] Tile_X5Y5_LUT4AB/S2MID[6] Tile_X5Y5_LUT4AB/S2MID[7]
+ Tile_X5Y5_LUT4AB/S2END[0] Tile_X5Y5_LUT4AB/S2END[1] Tile_X5Y5_LUT4AB/S2END[2] Tile_X5Y5_LUT4AB/S2END[3]
+ Tile_X5Y5_LUT4AB/S2END[4] Tile_X5Y5_LUT4AB/S2END[5] Tile_X5Y5_LUT4AB/S2END[6] Tile_X5Y5_LUT4AB/S2END[7]
+ Tile_X5Y4_LUT4AB/S2END[0] Tile_X5Y4_LUT4AB/S2END[1] Tile_X5Y4_LUT4AB/S2END[2] Tile_X5Y4_LUT4AB/S2END[3]
+ Tile_X5Y4_LUT4AB/S2END[4] Tile_X5Y4_LUT4AB/S2END[5] Tile_X5Y4_LUT4AB/S2END[6] Tile_X5Y4_LUT4AB/S2END[7]
+ Tile_X5Y4_LUT4AB/S2MID[0] Tile_X5Y4_LUT4AB/S2MID[1] Tile_X5Y4_LUT4AB/S2MID[2] Tile_X5Y4_LUT4AB/S2MID[3]
+ Tile_X5Y4_LUT4AB/S2MID[4] Tile_X5Y4_LUT4AB/S2MID[5] Tile_X5Y4_LUT4AB/S2MID[6] Tile_X5Y4_LUT4AB/S2MID[7]
+ Tile_X5Y5_LUT4AB/S4END[0] Tile_X5Y5_LUT4AB/S4END[10] Tile_X5Y5_LUT4AB/S4END[11]
+ Tile_X5Y5_LUT4AB/S4END[12] Tile_X5Y5_LUT4AB/S4END[13] Tile_X5Y5_LUT4AB/S4END[14]
+ Tile_X5Y5_LUT4AB/S4END[15] Tile_X5Y5_LUT4AB/S4END[1] Tile_X5Y5_LUT4AB/S4END[2] Tile_X5Y5_LUT4AB/S4END[3]
+ Tile_X5Y5_LUT4AB/S4END[4] Tile_X5Y5_LUT4AB/S4END[5] Tile_X5Y5_LUT4AB/S4END[6] Tile_X5Y5_LUT4AB/S4END[7]
+ Tile_X5Y5_LUT4AB/S4END[8] Tile_X5Y5_LUT4AB/S4END[9] Tile_X5Y4_LUT4AB/S4END[0] Tile_X5Y4_LUT4AB/S4END[10]
+ Tile_X5Y4_LUT4AB/S4END[11] Tile_X5Y4_LUT4AB/S4END[12] Tile_X5Y4_LUT4AB/S4END[13]
+ Tile_X5Y4_LUT4AB/S4END[14] Tile_X5Y4_LUT4AB/S4END[15] Tile_X5Y4_LUT4AB/S4END[1]
+ Tile_X5Y4_LUT4AB/S4END[2] Tile_X5Y4_LUT4AB/S4END[3] Tile_X5Y4_LUT4AB/S4END[4] Tile_X5Y4_LUT4AB/S4END[5]
+ Tile_X5Y4_LUT4AB/S4END[6] Tile_X5Y4_LUT4AB/S4END[7] Tile_X5Y4_LUT4AB/S4END[8] Tile_X5Y4_LUT4AB/S4END[9]
+ Tile_X5Y5_LUT4AB/SS4END[0] Tile_X5Y5_LUT4AB/SS4END[10] Tile_X5Y5_LUT4AB/SS4END[11]
+ Tile_X5Y5_LUT4AB/SS4END[12] Tile_X5Y5_LUT4AB/SS4END[13] Tile_X5Y5_LUT4AB/SS4END[14]
+ Tile_X5Y5_LUT4AB/SS4END[15] Tile_X5Y5_LUT4AB/SS4END[1] Tile_X5Y5_LUT4AB/SS4END[2]
+ Tile_X5Y5_LUT4AB/SS4END[3] Tile_X5Y5_LUT4AB/SS4END[4] Tile_X5Y5_LUT4AB/SS4END[5]
+ Tile_X5Y5_LUT4AB/SS4END[6] Tile_X5Y5_LUT4AB/SS4END[7] Tile_X5Y5_LUT4AB/SS4END[8]
+ Tile_X5Y5_LUT4AB/SS4END[9] Tile_X5Y4_LUT4AB/SS4END[0] Tile_X5Y4_LUT4AB/SS4END[10]
+ Tile_X5Y4_LUT4AB/SS4END[11] Tile_X5Y4_LUT4AB/SS4END[12] Tile_X5Y4_LUT4AB/SS4END[13]
+ Tile_X5Y4_LUT4AB/SS4END[14] Tile_X5Y4_LUT4AB/SS4END[15] Tile_X5Y4_LUT4AB/SS4END[1]
+ Tile_X5Y4_LUT4AB/SS4END[2] Tile_X5Y4_LUT4AB/SS4END[3] Tile_X5Y4_LUT4AB/SS4END[4]
+ Tile_X5Y4_LUT4AB/SS4END[5] Tile_X5Y4_LUT4AB/SS4END[6] Tile_X5Y4_LUT4AB/SS4END[7]
+ Tile_X5Y4_LUT4AB/SS4END[8] Tile_X5Y4_LUT4AB/SS4END[9] Tile_X5Y4_LUT4AB/UserCLK Tile_X5Y3_LUT4AB/UserCLK
+ VGND VPWR Tile_X5Y4_LUT4AB/W1BEG[0] Tile_X5Y4_LUT4AB/W1BEG[1] Tile_X5Y4_LUT4AB/W1BEG[2]
+ Tile_X5Y4_LUT4AB/W1BEG[3] Tile_X6Y4_LUT4AB/W1BEG[0] Tile_X6Y4_LUT4AB/W1BEG[1] Tile_X6Y4_LUT4AB/W1BEG[2]
+ Tile_X6Y4_LUT4AB/W1BEG[3] Tile_X5Y4_LUT4AB/W2BEG[0] Tile_X5Y4_LUT4AB/W2BEG[1] Tile_X5Y4_LUT4AB/W2BEG[2]
+ Tile_X5Y4_LUT4AB/W2BEG[3] Tile_X5Y4_LUT4AB/W2BEG[4] Tile_X5Y4_LUT4AB/W2BEG[5] Tile_X5Y4_LUT4AB/W2BEG[6]
+ Tile_X5Y4_LUT4AB/W2BEG[7] Tile_X5Y4_LUT4AB/W2BEGb[0] Tile_X5Y4_LUT4AB/W2BEGb[1]
+ Tile_X5Y4_LUT4AB/W2BEGb[2] Tile_X5Y4_LUT4AB/W2BEGb[3] Tile_X5Y4_LUT4AB/W2BEGb[4]
+ Tile_X5Y4_LUT4AB/W2BEGb[5] Tile_X5Y4_LUT4AB/W2BEGb[6] Tile_X5Y4_LUT4AB/W2BEGb[7]
+ Tile_X5Y4_LUT4AB/W2END[0] Tile_X5Y4_LUT4AB/W2END[1] Tile_X5Y4_LUT4AB/W2END[2] Tile_X5Y4_LUT4AB/W2END[3]
+ Tile_X5Y4_LUT4AB/W2END[4] Tile_X5Y4_LUT4AB/W2END[5] Tile_X5Y4_LUT4AB/W2END[6] Tile_X5Y4_LUT4AB/W2END[7]
+ Tile_X6Y4_LUT4AB/W2BEG[0] Tile_X6Y4_LUT4AB/W2BEG[1] Tile_X6Y4_LUT4AB/W2BEG[2] Tile_X6Y4_LUT4AB/W2BEG[3]
+ Tile_X6Y4_LUT4AB/W2BEG[4] Tile_X6Y4_LUT4AB/W2BEG[5] Tile_X6Y4_LUT4AB/W2BEG[6] Tile_X6Y4_LUT4AB/W2BEG[7]
+ Tile_X5Y4_LUT4AB/W6BEG[0] Tile_X5Y4_LUT4AB/W6BEG[10] Tile_X5Y4_LUT4AB/W6BEG[11]
+ Tile_X5Y4_LUT4AB/W6BEG[1] Tile_X5Y4_LUT4AB/W6BEG[2] Tile_X5Y4_LUT4AB/W6BEG[3] Tile_X5Y4_LUT4AB/W6BEG[4]
+ Tile_X5Y4_LUT4AB/W6BEG[5] Tile_X5Y4_LUT4AB/W6BEG[6] Tile_X5Y4_LUT4AB/W6BEG[7] Tile_X5Y4_LUT4AB/W6BEG[8]
+ Tile_X5Y4_LUT4AB/W6BEG[9] Tile_X6Y4_LUT4AB/W6BEG[0] Tile_X6Y4_LUT4AB/W6BEG[10] Tile_X6Y4_LUT4AB/W6BEG[11]
+ Tile_X6Y4_LUT4AB/W6BEG[1] Tile_X6Y4_LUT4AB/W6BEG[2] Tile_X6Y4_LUT4AB/W6BEG[3] Tile_X6Y4_LUT4AB/W6BEG[4]
+ Tile_X6Y4_LUT4AB/W6BEG[5] Tile_X6Y4_LUT4AB/W6BEG[6] Tile_X6Y4_LUT4AB/W6BEG[7] Tile_X6Y4_LUT4AB/W6BEG[8]
+ Tile_X6Y4_LUT4AB/W6BEG[9] Tile_X5Y4_LUT4AB/WW4BEG[0] Tile_X5Y4_LUT4AB/WW4BEG[10]
+ Tile_X5Y4_LUT4AB/WW4BEG[11] Tile_X5Y4_LUT4AB/WW4BEG[12] Tile_X5Y4_LUT4AB/WW4BEG[13]
+ Tile_X5Y4_LUT4AB/WW4BEG[14] Tile_X5Y4_LUT4AB/WW4BEG[15] Tile_X5Y4_LUT4AB/WW4BEG[1]
+ Tile_X5Y4_LUT4AB/WW4BEG[2] Tile_X5Y4_LUT4AB/WW4BEG[3] Tile_X5Y4_LUT4AB/WW4BEG[4]
+ Tile_X5Y4_LUT4AB/WW4BEG[5] Tile_X5Y4_LUT4AB/WW4BEG[6] Tile_X5Y4_LUT4AB/WW4BEG[7]
+ Tile_X5Y4_LUT4AB/WW4BEG[8] Tile_X5Y4_LUT4AB/WW4BEG[9] Tile_X6Y4_LUT4AB/WW4BEG[0]
+ Tile_X6Y4_LUT4AB/WW4BEG[10] Tile_X6Y4_LUT4AB/WW4BEG[11] Tile_X6Y4_LUT4AB/WW4BEG[12]
+ Tile_X6Y4_LUT4AB/WW4BEG[13] Tile_X6Y4_LUT4AB/WW4BEG[14] Tile_X6Y4_LUT4AB/WW4BEG[15]
+ Tile_X6Y4_LUT4AB/WW4BEG[1] Tile_X6Y4_LUT4AB/WW4BEG[2] Tile_X6Y4_LUT4AB/WW4BEG[3]
+ Tile_X6Y4_LUT4AB/WW4BEG[4] Tile_X6Y4_LUT4AB/WW4BEG[5] Tile_X6Y4_LUT4AB/WW4BEG[6]
+ Tile_X6Y4_LUT4AB/WW4BEG[7] Tile_X6Y4_LUT4AB/WW4BEG[8] Tile_X6Y4_LUT4AB/WW4BEG[9]
+ LUT4AB
XTile_X4Y10_RegFile Tile_X5Y10_LUT4AB/E1END[0] Tile_X5Y10_LUT4AB/E1END[1] Tile_X5Y10_LUT4AB/E1END[2]
+ Tile_X5Y10_LUT4AB/E1END[3] Tile_X3Y10_LUT4AB/E1BEG[0] Tile_X3Y10_LUT4AB/E1BEG[1]
+ Tile_X3Y10_LUT4AB/E1BEG[2] Tile_X3Y10_LUT4AB/E1BEG[3] Tile_X5Y10_LUT4AB/E2MID[0]
+ Tile_X5Y10_LUT4AB/E2MID[1] Tile_X5Y10_LUT4AB/E2MID[2] Tile_X5Y10_LUT4AB/E2MID[3]
+ Tile_X5Y10_LUT4AB/E2MID[4] Tile_X5Y10_LUT4AB/E2MID[5] Tile_X5Y10_LUT4AB/E2MID[6]
+ Tile_X5Y10_LUT4AB/E2MID[7] Tile_X5Y10_LUT4AB/E2END[0] Tile_X5Y10_LUT4AB/E2END[1]
+ Tile_X5Y10_LUT4AB/E2END[2] Tile_X5Y10_LUT4AB/E2END[3] Tile_X5Y10_LUT4AB/E2END[4]
+ Tile_X5Y10_LUT4AB/E2END[5] Tile_X5Y10_LUT4AB/E2END[6] Tile_X5Y10_LUT4AB/E2END[7]
+ Tile_X4Y10_RegFile/E2END[0] Tile_X4Y10_RegFile/E2END[1] Tile_X4Y10_RegFile/E2END[2]
+ Tile_X4Y10_RegFile/E2END[3] Tile_X4Y10_RegFile/E2END[4] Tile_X4Y10_RegFile/E2END[5]
+ Tile_X4Y10_RegFile/E2END[6] Tile_X4Y10_RegFile/E2END[7] Tile_X3Y10_LUT4AB/E2BEG[0]
+ Tile_X3Y10_LUT4AB/E2BEG[1] Tile_X3Y10_LUT4AB/E2BEG[2] Tile_X3Y10_LUT4AB/E2BEG[3]
+ Tile_X3Y10_LUT4AB/E2BEG[4] Tile_X3Y10_LUT4AB/E2BEG[5] Tile_X3Y10_LUT4AB/E2BEG[6]
+ Tile_X3Y10_LUT4AB/E2BEG[7] Tile_X5Y10_LUT4AB/E6END[0] Tile_X5Y10_LUT4AB/E6END[10]
+ Tile_X5Y10_LUT4AB/E6END[11] Tile_X5Y10_LUT4AB/E6END[1] Tile_X5Y10_LUT4AB/E6END[2]
+ Tile_X5Y10_LUT4AB/E6END[3] Tile_X5Y10_LUT4AB/E6END[4] Tile_X5Y10_LUT4AB/E6END[5]
+ Tile_X5Y10_LUT4AB/E6END[6] Tile_X5Y10_LUT4AB/E6END[7] Tile_X5Y10_LUT4AB/E6END[8]
+ Tile_X5Y10_LUT4AB/E6END[9] Tile_X3Y10_LUT4AB/E6BEG[0] Tile_X3Y10_LUT4AB/E6BEG[10]
+ Tile_X3Y10_LUT4AB/E6BEG[11] Tile_X3Y10_LUT4AB/E6BEG[1] Tile_X3Y10_LUT4AB/E6BEG[2]
+ Tile_X3Y10_LUT4AB/E6BEG[3] Tile_X3Y10_LUT4AB/E6BEG[4] Tile_X3Y10_LUT4AB/E6BEG[5]
+ Tile_X3Y10_LUT4AB/E6BEG[6] Tile_X3Y10_LUT4AB/E6BEG[7] Tile_X3Y10_LUT4AB/E6BEG[8]
+ Tile_X3Y10_LUT4AB/E6BEG[9] Tile_X5Y10_LUT4AB/EE4END[0] Tile_X5Y10_LUT4AB/EE4END[10]
+ Tile_X5Y10_LUT4AB/EE4END[11] Tile_X5Y10_LUT4AB/EE4END[12] Tile_X5Y10_LUT4AB/EE4END[13]
+ Tile_X5Y10_LUT4AB/EE4END[14] Tile_X5Y10_LUT4AB/EE4END[15] Tile_X5Y10_LUT4AB/EE4END[1]
+ Tile_X5Y10_LUT4AB/EE4END[2] Tile_X5Y10_LUT4AB/EE4END[3] Tile_X5Y10_LUT4AB/EE4END[4]
+ Tile_X5Y10_LUT4AB/EE4END[5] Tile_X5Y10_LUT4AB/EE4END[6] Tile_X5Y10_LUT4AB/EE4END[7]
+ Tile_X5Y10_LUT4AB/EE4END[8] Tile_X5Y10_LUT4AB/EE4END[9] Tile_X3Y10_LUT4AB/EE4BEG[0]
+ Tile_X3Y10_LUT4AB/EE4BEG[10] Tile_X3Y10_LUT4AB/EE4BEG[11] Tile_X3Y10_LUT4AB/EE4BEG[12]
+ Tile_X3Y10_LUT4AB/EE4BEG[13] Tile_X3Y10_LUT4AB/EE4BEG[14] Tile_X3Y10_LUT4AB/EE4BEG[15]
+ Tile_X3Y10_LUT4AB/EE4BEG[1] Tile_X3Y10_LUT4AB/EE4BEG[2] Tile_X3Y10_LUT4AB/EE4BEG[3]
+ Tile_X3Y10_LUT4AB/EE4BEG[4] Tile_X3Y10_LUT4AB/EE4BEG[5] Tile_X3Y10_LUT4AB/EE4BEG[6]
+ Tile_X3Y10_LUT4AB/EE4BEG[7] Tile_X3Y10_LUT4AB/EE4BEG[8] Tile_X3Y10_LUT4AB/EE4BEG[9]
+ Tile_X4Y10_RegFile/FrameData[0] Tile_X4Y10_RegFile/FrameData[10] Tile_X4Y10_RegFile/FrameData[11]
+ Tile_X4Y10_RegFile/FrameData[12] Tile_X4Y10_RegFile/FrameData[13] Tile_X4Y10_RegFile/FrameData[14]
+ Tile_X4Y10_RegFile/FrameData[15] Tile_X4Y10_RegFile/FrameData[16] Tile_X4Y10_RegFile/FrameData[17]
+ Tile_X4Y10_RegFile/FrameData[18] Tile_X4Y10_RegFile/FrameData[19] Tile_X4Y10_RegFile/FrameData[1]
+ Tile_X4Y10_RegFile/FrameData[20] Tile_X4Y10_RegFile/FrameData[21] Tile_X4Y10_RegFile/FrameData[22]
+ Tile_X4Y10_RegFile/FrameData[23] Tile_X4Y10_RegFile/FrameData[24] Tile_X4Y10_RegFile/FrameData[25]
+ Tile_X4Y10_RegFile/FrameData[26] Tile_X4Y10_RegFile/FrameData[27] Tile_X4Y10_RegFile/FrameData[28]
+ Tile_X4Y10_RegFile/FrameData[29] Tile_X4Y10_RegFile/FrameData[2] Tile_X4Y10_RegFile/FrameData[30]
+ Tile_X4Y10_RegFile/FrameData[31] Tile_X4Y10_RegFile/FrameData[3] Tile_X4Y10_RegFile/FrameData[4]
+ Tile_X4Y10_RegFile/FrameData[5] Tile_X4Y10_RegFile/FrameData[6] Tile_X4Y10_RegFile/FrameData[7]
+ Tile_X4Y10_RegFile/FrameData[8] Tile_X4Y10_RegFile/FrameData[9] Tile_X5Y10_LUT4AB/FrameData[0]
+ Tile_X5Y10_LUT4AB/FrameData[10] Tile_X5Y10_LUT4AB/FrameData[11] Tile_X5Y10_LUT4AB/FrameData[12]
+ Tile_X5Y10_LUT4AB/FrameData[13] Tile_X5Y10_LUT4AB/FrameData[14] Tile_X5Y10_LUT4AB/FrameData[15]
+ Tile_X5Y10_LUT4AB/FrameData[16] Tile_X5Y10_LUT4AB/FrameData[17] Tile_X5Y10_LUT4AB/FrameData[18]
+ Tile_X5Y10_LUT4AB/FrameData[19] Tile_X5Y10_LUT4AB/FrameData[1] Tile_X5Y10_LUT4AB/FrameData[20]
+ Tile_X5Y10_LUT4AB/FrameData[21] Tile_X5Y10_LUT4AB/FrameData[22] Tile_X5Y10_LUT4AB/FrameData[23]
+ Tile_X5Y10_LUT4AB/FrameData[24] Tile_X5Y10_LUT4AB/FrameData[25] Tile_X5Y10_LUT4AB/FrameData[26]
+ Tile_X5Y10_LUT4AB/FrameData[27] Tile_X5Y10_LUT4AB/FrameData[28] Tile_X5Y10_LUT4AB/FrameData[29]
+ Tile_X5Y10_LUT4AB/FrameData[2] Tile_X5Y10_LUT4AB/FrameData[30] Tile_X5Y10_LUT4AB/FrameData[31]
+ Tile_X5Y10_LUT4AB/FrameData[3] Tile_X5Y10_LUT4AB/FrameData[4] Tile_X5Y10_LUT4AB/FrameData[5]
+ Tile_X5Y10_LUT4AB/FrameData[6] Tile_X5Y10_LUT4AB/FrameData[7] Tile_X5Y10_LUT4AB/FrameData[8]
+ Tile_X5Y10_LUT4AB/FrameData[9] Tile_X4Y10_RegFile/FrameStrobe[0] Tile_X4Y10_RegFile/FrameStrobe[10]
+ Tile_X4Y10_RegFile/FrameStrobe[11] Tile_X4Y10_RegFile/FrameStrobe[12] Tile_X4Y10_RegFile/FrameStrobe[13]
+ Tile_X4Y10_RegFile/FrameStrobe[14] Tile_X4Y10_RegFile/FrameStrobe[15] Tile_X4Y10_RegFile/FrameStrobe[16]
+ Tile_X4Y10_RegFile/FrameStrobe[17] Tile_X4Y10_RegFile/FrameStrobe[18] Tile_X4Y10_RegFile/FrameStrobe[19]
+ Tile_X4Y10_RegFile/FrameStrobe[1] Tile_X4Y10_RegFile/FrameStrobe[2] Tile_X4Y10_RegFile/FrameStrobe[3]
+ Tile_X4Y10_RegFile/FrameStrobe[4] Tile_X4Y10_RegFile/FrameStrobe[5] Tile_X4Y10_RegFile/FrameStrobe[6]
+ Tile_X4Y10_RegFile/FrameStrobe[7] Tile_X4Y10_RegFile/FrameStrobe[8] Tile_X4Y10_RegFile/FrameStrobe[9]
+ Tile_X4Y9_RegFile/FrameStrobe[0] Tile_X4Y9_RegFile/FrameStrobe[10] Tile_X4Y9_RegFile/FrameStrobe[11]
+ Tile_X4Y9_RegFile/FrameStrobe[12] Tile_X4Y9_RegFile/FrameStrobe[13] Tile_X4Y9_RegFile/FrameStrobe[14]
+ Tile_X4Y9_RegFile/FrameStrobe[15] Tile_X4Y9_RegFile/FrameStrobe[16] Tile_X4Y9_RegFile/FrameStrobe[17]
+ Tile_X4Y9_RegFile/FrameStrobe[18] Tile_X4Y9_RegFile/FrameStrobe[19] Tile_X4Y9_RegFile/FrameStrobe[1]
+ Tile_X4Y9_RegFile/FrameStrobe[2] Tile_X4Y9_RegFile/FrameStrobe[3] Tile_X4Y9_RegFile/FrameStrobe[4]
+ Tile_X4Y9_RegFile/FrameStrobe[5] Tile_X4Y9_RegFile/FrameStrobe[6] Tile_X4Y9_RegFile/FrameStrobe[7]
+ Tile_X4Y9_RegFile/FrameStrobe[8] Tile_X4Y9_RegFile/FrameStrobe[9] Tile_X4Y9_RegFile/N1END[0]
+ Tile_X4Y9_RegFile/N1END[1] Tile_X4Y9_RegFile/N1END[2] Tile_X4Y9_RegFile/N1END[3]
+ Tile_X4Y11_RegFile/N1BEG[0] Tile_X4Y11_RegFile/N1BEG[1] Tile_X4Y11_RegFile/N1BEG[2]
+ Tile_X4Y11_RegFile/N1BEG[3] Tile_X4Y9_RegFile/N2MID[0] Tile_X4Y9_RegFile/N2MID[1]
+ Tile_X4Y9_RegFile/N2MID[2] Tile_X4Y9_RegFile/N2MID[3] Tile_X4Y9_RegFile/N2MID[4]
+ Tile_X4Y9_RegFile/N2MID[5] Tile_X4Y9_RegFile/N2MID[6] Tile_X4Y9_RegFile/N2MID[7]
+ Tile_X4Y9_RegFile/N2END[0] Tile_X4Y9_RegFile/N2END[1] Tile_X4Y9_RegFile/N2END[2]
+ Tile_X4Y9_RegFile/N2END[3] Tile_X4Y9_RegFile/N2END[4] Tile_X4Y9_RegFile/N2END[5]
+ Tile_X4Y9_RegFile/N2END[6] Tile_X4Y9_RegFile/N2END[7] Tile_X4Y10_RegFile/N2END[0]
+ Tile_X4Y10_RegFile/N2END[1] Tile_X4Y10_RegFile/N2END[2] Tile_X4Y10_RegFile/N2END[3]
+ Tile_X4Y10_RegFile/N2END[4] Tile_X4Y10_RegFile/N2END[5] Tile_X4Y10_RegFile/N2END[6]
+ Tile_X4Y10_RegFile/N2END[7] Tile_X4Y11_RegFile/N2BEG[0] Tile_X4Y11_RegFile/N2BEG[1]
+ Tile_X4Y11_RegFile/N2BEG[2] Tile_X4Y11_RegFile/N2BEG[3] Tile_X4Y11_RegFile/N2BEG[4]
+ Tile_X4Y11_RegFile/N2BEG[5] Tile_X4Y11_RegFile/N2BEG[6] Tile_X4Y11_RegFile/N2BEG[7]
+ Tile_X4Y9_RegFile/N4END[0] Tile_X4Y9_RegFile/N4END[10] Tile_X4Y9_RegFile/N4END[11]
+ Tile_X4Y9_RegFile/N4END[12] Tile_X4Y9_RegFile/N4END[13] Tile_X4Y9_RegFile/N4END[14]
+ Tile_X4Y9_RegFile/N4END[15] Tile_X4Y9_RegFile/N4END[1] Tile_X4Y9_RegFile/N4END[2]
+ Tile_X4Y9_RegFile/N4END[3] Tile_X4Y9_RegFile/N4END[4] Tile_X4Y9_RegFile/N4END[5]
+ Tile_X4Y9_RegFile/N4END[6] Tile_X4Y9_RegFile/N4END[7] Tile_X4Y9_RegFile/N4END[8]
+ Tile_X4Y9_RegFile/N4END[9] Tile_X4Y11_RegFile/N4BEG[0] Tile_X4Y11_RegFile/N4BEG[10]
+ Tile_X4Y11_RegFile/N4BEG[11] Tile_X4Y11_RegFile/N4BEG[12] Tile_X4Y11_RegFile/N4BEG[13]
+ Tile_X4Y11_RegFile/N4BEG[14] Tile_X4Y11_RegFile/N4BEG[15] Tile_X4Y11_RegFile/N4BEG[1]
+ Tile_X4Y11_RegFile/N4BEG[2] Tile_X4Y11_RegFile/N4BEG[3] Tile_X4Y11_RegFile/N4BEG[4]
+ Tile_X4Y11_RegFile/N4BEG[5] Tile_X4Y11_RegFile/N4BEG[6] Tile_X4Y11_RegFile/N4BEG[7]
+ Tile_X4Y11_RegFile/N4BEG[8] Tile_X4Y11_RegFile/N4BEG[9] Tile_X4Y9_RegFile/NN4END[0]
+ Tile_X4Y9_RegFile/NN4END[10] Tile_X4Y9_RegFile/NN4END[11] Tile_X4Y9_RegFile/NN4END[12]
+ Tile_X4Y9_RegFile/NN4END[13] Tile_X4Y9_RegFile/NN4END[14] Tile_X4Y9_RegFile/NN4END[15]
+ Tile_X4Y9_RegFile/NN4END[1] Tile_X4Y9_RegFile/NN4END[2] Tile_X4Y9_RegFile/NN4END[3]
+ Tile_X4Y9_RegFile/NN4END[4] Tile_X4Y9_RegFile/NN4END[5] Tile_X4Y9_RegFile/NN4END[6]
+ Tile_X4Y9_RegFile/NN4END[7] Tile_X4Y9_RegFile/NN4END[8] Tile_X4Y9_RegFile/NN4END[9]
+ Tile_X4Y11_RegFile/NN4BEG[0] Tile_X4Y11_RegFile/NN4BEG[10] Tile_X4Y11_RegFile/NN4BEG[11]
+ Tile_X4Y11_RegFile/NN4BEG[12] Tile_X4Y11_RegFile/NN4BEG[13] Tile_X4Y11_RegFile/NN4BEG[14]
+ Tile_X4Y11_RegFile/NN4BEG[15] Tile_X4Y11_RegFile/NN4BEG[1] Tile_X4Y11_RegFile/NN4BEG[2]
+ Tile_X4Y11_RegFile/NN4BEG[3] Tile_X4Y11_RegFile/NN4BEG[4] Tile_X4Y11_RegFile/NN4BEG[5]
+ Tile_X4Y11_RegFile/NN4BEG[6] Tile_X4Y11_RegFile/NN4BEG[7] Tile_X4Y11_RegFile/NN4BEG[8]
+ Tile_X4Y11_RegFile/NN4BEG[9] Tile_X4Y11_RegFile/S1END[0] Tile_X4Y11_RegFile/S1END[1]
+ Tile_X4Y11_RegFile/S1END[2] Tile_X4Y11_RegFile/S1END[3] Tile_X4Y9_RegFile/S1BEG[0]
+ Tile_X4Y9_RegFile/S1BEG[1] Tile_X4Y9_RegFile/S1BEG[2] Tile_X4Y9_RegFile/S1BEG[3]
+ Tile_X4Y11_RegFile/S2MID[0] Tile_X4Y11_RegFile/S2MID[1] Tile_X4Y11_RegFile/S2MID[2]
+ Tile_X4Y11_RegFile/S2MID[3] Tile_X4Y11_RegFile/S2MID[4] Tile_X4Y11_RegFile/S2MID[5]
+ Tile_X4Y11_RegFile/S2MID[6] Tile_X4Y11_RegFile/S2MID[7] Tile_X4Y11_RegFile/S2END[0]
+ Tile_X4Y11_RegFile/S2END[1] Tile_X4Y11_RegFile/S2END[2] Tile_X4Y11_RegFile/S2END[3]
+ Tile_X4Y11_RegFile/S2END[4] Tile_X4Y11_RegFile/S2END[5] Tile_X4Y11_RegFile/S2END[6]
+ Tile_X4Y11_RegFile/S2END[7] Tile_X4Y9_RegFile/S2BEGb[0] Tile_X4Y9_RegFile/S2BEGb[1]
+ Tile_X4Y9_RegFile/S2BEGb[2] Tile_X4Y9_RegFile/S2BEGb[3] Tile_X4Y9_RegFile/S2BEGb[4]
+ Tile_X4Y9_RegFile/S2BEGb[5] Tile_X4Y9_RegFile/S2BEGb[6] Tile_X4Y9_RegFile/S2BEGb[7]
+ Tile_X4Y9_RegFile/S2BEG[0] Tile_X4Y9_RegFile/S2BEG[1] Tile_X4Y9_RegFile/S2BEG[2]
+ Tile_X4Y9_RegFile/S2BEG[3] Tile_X4Y9_RegFile/S2BEG[4] Tile_X4Y9_RegFile/S2BEG[5]
+ Tile_X4Y9_RegFile/S2BEG[6] Tile_X4Y9_RegFile/S2BEG[7] Tile_X4Y11_RegFile/S4END[0]
+ Tile_X4Y11_RegFile/S4END[10] Tile_X4Y11_RegFile/S4END[11] Tile_X4Y11_RegFile/S4END[12]
+ Tile_X4Y11_RegFile/S4END[13] Tile_X4Y11_RegFile/S4END[14] Tile_X4Y11_RegFile/S4END[15]
+ Tile_X4Y11_RegFile/S4END[1] Tile_X4Y11_RegFile/S4END[2] Tile_X4Y11_RegFile/S4END[3]
+ Tile_X4Y11_RegFile/S4END[4] Tile_X4Y11_RegFile/S4END[5] Tile_X4Y11_RegFile/S4END[6]
+ Tile_X4Y11_RegFile/S4END[7] Tile_X4Y11_RegFile/S4END[8] Tile_X4Y11_RegFile/S4END[9]
+ Tile_X4Y9_RegFile/S4BEG[0] Tile_X4Y9_RegFile/S4BEG[10] Tile_X4Y9_RegFile/S4BEG[11]
+ Tile_X4Y9_RegFile/S4BEG[12] Tile_X4Y9_RegFile/S4BEG[13] Tile_X4Y9_RegFile/S4BEG[14]
+ Tile_X4Y9_RegFile/S4BEG[15] Tile_X4Y9_RegFile/S4BEG[1] Tile_X4Y9_RegFile/S4BEG[2]
+ Tile_X4Y9_RegFile/S4BEG[3] Tile_X4Y9_RegFile/S4BEG[4] Tile_X4Y9_RegFile/S4BEG[5]
+ Tile_X4Y9_RegFile/S4BEG[6] Tile_X4Y9_RegFile/S4BEG[7] Tile_X4Y9_RegFile/S4BEG[8]
+ Tile_X4Y9_RegFile/S4BEG[9] Tile_X4Y11_RegFile/SS4END[0] Tile_X4Y11_RegFile/SS4END[10]
+ Tile_X4Y11_RegFile/SS4END[11] Tile_X4Y11_RegFile/SS4END[12] Tile_X4Y11_RegFile/SS4END[13]
+ Tile_X4Y11_RegFile/SS4END[14] Tile_X4Y11_RegFile/SS4END[15] Tile_X4Y11_RegFile/SS4END[1]
+ Tile_X4Y11_RegFile/SS4END[2] Tile_X4Y11_RegFile/SS4END[3] Tile_X4Y11_RegFile/SS4END[4]
+ Tile_X4Y11_RegFile/SS4END[5] Tile_X4Y11_RegFile/SS4END[6] Tile_X4Y11_RegFile/SS4END[7]
+ Tile_X4Y11_RegFile/SS4END[8] Tile_X4Y11_RegFile/SS4END[9] Tile_X4Y9_RegFile/SS4BEG[0]
+ Tile_X4Y9_RegFile/SS4BEG[10] Tile_X4Y9_RegFile/SS4BEG[11] Tile_X4Y9_RegFile/SS4BEG[12]
+ Tile_X4Y9_RegFile/SS4BEG[13] Tile_X4Y9_RegFile/SS4BEG[14] Tile_X4Y9_RegFile/SS4BEG[15]
+ Tile_X4Y9_RegFile/SS4BEG[1] Tile_X4Y9_RegFile/SS4BEG[2] Tile_X4Y9_RegFile/SS4BEG[3]
+ Tile_X4Y9_RegFile/SS4BEG[4] Tile_X4Y9_RegFile/SS4BEG[5] Tile_X4Y9_RegFile/SS4BEG[6]
+ Tile_X4Y9_RegFile/SS4BEG[7] Tile_X4Y9_RegFile/SS4BEG[8] Tile_X4Y9_RegFile/SS4BEG[9]
+ Tile_X4Y10_RegFile/UserCLK Tile_X4Y9_RegFile/UserCLK VGND VPWR Tile_X3Y10_LUT4AB/W1END[0]
+ Tile_X3Y10_LUT4AB/W1END[1] Tile_X3Y10_LUT4AB/W1END[2] Tile_X3Y10_LUT4AB/W1END[3]
+ Tile_X5Y10_LUT4AB/W1BEG[0] Tile_X5Y10_LUT4AB/W1BEG[1] Tile_X5Y10_LUT4AB/W1BEG[2]
+ Tile_X5Y10_LUT4AB/W1BEG[3] Tile_X3Y10_LUT4AB/W2MID[0] Tile_X3Y10_LUT4AB/W2MID[1]
+ Tile_X3Y10_LUT4AB/W2MID[2] Tile_X3Y10_LUT4AB/W2MID[3] Tile_X3Y10_LUT4AB/W2MID[4]
+ Tile_X3Y10_LUT4AB/W2MID[5] Tile_X3Y10_LUT4AB/W2MID[6] Tile_X3Y10_LUT4AB/W2MID[7]
+ Tile_X3Y10_LUT4AB/W2END[0] Tile_X3Y10_LUT4AB/W2END[1] Tile_X3Y10_LUT4AB/W2END[2]
+ Tile_X3Y10_LUT4AB/W2END[3] Tile_X3Y10_LUT4AB/W2END[4] Tile_X3Y10_LUT4AB/W2END[5]
+ Tile_X3Y10_LUT4AB/W2END[6] Tile_X3Y10_LUT4AB/W2END[7] Tile_X5Y10_LUT4AB/W2BEGb[0]
+ Tile_X5Y10_LUT4AB/W2BEGb[1] Tile_X5Y10_LUT4AB/W2BEGb[2] Tile_X5Y10_LUT4AB/W2BEGb[3]
+ Tile_X5Y10_LUT4AB/W2BEGb[4] Tile_X5Y10_LUT4AB/W2BEGb[5] Tile_X5Y10_LUT4AB/W2BEGb[6]
+ Tile_X5Y10_LUT4AB/W2BEGb[7] Tile_X5Y10_LUT4AB/W2BEG[0] Tile_X5Y10_LUT4AB/W2BEG[1]
+ Tile_X5Y10_LUT4AB/W2BEG[2] Tile_X5Y10_LUT4AB/W2BEG[3] Tile_X5Y10_LUT4AB/W2BEG[4]
+ Tile_X5Y10_LUT4AB/W2BEG[5] Tile_X5Y10_LUT4AB/W2BEG[6] Tile_X5Y10_LUT4AB/W2BEG[7]
+ Tile_X3Y10_LUT4AB/W6END[0] Tile_X3Y10_LUT4AB/W6END[10] Tile_X3Y10_LUT4AB/W6END[11]
+ Tile_X3Y10_LUT4AB/W6END[1] Tile_X3Y10_LUT4AB/W6END[2] Tile_X3Y10_LUT4AB/W6END[3]
+ Tile_X3Y10_LUT4AB/W6END[4] Tile_X3Y10_LUT4AB/W6END[5] Tile_X3Y10_LUT4AB/W6END[6]
+ Tile_X3Y10_LUT4AB/W6END[7] Tile_X3Y10_LUT4AB/W6END[8] Tile_X3Y10_LUT4AB/W6END[9]
+ Tile_X5Y10_LUT4AB/W6BEG[0] Tile_X5Y10_LUT4AB/W6BEG[10] Tile_X5Y10_LUT4AB/W6BEG[11]
+ Tile_X5Y10_LUT4AB/W6BEG[1] Tile_X5Y10_LUT4AB/W6BEG[2] Tile_X5Y10_LUT4AB/W6BEG[3]
+ Tile_X5Y10_LUT4AB/W6BEG[4] Tile_X5Y10_LUT4AB/W6BEG[5] Tile_X5Y10_LUT4AB/W6BEG[6]
+ Tile_X5Y10_LUT4AB/W6BEG[7] Tile_X5Y10_LUT4AB/W6BEG[8] Tile_X5Y10_LUT4AB/W6BEG[9]
+ Tile_X3Y10_LUT4AB/WW4END[0] Tile_X3Y10_LUT4AB/WW4END[10] Tile_X3Y10_LUT4AB/WW4END[11]
+ Tile_X3Y10_LUT4AB/WW4END[12] Tile_X3Y10_LUT4AB/WW4END[13] Tile_X3Y10_LUT4AB/WW4END[14]
+ Tile_X3Y10_LUT4AB/WW4END[15] Tile_X3Y10_LUT4AB/WW4END[1] Tile_X3Y10_LUT4AB/WW4END[2]
+ Tile_X3Y10_LUT4AB/WW4END[3] Tile_X3Y10_LUT4AB/WW4END[4] Tile_X3Y10_LUT4AB/WW4END[5]
+ Tile_X3Y10_LUT4AB/WW4END[6] Tile_X3Y10_LUT4AB/WW4END[7] Tile_X3Y10_LUT4AB/WW4END[8]
+ Tile_X3Y10_LUT4AB/WW4END[9] Tile_X5Y10_LUT4AB/WW4BEG[0] Tile_X5Y10_LUT4AB/WW4BEG[10]
+ Tile_X5Y10_LUT4AB/WW4BEG[11] Tile_X5Y10_LUT4AB/WW4BEG[12] Tile_X5Y10_LUT4AB/WW4BEG[13]
+ Tile_X5Y10_LUT4AB/WW4BEG[14] Tile_X5Y10_LUT4AB/WW4BEG[15] Tile_X5Y10_LUT4AB/WW4BEG[1]
+ Tile_X5Y10_LUT4AB/WW4BEG[2] Tile_X5Y10_LUT4AB/WW4BEG[3] Tile_X5Y10_LUT4AB/WW4BEG[4]
+ Tile_X5Y10_LUT4AB/WW4BEG[5] Tile_X5Y10_LUT4AB/WW4BEG[6] Tile_X5Y10_LUT4AB/WW4BEG[7]
+ Tile_X5Y10_LUT4AB/WW4BEG[8] Tile_X5Y10_LUT4AB/WW4BEG[9] RegFile
XTile_X8Y9_LUT4AB Tile_X8Y9_LUT4AB/Ci Tile_X8Y9_LUT4AB/Co Tile_X9Y9_LUT4AB/E1END[0]
+ Tile_X9Y9_LUT4AB/E1END[1] Tile_X9Y9_LUT4AB/E1END[2] Tile_X9Y9_LUT4AB/E1END[3] Tile_X8Y9_LUT4AB/E1END[0]
+ Tile_X8Y9_LUT4AB/E1END[1] Tile_X8Y9_LUT4AB/E1END[2] Tile_X8Y9_LUT4AB/E1END[3] Tile_X9Y9_LUT4AB/E2MID[0]
+ Tile_X9Y9_LUT4AB/E2MID[1] Tile_X9Y9_LUT4AB/E2MID[2] Tile_X9Y9_LUT4AB/E2MID[3] Tile_X9Y9_LUT4AB/E2MID[4]
+ Tile_X9Y9_LUT4AB/E2MID[5] Tile_X9Y9_LUT4AB/E2MID[6] Tile_X9Y9_LUT4AB/E2MID[7] Tile_X9Y9_LUT4AB/E2END[0]
+ Tile_X9Y9_LUT4AB/E2END[1] Tile_X9Y9_LUT4AB/E2END[2] Tile_X9Y9_LUT4AB/E2END[3] Tile_X9Y9_LUT4AB/E2END[4]
+ Tile_X9Y9_LUT4AB/E2END[5] Tile_X9Y9_LUT4AB/E2END[6] Tile_X9Y9_LUT4AB/E2END[7] Tile_X8Y9_LUT4AB/E2END[0]
+ Tile_X8Y9_LUT4AB/E2END[1] Tile_X8Y9_LUT4AB/E2END[2] Tile_X8Y9_LUT4AB/E2END[3] Tile_X8Y9_LUT4AB/E2END[4]
+ Tile_X8Y9_LUT4AB/E2END[5] Tile_X8Y9_LUT4AB/E2END[6] Tile_X8Y9_LUT4AB/E2END[7] Tile_X8Y9_LUT4AB/E2MID[0]
+ Tile_X8Y9_LUT4AB/E2MID[1] Tile_X8Y9_LUT4AB/E2MID[2] Tile_X8Y9_LUT4AB/E2MID[3] Tile_X8Y9_LUT4AB/E2MID[4]
+ Tile_X8Y9_LUT4AB/E2MID[5] Tile_X8Y9_LUT4AB/E2MID[6] Tile_X8Y9_LUT4AB/E2MID[7] Tile_X9Y9_LUT4AB/E6END[0]
+ Tile_X9Y9_LUT4AB/E6END[10] Tile_X9Y9_LUT4AB/E6END[11] Tile_X9Y9_LUT4AB/E6END[1]
+ Tile_X9Y9_LUT4AB/E6END[2] Tile_X9Y9_LUT4AB/E6END[3] Tile_X9Y9_LUT4AB/E6END[4] Tile_X9Y9_LUT4AB/E6END[5]
+ Tile_X9Y9_LUT4AB/E6END[6] Tile_X9Y9_LUT4AB/E6END[7] Tile_X9Y9_LUT4AB/E6END[8] Tile_X9Y9_LUT4AB/E6END[9]
+ Tile_X8Y9_LUT4AB/E6END[0] Tile_X8Y9_LUT4AB/E6END[10] Tile_X8Y9_LUT4AB/E6END[11]
+ Tile_X8Y9_LUT4AB/E6END[1] Tile_X8Y9_LUT4AB/E6END[2] Tile_X8Y9_LUT4AB/E6END[3] Tile_X8Y9_LUT4AB/E6END[4]
+ Tile_X8Y9_LUT4AB/E6END[5] Tile_X8Y9_LUT4AB/E6END[6] Tile_X8Y9_LUT4AB/E6END[7] Tile_X8Y9_LUT4AB/E6END[8]
+ Tile_X8Y9_LUT4AB/E6END[9] Tile_X9Y9_LUT4AB/EE4END[0] Tile_X9Y9_LUT4AB/EE4END[10]
+ Tile_X9Y9_LUT4AB/EE4END[11] Tile_X9Y9_LUT4AB/EE4END[12] Tile_X9Y9_LUT4AB/EE4END[13]
+ Tile_X9Y9_LUT4AB/EE4END[14] Tile_X9Y9_LUT4AB/EE4END[15] Tile_X9Y9_LUT4AB/EE4END[1]
+ Tile_X9Y9_LUT4AB/EE4END[2] Tile_X9Y9_LUT4AB/EE4END[3] Tile_X9Y9_LUT4AB/EE4END[4]
+ Tile_X9Y9_LUT4AB/EE4END[5] Tile_X9Y9_LUT4AB/EE4END[6] Tile_X9Y9_LUT4AB/EE4END[7]
+ Tile_X9Y9_LUT4AB/EE4END[8] Tile_X9Y9_LUT4AB/EE4END[9] Tile_X8Y9_LUT4AB/EE4END[0]
+ Tile_X8Y9_LUT4AB/EE4END[10] Tile_X8Y9_LUT4AB/EE4END[11] Tile_X8Y9_LUT4AB/EE4END[12]
+ Tile_X8Y9_LUT4AB/EE4END[13] Tile_X8Y9_LUT4AB/EE4END[14] Tile_X8Y9_LUT4AB/EE4END[15]
+ Tile_X8Y9_LUT4AB/EE4END[1] Tile_X8Y9_LUT4AB/EE4END[2] Tile_X8Y9_LUT4AB/EE4END[3]
+ Tile_X8Y9_LUT4AB/EE4END[4] Tile_X8Y9_LUT4AB/EE4END[5] Tile_X8Y9_LUT4AB/EE4END[6]
+ Tile_X8Y9_LUT4AB/EE4END[7] Tile_X8Y9_LUT4AB/EE4END[8] Tile_X8Y9_LUT4AB/EE4END[9]
+ Tile_X8Y9_LUT4AB/FrameData[0] Tile_X8Y9_LUT4AB/FrameData[10] Tile_X8Y9_LUT4AB/FrameData[11]
+ Tile_X8Y9_LUT4AB/FrameData[12] Tile_X8Y9_LUT4AB/FrameData[13] Tile_X8Y9_LUT4AB/FrameData[14]
+ Tile_X8Y9_LUT4AB/FrameData[15] Tile_X8Y9_LUT4AB/FrameData[16] Tile_X8Y9_LUT4AB/FrameData[17]
+ Tile_X8Y9_LUT4AB/FrameData[18] Tile_X8Y9_LUT4AB/FrameData[19] Tile_X8Y9_LUT4AB/FrameData[1]
+ Tile_X8Y9_LUT4AB/FrameData[20] Tile_X8Y9_LUT4AB/FrameData[21] Tile_X8Y9_LUT4AB/FrameData[22]
+ Tile_X8Y9_LUT4AB/FrameData[23] Tile_X8Y9_LUT4AB/FrameData[24] Tile_X8Y9_LUT4AB/FrameData[25]
+ Tile_X8Y9_LUT4AB/FrameData[26] Tile_X8Y9_LUT4AB/FrameData[27] Tile_X8Y9_LUT4AB/FrameData[28]
+ Tile_X8Y9_LUT4AB/FrameData[29] Tile_X8Y9_LUT4AB/FrameData[2] Tile_X8Y9_LUT4AB/FrameData[30]
+ Tile_X8Y9_LUT4AB/FrameData[31] Tile_X8Y9_LUT4AB/FrameData[3] Tile_X8Y9_LUT4AB/FrameData[4]
+ Tile_X8Y9_LUT4AB/FrameData[5] Tile_X8Y9_LUT4AB/FrameData[6] Tile_X8Y9_LUT4AB/FrameData[7]
+ Tile_X8Y9_LUT4AB/FrameData[8] Tile_X8Y9_LUT4AB/FrameData[9] Tile_X9Y9_LUT4AB/FrameData[0]
+ Tile_X9Y9_LUT4AB/FrameData[10] Tile_X9Y9_LUT4AB/FrameData[11] Tile_X9Y9_LUT4AB/FrameData[12]
+ Tile_X9Y9_LUT4AB/FrameData[13] Tile_X9Y9_LUT4AB/FrameData[14] Tile_X9Y9_LUT4AB/FrameData[15]
+ Tile_X9Y9_LUT4AB/FrameData[16] Tile_X9Y9_LUT4AB/FrameData[17] Tile_X9Y9_LUT4AB/FrameData[18]
+ Tile_X9Y9_LUT4AB/FrameData[19] Tile_X9Y9_LUT4AB/FrameData[1] Tile_X9Y9_LUT4AB/FrameData[20]
+ Tile_X9Y9_LUT4AB/FrameData[21] Tile_X9Y9_LUT4AB/FrameData[22] Tile_X9Y9_LUT4AB/FrameData[23]
+ Tile_X9Y9_LUT4AB/FrameData[24] Tile_X9Y9_LUT4AB/FrameData[25] Tile_X9Y9_LUT4AB/FrameData[26]
+ Tile_X9Y9_LUT4AB/FrameData[27] Tile_X9Y9_LUT4AB/FrameData[28] Tile_X9Y9_LUT4AB/FrameData[29]
+ Tile_X9Y9_LUT4AB/FrameData[2] Tile_X9Y9_LUT4AB/FrameData[30] Tile_X9Y9_LUT4AB/FrameData[31]
+ Tile_X9Y9_LUT4AB/FrameData[3] Tile_X9Y9_LUT4AB/FrameData[4] Tile_X9Y9_LUT4AB/FrameData[5]
+ Tile_X9Y9_LUT4AB/FrameData[6] Tile_X9Y9_LUT4AB/FrameData[7] Tile_X9Y9_LUT4AB/FrameData[8]
+ Tile_X9Y9_LUT4AB/FrameData[9] Tile_X8Y9_LUT4AB/FrameStrobe[0] Tile_X8Y9_LUT4AB/FrameStrobe[10]
+ Tile_X8Y9_LUT4AB/FrameStrobe[11] Tile_X8Y9_LUT4AB/FrameStrobe[12] Tile_X8Y9_LUT4AB/FrameStrobe[13]
+ Tile_X8Y9_LUT4AB/FrameStrobe[14] Tile_X8Y9_LUT4AB/FrameStrobe[15] Tile_X8Y9_LUT4AB/FrameStrobe[16]
+ Tile_X8Y9_LUT4AB/FrameStrobe[17] Tile_X8Y9_LUT4AB/FrameStrobe[18] Tile_X8Y9_LUT4AB/FrameStrobe[19]
+ Tile_X8Y9_LUT4AB/FrameStrobe[1] Tile_X8Y9_LUT4AB/FrameStrobe[2] Tile_X8Y9_LUT4AB/FrameStrobe[3]
+ Tile_X8Y9_LUT4AB/FrameStrobe[4] Tile_X8Y9_LUT4AB/FrameStrobe[5] Tile_X8Y9_LUT4AB/FrameStrobe[6]
+ Tile_X8Y9_LUT4AB/FrameStrobe[7] Tile_X8Y9_LUT4AB/FrameStrobe[8] Tile_X8Y9_LUT4AB/FrameStrobe[9]
+ Tile_X8Y8_LUT4AB/FrameStrobe[0] Tile_X8Y8_LUT4AB/FrameStrobe[10] Tile_X8Y8_LUT4AB/FrameStrobe[11]
+ Tile_X8Y8_LUT4AB/FrameStrobe[12] Tile_X8Y8_LUT4AB/FrameStrobe[13] Tile_X8Y8_LUT4AB/FrameStrobe[14]
+ Tile_X8Y8_LUT4AB/FrameStrobe[15] Tile_X8Y8_LUT4AB/FrameStrobe[16] Tile_X8Y8_LUT4AB/FrameStrobe[17]
+ Tile_X8Y8_LUT4AB/FrameStrobe[18] Tile_X8Y8_LUT4AB/FrameStrobe[19] Tile_X8Y8_LUT4AB/FrameStrobe[1]
+ Tile_X8Y8_LUT4AB/FrameStrobe[2] Tile_X8Y8_LUT4AB/FrameStrobe[3] Tile_X8Y8_LUT4AB/FrameStrobe[4]
+ Tile_X8Y8_LUT4AB/FrameStrobe[5] Tile_X8Y8_LUT4AB/FrameStrobe[6] Tile_X8Y8_LUT4AB/FrameStrobe[7]
+ Tile_X8Y8_LUT4AB/FrameStrobe[8] Tile_X8Y8_LUT4AB/FrameStrobe[9] Tile_X8Y9_LUT4AB/N1BEG[0]
+ Tile_X8Y9_LUT4AB/N1BEG[1] Tile_X8Y9_LUT4AB/N1BEG[2] Tile_X8Y9_LUT4AB/N1BEG[3] Tile_X8Y9_LUT4AB/N1END[0]
+ Tile_X8Y9_LUT4AB/N1END[1] Tile_X8Y9_LUT4AB/N1END[2] Tile_X8Y9_LUT4AB/N1END[3] Tile_X8Y9_LUT4AB/N2BEG[0]
+ Tile_X8Y9_LUT4AB/N2BEG[1] Tile_X8Y9_LUT4AB/N2BEG[2] Tile_X8Y9_LUT4AB/N2BEG[3] Tile_X8Y9_LUT4AB/N2BEG[4]
+ Tile_X8Y9_LUT4AB/N2BEG[5] Tile_X8Y9_LUT4AB/N2BEG[6] Tile_X8Y9_LUT4AB/N2BEG[7] Tile_X8Y8_LUT4AB/N2END[0]
+ Tile_X8Y8_LUT4AB/N2END[1] Tile_X8Y8_LUT4AB/N2END[2] Tile_X8Y8_LUT4AB/N2END[3] Tile_X8Y8_LUT4AB/N2END[4]
+ Tile_X8Y8_LUT4AB/N2END[5] Tile_X8Y8_LUT4AB/N2END[6] Tile_X8Y8_LUT4AB/N2END[7] Tile_X8Y9_LUT4AB/N2END[0]
+ Tile_X8Y9_LUT4AB/N2END[1] Tile_X8Y9_LUT4AB/N2END[2] Tile_X8Y9_LUT4AB/N2END[3] Tile_X8Y9_LUT4AB/N2END[4]
+ Tile_X8Y9_LUT4AB/N2END[5] Tile_X8Y9_LUT4AB/N2END[6] Tile_X8Y9_LUT4AB/N2END[7] Tile_X8Y9_LUT4AB/N2MID[0]
+ Tile_X8Y9_LUT4AB/N2MID[1] Tile_X8Y9_LUT4AB/N2MID[2] Tile_X8Y9_LUT4AB/N2MID[3] Tile_X8Y9_LUT4AB/N2MID[4]
+ Tile_X8Y9_LUT4AB/N2MID[5] Tile_X8Y9_LUT4AB/N2MID[6] Tile_X8Y9_LUT4AB/N2MID[7] Tile_X8Y9_LUT4AB/N4BEG[0]
+ Tile_X8Y9_LUT4AB/N4BEG[10] Tile_X8Y9_LUT4AB/N4BEG[11] Tile_X8Y9_LUT4AB/N4BEG[12]
+ Tile_X8Y9_LUT4AB/N4BEG[13] Tile_X8Y9_LUT4AB/N4BEG[14] Tile_X8Y9_LUT4AB/N4BEG[15]
+ Tile_X8Y9_LUT4AB/N4BEG[1] Tile_X8Y9_LUT4AB/N4BEG[2] Tile_X8Y9_LUT4AB/N4BEG[3] Tile_X8Y9_LUT4AB/N4BEG[4]
+ Tile_X8Y9_LUT4AB/N4BEG[5] Tile_X8Y9_LUT4AB/N4BEG[6] Tile_X8Y9_LUT4AB/N4BEG[7] Tile_X8Y9_LUT4AB/N4BEG[8]
+ Tile_X8Y9_LUT4AB/N4BEG[9] Tile_X8Y9_LUT4AB/N4END[0] Tile_X8Y9_LUT4AB/N4END[10] Tile_X8Y9_LUT4AB/N4END[11]
+ Tile_X8Y9_LUT4AB/N4END[12] Tile_X8Y9_LUT4AB/N4END[13] Tile_X8Y9_LUT4AB/N4END[14]
+ Tile_X8Y9_LUT4AB/N4END[15] Tile_X8Y9_LUT4AB/N4END[1] Tile_X8Y9_LUT4AB/N4END[2] Tile_X8Y9_LUT4AB/N4END[3]
+ Tile_X8Y9_LUT4AB/N4END[4] Tile_X8Y9_LUT4AB/N4END[5] Tile_X8Y9_LUT4AB/N4END[6] Tile_X8Y9_LUT4AB/N4END[7]
+ Tile_X8Y9_LUT4AB/N4END[8] Tile_X8Y9_LUT4AB/N4END[9] Tile_X8Y9_LUT4AB/NN4BEG[0] Tile_X8Y9_LUT4AB/NN4BEG[10]
+ Tile_X8Y9_LUT4AB/NN4BEG[11] Tile_X8Y9_LUT4AB/NN4BEG[12] Tile_X8Y9_LUT4AB/NN4BEG[13]
+ Tile_X8Y9_LUT4AB/NN4BEG[14] Tile_X8Y9_LUT4AB/NN4BEG[15] Tile_X8Y9_LUT4AB/NN4BEG[1]
+ Tile_X8Y9_LUT4AB/NN4BEG[2] Tile_X8Y9_LUT4AB/NN4BEG[3] Tile_X8Y9_LUT4AB/NN4BEG[4]
+ Tile_X8Y9_LUT4AB/NN4BEG[5] Tile_X8Y9_LUT4AB/NN4BEG[6] Tile_X8Y9_LUT4AB/NN4BEG[7]
+ Tile_X8Y9_LUT4AB/NN4BEG[8] Tile_X8Y9_LUT4AB/NN4BEG[9] Tile_X8Y9_LUT4AB/NN4END[0]
+ Tile_X8Y9_LUT4AB/NN4END[10] Tile_X8Y9_LUT4AB/NN4END[11] Tile_X8Y9_LUT4AB/NN4END[12]
+ Tile_X8Y9_LUT4AB/NN4END[13] Tile_X8Y9_LUT4AB/NN4END[14] Tile_X8Y9_LUT4AB/NN4END[15]
+ Tile_X8Y9_LUT4AB/NN4END[1] Tile_X8Y9_LUT4AB/NN4END[2] Tile_X8Y9_LUT4AB/NN4END[3]
+ Tile_X8Y9_LUT4AB/NN4END[4] Tile_X8Y9_LUT4AB/NN4END[5] Tile_X8Y9_LUT4AB/NN4END[6]
+ Tile_X8Y9_LUT4AB/NN4END[7] Tile_X8Y9_LUT4AB/NN4END[8] Tile_X8Y9_LUT4AB/NN4END[9]
+ Tile_X8Y9_LUT4AB/S1BEG[0] Tile_X8Y9_LUT4AB/S1BEG[1] Tile_X8Y9_LUT4AB/S1BEG[2] Tile_X8Y9_LUT4AB/S1BEG[3]
+ Tile_X8Y9_LUT4AB/S1END[0] Tile_X8Y9_LUT4AB/S1END[1] Tile_X8Y9_LUT4AB/S1END[2] Tile_X8Y9_LUT4AB/S1END[3]
+ Tile_X8Y9_LUT4AB/S2BEG[0] Tile_X8Y9_LUT4AB/S2BEG[1] Tile_X8Y9_LUT4AB/S2BEG[2] Tile_X8Y9_LUT4AB/S2BEG[3]
+ Tile_X8Y9_LUT4AB/S2BEG[4] Tile_X8Y9_LUT4AB/S2BEG[5] Tile_X8Y9_LUT4AB/S2BEG[6] Tile_X8Y9_LUT4AB/S2BEG[7]
+ Tile_X8Y9_LUT4AB/S2BEGb[0] Tile_X8Y9_LUT4AB/S2BEGb[1] Tile_X8Y9_LUT4AB/S2BEGb[2]
+ Tile_X8Y9_LUT4AB/S2BEGb[3] Tile_X8Y9_LUT4AB/S2BEGb[4] Tile_X8Y9_LUT4AB/S2BEGb[5]
+ Tile_X8Y9_LUT4AB/S2BEGb[6] Tile_X8Y9_LUT4AB/S2BEGb[7] Tile_X8Y9_LUT4AB/S2END[0]
+ Tile_X8Y9_LUT4AB/S2END[1] Tile_X8Y9_LUT4AB/S2END[2] Tile_X8Y9_LUT4AB/S2END[3] Tile_X8Y9_LUT4AB/S2END[4]
+ Tile_X8Y9_LUT4AB/S2END[5] Tile_X8Y9_LUT4AB/S2END[6] Tile_X8Y9_LUT4AB/S2END[7] Tile_X8Y9_LUT4AB/S2MID[0]
+ Tile_X8Y9_LUT4AB/S2MID[1] Tile_X8Y9_LUT4AB/S2MID[2] Tile_X8Y9_LUT4AB/S2MID[3] Tile_X8Y9_LUT4AB/S2MID[4]
+ Tile_X8Y9_LUT4AB/S2MID[5] Tile_X8Y9_LUT4AB/S2MID[6] Tile_X8Y9_LUT4AB/S2MID[7] Tile_X8Y9_LUT4AB/S4BEG[0]
+ Tile_X8Y9_LUT4AB/S4BEG[10] Tile_X8Y9_LUT4AB/S4BEG[11] Tile_X8Y9_LUT4AB/S4BEG[12]
+ Tile_X8Y9_LUT4AB/S4BEG[13] Tile_X8Y9_LUT4AB/S4BEG[14] Tile_X8Y9_LUT4AB/S4BEG[15]
+ Tile_X8Y9_LUT4AB/S4BEG[1] Tile_X8Y9_LUT4AB/S4BEG[2] Tile_X8Y9_LUT4AB/S4BEG[3] Tile_X8Y9_LUT4AB/S4BEG[4]
+ Tile_X8Y9_LUT4AB/S4BEG[5] Tile_X8Y9_LUT4AB/S4BEG[6] Tile_X8Y9_LUT4AB/S4BEG[7] Tile_X8Y9_LUT4AB/S4BEG[8]
+ Tile_X8Y9_LUT4AB/S4BEG[9] Tile_X8Y9_LUT4AB/S4END[0] Tile_X8Y9_LUT4AB/S4END[10] Tile_X8Y9_LUT4AB/S4END[11]
+ Tile_X8Y9_LUT4AB/S4END[12] Tile_X8Y9_LUT4AB/S4END[13] Tile_X8Y9_LUT4AB/S4END[14]
+ Tile_X8Y9_LUT4AB/S4END[15] Tile_X8Y9_LUT4AB/S4END[1] Tile_X8Y9_LUT4AB/S4END[2] Tile_X8Y9_LUT4AB/S4END[3]
+ Tile_X8Y9_LUT4AB/S4END[4] Tile_X8Y9_LUT4AB/S4END[5] Tile_X8Y9_LUT4AB/S4END[6] Tile_X8Y9_LUT4AB/S4END[7]
+ Tile_X8Y9_LUT4AB/S4END[8] Tile_X8Y9_LUT4AB/S4END[9] Tile_X8Y9_LUT4AB/SS4BEG[0] Tile_X8Y9_LUT4AB/SS4BEG[10]
+ Tile_X8Y9_LUT4AB/SS4BEG[11] Tile_X8Y9_LUT4AB/SS4BEG[12] Tile_X8Y9_LUT4AB/SS4BEG[13]
+ Tile_X8Y9_LUT4AB/SS4BEG[14] Tile_X8Y9_LUT4AB/SS4BEG[15] Tile_X8Y9_LUT4AB/SS4BEG[1]
+ Tile_X8Y9_LUT4AB/SS4BEG[2] Tile_X8Y9_LUT4AB/SS4BEG[3] Tile_X8Y9_LUT4AB/SS4BEG[4]
+ Tile_X8Y9_LUT4AB/SS4BEG[5] Tile_X8Y9_LUT4AB/SS4BEG[6] Tile_X8Y9_LUT4AB/SS4BEG[7]
+ Tile_X8Y9_LUT4AB/SS4BEG[8] Tile_X8Y9_LUT4AB/SS4BEG[9] Tile_X8Y9_LUT4AB/SS4END[0]
+ Tile_X8Y9_LUT4AB/SS4END[10] Tile_X8Y9_LUT4AB/SS4END[11] Tile_X8Y9_LUT4AB/SS4END[12]
+ Tile_X8Y9_LUT4AB/SS4END[13] Tile_X8Y9_LUT4AB/SS4END[14] Tile_X8Y9_LUT4AB/SS4END[15]
+ Tile_X8Y9_LUT4AB/SS4END[1] Tile_X8Y9_LUT4AB/SS4END[2] Tile_X8Y9_LUT4AB/SS4END[3]
+ Tile_X8Y9_LUT4AB/SS4END[4] Tile_X8Y9_LUT4AB/SS4END[5] Tile_X8Y9_LUT4AB/SS4END[6]
+ Tile_X8Y9_LUT4AB/SS4END[7] Tile_X8Y9_LUT4AB/SS4END[8] Tile_X8Y9_LUT4AB/SS4END[9]
+ Tile_X8Y9_LUT4AB/UserCLK Tile_X8Y8_LUT4AB/UserCLK VGND VPWR Tile_X8Y9_LUT4AB/W1BEG[0]
+ Tile_X8Y9_LUT4AB/W1BEG[1] Tile_X8Y9_LUT4AB/W1BEG[2] Tile_X8Y9_LUT4AB/W1BEG[3] Tile_X9Y9_LUT4AB/W1BEG[0]
+ Tile_X9Y9_LUT4AB/W1BEG[1] Tile_X9Y9_LUT4AB/W1BEG[2] Tile_X9Y9_LUT4AB/W1BEG[3] Tile_X8Y9_LUT4AB/W2BEG[0]
+ Tile_X8Y9_LUT4AB/W2BEG[1] Tile_X8Y9_LUT4AB/W2BEG[2] Tile_X8Y9_LUT4AB/W2BEG[3] Tile_X8Y9_LUT4AB/W2BEG[4]
+ Tile_X8Y9_LUT4AB/W2BEG[5] Tile_X8Y9_LUT4AB/W2BEG[6] Tile_X8Y9_LUT4AB/W2BEG[7] Tile_X8Y9_LUT4AB/W2BEGb[0]
+ Tile_X8Y9_LUT4AB/W2BEGb[1] Tile_X8Y9_LUT4AB/W2BEGb[2] Tile_X8Y9_LUT4AB/W2BEGb[3]
+ Tile_X8Y9_LUT4AB/W2BEGb[4] Tile_X8Y9_LUT4AB/W2BEGb[5] Tile_X8Y9_LUT4AB/W2BEGb[6]
+ Tile_X8Y9_LUT4AB/W2BEGb[7] Tile_X8Y9_LUT4AB/W2END[0] Tile_X8Y9_LUT4AB/W2END[1] Tile_X8Y9_LUT4AB/W2END[2]
+ Tile_X8Y9_LUT4AB/W2END[3] Tile_X8Y9_LUT4AB/W2END[4] Tile_X8Y9_LUT4AB/W2END[5] Tile_X8Y9_LUT4AB/W2END[6]
+ Tile_X8Y9_LUT4AB/W2END[7] Tile_X9Y9_LUT4AB/W2BEG[0] Tile_X9Y9_LUT4AB/W2BEG[1] Tile_X9Y9_LUT4AB/W2BEG[2]
+ Tile_X9Y9_LUT4AB/W2BEG[3] Tile_X9Y9_LUT4AB/W2BEG[4] Tile_X9Y9_LUT4AB/W2BEG[5] Tile_X9Y9_LUT4AB/W2BEG[6]
+ Tile_X9Y9_LUT4AB/W2BEG[7] Tile_X8Y9_LUT4AB/W6BEG[0] Tile_X8Y9_LUT4AB/W6BEG[10] Tile_X8Y9_LUT4AB/W6BEG[11]
+ Tile_X8Y9_LUT4AB/W6BEG[1] Tile_X8Y9_LUT4AB/W6BEG[2] Tile_X8Y9_LUT4AB/W6BEG[3] Tile_X8Y9_LUT4AB/W6BEG[4]
+ Tile_X8Y9_LUT4AB/W6BEG[5] Tile_X8Y9_LUT4AB/W6BEG[6] Tile_X8Y9_LUT4AB/W6BEG[7] Tile_X8Y9_LUT4AB/W6BEG[8]
+ Tile_X8Y9_LUT4AB/W6BEG[9] Tile_X9Y9_LUT4AB/W6BEG[0] Tile_X9Y9_LUT4AB/W6BEG[10] Tile_X9Y9_LUT4AB/W6BEG[11]
+ Tile_X9Y9_LUT4AB/W6BEG[1] Tile_X9Y9_LUT4AB/W6BEG[2] Tile_X9Y9_LUT4AB/W6BEG[3] Tile_X9Y9_LUT4AB/W6BEG[4]
+ Tile_X9Y9_LUT4AB/W6BEG[5] Tile_X9Y9_LUT4AB/W6BEG[6] Tile_X9Y9_LUT4AB/W6BEG[7] Tile_X9Y9_LUT4AB/W6BEG[8]
+ Tile_X9Y9_LUT4AB/W6BEG[9] Tile_X8Y9_LUT4AB/WW4BEG[0] Tile_X8Y9_LUT4AB/WW4BEG[10]
+ Tile_X8Y9_LUT4AB/WW4BEG[11] Tile_X8Y9_LUT4AB/WW4BEG[12] Tile_X8Y9_LUT4AB/WW4BEG[13]
+ Tile_X8Y9_LUT4AB/WW4BEG[14] Tile_X8Y9_LUT4AB/WW4BEG[15] Tile_X8Y9_LUT4AB/WW4BEG[1]
+ Tile_X8Y9_LUT4AB/WW4BEG[2] Tile_X8Y9_LUT4AB/WW4BEG[3] Tile_X8Y9_LUT4AB/WW4BEG[4]
+ Tile_X8Y9_LUT4AB/WW4BEG[5] Tile_X8Y9_LUT4AB/WW4BEG[6] Tile_X8Y9_LUT4AB/WW4BEG[7]
+ Tile_X8Y9_LUT4AB/WW4BEG[8] Tile_X8Y9_LUT4AB/WW4BEG[9] Tile_X9Y9_LUT4AB/WW4BEG[0]
+ Tile_X9Y9_LUT4AB/WW4BEG[10] Tile_X9Y9_LUT4AB/WW4BEG[11] Tile_X9Y9_LUT4AB/WW4BEG[12]
+ Tile_X9Y9_LUT4AB/WW4BEG[13] Tile_X9Y9_LUT4AB/WW4BEG[14] Tile_X9Y9_LUT4AB/WW4BEG[15]
+ Tile_X9Y9_LUT4AB/WW4BEG[1] Tile_X9Y9_LUT4AB/WW4BEG[2] Tile_X9Y9_LUT4AB/WW4BEG[3]
+ Tile_X9Y9_LUT4AB/WW4BEG[4] Tile_X9Y9_LUT4AB/WW4BEG[5] Tile_X9Y9_LUT4AB/WW4BEG[6]
+ Tile_X9Y9_LUT4AB/WW4BEG[7] Tile_X9Y9_LUT4AB/WW4BEG[8] Tile_X9Y9_LUT4AB/WW4BEG[9]
+ LUT4AB
XTile_X0Y12_W_IO Tile_X0Y12_A_I_top Tile_X0Y12_A_O_top Tile_X0Y12_A_T_top Tile_X0Y12_A_config_C_bit0
+ Tile_X0Y12_A_config_C_bit1 Tile_X0Y12_A_config_C_bit2 Tile_X0Y12_A_config_C_bit3
+ Tile_X0Y12_B_I_top Tile_X0Y12_B_O_top Tile_X0Y12_B_T_top Tile_X0Y12_B_config_C_bit0
+ Tile_X0Y12_B_config_C_bit1 Tile_X0Y12_B_config_C_bit2 Tile_X0Y12_B_config_C_bit3
+ Tile_X0Y12_W_IO/E1BEG[0] Tile_X0Y12_W_IO/E1BEG[1] Tile_X0Y12_W_IO/E1BEG[2] Tile_X0Y12_W_IO/E1BEG[3]
+ Tile_X0Y12_W_IO/E2BEG[0] Tile_X0Y12_W_IO/E2BEG[1] Tile_X0Y12_W_IO/E2BEG[2] Tile_X0Y12_W_IO/E2BEG[3]
+ Tile_X0Y12_W_IO/E2BEG[4] Tile_X0Y12_W_IO/E2BEG[5] Tile_X0Y12_W_IO/E2BEG[6] Tile_X0Y12_W_IO/E2BEG[7]
+ Tile_X0Y12_W_IO/E2BEGb[0] Tile_X0Y12_W_IO/E2BEGb[1] Tile_X0Y12_W_IO/E2BEGb[2] Tile_X0Y12_W_IO/E2BEGb[3]
+ Tile_X0Y12_W_IO/E2BEGb[4] Tile_X0Y12_W_IO/E2BEGb[5] Tile_X0Y12_W_IO/E2BEGb[6] Tile_X0Y12_W_IO/E2BEGb[7]
+ Tile_X0Y12_W_IO/E6BEG[0] Tile_X0Y12_W_IO/E6BEG[10] Tile_X0Y12_W_IO/E6BEG[11] Tile_X0Y12_W_IO/E6BEG[1]
+ Tile_X0Y12_W_IO/E6BEG[2] Tile_X0Y12_W_IO/E6BEG[3] Tile_X0Y12_W_IO/E6BEG[4] Tile_X0Y12_W_IO/E6BEG[5]
+ Tile_X0Y12_W_IO/E6BEG[6] Tile_X0Y12_W_IO/E6BEG[7] Tile_X0Y12_W_IO/E6BEG[8] Tile_X0Y12_W_IO/E6BEG[9]
+ Tile_X0Y12_W_IO/EE4BEG[0] Tile_X0Y12_W_IO/EE4BEG[10] Tile_X0Y12_W_IO/EE4BEG[11]
+ Tile_X0Y12_W_IO/EE4BEG[12] Tile_X0Y12_W_IO/EE4BEG[13] Tile_X0Y12_W_IO/EE4BEG[14]
+ Tile_X0Y12_W_IO/EE4BEG[15] Tile_X0Y12_W_IO/EE4BEG[1] Tile_X0Y12_W_IO/EE4BEG[2] Tile_X0Y12_W_IO/EE4BEG[3]
+ Tile_X0Y12_W_IO/EE4BEG[4] Tile_X0Y12_W_IO/EE4BEG[5] Tile_X0Y12_W_IO/EE4BEG[6] Tile_X0Y12_W_IO/EE4BEG[7]
+ Tile_X0Y12_W_IO/EE4BEG[8] Tile_X0Y12_W_IO/EE4BEG[9] FrameData[384] FrameData[394]
+ FrameData[395] FrameData[396] FrameData[397] FrameData[398] FrameData[399] FrameData[400]
+ FrameData[401] FrameData[402] FrameData[403] FrameData[385] FrameData[404] FrameData[405]
+ FrameData[406] FrameData[407] FrameData[408] FrameData[409] FrameData[410] FrameData[411]
+ FrameData[412] FrameData[413] FrameData[386] FrameData[414] FrameData[415] FrameData[387]
+ FrameData[388] FrameData[389] FrameData[390] FrameData[391] FrameData[392] FrameData[393]
+ Tile_X1Y12_LUT4AB/FrameData[0] Tile_X1Y12_LUT4AB/FrameData[10] Tile_X1Y12_LUT4AB/FrameData[11]
+ Tile_X1Y12_LUT4AB/FrameData[12] Tile_X1Y12_LUT4AB/FrameData[13] Tile_X1Y12_LUT4AB/FrameData[14]
+ Tile_X1Y12_LUT4AB/FrameData[15] Tile_X1Y12_LUT4AB/FrameData[16] Tile_X1Y12_LUT4AB/FrameData[17]
+ Tile_X1Y12_LUT4AB/FrameData[18] Tile_X1Y12_LUT4AB/FrameData[19] Tile_X1Y12_LUT4AB/FrameData[1]
+ Tile_X1Y12_LUT4AB/FrameData[20] Tile_X1Y12_LUT4AB/FrameData[21] Tile_X1Y12_LUT4AB/FrameData[22]
+ Tile_X1Y12_LUT4AB/FrameData[23] Tile_X1Y12_LUT4AB/FrameData[24] Tile_X1Y12_LUT4AB/FrameData[25]
+ Tile_X1Y12_LUT4AB/FrameData[26] Tile_X1Y12_LUT4AB/FrameData[27] Tile_X1Y12_LUT4AB/FrameData[28]
+ Tile_X1Y12_LUT4AB/FrameData[29] Tile_X1Y12_LUT4AB/FrameData[2] Tile_X1Y12_LUT4AB/FrameData[30]
+ Tile_X1Y12_LUT4AB/FrameData[31] Tile_X1Y12_LUT4AB/FrameData[3] Tile_X1Y12_LUT4AB/FrameData[4]
+ Tile_X1Y12_LUT4AB/FrameData[5] Tile_X1Y12_LUT4AB/FrameData[6] Tile_X1Y12_LUT4AB/FrameData[7]
+ Tile_X1Y12_LUT4AB/FrameData[8] Tile_X1Y12_LUT4AB/FrameData[9] Tile_X0Y12_W_IO/FrameStrobe[0]
+ Tile_X0Y12_W_IO/FrameStrobe[10] Tile_X0Y12_W_IO/FrameStrobe[11] Tile_X0Y12_W_IO/FrameStrobe[12]
+ Tile_X0Y12_W_IO/FrameStrobe[13] Tile_X0Y12_W_IO/FrameStrobe[14] Tile_X0Y12_W_IO/FrameStrobe[15]
+ Tile_X0Y12_W_IO/FrameStrobe[16] Tile_X0Y12_W_IO/FrameStrobe[17] Tile_X0Y12_W_IO/FrameStrobe[18]
+ Tile_X0Y12_W_IO/FrameStrobe[19] Tile_X0Y12_W_IO/FrameStrobe[1] Tile_X0Y12_W_IO/FrameStrobe[2]
+ Tile_X0Y12_W_IO/FrameStrobe[3] Tile_X0Y12_W_IO/FrameStrobe[4] Tile_X0Y12_W_IO/FrameStrobe[5]
+ Tile_X0Y12_W_IO/FrameStrobe[6] Tile_X0Y12_W_IO/FrameStrobe[7] Tile_X0Y12_W_IO/FrameStrobe[8]
+ Tile_X0Y12_W_IO/FrameStrobe[9] Tile_X0Y11_W_IO/FrameStrobe[0] Tile_X0Y11_W_IO/FrameStrobe[10]
+ Tile_X0Y11_W_IO/FrameStrobe[11] Tile_X0Y11_W_IO/FrameStrobe[12] Tile_X0Y11_W_IO/FrameStrobe[13]
+ Tile_X0Y11_W_IO/FrameStrobe[14] Tile_X0Y11_W_IO/FrameStrobe[15] Tile_X0Y11_W_IO/FrameStrobe[16]
+ Tile_X0Y11_W_IO/FrameStrobe[17] Tile_X0Y11_W_IO/FrameStrobe[18] Tile_X0Y11_W_IO/FrameStrobe[19]
+ Tile_X0Y11_W_IO/FrameStrobe[1] Tile_X0Y11_W_IO/FrameStrobe[2] Tile_X0Y11_W_IO/FrameStrobe[3]
+ Tile_X0Y11_W_IO/FrameStrobe[4] Tile_X0Y11_W_IO/FrameStrobe[5] Tile_X0Y11_W_IO/FrameStrobe[6]
+ Tile_X0Y11_W_IO/FrameStrobe[7] Tile_X0Y11_W_IO/FrameStrobe[8] Tile_X0Y11_W_IO/FrameStrobe[9]
+ Tile_X0Y12_W_IO/UserCLK Tile_X0Y11_W_IO/UserCLK VGND VPWR Tile_X0Y12_W_IO/W1END[0]
+ Tile_X0Y12_W_IO/W1END[1] Tile_X0Y12_W_IO/W1END[2] Tile_X0Y12_W_IO/W1END[3] Tile_X0Y12_W_IO/W2END[0]
+ Tile_X0Y12_W_IO/W2END[1] Tile_X0Y12_W_IO/W2END[2] Tile_X0Y12_W_IO/W2END[3] Tile_X0Y12_W_IO/W2END[4]
+ Tile_X0Y12_W_IO/W2END[5] Tile_X0Y12_W_IO/W2END[6] Tile_X0Y12_W_IO/W2END[7] Tile_X0Y12_W_IO/W2MID[0]
+ Tile_X0Y12_W_IO/W2MID[1] Tile_X0Y12_W_IO/W2MID[2] Tile_X0Y12_W_IO/W2MID[3] Tile_X0Y12_W_IO/W2MID[4]
+ Tile_X0Y12_W_IO/W2MID[5] Tile_X0Y12_W_IO/W2MID[6] Tile_X0Y12_W_IO/W2MID[7] Tile_X0Y12_W_IO/W6END[0]
+ Tile_X0Y12_W_IO/W6END[10] Tile_X0Y12_W_IO/W6END[11] Tile_X0Y12_W_IO/W6END[1] Tile_X0Y12_W_IO/W6END[2]
+ Tile_X0Y12_W_IO/W6END[3] Tile_X0Y12_W_IO/W6END[4] Tile_X0Y12_W_IO/W6END[5] Tile_X0Y12_W_IO/W6END[6]
+ Tile_X0Y12_W_IO/W6END[7] Tile_X0Y12_W_IO/W6END[8] Tile_X0Y12_W_IO/W6END[9] Tile_X0Y12_W_IO/WW4END[0]
+ Tile_X0Y12_W_IO/WW4END[10] Tile_X0Y12_W_IO/WW4END[11] Tile_X0Y12_W_IO/WW4END[12]
+ Tile_X0Y12_W_IO/WW4END[13] Tile_X0Y12_W_IO/WW4END[14] Tile_X0Y12_W_IO/WW4END[15]
+ Tile_X0Y12_W_IO/WW4END[1] Tile_X0Y12_W_IO/WW4END[2] Tile_X0Y12_W_IO/WW4END[3] Tile_X0Y12_W_IO/WW4END[4]
+ Tile_X0Y12_W_IO/WW4END[5] Tile_X0Y12_W_IO/WW4END[6] Tile_X0Y12_W_IO/WW4END[7] Tile_X0Y12_W_IO/WW4END[8]
+ Tile_X0Y12_W_IO/WW4END[9] W_IO
XTile_X10Y11_IHP_SRAM Tile_X10Y12_ADDR_SRAM0 Tile_X10Y12_ADDR_SRAM1 Tile_X10Y12_ADDR_SRAM2
+ Tile_X10Y12_ADDR_SRAM3 Tile_X10Y12_ADDR_SRAM4 Tile_X10Y12_ADDR_SRAM5 Tile_X10Y12_ADDR_SRAM6
+ Tile_X10Y12_ADDR_SRAM7 Tile_X10Y12_ADDR_SRAM8 Tile_X10Y12_ADDR_SRAM9 Tile_X10Y12_BM_SRAM0
+ Tile_X10Y12_BM_SRAM1 Tile_X10Y12_BM_SRAM10 Tile_X10Y12_BM_SRAM11 Tile_X10Y12_BM_SRAM12
+ Tile_X10Y12_BM_SRAM13 Tile_X10Y12_BM_SRAM14 Tile_X10Y12_BM_SRAM15 Tile_X10Y12_BM_SRAM16
+ Tile_X10Y12_BM_SRAM17 Tile_X10Y12_BM_SRAM18 Tile_X10Y12_BM_SRAM19 Tile_X10Y12_BM_SRAM2
+ Tile_X10Y12_BM_SRAM20 Tile_X10Y12_BM_SRAM21 Tile_X10Y12_BM_SRAM22 Tile_X10Y12_BM_SRAM23
+ Tile_X10Y12_BM_SRAM24 Tile_X10Y12_BM_SRAM25 Tile_X10Y12_BM_SRAM26 Tile_X10Y12_BM_SRAM27
+ Tile_X10Y12_BM_SRAM28 Tile_X10Y12_BM_SRAM29 Tile_X10Y12_BM_SRAM3 Tile_X10Y12_BM_SRAM30
+ Tile_X10Y12_BM_SRAM31 Tile_X10Y12_BM_SRAM4 Tile_X10Y12_BM_SRAM5 Tile_X10Y12_BM_SRAM6
+ Tile_X10Y12_BM_SRAM7 Tile_X10Y12_BM_SRAM8 Tile_X10Y12_BM_SRAM9 Tile_X10Y12_CLK_SRAM
+ Tile_X10Y12_CONFIGURED_top Tile_X10Y12_DIN_SRAM0 Tile_X10Y12_DIN_SRAM1 Tile_X10Y12_DIN_SRAM10
+ Tile_X10Y12_DIN_SRAM11 Tile_X10Y12_DIN_SRAM12 Tile_X10Y12_DIN_SRAM13 Tile_X10Y12_DIN_SRAM14
+ Tile_X10Y12_DIN_SRAM15 Tile_X10Y12_DIN_SRAM16 Tile_X10Y12_DIN_SRAM17 Tile_X10Y12_DIN_SRAM18
+ Tile_X10Y12_DIN_SRAM19 Tile_X10Y12_DIN_SRAM2 Tile_X10Y12_DIN_SRAM20 Tile_X10Y12_DIN_SRAM21
+ Tile_X10Y12_DIN_SRAM22 Tile_X10Y12_DIN_SRAM23 Tile_X10Y12_DIN_SRAM24 Tile_X10Y12_DIN_SRAM25
+ Tile_X10Y12_DIN_SRAM26 Tile_X10Y12_DIN_SRAM27 Tile_X10Y12_DIN_SRAM28 Tile_X10Y12_DIN_SRAM29
+ Tile_X10Y12_DIN_SRAM3 Tile_X10Y12_DIN_SRAM30 Tile_X10Y12_DIN_SRAM31 Tile_X10Y12_DIN_SRAM4
+ Tile_X10Y12_DIN_SRAM5 Tile_X10Y12_DIN_SRAM6 Tile_X10Y12_DIN_SRAM7 Tile_X10Y12_DIN_SRAM8
+ Tile_X10Y12_DIN_SRAM9 Tile_X10Y12_DOUT_SRAM0 Tile_X10Y12_DOUT_SRAM1 Tile_X10Y12_DOUT_SRAM10
+ Tile_X10Y12_DOUT_SRAM11 Tile_X10Y12_DOUT_SRAM12 Tile_X10Y12_DOUT_SRAM13 Tile_X10Y12_DOUT_SRAM14
+ Tile_X10Y12_DOUT_SRAM15 Tile_X10Y12_DOUT_SRAM16 Tile_X10Y12_DOUT_SRAM17 Tile_X10Y12_DOUT_SRAM18
+ Tile_X10Y12_DOUT_SRAM19 Tile_X10Y12_DOUT_SRAM2 Tile_X10Y12_DOUT_SRAM20 Tile_X10Y12_DOUT_SRAM21
+ Tile_X10Y12_DOUT_SRAM22 Tile_X10Y12_DOUT_SRAM23 Tile_X10Y12_DOUT_SRAM24 Tile_X10Y12_DOUT_SRAM25
+ Tile_X10Y12_DOUT_SRAM26 Tile_X10Y12_DOUT_SRAM27 Tile_X10Y12_DOUT_SRAM28 Tile_X10Y12_DOUT_SRAM29
+ Tile_X10Y12_DOUT_SRAM3 Tile_X10Y12_DOUT_SRAM30 Tile_X10Y12_DOUT_SRAM31 Tile_X10Y12_DOUT_SRAM4
+ Tile_X10Y12_DOUT_SRAM5 Tile_X10Y12_DOUT_SRAM6 Tile_X10Y12_DOUT_SRAM7 Tile_X10Y12_DOUT_SRAM8
+ Tile_X10Y12_DOUT_SRAM9 Tile_X10Y12_MEN_SRAM Tile_X10Y12_REN_SRAM Tile_X10Y12_TIE_HIGH_SRAM
+ Tile_X10Y12_TIE_LOW_SRAM Tile_X9Y11_LUT4AB/E1BEG[0] Tile_X9Y11_LUT4AB/E1BEG[1] Tile_X9Y11_LUT4AB/E1BEG[2]
+ Tile_X9Y11_LUT4AB/E1BEG[3] Tile_X9Y11_LUT4AB/E2BEGb[0] Tile_X9Y11_LUT4AB/E2BEGb[1]
+ Tile_X9Y11_LUT4AB/E2BEGb[2] Tile_X9Y11_LUT4AB/E2BEGb[3] Tile_X9Y11_LUT4AB/E2BEGb[4]
+ Tile_X9Y11_LUT4AB/E2BEGb[5] Tile_X9Y11_LUT4AB/E2BEGb[6] Tile_X9Y11_LUT4AB/E2BEGb[7]
+ Tile_X9Y11_LUT4AB/E2BEG[0] Tile_X9Y11_LUT4AB/E2BEG[1] Tile_X9Y11_LUT4AB/E2BEG[2]
+ Tile_X9Y11_LUT4AB/E2BEG[3] Tile_X9Y11_LUT4AB/E2BEG[4] Tile_X9Y11_LUT4AB/E2BEG[5]
+ Tile_X9Y11_LUT4AB/E2BEG[6] Tile_X9Y11_LUT4AB/E2BEG[7] Tile_X9Y11_LUT4AB/E6BEG[0]
+ Tile_X9Y11_LUT4AB/E6BEG[10] Tile_X9Y11_LUT4AB/E6BEG[11] Tile_X9Y11_LUT4AB/E6BEG[1]
+ Tile_X9Y11_LUT4AB/E6BEG[2] Tile_X9Y11_LUT4AB/E6BEG[3] Tile_X9Y11_LUT4AB/E6BEG[4]
+ Tile_X9Y11_LUT4AB/E6BEG[5] Tile_X9Y11_LUT4AB/E6BEG[6] Tile_X9Y11_LUT4AB/E6BEG[7]
+ Tile_X9Y11_LUT4AB/E6BEG[8] Tile_X9Y11_LUT4AB/E6BEG[9] Tile_X9Y11_LUT4AB/EE4BEG[0]
+ Tile_X9Y11_LUT4AB/EE4BEG[10] Tile_X9Y11_LUT4AB/EE4BEG[11] Tile_X9Y11_LUT4AB/EE4BEG[12]
+ Tile_X9Y11_LUT4AB/EE4BEG[13] Tile_X9Y11_LUT4AB/EE4BEG[14] Tile_X9Y11_LUT4AB/EE4BEG[15]
+ Tile_X9Y11_LUT4AB/EE4BEG[1] Tile_X9Y11_LUT4AB/EE4BEG[2] Tile_X9Y11_LUT4AB/EE4BEG[3]
+ Tile_X9Y11_LUT4AB/EE4BEG[4] Tile_X9Y11_LUT4AB/EE4BEG[5] Tile_X9Y11_LUT4AB/EE4BEG[6]
+ Tile_X9Y11_LUT4AB/EE4BEG[7] Tile_X9Y11_LUT4AB/EE4BEG[8] Tile_X9Y11_LUT4AB/EE4BEG[9]
+ Tile_X9Y11_LUT4AB/FrameData_O[0] Tile_X9Y11_LUT4AB/FrameData_O[10] Tile_X9Y11_LUT4AB/FrameData_O[11]
+ Tile_X9Y11_LUT4AB/FrameData_O[12] Tile_X9Y11_LUT4AB/FrameData_O[13] Tile_X9Y11_LUT4AB/FrameData_O[14]
+ Tile_X9Y11_LUT4AB/FrameData_O[15] Tile_X9Y11_LUT4AB/FrameData_O[16] Tile_X9Y11_LUT4AB/FrameData_O[17]
+ Tile_X9Y11_LUT4AB/FrameData_O[18] Tile_X9Y11_LUT4AB/FrameData_O[19] Tile_X9Y11_LUT4AB/FrameData_O[1]
+ Tile_X9Y11_LUT4AB/FrameData_O[20] Tile_X9Y11_LUT4AB/FrameData_O[21] Tile_X9Y11_LUT4AB/FrameData_O[22]
+ Tile_X9Y11_LUT4AB/FrameData_O[23] Tile_X9Y11_LUT4AB/FrameData_O[24] Tile_X9Y11_LUT4AB/FrameData_O[25]
+ Tile_X9Y11_LUT4AB/FrameData_O[26] Tile_X9Y11_LUT4AB/FrameData_O[27] Tile_X9Y11_LUT4AB/FrameData_O[28]
+ Tile_X9Y11_LUT4AB/FrameData_O[29] Tile_X9Y11_LUT4AB/FrameData_O[2] Tile_X9Y11_LUT4AB/FrameData_O[30]
+ Tile_X9Y11_LUT4AB/FrameData_O[31] Tile_X9Y11_LUT4AB/FrameData_O[3] Tile_X9Y11_LUT4AB/FrameData_O[4]
+ Tile_X9Y11_LUT4AB/FrameData_O[5] Tile_X9Y11_LUT4AB/FrameData_O[6] Tile_X9Y11_LUT4AB/FrameData_O[7]
+ Tile_X9Y11_LUT4AB/FrameData_O[8] Tile_X9Y11_LUT4AB/FrameData_O[9] Tile_X10Y11_IHP_SRAM/Tile_X0Y0_FrameData_O[0]
+ Tile_X10Y11_IHP_SRAM/Tile_X0Y0_FrameData_O[10] Tile_X10Y11_IHP_SRAM/Tile_X0Y0_FrameData_O[11]
+ Tile_X10Y11_IHP_SRAM/Tile_X0Y0_FrameData_O[12] Tile_X10Y11_IHP_SRAM/Tile_X0Y0_FrameData_O[13]
+ Tile_X10Y11_IHP_SRAM/Tile_X0Y0_FrameData_O[14] Tile_X10Y11_IHP_SRAM/Tile_X0Y0_FrameData_O[15]
+ Tile_X10Y11_IHP_SRAM/Tile_X0Y0_FrameData_O[16] Tile_X10Y11_IHP_SRAM/Tile_X0Y0_FrameData_O[17]
+ Tile_X10Y11_IHP_SRAM/Tile_X0Y0_FrameData_O[18] Tile_X10Y11_IHP_SRAM/Tile_X0Y0_FrameData_O[19]
+ Tile_X10Y11_IHP_SRAM/Tile_X0Y0_FrameData_O[1] Tile_X10Y11_IHP_SRAM/Tile_X0Y0_FrameData_O[20]
+ Tile_X10Y11_IHP_SRAM/Tile_X0Y0_FrameData_O[21] Tile_X10Y11_IHP_SRAM/Tile_X0Y0_FrameData_O[22]
+ Tile_X10Y11_IHP_SRAM/Tile_X0Y0_FrameData_O[23] Tile_X10Y11_IHP_SRAM/Tile_X0Y0_FrameData_O[24]
+ Tile_X10Y11_IHP_SRAM/Tile_X0Y0_FrameData_O[25] Tile_X10Y11_IHP_SRAM/Tile_X0Y0_FrameData_O[26]
+ Tile_X10Y11_IHP_SRAM/Tile_X0Y0_FrameData_O[27] Tile_X10Y11_IHP_SRAM/Tile_X0Y0_FrameData_O[28]
+ Tile_X10Y11_IHP_SRAM/Tile_X0Y0_FrameData_O[29] Tile_X10Y11_IHP_SRAM/Tile_X0Y0_FrameData_O[2]
+ Tile_X10Y11_IHP_SRAM/Tile_X0Y0_FrameData_O[30] Tile_X10Y11_IHP_SRAM/Tile_X0Y0_FrameData_O[31]
+ Tile_X10Y11_IHP_SRAM/Tile_X0Y0_FrameData_O[3] Tile_X10Y11_IHP_SRAM/Tile_X0Y0_FrameData_O[4]
+ Tile_X10Y11_IHP_SRAM/Tile_X0Y0_FrameData_O[5] Tile_X10Y11_IHP_SRAM/Tile_X0Y0_FrameData_O[6]
+ Tile_X10Y11_IHP_SRAM/Tile_X0Y0_FrameData_O[7] Tile_X10Y11_IHP_SRAM/Tile_X0Y0_FrameData_O[8]
+ Tile_X10Y11_IHP_SRAM/Tile_X0Y0_FrameData_O[9] Tile_X10Y9_IHP_SRAM/Tile_X0Y1_FrameStrobe[0]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y1_FrameStrobe[10] Tile_X10Y9_IHP_SRAM/Tile_X0Y1_FrameStrobe[11]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y1_FrameStrobe[12] Tile_X10Y9_IHP_SRAM/Tile_X0Y1_FrameStrobe[13]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y1_FrameStrobe[14] Tile_X10Y9_IHP_SRAM/Tile_X0Y1_FrameStrobe[15]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y1_FrameStrobe[16] Tile_X10Y9_IHP_SRAM/Tile_X0Y1_FrameStrobe[17]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y1_FrameStrobe[18] Tile_X10Y9_IHP_SRAM/Tile_X0Y1_FrameStrobe[19]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y1_FrameStrobe[1] Tile_X10Y9_IHP_SRAM/Tile_X0Y1_FrameStrobe[2]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y1_FrameStrobe[3] Tile_X10Y9_IHP_SRAM/Tile_X0Y1_FrameStrobe[4]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y1_FrameStrobe[5] Tile_X10Y9_IHP_SRAM/Tile_X0Y1_FrameStrobe[6]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y1_FrameStrobe[7] Tile_X10Y9_IHP_SRAM/Tile_X0Y1_FrameStrobe[8]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y1_FrameStrobe[9] Tile_X10Y9_IHP_SRAM/Tile_X0Y1_N1END[0]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y1_N1END[1] Tile_X10Y9_IHP_SRAM/Tile_X0Y1_N1END[2] Tile_X10Y9_IHP_SRAM/Tile_X0Y1_N1END[3]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y1_N2MID[0] Tile_X10Y9_IHP_SRAM/Tile_X0Y1_N2MID[1] Tile_X10Y9_IHP_SRAM/Tile_X0Y1_N2MID[2]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y1_N2MID[3] Tile_X10Y9_IHP_SRAM/Tile_X0Y1_N2MID[4] Tile_X10Y9_IHP_SRAM/Tile_X0Y1_N2MID[5]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y1_N2MID[6] Tile_X10Y9_IHP_SRAM/Tile_X0Y1_N2MID[7] Tile_X10Y9_IHP_SRAM/Tile_X0Y1_N2END[0]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y1_N2END[1] Tile_X10Y9_IHP_SRAM/Tile_X0Y1_N2END[2] Tile_X10Y9_IHP_SRAM/Tile_X0Y1_N2END[3]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y1_N2END[4] Tile_X10Y9_IHP_SRAM/Tile_X0Y1_N2END[5] Tile_X10Y9_IHP_SRAM/Tile_X0Y1_N2END[6]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y1_N2END[7] Tile_X10Y9_IHP_SRAM/Tile_X0Y1_N4END[0] Tile_X10Y9_IHP_SRAM/Tile_X0Y1_N4END[10]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y1_N4END[11] Tile_X10Y9_IHP_SRAM/Tile_X0Y1_N4END[12]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y1_N4END[13] Tile_X10Y9_IHP_SRAM/Tile_X0Y1_N4END[14]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y1_N4END[15] Tile_X10Y9_IHP_SRAM/Tile_X0Y1_N4END[1] Tile_X10Y9_IHP_SRAM/Tile_X0Y1_N4END[2]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y1_N4END[3] Tile_X10Y9_IHP_SRAM/Tile_X0Y1_N4END[4] Tile_X10Y9_IHP_SRAM/Tile_X0Y1_N4END[5]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y1_N4END[6] Tile_X10Y9_IHP_SRAM/Tile_X0Y1_N4END[7] Tile_X10Y9_IHP_SRAM/Tile_X0Y1_N4END[8]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y1_N4END[9] Tile_X10Y9_IHP_SRAM/Tile_X0Y1_S1BEG[0] Tile_X10Y9_IHP_SRAM/Tile_X0Y1_S1BEG[1]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y1_S1BEG[2] Tile_X10Y9_IHP_SRAM/Tile_X0Y1_S1BEG[3] Tile_X10Y9_IHP_SRAM/Tile_X0Y1_S2BEGb[0]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y1_S2BEGb[1] Tile_X10Y9_IHP_SRAM/Tile_X0Y1_S2BEGb[2]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y1_S2BEGb[3] Tile_X10Y9_IHP_SRAM/Tile_X0Y1_S2BEGb[4]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y1_S2BEGb[5] Tile_X10Y9_IHP_SRAM/Tile_X0Y1_S2BEGb[6]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y1_S2BEGb[7] Tile_X10Y9_IHP_SRAM/Tile_X0Y1_S2BEG[0] Tile_X10Y9_IHP_SRAM/Tile_X0Y1_S2BEG[1]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y1_S2BEG[2] Tile_X10Y9_IHP_SRAM/Tile_X0Y1_S2BEG[3] Tile_X10Y9_IHP_SRAM/Tile_X0Y1_S2BEG[4]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y1_S2BEG[5] Tile_X10Y9_IHP_SRAM/Tile_X0Y1_S2BEG[6] Tile_X10Y9_IHP_SRAM/Tile_X0Y1_S2BEG[7]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y1_S4BEG[0] Tile_X10Y9_IHP_SRAM/Tile_X0Y1_S4BEG[10] Tile_X10Y9_IHP_SRAM/Tile_X0Y1_S4BEG[11]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y1_S4BEG[12] Tile_X10Y9_IHP_SRAM/Tile_X0Y1_S4BEG[13]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y1_S4BEG[14] Tile_X10Y9_IHP_SRAM/Tile_X0Y1_S4BEG[15]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y1_S4BEG[1] Tile_X10Y9_IHP_SRAM/Tile_X0Y1_S4BEG[2] Tile_X10Y9_IHP_SRAM/Tile_X0Y1_S4BEG[3]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y1_S4BEG[4] Tile_X10Y9_IHP_SRAM/Tile_X0Y1_S4BEG[5] Tile_X10Y9_IHP_SRAM/Tile_X0Y1_S4BEG[6]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y1_S4BEG[7] Tile_X10Y9_IHP_SRAM/Tile_X0Y1_S4BEG[8] Tile_X10Y9_IHP_SRAM/Tile_X0Y1_S4BEG[9]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y1_UserCLK Tile_X9Y11_LUT4AB/W1END[0] Tile_X9Y11_LUT4AB/W1END[1]
+ Tile_X9Y11_LUT4AB/W1END[2] Tile_X9Y11_LUT4AB/W1END[3] Tile_X9Y11_LUT4AB/W2MID[0]
+ Tile_X9Y11_LUT4AB/W2MID[1] Tile_X9Y11_LUT4AB/W2MID[2] Tile_X9Y11_LUT4AB/W2MID[3]
+ Tile_X9Y11_LUT4AB/W2MID[4] Tile_X9Y11_LUT4AB/W2MID[5] Tile_X9Y11_LUT4AB/W2MID[6]
+ Tile_X9Y11_LUT4AB/W2MID[7] Tile_X9Y11_LUT4AB/W2END[0] Tile_X9Y11_LUT4AB/W2END[1]
+ Tile_X9Y11_LUT4AB/W2END[2] Tile_X9Y11_LUT4AB/W2END[3] Tile_X9Y11_LUT4AB/W2END[4]
+ Tile_X9Y11_LUT4AB/W2END[5] Tile_X9Y11_LUT4AB/W2END[6] Tile_X9Y11_LUT4AB/W2END[7]
+ Tile_X9Y11_LUT4AB/W6END[0] Tile_X9Y11_LUT4AB/W6END[10] Tile_X9Y11_LUT4AB/W6END[11]
+ Tile_X9Y11_LUT4AB/W6END[1] Tile_X9Y11_LUT4AB/W6END[2] Tile_X9Y11_LUT4AB/W6END[3]
+ Tile_X9Y11_LUT4AB/W6END[4] Tile_X9Y11_LUT4AB/W6END[5] Tile_X9Y11_LUT4AB/W6END[6]
+ Tile_X9Y11_LUT4AB/W6END[7] Tile_X9Y11_LUT4AB/W6END[8] Tile_X9Y11_LUT4AB/W6END[9]
+ Tile_X9Y11_LUT4AB/WW4END[0] Tile_X9Y11_LUT4AB/WW4END[10] Tile_X9Y11_LUT4AB/WW4END[11]
+ Tile_X9Y11_LUT4AB/WW4END[12] Tile_X9Y11_LUT4AB/WW4END[13] Tile_X9Y11_LUT4AB/WW4END[14]
+ Tile_X9Y11_LUT4AB/WW4END[15] Tile_X9Y11_LUT4AB/WW4END[1] Tile_X9Y11_LUT4AB/WW4END[2]
+ Tile_X9Y11_LUT4AB/WW4END[3] Tile_X9Y11_LUT4AB/WW4END[4] Tile_X9Y11_LUT4AB/WW4END[5]
+ Tile_X9Y11_LUT4AB/WW4END[6] Tile_X9Y11_LUT4AB/WW4END[7] Tile_X9Y11_LUT4AB/WW4END[8]
+ Tile_X9Y11_LUT4AB/WW4END[9] Tile_X9Y12_LUT4AB/E1BEG[0] Tile_X9Y12_LUT4AB/E1BEG[1]
+ Tile_X9Y12_LUT4AB/E1BEG[2] Tile_X9Y12_LUT4AB/E1BEG[3] Tile_X9Y12_LUT4AB/E2BEGb[0]
+ Tile_X9Y12_LUT4AB/E2BEGb[1] Tile_X9Y12_LUT4AB/E2BEGb[2] Tile_X9Y12_LUT4AB/E2BEGb[3]
+ Tile_X9Y12_LUT4AB/E2BEGb[4] Tile_X9Y12_LUT4AB/E2BEGb[5] Tile_X9Y12_LUT4AB/E2BEGb[6]
+ Tile_X9Y12_LUT4AB/E2BEGb[7] Tile_X9Y12_LUT4AB/E2BEG[0] Tile_X9Y12_LUT4AB/E2BEG[1]
+ Tile_X9Y12_LUT4AB/E2BEG[2] Tile_X9Y12_LUT4AB/E2BEG[3] Tile_X9Y12_LUT4AB/E2BEG[4]
+ Tile_X9Y12_LUT4AB/E2BEG[5] Tile_X9Y12_LUT4AB/E2BEG[6] Tile_X9Y12_LUT4AB/E2BEG[7]
+ Tile_X9Y12_LUT4AB/E6BEG[0] Tile_X9Y12_LUT4AB/E6BEG[10] Tile_X9Y12_LUT4AB/E6BEG[11]
+ Tile_X9Y12_LUT4AB/E6BEG[1] Tile_X9Y12_LUT4AB/E6BEG[2] Tile_X9Y12_LUT4AB/E6BEG[3]
+ Tile_X9Y12_LUT4AB/E6BEG[4] Tile_X9Y12_LUT4AB/E6BEG[5] Tile_X9Y12_LUT4AB/E6BEG[6]
+ Tile_X9Y12_LUT4AB/E6BEG[7] Tile_X9Y12_LUT4AB/E6BEG[8] Tile_X9Y12_LUT4AB/E6BEG[9]
+ Tile_X9Y12_LUT4AB/EE4BEG[0] Tile_X9Y12_LUT4AB/EE4BEG[10] Tile_X9Y12_LUT4AB/EE4BEG[11]
+ Tile_X9Y12_LUT4AB/EE4BEG[12] Tile_X9Y12_LUT4AB/EE4BEG[13] Tile_X9Y12_LUT4AB/EE4BEG[14]
+ Tile_X9Y12_LUT4AB/EE4BEG[15] Tile_X9Y12_LUT4AB/EE4BEG[1] Tile_X9Y12_LUT4AB/EE4BEG[2]
+ Tile_X9Y12_LUT4AB/EE4BEG[3] Tile_X9Y12_LUT4AB/EE4BEG[4] Tile_X9Y12_LUT4AB/EE4BEG[5]
+ Tile_X9Y12_LUT4AB/EE4BEG[6] Tile_X9Y12_LUT4AB/EE4BEG[7] Tile_X9Y12_LUT4AB/EE4BEG[8]
+ Tile_X9Y12_LUT4AB/EE4BEG[9] Tile_X9Y12_LUT4AB/FrameData_O[0] Tile_X9Y12_LUT4AB/FrameData_O[10]
+ Tile_X9Y12_LUT4AB/FrameData_O[11] Tile_X9Y12_LUT4AB/FrameData_O[12] Tile_X9Y12_LUT4AB/FrameData_O[13]
+ Tile_X9Y12_LUT4AB/FrameData_O[14] Tile_X9Y12_LUT4AB/FrameData_O[15] Tile_X9Y12_LUT4AB/FrameData_O[16]
+ Tile_X9Y12_LUT4AB/FrameData_O[17] Tile_X9Y12_LUT4AB/FrameData_O[18] Tile_X9Y12_LUT4AB/FrameData_O[19]
+ Tile_X9Y12_LUT4AB/FrameData_O[1] Tile_X9Y12_LUT4AB/FrameData_O[20] Tile_X9Y12_LUT4AB/FrameData_O[21]
+ Tile_X9Y12_LUT4AB/FrameData_O[22] Tile_X9Y12_LUT4AB/FrameData_O[23] Tile_X9Y12_LUT4AB/FrameData_O[24]
+ Tile_X9Y12_LUT4AB/FrameData_O[25] Tile_X9Y12_LUT4AB/FrameData_O[26] Tile_X9Y12_LUT4AB/FrameData_O[27]
+ Tile_X9Y12_LUT4AB/FrameData_O[28] Tile_X9Y12_LUT4AB/FrameData_O[29] Tile_X9Y12_LUT4AB/FrameData_O[2]
+ Tile_X9Y12_LUT4AB/FrameData_O[30] Tile_X9Y12_LUT4AB/FrameData_O[31] Tile_X9Y12_LUT4AB/FrameData_O[3]
+ Tile_X9Y12_LUT4AB/FrameData_O[4] Tile_X9Y12_LUT4AB/FrameData_O[5] Tile_X9Y12_LUT4AB/FrameData_O[6]
+ Tile_X9Y12_LUT4AB/FrameData_O[7] Tile_X9Y12_LUT4AB/FrameData_O[8] Tile_X9Y12_LUT4AB/FrameData_O[9]
+ Tile_X10Y11_IHP_SRAM/Tile_X0Y1_FrameData_O[0] Tile_X10Y11_IHP_SRAM/Tile_X0Y1_FrameData_O[10]
+ Tile_X10Y11_IHP_SRAM/Tile_X0Y1_FrameData_O[11] Tile_X10Y11_IHP_SRAM/Tile_X0Y1_FrameData_O[12]
+ Tile_X10Y11_IHP_SRAM/Tile_X0Y1_FrameData_O[13] Tile_X10Y11_IHP_SRAM/Tile_X0Y1_FrameData_O[14]
+ Tile_X10Y11_IHP_SRAM/Tile_X0Y1_FrameData_O[15] Tile_X10Y11_IHP_SRAM/Tile_X0Y1_FrameData_O[16]
+ Tile_X10Y11_IHP_SRAM/Tile_X0Y1_FrameData_O[17] Tile_X10Y11_IHP_SRAM/Tile_X0Y1_FrameData_O[18]
+ Tile_X10Y11_IHP_SRAM/Tile_X0Y1_FrameData_O[19] Tile_X10Y11_IHP_SRAM/Tile_X0Y1_FrameData_O[1]
+ Tile_X10Y11_IHP_SRAM/Tile_X0Y1_FrameData_O[20] Tile_X10Y11_IHP_SRAM/Tile_X0Y1_FrameData_O[21]
+ Tile_X10Y11_IHP_SRAM/Tile_X0Y1_FrameData_O[22] Tile_X10Y11_IHP_SRAM/Tile_X0Y1_FrameData_O[23]
+ Tile_X10Y11_IHP_SRAM/Tile_X0Y1_FrameData_O[24] Tile_X10Y11_IHP_SRAM/Tile_X0Y1_FrameData_O[25]
+ Tile_X10Y11_IHP_SRAM/Tile_X0Y1_FrameData_O[26] Tile_X10Y11_IHP_SRAM/Tile_X0Y1_FrameData_O[27]
+ Tile_X10Y11_IHP_SRAM/Tile_X0Y1_FrameData_O[28] Tile_X10Y11_IHP_SRAM/Tile_X0Y1_FrameData_O[29]
+ Tile_X10Y11_IHP_SRAM/Tile_X0Y1_FrameData_O[2] Tile_X10Y11_IHP_SRAM/Tile_X0Y1_FrameData_O[30]
+ Tile_X10Y11_IHP_SRAM/Tile_X0Y1_FrameData_O[31] Tile_X10Y11_IHP_SRAM/Tile_X0Y1_FrameData_O[3]
+ Tile_X10Y11_IHP_SRAM/Tile_X0Y1_FrameData_O[4] Tile_X10Y11_IHP_SRAM/Tile_X0Y1_FrameData_O[5]
+ Tile_X10Y11_IHP_SRAM/Tile_X0Y1_FrameData_O[6] Tile_X10Y11_IHP_SRAM/Tile_X0Y1_FrameData_O[7]
+ Tile_X10Y11_IHP_SRAM/Tile_X0Y1_FrameData_O[8] Tile_X10Y11_IHP_SRAM/Tile_X0Y1_FrameData_O[9]
+ Tile_X10Y11_IHP_SRAM/Tile_X0Y1_FrameStrobe[0] Tile_X10Y11_IHP_SRAM/Tile_X0Y1_FrameStrobe[10]
+ Tile_X10Y11_IHP_SRAM/Tile_X0Y1_FrameStrobe[11] Tile_X10Y11_IHP_SRAM/Tile_X0Y1_FrameStrobe[12]
+ Tile_X10Y11_IHP_SRAM/Tile_X0Y1_FrameStrobe[13] Tile_X10Y11_IHP_SRAM/Tile_X0Y1_FrameStrobe[14]
+ Tile_X10Y11_IHP_SRAM/Tile_X0Y1_FrameStrobe[15] Tile_X10Y11_IHP_SRAM/Tile_X0Y1_FrameStrobe[16]
+ Tile_X10Y11_IHP_SRAM/Tile_X0Y1_FrameStrobe[17] Tile_X10Y11_IHP_SRAM/Tile_X0Y1_FrameStrobe[18]
+ Tile_X10Y11_IHP_SRAM/Tile_X0Y1_FrameStrobe[19] Tile_X10Y11_IHP_SRAM/Tile_X0Y1_FrameStrobe[1]
+ Tile_X10Y11_IHP_SRAM/Tile_X0Y1_FrameStrobe[2] Tile_X10Y11_IHP_SRAM/Tile_X0Y1_FrameStrobe[3]
+ Tile_X10Y11_IHP_SRAM/Tile_X0Y1_FrameStrobe[4] Tile_X10Y11_IHP_SRAM/Tile_X0Y1_FrameStrobe[5]
+ Tile_X10Y11_IHP_SRAM/Tile_X0Y1_FrameStrobe[6] Tile_X10Y11_IHP_SRAM/Tile_X0Y1_FrameStrobe[7]
+ Tile_X10Y11_IHP_SRAM/Tile_X0Y1_FrameStrobe[8] Tile_X10Y11_IHP_SRAM/Tile_X0Y1_FrameStrobe[9]
+ Tile_X10Y13_IHP_SRAM/Tile_X0Y0_N1BEG[0] Tile_X10Y13_IHP_SRAM/Tile_X0Y0_N1BEG[1]
+ Tile_X10Y13_IHP_SRAM/Tile_X0Y0_N1BEG[2] Tile_X10Y13_IHP_SRAM/Tile_X0Y0_N1BEG[3]
+ Tile_X10Y11_IHP_SRAM/Tile_X0Y1_N2END[0] Tile_X10Y11_IHP_SRAM/Tile_X0Y1_N2END[1]
+ Tile_X10Y11_IHP_SRAM/Tile_X0Y1_N2END[2] Tile_X10Y11_IHP_SRAM/Tile_X0Y1_N2END[3]
+ Tile_X10Y11_IHP_SRAM/Tile_X0Y1_N2END[4] Tile_X10Y11_IHP_SRAM/Tile_X0Y1_N2END[5]
+ Tile_X10Y11_IHP_SRAM/Tile_X0Y1_N2END[6] Tile_X10Y11_IHP_SRAM/Tile_X0Y1_N2END[7]
+ Tile_X10Y13_IHP_SRAM/Tile_X0Y0_N2BEG[0] Tile_X10Y13_IHP_SRAM/Tile_X0Y0_N2BEG[1]
+ Tile_X10Y13_IHP_SRAM/Tile_X0Y0_N2BEG[2] Tile_X10Y13_IHP_SRAM/Tile_X0Y0_N2BEG[3]
+ Tile_X10Y13_IHP_SRAM/Tile_X0Y0_N2BEG[4] Tile_X10Y13_IHP_SRAM/Tile_X0Y0_N2BEG[5]
+ Tile_X10Y13_IHP_SRAM/Tile_X0Y0_N2BEG[6] Tile_X10Y13_IHP_SRAM/Tile_X0Y0_N2BEG[7]
+ Tile_X10Y13_IHP_SRAM/Tile_X0Y0_N4BEG[0] Tile_X10Y13_IHP_SRAM/Tile_X0Y0_N4BEG[10]
+ Tile_X10Y13_IHP_SRAM/Tile_X0Y0_N4BEG[11] Tile_X10Y13_IHP_SRAM/Tile_X0Y0_N4BEG[12]
+ Tile_X10Y13_IHP_SRAM/Tile_X0Y0_N4BEG[13] Tile_X10Y13_IHP_SRAM/Tile_X0Y0_N4BEG[14]
+ Tile_X10Y13_IHP_SRAM/Tile_X0Y0_N4BEG[15] Tile_X10Y13_IHP_SRAM/Tile_X0Y0_N4BEG[1]
+ Tile_X10Y13_IHP_SRAM/Tile_X0Y0_N4BEG[2] Tile_X10Y13_IHP_SRAM/Tile_X0Y0_N4BEG[3]
+ Tile_X10Y13_IHP_SRAM/Tile_X0Y0_N4BEG[4] Tile_X10Y13_IHP_SRAM/Tile_X0Y0_N4BEG[5]
+ Tile_X10Y13_IHP_SRAM/Tile_X0Y0_N4BEG[6] Tile_X10Y13_IHP_SRAM/Tile_X0Y0_N4BEG[7]
+ Tile_X10Y13_IHP_SRAM/Tile_X0Y0_N4BEG[8] Tile_X10Y13_IHP_SRAM/Tile_X0Y0_N4BEG[9]
+ Tile_X10Y13_IHP_SRAM/Tile_X0Y0_S1END[0] Tile_X10Y13_IHP_SRAM/Tile_X0Y0_S1END[1]
+ Tile_X10Y13_IHP_SRAM/Tile_X0Y0_S1END[2] Tile_X10Y13_IHP_SRAM/Tile_X0Y0_S1END[3]
+ Tile_X10Y13_IHP_SRAM/Tile_X0Y0_S2MID[0] Tile_X10Y13_IHP_SRAM/Tile_X0Y0_S2MID[1]
+ Tile_X10Y13_IHP_SRAM/Tile_X0Y0_S2MID[2] Tile_X10Y13_IHP_SRAM/Tile_X0Y0_S2MID[3]
+ Tile_X10Y13_IHP_SRAM/Tile_X0Y0_S2MID[4] Tile_X10Y13_IHP_SRAM/Tile_X0Y0_S2MID[5]
+ Tile_X10Y13_IHP_SRAM/Tile_X0Y0_S2MID[6] Tile_X10Y13_IHP_SRAM/Tile_X0Y0_S2MID[7]
+ Tile_X10Y13_IHP_SRAM/Tile_X0Y0_S2END[0] Tile_X10Y13_IHP_SRAM/Tile_X0Y0_S2END[1]
+ Tile_X10Y13_IHP_SRAM/Tile_X0Y0_S2END[2] Tile_X10Y13_IHP_SRAM/Tile_X0Y0_S2END[3]
+ Tile_X10Y13_IHP_SRAM/Tile_X0Y0_S2END[4] Tile_X10Y13_IHP_SRAM/Tile_X0Y0_S2END[5]
+ Tile_X10Y13_IHP_SRAM/Tile_X0Y0_S2END[6] Tile_X10Y13_IHP_SRAM/Tile_X0Y0_S2END[7]
+ Tile_X10Y13_IHP_SRAM/Tile_X0Y0_S4END[0] Tile_X10Y13_IHP_SRAM/Tile_X0Y0_S4END[10]
+ Tile_X10Y13_IHP_SRAM/Tile_X0Y0_S4END[11] Tile_X10Y13_IHP_SRAM/Tile_X0Y0_S4END[12]
+ Tile_X10Y13_IHP_SRAM/Tile_X0Y0_S4END[13] Tile_X10Y13_IHP_SRAM/Tile_X0Y0_S4END[14]
+ Tile_X10Y13_IHP_SRAM/Tile_X0Y0_S4END[15] Tile_X10Y13_IHP_SRAM/Tile_X0Y0_S4END[1]
+ Tile_X10Y13_IHP_SRAM/Tile_X0Y0_S4END[2] Tile_X10Y13_IHP_SRAM/Tile_X0Y0_S4END[3]
+ Tile_X10Y13_IHP_SRAM/Tile_X0Y0_S4END[4] Tile_X10Y13_IHP_SRAM/Tile_X0Y0_S4END[5]
+ Tile_X10Y13_IHP_SRAM/Tile_X0Y0_S4END[6] Tile_X10Y13_IHP_SRAM/Tile_X0Y0_S4END[7]
+ Tile_X10Y13_IHP_SRAM/Tile_X0Y0_S4END[8] Tile_X10Y13_IHP_SRAM/Tile_X0Y0_S4END[9]
+ Tile_X10Y11_IHP_SRAM/Tile_X0Y1_UserCLK Tile_X9Y12_LUT4AB/W1END[0] Tile_X9Y12_LUT4AB/W1END[1]
+ Tile_X9Y12_LUT4AB/W1END[2] Tile_X9Y12_LUT4AB/W1END[3] Tile_X9Y12_LUT4AB/W2MID[0]
+ Tile_X9Y12_LUT4AB/W2MID[1] Tile_X9Y12_LUT4AB/W2MID[2] Tile_X9Y12_LUT4AB/W2MID[3]
+ Tile_X9Y12_LUT4AB/W2MID[4] Tile_X9Y12_LUT4AB/W2MID[5] Tile_X9Y12_LUT4AB/W2MID[6]
+ Tile_X9Y12_LUT4AB/W2MID[7] Tile_X9Y12_LUT4AB/W2END[0] Tile_X9Y12_LUT4AB/W2END[1]
+ Tile_X9Y12_LUT4AB/W2END[2] Tile_X9Y12_LUT4AB/W2END[3] Tile_X9Y12_LUT4AB/W2END[4]
+ Tile_X9Y12_LUT4AB/W2END[5] Tile_X9Y12_LUT4AB/W2END[6] Tile_X9Y12_LUT4AB/W2END[7]
+ Tile_X9Y12_LUT4AB/W6END[0] Tile_X9Y12_LUT4AB/W6END[10] Tile_X9Y12_LUT4AB/W6END[11]
+ Tile_X9Y12_LUT4AB/W6END[1] Tile_X9Y12_LUT4AB/W6END[2] Tile_X9Y12_LUT4AB/W6END[3]
+ Tile_X9Y12_LUT4AB/W6END[4] Tile_X9Y12_LUT4AB/W6END[5] Tile_X9Y12_LUT4AB/W6END[6]
+ Tile_X9Y12_LUT4AB/W6END[7] Tile_X9Y12_LUT4AB/W6END[8] Tile_X9Y12_LUT4AB/W6END[9]
+ Tile_X9Y12_LUT4AB/WW4END[0] Tile_X9Y12_LUT4AB/WW4END[10] Tile_X9Y12_LUT4AB/WW4END[11]
+ Tile_X9Y12_LUT4AB/WW4END[12] Tile_X9Y12_LUT4AB/WW4END[13] Tile_X9Y12_LUT4AB/WW4END[14]
+ Tile_X9Y12_LUT4AB/WW4END[15] Tile_X9Y12_LUT4AB/WW4END[1] Tile_X9Y12_LUT4AB/WW4END[2]
+ Tile_X9Y12_LUT4AB/WW4END[3] Tile_X9Y12_LUT4AB/WW4END[4] Tile_X9Y12_LUT4AB/WW4END[5]
+ Tile_X9Y12_LUT4AB/WW4END[6] Tile_X9Y12_LUT4AB/WW4END[7] Tile_X9Y12_LUT4AB/WW4END[8]
+ Tile_X9Y12_LUT4AB/WW4END[9] VGND VPWR Tile_X10Y12_WEN_SRAM IHP_SRAM
XTile_X7Y3_DSP Tile_X8Y3_LUT4AB/E1END[0] Tile_X8Y3_LUT4AB/E1END[1] Tile_X8Y3_LUT4AB/E1END[2]
+ Tile_X8Y3_LUT4AB/E1END[3] Tile_X6Y3_LUT4AB/E1BEG[0] Tile_X6Y3_LUT4AB/E1BEG[1] Tile_X6Y3_LUT4AB/E1BEG[2]
+ Tile_X6Y3_LUT4AB/E1BEG[3] Tile_X8Y3_LUT4AB/E2MID[0] Tile_X8Y3_LUT4AB/E2MID[1] Tile_X8Y3_LUT4AB/E2MID[2]
+ Tile_X8Y3_LUT4AB/E2MID[3] Tile_X8Y3_LUT4AB/E2MID[4] Tile_X8Y3_LUT4AB/E2MID[5] Tile_X8Y3_LUT4AB/E2MID[6]
+ Tile_X8Y3_LUT4AB/E2MID[7] Tile_X8Y3_LUT4AB/E2END[0] Tile_X8Y3_LUT4AB/E2END[1] Tile_X8Y3_LUT4AB/E2END[2]
+ Tile_X8Y3_LUT4AB/E2END[3] Tile_X8Y3_LUT4AB/E2END[4] Tile_X8Y3_LUT4AB/E2END[5] Tile_X8Y3_LUT4AB/E2END[6]
+ Tile_X8Y3_LUT4AB/E2END[7] Tile_X6Y3_LUT4AB/E2BEGb[0] Tile_X6Y3_LUT4AB/E2BEGb[1]
+ Tile_X6Y3_LUT4AB/E2BEGb[2] Tile_X6Y3_LUT4AB/E2BEGb[3] Tile_X6Y3_LUT4AB/E2BEGb[4]
+ Tile_X6Y3_LUT4AB/E2BEGb[5] Tile_X6Y3_LUT4AB/E2BEGb[6] Tile_X6Y3_LUT4AB/E2BEGb[7]
+ Tile_X6Y3_LUT4AB/E2BEG[0] Tile_X6Y3_LUT4AB/E2BEG[1] Tile_X6Y3_LUT4AB/E2BEG[2] Tile_X6Y3_LUT4AB/E2BEG[3]
+ Tile_X6Y3_LUT4AB/E2BEG[4] Tile_X6Y3_LUT4AB/E2BEG[5] Tile_X6Y3_LUT4AB/E2BEG[6] Tile_X6Y3_LUT4AB/E2BEG[7]
+ Tile_X8Y3_LUT4AB/E6END[0] Tile_X8Y3_LUT4AB/E6END[10] Tile_X8Y3_LUT4AB/E6END[11]
+ Tile_X8Y3_LUT4AB/E6END[1] Tile_X8Y3_LUT4AB/E6END[2] Tile_X8Y3_LUT4AB/E6END[3] Tile_X8Y3_LUT4AB/E6END[4]
+ Tile_X8Y3_LUT4AB/E6END[5] Tile_X8Y3_LUT4AB/E6END[6] Tile_X8Y3_LUT4AB/E6END[7] Tile_X8Y3_LUT4AB/E6END[8]
+ Tile_X8Y3_LUT4AB/E6END[9] Tile_X6Y3_LUT4AB/E6BEG[0] Tile_X6Y3_LUT4AB/E6BEG[10] Tile_X6Y3_LUT4AB/E6BEG[11]
+ Tile_X6Y3_LUT4AB/E6BEG[1] Tile_X6Y3_LUT4AB/E6BEG[2] Tile_X6Y3_LUT4AB/E6BEG[3] Tile_X6Y3_LUT4AB/E6BEG[4]
+ Tile_X6Y3_LUT4AB/E6BEG[5] Tile_X6Y3_LUT4AB/E6BEG[6] Tile_X6Y3_LUT4AB/E6BEG[7] Tile_X6Y3_LUT4AB/E6BEG[8]
+ Tile_X6Y3_LUT4AB/E6BEG[9] Tile_X8Y3_LUT4AB/EE4END[0] Tile_X8Y3_LUT4AB/EE4END[10]
+ Tile_X8Y3_LUT4AB/EE4END[11] Tile_X8Y3_LUT4AB/EE4END[12] Tile_X8Y3_LUT4AB/EE4END[13]
+ Tile_X8Y3_LUT4AB/EE4END[14] Tile_X8Y3_LUT4AB/EE4END[15] Tile_X8Y3_LUT4AB/EE4END[1]
+ Tile_X8Y3_LUT4AB/EE4END[2] Tile_X8Y3_LUT4AB/EE4END[3] Tile_X8Y3_LUT4AB/EE4END[4]
+ Tile_X8Y3_LUT4AB/EE4END[5] Tile_X8Y3_LUT4AB/EE4END[6] Tile_X8Y3_LUT4AB/EE4END[7]
+ Tile_X8Y3_LUT4AB/EE4END[8] Tile_X8Y3_LUT4AB/EE4END[9] Tile_X6Y3_LUT4AB/EE4BEG[0]
+ Tile_X6Y3_LUT4AB/EE4BEG[10] Tile_X6Y3_LUT4AB/EE4BEG[11] Tile_X6Y3_LUT4AB/EE4BEG[12]
+ Tile_X6Y3_LUT4AB/EE4BEG[13] Tile_X6Y3_LUT4AB/EE4BEG[14] Tile_X6Y3_LUT4AB/EE4BEG[15]
+ Tile_X6Y3_LUT4AB/EE4BEG[1] Tile_X6Y3_LUT4AB/EE4BEG[2] Tile_X6Y3_LUT4AB/EE4BEG[3]
+ Tile_X6Y3_LUT4AB/EE4BEG[4] Tile_X6Y3_LUT4AB/EE4BEG[5] Tile_X6Y3_LUT4AB/EE4BEG[6]
+ Tile_X6Y3_LUT4AB/EE4BEG[7] Tile_X6Y3_LUT4AB/EE4BEG[8] Tile_X6Y3_LUT4AB/EE4BEG[9]
+ Tile_X6Y3_LUT4AB/FrameData_O[0] Tile_X6Y3_LUT4AB/FrameData_O[10] Tile_X6Y3_LUT4AB/FrameData_O[11]
+ Tile_X6Y3_LUT4AB/FrameData_O[12] Tile_X6Y3_LUT4AB/FrameData_O[13] Tile_X6Y3_LUT4AB/FrameData_O[14]
+ Tile_X6Y3_LUT4AB/FrameData_O[15] Tile_X6Y3_LUT4AB/FrameData_O[16] Tile_X6Y3_LUT4AB/FrameData_O[17]
+ Tile_X6Y3_LUT4AB/FrameData_O[18] Tile_X6Y3_LUT4AB/FrameData_O[19] Tile_X6Y3_LUT4AB/FrameData_O[1]
+ Tile_X6Y3_LUT4AB/FrameData_O[20] Tile_X6Y3_LUT4AB/FrameData_O[21] Tile_X6Y3_LUT4AB/FrameData_O[22]
+ Tile_X6Y3_LUT4AB/FrameData_O[23] Tile_X6Y3_LUT4AB/FrameData_O[24] Tile_X6Y3_LUT4AB/FrameData_O[25]
+ Tile_X6Y3_LUT4AB/FrameData_O[26] Tile_X6Y3_LUT4AB/FrameData_O[27] Tile_X6Y3_LUT4AB/FrameData_O[28]
+ Tile_X6Y3_LUT4AB/FrameData_O[29] Tile_X6Y3_LUT4AB/FrameData_O[2] Tile_X6Y3_LUT4AB/FrameData_O[30]
+ Tile_X6Y3_LUT4AB/FrameData_O[31] Tile_X6Y3_LUT4AB/FrameData_O[3] Tile_X6Y3_LUT4AB/FrameData_O[4]
+ Tile_X6Y3_LUT4AB/FrameData_O[5] Tile_X6Y3_LUT4AB/FrameData_O[6] Tile_X6Y3_LUT4AB/FrameData_O[7]
+ Tile_X6Y3_LUT4AB/FrameData_O[8] Tile_X6Y3_LUT4AB/FrameData_O[9] Tile_X8Y3_LUT4AB/FrameData[0]
+ Tile_X8Y3_LUT4AB/FrameData[10] Tile_X8Y3_LUT4AB/FrameData[11] Tile_X8Y3_LUT4AB/FrameData[12]
+ Tile_X8Y3_LUT4AB/FrameData[13] Tile_X8Y3_LUT4AB/FrameData[14] Tile_X8Y3_LUT4AB/FrameData[15]
+ Tile_X8Y3_LUT4AB/FrameData[16] Tile_X8Y3_LUT4AB/FrameData[17] Tile_X8Y3_LUT4AB/FrameData[18]
+ Tile_X8Y3_LUT4AB/FrameData[19] Tile_X8Y3_LUT4AB/FrameData[1] Tile_X8Y3_LUT4AB/FrameData[20]
+ Tile_X8Y3_LUT4AB/FrameData[21] Tile_X8Y3_LUT4AB/FrameData[22] Tile_X8Y3_LUT4AB/FrameData[23]
+ Tile_X8Y3_LUT4AB/FrameData[24] Tile_X8Y3_LUT4AB/FrameData[25] Tile_X8Y3_LUT4AB/FrameData[26]
+ Tile_X8Y3_LUT4AB/FrameData[27] Tile_X8Y3_LUT4AB/FrameData[28] Tile_X8Y3_LUT4AB/FrameData[29]
+ Tile_X8Y3_LUT4AB/FrameData[2] Tile_X8Y3_LUT4AB/FrameData[30] Tile_X8Y3_LUT4AB/FrameData[31]
+ Tile_X8Y3_LUT4AB/FrameData[3] Tile_X8Y3_LUT4AB/FrameData[4] Tile_X8Y3_LUT4AB/FrameData[5]
+ Tile_X8Y3_LUT4AB/FrameData[6] Tile_X8Y3_LUT4AB/FrameData[7] Tile_X8Y3_LUT4AB/FrameData[8]
+ Tile_X8Y3_LUT4AB/FrameData[9] Tile_X7Y1_DSP/Tile_X0Y1_FrameStrobe[0] Tile_X7Y1_DSP/Tile_X0Y1_FrameStrobe[10]
+ Tile_X7Y1_DSP/Tile_X0Y1_FrameStrobe[11] Tile_X7Y1_DSP/Tile_X0Y1_FrameStrobe[12]
+ Tile_X7Y1_DSP/Tile_X0Y1_FrameStrobe[13] Tile_X7Y1_DSP/Tile_X0Y1_FrameStrobe[14]
+ Tile_X7Y1_DSP/Tile_X0Y1_FrameStrobe[15] Tile_X7Y1_DSP/Tile_X0Y1_FrameStrobe[16]
+ Tile_X7Y1_DSP/Tile_X0Y1_FrameStrobe[17] Tile_X7Y1_DSP/Tile_X0Y1_FrameStrobe[18]
+ Tile_X7Y1_DSP/Tile_X0Y1_FrameStrobe[19] Tile_X7Y1_DSP/Tile_X0Y1_FrameStrobe[1] Tile_X7Y1_DSP/Tile_X0Y1_FrameStrobe[2]
+ Tile_X7Y1_DSP/Tile_X0Y1_FrameStrobe[3] Tile_X7Y1_DSP/Tile_X0Y1_FrameStrobe[4] Tile_X7Y1_DSP/Tile_X0Y1_FrameStrobe[5]
+ Tile_X7Y1_DSP/Tile_X0Y1_FrameStrobe[6] Tile_X7Y1_DSP/Tile_X0Y1_FrameStrobe[7] Tile_X7Y1_DSP/Tile_X0Y1_FrameStrobe[8]
+ Tile_X7Y1_DSP/Tile_X0Y1_FrameStrobe[9] Tile_X7Y3_DSP/Tile_X0Y0_N1BEG[0] Tile_X7Y3_DSP/Tile_X0Y0_N1BEG[1]
+ Tile_X7Y3_DSP/Tile_X0Y0_N1BEG[2] Tile_X7Y3_DSP/Tile_X0Y0_N1BEG[3] Tile_X7Y3_DSP/Tile_X0Y0_N2BEG[0]
+ Tile_X7Y3_DSP/Tile_X0Y0_N2BEG[1] Tile_X7Y3_DSP/Tile_X0Y0_N2BEG[2] Tile_X7Y3_DSP/Tile_X0Y0_N2BEG[3]
+ Tile_X7Y3_DSP/Tile_X0Y0_N2BEG[4] Tile_X7Y3_DSP/Tile_X0Y0_N2BEG[5] Tile_X7Y3_DSP/Tile_X0Y0_N2BEG[6]
+ Tile_X7Y3_DSP/Tile_X0Y0_N2BEG[7] Tile_X7Y1_DSP/Tile_X0Y1_N2END[0] Tile_X7Y1_DSP/Tile_X0Y1_N2END[1]
+ Tile_X7Y1_DSP/Tile_X0Y1_N2END[2] Tile_X7Y1_DSP/Tile_X0Y1_N2END[3] Tile_X7Y1_DSP/Tile_X0Y1_N2END[4]
+ Tile_X7Y1_DSP/Tile_X0Y1_N2END[5] Tile_X7Y1_DSP/Tile_X0Y1_N2END[6] Tile_X7Y1_DSP/Tile_X0Y1_N2END[7]
+ Tile_X7Y3_DSP/Tile_X0Y0_N4BEG[0] Tile_X7Y3_DSP/Tile_X0Y0_N4BEG[10] Tile_X7Y3_DSP/Tile_X0Y0_N4BEG[11]
+ Tile_X7Y3_DSP/Tile_X0Y0_N4BEG[12] Tile_X7Y3_DSP/Tile_X0Y0_N4BEG[13] Tile_X7Y3_DSP/Tile_X0Y0_N4BEG[14]
+ Tile_X7Y3_DSP/Tile_X0Y0_N4BEG[15] Tile_X7Y3_DSP/Tile_X0Y0_N4BEG[1] Tile_X7Y3_DSP/Tile_X0Y0_N4BEG[2]
+ Tile_X7Y3_DSP/Tile_X0Y0_N4BEG[3] Tile_X7Y3_DSP/Tile_X0Y0_N4BEG[4] Tile_X7Y3_DSP/Tile_X0Y0_N4BEG[5]
+ Tile_X7Y3_DSP/Tile_X0Y0_N4BEG[6] Tile_X7Y3_DSP/Tile_X0Y0_N4BEG[7] Tile_X7Y3_DSP/Tile_X0Y0_N4BEG[8]
+ Tile_X7Y3_DSP/Tile_X0Y0_N4BEG[9] Tile_X7Y3_DSP/Tile_X0Y0_NN4BEG[0] Tile_X7Y3_DSP/Tile_X0Y0_NN4BEG[10]
+ Tile_X7Y3_DSP/Tile_X0Y0_NN4BEG[11] Tile_X7Y3_DSP/Tile_X0Y0_NN4BEG[12] Tile_X7Y3_DSP/Tile_X0Y0_NN4BEG[13]
+ Tile_X7Y3_DSP/Tile_X0Y0_NN4BEG[14] Tile_X7Y3_DSP/Tile_X0Y0_NN4BEG[15] Tile_X7Y3_DSP/Tile_X0Y0_NN4BEG[1]
+ Tile_X7Y3_DSP/Tile_X0Y0_NN4BEG[2] Tile_X7Y3_DSP/Tile_X0Y0_NN4BEG[3] Tile_X7Y3_DSP/Tile_X0Y0_NN4BEG[4]
+ Tile_X7Y3_DSP/Tile_X0Y0_NN4BEG[5] Tile_X7Y3_DSP/Tile_X0Y0_NN4BEG[6] Tile_X7Y3_DSP/Tile_X0Y0_NN4BEG[7]
+ Tile_X7Y3_DSP/Tile_X0Y0_NN4BEG[8] Tile_X7Y3_DSP/Tile_X0Y0_NN4BEG[9] Tile_X7Y3_DSP/Tile_X0Y0_S1END[0]
+ Tile_X7Y3_DSP/Tile_X0Y0_S1END[1] Tile_X7Y3_DSP/Tile_X0Y0_S1END[2] Tile_X7Y3_DSP/Tile_X0Y0_S1END[3]
+ Tile_X7Y3_DSP/Tile_X0Y0_S2END[0] Tile_X7Y3_DSP/Tile_X0Y0_S2END[1] Tile_X7Y3_DSP/Tile_X0Y0_S2END[2]
+ Tile_X7Y3_DSP/Tile_X0Y0_S2END[3] Tile_X7Y3_DSP/Tile_X0Y0_S2END[4] Tile_X7Y3_DSP/Tile_X0Y0_S2END[5]
+ Tile_X7Y3_DSP/Tile_X0Y0_S2END[6] Tile_X7Y3_DSP/Tile_X0Y0_S2END[7] Tile_X7Y3_DSP/Tile_X0Y0_S2MID[0]
+ Tile_X7Y3_DSP/Tile_X0Y0_S2MID[1] Tile_X7Y3_DSP/Tile_X0Y0_S2MID[2] Tile_X7Y3_DSP/Tile_X0Y0_S2MID[3]
+ Tile_X7Y3_DSP/Tile_X0Y0_S2MID[4] Tile_X7Y3_DSP/Tile_X0Y0_S2MID[5] Tile_X7Y3_DSP/Tile_X0Y0_S2MID[6]
+ Tile_X7Y3_DSP/Tile_X0Y0_S2MID[7] Tile_X7Y3_DSP/Tile_X0Y0_S4END[0] Tile_X7Y3_DSP/Tile_X0Y0_S4END[10]
+ Tile_X7Y3_DSP/Tile_X0Y0_S4END[11] Tile_X7Y3_DSP/Tile_X0Y0_S4END[12] Tile_X7Y3_DSP/Tile_X0Y0_S4END[13]
+ Tile_X7Y3_DSP/Tile_X0Y0_S4END[14] Tile_X7Y3_DSP/Tile_X0Y0_S4END[15] Tile_X7Y3_DSP/Tile_X0Y0_S4END[1]
+ Tile_X7Y3_DSP/Tile_X0Y0_S4END[2] Tile_X7Y3_DSP/Tile_X0Y0_S4END[3] Tile_X7Y3_DSP/Tile_X0Y0_S4END[4]
+ Tile_X7Y3_DSP/Tile_X0Y0_S4END[5] Tile_X7Y3_DSP/Tile_X0Y0_S4END[6] Tile_X7Y3_DSP/Tile_X0Y0_S4END[7]
+ Tile_X7Y3_DSP/Tile_X0Y0_S4END[8] Tile_X7Y3_DSP/Tile_X0Y0_S4END[9] Tile_X7Y3_DSP/Tile_X0Y0_SS4END[0]
+ Tile_X7Y3_DSP/Tile_X0Y0_SS4END[10] Tile_X7Y3_DSP/Tile_X0Y0_SS4END[11] Tile_X7Y3_DSP/Tile_X0Y0_SS4END[12]
+ Tile_X7Y3_DSP/Tile_X0Y0_SS4END[13] Tile_X7Y3_DSP/Tile_X0Y0_SS4END[14] Tile_X7Y3_DSP/Tile_X0Y0_SS4END[15]
+ Tile_X7Y3_DSP/Tile_X0Y0_SS4END[1] Tile_X7Y3_DSP/Tile_X0Y0_SS4END[2] Tile_X7Y3_DSP/Tile_X0Y0_SS4END[3]
+ Tile_X7Y3_DSP/Tile_X0Y0_SS4END[4] Tile_X7Y3_DSP/Tile_X0Y0_SS4END[5] Tile_X7Y3_DSP/Tile_X0Y0_SS4END[6]
+ Tile_X7Y3_DSP/Tile_X0Y0_SS4END[7] Tile_X7Y3_DSP/Tile_X0Y0_SS4END[8] Tile_X7Y3_DSP/Tile_X0Y0_SS4END[9]
+ Tile_X7Y1_DSP/Tile_X0Y1_UserCLK Tile_X6Y3_LUT4AB/W1END[0] Tile_X6Y3_LUT4AB/W1END[1]
+ Tile_X6Y3_LUT4AB/W1END[2] Tile_X6Y3_LUT4AB/W1END[3] Tile_X8Y3_LUT4AB/W1BEG[0] Tile_X8Y3_LUT4AB/W1BEG[1]
+ Tile_X8Y3_LUT4AB/W1BEG[2] Tile_X8Y3_LUT4AB/W1BEG[3] Tile_X6Y3_LUT4AB/W2MID[0] Tile_X6Y3_LUT4AB/W2MID[1]
+ Tile_X6Y3_LUT4AB/W2MID[2] Tile_X6Y3_LUT4AB/W2MID[3] Tile_X6Y3_LUT4AB/W2MID[4] Tile_X6Y3_LUT4AB/W2MID[5]
+ Tile_X6Y3_LUT4AB/W2MID[6] Tile_X6Y3_LUT4AB/W2MID[7] Tile_X6Y3_LUT4AB/W2END[0] Tile_X6Y3_LUT4AB/W2END[1]
+ Tile_X6Y3_LUT4AB/W2END[2] Tile_X6Y3_LUT4AB/W2END[3] Tile_X6Y3_LUT4AB/W2END[4] Tile_X6Y3_LUT4AB/W2END[5]
+ Tile_X6Y3_LUT4AB/W2END[6] Tile_X6Y3_LUT4AB/W2END[7] Tile_X8Y3_LUT4AB/W2BEGb[0] Tile_X8Y3_LUT4AB/W2BEGb[1]
+ Tile_X8Y3_LUT4AB/W2BEGb[2] Tile_X8Y3_LUT4AB/W2BEGb[3] Tile_X8Y3_LUT4AB/W2BEGb[4]
+ Tile_X8Y3_LUT4AB/W2BEGb[5] Tile_X8Y3_LUT4AB/W2BEGb[6] Tile_X8Y3_LUT4AB/W2BEGb[7]
+ Tile_X8Y3_LUT4AB/W2BEG[0] Tile_X8Y3_LUT4AB/W2BEG[1] Tile_X8Y3_LUT4AB/W2BEG[2] Tile_X8Y3_LUT4AB/W2BEG[3]
+ Tile_X8Y3_LUT4AB/W2BEG[4] Tile_X8Y3_LUT4AB/W2BEG[5] Tile_X8Y3_LUT4AB/W2BEG[6] Tile_X8Y3_LUT4AB/W2BEG[7]
+ Tile_X6Y3_LUT4AB/W6END[0] Tile_X6Y3_LUT4AB/W6END[10] Tile_X6Y3_LUT4AB/W6END[11]
+ Tile_X6Y3_LUT4AB/W6END[1] Tile_X6Y3_LUT4AB/W6END[2] Tile_X6Y3_LUT4AB/W6END[3] Tile_X6Y3_LUT4AB/W6END[4]
+ Tile_X6Y3_LUT4AB/W6END[5] Tile_X6Y3_LUT4AB/W6END[6] Tile_X6Y3_LUT4AB/W6END[7] Tile_X6Y3_LUT4AB/W6END[8]
+ Tile_X6Y3_LUT4AB/W6END[9] Tile_X8Y3_LUT4AB/W6BEG[0] Tile_X8Y3_LUT4AB/W6BEG[10] Tile_X8Y3_LUT4AB/W6BEG[11]
+ Tile_X8Y3_LUT4AB/W6BEG[1] Tile_X8Y3_LUT4AB/W6BEG[2] Tile_X8Y3_LUT4AB/W6BEG[3] Tile_X8Y3_LUT4AB/W6BEG[4]
+ Tile_X8Y3_LUT4AB/W6BEG[5] Tile_X8Y3_LUT4AB/W6BEG[6] Tile_X8Y3_LUT4AB/W6BEG[7] Tile_X8Y3_LUT4AB/W6BEG[8]
+ Tile_X8Y3_LUT4AB/W6BEG[9] Tile_X6Y3_LUT4AB/WW4END[0] Tile_X6Y3_LUT4AB/WW4END[10]
+ Tile_X6Y3_LUT4AB/WW4END[11] Tile_X6Y3_LUT4AB/WW4END[12] Tile_X6Y3_LUT4AB/WW4END[13]
+ Tile_X6Y3_LUT4AB/WW4END[14] Tile_X6Y3_LUT4AB/WW4END[15] Tile_X6Y3_LUT4AB/WW4END[1]
+ Tile_X6Y3_LUT4AB/WW4END[2] Tile_X6Y3_LUT4AB/WW4END[3] Tile_X6Y3_LUT4AB/WW4END[4]
+ Tile_X6Y3_LUT4AB/WW4END[5] Tile_X6Y3_LUT4AB/WW4END[6] Tile_X6Y3_LUT4AB/WW4END[7]
+ Tile_X6Y3_LUT4AB/WW4END[8] Tile_X6Y3_LUT4AB/WW4END[9] Tile_X8Y3_LUT4AB/WW4BEG[0]
+ Tile_X8Y3_LUT4AB/WW4BEG[10] Tile_X8Y3_LUT4AB/WW4BEG[11] Tile_X8Y3_LUT4AB/WW4BEG[12]
+ Tile_X8Y3_LUT4AB/WW4BEG[13] Tile_X8Y3_LUT4AB/WW4BEG[14] Tile_X8Y3_LUT4AB/WW4BEG[15]
+ Tile_X8Y3_LUT4AB/WW4BEG[1] Tile_X8Y3_LUT4AB/WW4BEG[2] Tile_X8Y3_LUT4AB/WW4BEG[3]
+ Tile_X8Y3_LUT4AB/WW4BEG[4] Tile_X8Y3_LUT4AB/WW4BEG[5] Tile_X8Y3_LUT4AB/WW4BEG[6]
+ Tile_X8Y3_LUT4AB/WW4BEG[7] Tile_X8Y3_LUT4AB/WW4BEG[8] Tile_X8Y3_LUT4AB/WW4BEG[9]
+ Tile_X8Y4_LUT4AB/E1END[0] Tile_X8Y4_LUT4AB/E1END[1] Tile_X8Y4_LUT4AB/E1END[2] Tile_X8Y4_LUT4AB/E1END[3]
+ Tile_X6Y4_LUT4AB/E1BEG[0] Tile_X6Y4_LUT4AB/E1BEG[1] Tile_X6Y4_LUT4AB/E1BEG[2] Tile_X6Y4_LUT4AB/E1BEG[3]
+ Tile_X8Y4_LUT4AB/E2MID[0] Tile_X8Y4_LUT4AB/E2MID[1] Tile_X8Y4_LUT4AB/E2MID[2] Tile_X8Y4_LUT4AB/E2MID[3]
+ Tile_X8Y4_LUT4AB/E2MID[4] Tile_X8Y4_LUT4AB/E2MID[5] Tile_X8Y4_LUT4AB/E2MID[6] Tile_X8Y4_LUT4AB/E2MID[7]
+ Tile_X8Y4_LUT4AB/E2END[0] Tile_X8Y4_LUT4AB/E2END[1] Tile_X8Y4_LUT4AB/E2END[2] Tile_X8Y4_LUT4AB/E2END[3]
+ Tile_X8Y4_LUT4AB/E2END[4] Tile_X8Y4_LUT4AB/E2END[5] Tile_X8Y4_LUT4AB/E2END[6] Tile_X8Y4_LUT4AB/E2END[7]
+ Tile_X6Y4_LUT4AB/E2BEGb[0] Tile_X6Y4_LUT4AB/E2BEGb[1] Tile_X6Y4_LUT4AB/E2BEGb[2]
+ Tile_X6Y4_LUT4AB/E2BEGb[3] Tile_X6Y4_LUT4AB/E2BEGb[4] Tile_X6Y4_LUT4AB/E2BEGb[5]
+ Tile_X6Y4_LUT4AB/E2BEGb[6] Tile_X6Y4_LUT4AB/E2BEGb[7] Tile_X6Y4_LUT4AB/E2BEG[0]
+ Tile_X6Y4_LUT4AB/E2BEG[1] Tile_X6Y4_LUT4AB/E2BEG[2] Tile_X6Y4_LUT4AB/E2BEG[3] Tile_X6Y4_LUT4AB/E2BEG[4]
+ Tile_X6Y4_LUT4AB/E2BEG[5] Tile_X6Y4_LUT4AB/E2BEG[6] Tile_X6Y4_LUT4AB/E2BEG[7] Tile_X8Y4_LUT4AB/E6END[0]
+ Tile_X8Y4_LUT4AB/E6END[10] Tile_X8Y4_LUT4AB/E6END[11] Tile_X8Y4_LUT4AB/E6END[1]
+ Tile_X8Y4_LUT4AB/E6END[2] Tile_X8Y4_LUT4AB/E6END[3] Tile_X8Y4_LUT4AB/E6END[4] Tile_X8Y4_LUT4AB/E6END[5]
+ Tile_X8Y4_LUT4AB/E6END[6] Tile_X8Y4_LUT4AB/E6END[7] Tile_X8Y4_LUT4AB/E6END[8] Tile_X8Y4_LUT4AB/E6END[9]
+ Tile_X6Y4_LUT4AB/E6BEG[0] Tile_X6Y4_LUT4AB/E6BEG[10] Tile_X6Y4_LUT4AB/E6BEG[11]
+ Tile_X6Y4_LUT4AB/E6BEG[1] Tile_X6Y4_LUT4AB/E6BEG[2] Tile_X6Y4_LUT4AB/E6BEG[3] Tile_X6Y4_LUT4AB/E6BEG[4]
+ Tile_X6Y4_LUT4AB/E6BEG[5] Tile_X6Y4_LUT4AB/E6BEG[6] Tile_X6Y4_LUT4AB/E6BEG[7] Tile_X6Y4_LUT4AB/E6BEG[8]
+ Tile_X6Y4_LUT4AB/E6BEG[9] Tile_X8Y4_LUT4AB/EE4END[0] Tile_X8Y4_LUT4AB/EE4END[10]
+ Tile_X8Y4_LUT4AB/EE4END[11] Tile_X8Y4_LUT4AB/EE4END[12] Tile_X8Y4_LUT4AB/EE4END[13]
+ Tile_X8Y4_LUT4AB/EE4END[14] Tile_X8Y4_LUT4AB/EE4END[15] Tile_X8Y4_LUT4AB/EE4END[1]
+ Tile_X8Y4_LUT4AB/EE4END[2] Tile_X8Y4_LUT4AB/EE4END[3] Tile_X8Y4_LUT4AB/EE4END[4]
+ Tile_X8Y4_LUT4AB/EE4END[5] Tile_X8Y4_LUT4AB/EE4END[6] Tile_X8Y4_LUT4AB/EE4END[7]
+ Tile_X8Y4_LUT4AB/EE4END[8] Tile_X8Y4_LUT4AB/EE4END[9] Tile_X6Y4_LUT4AB/EE4BEG[0]
+ Tile_X6Y4_LUT4AB/EE4BEG[10] Tile_X6Y4_LUT4AB/EE4BEG[11] Tile_X6Y4_LUT4AB/EE4BEG[12]
+ Tile_X6Y4_LUT4AB/EE4BEG[13] Tile_X6Y4_LUT4AB/EE4BEG[14] Tile_X6Y4_LUT4AB/EE4BEG[15]
+ Tile_X6Y4_LUT4AB/EE4BEG[1] Tile_X6Y4_LUT4AB/EE4BEG[2] Tile_X6Y4_LUT4AB/EE4BEG[3]
+ Tile_X6Y4_LUT4AB/EE4BEG[4] Tile_X6Y4_LUT4AB/EE4BEG[5] Tile_X6Y4_LUT4AB/EE4BEG[6]
+ Tile_X6Y4_LUT4AB/EE4BEG[7] Tile_X6Y4_LUT4AB/EE4BEG[8] Tile_X6Y4_LUT4AB/EE4BEG[9]
+ Tile_X6Y4_LUT4AB/FrameData_O[0] Tile_X6Y4_LUT4AB/FrameData_O[10] Tile_X6Y4_LUT4AB/FrameData_O[11]
+ Tile_X6Y4_LUT4AB/FrameData_O[12] Tile_X6Y4_LUT4AB/FrameData_O[13] Tile_X6Y4_LUT4AB/FrameData_O[14]
+ Tile_X6Y4_LUT4AB/FrameData_O[15] Tile_X6Y4_LUT4AB/FrameData_O[16] Tile_X6Y4_LUT4AB/FrameData_O[17]
+ Tile_X6Y4_LUT4AB/FrameData_O[18] Tile_X6Y4_LUT4AB/FrameData_O[19] Tile_X6Y4_LUT4AB/FrameData_O[1]
+ Tile_X6Y4_LUT4AB/FrameData_O[20] Tile_X6Y4_LUT4AB/FrameData_O[21] Tile_X6Y4_LUT4AB/FrameData_O[22]
+ Tile_X6Y4_LUT4AB/FrameData_O[23] Tile_X6Y4_LUT4AB/FrameData_O[24] Tile_X6Y4_LUT4AB/FrameData_O[25]
+ Tile_X6Y4_LUT4AB/FrameData_O[26] Tile_X6Y4_LUT4AB/FrameData_O[27] Tile_X6Y4_LUT4AB/FrameData_O[28]
+ Tile_X6Y4_LUT4AB/FrameData_O[29] Tile_X6Y4_LUT4AB/FrameData_O[2] Tile_X6Y4_LUT4AB/FrameData_O[30]
+ Tile_X6Y4_LUT4AB/FrameData_O[31] Tile_X6Y4_LUT4AB/FrameData_O[3] Tile_X6Y4_LUT4AB/FrameData_O[4]
+ Tile_X6Y4_LUT4AB/FrameData_O[5] Tile_X6Y4_LUT4AB/FrameData_O[6] Tile_X6Y4_LUT4AB/FrameData_O[7]
+ Tile_X6Y4_LUT4AB/FrameData_O[8] Tile_X6Y4_LUT4AB/FrameData_O[9] Tile_X8Y4_LUT4AB/FrameData[0]
+ Tile_X8Y4_LUT4AB/FrameData[10] Tile_X8Y4_LUT4AB/FrameData[11] Tile_X8Y4_LUT4AB/FrameData[12]
+ Tile_X8Y4_LUT4AB/FrameData[13] Tile_X8Y4_LUT4AB/FrameData[14] Tile_X8Y4_LUT4AB/FrameData[15]
+ Tile_X8Y4_LUT4AB/FrameData[16] Tile_X8Y4_LUT4AB/FrameData[17] Tile_X8Y4_LUT4AB/FrameData[18]
+ Tile_X8Y4_LUT4AB/FrameData[19] Tile_X8Y4_LUT4AB/FrameData[1] Tile_X8Y4_LUT4AB/FrameData[20]
+ Tile_X8Y4_LUT4AB/FrameData[21] Tile_X8Y4_LUT4AB/FrameData[22] Tile_X8Y4_LUT4AB/FrameData[23]
+ Tile_X8Y4_LUT4AB/FrameData[24] Tile_X8Y4_LUT4AB/FrameData[25] Tile_X8Y4_LUT4AB/FrameData[26]
+ Tile_X8Y4_LUT4AB/FrameData[27] Tile_X8Y4_LUT4AB/FrameData[28] Tile_X8Y4_LUT4AB/FrameData[29]
+ Tile_X8Y4_LUT4AB/FrameData[2] Tile_X8Y4_LUT4AB/FrameData[30] Tile_X8Y4_LUT4AB/FrameData[31]
+ Tile_X8Y4_LUT4AB/FrameData[3] Tile_X8Y4_LUT4AB/FrameData[4] Tile_X8Y4_LUT4AB/FrameData[5]
+ Tile_X8Y4_LUT4AB/FrameData[6] Tile_X8Y4_LUT4AB/FrameData[7] Tile_X8Y4_LUT4AB/FrameData[8]
+ Tile_X8Y4_LUT4AB/FrameData[9] Tile_X7Y3_DSP/Tile_X0Y1_FrameStrobe[0] Tile_X7Y3_DSP/Tile_X0Y1_FrameStrobe[10]
+ Tile_X7Y3_DSP/Tile_X0Y1_FrameStrobe[11] Tile_X7Y3_DSP/Tile_X0Y1_FrameStrobe[12]
+ Tile_X7Y3_DSP/Tile_X0Y1_FrameStrobe[13] Tile_X7Y3_DSP/Tile_X0Y1_FrameStrobe[14]
+ Tile_X7Y3_DSP/Tile_X0Y1_FrameStrobe[15] Tile_X7Y3_DSP/Tile_X0Y1_FrameStrobe[16]
+ Tile_X7Y3_DSP/Tile_X0Y1_FrameStrobe[17] Tile_X7Y3_DSP/Tile_X0Y1_FrameStrobe[18]
+ Tile_X7Y3_DSP/Tile_X0Y1_FrameStrobe[19] Tile_X7Y3_DSP/Tile_X0Y1_FrameStrobe[1] Tile_X7Y3_DSP/Tile_X0Y1_FrameStrobe[2]
+ Tile_X7Y3_DSP/Tile_X0Y1_FrameStrobe[3] Tile_X7Y3_DSP/Tile_X0Y1_FrameStrobe[4] Tile_X7Y3_DSP/Tile_X0Y1_FrameStrobe[5]
+ Tile_X7Y3_DSP/Tile_X0Y1_FrameStrobe[6] Tile_X7Y3_DSP/Tile_X0Y1_FrameStrobe[7] Tile_X7Y3_DSP/Tile_X0Y1_FrameStrobe[8]
+ Tile_X7Y3_DSP/Tile_X0Y1_FrameStrobe[9] Tile_X7Y5_DSP/Tile_X0Y0_N1BEG[0] Tile_X7Y5_DSP/Tile_X0Y0_N1BEG[1]
+ Tile_X7Y5_DSP/Tile_X0Y0_N1BEG[2] Tile_X7Y5_DSP/Tile_X0Y0_N1BEG[3] Tile_X7Y3_DSP/Tile_X0Y1_N2END[0]
+ Tile_X7Y3_DSP/Tile_X0Y1_N2END[1] Tile_X7Y3_DSP/Tile_X0Y1_N2END[2] Tile_X7Y3_DSP/Tile_X0Y1_N2END[3]
+ Tile_X7Y3_DSP/Tile_X0Y1_N2END[4] Tile_X7Y3_DSP/Tile_X0Y1_N2END[5] Tile_X7Y3_DSP/Tile_X0Y1_N2END[6]
+ Tile_X7Y3_DSP/Tile_X0Y1_N2END[7] Tile_X7Y5_DSP/Tile_X0Y0_N2BEG[0] Tile_X7Y5_DSP/Tile_X0Y0_N2BEG[1]
+ Tile_X7Y5_DSP/Tile_X0Y0_N2BEG[2] Tile_X7Y5_DSP/Tile_X0Y0_N2BEG[3] Tile_X7Y5_DSP/Tile_X0Y0_N2BEG[4]
+ Tile_X7Y5_DSP/Tile_X0Y0_N2BEG[5] Tile_X7Y5_DSP/Tile_X0Y0_N2BEG[6] Tile_X7Y5_DSP/Tile_X0Y0_N2BEG[7]
+ Tile_X7Y5_DSP/Tile_X0Y0_N4BEG[0] Tile_X7Y5_DSP/Tile_X0Y0_N4BEG[10] Tile_X7Y5_DSP/Tile_X0Y0_N4BEG[11]
+ Tile_X7Y5_DSP/Tile_X0Y0_N4BEG[12] Tile_X7Y5_DSP/Tile_X0Y0_N4BEG[13] Tile_X7Y5_DSP/Tile_X0Y0_N4BEG[14]
+ Tile_X7Y5_DSP/Tile_X0Y0_N4BEG[15] Tile_X7Y5_DSP/Tile_X0Y0_N4BEG[1] Tile_X7Y5_DSP/Tile_X0Y0_N4BEG[2]
+ Tile_X7Y5_DSP/Tile_X0Y0_N4BEG[3] Tile_X7Y5_DSP/Tile_X0Y0_N4BEG[4] Tile_X7Y5_DSP/Tile_X0Y0_N4BEG[5]
+ Tile_X7Y5_DSP/Tile_X0Y0_N4BEG[6] Tile_X7Y5_DSP/Tile_X0Y0_N4BEG[7] Tile_X7Y5_DSP/Tile_X0Y0_N4BEG[8]
+ Tile_X7Y5_DSP/Tile_X0Y0_N4BEG[9] Tile_X7Y5_DSP/Tile_X0Y0_NN4BEG[0] Tile_X7Y5_DSP/Tile_X0Y0_NN4BEG[10]
+ Tile_X7Y5_DSP/Tile_X0Y0_NN4BEG[11] Tile_X7Y5_DSP/Tile_X0Y0_NN4BEG[12] Tile_X7Y5_DSP/Tile_X0Y0_NN4BEG[13]
+ Tile_X7Y5_DSP/Tile_X0Y0_NN4BEG[14] Tile_X7Y5_DSP/Tile_X0Y0_NN4BEG[15] Tile_X7Y5_DSP/Tile_X0Y0_NN4BEG[1]
+ Tile_X7Y5_DSP/Tile_X0Y0_NN4BEG[2] Tile_X7Y5_DSP/Tile_X0Y0_NN4BEG[3] Tile_X7Y5_DSP/Tile_X0Y0_NN4BEG[4]
+ Tile_X7Y5_DSP/Tile_X0Y0_NN4BEG[5] Tile_X7Y5_DSP/Tile_X0Y0_NN4BEG[6] Tile_X7Y5_DSP/Tile_X0Y0_NN4BEG[7]
+ Tile_X7Y5_DSP/Tile_X0Y0_NN4BEG[8] Tile_X7Y5_DSP/Tile_X0Y0_NN4BEG[9] Tile_X7Y5_DSP/Tile_X0Y0_S1END[0]
+ Tile_X7Y5_DSP/Tile_X0Y0_S1END[1] Tile_X7Y5_DSP/Tile_X0Y0_S1END[2] Tile_X7Y5_DSP/Tile_X0Y0_S1END[3]
+ Tile_X7Y5_DSP/Tile_X0Y0_S2MID[0] Tile_X7Y5_DSP/Tile_X0Y0_S2MID[1] Tile_X7Y5_DSP/Tile_X0Y0_S2MID[2]
+ Tile_X7Y5_DSP/Tile_X0Y0_S2MID[3] Tile_X7Y5_DSP/Tile_X0Y0_S2MID[4] Tile_X7Y5_DSP/Tile_X0Y0_S2MID[5]
+ Tile_X7Y5_DSP/Tile_X0Y0_S2MID[6] Tile_X7Y5_DSP/Tile_X0Y0_S2MID[7] Tile_X7Y5_DSP/Tile_X0Y0_S2END[0]
+ Tile_X7Y5_DSP/Tile_X0Y0_S2END[1] Tile_X7Y5_DSP/Tile_X0Y0_S2END[2] Tile_X7Y5_DSP/Tile_X0Y0_S2END[3]
+ Tile_X7Y5_DSP/Tile_X0Y0_S2END[4] Tile_X7Y5_DSP/Tile_X0Y0_S2END[5] Tile_X7Y5_DSP/Tile_X0Y0_S2END[6]
+ Tile_X7Y5_DSP/Tile_X0Y0_S2END[7] Tile_X7Y5_DSP/Tile_X0Y0_S4END[0] Tile_X7Y5_DSP/Tile_X0Y0_S4END[10]
+ Tile_X7Y5_DSP/Tile_X0Y0_S4END[11] Tile_X7Y5_DSP/Tile_X0Y0_S4END[12] Tile_X7Y5_DSP/Tile_X0Y0_S4END[13]
+ Tile_X7Y5_DSP/Tile_X0Y0_S4END[14] Tile_X7Y5_DSP/Tile_X0Y0_S4END[15] Tile_X7Y5_DSP/Tile_X0Y0_S4END[1]
+ Tile_X7Y5_DSP/Tile_X0Y0_S4END[2] Tile_X7Y5_DSP/Tile_X0Y0_S4END[3] Tile_X7Y5_DSP/Tile_X0Y0_S4END[4]
+ Tile_X7Y5_DSP/Tile_X0Y0_S4END[5] Tile_X7Y5_DSP/Tile_X0Y0_S4END[6] Tile_X7Y5_DSP/Tile_X0Y0_S4END[7]
+ Tile_X7Y5_DSP/Tile_X0Y0_S4END[8] Tile_X7Y5_DSP/Tile_X0Y0_S4END[9] Tile_X7Y5_DSP/Tile_X0Y0_SS4END[0]
+ Tile_X7Y5_DSP/Tile_X0Y0_SS4END[10] Tile_X7Y5_DSP/Tile_X0Y0_SS4END[11] Tile_X7Y5_DSP/Tile_X0Y0_SS4END[12]
+ Tile_X7Y5_DSP/Tile_X0Y0_SS4END[13] Tile_X7Y5_DSP/Tile_X0Y0_SS4END[14] Tile_X7Y5_DSP/Tile_X0Y0_SS4END[15]
+ Tile_X7Y5_DSP/Tile_X0Y0_SS4END[1] Tile_X7Y5_DSP/Tile_X0Y0_SS4END[2] Tile_X7Y5_DSP/Tile_X0Y0_SS4END[3]
+ Tile_X7Y5_DSP/Tile_X0Y0_SS4END[4] Tile_X7Y5_DSP/Tile_X0Y0_SS4END[5] Tile_X7Y5_DSP/Tile_X0Y0_SS4END[6]
+ Tile_X7Y5_DSP/Tile_X0Y0_SS4END[7] Tile_X7Y5_DSP/Tile_X0Y0_SS4END[8] Tile_X7Y5_DSP/Tile_X0Y0_SS4END[9]
+ Tile_X7Y3_DSP/Tile_X0Y1_UserCLK Tile_X6Y4_LUT4AB/W1END[0] Tile_X6Y4_LUT4AB/W1END[1]
+ Tile_X6Y4_LUT4AB/W1END[2] Tile_X6Y4_LUT4AB/W1END[3] Tile_X8Y4_LUT4AB/W1BEG[0] Tile_X8Y4_LUT4AB/W1BEG[1]
+ Tile_X8Y4_LUT4AB/W1BEG[2] Tile_X8Y4_LUT4AB/W1BEG[3] Tile_X6Y4_LUT4AB/W2MID[0] Tile_X6Y4_LUT4AB/W2MID[1]
+ Tile_X6Y4_LUT4AB/W2MID[2] Tile_X6Y4_LUT4AB/W2MID[3] Tile_X6Y4_LUT4AB/W2MID[4] Tile_X6Y4_LUT4AB/W2MID[5]
+ Tile_X6Y4_LUT4AB/W2MID[6] Tile_X6Y4_LUT4AB/W2MID[7] Tile_X6Y4_LUT4AB/W2END[0] Tile_X6Y4_LUT4AB/W2END[1]
+ Tile_X6Y4_LUT4AB/W2END[2] Tile_X6Y4_LUT4AB/W2END[3] Tile_X6Y4_LUT4AB/W2END[4] Tile_X6Y4_LUT4AB/W2END[5]
+ Tile_X6Y4_LUT4AB/W2END[6] Tile_X6Y4_LUT4AB/W2END[7] Tile_X8Y4_LUT4AB/W2BEGb[0] Tile_X8Y4_LUT4AB/W2BEGb[1]
+ Tile_X8Y4_LUT4AB/W2BEGb[2] Tile_X8Y4_LUT4AB/W2BEGb[3] Tile_X8Y4_LUT4AB/W2BEGb[4]
+ Tile_X8Y4_LUT4AB/W2BEGb[5] Tile_X8Y4_LUT4AB/W2BEGb[6] Tile_X8Y4_LUT4AB/W2BEGb[7]
+ Tile_X8Y4_LUT4AB/W2BEG[0] Tile_X8Y4_LUT4AB/W2BEG[1] Tile_X8Y4_LUT4AB/W2BEG[2] Tile_X8Y4_LUT4AB/W2BEG[3]
+ Tile_X8Y4_LUT4AB/W2BEG[4] Tile_X8Y4_LUT4AB/W2BEG[5] Tile_X8Y4_LUT4AB/W2BEG[6] Tile_X8Y4_LUT4AB/W2BEG[7]
+ Tile_X6Y4_LUT4AB/W6END[0] Tile_X6Y4_LUT4AB/W6END[10] Tile_X6Y4_LUT4AB/W6END[11]
+ Tile_X6Y4_LUT4AB/W6END[1] Tile_X6Y4_LUT4AB/W6END[2] Tile_X6Y4_LUT4AB/W6END[3] Tile_X6Y4_LUT4AB/W6END[4]
+ Tile_X6Y4_LUT4AB/W6END[5] Tile_X6Y4_LUT4AB/W6END[6] Tile_X6Y4_LUT4AB/W6END[7] Tile_X6Y4_LUT4AB/W6END[8]
+ Tile_X6Y4_LUT4AB/W6END[9] Tile_X8Y4_LUT4AB/W6BEG[0] Tile_X8Y4_LUT4AB/W6BEG[10] Tile_X8Y4_LUT4AB/W6BEG[11]
+ Tile_X8Y4_LUT4AB/W6BEG[1] Tile_X8Y4_LUT4AB/W6BEG[2] Tile_X8Y4_LUT4AB/W6BEG[3] Tile_X8Y4_LUT4AB/W6BEG[4]
+ Tile_X8Y4_LUT4AB/W6BEG[5] Tile_X8Y4_LUT4AB/W6BEG[6] Tile_X8Y4_LUT4AB/W6BEG[7] Tile_X8Y4_LUT4AB/W6BEG[8]
+ Tile_X8Y4_LUT4AB/W6BEG[9] Tile_X6Y4_LUT4AB/WW4END[0] Tile_X6Y4_LUT4AB/WW4END[10]
+ Tile_X6Y4_LUT4AB/WW4END[11] Tile_X6Y4_LUT4AB/WW4END[12] Tile_X6Y4_LUT4AB/WW4END[13]
+ Tile_X6Y4_LUT4AB/WW4END[14] Tile_X6Y4_LUT4AB/WW4END[15] Tile_X6Y4_LUT4AB/WW4END[1]
+ Tile_X6Y4_LUT4AB/WW4END[2] Tile_X6Y4_LUT4AB/WW4END[3] Tile_X6Y4_LUT4AB/WW4END[4]
+ Tile_X6Y4_LUT4AB/WW4END[5] Tile_X6Y4_LUT4AB/WW4END[6] Tile_X6Y4_LUT4AB/WW4END[7]
+ Tile_X6Y4_LUT4AB/WW4END[8] Tile_X6Y4_LUT4AB/WW4END[9] Tile_X8Y4_LUT4AB/WW4BEG[0]
+ Tile_X8Y4_LUT4AB/WW4BEG[10] Tile_X8Y4_LUT4AB/WW4BEG[11] Tile_X8Y4_LUT4AB/WW4BEG[12]
+ Tile_X8Y4_LUT4AB/WW4BEG[13] Tile_X8Y4_LUT4AB/WW4BEG[14] Tile_X8Y4_LUT4AB/WW4BEG[15]
+ Tile_X8Y4_LUT4AB/WW4BEG[1] Tile_X8Y4_LUT4AB/WW4BEG[2] Tile_X8Y4_LUT4AB/WW4BEG[3]
+ Tile_X8Y4_LUT4AB/WW4BEG[4] Tile_X8Y4_LUT4AB/WW4BEG[5] Tile_X8Y4_LUT4AB/WW4BEG[6]
+ Tile_X8Y4_LUT4AB/WW4BEG[7] Tile_X8Y4_LUT4AB/WW4BEG[8] Tile_X8Y4_LUT4AB/WW4BEG[9]
+ VGND VPWR DSP
XTile_X1Y3_LUT4AB Tile_X1Y4_LUT4AB/Co Tile_X1Y3_LUT4AB/Co Tile_X2Y3_LUT4AB/E1END[0]
+ Tile_X2Y3_LUT4AB/E1END[1] Tile_X2Y3_LUT4AB/E1END[2] Tile_X2Y3_LUT4AB/E1END[3] Tile_X0Y3_W_IO/E1BEG[0]
+ Tile_X0Y3_W_IO/E1BEG[1] Tile_X0Y3_W_IO/E1BEG[2] Tile_X0Y3_W_IO/E1BEG[3] Tile_X2Y3_LUT4AB/E2MID[0]
+ Tile_X2Y3_LUT4AB/E2MID[1] Tile_X2Y3_LUT4AB/E2MID[2] Tile_X2Y3_LUT4AB/E2MID[3] Tile_X2Y3_LUT4AB/E2MID[4]
+ Tile_X2Y3_LUT4AB/E2MID[5] Tile_X2Y3_LUT4AB/E2MID[6] Tile_X2Y3_LUT4AB/E2MID[7] Tile_X2Y3_LUT4AB/E2END[0]
+ Tile_X2Y3_LUT4AB/E2END[1] Tile_X2Y3_LUT4AB/E2END[2] Tile_X2Y3_LUT4AB/E2END[3] Tile_X2Y3_LUT4AB/E2END[4]
+ Tile_X2Y3_LUT4AB/E2END[5] Tile_X2Y3_LUT4AB/E2END[6] Tile_X2Y3_LUT4AB/E2END[7] Tile_X0Y3_W_IO/E2BEGb[0]
+ Tile_X0Y3_W_IO/E2BEGb[1] Tile_X0Y3_W_IO/E2BEGb[2] Tile_X0Y3_W_IO/E2BEGb[3] Tile_X0Y3_W_IO/E2BEGb[4]
+ Tile_X0Y3_W_IO/E2BEGb[5] Tile_X0Y3_W_IO/E2BEGb[6] Tile_X0Y3_W_IO/E2BEGb[7] Tile_X0Y3_W_IO/E2BEG[0]
+ Tile_X0Y3_W_IO/E2BEG[1] Tile_X0Y3_W_IO/E2BEG[2] Tile_X0Y3_W_IO/E2BEG[3] Tile_X0Y3_W_IO/E2BEG[4]
+ Tile_X0Y3_W_IO/E2BEG[5] Tile_X0Y3_W_IO/E2BEG[6] Tile_X0Y3_W_IO/E2BEG[7] Tile_X2Y3_LUT4AB/E6END[0]
+ Tile_X2Y3_LUT4AB/E6END[10] Tile_X2Y3_LUT4AB/E6END[11] Tile_X2Y3_LUT4AB/E6END[1]
+ Tile_X2Y3_LUT4AB/E6END[2] Tile_X2Y3_LUT4AB/E6END[3] Tile_X2Y3_LUT4AB/E6END[4] Tile_X2Y3_LUT4AB/E6END[5]
+ Tile_X2Y3_LUT4AB/E6END[6] Tile_X2Y3_LUT4AB/E6END[7] Tile_X2Y3_LUT4AB/E6END[8] Tile_X2Y3_LUT4AB/E6END[9]
+ Tile_X0Y3_W_IO/E6BEG[0] Tile_X0Y3_W_IO/E6BEG[10] Tile_X0Y3_W_IO/E6BEG[11] Tile_X0Y3_W_IO/E6BEG[1]
+ Tile_X0Y3_W_IO/E6BEG[2] Tile_X0Y3_W_IO/E6BEG[3] Tile_X0Y3_W_IO/E6BEG[4] Tile_X0Y3_W_IO/E6BEG[5]
+ Tile_X0Y3_W_IO/E6BEG[6] Tile_X0Y3_W_IO/E6BEG[7] Tile_X0Y3_W_IO/E6BEG[8] Tile_X0Y3_W_IO/E6BEG[9]
+ Tile_X2Y3_LUT4AB/EE4END[0] Tile_X2Y3_LUT4AB/EE4END[10] Tile_X2Y3_LUT4AB/EE4END[11]
+ Tile_X2Y3_LUT4AB/EE4END[12] Tile_X2Y3_LUT4AB/EE4END[13] Tile_X2Y3_LUT4AB/EE4END[14]
+ Tile_X2Y3_LUT4AB/EE4END[15] Tile_X2Y3_LUT4AB/EE4END[1] Tile_X2Y3_LUT4AB/EE4END[2]
+ Tile_X2Y3_LUT4AB/EE4END[3] Tile_X2Y3_LUT4AB/EE4END[4] Tile_X2Y3_LUT4AB/EE4END[5]
+ Tile_X2Y3_LUT4AB/EE4END[6] Tile_X2Y3_LUT4AB/EE4END[7] Tile_X2Y3_LUT4AB/EE4END[8]
+ Tile_X2Y3_LUT4AB/EE4END[9] Tile_X0Y3_W_IO/EE4BEG[0] Tile_X0Y3_W_IO/EE4BEG[10] Tile_X0Y3_W_IO/EE4BEG[11]
+ Tile_X0Y3_W_IO/EE4BEG[12] Tile_X0Y3_W_IO/EE4BEG[13] Tile_X0Y3_W_IO/EE4BEG[14] Tile_X0Y3_W_IO/EE4BEG[15]
+ Tile_X0Y3_W_IO/EE4BEG[1] Tile_X0Y3_W_IO/EE4BEG[2] Tile_X0Y3_W_IO/EE4BEG[3] Tile_X0Y3_W_IO/EE4BEG[4]
+ Tile_X0Y3_W_IO/EE4BEG[5] Tile_X0Y3_W_IO/EE4BEG[6] Tile_X0Y3_W_IO/EE4BEG[7] Tile_X0Y3_W_IO/EE4BEG[8]
+ Tile_X0Y3_W_IO/EE4BEG[9] Tile_X1Y3_LUT4AB/FrameData[0] Tile_X1Y3_LUT4AB/FrameData[10]
+ Tile_X1Y3_LUT4AB/FrameData[11] Tile_X1Y3_LUT4AB/FrameData[12] Tile_X1Y3_LUT4AB/FrameData[13]
+ Tile_X1Y3_LUT4AB/FrameData[14] Tile_X1Y3_LUT4AB/FrameData[15] Tile_X1Y3_LUT4AB/FrameData[16]
+ Tile_X1Y3_LUT4AB/FrameData[17] Tile_X1Y3_LUT4AB/FrameData[18] Tile_X1Y3_LUT4AB/FrameData[19]
+ Tile_X1Y3_LUT4AB/FrameData[1] Tile_X1Y3_LUT4AB/FrameData[20] Tile_X1Y3_LUT4AB/FrameData[21]
+ Tile_X1Y3_LUT4AB/FrameData[22] Tile_X1Y3_LUT4AB/FrameData[23] Tile_X1Y3_LUT4AB/FrameData[24]
+ Tile_X1Y3_LUT4AB/FrameData[25] Tile_X1Y3_LUT4AB/FrameData[26] Tile_X1Y3_LUT4AB/FrameData[27]
+ Tile_X1Y3_LUT4AB/FrameData[28] Tile_X1Y3_LUT4AB/FrameData[29] Tile_X1Y3_LUT4AB/FrameData[2]
+ Tile_X1Y3_LUT4AB/FrameData[30] Tile_X1Y3_LUT4AB/FrameData[31] Tile_X1Y3_LUT4AB/FrameData[3]
+ Tile_X1Y3_LUT4AB/FrameData[4] Tile_X1Y3_LUT4AB/FrameData[5] Tile_X1Y3_LUT4AB/FrameData[6]
+ Tile_X1Y3_LUT4AB/FrameData[7] Tile_X1Y3_LUT4AB/FrameData[8] Tile_X1Y3_LUT4AB/FrameData[9]
+ Tile_X2Y3_LUT4AB/FrameData[0] Tile_X2Y3_LUT4AB/FrameData[10] Tile_X2Y3_LUT4AB/FrameData[11]
+ Tile_X2Y3_LUT4AB/FrameData[12] Tile_X2Y3_LUT4AB/FrameData[13] Tile_X2Y3_LUT4AB/FrameData[14]
+ Tile_X2Y3_LUT4AB/FrameData[15] Tile_X2Y3_LUT4AB/FrameData[16] Tile_X2Y3_LUT4AB/FrameData[17]
+ Tile_X2Y3_LUT4AB/FrameData[18] Tile_X2Y3_LUT4AB/FrameData[19] Tile_X2Y3_LUT4AB/FrameData[1]
+ Tile_X2Y3_LUT4AB/FrameData[20] Tile_X2Y3_LUT4AB/FrameData[21] Tile_X2Y3_LUT4AB/FrameData[22]
+ Tile_X2Y3_LUT4AB/FrameData[23] Tile_X2Y3_LUT4AB/FrameData[24] Tile_X2Y3_LUT4AB/FrameData[25]
+ Tile_X2Y3_LUT4AB/FrameData[26] Tile_X2Y3_LUT4AB/FrameData[27] Tile_X2Y3_LUT4AB/FrameData[28]
+ Tile_X2Y3_LUT4AB/FrameData[29] Tile_X2Y3_LUT4AB/FrameData[2] Tile_X2Y3_LUT4AB/FrameData[30]
+ Tile_X2Y3_LUT4AB/FrameData[31] Tile_X2Y3_LUT4AB/FrameData[3] Tile_X2Y3_LUT4AB/FrameData[4]
+ Tile_X2Y3_LUT4AB/FrameData[5] Tile_X2Y3_LUT4AB/FrameData[6] Tile_X2Y3_LUT4AB/FrameData[7]
+ Tile_X2Y3_LUT4AB/FrameData[8] Tile_X2Y3_LUT4AB/FrameData[9] Tile_X1Y3_LUT4AB/FrameStrobe[0]
+ Tile_X1Y3_LUT4AB/FrameStrobe[10] Tile_X1Y3_LUT4AB/FrameStrobe[11] Tile_X1Y3_LUT4AB/FrameStrobe[12]
+ Tile_X1Y3_LUT4AB/FrameStrobe[13] Tile_X1Y3_LUT4AB/FrameStrobe[14] Tile_X1Y3_LUT4AB/FrameStrobe[15]
+ Tile_X1Y3_LUT4AB/FrameStrobe[16] Tile_X1Y3_LUT4AB/FrameStrobe[17] Tile_X1Y3_LUT4AB/FrameStrobe[18]
+ Tile_X1Y3_LUT4AB/FrameStrobe[19] Tile_X1Y3_LUT4AB/FrameStrobe[1] Tile_X1Y3_LUT4AB/FrameStrobe[2]
+ Tile_X1Y3_LUT4AB/FrameStrobe[3] Tile_X1Y3_LUT4AB/FrameStrobe[4] Tile_X1Y3_LUT4AB/FrameStrobe[5]
+ Tile_X1Y3_LUT4AB/FrameStrobe[6] Tile_X1Y3_LUT4AB/FrameStrobe[7] Tile_X1Y3_LUT4AB/FrameStrobe[8]
+ Tile_X1Y3_LUT4AB/FrameStrobe[9] Tile_X1Y2_LUT4AB/FrameStrobe[0] Tile_X1Y2_LUT4AB/FrameStrobe[10]
+ Tile_X1Y2_LUT4AB/FrameStrobe[11] Tile_X1Y2_LUT4AB/FrameStrobe[12] Tile_X1Y2_LUT4AB/FrameStrobe[13]
+ Tile_X1Y2_LUT4AB/FrameStrobe[14] Tile_X1Y2_LUT4AB/FrameStrobe[15] Tile_X1Y2_LUT4AB/FrameStrobe[16]
+ Tile_X1Y2_LUT4AB/FrameStrobe[17] Tile_X1Y2_LUT4AB/FrameStrobe[18] Tile_X1Y2_LUT4AB/FrameStrobe[19]
+ Tile_X1Y2_LUT4AB/FrameStrobe[1] Tile_X1Y2_LUT4AB/FrameStrobe[2] Tile_X1Y2_LUT4AB/FrameStrobe[3]
+ Tile_X1Y2_LUT4AB/FrameStrobe[4] Tile_X1Y2_LUT4AB/FrameStrobe[5] Tile_X1Y2_LUT4AB/FrameStrobe[6]
+ Tile_X1Y2_LUT4AB/FrameStrobe[7] Tile_X1Y2_LUT4AB/FrameStrobe[8] Tile_X1Y2_LUT4AB/FrameStrobe[9]
+ Tile_X1Y3_LUT4AB/N1BEG[0] Tile_X1Y3_LUT4AB/N1BEG[1] Tile_X1Y3_LUT4AB/N1BEG[2] Tile_X1Y3_LUT4AB/N1BEG[3]
+ Tile_X1Y4_LUT4AB/N1BEG[0] Tile_X1Y4_LUT4AB/N1BEG[1] Tile_X1Y4_LUT4AB/N1BEG[2] Tile_X1Y4_LUT4AB/N1BEG[3]
+ Tile_X1Y3_LUT4AB/N2BEG[0] Tile_X1Y3_LUT4AB/N2BEG[1] Tile_X1Y3_LUT4AB/N2BEG[2] Tile_X1Y3_LUT4AB/N2BEG[3]
+ Tile_X1Y3_LUT4AB/N2BEG[4] Tile_X1Y3_LUT4AB/N2BEG[5] Tile_X1Y3_LUT4AB/N2BEG[6] Tile_X1Y3_LUT4AB/N2BEG[7]
+ Tile_X1Y2_LUT4AB/N2END[0] Tile_X1Y2_LUT4AB/N2END[1] Tile_X1Y2_LUT4AB/N2END[2] Tile_X1Y2_LUT4AB/N2END[3]
+ Tile_X1Y2_LUT4AB/N2END[4] Tile_X1Y2_LUT4AB/N2END[5] Tile_X1Y2_LUT4AB/N2END[6] Tile_X1Y2_LUT4AB/N2END[7]
+ Tile_X1Y3_LUT4AB/N2END[0] Tile_X1Y3_LUT4AB/N2END[1] Tile_X1Y3_LUT4AB/N2END[2] Tile_X1Y3_LUT4AB/N2END[3]
+ Tile_X1Y3_LUT4AB/N2END[4] Tile_X1Y3_LUT4AB/N2END[5] Tile_X1Y3_LUT4AB/N2END[6] Tile_X1Y3_LUT4AB/N2END[7]
+ Tile_X1Y4_LUT4AB/N2BEG[0] Tile_X1Y4_LUT4AB/N2BEG[1] Tile_X1Y4_LUT4AB/N2BEG[2] Tile_X1Y4_LUT4AB/N2BEG[3]
+ Tile_X1Y4_LUT4AB/N2BEG[4] Tile_X1Y4_LUT4AB/N2BEG[5] Tile_X1Y4_LUT4AB/N2BEG[6] Tile_X1Y4_LUT4AB/N2BEG[7]
+ Tile_X1Y3_LUT4AB/N4BEG[0] Tile_X1Y3_LUT4AB/N4BEG[10] Tile_X1Y3_LUT4AB/N4BEG[11]
+ Tile_X1Y3_LUT4AB/N4BEG[12] Tile_X1Y3_LUT4AB/N4BEG[13] Tile_X1Y3_LUT4AB/N4BEG[14]
+ Tile_X1Y3_LUT4AB/N4BEG[15] Tile_X1Y3_LUT4AB/N4BEG[1] Tile_X1Y3_LUT4AB/N4BEG[2] Tile_X1Y3_LUT4AB/N4BEG[3]
+ Tile_X1Y3_LUT4AB/N4BEG[4] Tile_X1Y3_LUT4AB/N4BEG[5] Tile_X1Y3_LUT4AB/N4BEG[6] Tile_X1Y3_LUT4AB/N4BEG[7]
+ Tile_X1Y3_LUT4AB/N4BEG[8] Tile_X1Y3_LUT4AB/N4BEG[9] Tile_X1Y4_LUT4AB/N4BEG[0] Tile_X1Y4_LUT4AB/N4BEG[10]
+ Tile_X1Y4_LUT4AB/N4BEG[11] Tile_X1Y4_LUT4AB/N4BEG[12] Tile_X1Y4_LUT4AB/N4BEG[13]
+ Tile_X1Y4_LUT4AB/N4BEG[14] Tile_X1Y4_LUT4AB/N4BEG[15] Tile_X1Y4_LUT4AB/N4BEG[1]
+ Tile_X1Y4_LUT4AB/N4BEG[2] Tile_X1Y4_LUT4AB/N4BEG[3] Tile_X1Y4_LUT4AB/N4BEG[4] Tile_X1Y4_LUT4AB/N4BEG[5]
+ Tile_X1Y4_LUT4AB/N4BEG[6] Tile_X1Y4_LUT4AB/N4BEG[7] Tile_X1Y4_LUT4AB/N4BEG[8] Tile_X1Y4_LUT4AB/N4BEG[9]
+ Tile_X1Y3_LUT4AB/NN4BEG[0] Tile_X1Y3_LUT4AB/NN4BEG[10] Tile_X1Y3_LUT4AB/NN4BEG[11]
+ Tile_X1Y3_LUT4AB/NN4BEG[12] Tile_X1Y3_LUT4AB/NN4BEG[13] Tile_X1Y3_LUT4AB/NN4BEG[14]
+ Tile_X1Y3_LUT4AB/NN4BEG[15] Tile_X1Y3_LUT4AB/NN4BEG[1] Tile_X1Y3_LUT4AB/NN4BEG[2]
+ Tile_X1Y3_LUT4AB/NN4BEG[3] Tile_X1Y3_LUT4AB/NN4BEG[4] Tile_X1Y3_LUT4AB/NN4BEG[5]
+ Tile_X1Y3_LUT4AB/NN4BEG[6] Tile_X1Y3_LUT4AB/NN4BEG[7] Tile_X1Y3_LUT4AB/NN4BEG[8]
+ Tile_X1Y3_LUT4AB/NN4BEG[9] Tile_X1Y4_LUT4AB/NN4BEG[0] Tile_X1Y4_LUT4AB/NN4BEG[10]
+ Tile_X1Y4_LUT4AB/NN4BEG[11] Tile_X1Y4_LUT4AB/NN4BEG[12] Tile_X1Y4_LUT4AB/NN4BEG[13]
+ Tile_X1Y4_LUT4AB/NN4BEG[14] Tile_X1Y4_LUT4AB/NN4BEG[15] Tile_X1Y4_LUT4AB/NN4BEG[1]
+ Tile_X1Y4_LUT4AB/NN4BEG[2] Tile_X1Y4_LUT4AB/NN4BEG[3] Tile_X1Y4_LUT4AB/NN4BEG[4]
+ Tile_X1Y4_LUT4AB/NN4BEG[5] Tile_X1Y4_LUT4AB/NN4BEG[6] Tile_X1Y4_LUT4AB/NN4BEG[7]
+ Tile_X1Y4_LUT4AB/NN4BEG[8] Tile_X1Y4_LUT4AB/NN4BEG[9] Tile_X1Y4_LUT4AB/S1END[0]
+ Tile_X1Y4_LUT4AB/S1END[1] Tile_X1Y4_LUT4AB/S1END[2] Tile_X1Y4_LUT4AB/S1END[3] Tile_X1Y3_LUT4AB/S1END[0]
+ Tile_X1Y3_LUT4AB/S1END[1] Tile_X1Y3_LUT4AB/S1END[2] Tile_X1Y3_LUT4AB/S1END[3] Tile_X1Y4_LUT4AB/S2MID[0]
+ Tile_X1Y4_LUT4AB/S2MID[1] Tile_X1Y4_LUT4AB/S2MID[2] Tile_X1Y4_LUT4AB/S2MID[3] Tile_X1Y4_LUT4AB/S2MID[4]
+ Tile_X1Y4_LUT4AB/S2MID[5] Tile_X1Y4_LUT4AB/S2MID[6] Tile_X1Y4_LUT4AB/S2MID[7] Tile_X1Y4_LUT4AB/S2END[0]
+ Tile_X1Y4_LUT4AB/S2END[1] Tile_X1Y4_LUT4AB/S2END[2] Tile_X1Y4_LUT4AB/S2END[3] Tile_X1Y4_LUT4AB/S2END[4]
+ Tile_X1Y4_LUT4AB/S2END[5] Tile_X1Y4_LUT4AB/S2END[6] Tile_X1Y4_LUT4AB/S2END[7] Tile_X1Y3_LUT4AB/S2END[0]
+ Tile_X1Y3_LUT4AB/S2END[1] Tile_X1Y3_LUT4AB/S2END[2] Tile_X1Y3_LUT4AB/S2END[3] Tile_X1Y3_LUT4AB/S2END[4]
+ Tile_X1Y3_LUT4AB/S2END[5] Tile_X1Y3_LUT4AB/S2END[6] Tile_X1Y3_LUT4AB/S2END[7] Tile_X1Y3_LUT4AB/S2MID[0]
+ Tile_X1Y3_LUT4AB/S2MID[1] Tile_X1Y3_LUT4AB/S2MID[2] Tile_X1Y3_LUT4AB/S2MID[3] Tile_X1Y3_LUT4AB/S2MID[4]
+ Tile_X1Y3_LUT4AB/S2MID[5] Tile_X1Y3_LUT4AB/S2MID[6] Tile_X1Y3_LUT4AB/S2MID[7] Tile_X1Y4_LUT4AB/S4END[0]
+ Tile_X1Y4_LUT4AB/S4END[10] Tile_X1Y4_LUT4AB/S4END[11] Tile_X1Y4_LUT4AB/S4END[12]
+ Tile_X1Y4_LUT4AB/S4END[13] Tile_X1Y4_LUT4AB/S4END[14] Tile_X1Y4_LUT4AB/S4END[15]
+ Tile_X1Y4_LUT4AB/S4END[1] Tile_X1Y4_LUT4AB/S4END[2] Tile_X1Y4_LUT4AB/S4END[3] Tile_X1Y4_LUT4AB/S4END[4]
+ Tile_X1Y4_LUT4AB/S4END[5] Tile_X1Y4_LUT4AB/S4END[6] Tile_X1Y4_LUT4AB/S4END[7] Tile_X1Y4_LUT4AB/S4END[8]
+ Tile_X1Y4_LUT4AB/S4END[9] Tile_X1Y3_LUT4AB/S4END[0] Tile_X1Y3_LUT4AB/S4END[10] Tile_X1Y3_LUT4AB/S4END[11]
+ Tile_X1Y3_LUT4AB/S4END[12] Tile_X1Y3_LUT4AB/S4END[13] Tile_X1Y3_LUT4AB/S4END[14]
+ Tile_X1Y3_LUT4AB/S4END[15] Tile_X1Y3_LUT4AB/S4END[1] Tile_X1Y3_LUT4AB/S4END[2] Tile_X1Y3_LUT4AB/S4END[3]
+ Tile_X1Y3_LUT4AB/S4END[4] Tile_X1Y3_LUT4AB/S4END[5] Tile_X1Y3_LUT4AB/S4END[6] Tile_X1Y3_LUT4AB/S4END[7]
+ Tile_X1Y3_LUT4AB/S4END[8] Tile_X1Y3_LUT4AB/S4END[9] Tile_X1Y4_LUT4AB/SS4END[0] Tile_X1Y4_LUT4AB/SS4END[10]
+ Tile_X1Y4_LUT4AB/SS4END[11] Tile_X1Y4_LUT4AB/SS4END[12] Tile_X1Y4_LUT4AB/SS4END[13]
+ Tile_X1Y4_LUT4AB/SS4END[14] Tile_X1Y4_LUT4AB/SS4END[15] Tile_X1Y4_LUT4AB/SS4END[1]
+ Tile_X1Y4_LUT4AB/SS4END[2] Tile_X1Y4_LUT4AB/SS4END[3] Tile_X1Y4_LUT4AB/SS4END[4]
+ Tile_X1Y4_LUT4AB/SS4END[5] Tile_X1Y4_LUT4AB/SS4END[6] Tile_X1Y4_LUT4AB/SS4END[7]
+ Tile_X1Y4_LUT4AB/SS4END[8] Tile_X1Y4_LUT4AB/SS4END[9] Tile_X1Y3_LUT4AB/SS4END[0]
+ Tile_X1Y3_LUT4AB/SS4END[10] Tile_X1Y3_LUT4AB/SS4END[11] Tile_X1Y3_LUT4AB/SS4END[12]
+ Tile_X1Y3_LUT4AB/SS4END[13] Tile_X1Y3_LUT4AB/SS4END[14] Tile_X1Y3_LUT4AB/SS4END[15]
+ Tile_X1Y3_LUT4AB/SS4END[1] Tile_X1Y3_LUT4AB/SS4END[2] Tile_X1Y3_LUT4AB/SS4END[3]
+ Tile_X1Y3_LUT4AB/SS4END[4] Tile_X1Y3_LUT4AB/SS4END[5] Tile_X1Y3_LUT4AB/SS4END[6]
+ Tile_X1Y3_LUT4AB/SS4END[7] Tile_X1Y3_LUT4AB/SS4END[8] Tile_X1Y3_LUT4AB/SS4END[9]
+ Tile_X1Y3_LUT4AB/UserCLK Tile_X1Y2_LUT4AB/UserCLK VGND VPWR Tile_X0Y3_W_IO/W1END[0]
+ Tile_X0Y3_W_IO/W1END[1] Tile_X0Y3_W_IO/W1END[2] Tile_X0Y3_W_IO/W1END[3] Tile_X2Y3_LUT4AB/W1BEG[0]
+ Tile_X2Y3_LUT4AB/W1BEG[1] Tile_X2Y3_LUT4AB/W1BEG[2] Tile_X2Y3_LUT4AB/W1BEG[3] Tile_X0Y3_W_IO/W2MID[0]
+ Tile_X0Y3_W_IO/W2MID[1] Tile_X0Y3_W_IO/W2MID[2] Tile_X0Y3_W_IO/W2MID[3] Tile_X0Y3_W_IO/W2MID[4]
+ Tile_X0Y3_W_IO/W2MID[5] Tile_X0Y3_W_IO/W2MID[6] Tile_X0Y3_W_IO/W2MID[7] Tile_X0Y3_W_IO/W2END[0]
+ Tile_X0Y3_W_IO/W2END[1] Tile_X0Y3_W_IO/W2END[2] Tile_X0Y3_W_IO/W2END[3] Tile_X0Y3_W_IO/W2END[4]
+ Tile_X0Y3_W_IO/W2END[5] Tile_X0Y3_W_IO/W2END[6] Tile_X0Y3_W_IO/W2END[7] Tile_X1Y3_LUT4AB/W2END[0]
+ Tile_X1Y3_LUT4AB/W2END[1] Tile_X1Y3_LUT4AB/W2END[2] Tile_X1Y3_LUT4AB/W2END[3] Tile_X1Y3_LUT4AB/W2END[4]
+ Tile_X1Y3_LUT4AB/W2END[5] Tile_X1Y3_LUT4AB/W2END[6] Tile_X1Y3_LUT4AB/W2END[7] Tile_X2Y3_LUT4AB/W2BEG[0]
+ Tile_X2Y3_LUT4AB/W2BEG[1] Tile_X2Y3_LUT4AB/W2BEG[2] Tile_X2Y3_LUT4AB/W2BEG[3] Tile_X2Y3_LUT4AB/W2BEG[4]
+ Tile_X2Y3_LUT4AB/W2BEG[5] Tile_X2Y3_LUT4AB/W2BEG[6] Tile_X2Y3_LUT4AB/W2BEG[7] Tile_X0Y3_W_IO/W6END[0]
+ Tile_X0Y3_W_IO/W6END[10] Tile_X0Y3_W_IO/W6END[11] Tile_X0Y3_W_IO/W6END[1] Tile_X0Y3_W_IO/W6END[2]
+ Tile_X0Y3_W_IO/W6END[3] Tile_X0Y3_W_IO/W6END[4] Tile_X0Y3_W_IO/W6END[5] Tile_X0Y3_W_IO/W6END[6]
+ Tile_X0Y3_W_IO/W6END[7] Tile_X0Y3_W_IO/W6END[8] Tile_X0Y3_W_IO/W6END[9] Tile_X2Y3_LUT4AB/W6BEG[0]
+ Tile_X2Y3_LUT4AB/W6BEG[10] Tile_X2Y3_LUT4AB/W6BEG[11] Tile_X2Y3_LUT4AB/W6BEG[1]
+ Tile_X2Y3_LUT4AB/W6BEG[2] Tile_X2Y3_LUT4AB/W6BEG[3] Tile_X2Y3_LUT4AB/W6BEG[4] Tile_X2Y3_LUT4AB/W6BEG[5]
+ Tile_X2Y3_LUT4AB/W6BEG[6] Tile_X2Y3_LUT4AB/W6BEG[7] Tile_X2Y3_LUT4AB/W6BEG[8] Tile_X2Y3_LUT4AB/W6BEG[9]
+ Tile_X0Y3_W_IO/WW4END[0] Tile_X0Y3_W_IO/WW4END[10] Tile_X0Y3_W_IO/WW4END[11] Tile_X0Y3_W_IO/WW4END[12]
+ Tile_X0Y3_W_IO/WW4END[13] Tile_X0Y3_W_IO/WW4END[14] Tile_X0Y3_W_IO/WW4END[15] Tile_X0Y3_W_IO/WW4END[1]
+ Tile_X0Y3_W_IO/WW4END[2] Tile_X0Y3_W_IO/WW4END[3] Tile_X0Y3_W_IO/WW4END[4] Tile_X0Y3_W_IO/WW4END[5]
+ Tile_X0Y3_W_IO/WW4END[6] Tile_X0Y3_W_IO/WW4END[7] Tile_X0Y3_W_IO/WW4END[8] Tile_X0Y3_W_IO/WW4END[9]
+ Tile_X2Y3_LUT4AB/WW4BEG[0] Tile_X2Y3_LUT4AB/WW4BEG[10] Tile_X2Y3_LUT4AB/WW4BEG[11]
+ Tile_X2Y3_LUT4AB/WW4BEG[12] Tile_X2Y3_LUT4AB/WW4BEG[13] Tile_X2Y3_LUT4AB/WW4BEG[14]
+ Tile_X2Y3_LUT4AB/WW4BEG[15] Tile_X2Y3_LUT4AB/WW4BEG[1] Tile_X2Y3_LUT4AB/WW4BEG[2]
+ Tile_X2Y3_LUT4AB/WW4BEG[3] Tile_X2Y3_LUT4AB/WW4BEG[4] Tile_X2Y3_LUT4AB/WW4BEG[5]
+ Tile_X2Y3_LUT4AB/WW4BEG[6] Tile_X2Y3_LUT4AB/WW4BEG[7] Tile_X2Y3_LUT4AB/WW4BEG[8]
+ Tile_X2Y3_LUT4AB/WW4BEG[9] LUT4AB
XTile_X6Y12_LUT4AB Tile_X6Y13_LUT4AB/Co Tile_X6Y12_LUT4AB/Co Tile_X6Y12_LUT4AB/E1BEG[0]
+ Tile_X6Y12_LUT4AB/E1BEG[1] Tile_X6Y12_LUT4AB/E1BEG[2] Tile_X6Y12_LUT4AB/E1BEG[3]
+ Tile_X6Y12_LUT4AB/E1END[0] Tile_X6Y12_LUT4AB/E1END[1] Tile_X6Y12_LUT4AB/E1END[2]
+ Tile_X6Y12_LUT4AB/E1END[3] Tile_X6Y12_LUT4AB/E2BEG[0] Tile_X6Y12_LUT4AB/E2BEG[1]
+ Tile_X6Y12_LUT4AB/E2BEG[2] Tile_X6Y12_LUT4AB/E2BEG[3] Tile_X6Y12_LUT4AB/E2BEG[4]
+ Tile_X6Y12_LUT4AB/E2BEG[5] Tile_X6Y12_LUT4AB/E2BEG[6] Tile_X6Y12_LUT4AB/E2BEG[7]
+ Tile_X6Y12_LUT4AB/E2BEGb[0] Tile_X6Y12_LUT4AB/E2BEGb[1] Tile_X6Y12_LUT4AB/E2BEGb[2]
+ Tile_X6Y12_LUT4AB/E2BEGb[3] Tile_X6Y12_LUT4AB/E2BEGb[4] Tile_X6Y12_LUT4AB/E2BEGb[5]
+ Tile_X6Y12_LUT4AB/E2BEGb[6] Tile_X6Y12_LUT4AB/E2BEGb[7] Tile_X6Y12_LUT4AB/E2END[0]
+ Tile_X6Y12_LUT4AB/E2END[1] Tile_X6Y12_LUT4AB/E2END[2] Tile_X6Y12_LUT4AB/E2END[3]
+ Tile_X6Y12_LUT4AB/E2END[4] Tile_X6Y12_LUT4AB/E2END[5] Tile_X6Y12_LUT4AB/E2END[6]
+ Tile_X6Y12_LUT4AB/E2END[7] Tile_X6Y12_LUT4AB/E2MID[0] Tile_X6Y12_LUT4AB/E2MID[1]
+ Tile_X6Y12_LUT4AB/E2MID[2] Tile_X6Y12_LUT4AB/E2MID[3] Tile_X6Y12_LUT4AB/E2MID[4]
+ Tile_X6Y12_LUT4AB/E2MID[5] Tile_X6Y12_LUT4AB/E2MID[6] Tile_X6Y12_LUT4AB/E2MID[7]
+ Tile_X6Y12_LUT4AB/E6BEG[0] Tile_X6Y12_LUT4AB/E6BEG[10] Tile_X6Y12_LUT4AB/E6BEG[11]
+ Tile_X6Y12_LUT4AB/E6BEG[1] Tile_X6Y12_LUT4AB/E6BEG[2] Tile_X6Y12_LUT4AB/E6BEG[3]
+ Tile_X6Y12_LUT4AB/E6BEG[4] Tile_X6Y12_LUT4AB/E6BEG[5] Tile_X6Y12_LUT4AB/E6BEG[6]
+ Tile_X6Y12_LUT4AB/E6BEG[7] Tile_X6Y12_LUT4AB/E6BEG[8] Tile_X6Y12_LUT4AB/E6BEG[9]
+ Tile_X6Y12_LUT4AB/E6END[0] Tile_X6Y12_LUT4AB/E6END[10] Tile_X6Y12_LUT4AB/E6END[11]
+ Tile_X6Y12_LUT4AB/E6END[1] Tile_X6Y12_LUT4AB/E6END[2] Tile_X6Y12_LUT4AB/E6END[3]
+ Tile_X6Y12_LUT4AB/E6END[4] Tile_X6Y12_LUT4AB/E6END[5] Tile_X6Y12_LUT4AB/E6END[6]
+ Tile_X6Y12_LUT4AB/E6END[7] Tile_X6Y12_LUT4AB/E6END[8] Tile_X6Y12_LUT4AB/E6END[9]
+ Tile_X6Y12_LUT4AB/EE4BEG[0] Tile_X6Y12_LUT4AB/EE4BEG[10] Tile_X6Y12_LUT4AB/EE4BEG[11]
+ Tile_X6Y12_LUT4AB/EE4BEG[12] Tile_X6Y12_LUT4AB/EE4BEG[13] Tile_X6Y12_LUT4AB/EE4BEG[14]
+ Tile_X6Y12_LUT4AB/EE4BEG[15] Tile_X6Y12_LUT4AB/EE4BEG[1] Tile_X6Y12_LUT4AB/EE4BEG[2]
+ Tile_X6Y12_LUT4AB/EE4BEG[3] Tile_X6Y12_LUT4AB/EE4BEG[4] Tile_X6Y12_LUT4AB/EE4BEG[5]
+ Tile_X6Y12_LUT4AB/EE4BEG[6] Tile_X6Y12_LUT4AB/EE4BEG[7] Tile_X6Y12_LUT4AB/EE4BEG[8]
+ Tile_X6Y12_LUT4AB/EE4BEG[9] Tile_X6Y12_LUT4AB/EE4END[0] Tile_X6Y12_LUT4AB/EE4END[10]
+ Tile_X6Y12_LUT4AB/EE4END[11] Tile_X6Y12_LUT4AB/EE4END[12] Tile_X6Y12_LUT4AB/EE4END[13]
+ Tile_X6Y12_LUT4AB/EE4END[14] Tile_X6Y12_LUT4AB/EE4END[15] Tile_X6Y12_LUT4AB/EE4END[1]
+ Tile_X6Y12_LUT4AB/EE4END[2] Tile_X6Y12_LUT4AB/EE4END[3] Tile_X6Y12_LUT4AB/EE4END[4]
+ Tile_X6Y12_LUT4AB/EE4END[5] Tile_X6Y12_LUT4AB/EE4END[6] Tile_X6Y12_LUT4AB/EE4END[7]
+ Tile_X6Y12_LUT4AB/EE4END[8] Tile_X6Y12_LUT4AB/EE4END[9] Tile_X6Y12_LUT4AB/FrameData[0]
+ Tile_X6Y12_LUT4AB/FrameData[10] Tile_X6Y12_LUT4AB/FrameData[11] Tile_X6Y12_LUT4AB/FrameData[12]
+ Tile_X6Y12_LUT4AB/FrameData[13] Tile_X6Y12_LUT4AB/FrameData[14] Tile_X6Y12_LUT4AB/FrameData[15]
+ Tile_X6Y12_LUT4AB/FrameData[16] Tile_X6Y12_LUT4AB/FrameData[17] Tile_X6Y12_LUT4AB/FrameData[18]
+ Tile_X6Y12_LUT4AB/FrameData[19] Tile_X6Y12_LUT4AB/FrameData[1] Tile_X6Y12_LUT4AB/FrameData[20]
+ Tile_X6Y12_LUT4AB/FrameData[21] Tile_X6Y12_LUT4AB/FrameData[22] Tile_X6Y12_LUT4AB/FrameData[23]
+ Tile_X6Y12_LUT4AB/FrameData[24] Tile_X6Y12_LUT4AB/FrameData[25] Tile_X6Y12_LUT4AB/FrameData[26]
+ Tile_X6Y12_LUT4AB/FrameData[27] Tile_X6Y12_LUT4AB/FrameData[28] Tile_X6Y12_LUT4AB/FrameData[29]
+ Tile_X6Y12_LUT4AB/FrameData[2] Tile_X6Y12_LUT4AB/FrameData[30] Tile_X6Y12_LUT4AB/FrameData[31]
+ Tile_X6Y12_LUT4AB/FrameData[3] Tile_X6Y12_LUT4AB/FrameData[4] Tile_X6Y12_LUT4AB/FrameData[5]
+ Tile_X6Y12_LUT4AB/FrameData[6] Tile_X6Y12_LUT4AB/FrameData[7] Tile_X6Y12_LUT4AB/FrameData[8]
+ Tile_X6Y12_LUT4AB/FrameData[9] Tile_X6Y12_LUT4AB/FrameData_O[0] Tile_X6Y12_LUT4AB/FrameData_O[10]
+ Tile_X6Y12_LUT4AB/FrameData_O[11] Tile_X6Y12_LUT4AB/FrameData_O[12] Tile_X6Y12_LUT4AB/FrameData_O[13]
+ Tile_X6Y12_LUT4AB/FrameData_O[14] Tile_X6Y12_LUT4AB/FrameData_O[15] Tile_X6Y12_LUT4AB/FrameData_O[16]
+ Tile_X6Y12_LUT4AB/FrameData_O[17] Tile_X6Y12_LUT4AB/FrameData_O[18] Tile_X6Y12_LUT4AB/FrameData_O[19]
+ Tile_X6Y12_LUT4AB/FrameData_O[1] Tile_X6Y12_LUT4AB/FrameData_O[20] Tile_X6Y12_LUT4AB/FrameData_O[21]
+ Tile_X6Y12_LUT4AB/FrameData_O[22] Tile_X6Y12_LUT4AB/FrameData_O[23] Tile_X6Y12_LUT4AB/FrameData_O[24]
+ Tile_X6Y12_LUT4AB/FrameData_O[25] Tile_X6Y12_LUT4AB/FrameData_O[26] Tile_X6Y12_LUT4AB/FrameData_O[27]
+ Tile_X6Y12_LUT4AB/FrameData_O[28] Tile_X6Y12_LUT4AB/FrameData_O[29] Tile_X6Y12_LUT4AB/FrameData_O[2]
+ Tile_X6Y12_LUT4AB/FrameData_O[30] Tile_X6Y12_LUT4AB/FrameData_O[31] Tile_X6Y12_LUT4AB/FrameData_O[3]
+ Tile_X6Y12_LUT4AB/FrameData_O[4] Tile_X6Y12_LUT4AB/FrameData_O[5] Tile_X6Y12_LUT4AB/FrameData_O[6]
+ Tile_X6Y12_LUT4AB/FrameData_O[7] Tile_X6Y12_LUT4AB/FrameData_O[8] Tile_X6Y12_LUT4AB/FrameData_O[9]
+ Tile_X6Y12_LUT4AB/FrameStrobe[0] Tile_X6Y12_LUT4AB/FrameStrobe[10] Tile_X6Y12_LUT4AB/FrameStrobe[11]
+ Tile_X6Y12_LUT4AB/FrameStrobe[12] Tile_X6Y12_LUT4AB/FrameStrobe[13] Tile_X6Y12_LUT4AB/FrameStrobe[14]
+ Tile_X6Y12_LUT4AB/FrameStrobe[15] Tile_X6Y12_LUT4AB/FrameStrobe[16] Tile_X6Y12_LUT4AB/FrameStrobe[17]
+ Tile_X6Y12_LUT4AB/FrameStrobe[18] Tile_X6Y12_LUT4AB/FrameStrobe[19] Tile_X6Y12_LUT4AB/FrameStrobe[1]
+ Tile_X6Y12_LUT4AB/FrameStrobe[2] Tile_X6Y12_LUT4AB/FrameStrobe[3] Tile_X6Y12_LUT4AB/FrameStrobe[4]
+ Tile_X6Y12_LUT4AB/FrameStrobe[5] Tile_X6Y12_LUT4AB/FrameStrobe[6] Tile_X6Y12_LUT4AB/FrameStrobe[7]
+ Tile_X6Y12_LUT4AB/FrameStrobe[8] Tile_X6Y12_LUT4AB/FrameStrobe[9] Tile_X6Y11_LUT4AB/FrameStrobe[0]
+ Tile_X6Y11_LUT4AB/FrameStrobe[10] Tile_X6Y11_LUT4AB/FrameStrobe[11] Tile_X6Y11_LUT4AB/FrameStrobe[12]
+ Tile_X6Y11_LUT4AB/FrameStrobe[13] Tile_X6Y11_LUT4AB/FrameStrobe[14] Tile_X6Y11_LUT4AB/FrameStrobe[15]
+ Tile_X6Y11_LUT4AB/FrameStrobe[16] Tile_X6Y11_LUT4AB/FrameStrobe[17] Tile_X6Y11_LUT4AB/FrameStrobe[18]
+ Tile_X6Y11_LUT4AB/FrameStrobe[19] Tile_X6Y11_LUT4AB/FrameStrobe[1] Tile_X6Y11_LUT4AB/FrameStrobe[2]
+ Tile_X6Y11_LUT4AB/FrameStrobe[3] Tile_X6Y11_LUT4AB/FrameStrobe[4] Tile_X6Y11_LUT4AB/FrameStrobe[5]
+ Tile_X6Y11_LUT4AB/FrameStrobe[6] Tile_X6Y11_LUT4AB/FrameStrobe[7] Tile_X6Y11_LUT4AB/FrameStrobe[8]
+ Tile_X6Y11_LUT4AB/FrameStrobe[9] Tile_X6Y12_LUT4AB/N1BEG[0] Tile_X6Y12_LUT4AB/N1BEG[1]
+ Tile_X6Y12_LUT4AB/N1BEG[2] Tile_X6Y12_LUT4AB/N1BEG[3] Tile_X6Y13_LUT4AB/N1BEG[0]
+ Tile_X6Y13_LUT4AB/N1BEG[1] Tile_X6Y13_LUT4AB/N1BEG[2] Tile_X6Y13_LUT4AB/N1BEG[3]
+ Tile_X6Y12_LUT4AB/N2BEG[0] Tile_X6Y12_LUT4AB/N2BEG[1] Tile_X6Y12_LUT4AB/N2BEG[2]
+ Tile_X6Y12_LUT4AB/N2BEG[3] Tile_X6Y12_LUT4AB/N2BEG[4] Tile_X6Y12_LUT4AB/N2BEG[5]
+ Tile_X6Y12_LUT4AB/N2BEG[6] Tile_X6Y12_LUT4AB/N2BEG[7] Tile_X6Y11_LUT4AB/N2END[0]
+ Tile_X6Y11_LUT4AB/N2END[1] Tile_X6Y11_LUT4AB/N2END[2] Tile_X6Y11_LUT4AB/N2END[3]
+ Tile_X6Y11_LUT4AB/N2END[4] Tile_X6Y11_LUT4AB/N2END[5] Tile_X6Y11_LUT4AB/N2END[6]
+ Tile_X6Y11_LUT4AB/N2END[7] Tile_X6Y12_LUT4AB/N2END[0] Tile_X6Y12_LUT4AB/N2END[1]
+ Tile_X6Y12_LUT4AB/N2END[2] Tile_X6Y12_LUT4AB/N2END[3] Tile_X6Y12_LUT4AB/N2END[4]
+ Tile_X6Y12_LUT4AB/N2END[5] Tile_X6Y12_LUT4AB/N2END[6] Tile_X6Y12_LUT4AB/N2END[7]
+ Tile_X6Y13_LUT4AB/N2BEG[0] Tile_X6Y13_LUT4AB/N2BEG[1] Tile_X6Y13_LUT4AB/N2BEG[2]
+ Tile_X6Y13_LUT4AB/N2BEG[3] Tile_X6Y13_LUT4AB/N2BEG[4] Tile_X6Y13_LUT4AB/N2BEG[5]
+ Tile_X6Y13_LUT4AB/N2BEG[6] Tile_X6Y13_LUT4AB/N2BEG[7] Tile_X6Y12_LUT4AB/N4BEG[0]
+ Tile_X6Y12_LUT4AB/N4BEG[10] Tile_X6Y12_LUT4AB/N4BEG[11] Tile_X6Y12_LUT4AB/N4BEG[12]
+ Tile_X6Y12_LUT4AB/N4BEG[13] Tile_X6Y12_LUT4AB/N4BEG[14] Tile_X6Y12_LUT4AB/N4BEG[15]
+ Tile_X6Y12_LUT4AB/N4BEG[1] Tile_X6Y12_LUT4AB/N4BEG[2] Tile_X6Y12_LUT4AB/N4BEG[3]
+ Tile_X6Y12_LUT4AB/N4BEG[4] Tile_X6Y12_LUT4AB/N4BEG[5] Tile_X6Y12_LUT4AB/N4BEG[6]
+ Tile_X6Y12_LUT4AB/N4BEG[7] Tile_X6Y12_LUT4AB/N4BEG[8] Tile_X6Y12_LUT4AB/N4BEG[9]
+ Tile_X6Y13_LUT4AB/N4BEG[0] Tile_X6Y13_LUT4AB/N4BEG[10] Tile_X6Y13_LUT4AB/N4BEG[11]
+ Tile_X6Y13_LUT4AB/N4BEG[12] Tile_X6Y13_LUT4AB/N4BEG[13] Tile_X6Y13_LUT4AB/N4BEG[14]
+ Tile_X6Y13_LUT4AB/N4BEG[15] Tile_X6Y13_LUT4AB/N4BEG[1] Tile_X6Y13_LUT4AB/N4BEG[2]
+ Tile_X6Y13_LUT4AB/N4BEG[3] Tile_X6Y13_LUT4AB/N4BEG[4] Tile_X6Y13_LUT4AB/N4BEG[5]
+ Tile_X6Y13_LUT4AB/N4BEG[6] Tile_X6Y13_LUT4AB/N4BEG[7] Tile_X6Y13_LUT4AB/N4BEG[8]
+ Tile_X6Y13_LUT4AB/N4BEG[9] Tile_X6Y12_LUT4AB/NN4BEG[0] Tile_X6Y12_LUT4AB/NN4BEG[10]
+ Tile_X6Y12_LUT4AB/NN4BEG[11] Tile_X6Y12_LUT4AB/NN4BEG[12] Tile_X6Y12_LUT4AB/NN4BEG[13]
+ Tile_X6Y12_LUT4AB/NN4BEG[14] Tile_X6Y12_LUT4AB/NN4BEG[15] Tile_X6Y12_LUT4AB/NN4BEG[1]
+ Tile_X6Y12_LUT4AB/NN4BEG[2] Tile_X6Y12_LUT4AB/NN4BEG[3] Tile_X6Y12_LUT4AB/NN4BEG[4]
+ Tile_X6Y12_LUT4AB/NN4BEG[5] Tile_X6Y12_LUT4AB/NN4BEG[6] Tile_X6Y12_LUT4AB/NN4BEG[7]
+ Tile_X6Y12_LUT4AB/NN4BEG[8] Tile_X6Y12_LUT4AB/NN4BEG[9] Tile_X6Y13_LUT4AB/NN4BEG[0]
+ Tile_X6Y13_LUT4AB/NN4BEG[10] Tile_X6Y13_LUT4AB/NN4BEG[11] Tile_X6Y13_LUT4AB/NN4BEG[12]
+ Tile_X6Y13_LUT4AB/NN4BEG[13] Tile_X6Y13_LUT4AB/NN4BEG[14] Tile_X6Y13_LUT4AB/NN4BEG[15]
+ Tile_X6Y13_LUT4AB/NN4BEG[1] Tile_X6Y13_LUT4AB/NN4BEG[2] Tile_X6Y13_LUT4AB/NN4BEG[3]
+ Tile_X6Y13_LUT4AB/NN4BEG[4] Tile_X6Y13_LUT4AB/NN4BEG[5] Tile_X6Y13_LUT4AB/NN4BEG[6]
+ Tile_X6Y13_LUT4AB/NN4BEG[7] Tile_X6Y13_LUT4AB/NN4BEG[8] Tile_X6Y13_LUT4AB/NN4BEG[9]
+ Tile_X6Y13_LUT4AB/S1END[0] Tile_X6Y13_LUT4AB/S1END[1] Tile_X6Y13_LUT4AB/S1END[2]
+ Tile_X6Y13_LUT4AB/S1END[3] Tile_X6Y12_LUT4AB/S1END[0] Tile_X6Y12_LUT4AB/S1END[1]
+ Tile_X6Y12_LUT4AB/S1END[2] Tile_X6Y12_LUT4AB/S1END[3] Tile_X6Y13_LUT4AB/S2MID[0]
+ Tile_X6Y13_LUT4AB/S2MID[1] Tile_X6Y13_LUT4AB/S2MID[2] Tile_X6Y13_LUT4AB/S2MID[3]
+ Tile_X6Y13_LUT4AB/S2MID[4] Tile_X6Y13_LUT4AB/S2MID[5] Tile_X6Y13_LUT4AB/S2MID[6]
+ Tile_X6Y13_LUT4AB/S2MID[7] Tile_X6Y13_LUT4AB/S2END[0] Tile_X6Y13_LUT4AB/S2END[1]
+ Tile_X6Y13_LUT4AB/S2END[2] Tile_X6Y13_LUT4AB/S2END[3] Tile_X6Y13_LUT4AB/S2END[4]
+ Tile_X6Y13_LUT4AB/S2END[5] Tile_X6Y13_LUT4AB/S2END[6] Tile_X6Y13_LUT4AB/S2END[7]
+ Tile_X6Y12_LUT4AB/S2END[0] Tile_X6Y12_LUT4AB/S2END[1] Tile_X6Y12_LUT4AB/S2END[2]
+ Tile_X6Y12_LUT4AB/S2END[3] Tile_X6Y12_LUT4AB/S2END[4] Tile_X6Y12_LUT4AB/S2END[5]
+ Tile_X6Y12_LUT4AB/S2END[6] Tile_X6Y12_LUT4AB/S2END[7] Tile_X6Y12_LUT4AB/S2MID[0]
+ Tile_X6Y12_LUT4AB/S2MID[1] Tile_X6Y12_LUT4AB/S2MID[2] Tile_X6Y12_LUT4AB/S2MID[3]
+ Tile_X6Y12_LUT4AB/S2MID[4] Tile_X6Y12_LUT4AB/S2MID[5] Tile_X6Y12_LUT4AB/S2MID[6]
+ Tile_X6Y12_LUT4AB/S2MID[7] Tile_X6Y13_LUT4AB/S4END[0] Tile_X6Y13_LUT4AB/S4END[10]
+ Tile_X6Y13_LUT4AB/S4END[11] Tile_X6Y13_LUT4AB/S4END[12] Tile_X6Y13_LUT4AB/S4END[13]
+ Tile_X6Y13_LUT4AB/S4END[14] Tile_X6Y13_LUT4AB/S4END[15] Tile_X6Y13_LUT4AB/S4END[1]
+ Tile_X6Y13_LUT4AB/S4END[2] Tile_X6Y13_LUT4AB/S4END[3] Tile_X6Y13_LUT4AB/S4END[4]
+ Tile_X6Y13_LUT4AB/S4END[5] Tile_X6Y13_LUT4AB/S4END[6] Tile_X6Y13_LUT4AB/S4END[7]
+ Tile_X6Y13_LUT4AB/S4END[8] Tile_X6Y13_LUT4AB/S4END[9] Tile_X6Y12_LUT4AB/S4END[0]
+ Tile_X6Y12_LUT4AB/S4END[10] Tile_X6Y12_LUT4AB/S4END[11] Tile_X6Y12_LUT4AB/S4END[12]
+ Tile_X6Y12_LUT4AB/S4END[13] Tile_X6Y12_LUT4AB/S4END[14] Tile_X6Y12_LUT4AB/S4END[15]
+ Tile_X6Y12_LUT4AB/S4END[1] Tile_X6Y12_LUT4AB/S4END[2] Tile_X6Y12_LUT4AB/S4END[3]
+ Tile_X6Y12_LUT4AB/S4END[4] Tile_X6Y12_LUT4AB/S4END[5] Tile_X6Y12_LUT4AB/S4END[6]
+ Tile_X6Y12_LUT4AB/S4END[7] Tile_X6Y12_LUT4AB/S4END[8] Tile_X6Y12_LUT4AB/S4END[9]
+ Tile_X6Y13_LUT4AB/SS4END[0] Tile_X6Y13_LUT4AB/SS4END[10] Tile_X6Y13_LUT4AB/SS4END[11]
+ Tile_X6Y13_LUT4AB/SS4END[12] Tile_X6Y13_LUT4AB/SS4END[13] Tile_X6Y13_LUT4AB/SS4END[14]
+ Tile_X6Y13_LUT4AB/SS4END[15] Tile_X6Y13_LUT4AB/SS4END[1] Tile_X6Y13_LUT4AB/SS4END[2]
+ Tile_X6Y13_LUT4AB/SS4END[3] Tile_X6Y13_LUT4AB/SS4END[4] Tile_X6Y13_LUT4AB/SS4END[5]
+ Tile_X6Y13_LUT4AB/SS4END[6] Tile_X6Y13_LUT4AB/SS4END[7] Tile_X6Y13_LUT4AB/SS4END[8]
+ Tile_X6Y13_LUT4AB/SS4END[9] Tile_X6Y12_LUT4AB/SS4END[0] Tile_X6Y12_LUT4AB/SS4END[10]
+ Tile_X6Y12_LUT4AB/SS4END[11] Tile_X6Y12_LUT4AB/SS4END[12] Tile_X6Y12_LUT4AB/SS4END[13]
+ Tile_X6Y12_LUT4AB/SS4END[14] Tile_X6Y12_LUT4AB/SS4END[15] Tile_X6Y12_LUT4AB/SS4END[1]
+ Tile_X6Y12_LUT4AB/SS4END[2] Tile_X6Y12_LUT4AB/SS4END[3] Tile_X6Y12_LUT4AB/SS4END[4]
+ Tile_X6Y12_LUT4AB/SS4END[5] Tile_X6Y12_LUT4AB/SS4END[6] Tile_X6Y12_LUT4AB/SS4END[7]
+ Tile_X6Y12_LUT4AB/SS4END[8] Tile_X6Y12_LUT4AB/SS4END[9] Tile_X6Y12_LUT4AB/UserCLK
+ Tile_X6Y11_LUT4AB/UserCLK VGND VPWR Tile_X6Y12_LUT4AB/W1BEG[0] Tile_X6Y12_LUT4AB/W1BEG[1]
+ Tile_X6Y12_LUT4AB/W1BEG[2] Tile_X6Y12_LUT4AB/W1BEG[3] Tile_X6Y12_LUT4AB/W1END[0]
+ Tile_X6Y12_LUT4AB/W1END[1] Tile_X6Y12_LUT4AB/W1END[2] Tile_X6Y12_LUT4AB/W1END[3]
+ Tile_X6Y12_LUT4AB/W2BEG[0] Tile_X6Y12_LUT4AB/W2BEG[1] Tile_X6Y12_LUT4AB/W2BEG[2]
+ Tile_X6Y12_LUT4AB/W2BEG[3] Tile_X6Y12_LUT4AB/W2BEG[4] Tile_X6Y12_LUT4AB/W2BEG[5]
+ Tile_X6Y12_LUT4AB/W2BEG[6] Tile_X6Y12_LUT4AB/W2BEG[7] Tile_X5Y12_LUT4AB/W2END[0]
+ Tile_X5Y12_LUT4AB/W2END[1] Tile_X5Y12_LUT4AB/W2END[2] Tile_X5Y12_LUT4AB/W2END[3]
+ Tile_X5Y12_LUT4AB/W2END[4] Tile_X5Y12_LUT4AB/W2END[5] Tile_X5Y12_LUT4AB/W2END[6]
+ Tile_X5Y12_LUT4AB/W2END[7] Tile_X6Y12_LUT4AB/W2END[0] Tile_X6Y12_LUT4AB/W2END[1]
+ Tile_X6Y12_LUT4AB/W2END[2] Tile_X6Y12_LUT4AB/W2END[3] Tile_X6Y12_LUT4AB/W2END[4]
+ Tile_X6Y12_LUT4AB/W2END[5] Tile_X6Y12_LUT4AB/W2END[6] Tile_X6Y12_LUT4AB/W2END[7]
+ Tile_X6Y12_LUT4AB/W2MID[0] Tile_X6Y12_LUT4AB/W2MID[1] Tile_X6Y12_LUT4AB/W2MID[2]
+ Tile_X6Y12_LUT4AB/W2MID[3] Tile_X6Y12_LUT4AB/W2MID[4] Tile_X6Y12_LUT4AB/W2MID[5]
+ Tile_X6Y12_LUT4AB/W2MID[6] Tile_X6Y12_LUT4AB/W2MID[7] Tile_X6Y12_LUT4AB/W6BEG[0]
+ Tile_X6Y12_LUT4AB/W6BEG[10] Tile_X6Y12_LUT4AB/W6BEG[11] Tile_X6Y12_LUT4AB/W6BEG[1]
+ Tile_X6Y12_LUT4AB/W6BEG[2] Tile_X6Y12_LUT4AB/W6BEG[3] Tile_X6Y12_LUT4AB/W6BEG[4]
+ Tile_X6Y12_LUT4AB/W6BEG[5] Tile_X6Y12_LUT4AB/W6BEG[6] Tile_X6Y12_LUT4AB/W6BEG[7]
+ Tile_X6Y12_LUT4AB/W6BEG[8] Tile_X6Y12_LUT4AB/W6BEG[9] Tile_X6Y12_LUT4AB/W6END[0]
+ Tile_X6Y12_LUT4AB/W6END[10] Tile_X6Y12_LUT4AB/W6END[11] Tile_X6Y12_LUT4AB/W6END[1]
+ Tile_X6Y12_LUT4AB/W6END[2] Tile_X6Y12_LUT4AB/W6END[3] Tile_X6Y12_LUT4AB/W6END[4]
+ Tile_X6Y12_LUT4AB/W6END[5] Tile_X6Y12_LUT4AB/W6END[6] Tile_X6Y12_LUT4AB/W6END[7]
+ Tile_X6Y12_LUT4AB/W6END[8] Tile_X6Y12_LUT4AB/W6END[9] Tile_X6Y12_LUT4AB/WW4BEG[0]
+ Tile_X6Y12_LUT4AB/WW4BEG[10] Tile_X6Y12_LUT4AB/WW4BEG[11] Tile_X6Y12_LUT4AB/WW4BEG[12]
+ Tile_X6Y12_LUT4AB/WW4BEG[13] Tile_X6Y12_LUT4AB/WW4BEG[14] Tile_X6Y12_LUT4AB/WW4BEG[15]
+ Tile_X6Y12_LUT4AB/WW4BEG[1] Tile_X6Y12_LUT4AB/WW4BEG[2] Tile_X6Y12_LUT4AB/WW4BEG[3]
+ Tile_X6Y12_LUT4AB/WW4BEG[4] Tile_X6Y12_LUT4AB/WW4BEG[5] Tile_X6Y12_LUT4AB/WW4BEG[6]
+ Tile_X6Y12_LUT4AB/WW4BEG[7] Tile_X6Y12_LUT4AB/WW4BEG[8] Tile_X6Y12_LUT4AB/WW4BEG[9]
+ Tile_X6Y12_LUT4AB/WW4END[0] Tile_X6Y12_LUT4AB/WW4END[10] Tile_X6Y12_LUT4AB/WW4END[11]
+ Tile_X6Y12_LUT4AB/WW4END[12] Tile_X6Y12_LUT4AB/WW4END[13] Tile_X6Y12_LUT4AB/WW4END[14]
+ Tile_X6Y12_LUT4AB/WW4END[15] Tile_X6Y12_LUT4AB/WW4END[1] Tile_X6Y12_LUT4AB/WW4END[2]
+ Tile_X6Y12_LUT4AB/WW4END[3] Tile_X6Y12_LUT4AB/WW4END[4] Tile_X6Y12_LUT4AB/WW4END[5]
+ Tile_X6Y12_LUT4AB/WW4END[6] Tile_X6Y12_LUT4AB/WW4END[7] Tile_X6Y12_LUT4AB/WW4END[8]
+ Tile_X6Y12_LUT4AB/WW4END[9] LUT4AB
XTile_X1Y11_LUT4AB Tile_X1Y12_LUT4AB/Co Tile_X1Y11_LUT4AB/Co Tile_X2Y11_LUT4AB/E1END[0]
+ Tile_X2Y11_LUT4AB/E1END[1] Tile_X2Y11_LUT4AB/E1END[2] Tile_X2Y11_LUT4AB/E1END[3]
+ Tile_X0Y11_W_IO/E1BEG[0] Tile_X0Y11_W_IO/E1BEG[1] Tile_X0Y11_W_IO/E1BEG[2] Tile_X0Y11_W_IO/E1BEG[3]
+ Tile_X2Y11_LUT4AB/E2MID[0] Tile_X2Y11_LUT4AB/E2MID[1] Tile_X2Y11_LUT4AB/E2MID[2]
+ Tile_X2Y11_LUT4AB/E2MID[3] Tile_X2Y11_LUT4AB/E2MID[4] Tile_X2Y11_LUT4AB/E2MID[5]
+ Tile_X2Y11_LUT4AB/E2MID[6] Tile_X2Y11_LUT4AB/E2MID[7] Tile_X2Y11_LUT4AB/E2END[0]
+ Tile_X2Y11_LUT4AB/E2END[1] Tile_X2Y11_LUT4AB/E2END[2] Tile_X2Y11_LUT4AB/E2END[3]
+ Tile_X2Y11_LUT4AB/E2END[4] Tile_X2Y11_LUT4AB/E2END[5] Tile_X2Y11_LUT4AB/E2END[6]
+ Tile_X2Y11_LUT4AB/E2END[7] Tile_X0Y11_W_IO/E2BEGb[0] Tile_X0Y11_W_IO/E2BEGb[1] Tile_X0Y11_W_IO/E2BEGb[2]
+ Tile_X0Y11_W_IO/E2BEGb[3] Tile_X0Y11_W_IO/E2BEGb[4] Tile_X0Y11_W_IO/E2BEGb[5] Tile_X0Y11_W_IO/E2BEGb[6]
+ Tile_X0Y11_W_IO/E2BEGb[7] Tile_X0Y11_W_IO/E2BEG[0] Tile_X0Y11_W_IO/E2BEG[1] Tile_X0Y11_W_IO/E2BEG[2]
+ Tile_X0Y11_W_IO/E2BEG[3] Tile_X0Y11_W_IO/E2BEG[4] Tile_X0Y11_W_IO/E2BEG[5] Tile_X0Y11_W_IO/E2BEG[6]
+ Tile_X0Y11_W_IO/E2BEG[7] Tile_X2Y11_LUT4AB/E6END[0] Tile_X2Y11_LUT4AB/E6END[10]
+ Tile_X2Y11_LUT4AB/E6END[11] Tile_X2Y11_LUT4AB/E6END[1] Tile_X2Y11_LUT4AB/E6END[2]
+ Tile_X2Y11_LUT4AB/E6END[3] Tile_X2Y11_LUT4AB/E6END[4] Tile_X2Y11_LUT4AB/E6END[5]
+ Tile_X2Y11_LUT4AB/E6END[6] Tile_X2Y11_LUT4AB/E6END[7] Tile_X2Y11_LUT4AB/E6END[8]
+ Tile_X2Y11_LUT4AB/E6END[9] Tile_X0Y11_W_IO/E6BEG[0] Tile_X0Y11_W_IO/E6BEG[10] Tile_X0Y11_W_IO/E6BEG[11]
+ Tile_X0Y11_W_IO/E6BEG[1] Tile_X0Y11_W_IO/E6BEG[2] Tile_X0Y11_W_IO/E6BEG[3] Tile_X0Y11_W_IO/E6BEG[4]
+ Tile_X0Y11_W_IO/E6BEG[5] Tile_X0Y11_W_IO/E6BEG[6] Tile_X0Y11_W_IO/E6BEG[7] Tile_X0Y11_W_IO/E6BEG[8]
+ Tile_X0Y11_W_IO/E6BEG[9] Tile_X2Y11_LUT4AB/EE4END[0] Tile_X2Y11_LUT4AB/EE4END[10]
+ Tile_X2Y11_LUT4AB/EE4END[11] Tile_X2Y11_LUT4AB/EE4END[12] Tile_X2Y11_LUT4AB/EE4END[13]
+ Tile_X2Y11_LUT4AB/EE4END[14] Tile_X2Y11_LUT4AB/EE4END[15] Tile_X2Y11_LUT4AB/EE4END[1]
+ Tile_X2Y11_LUT4AB/EE4END[2] Tile_X2Y11_LUT4AB/EE4END[3] Tile_X2Y11_LUT4AB/EE4END[4]
+ Tile_X2Y11_LUT4AB/EE4END[5] Tile_X2Y11_LUT4AB/EE4END[6] Tile_X2Y11_LUT4AB/EE4END[7]
+ Tile_X2Y11_LUT4AB/EE4END[8] Tile_X2Y11_LUT4AB/EE4END[9] Tile_X0Y11_W_IO/EE4BEG[0]
+ Tile_X0Y11_W_IO/EE4BEG[10] Tile_X0Y11_W_IO/EE4BEG[11] Tile_X0Y11_W_IO/EE4BEG[12]
+ Tile_X0Y11_W_IO/EE4BEG[13] Tile_X0Y11_W_IO/EE4BEG[14] Tile_X0Y11_W_IO/EE4BEG[15]
+ Tile_X0Y11_W_IO/EE4BEG[1] Tile_X0Y11_W_IO/EE4BEG[2] Tile_X0Y11_W_IO/EE4BEG[3] Tile_X0Y11_W_IO/EE4BEG[4]
+ Tile_X0Y11_W_IO/EE4BEG[5] Tile_X0Y11_W_IO/EE4BEG[6] Tile_X0Y11_W_IO/EE4BEG[7] Tile_X0Y11_W_IO/EE4BEG[8]
+ Tile_X0Y11_W_IO/EE4BEG[9] Tile_X1Y11_LUT4AB/FrameData[0] Tile_X1Y11_LUT4AB/FrameData[10]
+ Tile_X1Y11_LUT4AB/FrameData[11] Tile_X1Y11_LUT4AB/FrameData[12] Tile_X1Y11_LUT4AB/FrameData[13]
+ Tile_X1Y11_LUT4AB/FrameData[14] Tile_X1Y11_LUT4AB/FrameData[15] Tile_X1Y11_LUT4AB/FrameData[16]
+ Tile_X1Y11_LUT4AB/FrameData[17] Tile_X1Y11_LUT4AB/FrameData[18] Tile_X1Y11_LUT4AB/FrameData[19]
+ Tile_X1Y11_LUT4AB/FrameData[1] Tile_X1Y11_LUT4AB/FrameData[20] Tile_X1Y11_LUT4AB/FrameData[21]
+ Tile_X1Y11_LUT4AB/FrameData[22] Tile_X1Y11_LUT4AB/FrameData[23] Tile_X1Y11_LUT4AB/FrameData[24]
+ Tile_X1Y11_LUT4AB/FrameData[25] Tile_X1Y11_LUT4AB/FrameData[26] Tile_X1Y11_LUT4AB/FrameData[27]
+ Tile_X1Y11_LUT4AB/FrameData[28] Tile_X1Y11_LUT4AB/FrameData[29] Tile_X1Y11_LUT4AB/FrameData[2]
+ Tile_X1Y11_LUT4AB/FrameData[30] Tile_X1Y11_LUT4AB/FrameData[31] Tile_X1Y11_LUT4AB/FrameData[3]
+ Tile_X1Y11_LUT4AB/FrameData[4] Tile_X1Y11_LUT4AB/FrameData[5] Tile_X1Y11_LUT4AB/FrameData[6]
+ Tile_X1Y11_LUT4AB/FrameData[7] Tile_X1Y11_LUT4AB/FrameData[8] Tile_X1Y11_LUT4AB/FrameData[9]
+ Tile_X2Y11_LUT4AB/FrameData[0] Tile_X2Y11_LUT4AB/FrameData[10] Tile_X2Y11_LUT4AB/FrameData[11]
+ Tile_X2Y11_LUT4AB/FrameData[12] Tile_X2Y11_LUT4AB/FrameData[13] Tile_X2Y11_LUT4AB/FrameData[14]
+ Tile_X2Y11_LUT4AB/FrameData[15] Tile_X2Y11_LUT4AB/FrameData[16] Tile_X2Y11_LUT4AB/FrameData[17]
+ Tile_X2Y11_LUT4AB/FrameData[18] Tile_X2Y11_LUT4AB/FrameData[19] Tile_X2Y11_LUT4AB/FrameData[1]
+ Tile_X2Y11_LUT4AB/FrameData[20] Tile_X2Y11_LUT4AB/FrameData[21] Tile_X2Y11_LUT4AB/FrameData[22]
+ Tile_X2Y11_LUT4AB/FrameData[23] Tile_X2Y11_LUT4AB/FrameData[24] Tile_X2Y11_LUT4AB/FrameData[25]
+ Tile_X2Y11_LUT4AB/FrameData[26] Tile_X2Y11_LUT4AB/FrameData[27] Tile_X2Y11_LUT4AB/FrameData[28]
+ Tile_X2Y11_LUT4AB/FrameData[29] Tile_X2Y11_LUT4AB/FrameData[2] Tile_X2Y11_LUT4AB/FrameData[30]
+ Tile_X2Y11_LUT4AB/FrameData[31] Tile_X2Y11_LUT4AB/FrameData[3] Tile_X2Y11_LUT4AB/FrameData[4]
+ Tile_X2Y11_LUT4AB/FrameData[5] Tile_X2Y11_LUT4AB/FrameData[6] Tile_X2Y11_LUT4AB/FrameData[7]
+ Tile_X2Y11_LUT4AB/FrameData[8] Tile_X2Y11_LUT4AB/FrameData[9] Tile_X1Y11_LUT4AB/FrameStrobe[0]
+ Tile_X1Y11_LUT4AB/FrameStrobe[10] Tile_X1Y11_LUT4AB/FrameStrobe[11] Tile_X1Y11_LUT4AB/FrameStrobe[12]
+ Tile_X1Y11_LUT4AB/FrameStrobe[13] Tile_X1Y11_LUT4AB/FrameStrobe[14] Tile_X1Y11_LUT4AB/FrameStrobe[15]
+ Tile_X1Y11_LUT4AB/FrameStrobe[16] Tile_X1Y11_LUT4AB/FrameStrobe[17] Tile_X1Y11_LUT4AB/FrameStrobe[18]
+ Tile_X1Y11_LUT4AB/FrameStrobe[19] Tile_X1Y11_LUT4AB/FrameStrobe[1] Tile_X1Y11_LUT4AB/FrameStrobe[2]
+ Tile_X1Y11_LUT4AB/FrameStrobe[3] Tile_X1Y11_LUT4AB/FrameStrobe[4] Tile_X1Y11_LUT4AB/FrameStrobe[5]
+ Tile_X1Y11_LUT4AB/FrameStrobe[6] Tile_X1Y11_LUT4AB/FrameStrobe[7] Tile_X1Y11_LUT4AB/FrameStrobe[8]
+ Tile_X1Y11_LUT4AB/FrameStrobe[9] Tile_X1Y10_LUT4AB/FrameStrobe[0] Tile_X1Y10_LUT4AB/FrameStrobe[10]
+ Tile_X1Y10_LUT4AB/FrameStrobe[11] Tile_X1Y10_LUT4AB/FrameStrobe[12] Tile_X1Y10_LUT4AB/FrameStrobe[13]
+ Tile_X1Y10_LUT4AB/FrameStrobe[14] Tile_X1Y10_LUT4AB/FrameStrobe[15] Tile_X1Y10_LUT4AB/FrameStrobe[16]
+ Tile_X1Y10_LUT4AB/FrameStrobe[17] Tile_X1Y10_LUT4AB/FrameStrobe[18] Tile_X1Y10_LUT4AB/FrameStrobe[19]
+ Tile_X1Y10_LUT4AB/FrameStrobe[1] Tile_X1Y10_LUT4AB/FrameStrobe[2] Tile_X1Y10_LUT4AB/FrameStrobe[3]
+ Tile_X1Y10_LUT4AB/FrameStrobe[4] Tile_X1Y10_LUT4AB/FrameStrobe[5] Tile_X1Y10_LUT4AB/FrameStrobe[6]
+ Tile_X1Y10_LUT4AB/FrameStrobe[7] Tile_X1Y10_LUT4AB/FrameStrobe[8] Tile_X1Y10_LUT4AB/FrameStrobe[9]
+ Tile_X1Y11_LUT4AB/N1BEG[0] Tile_X1Y11_LUT4AB/N1BEG[1] Tile_X1Y11_LUT4AB/N1BEG[2]
+ Tile_X1Y11_LUT4AB/N1BEG[3] Tile_X1Y12_LUT4AB/N1BEG[0] Tile_X1Y12_LUT4AB/N1BEG[1]
+ Tile_X1Y12_LUT4AB/N1BEG[2] Tile_X1Y12_LUT4AB/N1BEG[3] Tile_X1Y11_LUT4AB/N2BEG[0]
+ Tile_X1Y11_LUT4AB/N2BEG[1] Tile_X1Y11_LUT4AB/N2BEG[2] Tile_X1Y11_LUT4AB/N2BEG[3]
+ Tile_X1Y11_LUT4AB/N2BEG[4] Tile_X1Y11_LUT4AB/N2BEG[5] Tile_X1Y11_LUT4AB/N2BEG[6]
+ Tile_X1Y11_LUT4AB/N2BEG[7] Tile_X1Y10_LUT4AB/N2END[0] Tile_X1Y10_LUT4AB/N2END[1]
+ Tile_X1Y10_LUT4AB/N2END[2] Tile_X1Y10_LUT4AB/N2END[3] Tile_X1Y10_LUT4AB/N2END[4]
+ Tile_X1Y10_LUT4AB/N2END[5] Tile_X1Y10_LUT4AB/N2END[6] Tile_X1Y10_LUT4AB/N2END[7]
+ Tile_X1Y11_LUT4AB/N2END[0] Tile_X1Y11_LUT4AB/N2END[1] Tile_X1Y11_LUT4AB/N2END[2]
+ Tile_X1Y11_LUT4AB/N2END[3] Tile_X1Y11_LUT4AB/N2END[4] Tile_X1Y11_LUT4AB/N2END[5]
+ Tile_X1Y11_LUT4AB/N2END[6] Tile_X1Y11_LUT4AB/N2END[7] Tile_X1Y12_LUT4AB/N2BEG[0]
+ Tile_X1Y12_LUT4AB/N2BEG[1] Tile_X1Y12_LUT4AB/N2BEG[2] Tile_X1Y12_LUT4AB/N2BEG[3]
+ Tile_X1Y12_LUT4AB/N2BEG[4] Tile_X1Y12_LUT4AB/N2BEG[5] Tile_X1Y12_LUT4AB/N2BEG[6]
+ Tile_X1Y12_LUT4AB/N2BEG[7] Tile_X1Y11_LUT4AB/N4BEG[0] Tile_X1Y11_LUT4AB/N4BEG[10]
+ Tile_X1Y11_LUT4AB/N4BEG[11] Tile_X1Y11_LUT4AB/N4BEG[12] Tile_X1Y11_LUT4AB/N4BEG[13]
+ Tile_X1Y11_LUT4AB/N4BEG[14] Tile_X1Y11_LUT4AB/N4BEG[15] Tile_X1Y11_LUT4AB/N4BEG[1]
+ Tile_X1Y11_LUT4AB/N4BEG[2] Tile_X1Y11_LUT4AB/N4BEG[3] Tile_X1Y11_LUT4AB/N4BEG[4]
+ Tile_X1Y11_LUT4AB/N4BEG[5] Tile_X1Y11_LUT4AB/N4BEG[6] Tile_X1Y11_LUT4AB/N4BEG[7]
+ Tile_X1Y11_LUT4AB/N4BEG[8] Tile_X1Y11_LUT4AB/N4BEG[9] Tile_X1Y12_LUT4AB/N4BEG[0]
+ Tile_X1Y12_LUT4AB/N4BEG[10] Tile_X1Y12_LUT4AB/N4BEG[11] Tile_X1Y12_LUT4AB/N4BEG[12]
+ Tile_X1Y12_LUT4AB/N4BEG[13] Tile_X1Y12_LUT4AB/N4BEG[14] Tile_X1Y12_LUT4AB/N4BEG[15]
+ Tile_X1Y12_LUT4AB/N4BEG[1] Tile_X1Y12_LUT4AB/N4BEG[2] Tile_X1Y12_LUT4AB/N4BEG[3]
+ Tile_X1Y12_LUT4AB/N4BEG[4] Tile_X1Y12_LUT4AB/N4BEG[5] Tile_X1Y12_LUT4AB/N4BEG[6]
+ Tile_X1Y12_LUT4AB/N4BEG[7] Tile_X1Y12_LUT4AB/N4BEG[8] Tile_X1Y12_LUT4AB/N4BEG[9]
+ Tile_X1Y11_LUT4AB/NN4BEG[0] Tile_X1Y11_LUT4AB/NN4BEG[10] Tile_X1Y11_LUT4AB/NN4BEG[11]
+ Tile_X1Y11_LUT4AB/NN4BEG[12] Tile_X1Y11_LUT4AB/NN4BEG[13] Tile_X1Y11_LUT4AB/NN4BEG[14]
+ Tile_X1Y11_LUT4AB/NN4BEG[15] Tile_X1Y11_LUT4AB/NN4BEG[1] Tile_X1Y11_LUT4AB/NN4BEG[2]
+ Tile_X1Y11_LUT4AB/NN4BEG[3] Tile_X1Y11_LUT4AB/NN4BEG[4] Tile_X1Y11_LUT4AB/NN4BEG[5]
+ Tile_X1Y11_LUT4AB/NN4BEG[6] Tile_X1Y11_LUT4AB/NN4BEG[7] Tile_X1Y11_LUT4AB/NN4BEG[8]
+ Tile_X1Y11_LUT4AB/NN4BEG[9] Tile_X1Y12_LUT4AB/NN4BEG[0] Tile_X1Y12_LUT4AB/NN4BEG[10]
+ Tile_X1Y12_LUT4AB/NN4BEG[11] Tile_X1Y12_LUT4AB/NN4BEG[12] Tile_X1Y12_LUT4AB/NN4BEG[13]
+ Tile_X1Y12_LUT4AB/NN4BEG[14] Tile_X1Y12_LUT4AB/NN4BEG[15] Tile_X1Y12_LUT4AB/NN4BEG[1]
+ Tile_X1Y12_LUT4AB/NN4BEG[2] Tile_X1Y12_LUT4AB/NN4BEG[3] Tile_X1Y12_LUT4AB/NN4BEG[4]
+ Tile_X1Y12_LUT4AB/NN4BEG[5] Tile_X1Y12_LUT4AB/NN4BEG[6] Tile_X1Y12_LUT4AB/NN4BEG[7]
+ Tile_X1Y12_LUT4AB/NN4BEG[8] Tile_X1Y12_LUT4AB/NN4BEG[9] Tile_X1Y12_LUT4AB/S1END[0]
+ Tile_X1Y12_LUT4AB/S1END[1] Tile_X1Y12_LUT4AB/S1END[2] Tile_X1Y12_LUT4AB/S1END[3]
+ Tile_X1Y11_LUT4AB/S1END[0] Tile_X1Y11_LUT4AB/S1END[1] Tile_X1Y11_LUT4AB/S1END[2]
+ Tile_X1Y11_LUT4AB/S1END[3] Tile_X1Y12_LUT4AB/S2MID[0] Tile_X1Y12_LUT4AB/S2MID[1]
+ Tile_X1Y12_LUT4AB/S2MID[2] Tile_X1Y12_LUT4AB/S2MID[3] Tile_X1Y12_LUT4AB/S2MID[4]
+ Tile_X1Y12_LUT4AB/S2MID[5] Tile_X1Y12_LUT4AB/S2MID[6] Tile_X1Y12_LUT4AB/S2MID[7]
+ Tile_X1Y12_LUT4AB/S2END[0] Tile_X1Y12_LUT4AB/S2END[1] Tile_X1Y12_LUT4AB/S2END[2]
+ Tile_X1Y12_LUT4AB/S2END[3] Tile_X1Y12_LUT4AB/S2END[4] Tile_X1Y12_LUT4AB/S2END[5]
+ Tile_X1Y12_LUT4AB/S2END[6] Tile_X1Y12_LUT4AB/S2END[7] Tile_X1Y11_LUT4AB/S2END[0]
+ Tile_X1Y11_LUT4AB/S2END[1] Tile_X1Y11_LUT4AB/S2END[2] Tile_X1Y11_LUT4AB/S2END[3]
+ Tile_X1Y11_LUT4AB/S2END[4] Tile_X1Y11_LUT4AB/S2END[5] Tile_X1Y11_LUT4AB/S2END[6]
+ Tile_X1Y11_LUT4AB/S2END[7] Tile_X1Y11_LUT4AB/S2MID[0] Tile_X1Y11_LUT4AB/S2MID[1]
+ Tile_X1Y11_LUT4AB/S2MID[2] Tile_X1Y11_LUT4AB/S2MID[3] Tile_X1Y11_LUT4AB/S2MID[4]
+ Tile_X1Y11_LUT4AB/S2MID[5] Tile_X1Y11_LUT4AB/S2MID[6] Tile_X1Y11_LUT4AB/S2MID[7]
+ Tile_X1Y12_LUT4AB/S4END[0] Tile_X1Y12_LUT4AB/S4END[10] Tile_X1Y12_LUT4AB/S4END[11]
+ Tile_X1Y12_LUT4AB/S4END[12] Tile_X1Y12_LUT4AB/S4END[13] Tile_X1Y12_LUT4AB/S4END[14]
+ Tile_X1Y12_LUT4AB/S4END[15] Tile_X1Y12_LUT4AB/S4END[1] Tile_X1Y12_LUT4AB/S4END[2]
+ Tile_X1Y12_LUT4AB/S4END[3] Tile_X1Y12_LUT4AB/S4END[4] Tile_X1Y12_LUT4AB/S4END[5]
+ Tile_X1Y12_LUT4AB/S4END[6] Tile_X1Y12_LUT4AB/S4END[7] Tile_X1Y12_LUT4AB/S4END[8]
+ Tile_X1Y12_LUT4AB/S4END[9] Tile_X1Y11_LUT4AB/S4END[0] Tile_X1Y11_LUT4AB/S4END[10]
+ Tile_X1Y11_LUT4AB/S4END[11] Tile_X1Y11_LUT4AB/S4END[12] Tile_X1Y11_LUT4AB/S4END[13]
+ Tile_X1Y11_LUT4AB/S4END[14] Tile_X1Y11_LUT4AB/S4END[15] Tile_X1Y11_LUT4AB/S4END[1]
+ Tile_X1Y11_LUT4AB/S4END[2] Tile_X1Y11_LUT4AB/S4END[3] Tile_X1Y11_LUT4AB/S4END[4]
+ Tile_X1Y11_LUT4AB/S4END[5] Tile_X1Y11_LUT4AB/S4END[6] Tile_X1Y11_LUT4AB/S4END[7]
+ Tile_X1Y11_LUT4AB/S4END[8] Tile_X1Y11_LUT4AB/S4END[9] Tile_X1Y12_LUT4AB/SS4END[0]
+ Tile_X1Y12_LUT4AB/SS4END[10] Tile_X1Y12_LUT4AB/SS4END[11] Tile_X1Y12_LUT4AB/SS4END[12]
+ Tile_X1Y12_LUT4AB/SS4END[13] Tile_X1Y12_LUT4AB/SS4END[14] Tile_X1Y12_LUT4AB/SS4END[15]
+ Tile_X1Y12_LUT4AB/SS4END[1] Tile_X1Y12_LUT4AB/SS4END[2] Tile_X1Y12_LUT4AB/SS4END[3]
+ Tile_X1Y12_LUT4AB/SS4END[4] Tile_X1Y12_LUT4AB/SS4END[5] Tile_X1Y12_LUT4AB/SS4END[6]
+ Tile_X1Y12_LUT4AB/SS4END[7] Tile_X1Y12_LUT4AB/SS4END[8] Tile_X1Y12_LUT4AB/SS4END[9]
+ Tile_X1Y11_LUT4AB/SS4END[0] Tile_X1Y11_LUT4AB/SS4END[10] Tile_X1Y11_LUT4AB/SS4END[11]
+ Tile_X1Y11_LUT4AB/SS4END[12] Tile_X1Y11_LUT4AB/SS4END[13] Tile_X1Y11_LUT4AB/SS4END[14]
+ Tile_X1Y11_LUT4AB/SS4END[15] Tile_X1Y11_LUT4AB/SS4END[1] Tile_X1Y11_LUT4AB/SS4END[2]
+ Tile_X1Y11_LUT4AB/SS4END[3] Tile_X1Y11_LUT4AB/SS4END[4] Tile_X1Y11_LUT4AB/SS4END[5]
+ Tile_X1Y11_LUT4AB/SS4END[6] Tile_X1Y11_LUT4AB/SS4END[7] Tile_X1Y11_LUT4AB/SS4END[8]
+ Tile_X1Y11_LUT4AB/SS4END[9] Tile_X1Y11_LUT4AB/UserCLK Tile_X1Y10_LUT4AB/UserCLK
+ VGND VPWR Tile_X0Y11_W_IO/W1END[0] Tile_X0Y11_W_IO/W1END[1] Tile_X0Y11_W_IO/W1END[2]
+ Tile_X0Y11_W_IO/W1END[3] Tile_X2Y11_LUT4AB/W1BEG[0] Tile_X2Y11_LUT4AB/W1BEG[1] Tile_X2Y11_LUT4AB/W1BEG[2]
+ Tile_X2Y11_LUT4AB/W1BEG[3] Tile_X0Y11_W_IO/W2MID[0] Tile_X0Y11_W_IO/W2MID[1] Tile_X0Y11_W_IO/W2MID[2]
+ Tile_X0Y11_W_IO/W2MID[3] Tile_X0Y11_W_IO/W2MID[4] Tile_X0Y11_W_IO/W2MID[5] Tile_X0Y11_W_IO/W2MID[6]
+ Tile_X0Y11_W_IO/W2MID[7] Tile_X0Y11_W_IO/W2END[0] Tile_X0Y11_W_IO/W2END[1] Tile_X0Y11_W_IO/W2END[2]
+ Tile_X0Y11_W_IO/W2END[3] Tile_X0Y11_W_IO/W2END[4] Tile_X0Y11_W_IO/W2END[5] Tile_X0Y11_W_IO/W2END[6]
+ Tile_X0Y11_W_IO/W2END[7] Tile_X1Y11_LUT4AB/W2END[0] Tile_X1Y11_LUT4AB/W2END[1] Tile_X1Y11_LUT4AB/W2END[2]
+ Tile_X1Y11_LUT4AB/W2END[3] Tile_X1Y11_LUT4AB/W2END[4] Tile_X1Y11_LUT4AB/W2END[5]
+ Tile_X1Y11_LUT4AB/W2END[6] Tile_X1Y11_LUT4AB/W2END[7] Tile_X2Y11_LUT4AB/W2BEG[0]
+ Tile_X2Y11_LUT4AB/W2BEG[1] Tile_X2Y11_LUT4AB/W2BEG[2] Tile_X2Y11_LUT4AB/W2BEG[3]
+ Tile_X2Y11_LUT4AB/W2BEG[4] Tile_X2Y11_LUT4AB/W2BEG[5] Tile_X2Y11_LUT4AB/W2BEG[6]
+ Tile_X2Y11_LUT4AB/W2BEG[7] Tile_X0Y11_W_IO/W6END[0] Tile_X0Y11_W_IO/W6END[10] Tile_X0Y11_W_IO/W6END[11]
+ Tile_X0Y11_W_IO/W6END[1] Tile_X0Y11_W_IO/W6END[2] Tile_X0Y11_W_IO/W6END[3] Tile_X0Y11_W_IO/W6END[4]
+ Tile_X0Y11_W_IO/W6END[5] Tile_X0Y11_W_IO/W6END[6] Tile_X0Y11_W_IO/W6END[7] Tile_X0Y11_W_IO/W6END[8]
+ Tile_X0Y11_W_IO/W6END[9] Tile_X2Y11_LUT4AB/W6BEG[0] Tile_X2Y11_LUT4AB/W6BEG[10]
+ Tile_X2Y11_LUT4AB/W6BEG[11] Tile_X2Y11_LUT4AB/W6BEG[1] Tile_X2Y11_LUT4AB/W6BEG[2]
+ Tile_X2Y11_LUT4AB/W6BEG[3] Tile_X2Y11_LUT4AB/W6BEG[4] Tile_X2Y11_LUT4AB/W6BEG[5]
+ Tile_X2Y11_LUT4AB/W6BEG[6] Tile_X2Y11_LUT4AB/W6BEG[7] Tile_X2Y11_LUT4AB/W6BEG[8]
+ Tile_X2Y11_LUT4AB/W6BEG[9] Tile_X0Y11_W_IO/WW4END[0] Tile_X0Y11_W_IO/WW4END[10]
+ Tile_X0Y11_W_IO/WW4END[11] Tile_X0Y11_W_IO/WW4END[12] Tile_X0Y11_W_IO/WW4END[13]
+ Tile_X0Y11_W_IO/WW4END[14] Tile_X0Y11_W_IO/WW4END[15] Tile_X0Y11_W_IO/WW4END[1]
+ Tile_X0Y11_W_IO/WW4END[2] Tile_X0Y11_W_IO/WW4END[3] Tile_X0Y11_W_IO/WW4END[4] Tile_X0Y11_W_IO/WW4END[5]
+ Tile_X0Y11_W_IO/WW4END[6] Tile_X0Y11_W_IO/WW4END[7] Tile_X0Y11_W_IO/WW4END[8] Tile_X0Y11_W_IO/WW4END[9]
+ Tile_X2Y11_LUT4AB/WW4BEG[0] Tile_X2Y11_LUT4AB/WW4BEG[10] Tile_X2Y11_LUT4AB/WW4BEG[11]
+ Tile_X2Y11_LUT4AB/WW4BEG[12] Tile_X2Y11_LUT4AB/WW4BEG[13] Tile_X2Y11_LUT4AB/WW4BEG[14]
+ Tile_X2Y11_LUT4AB/WW4BEG[15] Tile_X2Y11_LUT4AB/WW4BEG[1] Tile_X2Y11_LUT4AB/WW4BEG[2]
+ Tile_X2Y11_LUT4AB/WW4BEG[3] Tile_X2Y11_LUT4AB/WW4BEG[4] Tile_X2Y11_LUT4AB/WW4BEG[5]
+ Tile_X2Y11_LUT4AB/WW4BEG[6] Tile_X2Y11_LUT4AB/WW4BEG[7] Tile_X2Y11_LUT4AB/WW4BEG[8]
+ Tile_X2Y11_LUT4AB/WW4BEG[9] LUT4AB
XTile_X3Y1_LUT4AB Tile_X3Y2_LUT4AB/Co Tile_X3Y1_LUT4AB/Co Tile_X3Y1_LUT4AB/E1BEG[0]
+ Tile_X3Y1_LUT4AB/E1BEG[1] Tile_X3Y1_LUT4AB/E1BEG[2] Tile_X3Y1_LUT4AB/E1BEG[3] Tile_X3Y1_LUT4AB/E1END[0]
+ Tile_X3Y1_LUT4AB/E1END[1] Tile_X3Y1_LUT4AB/E1END[2] Tile_X3Y1_LUT4AB/E1END[3] Tile_X3Y1_LUT4AB/E2BEG[0]
+ Tile_X3Y1_LUT4AB/E2BEG[1] Tile_X3Y1_LUT4AB/E2BEG[2] Tile_X3Y1_LUT4AB/E2BEG[3] Tile_X3Y1_LUT4AB/E2BEG[4]
+ Tile_X3Y1_LUT4AB/E2BEG[5] Tile_X3Y1_LUT4AB/E2BEG[6] Tile_X3Y1_LUT4AB/E2BEG[7] Tile_X4Y1_RegFile/E2END[0]
+ Tile_X4Y1_RegFile/E2END[1] Tile_X4Y1_RegFile/E2END[2] Tile_X4Y1_RegFile/E2END[3]
+ Tile_X4Y1_RegFile/E2END[4] Tile_X4Y1_RegFile/E2END[5] Tile_X4Y1_RegFile/E2END[6]
+ Tile_X4Y1_RegFile/E2END[7] Tile_X3Y1_LUT4AB/E2END[0] Tile_X3Y1_LUT4AB/E2END[1] Tile_X3Y1_LUT4AB/E2END[2]
+ Tile_X3Y1_LUT4AB/E2END[3] Tile_X3Y1_LUT4AB/E2END[4] Tile_X3Y1_LUT4AB/E2END[5] Tile_X3Y1_LUT4AB/E2END[6]
+ Tile_X3Y1_LUT4AB/E2END[7] Tile_X3Y1_LUT4AB/E2MID[0] Tile_X3Y1_LUT4AB/E2MID[1] Tile_X3Y1_LUT4AB/E2MID[2]
+ Tile_X3Y1_LUT4AB/E2MID[3] Tile_X3Y1_LUT4AB/E2MID[4] Tile_X3Y1_LUT4AB/E2MID[5] Tile_X3Y1_LUT4AB/E2MID[6]
+ Tile_X3Y1_LUT4AB/E2MID[7] Tile_X3Y1_LUT4AB/E6BEG[0] Tile_X3Y1_LUT4AB/E6BEG[10] Tile_X3Y1_LUT4AB/E6BEG[11]
+ Tile_X3Y1_LUT4AB/E6BEG[1] Tile_X3Y1_LUT4AB/E6BEG[2] Tile_X3Y1_LUT4AB/E6BEG[3] Tile_X3Y1_LUT4AB/E6BEG[4]
+ Tile_X3Y1_LUT4AB/E6BEG[5] Tile_X3Y1_LUT4AB/E6BEG[6] Tile_X3Y1_LUT4AB/E6BEG[7] Tile_X3Y1_LUT4AB/E6BEG[8]
+ Tile_X3Y1_LUT4AB/E6BEG[9] Tile_X3Y1_LUT4AB/E6END[0] Tile_X3Y1_LUT4AB/E6END[10] Tile_X3Y1_LUT4AB/E6END[11]
+ Tile_X3Y1_LUT4AB/E6END[1] Tile_X3Y1_LUT4AB/E6END[2] Tile_X3Y1_LUT4AB/E6END[3] Tile_X3Y1_LUT4AB/E6END[4]
+ Tile_X3Y1_LUT4AB/E6END[5] Tile_X3Y1_LUT4AB/E6END[6] Tile_X3Y1_LUT4AB/E6END[7] Tile_X3Y1_LUT4AB/E6END[8]
+ Tile_X3Y1_LUT4AB/E6END[9] Tile_X3Y1_LUT4AB/EE4BEG[0] Tile_X3Y1_LUT4AB/EE4BEG[10]
+ Tile_X3Y1_LUT4AB/EE4BEG[11] Tile_X3Y1_LUT4AB/EE4BEG[12] Tile_X3Y1_LUT4AB/EE4BEG[13]
+ Tile_X3Y1_LUT4AB/EE4BEG[14] Tile_X3Y1_LUT4AB/EE4BEG[15] Tile_X3Y1_LUT4AB/EE4BEG[1]
+ Tile_X3Y1_LUT4AB/EE4BEG[2] Tile_X3Y1_LUT4AB/EE4BEG[3] Tile_X3Y1_LUT4AB/EE4BEG[4]
+ Tile_X3Y1_LUT4AB/EE4BEG[5] Tile_X3Y1_LUT4AB/EE4BEG[6] Tile_X3Y1_LUT4AB/EE4BEG[7]
+ Tile_X3Y1_LUT4AB/EE4BEG[8] Tile_X3Y1_LUT4AB/EE4BEG[9] Tile_X3Y1_LUT4AB/EE4END[0]
+ Tile_X3Y1_LUT4AB/EE4END[10] Tile_X3Y1_LUT4AB/EE4END[11] Tile_X3Y1_LUT4AB/EE4END[12]
+ Tile_X3Y1_LUT4AB/EE4END[13] Tile_X3Y1_LUT4AB/EE4END[14] Tile_X3Y1_LUT4AB/EE4END[15]
+ Tile_X3Y1_LUT4AB/EE4END[1] Tile_X3Y1_LUT4AB/EE4END[2] Tile_X3Y1_LUT4AB/EE4END[3]
+ Tile_X3Y1_LUT4AB/EE4END[4] Tile_X3Y1_LUT4AB/EE4END[5] Tile_X3Y1_LUT4AB/EE4END[6]
+ Tile_X3Y1_LUT4AB/EE4END[7] Tile_X3Y1_LUT4AB/EE4END[8] Tile_X3Y1_LUT4AB/EE4END[9]
+ Tile_X3Y1_LUT4AB/FrameData[0] Tile_X3Y1_LUT4AB/FrameData[10] Tile_X3Y1_LUT4AB/FrameData[11]
+ Tile_X3Y1_LUT4AB/FrameData[12] Tile_X3Y1_LUT4AB/FrameData[13] Tile_X3Y1_LUT4AB/FrameData[14]
+ Tile_X3Y1_LUT4AB/FrameData[15] Tile_X3Y1_LUT4AB/FrameData[16] Tile_X3Y1_LUT4AB/FrameData[17]
+ Tile_X3Y1_LUT4AB/FrameData[18] Tile_X3Y1_LUT4AB/FrameData[19] Tile_X3Y1_LUT4AB/FrameData[1]
+ Tile_X3Y1_LUT4AB/FrameData[20] Tile_X3Y1_LUT4AB/FrameData[21] Tile_X3Y1_LUT4AB/FrameData[22]
+ Tile_X3Y1_LUT4AB/FrameData[23] Tile_X3Y1_LUT4AB/FrameData[24] Tile_X3Y1_LUT4AB/FrameData[25]
+ Tile_X3Y1_LUT4AB/FrameData[26] Tile_X3Y1_LUT4AB/FrameData[27] Tile_X3Y1_LUT4AB/FrameData[28]
+ Tile_X3Y1_LUT4AB/FrameData[29] Tile_X3Y1_LUT4AB/FrameData[2] Tile_X3Y1_LUT4AB/FrameData[30]
+ Tile_X3Y1_LUT4AB/FrameData[31] Tile_X3Y1_LUT4AB/FrameData[3] Tile_X3Y1_LUT4AB/FrameData[4]
+ Tile_X3Y1_LUT4AB/FrameData[5] Tile_X3Y1_LUT4AB/FrameData[6] Tile_X3Y1_LUT4AB/FrameData[7]
+ Tile_X3Y1_LUT4AB/FrameData[8] Tile_X3Y1_LUT4AB/FrameData[9] Tile_X4Y1_RegFile/FrameData[0]
+ Tile_X4Y1_RegFile/FrameData[10] Tile_X4Y1_RegFile/FrameData[11] Tile_X4Y1_RegFile/FrameData[12]
+ Tile_X4Y1_RegFile/FrameData[13] Tile_X4Y1_RegFile/FrameData[14] Tile_X4Y1_RegFile/FrameData[15]
+ Tile_X4Y1_RegFile/FrameData[16] Tile_X4Y1_RegFile/FrameData[17] Tile_X4Y1_RegFile/FrameData[18]
+ Tile_X4Y1_RegFile/FrameData[19] Tile_X4Y1_RegFile/FrameData[1] Tile_X4Y1_RegFile/FrameData[20]
+ Tile_X4Y1_RegFile/FrameData[21] Tile_X4Y1_RegFile/FrameData[22] Tile_X4Y1_RegFile/FrameData[23]
+ Tile_X4Y1_RegFile/FrameData[24] Tile_X4Y1_RegFile/FrameData[25] Tile_X4Y1_RegFile/FrameData[26]
+ Tile_X4Y1_RegFile/FrameData[27] Tile_X4Y1_RegFile/FrameData[28] Tile_X4Y1_RegFile/FrameData[29]
+ Tile_X4Y1_RegFile/FrameData[2] Tile_X4Y1_RegFile/FrameData[30] Tile_X4Y1_RegFile/FrameData[31]
+ Tile_X4Y1_RegFile/FrameData[3] Tile_X4Y1_RegFile/FrameData[4] Tile_X4Y1_RegFile/FrameData[5]
+ Tile_X4Y1_RegFile/FrameData[6] Tile_X4Y1_RegFile/FrameData[7] Tile_X4Y1_RegFile/FrameData[8]
+ Tile_X4Y1_RegFile/FrameData[9] Tile_X3Y1_LUT4AB/FrameStrobe[0] Tile_X3Y1_LUT4AB/FrameStrobe[10]
+ Tile_X3Y1_LUT4AB/FrameStrobe[11] Tile_X3Y1_LUT4AB/FrameStrobe[12] Tile_X3Y1_LUT4AB/FrameStrobe[13]
+ Tile_X3Y1_LUT4AB/FrameStrobe[14] Tile_X3Y1_LUT4AB/FrameStrobe[15] Tile_X3Y1_LUT4AB/FrameStrobe[16]
+ Tile_X3Y1_LUT4AB/FrameStrobe[17] Tile_X3Y1_LUT4AB/FrameStrobe[18] Tile_X3Y1_LUT4AB/FrameStrobe[19]
+ Tile_X3Y1_LUT4AB/FrameStrobe[1] Tile_X3Y1_LUT4AB/FrameStrobe[2] Tile_X3Y1_LUT4AB/FrameStrobe[3]
+ Tile_X3Y1_LUT4AB/FrameStrobe[4] Tile_X3Y1_LUT4AB/FrameStrobe[5] Tile_X3Y1_LUT4AB/FrameStrobe[6]
+ Tile_X3Y1_LUT4AB/FrameStrobe[7] Tile_X3Y1_LUT4AB/FrameStrobe[8] Tile_X3Y1_LUT4AB/FrameStrobe[9]
+ Tile_X3Y1_LUT4AB/FrameStrobe_O[0] Tile_X3Y1_LUT4AB/FrameStrobe_O[10] Tile_X3Y1_LUT4AB/FrameStrobe_O[11]
+ Tile_X3Y1_LUT4AB/FrameStrobe_O[12] Tile_X3Y1_LUT4AB/FrameStrobe_O[13] Tile_X3Y1_LUT4AB/FrameStrobe_O[14]
+ Tile_X3Y1_LUT4AB/FrameStrobe_O[15] Tile_X3Y1_LUT4AB/FrameStrobe_O[16] Tile_X3Y1_LUT4AB/FrameStrobe_O[17]
+ Tile_X3Y1_LUT4AB/FrameStrobe_O[18] Tile_X3Y1_LUT4AB/FrameStrobe_O[19] Tile_X3Y1_LUT4AB/FrameStrobe_O[1]
+ Tile_X3Y1_LUT4AB/FrameStrobe_O[2] Tile_X3Y1_LUT4AB/FrameStrobe_O[3] Tile_X3Y1_LUT4AB/FrameStrobe_O[4]
+ Tile_X3Y1_LUT4AB/FrameStrobe_O[5] Tile_X3Y1_LUT4AB/FrameStrobe_O[6] Tile_X3Y1_LUT4AB/FrameStrobe_O[7]
+ Tile_X3Y1_LUT4AB/FrameStrobe_O[8] Tile_X3Y1_LUT4AB/FrameStrobe_O[9] Tile_X3Y1_LUT4AB/N1BEG[0]
+ Tile_X3Y1_LUT4AB/N1BEG[1] Tile_X3Y1_LUT4AB/N1BEG[2] Tile_X3Y1_LUT4AB/N1BEG[3] Tile_X3Y2_LUT4AB/N1BEG[0]
+ Tile_X3Y2_LUT4AB/N1BEG[1] Tile_X3Y2_LUT4AB/N1BEG[2] Tile_X3Y2_LUT4AB/N1BEG[3] Tile_X3Y1_LUT4AB/N2BEG[0]
+ Tile_X3Y1_LUT4AB/N2BEG[1] Tile_X3Y1_LUT4AB/N2BEG[2] Tile_X3Y1_LUT4AB/N2BEG[3] Tile_X3Y1_LUT4AB/N2BEG[4]
+ Tile_X3Y1_LUT4AB/N2BEG[5] Tile_X3Y1_LUT4AB/N2BEG[6] Tile_X3Y1_LUT4AB/N2BEG[7] Tile_X3Y1_LUT4AB/N2BEGb[0]
+ Tile_X3Y1_LUT4AB/N2BEGb[1] Tile_X3Y1_LUT4AB/N2BEGb[2] Tile_X3Y1_LUT4AB/N2BEGb[3]
+ Tile_X3Y1_LUT4AB/N2BEGb[4] Tile_X3Y1_LUT4AB/N2BEGb[5] Tile_X3Y1_LUT4AB/N2BEGb[6]
+ Tile_X3Y1_LUT4AB/N2BEGb[7] Tile_X3Y1_LUT4AB/N2END[0] Tile_X3Y1_LUT4AB/N2END[1] Tile_X3Y1_LUT4AB/N2END[2]
+ Tile_X3Y1_LUT4AB/N2END[3] Tile_X3Y1_LUT4AB/N2END[4] Tile_X3Y1_LUT4AB/N2END[5] Tile_X3Y1_LUT4AB/N2END[6]
+ Tile_X3Y1_LUT4AB/N2END[7] Tile_X3Y2_LUT4AB/N2BEG[0] Tile_X3Y2_LUT4AB/N2BEG[1] Tile_X3Y2_LUT4AB/N2BEG[2]
+ Tile_X3Y2_LUT4AB/N2BEG[3] Tile_X3Y2_LUT4AB/N2BEG[4] Tile_X3Y2_LUT4AB/N2BEG[5] Tile_X3Y2_LUT4AB/N2BEG[6]
+ Tile_X3Y2_LUT4AB/N2BEG[7] Tile_X3Y1_LUT4AB/N4BEG[0] Tile_X3Y1_LUT4AB/N4BEG[10] Tile_X3Y1_LUT4AB/N4BEG[11]
+ Tile_X3Y1_LUT4AB/N4BEG[12] Tile_X3Y1_LUT4AB/N4BEG[13] Tile_X3Y1_LUT4AB/N4BEG[14]
+ Tile_X3Y1_LUT4AB/N4BEG[15] Tile_X3Y1_LUT4AB/N4BEG[1] Tile_X3Y1_LUT4AB/N4BEG[2] Tile_X3Y1_LUT4AB/N4BEG[3]
+ Tile_X3Y1_LUT4AB/N4BEG[4] Tile_X3Y1_LUT4AB/N4BEG[5] Tile_X3Y1_LUT4AB/N4BEG[6] Tile_X3Y1_LUT4AB/N4BEG[7]
+ Tile_X3Y1_LUT4AB/N4BEG[8] Tile_X3Y1_LUT4AB/N4BEG[9] Tile_X3Y2_LUT4AB/N4BEG[0] Tile_X3Y2_LUT4AB/N4BEG[10]
+ Tile_X3Y2_LUT4AB/N4BEG[11] Tile_X3Y2_LUT4AB/N4BEG[12] Tile_X3Y2_LUT4AB/N4BEG[13]
+ Tile_X3Y2_LUT4AB/N4BEG[14] Tile_X3Y2_LUT4AB/N4BEG[15] Tile_X3Y2_LUT4AB/N4BEG[1]
+ Tile_X3Y2_LUT4AB/N4BEG[2] Tile_X3Y2_LUT4AB/N4BEG[3] Tile_X3Y2_LUT4AB/N4BEG[4] Tile_X3Y2_LUT4AB/N4BEG[5]
+ Tile_X3Y2_LUT4AB/N4BEG[6] Tile_X3Y2_LUT4AB/N4BEG[7] Tile_X3Y2_LUT4AB/N4BEG[8] Tile_X3Y2_LUT4AB/N4BEG[9]
+ Tile_X3Y1_LUT4AB/NN4BEG[0] Tile_X3Y1_LUT4AB/NN4BEG[10] Tile_X3Y1_LUT4AB/NN4BEG[11]
+ Tile_X3Y1_LUT4AB/NN4BEG[12] Tile_X3Y1_LUT4AB/NN4BEG[13] Tile_X3Y1_LUT4AB/NN4BEG[14]
+ Tile_X3Y1_LUT4AB/NN4BEG[15] Tile_X3Y1_LUT4AB/NN4BEG[1] Tile_X3Y1_LUT4AB/NN4BEG[2]
+ Tile_X3Y1_LUT4AB/NN4BEG[3] Tile_X3Y1_LUT4AB/NN4BEG[4] Tile_X3Y1_LUT4AB/NN4BEG[5]
+ Tile_X3Y1_LUT4AB/NN4BEG[6] Tile_X3Y1_LUT4AB/NN4BEG[7] Tile_X3Y1_LUT4AB/NN4BEG[8]
+ Tile_X3Y1_LUT4AB/NN4BEG[9] Tile_X3Y2_LUT4AB/NN4BEG[0] Tile_X3Y2_LUT4AB/NN4BEG[10]
+ Tile_X3Y2_LUT4AB/NN4BEG[11] Tile_X3Y2_LUT4AB/NN4BEG[12] Tile_X3Y2_LUT4AB/NN4BEG[13]
+ Tile_X3Y2_LUT4AB/NN4BEG[14] Tile_X3Y2_LUT4AB/NN4BEG[15] Tile_X3Y2_LUT4AB/NN4BEG[1]
+ Tile_X3Y2_LUT4AB/NN4BEG[2] Tile_X3Y2_LUT4AB/NN4BEG[3] Tile_X3Y2_LUT4AB/NN4BEG[4]
+ Tile_X3Y2_LUT4AB/NN4BEG[5] Tile_X3Y2_LUT4AB/NN4BEG[6] Tile_X3Y2_LUT4AB/NN4BEG[7]
+ Tile_X3Y2_LUT4AB/NN4BEG[8] Tile_X3Y2_LUT4AB/NN4BEG[9] Tile_X3Y2_LUT4AB/S1END[0]
+ Tile_X3Y2_LUT4AB/S1END[1] Tile_X3Y2_LUT4AB/S1END[2] Tile_X3Y2_LUT4AB/S1END[3] Tile_X3Y1_LUT4AB/S1END[0]
+ Tile_X3Y1_LUT4AB/S1END[1] Tile_X3Y1_LUT4AB/S1END[2] Tile_X3Y1_LUT4AB/S1END[3] Tile_X3Y2_LUT4AB/S2MID[0]
+ Tile_X3Y2_LUT4AB/S2MID[1] Tile_X3Y2_LUT4AB/S2MID[2] Tile_X3Y2_LUT4AB/S2MID[3] Tile_X3Y2_LUT4AB/S2MID[4]
+ Tile_X3Y2_LUT4AB/S2MID[5] Tile_X3Y2_LUT4AB/S2MID[6] Tile_X3Y2_LUT4AB/S2MID[7] Tile_X3Y2_LUT4AB/S2END[0]
+ Tile_X3Y2_LUT4AB/S2END[1] Tile_X3Y2_LUT4AB/S2END[2] Tile_X3Y2_LUT4AB/S2END[3] Tile_X3Y2_LUT4AB/S2END[4]
+ Tile_X3Y2_LUT4AB/S2END[5] Tile_X3Y2_LUT4AB/S2END[6] Tile_X3Y2_LUT4AB/S2END[7] Tile_X3Y1_LUT4AB/S2END[0]
+ Tile_X3Y1_LUT4AB/S2END[1] Tile_X3Y1_LUT4AB/S2END[2] Tile_X3Y1_LUT4AB/S2END[3] Tile_X3Y1_LUT4AB/S2END[4]
+ Tile_X3Y1_LUT4AB/S2END[5] Tile_X3Y1_LUT4AB/S2END[6] Tile_X3Y1_LUT4AB/S2END[7] Tile_X3Y1_LUT4AB/S2MID[0]
+ Tile_X3Y1_LUT4AB/S2MID[1] Tile_X3Y1_LUT4AB/S2MID[2] Tile_X3Y1_LUT4AB/S2MID[3] Tile_X3Y1_LUT4AB/S2MID[4]
+ Tile_X3Y1_LUT4AB/S2MID[5] Tile_X3Y1_LUT4AB/S2MID[6] Tile_X3Y1_LUT4AB/S2MID[7] Tile_X3Y2_LUT4AB/S4END[0]
+ Tile_X3Y2_LUT4AB/S4END[10] Tile_X3Y2_LUT4AB/S4END[11] Tile_X3Y2_LUT4AB/S4END[12]
+ Tile_X3Y2_LUT4AB/S4END[13] Tile_X3Y2_LUT4AB/S4END[14] Tile_X3Y2_LUT4AB/S4END[15]
+ Tile_X3Y2_LUT4AB/S4END[1] Tile_X3Y2_LUT4AB/S4END[2] Tile_X3Y2_LUT4AB/S4END[3] Tile_X3Y2_LUT4AB/S4END[4]
+ Tile_X3Y2_LUT4AB/S4END[5] Tile_X3Y2_LUT4AB/S4END[6] Tile_X3Y2_LUT4AB/S4END[7] Tile_X3Y2_LUT4AB/S4END[8]
+ Tile_X3Y2_LUT4AB/S4END[9] Tile_X3Y1_LUT4AB/S4END[0] Tile_X3Y1_LUT4AB/S4END[10] Tile_X3Y1_LUT4AB/S4END[11]
+ Tile_X3Y1_LUT4AB/S4END[12] Tile_X3Y1_LUT4AB/S4END[13] Tile_X3Y1_LUT4AB/S4END[14]
+ Tile_X3Y1_LUT4AB/S4END[15] Tile_X3Y1_LUT4AB/S4END[1] Tile_X3Y1_LUT4AB/S4END[2] Tile_X3Y1_LUT4AB/S4END[3]
+ Tile_X3Y1_LUT4AB/S4END[4] Tile_X3Y1_LUT4AB/S4END[5] Tile_X3Y1_LUT4AB/S4END[6] Tile_X3Y1_LUT4AB/S4END[7]
+ Tile_X3Y1_LUT4AB/S4END[8] Tile_X3Y1_LUT4AB/S4END[9] Tile_X3Y2_LUT4AB/SS4END[0] Tile_X3Y2_LUT4AB/SS4END[10]
+ Tile_X3Y2_LUT4AB/SS4END[11] Tile_X3Y2_LUT4AB/SS4END[12] Tile_X3Y2_LUT4AB/SS4END[13]
+ Tile_X3Y2_LUT4AB/SS4END[14] Tile_X3Y2_LUT4AB/SS4END[15] Tile_X3Y2_LUT4AB/SS4END[1]
+ Tile_X3Y2_LUT4AB/SS4END[2] Tile_X3Y2_LUT4AB/SS4END[3] Tile_X3Y2_LUT4AB/SS4END[4]
+ Tile_X3Y2_LUT4AB/SS4END[5] Tile_X3Y2_LUT4AB/SS4END[6] Tile_X3Y2_LUT4AB/SS4END[7]
+ Tile_X3Y2_LUT4AB/SS4END[8] Tile_X3Y2_LUT4AB/SS4END[9] Tile_X3Y1_LUT4AB/SS4END[0]
+ Tile_X3Y1_LUT4AB/SS4END[10] Tile_X3Y1_LUT4AB/SS4END[11] Tile_X3Y1_LUT4AB/SS4END[12]
+ Tile_X3Y1_LUT4AB/SS4END[13] Tile_X3Y1_LUT4AB/SS4END[14] Tile_X3Y1_LUT4AB/SS4END[15]
+ Tile_X3Y1_LUT4AB/SS4END[1] Tile_X3Y1_LUT4AB/SS4END[2] Tile_X3Y1_LUT4AB/SS4END[3]
+ Tile_X3Y1_LUT4AB/SS4END[4] Tile_X3Y1_LUT4AB/SS4END[5] Tile_X3Y1_LUT4AB/SS4END[6]
+ Tile_X3Y1_LUT4AB/SS4END[7] Tile_X3Y1_LUT4AB/SS4END[8] Tile_X3Y1_LUT4AB/SS4END[9]
+ Tile_X3Y1_LUT4AB/UserCLK Tile_X3Y1_LUT4AB/UserCLKo VGND VPWR Tile_X3Y1_LUT4AB/W1BEG[0]
+ Tile_X3Y1_LUT4AB/W1BEG[1] Tile_X3Y1_LUT4AB/W1BEG[2] Tile_X3Y1_LUT4AB/W1BEG[3] Tile_X3Y1_LUT4AB/W1END[0]
+ Tile_X3Y1_LUT4AB/W1END[1] Tile_X3Y1_LUT4AB/W1END[2] Tile_X3Y1_LUT4AB/W1END[3] Tile_X3Y1_LUT4AB/W2BEG[0]
+ Tile_X3Y1_LUT4AB/W2BEG[1] Tile_X3Y1_LUT4AB/W2BEG[2] Tile_X3Y1_LUT4AB/W2BEG[3] Tile_X3Y1_LUT4AB/W2BEG[4]
+ Tile_X3Y1_LUT4AB/W2BEG[5] Tile_X3Y1_LUT4AB/W2BEG[6] Tile_X3Y1_LUT4AB/W2BEG[7] Tile_X2Y1_LUT4AB/W2END[0]
+ Tile_X2Y1_LUT4AB/W2END[1] Tile_X2Y1_LUT4AB/W2END[2] Tile_X2Y1_LUT4AB/W2END[3] Tile_X2Y1_LUT4AB/W2END[4]
+ Tile_X2Y1_LUT4AB/W2END[5] Tile_X2Y1_LUT4AB/W2END[6] Tile_X2Y1_LUT4AB/W2END[7] Tile_X3Y1_LUT4AB/W2END[0]
+ Tile_X3Y1_LUT4AB/W2END[1] Tile_X3Y1_LUT4AB/W2END[2] Tile_X3Y1_LUT4AB/W2END[3] Tile_X3Y1_LUT4AB/W2END[4]
+ Tile_X3Y1_LUT4AB/W2END[5] Tile_X3Y1_LUT4AB/W2END[6] Tile_X3Y1_LUT4AB/W2END[7] Tile_X3Y1_LUT4AB/W2MID[0]
+ Tile_X3Y1_LUT4AB/W2MID[1] Tile_X3Y1_LUT4AB/W2MID[2] Tile_X3Y1_LUT4AB/W2MID[3] Tile_X3Y1_LUT4AB/W2MID[4]
+ Tile_X3Y1_LUT4AB/W2MID[5] Tile_X3Y1_LUT4AB/W2MID[6] Tile_X3Y1_LUT4AB/W2MID[7] Tile_X3Y1_LUT4AB/W6BEG[0]
+ Tile_X3Y1_LUT4AB/W6BEG[10] Tile_X3Y1_LUT4AB/W6BEG[11] Tile_X3Y1_LUT4AB/W6BEG[1]
+ Tile_X3Y1_LUT4AB/W6BEG[2] Tile_X3Y1_LUT4AB/W6BEG[3] Tile_X3Y1_LUT4AB/W6BEG[4] Tile_X3Y1_LUT4AB/W6BEG[5]
+ Tile_X3Y1_LUT4AB/W6BEG[6] Tile_X3Y1_LUT4AB/W6BEG[7] Tile_X3Y1_LUT4AB/W6BEG[8] Tile_X3Y1_LUT4AB/W6BEG[9]
+ Tile_X3Y1_LUT4AB/W6END[0] Tile_X3Y1_LUT4AB/W6END[10] Tile_X3Y1_LUT4AB/W6END[11]
+ Tile_X3Y1_LUT4AB/W6END[1] Tile_X3Y1_LUT4AB/W6END[2] Tile_X3Y1_LUT4AB/W6END[3] Tile_X3Y1_LUT4AB/W6END[4]
+ Tile_X3Y1_LUT4AB/W6END[5] Tile_X3Y1_LUT4AB/W6END[6] Tile_X3Y1_LUT4AB/W6END[7] Tile_X3Y1_LUT4AB/W6END[8]
+ Tile_X3Y1_LUT4AB/W6END[9] Tile_X3Y1_LUT4AB/WW4BEG[0] Tile_X3Y1_LUT4AB/WW4BEG[10]
+ Tile_X3Y1_LUT4AB/WW4BEG[11] Tile_X3Y1_LUT4AB/WW4BEG[12] Tile_X3Y1_LUT4AB/WW4BEG[13]
+ Tile_X3Y1_LUT4AB/WW4BEG[14] Tile_X3Y1_LUT4AB/WW4BEG[15] Tile_X3Y1_LUT4AB/WW4BEG[1]
+ Tile_X3Y1_LUT4AB/WW4BEG[2] Tile_X3Y1_LUT4AB/WW4BEG[3] Tile_X3Y1_LUT4AB/WW4BEG[4]
+ Tile_X3Y1_LUT4AB/WW4BEG[5] Tile_X3Y1_LUT4AB/WW4BEG[6] Tile_X3Y1_LUT4AB/WW4BEG[7]
+ Tile_X3Y1_LUT4AB/WW4BEG[8] Tile_X3Y1_LUT4AB/WW4BEG[9] Tile_X3Y1_LUT4AB/WW4END[0]
+ Tile_X3Y1_LUT4AB/WW4END[10] Tile_X3Y1_LUT4AB/WW4END[11] Tile_X3Y1_LUT4AB/WW4END[12]
+ Tile_X3Y1_LUT4AB/WW4END[13] Tile_X3Y1_LUT4AB/WW4END[14] Tile_X3Y1_LUT4AB/WW4END[15]
+ Tile_X3Y1_LUT4AB/WW4END[1] Tile_X3Y1_LUT4AB/WW4END[2] Tile_X3Y1_LUT4AB/WW4END[3]
+ Tile_X3Y1_LUT4AB/WW4END[4] Tile_X3Y1_LUT4AB/WW4END[5] Tile_X3Y1_LUT4AB/WW4END[6]
+ Tile_X3Y1_LUT4AB/WW4END[7] Tile_X3Y1_LUT4AB/WW4END[8] Tile_X3Y1_LUT4AB/WW4END[9]
+ LUT4AB
XTile_X0Y4_W_IO Tile_X0Y4_A_I_top Tile_X0Y4_A_O_top Tile_X0Y4_A_T_top Tile_X0Y4_A_config_C_bit0
+ Tile_X0Y4_A_config_C_bit1 Tile_X0Y4_A_config_C_bit2 Tile_X0Y4_A_config_C_bit3 Tile_X0Y4_B_I_top
+ Tile_X0Y4_B_O_top Tile_X0Y4_B_T_top Tile_X0Y4_B_config_C_bit0 Tile_X0Y4_B_config_C_bit1
+ Tile_X0Y4_B_config_C_bit2 Tile_X0Y4_B_config_C_bit3 Tile_X0Y4_W_IO/E1BEG[0] Tile_X0Y4_W_IO/E1BEG[1]
+ Tile_X0Y4_W_IO/E1BEG[2] Tile_X0Y4_W_IO/E1BEG[3] Tile_X0Y4_W_IO/E2BEG[0] Tile_X0Y4_W_IO/E2BEG[1]
+ Tile_X0Y4_W_IO/E2BEG[2] Tile_X0Y4_W_IO/E2BEG[3] Tile_X0Y4_W_IO/E2BEG[4] Tile_X0Y4_W_IO/E2BEG[5]
+ Tile_X0Y4_W_IO/E2BEG[6] Tile_X0Y4_W_IO/E2BEG[7] Tile_X0Y4_W_IO/E2BEGb[0] Tile_X0Y4_W_IO/E2BEGb[1]
+ Tile_X0Y4_W_IO/E2BEGb[2] Tile_X0Y4_W_IO/E2BEGb[3] Tile_X0Y4_W_IO/E2BEGb[4] Tile_X0Y4_W_IO/E2BEGb[5]
+ Tile_X0Y4_W_IO/E2BEGb[6] Tile_X0Y4_W_IO/E2BEGb[7] Tile_X0Y4_W_IO/E6BEG[0] Tile_X0Y4_W_IO/E6BEG[10]
+ Tile_X0Y4_W_IO/E6BEG[11] Tile_X0Y4_W_IO/E6BEG[1] Tile_X0Y4_W_IO/E6BEG[2] Tile_X0Y4_W_IO/E6BEG[3]
+ Tile_X0Y4_W_IO/E6BEG[4] Tile_X0Y4_W_IO/E6BEG[5] Tile_X0Y4_W_IO/E6BEG[6] Tile_X0Y4_W_IO/E6BEG[7]
+ Tile_X0Y4_W_IO/E6BEG[8] Tile_X0Y4_W_IO/E6BEG[9] Tile_X0Y4_W_IO/EE4BEG[0] Tile_X0Y4_W_IO/EE4BEG[10]
+ Tile_X0Y4_W_IO/EE4BEG[11] Tile_X0Y4_W_IO/EE4BEG[12] Tile_X0Y4_W_IO/EE4BEG[13] Tile_X0Y4_W_IO/EE4BEG[14]
+ Tile_X0Y4_W_IO/EE4BEG[15] Tile_X0Y4_W_IO/EE4BEG[1] Tile_X0Y4_W_IO/EE4BEG[2] Tile_X0Y4_W_IO/EE4BEG[3]
+ Tile_X0Y4_W_IO/EE4BEG[4] Tile_X0Y4_W_IO/EE4BEG[5] Tile_X0Y4_W_IO/EE4BEG[6] Tile_X0Y4_W_IO/EE4BEG[7]
+ Tile_X0Y4_W_IO/EE4BEG[8] Tile_X0Y4_W_IO/EE4BEG[9] FrameData[128] FrameData[138]
+ FrameData[139] FrameData[140] FrameData[141] FrameData[142] FrameData[143] FrameData[144]
+ FrameData[145] FrameData[146] FrameData[147] FrameData[129] FrameData[148] FrameData[149]
+ FrameData[150] FrameData[151] FrameData[152] FrameData[153] FrameData[154] FrameData[155]
+ FrameData[156] FrameData[157] FrameData[130] FrameData[158] FrameData[159] FrameData[131]
+ FrameData[132] FrameData[133] FrameData[134] FrameData[135] FrameData[136] FrameData[137]
+ Tile_X1Y4_LUT4AB/FrameData[0] Tile_X1Y4_LUT4AB/FrameData[10] Tile_X1Y4_LUT4AB/FrameData[11]
+ Tile_X1Y4_LUT4AB/FrameData[12] Tile_X1Y4_LUT4AB/FrameData[13] Tile_X1Y4_LUT4AB/FrameData[14]
+ Tile_X1Y4_LUT4AB/FrameData[15] Tile_X1Y4_LUT4AB/FrameData[16] Tile_X1Y4_LUT4AB/FrameData[17]
+ Tile_X1Y4_LUT4AB/FrameData[18] Tile_X1Y4_LUT4AB/FrameData[19] Tile_X1Y4_LUT4AB/FrameData[1]
+ Tile_X1Y4_LUT4AB/FrameData[20] Tile_X1Y4_LUT4AB/FrameData[21] Tile_X1Y4_LUT4AB/FrameData[22]
+ Tile_X1Y4_LUT4AB/FrameData[23] Tile_X1Y4_LUT4AB/FrameData[24] Tile_X1Y4_LUT4AB/FrameData[25]
+ Tile_X1Y4_LUT4AB/FrameData[26] Tile_X1Y4_LUT4AB/FrameData[27] Tile_X1Y4_LUT4AB/FrameData[28]
+ Tile_X1Y4_LUT4AB/FrameData[29] Tile_X1Y4_LUT4AB/FrameData[2] Tile_X1Y4_LUT4AB/FrameData[30]
+ Tile_X1Y4_LUT4AB/FrameData[31] Tile_X1Y4_LUT4AB/FrameData[3] Tile_X1Y4_LUT4AB/FrameData[4]
+ Tile_X1Y4_LUT4AB/FrameData[5] Tile_X1Y4_LUT4AB/FrameData[6] Tile_X1Y4_LUT4AB/FrameData[7]
+ Tile_X1Y4_LUT4AB/FrameData[8] Tile_X1Y4_LUT4AB/FrameData[9] Tile_X0Y4_W_IO/FrameStrobe[0]
+ Tile_X0Y4_W_IO/FrameStrobe[10] Tile_X0Y4_W_IO/FrameStrobe[11] Tile_X0Y4_W_IO/FrameStrobe[12]
+ Tile_X0Y4_W_IO/FrameStrobe[13] Tile_X0Y4_W_IO/FrameStrobe[14] Tile_X0Y4_W_IO/FrameStrobe[15]
+ Tile_X0Y4_W_IO/FrameStrobe[16] Tile_X0Y4_W_IO/FrameStrobe[17] Tile_X0Y4_W_IO/FrameStrobe[18]
+ Tile_X0Y4_W_IO/FrameStrobe[19] Tile_X0Y4_W_IO/FrameStrobe[1] Tile_X0Y4_W_IO/FrameStrobe[2]
+ Tile_X0Y4_W_IO/FrameStrobe[3] Tile_X0Y4_W_IO/FrameStrobe[4] Tile_X0Y4_W_IO/FrameStrobe[5]
+ Tile_X0Y4_W_IO/FrameStrobe[6] Tile_X0Y4_W_IO/FrameStrobe[7] Tile_X0Y4_W_IO/FrameStrobe[8]
+ Tile_X0Y4_W_IO/FrameStrobe[9] Tile_X0Y3_W_IO/FrameStrobe[0] Tile_X0Y3_W_IO/FrameStrobe[10]
+ Tile_X0Y3_W_IO/FrameStrobe[11] Tile_X0Y3_W_IO/FrameStrobe[12] Tile_X0Y3_W_IO/FrameStrobe[13]
+ Tile_X0Y3_W_IO/FrameStrobe[14] Tile_X0Y3_W_IO/FrameStrobe[15] Tile_X0Y3_W_IO/FrameStrobe[16]
+ Tile_X0Y3_W_IO/FrameStrobe[17] Tile_X0Y3_W_IO/FrameStrobe[18] Tile_X0Y3_W_IO/FrameStrobe[19]
+ Tile_X0Y3_W_IO/FrameStrobe[1] Tile_X0Y3_W_IO/FrameStrobe[2] Tile_X0Y3_W_IO/FrameStrobe[3]
+ Tile_X0Y3_W_IO/FrameStrobe[4] Tile_X0Y3_W_IO/FrameStrobe[5] Tile_X0Y3_W_IO/FrameStrobe[6]
+ Tile_X0Y3_W_IO/FrameStrobe[7] Tile_X0Y3_W_IO/FrameStrobe[8] Tile_X0Y3_W_IO/FrameStrobe[9]
+ Tile_X0Y4_W_IO/UserCLK Tile_X0Y3_W_IO/UserCLK VGND VPWR Tile_X0Y4_W_IO/W1END[0]
+ Tile_X0Y4_W_IO/W1END[1] Tile_X0Y4_W_IO/W1END[2] Tile_X0Y4_W_IO/W1END[3] Tile_X0Y4_W_IO/W2END[0]
+ Tile_X0Y4_W_IO/W2END[1] Tile_X0Y4_W_IO/W2END[2] Tile_X0Y4_W_IO/W2END[3] Tile_X0Y4_W_IO/W2END[4]
+ Tile_X0Y4_W_IO/W2END[5] Tile_X0Y4_W_IO/W2END[6] Tile_X0Y4_W_IO/W2END[7] Tile_X0Y4_W_IO/W2MID[0]
+ Tile_X0Y4_W_IO/W2MID[1] Tile_X0Y4_W_IO/W2MID[2] Tile_X0Y4_W_IO/W2MID[3] Tile_X0Y4_W_IO/W2MID[4]
+ Tile_X0Y4_W_IO/W2MID[5] Tile_X0Y4_W_IO/W2MID[6] Tile_X0Y4_W_IO/W2MID[7] Tile_X0Y4_W_IO/W6END[0]
+ Tile_X0Y4_W_IO/W6END[10] Tile_X0Y4_W_IO/W6END[11] Tile_X0Y4_W_IO/W6END[1] Tile_X0Y4_W_IO/W6END[2]
+ Tile_X0Y4_W_IO/W6END[3] Tile_X0Y4_W_IO/W6END[4] Tile_X0Y4_W_IO/W6END[5] Tile_X0Y4_W_IO/W6END[6]
+ Tile_X0Y4_W_IO/W6END[7] Tile_X0Y4_W_IO/W6END[8] Tile_X0Y4_W_IO/W6END[9] Tile_X0Y4_W_IO/WW4END[0]
+ Tile_X0Y4_W_IO/WW4END[10] Tile_X0Y4_W_IO/WW4END[11] Tile_X0Y4_W_IO/WW4END[12] Tile_X0Y4_W_IO/WW4END[13]
+ Tile_X0Y4_W_IO/WW4END[14] Tile_X0Y4_W_IO/WW4END[15] Tile_X0Y4_W_IO/WW4END[1] Tile_X0Y4_W_IO/WW4END[2]
+ Tile_X0Y4_W_IO/WW4END[3] Tile_X0Y4_W_IO/WW4END[4] Tile_X0Y4_W_IO/WW4END[5] Tile_X0Y4_W_IO/WW4END[6]
+ Tile_X0Y4_W_IO/WW4END[7] Tile_X0Y4_W_IO/WW4END[8] Tile_X0Y4_W_IO/WW4END[9] W_IO
XTile_X6Y6_LUT4AB Tile_X6Y7_LUT4AB/Co Tile_X6Y6_LUT4AB/Co Tile_X6Y6_LUT4AB/E1BEG[0]
+ Tile_X6Y6_LUT4AB/E1BEG[1] Tile_X6Y6_LUT4AB/E1BEG[2] Tile_X6Y6_LUT4AB/E1BEG[3] Tile_X6Y6_LUT4AB/E1END[0]
+ Tile_X6Y6_LUT4AB/E1END[1] Tile_X6Y6_LUT4AB/E1END[2] Tile_X6Y6_LUT4AB/E1END[3] Tile_X6Y6_LUT4AB/E2BEG[0]
+ Tile_X6Y6_LUT4AB/E2BEG[1] Tile_X6Y6_LUT4AB/E2BEG[2] Tile_X6Y6_LUT4AB/E2BEG[3] Tile_X6Y6_LUT4AB/E2BEG[4]
+ Tile_X6Y6_LUT4AB/E2BEG[5] Tile_X6Y6_LUT4AB/E2BEG[6] Tile_X6Y6_LUT4AB/E2BEG[7] Tile_X6Y6_LUT4AB/E2BEGb[0]
+ Tile_X6Y6_LUT4AB/E2BEGb[1] Tile_X6Y6_LUT4AB/E2BEGb[2] Tile_X6Y6_LUT4AB/E2BEGb[3]
+ Tile_X6Y6_LUT4AB/E2BEGb[4] Tile_X6Y6_LUT4AB/E2BEGb[5] Tile_X6Y6_LUT4AB/E2BEGb[6]
+ Tile_X6Y6_LUT4AB/E2BEGb[7] Tile_X6Y6_LUT4AB/E2END[0] Tile_X6Y6_LUT4AB/E2END[1] Tile_X6Y6_LUT4AB/E2END[2]
+ Tile_X6Y6_LUT4AB/E2END[3] Tile_X6Y6_LUT4AB/E2END[4] Tile_X6Y6_LUT4AB/E2END[5] Tile_X6Y6_LUT4AB/E2END[6]
+ Tile_X6Y6_LUT4AB/E2END[7] Tile_X6Y6_LUT4AB/E2MID[0] Tile_X6Y6_LUT4AB/E2MID[1] Tile_X6Y6_LUT4AB/E2MID[2]
+ Tile_X6Y6_LUT4AB/E2MID[3] Tile_X6Y6_LUT4AB/E2MID[4] Tile_X6Y6_LUT4AB/E2MID[5] Tile_X6Y6_LUT4AB/E2MID[6]
+ Tile_X6Y6_LUT4AB/E2MID[7] Tile_X6Y6_LUT4AB/E6BEG[0] Tile_X6Y6_LUT4AB/E6BEG[10] Tile_X6Y6_LUT4AB/E6BEG[11]
+ Tile_X6Y6_LUT4AB/E6BEG[1] Tile_X6Y6_LUT4AB/E6BEG[2] Tile_X6Y6_LUT4AB/E6BEG[3] Tile_X6Y6_LUT4AB/E6BEG[4]
+ Tile_X6Y6_LUT4AB/E6BEG[5] Tile_X6Y6_LUT4AB/E6BEG[6] Tile_X6Y6_LUT4AB/E6BEG[7] Tile_X6Y6_LUT4AB/E6BEG[8]
+ Tile_X6Y6_LUT4AB/E6BEG[9] Tile_X6Y6_LUT4AB/E6END[0] Tile_X6Y6_LUT4AB/E6END[10] Tile_X6Y6_LUT4AB/E6END[11]
+ Tile_X6Y6_LUT4AB/E6END[1] Tile_X6Y6_LUT4AB/E6END[2] Tile_X6Y6_LUT4AB/E6END[3] Tile_X6Y6_LUT4AB/E6END[4]
+ Tile_X6Y6_LUT4AB/E6END[5] Tile_X6Y6_LUT4AB/E6END[6] Tile_X6Y6_LUT4AB/E6END[7] Tile_X6Y6_LUT4AB/E6END[8]
+ Tile_X6Y6_LUT4AB/E6END[9] Tile_X6Y6_LUT4AB/EE4BEG[0] Tile_X6Y6_LUT4AB/EE4BEG[10]
+ Tile_X6Y6_LUT4AB/EE4BEG[11] Tile_X6Y6_LUT4AB/EE4BEG[12] Tile_X6Y6_LUT4AB/EE4BEG[13]
+ Tile_X6Y6_LUT4AB/EE4BEG[14] Tile_X6Y6_LUT4AB/EE4BEG[15] Tile_X6Y6_LUT4AB/EE4BEG[1]
+ Tile_X6Y6_LUT4AB/EE4BEG[2] Tile_X6Y6_LUT4AB/EE4BEG[3] Tile_X6Y6_LUT4AB/EE4BEG[4]
+ Tile_X6Y6_LUT4AB/EE4BEG[5] Tile_X6Y6_LUT4AB/EE4BEG[6] Tile_X6Y6_LUT4AB/EE4BEG[7]
+ Tile_X6Y6_LUT4AB/EE4BEG[8] Tile_X6Y6_LUT4AB/EE4BEG[9] Tile_X6Y6_LUT4AB/EE4END[0]
+ Tile_X6Y6_LUT4AB/EE4END[10] Tile_X6Y6_LUT4AB/EE4END[11] Tile_X6Y6_LUT4AB/EE4END[12]
+ Tile_X6Y6_LUT4AB/EE4END[13] Tile_X6Y6_LUT4AB/EE4END[14] Tile_X6Y6_LUT4AB/EE4END[15]
+ Tile_X6Y6_LUT4AB/EE4END[1] Tile_X6Y6_LUT4AB/EE4END[2] Tile_X6Y6_LUT4AB/EE4END[3]
+ Tile_X6Y6_LUT4AB/EE4END[4] Tile_X6Y6_LUT4AB/EE4END[5] Tile_X6Y6_LUT4AB/EE4END[6]
+ Tile_X6Y6_LUT4AB/EE4END[7] Tile_X6Y6_LUT4AB/EE4END[8] Tile_X6Y6_LUT4AB/EE4END[9]
+ Tile_X6Y6_LUT4AB/FrameData[0] Tile_X6Y6_LUT4AB/FrameData[10] Tile_X6Y6_LUT4AB/FrameData[11]
+ Tile_X6Y6_LUT4AB/FrameData[12] Tile_X6Y6_LUT4AB/FrameData[13] Tile_X6Y6_LUT4AB/FrameData[14]
+ Tile_X6Y6_LUT4AB/FrameData[15] Tile_X6Y6_LUT4AB/FrameData[16] Tile_X6Y6_LUT4AB/FrameData[17]
+ Tile_X6Y6_LUT4AB/FrameData[18] Tile_X6Y6_LUT4AB/FrameData[19] Tile_X6Y6_LUT4AB/FrameData[1]
+ Tile_X6Y6_LUT4AB/FrameData[20] Tile_X6Y6_LUT4AB/FrameData[21] Tile_X6Y6_LUT4AB/FrameData[22]
+ Tile_X6Y6_LUT4AB/FrameData[23] Tile_X6Y6_LUT4AB/FrameData[24] Tile_X6Y6_LUT4AB/FrameData[25]
+ Tile_X6Y6_LUT4AB/FrameData[26] Tile_X6Y6_LUT4AB/FrameData[27] Tile_X6Y6_LUT4AB/FrameData[28]
+ Tile_X6Y6_LUT4AB/FrameData[29] Tile_X6Y6_LUT4AB/FrameData[2] Tile_X6Y6_LUT4AB/FrameData[30]
+ Tile_X6Y6_LUT4AB/FrameData[31] Tile_X6Y6_LUT4AB/FrameData[3] Tile_X6Y6_LUT4AB/FrameData[4]
+ Tile_X6Y6_LUT4AB/FrameData[5] Tile_X6Y6_LUT4AB/FrameData[6] Tile_X6Y6_LUT4AB/FrameData[7]
+ Tile_X6Y6_LUT4AB/FrameData[8] Tile_X6Y6_LUT4AB/FrameData[9] Tile_X6Y6_LUT4AB/FrameData_O[0]
+ Tile_X6Y6_LUT4AB/FrameData_O[10] Tile_X6Y6_LUT4AB/FrameData_O[11] Tile_X6Y6_LUT4AB/FrameData_O[12]
+ Tile_X6Y6_LUT4AB/FrameData_O[13] Tile_X6Y6_LUT4AB/FrameData_O[14] Tile_X6Y6_LUT4AB/FrameData_O[15]
+ Tile_X6Y6_LUT4AB/FrameData_O[16] Tile_X6Y6_LUT4AB/FrameData_O[17] Tile_X6Y6_LUT4AB/FrameData_O[18]
+ Tile_X6Y6_LUT4AB/FrameData_O[19] Tile_X6Y6_LUT4AB/FrameData_O[1] Tile_X6Y6_LUT4AB/FrameData_O[20]
+ Tile_X6Y6_LUT4AB/FrameData_O[21] Tile_X6Y6_LUT4AB/FrameData_O[22] Tile_X6Y6_LUT4AB/FrameData_O[23]
+ Tile_X6Y6_LUT4AB/FrameData_O[24] Tile_X6Y6_LUT4AB/FrameData_O[25] Tile_X6Y6_LUT4AB/FrameData_O[26]
+ Tile_X6Y6_LUT4AB/FrameData_O[27] Tile_X6Y6_LUT4AB/FrameData_O[28] Tile_X6Y6_LUT4AB/FrameData_O[29]
+ Tile_X6Y6_LUT4AB/FrameData_O[2] Tile_X6Y6_LUT4AB/FrameData_O[30] Tile_X6Y6_LUT4AB/FrameData_O[31]
+ Tile_X6Y6_LUT4AB/FrameData_O[3] Tile_X6Y6_LUT4AB/FrameData_O[4] Tile_X6Y6_LUT4AB/FrameData_O[5]
+ Tile_X6Y6_LUT4AB/FrameData_O[6] Tile_X6Y6_LUT4AB/FrameData_O[7] Tile_X6Y6_LUT4AB/FrameData_O[8]
+ Tile_X6Y6_LUT4AB/FrameData_O[9] Tile_X6Y6_LUT4AB/FrameStrobe[0] Tile_X6Y6_LUT4AB/FrameStrobe[10]
+ Tile_X6Y6_LUT4AB/FrameStrobe[11] Tile_X6Y6_LUT4AB/FrameStrobe[12] Tile_X6Y6_LUT4AB/FrameStrobe[13]
+ Tile_X6Y6_LUT4AB/FrameStrobe[14] Tile_X6Y6_LUT4AB/FrameStrobe[15] Tile_X6Y6_LUT4AB/FrameStrobe[16]
+ Tile_X6Y6_LUT4AB/FrameStrobe[17] Tile_X6Y6_LUT4AB/FrameStrobe[18] Tile_X6Y6_LUT4AB/FrameStrobe[19]
+ Tile_X6Y6_LUT4AB/FrameStrobe[1] Tile_X6Y6_LUT4AB/FrameStrobe[2] Tile_X6Y6_LUT4AB/FrameStrobe[3]
+ Tile_X6Y6_LUT4AB/FrameStrobe[4] Tile_X6Y6_LUT4AB/FrameStrobe[5] Tile_X6Y6_LUT4AB/FrameStrobe[6]
+ Tile_X6Y6_LUT4AB/FrameStrobe[7] Tile_X6Y6_LUT4AB/FrameStrobe[8] Tile_X6Y6_LUT4AB/FrameStrobe[9]
+ Tile_X6Y5_LUT4AB/FrameStrobe[0] Tile_X6Y5_LUT4AB/FrameStrobe[10] Tile_X6Y5_LUT4AB/FrameStrobe[11]
+ Tile_X6Y5_LUT4AB/FrameStrobe[12] Tile_X6Y5_LUT4AB/FrameStrobe[13] Tile_X6Y5_LUT4AB/FrameStrobe[14]
+ Tile_X6Y5_LUT4AB/FrameStrobe[15] Tile_X6Y5_LUT4AB/FrameStrobe[16] Tile_X6Y5_LUT4AB/FrameStrobe[17]
+ Tile_X6Y5_LUT4AB/FrameStrobe[18] Tile_X6Y5_LUT4AB/FrameStrobe[19] Tile_X6Y5_LUT4AB/FrameStrobe[1]
+ Tile_X6Y5_LUT4AB/FrameStrobe[2] Tile_X6Y5_LUT4AB/FrameStrobe[3] Tile_X6Y5_LUT4AB/FrameStrobe[4]
+ Tile_X6Y5_LUT4AB/FrameStrobe[5] Tile_X6Y5_LUT4AB/FrameStrobe[6] Tile_X6Y5_LUT4AB/FrameStrobe[7]
+ Tile_X6Y5_LUT4AB/FrameStrobe[8] Tile_X6Y5_LUT4AB/FrameStrobe[9] Tile_X6Y6_LUT4AB/N1BEG[0]
+ Tile_X6Y6_LUT4AB/N1BEG[1] Tile_X6Y6_LUT4AB/N1BEG[2] Tile_X6Y6_LUT4AB/N1BEG[3] Tile_X6Y7_LUT4AB/N1BEG[0]
+ Tile_X6Y7_LUT4AB/N1BEG[1] Tile_X6Y7_LUT4AB/N1BEG[2] Tile_X6Y7_LUT4AB/N1BEG[3] Tile_X6Y6_LUT4AB/N2BEG[0]
+ Tile_X6Y6_LUT4AB/N2BEG[1] Tile_X6Y6_LUT4AB/N2BEG[2] Tile_X6Y6_LUT4AB/N2BEG[3] Tile_X6Y6_LUT4AB/N2BEG[4]
+ Tile_X6Y6_LUT4AB/N2BEG[5] Tile_X6Y6_LUT4AB/N2BEG[6] Tile_X6Y6_LUT4AB/N2BEG[7] Tile_X6Y5_LUT4AB/N2END[0]
+ Tile_X6Y5_LUT4AB/N2END[1] Tile_X6Y5_LUT4AB/N2END[2] Tile_X6Y5_LUT4AB/N2END[3] Tile_X6Y5_LUT4AB/N2END[4]
+ Tile_X6Y5_LUT4AB/N2END[5] Tile_X6Y5_LUT4AB/N2END[6] Tile_X6Y5_LUT4AB/N2END[7] Tile_X6Y6_LUT4AB/N2END[0]
+ Tile_X6Y6_LUT4AB/N2END[1] Tile_X6Y6_LUT4AB/N2END[2] Tile_X6Y6_LUT4AB/N2END[3] Tile_X6Y6_LUT4AB/N2END[4]
+ Tile_X6Y6_LUT4AB/N2END[5] Tile_X6Y6_LUT4AB/N2END[6] Tile_X6Y6_LUT4AB/N2END[7] Tile_X6Y7_LUT4AB/N2BEG[0]
+ Tile_X6Y7_LUT4AB/N2BEG[1] Tile_X6Y7_LUT4AB/N2BEG[2] Tile_X6Y7_LUT4AB/N2BEG[3] Tile_X6Y7_LUT4AB/N2BEG[4]
+ Tile_X6Y7_LUT4AB/N2BEG[5] Tile_X6Y7_LUT4AB/N2BEG[6] Tile_X6Y7_LUT4AB/N2BEG[7] Tile_X6Y6_LUT4AB/N4BEG[0]
+ Tile_X6Y6_LUT4AB/N4BEG[10] Tile_X6Y6_LUT4AB/N4BEG[11] Tile_X6Y6_LUT4AB/N4BEG[12]
+ Tile_X6Y6_LUT4AB/N4BEG[13] Tile_X6Y6_LUT4AB/N4BEG[14] Tile_X6Y6_LUT4AB/N4BEG[15]
+ Tile_X6Y6_LUT4AB/N4BEG[1] Tile_X6Y6_LUT4AB/N4BEG[2] Tile_X6Y6_LUT4AB/N4BEG[3] Tile_X6Y6_LUT4AB/N4BEG[4]
+ Tile_X6Y6_LUT4AB/N4BEG[5] Tile_X6Y6_LUT4AB/N4BEG[6] Tile_X6Y6_LUT4AB/N4BEG[7] Tile_X6Y6_LUT4AB/N4BEG[8]
+ Tile_X6Y6_LUT4AB/N4BEG[9] Tile_X6Y7_LUT4AB/N4BEG[0] Tile_X6Y7_LUT4AB/N4BEG[10] Tile_X6Y7_LUT4AB/N4BEG[11]
+ Tile_X6Y7_LUT4AB/N4BEG[12] Tile_X6Y7_LUT4AB/N4BEG[13] Tile_X6Y7_LUT4AB/N4BEG[14]
+ Tile_X6Y7_LUT4AB/N4BEG[15] Tile_X6Y7_LUT4AB/N4BEG[1] Tile_X6Y7_LUT4AB/N4BEG[2] Tile_X6Y7_LUT4AB/N4BEG[3]
+ Tile_X6Y7_LUT4AB/N4BEG[4] Tile_X6Y7_LUT4AB/N4BEG[5] Tile_X6Y7_LUT4AB/N4BEG[6] Tile_X6Y7_LUT4AB/N4BEG[7]
+ Tile_X6Y7_LUT4AB/N4BEG[8] Tile_X6Y7_LUT4AB/N4BEG[9] Tile_X6Y6_LUT4AB/NN4BEG[0] Tile_X6Y6_LUT4AB/NN4BEG[10]
+ Tile_X6Y6_LUT4AB/NN4BEG[11] Tile_X6Y6_LUT4AB/NN4BEG[12] Tile_X6Y6_LUT4AB/NN4BEG[13]
+ Tile_X6Y6_LUT4AB/NN4BEG[14] Tile_X6Y6_LUT4AB/NN4BEG[15] Tile_X6Y6_LUT4AB/NN4BEG[1]
+ Tile_X6Y6_LUT4AB/NN4BEG[2] Tile_X6Y6_LUT4AB/NN4BEG[3] Tile_X6Y6_LUT4AB/NN4BEG[4]
+ Tile_X6Y6_LUT4AB/NN4BEG[5] Tile_X6Y6_LUT4AB/NN4BEG[6] Tile_X6Y6_LUT4AB/NN4BEG[7]
+ Tile_X6Y6_LUT4AB/NN4BEG[8] Tile_X6Y6_LUT4AB/NN4BEG[9] Tile_X6Y7_LUT4AB/NN4BEG[0]
+ Tile_X6Y7_LUT4AB/NN4BEG[10] Tile_X6Y7_LUT4AB/NN4BEG[11] Tile_X6Y7_LUT4AB/NN4BEG[12]
+ Tile_X6Y7_LUT4AB/NN4BEG[13] Tile_X6Y7_LUT4AB/NN4BEG[14] Tile_X6Y7_LUT4AB/NN4BEG[15]
+ Tile_X6Y7_LUT4AB/NN4BEG[1] Tile_X6Y7_LUT4AB/NN4BEG[2] Tile_X6Y7_LUT4AB/NN4BEG[3]
+ Tile_X6Y7_LUT4AB/NN4BEG[4] Tile_X6Y7_LUT4AB/NN4BEG[5] Tile_X6Y7_LUT4AB/NN4BEG[6]
+ Tile_X6Y7_LUT4AB/NN4BEG[7] Tile_X6Y7_LUT4AB/NN4BEG[8] Tile_X6Y7_LUT4AB/NN4BEG[9]
+ Tile_X6Y7_LUT4AB/S1END[0] Tile_X6Y7_LUT4AB/S1END[1] Tile_X6Y7_LUT4AB/S1END[2] Tile_X6Y7_LUT4AB/S1END[3]
+ Tile_X6Y6_LUT4AB/S1END[0] Tile_X6Y6_LUT4AB/S1END[1] Tile_X6Y6_LUT4AB/S1END[2] Tile_X6Y6_LUT4AB/S1END[3]
+ Tile_X6Y7_LUT4AB/S2MID[0] Tile_X6Y7_LUT4AB/S2MID[1] Tile_X6Y7_LUT4AB/S2MID[2] Tile_X6Y7_LUT4AB/S2MID[3]
+ Tile_X6Y7_LUT4AB/S2MID[4] Tile_X6Y7_LUT4AB/S2MID[5] Tile_X6Y7_LUT4AB/S2MID[6] Tile_X6Y7_LUT4AB/S2MID[7]
+ Tile_X6Y7_LUT4AB/S2END[0] Tile_X6Y7_LUT4AB/S2END[1] Tile_X6Y7_LUT4AB/S2END[2] Tile_X6Y7_LUT4AB/S2END[3]
+ Tile_X6Y7_LUT4AB/S2END[4] Tile_X6Y7_LUT4AB/S2END[5] Tile_X6Y7_LUT4AB/S2END[6] Tile_X6Y7_LUT4AB/S2END[7]
+ Tile_X6Y6_LUT4AB/S2END[0] Tile_X6Y6_LUT4AB/S2END[1] Tile_X6Y6_LUT4AB/S2END[2] Tile_X6Y6_LUT4AB/S2END[3]
+ Tile_X6Y6_LUT4AB/S2END[4] Tile_X6Y6_LUT4AB/S2END[5] Tile_X6Y6_LUT4AB/S2END[6] Tile_X6Y6_LUT4AB/S2END[7]
+ Tile_X6Y6_LUT4AB/S2MID[0] Tile_X6Y6_LUT4AB/S2MID[1] Tile_X6Y6_LUT4AB/S2MID[2] Tile_X6Y6_LUT4AB/S2MID[3]
+ Tile_X6Y6_LUT4AB/S2MID[4] Tile_X6Y6_LUT4AB/S2MID[5] Tile_X6Y6_LUT4AB/S2MID[6] Tile_X6Y6_LUT4AB/S2MID[7]
+ Tile_X6Y7_LUT4AB/S4END[0] Tile_X6Y7_LUT4AB/S4END[10] Tile_X6Y7_LUT4AB/S4END[11]
+ Tile_X6Y7_LUT4AB/S4END[12] Tile_X6Y7_LUT4AB/S4END[13] Tile_X6Y7_LUT4AB/S4END[14]
+ Tile_X6Y7_LUT4AB/S4END[15] Tile_X6Y7_LUT4AB/S4END[1] Tile_X6Y7_LUT4AB/S4END[2] Tile_X6Y7_LUT4AB/S4END[3]
+ Tile_X6Y7_LUT4AB/S4END[4] Tile_X6Y7_LUT4AB/S4END[5] Tile_X6Y7_LUT4AB/S4END[6] Tile_X6Y7_LUT4AB/S4END[7]
+ Tile_X6Y7_LUT4AB/S4END[8] Tile_X6Y7_LUT4AB/S4END[9] Tile_X6Y6_LUT4AB/S4END[0] Tile_X6Y6_LUT4AB/S4END[10]
+ Tile_X6Y6_LUT4AB/S4END[11] Tile_X6Y6_LUT4AB/S4END[12] Tile_X6Y6_LUT4AB/S4END[13]
+ Tile_X6Y6_LUT4AB/S4END[14] Tile_X6Y6_LUT4AB/S4END[15] Tile_X6Y6_LUT4AB/S4END[1]
+ Tile_X6Y6_LUT4AB/S4END[2] Tile_X6Y6_LUT4AB/S4END[3] Tile_X6Y6_LUT4AB/S4END[4] Tile_X6Y6_LUT4AB/S4END[5]
+ Tile_X6Y6_LUT4AB/S4END[6] Tile_X6Y6_LUT4AB/S4END[7] Tile_X6Y6_LUT4AB/S4END[8] Tile_X6Y6_LUT4AB/S4END[9]
+ Tile_X6Y7_LUT4AB/SS4END[0] Tile_X6Y7_LUT4AB/SS4END[10] Tile_X6Y7_LUT4AB/SS4END[11]
+ Tile_X6Y7_LUT4AB/SS4END[12] Tile_X6Y7_LUT4AB/SS4END[13] Tile_X6Y7_LUT4AB/SS4END[14]
+ Tile_X6Y7_LUT4AB/SS4END[15] Tile_X6Y7_LUT4AB/SS4END[1] Tile_X6Y7_LUT4AB/SS4END[2]
+ Tile_X6Y7_LUT4AB/SS4END[3] Tile_X6Y7_LUT4AB/SS4END[4] Tile_X6Y7_LUT4AB/SS4END[5]
+ Tile_X6Y7_LUT4AB/SS4END[6] Tile_X6Y7_LUT4AB/SS4END[7] Tile_X6Y7_LUT4AB/SS4END[8]
+ Tile_X6Y7_LUT4AB/SS4END[9] Tile_X6Y6_LUT4AB/SS4END[0] Tile_X6Y6_LUT4AB/SS4END[10]
+ Tile_X6Y6_LUT4AB/SS4END[11] Tile_X6Y6_LUT4AB/SS4END[12] Tile_X6Y6_LUT4AB/SS4END[13]
+ Tile_X6Y6_LUT4AB/SS4END[14] Tile_X6Y6_LUT4AB/SS4END[15] Tile_X6Y6_LUT4AB/SS4END[1]
+ Tile_X6Y6_LUT4AB/SS4END[2] Tile_X6Y6_LUT4AB/SS4END[3] Tile_X6Y6_LUT4AB/SS4END[4]
+ Tile_X6Y6_LUT4AB/SS4END[5] Tile_X6Y6_LUT4AB/SS4END[6] Tile_X6Y6_LUT4AB/SS4END[7]
+ Tile_X6Y6_LUT4AB/SS4END[8] Tile_X6Y6_LUT4AB/SS4END[9] Tile_X6Y6_LUT4AB/UserCLK Tile_X6Y5_LUT4AB/UserCLK
+ VGND VPWR Tile_X6Y6_LUT4AB/W1BEG[0] Tile_X6Y6_LUT4AB/W1BEG[1] Tile_X6Y6_LUT4AB/W1BEG[2]
+ Tile_X6Y6_LUT4AB/W1BEG[3] Tile_X6Y6_LUT4AB/W1END[0] Tile_X6Y6_LUT4AB/W1END[1] Tile_X6Y6_LUT4AB/W1END[2]
+ Tile_X6Y6_LUT4AB/W1END[3] Tile_X6Y6_LUT4AB/W2BEG[0] Tile_X6Y6_LUT4AB/W2BEG[1] Tile_X6Y6_LUT4AB/W2BEG[2]
+ Tile_X6Y6_LUT4AB/W2BEG[3] Tile_X6Y6_LUT4AB/W2BEG[4] Tile_X6Y6_LUT4AB/W2BEG[5] Tile_X6Y6_LUT4AB/W2BEG[6]
+ Tile_X6Y6_LUT4AB/W2BEG[7] Tile_X5Y6_LUT4AB/W2END[0] Tile_X5Y6_LUT4AB/W2END[1] Tile_X5Y6_LUT4AB/W2END[2]
+ Tile_X5Y6_LUT4AB/W2END[3] Tile_X5Y6_LUT4AB/W2END[4] Tile_X5Y6_LUT4AB/W2END[5] Tile_X5Y6_LUT4AB/W2END[6]
+ Tile_X5Y6_LUT4AB/W2END[7] Tile_X6Y6_LUT4AB/W2END[0] Tile_X6Y6_LUT4AB/W2END[1] Tile_X6Y6_LUT4AB/W2END[2]
+ Tile_X6Y6_LUT4AB/W2END[3] Tile_X6Y6_LUT4AB/W2END[4] Tile_X6Y6_LUT4AB/W2END[5] Tile_X6Y6_LUT4AB/W2END[6]
+ Tile_X6Y6_LUT4AB/W2END[7] Tile_X6Y6_LUT4AB/W2MID[0] Tile_X6Y6_LUT4AB/W2MID[1] Tile_X6Y6_LUT4AB/W2MID[2]
+ Tile_X6Y6_LUT4AB/W2MID[3] Tile_X6Y6_LUT4AB/W2MID[4] Tile_X6Y6_LUT4AB/W2MID[5] Tile_X6Y6_LUT4AB/W2MID[6]
+ Tile_X6Y6_LUT4AB/W2MID[7] Tile_X6Y6_LUT4AB/W6BEG[0] Tile_X6Y6_LUT4AB/W6BEG[10] Tile_X6Y6_LUT4AB/W6BEG[11]
+ Tile_X6Y6_LUT4AB/W6BEG[1] Tile_X6Y6_LUT4AB/W6BEG[2] Tile_X6Y6_LUT4AB/W6BEG[3] Tile_X6Y6_LUT4AB/W6BEG[4]
+ Tile_X6Y6_LUT4AB/W6BEG[5] Tile_X6Y6_LUT4AB/W6BEG[6] Tile_X6Y6_LUT4AB/W6BEG[7] Tile_X6Y6_LUT4AB/W6BEG[8]
+ Tile_X6Y6_LUT4AB/W6BEG[9] Tile_X6Y6_LUT4AB/W6END[0] Tile_X6Y6_LUT4AB/W6END[10] Tile_X6Y6_LUT4AB/W6END[11]
+ Tile_X6Y6_LUT4AB/W6END[1] Tile_X6Y6_LUT4AB/W6END[2] Tile_X6Y6_LUT4AB/W6END[3] Tile_X6Y6_LUT4AB/W6END[4]
+ Tile_X6Y6_LUT4AB/W6END[5] Tile_X6Y6_LUT4AB/W6END[6] Tile_X6Y6_LUT4AB/W6END[7] Tile_X6Y6_LUT4AB/W6END[8]
+ Tile_X6Y6_LUT4AB/W6END[9] Tile_X6Y6_LUT4AB/WW4BEG[0] Tile_X6Y6_LUT4AB/WW4BEG[10]
+ Tile_X6Y6_LUT4AB/WW4BEG[11] Tile_X6Y6_LUT4AB/WW4BEG[12] Tile_X6Y6_LUT4AB/WW4BEG[13]
+ Tile_X6Y6_LUT4AB/WW4BEG[14] Tile_X6Y6_LUT4AB/WW4BEG[15] Tile_X6Y6_LUT4AB/WW4BEG[1]
+ Tile_X6Y6_LUT4AB/WW4BEG[2] Tile_X6Y6_LUT4AB/WW4BEG[3] Tile_X6Y6_LUT4AB/WW4BEG[4]
+ Tile_X6Y6_LUT4AB/WW4BEG[5] Tile_X6Y6_LUT4AB/WW4BEG[6] Tile_X6Y6_LUT4AB/WW4BEG[7]
+ Tile_X6Y6_LUT4AB/WW4BEG[8] Tile_X6Y6_LUT4AB/WW4BEG[9] Tile_X6Y6_LUT4AB/WW4END[0]
+ Tile_X6Y6_LUT4AB/WW4END[10] Tile_X6Y6_LUT4AB/WW4END[11] Tile_X6Y6_LUT4AB/WW4END[12]
+ Tile_X6Y6_LUT4AB/WW4END[13] Tile_X6Y6_LUT4AB/WW4END[14] Tile_X6Y6_LUT4AB/WW4END[15]
+ Tile_X6Y6_LUT4AB/WW4END[1] Tile_X6Y6_LUT4AB/WW4END[2] Tile_X6Y6_LUT4AB/WW4END[3]
+ Tile_X6Y6_LUT4AB/WW4END[4] Tile_X6Y6_LUT4AB/WW4END[5] Tile_X6Y6_LUT4AB/WW4END[6]
+ Tile_X6Y6_LUT4AB/WW4END[7] Tile_X6Y6_LUT4AB/WW4END[8] Tile_X6Y6_LUT4AB/WW4END[9]
+ LUT4AB
XTile_X2Y5_LUT4AB Tile_X2Y6_LUT4AB/Co Tile_X2Y5_LUT4AB/Co Tile_X3Y5_LUT4AB/E1END[0]
+ Tile_X3Y5_LUT4AB/E1END[1] Tile_X3Y5_LUT4AB/E1END[2] Tile_X3Y5_LUT4AB/E1END[3] Tile_X2Y5_LUT4AB/E1END[0]
+ Tile_X2Y5_LUT4AB/E1END[1] Tile_X2Y5_LUT4AB/E1END[2] Tile_X2Y5_LUT4AB/E1END[3] Tile_X3Y5_LUT4AB/E2MID[0]
+ Tile_X3Y5_LUT4AB/E2MID[1] Tile_X3Y5_LUT4AB/E2MID[2] Tile_X3Y5_LUT4AB/E2MID[3] Tile_X3Y5_LUT4AB/E2MID[4]
+ Tile_X3Y5_LUT4AB/E2MID[5] Tile_X3Y5_LUT4AB/E2MID[6] Tile_X3Y5_LUT4AB/E2MID[7] Tile_X3Y5_LUT4AB/E2END[0]
+ Tile_X3Y5_LUT4AB/E2END[1] Tile_X3Y5_LUT4AB/E2END[2] Tile_X3Y5_LUT4AB/E2END[3] Tile_X3Y5_LUT4AB/E2END[4]
+ Tile_X3Y5_LUT4AB/E2END[5] Tile_X3Y5_LUT4AB/E2END[6] Tile_X3Y5_LUT4AB/E2END[7] Tile_X2Y5_LUT4AB/E2END[0]
+ Tile_X2Y5_LUT4AB/E2END[1] Tile_X2Y5_LUT4AB/E2END[2] Tile_X2Y5_LUT4AB/E2END[3] Tile_X2Y5_LUT4AB/E2END[4]
+ Tile_X2Y5_LUT4AB/E2END[5] Tile_X2Y5_LUT4AB/E2END[6] Tile_X2Y5_LUT4AB/E2END[7] Tile_X2Y5_LUT4AB/E2MID[0]
+ Tile_X2Y5_LUT4AB/E2MID[1] Tile_X2Y5_LUT4AB/E2MID[2] Tile_X2Y5_LUT4AB/E2MID[3] Tile_X2Y5_LUT4AB/E2MID[4]
+ Tile_X2Y5_LUT4AB/E2MID[5] Tile_X2Y5_LUT4AB/E2MID[6] Tile_X2Y5_LUT4AB/E2MID[7] Tile_X3Y5_LUT4AB/E6END[0]
+ Tile_X3Y5_LUT4AB/E6END[10] Tile_X3Y5_LUT4AB/E6END[11] Tile_X3Y5_LUT4AB/E6END[1]
+ Tile_X3Y5_LUT4AB/E6END[2] Tile_X3Y5_LUT4AB/E6END[3] Tile_X3Y5_LUT4AB/E6END[4] Tile_X3Y5_LUT4AB/E6END[5]
+ Tile_X3Y5_LUT4AB/E6END[6] Tile_X3Y5_LUT4AB/E6END[7] Tile_X3Y5_LUT4AB/E6END[8] Tile_X3Y5_LUT4AB/E6END[9]
+ Tile_X2Y5_LUT4AB/E6END[0] Tile_X2Y5_LUT4AB/E6END[10] Tile_X2Y5_LUT4AB/E6END[11]
+ Tile_X2Y5_LUT4AB/E6END[1] Tile_X2Y5_LUT4AB/E6END[2] Tile_X2Y5_LUT4AB/E6END[3] Tile_X2Y5_LUT4AB/E6END[4]
+ Tile_X2Y5_LUT4AB/E6END[5] Tile_X2Y5_LUT4AB/E6END[6] Tile_X2Y5_LUT4AB/E6END[7] Tile_X2Y5_LUT4AB/E6END[8]
+ Tile_X2Y5_LUT4AB/E6END[9] Tile_X3Y5_LUT4AB/EE4END[0] Tile_X3Y5_LUT4AB/EE4END[10]
+ Tile_X3Y5_LUT4AB/EE4END[11] Tile_X3Y5_LUT4AB/EE4END[12] Tile_X3Y5_LUT4AB/EE4END[13]
+ Tile_X3Y5_LUT4AB/EE4END[14] Tile_X3Y5_LUT4AB/EE4END[15] Tile_X3Y5_LUT4AB/EE4END[1]
+ Tile_X3Y5_LUT4AB/EE4END[2] Tile_X3Y5_LUT4AB/EE4END[3] Tile_X3Y5_LUT4AB/EE4END[4]
+ Tile_X3Y5_LUT4AB/EE4END[5] Tile_X3Y5_LUT4AB/EE4END[6] Tile_X3Y5_LUT4AB/EE4END[7]
+ Tile_X3Y5_LUT4AB/EE4END[8] Tile_X3Y5_LUT4AB/EE4END[9] Tile_X2Y5_LUT4AB/EE4END[0]
+ Tile_X2Y5_LUT4AB/EE4END[10] Tile_X2Y5_LUT4AB/EE4END[11] Tile_X2Y5_LUT4AB/EE4END[12]
+ Tile_X2Y5_LUT4AB/EE4END[13] Tile_X2Y5_LUT4AB/EE4END[14] Tile_X2Y5_LUT4AB/EE4END[15]
+ Tile_X2Y5_LUT4AB/EE4END[1] Tile_X2Y5_LUT4AB/EE4END[2] Tile_X2Y5_LUT4AB/EE4END[3]
+ Tile_X2Y5_LUT4AB/EE4END[4] Tile_X2Y5_LUT4AB/EE4END[5] Tile_X2Y5_LUT4AB/EE4END[6]
+ Tile_X2Y5_LUT4AB/EE4END[7] Tile_X2Y5_LUT4AB/EE4END[8] Tile_X2Y5_LUT4AB/EE4END[9]
+ Tile_X2Y5_LUT4AB/FrameData[0] Tile_X2Y5_LUT4AB/FrameData[10] Tile_X2Y5_LUT4AB/FrameData[11]
+ Tile_X2Y5_LUT4AB/FrameData[12] Tile_X2Y5_LUT4AB/FrameData[13] Tile_X2Y5_LUT4AB/FrameData[14]
+ Tile_X2Y5_LUT4AB/FrameData[15] Tile_X2Y5_LUT4AB/FrameData[16] Tile_X2Y5_LUT4AB/FrameData[17]
+ Tile_X2Y5_LUT4AB/FrameData[18] Tile_X2Y5_LUT4AB/FrameData[19] Tile_X2Y5_LUT4AB/FrameData[1]
+ Tile_X2Y5_LUT4AB/FrameData[20] Tile_X2Y5_LUT4AB/FrameData[21] Tile_X2Y5_LUT4AB/FrameData[22]
+ Tile_X2Y5_LUT4AB/FrameData[23] Tile_X2Y5_LUT4AB/FrameData[24] Tile_X2Y5_LUT4AB/FrameData[25]
+ Tile_X2Y5_LUT4AB/FrameData[26] Tile_X2Y5_LUT4AB/FrameData[27] Tile_X2Y5_LUT4AB/FrameData[28]
+ Tile_X2Y5_LUT4AB/FrameData[29] Tile_X2Y5_LUT4AB/FrameData[2] Tile_X2Y5_LUT4AB/FrameData[30]
+ Tile_X2Y5_LUT4AB/FrameData[31] Tile_X2Y5_LUT4AB/FrameData[3] Tile_X2Y5_LUT4AB/FrameData[4]
+ Tile_X2Y5_LUT4AB/FrameData[5] Tile_X2Y5_LUT4AB/FrameData[6] Tile_X2Y5_LUT4AB/FrameData[7]
+ Tile_X2Y5_LUT4AB/FrameData[8] Tile_X2Y5_LUT4AB/FrameData[9] Tile_X3Y5_LUT4AB/FrameData[0]
+ Tile_X3Y5_LUT4AB/FrameData[10] Tile_X3Y5_LUT4AB/FrameData[11] Tile_X3Y5_LUT4AB/FrameData[12]
+ Tile_X3Y5_LUT4AB/FrameData[13] Tile_X3Y5_LUT4AB/FrameData[14] Tile_X3Y5_LUT4AB/FrameData[15]
+ Tile_X3Y5_LUT4AB/FrameData[16] Tile_X3Y5_LUT4AB/FrameData[17] Tile_X3Y5_LUT4AB/FrameData[18]
+ Tile_X3Y5_LUT4AB/FrameData[19] Tile_X3Y5_LUT4AB/FrameData[1] Tile_X3Y5_LUT4AB/FrameData[20]
+ Tile_X3Y5_LUT4AB/FrameData[21] Tile_X3Y5_LUT4AB/FrameData[22] Tile_X3Y5_LUT4AB/FrameData[23]
+ Tile_X3Y5_LUT4AB/FrameData[24] Tile_X3Y5_LUT4AB/FrameData[25] Tile_X3Y5_LUT4AB/FrameData[26]
+ Tile_X3Y5_LUT4AB/FrameData[27] Tile_X3Y5_LUT4AB/FrameData[28] Tile_X3Y5_LUT4AB/FrameData[29]
+ Tile_X3Y5_LUT4AB/FrameData[2] Tile_X3Y5_LUT4AB/FrameData[30] Tile_X3Y5_LUT4AB/FrameData[31]
+ Tile_X3Y5_LUT4AB/FrameData[3] Tile_X3Y5_LUT4AB/FrameData[4] Tile_X3Y5_LUT4AB/FrameData[5]
+ Tile_X3Y5_LUT4AB/FrameData[6] Tile_X3Y5_LUT4AB/FrameData[7] Tile_X3Y5_LUT4AB/FrameData[8]
+ Tile_X3Y5_LUT4AB/FrameData[9] Tile_X2Y5_LUT4AB/FrameStrobe[0] Tile_X2Y5_LUT4AB/FrameStrobe[10]
+ Tile_X2Y5_LUT4AB/FrameStrobe[11] Tile_X2Y5_LUT4AB/FrameStrobe[12] Tile_X2Y5_LUT4AB/FrameStrobe[13]
+ Tile_X2Y5_LUT4AB/FrameStrobe[14] Tile_X2Y5_LUT4AB/FrameStrobe[15] Tile_X2Y5_LUT4AB/FrameStrobe[16]
+ Tile_X2Y5_LUT4AB/FrameStrobe[17] Tile_X2Y5_LUT4AB/FrameStrobe[18] Tile_X2Y5_LUT4AB/FrameStrobe[19]
+ Tile_X2Y5_LUT4AB/FrameStrobe[1] Tile_X2Y5_LUT4AB/FrameStrobe[2] Tile_X2Y5_LUT4AB/FrameStrobe[3]
+ Tile_X2Y5_LUT4AB/FrameStrobe[4] Tile_X2Y5_LUT4AB/FrameStrobe[5] Tile_X2Y5_LUT4AB/FrameStrobe[6]
+ Tile_X2Y5_LUT4AB/FrameStrobe[7] Tile_X2Y5_LUT4AB/FrameStrobe[8] Tile_X2Y5_LUT4AB/FrameStrobe[9]
+ Tile_X2Y4_LUT4AB/FrameStrobe[0] Tile_X2Y4_LUT4AB/FrameStrobe[10] Tile_X2Y4_LUT4AB/FrameStrobe[11]
+ Tile_X2Y4_LUT4AB/FrameStrobe[12] Tile_X2Y4_LUT4AB/FrameStrobe[13] Tile_X2Y4_LUT4AB/FrameStrobe[14]
+ Tile_X2Y4_LUT4AB/FrameStrobe[15] Tile_X2Y4_LUT4AB/FrameStrobe[16] Tile_X2Y4_LUT4AB/FrameStrobe[17]
+ Tile_X2Y4_LUT4AB/FrameStrobe[18] Tile_X2Y4_LUT4AB/FrameStrobe[19] Tile_X2Y4_LUT4AB/FrameStrobe[1]
+ Tile_X2Y4_LUT4AB/FrameStrobe[2] Tile_X2Y4_LUT4AB/FrameStrobe[3] Tile_X2Y4_LUT4AB/FrameStrobe[4]
+ Tile_X2Y4_LUT4AB/FrameStrobe[5] Tile_X2Y4_LUT4AB/FrameStrobe[6] Tile_X2Y4_LUT4AB/FrameStrobe[7]
+ Tile_X2Y4_LUT4AB/FrameStrobe[8] Tile_X2Y4_LUT4AB/FrameStrobe[9] Tile_X2Y5_LUT4AB/N1BEG[0]
+ Tile_X2Y5_LUT4AB/N1BEG[1] Tile_X2Y5_LUT4AB/N1BEG[2] Tile_X2Y5_LUT4AB/N1BEG[3] Tile_X2Y6_LUT4AB/N1BEG[0]
+ Tile_X2Y6_LUT4AB/N1BEG[1] Tile_X2Y6_LUT4AB/N1BEG[2] Tile_X2Y6_LUT4AB/N1BEG[3] Tile_X2Y5_LUT4AB/N2BEG[0]
+ Tile_X2Y5_LUT4AB/N2BEG[1] Tile_X2Y5_LUT4AB/N2BEG[2] Tile_X2Y5_LUT4AB/N2BEG[3] Tile_X2Y5_LUT4AB/N2BEG[4]
+ Tile_X2Y5_LUT4AB/N2BEG[5] Tile_X2Y5_LUT4AB/N2BEG[6] Tile_X2Y5_LUT4AB/N2BEG[7] Tile_X2Y4_LUT4AB/N2END[0]
+ Tile_X2Y4_LUT4AB/N2END[1] Tile_X2Y4_LUT4AB/N2END[2] Tile_X2Y4_LUT4AB/N2END[3] Tile_X2Y4_LUT4AB/N2END[4]
+ Tile_X2Y4_LUT4AB/N2END[5] Tile_X2Y4_LUT4AB/N2END[6] Tile_X2Y4_LUT4AB/N2END[7] Tile_X2Y5_LUT4AB/N2END[0]
+ Tile_X2Y5_LUT4AB/N2END[1] Tile_X2Y5_LUT4AB/N2END[2] Tile_X2Y5_LUT4AB/N2END[3] Tile_X2Y5_LUT4AB/N2END[4]
+ Tile_X2Y5_LUT4AB/N2END[5] Tile_X2Y5_LUT4AB/N2END[6] Tile_X2Y5_LUT4AB/N2END[7] Tile_X2Y6_LUT4AB/N2BEG[0]
+ Tile_X2Y6_LUT4AB/N2BEG[1] Tile_X2Y6_LUT4AB/N2BEG[2] Tile_X2Y6_LUT4AB/N2BEG[3] Tile_X2Y6_LUT4AB/N2BEG[4]
+ Tile_X2Y6_LUT4AB/N2BEG[5] Tile_X2Y6_LUT4AB/N2BEG[6] Tile_X2Y6_LUT4AB/N2BEG[7] Tile_X2Y5_LUT4AB/N4BEG[0]
+ Tile_X2Y5_LUT4AB/N4BEG[10] Tile_X2Y5_LUT4AB/N4BEG[11] Tile_X2Y5_LUT4AB/N4BEG[12]
+ Tile_X2Y5_LUT4AB/N4BEG[13] Tile_X2Y5_LUT4AB/N4BEG[14] Tile_X2Y5_LUT4AB/N4BEG[15]
+ Tile_X2Y5_LUT4AB/N4BEG[1] Tile_X2Y5_LUT4AB/N4BEG[2] Tile_X2Y5_LUT4AB/N4BEG[3] Tile_X2Y5_LUT4AB/N4BEG[4]
+ Tile_X2Y5_LUT4AB/N4BEG[5] Tile_X2Y5_LUT4AB/N4BEG[6] Tile_X2Y5_LUT4AB/N4BEG[7] Tile_X2Y5_LUT4AB/N4BEG[8]
+ Tile_X2Y5_LUT4AB/N4BEG[9] Tile_X2Y6_LUT4AB/N4BEG[0] Tile_X2Y6_LUT4AB/N4BEG[10] Tile_X2Y6_LUT4AB/N4BEG[11]
+ Tile_X2Y6_LUT4AB/N4BEG[12] Tile_X2Y6_LUT4AB/N4BEG[13] Tile_X2Y6_LUT4AB/N4BEG[14]
+ Tile_X2Y6_LUT4AB/N4BEG[15] Tile_X2Y6_LUT4AB/N4BEG[1] Tile_X2Y6_LUT4AB/N4BEG[2] Tile_X2Y6_LUT4AB/N4BEG[3]
+ Tile_X2Y6_LUT4AB/N4BEG[4] Tile_X2Y6_LUT4AB/N4BEG[5] Tile_X2Y6_LUT4AB/N4BEG[6] Tile_X2Y6_LUT4AB/N4BEG[7]
+ Tile_X2Y6_LUT4AB/N4BEG[8] Tile_X2Y6_LUT4AB/N4BEG[9] Tile_X2Y5_LUT4AB/NN4BEG[0] Tile_X2Y5_LUT4AB/NN4BEG[10]
+ Tile_X2Y5_LUT4AB/NN4BEG[11] Tile_X2Y5_LUT4AB/NN4BEG[12] Tile_X2Y5_LUT4AB/NN4BEG[13]
+ Tile_X2Y5_LUT4AB/NN4BEG[14] Tile_X2Y5_LUT4AB/NN4BEG[15] Tile_X2Y5_LUT4AB/NN4BEG[1]
+ Tile_X2Y5_LUT4AB/NN4BEG[2] Tile_X2Y5_LUT4AB/NN4BEG[3] Tile_X2Y5_LUT4AB/NN4BEG[4]
+ Tile_X2Y5_LUT4AB/NN4BEG[5] Tile_X2Y5_LUT4AB/NN4BEG[6] Tile_X2Y5_LUT4AB/NN4BEG[7]
+ Tile_X2Y5_LUT4AB/NN4BEG[8] Tile_X2Y5_LUT4AB/NN4BEG[9] Tile_X2Y6_LUT4AB/NN4BEG[0]
+ Tile_X2Y6_LUT4AB/NN4BEG[10] Tile_X2Y6_LUT4AB/NN4BEG[11] Tile_X2Y6_LUT4AB/NN4BEG[12]
+ Tile_X2Y6_LUT4AB/NN4BEG[13] Tile_X2Y6_LUT4AB/NN4BEG[14] Tile_X2Y6_LUT4AB/NN4BEG[15]
+ Tile_X2Y6_LUT4AB/NN4BEG[1] Tile_X2Y6_LUT4AB/NN4BEG[2] Tile_X2Y6_LUT4AB/NN4BEG[3]
+ Tile_X2Y6_LUT4AB/NN4BEG[4] Tile_X2Y6_LUT4AB/NN4BEG[5] Tile_X2Y6_LUT4AB/NN4BEG[6]
+ Tile_X2Y6_LUT4AB/NN4BEG[7] Tile_X2Y6_LUT4AB/NN4BEG[8] Tile_X2Y6_LUT4AB/NN4BEG[9]
+ Tile_X2Y6_LUT4AB/S1END[0] Tile_X2Y6_LUT4AB/S1END[1] Tile_X2Y6_LUT4AB/S1END[2] Tile_X2Y6_LUT4AB/S1END[3]
+ Tile_X2Y5_LUT4AB/S1END[0] Tile_X2Y5_LUT4AB/S1END[1] Tile_X2Y5_LUT4AB/S1END[2] Tile_X2Y5_LUT4AB/S1END[3]
+ Tile_X2Y6_LUT4AB/S2MID[0] Tile_X2Y6_LUT4AB/S2MID[1] Tile_X2Y6_LUT4AB/S2MID[2] Tile_X2Y6_LUT4AB/S2MID[3]
+ Tile_X2Y6_LUT4AB/S2MID[4] Tile_X2Y6_LUT4AB/S2MID[5] Tile_X2Y6_LUT4AB/S2MID[6] Tile_X2Y6_LUT4AB/S2MID[7]
+ Tile_X2Y6_LUT4AB/S2END[0] Tile_X2Y6_LUT4AB/S2END[1] Tile_X2Y6_LUT4AB/S2END[2] Tile_X2Y6_LUT4AB/S2END[3]
+ Tile_X2Y6_LUT4AB/S2END[4] Tile_X2Y6_LUT4AB/S2END[5] Tile_X2Y6_LUT4AB/S2END[6] Tile_X2Y6_LUT4AB/S2END[7]
+ Tile_X2Y5_LUT4AB/S2END[0] Tile_X2Y5_LUT4AB/S2END[1] Tile_X2Y5_LUT4AB/S2END[2] Tile_X2Y5_LUT4AB/S2END[3]
+ Tile_X2Y5_LUT4AB/S2END[4] Tile_X2Y5_LUT4AB/S2END[5] Tile_X2Y5_LUT4AB/S2END[6] Tile_X2Y5_LUT4AB/S2END[7]
+ Tile_X2Y5_LUT4AB/S2MID[0] Tile_X2Y5_LUT4AB/S2MID[1] Tile_X2Y5_LUT4AB/S2MID[2] Tile_X2Y5_LUT4AB/S2MID[3]
+ Tile_X2Y5_LUT4AB/S2MID[4] Tile_X2Y5_LUT4AB/S2MID[5] Tile_X2Y5_LUT4AB/S2MID[6] Tile_X2Y5_LUT4AB/S2MID[7]
+ Tile_X2Y6_LUT4AB/S4END[0] Tile_X2Y6_LUT4AB/S4END[10] Tile_X2Y6_LUT4AB/S4END[11]
+ Tile_X2Y6_LUT4AB/S4END[12] Tile_X2Y6_LUT4AB/S4END[13] Tile_X2Y6_LUT4AB/S4END[14]
+ Tile_X2Y6_LUT4AB/S4END[15] Tile_X2Y6_LUT4AB/S4END[1] Tile_X2Y6_LUT4AB/S4END[2] Tile_X2Y6_LUT4AB/S4END[3]
+ Tile_X2Y6_LUT4AB/S4END[4] Tile_X2Y6_LUT4AB/S4END[5] Tile_X2Y6_LUT4AB/S4END[6] Tile_X2Y6_LUT4AB/S4END[7]
+ Tile_X2Y6_LUT4AB/S4END[8] Tile_X2Y6_LUT4AB/S4END[9] Tile_X2Y5_LUT4AB/S4END[0] Tile_X2Y5_LUT4AB/S4END[10]
+ Tile_X2Y5_LUT4AB/S4END[11] Tile_X2Y5_LUT4AB/S4END[12] Tile_X2Y5_LUT4AB/S4END[13]
+ Tile_X2Y5_LUT4AB/S4END[14] Tile_X2Y5_LUT4AB/S4END[15] Tile_X2Y5_LUT4AB/S4END[1]
+ Tile_X2Y5_LUT4AB/S4END[2] Tile_X2Y5_LUT4AB/S4END[3] Tile_X2Y5_LUT4AB/S4END[4] Tile_X2Y5_LUT4AB/S4END[5]
+ Tile_X2Y5_LUT4AB/S4END[6] Tile_X2Y5_LUT4AB/S4END[7] Tile_X2Y5_LUT4AB/S4END[8] Tile_X2Y5_LUT4AB/S4END[9]
+ Tile_X2Y6_LUT4AB/SS4END[0] Tile_X2Y6_LUT4AB/SS4END[10] Tile_X2Y6_LUT4AB/SS4END[11]
+ Tile_X2Y6_LUT4AB/SS4END[12] Tile_X2Y6_LUT4AB/SS4END[13] Tile_X2Y6_LUT4AB/SS4END[14]
+ Tile_X2Y6_LUT4AB/SS4END[15] Tile_X2Y6_LUT4AB/SS4END[1] Tile_X2Y6_LUT4AB/SS4END[2]
+ Tile_X2Y6_LUT4AB/SS4END[3] Tile_X2Y6_LUT4AB/SS4END[4] Tile_X2Y6_LUT4AB/SS4END[5]
+ Tile_X2Y6_LUT4AB/SS4END[6] Tile_X2Y6_LUT4AB/SS4END[7] Tile_X2Y6_LUT4AB/SS4END[8]
+ Tile_X2Y6_LUT4AB/SS4END[9] Tile_X2Y5_LUT4AB/SS4END[0] Tile_X2Y5_LUT4AB/SS4END[10]
+ Tile_X2Y5_LUT4AB/SS4END[11] Tile_X2Y5_LUT4AB/SS4END[12] Tile_X2Y5_LUT4AB/SS4END[13]
+ Tile_X2Y5_LUT4AB/SS4END[14] Tile_X2Y5_LUT4AB/SS4END[15] Tile_X2Y5_LUT4AB/SS4END[1]
+ Tile_X2Y5_LUT4AB/SS4END[2] Tile_X2Y5_LUT4AB/SS4END[3] Tile_X2Y5_LUT4AB/SS4END[4]
+ Tile_X2Y5_LUT4AB/SS4END[5] Tile_X2Y5_LUT4AB/SS4END[6] Tile_X2Y5_LUT4AB/SS4END[7]
+ Tile_X2Y5_LUT4AB/SS4END[8] Tile_X2Y5_LUT4AB/SS4END[9] Tile_X2Y5_LUT4AB/UserCLK Tile_X2Y4_LUT4AB/UserCLK
+ VGND VPWR Tile_X2Y5_LUT4AB/W1BEG[0] Tile_X2Y5_LUT4AB/W1BEG[1] Tile_X2Y5_LUT4AB/W1BEG[2]
+ Tile_X2Y5_LUT4AB/W1BEG[3] Tile_X3Y5_LUT4AB/W1BEG[0] Tile_X3Y5_LUT4AB/W1BEG[1] Tile_X3Y5_LUT4AB/W1BEG[2]
+ Tile_X3Y5_LUT4AB/W1BEG[3] Tile_X2Y5_LUT4AB/W2BEG[0] Tile_X2Y5_LUT4AB/W2BEG[1] Tile_X2Y5_LUT4AB/W2BEG[2]
+ Tile_X2Y5_LUT4AB/W2BEG[3] Tile_X2Y5_LUT4AB/W2BEG[4] Tile_X2Y5_LUT4AB/W2BEG[5] Tile_X2Y5_LUT4AB/W2BEG[6]
+ Tile_X2Y5_LUT4AB/W2BEG[7] Tile_X1Y5_LUT4AB/W2END[0] Tile_X1Y5_LUT4AB/W2END[1] Tile_X1Y5_LUT4AB/W2END[2]
+ Tile_X1Y5_LUT4AB/W2END[3] Tile_X1Y5_LUT4AB/W2END[4] Tile_X1Y5_LUT4AB/W2END[5] Tile_X1Y5_LUT4AB/W2END[6]
+ Tile_X1Y5_LUT4AB/W2END[7] Tile_X2Y5_LUT4AB/W2END[0] Tile_X2Y5_LUT4AB/W2END[1] Tile_X2Y5_LUT4AB/W2END[2]
+ Tile_X2Y5_LUT4AB/W2END[3] Tile_X2Y5_LUT4AB/W2END[4] Tile_X2Y5_LUT4AB/W2END[5] Tile_X2Y5_LUT4AB/W2END[6]
+ Tile_X2Y5_LUT4AB/W2END[7] Tile_X3Y5_LUT4AB/W2BEG[0] Tile_X3Y5_LUT4AB/W2BEG[1] Tile_X3Y5_LUT4AB/W2BEG[2]
+ Tile_X3Y5_LUT4AB/W2BEG[3] Tile_X3Y5_LUT4AB/W2BEG[4] Tile_X3Y5_LUT4AB/W2BEG[5] Tile_X3Y5_LUT4AB/W2BEG[6]
+ Tile_X3Y5_LUT4AB/W2BEG[7] Tile_X2Y5_LUT4AB/W6BEG[0] Tile_X2Y5_LUT4AB/W6BEG[10] Tile_X2Y5_LUT4AB/W6BEG[11]
+ Tile_X2Y5_LUT4AB/W6BEG[1] Tile_X2Y5_LUT4AB/W6BEG[2] Tile_X2Y5_LUT4AB/W6BEG[3] Tile_X2Y5_LUT4AB/W6BEG[4]
+ Tile_X2Y5_LUT4AB/W6BEG[5] Tile_X2Y5_LUT4AB/W6BEG[6] Tile_X2Y5_LUT4AB/W6BEG[7] Tile_X2Y5_LUT4AB/W6BEG[8]
+ Tile_X2Y5_LUT4AB/W6BEG[9] Tile_X3Y5_LUT4AB/W6BEG[0] Tile_X3Y5_LUT4AB/W6BEG[10] Tile_X3Y5_LUT4AB/W6BEG[11]
+ Tile_X3Y5_LUT4AB/W6BEG[1] Tile_X3Y5_LUT4AB/W6BEG[2] Tile_X3Y5_LUT4AB/W6BEG[3] Tile_X3Y5_LUT4AB/W6BEG[4]
+ Tile_X3Y5_LUT4AB/W6BEG[5] Tile_X3Y5_LUT4AB/W6BEG[6] Tile_X3Y5_LUT4AB/W6BEG[7] Tile_X3Y5_LUT4AB/W6BEG[8]
+ Tile_X3Y5_LUT4AB/W6BEG[9] Tile_X2Y5_LUT4AB/WW4BEG[0] Tile_X2Y5_LUT4AB/WW4BEG[10]
+ Tile_X2Y5_LUT4AB/WW4BEG[11] Tile_X2Y5_LUT4AB/WW4BEG[12] Tile_X2Y5_LUT4AB/WW4BEG[13]
+ Tile_X2Y5_LUT4AB/WW4BEG[14] Tile_X2Y5_LUT4AB/WW4BEG[15] Tile_X2Y5_LUT4AB/WW4BEG[1]
+ Tile_X2Y5_LUT4AB/WW4BEG[2] Tile_X2Y5_LUT4AB/WW4BEG[3] Tile_X2Y5_LUT4AB/WW4BEG[4]
+ Tile_X2Y5_LUT4AB/WW4BEG[5] Tile_X2Y5_LUT4AB/WW4BEG[6] Tile_X2Y5_LUT4AB/WW4BEG[7]
+ Tile_X2Y5_LUT4AB/WW4BEG[8] Tile_X2Y5_LUT4AB/WW4BEG[9] Tile_X3Y5_LUT4AB/WW4BEG[0]
+ Tile_X3Y5_LUT4AB/WW4BEG[10] Tile_X3Y5_LUT4AB/WW4BEG[11] Tile_X3Y5_LUT4AB/WW4BEG[12]
+ Tile_X3Y5_LUT4AB/WW4BEG[13] Tile_X3Y5_LUT4AB/WW4BEG[14] Tile_X3Y5_LUT4AB/WW4BEG[15]
+ Tile_X3Y5_LUT4AB/WW4BEG[1] Tile_X3Y5_LUT4AB/WW4BEG[2] Tile_X3Y5_LUT4AB/WW4BEG[3]
+ Tile_X3Y5_LUT4AB/WW4BEG[4] Tile_X3Y5_LUT4AB/WW4BEG[5] Tile_X3Y5_LUT4AB/WW4BEG[6]
+ Tile_X3Y5_LUT4AB/WW4BEG[7] Tile_X3Y5_LUT4AB/WW4BEG[8] Tile_X3Y5_LUT4AB/WW4BEG[9]
+ LUT4AB
XTile_X5Y11_LUT4AB Tile_X5Y12_LUT4AB/Co Tile_X5Y11_LUT4AB/Co Tile_X6Y11_LUT4AB/E1END[0]
+ Tile_X6Y11_LUT4AB/E1END[1] Tile_X6Y11_LUT4AB/E1END[2] Tile_X6Y11_LUT4AB/E1END[3]
+ Tile_X5Y11_LUT4AB/E1END[0] Tile_X5Y11_LUT4AB/E1END[1] Tile_X5Y11_LUT4AB/E1END[2]
+ Tile_X5Y11_LUT4AB/E1END[3] Tile_X6Y11_LUT4AB/E2MID[0] Tile_X6Y11_LUT4AB/E2MID[1]
+ Tile_X6Y11_LUT4AB/E2MID[2] Tile_X6Y11_LUT4AB/E2MID[3] Tile_X6Y11_LUT4AB/E2MID[4]
+ Tile_X6Y11_LUT4AB/E2MID[5] Tile_X6Y11_LUT4AB/E2MID[6] Tile_X6Y11_LUT4AB/E2MID[7]
+ Tile_X6Y11_LUT4AB/E2END[0] Tile_X6Y11_LUT4AB/E2END[1] Tile_X6Y11_LUT4AB/E2END[2]
+ Tile_X6Y11_LUT4AB/E2END[3] Tile_X6Y11_LUT4AB/E2END[4] Tile_X6Y11_LUT4AB/E2END[5]
+ Tile_X6Y11_LUT4AB/E2END[6] Tile_X6Y11_LUT4AB/E2END[7] Tile_X5Y11_LUT4AB/E2END[0]
+ Tile_X5Y11_LUT4AB/E2END[1] Tile_X5Y11_LUT4AB/E2END[2] Tile_X5Y11_LUT4AB/E2END[3]
+ Tile_X5Y11_LUT4AB/E2END[4] Tile_X5Y11_LUT4AB/E2END[5] Tile_X5Y11_LUT4AB/E2END[6]
+ Tile_X5Y11_LUT4AB/E2END[7] Tile_X5Y11_LUT4AB/E2MID[0] Tile_X5Y11_LUT4AB/E2MID[1]
+ Tile_X5Y11_LUT4AB/E2MID[2] Tile_X5Y11_LUT4AB/E2MID[3] Tile_X5Y11_LUT4AB/E2MID[4]
+ Tile_X5Y11_LUT4AB/E2MID[5] Tile_X5Y11_LUT4AB/E2MID[6] Tile_X5Y11_LUT4AB/E2MID[7]
+ Tile_X6Y11_LUT4AB/E6END[0] Tile_X6Y11_LUT4AB/E6END[10] Tile_X6Y11_LUT4AB/E6END[11]
+ Tile_X6Y11_LUT4AB/E6END[1] Tile_X6Y11_LUT4AB/E6END[2] Tile_X6Y11_LUT4AB/E6END[3]
+ Tile_X6Y11_LUT4AB/E6END[4] Tile_X6Y11_LUT4AB/E6END[5] Tile_X6Y11_LUT4AB/E6END[6]
+ Tile_X6Y11_LUT4AB/E6END[7] Tile_X6Y11_LUT4AB/E6END[8] Tile_X6Y11_LUT4AB/E6END[9]
+ Tile_X5Y11_LUT4AB/E6END[0] Tile_X5Y11_LUT4AB/E6END[10] Tile_X5Y11_LUT4AB/E6END[11]
+ Tile_X5Y11_LUT4AB/E6END[1] Tile_X5Y11_LUT4AB/E6END[2] Tile_X5Y11_LUT4AB/E6END[3]
+ Tile_X5Y11_LUT4AB/E6END[4] Tile_X5Y11_LUT4AB/E6END[5] Tile_X5Y11_LUT4AB/E6END[6]
+ Tile_X5Y11_LUT4AB/E6END[7] Tile_X5Y11_LUT4AB/E6END[8] Tile_X5Y11_LUT4AB/E6END[9]
+ Tile_X6Y11_LUT4AB/EE4END[0] Tile_X6Y11_LUT4AB/EE4END[10] Tile_X6Y11_LUT4AB/EE4END[11]
+ Tile_X6Y11_LUT4AB/EE4END[12] Tile_X6Y11_LUT4AB/EE4END[13] Tile_X6Y11_LUT4AB/EE4END[14]
+ Tile_X6Y11_LUT4AB/EE4END[15] Tile_X6Y11_LUT4AB/EE4END[1] Tile_X6Y11_LUT4AB/EE4END[2]
+ Tile_X6Y11_LUT4AB/EE4END[3] Tile_X6Y11_LUT4AB/EE4END[4] Tile_X6Y11_LUT4AB/EE4END[5]
+ Tile_X6Y11_LUT4AB/EE4END[6] Tile_X6Y11_LUT4AB/EE4END[7] Tile_X6Y11_LUT4AB/EE4END[8]
+ Tile_X6Y11_LUT4AB/EE4END[9] Tile_X5Y11_LUT4AB/EE4END[0] Tile_X5Y11_LUT4AB/EE4END[10]
+ Tile_X5Y11_LUT4AB/EE4END[11] Tile_X5Y11_LUT4AB/EE4END[12] Tile_X5Y11_LUT4AB/EE4END[13]
+ Tile_X5Y11_LUT4AB/EE4END[14] Tile_X5Y11_LUT4AB/EE4END[15] Tile_X5Y11_LUT4AB/EE4END[1]
+ Tile_X5Y11_LUT4AB/EE4END[2] Tile_X5Y11_LUT4AB/EE4END[3] Tile_X5Y11_LUT4AB/EE4END[4]
+ Tile_X5Y11_LUT4AB/EE4END[5] Tile_X5Y11_LUT4AB/EE4END[6] Tile_X5Y11_LUT4AB/EE4END[7]
+ Tile_X5Y11_LUT4AB/EE4END[8] Tile_X5Y11_LUT4AB/EE4END[9] Tile_X5Y11_LUT4AB/FrameData[0]
+ Tile_X5Y11_LUT4AB/FrameData[10] Tile_X5Y11_LUT4AB/FrameData[11] Tile_X5Y11_LUT4AB/FrameData[12]
+ Tile_X5Y11_LUT4AB/FrameData[13] Tile_X5Y11_LUT4AB/FrameData[14] Tile_X5Y11_LUT4AB/FrameData[15]
+ Tile_X5Y11_LUT4AB/FrameData[16] Tile_X5Y11_LUT4AB/FrameData[17] Tile_X5Y11_LUT4AB/FrameData[18]
+ Tile_X5Y11_LUT4AB/FrameData[19] Tile_X5Y11_LUT4AB/FrameData[1] Tile_X5Y11_LUT4AB/FrameData[20]
+ Tile_X5Y11_LUT4AB/FrameData[21] Tile_X5Y11_LUT4AB/FrameData[22] Tile_X5Y11_LUT4AB/FrameData[23]
+ Tile_X5Y11_LUT4AB/FrameData[24] Tile_X5Y11_LUT4AB/FrameData[25] Tile_X5Y11_LUT4AB/FrameData[26]
+ Tile_X5Y11_LUT4AB/FrameData[27] Tile_X5Y11_LUT4AB/FrameData[28] Tile_X5Y11_LUT4AB/FrameData[29]
+ Tile_X5Y11_LUT4AB/FrameData[2] Tile_X5Y11_LUT4AB/FrameData[30] Tile_X5Y11_LUT4AB/FrameData[31]
+ Tile_X5Y11_LUT4AB/FrameData[3] Tile_X5Y11_LUT4AB/FrameData[4] Tile_X5Y11_LUT4AB/FrameData[5]
+ Tile_X5Y11_LUT4AB/FrameData[6] Tile_X5Y11_LUT4AB/FrameData[7] Tile_X5Y11_LUT4AB/FrameData[8]
+ Tile_X5Y11_LUT4AB/FrameData[9] Tile_X6Y11_LUT4AB/FrameData[0] Tile_X6Y11_LUT4AB/FrameData[10]
+ Tile_X6Y11_LUT4AB/FrameData[11] Tile_X6Y11_LUT4AB/FrameData[12] Tile_X6Y11_LUT4AB/FrameData[13]
+ Tile_X6Y11_LUT4AB/FrameData[14] Tile_X6Y11_LUT4AB/FrameData[15] Tile_X6Y11_LUT4AB/FrameData[16]
+ Tile_X6Y11_LUT4AB/FrameData[17] Tile_X6Y11_LUT4AB/FrameData[18] Tile_X6Y11_LUT4AB/FrameData[19]
+ Tile_X6Y11_LUT4AB/FrameData[1] Tile_X6Y11_LUT4AB/FrameData[20] Tile_X6Y11_LUT4AB/FrameData[21]
+ Tile_X6Y11_LUT4AB/FrameData[22] Tile_X6Y11_LUT4AB/FrameData[23] Tile_X6Y11_LUT4AB/FrameData[24]
+ Tile_X6Y11_LUT4AB/FrameData[25] Tile_X6Y11_LUT4AB/FrameData[26] Tile_X6Y11_LUT4AB/FrameData[27]
+ Tile_X6Y11_LUT4AB/FrameData[28] Tile_X6Y11_LUT4AB/FrameData[29] Tile_X6Y11_LUT4AB/FrameData[2]
+ Tile_X6Y11_LUT4AB/FrameData[30] Tile_X6Y11_LUT4AB/FrameData[31] Tile_X6Y11_LUT4AB/FrameData[3]
+ Tile_X6Y11_LUT4AB/FrameData[4] Tile_X6Y11_LUT4AB/FrameData[5] Tile_X6Y11_LUT4AB/FrameData[6]
+ Tile_X6Y11_LUT4AB/FrameData[7] Tile_X6Y11_LUT4AB/FrameData[8] Tile_X6Y11_LUT4AB/FrameData[9]
+ Tile_X5Y11_LUT4AB/FrameStrobe[0] Tile_X5Y11_LUT4AB/FrameStrobe[10] Tile_X5Y11_LUT4AB/FrameStrobe[11]
+ Tile_X5Y11_LUT4AB/FrameStrobe[12] Tile_X5Y11_LUT4AB/FrameStrobe[13] Tile_X5Y11_LUT4AB/FrameStrobe[14]
+ Tile_X5Y11_LUT4AB/FrameStrobe[15] Tile_X5Y11_LUT4AB/FrameStrobe[16] Tile_X5Y11_LUT4AB/FrameStrobe[17]
+ Tile_X5Y11_LUT4AB/FrameStrobe[18] Tile_X5Y11_LUT4AB/FrameStrobe[19] Tile_X5Y11_LUT4AB/FrameStrobe[1]
+ Tile_X5Y11_LUT4AB/FrameStrobe[2] Tile_X5Y11_LUT4AB/FrameStrobe[3] Tile_X5Y11_LUT4AB/FrameStrobe[4]
+ Tile_X5Y11_LUT4AB/FrameStrobe[5] Tile_X5Y11_LUT4AB/FrameStrobe[6] Tile_X5Y11_LUT4AB/FrameStrobe[7]
+ Tile_X5Y11_LUT4AB/FrameStrobe[8] Tile_X5Y11_LUT4AB/FrameStrobe[9] Tile_X5Y10_LUT4AB/FrameStrobe[0]
+ Tile_X5Y10_LUT4AB/FrameStrobe[10] Tile_X5Y10_LUT4AB/FrameStrobe[11] Tile_X5Y10_LUT4AB/FrameStrobe[12]
+ Tile_X5Y10_LUT4AB/FrameStrobe[13] Tile_X5Y10_LUT4AB/FrameStrobe[14] Tile_X5Y10_LUT4AB/FrameStrobe[15]
+ Tile_X5Y10_LUT4AB/FrameStrobe[16] Tile_X5Y10_LUT4AB/FrameStrobe[17] Tile_X5Y10_LUT4AB/FrameStrobe[18]
+ Tile_X5Y10_LUT4AB/FrameStrobe[19] Tile_X5Y10_LUT4AB/FrameStrobe[1] Tile_X5Y10_LUT4AB/FrameStrobe[2]
+ Tile_X5Y10_LUT4AB/FrameStrobe[3] Tile_X5Y10_LUT4AB/FrameStrobe[4] Tile_X5Y10_LUT4AB/FrameStrobe[5]
+ Tile_X5Y10_LUT4AB/FrameStrobe[6] Tile_X5Y10_LUT4AB/FrameStrobe[7] Tile_X5Y10_LUT4AB/FrameStrobe[8]
+ Tile_X5Y10_LUT4AB/FrameStrobe[9] Tile_X5Y11_LUT4AB/N1BEG[0] Tile_X5Y11_LUT4AB/N1BEG[1]
+ Tile_X5Y11_LUT4AB/N1BEG[2] Tile_X5Y11_LUT4AB/N1BEG[3] Tile_X5Y12_LUT4AB/N1BEG[0]
+ Tile_X5Y12_LUT4AB/N1BEG[1] Tile_X5Y12_LUT4AB/N1BEG[2] Tile_X5Y12_LUT4AB/N1BEG[3]
+ Tile_X5Y11_LUT4AB/N2BEG[0] Tile_X5Y11_LUT4AB/N2BEG[1] Tile_X5Y11_LUT4AB/N2BEG[2]
+ Tile_X5Y11_LUT4AB/N2BEG[3] Tile_X5Y11_LUT4AB/N2BEG[4] Tile_X5Y11_LUT4AB/N2BEG[5]
+ Tile_X5Y11_LUT4AB/N2BEG[6] Tile_X5Y11_LUT4AB/N2BEG[7] Tile_X5Y10_LUT4AB/N2END[0]
+ Tile_X5Y10_LUT4AB/N2END[1] Tile_X5Y10_LUT4AB/N2END[2] Tile_X5Y10_LUT4AB/N2END[3]
+ Tile_X5Y10_LUT4AB/N2END[4] Tile_X5Y10_LUT4AB/N2END[5] Tile_X5Y10_LUT4AB/N2END[6]
+ Tile_X5Y10_LUT4AB/N2END[7] Tile_X5Y11_LUT4AB/N2END[0] Tile_X5Y11_LUT4AB/N2END[1]
+ Tile_X5Y11_LUT4AB/N2END[2] Tile_X5Y11_LUT4AB/N2END[3] Tile_X5Y11_LUT4AB/N2END[4]
+ Tile_X5Y11_LUT4AB/N2END[5] Tile_X5Y11_LUT4AB/N2END[6] Tile_X5Y11_LUT4AB/N2END[7]
+ Tile_X5Y12_LUT4AB/N2BEG[0] Tile_X5Y12_LUT4AB/N2BEG[1] Tile_X5Y12_LUT4AB/N2BEG[2]
+ Tile_X5Y12_LUT4AB/N2BEG[3] Tile_X5Y12_LUT4AB/N2BEG[4] Tile_X5Y12_LUT4AB/N2BEG[5]
+ Tile_X5Y12_LUT4AB/N2BEG[6] Tile_X5Y12_LUT4AB/N2BEG[7] Tile_X5Y11_LUT4AB/N4BEG[0]
+ Tile_X5Y11_LUT4AB/N4BEG[10] Tile_X5Y11_LUT4AB/N4BEG[11] Tile_X5Y11_LUT4AB/N4BEG[12]
+ Tile_X5Y11_LUT4AB/N4BEG[13] Tile_X5Y11_LUT4AB/N4BEG[14] Tile_X5Y11_LUT4AB/N4BEG[15]
+ Tile_X5Y11_LUT4AB/N4BEG[1] Tile_X5Y11_LUT4AB/N4BEG[2] Tile_X5Y11_LUT4AB/N4BEG[3]
+ Tile_X5Y11_LUT4AB/N4BEG[4] Tile_X5Y11_LUT4AB/N4BEG[5] Tile_X5Y11_LUT4AB/N4BEG[6]
+ Tile_X5Y11_LUT4AB/N4BEG[7] Tile_X5Y11_LUT4AB/N4BEG[8] Tile_X5Y11_LUT4AB/N4BEG[9]
+ Tile_X5Y12_LUT4AB/N4BEG[0] Tile_X5Y12_LUT4AB/N4BEG[10] Tile_X5Y12_LUT4AB/N4BEG[11]
+ Tile_X5Y12_LUT4AB/N4BEG[12] Tile_X5Y12_LUT4AB/N4BEG[13] Tile_X5Y12_LUT4AB/N4BEG[14]
+ Tile_X5Y12_LUT4AB/N4BEG[15] Tile_X5Y12_LUT4AB/N4BEG[1] Tile_X5Y12_LUT4AB/N4BEG[2]
+ Tile_X5Y12_LUT4AB/N4BEG[3] Tile_X5Y12_LUT4AB/N4BEG[4] Tile_X5Y12_LUT4AB/N4BEG[5]
+ Tile_X5Y12_LUT4AB/N4BEG[6] Tile_X5Y12_LUT4AB/N4BEG[7] Tile_X5Y12_LUT4AB/N4BEG[8]
+ Tile_X5Y12_LUT4AB/N4BEG[9] Tile_X5Y11_LUT4AB/NN4BEG[0] Tile_X5Y11_LUT4AB/NN4BEG[10]
+ Tile_X5Y11_LUT4AB/NN4BEG[11] Tile_X5Y11_LUT4AB/NN4BEG[12] Tile_X5Y11_LUT4AB/NN4BEG[13]
+ Tile_X5Y11_LUT4AB/NN4BEG[14] Tile_X5Y11_LUT4AB/NN4BEG[15] Tile_X5Y11_LUT4AB/NN4BEG[1]
+ Tile_X5Y11_LUT4AB/NN4BEG[2] Tile_X5Y11_LUT4AB/NN4BEG[3] Tile_X5Y11_LUT4AB/NN4BEG[4]
+ Tile_X5Y11_LUT4AB/NN4BEG[5] Tile_X5Y11_LUT4AB/NN4BEG[6] Tile_X5Y11_LUT4AB/NN4BEG[7]
+ Tile_X5Y11_LUT4AB/NN4BEG[8] Tile_X5Y11_LUT4AB/NN4BEG[9] Tile_X5Y12_LUT4AB/NN4BEG[0]
+ Tile_X5Y12_LUT4AB/NN4BEG[10] Tile_X5Y12_LUT4AB/NN4BEG[11] Tile_X5Y12_LUT4AB/NN4BEG[12]
+ Tile_X5Y12_LUT4AB/NN4BEG[13] Tile_X5Y12_LUT4AB/NN4BEG[14] Tile_X5Y12_LUT4AB/NN4BEG[15]
+ Tile_X5Y12_LUT4AB/NN4BEG[1] Tile_X5Y12_LUT4AB/NN4BEG[2] Tile_X5Y12_LUT4AB/NN4BEG[3]
+ Tile_X5Y12_LUT4AB/NN4BEG[4] Tile_X5Y12_LUT4AB/NN4BEG[5] Tile_X5Y12_LUT4AB/NN4BEG[6]
+ Tile_X5Y12_LUT4AB/NN4BEG[7] Tile_X5Y12_LUT4AB/NN4BEG[8] Tile_X5Y12_LUT4AB/NN4BEG[9]
+ Tile_X5Y12_LUT4AB/S1END[0] Tile_X5Y12_LUT4AB/S1END[1] Tile_X5Y12_LUT4AB/S1END[2]
+ Tile_X5Y12_LUT4AB/S1END[3] Tile_X5Y11_LUT4AB/S1END[0] Tile_X5Y11_LUT4AB/S1END[1]
+ Tile_X5Y11_LUT4AB/S1END[2] Tile_X5Y11_LUT4AB/S1END[3] Tile_X5Y12_LUT4AB/S2MID[0]
+ Tile_X5Y12_LUT4AB/S2MID[1] Tile_X5Y12_LUT4AB/S2MID[2] Tile_X5Y12_LUT4AB/S2MID[3]
+ Tile_X5Y12_LUT4AB/S2MID[4] Tile_X5Y12_LUT4AB/S2MID[5] Tile_X5Y12_LUT4AB/S2MID[6]
+ Tile_X5Y12_LUT4AB/S2MID[7] Tile_X5Y12_LUT4AB/S2END[0] Tile_X5Y12_LUT4AB/S2END[1]
+ Tile_X5Y12_LUT4AB/S2END[2] Tile_X5Y12_LUT4AB/S2END[3] Tile_X5Y12_LUT4AB/S2END[4]
+ Tile_X5Y12_LUT4AB/S2END[5] Tile_X5Y12_LUT4AB/S2END[6] Tile_X5Y12_LUT4AB/S2END[7]
+ Tile_X5Y11_LUT4AB/S2END[0] Tile_X5Y11_LUT4AB/S2END[1] Tile_X5Y11_LUT4AB/S2END[2]
+ Tile_X5Y11_LUT4AB/S2END[3] Tile_X5Y11_LUT4AB/S2END[4] Tile_X5Y11_LUT4AB/S2END[5]
+ Tile_X5Y11_LUT4AB/S2END[6] Tile_X5Y11_LUT4AB/S2END[7] Tile_X5Y11_LUT4AB/S2MID[0]
+ Tile_X5Y11_LUT4AB/S2MID[1] Tile_X5Y11_LUT4AB/S2MID[2] Tile_X5Y11_LUT4AB/S2MID[3]
+ Tile_X5Y11_LUT4AB/S2MID[4] Tile_X5Y11_LUT4AB/S2MID[5] Tile_X5Y11_LUT4AB/S2MID[6]
+ Tile_X5Y11_LUT4AB/S2MID[7] Tile_X5Y12_LUT4AB/S4END[0] Tile_X5Y12_LUT4AB/S4END[10]
+ Tile_X5Y12_LUT4AB/S4END[11] Tile_X5Y12_LUT4AB/S4END[12] Tile_X5Y12_LUT4AB/S4END[13]
+ Tile_X5Y12_LUT4AB/S4END[14] Tile_X5Y12_LUT4AB/S4END[15] Tile_X5Y12_LUT4AB/S4END[1]
+ Tile_X5Y12_LUT4AB/S4END[2] Tile_X5Y12_LUT4AB/S4END[3] Tile_X5Y12_LUT4AB/S4END[4]
+ Tile_X5Y12_LUT4AB/S4END[5] Tile_X5Y12_LUT4AB/S4END[6] Tile_X5Y12_LUT4AB/S4END[7]
+ Tile_X5Y12_LUT4AB/S4END[8] Tile_X5Y12_LUT4AB/S4END[9] Tile_X5Y11_LUT4AB/S4END[0]
+ Tile_X5Y11_LUT4AB/S4END[10] Tile_X5Y11_LUT4AB/S4END[11] Tile_X5Y11_LUT4AB/S4END[12]
+ Tile_X5Y11_LUT4AB/S4END[13] Tile_X5Y11_LUT4AB/S4END[14] Tile_X5Y11_LUT4AB/S4END[15]
+ Tile_X5Y11_LUT4AB/S4END[1] Tile_X5Y11_LUT4AB/S4END[2] Tile_X5Y11_LUT4AB/S4END[3]
+ Tile_X5Y11_LUT4AB/S4END[4] Tile_X5Y11_LUT4AB/S4END[5] Tile_X5Y11_LUT4AB/S4END[6]
+ Tile_X5Y11_LUT4AB/S4END[7] Tile_X5Y11_LUT4AB/S4END[8] Tile_X5Y11_LUT4AB/S4END[9]
+ Tile_X5Y12_LUT4AB/SS4END[0] Tile_X5Y12_LUT4AB/SS4END[10] Tile_X5Y12_LUT4AB/SS4END[11]
+ Tile_X5Y12_LUT4AB/SS4END[12] Tile_X5Y12_LUT4AB/SS4END[13] Tile_X5Y12_LUT4AB/SS4END[14]
+ Tile_X5Y12_LUT4AB/SS4END[15] Tile_X5Y12_LUT4AB/SS4END[1] Tile_X5Y12_LUT4AB/SS4END[2]
+ Tile_X5Y12_LUT4AB/SS4END[3] Tile_X5Y12_LUT4AB/SS4END[4] Tile_X5Y12_LUT4AB/SS4END[5]
+ Tile_X5Y12_LUT4AB/SS4END[6] Tile_X5Y12_LUT4AB/SS4END[7] Tile_X5Y12_LUT4AB/SS4END[8]
+ Tile_X5Y12_LUT4AB/SS4END[9] Tile_X5Y11_LUT4AB/SS4END[0] Tile_X5Y11_LUT4AB/SS4END[10]
+ Tile_X5Y11_LUT4AB/SS4END[11] Tile_X5Y11_LUT4AB/SS4END[12] Tile_X5Y11_LUT4AB/SS4END[13]
+ Tile_X5Y11_LUT4AB/SS4END[14] Tile_X5Y11_LUT4AB/SS4END[15] Tile_X5Y11_LUT4AB/SS4END[1]
+ Tile_X5Y11_LUT4AB/SS4END[2] Tile_X5Y11_LUT4AB/SS4END[3] Tile_X5Y11_LUT4AB/SS4END[4]
+ Tile_X5Y11_LUT4AB/SS4END[5] Tile_X5Y11_LUT4AB/SS4END[6] Tile_X5Y11_LUT4AB/SS4END[7]
+ Tile_X5Y11_LUT4AB/SS4END[8] Tile_X5Y11_LUT4AB/SS4END[9] Tile_X5Y11_LUT4AB/UserCLK
+ Tile_X5Y10_LUT4AB/UserCLK VGND VPWR Tile_X5Y11_LUT4AB/W1BEG[0] Tile_X5Y11_LUT4AB/W1BEG[1]
+ Tile_X5Y11_LUT4AB/W1BEG[2] Tile_X5Y11_LUT4AB/W1BEG[3] Tile_X6Y11_LUT4AB/W1BEG[0]
+ Tile_X6Y11_LUT4AB/W1BEG[1] Tile_X6Y11_LUT4AB/W1BEG[2] Tile_X6Y11_LUT4AB/W1BEG[3]
+ Tile_X5Y11_LUT4AB/W2BEG[0] Tile_X5Y11_LUT4AB/W2BEG[1] Tile_X5Y11_LUT4AB/W2BEG[2]
+ Tile_X5Y11_LUT4AB/W2BEG[3] Tile_X5Y11_LUT4AB/W2BEG[4] Tile_X5Y11_LUT4AB/W2BEG[5]
+ Tile_X5Y11_LUT4AB/W2BEG[6] Tile_X5Y11_LUT4AB/W2BEG[7] Tile_X5Y11_LUT4AB/W2BEGb[0]
+ Tile_X5Y11_LUT4AB/W2BEGb[1] Tile_X5Y11_LUT4AB/W2BEGb[2] Tile_X5Y11_LUT4AB/W2BEGb[3]
+ Tile_X5Y11_LUT4AB/W2BEGb[4] Tile_X5Y11_LUT4AB/W2BEGb[5] Tile_X5Y11_LUT4AB/W2BEGb[6]
+ Tile_X5Y11_LUT4AB/W2BEGb[7] Tile_X5Y11_LUT4AB/W2END[0] Tile_X5Y11_LUT4AB/W2END[1]
+ Tile_X5Y11_LUT4AB/W2END[2] Tile_X5Y11_LUT4AB/W2END[3] Tile_X5Y11_LUT4AB/W2END[4]
+ Tile_X5Y11_LUT4AB/W2END[5] Tile_X5Y11_LUT4AB/W2END[6] Tile_X5Y11_LUT4AB/W2END[7]
+ Tile_X6Y11_LUT4AB/W2BEG[0] Tile_X6Y11_LUT4AB/W2BEG[1] Tile_X6Y11_LUT4AB/W2BEG[2]
+ Tile_X6Y11_LUT4AB/W2BEG[3] Tile_X6Y11_LUT4AB/W2BEG[4] Tile_X6Y11_LUT4AB/W2BEG[5]
+ Tile_X6Y11_LUT4AB/W2BEG[6] Tile_X6Y11_LUT4AB/W2BEG[7] Tile_X5Y11_LUT4AB/W6BEG[0]
+ Tile_X5Y11_LUT4AB/W6BEG[10] Tile_X5Y11_LUT4AB/W6BEG[11] Tile_X5Y11_LUT4AB/W6BEG[1]
+ Tile_X5Y11_LUT4AB/W6BEG[2] Tile_X5Y11_LUT4AB/W6BEG[3] Tile_X5Y11_LUT4AB/W6BEG[4]
+ Tile_X5Y11_LUT4AB/W6BEG[5] Tile_X5Y11_LUT4AB/W6BEG[6] Tile_X5Y11_LUT4AB/W6BEG[7]
+ Tile_X5Y11_LUT4AB/W6BEG[8] Tile_X5Y11_LUT4AB/W6BEG[9] Tile_X6Y11_LUT4AB/W6BEG[0]
+ Tile_X6Y11_LUT4AB/W6BEG[10] Tile_X6Y11_LUT4AB/W6BEG[11] Tile_X6Y11_LUT4AB/W6BEG[1]
+ Tile_X6Y11_LUT4AB/W6BEG[2] Tile_X6Y11_LUT4AB/W6BEG[3] Tile_X6Y11_LUT4AB/W6BEG[4]
+ Tile_X6Y11_LUT4AB/W6BEG[5] Tile_X6Y11_LUT4AB/W6BEG[6] Tile_X6Y11_LUT4AB/W6BEG[7]
+ Tile_X6Y11_LUT4AB/W6BEG[8] Tile_X6Y11_LUT4AB/W6BEG[9] Tile_X5Y11_LUT4AB/WW4BEG[0]
+ Tile_X5Y11_LUT4AB/WW4BEG[10] Tile_X5Y11_LUT4AB/WW4BEG[11] Tile_X5Y11_LUT4AB/WW4BEG[12]
+ Tile_X5Y11_LUT4AB/WW4BEG[13] Tile_X5Y11_LUT4AB/WW4BEG[14] Tile_X5Y11_LUT4AB/WW4BEG[15]
+ Tile_X5Y11_LUT4AB/WW4BEG[1] Tile_X5Y11_LUT4AB/WW4BEG[2] Tile_X5Y11_LUT4AB/WW4BEG[3]
+ Tile_X5Y11_LUT4AB/WW4BEG[4] Tile_X5Y11_LUT4AB/WW4BEG[5] Tile_X5Y11_LUT4AB/WW4BEG[6]
+ Tile_X5Y11_LUT4AB/WW4BEG[7] Tile_X5Y11_LUT4AB/WW4BEG[8] Tile_X5Y11_LUT4AB/WW4BEG[9]
+ Tile_X6Y11_LUT4AB/WW4BEG[0] Tile_X6Y11_LUT4AB/WW4BEG[10] Tile_X6Y11_LUT4AB/WW4BEG[11]
+ Tile_X6Y11_LUT4AB/WW4BEG[12] Tile_X6Y11_LUT4AB/WW4BEG[13] Tile_X6Y11_LUT4AB/WW4BEG[14]
+ Tile_X6Y11_LUT4AB/WW4BEG[15] Tile_X6Y11_LUT4AB/WW4BEG[1] Tile_X6Y11_LUT4AB/WW4BEG[2]
+ Tile_X6Y11_LUT4AB/WW4BEG[3] Tile_X6Y11_LUT4AB/WW4BEG[4] Tile_X6Y11_LUT4AB/WW4BEG[5]
+ Tile_X6Y11_LUT4AB/WW4BEG[6] Tile_X6Y11_LUT4AB/WW4BEG[7] Tile_X6Y11_LUT4AB/WW4BEG[8]
+ Tile_X6Y11_LUT4AB/WW4BEG[9] LUT4AB
XTile_X1Y9_LUT4AB Tile_X1Y9_LUT4AB/Ci Tile_X1Y9_LUT4AB/Co Tile_X2Y9_LUT4AB/E1END[0]
+ Tile_X2Y9_LUT4AB/E1END[1] Tile_X2Y9_LUT4AB/E1END[2] Tile_X2Y9_LUT4AB/E1END[3] Tile_X0Y9_W_IO/E1BEG[0]
+ Tile_X0Y9_W_IO/E1BEG[1] Tile_X0Y9_W_IO/E1BEG[2] Tile_X0Y9_W_IO/E1BEG[3] Tile_X2Y9_LUT4AB/E2MID[0]
+ Tile_X2Y9_LUT4AB/E2MID[1] Tile_X2Y9_LUT4AB/E2MID[2] Tile_X2Y9_LUT4AB/E2MID[3] Tile_X2Y9_LUT4AB/E2MID[4]
+ Tile_X2Y9_LUT4AB/E2MID[5] Tile_X2Y9_LUT4AB/E2MID[6] Tile_X2Y9_LUT4AB/E2MID[7] Tile_X2Y9_LUT4AB/E2END[0]
+ Tile_X2Y9_LUT4AB/E2END[1] Tile_X2Y9_LUT4AB/E2END[2] Tile_X2Y9_LUT4AB/E2END[3] Tile_X2Y9_LUT4AB/E2END[4]
+ Tile_X2Y9_LUT4AB/E2END[5] Tile_X2Y9_LUT4AB/E2END[6] Tile_X2Y9_LUT4AB/E2END[7] Tile_X0Y9_W_IO/E2BEGb[0]
+ Tile_X0Y9_W_IO/E2BEGb[1] Tile_X0Y9_W_IO/E2BEGb[2] Tile_X0Y9_W_IO/E2BEGb[3] Tile_X0Y9_W_IO/E2BEGb[4]
+ Tile_X0Y9_W_IO/E2BEGb[5] Tile_X0Y9_W_IO/E2BEGb[6] Tile_X0Y9_W_IO/E2BEGb[7] Tile_X0Y9_W_IO/E2BEG[0]
+ Tile_X0Y9_W_IO/E2BEG[1] Tile_X0Y9_W_IO/E2BEG[2] Tile_X0Y9_W_IO/E2BEG[3] Tile_X0Y9_W_IO/E2BEG[4]
+ Tile_X0Y9_W_IO/E2BEG[5] Tile_X0Y9_W_IO/E2BEG[6] Tile_X0Y9_W_IO/E2BEG[7] Tile_X2Y9_LUT4AB/E6END[0]
+ Tile_X2Y9_LUT4AB/E6END[10] Tile_X2Y9_LUT4AB/E6END[11] Tile_X2Y9_LUT4AB/E6END[1]
+ Tile_X2Y9_LUT4AB/E6END[2] Tile_X2Y9_LUT4AB/E6END[3] Tile_X2Y9_LUT4AB/E6END[4] Tile_X2Y9_LUT4AB/E6END[5]
+ Tile_X2Y9_LUT4AB/E6END[6] Tile_X2Y9_LUT4AB/E6END[7] Tile_X2Y9_LUT4AB/E6END[8] Tile_X2Y9_LUT4AB/E6END[9]
+ Tile_X0Y9_W_IO/E6BEG[0] Tile_X0Y9_W_IO/E6BEG[10] Tile_X0Y9_W_IO/E6BEG[11] Tile_X0Y9_W_IO/E6BEG[1]
+ Tile_X0Y9_W_IO/E6BEG[2] Tile_X0Y9_W_IO/E6BEG[3] Tile_X0Y9_W_IO/E6BEG[4] Tile_X0Y9_W_IO/E6BEG[5]
+ Tile_X0Y9_W_IO/E6BEG[6] Tile_X0Y9_W_IO/E6BEG[7] Tile_X0Y9_W_IO/E6BEG[8] Tile_X0Y9_W_IO/E6BEG[9]
+ Tile_X2Y9_LUT4AB/EE4END[0] Tile_X2Y9_LUT4AB/EE4END[10] Tile_X2Y9_LUT4AB/EE4END[11]
+ Tile_X2Y9_LUT4AB/EE4END[12] Tile_X2Y9_LUT4AB/EE4END[13] Tile_X2Y9_LUT4AB/EE4END[14]
+ Tile_X2Y9_LUT4AB/EE4END[15] Tile_X2Y9_LUT4AB/EE4END[1] Tile_X2Y9_LUT4AB/EE4END[2]
+ Tile_X2Y9_LUT4AB/EE4END[3] Tile_X2Y9_LUT4AB/EE4END[4] Tile_X2Y9_LUT4AB/EE4END[5]
+ Tile_X2Y9_LUT4AB/EE4END[6] Tile_X2Y9_LUT4AB/EE4END[7] Tile_X2Y9_LUT4AB/EE4END[8]
+ Tile_X2Y9_LUT4AB/EE4END[9] Tile_X0Y9_W_IO/EE4BEG[0] Tile_X0Y9_W_IO/EE4BEG[10] Tile_X0Y9_W_IO/EE4BEG[11]
+ Tile_X0Y9_W_IO/EE4BEG[12] Tile_X0Y9_W_IO/EE4BEG[13] Tile_X0Y9_W_IO/EE4BEG[14] Tile_X0Y9_W_IO/EE4BEG[15]
+ Tile_X0Y9_W_IO/EE4BEG[1] Tile_X0Y9_W_IO/EE4BEG[2] Tile_X0Y9_W_IO/EE4BEG[3] Tile_X0Y9_W_IO/EE4BEG[4]
+ Tile_X0Y9_W_IO/EE4BEG[5] Tile_X0Y9_W_IO/EE4BEG[6] Tile_X0Y9_W_IO/EE4BEG[7] Tile_X0Y9_W_IO/EE4BEG[8]
+ Tile_X0Y9_W_IO/EE4BEG[9] Tile_X1Y9_LUT4AB/FrameData[0] Tile_X1Y9_LUT4AB/FrameData[10]
+ Tile_X1Y9_LUT4AB/FrameData[11] Tile_X1Y9_LUT4AB/FrameData[12] Tile_X1Y9_LUT4AB/FrameData[13]
+ Tile_X1Y9_LUT4AB/FrameData[14] Tile_X1Y9_LUT4AB/FrameData[15] Tile_X1Y9_LUT4AB/FrameData[16]
+ Tile_X1Y9_LUT4AB/FrameData[17] Tile_X1Y9_LUT4AB/FrameData[18] Tile_X1Y9_LUT4AB/FrameData[19]
+ Tile_X1Y9_LUT4AB/FrameData[1] Tile_X1Y9_LUT4AB/FrameData[20] Tile_X1Y9_LUT4AB/FrameData[21]
+ Tile_X1Y9_LUT4AB/FrameData[22] Tile_X1Y9_LUT4AB/FrameData[23] Tile_X1Y9_LUT4AB/FrameData[24]
+ Tile_X1Y9_LUT4AB/FrameData[25] Tile_X1Y9_LUT4AB/FrameData[26] Tile_X1Y9_LUT4AB/FrameData[27]
+ Tile_X1Y9_LUT4AB/FrameData[28] Tile_X1Y9_LUT4AB/FrameData[29] Tile_X1Y9_LUT4AB/FrameData[2]
+ Tile_X1Y9_LUT4AB/FrameData[30] Tile_X1Y9_LUT4AB/FrameData[31] Tile_X1Y9_LUT4AB/FrameData[3]
+ Tile_X1Y9_LUT4AB/FrameData[4] Tile_X1Y9_LUT4AB/FrameData[5] Tile_X1Y9_LUT4AB/FrameData[6]
+ Tile_X1Y9_LUT4AB/FrameData[7] Tile_X1Y9_LUT4AB/FrameData[8] Tile_X1Y9_LUT4AB/FrameData[9]
+ Tile_X2Y9_LUT4AB/FrameData[0] Tile_X2Y9_LUT4AB/FrameData[10] Tile_X2Y9_LUT4AB/FrameData[11]
+ Tile_X2Y9_LUT4AB/FrameData[12] Tile_X2Y9_LUT4AB/FrameData[13] Tile_X2Y9_LUT4AB/FrameData[14]
+ Tile_X2Y9_LUT4AB/FrameData[15] Tile_X2Y9_LUT4AB/FrameData[16] Tile_X2Y9_LUT4AB/FrameData[17]
+ Tile_X2Y9_LUT4AB/FrameData[18] Tile_X2Y9_LUT4AB/FrameData[19] Tile_X2Y9_LUT4AB/FrameData[1]
+ Tile_X2Y9_LUT4AB/FrameData[20] Tile_X2Y9_LUT4AB/FrameData[21] Tile_X2Y9_LUT4AB/FrameData[22]
+ Tile_X2Y9_LUT4AB/FrameData[23] Tile_X2Y9_LUT4AB/FrameData[24] Tile_X2Y9_LUT4AB/FrameData[25]
+ Tile_X2Y9_LUT4AB/FrameData[26] Tile_X2Y9_LUT4AB/FrameData[27] Tile_X2Y9_LUT4AB/FrameData[28]
+ Tile_X2Y9_LUT4AB/FrameData[29] Tile_X2Y9_LUT4AB/FrameData[2] Tile_X2Y9_LUT4AB/FrameData[30]
+ Tile_X2Y9_LUT4AB/FrameData[31] Tile_X2Y9_LUT4AB/FrameData[3] Tile_X2Y9_LUT4AB/FrameData[4]
+ Tile_X2Y9_LUT4AB/FrameData[5] Tile_X2Y9_LUT4AB/FrameData[6] Tile_X2Y9_LUT4AB/FrameData[7]
+ Tile_X2Y9_LUT4AB/FrameData[8] Tile_X2Y9_LUT4AB/FrameData[9] Tile_X1Y9_LUT4AB/FrameStrobe[0]
+ Tile_X1Y9_LUT4AB/FrameStrobe[10] Tile_X1Y9_LUT4AB/FrameStrobe[11] Tile_X1Y9_LUT4AB/FrameStrobe[12]
+ Tile_X1Y9_LUT4AB/FrameStrobe[13] Tile_X1Y9_LUT4AB/FrameStrobe[14] Tile_X1Y9_LUT4AB/FrameStrobe[15]
+ Tile_X1Y9_LUT4AB/FrameStrobe[16] Tile_X1Y9_LUT4AB/FrameStrobe[17] Tile_X1Y9_LUT4AB/FrameStrobe[18]
+ Tile_X1Y9_LUT4AB/FrameStrobe[19] Tile_X1Y9_LUT4AB/FrameStrobe[1] Tile_X1Y9_LUT4AB/FrameStrobe[2]
+ Tile_X1Y9_LUT4AB/FrameStrobe[3] Tile_X1Y9_LUT4AB/FrameStrobe[4] Tile_X1Y9_LUT4AB/FrameStrobe[5]
+ Tile_X1Y9_LUT4AB/FrameStrobe[6] Tile_X1Y9_LUT4AB/FrameStrobe[7] Tile_X1Y9_LUT4AB/FrameStrobe[8]
+ Tile_X1Y9_LUT4AB/FrameStrobe[9] Tile_X1Y8_LUT4AB/FrameStrobe[0] Tile_X1Y8_LUT4AB/FrameStrobe[10]
+ Tile_X1Y8_LUT4AB/FrameStrobe[11] Tile_X1Y8_LUT4AB/FrameStrobe[12] Tile_X1Y8_LUT4AB/FrameStrobe[13]
+ Tile_X1Y8_LUT4AB/FrameStrobe[14] Tile_X1Y8_LUT4AB/FrameStrobe[15] Tile_X1Y8_LUT4AB/FrameStrobe[16]
+ Tile_X1Y8_LUT4AB/FrameStrobe[17] Tile_X1Y8_LUT4AB/FrameStrobe[18] Tile_X1Y8_LUT4AB/FrameStrobe[19]
+ Tile_X1Y8_LUT4AB/FrameStrobe[1] Tile_X1Y8_LUT4AB/FrameStrobe[2] Tile_X1Y8_LUT4AB/FrameStrobe[3]
+ Tile_X1Y8_LUT4AB/FrameStrobe[4] Tile_X1Y8_LUT4AB/FrameStrobe[5] Tile_X1Y8_LUT4AB/FrameStrobe[6]
+ Tile_X1Y8_LUT4AB/FrameStrobe[7] Tile_X1Y8_LUT4AB/FrameStrobe[8] Tile_X1Y8_LUT4AB/FrameStrobe[9]
+ Tile_X1Y9_LUT4AB/N1BEG[0] Tile_X1Y9_LUT4AB/N1BEG[1] Tile_X1Y9_LUT4AB/N1BEG[2] Tile_X1Y9_LUT4AB/N1BEG[3]
+ Tile_X1Y9_LUT4AB/N1END[0] Tile_X1Y9_LUT4AB/N1END[1] Tile_X1Y9_LUT4AB/N1END[2] Tile_X1Y9_LUT4AB/N1END[3]
+ Tile_X1Y9_LUT4AB/N2BEG[0] Tile_X1Y9_LUT4AB/N2BEG[1] Tile_X1Y9_LUT4AB/N2BEG[2] Tile_X1Y9_LUT4AB/N2BEG[3]
+ Tile_X1Y9_LUT4AB/N2BEG[4] Tile_X1Y9_LUT4AB/N2BEG[5] Tile_X1Y9_LUT4AB/N2BEG[6] Tile_X1Y9_LUT4AB/N2BEG[7]
+ Tile_X1Y8_LUT4AB/N2END[0] Tile_X1Y8_LUT4AB/N2END[1] Tile_X1Y8_LUT4AB/N2END[2] Tile_X1Y8_LUT4AB/N2END[3]
+ Tile_X1Y8_LUT4AB/N2END[4] Tile_X1Y8_LUT4AB/N2END[5] Tile_X1Y8_LUT4AB/N2END[6] Tile_X1Y8_LUT4AB/N2END[7]
+ Tile_X1Y9_LUT4AB/N2END[0] Tile_X1Y9_LUT4AB/N2END[1] Tile_X1Y9_LUT4AB/N2END[2] Tile_X1Y9_LUT4AB/N2END[3]
+ Tile_X1Y9_LUT4AB/N2END[4] Tile_X1Y9_LUT4AB/N2END[5] Tile_X1Y9_LUT4AB/N2END[6] Tile_X1Y9_LUT4AB/N2END[7]
+ Tile_X1Y9_LUT4AB/N2MID[0] Tile_X1Y9_LUT4AB/N2MID[1] Tile_X1Y9_LUT4AB/N2MID[2] Tile_X1Y9_LUT4AB/N2MID[3]
+ Tile_X1Y9_LUT4AB/N2MID[4] Tile_X1Y9_LUT4AB/N2MID[5] Tile_X1Y9_LUT4AB/N2MID[6] Tile_X1Y9_LUT4AB/N2MID[7]
+ Tile_X1Y9_LUT4AB/N4BEG[0] Tile_X1Y9_LUT4AB/N4BEG[10] Tile_X1Y9_LUT4AB/N4BEG[11]
+ Tile_X1Y9_LUT4AB/N4BEG[12] Tile_X1Y9_LUT4AB/N4BEG[13] Tile_X1Y9_LUT4AB/N4BEG[14]
+ Tile_X1Y9_LUT4AB/N4BEG[15] Tile_X1Y9_LUT4AB/N4BEG[1] Tile_X1Y9_LUT4AB/N4BEG[2] Tile_X1Y9_LUT4AB/N4BEG[3]
+ Tile_X1Y9_LUT4AB/N4BEG[4] Tile_X1Y9_LUT4AB/N4BEG[5] Tile_X1Y9_LUT4AB/N4BEG[6] Tile_X1Y9_LUT4AB/N4BEG[7]
+ Tile_X1Y9_LUT4AB/N4BEG[8] Tile_X1Y9_LUT4AB/N4BEG[9] Tile_X1Y9_LUT4AB/N4END[0] Tile_X1Y9_LUT4AB/N4END[10]
+ Tile_X1Y9_LUT4AB/N4END[11] Tile_X1Y9_LUT4AB/N4END[12] Tile_X1Y9_LUT4AB/N4END[13]
+ Tile_X1Y9_LUT4AB/N4END[14] Tile_X1Y9_LUT4AB/N4END[15] Tile_X1Y9_LUT4AB/N4END[1]
+ Tile_X1Y9_LUT4AB/N4END[2] Tile_X1Y9_LUT4AB/N4END[3] Tile_X1Y9_LUT4AB/N4END[4] Tile_X1Y9_LUT4AB/N4END[5]
+ Tile_X1Y9_LUT4AB/N4END[6] Tile_X1Y9_LUT4AB/N4END[7] Tile_X1Y9_LUT4AB/N4END[8] Tile_X1Y9_LUT4AB/N4END[9]
+ Tile_X1Y9_LUT4AB/NN4BEG[0] Tile_X1Y9_LUT4AB/NN4BEG[10] Tile_X1Y9_LUT4AB/NN4BEG[11]
+ Tile_X1Y9_LUT4AB/NN4BEG[12] Tile_X1Y9_LUT4AB/NN4BEG[13] Tile_X1Y9_LUT4AB/NN4BEG[14]
+ Tile_X1Y9_LUT4AB/NN4BEG[15] Tile_X1Y9_LUT4AB/NN4BEG[1] Tile_X1Y9_LUT4AB/NN4BEG[2]
+ Tile_X1Y9_LUT4AB/NN4BEG[3] Tile_X1Y9_LUT4AB/NN4BEG[4] Tile_X1Y9_LUT4AB/NN4BEG[5]
+ Tile_X1Y9_LUT4AB/NN4BEG[6] Tile_X1Y9_LUT4AB/NN4BEG[7] Tile_X1Y9_LUT4AB/NN4BEG[8]
+ Tile_X1Y9_LUT4AB/NN4BEG[9] Tile_X1Y9_LUT4AB/NN4END[0] Tile_X1Y9_LUT4AB/NN4END[10]
+ Tile_X1Y9_LUT4AB/NN4END[11] Tile_X1Y9_LUT4AB/NN4END[12] Tile_X1Y9_LUT4AB/NN4END[13]
+ Tile_X1Y9_LUT4AB/NN4END[14] Tile_X1Y9_LUT4AB/NN4END[15] Tile_X1Y9_LUT4AB/NN4END[1]
+ Tile_X1Y9_LUT4AB/NN4END[2] Tile_X1Y9_LUT4AB/NN4END[3] Tile_X1Y9_LUT4AB/NN4END[4]
+ Tile_X1Y9_LUT4AB/NN4END[5] Tile_X1Y9_LUT4AB/NN4END[6] Tile_X1Y9_LUT4AB/NN4END[7]
+ Tile_X1Y9_LUT4AB/NN4END[8] Tile_X1Y9_LUT4AB/NN4END[9] Tile_X1Y9_LUT4AB/S1BEG[0]
+ Tile_X1Y9_LUT4AB/S1BEG[1] Tile_X1Y9_LUT4AB/S1BEG[2] Tile_X1Y9_LUT4AB/S1BEG[3] Tile_X1Y9_LUT4AB/S1END[0]
+ Tile_X1Y9_LUT4AB/S1END[1] Tile_X1Y9_LUT4AB/S1END[2] Tile_X1Y9_LUT4AB/S1END[3] Tile_X1Y9_LUT4AB/S2BEG[0]
+ Tile_X1Y9_LUT4AB/S2BEG[1] Tile_X1Y9_LUT4AB/S2BEG[2] Tile_X1Y9_LUT4AB/S2BEG[3] Tile_X1Y9_LUT4AB/S2BEG[4]
+ Tile_X1Y9_LUT4AB/S2BEG[5] Tile_X1Y9_LUT4AB/S2BEG[6] Tile_X1Y9_LUT4AB/S2BEG[7] Tile_X1Y9_LUT4AB/S2BEGb[0]
+ Tile_X1Y9_LUT4AB/S2BEGb[1] Tile_X1Y9_LUT4AB/S2BEGb[2] Tile_X1Y9_LUT4AB/S2BEGb[3]
+ Tile_X1Y9_LUT4AB/S2BEGb[4] Tile_X1Y9_LUT4AB/S2BEGb[5] Tile_X1Y9_LUT4AB/S2BEGb[6]
+ Tile_X1Y9_LUT4AB/S2BEGb[7] Tile_X1Y9_LUT4AB/S2END[0] Tile_X1Y9_LUT4AB/S2END[1] Tile_X1Y9_LUT4AB/S2END[2]
+ Tile_X1Y9_LUT4AB/S2END[3] Tile_X1Y9_LUT4AB/S2END[4] Tile_X1Y9_LUT4AB/S2END[5] Tile_X1Y9_LUT4AB/S2END[6]
+ Tile_X1Y9_LUT4AB/S2END[7] Tile_X1Y9_LUT4AB/S2MID[0] Tile_X1Y9_LUT4AB/S2MID[1] Tile_X1Y9_LUT4AB/S2MID[2]
+ Tile_X1Y9_LUT4AB/S2MID[3] Tile_X1Y9_LUT4AB/S2MID[4] Tile_X1Y9_LUT4AB/S2MID[5] Tile_X1Y9_LUT4AB/S2MID[6]
+ Tile_X1Y9_LUT4AB/S2MID[7] Tile_X1Y9_LUT4AB/S4BEG[0] Tile_X1Y9_LUT4AB/S4BEG[10] Tile_X1Y9_LUT4AB/S4BEG[11]
+ Tile_X1Y9_LUT4AB/S4BEG[12] Tile_X1Y9_LUT4AB/S4BEG[13] Tile_X1Y9_LUT4AB/S4BEG[14]
+ Tile_X1Y9_LUT4AB/S4BEG[15] Tile_X1Y9_LUT4AB/S4BEG[1] Tile_X1Y9_LUT4AB/S4BEG[2] Tile_X1Y9_LUT4AB/S4BEG[3]
+ Tile_X1Y9_LUT4AB/S4BEG[4] Tile_X1Y9_LUT4AB/S4BEG[5] Tile_X1Y9_LUT4AB/S4BEG[6] Tile_X1Y9_LUT4AB/S4BEG[7]
+ Tile_X1Y9_LUT4AB/S4BEG[8] Tile_X1Y9_LUT4AB/S4BEG[9] Tile_X1Y9_LUT4AB/S4END[0] Tile_X1Y9_LUT4AB/S4END[10]
+ Tile_X1Y9_LUT4AB/S4END[11] Tile_X1Y9_LUT4AB/S4END[12] Tile_X1Y9_LUT4AB/S4END[13]
+ Tile_X1Y9_LUT4AB/S4END[14] Tile_X1Y9_LUT4AB/S4END[15] Tile_X1Y9_LUT4AB/S4END[1]
+ Tile_X1Y9_LUT4AB/S4END[2] Tile_X1Y9_LUT4AB/S4END[3] Tile_X1Y9_LUT4AB/S4END[4] Tile_X1Y9_LUT4AB/S4END[5]
+ Tile_X1Y9_LUT4AB/S4END[6] Tile_X1Y9_LUT4AB/S4END[7] Tile_X1Y9_LUT4AB/S4END[8] Tile_X1Y9_LUT4AB/S4END[9]
+ Tile_X1Y9_LUT4AB/SS4BEG[0] Tile_X1Y9_LUT4AB/SS4BEG[10] Tile_X1Y9_LUT4AB/SS4BEG[11]
+ Tile_X1Y9_LUT4AB/SS4BEG[12] Tile_X1Y9_LUT4AB/SS4BEG[13] Tile_X1Y9_LUT4AB/SS4BEG[14]
+ Tile_X1Y9_LUT4AB/SS4BEG[15] Tile_X1Y9_LUT4AB/SS4BEG[1] Tile_X1Y9_LUT4AB/SS4BEG[2]
+ Tile_X1Y9_LUT4AB/SS4BEG[3] Tile_X1Y9_LUT4AB/SS4BEG[4] Tile_X1Y9_LUT4AB/SS4BEG[5]
+ Tile_X1Y9_LUT4AB/SS4BEG[6] Tile_X1Y9_LUT4AB/SS4BEG[7] Tile_X1Y9_LUT4AB/SS4BEG[8]
+ Tile_X1Y9_LUT4AB/SS4BEG[9] Tile_X1Y9_LUT4AB/SS4END[0] Tile_X1Y9_LUT4AB/SS4END[10]
+ Tile_X1Y9_LUT4AB/SS4END[11] Tile_X1Y9_LUT4AB/SS4END[12] Tile_X1Y9_LUT4AB/SS4END[13]
+ Tile_X1Y9_LUT4AB/SS4END[14] Tile_X1Y9_LUT4AB/SS4END[15] Tile_X1Y9_LUT4AB/SS4END[1]
+ Tile_X1Y9_LUT4AB/SS4END[2] Tile_X1Y9_LUT4AB/SS4END[3] Tile_X1Y9_LUT4AB/SS4END[4]
+ Tile_X1Y9_LUT4AB/SS4END[5] Tile_X1Y9_LUT4AB/SS4END[6] Tile_X1Y9_LUT4AB/SS4END[7]
+ Tile_X1Y9_LUT4AB/SS4END[8] Tile_X1Y9_LUT4AB/SS4END[9] Tile_X1Y9_LUT4AB/UserCLK Tile_X1Y8_LUT4AB/UserCLK
+ VGND VPWR Tile_X0Y9_W_IO/W1END[0] Tile_X0Y9_W_IO/W1END[1] Tile_X0Y9_W_IO/W1END[2]
+ Tile_X0Y9_W_IO/W1END[3] Tile_X2Y9_LUT4AB/W1BEG[0] Tile_X2Y9_LUT4AB/W1BEG[1] Tile_X2Y9_LUT4AB/W1BEG[2]
+ Tile_X2Y9_LUT4AB/W1BEG[3] Tile_X0Y9_W_IO/W2MID[0] Tile_X0Y9_W_IO/W2MID[1] Tile_X0Y9_W_IO/W2MID[2]
+ Tile_X0Y9_W_IO/W2MID[3] Tile_X0Y9_W_IO/W2MID[4] Tile_X0Y9_W_IO/W2MID[5] Tile_X0Y9_W_IO/W2MID[6]
+ Tile_X0Y9_W_IO/W2MID[7] Tile_X0Y9_W_IO/W2END[0] Tile_X0Y9_W_IO/W2END[1] Tile_X0Y9_W_IO/W2END[2]
+ Tile_X0Y9_W_IO/W2END[3] Tile_X0Y9_W_IO/W2END[4] Tile_X0Y9_W_IO/W2END[5] Tile_X0Y9_W_IO/W2END[6]
+ Tile_X0Y9_W_IO/W2END[7] Tile_X1Y9_LUT4AB/W2END[0] Tile_X1Y9_LUT4AB/W2END[1] Tile_X1Y9_LUT4AB/W2END[2]
+ Tile_X1Y9_LUT4AB/W2END[3] Tile_X1Y9_LUT4AB/W2END[4] Tile_X1Y9_LUT4AB/W2END[5] Tile_X1Y9_LUT4AB/W2END[6]
+ Tile_X1Y9_LUT4AB/W2END[7] Tile_X2Y9_LUT4AB/W2BEG[0] Tile_X2Y9_LUT4AB/W2BEG[1] Tile_X2Y9_LUT4AB/W2BEG[2]
+ Tile_X2Y9_LUT4AB/W2BEG[3] Tile_X2Y9_LUT4AB/W2BEG[4] Tile_X2Y9_LUT4AB/W2BEG[5] Tile_X2Y9_LUT4AB/W2BEG[6]
+ Tile_X2Y9_LUT4AB/W2BEG[7] Tile_X0Y9_W_IO/W6END[0] Tile_X0Y9_W_IO/W6END[10] Tile_X0Y9_W_IO/W6END[11]
+ Tile_X0Y9_W_IO/W6END[1] Tile_X0Y9_W_IO/W6END[2] Tile_X0Y9_W_IO/W6END[3] Tile_X0Y9_W_IO/W6END[4]
+ Tile_X0Y9_W_IO/W6END[5] Tile_X0Y9_W_IO/W6END[6] Tile_X0Y9_W_IO/W6END[7] Tile_X0Y9_W_IO/W6END[8]
+ Tile_X0Y9_W_IO/W6END[9] Tile_X2Y9_LUT4AB/W6BEG[0] Tile_X2Y9_LUT4AB/W6BEG[10] Tile_X2Y9_LUT4AB/W6BEG[11]
+ Tile_X2Y9_LUT4AB/W6BEG[1] Tile_X2Y9_LUT4AB/W6BEG[2] Tile_X2Y9_LUT4AB/W6BEG[3] Tile_X2Y9_LUT4AB/W6BEG[4]
+ Tile_X2Y9_LUT4AB/W6BEG[5] Tile_X2Y9_LUT4AB/W6BEG[6] Tile_X2Y9_LUT4AB/W6BEG[7] Tile_X2Y9_LUT4AB/W6BEG[8]
+ Tile_X2Y9_LUT4AB/W6BEG[9] Tile_X0Y9_W_IO/WW4END[0] Tile_X0Y9_W_IO/WW4END[10] Tile_X0Y9_W_IO/WW4END[11]
+ Tile_X0Y9_W_IO/WW4END[12] Tile_X0Y9_W_IO/WW4END[13] Tile_X0Y9_W_IO/WW4END[14] Tile_X0Y9_W_IO/WW4END[15]
+ Tile_X0Y9_W_IO/WW4END[1] Tile_X0Y9_W_IO/WW4END[2] Tile_X0Y9_W_IO/WW4END[3] Tile_X0Y9_W_IO/WW4END[4]
+ Tile_X0Y9_W_IO/WW4END[5] Tile_X0Y9_W_IO/WW4END[6] Tile_X0Y9_W_IO/WW4END[7] Tile_X0Y9_W_IO/WW4END[8]
+ Tile_X0Y9_W_IO/WW4END[9] Tile_X2Y9_LUT4AB/WW4BEG[0] Tile_X2Y9_LUT4AB/WW4BEG[10]
+ Tile_X2Y9_LUT4AB/WW4BEG[11] Tile_X2Y9_LUT4AB/WW4BEG[12] Tile_X2Y9_LUT4AB/WW4BEG[13]
+ Tile_X2Y9_LUT4AB/WW4BEG[14] Tile_X2Y9_LUT4AB/WW4BEG[15] Tile_X2Y9_LUT4AB/WW4BEG[1]
+ Tile_X2Y9_LUT4AB/WW4BEG[2] Tile_X2Y9_LUT4AB/WW4BEG[3] Tile_X2Y9_LUT4AB/WW4BEG[4]
+ Tile_X2Y9_LUT4AB/WW4BEG[5] Tile_X2Y9_LUT4AB/WW4BEG[6] Tile_X2Y9_LUT4AB/WW4BEG[7]
+ Tile_X2Y9_LUT4AB/WW4BEG[8] Tile_X2Y9_LUT4AB/WW4BEG[9] LUT4AB
XTile_X8Y4_LUT4AB Tile_X8Y5_LUT4AB/Co Tile_X8Y4_LUT4AB/Co Tile_X9Y4_LUT4AB/E1END[0]
+ Tile_X9Y4_LUT4AB/E1END[1] Tile_X9Y4_LUT4AB/E1END[2] Tile_X9Y4_LUT4AB/E1END[3] Tile_X8Y4_LUT4AB/E1END[0]
+ Tile_X8Y4_LUT4AB/E1END[1] Tile_X8Y4_LUT4AB/E1END[2] Tile_X8Y4_LUT4AB/E1END[3] Tile_X9Y4_LUT4AB/E2MID[0]
+ Tile_X9Y4_LUT4AB/E2MID[1] Tile_X9Y4_LUT4AB/E2MID[2] Tile_X9Y4_LUT4AB/E2MID[3] Tile_X9Y4_LUT4AB/E2MID[4]
+ Tile_X9Y4_LUT4AB/E2MID[5] Tile_X9Y4_LUT4AB/E2MID[6] Tile_X9Y4_LUT4AB/E2MID[7] Tile_X9Y4_LUT4AB/E2END[0]
+ Tile_X9Y4_LUT4AB/E2END[1] Tile_X9Y4_LUT4AB/E2END[2] Tile_X9Y4_LUT4AB/E2END[3] Tile_X9Y4_LUT4AB/E2END[4]
+ Tile_X9Y4_LUT4AB/E2END[5] Tile_X9Y4_LUT4AB/E2END[6] Tile_X9Y4_LUT4AB/E2END[7] Tile_X8Y4_LUT4AB/E2END[0]
+ Tile_X8Y4_LUT4AB/E2END[1] Tile_X8Y4_LUT4AB/E2END[2] Tile_X8Y4_LUT4AB/E2END[3] Tile_X8Y4_LUT4AB/E2END[4]
+ Tile_X8Y4_LUT4AB/E2END[5] Tile_X8Y4_LUT4AB/E2END[6] Tile_X8Y4_LUT4AB/E2END[7] Tile_X8Y4_LUT4AB/E2MID[0]
+ Tile_X8Y4_LUT4AB/E2MID[1] Tile_X8Y4_LUT4AB/E2MID[2] Tile_X8Y4_LUT4AB/E2MID[3] Tile_X8Y4_LUT4AB/E2MID[4]
+ Tile_X8Y4_LUT4AB/E2MID[5] Tile_X8Y4_LUT4AB/E2MID[6] Tile_X8Y4_LUT4AB/E2MID[7] Tile_X9Y4_LUT4AB/E6END[0]
+ Tile_X9Y4_LUT4AB/E6END[10] Tile_X9Y4_LUT4AB/E6END[11] Tile_X9Y4_LUT4AB/E6END[1]
+ Tile_X9Y4_LUT4AB/E6END[2] Tile_X9Y4_LUT4AB/E6END[3] Tile_X9Y4_LUT4AB/E6END[4] Tile_X9Y4_LUT4AB/E6END[5]
+ Tile_X9Y4_LUT4AB/E6END[6] Tile_X9Y4_LUT4AB/E6END[7] Tile_X9Y4_LUT4AB/E6END[8] Tile_X9Y4_LUT4AB/E6END[9]
+ Tile_X8Y4_LUT4AB/E6END[0] Tile_X8Y4_LUT4AB/E6END[10] Tile_X8Y4_LUT4AB/E6END[11]
+ Tile_X8Y4_LUT4AB/E6END[1] Tile_X8Y4_LUT4AB/E6END[2] Tile_X8Y4_LUT4AB/E6END[3] Tile_X8Y4_LUT4AB/E6END[4]
+ Tile_X8Y4_LUT4AB/E6END[5] Tile_X8Y4_LUT4AB/E6END[6] Tile_X8Y4_LUT4AB/E6END[7] Tile_X8Y4_LUT4AB/E6END[8]
+ Tile_X8Y4_LUT4AB/E6END[9] Tile_X9Y4_LUT4AB/EE4END[0] Tile_X9Y4_LUT4AB/EE4END[10]
+ Tile_X9Y4_LUT4AB/EE4END[11] Tile_X9Y4_LUT4AB/EE4END[12] Tile_X9Y4_LUT4AB/EE4END[13]
+ Tile_X9Y4_LUT4AB/EE4END[14] Tile_X9Y4_LUT4AB/EE4END[15] Tile_X9Y4_LUT4AB/EE4END[1]
+ Tile_X9Y4_LUT4AB/EE4END[2] Tile_X9Y4_LUT4AB/EE4END[3] Tile_X9Y4_LUT4AB/EE4END[4]
+ Tile_X9Y4_LUT4AB/EE4END[5] Tile_X9Y4_LUT4AB/EE4END[6] Tile_X9Y4_LUT4AB/EE4END[7]
+ Tile_X9Y4_LUT4AB/EE4END[8] Tile_X9Y4_LUT4AB/EE4END[9] Tile_X8Y4_LUT4AB/EE4END[0]
+ Tile_X8Y4_LUT4AB/EE4END[10] Tile_X8Y4_LUT4AB/EE4END[11] Tile_X8Y4_LUT4AB/EE4END[12]
+ Tile_X8Y4_LUT4AB/EE4END[13] Tile_X8Y4_LUT4AB/EE4END[14] Tile_X8Y4_LUT4AB/EE4END[15]
+ Tile_X8Y4_LUT4AB/EE4END[1] Tile_X8Y4_LUT4AB/EE4END[2] Tile_X8Y4_LUT4AB/EE4END[3]
+ Tile_X8Y4_LUT4AB/EE4END[4] Tile_X8Y4_LUT4AB/EE4END[5] Tile_X8Y4_LUT4AB/EE4END[6]
+ Tile_X8Y4_LUT4AB/EE4END[7] Tile_X8Y4_LUT4AB/EE4END[8] Tile_X8Y4_LUT4AB/EE4END[9]
+ Tile_X8Y4_LUT4AB/FrameData[0] Tile_X8Y4_LUT4AB/FrameData[10] Tile_X8Y4_LUT4AB/FrameData[11]
+ Tile_X8Y4_LUT4AB/FrameData[12] Tile_X8Y4_LUT4AB/FrameData[13] Tile_X8Y4_LUT4AB/FrameData[14]
+ Tile_X8Y4_LUT4AB/FrameData[15] Tile_X8Y4_LUT4AB/FrameData[16] Tile_X8Y4_LUT4AB/FrameData[17]
+ Tile_X8Y4_LUT4AB/FrameData[18] Tile_X8Y4_LUT4AB/FrameData[19] Tile_X8Y4_LUT4AB/FrameData[1]
+ Tile_X8Y4_LUT4AB/FrameData[20] Tile_X8Y4_LUT4AB/FrameData[21] Tile_X8Y4_LUT4AB/FrameData[22]
+ Tile_X8Y4_LUT4AB/FrameData[23] Tile_X8Y4_LUT4AB/FrameData[24] Tile_X8Y4_LUT4AB/FrameData[25]
+ Tile_X8Y4_LUT4AB/FrameData[26] Tile_X8Y4_LUT4AB/FrameData[27] Tile_X8Y4_LUT4AB/FrameData[28]
+ Tile_X8Y4_LUT4AB/FrameData[29] Tile_X8Y4_LUT4AB/FrameData[2] Tile_X8Y4_LUT4AB/FrameData[30]
+ Tile_X8Y4_LUT4AB/FrameData[31] Tile_X8Y4_LUT4AB/FrameData[3] Tile_X8Y4_LUT4AB/FrameData[4]
+ Tile_X8Y4_LUT4AB/FrameData[5] Tile_X8Y4_LUT4AB/FrameData[6] Tile_X8Y4_LUT4AB/FrameData[7]
+ Tile_X8Y4_LUT4AB/FrameData[8] Tile_X8Y4_LUT4AB/FrameData[9] Tile_X9Y4_LUT4AB/FrameData[0]
+ Tile_X9Y4_LUT4AB/FrameData[10] Tile_X9Y4_LUT4AB/FrameData[11] Tile_X9Y4_LUT4AB/FrameData[12]
+ Tile_X9Y4_LUT4AB/FrameData[13] Tile_X9Y4_LUT4AB/FrameData[14] Tile_X9Y4_LUT4AB/FrameData[15]
+ Tile_X9Y4_LUT4AB/FrameData[16] Tile_X9Y4_LUT4AB/FrameData[17] Tile_X9Y4_LUT4AB/FrameData[18]
+ Tile_X9Y4_LUT4AB/FrameData[19] Tile_X9Y4_LUT4AB/FrameData[1] Tile_X9Y4_LUT4AB/FrameData[20]
+ Tile_X9Y4_LUT4AB/FrameData[21] Tile_X9Y4_LUT4AB/FrameData[22] Tile_X9Y4_LUT4AB/FrameData[23]
+ Tile_X9Y4_LUT4AB/FrameData[24] Tile_X9Y4_LUT4AB/FrameData[25] Tile_X9Y4_LUT4AB/FrameData[26]
+ Tile_X9Y4_LUT4AB/FrameData[27] Tile_X9Y4_LUT4AB/FrameData[28] Tile_X9Y4_LUT4AB/FrameData[29]
+ Tile_X9Y4_LUT4AB/FrameData[2] Tile_X9Y4_LUT4AB/FrameData[30] Tile_X9Y4_LUT4AB/FrameData[31]
+ Tile_X9Y4_LUT4AB/FrameData[3] Tile_X9Y4_LUT4AB/FrameData[4] Tile_X9Y4_LUT4AB/FrameData[5]
+ Tile_X9Y4_LUT4AB/FrameData[6] Tile_X9Y4_LUT4AB/FrameData[7] Tile_X9Y4_LUT4AB/FrameData[8]
+ Tile_X9Y4_LUT4AB/FrameData[9] Tile_X8Y4_LUT4AB/FrameStrobe[0] Tile_X8Y4_LUT4AB/FrameStrobe[10]
+ Tile_X8Y4_LUT4AB/FrameStrobe[11] Tile_X8Y4_LUT4AB/FrameStrobe[12] Tile_X8Y4_LUT4AB/FrameStrobe[13]
+ Tile_X8Y4_LUT4AB/FrameStrobe[14] Tile_X8Y4_LUT4AB/FrameStrobe[15] Tile_X8Y4_LUT4AB/FrameStrobe[16]
+ Tile_X8Y4_LUT4AB/FrameStrobe[17] Tile_X8Y4_LUT4AB/FrameStrobe[18] Tile_X8Y4_LUT4AB/FrameStrobe[19]
+ Tile_X8Y4_LUT4AB/FrameStrobe[1] Tile_X8Y4_LUT4AB/FrameStrobe[2] Tile_X8Y4_LUT4AB/FrameStrobe[3]
+ Tile_X8Y4_LUT4AB/FrameStrobe[4] Tile_X8Y4_LUT4AB/FrameStrobe[5] Tile_X8Y4_LUT4AB/FrameStrobe[6]
+ Tile_X8Y4_LUT4AB/FrameStrobe[7] Tile_X8Y4_LUT4AB/FrameStrobe[8] Tile_X8Y4_LUT4AB/FrameStrobe[9]
+ Tile_X8Y3_LUT4AB/FrameStrobe[0] Tile_X8Y3_LUT4AB/FrameStrobe[10] Tile_X8Y3_LUT4AB/FrameStrobe[11]
+ Tile_X8Y3_LUT4AB/FrameStrobe[12] Tile_X8Y3_LUT4AB/FrameStrobe[13] Tile_X8Y3_LUT4AB/FrameStrobe[14]
+ Tile_X8Y3_LUT4AB/FrameStrobe[15] Tile_X8Y3_LUT4AB/FrameStrobe[16] Tile_X8Y3_LUT4AB/FrameStrobe[17]
+ Tile_X8Y3_LUT4AB/FrameStrobe[18] Tile_X8Y3_LUT4AB/FrameStrobe[19] Tile_X8Y3_LUT4AB/FrameStrobe[1]
+ Tile_X8Y3_LUT4AB/FrameStrobe[2] Tile_X8Y3_LUT4AB/FrameStrobe[3] Tile_X8Y3_LUT4AB/FrameStrobe[4]
+ Tile_X8Y3_LUT4AB/FrameStrobe[5] Tile_X8Y3_LUT4AB/FrameStrobe[6] Tile_X8Y3_LUT4AB/FrameStrobe[7]
+ Tile_X8Y3_LUT4AB/FrameStrobe[8] Tile_X8Y3_LUT4AB/FrameStrobe[9] Tile_X8Y4_LUT4AB/N1BEG[0]
+ Tile_X8Y4_LUT4AB/N1BEG[1] Tile_X8Y4_LUT4AB/N1BEG[2] Tile_X8Y4_LUT4AB/N1BEG[3] Tile_X8Y5_LUT4AB/N1BEG[0]
+ Tile_X8Y5_LUT4AB/N1BEG[1] Tile_X8Y5_LUT4AB/N1BEG[2] Tile_X8Y5_LUT4AB/N1BEG[3] Tile_X8Y4_LUT4AB/N2BEG[0]
+ Tile_X8Y4_LUT4AB/N2BEG[1] Tile_X8Y4_LUT4AB/N2BEG[2] Tile_X8Y4_LUT4AB/N2BEG[3] Tile_X8Y4_LUT4AB/N2BEG[4]
+ Tile_X8Y4_LUT4AB/N2BEG[5] Tile_X8Y4_LUT4AB/N2BEG[6] Tile_X8Y4_LUT4AB/N2BEG[7] Tile_X8Y3_LUT4AB/N2END[0]
+ Tile_X8Y3_LUT4AB/N2END[1] Tile_X8Y3_LUT4AB/N2END[2] Tile_X8Y3_LUT4AB/N2END[3] Tile_X8Y3_LUT4AB/N2END[4]
+ Tile_X8Y3_LUT4AB/N2END[5] Tile_X8Y3_LUT4AB/N2END[6] Tile_X8Y3_LUT4AB/N2END[7] Tile_X8Y4_LUT4AB/N2END[0]
+ Tile_X8Y4_LUT4AB/N2END[1] Tile_X8Y4_LUT4AB/N2END[2] Tile_X8Y4_LUT4AB/N2END[3] Tile_X8Y4_LUT4AB/N2END[4]
+ Tile_X8Y4_LUT4AB/N2END[5] Tile_X8Y4_LUT4AB/N2END[6] Tile_X8Y4_LUT4AB/N2END[7] Tile_X8Y5_LUT4AB/N2BEG[0]
+ Tile_X8Y5_LUT4AB/N2BEG[1] Tile_X8Y5_LUT4AB/N2BEG[2] Tile_X8Y5_LUT4AB/N2BEG[3] Tile_X8Y5_LUT4AB/N2BEG[4]
+ Tile_X8Y5_LUT4AB/N2BEG[5] Tile_X8Y5_LUT4AB/N2BEG[6] Tile_X8Y5_LUT4AB/N2BEG[7] Tile_X8Y4_LUT4AB/N4BEG[0]
+ Tile_X8Y4_LUT4AB/N4BEG[10] Tile_X8Y4_LUT4AB/N4BEG[11] Tile_X8Y4_LUT4AB/N4BEG[12]
+ Tile_X8Y4_LUT4AB/N4BEG[13] Tile_X8Y4_LUT4AB/N4BEG[14] Tile_X8Y4_LUT4AB/N4BEG[15]
+ Tile_X8Y4_LUT4AB/N4BEG[1] Tile_X8Y4_LUT4AB/N4BEG[2] Tile_X8Y4_LUT4AB/N4BEG[3] Tile_X8Y4_LUT4AB/N4BEG[4]
+ Tile_X8Y4_LUT4AB/N4BEG[5] Tile_X8Y4_LUT4AB/N4BEG[6] Tile_X8Y4_LUT4AB/N4BEG[7] Tile_X8Y4_LUT4AB/N4BEG[8]
+ Tile_X8Y4_LUT4AB/N4BEG[9] Tile_X8Y5_LUT4AB/N4BEG[0] Tile_X8Y5_LUT4AB/N4BEG[10] Tile_X8Y5_LUT4AB/N4BEG[11]
+ Tile_X8Y5_LUT4AB/N4BEG[12] Tile_X8Y5_LUT4AB/N4BEG[13] Tile_X8Y5_LUT4AB/N4BEG[14]
+ Tile_X8Y5_LUT4AB/N4BEG[15] Tile_X8Y5_LUT4AB/N4BEG[1] Tile_X8Y5_LUT4AB/N4BEG[2] Tile_X8Y5_LUT4AB/N4BEG[3]
+ Tile_X8Y5_LUT4AB/N4BEG[4] Tile_X8Y5_LUT4AB/N4BEG[5] Tile_X8Y5_LUT4AB/N4BEG[6] Tile_X8Y5_LUT4AB/N4BEG[7]
+ Tile_X8Y5_LUT4AB/N4BEG[8] Tile_X8Y5_LUT4AB/N4BEG[9] Tile_X8Y4_LUT4AB/NN4BEG[0] Tile_X8Y4_LUT4AB/NN4BEG[10]
+ Tile_X8Y4_LUT4AB/NN4BEG[11] Tile_X8Y4_LUT4AB/NN4BEG[12] Tile_X8Y4_LUT4AB/NN4BEG[13]
+ Tile_X8Y4_LUT4AB/NN4BEG[14] Tile_X8Y4_LUT4AB/NN4BEG[15] Tile_X8Y4_LUT4AB/NN4BEG[1]
+ Tile_X8Y4_LUT4AB/NN4BEG[2] Tile_X8Y4_LUT4AB/NN4BEG[3] Tile_X8Y4_LUT4AB/NN4BEG[4]
+ Tile_X8Y4_LUT4AB/NN4BEG[5] Tile_X8Y4_LUT4AB/NN4BEG[6] Tile_X8Y4_LUT4AB/NN4BEG[7]
+ Tile_X8Y4_LUT4AB/NN4BEG[8] Tile_X8Y4_LUT4AB/NN4BEG[9] Tile_X8Y5_LUT4AB/NN4BEG[0]
+ Tile_X8Y5_LUT4AB/NN4BEG[10] Tile_X8Y5_LUT4AB/NN4BEG[11] Tile_X8Y5_LUT4AB/NN4BEG[12]
+ Tile_X8Y5_LUT4AB/NN4BEG[13] Tile_X8Y5_LUT4AB/NN4BEG[14] Tile_X8Y5_LUT4AB/NN4BEG[15]
+ Tile_X8Y5_LUT4AB/NN4BEG[1] Tile_X8Y5_LUT4AB/NN4BEG[2] Tile_X8Y5_LUT4AB/NN4BEG[3]
+ Tile_X8Y5_LUT4AB/NN4BEG[4] Tile_X8Y5_LUT4AB/NN4BEG[5] Tile_X8Y5_LUT4AB/NN4BEG[6]
+ Tile_X8Y5_LUT4AB/NN4BEG[7] Tile_X8Y5_LUT4AB/NN4BEG[8] Tile_X8Y5_LUT4AB/NN4BEG[9]
+ Tile_X8Y5_LUT4AB/S1END[0] Tile_X8Y5_LUT4AB/S1END[1] Tile_X8Y5_LUT4AB/S1END[2] Tile_X8Y5_LUT4AB/S1END[3]
+ Tile_X8Y4_LUT4AB/S1END[0] Tile_X8Y4_LUT4AB/S1END[1] Tile_X8Y4_LUT4AB/S1END[2] Tile_X8Y4_LUT4AB/S1END[3]
+ Tile_X8Y5_LUT4AB/S2MID[0] Tile_X8Y5_LUT4AB/S2MID[1] Tile_X8Y5_LUT4AB/S2MID[2] Tile_X8Y5_LUT4AB/S2MID[3]
+ Tile_X8Y5_LUT4AB/S2MID[4] Tile_X8Y5_LUT4AB/S2MID[5] Tile_X8Y5_LUT4AB/S2MID[6] Tile_X8Y5_LUT4AB/S2MID[7]
+ Tile_X8Y5_LUT4AB/S2END[0] Tile_X8Y5_LUT4AB/S2END[1] Tile_X8Y5_LUT4AB/S2END[2] Tile_X8Y5_LUT4AB/S2END[3]
+ Tile_X8Y5_LUT4AB/S2END[4] Tile_X8Y5_LUT4AB/S2END[5] Tile_X8Y5_LUT4AB/S2END[6] Tile_X8Y5_LUT4AB/S2END[7]
+ Tile_X8Y4_LUT4AB/S2END[0] Tile_X8Y4_LUT4AB/S2END[1] Tile_X8Y4_LUT4AB/S2END[2] Tile_X8Y4_LUT4AB/S2END[3]
+ Tile_X8Y4_LUT4AB/S2END[4] Tile_X8Y4_LUT4AB/S2END[5] Tile_X8Y4_LUT4AB/S2END[6] Tile_X8Y4_LUT4AB/S2END[7]
+ Tile_X8Y4_LUT4AB/S2MID[0] Tile_X8Y4_LUT4AB/S2MID[1] Tile_X8Y4_LUT4AB/S2MID[2] Tile_X8Y4_LUT4AB/S2MID[3]
+ Tile_X8Y4_LUT4AB/S2MID[4] Tile_X8Y4_LUT4AB/S2MID[5] Tile_X8Y4_LUT4AB/S2MID[6] Tile_X8Y4_LUT4AB/S2MID[7]
+ Tile_X8Y5_LUT4AB/S4END[0] Tile_X8Y5_LUT4AB/S4END[10] Tile_X8Y5_LUT4AB/S4END[11]
+ Tile_X8Y5_LUT4AB/S4END[12] Tile_X8Y5_LUT4AB/S4END[13] Tile_X8Y5_LUT4AB/S4END[14]
+ Tile_X8Y5_LUT4AB/S4END[15] Tile_X8Y5_LUT4AB/S4END[1] Tile_X8Y5_LUT4AB/S4END[2] Tile_X8Y5_LUT4AB/S4END[3]
+ Tile_X8Y5_LUT4AB/S4END[4] Tile_X8Y5_LUT4AB/S4END[5] Tile_X8Y5_LUT4AB/S4END[6] Tile_X8Y5_LUT4AB/S4END[7]
+ Tile_X8Y5_LUT4AB/S4END[8] Tile_X8Y5_LUT4AB/S4END[9] Tile_X8Y4_LUT4AB/S4END[0] Tile_X8Y4_LUT4AB/S4END[10]
+ Tile_X8Y4_LUT4AB/S4END[11] Tile_X8Y4_LUT4AB/S4END[12] Tile_X8Y4_LUT4AB/S4END[13]
+ Tile_X8Y4_LUT4AB/S4END[14] Tile_X8Y4_LUT4AB/S4END[15] Tile_X8Y4_LUT4AB/S4END[1]
+ Tile_X8Y4_LUT4AB/S4END[2] Tile_X8Y4_LUT4AB/S4END[3] Tile_X8Y4_LUT4AB/S4END[4] Tile_X8Y4_LUT4AB/S4END[5]
+ Tile_X8Y4_LUT4AB/S4END[6] Tile_X8Y4_LUT4AB/S4END[7] Tile_X8Y4_LUT4AB/S4END[8] Tile_X8Y4_LUT4AB/S4END[9]
+ Tile_X8Y5_LUT4AB/SS4END[0] Tile_X8Y5_LUT4AB/SS4END[10] Tile_X8Y5_LUT4AB/SS4END[11]
+ Tile_X8Y5_LUT4AB/SS4END[12] Tile_X8Y5_LUT4AB/SS4END[13] Tile_X8Y5_LUT4AB/SS4END[14]
+ Tile_X8Y5_LUT4AB/SS4END[15] Tile_X8Y5_LUT4AB/SS4END[1] Tile_X8Y5_LUT4AB/SS4END[2]
+ Tile_X8Y5_LUT4AB/SS4END[3] Tile_X8Y5_LUT4AB/SS4END[4] Tile_X8Y5_LUT4AB/SS4END[5]
+ Tile_X8Y5_LUT4AB/SS4END[6] Tile_X8Y5_LUT4AB/SS4END[7] Tile_X8Y5_LUT4AB/SS4END[8]
+ Tile_X8Y5_LUT4AB/SS4END[9] Tile_X8Y4_LUT4AB/SS4END[0] Tile_X8Y4_LUT4AB/SS4END[10]
+ Tile_X8Y4_LUT4AB/SS4END[11] Tile_X8Y4_LUT4AB/SS4END[12] Tile_X8Y4_LUT4AB/SS4END[13]
+ Tile_X8Y4_LUT4AB/SS4END[14] Tile_X8Y4_LUT4AB/SS4END[15] Tile_X8Y4_LUT4AB/SS4END[1]
+ Tile_X8Y4_LUT4AB/SS4END[2] Tile_X8Y4_LUT4AB/SS4END[3] Tile_X8Y4_LUT4AB/SS4END[4]
+ Tile_X8Y4_LUT4AB/SS4END[5] Tile_X8Y4_LUT4AB/SS4END[6] Tile_X8Y4_LUT4AB/SS4END[7]
+ Tile_X8Y4_LUT4AB/SS4END[8] Tile_X8Y4_LUT4AB/SS4END[9] Tile_X8Y4_LUT4AB/UserCLK Tile_X8Y3_LUT4AB/UserCLK
+ VGND VPWR Tile_X8Y4_LUT4AB/W1BEG[0] Tile_X8Y4_LUT4AB/W1BEG[1] Tile_X8Y4_LUT4AB/W1BEG[2]
+ Tile_X8Y4_LUT4AB/W1BEG[3] Tile_X9Y4_LUT4AB/W1BEG[0] Tile_X9Y4_LUT4AB/W1BEG[1] Tile_X9Y4_LUT4AB/W1BEG[2]
+ Tile_X9Y4_LUT4AB/W1BEG[3] Tile_X8Y4_LUT4AB/W2BEG[0] Tile_X8Y4_LUT4AB/W2BEG[1] Tile_X8Y4_LUT4AB/W2BEG[2]
+ Tile_X8Y4_LUT4AB/W2BEG[3] Tile_X8Y4_LUT4AB/W2BEG[4] Tile_X8Y4_LUT4AB/W2BEG[5] Tile_X8Y4_LUT4AB/W2BEG[6]
+ Tile_X8Y4_LUT4AB/W2BEG[7] Tile_X8Y4_LUT4AB/W2BEGb[0] Tile_X8Y4_LUT4AB/W2BEGb[1]
+ Tile_X8Y4_LUT4AB/W2BEGb[2] Tile_X8Y4_LUT4AB/W2BEGb[3] Tile_X8Y4_LUT4AB/W2BEGb[4]
+ Tile_X8Y4_LUT4AB/W2BEGb[5] Tile_X8Y4_LUT4AB/W2BEGb[6] Tile_X8Y4_LUT4AB/W2BEGb[7]
+ Tile_X8Y4_LUT4AB/W2END[0] Tile_X8Y4_LUT4AB/W2END[1] Tile_X8Y4_LUT4AB/W2END[2] Tile_X8Y4_LUT4AB/W2END[3]
+ Tile_X8Y4_LUT4AB/W2END[4] Tile_X8Y4_LUT4AB/W2END[5] Tile_X8Y4_LUT4AB/W2END[6] Tile_X8Y4_LUT4AB/W2END[7]
+ Tile_X9Y4_LUT4AB/W2BEG[0] Tile_X9Y4_LUT4AB/W2BEG[1] Tile_X9Y4_LUT4AB/W2BEG[2] Tile_X9Y4_LUT4AB/W2BEG[3]
+ Tile_X9Y4_LUT4AB/W2BEG[4] Tile_X9Y4_LUT4AB/W2BEG[5] Tile_X9Y4_LUT4AB/W2BEG[6] Tile_X9Y4_LUT4AB/W2BEG[7]
+ Tile_X8Y4_LUT4AB/W6BEG[0] Tile_X8Y4_LUT4AB/W6BEG[10] Tile_X8Y4_LUT4AB/W6BEG[11]
+ Tile_X8Y4_LUT4AB/W6BEG[1] Tile_X8Y4_LUT4AB/W6BEG[2] Tile_X8Y4_LUT4AB/W6BEG[3] Tile_X8Y4_LUT4AB/W6BEG[4]
+ Tile_X8Y4_LUT4AB/W6BEG[5] Tile_X8Y4_LUT4AB/W6BEG[6] Tile_X8Y4_LUT4AB/W6BEG[7] Tile_X8Y4_LUT4AB/W6BEG[8]
+ Tile_X8Y4_LUT4AB/W6BEG[9] Tile_X9Y4_LUT4AB/W6BEG[0] Tile_X9Y4_LUT4AB/W6BEG[10] Tile_X9Y4_LUT4AB/W6BEG[11]
+ Tile_X9Y4_LUT4AB/W6BEG[1] Tile_X9Y4_LUT4AB/W6BEG[2] Tile_X9Y4_LUT4AB/W6BEG[3] Tile_X9Y4_LUT4AB/W6BEG[4]
+ Tile_X9Y4_LUT4AB/W6BEG[5] Tile_X9Y4_LUT4AB/W6BEG[6] Tile_X9Y4_LUT4AB/W6BEG[7] Tile_X9Y4_LUT4AB/W6BEG[8]
+ Tile_X9Y4_LUT4AB/W6BEG[9] Tile_X8Y4_LUT4AB/WW4BEG[0] Tile_X8Y4_LUT4AB/WW4BEG[10]
+ Tile_X8Y4_LUT4AB/WW4BEG[11] Tile_X8Y4_LUT4AB/WW4BEG[12] Tile_X8Y4_LUT4AB/WW4BEG[13]
+ Tile_X8Y4_LUT4AB/WW4BEG[14] Tile_X8Y4_LUT4AB/WW4BEG[15] Tile_X8Y4_LUT4AB/WW4BEG[1]
+ Tile_X8Y4_LUT4AB/WW4BEG[2] Tile_X8Y4_LUT4AB/WW4BEG[3] Tile_X8Y4_LUT4AB/WW4BEG[4]
+ Tile_X8Y4_LUT4AB/WW4BEG[5] Tile_X8Y4_LUT4AB/WW4BEG[6] Tile_X8Y4_LUT4AB/WW4BEG[7]
+ Tile_X8Y4_LUT4AB/WW4BEG[8] Tile_X8Y4_LUT4AB/WW4BEG[9] Tile_X9Y4_LUT4AB/WW4BEG[0]
+ Tile_X9Y4_LUT4AB/WW4BEG[10] Tile_X9Y4_LUT4AB/WW4BEG[11] Tile_X9Y4_LUT4AB/WW4BEG[12]
+ Tile_X9Y4_LUT4AB/WW4BEG[13] Tile_X9Y4_LUT4AB/WW4BEG[14] Tile_X9Y4_LUT4AB/WW4BEG[15]
+ Tile_X9Y4_LUT4AB/WW4BEG[1] Tile_X9Y4_LUT4AB/WW4BEG[2] Tile_X9Y4_LUT4AB/WW4BEG[3]
+ Tile_X9Y4_LUT4AB/WW4BEG[4] Tile_X9Y4_LUT4AB/WW4BEG[5] Tile_X9Y4_LUT4AB/WW4BEG[6]
+ Tile_X9Y4_LUT4AB/WW4BEG[7] Tile_X9Y4_LUT4AB/WW4BEG[8] Tile_X9Y4_LUT4AB/WW4BEG[9]
+ LUT4AB
XTile_X3Y14_LUT4AB Tile_X3Y14_LUT4AB/Ci Tile_X3Y14_LUT4AB/Co Tile_X3Y14_LUT4AB/E1BEG[0]
+ Tile_X3Y14_LUT4AB/E1BEG[1] Tile_X3Y14_LUT4AB/E1BEG[2] Tile_X3Y14_LUT4AB/E1BEG[3]
+ Tile_X3Y14_LUT4AB/E1END[0] Tile_X3Y14_LUT4AB/E1END[1] Tile_X3Y14_LUT4AB/E1END[2]
+ Tile_X3Y14_LUT4AB/E1END[3] Tile_X3Y14_LUT4AB/E2BEG[0] Tile_X3Y14_LUT4AB/E2BEG[1]
+ Tile_X3Y14_LUT4AB/E2BEG[2] Tile_X3Y14_LUT4AB/E2BEG[3] Tile_X3Y14_LUT4AB/E2BEG[4]
+ Tile_X3Y14_LUT4AB/E2BEG[5] Tile_X3Y14_LUT4AB/E2BEG[6] Tile_X3Y14_LUT4AB/E2BEG[7]
+ Tile_X4Y14_RegFile/E2END[0] Tile_X4Y14_RegFile/E2END[1] Tile_X4Y14_RegFile/E2END[2]
+ Tile_X4Y14_RegFile/E2END[3] Tile_X4Y14_RegFile/E2END[4] Tile_X4Y14_RegFile/E2END[5]
+ Tile_X4Y14_RegFile/E2END[6] Tile_X4Y14_RegFile/E2END[7] Tile_X3Y14_LUT4AB/E2END[0]
+ Tile_X3Y14_LUT4AB/E2END[1] Tile_X3Y14_LUT4AB/E2END[2] Tile_X3Y14_LUT4AB/E2END[3]
+ Tile_X3Y14_LUT4AB/E2END[4] Tile_X3Y14_LUT4AB/E2END[5] Tile_X3Y14_LUT4AB/E2END[6]
+ Tile_X3Y14_LUT4AB/E2END[7] Tile_X3Y14_LUT4AB/E2MID[0] Tile_X3Y14_LUT4AB/E2MID[1]
+ Tile_X3Y14_LUT4AB/E2MID[2] Tile_X3Y14_LUT4AB/E2MID[3] Tile_X3Y14_LUT4AB/E2MID[4]
+ Tile_X3Y14_LUT4AB/E2MID[5] Tile_X3Y14_LUT4AB/E2MID[6] Tile_X3Y14_LUT4AB/E2MID[7]
+ Tile_X3Y14_LUT4AB/E6BEG[0] Tile_X3Y14_LUT4AB/E6BEG[10] Tile_X3Y14_LUT4AB/E6BEG[11]
+ Tile_X3Y14_LUT4AB/E6BEG[1] Tile_X3Y14_LUT4AB/E6BEG[2] Tile_X3Y14_LUT4AB/E6BEG[3]
+ Tile_X3Y14_LUT4AB/E6BEG[4] Tile_X3Y14_LUT4AB/E6BEG[5] Tile_X3Y14_LUT4AB/E6BEG[6]
+ Tile_X3Y14_LUT4AB/E6BEG[7] Tile_X3Y14_LUT4AB/E6BEG[8] Tile_X3Y14_LUT4AB/E6BEG[9]
+ Tile_X3Y14_LUT4AB/E6END[0] Tile_X3Y14_LUT4AB/E6END[10] Tile_X3Y14_LUT4AB/E6END[11]
+ Tile_X3Y14_LUT4AB/E6END[1] Tile_X3Y14_LUT4AB/E6END[2] Tile_X3Y14_LUT4AB/E6END[3]
+ Tile_X3Y14_LUT4AB/E6END[4] Tile_X3Y14_LUT4AB/E6END[5] Tile_X3Y14_LUT4AB/E6END[6]
+ Tile_X3Y14_LUT4AB/E6END[7] Tile_X3Y14_LUT4AB/E6END[8] Tile_X3Y14_LUT4AB/E6END[9]
+ Tile_X3Y14_LUT4AB/EE4BEG[0] Tile_X3Y14_LUT4AB/EE4BEG[10] Tile_X3Y14_LUT4AB/EE4BEG[11]
+ Tile_X3Y14_LUT4AB/EE4BEG[12] Tile_X3Y14_LUT4AB/EE4BEG[13] Tile_X3Y14_LUT4AB/EE4BEG[14]
+ Tile_X3Y14_LUT4AB/EE4BEG[15] Tile_X3Y14_LUT4AB/EE4BEG[1] Tile_X3Y14_LUT4AB/EE4BEG[2]
+ Tile_X3Y14_LUT4AB/EE4BEG[3] Tile_X3Y14_LUT4AB/EE4BEG[4] Tile_X3Y14_LUT4AB/EE4BEG[5]
+ Tile_X3Y14_LUT4AB/EE4BEG[6] Tile_X3Y14_LUT4AB/EE4BEG[7] Tile_X3Y14_LUT4AB/EE4BEG[8]
+ Tile_X3Y14_LUT4AB/EE4BEG[9] Tile_X3Y14_LUT4AB/EE4END[0] Tile_X3Y14_LUT4AB/EE4END[10]
+ Tile_X3Y14_LUT4AB/EE4END[11] Tile_X3Y14_LUT4AB/EE4END[12] Tile_X3Y14_LUT4AB/EE4END[13]
+ Tile_X3Y14_LUT4AB/EE4END[14] Tile_X3Y14_LUT4AB/EE4END[15] Tile_X3Y14_LUT4AB/EE4END[1]
+ Tile_X3Y14_LUT4AB/EE4END[2] Tile_X3Y14_LUT4AB/EE4END[3] Tile_X3Y14_LUT4AB/EE4END[4]
+ Tile_X3Y14_LUT4AB/EE4END[5] Tile_X3Y14_LUT4AB/EE4END[6] Tile_X3Y14_LUT4AB/EE4END[7]
+ Tile_X3Y14_LUT4AB/EE4END[8] Tile_X3Y14_LUT4AB/EE4END[9] Tile_X3Y14_LUT4AB/FrameData[0]
+ Tile_X3Y14_LUT4AB/FrameData[10] Tile_X3Y14_LUT4AB/FrameData[11] Tile_X3Y14_LUT4AB/FrameData[12]
+ Tile_X3Y14_LUT4AB/FrameData[13] Tile_X3Y14_LUT4AB/FrameData[14] Tile_X3Y14_LUT4AB/FrameData[15]
+ Tile_X3Y14_LUT4AB/FrameData[16] Tile_X3Y14_LUT4AB/FrameData[17] Tile_X3Y14_LUT4AB/FrameData[18]
+ Tile_X3Y14_LUT4AB/FrameData[19] Tile_X3Y14_LUT4AB/FrameData[1] Tile_X3Y14_LUT4AB/FrameData[20]
+ Tile_X3Y14_LUT4AB/FrameData[21] Tile_X3Y14_LUT4AB/FrameData[22] Tile_X3Y14_LUT4AB/FrameData[23]
+ Tile_X3Y14_LUT4AB/FrameData[24] Tile_X3Y14_LUT4AB/FrameData[25] Tile_X3Y14_LUT4AB/FrameData[26]
+ Tile_X3Y14_LUT4AB/FrameData[27] Tile_X3Y14_LUT4AB/FrameData[28] Tile_X3Y14_LUT4AB/FrameData[29]
+ Tile_X3Y14_LUT4AB/FrameData[2] Tile_X3Y14_LUT4AB/FrameData[30] Tile_X3Y14_LUT4AB/FrameData[31]
+ Tile_X3Y14_LUT4AB/FrameData[3] Tile_X3Y14_LUT4AB/FrameData[4] Tile_X3Y14_LUT4AB/FrameData[5]
+ Tile_X3Y14_LUT4AB/FrameData[6] Tile_X3Y14_LUT4AB/FrameData[7] Tile_X3Y14_LUT4AB/FrameData[8]
+ Tile_X3Y14_LUT4AB/FrameData[9] Tile_X4Y14_RegFile/FrameData[0] Tile_X4Y14_RegFile/FrameData[10]
+ Tile_X4Y14_RegFile/FrameData[11] Tile_X4Y14_RegFile/FrameData[12] Tile_X4Y14_RegFile/FrameData[13]
+ Tile_X4Y14_RegFile/FrameData[14] Tile_X4Y14_RegFile/FrameData[15] Tile_X4Y14_RegFile/FrameData[16]
+ Tile_X4Y14_RegFile/FrameData[17] Tile_X4Y14_RegFile/FrameData[18] Tile_X4Y14_RegFile/FrameData[19]
+ Tile_X4Y14_RegFile/FrameData[1] Tile_X4Y14_RegFile/FrameData[20] Tile_X4Y14_RegFile/FrameData[21]
+ Tile_X4Y14_RegFile/FrameData[22] Tile_X4Y14_RegFile/FrameData[23] Tile_X4Y14_RegFile/FrameData[24]
+ Tile_X4Y14_RegFile/FrameData[25] Tile_X4Y14_RegFile/FrameData[26] Tile_X4Y14_RegFile/FrameData[27]
+ Tile_X4Y14_RegFile/FrameData[28] Tile_X4Y14_RegFile/FrameData[29] Tile_X4Y14_RegFile/FrameData[2]
+ Tile_X4Y14_RegFile/FrameData[30] Tile_X4Y14_RegFile/FrameData[31] Tile_X4Y14_RegFile/FrameData[3]
+ Tile_X4Y14_RegFile/FrameData[4] Tile_X4Y14_RegFile/FrameData[5] Tile_X4Y14_RegFile/FrameData[6]
+ Tile_X4Y14_RegFile/FrameData[7] Tile_X4Y14_RegFile/FrameData[8] Tile_X4Y14_RegFile/FrameData[9]
+ Tile_X3Y14_LUT4AB/FrameStrobe[0] Tile_X3Y14_LUT4AB/FrameStrobe[10] Tile_X3Y14_LUT4AB/FrameStrobe[11]
+ Tile_X3Y14_LUT4AB/FrameStrobe[12] Tile_X3Y14_LUT4AB/FrameStrobe[13] Tile_X3Y14_LUT4AB/FrameStrobe[14]
+ Tile_X3Y14_LUT4AB/FrameStrobe[15] Tile_X3Y14_LUT4AB/FrameStrobe[16] Tile_X3Y14_LUT4AB/FrameStrobe[17]
+ Tile_X3Y14_LUT4AB/FrameStrobe[18] Tile_X3Y14_LUT4AB/FrameStrobe[19] Tile_X3Y14_LUT4AB/FrameStrobe[1]
+ Tile_X3Y14_LUT4AB/FrameStrobe[2] Tile_X3Y14_LUT4AB/FrameStrobe[3] Tile_X3Y14_LUT4AB/FrameStrobe[4]
+ Tile_X3Y14_LUT4AB/FrameStrobe[5] Tile_X3Y14_LUT4AB/FrameStrobe[6] Tile_X3Y14_LUT4AB/FrameStrobe[7]
+ Tile_X3Y14_LUT4AB/FrameStrobe[8] Tile_X3Y14_LUT4AB/FrameStrobe[9] Tile_X3Y13_LUT4AB/FrameStrobe[0]
+ Tile_X3Y13_LUT4AB/FrameStrobe[10] Tile_X3Y13_LUT4AB/FrameStrobe[11] Tile_X3Y13_LUT4AB/FrameStrobe[12]
+ Tile_X3Y13_LUT4AB/FrameStrobe[13] Tile_X3Y13_LUT4AB/FrameStrobe[14] Tile_X3Y13_LUT4AB/FrameStrobe[15]
+ Tile_X3Y13_LUT4AB/FrameStrobe[16] Tile_X3Y13_LUT4AB/FrameStrobe[17] Tile_X3Y13_LUT4AB/FrameStrobe[18]
+ Tile_X3Y13_LUT4AB/FrameStrobe[19] Tile_X3Y13_LUT4AB/FrameStrobe[1] Tile_X3Y13_LUT4AB/FrameStrobe[2]
+ Tile_X3Y13_LUT4AB/FrameStrobe[3] Tile_X3Y13_LUT4AB/FrameStrobe[4] Tile_X3Y13_LUT4AB/FrameStrobe[5]
+ Tile_X3Y13_LUT4AB/FrameStrobe[6] Tile_X3Y13_LUT4AB/FrameStrobe[7] Tile_X3Y13_LUT4AB/FrameStrobe[8]
+ Tile_X3Y13_LUT4AB/FrameStrobe[9] Tile_X3Y14_LUT4AB/N1BEG[0] Tile_X3Y14_LUT4AB/N1BEG[1]
+ Tile_X3Y14_LUT4AB/N1BEG[2] Tile_X3Y14_LUT4AB/N1BEG[3] Tile_X3Y14_LUT4AB/N1END[0]
+ Tile_X3Y14_LUT4AB/N1END[1] Tile_X3Y14_LUT4AB/N1END[2] Tile_X3Y14_LUT4AB/N1END[3]
+ Tile_X3Y14_LUT4AB/N2BEG[0] Tile_X3Y14_LUT4AB/N2BEG[1] Tile_X3Y14_LUT4AB/N2BEG[2]
+ Tile_X3Y14_LUT4AB/N2BEG[3] Tile_X3Y14_LUT4AB/N2BEG[4] Tile_X3Y14_LUT4AB/N2BEG[5]
+ Tile_X3Y14_LUT4AB/N2BEG[6] Tile_X3Y14_LUT4AB/N2BEG[7] Tile_X3Y13_LUT4AB/N2END[0]
+ Tile_X3Y13_LUT4AB/N2END[1] Tile_X3Y13_LUT4AB/N2END[2] Tile_X3Y13_LUT4AB/N2END[3]
+ Tile_X3Y13_LUT4AB/N2END[4] Tile_X3Y13_LUT4AB/N2END[5] Tile_X3Y13_LUT4AB/N2END[6]
+ Tile_X3Y13_LUT4AB/N2END[7] Tile_X3Y14_LUT4AB/N2END[0] Tile_X3Y14_LUT4AB/N2END[1]
+ Tile_X3Y14_LUT4AB/N2END[2] Tile_X3Y14_LUT4AB/N2END[3] Tile_X3Y14_LUT4AB/N2END[4]
+ Tile_X3Y14_LUT4AB/N2END[5] Tile_X3Y14_LUT4AB/N2END[6] Tile_X3Y14_LUT4AB/N2END[7]
+ Tile_X3Y14_LUT4AB/N2MID[0] Tile_X3Y14_LUT4AB/N2MID[1] Tile_X3Y14_LUT4AB/N2MID[2]
+ Tile_X3Y14_LUT4AB/N2MID[3] Tile_X3Y14_LUT4AB/N2MID[4] Tile_X3Y14_LUT4AB/N2MID[5]
+ Tile_X3Y14_LUT4AB/N2MID[6] Tile_X3Y14_LUT4AB/N2MID[7] Tile_X3Y14_LUT4AB/N4BEG[0]
+ Tile_X3Y14_LUT4AB/N4BEG[10] Tile_X3Y14_LUT4AB/N4BEG[11] Tile_X3Y14_LUT4AB/N4BEG[12]
+ Tile_X3Y14_LUT4AB/N4BEG[13] Tile_X3Y14_LUT4AB/N4BEG[14] Tile_X3Y14_LUT4AB/N4BEG[15]
+ Tile_X3Y14_LUT4AB/N4BEG[1] Tile_X3Y14_LUT4AB/N4BEG[2] Tile_X3Y14_LUT4AB/N4BEG[3]
+ Tile_X3Y14_LUT4AB/N4BEG[4] Tile_X3Y14_LUT4AB/N4BEG[5] Tile_X3Y14_LUT4AB/N4BEG[6]
+ Tile_X3Y14_LUT4AB/N4BEG[7] Tile_X3Y14_LUT4AB/N4BEG[8] Tile_X3Y14_LUT4AB/N4BEG[9]
+ Tile_X3Y14_LUT4AB/N4END[0] Tile_X3Y14_LUT4AB/N4END[10] Tile_X3Y14_LUT4AB/N4END[11]
+ Tile_X3Y14_LUT4AB/N4END[12] Tile_X3Y14_LUT4AB/N4END[13] Tile_X3Y14_LUT4AB/N4END[14]
+ Tile_X3Y14_LUT4AB/N4END[15] Tile_X3Y14_LUT4AB/N4END[1] Tile_X3Y14_LUT4AB/N4END[2]
+ Tile_X3Y14_LUT4AB/N4END[3] Tile_X3Y14_LUT4AB/N4END[4] Tile_X3Y14_LUT4AB/N4END[5]
+ Tile_X3Y14_LUT4AB/N4END[6] Tile_X3Y14_LUT4AB/N4END[7] Tile_X3Y14_LUT4AB/N4END[8]
+ Tile_X3Y14_LUT4AB/N4END[9] Tile_X3Y14_LUT4AB/NN4BEG[0] Tile_X3Y14_LUT4AB/NN4BEG[10]
+ Tile_X3Y14_LUT4AB/NN4BEG[11] Tile_X3Y14_LUT4AB/NN4BEG[12] Tile_X3Y14_LUT4AB/NN4BEG[13]
+ Tile_X3Y14_LUT4AB/NN4BEG[14] Tile_X3Y14_LUT4AB/NN4BEG[15] Tile_X3Y14_LUT4AB/NN4BEG[1]
+ Tile_X3Y14_LUT4AB/NN4BEG[2] Tile_X3Y14_LUT4AB/NN4BEG[3] Tile_X3Y14_LUT4AB/NN4BEG[4]
+ Tile_X3Y14_LUT4AB/NN4BEG[5] Tile_X3Y14_LUT4AB/NN4BEG[6] Tile_X3Y14_LUT4AB/NN4BEG[7]
+ Tile_X3Y14_LUT4AB/NN4BEG[8] Tile_X3Y14_LUT4AB/NN4BEG[9] Tile_X3Y14_LUT4AB/NN4END[0]
+ Tile_X3Y14_LUT4AB/NN4END[10] Tile_X3Y14_LUT4AB/NN4END[11] Tile_X3Y14_LUT4AB/NN4END[12]
+ Tile_X3Y14_LUT4AB/NN4END[13] Tile_X3Y14_LUT4AB/NN4END[14] Tile_X3Y14_LUT4AB/NN4END[15]
+ Tile_X3Y14_LUT4AB/NN4END[1] Tile_X3Y14_LUT4AB/NN4END[2] Tile_X3Y14_LUT4AB/NN4END[3]
+ Tile_X3Y14_LUT4AB/NN4END[4] Tile_X3Y14_LUT4AB/NN4END[5] Tile_X3Y14_LUT4AB/NN4END[6]
+ Tile_X3Y14_LUT4AB/NN4END[7] Tile_X3Y14_LUT4AB/NN4END[8] Tile_X3Y14_LUT4AB/NN4END[9]
+ Tile_X3Y14_LUT4AB/S1BEG[0] Tile_X3Y14_LUT4AB/S1BEG[1] Tile_X3Y14_LUT4AB/S1BEG[2]
+ Tile_X3Y14_LUT4AB/S1BEG[3] Tile_X3Y14_LUT4AB/S1END[0] Tile_X3Y14_LUT4AB/S1END[1]
+ Tile_X3Y14_LUT4AB/S1END[2] Tile_X3Y14_LUT4AB/S1END[3] Tile_X3Y14_LUT4AB/S2BEG[0]
+ Tile_X3Y14_LUT4AB/S2BEG[1] Tile_X3Y14_LUT4AB/S2BEG[2] Tile_X3Y14_LUT4AB/S2BEG[3]
+ Tile_X3Y14_LUT4AB/S2BEG[4] Tile_X3Y14_LUT4AB/S2BEG[5] Tile_X3Y14_LUT4AB/S2BEG[6]
+ Tile_X3Y14_LUT4AB/S2BEG[7] Tile_X3Y14_LUT4AB/S2BEGb[0] Tile_X3Y14_LUT4AB/S2BEGb[1]
+ Tile_X3Y14_LUT4AB/S2BEGb[2] Tile_X3Y14_LUT4AB/S2BEGb[3] Tile_X3Y14_LUT4AB/S2BEGb[4]
+ Tile_X3Y14_LUT4AB/S2BEGb[5] Tile_X3Y14_LUT4AB/S2BEGb[6] Tile_X3Y14_LUT4AB/S2BEGb[7]
+ Tile_X3Y14_LUT4AB/S2END[0] Tile_X3Y14_LUT4AB/S2END[1] Tile_X3Y14_LUT4AB/S2END[2]
+ Tile_X3Y14_LUT4AB/S2END[3] Tile_X3Y14_LUT4AB/S2END[4] Tile_X3Y14_LUT4AB/S2END[5]
+ Tile_X3Y14_LUT4AB/S2END[6] Tile_X3Y14_LUT4AB/S2END[7] Tile_X3Y14_LUT4AB/S2MID[0]
+ Tile_X3Y14_LUT4AB/S2MID[1] Tile_X3Y14_LUT4AB/S2MID[2] Tile_X3Y14_LUT4AB/S2MID[3]
+ Tile_X3Y14_LUT4AB/S2MID[4] Tile_X3Y14_LUT4AB/S2MID[5] Tile_X3Y14_LUT4AB/S2MID[6]
+ Tile_X3Y14_LUT4AB/S2MID[7] Tile_X3Y14_LUT4AB/S4BEG[0] Tile_X3Y14_LUT4AB/S4BEG[10]
+ Tile_X3Y14_LUT4AB/S4BEG[11] Tile_X3Y14_LUT4AB/S4BEG[12] Tile_X3Y14_LUT4AB/S4BEG[13]
+ Tile_X3Y14_LUT4AB/S4BEG[14] Tile_X3Y14_LUT4AB/S4BEG[15] Tile_X3Y14_LUT4AB/S4BEG[1]
+ Tile_X3Y14_LUT4AB/S4BEG[2] Tile_X3Y14_LUT4AB/S4BEG[3] Tile_X3Y14_LUT4AB/S4BEG[4]
+ Tile_X3Y14_LUT4AB/S4BEG[5] Tile_X3Y14_LUT4AB/S4BEG[6] Tile_X3Y14_LUT4AB/S4BEG[7]
+ Tile_X3Y14_LUT4AB/S4BEG[8] Tile_X3Y14_LUT4AB/S4BEG[9] Tile_X3Y14_LUT4AB/S4END[0]
+ Tile_X3Y14_LUT4AB/S4END[10] Tile_X3Y14_LUT4AB/S4END[11] Tile_X3Y14_LUT4AB/S4END[12]
+ Tile_X3Y14_LUT4AB/S4END[13] Tile_X3Y14_LUT4AB/S4END[14] Tile_X3Y14_LUT4AB/S4END[15]
+ Tile_X3Y14_LUT4AB/S4END[1] Tile_X3Y14_LUT4AB/S4END[2] Tile_X3Y14_LUT4AB/S4END[3]
+ Tile_X3Y14_LUT4AB/S4END[4] Tile_X3Y14_LUT4AB/S4END[5] Tile_X3Y14_LUT4AB/S4END[6]
+ Tile_X3Y14_LUT4AB/S4END[7] Tile_X3Y14_LUT4AB/S4END[8] Tile_X3Y14_LUT4AB/S4END[9]
+ Tile_X3Y14_LUT4AB/SS4BEG[0] Tile_X3Y14_LUT4AB/SS4BEG[10] Tile_X3Y14_LUT4AB/SS4BEG[11]
+ Tile_X3Y14_LUT4AB/SS4BEG[12] Tile_X3Y14_LUT4AB/SS4BEG[13] Tile_X3Y14_LUT4AB/SS4BEG[14]
+ Tile_X3Y14_LUT4AB/SS4BEG[15] Tile_X3Y14_LUT4AB/SS4BEG[1] Tile_X3Y14_LUT4AB/SS4BEG[2]
+ Tile_X3Y14_LUT4AB/SS4BEG[3] Tile_X3Y14_LUT4AB/SS4BEG[4] Tile_X3Y14_LUT4AB/SS4BEG[5]
+ Tile_X3Y14_LUT4AB/SS4BEG[6] Tile_X3Y14_LUT4AB/SS4BEG[7] Tile_X3Y14_LUT4AB/SS4BEG[8]
+ Tile_X3Y14_LUT4AB/SS4BEG[9] Tile_X3Y14_LUT4AB/SS4END[0] Tile_X3Y14_LUT4AB/SS4END[10]
+ Tile_X3Y14_LUT4AB/SS4END[11] Tile_X3Y14_LUT4AB/SS4END[12] Tile_X3Y14_LUT4AB/SS4END[13]
+ Tile_X3Y14_LUT4AB/SS4END[14] Tile_X3Y14_LUT4AB/SS4END[15] Tile_X3Y14_LUT4AB/SS4END[1]
+ Tile_X3Y14_LUT4AB/SS4END[2] Tile_X3Y14_LUT4AB/SS4END[3] Tile_X3Y14_LUT4AB/SS4END[4]
+ Tile_X3Y14_LUT4AB/SS4END[5] Tile_X3Y14_LUT4AB/SS4END[6] Tile_X3Y14_LUT4AB/SS4END[7]
+ Tile_X3Y14_LUT4AB/SS4END[8] Tile_X3Y14_LUT4AB/SS4END[9] Tile_X3Y14_LUT4AB/UserCLK
+ Tile_X3Y13_LUT4AB/UserCLK VGND VPWR Tile_X3Y14_LUT4AB/W1BEG[0] Tile_X3Y14_LUT4AB/W1BEG[1]
+ Tile_X3Y14_LUT4AB/W1BEG[2] Tile_X3Y14_LUT4AB/W1BEG[3] Tile_X3Y14_LUT4AB/W1END[0]
+ Tile_X3Y14_LUT4AB/W1END[1] Tile_X3Y14_LUT4AB/W1END[2] Tile_X3Y14_LUT4AB/W1END[3]
+ Tile_X3Y14_LUT4AB/W2BEG[0] Tile_X3Y14_LUT4AB/W2BEG[1] Tile_X3Y14_LUT4AB/W2BEG[2]
+ Tile_X3Y14_LUT4AB/W2BEG[3] Tile_X3Y14_LUT4AB/W2BEG[4] Tile_X3Y14_LUT4AB/W2BEG[5]
+ Tile_X3Y14_LUT4AB/W2BEG[6] Tile_X3Y14_LUT4AB/W2BEG[7] Tile_X2Y14_LUT4AB/W2END[0]
+ Tile_X2Y14_LUT4AB/W2END[1] Tile_X2Y14_LUT4AB/W2END[2] Tile_X2Y14_LUT4AB/W2END[3]
+ Tile_X2Y14_LUT4AB/W2END[4] Tile_X2Y14_LUT4AB/W2END[5] Tile_X2Y14_LUT4AB/W2END[6]
+ Tile_X2Y14_LUT4AB/W2END[7] Tile_X3Y14_LUT4AB/W2END[0] Tile_X3Y14_LUT4AB/W2END[1]
+ Tile_X3Y14_LUT4AB/W2END[2] Tile_X3Y14_LUT4AB/W2END[3] Tile_X3Y14_LUT4AB/W2END[4]
+ Tile_X3Y14_LUT4AB/W2END[5] Tile_X3Y14_LUT4AB/W2END[6] Tile_X3Y14_LUT4AB/W2END[7]
+ Tile_X3Y14_LUT4AB/W2MID[0] Tile_X3Y14_LUT4AB/W2MID[1] Tile_X3Y14_LUT4AB/W2MID[2]
+ Tile_X3Y14_LUT4AB/W2MID[3] Tile_X3Y14_LUT4AB/W2MID[4] Tile_X3Y14_LUT4AB/W2MID[5]
+ Tile_X3Y14_LUT4AB/W2MID[6] Tile_X3Y14_LUT4AB/W2MID[7] Tile_X3Y14_LUT4AB/W6BEG[0]
+ Tile_X3Y14_LUT4AB/W6BEG[10] Tile_X3Y14_LUT4AB/W6BEG[11] Tile_X3Y14_LUT4AB/W6BEG[1]
+ Tile_X3Y14_LUT4AB/W6BEG[2] Tile_X3Y14_LUT4AB/W6BEG[3] Tile_X3Y14_LUT4AB/W6BEG[4]
+ Tile_X3Y14_LUT4AB/W6BEG[5] Tile_X3Y14_LUT4AB/W6BEG[6] Tile_X3Y14_LUT4AB/W6BEG[7]
+ Tile_X3Y14_LUT4AB/W6BEG[8] Tile_X3Y14_LUT4AB/W6BEG[9] Tile_X3Y14_LUT4AB/W6END[0]
+ Tile_X3Y14_LUT4AB/W6END[10] Tile_X3Y14_LUT4AB/W6END[11] Tile_X3Y14_LUT4AB/W6END[1]
+ Tile_X3Y14_LUT4AB/W6END[2] Tile_X3Y14_LUT4AB/W6END[3] Tile_X3Y14_LUT4AB/W6END[4]
+ Tile_X3Y14_LUT4AB/W6END[5] Tile_X3Y14_LUT4AB/W6END[6] Tile_X3Y14_LUT4AB/W6END[7]
+ Tile_X3Y14_LUT4AB/W6END[8] Tile_X3Y14_LUT4AB/W6END[9] Tile_X3Y14_LUT4AB/WW4BEG[0]
+ Tile_X3Y14_LUT4AB/WW4BEG[10] Tile_X3Y14_LUT4AB/WW4BEG[11] Tile_X3Y14_LUT4AB/WW4BEG[12]
+ Tile_X3Y14_LUT4AB/WW4BEG[13] Tile_X3Y14_LUT4AB/WW4BEG[14] Tile_X3Y14_LUT4AB/WW4BEG[15]
+ Tile_X3Y14_LUT4AB/WW4BEG[1] Tile_X3Y14_LUT4AB/WW4BEG[2] Tile_X3Y14_LUT4AB/WW4BEG[3]
+ Tile_X3Y14_LUT4AB/WW4BEG[4] Tile_X3Y14_LUT4AB/WW4BEG[5] Tile_X3Y14_LUT4AB/WW4BEG[6]
+ Tile_X3Y14_LUT4AB/WW4BEG[7] Tile_X3Y14_LUT4AB/WW4BEG[8] Tile_X3Y14_LUT4AB/WW4BEG[9]
+ Tile_X3Y14_LUT4AB/WW4END[0] Tile_X3Y14_LUT4AB/WW4END[10] Tile_X3Y14_LUT4AB/WW4END[11]
+ Tile_X3Y14_LUT4AB/WW4END[12] Tile_X3Y14_LUT4AB/WW4END[13] Tile_X3Y14_LUT4AB/WW4END[14]
+ Tile_X3Y14_LUT4AB/WW4END[15] Tile_X3Y14_LUT4AB/WW4END[1] Tile_X3Y14_LUT4AB/WW4END[2]
+ Tile_X3Y14_LUT4AB/WW4END[3] Tile_X3Y14_LUT4AB/WW4END[4] Tile_X3Y14_LUT4AB/WW4END[5]
+ Tile_X3Y14_LUT4AB/WW4END[6] Tile_X3Y14_LUT4AB/WW4END[7] Tile_X3Y14_LUT4AB/WW4END[8]
+ Tile_X3Y14_LUT4AB/WW4END[9] LUT4AB
XTile_X9Y11_LUT4AB Tile_X9Y12_LUT4AB/Co Tile_X9Y11_LUT4AB/Co Tile_X9Y11_LUT4AB/E1BEG[0]
+ Tile_X9Y11_LUT4AB/E1BEG[1] Tile_X9Y11_LUT4AB/E1BEG[2] Tile_X9Y11_LUT4AB/E1BEG[3]
+ Tile_X9Y11_LUT4AB/E1END[0] Tile_X9Y11_LUT4AB/E1END[1] Tile_X9Y11_LUT4AB/E1END[2]
+ Tile_X9Y11_LUT4AB/E1END[3] Tile_X9Y11_LUT4AB/E2BEG[0] Tile_X9Y11_LUT4AB/E2BEG[1]
+ Tile_X9Y11_LUT4AB/E2BEG[2] Tile_X9Y11_LUT4AB/E2BEG[3] Tile_X9Y11_LUT4AB/E2BEG[4]
+ Tile_X9Y11_LUT4AB/E2BEG[5] Tile_X9Y11_LUT4AB/E2BEG[6] Tile_X9Y11_LUT4AB/E2BEG[7]
+ Tile_X9Y11_LUT4AB/E2BEGb[0] Tile_X9Y11_LUT4AB/E2BEGb[1] Tile_X9Y11_LUT4AB/E2BEGb[2]
+ Tile_X9Y11_LUT4AB/E2BEGb[3] Tile_X9Y11_LUT4AB/E2BEGb[4] Tile_X9Y11_LUT4AB/E2BEGb[5]
+ Tile_X9Y11_LUT4AB/E2BEGb[6] Tile_X9Y11_LUT4AB/E2BEGb[7] Tile_X9Y11_LUT4AB/E2END[0]
+ Tile_X9Y11_LUT4AB/E2END[1] Tile_X9Y11_LUT4AB/E2END[2] Tile_X9Y11_LUT4AB/E2END[3]
+ Tile_X9Y11_LUT4AB/E2END[4] Tile_X9Y11_LUT4AB/E2END[5] Tile_X9Y11_LUT4AB/E2END[6]
+ Tile_X9Y11_LUT4AB/E2END[7] Tile_X9Y11_LUT4AB/E2MID[0] Tile_X9Y11_LUT4AB/E2MID[1]
+ Tile_X9Y11_LUT4AB/E2MID[2] Tile_X9Y11_LUT4AB/E2MID[3] Tile_X9Y11_LUT4AB/E2MID[4]
+ Tile_X9Y11_LUT4AB/E2MID[5] Tile_X9Y11_LUT4AB/E2MID[6] Tile_X9Y11_LUT4AB/E2MID[7]
+ Tile_X9Y11_LUT4AB/E6BEG[0] Tile_X9Y11_LUT4AB/E6BEG[10] Tile_X9Y11_LUT4AB/E6BEG[11]
+ Tile_X9Y11_LUT4AB/E6BEG[1] Tile_X9Y11_LUT4AB/E6BEG[2] Tile_X9Y11_LUT4AB/E6BEG[3]
+ Tile_X9Y11_LUT4AB/E6BEG[4] Tile_X9Y11_LUT4AB/E6BEG[5] Tile_X9Y11_LUT4AB/E6BEG[6]
+ Tile_X9Y11_LUT4AB/E6BEG[7] Tile_X9Y11_LUT4AB/E6BEG[8] Tile_X9Y11_LUT4AB/E6BEG[9]
+ Tile_X9Y11_LUT4AB/E6END[0] Tile_X9Y11_LUT4AB/E6END[10] Tile_X9Y11_LUT4AB/E6END[11]
+ Tile_X9Y11_LUT4AB/E6END[1] Tile_X9Y11_LUT4AB/E6END[2] Tile_X9Y11_LUT4AB/E6END[3]
+ Tile_X9Y11_LUT4AB/E6END[4] Tile_X9Y11_LUT4AB/E6END[5] Tile_X9Y11_LUT4AB/E6END[6]
+ Tile_X9Y11_LUT4AB/E6END[7] Tile_X9Y11_LUT4AB/E6END[8] Tile_X9Y11_LUT4AB/E6END[9]
+ Tile_X9Y11_LUT4AB/EE4BEG[0] Tile_X9Y11_LUT4AB/EE4BEG[10] Tile_X9Y11_LUT4AB/EE4BEG[11]
+ Tile_X9Y11_LUT4AB/EE4BEG[12] Tile_X9Y11_LUT4AB/EE4BEG[13] Tile_X9Y11_LUT4AB/EE4BEG[14]
+ Tile_X9Y11_LUT4AB/EE4BEG[15] Tile_X9Y11_LUT4AB/EE4BEG[1] Tile_X9Y11_LUT4AB/EE4BEG[2]
+ Tile_X9Y11_LUT4AB/EE4BEG[3] Tile_X9Y11_LUT4AB/EE4BEG[4] Tile_X9Y11_LUT4AB/EE4BEG[5]
+ Tile_X9Y11_LUT4AB/EE4BEG[6] Tile_X9Y11_LUT4AB/EE4BEG[7] Tile_X9Y11_LUT4AB/EE4BEG[8]
+ Tile_X9Y11_LUT4AB/EE4BEG[9] Tile_X9Y11_LUT4AB/EE4END[0] Tile_X9Y11_LUT4AB/EE4END[10]
+ Tile_X9Y11_LUT4AB/EE4END[11] Tile_X9Y11_LUT4AB/EE4END[12] Tile_X9Y11_LUT4AB/EE4END[13]
+ Tile_X9Y11_LUT4AB/EE4END[14] Tile_X9Y11_LUT4AB/EE4END[15] Tile_X9Y11_LUT4AB/EE4END[1]
+ Tile_X9Y11_LUT4AB/EE4END[2] Tile_X9Y11_LUT4AB/EE4END[3] Tile_X9Y11_LUT4AB/EE4END[4]
+ Tile_X9Y11_LUT4AB/EE4END[5] Tile_X9Y11_LUT4AB/EE4END[6] Tile_X9Y11_LUT4AB/EE4END[7]
+ Tile_X9Y11_LUT4AB/EE4END[8] Tile_X9Y11_LUT4AB/EE4END[9] Tile_X9Y11_LUT4AB/FrameData[0]
+ Tile_X9Y11_LUT4AB/FrameData[10] Tile_X9Y11_LUT4AB/FrameData[11] Tile_X9Y11_LUT4AB/FrameData[12]
+ Tile_X9Y11_LUT4AB/FrameData[13] Tile_X9Y11_LUT4AB/FrameData[14] Tile_X9Y11_LUT4AB/FrameData[15]
+ Tile_X9Y11_LUT4AB/FrameData[16] Tile_X9Y11_LUT4AB/FrameData[17] Tile_X9Y11_LUT4AB/FrameData[18]
+ Tile_X9Y11_LUT4AB/FrameData[19] Tile_X9Y11_LUT4AB/FrameData[1] Tile_X9Y11_LUT4AB/FrameData[20]
+ Tile_X9Y11_LUT4AB/FrameData[21] Tile_X9Y11_LUT4AB/FrameData[22] Tile_X9Y11_LUT4AB/FrameData[23]
+ Tile_X9Y11_LUT4AB/FrameData[24] Tile_X9Y11_LUT4AB/FrameData[25] Tile_X9Y11_LUT4AB/FrameData[26]
+ Tile_X9Y11_LUT4AB/FrameData[27] Tile_X9Y11_LUT4AB/FrameData[28] Tile_X9Y11_LUT4AB/FrameData[29]
+ Tile_X9Y11_LUT4AB/FrameData[2] Tile_X9Y11_LUT4AB/FrameData[30] Tile_X9Y11_LUT4AB/FrameData[31]
+ Tile_X9Y11_LUT4AB/FrameData[3] Tile_X9Y11_LUT4AB/FrameData[4] Tile_X9Y11_LUT4AB/FrameData[5]
+ Tile_X9Y11_LUT4AB/FrameData[6] Tile_X9Y11_LUT4AB/FrameData[7] Tile_X9Y11_LUT4AB/FrameData[8]
+ Tile_X9Y11_LUT4AB/FrameData[9] Tile_X9Y11_LUT4AB/FrameData_O[0] Tile_X9Y11_LUT4AB/FrameData_O[10]
+ Tile_X9Y11_LUT4AB/FrameData_O[11] Tile_X9Y11_LUT4AB/FrameData_O[12] Tile_X9Y11_LUT4AB/FrameData_O[13]
+ Tile_X9Y11_LUT4AB/FrameData_O[14] Tile_X9Y11_LUT4AB/FrameData_O[15] Tile_X9Y11_LUT4AB/FrameData_O[16]
+ Tile_X9Y11_LUT4AB/FrameData_O[17] Tile_X9Y11_LUT4AB/FrameData_O[18] Tile_X9Y11_LUT4AB/FrameData_O[19]
+ Tile_X9Y11_LUT4AB/FrameData_O[1] Tile_X9Y11_LUT4AB/FrameData_O[20] Tile_X9Y11_LUT4AB/FrameData_O[21]
+ Tile_X9Y11_LUT4AB/FrameData_O[22] Tile_X9Y11_LUT4AB/FrameData_O[23] Tile_X9Y11_LUT4AB/FrameData_O[24]
+ Tile_X9Y11_LUT4AB/FrameData_O[25] Tile_X9Y11_LUT4AB/FrameData_O[26] Tile_X9Y11_LUT4AB/FrameData_O[27]
+ Tile_X9Y11_LUT4AB/FrameData_O[28] Tile_X9Y11_LUT4AB/FrameData_O[29] Tile_X9Y11_LUT4AB/FrameData_O[2]
+ Tile_X9Y11_LUT4AB/FrameData_O[30] Tile_X9Y11_LUT4AB/FrameData_O[31] Tile_X9Y11_LUT4AB/FrameData_O[3]
+ Tile_X9Y11_LUT4AB/FrameData_O[4] Tile_X9Y11_LUT4AB/FrameData_O[5] Tile_X9Y11_LUT4AB/FrameData_O[6]
+ Tile_X9Y11_LUT4AB/FrameData_O[7] Tile_X9Y11_LUT4AB/FrameData_O[8] Tile_X9Y11_LUT4AB/FrameData_O[9]
+ Tile_X9Y11_LUT4AB/FrameStrobe[0] Tile_X9Y11_LUT4AB/FrameStrobe[10] Tile_X9Y11_LUT4AB/FrameStrobe[11]
+ Tile_X9Y11_LUT4AB/FrameStrobe[12] Tile_X9Y11_LUT4AB/FrameStrobe[13] Tile_X9Y11_LUT4AB/FrameStrobe[14]
+ Tile_X9Y11_LUT4AB/FrameStrobe[15] Tile_X9Y11_LUT4AB/FrameStrobe[16] Tile_X9Y11_LUT4AB/FrameStrobe[17]
+ Tile_X9Y11_LUT4AB/FrameStrobe[18] Tile_X9Y11_LUT4AB/FrameStrobe[19] Tile_X9Y11_LUT4AB/FrameStrobe[1]
+ Tile_X9Y11_LUT4AB/FrameStrobe[2] Tile_X9Y11_LUT4AB/FrameStrobe[3] Tile_X9Y11_LUT4AB/FrameStrobe[4]
+ Tile_X9Y11_LUT4AB/FrameStrobe[5] Tile_X9Y11_LUT4AB/FrameStrobe[6] Tile_X9Y11_LUT4AB/FrameStrobe[7]
+ Tile_X9Y11_LUT4AB/FrameStrobe[8] Tile_X9Y11_LUT4AB/FrameStrobe[9] Tile_X9Y10_LUT4AB/FrameStrobe[0]
+ Tile_X9Y10_LUT4AB/FrameStrobe[10] Tile_X9Y10_LUT4AB/FrameStrobe[11] Tile_X9Y10_LUT4AB/FrameStrobe[12]
+ Tile_X9Y10_LUT4AB/FrameStrobe[13] Tile_X9Y10_LUT4AB/FrameStrobe[14] Tile_X9Y10_LUT4AB/FrameStrobe[15]
+ Tile_X9Y10_LUT4AB/FrameStrobe[16] Tile_X9Y10_LUT4AB/FrameStrobe[17] Tile_X9Y10_LUT4AB/FrameStrobe[18]
+ Tile_X9Y10_LUT4AB/FrameStrobe[19] Tile_X9Y10_LUT4AB/FrameStrobe[1] Tile_X9Y10_LUT4AB/FrameStrobe[2]
+ Tile_X9Y10_LUT4AB/FrameStrobe[3] Tile_X9Y10_LUT4AB/FrameStrobe[4] Tile_X9Y10_LUT4AB/FrameStrobe[5]
+ Tile_X9Y10_LUT4AB/FrameStrobe[6] Tile_X9Y10_LUT4AB/FrameStrobe[7] Tile_X9Y10_LUT4AB/FrameStrobe[8]
+ Tile_X9Y10_LUT4AB/FrameStrobe[9] Tile_X9Y11_LUT4AB/N1BEG[0] Tile_X9Y11_LUT4AB/N1BEG[1]
+ Tile_X9Y11_LUT4AB/N1BEG[2] Tile_X9Y11_LUT4AB/N1BEG[3] Tile_X9Y12_LUT4AB/N1BEG[0]
+ Tile_X9Y12_LUT4AB/N1BEG[1] Tile_X9Y12_LUT4AB/N1BEG[2] Tile_X9Y12_LUT4AB/N1BEG[3]
+ Tile_X9Y11_LUT4AB/N2BEG[0] Tile_X9Y11_LUT4AB/N2BEG[1] Tile_X9Y11_LUT4AB/N2BEG[2]
+ Tile_X9Y11_LUT4AB/N2BEG[3] Tile_X9Y11_LUT4AB/N2BEG[4] Tile_X9Y11_LUT4AB/N2BEG[5]
+ Tile_X9Y11_LUT4AB/N2BEG[6] Tile_X9Y11_LUT4AB/N2BEG[7] Tile_X9Y10_LUT4AB/N2END[0]
+ Tile_X9Y10_LUT4AB/N2END[1] Tile_X9Y10_LUT4AB/N2END[2] Tile_X9Y10_LUT4AB/N2END[3]
+ Tile_X9Y10_LUT4AB/N2END[4] Tile_X9Y10_LUT4AB/N2END[5] Tile_X9Y10_LUT4AB/N2END[6]
+ Tile_X9Y10_LUT4AB/N2END[7] Tile_X9Y11_LUT4AB/N2END[0] Tile_X9Y11_LUT4AB/N2END[1]
+ Tile_X9Y11_LUT4AB/N2END[2] Tile_X9Y11_LUT4AB/N2END[3] Tile_X9Y11_LUT4AB/N2END[4]
+ Tile_X9Y11_LUT4AB/N2END[5] Tile_X9Y11_LUT4AB/N2END[6] Tile_X9Y11_LUT4AB/N2END[7]
+ Tile_X9Y12_LUT4AB/N2BEG[0] Tile_X9Y12_LUT4AB/N2BEG[1] Tile_X9Y12_LUT4AB/N2BEG[2]
+ Tile_X9Y12_LUT4AB/N2BEG[3] Tile_X9Y12_LUT4AB/N2BEG[4] Tile_X9Y12_LUT4AB/N2BEG[5]
+ Tile_X9Y12_LUT4AB/N2BEG[6] Tile_X9Y12_LUT4AB/N2BEG[7] Tile_X9Y11_LUT4AB/N4BEG[0]
+ Tile_X9Y11_LUT4AB/N4BEG[10] Tile_X9Y11_LUT4AB/N4BEG[11] Tile_X9Y11_LUT4AB/N4BEG[12]
+ Tile_X9Y11_LUT4AB/N4BEG[13] Tile_X9Y11_LUT4AB/N4BEG[14] Tile_X9Y11_LUT4AB/N4BEG[15]
+ Tile_X9Y11_LUT4AB/N4BEG[1] Tile_X9Y11_LUT4AB/N4BEG[2] Tile_X9Y11_LUT4AB/N4BEG[3]
+ Tile_X9Y11_LUT4AB/N4BEG[4] Tile_X9Y11_LUT4AB/N4BEG[5] Tile_X9Y11_LUT4AB/N4BEG[6]
+ Tile_X9Y11_LUT4AB/N4BEG[7] Tile_X9Y11_LUT4AB/N4BEG[8] Tile_X9Y11_LUT4AB/N4BEG[9]
+ Tile_X9Y12_LUT4AB/N4BEG[0] Tile_X9Y12_LUT4AB/N4BEG[10] Tile_X9Y12_LUT4AB/N4BEG[11]
+ Tile_X9Y12_LUT4AB/N4BEG[12] Tile_X9Y12_LUT4AB/N4BEG[13] Tile_X9Y12_LUT4AB/N4BEG[14]
+ Tile_X9Y12_LUT4AB/N4BEG[15] Tile_X9Y12_LUT4AB/N4BEG[1] Tile_X9Y12_LUT4AB/N4BEG[2]
+ Tile_X9Y12_LUT4AB/N4BEG[3] Tile_X9Y12_LUT4AB/N4BEG[4] Tile_X9Y12_LUT4AB/N4BEG[5]
+ Tile_X9Y12_LUT4AB/N4BEG[6] Tile_X9Y12_LUT4AB/N4BEG[7] Tile_X9Y12_LUT4AB/N4BEG[8]
+ Tile_X9Y12_LUT4AB/N4BEG[9] Tile_X9Y11_LUT4AB/NN4BEG[0] Tile_X9Y11_LUT4AB/NN4BEG[10]
+ Tile_X9Y11_LUT4AB/NN4BEG[11] Tile_X9Y11_LUT4AB/NN4BEG[12] Tile_X9Y11_LUT4AB/NN4BEG[13]
+ Tile_X9Y11_LUT4AB/NN4BEG[14] Tile_X9Y11_LUT4AB/NN4BEG[15] Tile_X9Y11_LUT4AB/NN4BEG[1]
+ Tile_X9Y11_LUT4AB/NN4BEG[2] Tile_X9Y11_LUT4AB/NN4BEG[3] Tile_X9Y11_LUT4AB/NN4BEG[4]
+ Tile_X9Y11_LUT4AB/NN4BEG[5] Tile_X9Y11_LUT4AB/NN4BEG[6] Tile_X9Y11_LUT4AB/NN4BEG[7]
+ Tile_X9Y11_LUT4AB/NN4BEG[8] Tile_X9Y11_LUT4AB/NN4BEG[9] Tile_X9Y12_LUT4AB/NN4BEG[0]
+ Tile_X9Y12_LUT4AB/NN4BEG[10] Tile_X9Y12_LUT4AB/NN4BEG[11] Tile_X9Y12_LUT4AB/NN4BEG[12]
+ Tile_X9Y12_LUT4AB/NN4BEG[13] Tile_X9Y12_LUT4AB/NN4BEG[14] Tile_X9Y12_LUT4AB/NN4BEG[15]
+ Tile_X9Y12_LUT4AB/NN4BEG[1] Tile_X9Y12_LUT4AB/NN4BEG[2] Tile_X9Y12_LUT4AB/NN4BEG[3]
+ Tile_X9Y12_LUT4AB/NN4BEG[4] Tile_X9Y12_LUT4AB/NN4BEG[5] Tile_X9Y12_LUT4AB/NN4BEG[6]
+ Tile_X9Y12_LUT4AB/NN4BEG[7] Tile_X9Y12_LUT4AB/NN4BEG[8] Tile_X9Y12_LUT4AB/NN4BEG[9]
+ Tile_X9Y12_LUT4AB/S1END[0] Tile_X9Y12_LUT4AB/S1END[1] Tile_X9Y12_LUT4AB/S1END[2]
+ Tile_X9Y12_LUT4AB/S1END[3] Tile_X9Y11_LUT4AB/S1END[0] Tile_X9Y11_LUT4AB/S1END[1]
+ Tile_X9Y11_LUT4AB/S1END[2] Tile_X9Y11_LUT4AB/S1END[3] Tile_X9Y12_LUT4AB/S2MID[0]
+ Tile_X9Y12_LUT4AB/S2MID[1] Tile_X9Y12_LUT4AB/S2MID[2] Tile_X9Y12_LUT4AB/S2MID[3]
+ Tile_X9Y12_LUT4AB/S2MID[4] Tile_X9Y12_LUT4AB/S2MID[5] Tile_X9Y12_LUT4AB/S2MID[6]
+ Tile_X9Y12_LUT4AB/S2MID[7] Tile_X9Y12_LUT4AB/S2END[0] Tile_X9Y12_LUT4AB/S2END[1]
+ Tile_X9Y12_LUT4AB/S2END[2] Tile_X9Y12_LUT4AB/S2END[3] Tile_X9Y12_LUT4AB/S2END[4]
+ Tile_X9Y12_LUT4AB/S2END[5] Tile_X9Y12_LUT4AB/S2END[6] Tile_X9Y12_LUT4AB/S2END[7]
+ Tile_X9Y11_LUT4AB/S2END[0] Tile_X9Y11_LUT4AB/S2END[1] Tile_X9Y11_LUT4AB/S2END[2]
+ Tile_X9Y11_LUT4AB/S2END[3] Tile_X9Y11_LUT4AB/S2END[4] Tile_X9Y11_LUT4AB/S2END[5]
+ Tile_X9Y11_LUT4AB/S2END[6] Tile_X9Y11_LUT4AB/S2END[7] Tile_X9Y11_LUT4AB/S2MID[0]
+ Tile_X9Y11_LUT4AB/S2MID[1] Tile_X9Y11_LUT4AB/S2MID[2] Tile_X9Y11_LUT4AB/S2MID[3]
+ Tile_X9Y11_LUT4AB/S2MID[4] Tile_X9Y11_LUT4AB/S2MID[5] Tile_X9Y11_LUT4AB/S2MID[6]
+ Tile_X9Y11_LUT4AB/S2MID[7] Tile_X9Y12_LUT4AB/S4END[0] Tile_X9Y12_LUT4AB/S4END[10]
+ Tile_X9Y12_LUT4AB/S4END[11] Tile_X9Y12_LUT4AB/S4END[12] Tile_X9Y12_LUT4AB/S4END[13]
+ Tile_X9Y12_LUT4AB/S4END[14] Tile_X9Y12_LUT4AB/S4END[15] Tile_X9Y12_LUT4AB/S4END[1]
+ Tile_X9Y12_LUT4AB/S4END[2] Tile_X9Y12_LUT4AB/S4END[3] Tile_X9Y12_LUT4AB/S4END[4]
+ Tile_X9Y12_LUT4AB/S4END[5] Tile_X9Y12_LUT4AB/S4END[6] Tile_X9Y12_LUT4AB/S4END[7]
+ Tile_X9Y12_LUT4AB/S4END[8] Tile_X9Y12_LUT4AB/S4END[9] Tile_X9Y11_LUT4AB/S4END[0]
+ Tile_X9Y11_LUT4AB/S4END[10] Tile_X9Y11_LUT4AB/S4END[11] Tile_X9Y11_LUT4AB/S4END[12]
+ Tile_X9Y11_LUT4AB/S4END[13] Tile_X9Y11_LUT4AB/S4END[14] Tile_X9Y11_LUT4AB/S4END[15]
+ Tile_X9Y11_LUT4AB/S4END[1] Tile_X9Y11_LUT4AB/S4END[2] Tile_X9Y11_LUT4AB/S4END[3]
+ Tile_X9Y11_LUT4AB/S4END[4] Tile_X9Y11_LUT4AB/S4END[5] Tile_X9Y11_LUT4AB/S4END[6]
+ Tile_X9Y11_LUT4AB/S4END[7] Tile_X9Y11_LUT4AB/S4END[8] Tile_X9Y11_LUT4AB/S4END[9]
+ Tile_X9Y12_LUT4AB/SS4END[0] Tile_X9Y12_LUT4AB/SS4END[10] Tile_X9Y12_LUT4AB/SS4END[11]
+ Tile_X9Y12_LUT4AB/SS4END[12] Tile_X9Y12_LUT4AB/SS4END[13] Tile_X9Y12_LUT4AB/SS4END[14]
+ Tile_X9Y12_LUT4AB/SS4END[15] Tile_X9Y12_LUT4AB/SS4END[1] Tile_X9Y12_LUT4AB/SS4END[2]
+ Tile_X9Y12_LUT4AB/SS4END[3] Tile_X9Y12_LUT4AB/SS4END[4] Tile_X9Y12_LUT4AB/SS4END[5]
+ Tile_X9Y12_LUT4AB/SS4END[6] Tile_X9Y12_LUT4AB/SS4END[7] Tile_X9Y12_LUT4AB/SS4END[8]
+ Tile_X9Y12_LUT4AB/SS4END[9] Tile_X9Y11_LUT4AB/SS4END[0] Tile_X9Y11_LUT4AB/SS4END[10]
+ Tile_X9Y11_LUT4AB/SS4END[11] Tile_X9Y11_LUT4AB/SS4END[12] Tile_X9Y11_LUT4AB/SS4END[13]
+ Tile_X9Y11_LUT4AB/SS4END[14] Tile_X9Y11_LUT4AB/SS4END[15] Tile_X9Y11_LUT4AB/SS4END[1]
+ Tile_X9Y11_LUT4AB/SS4END[2] Tile_X9Y11_LUT4AB/SS4END[3] Tile_X9Y11_LUT4AB/SS4END[4]
+ Tile_X9Y11_LUT4AB/SS4END[5] Tile_X9Y11_LUT4AB/SS4END[6] Tile_X9Y11_LUT4AB/SS4END[7]
+ Tile_X9Y11_LUT4AB/SS4END[8] Tile_X9Y11_LUT4AB/SS4END[9] Tile_X9Y11_LUT4AB/UserCLK
+ Tile_X9Y10_LUT4AB/UserCLK VGND VPWR Tile_X9Y11_LUT4AB/W1BEG[0] Tile_X9Y11_LUT4AB/W1BEG[1]
+ Tile_X9Y11_LUT4AB/W1BEG[2] Tile_X9Y11_LUT4AB/W1BEG[3] Tile_X9Y11_LUT4AB/W1END[0]
+ Tile_X9Y11_LUT4AB/W1END[1] Tile_X9Y11_LUT4AB/W1END[2] Tile_X9Y11_LUT4AB/W1END[3]
+ Tile_X9Y11_LUT4AB/W2BEG[0] Tile_X9Y11_LUT4AB/W2BEG[1] Tile_X9Y11_LUT4AB/W2BEG[2]
+ Tile_X9Y11_LUT4AB/W2BEG[3] Tile_X9Y11_LUT4AB/W2BEG[4] Tile_X9Y11_LUT4AB/W2BEG[5]
+ Tile_X9Y11_LUT4AB/W2BEG[6] Tile_X9Y11_LUT4AB/W2BEG[7] Tile_X8Y11_LUT4AB/W2END[0]
+ Tile_X8Y11_LUT4AB/W2END[1] Tile_X8Y11_LUT4AB/W2END[2] Tile_X8Y11_LUT4AB/W2END[3]
+ Tile_X8Y11_LUT4AB/W2END[4] Tile_X8Y11_LUT4AB/W2END[5] Tile_X8Y11_LUT4AB/W2END[6]
+ Tile_X8Y11_LUT4AB/W2END[7] Tile_X9Y11_LUT4AB/W2END[0] Tile_X9Y11_LUT4AB/W2END[1]
+ Tile_X9Y11_LUT4AB/W2END[2] Tile_X9Y11_LUT4AB/W2END[3] Tile_X9Y11_LUT4AB/W2END[4]
+ Tile_X9Y11_LUT4AB/W2END[5] Tile_X9Y11_LUT4AB/W2END[6] Tile_X9Y11_LUT4AB/W2END[7]
+ Tile_X9Y11_LUT4AB/W2MID[0] Tile_X9Y11_LUT4AB/W2MID[1] Tile_X9Y11_LUT4AB/W2MID[2]
+ Tile_X9Y11_LUT4AB/W2MID[3] Tile_X9Y11_LUT4AB/W2MID[4] Tile_X9Y11_LUT4AB/W2MID[5]
+ Tile_X9Y11_LUT4AB/W2MID[6] Tile_X9Y11_LUT4AB/W2MID[7] Tile_X9Y11_LUT4AB/W6BEG[0]
+ Tile_X9Y11_LUT4AB/W6BEG[10] Tile_X9Y11_LUT4AB/W6BEG[11] Tile_X9Y11_LUT4AB/W6BEG[1]
+ Tile_X9Y11_LUT4AB/W6BEG[2] Tile_X9Y11_LUT4AB/W6BEG[3] Tile_X9Y11_LUT4AB/W6BEG[4]
+ Tile_X9Y11_LUT4AB/W6BEG[5] Tile_X9Y11_LUT4AB/W6BEG[6] Tile_X9Y11_LUT4AB/W6BEG[7]
+ Tile_X9Y11_LUT4AB/W6BEG[8] Tile_X9Y11_LUT4AB/W6BEG[9] Tile_X9Y11_LUT4AB/W6END[0]
+ Tile_X9Y11_LUT4AB/W6END[10] Tile_X9Y11_LUT4AB/W6END[11] Tile_X9Y11_LUT4AB/W6END[1]
+ Tile_X9Y11_LUT4AB/W6END[2] Tile_X9Y11_LUT4AB/W6END[3] Tile_X9Y11_LUT4AB/W6END[4]
+ Tile_X9Y11_LUT4AB/W6END[5] Tile_X9Y11_LUT4AB/W6END[6] Tile_X9Y11_LUT4AB/W6END[7]
+ Tile_X9Y11_LUT4AB/W6END[8] Tile_X9Y11_LUT4AB/W6END[9] Tile_X9Y11_LUT4AB/WW4BEG[0]
+ Tile_X9Y11_LUT4AB/WW4BEG[10] Tile_X9Y11_LUT4AB/WW4BEG[11] Tile_X9Y11_LUT4AB/WW4BEG[12]
+ Tile_X9Y11_LUT4AB/WW4BEG[13] Tile_X9Y11_LUT4AB/WW4BEG[14] Tile_X9Y11_LUT4AB/WW4BEG[15]
+ Tile_X9Y11_LUT4AB/WW4BEG[1] Tile_X9Y11_LUT4AB/WW4BEG[2] Tile_X9Y11_LUT4AB/WW4BEG[3]
+ Tile_X9Y11_LUT4AB/WW4BEG[4] Tile_X9Y11_LUT4AB/WW4BEG[5] Tile_X9Y11_LUT4AB/WW4BEG[6]
+ Tile_X9Y11_LUT4AB/WW4BEG[7] Tile_X9Y11_LUT4AB/WW4BEG[8] Tile_X9Y11_LUT4AB/WW4BEG[9]
+ Tile_X9Y11_LUT4AB/WW4END[0] Tile_X9Y11_LUT4AB/WW4END[10] Tile_X9Y11_LUT4AB/WW4END[11]
+ Tile_X9Y11_LUT4AB/WW4END[12] Tile_X9Y11_LUT4AB/WW4END[13] Tile_X9Y11_LUT4AB/WW4END[14]
+ Tile_X9Y11_LUT4AB/WW4END[15] Tile_X9Y11_LUT4AB/WW4END[1] Tile_X9Y11_LUT4AB/WW4END[2]
+ Tile_X9Y11_LUT4AB/WW4END[3] Tile_X9Y11_LUT4AB/WW4END[4] Tile_X9Y11_LUT4AB/WW4END[5]
+ Tile_X9Y11_LUT4AB/WW4END[6] Tile_X9Y11_LUT4AB/WW4END[7] Tile_X9Y11_LUT4AB/WW4END[8]
+ Tile_X9Y11_LUT4AB/WW4END[9] LUT4AB
XTile_X3Y7_LUT4AB Tile_X3Y8_LUT4AB/Co Tile_X3Y7_LUT4AB/Co Tile_X3Y7_LUT4AB/E1BEG[0]
+ Tile_X3Y7_LUT4AB/E1BEG[1] Tile_X3Y7_LUT4AB/E1BEG[2] Tile_X3Y7_LUT4AB/E1BEG[3] Tile_X3Y7_LUT4AB/E1END[0]
+ Tile_X3Y7_LUT4AB/E1END[1] Tile_X3Y7_LUT4AB/E1END[2] Tile_X3Y7_LUT4AB/E1END[3] Tile_X3Y7_LUT4AB/E2BEG[0]
+ Tile_X3Y7_LUT4AB/E2BEG[1] Tile_X3Y7_LUT4AB/E2BEG[2] Tile_X3Y7_LUT4AB/E2BEG[3] Tile_X3Y7_LUT4AB/E2BEG[4]
+ Tile_X3Y7_LUT4AB/E2BEG[5] Tile_X3Y7_LUT4AB/E2BEG[6] Tile_X3Y7_LUT4AB/E2BEG[7] Tile_X4Y7_RegFile/E2END[0]
+ Tile_X4Y7_RegFile/E2END[1] Tile_X4Y7_RegFile/E2END[2] Tile_X4Y7_RegFile/E2END[3]
+ Tile_X4Y7_RegFile/E2END[4] Tile_X4Y7_RegFile/E2END[5] Tile_X4Y7_RegFile/E2END[6]
+ Tile_X4Y7_RegFile/E2END[7] Tile_X3Y7_LUT4AB/E2END[0] Tile_X3Y7_LUT4AB/E2END[1] Tile_X3Y7_LUT4AB/E2END[2]
+ Tile_X3Y7_LUT4AB/E2END[3] Tile_X3Y7_LUT4AB/E2END[4] Tile_X3Y7_LUT4AB/E2END[5] Tile_X3Y7_LUT4AB/E2END[6]
+ Tile_X3Y7_LUT4AB/E2END[7] Tile_X3Y7_LUT4AB/E2MID[0] Tile_X3Y7_LUT4AB/E2MID[1] Tile_X3Y7_LUT4AB/E2MID[2]
+ Tile_X3Y7_LUT4AB/E2MID[3] Tile_X3Y7_LUT4AB/E2MID[4] Tile_X3Y7_LUT4AB/E2MID[5] Tile_X3Y7_LUT4AB/E2MID[6]
+ Tile_X3Y7_LUT4AB/E2MID[7] Tile_X3Y7_LUT4AB/E6BEG[0] Tile_X3Y7_LUT4AB/E6BEG[10] Tile_X3Y7_LUT4AB/E6BEG[11]
+ Tile_X3Y7_LUT4AB/E6BEG[1] Tile_X3Y7_LUT4AB/E6BEG[2] Tile_X3Y7_LUT4AB/E6BEG[3] Tile_X3Y7_LUT4AB/E6BEG[4]
+ Tile_X3Y7_LUT4AB/E6BEG[5] Tile_X3Y7_LUT4AB/E6BEG[6] Tile_X3Y7_LUT4AB/E6BEG[7] Tile_X3Y7_LUT4AB/E6BEG[8]
+ Tile_X3Y7_LUT4AB/E6BEG[9] Tile_X3Y7_LUT4AB/E6END[0] Tile_X3Y7_LUT4AB/E6END[10] Tile_X3Y7_LUT4AB/E6END[11]
+ Tile_X3Y7_LUT4AB/E6END[1] Tile_X3Y7_LUT4AB/E6END[2] Tile_X3Y7_LUT4AB/E6END[3] Tile_X3Y7_LUT4AB/E6END[4]
+ Tile_X3Y7_LUT4AB/E6END[5] Tile_X3Y7_LUT4AB/E6END[6] Tile_X3Y7_LUT4AB/E6END[7] Tile_X3Y7_LUT4AB/E6END[8]
+ Tile_X3Y7_LUT4AB/E6END[9] Tile_X3Y7_LUT4AB/EE4BEG[0] Tile_X3Y7_LUT4AB/EE4BEG[10]
+ Tile_X3Y7_LUT4AB/EE4BEG[11] Tile_X3Y7_LUT4AB/EE4BEG[12] Tile_X3Y7_LUT4AB/EE4BEG[13]
+ Tile_X3Y7_LUT4AB/EE4BEG[14] Tile_X3Y7_LUT4AB/EE4BEG[15] Tile_X3Y7_LUT4AB/EE4BEG[1]
+ Tile_X3Y7_LUT4AB/EE4BEG[2] Tile_X3Y7_LUT4AB/EE4BEG[3] Tile_X3Y7_LUT4AB/EE4BEG[4]
+ Tile_X3Y7_LUT4AB/EE4BEG[5] Tile_X3Y7_LUT4AB/EE4BEG[6] Tile_X3Y7_LUT4AB/EE4BEG[7]
+ Tile_X3Y7_LUT4AB/EE4BEG[8] Tile_X3Y7_LUT4AB/EE4BEG[9] Tile_X3Y7_LUT4AB/EE4END[0]
+ Tile_X3Y7_LUT4AB/EE4END[10] Tile_X3Y7_LUT4AB/EE4END[11] Tile_X3Y7_LUT4AB/EE4END[12]
+ Tile_X3Y7_LUT4AB/EE4END[13] Tile_X3Y7_LUT4AB/EE4END[14] Tile_X3Y7_LUT4AB/EE4END[15]
+ Tile_X3Y7_LUT4AB/EE4END[1] Tile_X3Y7_LUT4AB/EE4END[2] Tile_X3Y7_LUT4AB/EE4END[3]
+ Tile_X3Y7_LUT4AB/EE4END[4] Tile_X3Y7_LUT4AB/EE4END[5] Tile_X3Y7_LUT4AB/EE4END[6]
+ Tile_X3Y7_LUT4AB/EE4END[7] Tile_X3Y7_LUT4AB/EE4END[8] Tile_X3Y7_LUT4AB/EE4END[9]
+ Tile_X3Y7_LUT4AB/FrameData[0] Tile_X3Y7_LUT4AB/FrameData[10] Tile_X3Y7_LUT4AB/FrameData[11]
+ Tile_X3Y7_LUT4AB/FrameData[12] Tile_X3Y7_LUT4AB/FrameData[13] Tile_X3Y7_LUT4AB/FrameData[14]
+ Tile_X3Y7_LUT4AB/FrameData[15] Tile_X3Y7_LUT4AB/FrameData[16] Tile_X3Y7_LUT4AB/FrameData[17]
+ Tile_X3Y7_LUT4AB/FrameData[18] Tile_X3Y7_LUT4AB/FrameData[19] Tile_X3Y7_LUT4AB/FrameData[1]
+ Tile_X3Y7_LUT4AB/FrameData[20] Tile_X3Y7_LUT4AB/FrameData[21] Tile_X3Y7_LUT4AB/FrameData[22]
+ Tile_X3Y7_LUT4AB/FrameData[23] Tile_X3Y7_LUT4AB/FrameData[24] Tile_X3Y7_LUT4AB/FrameData[25]
+ Tile_X3Y7_LUT4AB/FrameData[26] Tile_X3Y7_LUT4AB/FrameData[27] Tile_X3Y7_LUT4AB/FrameData[28]
+ Tile_X3Y7_LUT4AB/FrameData[29] Tile_X3Y7_LUT4AB/FrameData[2] Tile_X3Y7_LUT4AB/FrameData[30]
+ Tile_X3Y7_LUT4AB/FrameData[31] Tile_X3Y7_LUT4AB/FrameData[3] Tile_X3Y7_LUT4AB/FrameData[4]
+ Tile_X3Y7_LUT4AB/FrameData[5] Tile_X3Y7_LUT4AB/FrameData[6] Tile_X3Y7_LUT4AB/FrameData[7]
+ Tile_X3Y7_LUT4AB/FrameData[8] Tile_X3Y7_LUT4AB/FrameData[9] Tile_X4Y7_RegFile/FrameData[0]
+ Tile_X4Y7_RegFile/FrameData[10] Tile_X4Y7_RegFile/FrameData[11] Tile_X4Y7_RegFile/FrameData[12]
+ Tile_X4Y7_RegFile/FrameData[13] Tile_X4Y7_RegFile/FrameData[14] Tile_X4Y7_RegFile/FrameData[15]
+ Tile_X4Y7_RegFile/FrameData[16] Tile_X4Y7_RegFile/FrameData[17] Tile_X4Y7_RegFile/FrameData[18]
+ Tile_X4Y7_RegFile/FrameData[19] Tile_X4Y7_RegFile/FrameData[1] Tile_X4Y7_RegFile/FrameData[20]
+ Tile_X4Y7_RegFile/FrameData[21] Tile_X4Y7_RegFile/FrameData[22] Tile_X4Y7_RegFile/FrameData[23]
+ Tile_X4Y7_RegFile/FrameData[24] Tile_X4Y7_RegFile/FrameData[25] Tile_X4Y7_RegFile/FrameData[26]
+ Tile_X4Y7_RegFile/FrameData[27] Tile_X4Y7_RegFile/FrameData[28] Tile_X4Y7_RegFile/FrameData[29]
+ Tile_X4Y7_RegFile/FrameData[2] Tile_X4Y7_RegFile/FrameData[30] Tile_X4Y7_RegFile/FrameData[31]
+ Tile_X4Y7_RegFile/FrameData[3] Tile_X4Y7_RegFile/FrameData[4] Tile_X4Y7_RegFile/FrameData[5]
+ Tile_X4Y7_RegFile/FrameData[6] Tile_X4Y7_RegFile/FrameData[7] Tile_X4Y7_RegFile/FrameData[8]
+ Tile_X4Y7_RegFile/FrameData[9] Tile_X3Y7_LUT4AB/FrameStrobe[0] Tile_X3Y7_LUT4AB/FrameStrobe[10]
+ Tile_X3Y7_LUT4AB/FrameStrobe[11] Tile_X3Y7_LUT4AB/FrameStrobe[12] Tile_X3Y7_LUT4AB/FrameStrobe[13]
+ Tile_X3Y7_LUT4AB/FrameStrobe[14] Tile_X3Y7_LUT4AB/FrameStrobe[15] Tile_X3Y7_LUT4AB/FrameStrobe[16]
+ Tile_X3Y7_LUT4AB/FrameStrobe[17] Tile_X3Y7_LUT4AB/FrameStrobe[18] Tile_X3Y7_LUT4AB/FrameStrobe[19]
+ Tile_X3Y7_LUT4AB/FrameStrobe[1] Tile_X3Y7_LUT4AB/FrameStrobe[2] Tile_X3Y7_LUT4AB/FrameStrobe[3]
+ Tile_X3Y7_LUT4AB/FrameStrobe[4] Tile_X3Y7_LUT4AB/FrameStrobe[5] Tile_X3Y7_LUT4AB/FrameStrobe[6]
+ Tile_X3Y7_LUT4AB/FrameStrobe[7] Tile_X3Y7_LUT4AB/FrameStrobe[8] Tile_X3Y7_LUT4AB/FrameStrobe[9]
+ Tile_X3Y6_LUT4AB/FrameStrobe[0] Tile_X3Y6_LUT4AB/FrameStrobe[10] Tile_X3Y6_LUT4AB/FrameStrobe[11]
+ Tile_X3Y6_LUT4AB/FrameStrobe[12] Tile_X3Y6_LUT4AB/FrameStrobe[13] Tile_X3Y6_LUT4AB/FrameStrobe[14]
+ Tile_X3Y6_LUT4AB/FrameStrobe[15] Tile_X3Y6_LUT4AB/FrameStrobe[16] Tile_X3Y6_LUT4AB/FrameStrobe[17]
+ Tile_X3Y6_LUT4AB/FrameStrobe[18] Tile_X3Y6_LUT4AB/FrameStrobe[19] Tile_X3Y6_LUT4AB/FrameStrobe[1]
+ Tile_X3Y6_LUT4AB/FrameStrobe[2] Tile_X3Y6_LUT4AB/FrameStrobe[3] Tile_X3Y6_LUT4AB/FrameStrobe[4]
+ Tile_X3Y6_LUT4AB/FrameStrobe[5] Tile_X3Y6_LUT4AB/FrameStrobe[6] Tile_X3Y6_LUT4AB/FrameStrobe[7]
+ Tile_X3Y6_LUT4AB/FrameStrobe[8] Tile_X3Y6_LUT4AB/FrameStrobe[9] Tile_X3Y7_LUT4AB/N1BEG[0]
+ Tile_X3Y7_LUT4AB/N1BEG[1] Tile_X3Y7_LUT4AB/N1BEG[2] Tile_X3Y7_LUT4AB/N1BEG[3] Tile_X3Y8_LUT4AB/N1BEG[0]
+ Tile_X3Y8_LUT4AB/N1BEG[1] Tile_X3Y8_LUT4AB/N1BEG[2] Tile_X3Y8_LUT4AB/N1BEG[3] Tile_X3Y7_LUT4AB/N2BEG[0]
+ Tile_X3Y7_LUT4AB/N2BEG[1] Tile_X3Y7_LUT4AB/N2BEG[2] Tile_X3Y7_LUT4AB/N2BEG[3] Tile_X3Y7_LUT4AB/N2BEG[4]
+ Tile_X3Y7_LUT4AB/N2BEG[5] Tile_X3Y7_LUT4AB/N2BEG[6] Tile_X3Y7_LUT4AB/N2BEG[7] Tile_X3Y6_LUT4AB/N2END[0]
+ Tile_X3Y6_LUT4AB/N2END[1] Tile_X3Y6_LUT4AB/N2END[2] Tile_X3Y6_LUT4AB/N2END[3] Tile_X3Y6_LUT4AB/N2END[4]
+ Tile_X3Y6_LUT4AB/N2END[5] Tile_X3Y6_LUT4AB/N2END[6] Tile_X3Y6_LUT4AB/N2END[7] Tile_X3Y7_LUT4AB/N2END[0]
+ Tile_X3Y7_LUT4AB/N2END[1] Tile_X3Y7_LUT4AB/N2END[2] Tile_X3Y7_LUT4AB/N2END[3] Tile_X3Y7_LUT4AB/N2END[4]
+ Tile_X3Y7_LUT4AB/N2END[5] Tile_X3Y7_LUT4AB/N2END[6] Tile_X3Y7_LUT4AB/N2END[7] Tile_X3Y8_LUT4AB/N2BEG[0]
+ Tile_X3Y8_LUT4AB/N2BEG[1] Tile_X3Y8_LUT4AB/N2BEG[2] Tile_X3Y8_LUT4AB/N2BEG[3] Tile_X3Y8_LUT4AB/N2BEG[4]
+ Tile_X3Y8_LUT4AB/N2BEG[5] Tile_X3Y8_LUT4AB/N2BEG[6] Tile_X3Y8_LUT4AB/N2BEG[7] Tile_X3Y7_LUT4AB/N4BEG[0]
+ Tile_X3Y7_LUT4AB/N4BEG[10] Tile_X3Y7_LUT4AB/N4BEG[11] Tile_X3Y7_LUT4AB/N4BEG[12]
+ Tile_X3Y7_LUT4AB/N4BEG[13] Tile_X3Y7_LUT4AB/N4BEG[14] Tile_X3Y7_LUT4AB/N4BEG[15]
+ Tile_X3Y7_LUT4AB/N4BEG[1] Tile_X3Y7_LUT4AB/N4BEG[2] Tile_X3Y7_LUT4AB/N4BEG[3] Tile_X3Y7_LUT4AB/N4BEG[4]
+ Tile_X3Y7_LUT4AB/N4BEG[5] Tile_X3Y7_LUT4AB/N4BEG[6] Tile_X3Y7_LUT4AB/N4BEG[7] Tile_X3Y7_LUT4AB/N4BEG[8]
+ Tile_X3Y7_LUT4AB/N4BEG[9] Tile_X3Y8_LUT4AB/N4BEG[0] Tile_X3Y8_LUT4AB/N4BEG[10] Tile_X3Y8_LUT4AB/N4BEG[11]
+ Tile_X3Y8_LUT4AB/N4BEG[12] Tile_X3Y8_LUT4AB/N4BEG[13] Tile_X3Y8_LUT4AB/N4BEG[14]
+ Tile_X3Y8_LUT4AB/N4BEG[15] Tile_X3Y8_LUT4AB/N4BEG[1] Tile_X3Y8_LUT4AB/N4BEG[2] Tile_X3Y8_LUT4AB/N4BEG[3]
+ Tile_X3Y8_LUT4AB/N4BEG[4] Tile_X3Y8_LUT4AB/N4BEG[5] Tile_X3Y8_LUT4AB/N4BEG[6] Tile_X3Y8_LUT4AB/N4BEG[7]
+ Tile_X3Y8_LUT4AB/N4BEG[8] Tile_X3Y8_LUT4AB/N4BEG[9] Tile_X3Y7_LUT4AB/NN4BEG[0] Tile_X3Y7_LUT4AB/NN4BEG[10]
+ Tile_X3Y7_LUT4AB/NN4BEG[11] Tile_X3Y7_LUT4AB/NN4BEG[12] Tile_X3Y7_LUT4AB/NN4BEG[13]
+ Tile_X3Y7_LUT4AB/NN4BEG[14] Tile_X3Y7_LUT4AB/NN4BEG[15] Tile_X3Y7_LUT4AB/NN4BEG[1]
+ Tile_X3Y7_LUT4AB/NN4BEG[2] Tile_X3Y7_LUT4AB/NN4BEG[3] Tile_X3Y7_LUT4AB/NN4BEG[4]
+ Tile_X3Y7_LUT4AB/NN4BEG[5] Tile_X3Y7_LUT4AB/NN4BEG[6] Tile_X3Y7_LUT4AB/NN4BEG[7]
+ Tile_X3Y7_LUT4AB/NN4BEG[8] Tile_X3Y7_LUT4AB/NN4BEG[9] Tile_X3Y8_LUT4AB/NN4BEG[0]
+ Tile_X3Y8_LUT4AB/NN4BEG[10] Tile_X3Y8_LUT4AB/NN4BEG[11] Tile_X3Y8_LUT4AB/NN4BEG[12]
+ Tile_X3Y8_LUT4AB/NN4BEG[13] Tile_X3Y8_LUT4AB/NN4BEG[14] Tile_X3Y8_LUT4AB/NN4BEG[15]
+ Tile_X3Y8_LUT4AB/NN4BEG[1] Tile_X3Y8_LUT4AB/NN4BEG[2] Tile_X3Y8_LUT4AB/NN4BEG[3]
+ Tile_X3Y8_LUT4AB/NN4BEG[4] Tile_X3Y8_LUT4AB/NN4BEG[5] Tile_X3Y8_LUT4AB/NN4BEG[6]
+ Tile_X3Y8_LUT4AB/NN4BEG[7] Tile_X3Y8_LUT4AB/NN4BEG[8] Tile_X3Y8_LUT4AB/NN4BEG[9]
+ Tile_X3Y8_LUT4AB/S1END[0] Tile_X3Y8_LUT4AB/S1END[1] Tile_X3Y8_LUT4AB/S1END[2] Tile_X3Y8_LUT4AB/S1END[3]
+ Tile_X3Y7_LUT4AB/S1END[0] Tile_X3Y7_LUT4AB/S1END[1] Tile_X3Y7_LUT4AB/S1END[2] Tile_X3Y7_LUT4AB/S1END[3]
+ Tile_X3Y8_LUT4AB/S2MID[0] Tile_X3Y8_LUT4AB/S2MID[1] Tile_X3Y8_LUT4AB/S2MID[2] Tile_X3Y8_LUT4AB/S2MID[3]
+ Tile_X3Y8_LUT4AB/S2MID[4] Tile_X3Y8_LUT4AB/S2MID[5] Tile_X3Y8_LUT4AB/S2MID[6] Tile_X3Y8_LUT4AB/S2MID[7]
+ Tile_X3Y8_LUT4AB/S2END[0] Tile_X3Y8_LUT4AB/S2END[1] Tile_X3Y8_LUT4AB/S2END[2] Tile_X3Y8_LUT4AB/S2END[3]
+ Tile_X3Y8_LUT4AB/S2END[4] Tile_X3Y8_LUT4AB/S2END[5] Tile_X3Y8_LUT4AB/S2END[6] Tile_X3Y8_LUT4AB/S2END[7]
+ Tile_X3Y7_LUT4AB/S2END[0] Tile_X3Y7_LUT4AB/S2END[1] Tile_X3Y7_LUT4AB/S2END[2] Tile_X3Y7_LUT4AB/S2END[3]
+ Tile_X3Y7_LUT4AB/S2END[4] Tile_X3Y7_LUT4AB/S2END[5] Tile_X3Y7_LUT4AB/S2END[6] Tile_X3Y7_LUT4AB/S2END[7]
+ Tile_X3Y7_LUT4AB/S2MID[0] Tile_X3Y7_LUT4AB/S2MID[1] Tile_X3Y7_LUT4AB/S2MID[2] Tile_X3Y7_LUT4AB/S2MID[3]
+ Tile_X3Y7_LUT4AB/S2MID[4] Tile_X3Y7_LUT4AB/S2MID[5] Tile_X3Y7_LUT4AB/S2MID[6] Tile_X3Y7_LUT4AB/S2MID[7]
+ Tile_X3Y8_LUT4AB/S4END[0] Tile_X3Y8_LUT4AB/S4END[10] Tile_X3Y8_LUT4AB/S4END[11]
+ Tile_X3Y8_LUT4AB/S4END[12] Tile_X3Y8_LUT4AB/S4END[13] Tile_X3Y8_LUT4AB/S4END[14]
+ Tile_X3Y8_LUT4AB/S4END[15] Tile_X3Y8_LUT4AB/S4END[1] Tile_X3Y8_LUT4AB/S4END[2] Tile_X3Y8_LUT4AB/S4END[3]
+ Tile_X3Y8_LUT4AB/S4END[4] Tile_X3Y8_LUT4AB/S4END[5] Tile_X3Y8_LUT4AB/S4END[6] Tile_X3Y8_LUT4AB/S4END[7]
+ Tile_X3Y8_LUT4AB/S4END[8] Tile_X3Y8_LUT4AB/S4END[9] Tile_X3Y7_LUT4AB/S4END[0] Tile_X3Y7_LUT4AB/S4END[10]
+ Tile_X3Y7_LUT4AB/S4END[11] Tile_X3Y7_LUT4AB/S4END[12] Tile_X3Y7_LUT4AB/S4END[13]
+ Tile_X3Y7_LUT4AB/S4END[14] Tile_X3Y7_LUT4AB/S4END[15] Tile_X3Y7_LUT4AB/S4END[1]
+ Tile_X3Y7_LUT4AB/S4END[2] Tile_X3Y7_LUT4AB/S4END[3] Tile_X3Y7_LUT4AB/S4END[4] Tile_X3Y7_LUT4AB/S4END[5]
+ Tile_X3Y7_LUT4AB/S4END[6] Tile_X3Y7_LUT4AB/S4END[7] Tile_X3Y7_LUT4AB/S4END[8] Tile_X3Y7_LUT4AB/S4END[9]
+ Tile_X3Y8_LUT4AB/SS4END[0] Tile_X3Y8_LUT4AB/SS4END[10] Tile_X3Y8_LUT4AB/SS4END[11]
+ Tile_X3Y8_LUT4AB/SS4END[12] Tile_X3Y8_LUT4AB/SS4END[13] Tile_X3Y8_LUT4AB/SS4END[14]
+ Tile_X3Y8_LUT4AB/SS4END[15] Tile_X3Y8_LUT4AB/SS4END[1] Tile_X3Y8_LUT4AB/SS4END[2]
+ Tile_X3Y8_LUT4AB/SS4END[3] Tile_X3Y8_LUT4AB/SS4END[4] Tile_X3Y8_LUT4AB/SS4END[5]
+ Tile_X3Y8_LUT4AB/SS4END[6] Tile_X3Y8_LUT4AB/SS4END[7] Tile_X3Y8_LUT4AB/SS4END[8]
+ Tile_X3Y8_LUT4AB/SS4END[9] Tile_X3Y7_LUT4AB/SS4END[0] Tile_X3Y7_LUT4AB/SS4END[10]
+ Tile_X3Y7_LUT4AB/SS4END[11] Tile_X3Y7_LUT4AB/SS4END[12] Tile_X3Y7_LUT4AB/SS4END[13]
+ Tile_X3Y7_LUT4AB/SS4END[14] Tile_X3Y7_LUT4AB/SS4END[15] Tile_X3Y7_LUT4AB/SS4END[1]
+ Tile_X3Y7_LUT4AB/SS4END[2] Tile_X3Y7_LUT4AB/SS4END[3] Tile_X3Y7_LUT4AB/SS4END[4]
+ Tile_X3Y7_LUT4AB/SS4END[5] Tile_X3Y7_LUT4AB/SS4END[6] Tile_X3Y7_LUT4AB/SS4END[7]
+ Tile_X3Y7_LUT4AB/SS4END[8] Tile_X3Y7_LUT4AB/SS4END[9] Tile_X3Y7_LUT4AB/UserCLK Tile_X3Y6_LUT4AB/UserCLK
+ VGND VPWR Tile_X3Y7_LUT4AB/W1BEG[0] Tile_X3Y7_LUT4AB/W1BEG[1] Tile_X3Y7_LUT4AB/W1BEG[2]
+ Tile_X3Y7_LUT4AB/W1BEG[3] Tile_X3Y7_LUT4AB/W1END[0] Tile_X3Y7_LUT4AB/W1END[1] Tile_X3Y7_LUT4AB/W1END[2]
+ Tile_X3Y7_LUT4AB/W1END[3] Tile_X3Y7_LUT4AB/W2BEG[0] Tile_X3Y7_LUT4AB/W2BEG[1] Tile_X3Y7_LUT4AB/W2BEG[2]
+ Tile_X3Y7_LUT4AB/W2BEG[3] Tile_X3Y7_LUT4AB/W2BEG[4] Tile_X3Y7_LUT4AB/W2BEG[5] Tile_X3Y7_LUT4AB/W2BEG[6]
+ Tile_X3Y7_LUT4AB/W2BEG[7] Tile_X2Y7_LUT4AB/W2END[0] Tile_X2Y7_LUT4AB/W2END[1] Tile_X2Y7_LUT4AB/W2END[2]
+ Tile_X2Y7_LUT4AB/W2END[3] Tile_X2Y7_LUT4AB/W2END[4] Tile_X2Y7_LUT4AB/W2END[5] Tile_X2Y7_LUT4AB/W2END[6]
+ Tile_X2Y7_LUT4AB/W2END[7] Tile_X3Y7_LUT4AB/W2END[0] Tile_X3Y7_LUT4AB/W2END[1] Tile_X3Y7_LUT4AB/W2END[2]
+ Tile_X3Y7_LUT4AB/W2END[3] Tile_X3Y7_LUT4AB/W2END[4] Tile_X3Y7_LUT4AB/W2END[5] Tile_X3Y7_LUT4AB/W2END[6]
+ Tile_X3Y7_LUT4AB/W2END[7] Tile_X3Y7_LUT4AB/W2MID[0] Tile_X3Y7_LUT4AB/W2MID[1] Tile_X3Y7_LUT4AB/W2MID[2]
+ Tile_X3Y7_LUT4AB/W2MID[3] Tile_X3Y7_LUT4AB/W2MID[4] Tile_X3Y7_LUT4AB/W2MID[5] Tile_X3Y7_LUT4AB/W2MID[6]
+ Tile_X3Y7_LUT4AB/W2MID[7] Tile_X3Y7_LUT4AB/W6BEG[0] Tile_X3Y7_LUT4AB/W6BEG[10] Tile_X3Y7_LUT4AB/W6BEG[11]
+ Tile_X3Y7_LUT4AB/W6BEG[1] Tile_X3Y7_LUT4AB/W6BEG[2] Tile_X3Y7_LUT4AB/W6BEG[3] Tile_X3Y7_LUT4AB/W6BEG[4]
+ Tile_X3Y7_LUT4AB/W6BEG[5] Tile_X3Y7_LUT4AB/W6BEG[6] Tile_X3Y7_LUT4AB/W6BEG[7] Tile_X3Y7_LUT4AB/W6BEG[8]
+ Tile_X3Y7_LUT4AB/W6BEG[9] Tile_X3Y7_LUT4AB/W6END[0] Tile_X3Y7_LUT4AB/W6END[10] Tile_X3Y7_LUT4AB/W6END[11]
+ Tile_X3Y7_LUT4AB/W6END[1] Tile_X3Y7_LUT4AB/W6END[2] Tile_X3Y7_LUT4AB/W6END[3] Tile_X3Y7_LUT4AB/W6END[4]
+ Tile_X3Y7_LUT4AB/W6END[5] Tile_X3Y7_LUT4AB/W6END[6] Tile_X3Y7_LUT4AB/W6END[7] Tile_X3Y7_LUT4AB/W6END[8]
+ Tile_X3Y7_LUT4AB/W6END[9] Tile_X3Y7_LUT4AB/WW4BEG[0] Tile_X3Y7_LUT4AB/WW4BEG[10]
+ Tile_X3Y7_LUT4AB/WW4BEG[11] Tile_X3Y7_LUT4AB/WW4BEG[12] Tile_X3Y7_LUT4AB/WW4BEG[13]
+ Tile_X3Y7_LUT4AB/WW4BEG[14] Tile_X3Y7_LUT4AB/WW4BEG[15] Tile_X3Y7_LUT4AB/WW4BEG[1]
+ Tile_X3Y7_LUT4AB/WW4BEG[2] Tile_X3Y7_LUT4AB/WW4BEG[3] Tile_X3Y7_LUT4AB/WW4BEG[4]
+ Tile_X3Y7_LUT4AB/WW4BEG[5] Tile_X3Y7_LUT4AB/WW4BEG[6] Tile_X3Y7_LUT4AB/WW4BEG[7]
+ Tile_X3Y7_LUT4AB/WW4BEG[8] Tile_X3Y7_LUT4AB/WW4BEG[9] Tile_X3Y7_LUT4AB/WW4END[0]
+ Tile_X3Y7_LUT4AB/WW4END[10] Tile_X3Y7_LUT4AB/WW4END[11] Tile_X3Y7_LUT4AB/WW4END[12]
+ Tile_X3Y7_LUT4AB/WW4END[13] Tile_X3Y7_LUT4AB/WW4END[14] Tile_X3Y7_LUT4AB/WW4END[15]
+ Tile_X3Y7_LUT4AB/WW4END[1] Tile_X3Y7_LUT4AB/WW4END[2] Tile_X3Y7_LUT4AB/WW4END[3]
+ Tile_X3Y7_LUT4AB/WW4END[4] Tile_X3Y7_LUT4AB/WW4END[5] Tile_X3Y7_LUT4AB/WW4END[6]
+ Tile_X3Y7_LUT4AB/WW4END[7] Tile_X3Y7_LUT4AB/WW4END[8] Tile_X3Y7_LUT4AB/WW4END[9]
+ LUT4AB
XTile_X0Y7_W_IO Tile_X0Y7_A_I_top Tile_X0Y7_A_O_top Tile_X0Y7_A_T_top Tile_X0Y7_A_config_C_bit0
+ Tile_X0Y7_A_config_C_bit1 Tile_X0Y7_A_config_C_bit2 Tile_X0Y7_A_config_C_bit3 Tile_X0Y7_B_I_top
+ Tile_X0Y7_B_O_top Tile_X0Y7_B_T_top Tile_X0Y7_B_config_C_bit0 Tile_X0Y7_B_config_C_bit1
+ Tile_X0Y7_B_config_C_bit2 Tile_X0Y7_B_config_C_bit3 Tile_X0Y7_W_IO/E1BEG[0] Tile_X0Y7_W_IO/E1BEG[1]
+ Tile_X0Y7_W_IO/E1BEG[2] Tile_X0Y7_W_IO/E1BEG[3] Tile_X0Y7_W_IO/E2BEG[0] Tile_X0Y7_W_IO/E2BEG[1]
+ Tile_X0Y7_W_IO/E2BEG[2] Tile_X0Y7_W_IO/E2BEG[3] Tile_X0Y7_W_IO/E2BEG[4] Tile_X0Y7_W_IO/E2BEG[5]
+ Tile_X0Y7_W_IO/E2BEG[6] Tile_X0Y7_W_IO/E2BEG[7] Tile_X0Y7_W_IO/E2BEGb[0] Tile_X0Y7_W_IO/E2BEGb[1]
+ Tile_X0Y7_W_IO/E2BEGb[2] Tile_X0Y7_W_IO/E2BEGb[3] Tile_X0Y7_W_IO/E2BEGb[4] Tile_X0Y7_W_IO/E2BEGb[5]
+ Tile_X0Y7_W_IO/E2BEGb[6] Tile_X0Y7_W_IO/E2BEGb[7] Tile_X0Y7_W_IO/E6BEG[0] Tile_X0Y7_W_IO/E6BEG[10]
+ Tile_X0Y7_W_IO/E6BEG[11] Tile_X0Y7_W_IO/E6BEG[1] Tile_X0Y7_W_IO/E6BEG[2] Tile_X0Y7_W_IO/E6BEG[3]
+ Tile_X0Y7_W_IO/E6BEG[4] Tile_X0Y7_W_IO/E6BEG[5] Tile_X0Y7_W_IO/E6BEG[6] Tile_X0Y7_W_IO/E6BEG[7]
+ Tile_X0Y7_W_IO/E6BEG[8] Tile_X0Y7_W_IO/E6BEG[9] Tile_X0Y7_W_IO/EE4BEG[0] Tile_X0Y7_W_IO/EE4BEG[10]
+ Tile_X0Y7_W_IO/EE4BEG[11] Tile_X0Y7_W_IO/EE4BEG[12] Tile_X0Y7_W_IO/EE4BEG[13] Tile_X0Y7_W_IO/EE4BEG[14]
+ Tile_X0Y7_W_IO/EE4BEG[15] Tile_X0Y7_W_IO/EE4BEG[1] Tile_X0Y7_W_IO/EE4BEG[2] Tile_X0Y7_W_IO/EE4BEG[3]
+ Tile_X0Y7_W_IO/EE4BEG[4] Tile_X0Y7_W_IO/EE4BEG[5] Tile_X0Y7_W_IO/EE4BEG[6] Tile_X0Y7_W_IO/EE4BEG[7]
+ Tile_X0Y7_W_IO/EE4BEG[8] Tile_X0Y7_W_IO/EE4BEG[9] FrameData[224] FrameData[234]
+ FrameData[235] FrameData[236] FrameData[237] FrameData[238] FrameData[239] FrameData[240]
+ FrameData[241] FrameData[242] FrameData[243] FrameData[225] FrameData[244] FrameData[245]
+ FrameData[246] FrameData[247] FrameData[248] FrameData[249] FrameData[250] FrameData[251]
+ FrameData[252] FrameData[253] FrameData[226] FrameData[254] FrameData[255] FrameData[227]
+ FrameData[228] FrameData[229] FrameData[230] FrameData[231] FrameData[232] FrameData[233]
+ Tile_X1Y7_LUT4AB/FrameData[0] Tile_X1Y7_LUT4AB/FrameData[10] Tile_X1Y7_LUT4AB/FrameData[11]
+ Tile_X1Y7_LUT4AB/FrameData[12] Tile_X1Y7_LUT4AB/FrameData[13] Tile_X1Y7_LUT4AB/FrameData[14]
+ Tile_X1Y7_LUT4AB/FrameData[15] Tile_X1Y7_LUT4AB/FrameData[16] Tile_X1Y7_LUT4AB/FrameData[17]
+ Tile_X1Y7_LUT4AB/FrameData[18] Tile_X1Y7_LUT4AB/FrameData[19] Tile_X1Y7_LUT4AB/FrameData[1]
+ Tile_X1Y7_LUT4AB/FrameData[20] Tile_X1Y7_LUT4AB/FrameData[21] Tile_X1Y7_LUT4AB/FrameData[22]
+ Tile_X1Y7_LUT4AB/FrameData[23] Tile_X1Y7_LUT4AB/FrameData[24] Tile_X1Y7_LUT4AB/FrameData[25]
+ Tile_X1Y7_LUT4AB/FrameData[26] Tile_X1Y7_LUT4AB/FrameData[27] Tile_X1Y7_LUT4AB/FrameData[28]
+ Tile_X1Y7_LUT4AB/FrameData[29] Tile_X1Y7_LUT4AB/FrameData[2] Tile_X1Y7_LUT4AB/FrameData[30]
+ Tile_X1Y7_LUT4AB/FrameData[31] Tile_X1Y7_LUT4AB/FrameData[3] Tile_X1Y7_LUT4AB/FrameData[4]
+ Tile_X1Y7_LUT4AB/FrameData[5] Tile_X1Y7_LUT4AB/FrameData[6] Tile_X1Y7_LUT4AB/FrameData[7]
+ Tile_X1Y7_LUT4AB/FrameData[8] Tile_X1Y7_LUT4AB/FrameData[9] Tile_X0Y7_W_IO/FrameStrobe[0]
+ Tile_X0Y7_W_IO/FrameStrobe[10] Tile_X0Y7_W_IO/FrameStrobe[11] Tile_X0Y7_W_IO/FrameStrobe[12]
+ Tile_X0Y7_W_IO/FrameStrobe[13] Tile_X0Y7_W_IO/FrameStrobe[14] Tile_X0Y7_W_IO/FrameStrobe[15]
+ Tile_X0Y7_W_IO/FrameStrobe[16] Tile_X0Y7_W_IO/FrameStrobe[17] Tile_X0Y7_W_IO/FrameStrobe[18]
+ Tile_X0Y7_W_IO/FrameStrobe[19] Tile_X0Y7_W_IO/FrameStrobe[1] Tile_X0Y7_W_IO/FrameStrobe[2]
+ Tile_X0Y7_W_IO/FrameStrobe[3] Tile_X0Y7_W_IO/FrameStrobe[4] Tile_X0Y7_W_IO/FrameStrobe[5]
+ Tile_X0Y7_W_IO/FrameStrobe[6] Tile_X0Y7_W_IO/FrameStrobe[7] Tile_X0Y7_W_IO/FrameStrobe[8]
+ Tile_X0Y7_W_IO/FrameStrobe[9] Tile_X0Y6_W_IO/FrameStrobe[0] Tile_X0Y6_W_IO/FrameStrobe[10]
+ Tile_X0Y6_W_IO/FrameStrobe[11] Tile_X0Y6_W_IO/FrameStrobe[12] Tile_X0Y6_W_IO/FrameStrobe[13]
+ Tile_X0Y6_W_IO/FrameStrobe[14] Tile_X0Y6_W_IO/FrameStrobe[15] Tile_X0Y6_W_IO/FrameStrobe[16]
+ Tile_X0Y6_W_IO/FrameStrobe[17] Tile_X0Y6_W_IO/FrameStrobe[18] Tile_X0Y6_W_IO/FrameStrobe[19]
+ Tile_X0Y6_W_IO/FrameStrobe[1] Tile_X0Y6_W_IO/FrameStrobe[2] Tile_X0Y6_W_IO/FrameStrobe[3]
+ Tile_X0Y6_W_IO/FrameStrobe[4] Tile_X0Y6_W_IO/FrameStrobe[5] Tile_X0Y6_W_IO/FrameStrobe[6]
+ Tile_X0Y6_W_IO/FrameStrobe[7] Tile_X0Y6_W_IO/FrameStrobe[8] Tile_X0Y6_W_IO/FrameStrobe[9]
+ Tile_X0Y7_W_IO/UserCLK Tile_X0Y6_W_IO/UserCLK VGND VPWR Tile_X0Y7_W_IO/W1END[0]
+ Tile_X0Y7_W_IO/W1END[1] Tile_X0Y7_W_IO/W1END[2] Tile_X0Y7_W_IO/W1END[3] Tile_X0Y7_W_IO/W2END[0]
+ Tile_X0Y7_W_IO/W2END[1] Tile_X0Y7_W_IO/W2END[2] Tile_X0Y7_W_IO/W2END[3] Tile_X0Y7_W_IO/W2END[4]
+ Tile_X0Y7_W_IO/W2END[5] Tile_X0Y7_W_IO/W2END[6] Tile_X0Y7_W_IO/W2END[7] Tile_X0Y7_W_IO/W2MID[0]
+ Tile_X0Y7_W_IO/W2MID[1] Tile_X0Y7_W_IO/W2MID[2] Tile_X0Y7_W_IO/W2MID[3] Tile_X0Y7_W_IO/W2MID[4]
+ Tile_X0Y7_W_IO/W2MID[5] Tile_X0Y7_W_IO/W2MID[6] Tile_X0Y7_W_IO/W2MID[7] Tile_X0Y7_W_IO/W6END[0]
+ Tile_X0Y7_W_IO/W6END[10] Tile_X0Y7_W_IO/W6END[11] Tile_X0Y7_W_IO/W6END[1] Tile_X0Y7_W_IO/W6END[2]
+ Tile_X0Y7_W_IO/W6END[3] Tile_X0Y7_W_IO/W6END[4] Tile_X0Y7_W_IO/W6END[5] Tile_X0Y7_W_IO/W6END[6]
+ Tile_X0Y7_W_IO/W6END[7] Tile_X0Y7_W_IO/W6END[8] Tile_X0Y7_W_IO/W6END[9] Tile_X0Y7_W_IO/WW4END[0]
+ Tile_X0Y7_W_IO/WW4END[10] Tile_X0Y7_W_IO/WW4END[11] Tile_X0Y7_W_IO/WW4END[12] Tile_X0Y7_W_IO/WW4END[13]
+ Tile_X0Y7_W_IO/WW4END[14] Tile_X0Y7_W_IO/WW4END[15] Tile_X0Y7_W_IO/WW4END[1] Tile_X0Y7_W_IO/WW4END[2]
+ Tile_X0Y7_W_IO/WW4END[3] Tile_X0Y7_W_IO/WW4END[4] Tile_X0Y7_W_IO/WW4END[5] Tile_X0Y7_W_IO/WW4END[6]
+ Tile_X0Y7_W_IO/WW4END[7] Tile_X0Y7_W_IO/WW4END[8] Tile_X0Y7_W_IO/WW4END[9] W_IO
XTile_X9Y15_S_CPU_IF Tile_X9Y14_LUT4AB/Ci Tile_X9Y15_S_CPU_IF/FrameData[0] Tile_X9Y15_S_CPU_IF/FrameData[10]
+ Tile_X9Y15_S_CPU_IF/FrameData[11] Tile_X9Y15_S_CPU_IF/FrameData[12] Tile_X9Y15_S_CPU_IF/FrameData[13]
+ Tile_X9Y15_S_CPU_IF/FrameData[14] Tile_X9Y15_S_CPU_IF/FrameData[15] Tile_X9Y15_S_CPU_IF/FrameData[16]
+ Tile_X9Y15_S_CPU_IF/FrameData[17] Tile_X9Y15_S_CPU_IF/FrameData[18] Tile_X9Y15_S_CPU_IF/FrameData[19]
+ Tile_X9Y15_S_CPU_IF/FrameData[1] Tile_X9Y15_S_CPU_IF/FrameData[20] Tile_X9Y15_S_CPU_IF/FrameData[21]
+ Tile_X9Y15_S_CPU_IF/FrameData[22] Tile_X9Y15_S_CPU_IF/FrameData[23] Tile_X9Y15_S_CPU_IF/FrameData[24]
+ Tile_X9Y15_S_CPU_IF/FrameData[25] Tile_X9Y15_S_CPU_IF/FrameData[26] Tile_X9Y15_S_CPU_IF/FrameData[27]
+ Tile_X9Y15_S_CPU_IF/FrameData[28] Tile_X9Y15_S_CPU_IF/FrameData[29] Tile_X9Y15_S_CPU_IF/FrameData[2]
+ Tile_X9Y15_S_CPU_IF/FrameData[30] Tile_X9Y15_S_CPU_IF/FrameData[31] Tile_X9Y15_S_CPU_IF/FrameData[3]
+ Tile_X9Y15_S_CPU_IF/FrameData[4] Tile_X9Y15_S_CPU_IF/FrameData[5] Tile_X9Y15_S_CPU_IF/FrameData[6]
+ Tile_X9Y15_S_CPU_IF/FrameData[7] Tile_X9Y15_S_CPU_IF/FrameData[8] Tile_X9Y15_S_CPU_IF/FrameData[9]
+ Tile_X9Y15_S_CPU_IF/FrameData_O[0] Tile_X9Y15_S_CPU_IF/FrameData_O[10] Tile_X9Y15_S_CPU_IF/FrameData_O[11]
+ Tile_X9Y15_S_CPU_IF/FrameData_O[12] Tile_X9Y15_S_CPU_IF/FrameData_O[13] Tile_X9Y15_S_CPU_IF/FrameData_O[14]
+ Tile_X9Y15_S_CPU_IF/FrameData_O[15] Tile_X9Y15_S_CPU_IF/FrameData_O[16] Tile_X9Y15_S_CPU_IF/FrameData_O[17]
+ Tile_X9Y15_S_CPU_IF/FrameData_O[18] Tile_X9Y15_S_CPU_IF/FrameData_O[19] Tile_X9Y15_S_CPU_IF/FrameData_O[1]
+ Tile_X9Y15_S_CPU_IF/FrameData_O[20] Tile_X9Y15_S_CPU_IF/FrameData_O[21] Tile_X9Y15_S_CPU_IF/FrameData_O[22]
+ Tile_X9Y15_S_CPU_IF/FrameData_O[23] Tile_X9Y15_S_CPU_IF/FrameData_O[24] Tile_X9Y15_S_CPU_IF/FrameData_O[25]
+ Tile_X9Y15_S_CPU_IF/FrameData_O[26] Tile_X9Y15_S_CPU_IF/FrameData_O[27] Tile_X9Y15_S_CPU_IF/FrameData_O[28]
+ Tile_X9Y15_S_CPU_IF/FrameData_O[29] Tile_X9Y15_S_CPU_IF/FrameData_O[2] Tile_X9Y15_S_CPU_IF/FrameData_O[30]
+ Tile_X9Y15_S_CPU_IF/FrameData_O[31] Tile_X9Y15_S_CPU_IF/FrameData_O[3] Tile_X9Y15_S_CPU_IF/FrameData_O[4]
+ Tile_X9Y15_S_CPU_IF/FrameData_O[5] Tile_X9Y15_S_CPU_IF/FrameData_O[6] Tile_X9Y15_S_CPU_IF/FrameData_O[7]
+ Tile_X9Y15_S_CPU_IF/FrameData_O[8] Tile_X9Y15_S_CPU_IF/FrameData_O[9] FrameStrobe[180]
+ FrameStrobe[190] FrameStrobe[191] FrameStrobe[192] FrameStrobe[193] FrameStrobe[194]
+ FrameStrobe[195] FrameStrobe[196] FrameStrobe[197] FrameStrobe[198] FrameStrobe[199]
+ FrameStrobe[181] FrameStrobe[182] FrameStrobe[183] FrameStrobe[184] FrameStrobe[185]
+ FrameStrobe[186] FrameStrobe[187] FrameStrobe[188] FrameStrobe[189] Tile_X9Y14_LUT4AB/FrameStrobe[0]
+ Tile_X9Y14_LUT4AB/FrameStrobe[10] Tile_X9Y14_LUT4AB/FrameStrobe[11] Tile_X9Y14_LUT4AB/FrameStrobe[12]
+ Tile_X9Y14_LUT4AB/FrameStrobe[13] Tile_X9Y14_LUT4AB/FrameStrobe[14] Tile_X9Y14_LUT4AB/FrameStrobe[15]
+ Tile_X9Y14_LUT4AB/FrameStrobe[16] Tile_X9Y14_LUT4AB/FrameStrobe[17] Tile_X9Y14_LUT4AB/FrameStrobe[18]
+ Tile_X9Y14_LUT4AB/FrameStrobe[19] Tile_X9Y14_LUT4AB/FrameStrobe[1] Tile_X9Y14_LUT4AB/FrameStrobe[2]
+ Tile_X9Y14_LUT4AB/FrameStrobe[3] Tile_X9Y14_LUT4AB/FrameStrobe[4] Tile_X9Y14_LUT4AB/FrameStrobe[5]
+ Tile_X9Y14_LUT4AB/FrameStrobe[6] Tile_X9Y14_LUT4AB/FrameStrobe[7] Tile_X9Y14_LUT4AB/FrameStrobe[8]
+ Tile_X9Y14_LUT4AB/FrameStrobe[9] Tile_X9Y15_I_top0 Tile_X9Y15_I_top1 Tile_X9Y15_I_top10
+ Tile_X9Y15_I_top11 Tile_X9Y15_I_top12 Tile_X9Y15_I_top13 Tile_X9Y15_I_top14 Tile_X9Y15_I_top15
+ Tile_X9Y15_I_top2 Tile_X9Y15_I_top3 Tile_X9Y15_I_top4 Tile_X9Y15_I_top5 Tile_X9Y15_I_top6
+ Tile_X9Y15_I_top7 Tile_X9Y15_I_top8 Tile_X9Y15_I_top9 Tile_X9Y14_LUT4AB/N1END[0]
+ Tile_X9Y14_LUT4AB/N1END[1] Tile_X9Y14_LUT4AB/N1END[2] Tile_X9Y14_LUT4AB/N1END[3]
+ Tile_X9Y14_LUT4AB/N2MID[0] Tile_X9Y14_LUT4AB/N2MID[1] Tile_X9Y14_LUT4AB/N2MID[2]
+ Tile_X9Y14_LUT4AB/N2MID[3] Tile_X9Y14_LUT4AB/N2MID[4] Tile_X9Y14_LUT4AB/N2MID[5]
+ Tile_X9Y14_LUT4AB/N2MID[6] Tile_X9Y14_LUT4AB/N2MID[7] Tile_X9Y14_LUT4AB/N2END[0]
+ Tile_X9Y14_LUT4AB/N2END[1] Tile_X9Y14_LUT4AB/N2END[2] Tile_X9Y14_LUT4AB/N2END[3]
+ Tile_X9Y14_LUT4AB/N2END[4] Tile_X9Y14_LUT4AB/N2END[5] Tile_X9Y14_LUT4AB/N2END[6]
+ Tile_X9Y14_LUT4AB/N2END[7] Tile_X9Y14_LUT4AB/N4END[0] Tile_X9Y14_LUT4AB/N4END[10]
+ Tile_X9Y14_LUT4AB/N4END[11] Tile_X9Y14_LUT4AB/N4END[12] Tile_X9Y14_LUT4AB/N4END[13]
+ Tile_X9Y14_LUT4AB/N4END[14] Tile_X9Y14_LUT4AB/N4END[15] Tile_X9Y14_LUT4AB/N4END[1]
+ Tile_X9Y14_LUT4AB/N4END[2] Tile_X9Y14_LUT4AB/N4END[3] Tile_X9Y14_LUT4AB/N4END[4]
+ Tile_X9Y14_LUT4AB/N4END[5] Tile_X9Y14_LUT4AB/N4END[6] Tile_X9Y14_LUT4AB/N4END[7]
+ Tile_X9Y14_LUT4AB/N4END[8] Tile_X9Y14_LUT4AB/N4END[9] Tile_X9Y14_LUT4AB/NN4END[0]
+ Tile_X9Y14_LUT4AB/NN4END[10] Tile_X9Y14_LUT4AB/NN4END[11] Tile_X9Y14_LUT4AB/NN4END[12]
+ Tile_X9Y14_LUT4AB/NN4END[13] Tile_X9Y14_LUT4AB/NN4END[14] Tile_X9Y14_LUT4AB/NN4END[15]
+ Tile_X9Y14_LUT4AB/NN4END[1] Tile_X9Y14_LUT4AB/NN4END[2] Tile_X9Y14_LUT4AB/NN4END[3]
+ Tile_X9Y14_LUT4AB/NN4END[4] Tile_X9Y14_LUT4AB/NN4END[5] Tile_X9Y14_LUT4AB/NN4END[6]
+ Tile_X9Y14_LUT4AB/NN4END[7] Tile_X9Y14_LUT4AB/NN4END[8] Tile_X9Y14_LUT4AB/NN4END[9]
+ Tile_X9Y15_O_top0 Tile_X9Y15_O_top1 Tile_X9Y15_O_top10 Tile_X9Y15_O_top11 Tile_X9Y15_O_top12
+ Tile_X9Y15_O_top13 Tile_X9Y15_O_top14 Tile_X9Y15_O_top15 Tile_X9Y15_O_top2 Tile_X9Y15_O_top3
+ Tile_X9Y15_O_top4 Tile_X9Y15_O_top5 Tile_X9Y15_O_top6 Tile_X9Y15_O_top7 Tile_X9Y15_O_top8
+ Tile_X9Y15_O_top9 Tile_X9Y14_LUT4AB/S1BEG[0] Tile_X9Y14_LUT4AB/S1BEG[1] Tile_X9Y14_LUT4AB/S1BEG[2]
+ Tile_X9Y14_LUT4AB/S1BEG[3] Tile_X9Y14_LUT4AB/S2BEGb[0] Tile_X9Y14_LUT4AB/S2BEGb[1]
+ Tile_X9Y14_LUT4AB/S2BEGb[2] Tile_X9Y14_LUT4AB/S2BEGb[3] Tile_X9Y14_LUT4AB/S2BEGb[4]
+ Tile_X9Y14_LUT4AB/S2BEGb[5] Tile_X9Y14_LUT4AB/S2BEGb[6] Tile_X9Y14_LUT4AB/S2BEGb[7]
+ Tile_X9Y14_LUT4AB/S2BEG[0] Tile_X9Y14_LUT4AB/S2BEG[1] Tile_X9Y14_LUT4AB/S2BEG[2]
+ Tile_X9Y14_LUT4AB/S2BEG[3] Tile_X9Y14_LUT4AB/S2BEG[4] Tile_X9Y14_LUT4AB/S2BEG[5]
+ Tile_X9Y14_LUT4AB/S2BEG[6] Tile_X9Y14_LUT4AB/S2BEG[7] Tile_X9Y14_LUT4AB/S4BEG[0]
+ Tile_X9Y14_LUT4AB/S4BEG[10] Tile_X9Y14_LUT4AB/S4BEG[11] Tile_X9Y14_LUT4AB/S4BEG[12]
+ Tile_X9Y14_LUT4AB/S4BEG[13] Tile_X9Y14_LUT4AB/S4BEG[14] Tile_X9Y14_LUT4AB/S4BEG[15]
+ Tile_X9Y14_LUT4AB/S4BEG[1] Tile_X9Y14_LUT4AB/S4BEG[2] Tile_X9Y14_LUT4AB/S4BEG[3]
+ Tile_X9Y14_LUT4AB/S4BEG[4] Tile_X9Y14_LUT4AB/S4BEG[5] Tile_X9Y14_LUT4AB/S4BEG[6]
+ Tile_X9Y14_LUT4AB/S4BEG[7] Tile_X9Y14_LUT4AB/S4BEG[8] Tile_X9Y14_LUT4AB/S4BEG[9]
+ Tile_X9Y14_LUT4AB/SS4BEG[0] Tile_X9Y14_LUT4AB/SS4BEG[10] Tile_X9Y14_LUT4AB/SS4BEG[11]
+ Tile_X9Y14_LUT4AB/SS4BEG[12] Tile_X9Y14_LUT4AB/SS4BEG[13] Tile_X9Y14_LUT4AB/SS4BEG[14]
+ Tile_X9Y14_LUT4AB/SS4BEG[15] Tile_X9Y14_LUT4AB/SS4BEG[1] Tile_X9Y14_LUT4AB/SS4BEG[2]
+ Tile_X9Y14_LUT4AB/SS4BEG[3] Tile_X9Y14_LUT4AB/SS4BEG[4] Tile_X9Y14_LUT4AB/SS4BEG[5]
+ Tile_X9Y14_LUT4AB/SS4BEG[6] Tile_X9Y14_LUT4AB/SS4BEG[7] Tile_X9Y14_LUT4AB/SS4BEG[8]
+ Tile_X9Y14_LUT4AB/SS4BEG[9] UserCLK Tile_X9Y14_LUT4AB/UserCLK VGND VPWR S_CPU_IF
XTile_X4Y8_RegFile Tile_X5Y8_LUT4AB/E1END[0] Tile_X5Y8_LUT4AB/E1END[1] Tile_X5Y8_LUT4AB/E1END[2]
+ Tile_X5Y8_LUT4AB/E1END[3] Tile_X3Y8_LUT4AB/E1BEG[0] Tile_X3Y8_LUT4AB/E1BEG[1] Tile_X3Y8_LUT4AB/E1BEG[2]
+ Tile_X3Y8_LUT4AB/E1BEG[3] Tile_X5Y8_LUT4AB/E2MID[0] Tile_X5Y8_LUT4AB/E2MID[1] Tile_X5Y8_LUT4AB/E2MID[2]
+ Tile_X5Y8_LUT4AB/E2MID[3] Tile_X5Y8_LUT4AB/E2MID[4] Tile_X5Y8_LUT4AB/E2MID[5] Tile_X5Y8_LUT4AB/E2MID[6]
+ Tile_X5Y8_LUT4AB/E2MID[7] Tile_X5Y8_LUT4AB/E2END[0] Tile_X5Y8_LUT4AB/E2END[1] Tile_X5Y8_LUT4AB/E2END[2]
+ Tile_X5Y8_LUT4AB/E2END[3] Tile_X5Y8_LUT4AB/E2END[4] Tile_X5Y8_LUT4AB/E2END[5] Tile_X5Y8_LUT4AB/E2END[6]
+ Tile_X5Y8_LUT4AB/E2END[7] Tile_X4Y8_RegFile/E2END[0] Tile_X4Y8_RegFile/E2END[1]
+ Tile_X4Y8_RegFile/E2END[2] Tile_X4Y8_RegFile/E2END[3] Tile_X4Y8_RegFile/E2END[4]
+ Tile_X4Y8_RegFile/E2END[5] Tile_X4Y8_RegFile/E2END[6] Tile_X4Y8_RegFile/E2END[7]
+ Tile_X3Y8_LUT4AB/E2BEG[0] Tile_X3Y8_LUT4AB/E2BEG[1] Tile_X3Y8_LUT4AB/E2BEG[2] Tile_X3Y8_LUT4AB/E2BEG[3]
+ Tile_X3Y8_LUT4AB/E2BEG[4] Tile_X3Y8_LUT4AB/E2BEG[5] Tile_X3Y8_LUT4AB/E2BEG[6] Tile_X3Y8_LUT4AB/E2BEG[7]
+ Tile_X5Y8_LUT4AB/E6END[0] Tile_X5Y8_LUT4AB/E6END[10] Tile_X5Y8_LUT4AB/E6END[11]
+ Tile_X5Y8_LUT4AB/E6END[1] Tile_X5Y8_LUT4AB/E6END[2] Tile_X5Y8_LUT4AB/E6END[3] Tile_X5Y8_LUT4AB/E6END[4]
+ Tile_X5Y8_LUT4AB/E6END[5] Tile_X5Y8_LUT4AB/E6END[6] Tile_X5Y8_LUT4AB/E6END[7] Tile_X5Y8_LUT4AB/E6END[8]
+ Tile_X5Y8_LUT4AB/E6END[9] Tile_X3Y8_LUT4AB/E6BEG[0] Tile_X3Y8_LUT4AB/E6BEG[10] Tile_X3Y8_LUT4AB/E6BEG[11]
+ Tile_X3Y8_LUT4AB/E6BEG[1] Tile_X3Y8_LUT4AB/E6BEG[2] Tile_X3Y8_LUT4AB/E6BEG[3] Tile_X3Y8_LUT4AB/E6BEG[4]
+ Tile_X3Y8_LUT4AB/E6BEG[5] Tile_X3Y8_LUT4AB/E6BEG[6] Tile_X3Y8_LUT4AB/E6BEG[7] Tile_X3Y8_LUT4AB/E6BEG[8]
+ Tile_X3Y8_LUT4AB/E6BEG[9] Tile_X5Y8_LUT4AB/EE4END[0] Tile_X5Y8_LUT4AB/EE4END[10]
+ Tile_X5Y8_LUT4AB/EE4END[11] Tile_X5Y8_LUT4AB/EE4END[12] Tile_X5Y8_LUT4AB/EE4END[13]
+ Tile_X5Y8_LUT4AB/EE4END[14] Tile_X5Y8_LUT4AB/EE4END[15] Tile_X5Y8_LUT4AB/EE4END[1]
+ Tile_X5Y8_LUT4AB/EE4END[2] Tile_X5Y8_LUT4AB/EE4END[3] Tile_X5Y8_LUT4AB/EE4END[4]
+ Tile_X5Y8_LUT4AB/EE4END[5] Tile_X5Y8_LUT4AB/EE4END[6] Tile_X5Y8_LUT4AB/EE4END[7]
+ Tile_X5Y8_LUT4AB/EE4END[8] Tile_X5Y8_LUT4AB/EE4END[9] Tile_X3Y8_LUT4AB/EE4BEG[0]
+ Tile_X3Y8_LUT4AB/EE4BEG[10] Tile_X3Y8_LUT4AB/EE4BEG[11] Tile_X3Y8_LUT4AB/EE4BEG[12]
+ Tile_X3Y8_LUT4AB/EE4BEG[13] Tile_X3Y8_LUT4AB/EE4BEG[14] Tile_X3Y8_LUT4AB/EE4BEG[15]
+ Tile_X3Y8_LUT4AB/EE4BEG[1] Tile_X3Y8_LUT4AB/EE4BEG[2] Tile_X3Y8_LUT4AB/EE4BEG[3]
+ Tile_X3Y8_LUT4AB/EE4BEG[4] Tile_X3Y8_LUT4AB/EE4BEG[5] Tile_X3Y8_LUT4AB/EE4BEG[6]
+ Tile_X3Y8_LUT4AB/EE4BEG[7] Tile_X3Y8_LUT4AB/EE4BEG[8] Tile_X3Y8_LUT4AB/EE4BEG[9]
+ Tile_X4Y8_RegFile/FrameData[0] Tile_X4Y8_RegFile/FrameData[10] Tile_X4Y8_RegFile/FrameData[11]
+ Tile_X4Y8_RegFile/FrameData[12] Tile_X4Y8_RegFile/FrameData[13] Tile_X4Y8_RegFile/FrameData[14]
+ Tile_X4Y8_RegFile/FrameData[15] Tile_X4Y8_RegFile/FrameData[16] Tile_X4Y8_RegFile/FrameData[17]
+ Tile_X4Y8_RegFile/FrameData[18] Tile_X4Y8_RegFile/FrameData[19] Tile_X4Y8_RegFile/FrameData[1]
+ Tile_X4Y8_RegFile/FrameData[20] Tile_X4Y8_RegFile/FrameData[21] Tile_X4Y8_RegFile/FrameData[22]
+ Tile_X4Y8_RegFile/FrameData[23] Tile_X4Y8_RegFile/FrameData[24] Tile_X4Y8_RegFile/FrameData[25]
+ Tile_X4Y8_RegFile/FrameData[26] Tile_X4Y8_RegFile/FrameData[27] Tile_X4Y8_RegFile/FrameData[28]
+ Tile_X4Y8_RegFile/FrameData[29] Tile_X4Y8_RegFile/FrameData[2] Tile_X4Y8_RegFile/FrameData[30]
+ Tile_X4Y8_RegFile/FrameData[31] Tile_X4Y8_RegFile/FrameData[3] Tile_X4Y8_RegFile/FrameData[4]
+ Tile_X4Y8_RegFile/FrameData[5] Tile_X4Y8_RegFile/FrameData[6] Tile_X4Y8_RegFile/FrameData[7]
+ Tile_X4Y8_RegFile/FrameData[8] Tile_X4Y8_RegFile/FrameData[9] Tile_X5Y8_LUT4AB/FrameData[0]
+ Tile_X5Y8_LUT4AB/FrameData[10] Tile_X5Y8_LUT4AB/FrameData[11] Tile_X5Y8_LUT4AB/FrameData[12]
+ Tile_X5Y8_LUT4AB/FrameData[13] Tile_X5Y8_LUT4AB/FrameData[14] Tile_X5Y8_LUT4AB/FrameData[15]
+ Tile_X5Y8_LUT4AB/FrameData[16] Tile_X5Y8_LUT4AB/FrameData[17] Tile_X5Y8_LUT4AB/FrameData[18]
+ Tile_X5Y8_LUT4AB/FrameData[19] Tile_X5Y8_LUT4AB/FrameData[1] Tile_X5Y8_LUT4AB/FrameData[20]
+ Tile_X5Y8_LUT4AB/FrameData[21] Tile_X5Y8_LUT4AB/FrameData[22] Tile_X5Y8_LUT4AB/FrameData[23]
+ Tile_X5Y8_LUT4AB/FrameData[24] Tile_X5Y8_LUT4AB/FrameData[25] Tile_X5Y8_LUT4AB/FrameData[26]
+ Tile_X5Y8_LUT4AB/FrameData[27] Tile_X5Y8_LUT4AB/FrameData[28] Tile_X5Y8_LUT4AB/FrameData[29]
+ Tile_X5Y8_LUT4AB/FrameData[2] Tile_X5Y8_LUT4AB/FrameData[30] Tile_X5Y8_LUT4AB/FrameData[31]
+ Tile_X5Y8_LUT4AB/FrameData[3] Tile_X5Y8_LUT4AB/FrameData[4] Tile_X5Y8_LUT4AB/FrameData[5]
+ Tile_X5Y8_LUT4AB/FrameData[6] Tile_X5Y8_LUT4AB/FrameData[7] Tile_X5Y8_LUT4AB/FrameData[8]
+ Tile_X5Y8_LUT4AB/FrameData[9] Tile_X4Y8_RegFile/FrameStrobe[0] Tile_X4Y8_RegFile/FrameStrobe[10]
+ Tile_X4Y8_RegFile/FrameStrobe[11] Tile_X4Y8_RegFile/FrameStrobe[12] Tile_X4Y8_RegFile/FrameStrobe[13]
+ Tile_X4Y8_RegFile/FrameStrobe[14] Tile_X4Y8_RegFile/FrameStrobe[15] Tile_X4Y8_RegFile/FrameStrobe[16]
+ Tile_X4Y8_RegFile/FrameStrobe[17] Tile_X4Y8_RegFile/FrameStrobe[18] Tile_X4Y8_RegFile/FrameStrobe[19]
+ Tile_X4Y8_RegFile/FrameStrobe[1] Tile_X4Y8_RegFile/FrameStrobe[2] Tile_X4Y8_RegFile/FrameStrobe[3]
+ Tile_X4Y8_RegFile/FrameStrobe[4] Tile_X4Y8_RegFile/FrameStrobe[5] Tile_X4Y8_RegFile/FrameStrobe[6]
+ Tile_X4Y8_RegFile/FrameStrobe[7] Tile_X4Y8_RegFile/FrameStrobe[8] Tile_X4Y8_RegFile/FrameStrobe[9]
+ Tile_X4Y7_RegFile/FrameStrobe[0] Tile_X4Y7_RegFile/FrameStrobe[10] Tile_X4Y7_RegFile/FrameStrobe[11]
+ Tile_X4Y7_RegFile/FrameStrobe[12] Tile_X4Y7_RegFile/FrameStrobe[13] Tile_X4Y7_RegFile/FrameStrobe[14]
+ Tile_X4Y7_RegFile/FrameStrobe[15] Tile_X4Y7_RegFile/FrameStrobe[16] Tile_X4Y7_RegFile/FrameStrobe[17]
+ Tile_X4Y7_RegFile/FrameStrobe[18] Tile_X4Y7_RegFile/FrameStrobe[19] Tile_X4Y7_RegFile/FrameStrobe[1]
+ Tile_X4Y7_RegFile/FrameStrobe[2] Tile_X4Y7_RegFile/FrameStrobe[3] Tile_X4Y7_RegFile/FrameStrobe[4]
+ Tile_X4Y7_RegFile/FrameStrobe[5] Tile_X4Y7_RegFile/FrameStrobe[6] Tile_X4Y7_RegFile/FrameStrobe[7]
+ Tile_X4Y7_RegFile/FrameStrobe[8] Tile_X4Y7_RegFile/FrameStrobe[9] Tile_X4Y8_RegFile/N1BEG[0]
+ Tile_X4Y8_RegFile/N1BEG[1] Tile_X4Y8_RegFile/N1BEG[2] Tile_X4Y8_RegFile/N1BEG[3]
+ Tile_X4Y9_RegFile/N1BEG[0] Tile_X4Y9_RegFile/N1BEG[1] Tile_X4Y9_RegFile/N1BEG[2]
+ Tile_X4Y9_RegFile/N1BEG[3] Tile_X4Y8_RegFile/N2BEG[0] Tile_X4Y8_RegFile/N2BEG[1]
+ Tile_X4Y8_RegFile/N2BEG[2] Tile_X4Y8_RegFile/N2BEG[3] Tile_X4Y8_RegFile/N2BEG[4]
+ Tile_X4Y8_RegFile/N2BEG[5] Tile_X4Y8_RegFile/N2BEG[6] Tile_X4Y8_RegFile/N2BEG[7]
+ Tile_X4Y7_RegFile/N2END[0] Tile_X4Y7_RegFile/N2END[1] Tile_X4Y7_RegFile/N2END[2]
+ Tile_X4Y7_RegFile/N2END[3] Tile_X4Y7_RegFile/N2END[4] Tile_X4Y7_RegFile/N2END[5]
+ Tile_X4Y7_RegFile/N2END[6] Tile_X4Y7_RegFile/N2END[7] Tile_X4Y8_RegFile/N2END[0]
+ Tile_X4Y8_RegFile/N2END[1] Tile_X4Y8_RegFile/N2END[2] Tile_X4Y8_RegFile/N2END[3]
+ Tile_X4Y8_RegFile/N2END[4] Tile_X4Y8_RegFile/N2END[5] Tile_X4Y8_RegFile/N2END[6]
+ Tile_X4Y8_RegFile/N2END[7] Tile_X4Y9_RegFile/N2BEG[0] Tile_X4Y9_RegFile/N2BEG[1]
+ Tile_X4Y9_RegFile/N2BEG[2] Tile_X4Y9_RegFile/N2BEG[3] Tile_X4Y9_RegFile/N2BEG[4]
+ Tile_X4Y9_RegFile/N2BEG[5] Tile_X4Y9_RegFile/N2BEG[6] Tile_X4Y9_RegFile/N2BEG[7]
+ Tile_X4Y8_RegFile/N4BEG[0] Tile_X4Y8_RegFile/N4BEG[10] Tile_X4Y8_RegFile/N4BEG[11]
+ Tile_X4Y8_RegFile/N4BEG[12] Tile_X4Y8_RegFile/N4BEG[13] Tile_X4Y8_RegFile/N4BEG[14]
+ Tile_X4Y8_RegFile/N4BEG[15] Tile_X4Y8_RegFile/N4BEG[1] Tile_X4Y8_RegFile/N4BEG[2]
+ Tile_X4Y8_RegFile/N4BEG[3] Tile_X4Y8_RegFile/N4BEG[4] Tile_X4Y8_RegFile/N4BEG[5]
+ Tile_X4Y8_RegFile/N4BEG[6] Tile_X4Y8_RegFile/N4BEG[7] Tile_X4Y8_RegFile/N4BEG[8]
+ Tile_X4Y8_RegFile/N4BEG[9] Tile_X4Y9_RegFile/N4BEG[0] Tile_X4Y9_RegFile/N4BEG[10]
+ Tile_X4Y9_RegFile/N4BEG[11] Tile_X4Y9_RegFile/N4BEG[12] Tile_X4Y9_RegFile/N4BEG[13]
+ Tile_X4Y9_RegFile/N4BEG[14] Tile_X4Y9_RegFile/N4BEG[15] Tile_X4Y9_RegFile/N4BEG[1]
+ Tile_X4Y9_RegFile/N4BEG[2] Tile_X4Y9_RegFile/N4BEG[3] Tile_X4Y9_RegFile/N4BEG[4]
+ Tile_X4Y9_RegFile/N4BEG[5] Tile_X4Y9_RegFile/N4BEG[6] Tile_X4Y9_RegFile/N4BEG[7]
+ Tile_X4Y9_RegFile/N4BEG[8] Tile_X4Y9_RegFile/N4BEG[9] Tile_X4Y8_RegFile/NN4BEG[0]
+ Tile_X4Y8_RegFile/NN4BEG[10] Tile_X4Y8_RegFile/NN4BEG[11] Tile_X4Y8_RegFile/NN4BEG[12]
+ Tile_X4Y8_RegFile/NN4BEG[13] Tile_X4Y8_RegFile/NN4BEG[14] Tile_X4Y8_RegFile/NN4BEG[15]
+ Tile_X4Y8_RegFile/NN4BEG[1] Tile_X4Y8_RegFile/NN4BEG[2] Tile_X4Y8_RegFile/NN4BEG[3]
+ Tile_X4Y8_RegFile/NN4BEG[4] Tile_X4Y8_RegFile/NN4BEG[5] Tile_X4Y8_RegFile/NN4BEG[6]
+ Tile_X4Y8_RegFile/NN4BEG[7] Tile_X4Y8_RegFile/NN4BEG[8] Tile_X4Y8_RegFile/NN4BEG[9]
+ Tile_X4Y9_RegFile/NN4BEG[0] Tile_X4Y9_RegFile/NN4BEG[10] Tile_X4Y9_RegFile/NN4BEG[11]
+ Tile_X4Y9_RegFile/NN4BEG[12] Tile_X4Y9_RegFile/NN4BEG[13] Tile_X4Y9_RegFile/NN4BEG[14]
+ Tile_X4Y9_RegFile/NN4BEG[15] Tile_X4Y9_RegFile/NN4BEG[1] Tile_X4Y9_RegFile/NN4BEG[2]
+ Tile_X4Y9_RegFile/NN4BEG[3] Tile_X4Y9_RegFile/NN4BEG[4] Tile_X4Y9_RegFile/NN4BEG[5]
+ Tile_X4Y9_RegFile/NN4BEG[6] Tile_X4Y9_RegFile/NN4BEG[7] Tile_X4Y9_RegFile/NN4BEG[8]
+ Tile_X4Y9_RegFile/NN4BEG[9] Tile_X4Y9_RegFile/S1END[0] Tile_X4Y9_RegFile/S1END[1]
+ Tile_X4Y9_RegFile/S1END[2] Tile_X4Y9_RegFile/S1END[3] Tile_X4Y8_RegFile/S1END[0]
+ Tile_X4Y8_RegFile/S1END[1] Tile_X4Y8_RegFile/S1END[2] Tile_X4Y8_RegFile/S1END[3]
+ Tile_X4Y9_RegFile/S2MID[0] Tile_X4Y9_RegFile/S2MID[1] Tile_X4Y9_RegFile/S2MID[2]
+ Tile_X4Y9_RegFile/S2MID[3] Tile_X4Y9_RegFile/S2MID[4] Tile_X4Y9_RegFile/S2MID[5]
+ Tile_X4Y9_RegFile/S2MID[6] Tile_X4Y9_RegFile/S2MID[7] Tile_X4Y9_RegFile/S2END[0]
+ Tile_X4Y9_RegFile/S2END[1] Tile_X4Y9_RegFile/S2END[2] Tile_X4Y9_RegFile/S2END[3]
+ Tile_X4Y9_RegFile/S2END[4] Tile_X4Y9_RegFile/S2END[5] Tile_X4Y9_RegFile/S2END[6]
+ Tile_X4Y9_RegFile/S2END[7] Tile_X4Y8_RegFile/S2END[0] Tile_X4Y8_RegFile/S2END[1]
+ Tile_X4Y8_RegFile/S2END[2] Tile_X4Y8_RegFile/S2END[3] Tile_X4Y8_RegFile/S2END[4]
+ Tile_X4Y8_RegFile/S2END[5] Tile_X4Y8_RegFile/S2END[6] Tile_X4Y8_RegFile/S2END[7]
+ Tile_X4Y8_RegFile/S2MID[0] Tile_X4Y8_RegFile/S2MID[1] Tile_X4Y8_RegFile/S2MID[2]
+ Tile_X4Y8_RegFile/S2MID[3] Tile_X4Y8_RegFile/S2MID[4] Tile_X4Y8_RegFile/S2MID[5]
+ Tile_X4Y8_RegFile/S2MID[6] Tile_X4Y8_RegFile/S2MID[7] Tile_X4Y9_RegFile/S4END[0]
+ Tile_X4Y9_RegFile/S4END[10] Tile_X4Y9_RegFile/S4END[11] Tile_X4Y9_RegFile/S4END[12]
+ Tile_X4Y9_RegFile/S4END[13] Tile_X4Y9_RegFile/S4END[14] Tile_X4Y9_RegFile/S4END[15]
+ Tile_X4Y9_RegFile/S4END[1] Tile_X4Y9_RegFile/S4END[2] Tile_X4Y9_RegFile/S4END[3]
+ Tile_X4Y9_RegFile/S4END[4] Tile_X4Y9_RegFile/S4END[5] Tile_X4Y9_RegFile/S4END[6]
+ Tile_X4Y9_RegFile/S4END[7] Tile_X4Y9_RegFile/S4END[8] Tile_X4Y9_RegFile/S4END[9]
+ Tile_X4Y8_RegFile/S4END[0] Tile_X4Y8_RegFile/S4END[10] Tile_X4Y8_RegFile/S4END[11]
+ Tile_X4Y8_RegFile/S4END[12] Tile_X4Y8_RegFile/S4END[13] Tile_X4Y8_RegFile/S4END[14]
+ Tile_X4Y8_RegFile/S4END[15] Tile_X4Y8_RegFile/S4END[1] Tile_X4Y8_RegFile/S4END[2]
+ Tile_X4Y8_RegFile/S4END[3] Tile_X4Y8_RegFile/S4END[4] Tile_X4Y8_RegFile/S4END[5]
+ Tile_X4Y8_RegFile/S4END[6] Tile_X4Y8_RegFile/S4END[7] Tile_X4Y8_RegFile/S4END[8]
+ Tile_X4Y8_RegFile/S4END[9] Tile_X4Y9_RegFile/SS4END[0] Tile_X4Y9_RegFile/SS4END[10]
+ Tile_X4Y9_RegFile/SS4END[11] Tile_X4Y9_RegFile/SS4END[12] Tile_X4Y9_RegFile/SS4END[13]
+ Tile_X4Y9_RegFile/SS4END[14] Tile_X4Y9_RegFile/SS4END[15] Tile_X4Y9_RegFile/SS4END[1]
+ Tile_X4Y9_RegFile/SS4END[2] Tile_X4Y9_RegFile/SS4END[3] Tile_X4Y9_RegFile/SS4END[4]
+ Tile_X4Y9_RegFile/SS4END[5] Tile_X4Y9_RegFile/SS4END[6] Tile_X4Y9_RegFile/SS4END[7]
+ Tile_X4Y9_RegFile/SS4END[8] Tile_X4Y9_RegFile/SS4END[9] Tile_X4Y8_RegFile/SS4END[0]
+ Tile_X4Y8_RegFile/SS4END[10] Tile_X4Y8_RegFile/SS4END[11] Tile_X4Y8_RegFile/SS4END[12]
+ Tile_X4Y8_RegFile/SS4END[13] Tile_X4Y8_RegFile/SS4END[14] Tile_X4Y8_RegFile/SS4END[15]
+ Tile_X4Y8_RegFile/SS4END[1] Tile_X4Y8_RegFile/SS4END[2] Tile_X4Y8_RegFile/SS4END[3]
+ Tile_X4Y8_RegFile/SS4END[4] Tile_X4Y8_RegFile/SS4END[5] Tile_X4Y8_RegFile/SS4END[6]
+ Tile_X4Y8_RegFile/SS4END[7] Tile_X4Y8_RegFile/SS4END[8] Tile_X4Y8_RegFile/SS4END[9]
+ Tile_X4Y8_RegFile/UserCLK Tile_X4Y7_RegFile/UserCLK VGND VPWR Tile_X3Y8_LUT4AB/W1END[0]
+ Tile_X3Y8_LUT4AB/W1END[1] Tile_X3Y8_LUT4AB/W1END[2] Tile_X3Y8_LUT4AB/W1END[3] Tile_X5Y8_LUT4AB/W1BEG[0]
+ Tile_X5Y8_LUT4AB/W1BEG[1] Tile_X5Y8_LUT4AB/W1BEG[2] Tile_X5Y8_LUT4AB/W1BEG[3] Tile_X3Y8_LUT4AB/W2MID[0]
+ Tile_X3Y8_LUT4AB/W2MID[1] Tile_X3Y8_LUT4AB/W2MID[2] Tile_X3Y8_LUT4AB/W2MID[3] Tile_X3Y8_LUT4AB/W2MID[4]
+ Tile_X3Y8_LUT4AB/W2MID[5] Tile_X3Y8_LUT4AB/W2MID[6] Tile_X3Y8_LUT4AB/W2MID[7] Tile_X3Y8_LUT4AB/W2END[0]
+ Tile_X3Y8_LUT4AB/W2END[1] Tile_X3Y8_LUT4AB/W2END[2] Tile_X3Y8_LUT4AB/W2END[3] Tile_X3Y8_LUT4AB/W2END[4]
+ Tile_X3Y8_LUT4AB/W2END[5] Tile_X3Y8_LUT4AB/W2END[6] Tile_X3Y8_LUT4AB/W2END[7] Tile_X5Y8_LUT4AB/W2BEGb[0]
+ Tile_X5Y8_LUT4AB/W2BEGb[1] Tile_X5Y8_LUT4AB/W2BEGb[2] Tile_X5Y8_LUT4AB/W2BEGb[3]
+ Tile_X5Y8_LUT4AB/W2BEGb[4] Tile_X5Y8_LUT4AB/W2BEGb[5] Tile_X5Y8_LUT4AB/W2BEGb[6]
+ Tile_X5Y8_LUT4AB/W2BEGb[7] Tile_X5Y8_LUT4AB/W2BEG[0] Tile_X5Y8_LUT4AB/W2BEG[1] Tile_X5Y8_LUT4AB/W2BEG[2]
+ Tile_X5Y8_LUT4AB/W2BEG[3] Tile_X5Y8_LUT4AB/W2BEG[4] Tile_X5Y8_LUT4AB/W2BEG[5] Tile_X5Y8_LUT4AB/W2BEG[6]
+ Tile_X5Y8_LUT4AB/W2BEG[7] Tile_X3Y8_LUT4AB/W6END[0] Tile_X3Y8_LUT4AB/W6END[10] Tile_X3Y8_LUT4AB/W6END[11]
+ Tile_X3Y8_LUT4AB/W6END[1] Tile_X3Y8_LUT4AB/W6END[2] Tile_X3Y8_LUT4AB/W6END[3] Tile_X3Y8_LUT4AB/W6END[4]
+ Tile_X3Y8_LUT4AB/W6END[5] Tile_X3Y8_LUT4AB/W6END[6] Tile_X3Y8_LUT4AB/W6END[7] Tile_X3Y8_LUT4AB/W6END[8]
+ Tile_X3Y8_LUT4AB/W6END[9] Tile_X5Y8_LUT4AB/W6BEG[0] Tile_X5Y8_LUT4AB/W6BEG[10] Tile_X5Y8_LUT4AB/W6BEG[11]
+ Tile_X5Y8_LUT4AB/W6BEG[1] Tile_X5Y8_LUT4AB/W6BEG[2] Tile_X5Y8_LUT4AB/W6BEG[3] Tile_X5Y8_LUT4AB/W6BEG[4]
+ Tile_X5Y8_LUT4AB/W6BEG[5] Tile_X5Y8_LUT4AB/W6BEG[6] Tile_X5Y8_LUT4AB/W6BEG[7] Tile_X5Y8_LUT4AB/W6BEG[8]
+ Tile_X5Y8_LUT4AB/W6BEG[9] Tile_X3Y8_LUT4AB/WW4END[0] Tile_X3Y8_LUT4AB/WW4END[10]
+ Tile_X3Y8_LUT4AB/WW4END[11] Tile_X3Y8_LUT4AB/WW4END[12] Tile_X3Y8_LUT4AB/WW4END[13]
+ Tile_X3Y8_LUT4AB/WW4END[14] Tile_X3Y8_LUT4AB/WW4END[15] Tile_X3Y8_LUT4AB/WW4END[1]
+ Tile_X3Y8_LUT4AB/WW4END[2] Tile_X3Y8_LUT4AB/WW4END[3] Tile_X3Y8_LUT4AB/WW4END[4]
+ Tile_X3Y8_LUT4AB/WW4END[5] Tile_X3Y8_LUT4AB/WW4END[6] Tile_X3Y8_LUT4AB/WW4END[7]
+ Tile_X3Y8_LUT4AB/WW4END[8] Tile_X3Y8_LUT4AB/WW4END[9] Tile_X5Y8_LUT4AB/WW4BEG[0]
+ Tile_X5Y8_LUT4AB/WW4BEG[10] Tile_X5Y8_LUT4AB/WW4BEG[11] Tile_X5Y8_LUT4AB/WW4BEG[12]
+ Tile_X5Y8_LUT4AB/WW4BEG[13] Tile_X5Y8_LUT4AB/WW4BEG[14] Tile_X5Y8_LUT4AB/WW4BEG[15]
+ Tile_X5Y8_LUT4AB/WW4BEG[1] Tile_X5Y8_LUT4AB/WW4BEG[2] Tile_X5Y8_LUT4AB/WW4BEG[3]
+ Tile_X5Y8_LUT4AB/WW4BEG[4] Tile_X5Y8_LUT4AB/WW4BEG[5] Tile_X5Y8_LUT4AB/WW4BEG[6]
+ Tile_X5Y8_LUT4AB/WW4BEG[7] Tile_X5Y8_LUT4AB/WW4BEG[8] Tile_X5Y8_LUT4AB/WW4BEG[9]
+ RegFile
XTile_X6Y1_LUT4AB Tile_X6Y2_LUT4AB/Co Tile_X6Y1_LUT4AB/Co Tile_X6Y1_LUT4AB/E1BEG[0]
+ Tile_X6Y1_LUT4AB/E1BEG[1] Tile_X6Y1_LUT4AB/E1BEG[2] Tile_X6Y1_LUT4AB/E1BEG[3] Tile_X6Y1_LUT4AB/E1END[0]
+ Tile_X6Y1_LUT4AB/E1END[1] Tile_X6Y1_LUT4AB/E1END[2] Tile_X6Y1_LUT4AB/E1END[3] Tile_X6Y1_LUT4AB/E2BEG[0]
+ Tile_X6Y1_LUT4AB/E2BEG[1] Tile_X6Y1_LUT4AB/E2BEG[2] Tile_X6Y1_LUT4AB/E2BEG[3] Tile_X6Y1_LUT4AB/E2BEG[4]
+ Tile_X6Y1_LUT4AB/E2BEG[5] Tile_X6Y1_LUT4AB/E2BEG[6] Tile_X6Y1_LUT4AB/E2BEG[7] Tile_X6Y1_LUT4AB/E2BEGb[0]
+ Tile_X6Y1_LUT4AB/E2BEGb[1] Tile_X6Y1_LUT4AB/E2BEGb[2] Tile_X6Y1_LUT4AB/E2BEGb[3]
+ Tile_X6Y1_LUT4AB/E2BEGb[4] Tile_X6Y1_LUT4AB/E2BEGb[5] Tile_X6Y1_LUT4AB/E2BEGb[6]
+ Tile_X6Y1_LUT4AB/E2BEGb[7] Tile_X6Y1_LUT4AB/E2END[0] Tile_X6Y1_LUT4AB/E2END[1] Tile_X6Y1_LUT4AB/E2END[2]
+ Tile_X6Y1_LUT4AB/E2END[3] Tile_X6Y1_LUT4AB/E2END[4] Tile_X6Y1_LUT4AB/E2END[5] Tile_X6Y1_LUT4AB/E2END[6]
+ Tile_X6Y1_LUT4AB/E2END[7] Tile_X6Y1_LUT4AB/E2MID[0] Tile_X6Y1_LUT4AB/E2MID[1] Tile_X6Y1_LUT4AB/E2MID[2]
+ Tile_X6Y1_LUT4AB/E2MID[3] Tile_X6Y1_LUT4AB/E2MID[4] Tile_X6Y1_LUT4AB/E2MID[5] Tile_X6Y1_LUT4AB/E2MID[6]
+ Tile_X6Y1_LUT4AB/E2MID[7] Tile_X6Y1_LUT4AB/E6BEG[0] Tile_X6Y1_LUT4AB/E6BEG[10] Tile_X6Y1_LUT4AB/E6BEG[11]
+ Tile_X6Y1_LUT4AB/E6BEG[1] Tile_X6Y1_LUT4AB/E6BEG[2] Tile_X6Y1_LUT4AB/E6BEG[3] Tile_X6Y1_LUT4AB/E6BEG[4]
+ Tile_X6Y1_LUT4AB/E6BEG[5] Tile_X6Y1_LUT4AB/E6BEG[6] Tile_X6Y1_LUT4AB/E6BEG[7] Tile_X6Y1_LUT4AB/E6BEG[8]
+ Tile_X6Y1_LUT4AB/E6BEG[9] Tile_X6Y1_LUT4AB/E6END[0] Tile_X6Y1_LUT4AB/E6END[10] Tile_X6Y1_LUT4AB/E6END[11]
+ Tile_X6Y1_LUT4AB/E6END[1] Tile_X6Y1_LUT4AB/E6END[2] Tile_X6Y1_LUT4AB/E6END[3] Tile_X6Y1_LUT4AB/E6END[4]
+ Tile_X6Y1_LUT4AB/E6END[5] Tile_X6Y1_LUT4AB/E6END[6] Tile_X6Y1_LUT4AB/E6END[7] Tile_X6Y1_LUT4AB/E6END[8]
+ Tile_X6Y1_LUT4AB/E6END[9] Tile_X6Y1_LUT4AB/EE4BEG[0] Tile_X6Y1_LUT4AB/EE4BEG[10]
+ Tile_X6Y1_LUT4AB/EE4BEG[11] Tile_X6Y1_LUT4AB/EE4BEG[12] Tile_X6Y1_LUT4AB/EE4BEG[13]
+ Tile_X6Y1_LUT4AB/EE4BEG[14] Tile_X6Y1_LUT4AB/EE4BEG[15] Tile_X6Y1_LUT4AB/EE4BEG[1]
+ Tile_X6Y1_LUT4AB/EE4BEG[2] Tile_X6Y1_LUT4AB/EE4BEG[3] Tile_X6Y1_LUT4AB/EE4BEG[4]
+ Tile_X6Y1_LUT4AB/EE4BEG[5] Tile_X6Y1_LUT4AB/EE4BEG[6] Tile_X6Y1_LUT4AB/EE4BEG[7]
+ Tile_X6Y1_LUT4AB/EE4BEG[8] Tile_X6Y1_LUT4AB/EE4BEG[9] Tile_X6Y1_LUT4AB/EE4END[0]
+ Tile_X6Y1_LUT4AB/EE4END[10] Tile_X6Y1_LUT4AB/EE4END[11] Tile_X6Y1_LUT4AB/EE4END[12]
+ Tile_X6Y1_LUT4AB/EE4END[13] Tile_X6Y1_LUT4AB/EE4END[14] Tile_X6Y1_LUT4AB/EE4END[15]
+ Tile_X6Y1_LUT4AB/EE4END[1] Tile_X6Y1_LUT4AB/EE4END[2] Tile_X6Y1_LUT4AB/EE4END[3]
+ Tile_X6Y1_LUT4AB/EE4END[4] Tile_X6Y1_LUT4AB/EE4END[5] Tile_X6Y1_LUT4AB/EE4END[6]
+ Tile_X6Y1_LUT4AB/EE4END[7] Tile_X6Y1_LUT4AB/EE4END[8] Tile_X6Y1_LUT4AB/EE4END[9]
+ Tile_X6Y1_LUT4AB/FrameData[0] Tile_X6Y1_LUT4AB/FrameData[10] Tile_X6Y1_LUT4AB/FrameData[11]
+ Tile_X6Y1_LUT4AB/FrameData[12] Tile_X6Y1_LUT4AB/FrameData[13] Tile_X6Y1_LUT4AB/FrameData[14]
+ Tile_X6Y1_LUT4AB/FrameData[15] Tile_X6Y1_LUT4AB/FrameData[16] Tile_X6Y1_LUT4AB/FrameData[17]
+ Tile_X6Y1_LUT4AB/FrameData[18] Tile_X6Y1_LUT4AB/FrameData[19] Tile_X6Y1_LUT4AB/FrameData[1]
+ Tile_X6Y1_LUT4AB/FrameData[20] Tile_X6Y1_LUT4AB/FrameData[21] Tile_X6Y1_LUT4AB/FrameData[22]
+ Tile_X6Y1_LUT4AB/FrameData[23] Tile_X6Y1_LUT4AB/FrameData[24] Tile_X6Y1_LUT4AB/FrameData[25]
+ Tile_X6Y1_LUT4AB/FrameData[26] Tile_X6Y1_LUT4AB/FrameData[27] Tile_X6Y1_LUT4AB/FrameData[28]
+ Tile_X6Y1_LUT4AB/FrameData[29] Tile_X6Y1_LUT4AB/FrameData[2] Tile_X6Y1_LUT4AB/FrameData[30]
+ Tile_X6Y1_LUT4AB/FrameData[31] Tile_X6Y1_LUT4AB/FrameData[3] Tile_X6Y1_LUT4AB/FrameData[4]
+ Tile_X6Y1_LUT4AB/FrameData[5] Tile_X6Y1_LUT4AB/FrameData[6] Tile_X6Y1_LUT4AB/FrameData[7]
+ Tile_X6Y1_LUT4AB/FrameData[8] Tile_X6Y1_LUT4AB/FrameData[9] Tile_X6Y1_LUT4AB/FrameData_O[0]
+ Tile_X6Y1_LUT4AB/FrameData_O[10] Tile_X6Y1_LUT4AB/FrameData_O[11] Tile_X6Y1_LUT4AB/FrameData_O[12]
+ Tile_X6Y1_LUT4AB/FrameData_O[13] Tile_X6Y1_LUT4AB/FrameData_O[14] Tile_X6Y1_LUT4AB/FrameData_O[15]
+ Tile_X6Y1_LUT4AB/FrameData_O[16] Tile_X6Y1_LUT4AB/FrameData_O[17] Tile_X6Y1_LUT4AB/FrameData_O[18]
+ Tile_X6Y1_LUT4AB/FrameData_O[19] Tile_X6Y1_LUT4AB/FrameData_O[1] Tile_X6Y1_LUT4AB/FrameData_O[20]
+ Tile_X6Y1_LUT4AB/FrameData_O[21] Tile_X6Y1_LUT4AB/FrameData_O[22] Tile_X6Y1_LUT4AB/FrameData_O[23]
+ Tile_X6Y1_LUT4AB/FrameData_O[24] Tile_X6Y1_LUT4AB/FrameData_O[25] Tile_X6Y1_LUT4AB/FrameData_O[26]
+ Tile_X6Y1_LUT4AB/FrameData_O[27] Tile_X6Y1_LUT4AB/FrameData_O[28] Tile_X6Y1_LUT4AB/FrameData_O[29]
+ Tile_X6Y1_LUT4AB/FrameData_O[2] Tile_X6Y1_LUT4AB/FrameData_O[30] Tile_X6Y1_LUT4AB/FrameData_O[31]
+ Tile_X6Y1_LUT4AB/FrameData_O[3] Tile_X6Y1_LUT4AB/FrameData_O[4] Tile_X6Y1_LUT4AB/FrameData_O[5]
+ Tile_X6Y1_LUT4AB/FrameData_O[6] Tile_X6Y1_LUT4AB/FrameData_O[7] Tile_X6Y1_LUT4AB/FrameData_O[8]
+ Tile_X6Y1_LUT4AB/FrameData_O[9] Tile_X6Y1_LUT4AB/FrameStrobe[0] Tile_X6Y1_LUT4AB/FrameStrobe[10]
+ Tile_X6Y1_LUT4AB/FrameStrobe[11] Tile_X6Y1_LUT4AB/FrameStrobe[12] Tile_X6Y1_LUT4AB/FrameStrobe[13]
+ Tile_X6Y1_LUT4AB/FrameStrobe[14] Tile_X6Y1_LUT4AB/FrameStrobe[15] Tile_X6Y1_LUT4AB/FrameStrobe[16]
+ Tile_X6Y1_LUT4AB/FrameStrobe[17] Tile_X6Y1_LUT4AB/FrameStrobe[18] Tile_X6Y1_LUT4AB/FrameStrobe[19]
+ Tile_X6Y1_LUT4AB/FrameStrobe[1] Tile_X6Y1_LUT4AB/FrameStrobe[2] Tile_X6Y1_LUT4AB/FrameStrobe[3]
+ Tile_X6Y1_LUT4AB/FrameStrobe[4] Tile_X6Y1_LUT4AB/FrameStrobe[5] Tile_X6Y1_LUT4AB/FrameStrobe[6]
+ Tile_X6Y1_LUT4AB/FrameStrobe[7] Tile_X6Y1_LUT4AB/FrameStrobe[8] Tile_X6Y1_LUT4AB/FrameStrobe[9]
+ Tile_X6Y1_LUT4AB/FrameStrobe_O[0] Tile_X6Y1_LUT4AB/FrameStrobe_O[10] Tile_X6Y1_LUT4AB/FrameStrobe_O[11]
+ Tile_X6Y1_LUT4AB/FrameStrobe_O[12] Tile_X6Y1_LUT4AB/FrameStrobe_O[13] Tile_X6Y1_LUT4AB/FrameStrobe_O[14]
+ Tile_X6Y1_LUT4AB/FrameStrobe_O[15] Tile_X6Y1_LUT4AB/FrameStrobe_O[16] Tile_X6Y1_LUT4AB/FrameStrobe_O[17]
+ Tile_X6Y1_LUT4AB/FrameStrobe_O[18] Tile_X6Y1_LUT4AB/FrameStrobe_O[19] Tile_X6Y1_LUT4AB/FrameStrobe_O[1]
+ Tile_X6Y1_LUT4AB/FrameStrobe_O[2] Tile_X6Y1_LUT4AB/FrameStrobe_O[3] Tile_X6Y1_LUT4AB/FrameStrobe_O[4]
+ Tile_X6Y1_LUT4AB/FrameStrobe_O[5] Tile_X6Y1_LUT4AB/FrameStrobe_O[6] Tile_X6Y1_LUT4AB/FrameStrobe_O[7]
+ Tile_X6Y1_LUT4AB/FrameStrobe_O[8] Tile_X6Y1_LUT4AB/FrameStrobe_O[9] Tile_X6Y1_LUT4AB/N1BEG[0]
+ Tile_X6Y1_LUT4AB/N1BEG[1] Tile_X6Y1_LUT4AB/N1BEG[2] Tile_X6Y1_LUT4AB/N1BEG[3] Tile_X6Y2_LUT4AB/N1BEG[0]
+ Tile_X6Y2_LUT4AB/N1BEG[1] Tile_X6Y2_LUT4AB/N1BEG[2] Tile_X6Y2_LUT4AB/N1BEG[3] Tile_X6Y1_LUT4AB/N2BEG[0]
+ Tile_X6Y1_LUT4AB/N2BEG[1] Tile_X6Y1_LUT4AB/N2BEG[2] Tile_X6Y1_LUT4AB/N2BEG[3] Tile_X6Y1_LUT4AB/N2BEG[4]
+ Tile_X6Y1_LUT4AB/N2BEG[5] Tile_X6Y1_LUT4AB/N2BEG[6] Tile_X6Y1_LUT4AB/N2BEG[7] Tile_X6Y1_LUT4AB/N2BEGb[0]
+ Tile_X6Y1_LUT4AB/N2BEGb[1] Tile_X6Y1_LUT4AB/N2BEGb[2] Tile_X6Y1_LUT4AB/N2BEGb[3]
+ Tile_X6Y1_LUT4AB/N2BEGb[4] Tile_X6Y1_LUT4AB/N2BEGb[5] Tile_X6Y1_LUT4AB/N2BEGb[6]
+ Tile_X6Y1_LUT4AB/N2BEGb[7] Tile_X6Y1_LUT4AB/N2END[0] Tile_X6Y1_LUT4AB/N2END[1] Tile_X6Y1_LUT4AB/N2END[2]
+ Tile_X6Y1_LUT4AB/N2END[3] Tile_X6Y1_LUT4AB/N2END[4] Tile_X6Y1_LUT4AB/N2END[5] Tile_X6Y1_LUT4AB/N2END[6]
+ Tile_X6Y1_LUT4AB/N2END[7] Tile_X6Y2_LUT4AB/N2BEG[0] Tile_X6Y2_LUT4AB/N2BEG[1] Tile_X6Y2_LUT4AB/N2BEG[2]
+ Tile_X6Y2_LUT4AB/N2BEG[3] Tile_X6Y2_LUT4AB/N2BEG[4] Tile_X6Y2_LUT4AB/N2BEG[5] Tile_X6Y2_LUT4AB/N2BEG[6]
+ Tile_X6Y2_LUT4AB/N2BEG[7] Tile_X6Y1_LUT4AB/N4BEG[0] Tile_X6Y1_LUT4AB/N4BEG[10] Tile_X6Y1_LUT4AB/N4BEG[11]
+ Tile_X6Y1_LUT4AB/N4BEG[12] Tile_X6Y1_LUT4AB/N4BEG[13] Tile_X6Y1_LUT4AB/N4BEG[14]
+ Tile_X6Y1_LUT4AB/N4BEG[15] Tile_X6Y1_LUT4AB/N4BEG[1] Tile_X6Y1_LUT4AB/N4BEG[2] Tile_X6Y1_LUT4AB/N4BEG[3]
+ Tile_X6Y1_LUT4AB/N4BEG[4] Tile_X6Y1_LUT4AB/N4BEG[5] Tile_X6Y1_LUT4AB/N4BEG[6] Tile_X6Y1_LUT4AB/N4BEG[7]
+ Tile_X6Y1_LUT4AB/N4BEG[8] Tile_X6Y1_LUT4AB/N4BEG[9] Tile_X6Y2_LUT4AB/N4BEG[0] Tile_X6Y2_LUT4AB/N4BEG[10]
+ Tile_X6Y2_LUT4AB/N4BEG[11] Tile_X6Y2_LUT4AB/N4BEG[12] Tile_X6Y2_LUT4AB/N4BEG[13]
+ Tile_X6Y2_LUT4AB/N4BEG[14] Tile_X6Y2_LUT4AB/N4BEG[15] Tile_X6Y2_LUT4AB/N4BEG[1]
+ Tile_X6Y2_LUT4AB/N4BEG[2] Tile_X6Y2_LUT4AB/N4BEG[3] Tile_X6Y2_LUT4AB/N4BEG[4] Tile_X6Y2_LUT4AB/N4BEG[5]
+ Tile_X6Y2_LUT4AB/N4BEG[6] Tile_X6Y2_LUT4AB/N4BEG[7] Tile_X6Y2_LUT4AB/N4BEG[8] Tile_X6Y2_LUT4AB/N4BEG[9]
+ Tile_X6Y1_LUT4AB/NN4BEG[0] Tile_X6Y1_LUT4AB/NN4BEG[10] Tile_X6Y1_LUT4AB/NN4BEG[11]
+ Tile_X6Y1_LUT4AB/NN4BEG[12] Tile_X6Y1_LUT4AB/NN4BEG[13] Tile_X6Y1_LUT4AB/NN4BEG[14]
+ Tile_X6Y1_LUT4AB/NN4BEG[15] Tile_X6Y1_LUT4AB/NN4BEG[1] Tile_X6Y1_LUT4AB/NN4BEG[2]
+ Tile_X6Y1_LUT4AB/NN4BEG[3] Tile_X6Y1_LUT4AB/NN4BEG[4] Tile_X6Y1_LUT4AB/NN4BEG[5]
+ Tile_X6Y1_LUT4AB/NN4BEG[6] Tile_X6Y1_LUT4AB/NN4BEG[7] Tile_X6Y1_LUT4AB/NN4BEG[8]
+ Tile_X6Y1_LUT4AB/NN4BEG[9] Tile_X6Y2_LUT4AB/NN4BEG[0] Tile_X6Y2_LUT4AB/NN4BEG[10]
+ Tile_X6Y2_LUT4AB/NN4BEG[11] Tile_X6Y2_LUT4AB/NN4BEG[12] Tile_X6Y2_LUT4AB/NN4BEG[13]
+ Tile_X6Y2_LUT4AB/NN4BEG[14] Tile_X6Y2_LUT4AB/NN4BEG[15] Tile_X6Y2_LUT4AB/NN4BEG[1]
+ Tile_X6Y2_LUT4AB/NN4BEG[2] Tile_X6Y2_LUT4AB/NN4BEG[3] Tile_X6Y2_LUT4AB/NN4BEG[4]
+ Tile_X6Y2_LUT4AB/NN4BEG[5] Tile_X6Y2_LUT4AB/NN4BEG[6] Tile_X6Y2_LUT4AB/NN4BEG[7]
+ Tile_X6Y2_LUT4AB/NN4BEG[8] Tile_X6Y2_LUT4AB/NN4BEG[9] Tile_X6Y2_LUT4AB/S1END[0]
+ Tile_X6Y2_LUT4AB/S1END[1] Tile_X6Y2_LUT4AB/S1END[2] Tile_X6Y2_LUT4AB/S1END[3] Tile_X6Y1_LUT4AB/S1END[0]
+ Tile_X6Y1_LUT4AB/S1END[1] Tile_X6Y1_LUT4AB/S1END[2] Tile_X6Y1_LUT4AB/S1END[3] Tile_X6Y2_LUT4AB/S2MID[0]
+ Tile_X6Y2_LUT4AB/S2MID[1] Tile_X6Y2_LUT4AB/S2MID[2] Tile_X6Y2_LUT4AB/S2MID[3] Tile_X6Y2_LUT4AB/S2MID[4]
+ Tile_X6Y2_LUT4AB/S2MID[5] Tile_X6Y2_LUT4AB/S2MID[6] Tile_X6Y2_LUT4AB/S2MID[7] Tile_X6Y2_LUT4AB/S2END[0]
+ Tile_X6Y2_LUT4AB/S2END[1] Tile_X6Y2_LUT4AB/S2END[2] Tile_X6Y2_LUT4AB/S2END[3] Tile_X6Y2_LUT4AB/S2END[4]
+ Tile_X6Y2_LUT4AB/S2END[5] Tile_X6Y2_LUT4AB/S2END[6] Tile_X6Y2_LUT4AB/S2END[7] Tile_X6Y1_LUT4AB/S2END[0]
+ Tile_X6Y1_LUT4AB/S2END[1] Tile_X6Y1_LUT4AB/S2END[2] Tile_X6Y1_LUT4AB/S2END[3] Tile_X6Y1_LUT4AB/S2END[4]
+ Tile_X6Y1_LUT4AB/S2END[5] Tile_X6Y1_LUT4AB/S2END[6] Tile_X6Y1_LUT4AB/S2END[7] Tile_X6Y1_LUT4AB/S2MID[0]
+ Tile_X6Y1_LUT4AB/S2MID[1] Tile_X6Y1_LUT4AB/S2MID[2] Tile_X6Y1_LUT4AB/S2MID[3] Tile_X6Y1_LUT4AB/S2MID[4]
+ Tile_X6Y1_LUT4AB/S2MID[5] Tile_X6Y1_LUT4AB/S2MID[6] Tile_X6Y1_LUT4AB/S2MID[7] Tile_X6Y2_LUT4AB/S4END[0]
+ Tile_X6Y2_LUT4AB/S4END[10] Tile_X6Y2_LUT4AB/S4END[11] Tile_X6Y2_LUT4AB/S4END[12]
+ Tile_X6Y2_LUT4AB/S4END[13] Tile_X6Y2_LUT4AB/S4END[14] Tile_X6Y2_LUT4AB/S4END[15]
+ Tile_X6Y2_LUT4AB/S4END[1] Tile_X6Y2_LUT4AB/S4END[2] Tile_X6Y2_LUT4AB/S4END[3] Tile_X6Y2_LUT4AB/S4END[4]
+ Tile_X6Y2_LUT4AB/S4END[5] Tile_X6Y2_LUT4AB/S4END[6] Tile_X6Y2_LUT4AB/S4END[7] Tile_X6Y2_LUT4AB/S4END[8]
+ Tile_X6Y2_LUT4AB/S4END[9] Tile_X6Y1_LUT4AB/S4END[0] Tile_X6Y1_LUT4AB/S4END[10] Tile_X6Y1_LUT4AB/S4END[11]
+ Tile_X6Y1_LUT4AB/S4END[12] Tile_X6Y1_LUT4AB/S4END[13] Tile_X6Y1_LUT4AB/S4END[14]
+ Tile_X6Y1_LUT4AB/S4END[15] Tile_X6Y1_LUT4AB/S4END[1] Tile_X6Y1_LUT4AB/S4END[2] Tile_X6Y1_LUT4AB/S4END[3]
+ Tile_X6Y1_LUT4AB/S4END[4] Tile_X6Y1_LUT4AB/S4END[5] Tile_X6Y1_LUT4AB/S4END[6] Tile_X6Y1_LUT4AB/S4END[7]
+ Tile_X6Y1_LUT4AB/S4END[8] Tile_X6Y1_LUT4AB/S4END[9] Tile_X6Y2_LUT4AB/SS4END[0] Tile_X6Y2_LUT4AB/SS4END[10]
+ Tile_X6Y2_LUT4AB/SS4END[11] Tile_X6Y2_LUT4AB/SS4END[12] Tile_X6Y2_LUT4AB/SS4END[13]
+ Tile_X6Y2_LUT4AB/SS4END[14] Tile_X6Y2_LUT4AB/SS4END[15] Tile_X6Y2_LUT4AB/SS4END[1]
+ Tile_X6Y2_LUT4AB/SS4END[2] Tile_X6Y2_LUT4AB/SS4END[3] Tile_X6Y2_LUT4AB/SS4END[4]
+ Tile_X6Y2_LUT4AB/SS4END[5] Tile_X6Y2_LUT4AB/SS4END[6] Tile_X6Y2_LUT4AB/SS4END[7]
+ Tile_X6Y2_LUT4AB/SS4END[8] Tile_X6Y2_LUT4AB/SS4END[9] Tile_X6Y1_LUT4AB/SS4END[0]
+ Tile_X6Y1_LUT4AB/SS4END[10] Tile_X6Y1_LUT4AB/SS4END[11] Tile_X6Y1_LUT4AB/SS4END[12]
+ Tile_X6Y1_LUT4AB/SS4END[13] Tile_X6Y1_LUT4AB/SS4END[14] Tile_X6Y1_LUT4AB/SS4END[15]
+ Tile_X6Y1_LUT4AB/SS4END[1] Tile_X6Y1_LUT4AB/SS4END[2] Tile_X6Y1_LUT4AB/SS4END[3]
+ Tile_X6Y1_LUT4AB/SS4END[4] Tile_X6Y1_LUT4AB/SS4END[5] Tile_X6Y1_LUT4AB/SS4END[6]
+ Tile_X6Y1_LUT4AB/SS4END[7] Tile_X6Y1_LUT4AB/SS4END[8] Tile_X6Y1_LUT4AB/SS4END[9]
+ Tile_X6Y1_LUT4AB/UserCLK Tile_X6Y1_LUT4AB/UserCLKo VGND VPWR Tile_X6Y1_LUT4AB/W1BEG[0]
+ Tile_X6Y1_LUT4AB/W1BEG[1] Tile_X6Y1_LUT4AB/W1BEG[2] Tile_X6Y1_LUT4AB/W1BEG[3] Tile_X6Y1_LUT4AB/W1END[0]
+ Tile_X6Y1_LUT4AB/W1END[1] Tile_X6Y1_LUT4AB/W1END[2] Tile_X6Y1_LUT4AB/W1END[3] Tile_X6Y1_LUT4AB/W2BEG[0]
+ Tile_X6Y1_LUT4AB/W2BEG[1] Tile_X6Y1_LUT4AB/W2BEG[2] Tile_X6Y1_LUT4AB/W2BEG[3] Tile_X6Y1_LUT4AB/W2BEG[4]
+ Tile_X6Y1_LUT4AB/W2BEG[5] Tile_X6Y1_LUT4AB/W2BEG[6] Tile_X6Y1_LUT4AB/W2BEG[7] Tile_X5Y1_LUT4AB/W2END[0]
+ Tile_X5Y1_LUT4AB/W2END[1] Tile_X5Y1_LUT4AB/W2END[2] Tile_X5Y1_LUT4AB/W2END[3] Tile_X5Y1_LUT4AB/W2END[4]
+ Tile_X5Y1_LUT4AB/W2END[5] Tile_X5Y1_LUT4AB/W2END[6] Tile_X5Y1_LUT4AB/W2END[7] Tile_X6Y1_LUT4AB/W2END[0]
+ Tile_X6Y1_LUT4AB/W2END[1] Tile_X6Y1_LUT4AB/W2END[2] Tile_X6Y1_LUT4AB/W2END[3] Tile_X6Y1_LUT4AB/W2END[4]
+ Tile_X6Y1_LUT4AB/W2END[5] Tile_X6Y1_LUT4AB/W2END[6] Tile_X6Y1_LUT4AB/W2END[7] Tile_X6Y1_LUT4AB/W2MID[0]
+ Tile_X6Y1_LUT4AB/W2MID[1] Tile_X6Y1_LUT4AB/W2MID[2] Tile_X6Y1_LUT4AB/W2MID[3] Tile_X6Y1_LUT4AB/W2MID[4]
+ Tile_X6Y1_LUT4AB/W2MID[5] Tile_X6Y1_LUT4AB/W2MID[6] Tile_X6Y1_LUT4AB/W2MID[7] Tile_X6Y1_LUT4AB/W6BEG[0]
+ Tile_X6Y1_LUT4AB/W6BEG[10] Tile_X6Y1_LUT4AB/W6BEG[11] Tile_X6Y1_LUT4AB/W6BEG[1]
+ Tile_X6Y1_LUT4AB/W6BEG[2] Tile_X6Y1_LUT4AB/W6BEG[3] Tile_X6Y1_LUT4AB/W6BEG[4] Tile_X6Y1_LUT4AB/W6BEG[5]
+ Tile_X6Y1_LUT4AB/W6BEG[6] Tile_X6Y1_LUT4AB/W6BEG[7] Tile_X6Y1_LUT4AB/W6BEG[8] Tile_X6Y1_LUT4AB/W6BEG[9]
+ Tile_X6Y1_LUT4AB/W6END[0] Tile_X6Y1_LUT4AB/W6END[10] Tile_X6Y1_LUT4AB/W6END[11]
+ Tile_X6Y1_LUT4AB/W6END[1] Tile_X6Y1_LUT4AB/W6END[2] Tile_X6Y1_LUT4AB/W6END[3] Tile_X6Y1_LUT4AB/W6END[4]
+ Tile_X6Y1_LUT4AB/W6END[5] Tile_X6Y1_LUT4AB/W6END[6] Tile_X6Y1_LUT4AB/W6END[7] Tile_X6Y1_LUT4AB/W6END[8]
+ Tile_X6Y1_LUT4AB/W6END[9] Tile_X6Y1_LUT4AB/WW4BEG[0] Tile_X6Y1_LUT4AB/WW4BEG[10]
+ Tile_X6Y1_LUT4AB/WW4BEG[11] Tile_X6Y1_LUT4AB/WW4BEG[12] Tile_X6Y1_LUT4AB/WW4BEG[13]
+ Tile_X6Y1_LUT4AB/WW4BEG[14] Tile_X6Y1_LUT4AB/WW4BEG[15] Tile_X6Y1_LUT4AB/WW4BEG[1]
+ Tile_X6Y1_LUT4AB/WW4BEG[2] Tile_X6Y1_LUT4AB/WW4BEG[3] Tile_X6Y1_LUT4AB/WW4BEG[4]
+ Tile_X6Y1_LUT4AB/WW4BEG[5] Tile_X6Y1_LUT4AB/WW4BEG[6] Tile_X6Y1_LUT4AB/WW4BEG[7]
+ Tile_X6Y1_LUT4AB/WW4BEG[8] Tile_X6Y1_LUT4AB/WW4BEG[9] Tile_X6Y1_LUT4AB/WW4END[0]
+ Tile_X6Y1_LUT4AB/WW4END[10] Tile_X6Y1_LUT4AB/WW4END[11] Tile_X6Y1_LUT4AB/WW4END[12]
+ Tile_X6Y1_LUT4AB/WW4END[13] Tile_X6Y1_LUT4AB/WW4END[14] Tile_X6Y1_LUT4AB/WW4END[15]
+ Tile_X6Y1_LUT4AB/WW4END[1] Tile_X6Y1_LUT4AB/WW4END[2] Tile_X6Y1_LUT4AB/WW4END[3]
+ Tile_X6Y1_LUT4AB/WW4END[4] Tile_X6Y1_LUT4AB/WW4END[5] Tile_X6Y1_LUT4AB/WW4END[6]
+ Tile_X6Y1_LUT4AB/WW4END[7] Tile_X6Y1_LUT4AB/WW4END[8] Tile_X6Y1_LUT4AB/WW4END[9]
+ LUT4AB
XTile_X9Y6_LUT4AB Tile_X9Y7_LUT4AB/Co Tile_X9Y6_LUT4AB/Co Tile_X9Y6_LUT4AB/E1BEG[0]
+ Tile_X9Y6_LUT4AB/E1BEG[1] Tile_X9Y6_LUT4AB/E1BEG[2] Tile_X9Y6_LUT4AB/E1BEG[3] Tile_X9Y6_LUT4AB/E1END[0]
+ Tile_X9Y6_LUT4AB/E1END[1] Tile_X9Y6_LUT4AB/E1END[2] Tile_X9Y6_LUT4AB/E1END[3] Tile_X9Y6_LUT4AB/E2BEG[0]
+ Tile_X9Y6_LUT4AB/E2BEG[1] Tile_X9Y6_LUT4AB/E2BEG[2] Tile_X9Y6_LUT4AB/E2BEG[3] Tile_X9Y6_LUT4AB/E2BEG[4]
+ Tile_X9Y6_LUT4AB/E2BEG[5] Tile_X9Y6_LUT4AB/E2BEG[6] Tile_X9Y6_LUT4AB/E2BEG[7] Tile_X9Y6_LUT4AB/E2BEGb[0]
+ Tile_X9Y6_LUT4AB/E2BEGb[1] Tile_X9Y6_LUT4AB/E2BEGb[2] Tile_X9Y6_LUT4AB/E2BEGb[3]
+ Tile_X9Y6_LUT4AB/E2BEGb[4] Tile_X9Y6_LUT4AB/E2BEGb[5] Tile_X9Y6_LUT4AB/E2BEGb[6]
+ Tile_X9Y6_LUT4AB/E2BEGb[7] Tile_X9Y6_LUT4AB/E2END[0] Tile_X9Y6_LUT4AB/E2END[1] Tile_X9Y6_LUT4AB/E2END[2]
+ Tile_X9Y6_LUT4AB/E2END[3] Tile_X9Y6_LUT4AB/E2END[4] Tile_X9Y6_LUT4AB/E2END[5] Tile_X9Y6_LUT4AB/E2END[6]
+ Tile_X9Y6_LUT4AB/E2END[7] Tile_X9Y6_LUT4AB/E2MID[0] Tile_X9Y6_LUT4AB/E2MID[1] Tile_X9Y6_LUT4AB/E2MID[2]
+ Tile_X9Y6_LUT4AB/E2MID[3] Tile_X9Y6_LUT4AB/E2MID[4] Tile_X9Y6_LUT4AB/E2MID[5] Tile_X9Y6_LUT4AB/E2MID[6]
+ Tile_X9Y6_LUT4AB/E2MID[7] Tile_X9Y6_LUT4AB/E6BEG[0] Tile_X9Y6_LUT4AB/E6BEG[10] Tile_X9Y6_LUT4AB/E6BEG[11]
+ Tile_X9Y6_LUT4AB/E6BEG[1] Tile_X9Y6_LUT4AB/E6BEG[2] Tile_X9Y6_LUT4AB/E6BEG[3] Tile_X9Y6_LUT4AB/E6BEG[4]
+ Tile_X9Y6_LUT4AB/E6BEG[5] Tile_X9Y6_LUT4AB/E6BEG[6] Tile_X9Y6_LUT4AB/E6BEG[7] Tile_X9Y6_LUT4AB/E6BEG[8]
+ Tile_X9Y6_LUT4AB/E6BEG[9] Tile_X9Y6_LUT4AB/E6END[0] Tile_X9Y6_LUT4AB/E6END[10] Tile_X9Y6_LUT4AB/E6END[11]
+ Tile_X9Y6_LUT4AB/E6END[1] Tile_X9Y6_LUT4AB/E6END[2] Tile_X9Y6_LUT4AB/E6END[3] Tile_X9Y6_LUT4AB/E6END[4]
+ Tile_X9Y6_LUT4AB/E6END[5] Tile_X9Y6_LUT4AB/E6END[6] Tile_X9Y6_LUT4AB/E6END[7] Tile_X9Y6_LUT4AB/E6END[8]
+ Tile_X9Y6_LUT4AB/E6END[9] Tile_X9Y6_LUT4AB/EE4BEG[0] Tile_X9Y6_LUT4AB/EE4BEG[10]
+ Tile_X9Y6_LUT4AB/EE4BEG[11] Tile_X9Y6_LUT4AB/EE4BEG[12] Tile_X9Y6_LUT4AB/EE4BEG[13]
+ Tile_X9Y6_LUT4AB/EE4BEG[14] Tile_X9Y6_LUT4AB/EE4BEG[15] Tile_X9Y6_LUT4AB/EE4BEG[1]
+ Tile_X9Y6_LUT4AB/EE4BEG[2] Tile_X9Y6_LUT4AB/EE4BEG[3] Tile_X9Y6_LUT4AB/EE4BEG[4]
+ Tile_X9Y6_LUT4AB/EE4BEG[5] Tile_X9Y6_LUT4AB/EE4BEG[6] Tile_X9Y6_LUT4AB/EE4BEG[7]
+ Tile_X9Y6_LUT4AB/EE4BEG[8] Tile_X9Y6_LUT4AB/EE4BEG[9] Tile_X9Y6_LUT4AB/EE4END[0]
+ Tile_X9Y6_LUT4AB/EE4END[10] Tile_X9Y6_LUT4AB/EE4END[11] Tile_X9Y6_LUT4AB/EE4END[12]
+ Tile_X9Y6_LUT4AB/EE4END[13] Tile_X9Y6_LUT4AB/EE4END[14] Tile_X9Y6_LUT4AB/EE4END[15]
+ Tile_X9Y6_LUT4AB/EE4END[1] Tile_X9Y6_LUT4AB/EE4END[2] Tile_X9Y6_LUT4AB/EE4END[3]
+ Tile_X9Y6_LUT4AB/EE4END[4] Tile_X9Y6_LUT4AB/EE4END[5] Tile_X9Y6_LUT4AB/EE4END[6]
+ Tile_X9Y6_LUT4AB/EE4END[7] Tile_X9Y6_LUT4AB/EE4END[8] Tile_X9Y6_LUT4AB/EE4END[9]
+ Tile_X9Y6_LUT4AB/FrameData[0] Tile_X9Y6_LUT4AB/FrameData[10] Tile_X9Y6_LUT4AB/FrameData[11]
+ Tile_X9Y6_LUT4AB/FrameData[12] Tile_X9Y6_LUT4AB/FrameData[13] Tile_X9Y6_LUT4AB/FrameData[14]
+ Tile_X9Y6_LUT4AB/FrameData[15] Tile_X9Y6_LUT4AB/FrameData[16] Tile_X9Y6_LUT4AB/FrameData[17]
+ Tile_X9Y6_LUT4AB/FrameData[18] Tile_X9Y6_LUT4AB/FrameData[19] Tile_X9Y6_LUT4AB/FrameData[1]
+ Tile_X9Y6_LUT4AB/FrameData[20] Tile_X9Y6_LUT4AB/FrameData[21] Tile_X9Y6_LUT4AB/FrameData[22]
+ Tile_X9Y6_LUT4AB/FrameData[23] Tile_X9Y6_LUT4AB/FrameData[24] Tile_X9Y6_LUT4AB/FrameData[25]
+ Tile_X9Y6_LUT4AB/FrameData[26] Tile_X9Y6_LUT4AB/FrameData[27] Tile_X9Y6_LUT4AB/FrameData[28]
+ Tile_X9Y6_LUT4AB/FrameData[29] Tile_X9Y6_LUT4AB/FrameData[2] Tile_X9Y6_LUT4AB/FrameData[30]
+ Tile_X9Y6_LUT4AB/FrameData[31] Tile_X9Y6_LUT4AB/FrameData[3] Tile_X9Y6_LUT4AB/FrameData[4]
+ Tile_X9Y6_LUT4AB/FrameData[5] Tile_X9Y6_LUT4AB/FrameData[6] Tile_X9Y6_LUT4AB/FrameData[7]
+ Tile_X9Y6_LUT4AB/FrameData[8] Tile_X9Y6_LUT4AB/FrameData[9] Tile_X9Y6_LUT4AB/FrameData_O[0]
+ Tile_X9Y6_LUT4AB/FrameData_O[10] Tile_X9Y6_LUT4AB/FrameData_O[11] Tile_X9Y6_LUT4AB/FrameData_O[12]
+ Tile_X9Y6_LUT4AB/FrameData_O[13] Tile_X9Y6_LUT4AB/FrameData_O[14] Tile_X9Y6_LUT4AB/FrameData_O[15]
+ Tile_X9Y6_LUT4AB/FrameData_O[16] Tile_X9Y6_LUT4AB/FrameData_O[17] Tile_X9Y6_LUT4AB/FrameData_O[18]
+ Tile_X9Y6_LUT4AB/FrameData_O[19] Tile_X9Y6_LUT4AB/FrameData_O[1] Tile_X9Y6_LUT4AB/FrameData_O[20]
+ Tile_X9Y6_LUT4AB/FrameData_O[21] Tile_X9Y6_LUT4AB/FrameData_O[22] Tile_X9Y6_LUT4AB/FrameData_O[23]
+ Tile_X9Y6_LUT4AB/FrameData_O[24] Tile_X9Y6_LUT4AB/FrameData_O[25] Tile_X9Y6_LUT4AB/FrameData_O[26]
+ Tile_X9Y6_LUT4AB/FrameData_O[27] Tile_X9Y6_LUT4AB/FrameData_O[28] Tile_X9Y6_LUT4AB/FrameData_O[29]
+ Tile_X9Y6_LUT4AB/FrameData_O[2] Tile_X9Y6_LUT4AB/FrameData_O[30] Tile_X9Y6_LUT4AB/FrameData_O[31]
+ Tile_X9Y6_LUT4AB/FrameData_O[3] Tile_X9Y6_LUT4AB/FrameData_O[4] Tile_X9Y6_LUT4AB/FrameData_O[5]
+ Tile_X9Y6_LUT4AB/FrameData_O[6] Tile_X9Y6_LUT4AB/FrameData_O[7] Tile_X9Y6_LUT4AB/FrameData_O[8]
+ Tile_X9Y6_LUT4AB/FrameData_O[9] Tile_X9Y6_LUT4AB/FrameStrobe[0] Tile_X9Y6_LUT4AB/FrameStrobe[10]
+ Tile_X9Y6_LUT4AB/FrameStrobe[11] Tile_X9Y6_LUT4AB/FrameStrobe[12] Tile_X9Y6_LUT4AB/FrameStrobe[13]
+ Tile_X9Y6_LUT4AB/FrameStrobe[14] Tile_X9Y6_LUT4AB/FrameStrobe[15] Tile_X9Y6_LUT4AB/FrameStrobe[16]
+ Tile_X9Y6_LUT4AB/FrameStrobe[17] Tile_X9Y6_LUT4AB/FrameStrobe[18] Tile_X9Y6_LUT4AB/FrameStrobe[19]
+ Tile_X9Y6_LUT4AB/FrameStrobe[1] Tile_X9Y6_LUT4AB/FrameStrobe[2] Tile_X9Y6_LUT4AB/FrameStrobe[3]
+ Tile_X9Y6_LUT4AB/FrameStrobe[4] Tile_X9Y6_LUT4AB/FrameStrobe[5] Tile_X9Y6_LUT4AB/FrameStrobe[6]
+ Tile_X9Y6_LUT4AB/FrameStrobe[7] Tile_X9Y6_LUT4AB/FrameStrobe[8] Tile_X9Y6_LUT4AB/FrameStrobe[9]
+ Tile_X9Y5_LUT4AB/FrameStrobe[0] Tile_X9Y5_LUT4AB/FrameStrobe[10] Tile_X9Y5_LUT4AB/FrameStrobe[11]
+ Tile_X9Y5_LUT4AB/FrameStrobe[12] Tile_X9Y5_LUT4AB/FrameStrobe[13] Tile_X9Y5_LUT4AB/FrameStrobe[14]
+ Tile_X9Y5_LUT4AB/FrameStrobe[15] Tile_X9Y5_LUT4AB/FrameStrobe[16] Tile_X9Y5_LUT4AB/FrameStrobe[17]
+ Tile_X9Y5_LUT4AB/FrameStrobe[18] Tile_X9Y5_LUT4AB/FrameStrobe[19] Tile_X9Y5_LUT4AB/FrameStrobe[1]
+ Tile_X9Y5_LUT4AB/FrameStrobe[2] Tile_X9Y5_LUT4AB/FrameStrobe[3] Tile_X9Y5_LUT4AB/FrameStrobe[4]
+ Tile_X9Y5_LUT4AB/FrameStrobe[5] Tile_X9Y5_LUT4AB/FrameStrobe[6] Tile_X9Y5_LUT4AB/FrameStrobe[7]
+ Tile_X9Y5_LUT4AB/FrameStrobe[8] Tile_X9Y5_LUT4AB/FrameStrobe[9] Tile_X9Y6_LUT4AB/N1BEG[0]
+ Tile_X9Y6_LUT4AB/N1BEG[1] Tile_X9Y6_LUT4AB/N1BEG[2] Tile_X9Y6_LUT4AB/N1BEG[3] Tile_X9Y7_LUT4AB/N1BEG[0]
+ Tile_X9Y7_LUT4AB/N1BEG[1] Tile_X9Y7_LUT4AB/N1BEG[2] Tile_X9Y7_LUT4AB/N1BEG[3] Tile_X9Y6_LUT4AB/N2BEG[0]
+ Tile_X9Y6_LUT4AB/N2BEG[1] Tile_X9Y6_LUT4AB/N2BEG[2] Tile_X9Y6_LUT4AB/N2BEG[3] Tile_X9Y6_LUT4AB/N2BEG[4]
+ Tile_X9Y6_LUT4AB/N2BEG[5] Tile_X9Y6_LUT4AB/N2BEG[6] Tile_X9Y6_LUT4AB/N2BEG[7] Tile_X9Y5_LUT4AB/N2END[0]
+ Tile_X9Y5_LUT4AB/N2END[1] Tile_X9Y5_LUT4AB/N2END[2] Tile_X9Y5_LUT4AB/N2END[3] Tile_X9Y5_LUT4AB/N2END[4]
+ Tile_X9Y5_LUT4AB/N2END[5] Tile_X9Y5_LUT4AB/N2END[6] Tile_X9Y5_LUT4AB/N2END[7] Tile_X9Y6_LUT4AB/N2END[0]
+ Tile_X9Y6_LUT4AB/N2END[1] Tile_X9Y6_LUT4AB/N2END[2] Tile_X9Y6_LUT4AB/N2END[3] Tile_X9Y6_LUT4AB/N2END[4]
+ Tile_X9Y6_LUT4AB/N2END[5] Tile_X9Y6_LUT4AB/N2END[6] Tile_X9Y6_LUT4AB/N2END[7] Tile_X9Y7_LUT4AB/N2BEG[0]
+ Tile_X9Y7_LUT4AB/N2BEG[1] Tile_X9Y7_LUT4AB/N2BEG[2] Tile_X9Y7_LUT4AB/N2BEG[3] Tile_X9Y7_LUT4AB/N2BEG[4]
+ Tile_X9Y7_LUT4AB/N2BEG[5] Tile_X9Y7_LUT4AB/N2BEG[6] Tile_X9Y7_LUT4AB/N2BEG[7] Tile_X9Y6_LUT4AB/N4BEG[0]
+ Tile_X9Y6_LUT4AB/N4BEG[10] Tile_X9Y6_LUT4AB/N4BEG[11] Tile_X9Y6_LUT4AB/N4BEG[12]
+ Tile_X9Y6_LUT4AB/N4BEG[13] Tile_X9Y6_LUT4AB/N4BEG[14] Tile_X9Y6_LUT4AB/N4BEG[15]
+ Tile_X9Y6_LUT4AB/N4BEG[1] Tile_X9Y6_LUT4AB/N4BEG[2] Tile_X9Y6_LUT4AB/N4BEG[3] Tile_X9Y6_LUT4AB/N4BEG[4]
+ Tile_X9Y6_LUT4AB/N4BEG[5] Tile_X9Y6_LUT4AB/N4BEG[6] Tile_X9Y6_LUT4AB/N4BEG[7] Tile_X9Y6_LUT4AB/N4BEG[8]
+ Tile_X9Y6_LUT4AB/N4BEG[9] Tile_X9Y7_LUT4AB/N4BEG[0] Tile_X9Y7_LUT4AB/N4BEG[10] Tile_X9Y7_LUT4AB/N4BEG[11]
+ Tile_X9Y7_LUT4AB/N4BEG[12] Tile_X9Y7_LUT4AB/N4BEG[13] Tile_X9Y7_LUT4AB/N4BEG[14]
+ Tile_X9Y7_LUT4AB/N4BEG[15] Tile_X9Y7_LUT4AB/N4BEG[1] Tile_X9Y7_LUT4AB/N4BEG[2] Tile_X9Y7_LUT4AB/N4BEG[3]
+ Tile_X9Y7_LUT4AB/N4BEG[4] Tile_X9Y7_LUT4AB/N4BEG[5] Tile_X9Y7_LUT4AB/N4BEG[6] Tile_X9Y7_LUT4AB/N4BEG[7]
+ Tile_X9Y7_LUT4AB/N4BEG[8] Tile_X9Y7_LUT4AB/N4BEG[9] Tile_X9Y6_LUT4AB/NN4BEG[0] Tile_X9Y6_LUT4AB/NN4BEG[10]
+ Tile_X9Y6_LUT4AB/NN4BEG[11] Tile_X9Y6_LUT4AB/NN4BEG[12] Tile_X9Y6_LUT4AB/NN4BEG[13]
+ Tile_X9Y6_LUT4AB/NN4BEG[14] Tile_X9Y6_LUT4AB/NN4BEG[15] Tile_X9Y6_LUT4AB/NN4BEG[1]
+ Tile_X9Y6_LUT4AB/NN4BEG[2] Tile_X9Y6_LUT4AB/NN4BEG[3] Tile_X9Y6_LUT4AB/NN4BEG[4]
+ Tile_X9Y6_LUT4AB/NN4BEG[5] Tile_X9Y6_LUT4AB/NN4BEG[6] Tile_X9Y6_LUT4AB/NN4BEG[7]
+ Tile_X9Y6_LUT4AB/NN4BEG[8] Tile_X9Y6_LUT4AB/NN4BEG[9] Tile_X9Y7_LUT4AB/NN4BEG[0]
+ Tile_X9Y7_LUT4AB/NN4BEG[10] Tile_X9Y7_LUT4AB/NN4BEG[11] Tile_X9Y7_LUT4AB/NN4BEG[12]
+ Tile_X9Y7_LUT4AB/NN4BEG[13] Tile_X9Y7_LUT4AB/NN4BEG[14] Tile_X9Y7_LUT4AB/NN4BEG[15]
+ Tile_X9Y7_LUT4AB/NN4BEG[1] Tile_X9Y7_LUT4AB/NN4BEG[2] Tile_X9Y7_LUT4AB/NN4BEG[3]
+ Tile_X9Y7_LUT4AB/NN4BEG[4] Tile_X9Y7_LUT4AB/NN4BEG[5] Tile_X9Y7_LUT4AB/NN4BEG[6]
+ Tile_X9Y7_LUT4AB/NN4BEG[7] Tile_X9Y7_LUT4AB/NN4BEG[8] Tile_X9Y7_LUT4AB/NN4BEG[9]
+ Tile_X9Y7_LUT4AB/S1END[0] Tile_X9Y7_LUT4AB/S1END[1] Tile_X9Y7_LUT4AB/S1END[2] Tile_X9Y7_LUT4AB/S1END[3]
+ Tile_X9Y6_LUT4AB/S1END[0] Tile_X9Y6_LUT4AB/S1END[1] Tile_X9Y6_LUT4AB/S1END[2] Tile_X9Y6_LUT4AB/S1END[3]
+ Tile_X9Y7_LUT4AB/S2MID[0] Tile_X9Y7_LUT4AB/S2MID[1] Tile_X9Y7_LUT4AB/S2MID[2] Tile_X9Y7_LUT4AB/S2MID[3]
+ Tile_X9Y7_LUT4AB/S2MID[4] Tile_X9Y7_LUT4AB/S2MID[5] Tile_X9Y7_LUT4AB/S2MID[6] Tile_X9Y7_LUT4AB/S2MID[7]
+ Tile_X9Y7_LUT4AB/S2END[0] Tile_X9Y7_LUT4AB/S2END[1] Tile_X9Y7_LUT4AB/S2END[2] Tile_X9Y7_LUT4AB/S2END[3]
+ Tile_X9Y7_LUT4AB/S2END[4] Tile_X9Y7_LUT4AB/S2END[5] Tile_X9Y7_LUT4AB/S2END[6] Tile_X9Y7_LUT4AB/S2END[7]
+ Tile_X9Y6_LUT4AB/S2END[0] Tile_X9Y6_LUT4AB/S2END[1] Tile_X9Y6_LUT4AB/S2END[2] Tile_X9Y6_LUT4AB/S2END[3]
+ Tile_X9Y6_LUT4AB/S2END[4] Tile_X9Y6_LUT4AB/S2END[5] Tile_X9Y6_LUT4AB/S2END[6] Tile_X9Y6_LUT4AB/S2END[7]
+ Tile_X9Y6_LUT4AB/S2MID[0] Tile_X9Y6_LUT4AB/S2MID[1] Tile_X9Y6_LUT4AB/S2MID[2] Tile_X9Y6_LUT4AB/S2MID[3]
+ Tile_X9Y6_LUT4AB/S2MID[4] Tile_X9Y6_LUT4AB/S2MID[5] Tile_X9Y6_LUT4AB/S2MID[6] Tile_X9Y6_LUT4AB/S2MID[7]
+ Tile_X9Y7_LUT4AB/S4END[0] Tile_X9Y7_LUT4AB/S4END[10] Tile_X9Y7_LUT4AB/S4END[11]
+ Tile_X9Y7_LUT4AB/S4END[12] Tile_X9Y7_LUT4AB/S4END[13] Tile_X9Y7_LUT4AB/S4END[14]
+ Tile_X9Y7_LUT4AB/S4END[15] Tile_X9Y7_LUT4AB/S4END[1] Tile_X9Y7_LUT4AB/S4END[2] Tile_X9Y7_LUT4AB/S4END[3]
+ Tile_X9Y7_LUT4AB/S4END[4] Tile_X9Y7_LUT4AB/S4END[5] Tile_X9Y7_LUT4AB/S4END[6] Tile_X9Y7_LUT4AB/S4END[7]
+ Tile_X9Y7_LUT4AB/S4END[8] Tile_X9Y7_LUT4AB/S4END[9] Tile_X9Y6_LUT4AB/S4END[0] Tile_X9Y6_LUT4AB/S4END[10]
+ Tile_X9Y6_LUT4AB/S4END[11] Tile_X9Y6_LUT4AB/S4END[12] Tile_X9Y6_LUT4AB/S4END[13]
+ Tile_X9Y6_LUT4AB/S4END[14] Tile_X9Y6_LUT4AB/S4END[15] Tile_X9Y6_LUT4AB/S4END[1]
+ Tile_X9Y6_LUT4AB/S4END[2] Tile_X9Y6_LUT4AB/S4END[3] Tile_X9Y6_LUT4AB/S4END[4] Tile_X9Y6_LUT4AB/S4END[5]
+ Tile_X9Y6_LUT4AB/S4END[6] Tile_X9Y6_LUT4AB/S4END[7] Tile_X9Y6_LUT4AB/S4END[8] Tile_X9Y6_LUT4AB/S4END[9]
+ Tile_X9Y7_LUT4AB/SS4END[0] Tile_X9Y7_LUT4AB/SS4END[10] Tile_X9Y7_LUT4AB/SS4END[11]
+ Tile_X9Y7_LUT4AB/SS4END[12] Tile_X9Y7_LUT4AB/SS4END[13] Tile_X9Y7_LUT4AB/SS4END[14]
+ Tile_X9Y7_LUT4AB/SS4END[15] Tile_X9Y7_LUT4AB/SS4END[1] Tile_X9Y7_LUT4AB/SS4END[2]
+ Tile_X9Y7_LUT4AB/SS4END[3] Tile_X9Y7_LUT4AB/SS4END[4] Tile_X9Y7_LUT4AB/SS4END[5]
+ Tile_X9Y7_LUT4AB/SS4END[6] Tile_X9Y7_LUT4AB/SS4END[7] Tile_X9Y7_LUT4AB/SS4END[8]
+ Tile_X9Y7_LUT4AB/SS4END[9] Tile_X9Y6_LUT4AB/SS4END[0] Tile_X9Y6_LUT4AB/SS4END[10]
+ Tile_X9Y6_LUT4AB/SS4END[11] Tile_X9Y6_LUT4AB/SS4END[12] Tile_X9Y6_LUT4AB/SS4END[13]
+ Tile_X9Y6_LUT4AB/SS4END[14] Tile_X9Y6_LUT4AB/SS4END[15] Tile_X9Y6_LUT4AB/SS4END[1]
+ Tile_X9Y6_LUT4AB/SS4END[2] Tile_X9Y6_LUT4AB/SS4END[3] Tile_X9Y6_LUT4AB/SS4END[4]
+ Tile_X9Y6_LUT4AB/SS4END[5] Tile_X9Y6_LUT4AB/SS4END[6] Tile_X9Y6_LUT4AB/SS4END[7]
+ Tile_X9Y6_LUT4AB/SS4END[8] Tile_X9Y6_LUT4AB/SS4END[9] Tile_X9Y6_LUT4AB/UserCLK Tile_X9Y5_LUT4AB/UserCLK
+ VGND VPWR Tile_X9Y6_LUT4AB/W1BEG[0] Tile_X9Y6_LUT4AB/W1BEG[1] Tile_X9Y6_LUT4AB/W1BEG[2]
+ Tile_X9Y6_LUT4AB/W1BEG[3] Tile_X9Y6_LUT4AB/W1END[0] Tile_X9Y6_LUT4AB/W1END[1] Tile_X9Y6_LUT4AB/W1END[2]
+ Tile_X9Y6_LUT4AB/W1END[3] Tile_X9Y6_LUT4AB/W2BEG[0] Tile_X9Y6_LUT4AB/W2BEG[1] Tile_X9Y6_LUT4AB/W2BEG[2]
+ Tile_X9Y6_LUT4AB/W2BEG[3] Tile_X9Y6_LUT4AB/W2BEG[4] Tile_X9Y6_LUT4AB/W2BEG[5] Tile_X9Y6_LUT4AB/W2BEG[6]
+ Tile_X9Y6_LUT4AB/W2BEG[7] Tile_X8Y6_LUT4AB/W2END[0] Tile_X8Y6_LUT4AB/W2END[1] Tile_X8Y6_LUT4AB/W2END[2]
+ Tile_X8Y6_LUT4AB/W2END[3] Tile_X8Y6_LUT4AB/W2END[4] Tile_X8Y6_LUT4AB/W2END[5] Tile_X8Y6_LUT4AB/W2END[6]
+ Tile_X8Y6_LUT4AB/W2END[7] Tile_X9Y6_LUT4AB/W2END[0] Tile_X9Y6_LUT4AB/W2END[1] Tile_X9Y6_LUT4AB/W2END[2]
+ Tile_X9Y6_LUT4AB/W2END[3] Tile_X9Y6_LUT4AB/W2END[4] Tile_X9Y6_LUT4AB/W2END[5] Tile_X9Y6_LUT4AB/W2END[6]
+ Tile_X9Y6_LUT4AB/W2END[7] Tile_X9Y6_LUT4AB/W2MID[0] Tile_X9Y6_LUT4AB/W2MID[1] Tile_X9Y6_LUT4AB/W2MID[2]
+ Tile_X9Y6_LUT4AB/W2MID[3] Tile_X9Y6_LUT4AB/W2MID[4] Tile_X9Y6_LUT4AB/W2MID[5] Tile_X9Y6_LUT4AB/W2MID[6]
+ Tile_X9Y6_LUT4AB/W2MID[7] Tile_X9Y6_LUT4AB/W6BEG[0] Tile_X9Y6_LUT4AB/W6BEG[10] Tile_X9Y6_LUT4AB/W6BEG[11]
+ Tile_X9Y6_LUT4AB/W6BEG[1] Tile_X9Y6_LUT4AB/W6BEG[2] Tile_X9Y6_LUT4AB/W6BEG[3] Tile_X9Y6_LUT4AB/W6BEG[4]
+ Tile_X9Y6_LUT4AB/W6BEG[5] Tile_X9Y6_LUT4AB/W6BEG[6] Tile_X9Y6_LUT4AB/W6BEG[7] Tile_X9Y6_LUT4AB/W6BEG[8]
+ Tile_X9Y6_LUT4AB/W6BEG[9] Tile_X9Y6_LUT4AB/W6END[0] Tile_X9Y6_LUT4AB/W6END[10] Tile_X9Y6_LUT4AB/W6END[11]
+ Tile_X9Y6_LUT4AB/W6END[1] Tile_X9Y6_LUT4AB/W6END[2] Tile_X9Y6_LUT4AB/W6END[3] Tile_X9Y6_LUT4AB/W6END[4]
+ Tile_X9Y6_LUT4AB/W6END[5] Tile_X9Y6_LUT4AB/W6END[6] Tile_X9Y6_LUT4AB/W6END[7] Tile_X9Y6_LUT4AB/W6END[8]
+ Tile_X9Y6_LUT4AB/W6END[9] Tile_X9Y6_LUT4AB/WW4BEG[0] Tile_X9Y6_LUT4AB/WW4BEG[10]
+ Tile_X9Y6_LUT4AB/WW4BEG[11] Tile_X9Y6_LUT4AB/WW4BEG[12] Tile_X9Y6_LUT4AB/WW4BEG[13]
+ Tile_X9Y6_LUT4AB/WW4BEG[14] Tile_X9Y6_LUT4AB/WW4BEG[15] Tile_X9Y6_LUT4AB/WW4BEG[1]
+ Tile_X9Y6_LUT4AB/WW4BEG[2] Tile_X9Y6_LUT4AB/WW4BEG[3] Tile_X9Y6_LUT4AB/WW4BEG[4]
+ Tile_X9Y6_LUT4AB/WW4BEG[5] Tile_X9Y6_LUT4AB/WW4BEG[6] Tile_X9Y6_LUT4AB/WW4BEG[7]
+ Tile_X9Y6_LUT4AB/WW4BEG[8] Tile_X9Y6_LUT4AB/WW4BEG[9] Tile_X9Y6_LUT4AB/WW4END[0]
+ Tile_X9Y6_LUT4AB/WW4END[10] Tile_X9Y6_LUT4AB/WW4END[11] Tile_X9Y6_LUT4AB/WW4END[12]
+ Tile_X9Y6_LUT4AB/WW4END[13] Tile_X9Y6_LUT4AB/WW4END[14] Tile_X9Y6_LUT4AB/WW4END[15]
+ Tile_X9Y6_LUT4AB/WW4END[1] Tile_X9Y6_LUT4AB/WW4END[2] Tile_X9Y6_LUT4AB/WW4END[3]
+ Tile_X9Y6_LUT4AB/WW4END[4] Tile_X9Y6_LUT4AB/WW4END[5] Tile_X9Y6_LUT4AB/WW4END[6]
+ Tile_X9Y6_LUT4AB/WW4END[7] Tile_X9Y6_LUT4AB/WW4END[8] Tile_X9Y6_LUT4AB/WW4END[9]
+ LUT4AB
XTile_X10Y0_N_term_IHP_SRAM Tile_X9Y0_N_term_single/FrameData_O[0] Tile_X9Y0_N_term_single/FrameData_O[10]
+ Tile_X9Y0_N_term_single/FrameData_O[11] Tile_X9Y0_N_term_single/FrameData_O[12]
+ Tile_X9Y0_N_term_single/FrameData_O[13] Tile_X9Y0_N_term_single/FrameData_O[14]
+ Tile_X9Y0_N_term_single/FrameData_O[15] Tile_X9Y0_N_term_single/FrameData_O[16]
+ Tile_X9Y0_N_term_single/FrameData_O[17] Tile_X9Y0_N_term_single/FrameData_O[18]
+ Tile_X9Y0_N_term_single/FrameData_O[19] Tile_X9Y0_N_term_single/FrameData_O[1] Tile_X9Y0_N_term_single/FrameData_O[20]
+ Tile_X9Y0_N_term_single/FrameData_O[21] Tile_X9Y0_N_term_single/FrameData_O[22]
+ Tile_X9Y0_N_term_single/FrameData_O[23] Tile_X9Y0_N_term_single/FrameData_O[24]
+ Tile_X9Y0_N_term_single/FrameData_O[25] Tile_X9Y0_N_term_single/FrameData_O[26]
+ Tile_X9Y0_N_term_single/FrameData_O[27] Tile_X9Y0_N_term_single/FrameData_O[28]
+ Tile_X9Y0_N_term_single/FrameData_O[29] Tile_X9Y0_N_term_single/FrameData_O[2] Tile_X9Y0_N_term_single/FrameData_O[30]
+ Tile_X9Y0_N_term_single/FrameData_O[31] Tile_X9Y0_N_term_single/FrameData_O[3] Tile_X9Y0_N_term_single/FrameData_O[4]
+ Tile_X9Y0_N_term_single/FrameData_O[5] Tile_X9Y0_N_term_single/FrameData_O[6] Tile_X9Y0_N_term_single/FrameData_O[7]
+ Tile_X9Y0_N_term_single/FrameData_O[8] Tile_X9Y0_N_term_single/FrameData_O[9] Tile_X10Y0_N_term_IHP_SRAM/FrameData_O[0]
+ Tile_X10Y0_N_term_IHP_SRAM/FrameData_O[10] Tile_X10Y0_N_term_IHP_SRAM/FrameData_O[11]
+ Tile_X10Y0_N_term_IHP_SRAM/FrameData_O[12] Tile_X10Y0_N_term_IHP_SRAM/FrameData_O[13]
+ Tile_X10Y0_N_term_IHP_SRAM/FrameData_O[14] Tile_X10Y0_N_term_IHP_SRAM/FrameData_O[15]
+ Tile_X10Y0_N_term_IHP_SRAM/FrameData_O[16] Tile_X10Y0_N_term_IHP_SRAM/FrameData_O[17]
+ Tile_X10Y0_N_term_IHP_SRAM/FrameData_O[18] Tile_X10Y0_N_term_IHP_SRAM/FrameData_O[19]
+ Tile_X10Y0_N_term_IHP_SRAM/FrameData_O[1] Tile_X10Y0_N_term_IHP_SRAM/FrameData_O[20]
+ Tile_X10Y0_N_term_IHP_SRAM/FrameData_O[21] Tile_X10Y0_N_term_IHP_SRAM/FrameData_O[22]
+ Tile_X10Y0_N_term_IHP_SRAM/FrameData_O[23] Tile_X10Y0_N_term_IHP_SRAM/FrameData_O[24]
+ Tile_X10Y0_N_term_IHP_SRAM/FrameData_O[25] Tile_X10Y0_N_term_IHP_SRAM/FrameData_O[26]
+ Tile_X10Y0_N_term_IHP_SRAM/FrameData_O[27] Tile_X10Y0_N_term_IHP_SRAM/FrameData_O[28]
+ Tile_X10Y0_N_term_IHP_SRAM/FrameData_O[29] Tile_X10Y0_N_term_IHP_SRAM/FrameData_O[2]
+ Tile_X10Y0_N_term_IHP_SRAM/FrameData_O[30] Tile_X10Y0_N_term_IHP_SRAM/FrameData_O[31]
+ Tile_X10Y0_N_term_IHP_SRAM/FrameData_O[3] Tile_X10Y0_N_term_IHP_SRAM/FrameData_O[4]
+ Tile_X10Y0_N_term_IHP_SRAM/FrameData_O[5] Tile_X10Y0_N_term_IHP_SRAM/FrameData_O[6]
+ Tile_X10Y0_N_term_IHP_SRAM/FrameData_O[7] Tile_X10Y0_N_term_IHP_SRAM/FrameData_O[8]
+ Tile_X10Y0_N_term_IHP_SRAM/FrameData_O[9] Tile_X10Y0_N_term_IHP_SRAM/FrameStrobe[0]
+ Tile_X10Y0_N_term_IHP_SRAM/FrameStrobe[10] Tile_X10Y0_N_term_IHP_SRAM/FrameStrobe[11]
+ Tile_X10Y0_N_term_IHP_SRAM/FrameStrobe[12] Tile_X10Y0_N_term_IHP_SRAM/FrameStrobe[13]
+ Tile_X10Y0_N_term_IHP_SRAM/FrameStrobe[14] Tile_X10Y0_N_term_IHP_SRAM/FrameStrobe[15]
+ Tile_X10Y0_N_term_IHP_SRAM/FrameStrobe[16] Tile_X10Y0_N_term_IHP_SRAM/FrameStrobe[17]
+ Tile_X10Y0_N_term_IHP_SRAM/FrameStrobe[18] Tile_X10Y0_N_term_IHP_SRAM/FrameStrobe[19]
+ Tile_X10Y0_N_term_IHP_SRAM/FrameStrobe[1] Tile_X10Y0_N_term_IHP_SRAM/FrameStrobe[2]
+ Tile_X10Y0_N_term_IHP_SRAM/FrameStrobe[3] Tile_X10Y0_N_term_IHP_SRAM/FrameStrobe[4]
+ Tile_X10Y0_N_term_IHP_SRAM/FrameStrobe[5] Tile_X10Y0_N_term_IHP_SRAM/FrameStrobe[6]
+ Tile_X10Y0_N_term_IHP_SRAM/FrameStrobe[7] Tile_X10Y0_N_term_IHP_SRAM/FrameStrobe[8]
+ Tile_X10Y0_N_term_IHP_SRAM/FrameStrobe[9] Tile_X10Y0_N_term_IHP_SRAM/FrameStrobe_O[0]
+ Tile_X10Y0_N_term_IHP_SRAM/FrameStrobe_O[10] Tile_X10Y0_N_term_IHP_SRAM/FrameStrobe_O[11]
+ Tile_X10Y0_N_term_IHP_SRAM/FrameStrobe_O[12] Tile_X10Y0_N_term_IHP_SRAM/FrameStrobe_O[13]
+ Tile_X10Y0_N_term_IHP_SRAM/FrameStrobe_O[14] Tile_X10Y0_N_term_IHP_SRAM/FrameStrobe_O[15]
+ Tile_X10Y0_N_term_IHP_SRAM/FrameStrobe_O[16] Tile_X10Y0_N_term_IHP_SRAM/FrameStrobe_O[17]
+ Tile_X10Y0_N_term_IHP_SRAM/FrameStrobe_O[18] Tile_X10Y0_N_term_IHP_SRAM/FrameStrobe_O[19]
+ Tile_X10Y0_N_term_IHP_SRAM/FrameStrobe_O[1] Tile_X10Y0_N_term_IHP_SRAM/FrameStrobe_O[2]
+ Tile_X10Y0_N_term_IHP_SRAM/FrameStrobe_O[3] Tile_X10Y0_N_term_IHP_SRAM/FrameStrobe_O[4]
+ Tile_X10Y0_N_term_IHP_SRAM/FrameStrobe_O[5] Tile_X10Y0_N_term_IHP_SRAM/FrameStrobe_O[6]
+ Tile_X10Y0_N_term_IHP_SRAM/FrameStrobe_O[7] Tile_X10Y0_N_term_IHP_SRAM/FrameStrobe_O[8]
+ Tile_X10Y0_N_term_IHP_SRAM/FrameStrobe_O[9] Tile_X10Y0_N_term_IHP_SRAM/N1END[0]
+ Tile_X10Y0_N_term_IHP_SRAM/N1END[1] Tile_X10Y0_N_term_IHP_SRAM/N1END[2] Tile_X10Y0_N_term_IHP_SRAM/N1END[3]
+ Tile_X10Y0_N_term_IHP_SRAM/N2END[0] Tile_X10Y0_N_term_IHP_SRAM/N2END[1] Tile_X10Y0_N_term_IHP_SRAM/N2END[2]
+ Tile_X10Y0_N_term_IHP_SRAM/N2END[3] Tile_X10Y0_N_term_IHP_SRAM/N2END[4] Tile_X10Y0_N_term_IHP_SRAM/N2END[5]
+ Tile_X10Y0_N_term_IHP_SRAM/N2END[6] Tile_X10Y0_N_term_IHP_SRAM/N2END[7] Tile_X10Y0_N_term_IHP_SRAM/N2MID[0]
+ Tile_X10Y0_N_term_IHP_SRAM/N2MID[1] Tile_X10Y0_N_term_IHP_SRAM/N2MID[2] Tile_X10Y0_N_term_IHP_SRAM/N2MID[3]
+ Tile_X10Y0_N_term_IHP_SRAM/N2MID[4] Tile_X10Y0_N_term_IHP_SRAM/N2MID[5] Tile_X10Y0_N_term_IHP_SRAM/N2MID[6]
+ Tile_X10Y0_N_term_IHP_SRAM/N2MID[7] Tile_X10Y0_N_term_IHP_SRAM/N4END[0] Tile_X10Y0_N_term_IHP_SRAM/N4END[10]
+ Tile_X10Y0_N_term_IHP_SRAM/N4END[11] Tile_X10Y0_N_term_IHP_SRAM/N4END[12] Tile_X10Y0_N_term_IHP_SRAM/N4END[13]
+ Tile_X10Y0_N_term_IHP_SRAM/N4END[14] Tile_X10Y0_N_term_IHP_SRAM/N4END[15] Tile_X10Y0_N_term_IHP_SRAM/N4END[1]
+ Tile_X10Y0_N_term_IHP_SRAM/N4END[2] Tile_X10Y0_N_term_IHP_SRAM/N4END[3] Tile_X10Y0_N_term_IHP_SRAM/N4END[4]
+ Tile_X10Y0_N_term_IHP_SRAM/N4END[5] Tile_X10Y0_N_term_IHP_SRAM/N4END[6] Tile_X10Y0_N_term_IHP_SRAM/N4END[7]
+ Tile_X10Y0_N_term_IHP_SRAM/N4END[8] Tile_X10Y0_N_term_IHP_SRAM/N4END[9] Tile_X10Y0_N_term_IHP_SRAM/S1BEG[0]
+ Tile_X10Y0_N_term_IHP_SRAM/S1BEG[1] Tile_X10Y0_N_term_IHP_SRAM/S1BEG[2] Tile_X10Y0_N_term_IHP_SRAM/S1BEG[3]
+ Tile_X10Y0_N_term_IHP_SRAM/S2BEG[0] Tile_X10Y0_N_term_IHP_SRAM/S2BEG[1] Tile_X10Y0_N_term_IHP_SRAM/S2BEG[2]
+ Tile_X10Y0_N_term_IHP_SRAM/S2BEG[3] Tile_X10Y0_N_term_IHP_SRAM/S2BEG[4] Tile_X10Y0_N_term_IHP_SRAM/S2BEG[5]
+ Tile_X10Y0_N_term_IHP_SRAM/S2BEG[6] Tile_X10Y0_N_term_IHP_SRAM/S2BEG[7] Tile_X10Y0_N_term_IHP_SRAM/S2BEGb[0]
+ Tile_X10Y0_N_term_IHP_SRAM/S2BEGb[1] Tile_X10Y0_N_term_IHP_SRAM/S2BEGb[2] Tile_X10Y0_N_term_IHP_SRAM/S2BEGb[3]
+ Tile_X10Y0_N_term_IHP_SRAM/S2BEGb[4] Tile_X10Y0_N_term_IHP_SRAM/S2BEGb[5] Tile_X10Y0_N_term_IHP_SRAM/S2BEGb[6]
+ Tile_X10Y0_N_term_IHP_SRAM/S2BEGb[7] Tile_X10Y0_N_term_IHP_SRAM/S4BEG[0] Tile_X10Y0_N_term_IHP_SRAM/S4BEG[10]
+ Tile_X10Y0_N_term_IHP_SRAM/S4BEG[11] Tile_X10Y0_N_term_IHP_SRAM/S4BEG[12] Tile_X10Y0_N_term_IHP_SRAM/S4BEG[13]
+ Tile_X10Y0_N_term_IHP_SRAM/S4BEG[14] Tile_X10Y0_N_term_IHP_SRAM/S4BEG[15] Tile_X10Y0_N_term_IHP_SRAM/S4BEG[1]
+ Tile_X10Y0_N_term_IHP_SRAM/S4BEG[2] Tile_X10Y0_N_term_IHP_SRAM/S4BEG[3] Tile_X10Y0_N_term_IHP_SRAM/S4BEG[4]
+ Tile_X10Y0_N_term_IHP_SRAM/S4BEG[5] Tile_X10Y0_N_term_IHP_SRAM/S4BEG[6] Tile_X10Y0_N_term_IHP_SRAM/S4BEG[7]
+ Tile_X10Y0_N_term_IHP_SRAM/S4BEG[8] Tile_X10Y0_N_term_IHP_SRAM/S4BEG[9] Tile_X10Y0_N_term_IHP_SRAM/UserCLK
+ Tile_X10Y0_N_term_IHP_SRAM/UserCLKo VGND VPWR N_term_IHP_SRAM
XTile_X2Y13_LUT4AB Tile_X2Y14_LUT4AB/Co Tile_X2Y13_LUT4AB/Co Tile_X3Y13_LUT4AB/E1END[0]
+ Tile_X3Y13_LUT4AB/E1END[1] Tile_X3Y13_LUT4AB/E1END[2] Tile_X3Y13_LUT4AB/E1END[3]
+ Tile_X2Y13_LUT4AB/E1END[0] Tile_X2Y13_LUT4AB/E1END[1] Tile_X2Y13_LUT4AB/E1END[2]
+ Tile_X2Y13_LUT4AB/E1END[3] Tile_X3Y13_LUT4AB/E2MID[0] Tile_X3Y13_LUT4AB/E2MID[1]
+ Tile_X3Y13_LUT4AB/E2MID[2] Tile_X3Y13_LUT4AB/E2MID[3] Tile_X3Y13_LUT4AB/E2MID[4]
+ Tile_X3Y13_LUT4AB/E2MID[5] Tile_X3Y13_LUT4AB/E2MID[6] Tile_X3Y13_LUT4AB/E2MID[7]
+ Tile_X3Y13_LUT4AB/E2END[0] Tile_X3Y13_LUT4AB/E2END[1] Tile_X3Y13_LUT4AB/E2END[2]
+ Tile_X3Y13_LUT4AB/E2END[3] Tile_X3Y13_LUT4AB/E2END[4] Tile_X3Y13_LUT4AB/E2END[5]
+ Tile_X3Y13_LUT4AB/E2END[6] Tile_X3Y13_LUT4AB/E2END[7] Tile_X2Y13_LUT4AB/E2END[0]
+ Tile_X2Y13_LUT4AB/E2END[1] Tile_X2Y13_LUT4AB/E2END[2] Tile_X2Y13_LUT4AB/E2END[3]
+ Tile_X2Y13_LUT4AB/E2END[4] Tile_X2Y13_LUT4AB/E2END[5] Tile_X2Y13_LUT4AB/E2END[6]
+ Tile_X2Y13_LUT4AB/E2END[7] Tile_X2Y13_LUT4AB/E2MID[0] Tile_X2Y13_LUT4AB/E2MID[1]
+ Tile_X2Y13_LUT4AB/E2MID[2] Tile_X2Y13_LUT4AB/E2MID[3] Tile_X2Y13_LUT4AB/E2MID[4]
+ Tile_X2Y13_LUT4AB/E2MID[5] Tile_X2Y13_LUT4AB/E2MID[6] Tile_X2Y13_LUT4AB/E2MID[7]
+ Tile_X3Y13_LUT4AB/E6END[0] Tile_X3Y13_LUT4AB/E6END[10] Tile_X3Y13_LUT4AB/E6END[11]
+ Tile_X3Y13_LUT4AB/E6END[1] Tile_X3Y13_LUT4AB/E6END[2] Tile_X3Y13_LUT4AB/E6END[3]
+ Tile_X3Y13_LUT4AB/E6END[4] Tile_X3Y13_LUT4AB/E6END[5] Tile_X3Y13_LUT4AB/E6END[6]
+ Tile_X3Y13_LUT4AB/E6END[7] Tile_X3Y13_LUT4AB/E6END[8] Tile_X3Y13_LUT4AB/E6END[9]
+ Tile_X2Y13_LUT4AB/E6END[0] Tile_X2Y13_LUT4AB/E6END[10] Tile_X2Y13_LUT4AB/E6END[11]
+ Tile_X2Y13_LUT4AB/E6END[1] Tile_X2Y13_LUT4AB/E6END[2] Tile_X2Y13_LUT4AB/E6END[3]
+ Tile_X2Y13_LUT4AB/E6END[4] Tile_X2Y13_LUT4AB/E6END[5] Tile_X2Y13_LUT4AB/E6END[6]
+ Tile_X2Y13_LUT4AB/E6END[7] Tile_X2Y13_LUT4AB/E6END[8] Tile_X2Y13_LUT4AB/E6END[9]
+ Tile_X3Y13_LUT4AB/EE4END[0] Tile_X3Y13_LUT4AB/EE4END[10] Tile_X3Y13_LUT4AB/EE4END[11]
+ Tile_X3Y13_LUT4AB/EE4END[12] Tile_X3Y13_LUT4AB/EE4END[13] Tile_X3Y13_LUT4AB/EE4END[14]
+ Tile_X3Y13_LUT4AB/EE4END[15] Tile_X3Y13_LUT4AB/EE4END[1] Tile_X3Y13_LUT4AB/EE4END[2]
+ Tile_X3Y13_LUT4AB/EE4END[3] Tile_X3Y13_LUT4AB/EE4END[4] Tile_X3Y13_LUT4AB/EE4END[5]
+ Tile_X3Y13_LUT4AB/EE4END[6] Tile_X3Y13_LUT4AB/EE4END[7] Tile_X3Y13_LUT4AB/EE4END[8]
+ Tile_X3Y13_LUT4AB/EE4END[9] Tile_X2Y13_LUT4AB/EE4END[0] Tile_X2Y13_LUT4AB/EE4END[10]
+ Tile_X2Y13_LUT4AB/EE4END[11] Tile_X2Y13_LUT4AB/EE4END[12] Tile_X2Y13_LUT4AB/EE4END[13]
+ Tile_X2Y13_LUT4AB/EE4END[14] Tile_X2Y13_LUT4AB/EE4END[15] Tile_X2Y13_LUT4AB/EE4END[1]
+ Tile_X2Y13_LUT4AB/EE4END[2] Tile_X2Y13_LUT4AB/EE4END[3] Tile_X2Y13_LUT4AB/EE4END[4]
+ Tile_X2Y13_LUT4AB/EE4END[5] Tile_X2Y13_LUT4AB/EE4END[6] Tile_X2Y13_LUT4AB/EE4END[7]
+ Tile_X2Y13_LUT4AB/EE4END[8] Tile_X2Y13_LUT4AB/EE4END[9] Tile_X2Y13_LUT4AB/FrameData[0]
+ Tile_X2Y13_LUT4AB/FrameData[10] Tile_X2Y13_LUT4AB/FrameData[11] Tile_X2Y13_LUT4AB/FrameData[12]
+ Tile_X2Y13_LUT4AB/FrameData[13] Tile_X2Y13_LUT4AB/FrameData[14] Tile_X2Y13_LUT4AB/FrameData[15]
+ Tile_X2Y13_LUT4AB/FrameData[16] Tile_X2Y13_LUT4AB/FrameData[17] Tile_X2Y13_LUT4AB/FrameData[18]
+ Tile_X2Y13_LUT4AB/FrameData[19] Tile_X2Y13_LUT4AB/FrameData[1] Tile_X2Y13_LUT4AB/FrameData[20]
+ Tile_X2Y13_LUT4AB/FrameData[21] Tile_X2Y13_LUT4AB/FrameData[22] Tile_X2Y13_LUT4AB/FrameData[23]
+ Tile_X2Y13_LUT4AB/FrameData[24] Tile_X2Y13_LUT4AB/FrameData[25] Tile_X2Y13_LUT4AB/FrameData[26]
+ Tile_X2Y13_LUT4AB/FrameData[27] Tile_X2Y13_LUT4AB/FrameData[28] Tile_X2Y13_LUT4AB/FrameData[29]
+ Tile_X2Y13_LUT4AB/FrameData[2] Tile_X2Y13_LUT4AB/FrameData[30] Tile_X2Y13_LUT4AB/FrameData[31]
+ Tile_X2Y13_LUT4AB/FrameData[3] Tile_X2Y13_LUT4AB/FrameData[4] Tile_X2Y13_LUT4AB/FrameData[5]
+ Tile_X2Y13_LUT4AB/FrameData[6] Tile_X2Y13_LUT4AB/FrameData[7] Tile_X2Y13_LUT4AB/FrameData[8]
+ Tile_X2Y13_LUT4AB/FrameData[9] Tile_X3Y13_LUT4AB/FrameData[0] Tile_X3Y13_LUT4AB/FrameData[10]
+ Tile_X3Y13_LUT4AB/FrameData[11] Tile_X3Y13_LUT4AB/FrameData[12] Tile_X3Y13_LUT4AB/FrameData[13]
+ Tile_X3Y13_LUT4AB/FrameData[14] Tile_X3Y13_LUT4AB/FrameData[15] Tile_X3Y13_LUT4AB/FrameData[16]
+ Tile_X3Y13_LUT4AB/FrameData[17] Tile_X3Y13_LUT4AB/FrameData[18] Tile_X3Y13_LUT4AB/FrameData[19]
+ Tile_X3Y13_LUT4AB/FrameData[1] Tile_X3Y13_LUT4AB/FrameData[20] Tile_X3Y13_LUT4AB/FrameData[21]
+ Tile_X3Y13_LUT4AB/FrameData[22] Tile_X3Y13_LUT4AB/FrameData[23] Tile_X3Y13_LUT4AB/FrameData[24]
+ Tile_X3Y13_LUT4AB/FrameData[25] Tile_X3Y13_LUT4AB/FrameData[26] Tile_X3Y13_LUT4AB/FrameData[27]
+ Tile_X3Y13_LUT4AB/FrameData[28] Tile_X3Y13_LUT4AB/FrameData[29] Tile_X3Y13_LUT4AB/FrameData[2]
+ Tile_X3Y13_LUT4AB/FrameData[30] Tile_X3Y13_LUT4AB/FrameData[31] Tile_X3Y13_LUT4AB/FrameData[3]
+ Tile_X3Y13_LUT4AB/FrameData[4] Tile_X3Y13_LUT4AB/FrameData[5] Tile_X3Y13_LUT4AB/FrameData[6]
+ Tile_X3Y13_LUT4AB/FrameData[7] Tile_X3Y13_LUT4AB/FrameData[8] Tile_X3Y13_LUT4AB/FrameData[9]
+ Tile_X2Y13_LUT4AB/FrameStrobe[0] Tile_X2Y13_LUT4AB/FrameStrobe[10] Tile_X2Y13_LUT4AB/FrameStrobe[11]
+ Tile_X2Y13_LUT4AB/FrameStrobe[12] Tile_X2Y13_LUT4AB/FrameStrobe[13] Tile_X2Y13_LUT4AB/FrameStrobe[14]
+ Tile_X2Y13_LUT4AB/FrameStrobe[15] Tile_X2Y13_LUT4AB/FrameStrobe[16] Tile_X2Y13_LUT4AB/FrameStrobe[17]
+ Tile_X2Y13_LUT4AB/FrameStrobe[18] Tile_X2Y13_LUT4AB/FrameStrobe[19] Tile_X2Y13_LUT4AB/FrameStrobe[1]
+ Tile_X2Y13_LUT4AB/FrameStrobe[2] Tile_X2Y13_LUT4AB/FrameStrobe[3] Tile_X2Y13_LUT4AB/FrameStrobe[4]
+ Tile_X2Y13_LUT4AB/FrameStrobe[5] Tile_X2Y13_LUT4AB/FrameStrobe[6] Tile_X2Y13_LUT4AB/FrameStrobe[7]
+ Tile_X2Y13_LUT4AB/FrameStrobe[8] Tile_X2Y13_LUT4AB/FrameStrobe[9] Tile_X2Y12_LUT4AB/FrameStrobe[0]
+ Tile_X2Y12_LUT4AB/FrameStrobe[10] Tile_X2Y12_LUT4AB/FrameStrobe[11] Tile_X2Y12_LUT4AB/FrameStrobe[12]
+ Tile_X2Y12_LUT4AB/FrameStrobe[13] Tile_X2Y12_LUT4AB/FrameStrobe[14] Tile_X2Y12_LUT4AB/FrameStrobe[15]
+ Tile_X2Y12_LUT4AB/FrameStrobe[16] Tile_X2Y12_LUT4AB/FrameStrobe[17] Tile_X2Y12_LUT4AB/FrameStrobe[18]
+ Tile_X2Y12_LUT4AB/FrameStrobe[19] Tile_X2Y12_LUT4AB/FrameStrobe[1] Tile_X2Y12_LUT4AB/FrameStrobe[2]
+ Tile_X2Y12_LUT4AB/FrameStrobe[3] Tile_X2Y12_LUT4AB/FrameStrobe[4] Tile_X2Y12_LUT4AB/FrameStrobe[5]
+ Tile_X2Y12_LUT4AB/FrameStrobe[6] Tile_X2Y12_LUT4AB/FrameStrobe[7] Tile_X2Y12_LUT4AB/FrameStrobe[8]
+ Tile_X2Y12_LUT4AB/FrameStrobe[9] Tile_X2Y13_LUT4AB/N1BEG[0] Tile_X2Y13_LUT4AB/N1BEG[1]
+ Tile_X2Y13_LUT4AB/N1BEG[2] Tile_X2Y13_LUT4AB/N1BEG[3] Tile_X2Y14_LUT4AB/N1BEG[0]
+ Tile_X2Y14_LUT4AB/N1BEG[1] Tile_X2Y14_LUT4AB/N1BEG[2] Tile_X2Y14_LUT4AB/N1BEG[3]
+ Tile_X2Y13_LUT4AB/N2BEG[0] Tile_X2Y13_LUT4AB/N2BEG[1] Tile_X2Y13_LUT4AB/N2BEG[2]
+ Tile_X2Y13_LUT4AB/N2BEG[3] Tile_X2Y13_LUT4AB/N2BEG[4] Tile_X2Y13_LUT4AB/N2BEG[5]
+ Tile_X2Y13_LUT4AB/N2BEG[6] Tile_X2Y13_LUT4AB/N2BEG[7] Tile_X2Y12_LUT4AB/N2END[0]
+ Tile_X2Y12_LUT4AB/N2END[1] Tile_X2Y12_LUT4AB/N2END[2] Tile_X2Y12_LUT4AB/N2END[3]
+ Tile_X2Y12_LUT4AB/N2END[4] Tile_X2Y12_LUT4AB/N2END[5] Tile_X2Y12_LUT4AB/N2END[6]
+ Tile_X2Y12_LUT4AB/N2END[7] Tile_X2Y13_LUT4AB/N2END[0] Tile_X2Y13_LUT4AB/N2END[1]
+ Tile_X2Y13_LUT4AB/N2END[2] Tile_X2Y13_LUT4AB/N2END[3] Tile_X2Y13_LUT4AB/N2END[4]
+ Tile_X2Y13_LUT4AB/N2END[5] Tile_X2Y13_LUT4AB/N2END[6] Tile_X2Y13_LUT4AB/N2END[7]
+ Tile_X2Y14_LUT4AB/N2BEG[0] Tile_X2Y14_LUT4AB/N2BEG[1] Tile_X2Y14_LUT4AB/N2BEG[2]
+ Tile_X2Y14_LUT4AB/N2BEG[3] Tile_X2Y14_LUT4AB/N2BEG[4] Tile_X2Y14_LUT4AB/N2BEG[5]
+ Tile_X2Y14_LUT4AB/N2BEG[6] Tile_X2Y14_LUT4AB/N2BEG[7] Tile_X2Y13_LUT4AB/N4BEG[0]
+ Tile_X2Y13_LUT4AB/N4BEG[10] Tile_X2Y13_LUT4AB/N4BEG[11] Tile_X2Y13_LUT4AB/N4BEG[12]
+ Tile_X2Y13_LUT4AB/N4BEG[13] Tile_X2Y13_LUT4AB/N4BEG[14] Tile_X2Y13_LUT4AB/N4BEG[15]
+ Tile_X2Y13_LUT4AB/N4BEG[1] Tile_X2Y13_LUT4AB/N4BEG[2] Tile_X2Y13_LUT4AB/N4BEG[3]
+ Tile_X2Y13_LUT4AB/N4BEG[4] Tile_X2Y13_LUT4AB/N4BEG[5] Tile_X2Y13_LUT4AB/N4BEG[6]
+ Tile_X2Y13_LUT4AB/N4BEG[7] Tile_X2Y13_LUT4AB/N4BEG[8] Tile_X2Y13_LUT4AB/N4BEG[9]
+ Tile_X2Y14_LUT4AB/N4BEG[0] Tile_X2Y14_LUT4AB/N4BEG[10] Tile_X2Y14_LUT4AB/N4BEG[11]
+ Tile_X2Y14_LUT4AB/N4BEG[12] Tile_X2Y14_LUT4AB/N4BEG[13] Tile_X2Y14_LUT4AB/N4BEG[14]
+ Tile_X2Y14_LUT4AB/N4BEG[15] Tile_X2Y14_LUT4AB/N4BEG[1] Tile_X2Y14_LUT4AB/N4BEG[2]
+ Tile_X2Y14_LUT4AB/N4BEG[3] Tile_X2Y14_LUT4AB/N4BEG[4] Tile_X2Y14_LUT4AB/N4BEG[5]
+ Tile_X2Y14_LUT4AB/N4BEG[6] Tile_X2Y14_LUT4AB/N4BEG[7] Tile_X2Y14_LUT4AB/N4BEG[8]
+ Tile_X2Y14_LUT4AB/N4BEG[9] Tile_X2Y13_LUT4AB/NN4BEG[0] Tile_X2Y13_LUT4AB/NN4BEG[10]
+ Tile_X2Y13_LUT4AB/NN4BEG[11] Tile_X2Y13_LUT4AB/NN4BEG[12] Tile_X2Y13_LUT4AB/NN4BEG[13]
+ Tile_X2Y13_LUT4AB/NN4BEG[14] Tile_X2Y13_LUT4AB/NN4BEG[15] Tile_X2Y13_LUT4AB/NN4BEG[1]
+ Tile_X2Y13_LUT4AB/NN4BEG[2] Tile_X2Y13_LUT4AB/NN4BEG[3] Tile_X2Y13_LUT4AB/NN4BEG[4]
+ Tile_X2Y13_LUT4AB/NN4BEG[5] Tile_X2Y13_LUT4AB/NN4BEG[6] Tile_X2Y13_LUT4AB/NN4BEG[7]
+ Tile_X2Y13_LUT4AB/NN4BEG[8] Tile_X2Y13_LUT4AB/NN4BEG[9] Tile_X2Y14_LUT4AB/NN4BEG[0]
+ Tile_X2Y14_LUT4AB/NN4BEG[10] Tile_X2Y14_LUT4AB/NN4BEG[11] Tile_X2Y14_LUT4AB/NN4BEG[12]
+ Tile_X2Y14_LUT4AB/NN4BEG[13] Tile_X2Y14_LUT4AB/NN4BEG[14] Tile_X2Y14_LUT4AB/NN4BEG[15]
+ Tile_X2Y14_LUT4AB/NN4BEG[1] Tile_X2Y14_LUT4AB/NN4BEG[2] Tile_X2Y14_LUT4AB/NN4BEG[3]
+ Tile_X2Y14_LUT4AB/NN4BEG[4] Tile_X2Y14_LUT4AB/NN4BEG[5] Tile_X2Y14_LUT4AB/NN4BEG[6]
+ Tile_X2Y14_LUT4AB/NN4BEG[7] Tile_X2Y14_LUT4AB/NN4BEG[8] Tile_X2Y14_LUT4AB/NN4BEG[9]
+ Tile_X2Y14_LUT4AB/S1END[0] Tile_X2Y14_LUT4AB/S1END[1] Tile_X2Y14_LUT4AB/S1END[2]
+ Tile_X2Y14_LUT4AB/S1END[3] Tile_X2Y13_LUT4AB/S1END[0] Tile_X2Y13_LUT4AB/S1END[1]
+ Tile_X2Y13_LUT4AB/S1END[2] Tile_X2Y13_LUT4AB/S1END[3] Tile_X2Y14_LUT4AB/S2MID[0]
+ Tile_X2Y14_LUT4AB/S2MID[1] Tile_X2Y14_LUT4AB/S2MID[2] Tile_X2Y14_LUT4AB/S2MID[3]
+ Tile_X2Y14_LUT4AB/S2MID[4] Tile_X2Y14_LUT4AB/S2MID[5] Tile_X2Y14_LUT4AB/S2MID[6]
+ Tile_X2Y14_LUT4AB/S2MID[7] Tile_X2Y14_LUT4AB/S2END[0] Tile_X2Y14_LUT4AB/S2END[1]
+ Tile_X2Y14_LUT4AB/S2END[2] Tile_X2Y14_LUT4AB/S2END[3] Tile_X2Y14_LUT4AB/S2END[4]
+ Tile_X2Y14_LUT4AB/S2END[5] Tile_X2Y14_LUT4AB/S2END[6] Tile_X2Y14_LUT4AB/S2END[7]
+ Tile_X2Y13_LUT4AB/S2END[0] Tile_X2Y13_LUT4AB/S2END[1] Tile_X2Y13_LUT4AB/S2END[2]
+ Tile_X2Y13_LUT4AB/S2END[3] Tile_X2Y13_LUT4AB/S2END[4] Tile_X2Y13_LUT4AB/S2END[5]
+ Tile_X2Y13_LUT4AB/S2END[6] Tile_X2Y13_LUT4AB/S2END[7] Tile_X2Y13_LUT4AB/S2MID[0]
+ Tile_X2Y13_LUT4AB/S2MID[1] Tile_X2Y13_LUT4AB/S2MID[2] Tile_X2Y13_LUT4AB/S2MID[3]
+ Tile_X2Y13_LUT4AB/S2MID[4] Tile_X2Y13_LUT4AB/S2MID[5] Tile_X2Y13_LUT4AB/S2MID[6]
+ Tile_X2Y13_LUT4AB/S2MID[7] Tile_X2Y14_LUT4AB/S4END[0] Tile_X2Y14_LUT4AB/S4END[10]
+ Tile_X2Y14_LUT4AB/S4END[11] Tile_X2Y14_LUT4AB/S4END[12] Tile_X2Y14_LUT4AB/S4END[13]
+ Tile_X2Y14_LUT4AB/S4END[14] Tile_X2Y14_LUT4AB/S4END[15] Tile_X2Y14_LUT4AB/S4END[1]
+ Tile_X2Y14_LUT4AB/S4END[2] Tile_X2Y14_LUT4AB/S4END[3] Tile_X2Y14_LUT4AB/S4END[4]
+ Tile_X2Y14_LUT4AB/S4END[5] Tile_X2Y14_LUT4AB/S4END[6] Tile_X2Y14_LUT4AB/S4END[7]
+ Tile_X2Y14_LUT4AB/S4END[8] Tile_X2Y14_LUT4AB/S4END[9] Tile_X2Y13_LUT4AB/S4END[0]
+ Tile_X2Y13_LUT4AB/S4END[10] Tile_X2Y13_LUT4AB/S4END[11] Tile_X2Y13_LUT4AB/S4END[12]
+ Tile_X2Y13_LUT4AB/S4END[13] Tile_X2Y13_LUT4AB/S4END[14] Tile_X2Y13_LUT4AB/S4END[15]
+ Tile_X2Y13_LUT4AB/S4END[1] Tile_X2Y13_LUT4AB/S4END[2] Tile_X2Y13_LUT4AB/S4END[3]
+ Tile_X2Y13_LUT4AB/S4END[4] Tile_X2Y13_LUT4AB/S4END[5] Tile_X2Y13_LUT4AB/S4END[6]
+ Tile_X2Y13_LUT4AB/S4END[7] Tile_X2Y13_LUT4AB/S4END[8] Tile_X2Y13_LUT4AB/S4END[9]
+ Tile_X2Y14_LUT4AB/SS4END[0] Tile_X2Y14_LUT4AB/SS4END[10] Tile_X2Y14_LUT4AB/SS4END[11]
+ Tile_X2Y14_LUT4AB/SS4END[12] Tile_X2Y14_LUT4AB/SS4END[13] Tile_X2Y14_LUT4AB/SS4END[14]
+ Tile_X2Y14_LUT4AB/SS4END[15] Tile_X2Y14_LUT4AB/SS4END[1] Tile_X2Y14_LUT4AB/SS4END[2]
+ Tile_X2Y14_LUT4AB/SS4END[3] Tile_X2Y14_LUT4AB/SS4END[4] Tile_X2Y14_LUT4AB/SS4END[5]
+ Tile_X2Y14_LUT4AB/SS4END[6] Tile_X2Y14_LUT4AB/SS4END[7] Tile_X2Y14_LUT4AB/SS4END[8]
+ Tile_X2Y14_LUT4AB/SS4END[9] Tile_X2Y13_LUT4AB/SS4END[0] Tile_X2Y13_LUT4AB/SS4END[10]
+ Tile_X2Y13_LUT4AB/SS4END[11] Tile_X2Y13_LUT4AB/SS4END[12] Tile_X2Y13_LUT4AB/SS4END[13]
+ Tile_X2Y13_LUT4AB/SS4END[14] Tile_X2Y13_LUT4AB/SS4END[15] Tile_X2Y13_LUT4AB/SS4END[1]
+ Tile_X2Y13_LUT4AB/SS4END[2] Tile_X2Y13_LUT4AB/SS4END[3] Tile_X2Y13_LUT4AB/SS4END[4]
+ Tile_X2Y13_LUT4AB/SS4END[5] Tile_X2Y13_LUT4AB/SS4END[6] Tile_X2Y13_LUT4AB/SS4END[7]
+ Tile_X2Y13_LUT4AB/SS4END[8] Tile_X2Y13_LUT4AB/SS4END[9] Tile_X2Y13_LUT4AB/UserCLK
+ Tile_X2Y12_LUT4AB/UserCLK VGND VPWR Tile_X2Y13_LUT4AB/W1BEG[0] Tile_X2Y13_LUT4AB/W1BEG[1]
+ Tile_X2Y13_LUT4AB/W1BEG[2] Tile_X2Y13_LUT4AB/W1BEG[3] Tile_X3Y13_LUT4AB/W1BEG[0]
+ Tile_X3Y13_LUT4AB/W1BEG[1] Tile_X3Y13_LUT4AB/W1BEG[2] Tile_X3Y13_LUT4AB/W1BEG[3]
+ Tile_X2Y13_LUT4AB/W2BEG[0] Tile_X2Y13_LUT4AB/W2BEG[1] Tile_X2Y13_LUT4AB/W2BEG[2]
+ Tile_X2Y13_LUT4AB/W2BEG[3] Tile_X2Y13_LUT4AB/W2BEG[4] Tile_X2Y13_LUT4AB/W2BEG[5]
+ Tile_X2Y13_LUT4AB/W2BEG[6] Tile_X2Y13_LUT4AB/W2BEG[7] Tile_X1Y13_LUT4AB/W2END[0]
+ Tile_X1Y13_LUT4AB/W2END[1] Tile_X1Y13_LUT4AB/W2END[2] Tile_X1Y13_LUT4AB/W2END[3]
+ Tile_X1Y13_LUT4AB/W2END[4] Tile_X1Y13_LUT4AB/W2END[5] Tile_X1Y13_LUT4AB/W2END[6]
+ Tile_X1Y13_LUT4AB/W2END[7] Tile_X2Y13_LUT4AB/W2END[0] Tile_X2Y13_LUT4AB/W2END[1]
+ Tile_X2Y13_LUT4AB/W2END[2] Tile_X2Y13_LUT4AB/W2END[3] Tile_X2Y13_LUT4AB/W2END[4]
+ Tile_X2Y13_LUT4AB/W2END[5] Tile_X2Y13_LUT4AB/W2END[6] Tile_X2Y13_LUT4AB/W2END[7]
+ Tile_X3Y13_LUT4AB/W2BEG[0] Tile_X3Y13_LUT4AB/W2BEG[1] Tile_X3Y13_LUT4AB/W2BEG[2]
+ Tile_X3Y13_LUT4AB/W2BEG[3] Tile_X3Y13_LUT4AB/W2BEG[4] Tile_X3Y13_LUT4AB/W2BEG[5]
+ Tile_X3Y13_LUT4AB/W2BEG[6] Tile_X3Y13_LUT4AB/W2BEG[7] Tile_X2Y13_LUT4AB/W6BEG[0]
+ Tile_X2Y13_LUT4AB/W6BEG[10] Tile_X2Y13_LUT4AB/W6BEG[11] Tile_X2Y13_LUT4AB/W6BEG[1]
+ Tile_X2Y13_LUT4AB/W6BEG[2] Tile_X2Y13_LUT4AB/W6BEG[3] Tile_X2Y13_LUT4AB/W6BEG[4]
+ Tile_X2Y13_LUT4AB/W6BEG[5] Tile_X2Y13_LUT4AB/W6BEG[6] Tile_X2Y13_LUT4AB/W6BEG[7]
+ Tile_X2Y13_LUT4AB/W6BEG[8] Tile_X2Y13_LUT4AB/W6BEG[9] Tile_X3Y13_LUT4AB/W6BEG[0]
+ Tile_X3Y13_LUT4AB/W6BEG[10] Tile_X3Y13_LUT4AB/W6BEG[11] Tile_X3Y13_LUT4AB/W6BEG[1]
+ Tile_X3Y13_LUT4AB/W6BEG[2] Tile_X3Y13_LUT4AB/W6BEG[3] Tile_X3Y13_LUT4AB/W6BEG[4]
+ Tile_X3Y13_LUT4AB/W6BEG[5] Tile_X3Y13_LUT4AB/W6BEG[6] Tile_X3Y13_LUT4AB/W6BEG[7]
+ Tile_X3Y13_LUT4AB/W6BEG[8] Tile_X3Y13_LUT4AB/W6BEG[9] Tile_X2Y13_LUT4AB/WW4BEG[0]
+ Tile_X2Y13_LUT4AB/WW4BEG[10] Tile_X2Y13_LUT4AB/WW4BEG[11] Tile_X2Y13_LUT4AB/WW4BEG[12]
+ Tile_X2Y13_LUT4AB/WW4BEG[13] Tile_X2Y13_LUT4AB/WW4BEG[14] Tile_X2Y13_LUT4AB/WW4BEG[15]
+ Tile_X2Y13_LUT4AB/WW4BEG[1] Tile_X2Y13_LUT4AB/WW4BEG[2] Tile_X2Y13_LUT4AB/WW4BEG[3]
+ Tile_X2Y13_LUT4AB/WW4BEG[4] Tile_X2Y13_LUT4AB/WW4BEG[5] Tile_X2Y13_LUT4AB/WW4BEG[6]
+ Tile_X2Y13_LUT4AB/WW4BEG[7] Tile_X2Y13_LUT4AB/WW4BEG[8] Tile_X2Y13_LUT4AB/WW4BEG[9]
+ Tile_X3Y13_LUT4AB/WW4BEG[0] Tile_X3Y13_LUT4AB/WW4BEG[10] Tile_X3Y13_LUT4AB/WW4BEG[11]
+ Tile_X3Y13_LUT4AB/WW4BEG[12] Tile_X3Y13_LUT4AB/WW4BEG[13] Tile_X3Y13_LUT4AB/WW4BEG[14]
+ Tile_X3Y13_LUT4AB/WW4BEG[15] Tile_X3Y13_LUT4AB/WW4BEG[1] Tile_X3Y13_LUT4AB/WW4BEG[2]
+ Tile_X3Y13_LUT4AB/WW4BEG[3] Tile_X3Y13_LUT4AB/WW4BEG[4] Tile_X3Y13_LUT4AB/WW4BEG[5]
+ Tile_X3Y13_LUT4AB/WW4BEG[6] Tile_X3Y13_LUT4AB/WW4BEG[7] Tile_X3Y13_LUT4AB/WW4BEG[8]
+ Tile_X3Y13_LUT4AB/WW4BEG[9] LUT4AB
XTile_X10Y3_IHP_SRAM Tile_X10Y4_ADDR_SRAM0 Tile_X10Y4_ADDR_SRAM1 Tile_X10Y4_ADDR_SRAM2
+ Tile_X10Y4_ADDR_SRAM3 Tile_X10Y4_ADDR_SRAM4 Tile_X10Y4_ADDR_SRAM5 Tile_X10Y4_ADDR_SRAM6
+ Tile_X10Y4_ADDR_SRAM7 Tile_X10Y4_ADDR_SRAM8 Tile_X10Y4_ADDR_SRAM9 Tile_X10Y4_BM_SRAM0
+ Tile_X10Y4_BM_SRAM1 Tile_X10Y4_BM_SRAM10 Tile_X10Y4_BM_SRAM11 Tile_X10Y4_BM_SRAM12
+ Tile_X10Y4_BM_SRAM13 Tile_X10Y4_BM_SRAM14 Tile_X10Y4_BM_SRAM15 Tile_X10Y4_BM_SRAM16
+ Tile_X10Y4_BM_SRAM17 Tile_X10Y4_BM_SRAM18 Tile_X10Y4_BM_SRAM19 Tile_X10Y4_BM_SRAM2
+ Tile_X10Y4_BM_SRAM20 Tile_X10Y4_BM_SRAM21 Tile_X10Y4_BM_SRAM22 Tile_X10Y4_BM_SRAM23
+ Tile_X10Y4_BM_SRAM24 Tile_X10Y4_BM_SRAM25 Tile_X10Y4_BM_SRAM26 Tile_X10Y4_BM_SRAM27
+ Tile_X10Y4_BM_SRAM28 Tile_X10Y4_BM_SRAM29 Tile_X10Y4_BM_SRAM3 Tile_X10Y4_BM_SRAM30
+ Tile_X10Y4_BM_SRAM31 Tile_X10Y4_BM_SRAM4 Tile_X10Y4_BM_SRAM5 Tile_X10Y4_BM_SRAM6
+ Tile_X10Y4_BM_SRAM7 Tile_X10Y4_BM_SRAM8 Tile_X10Y4_BM_SRAM9 Tile_X10Y4_CLK_SRAM
+ Tile_X10Y4_CONFIGURED_top Tile_X10Y4_DIN_SRAM0 Tile_X10Y4_DIN_SRAM1 Tile_X10Y4_DIN_SRAM10
+ Tile_X10Y4_DIN_SRAM11 Tile_X10Y4_DIN_SRAM12 Tile_X10Y4_DIN_SRAM13 Tile_X10Y4_DIN_SRAM14
+ Tile_X10Y4_DIN_SRAM15 Tile_X10Y4_DIN_SRAM16 Tile_X10Y4_DIN_SRAM17 Tile_X10Y4_DIN_SRAM18
+ Tile_X10Y4_DIN_SRAM19 Tile_X10Y4_DIN_SRAM2 Tile_X10Y4_DIN_SRAM20 Tile_X10Y4_DIN_SRAM21
+ Tile_X10Y4_DIN_SRAM22 Tile_X10Y4_DIN_SRAM23 Tile_X10Y4_DIN_SRAM24 Tile_X10Y4_DIN_SRAM25
+ Tile_X10Y4_DIN_SRAM26 Tile_X10Y4_DIN_SRAM27 Tile_X10Y4_DIN_SRAM28 Tile_X10Y4_DIN_SRAM29
+ Tile_X10Y4_DIN_SRAM3 Tile_X10Y4_DIN_SRAM30 Tile_X10Y4_DIN_SRAM31 Tile_X10Y4_DIN_SRAM4
+ Tile_X10Y4_DIN_SRAM5 Tile_X10Y4_DIN_SRAM6 Tile_X10Y4_DIN_SRAM7 Tile_X10Y4_DIN_SRAM8
+ Tile_X10Y4_DIN_SRAM9 Tile_X10Y4_DOUT_SRAM0 Tile_X10Y4_DOUT_SRAM1 Tile_X10Y4_DOUT_SRAM10
+ Tile_X10Y4_DOUT_SRAM11 Tile_X10Y4_DOUT_SRAM12 Tile_X10Y4_DOUT_SRAM13 Tile_X10Y4_DOUT_SRAM14
+ Tile_X10Y4_DOUT_SRAM15 Tile_X10Y4_DOUT_SRAM16 Tile_X10Y4_DOUT_SRAM17 Tile_X10Y4_DOUT_SRAM18
+ Tile_X10Y4_DOUT_SRAM19 Tile_X10Y4_DOUT_SRAM2 Tile_X10Y4_DOUT_SRAM20 Tile_X10Y4_DOUT_SRAM21
+ Tile_X10Y4_DOUT_SRAM22 Tile_X10Y4_DOUT_SRAM23 Tile_X10Y4_DOUT_SRAM24 Tile_X10Y4_DOUT_SRAM25
+ Tile_X10Y4_DOUT_SRAM26 Tile_X10Y4_DOUT_SRAM27 Tile_X10Y4_DOUT_SRAM28 Tile_X10Y4_DOUT_SRAM29
+ Tile_X10Y4_DOUT_SRAM3 Tile_X10Y4_DOUT_SRAM30 Tile_X10Y4_DOUT_SRAM31 Tile_X10Y4_DOUT_SRAM4
+ Tile_X10Y4_DOUT_SRAM5 Tile_X10Y4_DOUT_SRAM6 Tile_X10Y4_DOUT_SRAM7 Tile_X10Y4_DOUT_SRAM8
+ Tile_X10Y4_DOUT_SRAM9 Tile_X10Y4_MEN_SRAM Tile_X10Y4_REN_SRAM Tile_X10Y4_TIE_HIGH_SRAM
+ Tile_X10Y4_TIE_LOW_SRAM Tile_X9Y3_LUT4AB/E1BEG[0] Tile_X9Y3_LUT4AB/E1BEG[1] Tile_X9Y3_LUT4AB/E1BEG[2]
+ Tile_X9Y3_LUT4AB/E1BEG[3] Tile_X9Y3_LUT4AB/E2BEGb[0] Tile_X9Y3_LUT4AB/E2BEGb[1]
+ Tile_X9Y3_LUT4AB/E2BEGb[2] Tile_X9Y3_LUT4AB/E2BEGb[3] Tile_X9Y3_LUT4AB/E2BEGb[4]
+ Tile_X9Y3_LUT4AB/E2BEGb[5] Tile_X9Y3_LUT4AB/E2BEGb[6] Tile_X9Y3_LUT4AB/E2BEGb[7]
+ Tile_X9Y3_LUT4AB/E2BEG[0] Tile_X9Y3_LUT4AB/E2BEG[1] Tile_X9Y3_LUT4AB/E2BEG[2] Tile_X9Y3_LUT4AB/E2BEG[3]
+ Tile_X9Y3_LUT4AB/E2BEG[4] Tile_X9Y3_LUT4AB/E2BEG[5] Tile_X9Y3_LUT4AB/E2BEG[6] Tile_X9Y3_LUT4AB/E2BEG[7]
+ Tile_X9Y3_LUT4AB/E6BEG[0] Tile_X9Y3_LUT4AB/E6BEG[10] Tile_X9Y3_LUT4AB/E6BEG[11]
+ Tile_X9Y3_LUT4AB/E6BEG[1] Tile_X9Y3_LUT4AB/E6BEG[2] Tile_X9Y3_LUT4AB/E6BEG[3] Tile_X9Y3_LUT4AB/E6BEG[4]
+ Tile_X9Y3_LUT4AB/E6BEG[5] Tile_X9Y3_LUT4AB/E6BEG[6] Tile_X9Y3_LUT4AB/E6BEG[7] Tile_X9Y3_LUT4AB/E6BEG[8]
+ Tile_X9Y3_LUT4AB/E6BEG[9] Tile_X9Y3_LUT4AB/EE4BEG[0] Tile_X9Y3_LUT4AB/EE4BEG[10]
+ Tile_X9Y3_LUT4AB/EE4BEG[11] Tile_X9Y3_LUT4AB/EE4BEG[12] Tile_X9Y3_LUT4AB/EE4BEG[13]
+ Tile_X9Y3_LUT4AB/EE4BEG[14] Tile_X9Y3_LUT4AB/EE4BEG[15] Tile_X9Y3_LUT4AB/EE4BEG[1]
+ Tile_X9Y3_LUT4AB/EE4BEG[2] Tile_X9Y3_LUT4AB/EE4BEG[3] Tile_X9Y3_LUT4AB/EE4BEG[4]
+ Tile_X9Y3_LUT4AB/EE4BEG[5] Tile_X9Y3_LUT4AB/EE4BEG[6] Tile_X9Y3_LUT4AB/EE4BEG[7]
+ Tile_X9Y3_LUT4AB/EE4BEG[8] Tile_X9Y3_LUT4AB/EE4BEG[9] Tile_X9Y3_LUT4AB/FrameData_O[0]
+ Tile_X9Y3_LUT4AB/FrameData_O[10] Tile_X9Y3_LUT4AB/FrameData_O[11] Tile_X9Y3_LUT4AB/FrameData_O[12]
+ Tile_X9Y3_LUT4AB/FrameData_O[13] Tile_X9Y3_LUT4AB/FrameData_O[14] Tile_X9Y3_LUT4AB/FrameData_O[15]
+ Tile_X9Y3_LUT4AB/FrameData_O[16] Tile_X9Y3_LUT4AB/FrameData_O[17] Tile_X9Y3_LUT4AB/FrameData_O[18]
+ Tile_X9Y3_LUT4AB/FrameData_O[19] Tile_X9Y3_LUT4AB/FrameData_O[1] Tile_X9Y3_LUT4AB/FrameData_O[20]
+ Tile_X9Y3_LUT4AB/FrameData_O[21] Tile_X9Y3_LUT4AB/FrameData_O[22] Tile_X9Y3_LUT4AB/FrameData_O[23]
+ Tile_X9Y3_LUT4AB/FrameData_O[24] Tile_X9Y3_LUT4AB/FrameData_O[25] Tile_X9Y3_LUT4AB/FrameData_O[26]
+ Tile_X9Y3_LUT4AB/FrameData_O[27] Tile_X9Y3_LUT4AB/FrameData_O[28] Tile_X9Y3_LUT4AB/FrameData_O[29]
+ Tile_X9Y3_LUT4AB/FrameData_O[2] Tile_X9Y3_LUT4AB/FrameData_O[30] Tile_X9Y3_LUT4AB/FrameData_O[31]
+ Tile_X9Y3_LUT4AB/FrameData_O[3] Tile_X9Y3_LUT4AB/FrameData_O[4] Tile_X9Y3_LUT4AB/FrameData_O[5]
+ Tile_X9Y3_LUT4AB/FrameData_O[6] Tile_X9Y3_LUT4AB/FrameData_O[7] Tile_X9Y3_LUT4AB/FrameData_O[8]
+ Tile_X9Y3_LUT4AB/FrameData_O[9] Tile_X10Y3_IHP_SRAM/Tile_X0Y0_FrameData_O[0] Tile_X10Y3_IHP_SRAM/Tile_X0Y0_FrameData_O[10]
+ Tile_X10Y3_IHP_SRAM/Tile_X0Y0_FrameData_O[11] Tile_X10Y3_IHP_SRAM/Tile_X0Y0_FrameData_O[12]
+ Tile_X10Y3_IHP_SRAM/Tile_X0Y0_FrameData_O[13] Tile_X10Y3_IHP_SRAM/Tile_X0Y0_FrameData_O[14]
+ Tile_X10Y3_IHP_SRAM/Tile_X0Y0_FrameData_O[15] Tile_X10Y3_IHP_SRAM/Tile_X0Y0_FrameData_O[16]
+ Tile_X10Y3_IHP_SRAM/Tile_X0Y0_FrameData_O[17] Tile_X10Y3_IHP_SRAM/Tile_X0Y0_FrameData_O[18]
+ Tile_X10Y3_IHP_SRAM/Tile_X0Y0_FrameData_O[19] Tile_X10Y3_IHP_SRAM/Tile_X0Y0_FrameData_O[1]
+ Tile_X10Y3_IHP_SRAM/Tile_X0Y0_FrameData_O[20] Tile_X10Y3_IHP_SRAM/Tile_X0Y0_FrameData_O[21]
+ Tile_X10Y3_IHP_SRAM/Tile_X0Y0_FrameData_O[22] Tile_X10Y3_IHP_SRAM/Tile_X0Y0_FrameData_O[23]
+ Tile_X10Y3_IHP_SRAM/Tile_X0Y0_FrameData_O[24] Tile_X10Y3_IHP_SRAM/Tile_X0Y0_FrameData_O[25]
+ Tile_X10Y3_IHP_SRAM/Tile_X0Y0_FrameData_O[26] Tile_X10Y3_IHP_SRAM/Tile_X0Y0_FrameData_O[27]
+ Tile_X10Y3_IHP_SRAM/Tile_X0Y0_FrameData_O[28] Tile_X10Y3_IHP_SRAM/Tile_X0Y0_FrameData_O[29]
+ Tile_X10Y3_IHP_SRAM/Tile_X0Y0_FrameData_O[2] Tile_X10Y3_IHP_SRAM/Tile_X0Y0_FrameData_O[30]
+ Tile_X10Y3_IHP_SRAM/Tile_X0Y0_FrameData_O[31] Tile_X10Y3_IHP_SRAM/Tile_X0Y0_FrameData_O[3]
+ Tile_X10Y3_IHP_SRAM/Tile_X0Y0_FrameData_O[4] Tile_X10Y3_IHP_SRAM/Tile_X0Y0_FrameData_O[5]
+ Tile_X10Y3_IHP_SRAM/Tile_X0Y0_FrameData_O[6] Tile_X10Y3_IHP_SRAM/Tile_X0Y0_FrameData_O[7]
+ Tile_X10Y3_IHP_SRAM/Tile_X0Y0_FrameData_O[8] Tile_X10Y3_IHP_SRAM/Tile_X0Y0_FrameData_O[9]
+ Tile_X10Y1_IHP_SRAM/Tile_X0Y1_FrameStrobe[0] Tile_X10Y1_IHP_SRAM/Tile_X0Y1_FrameStrobe[10]
+ Tile_X10Y1_IHP_SRAM/Tile_X0Y1_FrameStrobe[11] Tile_X10Y1_IHP_SRAM/Tile_X0Y1_FrameStrobe[12]
+ Tile_X10Y1_IHP_SRAM/Tile_X0Y1_FrameStrobe[13] Tile_X10Y1_IHP_SRAM/Tile_X0Y1_FrameStrobe[14]
+ Tile_X10Y1_IHP_SRAM/Tile_X0Y1_FrameStrobe[15] Tile_X10Y1_IHP_SRAM/Tile_X0Y1_FrameStrobe[16]
+ Tile_X10Y1_IHP_SRAM/Tile_X0Y1_FrameStrobe[17] Tile_X10Y1_IHP_SRAM/Tile_X0Y1_FrameStrobe[18]
+ Tile_X10Y1_IHP_SRAM/Tile_X0Y1_FrameStrobe[19] Tile_X10Y1_IHP_SRAM/Tile_X0Y1_FrameStrobe[1]
+ Tile_X10Y1_IHP_SRAM/Tile_X0Y1_FrameStrobe[2] Tile_X10Y1_IHP_SRAM/Tile_X0Y1_FrameStrobe[3]
+ Tile_X10Y1_IHP_SRAM/Tile_X0Y1_FrameStrobe[4] Tile_X10Y1_IHP_SRAM/Tile_X0Y1_FrameStrobe[5]
+ Tile_X10Y1_IHP_SRAM/Tile_X0Y1_FrameStrobe[6] Tile_X10Y1_IHP_SRAM/Tile_X0Y1_FrameStrobe[7]
+ Tile_X10Y1_IHP_SRAM/Tile_X0Y1_FrameStrobe[8] Tile_X10Y1_IHP_SRAM/Tile_X0Y1_FrameStrobe[9]
+ Tile_X10Y3_IHP_SRAM/Tile_X0Y0_N1BEG[0] Tile_X10Y3_IHP_SRAM/Tile_X0Y0_N1BEG[1] Tile_X10Y3_IHP_SRAM/Tile_X0Y0_N1BEG[2]
+ Tile_X10Y3_IHP_SRAM/Tile_X0Y0_N1BEG[3] Tile_X10Y3_IHP_SRAM/Tile_X0Y0_N2BEG[0] Tile_X10Y3_IHP_SRAM/Tile_X0Y0_N2BEG[1]
+ Tile_X10Y3_IHP_SRAM/Tile_X0Y0_N2BEG[2] Tile_X10Y3_IHP_SRAM/Tile_X0Y0_N2BEG[3] Tile_X10Y3_IHP_SRAM/Tile_X0Y0_N2BEG[4]
+ Tile_X10Y3_IHP_SRAM/Tile_X0Y0_N2BEG[5] Tile_X10Y3_IHP_SRAM/Tile_X0Y0_N2BEG[6] Tile_X10Y3_IHP_SRAM/Tile_X0Y0_N2BEG[7]
+ Tile_X10Y1_IHP_SRAM/Tile_X0Y1_N2END[0] Tile_X10Y1_IHP_SRAM/Tile_X0Y1_N2END[1] Tile_X10Y1_IHP_SRAM/Tile_X0Y1_N2END[2]
+ Tile_X10Y1_IHP_SRAM/Tile_X0Y1_N2END[3] Tile_X10Y1_IHP_SRAM/Tile_X0Y1_N2END[4] Tile_X10Y1_IHP_SRAM/Tile_X0Y1_N2END[5]
+ Tile_X10Y1_IHP_SRAM/Tile_X0Y1_N2END[6] Tile_X10Y1_IHP_SRAM/Tile_X0Y1_N2END[7] Tile_X10Y3_IHP_SRAM/Tile_X0Y0_N4BEG[0]
+ Tile_X10Y3_IHP_SRAM/Tile_X0Y0_N4BEG[10] Tile_X10Y3_IHP_SRAM/Tile_X0Y0_N4BEG[11]
+ Tile_X10Y3_IHP_SRAM/Tile_X0Y0_N4BEG[12] Tile_X10Y3_IHP_SRAM/Tile_X0Y0_N4BEG[13]
+ Tile_X10Y3_IHP_SRAM/Tile_X0Y0_N4BEG[14] Tile_X10Y3_IHP_SRAM/Tile_X0Y0_N4BEG[15]
+ Tile_X10Y3_IHP_SRAM/Tile_X0Y0_N4BEG[1] Tile_X10Y3_IHP_SRAM/Tile_X0Y0_N4BEG[2] Tile_X10Y3_IHP_SRAM/Tile_X0Y0_N4BEG[3]
+ Tile_X10Y3_IHP_SRAM/Tile_X0Y0_N4BEG[4] Tile_X10Y3_IHP_SRAM/Tile_X0Y0_N4BEG[5] Tile_X10Y3_IHP_SRAM/Tile_X0Y0_N4BEG[6]
+ Tile_X10Y3_IHP_SRAM/Tile_X0Y0_N4BEG[7] Tile_X10Y3_IHP_SRAM/Tile_X0Y0_N4BEG[8] Tile_X10Y3_IHP_SRAM/Tile_X0Y0_N4BEG[9]
+ Tile_X10Y3_IHP_SRAM/Tile_X0Y0_S1END[0] Tile_X10Y3_IHP_SRAM/Tile_X0Y0_S1END[1] Tile_X10Y3_IHP_SRAM/Tile_X0Y0_S1END[2]
+ Tile_X10Y3_IHP_SRAM/Tile_X0Y0_S1END[3] Tile_X10Y3_IHP_SRAM/Tile_X0Y0_S2END[0] Tile_X10Y3_IHP_SRAM/Tile_X0Y0_S2END[1]
+ Tile_X10Y3_IHP_SRAM/Tile_X0Y0_S2END[2] Tile_X10Y3_IHP_SRAM/Tile_X0Y0_S2END[3] Tile_X10Y3_IHP_SRAM/Tile_X0Y0_S2END[4]
+ Tile_X10Y3_IHP_SRAM/Tile_X0Y0_S2END[5] Tile_X10Y3_IHP_SRAM/Tile_X0Y0_S2END[6] Tile_X10Y3_IHP_SRAM/Tile_X0Y0_S2END[7]
+ Tile_X10Y3_IHP_SRAM/Tile_X0Y0_S2MID[0] Tile_X10Y3_IHP_SRAM/Tile_X0Y0_S2MID[1] Tile_X10Y3_IHP_SRAM/Tile_X0Y0_S2MID[2]
+ Tile_X10Y3_IHP_SRAM/Tile_X0Y0_S2MID[3] Tile_X10Y3_IHP_SRAM/Tile_X0Y0_S2MID[4] Tile_X10Y3_IHP_SRAM/Tile_X0Y0_S2MID[5]
+ Tile_X10Y3_IHP_SRAM/Tile_X0Y0_S2MID[6] Tile_X10Y3_IHP_SRAM/Tile_X0Y0_S2MID[7] Tile_X10Y3_IHP_SRAM/Tile_X0Y0_S4END[0]
+ Tile_X10Y3_IHP_SRAM/Tile_X0Y0_S4END[10] Tile_X10Y3_IHP_SRAM/Tile_X0Y0_S4END[11]
+ Tile_X10Y3_IHP_SRAM/Tile_X0Y0_S4END[12] Tile_X10Y3_IHP_SRAM/Tile_X0Y0_S4END[13]
+ Tile_X10Y3_IHP_SRAM/Tile_X0Y0_S4END[14] Tile_X10Y3_IHP_SRAM/Tile_X0Y0_S4END[15]
+ Tile_X10Y3_IHP_SRAM/Tile_X0Y0_S4END[1] Tile_X10Y3_IHP_SRAM/Tile_X0Y0_S4END[2] Tile_X10Y3_IHP_SRAM/Tile_X0Y0_S4END[3]
+ Tile_X10Y3_IHP_SRAM/Tile_X0Y0_S4END[4] Tile_X10Y3_IHP_SRAM/Tile_X0Y0_S4END[5] Tile_X10Y3_IHP_SRAM/Tile_X0Y0_S4END[6]
+ Tile_X10Y3_IHP_SRAM/Tile_X0Y0_S4END[7] Tile_X10Y3_IHP_SRAM/Tile_X0Y0_S4END[8] Tile_X10Y3_IHP_SRAM/Tile_X0Y0_S4END[9]
+ Tile_X10Y1_IHP_SRAM/Tile_X0Y1_UserCLK Tile_X9Y3_LUT4AB/W1END[0] Tile_X9Y3_LUT4AB/W1END[1]
+ Tile_X9Y3_LUT4AB/W1END[2] Tile_X9Y3_LUT4AB/W1END[3] Tile_X9Y3_LUT4AB/W2MID[0] Tile_X9Y3_LUT4AB/W2MID[1]
+ Tile_X9Y3_LUT4AB/W2MID[2] Tile_X9Y3_LUT4AB/W2MID[3] Tile_X9Y3_LUT4AB/W2MID[4] Tile_X9Y3_LUT4AB/W2MID[5]
+ Tile_X9Y3_LUT4AB/W2MID[6] Tile_X9Y3_LUT4AB/W2MID[7] Tile_X9Y3_LUT4AB/W2END[0] Tile_X9Y3_LUT4AB/W2END[1]
+ Tile_X9Y3_LUT4AB/W2END[2] Tile_X9Y3_LUT4AB/W2END[3] Tile_X9Y3_LUT4AB/W2END[4] Tile_X9Y3_LUT4AB/W2END[5]
+ Tile_X9Y3_LUT4AB/W2END[6] Tile_X9Y3_LUT4AB/W2END[7] Tile_X9Y3_LUT4AB/W6END[0] Tile_X9Y3_LUT4AB/W6END[10]
+ Tile_X9Y3_LUT4AB/W6END[11] Tile_X9Y3_LUT4AB/W6END[1] Tile_X9Y3_LUT4AB/W6END[2] Tile_X9Y3_LUT4AB/W6END[3]
+ Tile_X9Y3_LUT4AB/W6END[4] Tile_X9Y3_LUT4AB/W6END[5] Tile_X9Y3_LUT4AB/W6END[6] Tile_X9Y3_LUT4AB/W6END[7]
+ Tile_X9Y3_LUT4AB/W6END[8] Tile_X9Y3_LUT4AB/W6END[9] Tile_X9Y3_LUT4AB/WW4END[0] Tile_X9Y3_LUT4AB/WW4END[10]
+ Tile_X9Y3_LUT4AB/WW4END[11] Tile_X9Y3_LUT4AB/WW4END[12] Tile_X9Y3_LUT4AB/WW4END[13]
+ Tile_X9Y3_LUT4AB/WW4END[14] Tile_X9Y3_LUT4AB/WW4END[15] Tile_X9Y3_LUT4AB/WW4END[1]
+ Tile_X9Y3_LUT4AB/WW4END[2] Tile_X9Y3_LUT4AB/WW4END[3] Tile_X9Y3_LUT4AB/WW4END[4]
+ Tile_X9Y3_LUT4AB/WW4END[5] Tile_X9Y3_LUT4AB/WW4END[6] Tile_X9Y3_LUT4AB/WW4END[7]
+ Tile_X9Y3_LUT4AB/WW4END[8] Tile_X9Y3_LUT4AB/WW4END[9] Tile_X9Y4_LUT4AB/E1BEG[0]
+ Tile_X9Y4_LUT4AB/E1BEG[1] Tile_X9Y4_LUT4AB/E1BEG[2] Tile_X9Y4_LUT4AB/E1BEG[3] Tile_X9Y4_LUT4AB/E2BEGb[0]
+ Tile_X9Y4_LUT4AB/E2BEGb[1] Tile_X9Y4_LUT4AB/E2BEGb[2] Tile_X9Y4_LUT4AB/E2BEGb[3]
+ Tile_X9Y4_LUT4AB/E2BEGb[4] Tile_X9Y4_LUT4AB/E2BEGb[5] Tile_X9Y4_LUT4AB/E2BEGb[6]
+ Tile_X9Y4_LUT4AB/E2BEGb[7] Tile_X9Y4_LUT4AB/E2BEG[0] Tile_X9Y4_LUT4AB/E2BEG[1] Tile_X9Y4_LUT4AB/E2BEG[2]
+ Tile_X9Y4_LUT4AB/E2BEG[3] Tile_X9Y4_LUT4AB/E2BEG[4] Tile_X9Y4_LUT4AB/E2BEG[5] Tile_X9Y4_LUT4AB/E2BEG[6]
+ Tile_X9Y4_LUT4AB/E2BEG[7] Tile_X9Y4_LUT4AB/E6BEG[0] Tile_X9Y4_LUT4AB/E6BEG[10] Tile_X9Y4_LUT4AB/E6BEG[11]
+ Tile_X9Y4_LUT4AB/E6BEG[1] Tile_X9Y4_LUT4AB/E6BEG[2] Tile_X9Y4_LUT4AB/E6BEG[3] Tile_X9Y4_LUT4AB/E6BEG[4]
+ Tile_X9Y4_LUT4AB/E6BEG[5] Tile_X9Y4_LUT4AB/E6BEG[6] Tile_X9Y4_LUT4AB/E6BEG[7] Tile_X9Y4_LUT4AB/E6BEG[8]
+ Tile_X9Y4_LUT4AB/E6BEG[9] Tile_X9Y4_LUT4AB/EE4BEG[0] Tile_X9Y4_LUT4AB/EE4BEG[10]
+ Tile_X9Y4_LUT4AB/EE4BEG[11] Tile_X9Y4_LUT4AB/EE4BEG[12] Tile_X9Y4_LUT4AB/EE4BEG[13]
+ Tile_X9Y4_LUT4AB/EE4BEG[14] Tile_X9Y4_LUT4AB/EE4BEG[15] Tile_X9Y4_LUT4AB/EE4BEG[1]
+ Tile_X9Y4_LUT4AB/EE4BEG[2] Tile_X9Y4_LUT4AB/EE4BEG[3] Tile_X9Y4_LUT4AB/EE4BEG[4]
+ Tile_X9Y4_LUT4AB/EE4BEG[5] Tile_X9Y4_LUT4AB/EE4BEG[6] Tile_X9Y4_LUT4AB/EE4BEG[7]
+ Tile_X9Y4_LUT4AB/EE4BEG[8] Tile_X9Y4_LUT4AB/EE4BEG[9] Tile_X9Y4_LUT4AB/FrameData_O[0]
+ Tile_X9Y4_LUT4AB/FrameData_O[10] Tile_X9Y4_LUT4AB/FrameData_O[11] Tile_X9Y4_LUT4AB/FrameData_O[12]
+ Tile_X9Y4_LUT4AB/FrameData_O[13] Tile_X9Y4_LUT4AB/FrameData_O[14] Tile_X9Y4_LUT4AB/FrameData_O[15]
+ Tile_X9Y4_LUT4AB/FrameData_O[16] Tile_X9Y4_LUT4AB/FrameData_O[17] Tile_X9Y4_LUT4AB/FrameData_O[18]
+ Tile_X9Y4_LUT4AB/FrameData_O[19] Tile_X9Y4_LUT4AB/FrameData_O[1] Tile_X9Y4_LUT4AB/FrameData_O[20]
+ Tile_X9Y4_LUT4AB/FrameData_O[21] Tile_X9Y4_LUT4AB/FrameData_O[22] Tile_X9Y4_LUT4AB/FrameData_O[23]
+ Tile_X9Y4_LUT4AB/FrameData_O[24] Tile_X9Y4_LUT4AB/FrameData_O[25] Tile_X9Y4_LUT4AB/FrameData_O[26]
+ Tile_X9Y4_LUT4AB/FrameData_O[27] Tile_X9Y4_LUT4AB/FrameData_O[28] Tile_X9Y4_LUT4AB/FrameData_O[29]
+ Tile_X9Y4_LUT4AB/FrameData_O[2] Tile_X9Y4_LUT4AB/FrameData_O[30] Tile_X9Y4_LUT4AB/FrameData_O[31]
+ Tile_X9Y4_LUT4AB/FrameData_O[3] Tile_X9Y4_LUT4AB/FrameData_O[4] Tile_X9Y4_LUT4AB/FrameData_O[5]
+ Tile_X9Y4_LUT4AB/FrameData_O[6] Tile_X9Y4_LUT4AB/FrameData_O[7] Tile_X9Y4_LUT4AB/FrameData_O[8]
+ Tile_X9Y4_LUT4AB/FrameData_O[9] Tile_X10Y3_IHP_SRAM/Tile_X0Y1_FrameData_O[0] Tile_X10Y3_IHP_SRAM/Tile_X0Y1_FrameData_O[10]
+ Tile_X10Y3_IHP_SRAM/Tile_X0Y1_FrameData_O[11] Tile_X10Y3_IHP_SRAM/Tile_X0Y1_FrameData_O[12]
+ Tile_X10Y3_IHP_SRAM/Tile_X0Y1_FrameData_O[13] Tile_X10Y3_IHP_SRAM/Tile_X0Y1_FrameData_O[14]
+ Tile_X10Y3_IHP_SRAM/Tile_X0Y1_FrameData_O[15] Tile_X10Y3_IHP_SRAM/Tile_X0Y1_FrameData_O[16]
+ Tile_X10Y3_IHP_SRAM/Tile_X0Y1_FrameData_O[17] Tile_X10Y3_IHP_SRAM/Tile_X0Y1_FrameData_O[18]
+ Tile_X10Y3_IHP_SRAM/Tile_X0Y1_FrameData_O[19] Tile_X10Y3_IHP_SRAM/Tile_X0Y1_FrameData_O[1]
+ Tile_X10Y3_IHP_SRAM/Tile_X0Y1_FrameData_O[20] Tile_X10Y3_IHP_SRAM/Tile_X0Y1_FrameData_O[21]
+ Tile_X10Y3_IHP_SRAM/Tile_X0Y1_FrameData_O[22] Tile_X10Y3_IHP_SRAM/Tile_X0Y1_FrameData_O[23]
+ Tile_X10Y3_IHP_SRAM/Tile_X0Y1_FrameData_O[24] Tile_X10Y3_IHP_SRAM/Tile_X0Y1_FrameData_O[25]
+ Tile_X10Y3_IHP_SRAM/Tile_X0Y1_FrameData_O[26] Tile_X10Y3_IHP_SRAM/Tile_X0Y1_FrameData_O[27]
+ Tile_X10Y3_IHP_SRAM/Tile_X0Y1_FrameData_O[28] Tile_X10Y3_IHP_SRAM/Tile_X0Y1_FrameData_O[29]
+ Tile_X10Y3_IHP_SRAM/Tile_X0Y1_FrameData_O[2] Tile_X10Y3_IHP_SRAM/Tile_X0Y1_FrameData_O[30]
+ Tile_X10Y3_IHP_SRAM/Tile_X0Y1_FrameData_O[31] Tile_X10Y3_IHP_SRAM/Tile_X0Y1_FrameData_O[3]
+ Tile_X10Y3_IHP_SRAM/Tile_X0Y1_FrameData_O[4] Tile_X10Y3_IHP_SRAM/Tile_X0Y1_FrameData_O[5]
+ Tile_X10Y3_IHP_SRAM/Tile_X0Y1_FrameData_O[6] Tile_X10Y3_IHP_SRAM/Tile_X0Y1_FrameData_O[7]
+ Tile_X10Y3_IHP_SRAM/Tile_X0Y1_FrameData_O[8] Tile_X10Y3_IHP_SRAM/Tile_X0Y1_FrameData_O[9]
+ Tile_X10Y3_IHP_SRAM/Tile_X0Y1_FrameStrobe[0] Tile_X10Y3_IHP_SRAM/Tile_X0Y1_FrameStrobe[10]
+ Tile_X10Y3_IHP_SRAM/Tile_X0Y1_FrameStrobe[11] Tile_X10Y3_IHP_SRAM/Tile_X0Y1_FrameStrobe[12]
+ Tile_X10Y3_IHP_SRAM/Tile_X0Y1_FrameStrobe[13] Tile_X10Y3_IHP_SRAM/Tile_X0Y1_FrameStrobe[14]
+ Tile_X10Y3_IHP_SRAM/Tile_X0Y1_FrameStrobe[15] Tile_X10Y3_IHP_SRAM/Tile_X0Y1_FrameStrobe[16]
+ Tile_X10Y3_IHP_SRAM/Tile_X0Y1_FrameStrobe[17] Tile_X10Y3_IHP_SRAM/Tile_X0Y1_FrameStrobe[18]
+ Tile_X10Y3_IHP_SRAM/Tile_X0Y1_FrameStrobe[19] Tile_X10Y3_IHP_SRAM/Tile_X0Y1_FrameStrobe[1]
+ Tile_X10Y3_IHP_SRAM/Tile_X0Y1_FrameStrobe[2] Tile_X10Y3_IHP_SRAM/Tile_X0Y1_FrameStrobe[3]
+ Tile_X10Y3_IHP_SRAM/Tile_X0Y1_FrameStrobe[4] Tile_X10Y3_IHP_SRAM/Tile_X0Y1_FrameStrobe[5]
+ Tile_X10Y3_IHP_SRAM/Tile_X0Y1_FrameStrobe[6] Tile_X10Y3_IHP_SRAM/Tile_X0Y1_FrameStrobe[7]
+ Tile_X10Y3_IHP_SRAM/Tile_X0Y1_FrameStrobe[8] Tile_X10Y3_IHP_SRAM/Tile_X0Y1_FrameStrobe[9]
+ Tile_X10Y5_IHP_SRAM/Tile_X0Y0_N1BEG[0] Tile_X10Y5_IHP_SRAM/Tile_X0Y0_N1BEG[1] Tile_X10Y5_IHP_SRAM/Tile_X0Y0_N1BEG[2]
+ Tile_X10Y5_IHP_SRAM/Tile_X0Y0_N1BEG[3] Tile_X10Y3_IHP_SRAM/Tile_X0Y1_N2END[0] Tile_X10Y3_IHP_SRAM/Tile_X0Y1_N2END[1]
+ Tile_X10Y3_IHP_SRAM/Tile_X0Y1_N2END[2] Tile_X10Y3_IHP_SRAM/Tile_X0Y1_N2END[3] Tile_X10Y3_IHP_SRAM/Tile_X0Y1_N2END[4]
+ Tile_X10Y3_IHP_SRAM/Tile_X0Y1_N2END[5] Tile_X10Y3_IHP_SRAM/Tile_X0Y1_N2END[6] Tile_X10Y3_IHP_SRAM/Tile_X0Y1_N2END[7]
+ Tile_X10Y5_IHP_SRAM/Tile_X0Y0_N2BEG[0] Tile_X10Y5_IHP_SRAM/Tile_X0Y0_N2BEG[1] Tile_X10Y5_IHP_SRAM/Tile_X0Y0_N2BEG[2]
+ Tile_X10Y5_IHP_SRAM/Tile_X0Y0_N2BEG[3] Tile_X10Y5_IHP_SRAM/Tile_X0Y0_N2BEG[4] Tile_X10Y5_IHP_SRAM/Tile_X0Y0_N2BEG[5]
+ Tile_X10Y5_IHP_SRAM/Tile_X0Y0_N2BEG[6] Tile_X10Y5_IHP_SRAM/Tile_X0Y0_N2BEG[7] Tile_X10Y5_IHP_SRAM/Tile_X0Y0_N4BEG[0]
+ Tile_X10Y5_IHP_SRAM/Tile_X0Y0_N4BEG[10] Tile_X10Y5_IHP_SRAM/Tile_X0Y0_N4BEG[11]
+ Tile_X10Y5_IHP_SRAM/Tile_X0Y0_N4BEG[12] Tile_X10Y5_IHP_SRAM/Tile_X0Y0_N4BEG[13]
+ Tile_X10Y5_IHP_SRAM/Tile_X0Y0_N4BEG[14] Tile_X10Y5_IHP_SRAM/Tile_X0Y0_N4BEG[15]
+ Tile_X10Y5_IHP_SRAM/Tile_X0Y0_N4BEG[1] Tile_X10Y5_IHP_SRAM/Tile_X0Y0_N4BEG[2] Tile_X10Y5_IHP_SRAM/Tile_X0Y0_N4BEG[3]
+ Tile_X10Y5_IHP_SRAM/Tile_X0Y0_N4BEG[4] Tile_X10Y5_IHP_SRAM/Tile_X0Y0_N4BEG[5] Tile_X10Y5_IHP_SRAM/Tile_X0Y0_N4BEG[6]
+ Tile_X10Y5_IHP_SRAM/Tile_X0Y0_N4BEG[7] Tile_X10Y5_IHP_SRAM/Tile_X0Y0_N4BEG[8] Tile_X10Y5_IHP_SRAM/Tile_X0Y0_N4BEG[9]
+ Tile_X10Y5_IHP_SRAM/Tile_X0Y0_S1END[0] Tile_X10Y5_IHP_SRAM/Tile_X0Y0_S1END[1] Tile_X10Y5_IHP_SRAM/Tile_X0Y0_S1END[2]
+ Tile_X10Y5_IHP_SRAM/Tile_X0Y0_S1END[3] Tile_X10Y5_IHP_SRAM/Tile_X0Y0_S2MID[0] Tile_X10Y5_IHP_SRAM/Tile_X0Y0_S2MID[1]
+ Tile_X10Y5_IHP_SRAM/Tile_X0Y0_S2MID[2] Tile_X10Y5_IHP_SRAM/Tile_X0Y0_S2MID[3] Tile_X10Y5_IHP_SRAM/Tile_X0Y0_S2MID[4]
+ Tile_X10Y5_IHP_SRAM/Tile_X0Y0_S2MID[5] Tile_X10Y5_IHP_SRAM/Tile_X0Y0_S2MID[6] Tile_X10Y5_IHP_SRAM/Tile_X0Y0_S2MID[7]
+ Tile_X10Y5_IHP_SRAM/Tile_X0Y0_S2END[0] Tile_X10Y5_IHP_SRAM/Tile_X0Y0_S2END[1] Tile_X10Y5_IHP_SRAM/Tile_X0Y0_S2END[2]
+ Tile_X10Y5_IHP_SRAM/Tile_X0Y0_S2END[3] Tile_X10Y5_IHP_SRAM/Tile_X0Y0_S2END[4] Tile_X10Y5_IHP_SRAM/Tile_X0Y0_S2END[5]
+ Tile_X10Y5_IHP_SRAM/Tile_X0Y0_S2END[6] Tile_X10Y5_IHP_SRAM/Tile_X0Y0_S2END[7] Tile_X10Y5_IHP_SRAM/Tile_X0Y0_S4END[0]
+ Tile_X10Y5_IHP_SRAM/Tile_X0Y0_S4END[10] Tile_X10Y5_IHP_SRAM/Tile_X0Y0_S4END[11]
+ Tile_X10Y5_IHP_SRAM/Tile_X0Y0_S4END[12] Tile_X10Y5_IHP_SRAM/Tile_X0Y0_S4END[13]
+ Tile_X10Y5_IHP_SRAM/Tile_X0Y0_S4END[14] Tile_X10Y5_IHP_SRAM/Tile_X0Y0_S4END[15]
+ Tile_X10Y5_IHP_SRAM/Tile_X0Y0_S4END[1] Tile_X10Y5_IHP_SRAM/Tile_X0Y0_S4END[2] Tile_X10Y5_IHP_SRAM/Tile_X0Y0_S4END[3]
+ Tile_X10Y5_IHP_SRAM/Tile_X0Y0_S4END[4] Tile_X10Y5_IHP_SRAM/Tile_X0Y0_S4END[5] Tile_X10Y5_IHP_SRAM/Tile_X0Y0_S4END[6]
+ Tile_X10Y5_IHP_SRAM/Tile_X0Y0_S4END[7] Tile_X10Y5_IHP_SRAM/Tile_X0Y0_S4END[8] Tile_X10Y5_IHP_SRAM/Tile_X0Y0_S4END[9]
+ Tile_X10Y3_IHP_SRAM/Tile_X0Y1_UserCLK Tile_X9Y4_LUT4AB/W1END[0] Tile_X9Y4_LUT4AB/W1END[1]
+ Tile_X9Y4_LUT4AB/W1END[2] Tile_X9Y4_LUT4AB/W1END[3] Tile_X9Y4_LUT4AB/W2MID[0] Tile_X9Y4_LUT4AB/W2MID[1]
+ Tile_X9Y4_LUT4AB/W2MID[2] Tile_X9Y4_LUT4AB/W2MID[3] Tile_X9Y4_LUT4AB/W2MID[4] Tile_X9Y4_LUT4AB/W2MID[5]
+ Tile_X9Y4_LUT4AB/W2MID[6] Tile_X9Y4_LUT4AB/W2MID[7] Tile_X9Y4_LUT4AB/W2END[0] Tile_X9Y4_LUT4AB/W2END[1]
+ Tile_X9Y4_LUT4AB/W2END[2] Tile_X9Y4_LUT4AB/W2END[3] Tile_X9Y4_LUT4AB/W2END[4] Tile_X9Y4_LUT4AB/W2END[5]
+ Tile_X9Y4_LUT4AB/W2END[6] Tile_X9Y4_LUT4AB/W2END[7] Tile_X9Y4_LUT4AB/W6END[0] Tile_X9Y4_LUT4AB/W6END[10]
+ Tile_X9Y4_LUT4AB/W6END[11] Tile_X9Y4_LUT4AB/W6END[1] Tile_X9Y4_LUT4AB/W6END[2] Tile_X9Y4_LUT4AB/W6END[3]
+ Tile_X9Y4_LUT4AB/W6END[4] Tile_X9Y4_LUT4AB/W6END[5] Tile_X9Y4_LUT4AB/W6END[6] Tile_X9Y4_LUT4AB/W6END[7]
+ Tile_X9Y4_LUT4AB/W6END[8] Tile_X9Y4_LUT4AB/W6END[9] Tile_X9Y4_LUT4AB/WW4END[0] Tile_X9Y4_LUT4AB/WW4END[10]
+ Tile_X9Y4_LUT4AB/WW4END[11] Tile_X9Y4_LUT4AB/WW4END[12] Tile_X9Y4_LUT4AB/WW4END[13]
+ Tile_X9Y4_LUT4AB/WW4END[14] Tile_X9Y4_LUT4AB/WW4END[15] Tile_X9Y4_LUT4AB/WW4END[1]
+ Tile_X9Y4_LUT4AB/WW4END[2] Tile_X9Y4_LUT4AB/WW4END[3] Tile_X9Y4_LUT4AB/WW4END[4]
+ Tile_X9Y4_LUT4AB/WW4END[5] Tile_X9Y4_LUT4AB/WW4END[6] Tile_X9Y4_LUT4AB/WW4END[7]
+ Tile_X9Y4_LUT4AB/WW4END[8] Tile_X9Y4_LUT4AB/WW4END[9] VGND VPWR Tile_X10Y4_WEN_SRAM
+ IHP_SRAM
XTile_X4Y4_RegFile Tile_X5Y4_LUT4AB/E1END[0] Tile_X5Y4_LUT4AB/E1END[1] Tile_X5Y4_LUT4AB/E1END[2]
+ Tile_X5Y4_LUT4AB/E1END[3] Tile_X3Y4_LUT4AB/E1BEG[0] Tile_X3Y4_LUT4AB/E1BEG[1] Tile_X3Y4_LUT4AB/E1BEG[2]
+ Tile_X3Y4_LUT4AB/E1BEG[3] Tile_X5Y4_LUT4AB/E2MID[0] Tile_X5Y4_LUT4AB/E2MID[1] Tile_X5Y4_LUT4AB/E2MID[2]
+ Tile_X5Y4_LUT4AB/E2MID[3] Tile_X5Y4_LUT4AB/E2MID[4] Tile_X5Y4_LUT4AB/E2MID[5] Tile_X5Y4_LUT4AB/E2MID[6]
+ Tile_X5Y4_LUT4AB/E2MID[7] Tile_X5Y4_LUT4AB/E2END[0] Tile_X5Y4_LUT4AB/E2END[1] Tile_X5Y4_LUT4AB/E2END[2]
+ Tile_X5Y4_LUT4AB/E2END[3] Tile_X5Y4_LUT4AB/E2END[4] Tile_X5Y4_LUT4AB/E2END[5] Tile_X5Y4_LUT4AB/E2END[6]
+ Tile_X5Y4_LUT4AB/E2END[7] Tile_X4Y4_RegFile/E2END[0] Tile_X4Y4_RegFile/E2END[1]
+ Tile_X4Y4_RegFile/E2END[2] Tile_X4Y4_RegFile/E2END[3] Tile_X4Y4_RegFile/E2END[4]
+ Tile_X4Y4_RegFile/E2END[5] Tile_X4Y4_RegFile/E2END[6] Tile_X4Y4_RegFile/E2END[7]
+ Tile_X3Y4_LUT4AB/E2BEG[0] Tile_X3Y4_LUT4AB/E2BEG[1] Tile_X3Y4_LUT4AB/E2BEG[2] Tile_X3Y4_LUT4AB/E2BEG[3]
+ Tile_X3Y4_LUT4AB/E2BEG[4] Tile_X3Y4_LUT4AB/E2BEG[5] Tile_X3Y4_LUT4AB/E2BEG[6] Tile_X3Y4_LUT4AB/E2BEG[7]
+ Tile_X5Y4_LUT4AB/E6END[0] Tile_X5Y4_LUT4AB/E6END[10] Tile_X5Y4_LUT4AB/E6END[11]
+ Tile_X5Y4_LUT4AB/E6END[1] Tile_X5Y4_LUT4AB/E6END[2] Tile_X5Y4_LUT4AB/E6END[3] Tile_X5Y4_LUT4AB/E6END[4]
+ Tile_X5Y4_LUT4AB/E6END[5] Tile_X5Y4_LUT4AB/E6END[6] Tile_X5Y4_LUT4AB/E6END[7] Tile_X5Y4_LUT4AB/E6END[8]
+ Tile_X5Y4_LUT4AB/E6END[9] Tile_X3Y4_LUT4AB/E6BEG[0] Tile_X3Y4_LUT4AB/E6BEG[10] Tile_X3Y4_LUT4AB/E6BEG[11]
+ Tile_X3Y4_LUT4AB/E6BEG[1] Tile_X3Y4_LUT4AB/E6BEG[2] Tile_X3Y4_LUT4AB/E6BEG[3] Tile_X3Y4_LUT4AB/E6BEG[4]
+ Tile_X3Y4_LUT4AB/E6BEG[5] Tile_X3Y4_LUT4AB/E6BEG[6] Tile_X3Y4_LUT4AB/E6BEG[7] Tile_X3Y4_LUT4AB/E6BEG[8]
+ Tile_X3Y4_LUT4AB/E6BEG[9] Tile_X5Y4_LUT4AB/EE4END[0] Tile_X5Y4_LUT4AB/EE4END[10]
+ Tile_X5Y4_LUT4AB/EE4END[11] Tile_X5Y4_LUT4AB/EE4END[12] Tile_X5Y4_LUT4AB/EE4END[13]
+ Tile_X5Y4_LUT4AB/EE4END[14] Tile_X5Y4_LUT4AB/EE4END[15] Tile_X5Y4_LUT4AB/EE4END[1]
+ Tile_X5Y4_LUT4AB/EE4END[2] Tile_X5Y4_LUT4AB/EE4END[3] Tile_X5Y4_LUT4AB/EE4END[4]
+ Tile_X5Y4_LUT4AB/EE4END[5] Tile_X5Y4_LUT4AB/EE4END[6] Tile_X5Y4_LUT4AB/EE4END[7]
+ Tile_X5Y4_LUT4AB/EE4END[8] Tile_X5Y4_LUT4AB/EE4END[9] Tile_X3Y4_LUT4AB/EE4BEG[0]
+ Tile_X3Y4_LUT4AB/EE4BEG[10] Tile_X3Y4_LUT4AB/EE4BEG[11] Tile_X3Y4_LUT4AB/EE4BEG[12]
+ Tile_X3Y4_LUT4AB/EE4BEG[13] Tile_X3Y4_LUT4AB/EE4BEG[14] Tile_X3Y4_LUT4AB/EE4BEG[15]
+ Tile_X3Y4_LUT4AB/EE4BEG[1] Tile_X3Y4_LUT4AB/EE4BEG[2] Tile_X3Y4_LUT4AB/EE4BEG[3]
+ Tile_X3Y4_LUT4AB/EE4BEG[4] Tile_X3Y4_LUT4AB/EE4BEG[5] Tile_X3Y4_LUT4AB/EE4BEG[6]
+ Tile_X3Y4_LUT4AB/EE4BEG[7] Tile_X3Y4_LUT4AB/EE4BEG[8] Tile_X3Y4_LUT4AB/EE4BEG[9]
+ Tile_X4Y4_RegFile/FrameData[0] Tile_X4Y4_RegFile/FrameData[10] Tile_X4Y4_RegFile/FrameData[11]
+ Tile_X4Y4_RegFile/FrameData[12] Tile_X4Y4_RegFile/FrameData[13] Tile_X4Y4_RegFile/FrameData[14]
+ Tile_X4Y4_RegFile/FrameData[15] Tile_X4Y4_RegFile/FrameData[16] Tile_X4Y4_RegFile/FrameData[17]
+ Tile_X4Y4_RegFile/FrameData[18] Tile_X4Y4_RegFile/FrameData[19] Tile_X4Y4_RegFile/FrameData[1]
+ Tile_X4Y4_RegFile/FrameData[20] Tile_X4Y4_RegFile/FrameData[21] Tile_X4Y4_RegFile/FrameData[22]
+ Tile_X4Y4_RegFile/FrameData[23] Tile_X4Y4_RegFile/FrameData[24] Tile_X4Y4_RegFile/FrameData[25]
+ Tile_X4Y4_RegFile/FrameData[26] Tile_X4Y4_RegFile/FrameData[27] Tile_X4Y4_RegFile/FrameData[28]
+ Tile_X4Y4_RegFile/FrameData[29] Tile_X4Y4_RegFile/FrameData[2] Tile_X4Y4_RegFile/FrameData[30]
+ Tile_X4Y4_RegFile/FrameData[31] Tile_X4Y4_RegFile/FrameData[3] Tile_X4Y4_RegFile/FrameData[4]
+ Tile_X4Y4_RegFile/FrameData[5] Tile_X4Y4_RegFile/FrameData[6] Tile_X4Y4_RegFile/FrameData[7]
+ Tile_X4Y4_RegFile/FrameData[8] Tile_X4Y4_RegFile/FrameData[9] Tile_X5Y4_LUT4AB/FrameData[0]
+ Tile_X5Y4_LUT4AB/FrameData[10] Tile_X5Y4_LUT4AB/FrameData[11] Tile_X5Y4_LUT4AB/FrameData[12]
+ Tile_X5Y4_LUT4AB/FrameData[13] Tile_X5Y4_LUT4AB/FrameData[14] Tile_X5Y4_LUT4AB/FrameData[15]
+ Tile_X5Y4_LUT4AB/FrameData[16] Tile_X5Y4_LUT4AB/FrameData[17] Tile_X5Y4_LUT4AB/FrameData[18]
+ Tile_X5Y4_LUT4AB/FrameData[19] Tile_X5Y4_LUT4AB/FrameData[1] Tile_X5Y4_LUT4AB/FrameData[20]
+ Tile_X5Y4_LUT4AB/FrameData[21] Tile_X5Y4_LUT4AB/FrameData[22] Tile_X5Y4_LUT4AB/FrameData[23]
+ Tile_X5Y4_LUT4AB/FrameData[24] Tile_X5Y4_LUT4AB/FrameData[25] Tile_X5Y4_LUT4AB/FrameData[26]
+ Tile_X5Y4_LUT4AB/FrameData[27] Tile_X5Y4_LUT4AB/FrameData[28] Tile_X5Y4_LUT4AB/FrameData[29]
+ Tile_X5Y4_LUT4AB/FrameData[2] Tile_X5Y4_LUT4AB/FrameData[30] Tile_X5Y4_LUT4AB/FrameData[31]
+ Tile_X5Y4_LUT4AB/FrameData[3] Tile_X5Y4_LUT4AB/FrameData[4] Tile_X5Y4_LUT4AB/FrameData[5]
+ Tile_X5Y4_LUT4AB/FrameData[6] Tile_X5Y4_LUT4AB/FrameData[7] Tile_X5Y4_LUT4AB/FrameData[8]
+ Tile_X5Y4_LUT4AB/FrameData[9] Tile_X4Y4_RegFile/FrameStrobe[0] Tile_X4Y4_RegFile/FrameStrobe[10]
+ Tile_X4Y4_RegFile/FrameStrobe[11] Tile_X4Y4_RegFile/FrameStrobe[12] Tile_X4Y4_RegFile/FrameStrobe[13]
+ Tile_X4Y4_RegFile/FrameStrobe[14] Tile_X4Y4_RegFile/FrameStrobe[15] Tile_X4Y4_RegFile/FrameStrobe[16]
+ Tile_X4Y4_RegFile/FrameStrobe[17] Tile_X4Y4_RegFile/FrameStrobe[18] Tile_X4Y4_RegFile/FrameStrobe[19]
+ Tile_X4Y4_RegFile/FrameStrobe[1] Tile_X4Y4_RegFile/FrameStrobe[2] Tile_X4Y4_RegFile/FrameStrobe[3]
+ Tile_X4Y4_RegFile/FrameStrobe[4] Tile_X4Y4_RegFile/FrameStrobe[5] Tile_X4Y4_RegFile/FrameStrobe[6]
+ Tile_X4Y4_RegFile/FrameStrobe[7] Tile_X4Y4_RegFile/FrameStrobe[8] Tile_X4Y4_RegFile/FrameStrobe[9]
+ Tile_X4Y3_RegFile/FrameStrobe[0] Tile_X4Y3_RegFile/FrameStrobe[10] Tile_X4Y3_RegFile/FrameStrobe[11]
+ Tile_X4Y3_RegFile/FrameStrobe[12] Tile_X4Y3_RegFile/FrameStrobe[13] Tile_X4Y3_RegFile/FrameStrobe[14]
+ Tile_X4Y3_RegFile/FrameStrobe[15] Tile_X4Y3_RegFile/FrameStrobe[16] Tile_X4Y3_RegFile/FrameStrobe[17]
+ Tile_X4Y3_RegFile/FrameStrobe[18] Tile_X4Y3_RegFile/FrameStrobe[19] Tile_X4Y3_RegFile/FrameStrobe[1]
+ Tile_X4Y3_RegFile/FrameStrobe[2] Tile_X4Y3_RegFile/FrameStrobe[3] Tile_X4Y3_RegFile/FrameStrobe[4]
+ Tile_X4Y3_RegFile/FrameStrobe[5] Tile_X4Y3_RegFile/FrameStrobe[6] Tile_X4Y3_RegFile/FrameStrobe[7]
+ Tile_X4Y3_RegFile/FrameStrobe[8] Tile_X4Y3_RegFile/FrameStrobe[9] Tile_X4Y4_RegFile/N1BEG[0]
+ Tile_X4Y4_RegFile/N1BEG[1] Tile_X4Y4_RegFile/N1BEG[2] Tile_X4Y4_RegFile/N1BEG[3]
+ Tile_X4Y5_RegFile/N1BEG[0] Tile_X4Y5_RegFile/N1BEG[1] Tile_X4Y5_RegFile/N1BEG[2]
+ Tile_X4Y5_RegFile/N1BEG[3] Tile_X4Y4_RegFile/N2BEG[0] Tile_X4Y4_RegFile/N2BEG[1]
+ Tile_X4Y4_RegFile/N2BEG[2] Tile_X4Y4_RegFile/N2BEG[3] Tile_X4Y4_RegFile/N2BEG[4]
+ Tile_X4Y4_RegFile/N2BEG[5] Tile_X4Y4_RegFile/N2BEG[6] Tile_X4Y4_RegFile/N2BEG[7]
+ Tile_X4Y3_RegFile/N2END[0] Tile_X4Y3_RegFile/N2END[1] Tile_X4Y3_RegFile/N2END[2]
+ Tile_X4Y3_RegFile/N2END[3] Tile_X4Y3_RegFile/N2END[4] Tile_X4Y3_RegFile/N2END[5]
+ Tile_X4Y3_RegFile/N2END[6] Tile_X4Y3_RegFile/N2END[7] Tile_X4Y4_RegFile/N2END[0]
+ Tile_X4Y4_RegFile/N2END[1] Tile_X4Y4_RegFile/N2END[2] Tile_X4Y4_RegFile/N2END[3]
+ Tile_X4Y4_RegFile/N2END[4] Tile_X4Y4_RegFile/N2END[5] Tile_X4Y4_RegFile/N2END[6]
+ Tile_X4Y4_RegFile/N2END[7] Tile_X4Y5_RegFile/N2BEG[0] Tile_X4Y5_RegFile/N2BEG[1]
+ Tile_X4Y5_RegFile/N2BEG[2] Tile_X4Y5_RegFile/N2BEG[3] Tile_X4Y5_RegFile/N2BEG[4]
+ Tile_X4Y5_RegFile/N2BEG[5] Tile_X4Y5_RegFile/N2BEG[6] Tile_X4Y5_RegFile/N2BEG[7]
+ Tile_X4Y4_RegFile/N4BEG[0] Tile_X4Y4_RegFile/N4BEG[10] Tile_X4Y4_RegFile/N4BEG[11]
+ Tile_X4Y4_RegFile/N4BEG[12] Tile_X4Y4_RegFile/N4BEG[13] Tile_X4Y4_RegFile/N4BEG[14]
+ Tile_X4Y4_RegFile/N4BEG[15] Tile_X4Y4_RegFile/N4BEG[1] Tile_X4Y4_RegFile/N4BEG[2]
+ Tile_X4Y4_RegFile/N4BEG[3] Tile_X4Y4_RegFile/N4BEG[4] Tile_X4Y4_RegFile/N4BEG[5]
+ Tile_X4Y4_RegFile/N4BEG[6] Tile_X4Y4_RegFile/N4BEG[7] Tile_X4Y4_RegFile/N4BEG[8]
+ Tile_X4Y4_RegFile/N4BEG[9] Tile_X4Y5_RegFile/N4BEG[0] Tile_X4Y5_RegFile/N4BEG[10]
+ Tile_X4Y5_RegFile/N4BEG[11] Tile_X4Y5_RegFile/N4BEG[12] Tile_X4Y5_RegFile/N4BEG[13]
+ Tile_X4Y5_RegFile/N4BEG[14] Tile_X4Y5_RegFile/N4BEG[15] Tile_X4Y5_RegFile/N4BEG[1]
+ Tile_X4Y5_RegFile/N4BEG[2] Tile_X4Y5_RegFile/N4BEG[3] Tile_X4Y5_RegFile/N4BEG[4]
+ Tile_X4Y5_RegFile/N4BEG[5] Tile_X4Y5_RegFile/N4BEG[6] Tile_X4Y5_RegFile/N4BEG[7]
+ Tile_X4Y5_RegFile/N4BEG[8] Tile_X4Y5_RegFile/N4BEG[9] Tile_X4Y4_RegFile/NN4BEG[0]
+ Tile_X4Y4_RegFile/NN4BEG[10] Tile_X4Y4_RegFile/NN4BEG[11] Tile_X4Y4_RegFile/NN4BEG[12]
+ Tile_X4Y4_RegFile/NN4BEG[13] Tile_X4Y4_RegFile/NN4BEG[14] Tile_X4Y4_RegFile/NN4BEG[15]
+ Tile_X4Y4_RegFile/NN4BEG[1] Tile_X4Y4_RegFile/NN4BEG[2] Tile_X4Y4_RegFile/NN4BEG[3]
+ Tile_X4Y4_RegFile/NN4BEG[4] Tile_X4Y4_RegFile/NN4BEG[5] Tile_X4Y4_RegFile/NN4BEG[6]
+ Tile_X4Y4_RegFile/NN4BEG[7] Tile_X4Y4_RegFile/NN4BEG[8] Tile_X4Y4_RegFile/NN4BEG[9]
+ Tile_X4Y5_RegFile/NN4BEG[0] Tile_X4Y5_RegFile/NN4BEG[10] Tile_X4Y5_RegFile/NN4BEG[11]
+ Tile_X4Y5_RegFile/NN4BEG[12] Tile_X4Y5_RegFile/NN4BEG[13] Tile_X4Y5_RegFile/NN4BEG[14]
+ Tile_X4Y5_RegFile/NN4BEG[15] Tile_X4Y5_RegFile/NN4BEG[1] Tile_X4Y5_RegFile/NN4BEG[2]
+ Tile_X4Y5_RegFile/NN4BEG[3] Tile_X4Y5_RegFile/NN4BEG[4] Tile_X4Y5_RegFile/NN4BEG[5]
+ Tile_X4Y5_RegFile/NN4BEG[6] Tile_X4Y5_RegFile/NN4BEG[7] Tile_X4Y5_RegFile/NN4BEG[8]
+ Tile_X4Y5_RegFile/NN4BEG[9] Tile_X4Y5_RegFile/S1END[0] Tile_X4Y5_RegFile/S1END[1]
+ Tile_X4Y5_RegFile/S1END[2] Tile_X4Y5_RegFile/S1END[3] Tile_X4Y4_RegFile/S1END[0]
+ Tile_X4Y4_RegFile/S1END[1] Tile_X4Y4_RegFile/S1END[2] Tile_X4Y4_RegFile/S1END[3]
+ Tile_X4Y5_RegFile/S2MID[0] Tile_X4Y5_RegFile/S2MID[1] Tile_X4Y5_RegFile/S2MID[2]
+ Tile_X4Y5_RegFile/S2MID[3] Tile_X4Y5_RegFile/S2MID[4] Tile_X4Y5_RegFile/S2MID[5]
+ Tile_X4Y5_RegFile/S2MID[6] Tile_X4Y5_RegFile/S2MID[7] Tile_X4Y5_RegFile/S2END[0]
+ Tile_X4Y5_RegFile/S2END[1] Tile_X4Y5_RegFile/S2END[2] Tile_X4Y5_RegFile/S2END[3]
+ Tile_X4Y5_RegFile/S2END[4] Tile_X4Y5_RegFile/S2END[5] Tile_X4Y5_RegFile/S2END[6]
+ Tile_X4Y5_RegFile/S2END[7] Tile_X4Y4_RegFile/S2END[0] Tile_X4Y4_RegFile/S2END[1]
+ Tile_X4Y4_RegFile/S2END[2] Tile_X4Y4_RegFile/S2END[3] Tile_X4Y4_RegFile/S2END[4]
+ Tile_X4Y4_RegFile/S2END[5] Tile_X4Y4_RegFile/S2END[6] Tile_X4Y4_RegFile/S2END[7]
+ Tile_X4Y4_RegFile/S2MID[0] Tile_X4Y4_RegFile/S2MID[1] Tile_X4Y4_RegFile/S2MID[2]
+ Tile_X4Y4_RegFile/S2MID[3] Tile_X4Y4_RegFile/S2MID[4] Tile_X4Y4_RegFile/S2MID[5]
+ Tile_X4Y4_RegFile/S2MID[6] Tile_X4Y4_RegFile/S2MID[7] Tile_X4Y5_RegFile/S4END[0]
+ Tile_X4Y5_RegFile/S4END[10] Tile_X4Y5_RegFile/S4END[11] Tile_X4Y5_RegFile/S4END[12]
+ Tile_X4Y5_RegFile/S4END[13] Tile_X4Y5_RegFile/S4END[14] Tile_X4Y5_RegFile/S4END[15]
+ Tile_X4Y5_RegFile/S4END[1] Tile_X4Y5_RegFile/S4END[2] Tile_X4Y5_RegFile/S4END[3]
+ Tile_X4Y5_RegFile/S4END[4] Tile_X4Y5_RegFile/S4END[5] Tile_X4Y5_RegFile/S4END[6]
+ Tile_X4Y5_RegFile/S4END[7] Tile_X4Y5_RegFile/S4END[8] Tile_X4Y5_RegFile/S4END[9]
+ Tile_X4Y4_RegFile/S4END[0] Tile_X4Y4_RegFile/S4END[10] Tile_X4Y4_RegFile/S4END[11]
+ Tile_X4Y4_RegFile/S4END[12] Tile_X4Y4_RegFile/S4END[13] Tile_X4Y4_RegFile/S4END[14]
+ Tile_X4Y4_RegFile/S4END[15] Tile_X4Y4_RegFile/S4END[1] Tile_X4Y4_RegFile/S4END[2]
+ Tile_X4Y4_RegFile/S4END[3] Tile_X4Y4_RegFile/S4END[4] Tile_X4Y4_RegFile/S4END[5]
+ Tile_X4Y4_RegFile/S4END[6] Tile_X4Y4_RegFile/S4END[7] Tile_X4Y4_RegFile/S4END[8]
+ Tile_X4Y4_RegFile/S4END[9] Tile_X4Y5_RegFile/SS4END[0] Tile_X4Y5_RegFile/SS4END[10]
+ Tile_X4Y5_RegFile/SS4END[11] Tile_X4Y5_RegFile/SS4END[12] Tile_X4Y5_RegFile/SS4END[13]
+ Tile_X4Y5_RegFile/SS4END[14] Tile_X4Y5_RegFile/SS4END[15] Tile_X4Y5_RegFile/SS4END[1]
+ Tile_X4Y5_RegFile/SS4END[2] Tile_X4Y5_RegFile/SS4END[3] Tile_X4Y5_RegFile/SS4END[4]
+ Tile_X4Y5_RegFile/SS4END[5] Tile_X4Y5_RegFile/SS4END[6] Tile_X4Y5_RegFile/SS4END[7]
+ Tile_X4Y5_RegFile/SS4END[8] Tile_X4Y5_RegFile/SS4END[9] Tile_X4Y4_RegFile/SS4END[0]
+ Tile_X4Y4_RegFile/SS4END[10] Tile_X4Y4_RegFile/SS4END[11] Tile_X4Y4_RegFile/SS4END[12]
+ Tile_X4Y4_RegFile/SS4END[13] Tile_X4Y4_RegFile/SS4END[14] Tile_X4Y4_RegFile/SS4END[15]
+ Tile_X4Y4_RegFile/SS4END[1] Tile_X4Y4_RegFile/SS4END[2] Tile_X4Y4_RegFile/SS4END[3]
+ Tile_X4Y4_RegFile/SS4END[4] Tile_X4Y4_RegFile/SS4END[5] Tile_X4Y4_RegFile/SS4END[6]
+ Tile_X4Y4_RegFile/SS4END[7] Tile_X4Y4_RegFile/SS4END[8] Tile_X4Y4_RegFile/SS4END[9]
+ Tile_X4Y4_RegFile/UserCLK Tile_X4Y3_RegFile/UserCLK VGND VPWR Tile_X3Y4_LUT4AB/W1END[0]
+ Tile_X3Y4_LUT4AB/W1END[1] Tile_X3Y4_LUT4AB/W1END[2] Tile_X3Y4_LUT4AB/W1END[3] Tile_X5Y4_LUT4AB/W1BEG[0]
+ Tile_X5Y4_LUT4AB/W1BEG[1] Tile_X5Y4_LUT4AB/W1BEG[2] Tile_X5Y4_LUT4AB/W1BEG[3] Tile_X3Y4_LUT4AB/W2MID[0]
+ Tile_X3Y4_LUT4AB/W2MID[1] Tile_X3Y4_LUT4AB/W2MID[2] Tile_X3Y4_LUT4AB/W2MID[3] Tile_X3Y4_LUT4AB/W2MID[4]
+ Tile_X3Y4_LUT4AB/W2MID[5] Tile_X3Y4_LUT4AB/W2MID[6] Tile_X3Y4_LUT4AB/W2MID[7] Tile_X3Y4_LUT4AB/W2END[0]
+ Tile_X3Y4_LUT4AB/W2END[1] Tile_X3Y4_LUT4AB/W2END[2] Tile_X3Y4_LUT4AB/W2END[3] Tile_X3Y4_LUT4AB/W2END[4]
+ Tile_X3Y4_LUT4AB/W2END[5] Tile_X3Y4_LUT4AB/W2END[6] Tile_X3Y4_LUT4AB/W2END[7] Tile_X5Y4_LUT4AB/W2BEGb[0]
+ Tile_X5Y4_LUT4AB/W2BEGb[1] Tile_X5Y4_LUT4AB/W2BEGb[2] Tile_X5Y4_LUT4AB/W2BEGb[3]
+ Tile_X5Y4_LUT4AB/W2BEGb[4] Tile_X5Y4_LUT4AB/W2BEGb[5] Tile_X5Y4_LUT4AB/W2BEGb[6]
+ Tile_X5Y4_LUT4AB/W2BEGb[7] Tile_X5Y4_LUT4AB/W2BEG[0] Tile_X5Y4_LUT4AB/W2BEG[1] Tile_X5Y4_LUT4AB/W2BEG[2]
+ Tile_X5Y4_LUT4AB/W2BEG[3] Tile_X5Y4_LUT4AB/W2BEG[4] Tile_X5Y4_LUT4AB/W2BEG[5] Tile_X5Y4_LUT4AB/W2BEG[6]
+ Tile_X5Y4_LUT4AB/W2BEG[7] Tile_X3Y4_LUT4AB/W6END[0] Tile_X3Y4_LUT4AB/W6END[10] Tile_X3Y4_LUT4AB/W6END[11]
+ Tile_X3Y4_LUT4AB/W6END[1] Tile_X3Y4_LUT4AB/W6END[2] Tile_X3Y4_LUT4AB/W6END[3] Tile_X3Y4_LUT4AB/W6END[4]
+ Tile_X3Y4_LUT4AB/W6END[5] Tile_X3Y4_LUT4AB/W6END[6] Tile_X3Y4_LUT4AB/W6END[7] Tile_X3Y4_LUT4AB/W6END[8]
+ Tile_X3Y4_LUT4AB/W6END[9] Tile_X5Y4_LUT4AB/W6BEG[0] Tile_X5Y4_LUT4AB/W6BEG[10] Tile_X5Y4_LUT4AB/W6BEG[11]
+ Tile_X5Y4_LUT4AB/W6BEG[1] Tile_X5Y4_LUT4AB/W6BEG[2] Tile_X5Y4_LUT4AB/W6BEG[3] Tile_X5Y4_LUT4AB/W6BEG[4]
+ Tile_X5Y4_LUT4AB/W6BEG[5] Tile_X5Y4_LUT4AB/W6BEG[6] Tile_X5Y4_LUT4AB/W6BEG[7] Tile_X5Y4_LUT4AB/W6BEG[8]
+ Tile_X5Y4_LUT4AB/W6BEG[9] Tile_X3Y4_LUT4AB/WW4END[0] Tile_X3Y4_LUT4AB/WW4END[10]
+ Tile_X3Y4_LUT4AB/WW4END[11] Tile_X3Y4_LUT4AB/WW4END[12] Tile_X3Y4_LUT4AB/WW4END[13]
+ Tile_X3Y4_LUT4AB/WW4END[14] Tile_X3Y4_LUT4AB/WW4END[15] Tile_X3Y4_LUT4AB/WW4END[1]
+ Tile_X3Y4_LUT4AB/WW4END[2] Tile_X3Y4_LUT4AB/WW4END[3] Tile_X3Y4_LUT4AB/WW4END[4]
+ Tile_X3Y4_LUT4AB/WW4END[5] Tile_X3Y4_LUT4AB/WW4END[6] Tile_X3Y4_LUT4AB/WW4END[7]
+ Tile_X3Y4_LUT4AB/WW4END[8] Tile_X3Y4_LUT4AB/WW4END[9] Tile_X5Y4_LUT4AB/WW4BEG[0]
+ Tile_X5Y4_LUT4AB/WW4BEG[10] Tile_X5Y4_LUT4AB/WW4BEG[11] Tile_X5Y4_LUT4AB/WW4BEG[12]
+ Tile_X5Y4_LUT4AB/WW4BEG[13] Tile_X5Y4_LUT4AB/WW4BEG[14] Tile_X5Y4_LUT4AB/WW4BEG[15]
+ Tile_X5Y4_LUT4AB/WW4BEG[1] Tile_X5Y4_LUT4AB/WW4BEG[2] Tile_X5Y4_LUT4AB/WW4BEG[3]
+ Tile_X5Y4_LUT4AB/WW4BEG[4] Tile_X5Y4_LUT4AB/WW4BEG[5] Tile_X5Y4_LUT4AB/WW4BEG[6]
+ Tile_X5Y4_LUT4AB/WW4BEG[7] Tile_X5Y4_LUT4AB/WW4BEG[8] Tile_X5Y4_LUT4AB/WW4BEG[9]
+ RegFile
XTile_X5Y5_LUT4AB Tile_X5Y6_LUT4AB/Co Tile_X5Y5_LUT4AB/Co Tile_X6Y5_LUT4AB/E1END[0]
+ Tile_X6Y5_LUT4AB/E1END[1] Tile_X6Y5_LUT4AB/E1END[2] Tile_X6Y5_LUT4AB/E1END[3] Tile_X5Y5_LUT4AB/E1END[0]
+ Tile_X5Y5_LUT4AB/E1END[1] Tile_X5Y5_LUT4AB/E1END[2] Tile_X5Y5_LUT4AB/E1END[3] Tile_X6Y5_LUT4AB/E2MID[0]
+ Tile_X6Y5_LUT4AB/E2MID[1] Tile_X6Y5_LUT4AB/E2MID[2] Tile_X6Y5_LUT4AB/E2MID[3] Tile_X6Y5_LUT4AB/E2MID[4]
+ Tile_X6Y5_LUT4AB/E2MID[5] Tile_X6Y5_LUT4AB/E2MID[6] Tile_X6Y5_LUT4AB/E2MID[7] Tile_X6Y5_LUT4AB/E2END[0]
+ Tile_X6Y5_LUT4AB/E2END[1] Tile_X6Y5_LUT4AB/E2END[2] Tile_X6Y5_LUT4AB/E2END[3] Tile_X6Y5_LUT4AB/E2END[4]
+ Tile_X6Y5_LUT4AB/E2END[5] Tile_X6Y5_LUT4AB/E2END[6] Tile_X6Y5_LUT4AB/E2END[7] Tile_X5Y5_LUT4AB/E2END[0]
+ Tile_X5Y5_LUT4AB/E2END[1] Tile_X5Y5_LUT4AB/E2END[2] Tile_X5Y5_LUT4AB/E2END[3] Tile_X5Y5_LUT4AB/E2END[4]
+ Tile_X5Y5_LUT4AB/E2END[5] Tile_X5Y5_LUT4AB/E2END[6] Tile_X5Y5_LUT4AB/E2END[7] Tile_X5Y5_LUT4AB/E2MID[0]
+ Tile_X5Y5_LUT4AB/E2MID[1] Tile_X5Y5_LUT4AB/E2MID[2] Tile_X5Y5_LUT4AB/E2MID[3] Tile_X5Y5_LUT4AB/E2MID[4]
+ Tile_X5Y5_LUT4AB/E2MID[5] Tile_X5Y5_LUT4AB/E2MID[6] Tile_X5Y5_LUT4AB/E2MID[7] Tile_X6Y5_LUT4AB/E6END[0]
+ Tile_X6Y5_LUT4AB/E6END[10] Tile_X6Y5_LUT4AB/E6END[11] Tile_X6Y5_LUT4AB/E6END[1]
+ Tile_X6Y5_LUT4AB/E6END[2] Tile_X6Y5_LUT4AB/E6END[3] Tile_X6Y5_LUT4AB/E6END[4] Tile_X6Y5_LUT4AB/E6END[5]
+ Tile_X6Y5_LUT4AB/E6END[6] Tile_X6Y5_LUT4AB/E6END[7] Tile_X6Y5_LUT4AB/E6END[8] Tile_X6Y5_LUT4AB/E6END[9]
+ Tile_X5Y5_LUT4AB/E6END[0] Tile_X5Y5_LUT4AB/E6END[10] Tile_X5Y5_LUT4AB/E6END[11]
+ Tile_X5Y5_LUT4AB/E6END[1] Tile_X5Y5_LUT4AB/E6END[2] Tile_X5Y5_LUT4AB/E6END[3] Tile_X5Y5_LUT4AB/E6END[4]
+ Tile_X5Y5_LUT4AB/E6END[5] Tile_X5Y5_LUT4AB/E6END[6] Tile_X5Y5_LUT4AB/E6END[7] Tile_X5Y5_LUT4AB/E6END[8]
+ Tile_X5Y5_LUT4AB/E6END[9] Tile_X6Y5_LUT4AB/EE4END[0] Tile_X6Y5_LUT4AB/EE4END[10]
+ Tile_X6Y5_LUT4AB/EE4END[11] Tile_X6Y5_LUT4AB/EE4END[12] Tile_X6Y5_LUT4AB/EE4END[13]
+ Tile_X6Y5_LUT4AB/EE4END[14] Tile_X6Y5_LUT4AB/EE4END[15] Tile_X6Y5_LUT4AB/EE4END[1]
+ Tile_X6Y5_LUT4AB/EE4END[2] Tile_X6Y5_LUT4AB/EE4END[3] Tile_X6Y5_LUT4AB/EE4END[4]
+ Tile_X6Y5_LUT4AB/EE4END[5] Tile_X6Y5_LUT4AB/EE4END[6] Tile_X6Y5_LUT4AB/EE4END[7]
+ Tile_X6Y5_LUT4AB/EE4END[8] Tile_X6Y5_LUT4AB/EE4END[9] Tile_X5Y5_LUT4AB/EE4END[0]
+ Tile_X5Y5_LUT4AB/EE4END[10] Tile_X5Y5_LUT4AB/EE4END[11] Tile_X5Y5_LUT4AB/EE4END[12]
+ Tile_X5Y5_LUT4AB/EE4END[13] Tile_X5Y5_LUT4AB/EE4END[14] Tile_X5Y5_LUT4AB/EE4END[15]
+ Tile_X5Y5_LUT4AB/EE4END[1] Tile_X5Y5_LUT4AB/EE4END[2] Tile_X5Y5_LUT4AB/EE4END[3]
+ Tile_X5Y5_LUT4AB/EE4END[4] Tile_X5Y5_LUT4AB/EE4END[5] Tile_X5Y5_LUT4AB/EE4END[6]
+ Tile_X5Y5_LUT4AB/EE4END[7] Tile_X5Y5_LUT4AB/EE4END[8] Tile_X5Y5_LUT4AB/EE4END[9]
+ Tile_X5Y5_LUT4AB/FrameData[0] Tile_X5Y5_LUT4AB/FrameData[10] Tile_X5Y5_LUT4AB/FrameData[11]
+ Tile_X5Y5_LUT4AB/FrameData[12] Tile_X5Y5_LUT4AB/FrameData[13] Tile_X5Y5_LUT4AB/FrameData[14]
+ Tile_X5Y5_LUT4AB/FrameData[15] Tile_X5Y5_LUT4AB/FrameData[16] Tile_X5Y5_LUT4AB/FrameData[17]
+ Tile_X5Y5_LUT4AB/FrameData[18] Tile_X5Y5_LUT4AB/FrameData[19] Tile_X5Y5_LUT4AB/FrameData[1]
+ Tile_X5Y5_LUT4AB/FrameData[20] Tile_X5Y5_LUT4AB/FrameData[21] Tile_X5Y5_LUT4AB/FrameData[22]
+ Tile_X5Y5_LUT4AB/FrameData[23] Tile_X5Y5_LUT4AB/FrameData[24] Tile_X5Y5_LUT4AB/FrameData[25]
+ Tile_X5Y5_LUT4AB/FrameData[26] Tile_X5Y5_LUT4AB/FrameData[27] Tile_X5Y5_LUT4AB/FrameData[28]
+ Tile_X5Y5_LUT4AB/FrameData[29] Tile_X5Y5_LUT4AB/FrameData[2] Tile_X5Y5_LUT4AB/FrameData[30]
+ Tile_X5Y5_LUT4AB/FrameData[31] Tile_X5Y5_LUT4AB/FrameData[3] Tile_X5Y5_LUT4AB/FrameData[4]
+ Tile_X5Y5_LUT4AB/FrameData[5] Tile_X5Y5_LUT4AB/FrameData[6] Tile_X5Y5_LUT4AB/FrameData[7]
+ Tile_X5Y5_LUT4AB/FrameData[8] Tile_X5Y5_LUT4AB/FrameData[9] Tile_X6Y5_LUT4AB/FrameData[0]
+ Tile_X6Y5_LUT4AB/FrameData[10] Tile_X6Y5_LUT4AB/FrameData[11] Tile_X6Y5_LUT4AB/FrameData[12]
+ Tile_X6Y5_LUT4AB/FrameData[13] Tile_X6Y5_LUT4AB/FrameData[14] Tile_X6Y5_LUT4AB/FrameData[15]
+ Tile_X6Y5_LUT4AB/FrameData[16] Tile_X6Y5_LUT4AB/FrameData[17] Tile_X6Y5_LUT4AB/FrameData[18]
+ Tile_X6Y5_LUT4AB/FrameData[19] Tile_X6Y5_LUT4AB/FrameData[1] Tile_X6Y5_LUT4AB/FrameData[20]
+ Tile_X6Y5_LUT4AB/FrameData[21] Tile_X6Y5_LUT4AB/FrameData[22] Tile_X6Y5_LUT4AB/FrameData[23]
+ Tile_X6Y5_LUT4AB/FrameData[24] Tile_X6Y5_LUT4AB/FrameData[25] Tile_X6Y5_LUT4AB/FrameData[26]
+ Tile_X6Y5_LUT4AB/FrameData[27] Tile_X6Y5_LUT4AB/FrameData[28] Tile_X6Y5_LUT4AB/FrameData[29]
+ Tile_X6Y5_LUT4AB/FrameData[2] Tile_X6Y5_LUT4AB/FrameData[30] Tile_X6Y5_LUT4AB/FrameData[31]
+ Tile_X6Y5_LUT4AB/FrameData[3] Tile_X6Y5_LUT4AB/FrameData[4] Tile_X6Y5_LUT4AB/FrameData[5]
+ Tile_X6Y5_LUT4AB/FrameData[6] Tile_X6Y5_LUT4AB/FrameData[7] Tile_X6Y5_LUT4AB/FrameData[8]
+ Tile_X6Y5_LUT4AB/FrameData[9] Tile_X5Y5_LUT4AB/FrameStrobe[0] Tile_X5Y5_LUT4AB/FrameStrobe[10]
+ Tile_X5Y5_LUT4AB/FrameStrobe[11] Tile_X5Y5_LUT4AB/FrameStrobe[12] Tile_X5Y5_LUT4AB/FrameStrobe[13]
+ Tile_X5Y5_LUT4AB/FrameStrobe[14] Tile_X5Y5_LUT4AB/FrameStrobe[15] Tile_X5Y5_LUT4AB/FrameStrobe[16]
+ Tile_X5Y5_LUT4AB/FrameStrobe[17] Tile_X5Y5_LUT4AB/FrameStrobe[18] Tile_X5Y5_LUT4AB/FrameStrobe[19]
+ Tile_X5Y5_LUT4AB/FrameStrobe[1] Tile_X5Y5_LUT4AB/FrameStrobe[2] Tile_X5Y5_LUT4AB/FrameStrobe[3]
+ Tile_X5Y5_LUT4AB/FrameStrobe[4] Tile_X5Y5_LUT4AB/FrameStrobe[5] Tile_X5Y5_LUT4AB/FrameStrobe[6]
+ Tile_X5Y5_LUT4AB/FrameStrobe[7] Tile_X5Y5_LUT4AB/FrameStrobe[8] Tile_X5Y5_LUT4AB/FrameStrobe[9]
+ Tile_X5Y4_LUT4AB/FrameStrobe[0] Tile_X5Y4_LUT4AB/FrameStrobe[10] Tile_X5Y4_LUT4AB/FrameStrobe[11]
+ Tile_X5Y4_LUT4AB/FrameStrobe[12] Tile_X5Y4_LUT4AB/FrameStrobe[13] Tile_X5Y4_LUT4AB/FrameStrobe[14]
+ Tile_X5Y4_LUT4AB/FrameStrobe[15] Tile_X5Y4_LUT4AB/FrameStrobe[16] Tile_X5Y4_LUT4AB/FrameStrobe[17]
+ Tile_X5Y4_LUT4AB/FrameStrobe[18] Tile_X5Y4_LUT4AB/FrameStrobe[19] Tile_X5Y4_LUT4AB/FrameStrobe[1]
+ Tile_X5Y4_LUT4AB/FrameStrobe[2] Tile_X5Y4_LUT4AB/FrameStrobe[3] Tile_X5Y4_LUT4AB/FrameStrobe[4]
+ Tile_X5Y4_LUT4AB/FrameStrobe[5] Tile_X5Y4_LUT4AB/FrameStrobe[6] Tile_X5Y4_LUT4AB/FrameStrobe[7]
+ Tile_X5Y4_LUT4AB/FrameStrobe[8] Tile_X5Y4_LUT4AB/FrameStrobe[9] Tile_X5Y5_LUT4AB/N1BEG[0]
+ Tile_X5Y5_LUT4AB/N1BEG[1] Tile_X5Y5_LUT4AB/N1BEG[2] Tile_X5Y5_LUT4AB/N1BEG[3] Tile_X5Y6_LUT4AB/N1BEG[0]
+ Tile_X5Y6_LUT4AB/N1BEG[1] Tile_X5Y6_LUT4AB/N1BEG[2] Tile_X5Y6_LUT4AB/N1BEG[3] Tile_X5Y5_LUT4AB/N2BEG[0]
+ Tile_X5Y5_LUT4AB/N2BEG[1] Tile_X5Y5_LUT4AB/N2BEG[2] Tile_X5Y5_LUT4AB/N2BEG[3] Tile_X5Y5_LUT4AB/N2BEG[4]
+ Tile_X5Y5_LUT4AB/N2BEG[5] Tile_X5Y5_LUT4AB/N2BEG[6] Tile_X5Y5_LUT4AB/N2BEG[7] Tile_X5Y4_LUT4AB/N2END[0]
+ Tile_X5Y4_LUT4AB/N2END[1] Tile_X5Y4_LUT4AB/N2END[2] Tile_X5Y4_LUT4AB/N2END[3] Tile_X5Y4_LUT4AB/N2END[4]
+ Tile_X5Y4_LUT4AB/N2END[5] Tile_X5Y4_LUT4AB/N2END[6] Tile_X5Y4_LUT4AB/N2END[7] Tile_X5Y5_LUT4AB/N2END[0]
+ Tile_X5Y5_LUT4AB/N2END[1] Tile_X5Y5_LUT4AB/N2END[2] Tile_X5Y5_LUT4AB/N2END[3] Tile_X5Y5_LUT4AB/N2END[4]
+ Tile_X5Y5_LUT4AB/N2END[5] Tile_X5Y5_LUT4AB/N2END[6] Tile_X5Y5_LUT4AB/N2END[7] Tile_X5Y6_LUT4AB/N2BEG[0]
+ Tile_X5Y6_LUT4AB/N2BEG[1] Tile_X5Y6_LUT4AB/N2BEG[2] Tile_X5Y6_LUT4AB/N2BEG[3] Tile_X5Y6_LUT4AB/N2BEG[4]
+ Tile_X5Y6_LUT4AB/N2BEG[5] Tile_X5Y6_LUT4AB/N2BEG[6] Tile_X5Y6_LUT4AB/N2BEG[7] Tile_X5Y5_LUT4AB/N4BEG[0]
+ Tile_X5Y5_LUT4AB/N4BEG[10] Tile_X5Y5_LUT4AB/N4BEG[11] Tile_X5Y5_LUT4AB/N4BEG[12]
+ Tile_X5Y5_LUT4AB/N4BEG[13] Tile_X5Y5_LUT4AB/N4BEG[14] Tile_X5Y5_LUT4AB/N4BEG[15]
+ Tile_X5Y5_LUT4AB/N4BEG[1] Tile_X5Y5_LUT4AB/N4BEG[2] Tile_X5Y5_LUT4AB/N4BEG[3] Tile_X5Y5_LUT4AB/N4BEG[4]
+ Tile_X5Y5_LUT4AB/N4BEG[5] Tile_X5Y5_LUT4AB/N4BEG[6] Tile_X5Y5_LUT4AB/N4BEG[7] Tile_X5Y5_LUT4AB/N4BEG[8]
+ Tile_X5Y5_LUT4AB/N4BEG[9] Tile_X5Y6_LUT4AB/N4BEG[0] Tile_X5Y6_LUT4AB/N4BEG[10] Tile_X5Y6_LUT4AB/N4BEG[11]
+ Tile_X5Y6_LUT4AB/N4BEG[12] Tile_X5Y6_LUT4AB/N4BEG[13] Tile_X5Y6_LUT4AB/N4BEG[14]
+ Tile_X5Y6_LUT4AB/N4BEG[15] Tile_X5Y6_LUT4AB/N4BEG[1] Tile_X5Y6_LUT4AB/N4BEG[2] Tile_X5Y6_LUT4AB/N4BEG[3]
+ Tile_X5Y6_LUT4AB/N4BEG[4] Tile_X5Y6_LUT4AB/N4BEG[5] Tile_X5Y6_LUT4AB/N4BEG[6] Tile_X5Y6_LUT4AB/N4BEG[7]
+ Tile_X5Y6_LUT4AB/N4BEG[8] Tile_X5Y6_LUT4AB/N4BEG[9] Tile_X5Y5_LUT4AB/NN4BEG[0] Tile_X5Y5_LUT4AB/NN4BEG[10]
+ Tile_X5Y5_LUT4AB/NN4BEG[11] Tile_X5Y5_LUT4AB/NN4BEG[12] Tile_X5Y5_LUT4AB/NN4BEG[13]
+ Tile_X5Y5_LUT4AB/NN4BEG[14] Tile_X5Y5_LUT4AB/NN4BEG[15] Tile_X5Y5_LUT4AB/NN4BEG[1]
+ Tile_X5Y5_LUT4AB/NN4BEG[2] Tile_X5Y5_LUT4AB/NN4BEG[3] Tile_X5Y5_LUT4AB/NN4BEG[4]
+ Tile_X5Y5_LUT4AB/NN4BEG[5] Tile_X5Y5_LUT4AB/NN4BEG[6] Tile_X5Y5_LUT4AB/NN4BEG[7]
+ Tile_X5Y5_LUT4AB/NN4BEG[8] Tile_X5Y5_LUT4AB/NN4BEG[9] Tile_X5Y6_LUT4AB/NN4BEG[0]
+ Tile_X5Y6_LUT4AB/NN4BEG[10] Tile_X5Y6_LUT4AB/NN4BEG[11] Tile_X5Y6_LUT4AB/NN4BEG[12]
+ Tile_X5Y6_LUT4AB/NN4BEG[13] Tile_X5Y6_LUT4AB/NN4BEG[14] Tile_X5Y6_LUT4AB/NN4BEG[15]
+ Tile_X5Y6_LUT4AB/NN4BEG[1] Tile_X5Y6_LUT4AB/NN4BEG[2] Tile_X5Y6_LUT4AB/NN4BEG[3]
+ Tile_X5Y6_LUT4AB/NN4BEG[4] Tile_X5Y6_LUT4AB/NN4BEG[5] Tile_X5Y6_LUT4AB/NN4BEG[6]
+ Tile_X5Y6_LUT4AB/NN4BEG[7] Tile_X5Y6_LUT4AB/NN4BEG[8] Tile_X5Y6_LUT4AB/NN4BEG[9]
+ Tile_X5Y6_LUT4AB/S1END[0] Tile_X5Y6_LUT4AB/S1END[1] Tile_X5Y6_LUT4AB/S1END[2] Tile_X5Y6_LUT4AB/S1END[3]
+ Tile_X5Y5_LUT4AB/S1END[0] Tile_X5Y5_LUT4AB/S1END[1] Tile_X5Y5_LUT4AB/S1END[2] Tile_X5Y5_LUT4AB/S1END[3]
+ Tile_X5Y6_LUT4AB/S2MID[0] Tile_X5Y6_LUT4AB/S2MID[1] Tile_X5Y6_LUT4AB/S2MID[2] Tile_X5Y6_LUT4AB/S2MID[3]
+ Tile_X5Y6_LUT4AB/S2MID[4] Tile_X5Y6_LUT4AB/S2MID[5] Tile_X5Y6_LUT4AB/S2MID[6] Tile_X5Y6_LUT4AB/S2MID[7]
+ Tile_X5Y6_LUT4AB/S2END[0] Tile_X5Y6_LUT4AB/S2END[1] Tile_X5Y6_LUT4AB/S2END[2] Tile_X5Y6_LUT4AB/S2END[3]
+ Tile_X5Y6_LUT4AB/S2END[4] Tile_X5Y6_LUT4AB/S2END[5] Tile_X5Y6_LUT4AB/S2END[6] Tile_X5Y6_LUT4AB/S2END[7]
+ Tile_X5Y5_LUT4AB/S2END[0] Tile_X5Y5_LUT4AB/S2END[1] Tile_X5Y5_LUT4AB/S2END[2] Tile_X5Y5_LUT4AB/S2END[3]
+ Tile_X5Y5_LUT4AB/S2END[4] Tile_X5Y5_LUT4AB/S2END[5] Tile_X5Y5_LUT4AB/S2END[6] Tile_X5Y5_LUT4AB/S2END[7]
+ Tile_X5Y5_LUT4AB/S2MID[0] Tile_X5Y5_LUT4AB/S2MID[1] Tile_X5Y5_LUT4AB/S2MID[2] Tile_X5Y5_LUT4AB/S2MID[3]
+ Tile_X5Y5_LUT4AB/S2MID[4] Tile_X5Y5_LUT4AB/S2MID[5] Tile_X5Y5_LUT4AB/S2MID[6] Tile_X5Y5_LUT4AB/S2MID[7]
+ Tile_X5Y6_LUT4AB/S4END[0] Tile_X5Y6_LUT4AB/S4END[10] Tile_X5Y6_LUT4AB/S4END[11]
+ Tile_X5Y6_LUT4AB/S4END[12] Tile_X5Y6_LUT4AB/S4END[13] Tile_X5Y6_LUT4AB/S4END[14]
+ Tile_X5Y6_LUT4AB/S4END[15] Tile_X5Y6_LUT4AB/S4END[1] Tile_X5Y6_LUT4AB/S4END[2] Tile_X5Y6_LUT4AB/S4END[3]
+ Tile_X5Y6_LUT4AB/S4END[4] Tile_X5Y6_LUT4AB/S4END[5] Tile_X5Y6_LUT4AB/S4END[6] Tile_X5Y6_LUT4AB/S4END[7]
+ Tile_X5Y6_LUT4AB/S4END[8] Tile_X5Y6_LUT4AB/S4END[9] Tile_X5Y5_LUT4AB/S4END[0] Tile_X5Y5_LUT4AB/S4END[10]
+ Tile_X5Y5_LUT4AB/S4END[11] Tile_X5Y5_LUT4AB/S4END[12] Tile_X5Y5_LUT4AB/S4END[13]
+ Tile_X5Y5_LUT4AB/S4END[14] Tile_X5Y5_LUT4AB/S4END[15] Tile_X5Y5_LUT4AB/S4END[1]
+ Tile_X5Y5_LUT4AB/S4END[2] Tile_X5Y5_LUT4AB/S4END[3] Tile_X5Y5_LUT4AB/S4END[4] Tile_X5Y5_LUT4AB/S4END[5]
+ Tile_X5Y5_LUT4AB/S4END[6] Tile_X5Y5_LUT4AB/S4END[7] Tile_X5Y5_LUT4AB/S4END[8] Tile_X5Y5_LUT4AB/S4END[9]
+ Tile_X5Y6_LUT4AB/SS4END[0] Tile_X5Y6_LUT4AB/SS4END[10] Tile_X5Y6_LUT4AB/SS4END[11]
+ Tile_X5Y6_LUT4AB/SS4END[12] Tile_X5Y6_LUT4AB/SS4END[13] Tile_X5Y6_LUT4AB/SS4END[14]
+ Tile_X5Y6_LUT4AB/SS4END[15] Tile_X5Y6_LUT4AB/SS4END[1] Tile_X5Y6_LUT4AB/SS4END[2]
+ Tile_X5Y6_LUT4AB/SS4END[3] Tile_X5Y6_LUT4AB/SS4END[4] Tile_X5Y6_LUT4AB/SS4END[5]
+ Tile_X5Y6_LUT4AB/SS4END[6] Tile_X5Y6_LUT4AB/SS4END[7] Tile_X5Y6_LUT4AB/SS4END[8]
+ Tile_X5Y6_LUT4AB/SS4END[9] Tile_X5Y5_LUT4AB/SS4END[0] Tile_X5Y5_LUT4AB/SS4END[10]
+ Tile_X5Y5_LUT4AB/SS4END[11] Tile_X5Y5_LUT4AB/SS4END[12] Tile_X5Y5_LUT4AB/SS4END[13]
+ Tile_X5Y5_LUT4AB/SS4END[14] Tile_X5Y5_LUT4AB/SS4END[15] Tile_X5Y5_LUT4AB/SS4END[1]
+ Tile_X5Y5_LUT4AB/SS4END[2] Tile_X5Y5_LUT4AB/SS4END[3] Tile_X5Y5_LUT4AB/SS4END[4]
+ Tile_X5Y5_LUT4AB/SS4END[5] Tile_X5Y5_LUT4AB/SS4END[6] Tile_X5Y5_LUT4AB/SS4END[7]
+ Tile_X5Y5_LUT4AB/SS4END[8] Tile_X5Y5_LUT4AB/SS4END[9] Tile_X5Y5_LUT4AB/UserCLK Tile_X5Y4_LUT4AB/UserCLK
+ VGND VPWR Tile_X5Y5_LUT4AB/W1BEG[0] Tile_X5Y5_LUT4AB/W1BEG[1] Tile_X5Y5_LUT4AB/W1BEG[2]
+ Tile_X5Y5_LUT4AB/W1BEG[3] Tile_X6Y5_LUT4AB/W1BEG[0] Tile_X6Y5_LUT4AB/W1BEG[1] Tile_X6Y5_LUT4AB/W1BEG[2]
+ Tile_X6Y5_LUT4AB/W1BEG[3] Tile_X5Y5_LUT4AB/W2BEG[0] Tile_X5Y5_LUT4AB/W2BEG[1] Tile_X5Y5_LUT4AB/W2BEG[2]
+ Tile_X5Y5_LUT4AB/W2BEG[3] Tile_X5Y5_LUT4AB/W2BEG[4] Tile_X5Y5_LUT4AB/W2BEG[5] Tile_X5Y5_LUT4AB/W2BEG[6]
+ Tile_X5Y5_LUT4AB/W2BEG[7] Tile_X5Y5_LUT4AB/W2BEGb[0] Tile_X5Y5_LUT4AB/W2BEGb[1]
+ Tile_X5Y5_LUT4AB/W2BEGb[2] Tile_X5Y5_LUT4AB/W2BEGb[3] Tile_X5Y5_LUT4AB/W2BEGb[4]
+ Tile_X5Y5_LUT4AB/W2BEGb[5] Tile_X5Y5_LUT4AB/W2BEGb[6] Tile_X5Y5_LUT4AB/W2BEGb[7]
+ Tile_X5Y5_LUT4AB/W2END[0] Tile_X5Y5_LUT4AB/W2END[1] Tile_X5Y5_LUT4AB/W2END[2] Tile_X5Y5_LUT4AB/W2END[3]
+ Tile_X5Y5_LUT4AB/W2END[4] Tile_X5Y5_LUT4AB/W2END[5] Tile_X5Y5_LUT4AB/W2END[6] Tile_X5Y5_LUT4AB/W2END[7]
+ Tile_X6Y5_LUT4AB/W2BEG[0] Tile_X6Y5_LUT4AB/W2BEG[1] Tile_X6Y5_LUT4AB/W2BEG[2] Tile_X6Y5_LUT4AB/W2BEG[3]
+ Tile_X6Y5_LUT4AB/W2BEG[4] Tile_X6Y5_LUT4AB/W2BEG[5] Tile_X6Y5_LUT4AB/W2BEG[6] Tile_X6Y5_LUT4AB/W2BEG[7]
+ Tile_X5Y5_LUT4AB/W6BEG[0] Tile_X5Y5_LUT4AB/W6BEG[10] Tile_X5Y5_LUT4AB/W6BEG[11]
+ Tile_X5Y5_LUT4AB/W6BEG[1] Tile_X5Y5_LUT4AB/W6BEG[2] Tile_X5Y5_LUT4AB/W6BEG[3] Tile_X5Y5_LUT4AB/W6BEG[4]
+ Tile_X5Y5_LUT4AB/W6BEG[5] Tile_X5Y5_LUT4AB/W6BEG[6] Tile_X5Y5_LUT4AB/W6BEG[7] Tile_X5Y5_LUT4AB/W6BEG[8]
+ Tile_X5Y5_LUT4AB/W6BEG[9] Tile_X6Y5_LUT4AB/W6BEG[0] Tile_X6Y5_LUT4AB/W6BEG[10] Tile_X6Y5_LUT4AB/W6BEG[11]
+ Tile_X6Y5_LUT4AB/W6BEG[1] Tile_X6Y5_LUT4AB/W6BEG[2] Tile_X6Y5_LUT4AB/W6BEG[3] Tile_X6Y5_LUT4AB/W6BEG[4]
+ Tile_X6Y5_LUT4AB/W6BEG[5] Tile_X6Y5_LUT4AB/W6BEG[6] Tile_X6Y5_LUT4AB/W6BEG[7] Tile_X6Y5_LUT4AB/W6BEG[8]
+ Tile_X6Y5_LUT4AB/W6BEG[9] Tile_X5Y5_LUT4AB/WW4BEG[0] Tile_X5Y5_LUT4AB/WW4BEG[10]
+ Tile_X5Y5_LUT4AB/WW4BEG[11] Tile_X5Y5_LUT4AB/WW4BEG[12] Tile_X5Y5_LUT4AB/WW4BEG[13]
+ Tile_X5Y5_LUT4AB/WW4BEG[14] Tile_X5Y5_LUT4AB/WW4BEG[15] Tile_X5Y5_LUT4AB/WW4BEG[1]
+ Tile_X5Y5_LUT4AB/WW4BEG[2] Tile_X5Y5_LUT4AB/WW4BEG[3] Tile_X5Y5_LUT4AB/WW4BEG[4]
+ Tile_X5Y5_LUT4AB/WW4BEG[5] Tile_X5Y5_LUT4AB/WW4BEG[6] Tile_X5Y5_LUT4AB/WW4BEG[7]
+ Tile_X5Y5_LUT4AB/WW4BEG[8] Tile_X5Y5_LUT4AB/WW4BEG[9] Tile_X6Y5_LUT4AB/WW4BEG[0]
+ Tile_X6Y5_LUT4AB/WW4BEG[10] Tile_X6Y5_LUT4AB/WW4BEG[11] Tile_X6Y5_LUT4AB/WW4BEG[12]
+ Tile_X6Y5_LUT4AB/WW4BEG[13] Tile_X6Y5_LUT4AB/WW4BEG[14] Tile_X6Y5_LUT4AB/WW4BEG[15]
+ Tile_X6Y5_LUT4AB/WW4BEG[1] Tile_X6Y5_LUT4AB/WW4BEG[2] Tile_X6Y5_LUT4AB/WW4BEG[3]
+ Tile_X6Y5_LUT4AB/WW4BEG[4] Tile_X6Y5_LUT4AB/WW4BEG[5] Tile_X6Y5_LUT4AB/WW4BEG[6]
+ Tile_X6Y5_LUT4AB/WW4BEG[7] Tile_X6Y5_LUT4AB/WW4BEG[8] Tile_X6Y5_LUT4AB/WW4BEG[9]
+ LUT4AB
XTile_X8Y15_S_CPU_IF Tile_X8Y14_LUT4AB/Ci Tile_X8Y15_S_CPU_IF/FrameData[0] Tile_X8Y15_S_CPU_IF/FrameData[10]
+ Tile_X8Y15_S_CPU_IF/FrameData[11] Tile_X8Y15_S_CPU_IF/FrameData[12] Tile_X8Y15_S_CPU_IF/FrameData[13]
+ Tile_X8Y15_S_CPU_IF/FrameData[14] Tile_X8Y15_S_CPU_IF/FrameData[15] Tile_X8Y15_S_CPU_IF/FrameData[16]
+ Tile_X8Y15_S_CPU_IF/FrameData[17] Tile_X8Y15_S_CPU_IF/FrameData[18] Tile_X8Y15_S_CPU_IF/FrameData[19]
+ Tile_X8Y15_S_CPU_IF/FrameData[1] Tile_X8Y15_S_CPU_IF/FrameData[20] Tile_X8Y15_S_CPU_IF/FrameData[21]
+ Tile_X8Y15_S_CPU_IF/FrameData[22] Tile_X8Y15_S_CPU_IF/FrameData[23] Tile_X8Y15_S_CPU_IF/FrameData[24]
+ Tile_X8Y15_S_CPU_IF/FrameData[25] Tile_X8Y15_S_CPU_IF/FrameData[26] Tile_X8Y15_S_CPU_IF/FrameData[27]
+ Tile_X8Y15_S_CPU_IF/FrameData[28] Tile_X8Y15_S_CPU_IF/FrameData[29] Tile_X8Y15_S_CPU_IF/FrameData[2]
+ Tile_X8Y15_S_CPU_IF/FrameData[30] Tile_X8Y15_S_CPU_IF/FrameData[31] Tile_X8Y15_S_CPU_IF/FrameData[3]
+ Tile_X8Y15_S_CPU_IF/FrameData[4] Tile_X8Y15_S_CPU_IF/FrameData[5] Tile_X8Y15_S_CPU_IF/FrameData[6]
+ Tile_X8Y15_S_CPU_IF/FrameData[7] Tile_X8Y15_S_CPU_IF/FrameData[8] Tile_X8Y15_S_CPU_IF/FrameData[9]
+ Tile_X9Y15_S_CPU_IF/FrameData[0] Tile_X9Y15_S_CPU_IF/FrameData[10] Tile_X9Y15_S_CPU_IF/FrameData[11]
+ Tile_X9Y15_S_CPU_IF/FrameData[12] Tile_X9Y15_S_CPU_IF/FrameData[13] Tile_X9Y15_S_CPU_IF/FrameData[14]
+ Tile_X9Y15_S_CPU_IF/FrameData[15] Tile_X9Y15_S_CPU_IF/FrameData[16] Tile_X9Y15_S_CPU_IF/FrameData[17]
+ Tile_X9Y15_S_CPU_IF/FrameData[18] Tile_X9Y15_S_CPU_IF/FrameData[19] Tile_X9Y15_S_CPU_IF/FrameData[1]
+ Tile_X9Y15_S_CPU_IF/FrameData[20] Tile_X9Y15_S_CPU_IF/FrameData[21] Tile_X9Y15_S_CPU_IF/FrameData[22]
+ Tile_X9Y15_S_CPU_IF/FrameData[23] Tile_X9Y15_S_CPU_IF/FrameData[24] Tile_X9Y15_S_CPU_IF/FrameData[25]
+ Tile_X9Y15_S_CPU_IF/FrameData[26] Tile_X9Y15_S_CPU_IF/FrameData[27] Tile_X9Y15_S_CPU_IF/FrameData[28]
+ Tile_X9Y15_S_CPU_IF/FrameData[29] Tile_X9Y15_S_CPU_IF/FrameData[2] Tile_X9Y15_S_CPU_IF/FrameData[30]
+ Tile_X9Y15_S_CPU_IF/FrameData[31] Tile_X9Y15_S_CPU_IF/FrameData[3] Tile_X9Y15_S_CPU_IF/FrameData[4]
+ Tile_X9Y15_S_CPU_IF/FrameData[5] Tile_X9Y15_S_CPU_IF/FrameData[6] Tile_X9Y15_S_CPU_IF/FrameData[7]
+ Tile_X9Y15_S_CPU_IF/FrameData[8] Tile_X9Y15_S_CPU_IF/FrameData[9] FrameStrobe[160]
+ FrameStrobe[170] FrameStrobe[171] FrameStrobe[172] FrameStrobe[173] FrameStrobe[174]
+ FrameStrobe[175] FrameStrobe[176] FrameStrobe[177] FrameStrobe[178] FrameStrobe[179]
+ FrameStrobe[161] FrameStrobe[162] FrameStrobe[163] FrameStrobe[164] FrameStrobe[165]
+ FrameStrobe[166] FrameStrobe[167] FrameStrobe[168] FrameStrobe[169] Tile_X8Y14_LUT4AB/FrameStrobe[0]
+ Tile_X8Y14_LUT4AB/FrameStrobe[10] Tile_X8Y14_LUT4AB/FrameStrobe[11] Tile_X8Y14_LUT4AB/FrameStrobe[12]
+ Tile_X8Y14_LUT4AB/FrameStrobe[13] Tile_X8Y14_LUT4AB/FrameStrobe[14] Tile_X8Y14_LUT4AB/FrameStrobe[15]
+ Tile_X8Y14_LUT4AB/FrameStrobe[16] Tile_X8Y14_LUT4AB/FrameStrobe[17] Tile_X8Y14_LUT4AB/FrameStrobe[18]
+ Tile_X8Y14_LUT4AB/FrameStrobe[19] Tile_X8Y14_LUT4AB/FrameStrobe[1] Tile_X8Y14_LUT4AB/FrameStrobe[2]
+ Tile_X8Y14_LUT4AB/FrameStrobe[3] Tile_X8Y14_LUT4AB/FrameStrobe[4] Tile_X8Y14_LUT4AB/FrameStrobe[5]
+ Tile_X8Y14_LUT4AB/FrameStrobe[6] Tile_X8Y14_LUT4AB/FrameStrobe[7] Tile_X8Y14_LUT4AB/FrameStrobe[8]
+ Tile_X8Y14_LUT4AB/FrameStrobe[9] Tile_X8Y15_I_top0 Tile_X8Y15_I_top1 Tile_X8Y15_I_top10
+ Tile_X8Y15_I_top11 Tile_X8Y15_I_top12 Tile_X8Y15_I_top13 Tile_X8Y15_I_top14 Tile_X8Y15_I_top15
+ Tile_X8Y15_I_top2 Tile_X8Y15_I_top3 Tile_X8Y15_I_top4 Tile_X8Y15_I_top5 Tile_X8Y15_I_top6
+ Tile_X8Y15_I_top7 Tile_X8Y15_I_top8 Tile_X8Y15_I_top9 Tile_X8Y14_LUT4AB/N1END[0]
+ Tile_X8Y14_LUT4AB/N1END[1] Tile_X8Y14_LUT4AB/N1END[2] Tile_X8Y14_LUT4AB/N1END[3]
+ Tile_X8Y14_LUT4AB/N2MID[0] Tile_X8Y14_LUT4AB/N2MID[1] Tile_X8Y14_LUT4AB/N2MID[2]
+ Tile_X8Y14_LUT4AB/N2MID[3] Tile_X8Y14_LUT4AB/N2MID[4] Tile_X8Y14_LUT4AB/N2MID[5]
+ Tile_X8Y14_LUT4AB/N2MID[6] Tile_X8Y14_LUT4AB/N2MID[7] Tile_X8Y14_LUT4AB/N2END[0]
+ Tile_X8Y14_LUT4AB/N2END[1] Tile_X8Y14_LUT4AB/N2END[2] Tile_X8Y14_LUT4AB/N2END[3]
+ Tile_X8Y14_LUT4AB/N2END[4] Tile_X8Y14_LUT4AB/N2END[5] Tile_X8Y14_LUT4AB/N2END[6]
+ Tile_X8Y14_LUT4AB/N2END[7] Tile_X8Y14_LUT4AB/N4END[0] Tile_X8Y14_LUT4AB/N4END[10]
+ Tile_X8Y14_LUT4AB/N4END[11] Tile_X8Y14_LUT4AB/N4END[12] Tile_X8Y14_LUT4AB/N4END[13]
+ Tile_X8Y14_LUT4AB/N4END[14] Tile_X8Y14_LUT4AB/N4END[15] Tile_X8Y14_LUT4AB/N4END[1]
+ Tile_X8Y14_LUT4AB/N4END[2] Tile_X8Y14_LUT4AB/N4END[3] Tile_X8Y14_LUT4AB/N4END[4]
+ Tile_X8Y14_LUT4AB/N4END[5] Tile_X8Y14_LUT4AB/N4END[6] Tile_X8Y14_LUT4AB/N4END[7]
+ Tile_X8Y14_LUT4AB/N4END[8] Tile_X8Y14_LUT4AB/N4END[9] Tile_X8Y14_LUT4AB/NN4END[0]
+ Tile_X8Y14_LUT4AB/NN4END[10] Tile_X8Y14_LUT4AB/NN4END[11] Tile_X8Y14_LUT4AB/NN4END[12]
+ Tile_X8Y14_LUT4AB/NN4END[13] Tile_X8Y14_LUT4AB/NN4END[14] Tile_X8Y14_LUT4AB/NN4END[15]
+ Tile_X8Y14_LUT4AB/NN4END[1] Tile_X8Y14_LUT4AB/NN4END[2] Tile_X8Y14_LUT4AB/NN4END[3]
+ Tile_X8Y14_LUT4AB/NN4END[4] Tile_X8Y14_LUT4AB/NN4END[5] Tile_X8Y14_LUT4AB/NN4END[6]
+ Tile_X8Y14_LUT4AB/NN4END[7] Tile_X8Y14_LUT4AB/NN4END[8] Tile_X8Y14_LUT4AB/NN4END[9]
+ Tile_X8Y15_O_top0 Tile_X8Y15_O_top1 Tile_X8Y15_O_top10 Tile_X8Y15_O_top11 Tile_X8Y15_O_top12
+ Tile_X8Y15_O_top13 Tile_X8Y15_O_top14 Tile_X8Y15_O_top15 Tile_X8Y15_O_top2 Tile_X8Y15_O_top3
+ Tile_X8Y15_O_top4 Tile_X8Y15_O_top5 Tile_X8Y15_O_top6 Tile_X8Y15_O_top7 Tile_X8Y15_O_top8
+ Tile_X8Y15_O_top9 Tile_X8Y14_LUT4AB/S1BEG[0] Tile_X8Y14_LUT4AB/S1BEG[1] Tile_X8Y14_LUT4AB/S1BEG[2]
+ Tile_X8Y14_LUT4AB/S1BEG[3] Tile_X8Y14_LUT4AB/S2BEGb[0] Tile_X8Y14_LUT4AB/S2BEGb[1]
+ Tile_X8Y14_LUT4AB/S2BEGb[2] Tile_X8Y14_LUT4AB/S2BEGb[3] Tile_X8Y14_LUT4AB/S2BEGb[4]
+ Tile_X8Y14_LUT4AB/S2BEGb[5] Tile_X8Y14_LUT4AB/S2BEGb[6] Tile_X8Y14_LUT4AB/S2BEGb[7]
+ Tile_X8Y14_LUT4AB/S2BEG[0] Tile_X8Y14_LUT4AB/S2BEG[1] Tile_X8Y14_LUT4AB/S2BEG[2]
+ Tile_X8Y14_LUT4AB/S2BEG[3] Tile_X8Y14_LUT4AB/S2BEG[4] Tile_X8Y14_LUT4AB/S2BEG[5]
+ Tile_X8Y14_LUT4AB/S2BEG[6] Tile_X8Y14_LUT4AB/S2BEG[7] Tile_X8Y14_LUT4AB/S4BEG[0]
+ Tile_X8Y14_LUT4AB/S4BEG[10] Tile_X8Y14_LUT4AB/S4BEG[11] Tile_X8Y14_LUT4AB/S4BEG[12]
+ Tile_X8Y14_LUT4AB/S4BEG[13] Tile_X8Y14_LUT4AB/S4BEG[14] Tile_X8Y14_LUT4AB/S4BEG[15]
+ Tile_X8Y14_LUT4AB/S4BEG[1] Tile_X8Y14_LUT4AB/S4BEG[2] Tile_X8Y14_LUT4AB/S4BEG[3]
+ Tile_X8Y14_LUT4AB/S4BEG[4] Tile_X8Y14_LUT4AB/S4BEG[5] Tile_X8Y14_LUT4AB/S4BEG[6]
+ Tile_X8Y14_LUT4AB/S4BEG[7] Tile_X8Y14_LUT4AB/S4BEG[8] Tile_X8Y14_LUT4AB/S4BEG[9]
+ Tile_X8Y14_LUT4AB/SS4BEG[0] Tile_X8Y14_LUT4AB/SS4BEG[10] Tile_X8Y14_LUT4AB/SS4BEG[11]
+ Tile_X8Y14_LUT4AB/SS4BEG[12] Tile_X8Y14_LUT4AB/SS4BEG[13] Tile_X8Y14_LUT4AB/SS4BEG[14]
+ Tile_X8Y14_LUT4AB/SS4BEG[15] Tile_X8Y14_LUT4AB/SS4BEG[1] Tile_X8Y14_LUT4AB/SS4BEG[2]
+ Tile_X8Y14_LUT4AB/SS4BEG[3] Tile_X8Y14_LUT4AB/SS4BEG[4] Tile_X8Y14_LUT4AB/SS4BEG[5]
+ Tile_X8Y14_LUT4AB/SS4BEG[6] Tile_X8Y14_LUT4AB/SS4BEG[7] Tile_X8Y14_LUT4AB/SS4BEG[8]
+ Tile_X8Y14_LUT4AB/SS4BEG[9] UserCLK Tile_X8Y14_LUT4AB/UserCLK VGND VPWR S_CPU_IF
XTile_X7Y9_DSP Tile_X8Y9_LUT4AB/E1END[0] Tile_X8Y9_LUT4AB/E1END[1] Tile_X8Y9_LUT4AB/E1END[2]
+ Tile_X8Y9_LUT4AB/E1END[3] Tile_X6Y9_LUT4AB/E1BEG[0] Tile_X6Y9_LUT4AB/E1BEG[1] Tile_X6Y9_LUT4AB/E1BEG[2]
+ Tile_X6Y9_LUT4AB/E1BEG[3] Tile_X8Y9_LUT4AB/E2MID[0] Tile_X8Y9_LUT4AB/E2MID[1] Tile_X8Y9_LUT4AB/E2MID[2]
+ Tile_X8Y9_LUT4AB/E2MID[3] Tile_X8Y9_LUT4AB/E2MID[4] Tile_X8Y9_LUT4AB/E2MID[5] Tile_X8Y9_LUT4AB/E2MID[6]
+ Tile_X8Y9_LUT4AB/E2MID[7] Tile_X8Y9_LUT4AB/E2END[0] Tile_X8Y9_LUT4AB/E2END[1] Tile_X8Y9_LUT4AB/E2END[2]
+ Tile_X8Y9_LUT4AB/E2END[3] Tile_X8Y9_LUT4AB/E2END[4] Tile_X8Y9_LUT4AB/E2END[5] Tile_X8Y9_LUT4AB/E2END[6]
+ Tile_X8Y9_LUT4AB/E2END[7] Tile_X6Y9_LUT4AB/E2BEGb[0] Tile_X6Y9_LUT4AB/E2BEGb[1]
+ Tile_X6Y9_LUT4AB/E2BEGb[2] Tile_X6Y9_LUT4AB/E2BEGb[3] Tile_X6Y9_LUT4AB/E2BEGb[4]
+ Tile_X6Y9_LUT4AB/E2BEGb[5] Tile_X6Y9_LUT4AB/E2BEGb[6] Tile_X6Y9_LUT4AB/E2BEGb[7]
+ Tile_X6Y9_LUT4AB/E2BEG[0] Tile_X6Y9_LUT4AB/E2BEG[1] Tile_X6Y9_LUT4AB/E2BEG[2] Tile_X6Y9_LUT4AB/E2BEG[3]
+ Tile_X6Y9_LUT4AB/E2BEG[4] Tile_X6Y9_LUT4AB/E2BEG[5] Tile_X6Y9_LUT4AB/E2BEG[6] Tile_X6Y9_LUT4AB/E2BEG[7]
+ Tile_X8Y9_LUT4AB/E6END[0] Tile_X8Y9_LUT4AB/E6END[10] Tile_X8Y9_LUT4AB/E6END[11]
+ Tile_X8Y9_LUT4AB/E6END[1] Tile_X8Y9_LUT4AB/E6END[2] Tile_X8Y9_LUT4AB/E6END[3] Tile_X8Y9_LUT4AB/E6END[4]
+ Tile_X8Y9_LUT4AB/E6END[5] Tile_X8Y9_LUT4AB/E6END[6] Tile_X8Y9_LUT4AB/E6END[7] Tile_X8Y9_LUT4AB/E6END[8]
+ Tile_X8Y9_LUT4AB/E6END[9] Tile_X6Y9_LUT4AB/E6BEG[0] Tile_X6Y9_LUT4AB/E6BEG[10] Tile_X6Y9_LUT4AB/E6BEG[11]
+ Tile_X6Y9_LUT4AB/E6BEG[1] Tile_X6Y9_LUT4AB/E6BEG[2] Tile_X6Y9_LUT4AB/E6BEG[3] Tile_X6Y9_LUT4AB/E6BEG[4]
+ Tile_X6Y9_LUT4AB/E6BEG[5] Tile_X6Y9_LUT4AB/E6BEG[6] Tile_X6Y9_LUT4AB/E6BEG[7] Tile_X6Y9_LUT4AB/E6BEG[8]
+ Tile_X6Y9_LUT4AB/E6BEG[9] Tile_X8Y9_LUT4AB/EE4END[0] Tile_X8Y9_LUT4AB/EE4END[10]
+ Tile_X8Y9_LUT4AB/EE4END[11] Tile_X8Y9_LUT4AB/EE4END[12] Tile_X8Y9_LUT4AB/EE4END[13]
+ Tile_X8Y9_LUT4AB/EE4END[14] Tile_X8Y9_LUT4AB/EE4END[15] Tile_X8Y9_LUT4AB/EE4END[1]
+ Tile_X8Y9_LUT4AB/EE4END[2] Tile_X8Y9_LUT4AB/EE4END[3] Tile_X8Y9_LUT4AB/EE4END[4]
+ Tile_X8Y9_LUT4AB/EE4END[5] Tile_X8Y9_LUT4AB/EE4END[6] Tile_X8Y9_LUT4AB/EE4END[7]
+ Tile_X8Y9_LUT4AB/EE4END[8] Tile_X8Y9_LUT4AB/EE4END[9] Tile_X6Y9_LUT4AB/EE4BEG[0]
+ Tile_X6Y9_LUT4AB/EE4BEG[10] Tile_X6Y9_LUT4AB/EE4BEG[11] Tile_X6Y9_LUT4AB/EE4BEG[12]
+ Tile_X6Y9_LUT4AB/EE4BEG[13] Tile_X6Y9_LUT4AB/EE4BEG[14] Tile_X6Y9_LUT4AB/EE4BEG[15]
+ Tile_X6Y9_LUT4AB/EE4BEG[1] Tile_X6Y9_LUT4AB/EE4BEG[2] Tile_X6Y9_LUT4AB/EE4BEG[3]
+ Tile_X6Y9_LUT4AB/EE4BEG[4] Tile_X6Y9_LUT4AB/EE4BEG[5] Tile_X6Y9_LUT4AB/EE4BEG[6]
+ Tile_X6Y9_LUT4AB/EE4BEG[7] Tile_X6Y9_LUT4AB/EE4BEG[8] Tile_X6Y9_LUT4AB/EE4BEG[9]
+ Tile_X6Y9_LUT4AB/FrameData_O[0] Tile_X6Y9_LUT4AB/FrameData_O[10] Tile_X6Y9_LUT4AB/FrameData_O[11]
+ Tile_X6Y9_LUT4AB/FrameData_O[12] Tile_X6Y9_LUT4AB/FrameData_O[13] Tile_X6Y9_LUT4AB/FrameData_O[14]
+ Tile_X6Y9_LUT4AB/FrameData_O[15] Tile_X6Y9_LUT4AB/FrameData_O[16] Tile_X6Y9_LUT4AB/FrameData_O[17]
+ Tile_X6Y9_LUT4AB/FrameData_O[18] Tile_X6Y9_LUT4AB/FrameData_O[19] Tile_X6Y9_LUT4AB/FrameData_O[1]
+ Tile_X6Y9_LUT4AB/FrameData_O[20] Tile_X6Y9_LUT4AB/FrameData_O[21] Tile_X6Y9_LUT4AB/FrameData_O[22]
+ Tile_X6Y9_LUT4AB/FrameData_O[23] Tile_X6Y9_LUT4AB/FrameData_O[24] Tile_X6Y9_LUT4AB/FrameData_O[25]
+ Tile_X6Y9_LUT4AB/FrameData_O[26] Tile_X6Y9_LUT4AB/FrameData_O[27] Tile_X6Y9_LUT4AB/FrameData_O[28]
+ Tile_X6Y9_LUT4AB/FrameData_O[29] Tile_X6Y9_LUT4AB/FrameData_O[2] Tile_X6Y9_LUT4AB/FrameData_O[30]
+ Tile_X6Y9_LUT4AB/FrameData_O[31] Tile_X6Y9_LUT4AB/FrameData_O[3] Tile_X6Y9_LUT4AB/FrameData_O[4]
+ Tile_X6Y9_LUT4AB/FrameData_O[5] Tile_X6Y9_LUT4AB/FrameData_O[6] Tile_X6Y9_LUT4AB/FrameData_O[7]
+ Tile_X6Y9_LUT4AB/FrameData_O[8] Tile_X6Y9_LUT4AB/FrameData_O[9] Tile_X8Y9_LUT4AB/FrameData[0]
+ Tile_X8Y9_LUT4AB/FrameData[10] Tile_X8Y9_LUT4AB/FrameData[11] Tile_X8Y9_LUT4AB/FrameData[12]
+ Tile_X8Y9_LUT4AB/FrameData[13] Tile_X8Y9_LUT4AB/FrameData[14] Tile_X8Y9_LUT4AB/FrameData[15]
+ Tile_X8Y9_LUT4AB/FrameData[16] Tile_X8Y9_LUT4AB/FrameData[17] Tile_X8Y9_LUT4AB/FrameData[18]
+ Tile_X8Y9_LUT4AB/FrameData[19] Tile_X8Y9_LUT4AB/FrameData[1] Tile_X8Y9_LUT4AB/FrameData[20]
+ Tile_X8Y9_LUT4AB/FrameData[21] Tile_X8Y9_LUT4AB/FrameData[22] Tile_X8Y9_LUT4AB/FrameData[23]
+ Tile_X8Y9_LUT4AB/FrameData[24] Tile_X8Y9_LUT4AB/FrameData[25] Tile_X8Y9_LUT4AB/FrameData[26]
+ Tile_X8Y9_LUT4AB/FrameData[27] Tile_X8Y9_LUT4AB/FrameData[28] Tile_X8Y9_LUT4AB/FrameData[29]
+ Tile_X8Y9_LUT4AB/FrameData[2] Tile_X8Y9_LUT4AB/FrameData[30] Tile_X8Y9_LUT4AB/FrameData[31]
+ Tile_X8Y9_LUT4AB/FrameData[3] Tile_X8Y9_LUT4AB/FrameData[4] Tile_X8Y9_LUT4AB/FrameData[5]
+ Tile_X8Y9_LUT4AB/FrameData[6] Tile_X8Y9_LUT4AB/FrameData[7] Tile_X8Y9_LUT4AB/FrameData[8]
+ Tile_X8Y9_LUT4AB/FrameData[9] Tile_X7Y7_DSP/Tile_X0Y1_FrameStrobe[0] Tile_X7Y7_DSP/Tile_X0Y1_FrameStrobe[10]
+ Tile_X7Y7_DSP/Tile_X0Y1_FrameStrobe[11] Tile_X7Y7_DSP/Tile_X0Y1_FrameStrobe[12]
+ Tile_X7Y7_DSP/Tile_X0Y1_FrameStrobe[13] Tile_X7Y7_DSP/Tile_X0Y1_FrameStrobe[14]
+ Tile_X7Y7_DSP/Tile_X0Y1_FrameStrobe[15] Tile_X7Y7_DSP/Tile_X0Y1_FrameStrobe[16]
+ Tile_X7Y7_DSP/Tile_X0Y1_FrameStrobe[17] Tile_X7Y7_DSP/Tile_X0Y1_FrameStrobe[18]
+ Tile_X7Y7_DSP/Tile_X0Y1_FrameStrobe[19] Tile_X7Y7_DSP/Tile_X0Y1_FrameStrobe[1] Tile_X7Y7_DSP/Tile_X0Y1_FrameStrobe[2]
+ Tile_X7Y7_DSP/Tile_X0Y1_FrameStrobe[3] Tile_X7Y7_DSP/Tile_X0Y1_FrameStrobe[4] Tile_X7Y7_DSP/Tile_X0Y1_FrameStrobe[5]
+ Tile_X7Y7_DSP/Tile_X0Y1_FrameStrobe[6] Tile_X7Y7_DSP/Tile_X0Y1_FrameStrobe[7] Tile_X7Y7_DSP/Tile_X0Y1_FrameStrobe[8]
+ Tile_X7Y7_DSP/Tile_X0Y1_FrameStrobe[9] Tile_X7Y9_DSP/Tile_X0Y0_N1BEG[0] Tile_X7Y9_DSP/Tile_X0Y0_N1BEG[1]
+ Tile_X7Y9_DSP/Tile_X0Y0_N1BEG[2] Tile_X7Y9_DSP/Tile_X0Y0_N1BEG[3] Tile_X7Y9_DSP/Tile_X0Y0_N2BEG[0]
+ Tile_X7Y9_DSP/Tile_X0Y0_N2BEG[1] Tile_X7Y9_DSP/Tile_X0Y0_N2BEG[2] Tile_X7Y9_DSP/Tile_X0Y0_N2BEG[3]
+ Tile_X7Y9_DSP/Tile_X0Y0_N2BEG[4] Tile_X7Y9_DSP/Tile_X0Y0_N2BEG[5] Tile_X7Y9_DSP/Tile_X0Y0_N2BEG[6]
+ Tile_X7Y9_DSP/Tile_X0Y0_N2BEG[7] Tile_X7Y7_DSP/Tile_X0Y1_N2END[0] Tile_X7Y7_DSP/Tile_X0Y1_N2END[1]
+ Tile_X7Y7_DSP/Tile_X0Y1_N2END[2] Tile_X7Y7_DSP/Tile_X0Y1_N2END[3] Tile_X7Y7_DSP/Tile_X0Y1_N2END[4]
+ Tile_X7Y7_DSP/Tile_X0Y1_N2END[5] Tile_X7Y7_DSP/Tile_X0Y1_N2END[6] Tile_X7Y7_DSP/Tile_X0Y1_N2END[7]
+ Tile_X7Y9_DSP/Tile_X0Y0_N4BEG[0] Tile_X7Y9_DSP/Tile_X0Y0_N4BEG[10] Tile_X7Y9_DSP/Tile_X0Y0_N4BEG[11]
+ Tile_X7Y9_DSP/Tile_X0Y0_N4BEG[12] Tile_X7Y9_DSP/Tile_X0Y0_N4BEG[13] Tile_X7Y9_DSP/Tile_X0Y0_N4BEG[14]
+ Tile_X7Y9_DSP/Tile_X0Y0_N4BEG[15] Tile_X7Y9_DSP/Tile_X0Y0_N4BEG[1] Tile_X7Y9_DSP/Tile_X0Y0_N4BEG[2]
+ Tile_X7Y9_DSP/Tile_X0Y0_N4BEG[3] Tile_X7Y9_DSP/Tile_X0Y0_N4BEG[4] Tile_X7Y9_DSP/Tile_X0Y0_N4BEG[5]
+ Tile_X7Y9_DSP/Tile_X0Y0_N4BEG[6] Tile_X7Y9_DSP/Tile_X0Y0_N4BEG[7] Tile_X7Y9_DSP/Tile_X0Y0_N4BEG[8]
+ Tile_X7Y9_DSP/Tile_X0Y0_N4BEG[9] Tile_X7Y9_DSP/Tile_X0Y0_NN4BEG[0] Tile_X7Y9_DSP/Tile_X0Y0_NN4BEG[10]
+ Tile_X7Y9_DSP/Tile_X0Y0_NN4BEG[11] Tile_X7Y9_DSP/Tile_X0Y0_NN4BEG[12] Tile_X7Y9_DSP/Tile_X0Y0_NN4BEG[13]
+ Tile_X7Y9_DSP/Tile_X0Y0_NN4BEG[14] Tile_X7Y9_DSP/Tile_X0Y0_NN4BEG[15] Tile_X7Y9_DSP/Tile_X0Y0_NN4BEG[1]
+ Tile_X7Y9_DSP/Tile_X0Y0_NN4BEG[2] Tile_X7Y9_DSP/Tile_X0Y0_NN4BEG[3] Tile_X7Y9_DSP/Tile_X0Y0_NN4BEG[4]
+ Tile_X7Y9_DSP/Tile_X0Y0_NN4BEG[5] Tile_X7Y9_DSP/Tile_X0Y0_NN4BEG[6] Tile_X7Y9_DSP/Tile_X0Y0_NN4BEG[7]
+ Tile_X7Y9_DSP/Tile_X0Y0_NN4BEG[8] Tile_X7Y9_DSP/Tile_X0Y0_NN4BEG[9] Tile_X7Y9_DSP/Tile_X0Y0_S1END[0]
+ Tile_X7Y9_DSP/Tile_X0Y0_S1END[1] Tile_X7Y9_DSP/Tile_X0Y0_S1END[2] Tile_X7Y9_DSP/Tile_X0Y0_S1END[3]
+ Tile_X7Y9_DSP/Tile_X0Y0_S2END[0] Tile_X7Y9_DSP/Tile_X0Y0_S2END[1] Tile_X7Y9_DSP/Tile_X0Y0_S2END[2]
+ Tile_X7Y9_DSP/Tile_X0Y0_S2END[3] Tile_X7Y9_DSP/Tile_X0Y0_S2END[4] Tile_X7Y9_DSP/Tile_X0Y0_S2END[5]
+ Tile_X7Y9_DSP/Tile_X0Y0_S2END[6] Tile_X7Y9_DSP/Tile_X0Y0_S2END[7] Tile_X7Y9_DSP/Tile_X0Y0_S2MID[0]
+ Tile_X7Y9_DSP/Tile_X0Y0_S2MID[1] Tile_X7Y9_DSP/Tile_X0Y0_S2MID[2] Tile_X7Y9_DSP/Tile_X0Y0_S2MID[3]
+ Tile_X7Y9_DSP/Tile_X0Y0_S2MID[4] Tile_X7Y9_DSP/Tile_X0Y0_S2MID[5] Tile_X7Y9_DSP/Tile_X0Y0_S2MID[6]
+ Tile_X7Y9_DSP/Tile_X0Y0_S2MID[7] Tile_X7Y9_DSP/Tile_X0Y0_S4END[0] Tile_X7Y9_DSP/Tile_X0Y0_S4END[10]
+ Tile_X7Y9_DSP/Tile_X0Y0_S4END[11] Tile_X7Y9_DSP/Tile_X0Y0_S4END[12] Tile_X7Y9_DSP/Tile_X0Y0_S4END[13]
+ Tile_X7Y9_DSP/Tile_X0Y0_S4END[14] Tile_X7Y9_DSP/Tile_X0Y0_S4END[15] Tile_X7Y9_DSP/Tile_X0Y0_S4END[1]
+ Tile_X7Y9_DSP/Tile_X0Y0_S4END[2] Tile_X7Y9_DSP/Tile_X0Y0_S4END[3] Tile_X7Y9_DSP/Tile_X0Y0_S4END[4]
+ Tile_X7Y9_DSP/Tile_X0Y0_S4END[5] Tile_X7Y9_DSP/Tile_X0Y0_S4END[6] Tile_X7Y9_DSP/Tile_X0Y0_S4END[7]
+ Tile_X7Y9_DSP/Tile_X0Y0_S4END[8] Tile_X7Y9_DSP/Tile_X0Y0_S4END[9] Tile_X7Y9_DSP/Tile_X0Y0_SS4END[0]
+ Tile_X7Y9_DSP/Tile_X0Y0_SS4END[10] Tile_X7Y9_DSP/Tile_X0Y0_SS4END[11] Tile_X7Y9_DSP/Tile_X0Y0_SS4END[12]
+ Tile_X7Y9_DSP/Tile_X0Y0_SS4END[13] Tile_X7Y9_DSP/Tile_X0Y0_SS4END[14] Tile_X7Y9_DSP/Tile_X0Y0_SS4END[15]
+ Tile_X7Y9_DSP/Tile_X0Y0_SS4END[1] Tile_X7Y9_DSP/Tile_X0Y0_SS4END[2] Tile_X7Y9_DSP/Tile_X0Y0_SS4END[3]
+ Tile_X7Y9_DSP/Tile_X0Y0_SS4END[4] Tile_X7Y9_DSP/Tile_X0Y0_SS4END[5] Tile_X7Y9_DSP/Tile_X0Y0_SS4END[6]
+ Tile_X7Y9_DSP/Tile_X0Y0_SS4END[7] Tile_X7Y9_DSP/Tile_X0Y0_SS4END[8] Tile_X7Y9_DSP/Tile_X0Y0_SS4END[9]
+ Tile_X7Y7_DSP/Tile_X0Y1_UserCLK Tile_X6Y9_LUT4AB/W1END[0] Tile_X6Y9_LUT4AB/W1END[1]
+ Tile_X6Y9_LUT4AB/W1END[2] Tile_X6Y9_LUT4AB/W1END[3] Tile_X8Y9_LUT4AB/W1BEG[0] Tile_X8Y9_LUT4AB/W1BEG[1]
+ Tile_X8Y9_LUT4AB/W1BEG[2] Tile_X8Y9_LUT4AB/W1BEG[3] Tile_X6Y9_LUT4AB/W2MID[0] Tile_X6Y9_LUT4AB/W2MID[1]
+ Tile_X6Y9_LUT4AB/W2MID[2] Tile_X6Y9_LUT4AB/W2MID[3] Tile_X6Y9_LUT4AB/W2MID[4] Tile_X6Y9_LUT4AB/W2MID[5]
+ Tile_X6Y9_LUT4AB/W2MID[6] Tile_X6Y9_LUT4AB/W2MID[7] Tile_X6Y9_LUT4AB/W2END[0] Tile_X6Y9_LUT4AB/W2END[1]
+ Tile_X6Y9_LUT4AB/W2END[2] Tile_X6Y9_LUT4AB/W2END[3] Tile_X6Y9_LUT4AB/W2END[4] Tile_X6Y9_LUT4AB/W2END[5]
+ Tile_X6Y9_LUT4AB/W2END[6] Tile_X6Y9_LUT4AB/W2END[7] Tile_X8Y9_LUT4AB/W2BEGb[0] Tile_X8Y9_LUT4AB/W2BEGb[1]
+ Tile_X8Y9_LUT4AB/W2BEGb[2] Tile_X8Y9_LUT4AB/W2BEGb[3] Tile_X8Y9_LUT4AB/W2BEGb[4]
+ Tile_X8Y9_LUT4AB/W2BEGb[5] Tile_X8Y9_LUT4AB/W2BEGb[6] Tile_X8Y9_LUT4AB/W2BEGb[7]
+ Tile_X8Y9_LUT4AB/W2BEG[0] Tile_X8Y9_LUT4AB/W2BEG[1] Tile_X8Y9_LUT4AB/W2BEG[2] Tile_X8Y9_LUT4AB/W2BEG[3]
+ Tile_X8Y9_LUT4AB/W2BEG[4] Tile_X8Y9_LUT4AB/W2BEG[5] Tile_X8Y9_LUT4AB/W2BEG[6] Tile_X8Y9_LUT4AB/W2BEG[7]
+ Tile_X6Y9_LUT4AB/W6END[0] Tile_X6Y9_LUT4AB/W6END[10] Tile_X6Y9_LUT4AB/W6END[11]
+ Tile_X6Y9_LUT4AB/W6END[1] Tile_X6Y9_LUT4AB/W6END[2] Tile_X6Y9_LUT4AB/W6END[3] Tile_X6Y9_LUT4AB/W6END[4]
+ Tile_X6Y9_LUT4AB/W6END[5] Tile_X6Y9_LUT4AB/W6END[6] Tile_X6Y9_LUT4AB/W6END[7] Tile_X6Y9_LUT4AB/W6END[8]
+ Tile_X6Y9_LUT4AB/W6END[9] Tile_X8Y9_LUT4AB/W6BEG[0] Tile_X8Y9_LUT4AB/W6BEG[10] Tile_X8Y9_LUT4AB/W6BEG[11]
+ Tile_X8Y9_LUT4AB/W6BEG[1] Tile_X8Y9_LUT4AB/W6BEG[2] Tile_X8Y9_LUT4AB/W6BEG[3] Tile_X8Y9_LUT4AB/W6BEG[4]
+ Tile_X8Y9_LUT4AB/W6BEG[5] Tile_X8Y9_LUT4AB/W6BEG[6] Tile_X8Y9_LUT4AB/W6BEG[7] Tile_X8Y9_LUT4AB/W6BEG[8]
+ Tile_X8Y9_LUT4AB/W6BEG[9] Tile_X6Y9_LUT4AB/WW4END[0] Tile_X6Y9_LUT4AB/WW4END[10]
+ Tile_X6Y9_LUT4AB/WW4END[11] Tile_X6Y9_LUT4AB/WW4END[12] Tile_X6Y9_LUT4AB/WW4END[13]
+ Tile_X6Y9_LUT4AB/WW4END[14] Tile_X6Y9_LUT4AB/WW4END[15] Tile_X6Y9_LUT4AB/WW4END[1]
+ Tile_X6Y9_LUT4AB/WW4END[2] Tile_X6Y9_LUT4AB/WW4END[3] Tile_X6Y9_LUT4AB/WW4END[4]
+ Tile_X6Y9_LUT4AB/WW4END[5] Tile_X6Y9_LUT4AB/WW4END[6] Tile_X6Y9_LUT4AB/WW4END[7]
+ Tile_X6Y9_LUT4AB/WW4END[8] Tile_X6Y9_LUT4AB/WW4END[9] Tile_X8Y9_LUT4AB/WW4BEG[0]
+ Tile_X8Y9_LUT4AB/WW4BEG[10] Tile_X8Y9_LUT4AB/WW4BEG[11] Tile_X8Y9_LUT4AB/WW4BEG[12]
+ Tile_X8Y9_LUT4AB/WW4BEG[13] Tile_X8Y9_LUT4AB/WW4BEG[14] Tile_X8Y9_LUT4AB/WW4BEG[15]
+ Tile_X8Y9_LUT4AB/WW4BEG[1] Tile_X8Y9_LUT4AB/WW4BEG[2] Tile_X8Y9_LUT4AB/WW4BEG[3]
+ Tile_X8Y9_LUT4AB/WW4BEG[4] Tile_X8Y9_LUT4AB/WW4BEG[5] Tile_X8Y9_LUT4AB/WW4BEG[6]
+ Tile_X8Y9_LUT4AB/WW4BEG[7] Tile_X8Y9_LUT4AB/WW4BEG[8] Tile_X8Y9_LUT4AB/WW4BEG[9]
+ Tile_X8Y10_LUT4AB/E1END[0] Tile_X8Y10_LUT4AB/E1END[1] Tile_X8Y10_LUT4AB/E1END[2]
+ Tile_X8Y10_LUT4AB/E1END[3] Tile_X6Y10_LUT4AB/E1BEG[0] Tile_X6Y10_LUT4AB/E1BEG[1]
+ Tile_X6Y10_LUT4AB/E1BEG[2] Tile_X6Y10_LUT4AB/E1BEG[3] Tile_X8Y10_LUT4AB/E2MID[0]
+ Tile_X8Y10_LUT4AB/E2MID[1] Tile_X8Y10_LUT4AB/E2MID[2] Tile_X8Y10_LUT4AB/E2MID[3]
+ Tile_X8Y10_LUT4AB/E2MID[4] Tile_X8Y10_LUT4AB/E2MID[5] Tile_X8Y10_LUT4AB/E2MID[6]
+ Tile_X8Y10_LUT4AB/E2MID[7] Tile_X8Y10_LUT4AB/E2END[0] Tile_X8Y10_LUT4AB/E2END[1]
+ Tile_X8Y10_LUT4AB/E2END[2] Tile_X8Y10_LUT4AB/E2END[3] Tile_X8Y10_LUT4AB/E2END[4]
+ Tile_X8Y10_LUT4AB/E2END[5] Tile_X8Y10_LUT4AB/E2END[6] Tile_X8Y10_LUT4AB/E2END[7]
+ Tile_X6Y10_LUT4AB/E2BEGb[0] Tile_X6Y10_LUT4AB/E2BEGb[1] Tile_X6Y10_LUT4AB/E2BEGb[2]
+ Tile_X6Y10_LUT4AB/E2BEGb[3] Tile_X6Y10_LUT4AB/E2BEGb[4] Tile_X6Y10_LUT4AB/E2BEGb[5]
+ Tile_X6Y10_LUT4AB/E2BEGb[6] Tile_X6Y10_LUT4AB/E2BEGb[7] Tile_X6Y10_LUT4AB/E2BEG[0]
+ Tile_X6Y10_LUT4AB/E2BEG[1] Tile_X6Y10_LUT4AB/E2BEG[2] Tile_X6Y10_LUT4AB/E2BEG[3]
+ Tile_X6Y10_LUT4AB/E2BEG[4] Tile_X6Y10_LUT4AB/E2BEG[5] Tile_X6Y10_LUT4AB/E2BEG[6]
+ Tile_X6Y10_LUT4AB/E2BEG[7] Tile_X8Y10_LUT4AB/E6END[0] Tile_X8Y10_LUT4AB/E6END[10]
+ Tile_X8Y10_LUT4AB/E6END[11] Tile_X8Y10_LUT4AB/E6END[1] Tile_X8Y10_LUT4AB/E6END[2]
+ Tile_X8Y10_LUT4AB/E6END[3] Tile_X8Y10_LUT4AB/E6END[4] Tile_X8Y10_LUT4AB/E6END[5]
+ Tile_X8Y10_LUT4AB/E6END[6] Tile_X8Y10_LUT4AB/E6END[7] Tile_X8Y10_LUT4AB/E6END[8]
+ Tile_X8Y10_LUT4AB/E6END[9] Tile_X6Y10_LUT4AB/E6BEG[0] Tile_X6Y10_LUT4AB/E6BEG[10]
+ Tile_X6Y10_LUT4AB/E6BEG[11] Tile_X6Y10_LUT4AB/E6BEG[1] Tile_X6Y10_LUT4AB/E6BEG[2]
+ Tile_X6Y10_LUT4AB/E6BEG[3] Tile_X6Y10_LUT4AB/E6BEG[4] Tile_X6Y10_LUT4AB/E6BEG[5]
+ Tile_X6Y10_LUT4AB/E6BEG[6] Tile_X6Y10_LUT4AB/E6BEG[7] Tile_X6Y10_LUT4AB/E6BEG[8]
+ Tile_X6Y10_LUT4AB/E6BEG[9] Tile_X8Y10_LUT4AB/EE4END[0] Tile_X8Y10_LUT4AB/EE4END[10]
+ Tile_X8Y10_LUT4AB/EE4END[11] Tile_X8Y10_LUT4AB/EE4END[12] Tile_X8Y10_LUT4AB/EE4END[13]
+ Tile_X8Y10_LUT4AB/EE4END[14] Tile_X8Y10_LUT4AB/EE4END[15] Tile_X8Y10_LUT4AB/EE4END[1]
+ Tile_X8Y10_LUT4AB/EE4END[2] Tile_X8Y10_LUT4AB/EE4END[3] Tile_X8Y10_LUT4AB/EE4END[4]
+ Tile_X8Y10_LUT4AB/EE4END[5] Tile_X8Y10_LUT4AB/EE4END[6] Tile_X8Y10_LUT4AB/EE4END[7]
+ Tile_X8Y10_LUT4AB/EE4END[8] Tile_X8Y10_LUT4AB/EE4END[9] Tile_X6Y10_LUT4AB/EE4BEG[0]
+ Tile_X6Y10_LUT4AB/EE4BEG[10] Tile_X6Y10_LUT4AB/EE4BEG[11] Tile_X6Y10_LUT4AB/EE4BEG[12]
+ Tile_X6Y10_LUT4AB/EE4BEG[13] Tile_X6Y10_LUT4AB/EE4BEG[14] Tile_X6Y10_LUT4AB/EE4BEG[15]
+ Tile_X6Y10_LUT4AB/EE4BEG[1] Tile_X6Y10_LUT4AB/EE4BEG[2] Tile_X6Y10_LUT4AB/EE4BEG[3]
+ Tile_X6Y10_LUT4AB/EE4BEG[4] Tile_X6Y10_LUT4AB/EE4BEG[5] Tile_X6Y10_LUT4AB/EE4BEG[6]
+ Tile_X6Y10_LUT4AB/EE4BEG[7] Tile_X6Y10_LUT4AB/EE4BEG[8] Tile_X6Y10_LUT4AB/EE4BEG[9]
+ Tile_X6Y10_LUT4AB/FrameData_O[0] Tile_X6Y10_LUT4AB/FrameData_O[10] Tile_X6Y10_LUT4AB/FrameData_O[11]
+ Tile_X6Y10_LUT4AB/FrameData_O[12] Tile_X6Y10_LUT4AB/FrameData_O[13] Tile_X6Y10_LUT4AB/FrameData_O[14]
+ Tile_X6Y10_LUT4AB/FrameData_O[15] Tile_X6Y10_LUT4AB/FrameData_O[16] Tile_X6Y10_LUT4AB/FrameData_O[17]
+ Tile_X6Y10_LUT4AB/FrameData_O[18] Tile_X6Y10_LUT4AB/FrameData_O[19] Tile_X6Y10_LUT4AB/FrameData_O[1]
+ Tile_X6Y10_LUT4AB/FrameData_O[20] Tile_X6Y10_LUT4AB/FrameData_O[21] Tile_X6Y10_LUT4AB/FrameData_O[22]
+ Tile_X6Y10_LUT4AB/FrameData_O[23] Tile_X6Y10_LUT4AB/FrameData_O[24] Tile_X6Y10_LUT4AB/FrameData_O[25]
+ Tile_X6Y10_LUT4AB/FrameData_O[26] Tile_X6Y10_LUT4AB/FrameData_O[27] Tile_X6Y10_LUT4AB/FrameData_O[28]
+ Tile_X6Y10_LUT4AB/FrameData_O[29] Tile_X6Y10_LUT4AB/FrameData_O[2] Tile_X6Y10_LUT4AB/FrameData_O[30]
+ Tile_X6Y10_LUT4AB/FrameData_O[31] Tile_X6Y10_LUT4AB/FrameData_O[3] Tile_X6Y10_LUT4AB/FrameData_O[4]
+ Tile_X6Y10_LUT4AB/FrameData_O[5] Tile_X6Y10_LUT4AB/FrameData_O[6] Tile_X6Y10_LUT4AB/FrameData_O[7]
+ Tile_X6Y10_LUT4AB/FrameData_O[8] Tile_X6Y10_LUT4AB/FrameData_O[9] Tile_X8Y10_LUT4AB/FrameData[0]
+ Tile_X8Y10_LUT4AB/FrameData[10] Tile_X8Y10_LUT4AB/FrameData[11] Tile_X8Y10_LUT4AB/FrameData[12]
+ Tile_X8Y10_LUT4AB/FrameData[13] Tile_X8Y10_LUT4AB/FrameData[14] Tile_X8Y10_LUT4AB/FrameData[15]
+ Tile_X8Y10_LUT4AB/FrameData[16] Tile_X8Y10_LUT4AB/FrameData[17] Tile_X8Y10_LUT4AB/FrameData[18]
+ Tile_X8Y10_LUT4AB/FrameData[19] Tile_X8Y10_LUT4AB/FrameData[1] Tile_X8Y10_LUT4AB/FrameData[20]
+ Tile_X8Y10_LUT4AB/FrameData[21] Tile_X8Y10_LUT4AB/FrameData[22] Tile_X8Y10_LUT4AB/FrameData[23]
+ Tile_X8Y10_LUT4AB/FrameData[24] Tile_X8Y10_LUT4AB/FrameData[25] Tile_X8Y10_LUT4AB/FrameData[26]
+ Tile_X8Y10_LUT4AB/FrameData[27] Tile_X8Y10_LUT4AB/FrameData[28] Tile_X8Y10_LUT4AB/FrameData[29]
+ Tile_X8Y10_LUT4AB/FrameData[2] Tile_X8Y10_LUT4AB/FrameData[30] Tile_X8Y10_LUT4AB/FrameData[31]
+ Tile_X8Y10_LUT4AB/FrameData[3] Tile_X8Y10_LUT4AB/FrameData[4] Tile_X8Y10_LUT4AB/FrameData[5]
+ Tile_X8Y10_LUT4AB/FrameData[6] Tile_X8Y10_LUT4AB/FrameData[7] Tile_X8Y10_LUT4AB/FrameData[8]
+ Tile_X8Y10_LUT4AB/FrameData[9] Tile_X7Y9_DSP/Tile_X0Y1_FrameStrobe[0] Tile_X7Y9_DSP/Tile_X0Y1_FrameStrobe[10]
+ Tile_X7Y9_DSP/Tile_X0Y1_FrameStrobe[11] Tile_X7Y9_DSP/Tile_X0Y1_FrameStrobe[12]
+ Tile_X7Y9_DSP/Tile_X0Y1_FrameStrobe[13] Tile_X7Y9_DSP/Tile_X0Y1_FrameStrobe[14]
+ Tile_X7Y9_DSP/Tile_X0Y1_FrameStrobe[15] Tile_X7Y9_DSP/Tile_X0Y1_FrameStrobe[16]
+ Tile_X7Y9_DSP/Tile_X0Y1_FrameStrobe[17] Tile_X7Y9_DSP/Tile_X0Y1_FrameStrobe[18]
+ Tile_X7Y9_DSP/Tile_X0Y1_FrameStrobe[19] Tile_X7Y9_DSP/Tile_X0Y1_FrameStrobe[1] Tile_X7Y9_DSP/Tile_X0Y1_FrameStrobe[2]
+ Tile_X7Y9_DSP/Tile_X0Y1_FrameStrobe[3] Tile_X7Y9_DSP/Tile_X0Y1_FrameStrobe[4] Tile_X7Y9_DSP/Tile_X0Y1_FrameStrobe[5]
+ Tile_X7Y9_DSP/Tile_X0Y1_FrameStrobe[6] Tile_X7Y9_DSP/Tile_X0Y1_FrameStrobe[7] Tile_X7Y9_DSP/Tile_X0Y1_FrameStrobe[8]
+ Tile_X7Y9_DSP/Tile_X0Y1_FrameStrobe[9] Tile_X7Y9_DSP/Tile_X0Y1_N1END[0] Tile_X7Y9_DSP/Tile_X0Y1_N1END[1]
+ Tile_X7Y9_DSP/Tile_X0Y1_N1END[2] Tile_X7Y9_DSP/Tile_X0Y1_N1END[3] Tile_X7Y9_DSP/Tile_X0Y1_N2END[0]
+ Tile_X7Y9_DSP/Tile_X0Y1_N2END[1] Tile_X7Y9_DSP/Tile_X0Y1_N2END[2] Tile_X7Y9_DSP/Tile_X0Y1_N2END[3]
+ Tile_X7Y9_DSP/Tile_X0Y1_N2END[4] Tile_X7Y9_DSP/Tile_X0Y1_N2END[5] Tile_X7Y9_DSP/Tile_X0Y1_N2END[6]
+ Tile_X7Y9_DSP/Tile_X0Y1_N2END[7] Tile_X7Y9_DSP/Tile_X0Y1_N2MID[0] Tile_X7Y9_DSP/Tile_X0Y1_N2MID[1]
+ Tile_X7Y9_DSP/Tile_X0Y1_N2MID[2] Tile_X7Y9_DSP/Tile_X0Y1_N2MID[3] Tile_X7Y9_DSP/Tile_X0Y1_N2MID[4]
+ Tile_X7Y9_DSP/Tile_X0Y1_N2MID[5] Tile_X7Y9_DSP/Tile_X0Y1_N2MID[6] Tile_X7Y9_DSP/Tile_X0Y1_N2MID[7]
+ Tile_X7Y9_DSP/Tile_X0Y1_N4END[0] Tile_X7Y9_DSP/Tile_X0Y1_N4END[10] Tile_X7Y9_DSP/Tile_X0Y1_N4END[11]
+ Tile_X7Y9_DSP/Tile_X0Y1_N4END[12] Tile_X7Y9_DSP/Tile_X0Y1_N4END[13] Tile_X7Y9_DSP/Tile_X0Y1_N4END[14]
+ Tile_X7Y9_DSP/Tile_X0Y1_N4END[15] Tile_X7Y9_DSP/Tile_X0Y1_N4END[1] Tile_X7Y9_DSP/Tile_X0Y1_N4END[2]
+ Tile_X7Y9_DSP/Tile_X0Y1_N4END[3] Tile_X7Y9_DSP/Tile_X0Y1_N4END[4] Tile_X7Y9_DSP/Tile_X0Y1_N4END[5]
+ Tile_X7Y9_DSP/Tile_X0Y1_N4END[6] Tile_X7Y9_DSP/Tile_X0Y1_N4END[7] Tile_X7Y9_DSP/Tile_X0Y1_N4END[8]
+ Tile_X7Y9_DSP/Tile_X0Y1_N4END[9] Tile_X7Y9_DSP/Tile_X0Y1_NN4END[0] Tile_X7Y9_DSP/Tile_X0Y1_NN4END[10]
+ Tile_X7Y9_DSP/Tile_X0Y1_NN4END[11] Tile_X7Y9_DSP/Tile_X0Y1_NN4END[12] Tile_X7Y9_DSP/Tile_X0Y1_NN4END[13]
+ Tile_X7Y9_DSP/Tile_X0Y1_NN4END[14] Tile_X7Y9_DSP/Tile_X0Y1_NN4END[15] Tile_X7Y9_DSP/Tile_X0Y1_NN4END[1]
+ Tile_X7Y9_DSP/Tile_X0Y1_NN4END[2] Tile_X7Y9_DSP/Tile_X0Y1_NN4END[3] Tile_X7Y9_DSP/Tile_X0Y1_NN4END[4]
+ Tile_X7Y9_DSP/Tile_X0Y1_NN4END[5] Tile_X7Y9_DSP/Tile_X0Y1_NN4END[6] Tile_X7Y9_DSP/Tile_X0Y1_NN4END[7]
+ Tile_X7Y9_DSP/Tile_X0Y1_NN4END[8] Tile_X7Y9_DSP/Tile_X0Y1_NN4END[9] Tile_X7Y9_DSP/Tile_X0Y1_S1BEG[0]
+ Tile_X7Y9_DSP/Tile_X0Y1_S1BEG[1] Tile_X7Y9_DSP/Tile_X0Y1_S1BEG[2] Tile_X7Y9_DSP/Tile_X0Y1_S1BEG[3]
+ Tile_X7Y9_DSP/Tile_X0Y1_S2BEG[0] Tile_X7Y9_DSP/Tile_X0Y1_S2BEG[1] Tile_X7Y9_DSP/Tile_X0Y1_S2BEG[2]
+ Tile_X7Y9_DSP/Tile_X0Y1_S2BEG[3] Tile_X7Y9_DSP/Tile_X0Y1_S2BEG[4] Tile_X7Y9_DSP/Tile_X0Y1_S2BEG[5]
+ Tile_X7Y9_DSP/Tile_X0Y1_S2BEG[6] Tile_X7Y9_DSP/Tile_X0Y1_S2BEG[7] Tile_X7Y9_DSP/Tile_X0Y1_S2BEGb[0]
+ Tile_X7Y9_DSP/Tile_X0Y1_S2BEGb[1] Tile_X7Y9_DSP/Tile_X0Y1_S2BEGb[2] Tile_X7Y9_DSP/Tile_X0Y1_S2BEGb[3]
+ Tile_X7Y9_DSP/Tile_X0Y1_S2BEGb[4] Tile_X7Y9_DSP/Tile_X0Y1_S2BEGb[5] Tile_X7Y9_DSP/Tile_X0Y1_S2BEGb[6]
+ Tile_X7Y9_DSP/Tile_X0Y1_S2BEGb[7] Tile_X7Y9_DSP/Tile_X0Y1_S4BEG[0] Tile_X7Y9_DSP/Tile_X0Y1_S4BEG[10]
+ Tile_X7Y9_DSP/Tile_X0Y1_S4BEG[11] Tile_X7Y9_DSP/Tile_X0Y1_S4BEG[12] Tile_X7Y9_DSP/Tile_X0Y1_S4BEG[13]
+ Tile_X7Y9_DSP/Tile_X0Y1_S4BEG[14] Tile_X7Y9_DSP/Tile_X0Y1_S4BEG[15] Tile_X7Y9_DSP/Tile_X0Y1_S4BEG[1]
+ Tile_X7Y9_DSP/Tile_X0Y1_S4BEG[2] Tile_X7Y9_DSP/Tile_X0Y1_S4BEG[3] Tile_X7Y9_DSP/Tile_X0Y1_S4BEG[4]
+ Tile_X7Y9_DSP/Tile_X0Y1_S4BEG[5] Tile_X7Y9_DSP/Tile_X0Y1_S4BEG[6] Tile_X7Y9_DSP/Tile_X0Y1_S4BEG[7]
+ Tile_X7Y9_DSP/Tile_X0Y1_S4BEG[8] Tile_X7Y9_DSP/Tile_X0Y1_S4BEG[9] Tile_X7Y9_DSP/Tile_X0Y1_SS4BEG[0]
+ Tile_X7Y9_DSP/Tile_X0Y1_SS4BEG[10] Tile_X7Y9_DSP/Tile_X0Y1_SS4BEG[11] Tile_X7Y9_DSP/Tile_X0Y1_SS4BEG[12]
+ Tile_X7Y9_DSP/Tile_X0Y1_SS4BEG[13] Tile_X7Y9_DSP/Tile_X0Y1_SS4BEG[14] Tile_X7Y9_DSP/Tile_X0Y1_SS4BEG[15]
+ Tile_X7Y9_DSP/Tile_X0Y1_SS4BEG[1] Tile_X7Y9_DSP/Tile_X0Y1_SS4BEG[2] Tile_X7Y9_DSP/Tile_X0Y1_SS4BEG[3]
+ Tile_X7Y9_DSP/Tile_X0Y1_SS4BEG[4] Tile_X7Y9_DSP/Tile_X0Y1_SS4BEG[5] Tile_X7Y9_DSP/Tile_X0Y1_SS4BEG[6]
+ Tile_X7Y9_DSP/Tile_X0Y1_SS4BEG[7] Tile_X7Y9_DSP/Tile_X0Y1_SS4BEG[8] Tile_X7Y9_DSP/Tile_X0Y1_SS4BEG[9]
+ Tile_X7Y9_DSP/Tile_X0Y1_UserCLK Tile_X6Y10_LUT4AB/W1END[0] Tile_X6Y10_LUT4AB/W1END[1]
+ Tile_X6Y10_LUT4AB/W1END[2] Tile_X6Y10_LUT4AB/W1END[3] Tile_X8Y10_LUT4AB/W1BEG[0]
+ Tile_X8Y10_LUT4AB/W1BEG[1] Tile_X8Y10_LUT4AB/W1BEG[2] Tile_X8Y10_LUT4AB/W1BEG[3]
+ Tile_X6Y10_LUT4AB/W2MID[0] Tile_X6Y10_LUT4AB/W2MID[1] Tile_X6Y10_LUT4AB/W2MID[2]
+ Tile_X6Y10_LUT4AB/W2MID[3] Tile_X6Y10_LUT4AB/W2MID[4] Tile_X6Y10_LUT4AB/W2MID[5]
+ Tile_X6Y10_LUT4AB/W2MID[6] Tile_X6Y10_LUT4AB/W2MID[7] Tile_X6Y10_LUT4AB/W2END[0]
+ Tile_X6Y10_LUT4AB/W2END[1] Tile_X6Y10_LUT4AB/W2END[2] Tile_X6Y10_LUT4AB/W2END[3]
+ Tile_X6Y10_LUT4AB/W2END[4] Tile_X6Y10_LUT4AB/W2END[5] Tile_X6Y10_LUT4AB/W2END[6]
+ Tile_X6Y10_LUT4AB/W2END[7] Tile_X8Y10_LUT4AB/W2BEGb[0] Tile_X8Y10_LUT4AB/W2BEGb[1]
+ Tile_X8Y10_LUT4AB/W2BEGb[2] Tile_X8Y10_LUT4AB/W2BEGb[3] Tile_X8Y10_LUT4AB/W2BEGb[4]
+ Tile_X8Y10_LUT4AB/W2BEGb[5] Tile_X8Y10_LUT4AB/W2BEGb[6] Tile_X8Y10_LUT4AB/W2BEGb[7]
+ Tile_X8Y10_LUT4AB/W2BEG[0] Tile_X8Y10_LUT4AB/W2BEG[1] Tile_X8Y10_LUT4AB/W2BEG[2]
+ Tile_X8Y10_LUT4AB/W2BEG[3] Tile_X8Y10_LUT4AB/W2BEG[4] Tile_X8Y10_LUT4AB/W2BEG[5]
+ Tile_X8Y10_LUT4AB/W2BEG[6] Tile_X8Y10_LUT4AB/W2BEG[7] Tile_X6Y10_LUT4AB/W6END[0]
+ Tile_X6Y10_LUT4AB/W6END[10] Tile_X6Y10_LUT4AB/W6END[11] Tile_X6Y10_LUT4AB/W6END[1]
+ Tile_X6Y10_LUT4AB/W6END[2] Tile_X6Y10_LUT4AB/W6END[3] Tile_X6Y10_LUT4AB/W6END[4]
+ Tile_X6Y10_LUT4AB/W6END[5] Tile_X6Y10_LUT4AB/W6END[6] Tile_X6Y10_LUT4AB/W6END[7]
+ Tile_X6Y10_LUT4AB/W6END[8] Tile_X6Y10_LUT4AB/W6END[9] Tile_X8Y10_LUT4AB/W6BEG[0]
+ Tile_X8Y10_LUT4AB/W6BEG[10] Tile_X8Y10_LUT4AB/W6BEG[11] Tile_X8Y10_LUT4AB/W6BEG[1]
+ Tile_X8Y10_LUT4AB/W6BEG[2] Tile_X8Y10_LUT4AB/W6BEG[3] Tile_X8Y10_LUT4AB/W6BEG[4]
+ Tile_X8Y10_LUT4AB/W6BEG[5] Tile_X8Y10_LUT4AB/W6BEG[6] Tile_X8Y10_LUT4AB/W6BEG[7]
+ Tile_X8Y10_LUT4AB/W6BEG[8] Tile_X8Y10_LUT4AB/W6BEG[9] Tile_X6Y10_LUT4AB/WW4END[0]
+ Tile_X6Y10_LUT4AB/WW4END[10] Tile_X6Y10_LUT4AB/WW4END[11] Tile_X6Y10_LUT4AB/WW4END[12]
+ Tile_X6Y10_LUT4AB/WW4END[13] Tile_X6Y10_LUT4AB/WW4END[14] Tile_X6Y10_LUT4AB/WW4END[15]
+ Tile_X6Y10_LUT4AB/WW4END[1] Tile_X6Y10_LUT4AB/WW4END[2] Tile_X6Y10_LUT4AB/WW4END[3]
+ Tile_X6Y10_LUT4AB/WW4END[4] Tile_X6Y10_LUT4AB/WW4END[5] Tile_X6Y10_LUT4AB/WW4END[6]
+ Tile_X6Y10_LUT4AB/WW4END[7] Tile_X6Y10_LUT4AB/WW4END[8] Tile_X6Y10_LUT4AB/WW4END[9]
+ Tile_X8Y10_LUT4AB/WW4BEG[0] Tile_X8Y10_LUT4AB/WW4BEG[10] Tile_X8Y10_LUT4AB/WW4BEG[11]
+ Tile_X8Y10_LUT4AB/WW4BEG[12] Tile_X8Y10_LUT4AB/WW4BEG[13] Tile_X8Y10_LUT4AB/WW4BEG[14]
+ Tile_X8Y10_LUT4AB/WW4BEG[15] Tile_X8Y10_LUT4AB/WW4BEG[1] Tile_X8Y10_LUT4AB/WW4BEG[2]
+ Tile_X8Y10_LUT4AB/WW4BEG[3] Tile_X8Y10_LUT4AB/WW4BEG[4] Tile_X8Y10_LUT4AB/WW4BEG[5]
+ Tile_X8Y10_LUT4AB/WW4BEG[6] Tile_X8Y10_LUT4AB/WW4BEG[7] Tile_X8Y10_LUT4AB/WW4BEG[8]
+ Tile_X8Y10_LUT4AB/WW4BEG[9] VGND VPWR DSP
XTile_X8Y10_LUT4AB Tile_X8Y11_LUT4AB/Co Tile_X8Y9_LUT4AB/Ci Tile_X9Y10_LUT4AB/E1END[0]
+ Tile_X9Y10_LUT4AB/E1END[1] Tile_X9Y10_LUT4AB/E1END[2] Tile_X9Y10_LUT4AB/E1END[3]
+ Tile_X8Y10_LUT4AB/E1END[0] Tile_X8Y10_LUT4AB/E1END[1] Tile_X8Y10_LUT4AB/E1END[2]
+ Tile_X8Y10_LUT4AB/E1END[3] Tile_X9Y10_LUT4AB/E2MID[0] Tile_X9Y10_LUT4AB/E2MID[1]
+ Tile_X9Y10_LUT4AB/E2MID[2] Tile_X9Y10_LUT4AB/E2MID[3] Tile_X9Y10_LUT4AB/E2MID[4]
+ Tile_X9Y10_LUT4AB/E2MID[5] Tile_X9Y10_LUT4AB/E2MID[6] Tile_X9Y10_LUT4AB/E2MID[7]
+ Tile_X9Y10_LUT4AB/E2END[0] Tile_X9Y10_LUT4AB/E2END[1] Tile_X9Y10_LUT4AB/E2END[2]
+ Tile_X9Y10_LUT4AB/E2END[3] Tile_X9Y10_LUT4AB/E2END[4] Tile_X9Y10_LUT4AB/E2END[5]
+ Tile_X9Y10_LUT4AB/E2END[6] Tile_X9Y10_LUT4AB/E2END[7] Tile_X8Y10_LUT4AB/E2END[0]
+ Tile_X8Y10_LUT4AB/E2END[1] Tile_X8Y10_LUT4AB/E2END[2] Tile_X8Y10_LUT4AB/E2END[3]
+ Tile_X8Y10_LUT4AB/E2END[4] Tile_X8Y10_LUT4AB/E2END[5] Tile_X8Y10_LUT4AB/E2END[6]
+ Tile_X8Y10_LUT4AB/E2END[7] Tile_X8Y10_LUT4AB/E2MID[0] Tile_X8Y10_LUT4AB/E2MID[1]
+ Tile_X8Y10_LUT4AB/E2MID[2] Tile_X8Y10_LUT4AB/E2MID[3] Tile_X8Y10_LUT4AB/E2MID[4]
+ Tile_X8Y10_LUT4AB/E2MID[5] Tile_X8Y10_LUT4AB/E2MID[6] Tile_X8Y10_LUT4AB/E2MID[7]
+ Tile_X9Y10_LUT4AB/E6END[0] Tile_X9Y10_LUT4AB/E6END[10] Tile_X9Y10_LUT4AB/E6END[11]
+ Tile_X9Y10_LUT4AB/E6END[1] Tile_X9Y10_LUT4AB/E6END[2] Tile_X9Y10_LUT4AB/E6END[3]
+ Tile_X9Y10_LUT4AB/E6END[4] Tile_X9Y10_LUT4AB/E6END[5] Tile_X9Y10_LUT4AB/E6END[6]
+ Tile_X9Y10_LUT4AB/E6END[7] Tile_X9Y10_LUT4AB/E6END[8] Tile_X9Y10_LUT4AB/E6END[9]
+ Tile_X8Y10_LUT4AB/E6END[0] Tile_X8Y10_LUT4AB/E6END[10] Tile_X8Y10_LUT4AB/E6END[11]
+ Tile_X8Y10_LUT4AB/E6END[1] Tile_X8Y10_LUT4AB/E6END[2] Tile_X8Y10_LUT4AB/E6END[3]
+ Tile_X8Y10_LUT4AB/E6END[4] Tile_X8Y10_LUT4AB/E6END[5] Tile_X8Y10_LUT4AB/E6END[6]
+ Tile_X8Y10_LUT4AB/E6END[7] Tile_X8Y10_LUT4AB/E6END[8] Tile_X8Y10_LUT4AB/E6END[9]
+ Tile_X9Y10_LUT4AB/EE4END[0] Tile_X9Y10_LUT4AB/EE4END[10] Tile_X9Y10_LUT4AB/EE4END[11]
+ Tile_X9Y10_LUT4AB/EE4END[12] Tile_X9Y10_LUT4AB/EE4END[13] Tile_X9Y10_LUT4AB/EE4END[14]
+ Tile_X9Y10_LUT4AB/EE4END[15] Tile_X9Y10_LUT4AB/EE4END[1] Tile_X9Y10_LUT4AB/EE4END[2]
+ Tile_X9Y10_LUT4AB/EE4END[3] Tile_X9Y10_LUT4AB/EE4END[4] Tile_X9Y10_LUT4AB/EE4END[5]
+ Tile_X9Y10_LUT4AB/EE4END[6] Tile_X9Y10_LUT4AB/EE4END[7] Tile_X9Y10_LUT4AB/EE4END[8]
+ Tile_X9Y10_LUT4AB/EE4END[9] Tile_X8Y10_LUT4AB/EE4END[0] Tile_X8Y10_LUT4AB/EE4END[10]
+ Tile_X8Y10_LUT4AB/EE4END[11] Tile_X8Y10_LUT4AB/EE4END[12] Tile_X8Y10_LUT4AB/EE4END[13]
+ Tile_X8Y10_LUT4AB/EE4END[14] Tile_X8Y10_LUT4AB/EE4END[15] Tile_X8Y10_LUT4AB/EE4END[1]
+ Tile_X8Y10_LUT4AB/EE4END[2] Tile_X8Y10_LUT4AB/EE4END[3] Tile_X8Y10_LUT4AB/EE4END[4]
+ Tile_X8Y10_LUT4AB/EE4END[5] Tile_X8Y10_LUT4AB/EE4END[6] Tile_X8Y10_LUT4AB/EE4END[7]
+ Tile_X8Y10_LUT4AB/EE4END[8] Tile_X8Y10_LUT4AB/EE4END[9] Tile_X8Y10_LUT4AB/FrameData[0]
+ Tile_X8Y10_LUT4AB/FrameData[10] Tile_X8Y10_LUT4AB/FrameData[11] Tile_X8Y10_LUT4AB/FrameData[12]
+ Tile_X8Y10_LUT4AB/FrameData[13] Tile_X8Y10_LUT4AB/FrameData[14] Tile_X8Y10_LUT4AB/FrameData[15]
+ Tile_X8Y10_LUT4AB/FrameData[16] Tile_X8Y10_LUT4AB/FrameData[17] Tile_X8Y10_LUT4AB/FrameData[18]
+ Tile_X8Y10_LUT4AB/FrameData[19] Tile_X8Y10_LUT4AB/FrameData[1] Tile_X8Y10_LUT4AB/FrameData[20]
+ Tile_X8Y10_LUT4AB/FrameData[21] Tile_X8Y10_LUT4AB/FrameData[22] Tile_X8Y10_LUT4AB/FrameData[23]
+ Tile_X8Y10_LUT4AB/FrameData[24] Tile_X8Y10_LUT4AB/FrameData[25] Tile_X8Y10_LUT4AB/FrameData[26]
+ Tile_X8Y10_LUT4AB/FrameData[27] Tile_X8Y10_LUT4AB/FrameData[28] Tile_X8Y10_LUT4AB/FrameData[29]
+ Tile_X8Y10_LUT4AB/FrameData[2] Tile_X8Y10_LUT4AB/FrameData[30] Tile_X8Y10_LUT4AB/FrameData[31]
+ Tile_X8Y10_LUT4AB/FrameData[3] Tile_X8Y10_LUT4AB/FrameData[4] Tile_X8Y10_LUT4AB/FrameData[5]
+ Tile_X8Y10_LUT4AB/FrameData[6] Tile_X8Y10_LUT4AB/FrameData[7] Tile_X8Y10_LUT4AB/FrameData[8]
+ Tile_X8Y10_LUT4AB/FrameData[9] Tile_X9Y10_LUT4AB/FrameData[0] Tile_X9Y10_LUT4AB/FrameData[10]
+ Tile_X9Y10_LUT4AB/FrameData[11] Tile_X9Y10_LUT4AB/FrameData[12] Tile_X9Y10_LUT4AB/FrameData[13]
+ Tile_X9Y10_LUT4AB/FrameData[14] Tile_X9Y10_LUT4AB/FrameData[15] Tile_X9Y10_LUT4AB/FrameData[16]
+ Tile_X9Y10_LUT4AB/FrameData[17] Tile_X9Y10_LUT4AB/FrameData[18] Tile_X9Y10_LUT4AB/FrameData[19]
+ Tile_X9Y10_LUT4AB/FrameData[1] Tile_X9Y10_LUT4AB/FrameData[20] Tile_X9Y10_LUT4AB/FrameData[21]
+ Tile_X9Y10_LUT4AB/FrameData[22] Tile_X9Y10_LUT4AB/FrameData[23] Tile_X9Y10_LUT4AB/FrameData[24]
+ Tile_X9Y10_LUT4AB/FrameData[25] Tile_X9Y10_LUT4AB/FrameData[26] Tile_X9Y10_LUT4AB/FrameData[27]
+ Tile_X9Y10_LUT4AB/FrameData[28] Tile_X9Y10_LUT4AB/FrameData[29] Tile_X9Y10_LUT4AB/FrameData[2]
+ Tile_X9Y10_LUT4AB/FrameData[30] Tile_X9Y10_LUT4AB/FrameData[31] Tile_X9Y10_LUT4AB/FrameData[3]
+ Tile_X9Y10_LUT4AB/FrameData[4] Tile_X9Y10_LUT4AB/FrameData[5] Tile_X9Y10_LUT4AB/FrameData[6]
+ Tile_X9Y10_LUT4AB/FrameData[7] Tile_X9Y10_LUT4AB/FrameData[8] Tile_X9Y10_LUT4AB/FrameData[9]
+ Tile_X8Y10_LUT4AB/FrameStrobe[0] Tile_X8Y10_LUT4AB/FrameStrobe[10] Tile_X8Y10_LUT4AB/FrameStrobe[11]
+ Tile_X8Y10_LUT4AB/FrameStrobe[12] Tile_X8Y10_LUT4AB/FrameStrobe[13] Tile_X8Y10_LUT4AB/FrameStrobe[14]
+ Tile_X8Y10_LUT4AB/FrameStrobe[15] Tile_X8Y10_LUT4AB/FrameStrobe[16] Tile_X8Y10_LUT4AB/FrameStrobe[17]
+ Tile_X8Y10_LUT4AB/FrameStrobe[18] Tile_X8Y10_LUT4AB/FrameStrobe[19] Tile_X8Y10_LUT4AB/FrameStrobe[1]
+ Tile_X8Y10_LUT4AB/FrameStrobe[2] Tile_X8Y10_LUT4AB/FrameStrobe[3] Tile_X8Y10_LUT4AB/FrameStrobe[4]
+ Tile_X8Y10_LUT4AB/FrameStrobe[5] Tile_X8Y10_LUT4AB/FrameStrobe[6] Tile_X8Y10_LUT4AB/FrameStrobe[7]
+ Tile_X8Y10_LUT4AB/FrameStrobe[8] Tile_X8Y10_LUT4AB/FrameStrobe[9] Tile_X8Y9_LUT4AB/FrameStrobe[0]
+ Tile_X8Y9_LUT4AB/FrameStrobe[10] Tile_X8Y9_LUT4AB/FrameStrobe[11] Tile_X8Y9_LUT4AB/FrameStrobe[12]
+ Tile_X8Y9_LUT4AB/FrameStrobe[13] Tile_X8Y9_LUT4AB/FrameStrobe[14] Tile_X8Y9_LUT4AB/FrameStrobe[15]
+ Tile_X8Y9_LUT4AB/FrameStrobe[16] Tile_X8Y9_LUT4AB/FrameStrobe[17] Tile_X8Y9_LUT4AB/FrameStrobe[18]
+ Tile_X8Y9_LUT4AB/FrameStrobe[19] Tile_X8Y9_LUT4AB/FrameStrobe[1] Tile_X8Y9_LUT4AB/FrameStrobe[2]
+ Tile_X8Y9_LUT4AB/FrameStrobe[3] Tile_X8Y9_LUT4AB/FrameStrobe[4] Tile_X8Y9_LUT4AB/FrameStrobe[5]
+ Tile_X8Y9_LUT4AB/FrameStrobe[6] Tile_X8Y9_LUT4AB/FrameStrobe[7] Tile_X8Y9_LUT4AB/FrameStrobe[8]
+ Tile_X8Y9_LUT4AB/FrameStrobe[9] Tile_X8Y9_LUT4AB/N1END[0] Tile_X8Y9_LUT4AB/N1END[1]
+ Tile_X8Y9_LUT4AB/N1END[2] Tile_X8Y9_LUT4AB/N1END[3] Tile_X8Y11_LUT4AB/N1BEG[0] Tile_X8Y11_LUT4AB/N1BEG[1]
+ Tile_X8Y11_LUT4AB/N1BEG[2] Tile_X8Y11_LUT4AB/N1BEG[3] Tile_X8Y9_LUT4AB/N2MID[0]
+ Tile_X8Y9_LUT4AB/N2MID[1] Tile_X8Y9_LUT4AB/N2MID[2] Tile_X8Y9_LUT4AB/N2MID[3] Tile_X8Y9_LUT4AB/N2MID[4]
+ Tile_X8Y9_LUT4AB/N2MID[5] Tile_X8Y9_LUT4AB/N2MID[6] Tile_X8Y9_LUT4AB/N2MID[7] Tile_X8Y9_LUT4AB/N2END[0]
+ Tile_X8Y9_LUT4AB/N2END[1] Tile_X8Y9_LUT4AB/N2END[2] Tile_X8Y9_LUT4AB/N2END[3] Tile_X8Y9_LUT4AB/N2END[4]
+ Tile_X8Y9_LUT4AB/N2END[5] Tile_X8Y9_LUT4AB/N2END[6] Tile_X8Y9_LUT4AB/N2END[7] Tile_X8Y10_LUT4AB/N2END[0]
+ Tile_X8Y10_LUT4AB/N2END[1] Tile_X8Y10_LUT4AB/N2END[2] Tile_X8Y10_LUT4AB/N2END[3]
+ Tile_X8Y10_LUT4AB/N2END[4] Tile_X8Y10_LUT4AB/N2END[5] Tile_X8Y10_LUT4AB/N2END[6]
+ Tile_X8Y10_LUT4AB/N2END[7] Tile_X8Y11_LUT4AB/N2BEG[0] Tile_X8Y11_LUT4AB/N2BEG[1]
+ Tile_X8Y11_LUT4AB/N2BEG[2] Tile_X8Y11_LUT4AB/N2BEG[3] Tile_X8Y11_LUT4AB/N2BEG[4]
+ Tile_X8Y11_LUT4AB/N2BEG[5] Tile_X8Y11_LUT4AB/N2BEG[6] Tile_X8Y11_LUT4AB/N2BEG[7]
+ Tile_X8Y9_LUT4AB/N4END[0] Tile_X8Y9_LUT4AB/N4END[10] Tile_X8Y9_LUT4AB/N4END[11]
+ Tile_X8Y9_LUT4AB/N4END[12] Tile_X8Y9_LUT4AB/N4END[13] Tile_X8Y9_LUT4AB/N4END[14]
+ Tile_X8Y9_LUT4AB/N4END[15] Tile_X8Y9_LUT4AB/N4END[1] Tile_X8Y9_LUT4AB/N4END[2] Tile_X8Y9_LUT4AB/N4END[3]
+ Tile_X8Y9_LUT4AB/N4END[4] Tile_X8Y9_LUT4AB/N4END[5] Tile_X8Y9_LUT4AB/N4END[6] Tile_X8Y9_LUT4AB/N4END[7]
+ Tile_X8Y9_LUT4AB/N4END[8] Tile_X8Y9_LUT4AB/N4END[9] Tile_X8Y11_LUT4AB/N4BEG[0] Tile_X8Y11_LUT4AB/N4BEG[10]
+ Tile_X8Y11_LUT4AB/N4BEG[11] Tile_X8Y11_LUT4AB/N4BEG[12] Tile_X8Y11_LUT4AB/N4BEG[13]
+ Tile_X8Y11_LUT4AB/N4BEG[14] Tile_X8Y11_LUT4AB/N4BEG[15] Tile_X8Y11_LUT4AB/N4BEG[1]
+ Tile_X8Y11_LUT4AB/N4BEG[2] Tile_X8Y11_LUT4AB/N4BEG[3] Tile_X8Y11_LUT4AB/N4BEG[4]
+ Tile_X8Y11_LUT4AB/N4BEG[5] Tile_X8Y11_LUT4AB/N4BEG[6] Tile_X8Y11_LUT4AB/N4BEG[7]
+ Tile_X8Y11_LUT4AB/N4BEG[8] Tile_X8Y11_LUT4AB/N4BEG[9] Tile_X8Y9_LUT4AB/NN4END[0]
+ Tile_X8Y9_LUT4AB/NN4END[10] Tile_X8Y9_LUT4AB/NN4END[11] Tile_X8Y9_LUT4AB/NN4END[12]
+ Tile_X8Y9_LUT4AB/NN4END[13] Tile_X8Y9_LUT4AB/NN4END[14] Tile_X8Y9_LUT4AB/NN4END[15]
+ Tile_X8Y9_LUT4AB/NN4END[1] Tile_X8Y9_LUT4AB/NN4END[2] Tile_X8Y9_LUT4AB/NN4END[3]
+ Tile_X8Y9_LUT4AB/NN4END[4] Tile_X8Y9_LUT4AB/NN4END[5] Tile_X8Y9_LUT4AB/NN4END[6]
+ Tile_X8Y9_LUT4AB/NN4END[7] Tile_X8Y9_LUT4AB/NN4END[8] Tile_X8Y9_LUT4AB/NN4END[9]
+ Tile_X8Y11_LUT4AB/NN4BEG[0] Tile_X8Y11_LUT4AB/NN4BEG[10] Tile_X8Y11_LUT4AB/NN4BEG[11]
+ Tile_X8Y11_LUT4AB/NN4BEG[12] Tile_X8Y11_LUT4AB/NN4BEG[13] Tile_X8Y11_LUT4AB/NN4BEG[14]
+ Tile_X8Y11_LUT4AB/NN4BEG[15] Tile_X8Y11_LUT4AB/NN4BEG[1] Tile_X8Y11_LUT4AB/NN4BEG[2]
+ Tile_X8Y11_LUT4AB/NN4BEG[3] Tile_X8Y11_LUT4AB/NN4BEG[4] Tile_X8Y11_LUT4AB/NN4BEG[5]
+ Tile_X8Y11_LUT4AB/NN4BEG[6] Tile_X8Y11_LUT4AB/NN4BEG[7] Tile_X8Y11_LUT4AB/NN4BEG[8]
+ Tile_X8Y11_LUT4AB/NN4BEG[9] Tile_X8Y11_LUT4AB/S1END[0] Tile_X8Y11_LUT4AB/S1END[1]
+ Tile_X8Y11_LUT4AB/S1END[2] Tile_X8Y11_LUT4AB/S1END[3] Tile_X8Y9_LUT4AB/S1BEG[0]
+ Tile_X8Y9_LUT4AB/S1BEG[1] Tile_X8Y9_LUT4AB/S1BEG[2] Tile_X8Y9_LUT4AB/S1BEG[3] Tile_X8Y11_LUT4AB/S2MID[0]
+ Tile_X8Y11_LUT4AB/S2MID[1] Tile_X8Y11_LUT4AB/S2MID[2] Tile_X8Y11_LUT4AB/S2MID[3]
+ Tile_X8Y11_LUT4AB/S2MID[4] Tile_X8Y11_LUT4AB/S2MID[5] Tile_X8Y11_LUT4AB/S2MID[6]
+ Tile_X8Y11_LUT4AB/S2MID[7] Tile_X8Y11_LUT4AB/S2END[0] Tile_X8Y11_LUT4AB/S2END[1]
+ Tile_X8Y11_LUT4AB/S2END[2] Tile_X8Y11_LUT4AB/S2END[3] Tile_X8Y11_LUT4AB/S2END[4]
+ Tile_X8Y11_LUT4AB/S2END[5] Tile_X8Y11_LUT4AB/S2END[6] Tile_X8Y11_LUT4AB/S2END[7]
+ Tile_X8Y9_LUT4AB/S2BEGb[0] Tile_X8Y9_LUT4AB/S2BEGb[1] Tile_X8Y9_LUT4AB/S2BEGb[2]
+ Tile_X8Y9_LUT4AB/S2BEGb[3] Tile_X8Y9_LUT4AB/S2BEGb[4] Tile_X8Y9_LUT4AB/S2BEGb[5]
+ Tile_X8Y9_LUT4AB/S2BEGb[6] Tile_X8Y9_LUT4AB/S2BEGb[7] Tile_X8Y9_LUT4AB/S2BEG[0]
+ Tile_X8Y9_LUT4AB/S2BEG[1] Tile_X8Y9_LUT4AB/S2BEG[2] Tile_X8Y9_LUT4AB/S2BEG[3] Tile_X8Y9_LUT4AB/S2BEG[4]
+ Tile_X8Y9_LUT4AB/S2BEG[5] Tile_X8Y9_LUT4AB/S2BEG[6] Tile_X8Y9_LUT4AB/S2BEG[7] Tile_X8Y11_LUT4AB/S4END[0]
+ Tile_X8Y11_LUT4AB/S4END[10] Tile_X8Y11_LUT4AB/S4END[11] Tile_X8Y11_LUT4AB/S4END[12]
+ Tile_X8Y11_LUT4AB/S4END[13] Tile_X8Y11_LUT4AB/S4END[14] Tile_X8Y11_LUT4AB/S4END[15]
+ Tile_X8Y11_LUT4AB/S4END[1] Tile_X8Y11_LUT4AB/S4END[2] Tile_X8Y11_LUT4AB/S4END[3]
+ Tile_X8Y11_LUT4AB/S4END[4] Tile_X8Y11_LUT4AB/S4END[5] Tile_X8Y11_LUT4AB/S4END[6]
+ Tile_X8Y11_LUT4AB/S4END[7] Tile_X8Y11_LUT4AB/S4END[8] Tile_X8Y11_LUT4AB/S4END[9]
+ Tile_X8Y9_LUT4AB/S4BEG[0] Tile_X8Y9_LUT4AB/S4BEG[10] Tile_X8Y9_LUT4AB/S4BEG[11]
+ Tile_X8Y9_LUT4AB/S4BEG[12] Tile_X8Y9_LUT4AB/S4BEG[13] Tile_X8Y9_LUT4AB/S4BEG[14]
+ Tile_X8Y9_LUT4AB/S4BEG[15] Tile_X8Y9_LUT4AB/S4BEG[1] Tile_X8Y9_LUT4AB/S4BEG[2] Tile_X8Y9_LUT4AB/S4BEG[3]
+ Tile_X8Y9_LUT4AB/S4BEG[4] Tile_X8Y9_LUT4AB/S4BEG[5] Tile_X8Y9_LUT4AB/S4BEG[6] Tile_X8Y9_LUT4AB/S4BEG[7]
+ Tile_X8Y9_LUT4AB/S4BEG[8] Tile_X8Y9_LUT4AB/S4BEG[9] Tile_X8Y11_LUT4AB/SS4END[0]
+ Tile_X8Y11_LUT4AB/SS4END[10] Tile_X8Y11_LUT4AB/SS4END[11] Tile_X8Y11_LUT4AB/SS4END[12]
+ Tile_X8Y11_LUT4AB/SS4END[13] Tile_X8Y11_LUT4AB/SS4END[14] Tile_X8Y11_LUT4AB/SS4END[15]
+ Tile_X8Y11_LUT4AB/SS4END[1] Tile_X8Y11_LUT4AB/SS4END[2] Tile_X8Y11_LUT4AB/SS4END[3]
+ Tile_X8Y11_LUT4AB/SS4END[4] Tile_X8Y11_LUT4AB/SS4END[5] Tile_X8Y11_LUT4AB/SS4END[6]
+ Tile_X8Y11_LUT4AB/SS4END[7] Tile_X8Y11_LUT4AB/SS4END[8] Tile_X8Y11_LUT4AB/SS4END[9]
+ Tile_X8Y9_LUT4AB/SS4BEG[0] Tile_X8Y9_LUT4AB/SS4BEG[10] Tile_X8Y9_LUT4AB/SS4BEG[11]
+ Tile_X8Y9_LUT4AB/SS4BEG[12] Tile_X8Y9_LUT4AB/SS4BEG[13] Tile_X8Y9_LUT4AB/SS4BEG[14]
+ Tile_X8Y9_LUT4AB/SS4BEG[15] Tile_X8Y9_LUT4AB/SS4BEG[1] Tile_X8Y9_LUT4AB/SS4BEG[2]
+ Tile_X8Y9_LUT4AB/SS4BEG[3] Tile_X8Y9_LUT4AB/SS4BEG[4] Tile_X8Y9_LUT4AB/SS4BEG[5]
+ Tile_X8Y9_LUT4AB/SS4BEG[6] Tile_X8Y9_LUT4AB/SS4BEG[7] Tile_X8Y9_LUT4AB/SS4BEG[8]
+ Tile_X8Y9_LUT4AB/SS4BEG[9] Tile_X8Y10_LUT4AB/UserCLK Tile_X8Y9_LUT4AB/UserCLK VGND
+ VPWR Tile_X8Y10_LUT4AB/W1BEG[0] Tile_X8Y10_LUT4AB/W1BEG[1] Tile_X8Y10_LUT4AB/W1BEG[2]
+ Tile_X8Y10_LUT4AB/W1BEG[3] Tile_X9Y10_LUT4AB/W1BEG[0] Tile_X9Y10_LUT4AB/W1BEG[1]
+ Tile_X9Y10_LUT4AB/W1BEG[2] Tile_X9Y10_LUT4AB/W1BEG[3] Tile_X8Y10_LUT4AB/W2BEG[0]
+ Tile_X8Y10_LUT4AB/W2BEG[1] Tile_X8Y10_LUT4AB/W2BEG[2] Tile_X8Y10_LUT4AB/W2BEG[3]
+ Tile_X8Y10_LUT4AB/W2BEG[4] Tile_X8Y10_LUT4AB/W2BEG[5] Tile_X8Y10_LUT4AB/W2BEG[6]
+ Tile_X8Y10_LUT4AB/W2BEG[7] Tile_X8Y10_LUT4AB/W2BEGb[0] Tile_X8Y10_LUT4AB/W2BEGb[1]
+ Tile_X8Y10_LUT4AB/W2BEGb[2] Tile_X8Y10_LUT4AB/W2BEGb[3] Tile_X8Y10_LUT4AB/W2BEGb[4]
+ Tile_X8Y10_LUT4AB/W2BEGb[5] Tile_X8Y10_LUT4AB/W2BEGb[6] Tile_X8Y10_LUT4AB/W2BEGb[7]
+ Tile_X8Y10_LUT4AB/W2END[0] Tile_X8Y10_LUT4AB/W2END[1] Tile_X8Y10_LUT4AB/W2END[2]
+ Tile_X8Y10_LUT4AB/W2END[3] Tile_X8Y10_LUT4AB/W2END[4] Tile_X8Y10_LUT4AB/W2END[5]
+ Tile_X8Y10_LUT4AB/W2END[6] Tile_X8Y10_LUT4AB/W2END[7] Tile_X9Y10_LUT4AB/W2BEG[0]
+ Tile_X9Y10_LUT4AB/W2BEG[1] Tile_X9Y10_LUT4AB/W2BEG[2] Tile_X9Y10_LUT4AB/W2BEG[3]
+ Tile_X9Y10_LUT4AB/W2BEG[4] Tile_X9Y10_LUT4AB/W2BEG[5] Tile_X9Y10_LUT4AB/W2BEG[6]
+ Tile_X9Y10_LUT4AB/W2BEG[7] Tile_X8Y10_LUT4AB/W6BEG[0] Tile_X8Y10_LUT4AB/W6BEG[10]
+ Tile_X8Y10_LUT4AB/W6BEG[11] Tile_X8Y10_LUT4AB/W6BEG[1] Tile_X8Y10_LUT4AB/W6BEG[2]
+ Tile_X8Y10_LUT4AB/W6BEG[3] Tile_X8Y10_LUT4AB/W6BEG[4] Tile_X8Y10_LUT4AB/W6BEG[5]
+ Tile_X8Y10_LUT4AB/W6BEG[6] Tile_X8Y10_LUT4AB/W6BEG[7] Tile_X8Y10_LUT4AB/W6BEG[8]
+ Tile_X8Y10_LUT4AB/W6BEG[9] Tile_X9Y10_LUT4AB/W6BEG[0] Tile_X9Y10_LUT4AB/W6BEG[10]
+ Tile_X9Y10_LUT4AB/W6BEG[11] Tile_X9Y10_LUT4AB/W6BEG[1] Tile_X9Y10_LUT4AB/W6BEG[2]
+ Tile_X9Y10_LUT4AB/W6BEG[3] Tile_X9Y10_LUT4AB/W6BEG[4] Tile_X9Y10_LUT4AB/W6BEG[5]
+ Tile_X9Y10_LUT4AB/W6BEG[6] Tile_X9Y10_LUT4AB/W6BEG[7] Tile_X9Y10_LUT4AB/W6BEG[8]
+ Tile_X9Y10_LUT4AB/W6BEG[9] Tile_X8Y10_LUT4AB/WW4BEG[0] Tile_X8Y10_LUT4AB/WW4BEG[10]
+ Tile_X8Y10_LUT4AB/WW4BEG[11] Tile_X8Y10_LUT4AB/WW4BEG[12] Tile_X8Y10_LUT4AB/WW4BEG[13]
+ Tile_X8Y10_LUT4AB/WW4BEG[14] Tile_X8Y10_LUT4AB/WW4BEG[15] Tile_X8Y10_LUT4AB/WW4BEG[1]
+ Tile_X8Y10_LUT4AB/WW4BEG[2] Tile_X8Y10_LUT4AB/WW4BEG[3] Tile_X8Y10_LUT4AB/WW4BEG[4]
+ Tile_X8Y10_LUT4AB/WW4BEG[5] Tile_X8Y10_LUT4AB/WW4BEG[6] Tile_X8Y10_LUT4AB/WW4BEG[7]
+ Tile_X8Y10_LUT4AB/WW4BEG[8] Tile_X8Y10_LUT4AB/WW4BEG[9] Tile_X9Y10_LUT4AB/WW4BEG[0]
+ Tile_X9Y10_LUT4AB/WW4BEG[10] Tile_X9Y10_LUT4AB/WW4BEG[11] Tile_X9Y10_LUT4AB/WW4BEG[12]
+ Tile_X9Y10_LUT4AB/WW4BEG[13] Tile_X9Y10_LUT4AB/WW4BEG[14] Tile_X9Y10_LUT4AB/WW4BEG[15]
+ Tile_X9Y10_LUT4AB/WW4BEG[1] Tile_X9Y10_LUT4AB/WW4BEG[2] Tile_X9Y10_LUT4AB/WW4BEG[3]
+ Tile_X9Y10_LUT4AB/WW4BEG[4] Tile_X9Y10_LUT4AB/WW4BEG[5] Tile_X9Y10_LUT4AB/WW4BEG[6]
+ Tile_X9Y10_LUT4AB/WW4BEG[7] Tile_X9Y10_LUT4AB/WW4BEG[8] Tile_X9Y10_LUT4AB/WW4BEG[9]
+ LUT4AB
XTile_X1Y4_LUT4AB Tile_X1Y5_LUT4AB/Co Tile_X1Y4_LUT4AB/Co Tile_X2Y4_LUT4AB/E1END[0]
+ Tile_X2Y4_LUT4AB/E1END[1] Tile_X2Y4_LUT4AB/E1END[2] Tile_X2Y4_LUT4AB/E1END[3] Tile_X0Y4_W_IO/E1BEG[0]
+ Tile_X0Y4_W_IO/E1BEG[1] Tile_X0Y4_W_IO/E1BEG[2] Tile_X0Y4_W_IO/E1BEG[3] Tile_X2Y4_LUT4AB/E2MID[0]
+ Tile_X2Y4_LUT4AB/E2MID[1] Tile_X2Y4_LUT4AB/E2MID[2] Tile_X2Y4_LUT4AB/E2MID[3] Tile_X2Y4_LUT4AB/E2MID[4]
+ Tile_X2Y4_LUT4AB/E2MID[5] Tile_X2Y4_LUT4AB/E2MID[6] Tile_X2Y4_LUT4AB/E2MID[7] Tile_X2Y4_LUT4AB/E2END[0]
+ Tile_X2Y4_LUT4AB/E2END[1] Tile_X2Y4_LUT4AB/E2END[2] Tile_X2Y4_LUT4AB/E2END[3] Tile_X2Y4_LUT4AB/E2END[4]
+ Tile_X2Y4_LUT4AB/E2END[5] Tile_X2Y4_LUT4AB/E2END[6] Tile_X2Y4_LUT4AB/E2END[7] Tile_X0Y4_W_IO/E2BEGb[0]
+ Tile_X0Y4_W_IO/E2BEGb[1] Tile_X0Y4_W_IO/E2BEGb[2] Tile_X0Y4_W_IO/E2BEGb[3] Tile_X0Y4_W_IO/E2BEGb[4]
+ Tile_X0Y4_W_IO/E2BEGb[5] Tile_X0Y4_W_IO/E2BEGb[6] Tile_X0Y4_W_IO/E2BEGb[7] Tile_X0Y4_W_IO/E2BEG[0]
+ Tile_X0Y4_W_IO/E2BEG[1] Tile_X0Y4_W_IO/E2BEG[2] Tile_X0Y4_W_IO/E2BEG[3] Tile_X0Y4_W_IO/E2BEG[4]
+ Tile_X0Y4_W_IO/E2BEG[5] Tile_X0Y4_W_IO/E2BEG[6] Tile_X0Y4_W_IO/E2BEG[7] Tile_X2Y4_LUT4AB/E6END[0]
+ Tile_X2Y4_LUT4AB/E6END[10] Tile_X2Y4_LUT4AB/E6END[11] Tile_X2Y4_LUT4AB/E6END[1]
+ Tile_X2Y4_LUT4AB/E6END[2] Tile_X2Y4_LUT4AB/E6END[3] Tile_X2Y4_LUT4AB/E6END[4] Tile_X2Y4_LUT4AB/E6END[5]
+ Tile_X2Y4_LUT4AB/E6END[6] Tile_X2Y4_LUT4AB/E6END[7] Tile_X2Y4_LUT4AB/E6END[8] Tile_X2Y4_LUT4AB/E6END[9]
+ Tile_X0Y4_W_IO/E6BEG[0] Tile_X0Y4_W_IO/E6BEG[10] Tile_X0Y4_W_IO/E6BEG[11] Tile_X0Y4_W_IO/E6BEG[1]
+ Tile_X0Y4_W_IO/E6BEG[2] Tile_X0Y4_W_IO/E6BEG[3] Tile_X0Y4_W_IO/E6BEG[4] Tile_X0Y4_W_IO/E6BEG[5]
+ Tile_X0Y4_W_IO/E6BEG[6] Tile_X0Y4_W_IO/E6BEG[7] Tile_X0Y4_W_IO/E6BEG[8] Tile_X0Y4_W_IO/E6BEG[9]
+ Tile_X2Y4_LUT4AB/EE4END[0] Tile_X2Y4_LUT4AB/EE4END[10] Tile_X2Y4_LUT4AB/EE4END[11]
+ Tile_X2Y4_LUT4AB/EE4END[12] Tile_X2Y4_LUT4AB/EE4END[13] Tile_X2Y4_LUT4AB/EE4END[14]
+ Tile_X2Y4_LUT4AB/EE4END[15] Tile_X2Y4_LUT4AB/EE4END[1] Tile_X2Y4_LUT4AB/EE4END[2]
+ Tile_X2Y4_LUT4AB/EE4END[3] Tile_X2Y4_LUT4AB/EE4END[4] Tile_X2Y4_LUT4AB/EE4END[5]
+ Tile_X2Y4_LUT4AB/EE4END[6] Tile_X2Y4_LUT4AB/EE4END[7] Tile_X2Y4_LUT4AB/EE4END[8]
+ Tile_X2Y4_LUT4AB/EE4END[9] Tile_X0Y4_W_IO/EE4BEG[0] Tile_X0Y4_W_IO/EE4BEG[10] Tile_X0Y4_W_IO/EE4BEG[11]
+ Tile_X0Y4_W_IO/EE4BEG[12] Tile_X0Y4_W_IO/EE4BEG[13] Tile_X0Y4_W_IO/EE4BEG[14] Tile_X0Y4_W_IO/EE4BEG[15]
+ Tile_X0Y4_W_IO/EE4BEG[1] Tile_X0Y4_W_IO/EE4BEG[2] Tile_X0Y4_W_IO/EE4BEG[3] Tile_X0Y4_W_IO/EE4BEG[4]
+ Tile_X0Y4_W_IO/EE4BEG[5] Tile_X0Y4_W_IO/EE4BEG[6] Tile_X0Y4_W_IO/EE4BEG[7] Tile_X0Y4_W_IO/EE4BEG[8]
+ Tile_X0Y4_W_IO/EE4BEG[9] Tile_X1Y4_LUT4AB/FrameData[0] Tile_X1Y4_LUT4AB/FrameData[10]
+ Tile_X1Y4_LUT4AB/FrameData[11] Tile_X1Y4_LUT4AB/FrameData[12] Tile_X1Y4_LUT4AB/FrameData[13]
+ Tile_X1Y4_LUT4AB/FrameData[14] Tile_X1Y4_LUT4AB/FrameData[15] Tile_X1Y4_LUT4AB/FrameData[16]
+ Tile_X1Y4_LUT4AB/FrameData[17] Tile_X1Y4_LUT4AB/FrameData[18] Tile_X1Y4_LUT4AB/FrameData[19]
+ Tile_X1Y4_LUT4AB/FrameData[1] Tile_X1Y4_LUT4AB/FrameData[20] Tile_X1Y4_LUT4AB/FrameData[21]
+ Tile_X1Y4_LUT4AB/FrameData[22] Tile_X1Y4_LUT4AB/FrameData[23] Tile_X1Y4_LUT4AB/FrameData[24]
+ Tile_X1Y4_LUT4AB/FrameData[25] Tile_X1Y4_LUT4AB/FrameData[26] Tile_X1Y4_LUT4AB/FrameData[27]
+ Tile_X1Y4_LUT4AB/FrameData[28] Tile_X1Y4_LUT4AB/FrameData[29] Tile_X1Y4_LUT4AB/FrameData[2]
+ Tile_X1Y4_LUT4AB/FrameData[30] Tile_X1Y4_LUT4AB/FrameData[31] Tile_X1Y4_LUT4AB/FrameData[3]
+ Tile_X1Y4_LUT4AB/FrameData[4] Tile_X1Y4_LUT4AB/FrameData[5] Tile_X1Y4_LUT4AB/FrameData[6]
+ Tile_X1Y4_LUT4AB/FrameData[7] Tile_X1Y4_LUT4AB/FrameData[8] Tile_X1Y4_LUT4AB/FrameData[9]
+ Tile_X2Y4_LUT4AB/FrameData[0] Tile_X2Y4_LUT4AB/FrameData[10] Tile_X2Y4_LUT4AB/FrameData[11]
+ Tile_X2Y4_LUT4AB/FrameData[12] Tile_X2Y4_LUT4AB/FrameData[13] Tile_X2Y4_LUT4AB/FrameData[14]
+ Tile_X2Y4_LUT4AB/FrameData[15] Tile_X2Y4_LUT4AB/FrameData[16] Tile_X2Y4_LUT4AB/FrameData[17]
+ Tile_X2Y4_LUT4AB/FrameData[18] Tile_X2Y4_LUT4AB/FrameData[19] Tile_X2Y4_LUT4AB/FrameData[1]
+ Tile_X2Y4_LUT4AB/FrameData[20] Tile_X2Y4_LUT4AB/FrameData[21] Tile_X2Y4_LUT4AB/FrameData[22]
+ Tile_X2Y4_LUT4AB/FrameData[23] Tile_X2Y4_LUT4AB/FrameData[24] Tile_X2Y4_LUT4AB/FrameData[25]
+ Tile_X2Y4_LUT4AB/FrameData[26] Tile_X2Y4_LUT4AB/FrameData[27] Tile_X2Y4_LUT4AB/FrameData[28]
+ Tile_X2Y4_LUT4AB/FrameData[29] Tile_X2Y4_LUT4AB/FrameData[2] Tile_X2Y4_LUT4AB/FrameData[30]
+ Tile_X2Y4_LUT4AB/FrameData[31] Tile_X2Y4_LUT4AB/FrameData[3] Tile_X2Y4_LUT4AB/FrameData[4]
+ Tile_X2Y4_LUT4AB/FrameData[5] Tile_X2Y4_LUT4AB/FrameData[6] Tile_X2Y4_LUT4AB/FrameData[7]
+ Tile_X2Y4_LUT4AB/FrameData[8] Tile_X2Y4_LUT4AB/FrameData[9] Tile_X1Y4_LUT4AB/FrameStrobe[0]
+ Tile_X1Y4_LUT4AB/FrameStrobe[10] Tile_X1Y4_LUT4AB/FrameStrobe[11] Tile_X1Y4_LUT4AB/FrameStrobe[12]
+ Tile_X1Y4_LUT4AB/FrameStrobe[13] Tile_X1Y4_LUT4AB/FrameStrobe[14] Tile_X1Y4_LUT4AB/FrameStrobe[15]
+ Tile_X1Y4_LUT4AB/FrameStrobe[16] Tile_X1Y4_LUT4AB/FrameStrobe[17] Tile_X1Y4_LUT4AB/FrameStrobe[18]
+ Tile_X1Y4_LUT4AB/FrameStrobe[19] Tile_X1Y4_LUT4AB/FrameStrobe[1] Tile_X1Y4_LUT4AB/FrameStrobe[2]
+ Tile_X1Y4_LUT4AB/FrameStrobe[3] Tile_X1Y4_LUT4AB/FrameStrobe[4] Tile_X1Y4_LUT4AB/FrameStrobe[5]
+ Tile_X1Y4_LUT4AB/FrameStrobe[6] Tile_X1Y4_LUT4AB/FrameStrobe[7] Tile_X1Y4_LUT4AB/FrameStrobe[8]
+ Tile_X1Y4_LUT4AB/FrameStrobe[9] Tile_X1Y3_LUT4AB/FrameStrobe[0] Tile_X1Y3_LUT4AB/FrameStrobe[10]
+ Tile_X1Y3_LUT4AB/FrameStrobe[11] Tile_X1Y3_LUT4AB/FrameStrobe[12] Tile_X1Y3_LUT4AB/FrameStrobe[13]
+ Tile_X1Y3_LUT4AB/FrameStrobe[14] Tile_X1Y3_LUT4AB/FrameStrobe[15] Tile_X1Y3_LUT4AB/FrameStrobe[16]
+ Tile_X1Y3_LUT4AB/FrameStrobe[17] Tile_X1Y3_LUT4AB/FrameStrobe[18] Tile_X1Y3_LUT4AB/FrameStrobe[19]
+ Tile_X1Y3_LUT4AB/FrameStrobe[1] Tile_X1Y3_LUT4AB/FrameStrobe[2] Tile_X1Y3_LUT4AB/FrameStrobe[3]
+ Tile_X1Y3_LUT4AB/FrameStrobe[4] Tile_X1Y3_LUT4AB/FrameStrobe[5] Tile_X1Y3_LUT4AB/FrameStrobe[6]
+ Tile_X1Y3_LUT4AB/FrameStrobe[7] Tile_X1Y3_LUT4AB/FrameStrobe[8] Tile_X1Y3_LUT4AB/FrameStrobe[9]
+ Tile_X1Y4_LUT4AB/N1BEG[0] Tile_X1Y4_LUT4AB/N1BEG[1] Tile_X1Y4_LUT4AB/N1BEG[2] Tile_X1Y4_LUT4AB/N1BEG[3]
+ Tile_X1Y5_LUT4AB/N1BEG[0] Tile_X1Y5_LUT4AB/N1BEG[1] Tile_X1Y5_LUT4AB/N1BEG[2] Tile_X1Y5_LUT4AB/N1BEG[3]
+ Tile_X1Y4_LUT4AB/N2BEG[0] Tile_X1Y4_LUT4AB/N2BEG[1] Tile_X1Y4_LUT4AB/N2BEG[2] Tile_X1Y4_LUT4AB/N2BEG[3]
+ Tile_X1Y4_LUT4AB/N2BEG[4] Tile_X1Y4_LUT4AB/N2BEG[5] Tile_X1Y4_LUT4AB/N2BEG[6] Tile_X1Y4_LUT4AB/N2BEG[7]
+ Tile_X1Y3_LUT4AB/N2END[0] Tile_X1Y3_LUT4AB/N2END[1] Tile_X1Y3_LUT4AB/N2END[2] Tile_X1Y3_LUT4AB/N2END[3]
+ Tile_X1Y3_LUT4AB/N2END[4] Tile_X1Y3_LUT4AB/N2END[5] Tile_X1Y3_LUT4AB/N2END[6] Tile_X1Y3_LUT4AB/N2END[7]
+ Tile_X1Y4_LUT4AB/N2END[0] Tile_X1Y4_LUT4AB/N2END[1] Tile_X1Y4_LUT4AB/N2END[2] Tile_X1Y4_LUT4AB/N2END[3]
+ Tile_X1Y4_LUT4AB/N2END[4] Tile_X1Y4_LUT4AB/N2END[5] Tile_X1Y4_LUT4AB/N2END[6] Tile_X1Y4_LUT4AB/N2END[7]
+ Tile_X1Y5_LUT4AB/N2BEG[0] Tile_X1Y5_LUT4AB/N2BEG[1] Tile_X1Y5_LUT4AB/N2BEG[2] Tile_X1Y5_LUT4AB/N2BEG[3]
+ Tile_X1Y5_LUT4AB/N2BEG[4] Tile_X1Y5_LUT4AB/N2BEG[5] Tile_X1Y5_LUT4AB/N2BEG[6] Tile_X1Y5_LUT4AB/N2BEG[7]
+ Tile_X1Y4_LUT4AB/N4BEG[0] Tile_X1Y4_LUT4AB/N4BEG[10] Tile_X1Y4_LUT4AB/N4BEG[11]
+ Tile_X1Y4_LUT4AB/N4BEG[12] Tile_X1Y4_LUT4AB/N4BEG[13] Tile_X1Y4_LUT4AB/N4BEG[14]
+ Tile_X1Y4_LUT4AB/N4BEG[15] Tile_X1Y4_LUT4AB/N4BEG[1] Tile_X1Y4_LUT4AB/N4BEG[2] Tile_X1Y4_LUT4AB/N4BEG[3]
+ Tile_X1Y4_LUT4AB/N4BEG[4] Tile_X1Y4_LUT4AB/N4BEG[5] Tile_X1Y4_LUT4AB/N4BEG[6] Tile_X1Y4_LUT4AB/N4BEG[7]
+ Tile_X1Y4_LUT4AB/N4BEG[8] Tile_X1Y4_LUT4AB/N4BEG[9] Tile_X1Y5_LUT4AB/N4BEG[0] Tile_X1Y5_LUT4AB/N4BEG[10]
+ Tile_X1Y5_LUT4AB/N4BEG[11] Tile_X1Y5_LUT4AB/N4BEG[12] Tile_X1Y5_LUT4AB/N4BEG[13]
+ Tile_X1Y5_LUT4AB/N4BEG[14] Tile_X1Y5_LUT4AB/N4BEG[15] Tile_X1Y5_LUT4AB/N4BEG[1]
+ Tile_X1Y5_LUT4AB/N4BEG[2] Tile_X1Y5_LUT4AB/N4BEG[3] Tile_X1Y5_LUT4AB/N4BEG[4] Tile_X1Y5_LUT4AB/N4BEG[5]
+ Tile_X1Y5_LUT4AB/N4BEG[6] Tile_X1Y5_LUT4AB/N4BEG[7] Tile_X1Y5_LUT4AB/N4BEG[8] Tile_X1Y5_LUT4AB/N4BEG[9]
+ Tile_X1Y4_LUT4AB/NN4BEG[0] Tile_X1Y4_LUT4AB/NN4BEG[10] Tile_X1Y4_LUT4AB/NN4BEG[11]
+ Tile_X1Y4_LUT4AB/NN4BEG[12] Tile_X1Y4_LUT4AB/NN4BEG[13] Tile_X1Y4_LUT4AB/NN4BEG[14]
+ Tile_X1Y4_LUT4AB/NN4BEG[15] Tile_X1Y4_LUT4AB/NN4BEG[1] Tile_X1Y4_LUT4AB/NN4BEG[2]
+ Tile_X1Y4_LUT4AB/NN4BEG[3] Tile_X1Y4_LUT4AB/NN4BEG[4] Tile_X1Y4_LUT4AB/NN4BEG[5]
+ Tile_X1Y4_LUT4AB/NN4BEG[6] Tile_X1Y4_LUT4AB/NN4BEG[7] Tile_X1Y4_LUT4AB/NN4BEG[8]
+ Tile_X1Y4_LUT4AB/NN4BEG[9] Tile_X1Y5_LUT4AB/NN4BEG[0] Tile_X1Y5_LUT4AB/NN4BEG[10]
+ Tile_X1Y5_LUT4AB/NN4BEG[11] Tile_X1Y5_LUT4AB/NN4BEG[12] Tile_X1Y5_LUT4AB/NN4BEG[13]
+ Tile_X1Y5_LUT4AB/NN4BEG[14] Tile_X1Y5_LUT4AB/NN4BEG[15] Tile_X1Y5_LUT4AB/NN4BEG[1]
+ Tile_X1Y5_LUT4AB/NN4BEG[2] Tile_X1Y5_LUT4AB/NN4BEG[3] Tile_X1Y5_LUT4AB/NN4BEG[4]
+ Tile_X1Y5_LUT4AB/NN4BEG[5] Tile_X1Y5_LUT4AB/NN4BEG[6] Tile_X1Y5_LUT4AB/NN4BEG[7]
+ Tile_X1Y5_LUT4AB/NN4BEG[8] Tile_X1Y5_LUT4AB/NN4BEG[9] Tile_X1Y5_LUT4AB/S1END[0]
+ Tile_X1Y5_LUT4AB/S1END[1] Tile_X1Y5_LUT4AB/S1END[2] Tile_X1Y5_LUT4AB/S1END[3] Tile_X1Y4_LUT4AB/S1END[0]
+ Tile_X1Y4_LUT4AB/S1END[1] Tile_X1Y4_LUT4AB/S1END[2] Tile_X1Y4_LUT4AB/S1END[3] Tile_X1Y5_LUT4AB/S2MID[0]
+ Tile_X1Y5_LUT4AB/S2MID[1] Tile_X1Y5_LUT4AB/S2MID[2] Tile_X1Y5_LUT4AB/S2MID[3] Tile_X1Y5_LUT4AB/S2MID[4]
+ Tile_X1Y5_LUT4AB/S2MID[5] Tile_X1Y5_LUT4AB/S2MID[6] Tile_X1Y5_LUT4AB/S2MID[7] Tile_X1Y5_LUT4AB/S2END[0]
+ Tile_X1Y5_LUT4AB/S2END[1] Tile_X1Y5_LUT4AB/S2END[2] Tile_X1Y5_LUT4AB/S2END[3] Tile_X1Y5_LUT4AB/S2END[4]
+ Tile_X1Y5_LUT4AB/S2END[5] Tile_X1Y5_LUT4AB/S2END[6] Tile_X1Y5_LUT4AB/S2END[7] Tile_X1Y4_LUT4AB/S2END[0]
+ Tile_X1Y4_LUT4AB/S2END[1] Tile_X1Y4_LUT4AB/S2END[2] Tile_X1Y4_LUT4AB/S2END[3] Tile_X1Y4_LUT4AB/S2END[4]
+ Tile_X1Y4_LUT4AB/S2END[5] Tile_X1Y4_LUT4AB/S2END[6] Tile_X1Y4_LUT4AB/S2END[7] Tile_X1Y4_LUT4AB/S2MID[0]
+ Tile_X1Y4_LUT4AB/S2MID[1] Tile_X1Y4_LUT4AB/S2MID[2] Tile_X1Y4_LUT4AB/S2MID[3] Tile_X1Y4_LUT4AB/S2MID[4]
+ Tile_X1Y4_LUT4AB/S2MID[5] Tile_X1Y4_LUT4AB/S2MID[6] Tile_X1Y4_LUT4AB/S2MID[7] Tile_X1Y5_LUT4AB/S4END[0]
+ Tile_X1Y5_LUT4AB/S4END[10] Tile_X1Y5_LUT4AB/S4END[11] Tile_X1Y5_LUT4AB/S4END[12]
+ Tile_X1Y5_LUT4AB/S4END[13] Tile_X1Y5_LUT4AB/S4END[14] Tile_X1Y5_LUT4AB/S4END[15]
+ Tile_X1Y5_LUT4AB/S4END[1] Tile_X1Y5_LUT4AB/S4END[2] Tile_X1Y5_LUT4AB/S4END[3] Tile_X1Y5_LUT4AB/S4END[4]
+ Tile_X1Y5_LUT4AB/S4END[5] Tile_X1Y5_LUT4AB/S4END[6] Tile_X1Y5_LUT4AB/S4END[7] Tile_X1Y5_LUT4AB/S4END[8]
+ Tile_X1Y5_LUT4AB/S4END[9] Tile_X1Y4_LUT4AB/S4END[0] Tile_X1Y4_LUT4AB/S4END[10] Tile_X1Y4_LUT4AB/S4END[11]
+ Tile_X1Y4_LUT4AB/S4END[12] Tile_X1Y4_LUT4AB/S4END[13] Tile_X1Y4_LUT4AB/S4END[14]
+ Tile_X1Y4_LUT4AB/S4END[15] Tile_X1Y4_LUT4AB/S4END[1] Tile_X1Y4_LUT4AB/S4END[2] Tile_X1Y4_LUT4AB/S4END[3]
+ Tile_X1Y4_LUT4AB/S4END[4] Tile_X1Y4_LUT4AB/S4END[5] Tile_X1Y4_LUT4AB/S4END[6] Tile_X1Y4_LUT4AB/S4END[7]
+ Tile_X1Y4_LUT4AB/S4END[8] Tile_X1Y4_LUT4AB/S4END[9] Tile_X1Y5_LUT4AB/SS4END[0] Tile_X1Y5_LUT4AB/SS4END[10]
+ Tile_X1Y5_LUT4AB/SS4END[11] Tile_X1Y5_LUT4AB/SS4END[12] Tile_X1Y5_LUT4AB/SS4END[13]
+ Tile_X1Y5_LUT4AB/SS4END[14] Tile_X1Y5_LUT4AB/SS4END[15] Tile_X1Y5_LUT4AB/SS4END[1]
+ Tile_X1Y5_LUT4AB/SS4END[2] Tile_X1Y5_LUT4AB/SS4END[3] Tile_X1Y5_LUT4AB/SS4END[4]
+ Tile_X1Y5_LUT4AB/SS4END[5] Tile_X1Y5_LUT4AB/SS4END[6] Tile_X1Y5_LUT4AB/SS4END[7]
+ Tile_X1Y5_LUT4AB/SS4END[8] Tile_X1Y5_LUT4AB/SS4END[9] Tile_X1Y4_LUT4AB/SS4END[0]
+ Tile_X1Y4_LUT4AB/SS4END[10] Tile_X1Y4_LUT4AB/SS4END[11] Tile_X1Y4_LUT4AB/SS4END[12]
+ Tile_X1Y4_LUT4AB/SS4END[13] Tile_X1Y4_LUT4AB/SS4END[14] Tile_X1Y4_LUT4AB/SS4END[15]
+ Tile_X1Y4_LUT4AB/SS4END[1] Tile_X1Y4_LUT4AB/SS4END[2] Tile_X1Y4_LUT4AB/SS4END[3]
+ Tile_X1Y4_LUT4AB/SS4END[4] Tile_X1Y4_LUT4AB/SS4END[5] Tile_X1Y4_LUT4AB/SS4END[6]
+ Tile_X1Y4_LUT4AB/SS4END[7] Tile_X1Y4_LUT4AB/SS4END[8] Tile_X1Y4_LUT4AB/SS4END[9]
+ Tile_X1Y4_LUT4AB/UserCLK Tile_X1Y3_LUT4AB/UserCLK VGND VPWR Tile_X0Y4_W_IO/W1END[0]
+ Tile_X0Y4_W_IO/W1END[1] Tile_X0Y4_W_IO/W1END[2] Tile_X0Y4_W_IO/W1END[3] Tile_X2Y4_LUT4AB/W1BEG[0]
+ Tile_X2Y4_LUT4AB/W1BEG[1] Tile_X2Y4_LUT4AB/W1BEG[2] Tile_X2Y4_LUT4AB/W1BEG[3] Tile_X0Y4_W_IO/W2MID[0]
+ Tile_X0Y4_W_IO/W2MID[1] Tile_X0Y4_W_IO/W2MID[2] Tile_X0Y4_W_IO/W2MID[3] Tile_X0Y4_W_IO/W2MID[4]
+ Tile_X0Y4_W_IO/W2MID[5] Tile_X0Y4_W_IO/W2MID[6] Tile_X0Y4_W_IO/W2MID[7] Tile_X0Y4_W_IO/W2END[0]
+ Tile_X0Y4_W_IO/W2END[1] Tile_X0Y4_W_IO/W2END[2] Tile_X0Y4_W_IO/W2END[3] Tile_X0Y4_W_IO/W2END[4]
+ Tile_X0Y4_W_IO/W2END[5] Tile_X0Y4_W_IO/W2END[6] Tile_X0Y4_W_IO/W2END[7] Tile_X1Y4_LUT4AB/W2END[0]
+ Tile_X1Y4_LUT4AB/W2END[1] Tile_X1Y4_LUT4AB/W2END[2] Tile_X1Y4_LUT4AB/W2END[3] Tile_X1Y4_LUT4AB/W2END[4]
+ Tile_X1Y4_LUT4AB/W2END[5] Tile_X1Y4_LUT4AB/W2END[6] Tile_X1Y4_LUT4AB/W2END[7] Tile_X2Y4_LUT4AB/W2BEG[0]
+ Tile_X2Y4_LUT4AB/W2BEG[1] Tile_X2Y4_LUT4AB/W2BEG[2] Tile_X2Y4_LUT4AB/W2BEG[3] Tile_X2Y4_LUT4AB/W2BEG[4]
+ Tile_X2Y4_LUT4AB/W2BEG[5] Tile_X2Y4_LUT4AB/W2BEG[6] Tile_X2Y4_LUT4AB/W2BEG[7] Tile_X0Y4_W_IO/W6END[0]
+ Tile_X0Y4_W_IO/W6END[10] Tile_X0Y4_W_IO/W6END[11] Tile_X0Y4_W_IO/W6END[1] Tile_X0Y4_W_IO/W6END[2]
+ Tile_X0Y4_W_IO/W6END[3] Tile_X0Y4_W_IO/W6END[4] Tile_X0Y4_W_IO/W6END[5] Tile_X0Y4_W_IO/W6END[6]
+ Tile_X0Y4_W_IO/W6END[7] Tile_X0Y4_W_IO/W6END[8] Tile_X0Y4_W_IO/W6END[9] Tile_X2Y4_LUT4AB/W6BEG[0]
+ Tile_X2Y4_LUT4AB/W6BEG[10] Tile_X2Y4_LUT4AB/W6BEG[11] Tile_X2Y4_LUT4AB/W6BEG[1]
+ Tile_X2Y4_LUT4AB/W6BEG[2] Tile_X2Y4_LUT4AB/W6BEG[3] Tile_X2Y4_LUT4AB/W6BEG[4] Tile_X2Y4_LUT4AB/W6BEG[5]
+ Tile_X2Y4_LUT4AB/W6BEG[6] Tile_X2Y4_LUT4AB/W6BEG[7] Tile_X2Y4_LUT4AB/W6BEG[8] Tile_X2Y4_LUT4AB/W6BEG[9]
+ Tile_X0Y4_W_IO/WW4END[0] Tile_X0Y4_W_IO/WW4END[10] Tile_X0Y4_W_IO/WW4END[11] Tile_X0Y4_W_IO/WW4END[12]
+ Tile_X0Y4_W_IO/WW4END[13] Tile_X0Y4_W_IO/WW4END[14] Tile_X0Y4_W_IO/WW4END[15] Tile_X0Y4_W_IO/WW4END[1]
+ Tile_X0Y4_W_IO/WW4END[2] Tile_X0Y4_W_IO/WW4END[3] Tile_X0Y4_W_IO/WW4END[4] Tile_X0Y4_W_IO/WW4END[5]
+ Tile_X0Y4_W_IO/WW4END[6] Tile_X0Y4_W_IO/WW4END[7] Tile_X0Y4_W_IO/WW4END[8] Tile_X0Y4_W_IO/WW4END[9]
+ Tile_X2Y4_LUT4AB/WW4BEG[0] Tile_X2Y4_LUT4AB/WW4BEG[10] Tile_X2Y4_LUT4AB/WW4BEG[11]
+ Tile_X2Y4_LUT4AB/WW4BEG[12] Tile_X2Y4_LUT4AB/WW4BEG[13] Tile_X2Y4_LUT4AB/WW4BEG[14]
+ Tile_X2Y4_LUT4AB/WW4BEG[15] Tile_X2Y4_LUT4AB/WW4BEG[1] Tile_X2Y4_LUT4AB/WW4BEG[2]
+ Tile_X2Y4_LUT4AB/WW4BEG[3] Tile_X2Y4_LUT4AB/WW4BEG[4] Tile_X2Y4_LUT4AB/WW4BEG[5]
+ Tile_X2Y4_LUT4AB/WW4BEG[6] Tile_X2Y4_LUT4AB/WW4BEG[7] Tile_X2Y4_LUT4AB/WW4BEG[8]
+ Tile_X2Y4_LUT4AB/WW4BEG[9] LUT4AB
XTile_X6Y13_LUT4AB Tile_X6Y14_LUT4AB/Co Tile_X6Y13_LUT4AB/Co Tile_X6Y13_LUT4AB/E1BEG[0]
+ Tile_X6Y13_LUT4AB/E1BEG[1] Tile_X6Y13_LUT4AB/E1BEG[2] Tile_X6Y13_LUT4AB/E1BEG[3]
+ Tile_X6Y13_LUT4AB/E1END[0] Tile_X6Y13_LUT4AB/E1END[1] Tile_X6Y13_LUT4AB/E1END[2]
+ Tile_X6Y13_LUT4AB/E1END[3] Tile_X6Y13_LUT4AB/E2BEG[0] Tile_X6Y13_LUT4AB/E2BEG[1]
+ Tile_X6Y13_LUT4AB/E2BEG[2] Tile_X6Y13_LUT4AB/E2BEG[3] Tile_X6Y13_LUT4AB/E2BEG[4]
+ Tile_X6Y13_LUT4AB/E2BEG[5] Tile_X6Y13_LUT4AB/E2BEG[6] Tile_X6Y13_LUT4AB/E2BEG[7]
+ Tile_X6Y13_LUT4AB/E2BEGb[0] Tile_X6Y13_LUT4AB/E2BEGb[1] Tile_X6Y13_LUT4AB/E2BEGb[2]
+ Tile_X6Y13_LUT4AB/E2BEGb[3] Tile_X6Y13_LUT4AB/E2BEGb[4] Tile_X6Y13_LUT4AB/E2BEGb[5]
+ Tile_X6Y13_LUT4AB/E2BEGb[6] Tile_X6Y13_LUT4AB/E2BEGb[7] Tile_X6Y13_LUT4AB/E2END[0]
+ Tile_X6Y13_LUT4AB/E2END[1] Tile_X6Y13_LUT4AB/E2END[2] Tile_X6Y13_LUT4AB/E2END[3]
+ Tile_X6Y13_LUT4AB/E2END[4] Tile_X6Y13_LUT4AB/E2END[5] Tile_X6Y13_LUT4AB/E2END[6]
+ Tile_X6Y13_LUT4AB/E2END[7] Tile_X6Y13_LUT4AB/E2MID[0] Tile_X6Y13_LUT4AB/E2MID[1]
+ Tile_X6Y13_LUT4AB/E2MID[2] Tile_X6Y13_LUT4AB/E2MID[3] Tile_X6Y13_LUT4AB/E2MID[4]
+ Tile_X6Y13_LUT4AB/E2MID[5] Tile_X6Y13_LUT4AB/E2MID[6] Tile_X6Y13_LUT4AB/E2MID[7]
+ Tile_X6Y13_LUT4AB/E6BEG[0] Tile_X6Y13_LUT4AB/E6BEG[10] Tile_X6Y13_LUT4AB/E6BEG[11]
+ Tile_X6Y13_LUT4AB/E6BEG[1] Tile_X6Y13_LUT4AB/E6BEG[2] Tile_X6Y13_LUT4AB/E6BEG[3]
+ Tile_X6Y13_LUT4AB/E6BEG[4] Tile_X6Y13_LUT4AB/E6BEG[5] Tile_X6Y13_LUT4AB/E6BEG[6]
+ Tile_X6Y13_LUT4AB/E6BEG[7] Tile_X6Y13_LUT4AB/E6BEG[8] Tile_X6Y13_LUT4AB/E6BEG[9]
+ Tile_X6Y13_LUT4AB/E6END[0] Tile_X6Y13_LUT4AB/E6END[10] Tile_X6Y13_LUT4AB/E6END[11]
+ Tile_X6Y13_LUT4AB/E6END[1] Tile_X6Y13_LUT4AB/E6END[2] Tile_X6Y13_LUT4AB/E6END[3]
+ Tile_X6Y13_LUT4AB/E6END[4] Tile_X6Y13_LUT4AB/E6END[5] Tile_X6Y13_LUT4AB/E6END[6]
+ Tile_X6Y13_LUT4AB/E6END[7] Tile_X6Y13_LUT4AB/E6END[8] Tile_X6Y13_LUT4AB/E6END[9]
+ Tile_X6Y13_LUT4AB/EE4BEG[0] Tile_X6Y13_LUT4AB/EE4BEG[10] Tile_X6Y13_LUT4AB/EE4BEG[11]
+ Tile_X6Y13_LUT4AB/EE4BEG[12] Tile_X6Y13_LUT4AB/EE4BEG[13] Tile_X6Y13_LUT4AB/EE4BEG[14]
+ Tile_X6Y13_LUT4AB/EE4BEG[15] Tile_X6Y13_LUT4AB/EE4BEG[1] Tile_X6Y13_LUT4AB/EE4BEG[2]
+ Tile_X6Y13_LUT4AB/EE4BEG[3] Tile_X6Y13_LUT4AB/EE4BEG[4] Tile_X6Y13_LUT4AB/EE4BEG[5]
+ Tile_X6Y13_LUT4AB/EE4BEG[6] Tile_X6Y13_LUT4AB/EE4BEG[7] Tile_X6Y13_LUT4AB/EE4BEG[8]
+ Tile_X6Y13_LUT4AB/EE4BEG[9] Tile_X6Y13_LUT4AB/EE4END[0] Tile_X6Y13_LUT4AB/EE4END[10]
+ Tile_X6Y13_LUT4AB/EE4END[11] Tile_X6Y13_LUT4AB/EE4END[12] Tile_X6Y13_LUT4AB/EE4END[13]
+ Tile_X6Y13_LUT4AB/EE4END[14] Tile_X6Y13_LUT4AB/EE4END[15] Tile_X6Y13_LUT4AB/EE4END[1]
+ Tile_X6Y13_LUT4AB/EE4END[2] Tile_X6Y13_LUT4AB/EE4END[3] Tile_X6Y13_LUT4AB/EE4END[4]
+ Tile_X6Y13_LUT4AB/EE4END[5] Tile_X6Y13_LUT4AB/EE4END[6] Tile_X6Y13_LUT4AB/EE4END[7]
+ Tile_X6Y13_LUT4AB/EE4END[8] Tile_X6Y13_LUT4AB/EE4END[9] Tile_X6Y13_LUT4AB/FrameData[0]
+ Tile_X6Y13_LUT4AB/FrameData[10] Tile_X6Y13_LUT4AB/FrameData[11] Tile_X6Y13_LUT4AB/FrameData[12]
+ Tile_X6Y13_LUT4AB/FrameData[13] Tile_X6Y13_LUT4AB/FrameData[14] Tile_X6Y13_LUT4AB/FrameData[15]
+ Tile_X6Y13_LUT4AB/FrameData[16] Tile_X6Y13_LUT4AB/FrameData[17] Tile_X6Y13_LUT4AB/FrameData[18]
+ Tile_X6Y13_LUT4AB/FrameData[19] Tile_X6Y13_LUT4AB/FrameData[1] Tile_X6Y13_LUT4AB/FrameData[20]
+ Tile_X6Y13_LUT4AB/FrameData[21] Tile_X6Y13_LUT4AB/FrameData[22] Tile_X6Y13_LUT4AB/FrameData[23]
+ Tile_X6Y13_LUT4AB/FrameData[24] Tile_X6Y13_LUT4AB/FrameData[25] Tile_X6Y13_LUT4AB/FrameData[26]
+ Tile_X6Y13_LUT4AB/FrameData[27] Tile_X6Y13_LUT4AB/FrameData[28] Tile_X6Y13_LUT4AB/FrameData[29]
+ Tile_X6Y13_LUT4AB/FrameData[2] Tile_X6Y13_LUT4AB/FrameData[30] Tile_X6Y13_LUT4AB/FrameData[31]
+ Tile_X6Y13_LUT4AB/FrameData[3] Tile_X6Y13_LUT4AB/FrameData[4] Tile_X6Y13_LUT4AB/FrameData[5]
+ Tile_X6Y13_LUT4AB/FrameData[6] Tile_X6Y13_LUT4AB/FrameData[7] Tile_X6Y13_LUT4AB/FrameData[8]
+ Tile_X6Y13_LUT4AB/FrameData[9] Tile_X6Y13_LUT4AB/FrameData_O[0] Tile_X6Y13_LUT4AB/FrameData_O[10]
+ Tile_X6Y13_LUT4AB/FrameData_O[11] Tile_X6Y13_LUT4AB/FrameData_O[12] Tile_X6Y13_LUT4AB/FrameData_O[13]
+ Tile_X6Y13_LUT4AB/FrameData_O[14] Tile_X6Y13_LUT4AB/FrameData_O[15] Tile_X6Y13_LUT4AB/FrameData_O[16]
+ Tile_X6Y13_LUT4AB/FrameData_O[17] Tile_X6Y13_LUT4AB/FrameData_O[18] Tile_X6Y13_LUT4AB/FrameData_O[19]
+ Tile_X6Y13_LUT4AB/FrameData_O[1] Tile_X6Y13_LUT4AB/FrameData_O[20] Tile_X6Y13_LUT4AB/FrameData_O[21]
+ Tile_X6Y13_LUT4AB/FrameData_O[22] Tile_X6Y13_LUT4AB/FrameData_O[23] Tile_X6Y13_LUT4AB/FrameData_O[24]
+ Tile_X6Y13_LUT4AB/FrameData_O[25] Tile_X6Y13_LUT4AB/FrameData_O[26] Tile_X6Y13_LUT4AB/FrameData_O[27]
+ Tile_X6Y13_LUT4AB/FrameData_O[28] Tile_X6Y13_LUT4AB/FrameData_O[29] Tile_X6Y13_LUT4AB/FrameData_O[2]
+ Tile_X6Y13_LUT4AB/FrameData_O[30] Tile_X6Y13_LUT4AB/FrameData_O[31] Tile_X6Y13_LUT4AB/FrameData_O[3]
+ Tile_X6Y13_LUT4AB/FrameData_O[4] Tile_X6Y13_LUT4AB/FrameData_O[5] Tile_X6Y13_LUT4AB/FrameData_O[6]
+ Tile_X6Y13_LUT4AB/FrameData_O[7] Tile_X6Y13_LUT4AB/FrameData_O[8] Tile_X6Y13_LUT4AB/FrameData_O[9]
+ Tile_X6Y13_LUT4AB/FrameStrobe[0] Tile_X6Y13_LUT4AB/FrameStrobe[10] Tile_X6Y13_LUT4AB/FrameStrobe[11]
+ Tile_X6Y13_LUT4AB/FrameStrobe[12] Tile_X6Y13_LUT4AB/FrameStrobe[13] Tile_X6Y13_LUT4AB/FrameStrobe[14]
+ Tile_X6Y13_LUT4AB/FrameStrobe[15] Tile_X6Y13_LUT4AB/FrameStrobe[16] Tile_X6Y13_LUT4AB/FrameStrobe[17]
+ Tile_X6Y13_LUT4AB/FrameStrobe[18] Tile_X6Y13_LUT4AB/FrameStrobe[19] Tile_X6Y13_LUT4AB/FrameStrobe[1]
+ Tile_X6Y13_LUT4AB/FrameStrobe[2] Tile_X6Y13_LUT4AB/FrameStrobe[3] Tile_X6Y13_LUT4AB/FrameStrobe[4]
+ Tile_X6Y13_LUT4AB/FrameStrobe[5] Tile_X6Y13_LUT4AB/FrameStrobe[6] Tile_X6Y13_LUT4AB/FrameStrobe[7]
+ Tile_X6Y13_LUT4AB/FrameStrobe[8] Tile_X6Y13_LUT4AB/FrameStrobe[9] Tile_X6Y12_LUT4AB/FrameStrobe[0]
+ Tile_X6Y12_LUT4AB/FrameStrobe[10] Tile_X6Y12_LUT4AB/FrameStrobe[11] Tile_X6Y12_LUT4AB/FrameStrobe[12]
+ Tile_X6Y12_LUT4AB/FrameStrobe[13] Tile_X6Y12_LUT4AB/FrameStrobe[14] Tile_X6Y12_LUT4AB/FrameStrobe[15]
+ Tile_X6Y12_LUT4AB/FrameStrobe[16] Tile_X6Y12_LUT4AB/FrameStrobe[17] Tile_X6Y12_LUT4AB/FrameStrobe[18]
+ Tile_X6Y12_LUT4AB/FrameStrobe[19] Tile_X6Y12_LUT4AB/FrameStrobe[1] Tile_X6Y12_LUT4AB/FrameStrobe[2]
+ Tile_X6Y12_LUT4AB/FrameStrobe[3] Tile_X6Y12_LUT4AB/FrameStrobe[4] Tile_X6Y12_LUT4AB/FrameStrobe[5]
+ Tile_X6Y12_LUT4AB/FrameStrobe[6] Tile_X6Y12_LUT4AB/FrameStrobe[7] Tile_X6Y12_LUT4AB/FrameStrobe[8]
+ Tile_X6Y12_LUT4AB/FrameStrobe[9] Tile_X6Y13_LUT4AB/N1BEG[0] Tile_X6Y13_LUT4AB/N1BEG[1]
+ Tile_X6Y13_LUT4AB/N1BEG[2] Tile_X6Y13_LUT4AB/N1BEG[3] Tile_X6Y14_LUT4AB/N1BEG[0]
+ Tile_X6Y14_LUT4AB/N1BEG[1] Tile_X6Y14_LUT4AB/N1BEG[2] Tile_X6Y14_LUT4AB/N1BEG[3]
+ Tile_X6Y13_LUT4AB/N2BEG[0] Tile_X6Y13_LUT4AB/N2BEG[1] Tile_X6Y13_LUT4AB/N2BEG[2]
+ Tile_X6Y13_LUT4AB/N2BEG[3] Tile_X6Y13_LUT4AB/N2BEG[4] Tile_X6Y13_LUT4AB/N2BEG[5]
+ Tile_X6Y13_LUT4AB/N2BEG[6] Tile_X6Y13_LUT4AB/N2BEG[7] Tile_X6Y12_LUT4AB/N2END[0]
+ Tile_X6Y12_LUT4AB/N2END[1] Tile_X6Y12_LUT4AB/N2END[2] Tile_X6Y12_LUT4AB/N2END[3]
+ Tile_X6Y12_LUT4AB/N2END[4] Tile_X6Y12_LUT4AB/N2END[5] Tile_X6Y12_LUT4AB/N2END[6]
+ Tile_X6Y12_LUT4AB/N2END[7] Tile_X6Y13_LUT4AB/N2END[0] Tile_X6Y13_LUT4AB/N2END[1]
+ Tile_X6Y13_LUT4AB/N2END[2] Tile_X6Y13_LUT4AB/N2END[3] Tile_X6Y13_LUT4AB/N2END[4]
+ Tile_X6Y13_LUT4AB/N2END[5] Tile_X6Y13_LUT4AB/N2END[6] Tile_X6Y13_LUT4AB/N2END[7]
+ Tile_X6Y14_LUT4AB/N2BEG[0] Tile_X6Y14_LUT4AB/N2BEG[1] Tile_X6Y14_LUT4AB/N2BEG[2]
+ Tile_X6Y14_LUT4AB/N2BEG[3] Tile_X6Y14_LUT4AB/N2BEG[4] Tile_X6Y14_LUT4AB/N2BEG[5]
+ Tile_X6Y14_LUT4AB/N2BEG[6] Tile_X6Y14_LUT4AB/N2BEG[7] Tile_X6Y13_LUT4AB/N4BEG[0]
+ Tile_X6Y13_LUT4AB/N4BEG[10] Tile_X6Y13_LUT4AB/N4BEG[11] Tile_X6Y13_LUT4AB/N4BEG[12]
+ Tile_X6Y13_LUT4AB/N4BEG[13] Tile_X6Y13_LUT4AB/N4BEG[14] Tile_X6Y13_LUT4AB/N4BEG[15]
+ Tile_X6Y13_LUT4AB/N4BEG[1] Tile_X6Y13_LUT4AB/N4BEG[2] Tile_X6Y13_LUT4AB/N4BEG[3]
+ Tile_X6Y13_LUT4AB/N4BEG[4] Tile_X6Y13_LUT4AB/N4BEG[5] Tile_X6Y13_LUT4AB/N4BEG[6]
+ Tile_X6Y13_LUT4AB/N4BEG[7] Tile_X6Y13_LUT4AB/N4BEG[8] Tile_X6Y13_LUT4AB/N4BEG[9]
+ Tile_X6Y14_LUT4AB/N4BEG[0] Tile_X6Y14_LUT4AB/N4BEG[10] Tile_X6Y14_LUT4AB/N4BEG[11]
+ Tile_X6Y14_LUT4AB/N4BEG[12] Tile_X6Y14_LUT4AB/N4BEG[13] Tile_X6Y14_LUT4AB/N4BEG[14]
+ Tile_X6Y14_LUT4AB/N4BEG[15] Tile_X6Y14_LUT4AB/N4BEG[1] Tile_X6Y14_LUT4AB/N4BEG[2]
+ Tile_X6Y14_LUT4AB/N4BEG[3] Tile_X6Y14_LUT4AB/N4BEG[4] Tile_X6Y14_LUT4AB/N4BEG[5]
+ Tile_X6Y14_LUT4AB/N4BEG[6] Tile_X6Y14_LUT4AB/N4BEG[7] Tile_X6Y14_LUT4AB/N4BEG[8]
+ Tile_X6Y14_LUT4AB/N4BEG[9] Tile_X6Y13_LUT4AB/NN4BEG[0] Tile_X6Y13_LUT4AB/NN4BEG[10]
+ Tile_X6Y13_LUT4AB/NN4BEG[11] Tile_X6Y13_LUT4AB/NN4BEG[12] Tile_X6Y13_LUT4AB/NN4BEG[13]
+ Tile_X6Y13_LUT4AB/NN4BEG[14] Tile_X6Y13_LUT4AB/NN4BEG[15] Tile_X6Y13_LUT4AB/NN4BEG[1]
+ Tile_X6Y13_LUT4AB/NN4BEG[2] Tile_X6Y13_LUT4AB/NN4BEG[3] Tile_X6Y13_LUT4AB/NN4BEG[4]
+ Tile_X6Y13_LUT4AB/NN4BEG[5] Tile_X6Y13_LUT4AB/NN4BEG[6] Tile_X6Y13_LUT4AB/NN4BEG[7]
+ Tile_X6Y13_LUT4AB/NN4BEG[8] Tile_X6Y13_LUT4AB/NN4BEG[9] Tile_X6Y14_LUT4AB/NN4BEG[0]
+ Tile_X6Y14_LUT4AB/NN4BEG[10] Tile_X6Y14_LUT4AB/NN4BEG[11] Tile_X6Y14_LUT4AB/NN4BEG[12]
+ Tile_X6Y14_LUT4AB/NN4BEG[13] Tile_X6Y14_LUT4AB/NN4BEG[14] Tile_X6Y14_LUT4AB/NN4BEG[15]
+ Tile_X6Y14_LUT4AB/NN4BEG[1] Tile_X6Y14_LUT4AB/NN4BEG[2] Tile_X6Y14_LUT4AB/NN4BEG[3]
+ Tile_X6Y14_LUT4AB/NN4BEG[4] Tile_X6Y14_LUT4AB/NN4BEG[5] Tile_X6Y14_LUT4AB/NN4BEG[6]
+ Tile_X6Y14_LUT4AB/NN4BEG[7] Tile_X6Y14_LUT4AB/NN4BEG[8] Tile_X6Y14_LUT4AB/NN4BEG[9]
+ Tile_X6Y14_LUT4AB/S1END[0] Tile_X6Y14_LUT4AB/S1END[1] Tile_X6Y14_LUT4AB/S1END[2]
+ Tile_X6Y14_LUT4AB/S1END[3] Tile_X6Y13_LUT4AB/S1END[0] Tile_X6Y13_LUT4AB/S1END[1]
+ Tile_X6Y13_LUT4AB/S1END[2] Tile_X6Y13_LUT4AB/S1END[3] Tile_X6Y14_LUT4AB/S2MID[0]
+ Tile_X6Y14_LUT4AB/S2MID[1] Tile_X6Y14_LUT4AB/S2MID[2] Tile_X6Y14_LUT4AB/S2MID[3]
+ Tile_X6Y14_LUT4AB/S2MID[4] Tile_X6Y14_LUT4AB/S2MID[5] Tile_X6Y14_LUT4AB/S2MID[6]
+ Tile_X6Y14_LUT4AB/S2MID[7] Tile_X6Y14_LUT4AB/S2END[0] Tile_X6Y14_LUT4AB/S2END[1]
+ Tile_X6Y14_LUT4AB/S2END[2] Tile_X6Y14_LUT4AB/S2END[3] Tile_X6Y14_LUT4AB/S2END[4]
+ Tile_X6Y14_LUT4AB/S2END[5] Tile_X6Y14_LUT4AB/S2END[6] Tile_X6Y14_LUT4AB/S2END[7]
+ Tile_X6Y13_LUT4AB/S2END[0] Tile_X6Y13_LUT4AB/S2END[1] Tile_X6Y13_LUT4AB/S2END[2]
+ Tile_X6Y13_LUT4AB/S2END[3] Tile_X6Y13_LUT4AB/S2END[4] Tile_X6Y13_LUT4AB/S2END[5]
+ Tile_X6Y13_LUT4AB/S2END[6] Tile_X6Y13_LUT4AB/S2END[7] Tile_X6Y13_LUT4AB/S2MID[0]
+ Tile_X6Y13_LUT4AB/S2MID[1] Tile_X6Y13_LUT4AB/S2MID[2] Tile_X6Y13_LUT4AB/S2MID[3]
+ Tile_X6Y13_LUT4AB/S2MID[4] Tile_X6Y13_LUT4AB/S2MID[5] Tile_X6Y13_LUT4AB/S2MID[6]
+ Tile_X6Y13_LUT4AB/S2MID[7] Tile_X6Y14_LUT4AB/S4END[0] Tile_X6Y14_LUT4AB/S4END[10]
+ Tile_X6Y14_LUT4AB/S4END[11] Tile_X6Y14_LUT4AB/S4END[12] Tile_X6Y14_LUT4AB/S4END[13]
+ Tile_X6Y14_LUT4AB/S4END[14] Tile_X6Y14_LUT4AB/S4END[15] Tile_X6Y14_LUT4AB/S4END[1]
+ Tile_X6Y14_LUT4AB/S4END[2] Tile_X6Y14_LUT4AB/S4END[3] Tile_X6Y14_LUT4AB/S4END[4]
+ Tile_X6Y14_LUT4AB/S4END[5] Tile_X6Y14_LUT4AB/S4END[6] Tile_X6Y14_LUT4AB/S4END[7]
+ Tile_X6Y14_LUT4AB/S4END[8] Tile_X6Y14_LUT4AB/S4END[9] Tile_X6Y13_LUT4AB/S4END[0]
+ Tile_X6Y13_LUT4AB/S4END[10] Tile_X6Y13_LUT4AB/S4END[11] Tile_X6Y13_LUT4AB/S4END[12]
+ Tile_X6Y13_LUT4AB/S4END[13] Tile_X6Y13_LUT4AB/S4END[14] Tile_X6Y13_LUT4AB/S4END[15]
+ Tile_X6Y13_LUT4AB/S4END[1] Tile_X6Y13_LUT4AB/S4END[2] Tile_X6Y13_LUT4AB/S4END[3]
+ Tile_X6Y13_LUT4AB/S4END[4] Tile_X6Y13_LUT4AB/S4END[5] Tile_X6Y13_LUT4AB/S4END[6]
+ Tile_X6Y13_LUT4AB/S4END[7] Tile_X6Y13_LUT4AB/S4END[8] Tile_X6Y13_LUT4AB/S4END[9]
+ Tile_X6Y14_LUT4AB/SS4END[0] Tile_X6Y14_LUT4AB/SS4END[10] Tile_X6Y14_LUT4AB/SS4END[11]
+ Tile_X6Y14_LUT4AB/SS4END[12] Tile_X6Y14_LUT4AB/SS4END[13] Tile_X6Y14_LUT4AB/SS4END[14]
+ Tile_X6Y14_LUT4AB/SS4END[15] Tile_X6Y14_LUT4AB/SS4END[1] Tile_X6Y14_LUT4AB/SS4END[2]
+ Tile_X6Y14_LUT4AB/SS4END[3] Tile_X6Y14_LUT4AB/SS4END[4] Tile_X6Y14_LUT4AB/SS4END[5]
+ Tile_X6Y14_LUT4AB/SS4END[6] Tile_X6Y14_LUT4AB/SS4END[7] Tile_X6Y14_LUT4AB/SS4END[8]
+ Tile_X6Y14_LUT4AB/SS4END[9] Tile_X6Y13_LUT4AB/SS4END[0] Tile_X6Y13_LUT4AB/SS4END[10]
+ Tile_X6Y13_LUT4AB/SS4END[11] Tile_X6Y13_LUT4AB/SS4END[12] Tile_X6Y13_LUT4AB/SS4END[13]
+ Tile_X6Y13_LUT4AB/SS4END[14] Tile_X6Y13_LUT4AB/SS4END[15] Tile_X6Y13_LUT4AB/SS4END[1]
+ Tile_X6Y13_LUT4AB/SS4END[2] Tile_X6Y13_LUT4AB/SS4END[3] Tile_X6Y13_LUT4AB/SS4END[4]
+ Tile_X6Y13_LUT4AB/SS4END[5] Tile_X6Y13_LUT4AB/SS4END[6] Tile_X6Y13_LUT4AB/SS4END[7]
+ Tile_X6Y13_LUT4AB/SS4END[8] Tile_X6Y13_LUT4AB/SS4END[9] Tile_X6Y13_LUT4AB/UserCLK
+ Tile_X6Y12_LUT4AB/UserCLK VGND VPWR Tile_X6Y13_LUT4AB/W1BEG[0] Tile_X6Y13_LUT4AB/W1BEG[1]
+ Tile_X6Y13_LUT4AB/W1BEG[2] Tile_X6Y13_LUT4AB/W1BEG[3] Tile_X6Y13_LUT4AB/W1END[0]
+ Tile_X6Y13_LUT4AB/W1END[1] Tile_X6Y13_LUT4AB/W1END[2] Tile_X6Y13_LUT4AB/W1END[3]
+ Tile_X6Y13_LUT4AB/W2BEG[0] Tile_X6Y13_LUT4AB/W2BEG[1] Tile_X6Y13_LUT4AB/W2BEG[2]
+ Tile_X6Y13_LUT4AB/W2BEG[3] Tile_X6Y13_LUT4AB/W2BEG[4] Tile_X6Y13_LUT4AB/W2BEG[5]
+ Tile_X6Y13_LUT4AB/W2BEG[6] Tile_X6Y13_LUT4AB/W2BEG[7] Tile_X5Y13_LUT4AB/W2END[0]
+ Tile_X5Y13_LUT4AB/W2END[1] Tile_X5Y13_LUT4AB/W2END[2] Tile_X5Y13_LUT4AB/W2END[3]
+ Tile_X5Y13_LUT4AB/W2END[4] Tile_X5Y13_LUT4AB/W2END[5] Tile_X5Y13_LUT4AB/W2END[6]
+ Tile_X5Y13_LUT4AB/W2END[7] Tile_X6Y13_LUT4AB/W2END[0] Tile_X6Y13_LUT4AB/W2END[1]
+ Tile_X6Y13_LUT4AB/W2END[2] Tile_X6Y13_LUT4AB/W2END[3] Tile_X6Y13_LUT4AB/W2END[4]
+ Tile_X6Y13_LUT4AB/W2END[5] Tile_X6Y13_LUT4AB/W2END[6] Tile_X6Y13_LUT4AB/W2END[7]
+ Tile_X6Y13_LUT4AB/W2MID[0] Tile_X6Y13_LUT4AB/W2MID[1] Tile_X6Y13_LUT4AB/W2MID[2]
+ Tile_X6Y13_LUT4AB/W2MID[3] Tile_X6Y13_LUT4AB/W2MID[4] Tile_X6Y13_LUT4AB/W2MID[5]
+ Tile_X6Y13_LUT4AB/W2MID[6] Tile_X6Y13_LUT4AB/W2MID[7] Tile_X6Y13_LUT4AB/W6BEG[0]
+ Tile_X6Y13_LUT4AB/W6BEG[10] Tile_X6Y13_LUT4AB/W6BEG[11] Tile_X6Y13_LUT4AB/W6BEG[1]
+ Tile_X6Y13_LUT4AB/W6BEG[2] Tile_X6Y13_LUT4AB/W6BEG[3] Tile_X6Y13_LUT4AB/W6BEG[4]
+ Tile_X6Y13_LUT4AB/W6BEG[5] Tile_X6Y13_LUT4AB/W6BEG[6] Tile_X6Y13_LUT4AB/W6BEG[7]
+ Tile_X6Y13_LUT4AB/W6BEG[8] Tile_X6Y13_LUT4AB/W6BEG[9] Tile_X6Y13_LUT4AB/W6END[0]
+ Tile_X6Y13_LUT4AB/W6END[10] Tile_X6Y13_LUT4AB/W6END[11] Tile_X6Y13_LUT4AB/W6END[1]
+ Tile_X6Y13_LUT4AB/W6END[2] Tile_X6Y13_LUT4AB/W6END[3] Tile_X6Y13_LUT4AB/W6END[4]
+ Tile_X6Y13_LUT4AB/W6END[5] Tile_X6Y13_LUT4AB/W6END[6] Tile_X6Y13_LUT4AB/W6END[7]
+ Tile_X6Y13_LUT4AB/W6END[8] Tile_X6Y13_LUT4AB/W6END[9] Tile_X6Y13_LUT4AB/WW4BEG[0]
+ Tile_X6Y13_LUT4AB/WW4BEG[10] Tile_X6Y13_LUT4AB/WW4BEG[11] Tile_X6Y13_LUT4AB/WW4BEG[12]
+ Tile_X6Y13_LUT4AB/WW4BEG[13] Tile_X6Y13_LUT4AB/WW4BEG[14] Tile_X6Y13_LUT4AB/WW4BEG[15]
+ Tile_X6Y13_LUT4AB/WW4BEG[1] Tile_X6Y13_LUT4AB/WW4BEG[2] Tile_X6Y13_LUT4AB/WW4BEG[3]
+ Tile_X6Y13_LUT4AB/WW4BEG[4] Tile_X6Y13_LUT4AB/WW4BEG[5] Tile_X6Y13_LUT4AB/WW4BEG[6]
+ Tile_X6Y13_LUT4AB/WW4BEG[7] Tile_X6Y13_LUT4AB/WW4BEG[8] Tile_X6Y13_LUT4AB/WW4BEG[9]
+ Tile_X6Y13_LUT4AB/WW4END[0] Tile_X6Y13_LUT4AB/WW4END[10] Tile_X6Y13_LUT4AB/WW4END[11]
+ Tile_X6Y13_LUT4AB/WW4END[12] Tile_X6Y13_LUT4AB/WW4END[13] Tile_X6Y13_LUT4AB/WW4END[14]
+ Tile_X6Y13_LUT4AB/WW4END[15] Tile_X6Y13_LUT4AB/WW4END[1] Tile_X6Y13_LUT4AB/WW4END[2]
+ Tile_X6Y13_LUT4AB/WW4END[3] Tile_X6Y13_LUT4AB/WW4END[4] Tile_X6Y13_LUT4AB/WW4END[5]
+ Tile_X6Y13_LUT4AB/WW4END[6] Tile_X6Y13_LUT4AB/WW4END[7] Tile_X6Y13_LUT4AB/WW4END[8]
+ Tile_X6Y13_LUT4AB/WW4END[9] LUT4AB
XTile_X5Y0_N_term_single Tile_X5Y1_LUT4AB/Co Tile_X5Y0_N_term_single/FrameData[0]
+ Tile_X5Y0_N_term_single/FrameData[10] Tile_X5Y0_N_term_single/FrameData[11] Tile_X5Y0_N_term_single/FrameData[12]
+ Tile_X5Y0_N_term_single/FrameData[13] Tile_X5Y0_N_term_single/FrameData[14] Tile_X5Y0_N_term_single/FrameData[15]
+ Tile_X5Y0_N_term_single/FrameData[16] Tile_X5Y0_N_term_single/FrameData[17] Tile_X5Y0_N_term_single/FrameData[18]
+ Tile_X5Y0_N_term_single/FrameData[19] Tile_X5Y0_N_term_single/FrameData[1] Tile_X5Y0_N_term_single/FrameData[20]
+ Tile_X5Y0_N_term_single/FrameData[21] Tile_X5Y0_N_term_single/FrameData[22] Tile_X5Y0_N_term_single/FrameData[23]
+ Tile_X5Y0_N_term_single/FrameData[24] Tile_X5Y0_N_term_single/FrameData[25] Tile_X5Y0_N_term_single/FrameData[26]
+ Tile_X5Y0_N_term_single/FrameData[27] Tile_X5Y0_N_term_single/FrameData[28] Tile_X5Y0_N_term_single/FrameData[29]
+ Tile_X5Y0_N_term_single/FrameData[2] Tile_X5Y0_N_term_single/FrameData[30] Tile_X5Y0_N_term_single/FrameData[31]
+ Tile_X5Y0_N_term_single/FrameData[3] Tile_X5Y0_N_term_single/FrameData[4] Tile_X5Y0_N_term_single/FrameData[5]
+ Tile_X5Y0_N_term_single/FrameData[6] Tile_X5Y0_N_term_single/FrameData[7] Tile_X5Y0_N_term_single/FrameData[8]
+ Tile_X5Y0_N_term_single/FrameData[9] Tile_X6Y0_N_term_single/FrameData[0] Tile_X6Y0_N_term_single/FrameData[10]
+ Tile_X6Y0_N_term_single/FrameData[11] Tile_X6Y0_N_term_single/FrameData[12] Tile_X6Y0_N_term_single/FrameData[13]
+ Tile_X6Y0_N_term_single/FrameData[14] Tile_X6Y0_N_term_single/FrameData[15] Tile_X6Y0_N_term_single/FrameData[16]
+ Tile_X6Y0_N_term_single/FrameData[17] Tile_X6Y0_N_term_single/FrameData[18] Tile_X6Y0_N_term_single/FrameData[19]
+ Tile_X6Y0_N_term_single/FrameData[1] Tile_X6Y0_N_term_single/FrameData[20] Tile_X6Y0_N_term_single/FrameData[21]
+ Tile_X6Y0_N_term_single/FrameData[22] Tile_X6Y0_N_term_single/FrameData[23] Tile_X6Y0_N_term_single/FrameData[24]
+ Tile_X6Y0_N_term_single/FrameData[25] Tile_X6Y0_N_term_single/FrameData[26] Tile_X6Y0_N_term_single/FrameData[27]
+ Tile_X6Y0_N_term_single/FrameData[28] Tile_X6Y0_N_term_single/FrameData[29] Tile_X6Y0_N_term_single/FrameData[2]
+ Tile_X6Y0_N_term_single/FrameData[30] Tile_X6Y0_N_term_single/FrameData[31] Tile_X6Y0_N_term_single/FrameData[3]
+ Tile_X6Y0_N_term_single/FrameData[4] Tile_X6Y0_N_term_single/FrameData[5] Tile_X6Y0_N_term_single/FrameData[6]
+ Tile_X6Y0_N_term_single/FrameData[7] Tile_X6Y0_N_term_single/FrameData[8] Tile_X6Y0_N_term_single/FrameData[9]
+ Tile_X5Y1_LUT4AB/FrameStrobe_O[0] Tile_X5Y1_LUT4AB/FrameStrobe_O[10] Tile_X5Y1_LUT4AB/FrameStrobe_O[11]
+ Tile_X5Y1_LUT4AB/FrameStrobe_O[12] Tile_X5Y1_LUT4AB/FrameStrobe_O[13] Tile_X5Y1_LUT4AB/FrameStrobe_O[14]
+ Tile_X5Y1_LUT4AB/FrameStrobe_O[15] Tile_X5Y1_LUT4AB/FrameStrobe_O[16] Tile_X5Y1_LUT4AB/FrameStrobe_O[17]
+ Tile_X5Y1_LUT4AB/FrameStrobe_O[18] Tile_X5Y1_LUT4AB/FrameStrobe_O[19] Tile_X5Y1_LUT4AB/FrameStrobe_O[1]
+ Tile_X5Y1_LUT4AB/FrameStrobe_O[2] Tile_X5Y1_LUT4AB/FrameStrobe_O[3] Tile_X5Y1_LUT4AB/FrameStrobe_O[4]
+ Tile_X5Y1_LUT4AB/FrameStrobe_O[5] Tile_X5Y1_LUT4AB/FrameStrobe_O[6] Tile_X5Y1_LUT4AB/FrameStrobe_O[7]
+ Tile_X5Y1_LUT4AB/FrameStrobe_O[8] Tile_X5Y1_LUT4AB/FrameStrobe_O[9] Tile_X5Y0_N_term_single/FrameStrobe_O[0]
+ Tile_X5Y0_N_term_single/FrameStrobe_O[10] Tile_X5Y0_N_term_single/FrameStrobe_O[11]
+ Tile_X5Y0_N_term_single/FrameStrobe_O[12] Tile_X5Y0_N_term_single/FrameStrobe_O[13]
+ Tile_X5Y0_N_term_single/FrameStrobe_O[14] Tile_X5Y0_N_term_single/FrameStrobe_O[15]
+ Tile_X5Y0_N_term_single/FrameStrobe_O[16] Tile_X5Y0_N_term_single/FrameStrobe_O[17]
+ Tile_X5Y0_N_term_single/FrameStrobe_O[18] Tile_X5Y0_N_term_single/FrameStrobe_O[19]
+ Tile_X5Y0_N_term_single/FrameStrobe_O[1] Tile_X5Y0_N_term_single/FrameStrobe_O[2]
+ Tile_X5Y0_N_term_single/FrameStrobe_O[3] Tile_X5Y0_N_term_single/FrameStrobe_O[4]
+ Tile_X5Y0_N_term_single/FrameStrobe_O[5] Tile_X5Y0_N_term_single/FrameStrobe_O[6]
+ Tile_X5Y0_N_term_single/FrameStrobe_O[7] Tile_X5Y0_N_term_single/FrameStrobe_O[8]
+ Tile_X5Y0_N_term_single/FrameStrobe_O[9] Tile_X5Y1_LUT4AB/N1BEG[0] Tile_X5Y1_LUT4AB/N1BEG[1]
+ Tile_X5Y1_LUT4AB/N1BEG[2] Tile_X5Y1_LUT4AB/N1BEG[3] Tile_X5Y1_LUT4AB/N2BEGb[0] Tile_X5Y1_LUT4AB/N2BEGb[1]
+ Tile_X5Y1_LUT4AB/N2BEGb[2] Tile_X5Y1_LUT4AB/N2BEGb[3] Tile_X5Y1_LUT4AB/N2BEGb[4]
+ Tile_X5Y1_LUT4AB/N2BEGb[5] Tile_X5Y1_LUT4AB/N2BEGb[6] Tile_X5Y1_LUT4AB/N2BEGb[7]
+ Tile_X5Y1_LUT4AB/N2BEG[0] Tile_X5Y1_LUT4AB/N2BEG[1] Tile_X5Y1_LUT4AB/N2BEG[2] Tile_X5Y1_LUT4AB/N2BEG[3]
+ Tile_X5Y1_LUT4AB/N2BEG[4] Tile_X5Y1_LUT4AB/N2BEG[5] Tile_X5Y1_LUT4AB/N2BEG[6] Tile_X5Y1_LUT4AB/N2BEG[7]
+ Tile_X5Y1_LUT4AB/N4BEG[0] Tile_X5Y1_LUT4AB/N4BEG[10] Tile_X5Y1_LUT4AB/N4BEG[11]
+ Tile_X5Y1_LUT4AB/N4BEG[12] Tile_X5Y1_LUT4AB/N4BEG[13] Tile_X5Y1_LUT4AB/N4BEG[14]
+ Tile_X5Y1_LUT4AB/N4BEG[15] Tile_X5Y1_LUT4AB/N4BEG[1] Tile_X5Y1_LUT4AB/N4BEG[2] Tile_X5Y1_LUT4AB/N4BEG[3]
+ Tile_X5Y1_LUT4AB/N4BEG[4] Tile_X5Y1_LUT4AB/N4BEG[5] Tile_X5Y1_LUT4AB/N4BEG[6] Tile_X5Y1_LUT4AB/N4BEG[7]
+ Tile_X5Y1_LUT4AB/N4BEG[8] Tile_X5Y1_LUT4AB/N4BEG[9] Tile_X5Y1_LUT4AB/NN4BEG[0] Tile_X5Y1_LUT4AB/NN4BEG[10]
+ Tile_X5Y1_LUT4AB/NN4BEG[11] Tile_X5Y1_LUT4AB/NN4BEG[12] Tile_X5Y1_LUT4AB/NN4BEG[13]
+ Tile_X5Y1_LUT4AB/NN4BEG[14] Tile_X5Y1_LUT4AB/NN4BEG[15] Tile_X5Y1_LUT4AB/NN4BEG[1]
+ Tile_X5Y1_LUT4AB/NN4BEG[2] Tile_X5Y1_LUT4AB/NN4BEG[3] Tile_X5Y1_LUT4AB/NN4BEG[4]
+ Tile_X5Y1_LUT4AB/NN4BEG[5] Tile_X5Y1_LUT4AB/NN4BEG[6] Tile_X5Y1_LUT4AB/NN4BEG[7]
+ Tile_X5Y1_LUT4AB/NN4BEG[8] Tile_X5Y1_LUT4AB/NN4BEG[9] Tile_X5Y1_LUT4AB/S1END[0]
+ Tile_X5Y1_LUT4AB/S1END[1] Tile_X5Y1_LUT4AB/S1END[2] Tile_X5Y1_LUT4AB/S1END[3] Tile_X5Y1_LUT4AB/S2MID[0]
+ Tile_X5Y1_LUT4AB/S2MID[1] Tile_X5Y1_LUT4AB/S2MID[2] Tile_X5Y1_LUT4AB/S2MID[3] Tile_X5Y1_LUT4AB/S2MID[4]
+ Tile_X5Y1_LUT4AB/S2MID[5] Tile_X5Y1_LUT4AB/S2MID[6] Tile_X5Y1_LUT4AB/S2MID[7] Tile_X5Y1_LUT4AB/S2END[0]
+ Tile_X5Y1_LUT4AB/S2END[1] Tile_X5Y1_LUT4AB/S2END[2] Tile_X5Y1_LUT4AB/S2END[3] Tile_X5Y1_LUT4AB/S2END[4]
+ Tile_X5Y1_LUT4AB/S2END[5] Tile_X5Y1_LUT4AB/S2END[6] Tile_X5Y1_LUT4AB/S2END[7] Tile_X5Y1_LUT4AB/S4END[0]
+ Tile_X5Y1_LUT4AB/S4END[10] Tile_X5Y1_LUT4AB/S4END[11] Tile_X5Y1_LUT4AB/S4END[12]
+ Tile_X5Y1_LUT4AB/S4END[13] Tile_X5Y1_LUT4AB/S4END[14] Tile_X5Y1_LUT4AB/S4END[15]
+ Tile_X5Y1_LUT4AB/S4END[1] Tile_X5Y1_LUT4AB/S4END[2] Tile_X5Y1_LUT4AB/S4END[3] Tile_X5Y1_LUT4AB/S4END[4]
+ Tile_X5Y1_LUT4AB/S4END[5] Tile_X5Y1_LUT4AB/S4END[6] Tile_X5Y1_LUT4AB/S4END[7] Tile_X5Y1_LUT4AB/S4END[8]
+ Tile_X5Y1_LUT4AB/S4END[9] Tile_X5Y1_LUT4AB/SS4END[0] Tile_X5Y1_LUT4AB/SS4END[10]
+ Tile_X5Y1_LUT4AB/SS4END[11] Tile_X5Y1_LUT4AB/SS4END[12] Tile_X5Y1_LUT4AB/SS4END[13]
+ Tile_X5Y1_LUT4AB/SS4END[14] Tile_X5Y1_LUT4AB/SS4END[15] Tile_X5Y1_LUT4AB/SS4END[1]
+ Tile_X5Y1_LUT4AB/SS4END[2] Tile_X5Y1_LUT4AB/SS4END[3] Tile_X5Y1_LUT4AB/SS4END[4]
+ Tile_X5Y1_LUT4AB/SS4END[5] Tile_X5Y1_LUT4AB/SS4END[6] Tile_X5Y1_LUT4AB/SS4END[7]
+ Tile_X5Y1_LUT4AB/SS4END[8] Tile_X5Y1_LUT4AB/SS4END[9] Tile_X5Y1_LUT4AB/UserCLKo
+ Tile_X5Y0_N_term_single/UserCLKo VGND VPWR N_term_single
XTile_X6Y15_S_CPU_IF Tile_X6Y14_LUT4AB/Ci Tile_X6Y15_S_CPU_IF/FrameData[0] Tile_X6Y15_S_CPU_IF/FrameData[10]
+ Tile_X6Y15_S_CPU_IF/FrameData[11] Tile_X6Y15_S_CPU_IF/FrameData[12] Tile_X6Y15_S_CPU_IF/FrameData[13]
+ Tile_X6Y15_S_CPU_IF/FrameData[14] Tile_X6Y15_S_CPU_IF/FrameData[15] Tile_X6Y15_S_CPU_IF/FrameData[16]
+ Tile_X6Y15_S_CPU_IF/FrameData[17] Tile_X6Y15_S_CPU_IF/FrameData[18] Tile_X6Y15_S_CPU_IF/FrameData[19]
+ Tile_X6Y15_S_CPU_IF/FrameData[1] Tile_X6Y15_S_CPU_IF/FrameData[20] Tile_X6Y15_S_CPU_IF/FrameData[21]
+ Tile_X6Y15_S_CPU_IF/FrameData[22] Tile_X6Y15_S_CPU_IF/FrameData[23] Tile_X6Y15_S_CPU_IF/FrameData[24]
+ Tile_X6Y15_S_CPU_IF/FrameData[25] Tile_X6Y15_S_CPU_IF/FrameData[26] Tile_X6Y15_S_CPU_IF/FrameData[27]
+ Tile_X6Y15_S_CPU_IF/FrameData[28] Tile_X6Y15_S_CPU_IF/FrameData[29] Tile_X6Y15_S_CPU_IF/FrameData[2]
+ Tile_X6Y15_S_CPU_IF/FrameData[30] Tile_X6Y15_S_CPU_IF/FrameData[31] Tile_X6Y15_S_CPU_IF/FrameData[3]
+ Tile_X6Y15_S_CPU_IF/FrameData[4] Tile_X6Y15_S_CPU_IF/FrameData[5] Tile_X6Y15_S_CPU_IF/FrameData[6]
+ Tile_X6Y15_S_CPU_IF/FrameData[7] Tile_X6Y15_S_CPU_IF/FrameData[8] Tile_X6Y15_S_CPU_IF/FrameData[9]
+ Tile_X7Y15_S_term_DSP/FrameData[0] Tile_X7Y15_S_term_DSP/FrameData[10] Tile_X7Y15_S_term_DSP/FrameData[11]
+ Tile_X7Y15_S_term_DSP/FrameData[12] Tile_X7Y15_S_term_DSP/FrameData[13] Tile_X7Y15_S_term_DSP/FrameData[14]
+ Tile_X7Y15_S_term_DSP/FrameData[15] Tile_X7Y15_S_term_DSP/FrameData[16] Tile_X7Y15_S_term_DSP/FrameData[17]
+ Tile_X7Y15_S_term_DSP/FrameData[18] Tile_X7Y15_S_term_DSP/FrameData[19] Tile_X7Y15_S_term_DSP/FrameData[1]
+ Tile_X7Y15_S_term_DSP/FrameData[20] Tile_X7Y15_S_term_DSP/FrameData[21] Tile_X7Y15_S_term_DSP/FrameData[22]
+ Tile_X7Y15_S_term_DSP/FrameData[23] Tile_X7Y15_S_term_DSP/FrameData[24] Tile_X7Y15_S_term_DSP/FrameData[25]
+ Tile_X7Y15_S_term_DSP/FrameData[26] Tile_X7Y15_S_term_DSP/FrameData[27] Tile_X7Y15_S_term_DSP/FrameData[28]
+ Tile_X7Y15_S_term_DSP/FrameData[29] Tile_X7Y15_S_term_DSP/FrameData[2] Tile_X7Y15_S_term_DSP/FrameData[30]
+ Tile_X7Y15_S_term_DSP/FrameData[31] Tile_X7Y15_S_term_DSP/FrameData[3] Tile_X7Y15_S_term_DSP/FrameData[4]
+ Tile_X7Y15_S_term_DSP/FrameData[5] Tile_X7Y15_S_term_DSP/FrameData[6] Tile_X7Y15_S_term_DSP/FrameData[7]
+ Tile_X7Y15_S_term_DSP/FrameData[8] Tile_X7Y15_S_term_DSP/FrameData[9] FrameStrobe[120]
+ FrameStrobe[130] FrameStrobe[131] FrameStrobe[132] FrameStrobe[133] FrameStrobe[134]
+ FrameStrobe[135] FrameStrobe[136] FrameStrobe[137] FrameStrobe[138] FrameStrobe[139]
+ FrameStrobe[121] FrameStrobe[122] FrameStrobe[123] FrameStrobe[124] FrameStrobe[125]
+ FrameStrobe[126] FrameStrobe[127] FrameStrobe[128] FrameStrobe[129] Tile_X6Y14_LUT4AB/FrameStrobe[0]
+ Tile_X6Y14_LUT4AB/FrameStrobe[10] Tile_X6Y14_LUT4AB/FrameStrobe[11] Tile_X6Y14_LUT4AB/FrameStrobe[12]
+ Tile_X6Y14_LUT4AB/FrameStrobe[13] Tile_X6Y14_LUT4AB/FrameStrobe[14] Tile_X6Y14_LUT4AB/FrameStrobe[15]
+ Tile_X6Y14_LUT4AB/FrameStrobe[16] Tile_X6Y14_LUT4AB/FrameStrobe[17] Tile_X6Y14_LUT4AB/FrameStrobe[18]
+ Tile_X6Y14_LUT4AB/FrameStrobe[19] Tile_X6Y14_LUT4AB/FrameStrobe[1] Tile_X6Y14_LUT4AB/FrameStrobe[2]
+ Tile_X6Y14_LUT4AB/FrameStrobe[3] Tile_X6Y14_LUT4AB/FrameStrobe[4] Tile_X6Y14_LUT4AB/FrameStrobe[5]
+ Tile_X6Y14_LUT4AB/FrameStrobe[6] Tile_X6Y14_LUT4AB/FrameStrobe[7] Tile_X6Y14_LUT4AB/FrameStrobe[8]
+ Tile_X6Y14_LUT4AB/FrameStrobe[9] Tile_X6Y15_I_top0 Tile_X6Y15_I_top1 Tile_X6Y15_I_top10
+ Tile_X6Y15_I_top11 Tile_X6Y15_I_top12 Tile_X6Y15_I_top13 Tile_X6Y15_I_top14 Tile_X6Y15_I_top15
+ Tile_X6Y15_I_top2 Tile_X6Y15_I_top3 Tile_X6Y15_I_top4 Tile_X6Y15_I_top5 Tile_X6Y15_I_top6
+ Tile_X6Y15_I_top7 Tile_X6Y15_I_top8 Tile_X6Y15_I_top9 Tile_X6Y14_LUT4AB/N1END[0]
+ Tile_X6Y14_LUT4AB/N1END[1] Tile_X6Y14_LUT4AB/N1END[2] Tile_X6Y14_LUT4AB/N1END[3]
+ Tile_X6Y14_LUT4AB/N2MID[0] Tile_X6Y14_LUT4AB/N2MID[1] Tile_X6Y14_LUT4AB/N2MID[2]
+ Tile_X6Y14_LUT4AB/N2MID[3] Tile_X6Y14_LUT4AB/N2MID[4] Tile_X6Y14_LUT4AB/N2MID[5]
+ Tile_X6Y14_LUT4AB/N2MID[6] Tile_X6Y14_LUT4AB/N2MID[7] Tile_X6Y14_LUT4AB/N2END[0]
+ Tile_X6Y14_LUT4AB/N2END[1] Tile_X6Y14_LUT4AB/N2END[2] Tile_X6Y14_LUT4AB/N2END[3]
+ Tile_X6Y14_LUT4AB/N2END[4] Tile_X6Y14_LUT4AB/N2END[5] Tile_X6Y14_LUT4AB/N2END[6]
+ Tile_X6Y14_LUT4AB/N2END[7] Tile_X6Y14_LUT4AB/N4END[0] Tile_X6Y14_LUT4AB/N4END[10]
+ Tile_X6Y14_LUT4AB/N4END[11] Tile_X6Y14_LUT4AB/N4END[12] Tile_X6Y14_LUT4AB/N4END[13]
+ Tile_X6Y14_LUT4AB/N4END[14] Tile_X6Y14_LUT4AB/N4END[15] Tile_X6Y14_LUT4AB/N4END[1]
+ Tile_X6Y14_LUT4AB/N4END[2] Tile_X6Y14_LUT4AB/N4END[3] Tile_X6Y14_LUT4AB/N4END[4]
+ Tile_X6Y14_LUT4AB/N4END[5] Tile_X6Y14_LUT4AB/N4END[6] Tile_X6Y14_LUT4AB/N4END[7]
+ Tile_X6Y14_LUT4AB/N4END[8] Tile_X6Y14_LUT4AB/N4END[9] Tile_X6Y14_LUT4AB/NN4END[0]
+ Tile_X6Y14_LUT4AB/NN4END[10] Tile_X6Y14_LUT4AB/NN4END[11] Tile_X6Y14_LUT4AB/NN4END[12]
+ Tile_X6Y14_LUT4AB/NN4END[13] Tile_X6Y14_LUT4AB/NN4END[14] Tile_X6Y14_LUT4AB/NN4END[15]
+ Tile_X6Y14_LUT4AB/NN4END[1] Tile_X6Y14_LUT4AB/NN4END[2] Tile_X6Y14_LUT4AB/NN4END[3]
+ Tile_X6Y14_LUT4AB/NN4END[4] Tile_X6Y14_LUT4AB/NN4END[5] Tile_X6Y14_LUT4AB/NN4END[6]
+ Tile_X6Y14_LUT4AB/NN4END[7] Tile_X6Y14_LUT4AB/NN4END[8] Tile_X6Y14_LUT4AB/NN4END[9]
+ Tile_X6Y15_O_top0 Tile_X6Y15_O_top1 Tile_X6Y15_O_top10 Tile_X6Y15_O_top11 Tile_X6Y15_O_top12
+ Tile_X6Y15_O_top13 Tile_X6Y15_O_top14 Tile_X6Y15_O_top15 Tile_X6Y15_O_top2 Tile_X6Y15_O_top3
+ Tile_X6Y15_O_top4 Tile_X6Y15_O_top5 Tile_X6Y15_O_top6 Tile_X6Y15_O_top7 Tile_X6Y15_O_top8
+ Tile_X6Y15_O_top9 Tile_X6Y14_LUT4AB/S1BEG[0] Tile_X6Y14_LUT4AB/S1BEG[1] Tile_X6Y14_LUT4AB/S1BEG[2]
+ Tile_X6Y14_LUT4AB/S1BEG[3] Tile_X6Y14_LUT4AB/S2BEGb[0] Tile_X6Y14_LUT4AB/S2BEGb[1]
+ Tile_X6Y14_LUT4AB/S2BEGb[2] Tile_X6Y14_LUT4AB/S2BEGb[3] Tile_X6Y14_LUT4AB/S2BEGb[4]
+ Tile_X6Y14_LUT4AB/S2BEGb[5] Tile_X6Y14_LUT4AB/S2BEGb[6] Tile_X6Y14_LUT4AB/S2BEGb[7]
+ Tile_X6Y14_LUT4AB/S2BEG[0] Tile_X6Y14_LUT4AB/S2BEG[1] Tile_X6Y14_LUT4AB/S2BEG[2]
+ Tile_X6Y14_LUT4AB/S2BEG[3] Tile_X6Y14_LUT4AB/S2BEG[4] Tile_X6Y14_LUT4AB/S2BEG[5]
+ Tile_X6Y14_LUT4AB/S2BEG[6] Tile_X6Y14_LUT4AB/S2BEG[7] Tile_X6Y14_LUT4AB/S4BEG[0]
+ Tile_X6Y14_LUT4AB/S4BEG[10] Tile_X6Y14_LUT4AB/S4BEG[11] Tile_X6Y14_LUT4AB/S4BEG[12]
+ Tile_X6Y14_LUT4AB/S4BEG[13] Tile_X6Y14_LUT4AB/S4BEG[14] Tile_X6Y14_LUT4AB/S4BEG[15]
+ Tile_X6Y14_LUT4AB/S4BEG[1] Tile_X6Y14_LUT4AB/S4BEG[2] Tile_X6Y14_LUT4AB/S4BEG[3]
+ Tile_X6Y14_LUT4AB/S4BEG[4] Tile_X6Y14_LUT4AB/S4BEG[5] Tile_X6Y14_LUT4AB/S4BEG[6]
+ Tile_X6Y14_LUT4AB/S4BEG[7] Tile_X6Y14_LUT4AB/S4BEG[8] Tile_X6Y14_LUT4AB/S4BEG[9]
+ Tile_X6Y14_LUT4AB/SS4BEG[0] Tile_X6Y14_LUT4AB/SS4BEG[10] Tile_X6Y14_LUT4AB/SS4BEG[11]
+ Tile_X6Y14_LUT4AB/SS4BEG[12] Tile_X6Y14_LUT4AB/SS4BEG[13] Tile_X6Y14_LUT4AB/SS4BEG[14]
+ Tile_X6Y14_LUT4AB/SS4BEG[15] Tile_X6Y14_LUT4AB/SS4BEG[1] Tile_X6Y14_LUT4AB/SS4BEG[2]
+ Tile_X6Y14_LUT4AB/SS4BEG[3] Tile_X6Y14_LUT4AB/SS4BEG[4] Tile_X6Y14_LUT4AB/SS4BEG[5]
+ Tile_X6Y14_LUT4AB/SS4BEG[6] Tile_X6Y14_LUT4AB/SS4BEG[7] Tile_X6Y14_LUT4AB/SS4BEG[8]
+ Tile_X6Y14_LUT4AB/SS4BEG[9] UserCLK Tile_X6Y14_LUT4AB/UserCLK VGND VPWR S_CPU_IF
XTile_X4Y13_RegFile Tile_X5Y13_LUT4AB/E1END[0] Tile_X5Y13_LUT4AB/E1END[1] Tile_X5Y13_LUT4AB/E1END[2]
+ Tile_X5Y13_LUT4AB/E1END[3] Tile_X3Y13_LUT4AB/E1BEG[0] Tile_X3Y13_LUT4AB/E1BEG[1]
+ Tile_X3Y13_LUT4AB/E1BEG[2] Tile_X3Y13_LUT4AB/E1BEG[3] Tile_X5Y13_LUT4AB/E2MID[0]
+ Tile_X5Y13_LUT4AB/E2MID[1] Tile_X5Y13_LUT4AB/E2MID[2] Tile_X5Y13_LUT4AB/E2MID[3]
+ Tile_X5Y13_LUT4AB/E2MID[4] Tile_X5Y13_LUT4AB/E2MID[5] Tile_X5Y13_LUT4AB/E2MID[6]
+ Tile_X5Y13_LUT4AB/E2MID[7] Tile_X5Y13_LUT4AB/E2END[0] Tile_X5Y13_LUT4AB/E2END[1]
+ Tile_X5Y13_LUT4AB/E2END[2] Tile_X5Y13_LUT4AB/E2END[3] Tile_X5Y13_LUT4AB/E2END[4]
+ Tile_X5Y13_LUT4AB/E2END[5] Tile_X5Y13_LUT4AB/E2END[6] Tile_X5Y13_LUT4AB/E2END[7]
+ Tile_X4Y13_RegFile/E2END[0] Tile_X4Y13_RegFile/E2END[1] Tile_X4Y13_RegFile/E2END[2]
+ Tile_X4Y13_RegFile/E2END[3] Tile_X4Y13_RegFile/E2END[4] Tile_X4Y13_RegFile/E2END[5]
+ Tile_X4Y13_RegFile/E2END[6] Tile_X4Y13_RegFile/E2END[7] Tile_X3Y13_LUT4AB/E2BEG[0]
+ Tile_X3Y13_LUT4AB/E2BEG[1] Tile_X3Y13_LUT4AB/E2BEG[2] Tile_X3Y13_LUT4AB/E2BEG[3]
+ Tile_X3Y13_LUT4AB/E2BEG[4] Tile_X3Y13_LUT4AB/E2BEG[5] Tile_X3Y13_LUT4AB/E2BEG[6]
+ Tile_X3Y13_LUT4AB/E2BEG[7] Tile_X5Y13_LUT4AB/E6END[0] Tile_X5Y13_LUT4AB/E6END[10]
+ Tile_X5Y13_LUT4AB/E6END[11] Tile_X5Y13_LUT4AB/E6END[1] Tile_X5Y13_LUT4AB/E6END[2]
+ Tile_X5Y13_LUT4AB/E6END[3] Tile_X5Y13_LUT4AB/E6END[4] Tile_X5Y13_LUT4AB/E6END[5]
+ Tile_X5Y13_LUT4AB/E6END[6] Tile_X5Y13_LUT4AB/E6END[7] Tile_X5Y13_LUT4AB/E6END[8]
+ Tile_X5Y13_LUT4AB/E6END[9] Tile_X3Y13_LUT4AB/E6BEG[0] Tile_X3Y13_LUT4AB/E6BEG[10]
+ Tile_X3Y13_LUT4AB/E6BEG[11] Tile_X3Y13_LUT4AB/E6BEG[1] Tile_X3Y13_LUT4AB/E6BEG[2]
+ Tile_X3Y13_LUT4AB/E6BEG[3] Tile_X3Y13_LUT4AB/E6BEG[4] Tile_X3Y13_LUT4AB/E6BEG[5]
+ Tile_X3Y13_LUT4AB/E6BEG[6] Tile_X3Y13_LUT4AB/E6BEG[7] Tile_X3Y13_LUT4AB/E6BEG[8]
+ Tile_X3Y13_LUT4AB/E6BEG[9] Tile_X5Y13_LUT4AB/EE4END[0] Tile_X5Y13_LUT4AB/EE4END[10]
+ Tile_X5Y13_LUT4AB/EE4END[11] Tile_X5Y13_LUT4AB/EE4END[12] Tile_X5Y13_LUT4AB/EE4END[13]
+ Tile_X5Y13_LUT4AB/EE4END[14] Tile_X5Y13_LUT4AB/EE4END[15] Tile_X5Y13_LUT4AB/EE4END[1]
+ Tile_X5Y13_LUT4AB/EE4END[2] Tile_X5Y13_LUT4AB/EE4END[3] Tile_X5Y13_LUT4AB/EE4END[4]
+ Tile_X5Y13_LUT4AB/EE4END[5] Tile_X5Y13_LUT4AB/EE4END[6] Tile_X5Y13_LUT4AB/EE4END[7]
+ Tile_X5Y13_LUT4AB/EE4END[8] Tile_X5Y13_LUT4AB/EE4END[9] Tile_X3Y13_LUT4AB/EE4BEG[0]
+ Tile_X3Y13_LUT4AB/EE4BEG[10] Tile_X3Y13_LUT4AB/EE4BEG[11] Tile_X3Y13_LUT4AB/EE4BEG[12]
+ Tile_X3Y13_LUT4AB/EE4BEG[13] Tile_X3Y13_LUT4AB/EE4BEG[14] Tile_X3Y13_LUT4AB/EE4BEG[15]
+ Tile_X3Y13_LUT4AB/EE4BEG[1] Tile_X3Y13_LUT4AB/EE4BEG[2] Tile_X3Y13_LUT4AB/EE4BEG[3]
+ Tile_X3Y13_LUT4AB/EE4BEG[4] Tile_X3Y13_LUT4AB/EE4BEG[5] Tile_X3Y13_LUT4AB/EE4BEG[6]
+ Tile_X3Y13_LUT4AB/EE4BEG[7] Tile_X3Y13_LUT4AB/EE4BEG[8] Tile_X3Y13_LUT4AB/EE4BEG[9]
+ Tile_X4Y13_RegFile/FrameData[0] Tile_X4Y13_RegFile/FrameData[10] Tile_X4Y13_RegFile/FrameData[11]
+ Tile_X4Y13_RegFile/FrameData[12] Tile_X4Y13_RegFile/FrameData[13] Tile_X4Y13_RegFile/FrameData[14]
+ Tile_X4Y13_RegFile/FrameData[15] Tile_X4Y13_RegFile/FrameData[16] Tile_X4Y13_RegFile/FrameData[17]
+ Tile_X4Y13_RegFile/FrameData[18] Tile_X4Y13_RegFile/FrameData[19] Tile_X4Y13_RegFile/FrameData[1]
+ Tile_X4Y13_RegFile/FrameData[20] Tile_X4Y13_RegFile/FrameData[21] Tile_X4Y13_RegFile/FrameData[22]
+ Tile_X4Y13_RegFile/FrameData[23] Tile_X4Y13_RegFile/FrameData[24] Tile_X4Y13_RegFile/FrameData[25]
+ Tile_X4Y13_RegFile/FrameData[26] Tile_X4Y13_RegFile/FrameData[27] Tile_X4Y13_RegFile/FrameData[28]
+ Tile_X4Y13_RegFile/FrameData[29] Tile_X4Y13_RegFile/FrameData[2] Tile_X4Y13_RegFile/FrameData[30]
+ Tile_X4Y13_RegFile/FrameData[31] Tile_X4Y13_RegFile/FrameData[3] Tile_X4Y13_RegFile/FrameData[4]
+ Tile_X4Y13_RegFile/FrameData[5] Tile_X4Y13_RegFile/FrameData[6] Tile_X4Y13_RegFile/FrameData[7]
+ Tile_X4Y13_RegFile/FrameData[8] Tile_X4Y13_RegFile/FrameData[9] Tile_X5Y13_LUT4AB/FrameData[0]
+ Tile_X5Y13_LUT4AB/FrameData[10] Tile_X5Y13_LUT4AB/FrameData[11] Tile_X5Y13_LUT4AB/FrameData[12]
+ Tile_X5Y13_LUT4AB/FrameData[13] Tile_X5Y13_LUT4AB/FrameData[14] Tile_X5Y13_LUT4AB/FrameData[15]
+ Tile_X5Y13_LUT4AB/FrameData[16] Tile_X5Y13_LUT4AB/FrameData[17] Tile_X5Y13_LUT4AB/FrameData[18]
+ Tile_X5Y13_LUT4AB/FrameData[19] Tile_X5Y13_LUT4AB/FrameData[1] Tile_X5Y13_LUT4AB/FrameData[20]
+ Tile_X5Y13_LUT4AB/FrameData[21] Tile_X5Y13_LUT4AB/FrameData[22] Tile_X5Y13_LUT4AB/FrameData[23]
+ Tile_X5Y13_LUT4AB/FrameData[24] Tile_X5Y13_LUT4AB/FrameData[25] Tile_X5Y13_LUT4AB/FrameData[26]
+ Tile_X5Y13_LUT4AB/FrameData[27] Tile_X5Y13_LUT4AB/FrameData[28] Tile_X5Y13_LUT4AB/FrameData[29]
+ Tile_X5Y13_LUT4AB/FrameData[2] Tile_X5Y13_LUT4AB/FrameData[30] Tile_X5Y13_LUT4AB/FrameData[31]
+ Tile_X5Y13_LUT4AB/FrameData[3] Tile_X5Y13_LUT4AB/FrameData[4] Tile_X5Y13_LUT4AB/FrameData[5]
+ Tile_X5Y13_LUT4AB/FrameData[6] Tile_X5Y13_LUT4AB/FrameData[7] Tile_X5Y13_LUT4AB/FrameData[8]
+ Tile_X5Y13_LUT4AB/FrameData[9] Tile_X4Y13_RegFile/FrameStrobe[0] Tile_X4Y13_RegFile/FrameStrobe[10]
+ Tile_X4Y13_RegFile/FrameStrobe[11] Tile_X4Y13_RegFile/FrameStrobe[12] Tile_X4Y13_RegFile/FrameStrobe[13]
+ Tile_X4Y13_RegFile/FrameStrobe[14] Tile_X4Y13_RegFile/FrameStrobe[15] Tile_X4Y13_RegFile/FrameStrobe[16]
+ Tile_X4Y13_RegFile/FrameStrobe[17] Tile_X4Y13_RegFile/FrameStrobe[18] Tile_X4Y13_RegFile/FrameStrobe[19]
+ Tile_X4Y13_RegFile/FrameStrobe[1] Tile_X4Y13_RegFile/FrameStrobe[2] Tile_X4Y13_RegFile/FrameStrobe[3]
+ Tile_X4Y13_RegFile/FrameStrobe[4] Tile_X4Y13_RegFile/FrameStrobe[5] Tile_X4Y13_RegFile/FrameStrobe[6]
+ Tile_X4Y13_RegFile/FrameStrobe[7] Tile_X4Y13_RegFile/FrameStrobe[8] Tile_X4Y13_RegFile/FrameStrobe[9]
+ Tile_X4Y12_RegFile/FrameStrobe[0] Tile_X4Y12_RegFile/FrameStrobe[10] Tile_X4Y12_RegFile/FrameStrobe[11]
+ Tile_X4Y12_RegFile/FrameStrobe[12] Tile_X4Y12_RegFile/FrameStrobe[13] Tile_X4Y12_RegFile/FrameStrobe[14]
+ Tile_X4Y12_RegFile/FrameStrobe[15] Tile_X4Y12_RegFile/FrameStrobe[16] Tile_X4Y12_RegFile/FrameStrobe[17]
+ Tile_X4Y12_RegFile/FrameStrobe[18] Tile_X4Y12_RegFile/FrameStrobe[19] Tile_X4Y12_RegFile/FrameStrobe[1]
+ Tile_X4Y12_RegFile/FrameStrobe[2] Tile_X4Y12_RegFile/FrameStrobe[3] Tile_X4Y12_RegFile/FrameStrobe[4]
+ Tile_X4Y12_RegFile/FrameStrobe[5] Tile_X4Y12_RegFile/FrameStrobe[6] Tile_X4Y12_RegFile/FrameStrobe[7]
+ Tile_X4Y12_RegFile/FrameStrobe[8] Tile_X4Y12_RegFile/FrameStrobe[9] Tile_X4Y13_RegFile/N1BEG[0]
+ Tile_X4Y13_RegFile/N1BEG[1] Tile_X4Y13_RegFile/N1BEG[2] Tile_X4Y13_RegFile/N1BEG[3]
+ Tile_X4Y14_RegFile/N1BEG[0] Tile_X4Y14_RegFile/N1BEG[1] Tile_X4Y14_RegFile/N1BEG[2]
+ Tile_X4Y14_RegFile/N1BEG[3] Tile_X4Y13_RegFile/N2BEG[0] Tile_X4Y13_RegFile/N2BEG[1]
+ Tile_X4Y13_RegFile/N2BEG[2] Tile_X4Y13_RegFile/N2BEG[3] Tile_X4Y13_RegFile/N2BEG[4]
+ Tile_X4Y13_RegFile/N2BEG[5] Tile_X4Y13_RegFile/N2BEG[6] Tile_X4Y13_RegFile/N2BEG[7]
+ Tile_X4Y12_RegFile/N2END[0] Tile_X4Y12_RegFile/N2END[1] Tile_X4Y12_RegFile/N2END[2]
+ Tile_X4Y12_RegFile/N2END[3] Tile_X4Y12_RegFile/N2END[4] Tile_X4Y12_RegFile/N2END[5]
+ Tile_X4Y12_RegFile/N2END[6] Tile_X4Y12_RegFile/N2END[7] Tile_X4Y13_RegFile/N2END[0]
+ Tile_X4Y13_RegFile/N2END[1] Tile_X4Y13_RegFile/N2END[2] Tile_X4Y13_RegFile/N2END[3]
+ Tile_X4Y13_RegFile/N2END[4] Tile_X4Y13_RegFile/N2END[5] Tile_X4Y13_RegFile/N2END[6]
+ Tile_X4Y13_RegFile/N2END[7] Tile_X4Y14_RegFile/N2BEG[0] Tile_X4Y14_RegFile/N2BEG[1]
+ Tile_X4Y14_RegFile/N2BEG[2] Tile_X4Y14_RegFile/N2BEG[3] Tile_X4Y14_RegFile/N2BEG[4]
+ Tile_X4Y14_RegFile/N2BEG[5] Tile_X4Y14_RegFile/N2BEG[6] Tile_X4Y14_RegFile/N2BEG[7]
+ Tile_X4Y13_RegFile/N4BEG[0] Tile_X4Y13_RegFile/N4BEG[10] Tile_X4Y13_RegFile/N4BEG[11]
+ Tile_X4Y13_RegFile/N4BEG[12] Tile_X4Y13_RegFile/N4BEG[13] Tile_X4Y13_RegFile/N4BEG[14]
+ Tile_X4Y13_RegFile/N4BEG[15] Tile_X4Y13_RegFile/N4BEG[1] Tile_X4Y13_RegFile/N4BEG[2]
+ Tile_X4Y13_RegFile/N4BEG[3] Tile_X4Y13_RegFile/N4BEG[4] Tile_X4Y13_RegFile/N4BEG[5]
+ Tile_X4Y13_RegFile/N4BEG[6] Tile_X4Y13_RegFile/N4BEG[7] Tile_X4Y13_RegFile/N4BEG[8]
+ Tile_X4Y13_RegFile/N4BEG[9] Tile_X4Y14_RegFile/N4BEG[0] Tile_X4Y14_RegFile/N4BEG[10]
+ Tile_X4Y14_RegFile/N4BEG[11] Tile_X4Y14_RegFile/N4BEG[12] Tile_X4Y14_RegFile/N4BEG[13]
+ Tile_X4Y14_RegFile/N4BEG[14] Tile_X4Y14_RegFile/N4BEG[15] Tile_X4Y14_RegFile/N4BEG[1]
+ Tile_X4Y14_RegFile/N4BEG[2] Tile_X4Y14_RegFile/N4BEG[3] Tile_X4Y14_RegFile/N4BEG[4]
+ Tile_X4Y14_RegFile/N4BEG[5] Tile_X4Y14_RegFile/N4BEG[6] Tile_X4Y14_RegFile/N4BEG[7]
+ Tile_X4Y14_RegFile/N4BEG[8] Tile_X4Y14_RegFile/N4BEG[9] Tile_X4Y13_RegFile/NN4BEG[0]
+ Tile_X4Y13_RegFile/NN4BEG[10] Tile_X4Y13_RegFile/NN4BEG[11] Tile_X4Y13_RegFile/NN4BEG[12]
+ Tile_X4Y13_RegFile/NN4BEG[13] Tile_X4Y13_RegFile/NN4BEG[14] Tile_X4Y13_RegFile/NN4BEG[15]
+ Tile_X4Y13_RegFile/NN4BEG[1] Tile_X4Y13_RegFile/NN4BEG[2] Tile_X4Y13_RegFile/NN4BEG[3]
+ Tile_X4Y13_RegFile/NN4BEG[4] Tile_X4Y13_RegFile/NN4BEG[5] Tile_X4Y13_RegFile/NN4BEG[6]
+ Tile_X4Y13_RegFile/NN4BEG[7] Tile_X4Y13_RegFile/NN4BEG[8] Tile_X4Y13_RegFile/NN4BEG[9]
+ Tile_X4Y14_RegFile/NN4BEG[0] Tile_X4Y14_RegFile/NN4BEG[10] Tile_X4Y14_RegFile/NN4BEG[11]
+ Tile_X4Y14_RegFile/NN4BEG[12] Tile_X4Y14_RegFile/NN4BEG[13] Tile_X4Y14_RegFile/NN4BEG[14]
+ Tile_X4Y14_RegFile/NN4BEG[15] Tile_X4Y14_RegFile/NN4BEG[1] Tile_X4Y14_RegFile/NN4BEG[2]
+ Tile_X4Y14_RegFile/NN4BEG[3] Tile_X4Y14_RegFile/NN4BEG[4] Tile_X4Y14_RegFile/NN4BEG[5]
+ Tile_X4Y14_RegFile/NN4BEG[6] Tile_X4Y14_RegFile/NN4BEG[7] Tile_X4Y14_RegFile/NN4BEG[8]
+ Tile_X4Y14_RegFile/NN4BEG[9] Tile_X4Y14_RegFile/S1END[0] Tile_X4Y14_RegFile/S1END[1]
+ Tile_X4Y14_RegFile/S1END[2] Tile_X4Y14_RegFile/S1END[3] Tile_X4Y13_RegFile/S1END[0]
+ Tile_X4Y13_RegFile/S1END[1] Tile_X4Y13_RegFile/S1END[2] Tile_X4Y13_RegFile/S1END[3]
+ Tile_X4Y14_RegFile/S2MID[0] Tile_X4Y14_RegFile/S2MID[1] Tile_X4Y14_RegFile/S2MID[2]
+ Tile_X4Y14_RegFile/S2MID[3] Tile_X4Y14_RegFile/S2MID[4] Tile_X4Y14_RegFile/S2MID[5]
+ Tile_X4Y14_RegFile/S2MID[6] Tile_X4Y14_RegFile/S2MID[7] Tile_X4Y14_RegFile/S2END[0]
+ Tile_X4Y14_RegFile/S2END[1] Tile_X4Y14_RegFile/S2END[2] Tile_X4Y14_RegFile/S2END[3]
+ Tile_X4Y14_RegFile/S2END[4] Tile_X4Y14_RegFile/S2END[5] Tile_X4Y14_RegFile/S2END[6]
+ Tile_X4Y14_RegFile/S2END[7] Tile_X4Y13_RegFile/S2END[0] Tile_X4Y13_RegFile/S2END[1]
+ Tile_X4Y13_RegFile/S2END[2] Tile_X4Y13_RegFile/S2END[3] Tile_X4Y13_RegFile/S2END[4]
+ Tile_X4Y13_RegFile/S2END[5] Tile_X4Y13_RegFile/S2END[6] Tile_X4Y13_RegFile/S2END[7]
+ Tile_X4Y13_RegFile/S2MID[0] Tile_X4Y13_RegFile/S2MID[1] Tile_X4Y13_RegFile/S2MID[2]
+ Tile_X4Y13_RegFile/S2MID[3] Tile_X4Y13_RegFile/S2MID[4] Tile_X4Y13_RegFile/S2MID[5]
+ Tile_X4Y13_RegFile/S2MID[6] Tile_X4Y13_RegFile/S2MID[7] Tile_X4Y14_RegFile/S4END[0]
+ Tile_X4Y14_RegFile/S4END[10] Tile_X4Y14_RegFile/S4END[11] Tile_X4Y14_RegFile/S4END[12]
+ Tile_X4Y14_RegFile/S4END[13] Tile_X4Y14_RegFile/S4END[14] Tile_X4Y14_RegFile/S4END[15]
+ Tile_X4Y14_RegFile/S4END[1] Tile_X4Y14_RegFile/S4END[2] Tile_X4Y14_RegFile/S4END[3]
+ Tile_X4Y14_RegFile/S4END[4] Tile_X4Y14_RegFile/S4END[5] Tile_X4Y14_RegFile/S4END[6]
+ Tile_X4Y14_RegFile/S4END[7] Tile_X4Y14_RegFile/S4END[8] Tile_X4Y14_RegFile/S4END[9]
+ Tile_X4Y13_RegFile/S4END[0] Tile_X4Y13_RegFile/S4END[10] Tile_X4Y13_RegFile/S4END[11]
+ Tile_X4Y13_RegFile/S4END[12] Tile_X4Y13_RegFile/S4END[13] Tile_X4Y13_RegFile/S4END[14]
+ Tile_X4Y13_RegFile/S4END[15] Tile_X4Y13_RegFile/S4END[1] Tile_X4Y13_RegFile/S4END[2]
+ Tile_X4Y13_RegFile/S4END[3] Tile_X4Y13_RegFile/S4END[4] Tile_X4Y13_RegFile/S4END[5]
+ Tile_X4Y13_RegFile/S4END[6] Tile_X4Y13_RegFile/S4END[7] Tile_X4Y13_RegFile/S4END[8]
+ Tile_X4Y13_RegFile/S4END[9] Tile_X4Y14_RegFile/SS4END[0] Tile_X4Y14_RegFile/SS4END[10]
+ Tile_X4Y14_RegFile/SS4END[11] Tile_X4Y14_RegFile/SS4END[12] Tile_X4Y14_RegFile/SS4END[13]
+ Tile_X4Y14_RegFile/SS4END[14] Tile_X4Y14_RegFile/SS4END[15] Tile_X4Y14_RegFile/SS4END[1]
+ Tile_X4Y14_RegFile/SS4END[2] Tile_X4Y14_RegFile/SS4END[3] Tile_X4Y14_RegFile/SS4END[4]
+ Tile_X4Y14_RegFile/SS4END[5] Tile_X4Y14_RegFile/SS4END[6] Tile_X4Y14_RegFile/SS4END[7]
+ Tile_X4Y14_RegFile/SS4END[8] Tile_X4Y14_RegFile/SS4END[9] Tile_X4Y13_RegFile/SS4END[0]
+ Tile_X4Y13_RegFile/SS4END[10] Tile_X4Y13_RegFile/SS4END[11] Tile_X4Y13_RegFile/SS4END[12]
+ Tile_X4Y13_RegFile/SS4END[13] Tile_X4Y13_RegFile/SS4END[14] Tile_X4Y13_RegFile/SS4END[15]
+ Tile_X4Y13_RegFile/SS4END[1] Tile_X4Y13_RegFile/SS4END[2] Tile_X4Y13_RegFile/SS4END[3]
+ Tile_X4Y13_RegFile/SS4END[4] Tile_X4Y13_RegFile/SS4END[5] Tile_X4Y13_RegFile/SS4END[6]
+ Tile_X4Y13_RegFile/SS4END[7] Tile_X4Y13_RegFile/SS4END[8] Tile_X4Y13_RegFile/SS4END[9]
+ Tile_X4Y13_RegFile/UserCLK Tile_X4Y12_RegFile/UserCLK VGND VPWR Tile_X3Y13_LUT4AB/W1END[0]
+ Tile_X3Y13_LUT4AB/W1END[1] Tile_X3Y13_LUT4AB/W1END[2] Tile_X3Y13_LUT4AB/W1END[3]
+ Tile_X5Y13_LUT4AB/W1BEG[0] Tile_X5Y13_LUT4AB/W1BEG[1] Tile_X5Y13_LUT4AB/W1BEG[2]
+ Tile_X5Y13_LUT4AB/W1BEG[3] Tile_X3Y13_LUT4AB/W2MID[0] Tile_X3Y13_LUT4AB/W2MID[1]
+ Tile_X3Y13_LUT4AB/W2MID[2] Tile_X3Y13_LUT4AB/W2MID[3] Tile_X3Y13_LUT4AB/W2MID[4]
+ Tile_X3Y13_LUT4AB/W2MID[5] Tile_X3Y13_LUT4AB/W2MID[6] Tile_X3Y13_LUT4AB/W2MID[7]
+ Tile_X3Y13_LUT4AB/W2END[0] Tile_X3Y13_LUT4AB/W2END[1] Tile_X3Y13_LUT4AB/W2END[2]
+ Tile_X3Y13_LUT4AB/W2END[3] Tile_X3Y13_LUT4AB/W2END[4] Tile_X3Y13_LUT4AB/W2END[5]
+ Tile_X3Y13_LUT4AB/W2END[6] Tile_X3Y13_LUT4AB/W2END[7] Tile_X5Y13_LUT4AB/W2BEGb[0]
+ Tile_X5Y13_LUT4AB/W2BEGb[1] Tile_X5Y13_LUT4AB/W2BEGb[2] Tile_X5Y13_LUT4AB/W2BEGb[3]
+ Tile_X5Y13_LUT4AB/W2BEGb[4] Tile_X5Y13_LUT4AB/W2BEGb[5] Tile_X5Y13_LUT4AB/W2BEGb[6]
+ Tile_X5Y13_LUT4AB/W2BEGb[7] Tile_X5Y13_LUT4AB/W2BEG[0] Tile_X5Y13_LUT4AB/W2BEG[1]
+ Tile_X5Y13_LUT4AB/W2BEG[2] Tile_X5Y13_LUT4AB/W2BEG[3] Tile_X5Y13_LUT4AB/W2BEG[4]
+ Tile_X5Y13_LUT4AB/W2BEG[5] Tile_X5Y13_LUT4AB/W2BEG[6] Tile_X5Y13_LUT4AB/W2BEG[7]
+ Tile_X3Y13_LUT4AB/W6END[0] Tile_X3Y13_LUT4AB/W6END[10] Tile_X3Y13_LUT4AB/W6END[11]
+ Tile_X3Y13_LUT4AB/W6END[1] Tile_X3Y13_LUT4AB/W6END[2] Tile_X3Y13_LUT4AB/W6END[3]
+ Tile_X3Y13_LUT4AB/W6END[4] Tile_X3Y13_LUT4AB/W6END[5] Tile_X3Y13_LUT4AB/W6END[6]
+ Tile_X3Y13_LUT4AB/W6END[7] Tile_X3Y13_LUT4AB/W6END[8] Tile_X3Y13_LUT4AB/W6END[9]
+ Tile_X5Y13_LUT4AB/W6BEG[0] Tile_X5Y13_LUT4AB/W6BEG[10] Tile_X5Y13_LUT4AB/W6BEG[11]
+ Tile_X5Y13_LUT4AB/W6BEG[1] Tile_X5Y13_LUT4AB/W6BEG[2] Tile_X5Y13_LUT4AB/W6BEG[3]
+ Tile_X5Y13_LUT4AB/W6BEG[4] Tile_X5Y13_LUT4AB/W6BEG[5] Tile_X5Y13_LUT4AB/W6BEG[6]
+ Tile_X5Y13_LUT4AB/W6BEG[7] Tile_X5Y13_LUT4AB/W6BEG[8] Tile_X5Y13_LUT4AB/W6BEG[9]
+ Tile_X3Y13_LUT4AB/WW4END[0] Tile_X3Y13_LUT4AB/WW4END[10] Tile_X3Y13_LUT4AB/WW4END[11]
+ Tile_X3Y13_LUT4AB/WW4END[12] Tile_X3Y13_LUT4AB/WW4END[13] Tile_X3Y13_LUT4AB/WW4END[14]
+ Tile_X3Y13_LUT4AB/WW4END[15] Tile_X3Y13_LUT4AB/WW4END[1] Tile_X3Y13_LUT4AB/WW4END[2]
+ Tile_X3Y13_LUT4AB/WW4END[3] Tile_X3Y13_LUT4AB/WW4END[4] Tile_X3Y13_LUT4AB/WW4END[5]
+ Tile_X3Y13_LUT4AB/WW4END[6] Tile_X3Y13_LUT4AB/WW4END[7] Tile_X3Y13_LUT4AB/WW4END[8]
+ Tile_X3Y13_LUT4AB/WW4END[9] Tile_X5Y13_LUT4AB/WW4BEG[0] Tile_X5Y13_LUT4AB/WW4BEG[10]
+ Tile_X5Y13_LUT4AB/WW4BEG[11] Tile_X5Y13_LUT4AB/WW4BEG[12] Tile_X5Y13_LUT4AB/WW4BEG[13]
+ Tile_X5Y13_LUT4AB/WW4BEG[14] Tile_X5Y13_LUT4AB/WW4BEG[15] Tile_X5Y13_LUT4AB/WW4BEG[1]
+ Tile_X5Y13_LUT4AB/WW4BEG[2] Tile_X5Y13_LUT4AB/WW4BEG[3] Tile_X5Y13_LUT4AB/WW4BEG[4]
+ Tile_X5Y13_LUT4AB/WW4BEG[5] Tile_X5Y13_LUT4AB/WW4BEG[6] Tile_X5Y13_LUT4AB/WW4BEG[7]
+ Tile_X5Y13_LUT4AB/WW4BEG[8] Tile_X5Y13_LUT4AB/WW4BEG[9] RegFile
XTile_X1Y12_LUT4AB Tile_X1Y13_LUT4AB/Co Tile_X1Y12_LUT4AB/Co Tile_X2Y12_LUT4AB/E1END[0]
+ Tile_X2Y12_LUT4AB/E1END[1] Tile_X2Y12_LUT4AB/E1END[2] Tile_X2Y12_LUT4AB/E1END[3]
+ Tile_X0Y12_W_IO/E1BEG[0] Tile_X0Y12_W_IO/E1BEG[1] Tile_X0Y12_W_IO/E1BEG[2] Tile_X0Y12_W_IO/E1BEG[3]
+ Tile_X2Y12_LUT4AB/E2MID[0] Tile_X2Y12_LUT4AB/E2MID[1] Tile_X2Y12_LUT4AB/E2MID[2]
+ Tile_X2Y12_LUT4AB/E2MID[3] Tile_X2Y12_LUT4AB/E2MID[4] Tile_X2Y12_LUT4AB/E2MID[5]
+ Tile_X2Y12_LUT4AB/E2MID[6] Tile_X2Y12_LUT4AB/E2MID[7] Tile_X2Y12_LUT4AB/E2END[0]
+ Tile_X2Y12_LUT4AB/E2END[1] Tile_X2Y12_LUT4AB/E2END[2] Tile_X2Y12_LUT4AB/E2END[3]
+ Tile_X2Y12_LUT4AB/E2END[4] Tile_X2Y12_LUT4AB/E2END[5] Tile_X2Y12_LUT4AB/E2END[6]
+ Tile_X2Y12_LUT4AB/E2END[7] Tile_X0Y12_W_IO/E2BEGb[0] Tile_X0Y12_W_IO/E2BEGb[1] Tile_X0Y12_W_IO/E2BEGb[2]
+ Tile_X0Y12_W_IO/E2BEGb[3] Tile_X0Y12_W_IO/E2BEGb[4] Tile_X0Y12_W_IO/E2BEGb[5] Tile_X0Y12_W_IO/E2BEGb[6]
+ Tile_X0Y12_W_IO/E2BEGb[7] Tile_X0Y12_W_IO/E2BEG[0] Tile_X0Y12_W_IO/E2BEG[1] Tile_X0Y12_W_IO/E2BEG[2]
+ Tile_X0Y12_W_IO/E2BEG[3] Tile_X0Y12_W_IO/E2BEG[4] Tile_X0Y12_W_IO/E2BEG[5] Tile_X0Y12_W_IO/E2BEG[6]
+ Tile_X0Y12_W_IO/E2BEG[7] Tile_X2Y12_LUT4AB/E6END[0] Tile_X2Y12_LUT4AB/E6END[10]
+ Tile_X2Y12_LUT4AB/E6END[11] Tile_X2Y12_LUT4AB/E6END[1] Tile_X2Y12_LUT4AB/E6END[2]
+ Tile_X2Y12_LUT4AB/E6END[3] Tile_X2Y12_LUT4AB/E6END[4] Tile_X2Y12_LUT4AB/E6END[5]
+ Tile_X2Y12_LUT4AB/E6END[6] Tile_X2Y12_LUT4AB/E6END[7] Tile_X2Y12_LUT4AB/E6END[8]
+ Tile_X2Y12_LUT4AB/E6END[9] Tile_X0Y12_W_IO/E6BEG[0] Tile_X0Y12_W_IO/E6BEG[10] Tile_X0Y12_W_IO/E6BEG[11]
+ Tile_X0Y12_W_IO/E6BEG[1] Tile_X0Y12_W_IO/E6BEG[2] Tile_X0Y12_W_IO/E6BEG[3] Tile_X0Y12_W_IO/E6BEG[4]
+ Tile_X0Y12_W_IO/E6BEG[5] Tile_X0Y12_W_IO/E6BEG[6] Tile_X0Y12_W_IO/E6BEG[7] Tile_X0Y12_W_IO/E6BEG[8]
+ Tile_X0Y12_W_IO/E6BEG[9] Tile_X2Y12_LUT4AB/EE4END[0] Tile_X2Y12_LUT4AB/EE4END[10]
+ Tile_X2Y12_LUT4AB/EE4END[11] Tile_X2Y12_LUT4AB/EE4END[12] Tile_X2Y12_LUT4AB/EE4END[13]
+ Tile_X2Y12_LUT4AB/EE4END[14] Tile_X2Y12_LUT4AB/EE4END[15] Tile_X2Y12_LUT4AB/EE4END[1]
+ Tile_X2Y12_LUT4AB/EE4END[2] Tile_X2Y12_LUT4AB/EE4END[3] Tile_X2Y12_LUT4AB/EE4END[4]
+ Tile_X2Y12_LUT4AB/EE4END[5] Tile_X2Y12_LUT4AB/EE4END[6] Tile_X2Y12_LUT4AB/EE4END[7]
+ Tile_X2Y12_LUT4AB/EE4END[8] Tile_X2Y12_LUT4AB/EE4END[9] Tile_X0Y12_W_IO/EE4BEG[0]
+ Tile_X0Y12_W_IO/EE4BEG[10] Tile_X0Y12_W_IO/EE4BEG[11] Tile_X0Y12_W_IO/EE4BEG[12]
+ Tile_X0Y12_W_IO/EE4BEG[13] Tile_X0Y12_W_IO/EE4BEG[14] Tile_X0Y12_W_IO/EE4BEG[15]
+ Tile_X0Y12_W_IO/EE4BEG[1] Tile_X0Y12_W_IO/EE4BEG[2] Tile_X0Y12_W_IO/EE4BEG[3] Tile_X0Y12_W_IO/EE4BEG[4]
+ Tile_X0Y12_W_IO/EE4BEG[5] Tile_X0Y12_W_IO/EE4BEG[6] Tile_X0Y12_W_IO/EE4BEG[7] Tile_X0Y12_W_IO/EE4BEG[8]
+ Tile_X0Y12_W_IO/EE4BEG[9] Tile_X1Y12_LUT4AB/FrameData[0] Tile_X1Y12_LUT4AB/FrameData[10]
+ Tile_X1Y12_LUT4AB/FrameData[11] Tile_X1Y12_LUT4AB/FrameData[12] Tile_X1Y12_LUT4AB/FrameData[13]
+ Tile_X1Y12_LUT4AB/FrameData[14] Tile_X1Y12_LUT4AB/FrameData[15] Tile_X1Y12_LUT4AB/FrameData[16]
+ Tile_X1Y12_LUT4AB/FrameData[17] Tile_X1Y12_LUT4AB/FrameData[18] Tile_X1Y12_LUT4AB/FrameData[19]
+ Tile_X1Y12_LUT4AB/FrameData[1] Tile_X1Y12_LUT4AB/FrameData[20] Tile_X1Y12_LUT4AB/FrameData[21]
+ Tile_X1Y12_LUT4AB/FrameData[22] Tile_X1Y12_LUT4AB/FrameData[23] Tile_X1Y12_LUT4AB/FrameData[24]
+ Tile_X1Y12_LUT4AB/FrameData[25] Tile_X1Y12_LUT4AB/FrameData[26] Tile_X1Y12_LUT4AB/FrameData[27]
+ Tile_X1Y12_LUT4AB/FrameData[28] Tile_X1Y12_LUT4AB/FrameData[29] Tile_X1Y12_LUT4AB/FrameData[2]
+ Tile_X1Y12_LUT4AB/FrameData[30] Tile_X1Y12_LUT4AB/FrameData[31] Tile_X1Y12_LUT4AB/FrameData[3]
+ Tile_X1Y12_LUT4AB/FrameData[4] Tile_X1Y12_LUT4AB/FrameData[5] Tile_X1Y12_LUT4AB/FrameData[6]
+ Tile_X1Y12_LUT4AB/FrameData[7] Tile_X1Y12_LUT4AB/FrameData[8] Tile_X1Y12_LUT4AB/FrameData[9]
+ Tile_X2Y12_LUT4AB/FrameData[0] Tile_X2Y12_LUT4AB/FrameData[10] Tile_X2Y12_LUT4AB/FrameData[11]
+ Tile_X2Y12_LUT4AB/FrameData[12] Tile_X2Y12_LUT4AB/FrameData[13] Tile_X2Y12_LUT4AB/FrameData[14]
+ Tile_X2Y12_LUT4AB/FrameData[15] Tile_X2Y12_LUT4AB/FrameData[16] Tile_X2Y12_LUT4AB/FrameData[17]
+ Tile_X2Y12_LUT4AB/FrameData[18] Tile_X2Y12_LUT4AB/FrameData[19] Tile_X2Y12_LUT4AB/FrameData[1]
+ Tile_X2Y12_LUT4AB/FrameData[20] Tile_X2Y12_LUT4AB/FrameData[21] Tile_X2Y12_LUT4AB/FrameData[22]
+ Tile_X2Y12_LUT4AB/FrameData[23] Tile_X2Y12_LUT4AB/FrameData[24] Tile_X2Y12_LUT4AB/FrameData[25]
+ Tile_X2Y12_LUT4AB/FrameData[26] Tile_X2Y12_LUT4AB/FrameData[27] Tile_X2Y12_LUT4AB/FrameData[28]
+ Tile_X2Y12_LUT4AB/FrameData[29] Tile_X2Y12_LUT4AB/FrameData[2] Tile_X2Y12_LUT4AB/FrameData[30]
+ Tile_X2Y12_LUT4AB/FrameData[31] Tile_X2Y12_LUT4AB/FrameData[3] Tile_X2Y12_LUT4AB/FrameData[4]
+ Tile_X2Y12_LUT4AB/FrameData[5] Tile_X2Y12_LUT4AB/FrameData[6] Tile_X2Y12_LUT4AB/FrameData[7]
+ Tile_X2Y12_LUT4AB/FrameData[8] Tile_X2Y12_LUT4AB/FrameData[9] Tile_X1Y12_LUT4AB/FrameStrobe[0]
+ Tile_X1Y12_LUT4AB/FrameStrobe[10] Tile_X1Y12_LUT4AB/FrameStrobe[11] Tile_X1Y12_LUT4AB/FrameStrobe[12]
+ Tile_X1Y12_LUT4AB/FrameStrobe[13] Tile_X1Y12_LUT4AB/FrameStrobe[14] Tile_X1Y12_LUT4AB/FrameStrobe[15]
+ Tile_X1Y12_LUT4AB/FrameStrobe[16] Tile_X1Y12_LUT4AB/FrameStrobe[17] Tile_X1Y12_LUT4AB/FrameStrobe[18]
+ Tile_X1Y12_LUT4AB/FrameStrobe[19] Tile_X1Y12_LUT4AB/FrameStrobe[1] Tile_X1Y12_LUT4AB/FrameStrobe[2]
+ Tile_X1Y12_LUT4AB/FrameStrobe[3] Tile_X1Y12_LUT4AB/FrameStrobe[4] Tile_X1Y12_LUT4AB/FrameStrobe[5]
+ Tile_X1Y12_LUT4AB/FrameStrobe[6] Tile_X1Y12_LUT4AB/FrameStrobe[7] Tile_X1Y12_LUT4AB/FrameStrobe[8]
+ Tile_X1Y12_LUT4AB/FrameStrobe[9] Tile_X1Y11_LUT4AB/FrameStrobe[0] Tile_X1Y11_LUT4AB/FrameStrobe[10]
+ Tile_X1Y11_LUT4AB/FrameStrobe[11] Tile_X1Y11_LUT4AB/FrameStrobe[12] Tile_X1Y11_LUT4AB/FrameStrobe[13]
+ Tile_X1Y11_LUT4AB/FrameStrobe[14] Tile_X1Y11_LUT4AB/FrameStrobe[15] Tile_X1Y11_LUT4AB/FrameStrobe[16]
+ Tile_X1Y11_LUT4AB/FrameStrobe[17] Tile_X1Y11_LUT4AB/FrameStrobe[18] Tile_X1Y11_LUT4AB/FrameStrobe[19]
+ Tile_X1Y11_LUT4AB/FrameStrobe[1] Tile_X1Y11_LUT4AB/FrameStrobe[2] Tile_X1Y11_LUT4AB/FrameStrobe[3]
+ Tile_X1Y11_LUT4AB/FrameStrobe[4] Tile_X1Y11_LUT4AB/FrameStrobe[5] Tile_X1Y11_LUT4AB/FrameStrobe[6]
+ Tile_X1Y11_LUT4AB/FrameStrobe[7] Tile_X1Y11_LUT4AB/FrameStrobe[8] Tile_X1Y11_LUT4AB/FrameStrobe[9]
+ Tile_X1Y12_LUT4AB/N1BEG[0] Tile_X1Y12_LUT4AB/N1BEG[1] Tile_X1Y12_LUT4AB/N1BEG[2]
+ Tile_X1Y12_LUT4AB/N1BEG[3] Tile_X1Y13_LUT4AB/N1BEG[0] Tile_X1Y13_LUT4AB/N1BEG[1]
+ Tile_X1Y13_LUT4AB/N1BEG[2] Tile_X1Y13_LUT4AB/N1BEG[3] Tile_X1Y12_LUT4AB/N2BEG[0]
+ Tile_X1Y12_LUT4AB/N2BEG[1] Tile_X1Y12_LUT4AB/N2BEG[2] Tile_X1Y12_LUT4AB/N2BEG[3]
+ Tile_X1Y12_LUT4AB/N2BEG[4] Tile_X1Y12_LUT4AB/N2BEG[5] Tile_X1Y12_LUT4AB/N2BEG[6]
+ Tile_X1Y12_LUT4AB/N2BEG[7] Tile_X1Y11_LUT4AB/N2END[0] Tile_X1Y11_LUT4AB/N2END[1]
+ Tile_X1Y11_LUT4AB/N2END[2] Tile_X1Y11_LUT4AB/N2END[3] Tile_X1Y11_LUT4AB/N2END[4]
+ Tile_X1Y11_LUT4AB/N2END[5] Tile_X1Y11_LUT4AB/N2END[6] Tile_X1Y11_LUT4AB/N2END[7]
+ Tile_X1Y12_LUT4AB/N2END[0] Tile_X1Y12_LUT4AB/N2END[1] Tile_X1Y12_LUT4AB/N2END[2]
+ Tile_X1Y12_LUT4AB/N2END[3] Tile_X1Y12_LUT4AB/N2END[4] Tile_X1Y12_LUT4AB/N2END[5]
+ Tile_X1Y12_LUT4AB/N2END[6] Tile_X1Y12_LUT4AB/N2END[7] Tile_X1Y13_LUT4AB/N2BEG[0]
+ Tile_X1Y13_LUT4AB/N2BEG[1] Tile_X1Y13_LUT4AB/N2BEG[2] Tile_X1Y13_LUT4AB/N2BEG[3]
+ Tile_X1Y13_LUT4AB/N2BEG[4] Tile_X1Y13_LUT4AB/N2BEG[5] Tile_X1Y13_LUT4AB/N2BEG[6]
+ Tile_X1Y13_LUT4AB/N2BEG[7] Tile_X1Y12_LUT4AB/N4BEG[0] Tile_X1Y12_LUT4AB/N4BEG[10]
+ Tile_X1Y12_LUT4AB/N4BEG[11] Tile_X1Y12_LUT4AB/N4BEG[12] Tile_X1Y12_LUT4AB/N4BEG[13]
+ Tile_X1Y12_LUT4AB/N4BEG[14] Tile_X1Y12_LUT4AB/N4BEG[15] Tile_X1Y12_LUT4AB/N4BEG[1]
+ Tile_X1Y12_LUT4AB/N4BEG[2] Tile_X1Y12_LUT4AB/N4BEG[3] Tile_X1Y12_LUT4AB/N4BEG[4]
+ Tile_X1Y12_LUT4AB/N4BEG[5] Tile_X1Y12_LUT4AB/N4BEG[6] Tile_X1Y12_LUT4AB/N4BEG[7]
+ Tile_X1Y12_LUT4AB/N4BEG[8] Tile_X1Y12_LUT4AB/N4BEG[9] Tile_X1Y13_LUT4AB/N4BEG[0]
+ Tile_X1Y13_LUT4AB/N4BEG[10] Tile_X1Y13_LUT4AB/N4BEG[11] Tile_X1Y13_LUT4AB/N4BEG[12]
+ Tile_X1Y13_LUT4AB/N4BEG[13] Tile_X1Y13_LUT4AB/N4BEG[14] Tile_X1Y13_LUT4AB/N4BEG[15]
+ Tile_X1Y13_LUT4AB/N4BEG[1] Tile_X1Y13_LUT4AB/N4BEG[2] Tile_X1Y13_LUT4AB/N4BEG[3]
+ Tile_X1Y13_LUT4AB/N4BEG[4] Tile_X1Y13_LUT4AB/N4BEG[5] Tile_X1Y13_LUT4AB/N4BEG[6]
+ Tile_X1Y13_LUT4AB/N4BEG[7] Tile_X1Y13_LUT4AB/N4BEG[8] Tile_X1Y13_LUT4AB/N4BEG[9]
+ Tile_X1Y12_LUT4AB/NN4BEG[0] Tile_X1Y12_LUT4AB/NN4BEG[10] Tile_X1Y12_LUT4AB/NN4BEG[11]
+ Tile_X1Y12_LUT4AB/NN4BEG[12] Tile_X1Y12_LUT4AB/NN4BEG[13] Tile_X1Y12_LUT4AB/NN4BEG[14]
+ Tile_X1Y12_LUT4AB/NN4BEG[15] Tile_X1Y12_LUT4AB/NN4BEG[1] Tile_X1Y12_LUT4AB/NN4BEG[2]
+ Tile_X1Y12_LUT4AB/NN4BEG[3] Tile_X1Y12_LUT4AB/NN4BEG[4] Tile_X1Y12_LUT4AB/NN4BEG[5]
+ Tile_X1Y12_LUT4AB/NN4BEG[6] Tile_X1Y12_LUT4AB/NN4BEG[7] Tile_X1Y12_LUT4AB/NN4BEG[8]
+ Tile_X1Y12_LUT4AB/NN4BEG[9] Tile_X1Y13_LUT4AB/NN4BEG[0] Tile_X1Y13_LUT4AB/NN4BEG[10]
+ Tile_X1Y13_LUT4AB/NN4BEG[11] Tile_X1Y13_LUT4AB/NN4BEG[12] Tile_X1Y13_LUT4AB/NN4BEG[13]
+ Tile_X1Y13_LUT4AB/NN4BEG[14] Tile_X1Y13_LUT4AB/NN4BEG[15] Tile_X1Y13_LUT4AB/NN4BEG[1]
+ Tile_X1Y13_LUT4AB/NN4BEG[2] Tile_X1Y13_LUT4AB/NN4BEG[3] Tile_X1Y13_LUT4AB/NN4BEG[4]
+ Tile_X1Y13_LUT4AB/NN4BEG[5] Tile_X1Y13_LUT4AB/NN4BEG[6] Tile_X1Y13_LUT4AB/NN4BEG[7]
+ Tile_X1Y13_LUT4AB/NN4BEG[8] Tile_X1Y13_LUT4AB/NN4BEG[9] Tile_X1Y13_LUT4AB/S1END[0]
+ Tile_X1Y13_LUT4AB/S1END[1] Tile_X1Y13_LUT4AB/S1END[2] Tile_X1Y13_LUT4AB/S1END[3]
+ Tile_X1Y12_LUT4AB/S1END[0] Tile_X1Y12_LUT4AB/S1END[1] Tile_X1Y12_LUT4AB/S1END[2]
+ Tile_X1Y12_LUT4AB/S1END[3] Tile_X1Y13_LUT4AB/S2MID[0] Tile_X1Y13_LUT4AB/S2MID[1]
+ Tile_X1Y13_LUT4AB/S2MID[2] Tile_X1Y13_LUT4AB/S2MID[3] Tile_X1Y13_LUT4AB/S2MID[4]
+ Tile_X1Y13_LUT4AB/S2MID[5] Tile_X1Y13_LUT4AB/S2MID[6] Tile_X1Y13_LUT4AB/S2MID[7]
+ Tile_X1Y13_LUT4AB/S2END[0] Tile_X1Y13_LUT4AB/S2END[1] Tile_X1Y13_LUT4AB/S2END[2]
+ Tile_X1Y13_LUT4AB/S2END[3] Tile_X1Y13_LUT4AB/S2END[4] Tile_X1Y13_LUT4AB/S2END[5]
+ Tile_X1Y13_LUT4AB/S2END[6] Tile_X1Y13_LUT4AB/S2END[7] Tile_X1Y12_LUT4AB/S2END[0]
+ Tile_X1Y12_LUT4AB/S2END[1] Tile_X1Y12_LUT4AB/S2END[2] Tile_X1Y12_LUT4AB/S2END[3]
+ Tile_X1Y12_LUT4AB/S2END[4] Tile_X1Y12_LUT4AB/S2END[5] Tile_X1Y12_LUT4AB/S2END[6]
+ Tile_X1Y12_LUT4AB/S2END[7] Tile_X1Y12_LUT4AB/S2MID[0] Tile_X1Y12_LUT4AB/S2MID[1]
+ Tile_X1Y12_LUT4AB/S2MID[2] Tile_X1Y12_LUT4AB/S2MID[3] Tile_X1Y12_LUT4AB/S2MID[4]
+ Tile_X1Y12_LUT4AB/S2MID[5] Tile_X1Y12_LUT4AB/S2MID[6] Tile_X1Y12_LUT4AB/S2MID[7]
+ Tile_X1Y13_LUT4AB/S4END[0] Tile_X1Y13_LUT4AB/S4END[10] Tile_X1Y13_LUT4AB/S4END[11]
+ Tile_X1Y13_LUT4AB/S4END[12] Tile_X1Y13_LUT4AB/S4END[13] Tile_X1Y13_LUT4AB/S4END[14]
+ Tile_X1Y13_LUT4AB/S4END[15] Tile_X1Y13_LUT4AB/S4END[1] Tile_X1Y13_LUT4AB/S4END[2]
+ Tile_X1Y13_LUT4AB/S4END[3] Tile_X1Y13_LUT4AB/S4END[4] Tile_X1Y13_LUT4AB/S4END[5]
+ Tile_X1Y13_LUT4AB/S4END[6] Tile_X1Y13_LUT4AB/S4END[7] Tile_X1Y13_LUT4AB/S4END[8]
+ Tile_X1Y13_LUT4AB/S4END[9] Tile_X1Y12_LUT4AB/S4END[0] Tile_X1Y12_LUT4AB/S4END[10]
+ Tile_X1Y12_LUT4AB/S4END[11] Tile_X1Y12_LUT4AB/S4END[12] Tile_X1Y12_LUT4AB/S4END[13]
+ Tile_X1Y12_LUT4AB/S4END[14] Tile_X1Y12_LUT4AB/S4END[15] Tile_X1Y12_LUT4AB/S4END[1]
+ Tile_X1Y12_LUT4AB/S4END[2] Tile_X1Y12_LUT4AB/S4END[3] Tile_X1Y12_LUT4AB/S4END[4]
+ Tile_X1Y12_LUT4AB/S4END[5] Tile_X1Y12_LUT4AB/S4END[6] Tile_X1Y12_LUT4AB/S4END[7]
+ Tile_X1Y12_LUT4AB/S4END[8] Tile_X1Y12_LUT4AB/S4END[9] Tile_X1Y13_LUT4AB/SS4END[0]
+ Tile_X1Y13_LUT4AB/SS4END[10] Tile_X1Y13_LUT4AB/SS4END[11] Tile_X1Y13_LUT4AB/SS4END[12]
+ Tile_X1Y13_LUT4AB/SS4END[13] Tile_X1Y13_LUT4AB/SS4END[14] Tile_X1Y13_LUT4AB/SS4END[15]
+ Tile_X1Y13_LUT4AB/SS4END[1] Tile_X1Y13_LUT4AB/SS4END[2] Tile_X1Y13_LUT4AB/SS4END[3]
+ Tile_X1Y13_LUT4AB/SS4END[4] Tile_X1Y13_LUT4AB/SS4END[5] Tile_X1Y13_LUT4AB/SS4END[6]
+ Tile_X1Y13_LUT4AB/SS4END[7] Tile_X1Y13_LUT4AB/SS4END[8] Tile_X1Y13_LUT4AB/SS4END[9]
+ Tile_X1Y12_LUT4AB/SS4END[0] Tile_X1Y12_LUT4AB/SS4END[10] Tile_X1Y12_LUT4AB/SS4END[11]
+ Tile_X1Y12_LUT4AB/SS4END[12] Tile_X1Y12_LUT4AB/SS4END[13] Tile_X1Y12_LUT4AB/SS4END[14]
+ Tile_X1Y12_LUT4AB/SS4END[15] Tile_X1Y12_LUT4AB/SS4END[1] Tile_X1Y12_LUT4AB/SS4END[2]
+ Tile_X1Y12_LUT4AB/SS4END[3] Tile_X1Y12_LUT4AB/SS4END[4] Tile_X1Y12_LUT4AB/SS4END[5]
+ Tile_X1Y12_LUT4AB/SS4END[6] Tile_X1Y12_LUT4AB/SS4END[7] Tile_X1Y12_LUT4AB/SS4END[8]
+ Tile_X1Y12_LUT4AB/SS4END[9] Tile_X1Y12_LUT4AB/UserCLK Tile_X1Y11_LUT4AB/UserCLK
+ VGND VPWR Tile_X0Y12_W_IO/W1END[0] Tile_X0Y12_W_IO/W1END[1] Tile_X0Y12_W_IO/W1END[2]
+ Tile_X0Y12_W_IO/W1END[3] Tile_X2Y12_LUT4AB/W1BEG[0] Tile_X2Y12_LUT4AB/W1BEG[1] Tile_X2Y12_LUT4AB/W1BEG[2]
+ Tile_X2Y12_LUT4AB/W1BEG[3] Tile_X0Y12_W_IO/W2MID[0] Tile_X0Y12_W_IO/W2MID[1] Tile_X0Y12_W_IO/W2MID[2]
+ Tile_X0Y12_W_IO/W2MID[3] Tile_X0Y12_W_IO/W2MID[4] Tile_X0Y12_W_IO/W2MID[5] Tile_X0Y12_W_IO/W2MID[6]
+ Tile_X0Y12_W_IO/W2MID[7] Tile_X0Y12_W_IO/W2END[0] Tile_X0Y12_W_IO/W2END[1] Tile_X0Y12_W_IO/W2END[2]
+ Tile_X0Y12_W_IO/W2END[3] Tile_X0Y12_W_IO/W2END[4] Tile_X0Y12_W_IO/W2END[5] Tile_X0Y12_W_IO/W2END[6]
+ Tile_X0Y12_W_IO/W2END[7] Tile_X1Y12_LUT4AB/W2END[0] Tile_X1Y12_LUT4AB/W2END[1] Tile_X1Y12_LUT4AB/W2END[2]
+ Tile_X1Y12_LUT4AB/W2END[3] Tile_X1Y12_LUT4AB/W2END[4] Tile_X1Y12_LUT4AB/W2END[5]
+ Tile_X1Y12_LUT4AB/W2END[6] Tile_X1Y12_LUT4AB/W2END[7] Tile_X2Y12_LUT4AB/W2BEG[0]
+ Tile_X2Y12_LUT4AB/W2BEG[1] Tile_X2Y12_LUT4AB/W2BEG[2] Tile_X2Y12_LUT4AB/W2BEG[3]
+ Tile_X2Y12_LUT4AB/W2BEG[4] Tile_X2Y12_LUT4AB/W2BEG[5] Tile_X2Y12_LUT4AB/W2BEG[6]
+ Tile_X2Y12_LUT4AB/W2BEG[7] Tile_X0Y12_W_IO/W6END[0] Tile_X0Y12_W_IO/W6END[10] Tile_X0Y12_W_IO/W6END[11]
+ Tile_X0Y12_W_IO/W6END[1] Tile_X0Y12_W_IO/W6END[2] Tile_X0Y12_W_IO/W6END[3] Tile_X0Y12_W_IO/W6END[4]
+ Tile_X0Y12_W_IO/W6END[5] Tile_X0Y12_W_IO/W6END[6] Tile_X0Y12_W_IO/W6END[7] Tile_X0Y12_W_IO/W6END[8]
+ Tile_X0Y12_W_IO/W6END[9] Tile_X2Y12_LUT4AB/W6BEG[0] Tile_X2Y12_LUT4AB/W6BEG[10]
+ Tile_X2Y12_LUT4AB/W6BEG[11] Tile_X2Y12_LUT4AB/W6BEG[1] Tile_X2Y12_LUT4AB/W6BEG[2]
+ Tile_X2Y12_LUT4AB/W6BEG[3] Tile_X2Y12_LUT4AB/W6BEG[4] Tile_X2Y12_LUT4AB/W6BEG[5]
+ Tile_X2Y12_LUT4AB/W6BEG[6] Tile_X2Y12_LUT4AB/W6BEG[7] Tile_X2Y12_LUT4AB/W6BEG[8]
+ Tile_X2Y12_LUT4AB/W6BEG[9] Tile_X0Y12_W_IO/WW4END[0] Tile_X0Y12_W_IO/WW4END[10]
+ Tile_X0Y12_W_IO/WW4END[11] Tile_X0Y12_W_IO/WW4END[12] Tile_X0Y12_W_IO/WW4END[13]
+ Tile_X0Y12_W_IO/WW4END[14] Tile_X0Y12_W_IO/WW4END[15] Tile_X0Y12_W_IO/WW4END[1]
+ Tile_X0Y12_W_IO/WW4END[2] Tile_X0Y12_W_IO/WW4END[3] Tile_X0Y12_W_IO/WW4END[4] Tile_X0Y12_W_IO/WW4END[5]
+ Tile_X0Y12_W_IO/WW4END[6] Tile_X0Y12_W_IO/WW4END[7] Tile_X0Y12_W_IO/WW4END[8] Tile_X0Y12_W_IO/WW4END[9]
+ Tile_X2Y12_LUT4AB/WW4BEG[0] Tile_X2Y12_LUT4AB/WW4BEG[10] Tile_X2Y12_LUT4AB/WW4BEG[11]
+ Tile_X2Y12_LUT4AB/WW4BEG[12] Tile_X2Y12_LUT4AB/WW4BEG[13] Tile_X2Y12_LUT4AB/WW4BEG[14]
+ Tile_X2Y12_LUT4AB/WW4BEG[15] Tile_X2Y12_LUT4AB/WW4BEG[1] Tile_X2Y12_LUT4AB/WW4BEG[2]
+ Tile_X2Y12_LUT4AB/WW4BEG[3] Tile_X2Y12_LUT4AB/WW4BEG[4] Tile_X2Y12_LUT4AB/WW4BEG[5]
+ Tile_X2Y12_LUT4AB/WW4BEG[6] Tile_X2Y12_LUT4AB/WW4BEG[7] Tile_X2Y12_LUT4AB/WW4BEG[8]
+ Tile_X2Y12_LUT4AB/WW4BEG[9] LUT4AB
XTile_X6Y7_LUT4AB Tile_X6Y8_LUT4AB/Co Tile_X6Y7_LUT4AB/Co Tile_X6Y7_LUT4AB/E1BEG[0]
+ Tile_X6Y7_LUT4AB/E1BEG[1] Tile_X6Y7_LUT4AB/E1BEG[2] Tile_X6Y7_LUT4AB/E1BEG[3] Tile_X6Y7_LUT4AB/E1END[0]
+ Tile_X6Y7_LUT4AB/E1END[1] Tile_X6Y7_LUT4AB/E1END[2] Tile_X6Y7_LUT4AB/E1END[3] Tile_X6Y7_LUT4AB/E2BEG[0]
+ Tile_X6Y7_LUT4AB/E2BEG[1] Tile_X6Y7_LUT4AB/E2BEG[2] Tile_X6Y7_LUT4AB/E2BEG[3] Tile_X6Y7_LUT4AB/E2BEG[4]
+ Tile_X6Y7_LUT4AB/E2BEG[5] Tile_X6Y7_LUT4AB/E2BEG[6] Tile_X6Y7_LUT4AB/E2BEG[7] Tile_X6Y7_LUT4AB/E2BEGb[0]
+ Tile_X6Y7_LUT4AB/E2BEGb[1] Tile_X6Y7_LUT4AB/E2BEGb[2] Tile_X6Y7_LUT4AB/E2BEGb[3]
+ Tile_X6Y7_LUT4AB/E2BEGb[4] Tile_X6Y7_LUT4AB/E2BEGb[5] Tile_X6Y7_LUT4AB/E2BEGb[6]
+ Tile_X6Y7_LUT4AB/E2BEGb[7] Tile_X6Y7_LUT4AB/E2END[0] Tile_X6Y7_LUT4AB/E2END[1] Tile_X6Y7_LUT4AB/E2END[2]
+ Tile_X6Y7_LUT4AB/E2END[3] Tile_X6Y7_LUT4AB/E2END[4] Tile_X6Y7_LUT4AB/E2END[5] Tile_X6Y7_LUT4AB/E2END[6]
+ Tile_X6Y7_LUT4AB/E2END[7] Tile_X6Y7_LUT4AB/E2MID[0] Tile_X6Y7_LUT4AB/E2MID[1] Tile_X6Y7_LUT4AB/E2MID[2]
+ Tile_X6Y7_LUT4AB/E2MID[3] Tile_X6Y7_LUT4AB/E2MID[4] Tile_X6Y7_LUT4AB/E2MID[5] Tile_X6Y7_LUT4AB/E2MID[6]
+ Tile_X6Y7_LUT4AB/E2MID[7] Tile_X6Y7_LUT4AB/E6BEG[0] Tile_X6Y7_LUT4AB/E6BEG[10] Tile_X6Y7_LUT4AB/E6BEG[11]
+ Tile_X6Y7_LUT4AB/E6BEG[1] Tile_X6Y7_LUT4AB/E6BEG[2] Tile_X6Y7_LUT4AB/E6BEG[3] Tile_X6Y7_LUT4AB/E6BEG[4]
+ Tile_X6Y7_LUT4AB/E6BEG[5] Tile_X6Y7_LUT4AB/E6BEG[6] Tile_X6Y7_LUT4AB/E6BEG[7] Tile_X6Y7_LUT4AB/E6BEG[8]
+ Tile_X6Y7_LUT4AB/E6BEG[9] Tile_X6Y7_LUT4AB/E6END[0] Tile_X6Y7_LUT4AB/E6END[10] Tile_X6Y7_LUT4AB/E6END[11]
+ Tile_X6Y7_LUT4AB/E6END[1] Tile_X6Y7_LUT4AB/E6END[2] Tile_X6Y7_LUT4AB/E6END[3] Tile_X6Y7_LUT4AB/E6END[4]
+ Tile_X6Y7_LUT4AB/E6END[5] Tile_X6Y7_LUT4AB/E6END[6] Tile_X6Y7_LUT4AB/E6END[7] Tile_X6Y7_LUT4AB/E6END[8]
+ Tile_X6Y7_LUT4AB/E6END[9] Tile_X6Y7_LUT4AB/EE4BEG[0] Tile_X6Y7_LUT4AB/EE4BEG[10]
+ Tile_X6Y7_LUT4AB/EE4BEG[11] Tile_X6Y7_LUT4AB/EE4BEG[12] Tile_X6Y7_LUT4AB/EE4BEG[13]
+ Tile_X6Y7_LUT4AB/EE4BEG[14] Tile_X6Y7_LUT4AB/EE4BEG[15] Tile_X6Y7_LUT4AB/EE4BEG[1]
+ Tile_X6Y7_LUT4AB/EE4BEG[2] Tile_X6Y7_LUT4AB/EE4BEG[3] Tile_X6Y7_LUT4AB/EE4BEG[4]
+ Tile_X6Y7_LUT4AB/EE4BEG[5] Tile_X6Y7_LUT4AB/EE4BEG[6] Tile_X6Y7_LUT4AB/EE4BEG[7]
+ Tile_X6Y7_LUT4AB/EE4BEG[8] Tile_X6Y7_LUT4AB/EE4BEG[9] Tile_X6Y7_LUT4AB/EE4END[0]
+ Tile_X6Y7_LUT4AB/EE4END[10] Tile_X6Y7_LUT4AB/EE4END[11] Tile_X6Y7_LUT4AB/EE4END[12]
+ Tile_X6Y7_LUT4AB/EE4END[13] Tile_X6Y7_LUT4AB/EE4END[14] Tile_X6Y7_LUT4AB/EE4END[15]
+ Tile_X6Y7_LUT4AB/EE4END[1] Tile_X6Y7_LUT4AB/EE4END[2] Tile_X6Y7_LUT4AB/EE4END[3]
+ Tile_X6Y7_LUT4AB/EE4END[4] Tile_X6Y7_LUT4AB/EE4END[5] Tile_X6Y7_LUT4AB/EE4END[6]
+ Tile_X6Y7_LUT4AB/EE4END[7] Tile_X6Y7_LUT4AB/EE4END[8] Tile_X6Y7_LUT4AB/EE4END[9]
+ Tile_X6Y7_LUT4AB/FrameData[0] Tile_X6Y7_LUT4AB/FrameData[10] Tile_X6Y7_LUT4AB/FrameData[11]
+ Tile_X6Y7_LUT4AB/FrameData[12] Tile_X6Y7_LUT4AB/FrameData[13] Tile_X6Y7_LUT4AB/FrameData[14]
+ Tile_X6Y7_LUT4AB/FrameData[15] Tile_X6Y7_LUT4AB/FrameData[16] Tile_X6Y7_LUT4AB/FrameData[17]
+ Tile_X6Y7_LUT4AB/FrameData[18] Tile_X6Y7_LUT4AB/FrameData[19] Tile_X6Y7_LUT4AB/FrameData[1]
+ Tile_X6Y7_LUT4AB/FrameData[20] Tile_X6Y7_LUT4AB/FrameData[21] Tile_X6Y7_LUT4AB/FrameData[22]
+ Tile_X6Y7_LUT4AB/FrameData[23] Tile_X6Y7_LUT4AB/FrameData[24] Tile_X6Y7_LUT4AB/FrameData[25]
+ Tile_X6Y7_LUT4AB/FrameData[26] Tile_X6Y7_LUT4AB/FrameData[27] Tile_X6Y7_LUT4AB/FrameData[28]
+ Tile_X6Y7_LUT4AB/FrameData[29] Tile_X6Y7_LUT4AB/FrameData[2] Tile_X6Y7_LUT4AB/FrameData[30]
+ Tile_X6Y7_LUT4AB/FrameData[31] Tile_X6Y7_LUT4AB/FrameData[3] Tile_X6Y7_LUT4AB/FrameData[4]
+ Tile_X6Y7_LUT4AB/FrameData[5] Tile_X6Y7_LUT4AB/FrameData[6] Tile_X6Y7_LUT4AB/FrameData[7]
+ Tile_X6Y7_LUT4AB/FrameData[8] Tile_X6Y7_LUT4AB/FrameData[9] Tile_X6Y7_LUT4AB/FrameData_O[0]
+ Tile_X6Y7_LUT4AB/FrameData_O[10] Tile_X6Y7_LUT4AB/FrameData_O[11] Tile_X6Y7_LUT4AB/FrameData_O[12]
+ Tile_X6Y7_LUT4AB/FrameData_O[13] Tile_X6Y7_LUT4AB/FrameData_O[14] Tile_X6Y7_LUT4AB/FrameData_O[15]
+ Tile_X6Y7_LUT4AB/FrameData_O[16] Tile_X6Y7_LUT4AB/FrameData_O[17] Tile_X6Y7_LUT4AB/FrameData_O[18]
+ Tile_X6Y7_LUT4AB/FrameData_O[19] Tile_X6Y7_LUT4AB/FrameData_O[1] Tile_X6Y7_LUT4AB/FrameData_O[20]
+ Tile_X6Y7_LUT4AB/FrameData_O[21] Tile_X6Y7_LUT4AB/FrameData_O[22] Tile_X6Y7_LUT4AB/FrameData_O[23]
+ Tile_X6Y7_LUT4AB/FrameData_O[24] Tile_X6Y7_LUT4AB/FrameData_O[25] Tile_X6Y7_LUT4AB/FrameData_O[26]
+ Tile_X6Y7_LUT4AB/FrameData_O[27] Tile_X6Y7_LUT4AB/FrameData_O[28] Tile_X6Y7_LUT4AB/FrameData_O[29]
+ Tile_X6Y7_LUT4AB/FrameData_O[2] Tile_X6Y7_LUT4AB/FrameData_O[30] Tile_X6Y7_LUT4AB/FrameData_O[31]
+ Tile_X6Y7_LUT4AB/FrameData_O[3] Tile_X6Y7_LUT4AB/FrameData_O[4] Tile_X6Y7_LUT4AB/FrameData_O[5]
+ Tile_X6Y7_LUT4AB/FrameData_O[6] Tile_X6Y7_LUT4AB/FrameData_O[7] Tile_X6Y7_LUT4AB/FrameData_O[8]
+ Tile_X6Y7_LUT4AB/FrameData_O[9] Tile_X6Y7_LUT4AB/FrameStrobe[0] Tile_X6Y7_LUT4AB/FrameStrobe[10]
+ Tile_X6Y7_LUT4AB/FrameStrobe[11] Tile_X6Y7_LUT4AB/FrameStrobe[12] Tile_X6Y7_LUT4AB/FrameStrobe[13]
+ Tile_X6Y7_LUT4AB/FrameStrobe[14] Tile_X6Y7_LUT4AB/FrameStrobe[15] Tile_X6Y7_LUT4AB/FrameStrobe[16]
+ Tile_X6Y7_LUT4AB/FrameStrobe[17] Tile_X6Y7_LUT4AB/FrameStrobe[18] Tile_X6Y7_LUT4AB/FrameStrobe[19]
+ Tile_X6Y7_LUT4AB/FrameStrobe[1] Tile_X6Y7_LUT4AB/FrameStrobe[2] Tile_X6Y7_LUT4AB/FrameStrobe[3]
+ Tile_X6Y7_LUT4AB/FrameStrobe[4] Tile_X6Y7_LUT4AB/FrameStrobe[5] Tile_X6Y7_LUT4AB/FrameStrobe[6]
+ Tile_X6Y7_LUT4AB/FrameStrobe[7] Tile_X6Y7_LUT4AB/FrameStrobe[8] Tile_X6Y7_LUT4AB/FrameStrobe[9]
+ Tile_X6Y6_LUT4AB/FrameStrobe[0] Tile_X6Y6_LUT4AB/FrameStrobe[10] Tile_X6Y6_LUT4AB/FrameStrobe[11]
+ Tile_X6Y6_LUT4AB/FrameStrobe[12] Tile_X6Y6_LUT4AB/FrameStrobe[13] Tile_X6Y6_LUT4AB/FrameStrobe[14]
+ Tile_X6Y6_LUT4AB/FrameStrobe[15] Tile_X6Y6_LUT4AB/FrameStrobe[16] Tile_X6Y6_LUT4AB/FrameStrobe[17]
+ Tile_X6Y6_LUT4AB/FrameStrobe[18] Tile_X6Y6_LUT4AB/FrameStrobe[19] Tile_X6Y6_LUT4AB/FrameStrobe[1]
+ Tile_X6Y6_LUT4AB/FrameStrobe[2] Tile_X6Y6_LUT4AB/FrameStrobe[3] Tile_X6Y6_LUT4AB/FrameStrobe[4]
+ Tile_X6Y6_LUT4AB/FrameStrobe[5] Tile_X6Y6_LUT4AB/FrameStrobe[6] Tile_X6Y6_LUT4AB/FrameStrobe[7]
+ Tile_X6Y6_LUT4AB/FrameStrobe[8] Tile_X6Y6_LUT4AB/FrameStrobe[9] Tile_X6Y7_LUT4AB/N1BEG[0]
+ Tile_X6Y7_LUT4AB/N1BEG[1] Tile_X6Y7_LUT4AB/N1BEG[2] Tile_X6Y7_LUT4AB/N1BEG[3] Tile_X6Y8_LUT4AB/N1BEG[0]
+ Tile_X6Y8_LUT4AB/N1BEG[1] Tile_X6Y8_LUT4AB/N1BEG[2] Tile_X6Y8_LUT4AB/N1BEG[3] Tile_X6Y7_LUT4AB/N2BEG[0]
+ Tile_X6Y7_LUT4AB/N2BEG[1] Tile_X6Y7_LUT4AB/N2BEG[2] Tile_X6Y7_LUT4AB/N2BEG[3] Tile_X6Y7_LUT4AB/N2BEG[4]
+ Tile_X6Y7_LUT4AB/N2BEG[5] Tile_X6Y7_LUT4AB/N2BEG[6] Tile_X6Y7_LUT4AB/N2BEG[7] Tile_X6Y6_LUT4AB/N2END[0]
+ Tile_X6Y6_LUT4AB/N2END[1] Tile_X6Y6_LUT4AB/N2END[2] Tile_X6Y6_LUT4AB/N2END[3] Tile_X6Y6_LUT4AB/N2END[4]
+ Tile_X6Y6_LUT4AB/N2END[5] Tile_X6Y6_LUT4AB/N2END[6] Tile_X6Y6_LUT4AB/N2END[7] Tile_X6Y7_LUT4AB/N2END[0]
+ Tile_X6Y7_LUT4AB/N2END[1] Tile_X6Y7_LUT4AB/N2END[2] Tile_X6Y7_LUT4AB/N2END[3] Tile_X6Y7_LUT4AB/N2END[4]
+ Tile_X6Y7_LUT4AB/N2END[5] Tile_X6Y7_LUT4AB/N2END[6] Tile_X6Y7_LUT4AB/N2END[7] Tile_X6Y8_LUT4AB/N2BEG[0]
+ Tile_X6Y8_LUT4AB/N2BEG[1] Tile_X6Y8_LUT4AB/N2BEG[2] Tile_X6Y8_LUT4AB/N2BEG[3] Tile_X6Y8_LUT4AB/N2BEG[4]
+ Tile_X6Y8_LUT4AB/N2BEG[5] Tile_X6Y8_LUT4AB/N2BEG[6] Tile_X6Y8_LUT4AB/N2BEG[7] Tile_X6Y7_LUT4AB/N4BEG[0]
+ Tile_X6Y7_LUT4AB/N4BEG[10] Tile_X6Y7_LUT4AB/N4BEG[11] Tile_X6Y7_LUT4AB/N4BEG[12]
+ Tile_X6Y7_LUT4AB/N4BEG[13] Tile_X6Y7_LUT4AB/N4BEG[14] Tile_X6Y7_LUT4AB/N4BEG[15]
+ Tile_X6Y7_LUT4AB/N4BEG[1] Tile_X6Y7_LUT4AB/N4BEG[2] Tile_X6Y7_LUT4AB/N4BEG[3] Tile_X6Y7_LUT4AB/N4BEG[4]
+ Tile_X6Y7_LUT4AB/N4BEG[5] Tile_X6Y7_LUT4AB/N4BEG[6] Tile_X6Y7_LUT4AB/N4BEG[7] Tile_X6Y7_LUT4AB/N4BEG[8]
+ Tile_X6Y7_LUT4AB/N4BEG[9] Tile_X6Y8_LUT4AB/N4BEG[0] Tile_X6Y8_LUT4AB/N4BEG[10] Tile_X6Y8_LUT4AB/N4BEG[11]
+ Tile_X6Y8_LUT4AB/N4BEG[12] Tile_X6Y8_LUT4AB/N4BEG[13] Tile_X6Y8_LUT4AB/N4BEG[14]
+ Tile_X6Y8_LUT4AB/N4BEG[15] Tile_X6Y8_LUT4AB/N4BEG[1] Tile_X6Y8_LUT4AB/N4BEG[2] Tile_X6Y8_LUT4AB/N4BEG[3]
+ Tile_X6Y8_LUT4AB/N4BEG[4] Tile_X6Y8_LUT4AB/N4BEG[5] Tile_X6Y8_LUT4AB/N4BEG[6] Tile_X6Y8_LUT4AB/N4BEG[7]
+ Tile_X6Y8_LUT4AB/N4BEG[8] Tile_X6Y8_LUT4AB/N4BEG[9] Tile_X6Y7_LUT4AB/NN4BEG[0] Tile_X6Y7_LUT4AB/NN4BEG[10]
+ Tile_X6Y7_LUT4AB/NN4BEG[11] Tile_X6Y7_LUT4AB/NN4BEG[12] Tile_X6Y7_LUT4AB/NN4BEG[13]
+ Tile_X6Y7_LUT4AB/NN4BEG[14] Tile_X6Y7_LUT4AB/NN4BEG[15] Tile_X6Y7_LUT4AB/NN4BEG[1]
+ Tile_X6Y7_LUT4AB/NN4BEG[2] Tile_X6Y7_LUT4AB/NN4BEG[3] Tile_X6Y7_LUT4AB/NN4BEG[4]
+ Tile_X6Y7_LUT4AB/NN4BEG[5] Tile_X6Y7_LUT4AB/NN4BEG[6] Tile_X6Y7_LUT4AB/NN4BEG[7]
+ Tile_X6Y7_LUT4AB/NN4BEG[8] Tile_X6Y7_LUT4AB/NN4BEG[9] Tile_X6Y8_LUT4AB/NN4BEG[0]
+ Tile_X6Y8_LUT4AB/NN4BEG[10] Tile_X6Y8_LUT4AB/NN4BEG[11] Tile_X6Y8_LUT4AB/NN4BEG[12]
+ Tile_X6Y8_LUT4AB/NN4BEG[13] Tile_X6Y8_LUT4AB/NN4BEG[14] Tile_X6Y8_LUT4AB/NN4BEG[15]
+ Tile_X6Y8_LUT4AB/NN4BEG[1] Tile_X6Y8_LUT4AB/NN4BEG[2] Tile_X6Y8_LUT4AB/NN4BEG[3]
+ Tile_X6Y8_LUT4AB/NN4BEG[4] Tile_X6Y8_LUT4AB/NN4BEG[5] Tile_X6Y8_LUT4AB/NN4BEG[6]
+ Tile_X6Y8_LUT4AB/NN4BEG[7] Tile_X6Y8_LUT4AB/NN4BEG[8] Tile_X6Y8_LUT4AB/NN4BEG[9]
+ Tile_X6Y8_LUT4AB/S1END[0] Tile_X6Y8_LUT4AB/S1END[1] Tile_X6Y8_LUT4AB/S1END[2] Tile_X6Y8_LUT4AB/S1END[3]
+ Tile_X6Y7_LUT4AB/S1END[0] Tile_X6Y7_LUT4AB/S1END[1] Tile_X6Y7_LUT4AB/S1END[2] Tile_X6Y7_LUT4AB/S1END[3]
+ Tile_X6Y8_LUT4AB/S2MID[0] Tile_X6Y8_LUT4AB/S2MID[1] Tile_X6Y8_LUT4AB/S2MID[2] Tile_X6Y8_LUT4AB/S2MID[3]
+ Tile_X6Y8_LUT4AB/S2MID[4] Tile_X6Y8_LUT4AB/S2MID[5] Tile_X6Y8_LUT4AB/S2MID[6] Tile_X6Y8_LUT4AB/S2MID[7]
+ Tile_X6Y8_LUT4AB/S2END[0] Tile_X6Y8_LUT4AB/S2END[1] Tile_X6Y8_LUT4AB/S2END[2] Tile_X6Y8_LUT4AB/S2END[3]
+ Tile_X6Y8_LUT4AB/S2END[4] Tile_X6Y8_LUT4AB/S2END[5] Tile_X6Y8_LUT4AB/S2END[6] Tile_X6Y8_LUT4AB/S2END[7]
+ Tile_X6Y7_LUT4AB/S2END[0] Tile_X6Y7_LUT4AB/S2END[1] Tile_X6Y7_LUT4AB/S2END[2] Tile_X6Y7_LUT4AB/S2END[3]
+ Tile_X6Y7_LUT4AB/S2END[4] Tile_X6Y7_LUT4AB/S2END[5] Tile_X6Y7_LUT4AB/S2END[6] Tile_X6Y7_LUT4AB/S2END[7]
+ Tile_X6Y7_LUT4AB/S2MID[0] Tile_X6Y7_LUT4AB/S2MID[1] Tile_X6Y7_LUT4AB/S2MID[2] Tile_X6Y7_LUT4AB/S2MID[3]
+ Tile_X6Y7_LUT4AB/S2MID[4] Tile_X6Y7_LUT4AB/S2MID[5] Tile_X6Y7_LUT4AB/S2MID[6] Tile_X6Y7_LUT4AB/S2MID[7]
+ Tile_X6Y8_LUT4AB/S4END[0] Tile_X6Y8_LUT4AB/S4END[10] Tile_X6Y8_LUT4AB/S4END[11]
+ Tile_X6Y8_LUT4AB/S4END[12] Tile_X6Y8_LUT4AB/S4END[13] Tile_X6Y8_LUT4AB/S4END[14]
+ Tile_X6Y8_LUT4AB/S4END[15] Tile_X6Y8_LUT4AB/S4END[1] Tile_X6Y8_LUT4AB/S4END[2] Tile_X6Y8_LUT4AB/S4END[3]
+ Tile_X6Y8_LUT4AB/S4END[4] Tile_X6Y8_LUT4AB/S4END[5] Tile_X6Y8_LUT4AB/S4END[6] Tile_X6Y8_LUT4AB/S4END[7]
+ Tile_X6Y8_LUT4AB/S4END[8] Tile_X6Y8_LUT4AB/S4END[9] Tile_X6Y7_LUT4AB/S4END[0] Tile_X6Y7_LUT4AB/S4END[10]
+ Tile_X6Y7_LUT4AB/S4END[11] Tile_X6Y7_LUT4AB/S4END[12] Tile_X6Y7_LUT4AB/S4END[13]
+ Tile_X6Y7_LUT4AB/S4END[14] Tile_X6Y7_LUT4AB/S4END[15] Tile_X6Y7_LUT4AB/S4END[1]
+ Tile_X6Y7_LUT4AB/S4END[2] Tile_X6Y7_LUT4AB/S4END[3] Tile_X6Y7_LUT4AB/S4END[4] Tile_X6Y7_LUT4AB/S4END[5]
+ Tile_X6Y7_LUT4AB/S4END[6] Tile_X6Y7_LUT4AB/S4END[7] Tile_X6Y7_LUT4AB/S4END[8] Tile_X6Y7_LUT4AB/S4END[9]
+ Tile_X6Y8_LUT4AB/SS4END[0] Tile_X6Y8_LUT4AB/SS4END[10] Tile_X6Y8_LUT4AB/SS4END[11]
+ Tile_X6Y8_LUT4AB/SS4END[12] Tile_X6Y8_LUT4AB/SS4END[13] Tile_X6Y8_LUT4AB/SS4END[14]
+ Tile_X6Y8_LUT4AB/SS4END[15] Tile_X6Y8_LUT4AB/SS4END[1] Tile_X6Y8_LUT4AB/SS4END[2]
+ Tile_X6Y8_LUT4AB/SS4END[3] Tile_X6Y8_LUT4AB/SS4END[4] Tile_X6Y8_LUT4AB/SS4END[5]
+ Tile_X6Y8_LUT4AB/SS4END[6] Tile_X6Y8_LUT4AB/SS4END[7] Tile_X6Y8_LUT4AB/SS4END[8]
+ Tile_X6Y8_LUT4AB/SS4END[9] Tile_X6Y7_LUT4AB/SS4END[0] Tile_X6Y7_LUT4AB/SS4END[10]
+ Tile_X6Y7_LUT4AB/SS4END[11] Tile_X6Y7_LUT4AB/SS4END[12] Tile_X6Y7_LUT4AB/SS4END[13]
+ Tile_X6Y7_LUT4AB/SS4END[14] Tile_X6Y7_LUT4AB/SS4END[15] Tile_X6Y7_LUT4AB/SS4END[1]
+ Tile_X6Y7_LUT4AB/SS4END[2] Tile_X6Y7_LUT4AB/SS4END[3] Tile_X6Y7_LUT4AB/SS4END[4]
+ Tile_X6Y7_LUT4AB/SS4END[5] Tile_X6Y7_LUT4AB/SS4END[6] Tile_X6Y7_LUT4AB/SS4END[7]
+ Tile_X6Y7_LUT4AB/SS4END[8] Tile_X6Y7_LUT4AB/SS4END[9] Tile_X6Y7_LUT4AB/UserCLK Tile_X6Y6_LUT4AB/UserCLK
+ VGND VPWR Tile_X6Y7_LUT4AB/W1BEG[0] Tile_X6Y7_LUT4AB/W1BEG[1] Tile_X6Y7_LUT4AB/W1BEG[2]
+ Tile_X6Y7_LUT4AB/W1BEG[3] Tile_X6Y7_LUT4AB/W1END[0] Tile_X6Y7_LUT4AB/W1END[1] Tile_X6Y7_LUT4AB/W1END[2]
+ Tile_X6Y7_LUT4AB/W1END[3] Tile_X6Y7_LUT4AB/W2BEG[0] Tile_X6Y7_LUT4AB/W2BEG[1] Tile_X6Y7_LUT4AB/W2BEG[2]
+ Tile_X6Y7_LUT4AB/W2BEG[3] Tile_X6Y7_LUT4AB/W2BEG[4] Tile_X6Y7_LUT4AB/W2BEG[5] Tile_X6Y7_LUT4AB/W2BEG[6]
+ Tile_X6Y7_LUT4AB/W2BEG[7] Tile_X5Y7_LUT4AB/W2END[0] Tile_X5Y7_LUT4AB/W2END[1] Tile_X5Y7_LUT4AB/W2END[2]
+ Tile_X5Y7_LUT4AB/W2END[3] Tile_X5Y7_LUT4AB/W2END[4] Tile_X5Y7_LUT4AB/W2END[5] Tile_X5Y7_LUT4AB/W2END[6]
+ Tile_X5Y7_LUT4AB/W2END[7] Tile_X6Y7_LUT4AB/W2END[0] Tile_X6Y7_LUT4AB/W2END[1] Tile_X6Y7_LUT4AB/W2END[2]
+ Tile_X6Y7_LUT4AB/W2END[3] Tile_X6Y7_LUT4AB/W2END[4] Tile_X6Y7_LUT4AB/W2END[5] Tile_X6Y7_LUT4AB/W2END[6]
+ Tile_X6Y7_LUT4AB/W2END[7] Tile_X6Y7_LUT4AB/W2MID[0] Tile_X6Y7_LUT4AB/W2MID[1] Tile_X6Y7_LUT4AB/W2MID[2]
+ Tile_X6Y7_LUT4AB/W2MID[3] Tile_X6Y7_LUT4AB/W2MID[4] Tile_X6Y7_LUT4AB/W2MID[5] Tile_X6Y7_LUT4AB/W2MID[6]
+ Tile_X6Y7_LUT4AB/W2MID[7] Tile_X6Y7_LUT4AB/W6BEG[0] Tile_X6Y7_LUT4AB/W6BEG[10] Tile_X6Y7_LUT4AB/W6BEG[11]
+ Tile_X6Y7_LUT4AB/W6BEG[1] Tile_X6Y7_LUT4AB/W6BEG[2] Tile_X6Y7_LUT4AB/W6BEG[3] Tile_X6Y7_LUT4AB/W6BEG[4]
+ Tile_X6Y7_LUT4AB/W6BEG[5] Tile_X6Y7_LUT4AB/W6BEG[6] Tile_X6Y7_LUT4AB/W6BEG[7] Tile_X6Y7_LUT4AB/W6BEG[8]
+ Tile_X6Y7_LUT4AB/W6BEG[9] Tile_X6Y7_LUT4AB/W6END[0] Tile_X6Y7_LUT4AB/W6END[10] Tile_X6Y7_LUT4AB/W6END[11]
+ Tile_X6Y7_LUT4AB/W6END[1] Tile_X6Y7_LUT4AB/W6END[2] Tile_X6Y7_LUT4AB/W6END[3] Tile_X6Y7_LUT4AB/W6END[4]
+ Tile_X6Y7_LUT4AB/W6END[5] Tile_X6Y7_LUT4AB/W6END[6] Tile_X6Y7_LUT4AB/W6END[7] Tile_X6Y7_LUT4AB/W6END[8]
+ Tile_X6Y7_LUT4AB/W6END[9] Tile_X6Y7_LUT4AB/WW4BEG[0] Tile_X6Y7_LUT4AB/WW4BEG[10]
+ Tile_X6Y7_LUT4AB/WW4BEG[11] Tile_X6Y7_LUT4AB/WW4BEG[12] Tile_X6Y7_LUT4AB/WW4BEG[13]
+ Tile_X6Y7_LUT4AB/WW4BEG[14] Tile_X6Y7_LUT4AB/WW4BEG[15] Tile_X6Y7_LUT4AB/WW4BEG[1]
+ Tile_X6Y7_LUT4AB/WW4BEG[2] Tile_X6Y7_LUT4AB/WW4BEG[3] Tile_X6Y7_LUT4AB/WW4BEG[4]
+ Tile_X6Y7_LUT4AB/WW4BEG[5] Tile_X6Y7_LUT4AB/WW4BEG[6] Tile_X6Y7_LUT4AB/WW4BEG[7]
+ Tile_X6Y7_LUT4AB/WW4BEG[8] Tile_X6Y7_LUT4AB/WW4BEG[9] Tile_X6Y7_LUT4AB/WW4END[0]
+ Tile_X6Y7_LUT4AB/WW4END[10] Tile_X6Y7_LUT4AB/WW4END[11] Tile_X6Y7_LUT4AB/WW4END[12]
+ Tile_X6Y7_LUT4AB/WW4END[13] Tile_X6Y7_LUT4AB/WW4END[14] Tile_X6Y7_LUT4AB/WW4END[15]
+ Tile_X6Y7_LUT4AB/WW4END[1] Tile_X6Y7_LUT4AB/WW4END[2] Tile_X6Y7_LUT4AB/WW4END[3]
+ Tile_X6Y7_LUT4AB/WW4END[4] Tile_X6Y7_LUT4AB/WW4END[5] Tile_X6Y7_LUT4AB/WW4END[6]
+ Tile_X6Y7_LUT4AB/WW4END[7] Tile_X6Y7_LUT4AB/WW4END[8] Tile_X6Y7_LUT4AB/WW4END[9]
+ LUT4AB
XTile_X3Y2_LUT4AB Tile_X3Y3_LUT4AB/Co Tile_X3Y2_LUT4AB/Co Tile_X3Y2_LUT4AB/E1BEG[0]
+ Tile_X3Y2_LUT4AB/E1BEG[1] Tile_X3Y2_LUT4AB/E1BEG[2] Tile_X3Y2_LUT4AB/E1BEG[3] Tile_X3Y2_LUT4AB/E1END[0]
+ Tile_X3Y2_LUT4AB/E1END[1] Tile_X3Y2_LUT4AB/E1END[2] Tile_X3Y2_LUT4AB/E1END[3] Tile_X3Y2_LUT4AB/E2BEG[0]
+ Tile_X3Y2_LUT4AB/E2BEG[1] Tile_X3Y2_LUT4AB/E2BEG[2] Tile_X3Y2_LUT4AB/E2BEG[3] Tile_X3Y2_LUT4AB/E2BEG[4]
+ Tile_X3Y2_LUT4AB/E2BEG[5] Tile_X3Y2_LUT4AB/E2BEG[6] Tile_X3Y2_LUT4AB/E2BEG[7] Tile_X4Y2_RegFile/E2END[0]
+ Tile_X4Y2_RegFile/E2END[1] Tile_X4Y2_RegFile/E2END[2] Tile_X4Y2_RegFile/E2END[3]
+ Tile_X4Y2_RegFile/E2END[4] Tile_X4Y2_RegFile/E2END[5] Tile_X4Y2_RegFile/E2END[6]
+ Tile_X4Y2_RegFile/E2END[7] Tile_X3Y2_LUT4AB/E2END[0] Tile_X3Y2_LUT4AB/E2END[1] Tile_X3Y2_LUT4AB/E2END[2]
+ Tile_X3Y2_LUT4AB/E2END[3] Tile_X3Y2_LUT4AB/E2END[4] Tile_X3Y2_LUT4AB/E2END[5] Tile_X3Y2_LUT4AB/E2END[6]
+ Tile_X3Y2_LUT4AB/E2END[7] Tile_X3Y2_LUT4AB/E2MID[0] Tile_X3Y2_LUT4AB/E2MID[1] Tile_X3Y2_LUT4AB/E2MID[2]
+ Tile_X3Y2_LUT4AB/E2MID[3] Tile_X3Y2_LUT4AB/E2MID[4] Tile_X3Y2_LUT4AB/E2MID[5] Tile_X3Y2_LUT4AB/E2MID[6]
+ Tile_X3Y2_LUT4AB/E2MID[7] Tile_X3Y2_LUT4AB/E6BEG[0] Tile_X3Y2_LUT4AB/E6BEG[10] Tile_X3Y2_LUT4AB/E6BEG[11]
+ Tile_X3Y2_LUT4AB/E6BEG[1] Tile_X3Y2_LUT4AB/E6BEG[2] Tile_X3Y2_LUT4AB/E6BEG[3] Tile_X3Y2_LUT4AB/E6BEG[4]
+ Tile_X3Y2_LUT4AB/E6BEG[5] Tile_X3Y2_LUT4AB/E6BEG[6] Tile_X3Y2_LUT4AB/E6BEG[7] Tile_X3Y2_LUT4AB/E6BEG[8]
+ Tile_X3Y2_LUT4AB/E6BEG[9] Tile_X3Y2_LUT4AB/E6END[0] Tile_X3Y2_LUT4AB/E6END[10] Tile_X3Y2_LUT4AB/E6END[11]
+ Tile_X3Y2_LUT4AB/E6END[1] Tile_X3Y2_LUT4AB/E6END[2] Tile_X3Y2_LUT4AB/E6END[3] Tile_X3Y2_LUT4AB/E6END[4]
+ Tile_X3Y2_LUT4AB/E6END[5] Tile_X3Y2_LUT4AB/E6END[6] Tile_X3Y2_LUT4AB/E6END[7] Tile_X3Y2_LUT4AB/E6END[8]
+ Tile_X3Y2_LUT4AB/E6END[9] Tile_X3Y2_LUT4AB/EE4BEG[0] Tile_X3Y2_LUT4AB/EE4BEG[10]
+ Tile_X3Y2_LUT4AB/EE4BEG[11] Tile_X3Y2_LUT4AB/EE4BEG[12] Tile_X3Y2_LUT4AB/EE4BEG[13]
+ Tile_X3Y2_LUT4AB/EE4BEG[14] Tile_X3Y2_LUT4AB/EE4BEG[15] Tile_X3Y2_LUT4AB/EE4BEG[1]
+ Tile_X3Y2_LUT4AB/EE4BEG[2] Tile_X3Y2_LUT4AB/EE4BEG[3] Tile_X3Y2_LUT4AB/EE4BEG[4]
+ Tile_X3Y2_LUT4AB/EE4BEG[5] Tile_X3Y2_LUT4AB/EE4BEG[6] Tile_X3Y2_LUT4AB/EE4BEG[7]
+ Tile_X3Y2_LUT4AB/EE4BEG[8] Tile_X3Y2_LUT4AB/EE4BEG[9] Tile_X3Y2_LUT4AB/EE4END[0]
+ Tile_X3Y2_LUT4AB/EE4END[10] Tile_X3Y2_LUT4AB/EE4END[11] Tile_X3Y2_LUT4AB/EE4END[12]
+ Tile_X3Y2_LUT4AB/EE4END[13] Tile_X3Y2_LUT4AB/EE4END[14] Tile_X3Y2_LUT4AB/EE4END[15]
+ Tile_X3Y2_LUT4AB/EE4END[1] Tile_X3Y2_LUT4AB/EE4END[2] Tile_X3Y2_LUT4AB/EE4END[3]
+ Tile_X3Y2_LUT4AB/EE4END[4] Tile_X3Y2_LUT4AB/EE4END[5] Tile_X3Y2_LUT4AB/EE4END[6]
+ Tile_X3Y2_LUT4AB/EE4END[7] Tile_X3Y2_LUT4AB/EE4END[8] Tile_X3Y2_LUT4AB/EE4END[9]
+ Tile_X3Y2_LUT4AB/FrameData[0] Tile_X3Y2_LUT4AB/FrameData[10] Tile_X3Y2_LUT4AB/FrameData[11]
+ Tile_X3Y2_LUT4AB/FrameData[12] Tile_X3Y2_LUT4AB/FrameData[13] Tile_X3Y2_LUT4AB/FrameData[14]
+ Tile_X3Y2_LUT4AB/FrameData[15] Tile_X3Y2_LUT4AB/FrameData[16] Tile_X3Y2_LUT4AB/FrameData[17]
+ Tile_X3Y2_LUT4AB/FrameData[18] Tile_X3Y2_LUT4AB/FrameData[19] Tile_X3Y2_LUT4AB/FrameData[1]
+ Tile_X3Y2_LUT4AB/FrameData[20] Tile_X3Y2_LUT4AB/FrameData[21] Tile_X3Y2_LUT4AB/FrameData[22]
+ Tile_X3Y2_LUT4AB/FrameData[23] Tile_X3Y2_LUT4AB/FrameData[24] Tile_X3Y2_LUT4AB/FrameData[25]
+ Tile_X3Y2_LUT4AB/FrameData[26] Tile_X3Y2_LUT4AB/FrameData[27] Tile_X3Y2_LUT4AB/FrameData[28]
+ Tile_X3Y2_LUT4AB/FrameData[29] Tile_X3Y2_LUT4AB/FrameData[2] Tile_X3Y2_LUT4AB/FrameData[30]
+ Tile_X3Y2_LUT4AB/FrameData[31] Tile_X3Y2_LUT4AB/FrameData[3] Tile_X3Y2_LUT4AB/FrameData[4]
+ Tile_X3Y2_LUT4AB/FrameData[5] Tile_X3Y2_LUT4AB/FrameData[6] Tile_X3Y2_LUT4AB/FrameData[7]
+ Tile_X3Y2_LUT4AB/FrameData[8] Tile_X3Y2_LUT4AB/FrameData[9] Tile_X4Y2_RegFile/FrameData[0]
+ Tile_X4Y2_RegFile/FrameData[10] Tile_X4Y2_RegFile/FrameData[11] Tile_X4Y2_RegFile/FrameData[12]
+ Tile_X4Y2_RegFile/FrameData[13] Tile_X4Y2_RegFile/FrameData[14] Tile_X4Y2_RegFile/FrameData[15]
+ Tile_X4Y2_RegFile/FrameData[16] Tile_X4Y2_RegFile/FrameData[17] Tile_X4Y2_RegFile/FrameData[18]
+ Tile_X4Y2_RegFile/FrameData[19] Tile_X4Y2_RegFile/FrameData[1] Tile_X4Y2_RegFile/FrameData[20]
+ Tile_X4Y2_RegFile/FrameData[21] Tile_X4Y2_RegFile/FrameData[22] Tile_X4Y2_RegFile/FrameData[23]
+ Tile_X4Y2_RegFile/FrameData[24] Tile_X4Y2_RegFile/FrameData[25] Tile_X4Y2_RegFile/FrameData[26]
+ Tile_X4Y2_RegFile/FrameData[27] Tile_X4Y2_RegFile/FrameData[28] Tile_X4Y2_RegFile/FrameData[29]
+ Tile_X4Y2_RegFile/FrameData[2] Tile_X4Y2_RegFile/FrameData[30] Tile_X4Y2_RegFile/FrameData[31]
+ Tile_X4Y2_RegFile/FrameData[3] Tile_X4Y2_RegFile/FrameData[4] Tile_X4Y2_RegFile/FrameData[5]
+ Tile_X4Y2_RegFile/FrameData[6] Tile_X4Y2_RegFile/FrameData[7] Tile_X4Y2_RegFile/FrameData[8]
+ Tile_X4Y2_RegFile/FrameData[9] Tile_X3Y2_LUT4AB/FrameStrobe[0] Tile_X3Y2_LUT4AB/FrameStrobe[10]
+ Tile_X3Y2_LUT4AB/FrameStrobe[11] Tile_X3Y2_LUT4AB/FrameStrobe[12] Tile_X3Y2_LUT4AB/FrameStrobe[13]
+ Tile_X3Y2_LUT4AB/FrameStrobe[14] Tile_X3Y2_LUT4AB/FrameStrobe[15] Tile_X3Y2_LUT4AB/FrameStrobe[16]
+ Tile_X3Y2_LUT4AB/FrameStrobe[17] Tile_X3Y2_LUT4AB/FrameStrobe[18] Tile_X3Y2_LUT4AB/FrameStrobe[19]
+ Tile_X3Y2_LUT4AB/FrameStrobe[1] Tile_X3Y2_LUT4AB/FrameStrobe[2] Tile_X3Y2_LUT4AB/FrameStrobe[3]
+ Tile_X3Y2_LUT4AB/FrameStrobe[4] Tile_X3Y2_LUT4AB/FrameStrobe[5] Tile_X3Y2_LUT4AB/FrameStrobe[6]
+ Tile_X3Y2_LUT4AB/FrameStrobe[7] Tile_X3Y2_LUT4AB/FrameStrobe[8] Tile_X3Y2_LUT4AB/FrameStrobe[9]
+ Tile_X3Y1_LUT4AB/FrameStrobe[0] Tile_X3Y1_LUT4AB/FrameStrobe[10] Tile_X3Y1_LUT4AB/FrameStrobe[11]
+ Tile_X3Y1_LUT4AB/FrameStrobe[12] Tile_X3Y1_LUT4AB/FrameStrobe[13] Tile_X3Y1_LUT4AB/FrameStrobe[14]
+ Tile_X3Y1_LUT4AB/FrameStrobe[15] Tile_X3Y1_LUT4AB/FrameStrobe[16] Tile_X3Y1_LUT4AB/FrameStrobe[17]
+ Tile_X3Y1_LUT4AB/FrameStrobe[18] Tile_X3Y1_LUT4AB/FrameStrobe[19] Tile_X3Y1_LUT4AB/FrameStrobe[1]
+ Tile_X3Y1_LUT4AB/FrameStrobe[2] Tile_X3Y1_LUT4AB/FrameStrobe[3] Tile_X3Y1_LUT4AB/FrameStrobe[4]
+ Tile_X3Y1_LUT4AB/FrameStrobe[5] Tile_X3Y1_LUT4AB/FrameStrobe[6] Tile_X3Y1_LUT4AB/FrameStrobe[7]
+ Tile_X3Y1_LUT4AB/FrameStrobe[8] Tile_X3Y1_LUT4AB/FrameStrobe[9] Tile_X3Y2_LUT4AB/N1BEG[0]
+ Tile_X3Y2_LUT4AB/N1BEG[1] Tile_X3Y2_LUT4AB/N1BEG[2] Tile_X3Y2_LUT4AB/N1BEG[3] Tile_X3Y3_LUT4AB/N1BEG[0]
+ Tile_X3Y3_LUT4AB/N1BEG[1] Tile_X3Y3_LUT4AB/N1BEG[2] Tile_X3Y3_LUT4AB/N1BEG[3] Tile_X3Y2_LUT4AB/N2BEG[0]
+ Tile_X3Y2_LUT4AB/N2BEG[1] Tile_X3Y2_LUT4AB/N2BEG[2] Tile_X3Y2_LUT4AB/N2BEG[3] Tile_X3Y2_LUT4AB/N2BEG[4]
+ Tile_X3Y2_LUT4AB/N2BEG[5] Tile_X3Y2_LUT4AB/N2BEG[6] Tile_X3Y2_LUT4AB/N2BEG[7] Tile_X3Y1_LUT4AB/N2END[0]
+ Tile_X3Y1_LUT4AB/N2END[1] Tile_X3Y1_LUT4AB/N2END[2] Tile_X3Y1_LUT4AB/N2END[3] Tile_X3Y1_LUT4AB/N2END[4]
+ Tile_X3Y1_LUT4AB/N2END[5] Tile_X3Y1_LUT4AB/N2END[6] Tile_X3Y1_LUT4AB/N2END[7] Tile_X3Y2_LUT4AB/N2END[0]
+ Tile_X3Y2_LUT4AB/N2END[1] Tile_X3Y2_LUT4AB/N2END[2] Tile_X3Y2_LUT4AB/N2END[3] Tile_X3Y2_LUT4AB/N2END[4]
+ Tile_X3Y2_LUT4AB/N2END[5] Tile_X3Y2_LUT4AB/N2END[6] Tile_X3Y2_LUT4AB/N2END[7] Tile_X3Y3_LUT4AB/N2BEG[0]
+ Tile_X3Y3_LUT4AB/N2BEG[1] Tile_X3Y3_LUT4AB/N2BEG[2] Tile_X3Y3_LUT4AB/N2BEG[3] Tile_X3Y3_LUT4AB/N2BEG[4]
+ Tile_X3Y3_LUT4AB/N2BEG[5] Tile_X3Y3_LUT4AB/N2BEG[6] Tile_X3Y3_LUT4AB/N2BEG[7] Tile_X3Y2_LUT4AB/N4BEG[0]
+ Tile_X3Y2_LUT4AB/N4BEG[10] Tile_X3Y2_LUT4AB/N4BEG[11] Tile_X3Y2_LUT4AB/N4BEG[12]
+ Tile_X3Y2_LUT4AB/N4BEG[13] Tile_X3Y2_LUT4AB/N4BEG[14] Tile_X3Y2_LUT4AB/N4BEG[15]
+ Tile_X3Y2_LUT4AB/N4BEG[1] Tile_X3Y2_LUT4AB/N4BEG[2] Tile_X3Y2_LUT4AB/N4BEG[3] Tile_X3Y2_LUT4AB/N4BEG[4]
+ Tile_X3Y2_LUT4AB/N4BEG[5] Tile_X3Y2_LUT4AB/N4BEG[6] Tile_X3Y2_LUT4AB/N4BEG[7] Tile_X3Y2_LUT4AB/N4BEG[8]
+ Tile_X3Y2_LUT4AB/N4BEG[9] Tile_X3Y3_LUT4AB/N4BEG[0] Tile_X3Y3_LUT4AB/N4BEG[10] Tile_X3Y3_LUT4AB/N4BEG[11]
+ Tile_X3Y3_LUT4AB/N4BEG[12] Tile_X3Y3_LUT4AB/N4BEG[13] Tile_X3Y3_LUT4AB/N4BEG[14]
+ Tile_X3Y3_LUT4AB/N4BEG[15] Tile_X3Y3_LUT4AB/N4BEG[1] Tile_X3Y3_LUT4AB/N4BEG[2] Tile_X3Y3_LUT4AB/N4BEG[3]
+ Tile_X3Y3_LUT4AB/N4BEG[4] Tile_X3Y3_LUT4AB/N4BEG[5] Tile_X3Y3_LUT4AB/N4BEG[6] Tile_X3Y3_LUT4AB/N4BEG[7]
+ Tile_X3Y3_LUT4AB/N4BEG[8] Tile_X3Y3_LUT4AB/N4BEG[9] Tile_X3Y2_LUT4AB/NN4BEG[0] Tile_X3Y2_LUT4AB/NN4BEG[10]
+ Tile_X3Y2_LUT4AB/NN4BEG[11] Tile_X3Y2_LUT4AB/NN4BEG[12] Tile_X3Y2_LUT4AB/NN4BEG[13]
+ Tile_X3Y2_LUT4AB/NN4BEG[14] Tile_X3Y2_LUT4AB/NN4BEG[15] Tile_X3Y2_LUT4AB/NN4BEG[1]
+ Tile_X3Y2_LUT4AB/NN4BEG[2] Tile_X3Y2_LUT4AB/NN4BEG[3] Tile_X3Y2_LUT4AB/NN4BEG[4]
+ Tile_X3Y2_LUT4AB/NN4BEG[5] Tile_X3Y2_LUT4AB/NN4BEG[6] Tile_X3Y2_LUT4AB/NN4BEG[7]
+ Tile_X3Y2_LUT4AB/NN4BEG[8] Tile_X3Y2_LUT4AB/NN4BEG[9] Tile_X3Y3_LUT4AB/NN4BEG[0]
+ Tile_X3Y3_LUT4AB/NN4BEG[10] Tile_X3Y3_LUT4AB/NN4BEG[11] Tile_X3Y3_LUT4AB/NN4BEG[12]
+ Tile_X3Y3_LUT4AB/NN4BEG[13] Tile_X3Y3_LUT4AB/NN4BEG[14] Tile_X3Y3_LUT4AB/NN4BEG[15]
+ Tile_X3Y3_LUT4AB/NN4BEG[1] Tile_X3Y3_LUT4AB/NN4BEG[2] Tile_X3Y3_LUT4AB/NN4BEG[3]
+ Tile_X3Y3_LUT4AB/NN4BEG[4] Tile_X3Y3_LUT4AB/NN4BEG[5] Tile_X3Y3_LUT4AB/NN4BEG[6]
+ Tile_X3Y3_LUT4AB/NN4BEG[7] Tile_X3Y3_LUT4AB/NN4BEG[8] Tile_X3Y3_LUT4AB/NN4BEG[9]
+ Tile_X3Y3_LUT4AB/S1END[0] Tile_X3Y3_LUT4AB/S1END[1] Tile_X3Y3_LUT4AB/S1END[2] Tile_X3Y3_LUT4AB/S1END[3]
+ Tile_X3Y2_LUT4AB/S1END[0] Tile_X3Y2_LUT4AB/S1END[1] Tile_X3Y2_LUT4AB/S1END[2] Tile_X3Y2_LUT4AB/S1END[3]
+ Tile_X3Y3_LUT4AB/S2MID[0] Tile_X3Y3_LUT4AB/S2MID[1] Tile_X3Y3_LUT4AB/S2MID[2] Tile_X3Y3_LUT4AB/S2MID[3]
+ Tile_X3Y3_LUT4AB/S2MID[4] Tile_X3Y3_LUT4AB/S2MID[5] Tile_X3Y3_LUT4AB/S2MID[6] Tile_X3Y3_LUT4AB/S2MID[7]
+ Tile_X3Y3_LUT4AB/S2END[0] Tile_X3Y3_LUT4AB/S2END[1] Tile_X3Y3_LUT4AB/S2END[2] Tile_X3Y3_LUT4AB/S2END[3]
+ Tile_X3Y3_LUT4AB/S2END[4] Tile_X3Y3_LUT4AB/S2END[5] Tile_X3Y3_LUT4AB/S2END[6] Tile_X3Y3_LUT4AB/S2END[7]
+ Tile_X3Y2_LUT4AB/S2END[0] Tile_X3Y2_LUT4AB/S2END[1] Tile_X3Y2_LUT4AB/S2END[2] Tile_X3Y2_LUT4AB/S2END[3]
+ Tile_X3Y2_LUT4AB/S2END[4] Tile_X3Y2_LUT4AB/S2END[5] Tile_X3Y2_LUT4AB/S2END[6] Tile_X3Y2_LUT4AB/S2END[7]
+ Tile_X3Y2_LUT4AB/S2MID[0] Tile_X3Y2_LUT4AB/S2MID[1] Tile_X3Y2_LUT4AB/S2MID[2] Tile_X3Y2_LUT4AB/S2MID[3]
+ Tile_X3Y2_LUT4AB/S2MID[4] Tile_X3Y2_LUT4AB/S2MID[5] Tile_X3Y2_LUT4AB/S2MID[6] Tile_X3Y2_LUT4AB/S2MID[7]
+ Tile_X3Y3_LUT4AB/S4END[0] Tile_X3Y3_LUT4AB/S4END[10] Tile_X3Y3_LUT4AB/S4END[11]
+ Tile_X3Y3_LUT4AB/S4END[12] Tile_X3Y3_LUT4AB/S4END[13] Tile_X3Y3_LUT4AB/S4END[14]
+ Tile_X3Y3_LUT4AB/S4END[15] Tile_X3Y3_LUT4AB/S4END[1] Tile_X3Y3_LUT4AB/S4END[2] Tile_X3Y3_LUT4AB/S4END[3]
+ Tile_X3Y3_LUT4AB/S4END[4] Tile_X3Y3_LUT4AB/S4END[5] Tile_X3Y3_LUT4AB/S4END[6] Tile_X3Y3_LUT4AB/S4END[7]
+ Tile_X3Y3_LUT4AB/S4END[8] Tile_X3Y3_LUT4AB/S4END[9] Tile_X3Y2_LUT4AB/S4END[0] Tile_X3Y2_LUT4AB/S4END[10]
+ Tile_X3Y2_LUT4AB/S4END[11] Tile_X3Y2_LUT4AB/S4END[12] Tile_X3Y2_LUT4AB/S4END[13]
+ Tile_X3Y2_LUT4AB/S4END[14] Tile_X3Y2_LUT4AB/S4END[15] Tile_X3Y2_LUT4AB/S4END[1]
+ Tile_X3Y2_LUT4AB/S4END[2] Tile_X3Y2_LUT4AB/S4END[3] Tile_X3Y2_LUT4AB/S4END[4] Tile_X3Y2_LUT4AB/S4END[5]
+ Tile_X3Y2_LUT4AB/S4END[6] Tile_X3Y2_LUT4AB/S4END[7] Tile_X3Y2_LUT4AB/S4END[8] Tile_X3Y2_LUT4AB/S4END[9]
+ Tile_X3Y3_LUT4AB/SS4END[0] Tile_X3Y3_LUT4AB/SS4END[10] Tile_X3Y3_LUT4AB/SS4END[11]
+ Tile_X3Y3_LUT4AB/SS4END[12] Tile_X3Y3_LUT4AB/SS4END[13] Tile_X3Y3_LUT4AB/SS4END[14]
+ Tile_X3Y3_LUT4AB/SS4END[15] Tile_X3Y3_LUT4AB/SS4END[1] Tile_X3Y3_LUT4AB/SS4END[2]
+ Tile_X3Y3_LUT4AB/SS4END[3] Tile_X3Y3_LUT4AB/SS4END[4] Tile_X3Y3_LUT4AB/SS4END[5]
+ Tile_X3Y3_LUT4AB/SS4END[6] Tile_X3Y3_LUT4AB/SS4END[7] Tile_X3Y3_LUT4AB/SS4END[8]
+ Tile_X3Y3_LUT4AB/SS4END[9] Tile_X3Y2_LUT4AB/SS4END[0] Tile_X3Y2_LUT4AB/SS4END[10]
+ Tile_X3Y2_LUT4AB/SS4END[11] Tile_X3Y2_LUT4AB/SS4END[12] Tile_X3Y2_LUT4AB/SS4END[13]
+ Tile_X3Y2_LUT4AB/SS4END[14] Tile_X3Y2_LUT4AB/SS4END[15] Tile_X3Y2_LUT4AB/SS4END[1]
+ Tile_X3Y2_LUT4AB/SS4END[2] Tile_X3Y2_LUT4AB/SS4END[3] Tile_X3Y2_LUT4AB/SS4END[4]
+ Tile_X3Y2_LUT4AB/SS4END[5] Tile_X3Y2_LUT4AB/SS4END[6] Tile_X3Y2_LUT4AB/SS4END[7]
+ Tile_X3Y2_LUT4AB/SS4END[8] Tile_X3Y2_LUT4AB/SS4END[9] Tile_X3Y2_LUT4AB/UserCLK Tile_X3Y1_LUT4AB/UserCLK
+ VGND VPWR Tile_X3Y2_LUT4AB/W1BEG[0] Tile_X3Y2_LUT4AB/W1BEG[1] Tile_X3Y2_LUT4AB/W1BEG[2]
+ Tile_X3Y2_LUT4AB/W1BEG[3] Tile_X3Y2_LUT4AB/W1END[0] Tile_X3Y2_LUT4AB/W1END[1] Tile_X3Y2_LUT4AB/W1END[2]
+ Tile_X3Y2_LUT4AB/W1END[3] Tile_X3Y2_LUT4AB/W2BEG[0] Tile_X3Y2_LUT4AB/W2BEG[1] Tile_X3Y2_LUT4AB/W2BEG[2]
+ Tile_X3Y2_LUT4AB/W2BEG[3] Tile_X3Y2_LUT4AB/W2BEG[4] Tile_X3Y2_LUT4AB/W2BEG[5] Tile_X3Y2_LUT4AB/W2BEG[6]
+ Tile_X3Y2_LUT4AB/W2BEG[7] Tile_X2Y2_LUT4AB/W2END[0] Tile_X2Y2_LUT4AB/W2END[1] Tile_X2Y2_LUT4AB/W2END[2]
+ Tile_X2Y2_LUT4AB/W2END[3] Tile_X2Y2_LUT4AB/W2END[4] Tile_X2Y2_LUT4AB/W2END[5] Tile_X2Y2_LUT4AB/W2END[6]
+ Tile_X2Y2_LUT4AB/W2END[7] Tile_X3Y2_LUT4AB/W2END[0] Tile_X3Y2_LUT4AB/W2END[1] Tile_X3Y2_LUT4AB/W2END[2]
+ Tile_X3Y2_LUT4AB/W2END[3] Tile_X3Y2_LUT4AB/W2END[4] Tile_X3Y2_LUT4AB/W2END[5] Tile_X3Y2_LUT4AB/W2END[6]
+ Tile_X3Y2_LUT4AB/W2END[7] Tile_X3Y2_LUT4AB/W2MID[0] Tile_X3Y2_LUT4AB/W2MID[1] Tile_X3Y2_LUT4AB/W2MID[2]
+ Tile_X3Y2_LUT4AB/W2MID[3] Tile_X3Y2_LUT4AB/W2MID[4] Tile_X3Y2_LUT4AB/W2MID[5] Tile_X3Y2_LUT4AB/W2MID[6]
+ Tile_X3Y2_LUT4AB/W2MID[7] Tile_X3Y2_LUT4AB/W6BEG[0] Tile_X3Y2_LUT4AB/W6BEG[10] Tile_X3Y2_LUT4AB/W6BEG[11]
+ Tile_X3Y2_LUT4AB/W6BEG[1] Tile_X3Y2_LUT4AB/W6BEG[2] Tile_X3Y2_LUT4AB/W6BEG[3] Tile_X3Y2_LUT4AB/W6BEG[4]
+ Tile_X3Y2_LUT4AB/W6BEG[5] Tile_X3Y2_LUT4AB/W6BEG[6] Tile_X3Y2_LUT4AB/W6BEG[7] Tile_X3Y2_LUT4AB/W6BEG[8]
+ Tile_X3Y2_LUT4AB/W6BEG[9] Tile_X3Y2_LUT4AB/W6END[0] Tile_X3Y2_LUT4AB/W6END[10] Tile_X3Y2_LUT4AB/W6END[11]
+ Tile_X3Y2_LUT4AB/W6END[1] Tile_X3Y2_LUT4AB/W6END[2] Tile_X3Y2_LUT4AB/W6END[3] Tile_X3Y2_LUT4AB/W6END[4]
+ Tile_X3Y2_LUT4AB/W6END[5] Tile_X3Y2_LUT4AB/W6END[6] Tile_X3Y2_LUT4AB/W6END[7] Tile_X3Y2_LUT4AB/W6END[8]
+ Tile_X3Y2_LUT4AB/W6END[9] Tile_X3Y2_LUT4AB/WW4BEG[0] Tile_X3Y2_LUT4AB/WW4BEG[10]
+ Tile_X3Y2_LUT4AB/WW4BEG[11] Tile_X3Y2_LUT4AB/WW4BEG[12] Tile_X3Y2_LUT4AB/WW4BEG[13]
+ Tile_X3Y2_LUT4AB/WW4BEG[14] Tile_X3Y2_LUT4AB/WW4BEG[15] Tile_X3Y2_LUT4AB/WW4BEG[1]
+ Tile_X3Y2_LUT4AB/WW4BEG[2] Tile_X3Y2_LUT4AB/WW4BEG[3] Tile_X3Y2_LUT4AB/WW4BEG[4]
+ Tile_X3Y2_LUT4AB/WW4BEG[5] Tile_X3Y2_LUT4AB/WW4BEG[6] Tile_X3Y2_LUT4AB/WW4BEG[7]
+ Tile_X3Y2_LUT4AB/WW4BEG[8] Tile_X3Y2_LUT4AB/WW4BEG[9] Tile_X3Y2_LUT4AB/WW4END[0]
+ Tile_X3Y2_LUT4AB/WW4END[10] Tile_X3Y2_LUT4AB/WW4END[11] Tile_X3Y2_LUT4AB/WW4END[12]
+ Tile_X3Y2_LUT4AB/WW4END[13] Tile_X3Y2_LUT4AB/WW4END[14] Tile_X3Y2_LUT4AB/WW4END[15]
+ Tile_X3Y2_LUT4AB/WW4END[1] Tile_X3Y2_LUT4AB/WW4END[2] Tile_X3Y2_LUT4AB/WW4END[3]
+ Tile_X3Y2_LUT4AB/WW4END[4] Tile_X3Y2_LUT4AB/WW4END[5] Tile_X3Y2_LUT4AB/WW4END[6]
+ Tile_X3Y2_LUT4AB/WW4END[7] Tile_X3Y2_LUT4AB/WW4END[8] Tile_X3Y2_LUT4AB/WW4END[9]
+ LUT4AB
XTile_X3Y15_S_CPU_IRQ Tile_X3Y15_CONFIGURED_top Tile_X3Y14_LUT4AB/Ci Tile_X3Y15_S_CPU_IRQ/FrameData[0]
+ Tile_X3Y15_S_CPU_IRQ/FrameData[10] Tile_X3Y15_S_CPU_IRQ/FrameData[11] Tile_X3Y15_S_CPU_IRQ/FrameData[12]
+ Tile_X3Y15_S_CPU_IRQ/FrameData[13] Tile_X3Y15_S_CPU_IRQ/FrameData[14] Tile_X3Y15_S_CPU_IRQ/FrameData[15]
+ Tile_X3Y15_S_CPU_IRQ/FrameData[16] Tile_X3Y15_S_CPU_IRQ/FrameData[17] Tile_X3Y15_S_CPU_IRQ/FrameData[18]
+ Tile_X3Y15_S_CPU_IRQ/FrameData[19] Tile_X3Y15_S_CPU_IRQ/FrameData[1] Tile_X3Y15_S_CPU_IRQ/FrameData[20]
+ Tile_X3Y15_S_CPU_IRQ/FrameData[21] Tile_X3Y15_S_CPU_IRQ/FrameData[22] Tile_X3Y15_S_CPU_IRQ/FrameData[23]
+ Tile_X3Y15_S_CPU_IRQ/FrameData[24] Tile_X3Y15_S_CPU_IRQ/FrameData[25] Tile_X3Y15_S_CPU_IRQ/FrameData[26]
+ Tile_X3Y15_S_CPU_IRQ/FrameData[27] Tile_X3Y15_S_CPU_IRQ/FrameData[28] Tile_X3Y15_S_CPU_IRQ/FrameData[29]
+ Tile_X3Y15_S_CPU_IRQ/FrameData[2] Tile_X3Y15_S_CPU_IRQ/FrameData[30] Tile_X3Y15_S_CPU_IRQ/FrameData[31]
+ Tile_X3Y15_S_CPU_IRQ/FrameData[3] Tile_X3Y15_S_CPU_IRQ/FrameData[4] Tile_X3Y15_S_CPU_IRQ/FrameData[5]
+ Tile_X3Y15_S_CPU_IRQ/FrameData[6] Tile_X3Y15_S_CPU_IRQ/FrameData[7] Tile_X3Y15_S_CPU_IRQ/FrameData[8]
+ Tile_X3Y15_S_CPU_IRQ/FrameData[9] Tile_X3Y15_S_CPU_IRQ/FrameData_O[0] Tile_X3Y15_S_CPU_IRQ/FrameData_O[10]
+ Tile_X3Y15_S_CPU_IRQ/FrameData_O[11] Tile_X3Y15_S_CPU_IRQ/FrameData_O[12] Tile_X3Y15_S_CPU_IRQ/FrameData_O[13]
+ Tile_X3Y15_S_CPU_IRQ/FrameData_O[14] Tile_X3Y15_S_CPU_IRQ/FrameData_O[15] Tile_X3Y15_S_CPU_IRQ/FrameData_O[16]
+ Tile_X3Y15_S_CPU_IRQ/FrameData_O[17] Tile_X3Y15_S_CPU_IRQ/FrameData_O[18] Tile_X3Y15_S_CPU_IRQ/FrameData_O[19]
+ Tile_X3Y15_S_CPU_IRQ/FrameData_O[1] Tile_X3Y15_S_CPU_IRQ/FrameData_O[20] Tile_X3Y15_S_CPU_IRQ/FrameData_O[21]
+ Tile_X3Y15_S_CPU_IRQ/FrameData_O[22] Tile_X3Y15_S_CPU_IRQ/FrameData_O[23] Tile_X3Y15_S_CPU_IRQ/FrameData_O[24]
+ Tile_X3Y15_S_CPU_IRQ/FrameData_O[25] Tile_X3Y15_S_CPU_IRQ/FrameData_O[26] Tile_X3Y15_S_CPU_IRQ/FrameData_O[27]
+ Tile_X3Y15_S_CPU_IRQ/FrameData_O[28] Tile_X3Y15_S_CPU_IRQ/FrameData_O[29] Tile_X3Y15_S_CPU_IRQ/FrameData_O[2]
+ Tile_X3Y15_S_CPU_IRQ/FrameData_O[30] Tile_X3Y15_S_CPU_IRQ/FrameData_O[31] Tile_X3Y15_S_CPU_IRQ/FrameData_O[3]
+ Tile_X3Y15_S_CPU_IRQ/FrameData_O[4] Tile_X3Y15_S_CPU_IRQ/FrameData_O[5] Tile_X3Y15_S_CPU_IRQ/FrameData_O[6]
+ Tile_X3Y15_S_CPU_IRQ/FrameData_O[7] Tile_X3Y15_S_CPU_IRQ/FrameData_O[8] Tile_X3Y15_S_CPU_IRQ/FrameData_O[9]
+ FrameStrobe[60] FrameStrobe[70] FrameStrobe[71] FrameStrobe[72] FrameStrobe[73]
+ FrameStrobe[74] FrameStrobe[75] FrameStrobe[76] FrameStrobe[77] FrameStrobe[78]
+ FrameStrobe[79] FrameStrobe[61] FrameStrobe[62] FrameStrobe[63] FrameStrobe[64]
+ FrameStrobe[65] FrameStrobe[66] FrameStrobe[67] FrameStrobe[68] FrameStrobe[69]
+ Tile_X3Y14_LUT4AB/FrameStrobe[0] Tile_X3Y14_LUT4AB/FrameStrobe[10] Tile_X3Y14_LUT4AB/FrameStrobe[11]
+ Tile_X3Y14_LUT4AB/FrameStrobe[12] Tile_X3Y14_LUT4AB/FrameStrobe[13] Tile_X3Y14_LUT4AB/FrameStrobe[14]
+ Tile_X3Y14_LUT4AB/FrameStrobe[15] Tile_X3Y14_LUT4AB/FrameStrobe[16] Tile_X3Y14_LUT4AB/FrameStrobe[17]
+ Tile_X3Y14_LUT4AB/FrameStrobe[18] Tile_X3Y14_LUT4AB/FrameStrobe[19] Tile_X3Y14_LUT4AB/FrameStrobe[1]
+ Tile_X3Y14_LUT4AB/FrameStrobe[2] Tile_X3Y14_LUT4AB/FrameStrobe[3] Tile_X3Y14_LUT4AB/FrameStrobe[4]
+ Tile_X3Y14_LUT4AB/FrameStrobe[5] Tile_X3Y14_LUT4AB/FrameStrobe[6] Tile_X3Y14_LUT4AB/FrameStrobe[7]
+ Tile_X3Y14_LUT4AB/FrameStrobe[8] Tile_X3Y14_LUT4AB/FrameStrobe[9] Tile_X3Y15_IRQ_top0
+ Tile_X3Y15_IRQ_top1 Tile_X3Y15_IRQ_top2 Tile_X3Y15_IRQ_top3 Tile_X3Y14_LUT4AB/N1END[0]
+ Tile_X3Y14_LUT4AB/N1END[1] Tile_X3Y14_LUT4AB/N1END[2] Tile_X3Y14_LUT4AB/N1END[3]
+ Tile_X3Y14_LUT4AB/N2MID[0] Tile_X3Y14_LUT4AB/N2MID[1] Tile_X3Y14_LUT4AB/N2MID[2]
+ Tile_X3Y14_LUT4AB/N2MID[3] Tile_X3Y14_LUT4AB/N2MID[4] Tile_X3Y14_LUT4AB/N2MID[5]
+ Tile_X3Y14_LUT4AB/N2MID[6] Tile_X3Y14_LUT4AB/N2MID[7] Tile_X3Y14_LUT4AB/N2END[0]
+ Tile_X3Y14_LUT4AB/N2END[1] Tile_X3Y14_LUT4AB/N2END[2] Tile_X3Y14_LUT4AB/N2END[3]
+ Tile_X3Y14_LUT4AB/N2END[4] Tile_X3Y14_LUT4AB/N2END[5] Tile_X3Y14_LUT4AB/N2END[6]
+ Tile_X3Y14_LUT4AB/N2END[7] Tile_X3Y14_LUT4AB/N4END[0] Tile_X3Y14_LUT4AB/N4END[10]
+ Tile_X3Y14_LUT4AB/N4END[11] Tile_X3Y14_LUT4AB/N4END[12] Tile_X3Y14_LUT4AB/N4END[13]
+ Tile_X3Y14_LUT4AB/N4END[14] Tile_X3Y14_LUT4AB/N4END[15] Tile_X3Y14_LUT4AB/N4END[1]
+ Tile_X3Y14_LUT4AB/N4END[2] Tile_X3Y14_LUT4AB/N4END[3] Tile_X3Y14_LUT4AB/N4END[4]
+ Tile_X3Y14_LUT4AB/N4END[5] Tile_X3Y14_LUT4AB/N4END[6] Tile_X3Y14_LUT4AB/N4END[7]
+ Tile_X3Y14_LUT4AB/N4END[8] Tile_X3Y14_LUT4AB/N4END[9] Tile_X3Y14_LUT4AB/NN4END[0]
+ Tile_X3Y14_LUT4AB/NN4END[10] Tile_X3Y14_LUT4AB/NN4END[11] Tile_X3Y14_LUT4AB/NN4END[12]
+ Tile_X3Y14_LUT4AB/NN4END[13] Tile_X3Y14_LUT4AB/NN4END[14] Tile_X3Y14_LUT4AB/NN4END[15]
+ Tile_X3Y14_LUT4AB/NN4END[1] Tile_X3Y14_LUT4AB/NN4END[2] Tile_X3Y14_LUT4AB/NN4END[3]
+ Tile_X3Y14_LUT4AB/NN4END[4] Tile_X3Y14_LUT4AB/NN4END[5] Tile_X3Y14_LUT4AB/NN4END[6]
+ Tile_X3Y14_LUT4AB/NN4END[7] Tile_X3Y14_LUT4AB/NN4END[8] Tile_X3Y14_LUT4AB/NN4END[9]
+ Tile_X3Y14_LUT4AB/S1BEG[0] Tile_X3Y14_LUT4AB/S1BEG[1] Tile_X3Y14_LUT4AB/S1BEG[2]
+ Tile_X3Y14_LUT4AB/S1BEG[3] Tile_X3Y14_LUT4AB/S2BEGb[0] Tile_X3Y14_LUT4AB/S2BEGb[1]
+ Tile_X3Y14_LUT4AB/S2BEGb[2] Tile_X3Y14_LUT4AB/S2BEGb[3] Tile_X3Y14_LUT4AB/S2BEGb[4]
+ Tile_X3Y14_LUT4AB/S2BEGb[5] Tile_X3Y14_LUT4AB/S2BEGb[6] Tile_X3Y14_LUT4AB/S2BEGb[7]
+ Tile_X3Y14_LUT4AB/S2BEG[0] Tile_X3Y14_LUT4AB/S2BEG[1] Tile_X3Y14_LUT4AB/S2BEG[2]
+ Tile_X3Y14_LUT4AB/S2BEG[3] Tile_X3Y14_LUT4AB/S2BEG[4] Tile_X3Y14_LUT4AB/S2BEG[5]
+ Tile_X3Y14_LUT4AB/S2BEG[6] Tile_X3Y14_LUT4AB/S2BEG[7] Tile_X3Y14_LUT4AB/S4BEG[0]
+ Tile_X3Y14_LUT4AB/S4BEG[10] Tile_X3Y14_LUT4AB/S4BEG[11] Tile_X3Y14_LUT4AB/S4BEG[12]
+ Tile_X3Y14_LUT4AB/S4BEG[13] Tile_X3Y14_LUT4AB/S4BEG[14] Tile_X3Y14_LUT4AB/S4BEG[15]
+ Tile_X3Y14_LUT4AB/S4BEG[1] Tile_X3Y14_LUT4AB/S4BEG[2] Tile_X3Y14_LUT4AB/S4BEG[3]
+ Tile_X3Y14_LUT4AB/S4BEG[4] Tile_X3Y14_LUT4AB/S4BEG[5] Tile_X3Y14_LUT4AB/S4BEG[6]
+ Tile_X3Y14_LUT4AB/S4BEG[7] Tile_X3Y14_LUT4AB/S4BEG[8] Tile_X3Y14_LUT4AB/S4BEG[9]
+ Tile_X3Y14_LUT4AB/SS4BEG[0] Tile_X3Y14_LUT4AB/SS4BEG[10] Tile_X3Y14_LUT4AB/SS4BEG[11]
+ Tile_X3Y14_LUT4AB/SS4BEG[12] Tile_X3Y14_LUT4AB/SS4BEG[13] Tile_X3Y14_LUT4AB/SS4BEG[14]
+ Tile_X3Y14_LUT4AB/SS4BEG[15] Tile_X3Y14_LUT4AB/SS4BEG[1] Tile_X3Y14_LUT4AB/SS4BEG[2]
+ Tile_X3Y14_LUT4AB/SS4BEG[3] Tile_X3Y14_LUT4AB/SS4BEG[4] Tile_X3Y14_LUT4AB/SS4BEG[5]
+ Tile_X3Y14_LUT4AB/SS4BEG[6] Tile_X3Y14_LUT4AB/SS4BEG[7] Tile_X3Y14_LUT4AB/SS4BEG[8]
+ Tile_X3Y14_LUT4AB/SS4BEG[9] UserCLK Tile_X3Y14_LUT4AB/UserCLK VGND VPWR S_CPU_IRQ
XTile_X5Y15_S_CPU_IF Tile_X5Y14_LUT4AB/Ci Tile_X5Y15_S_CPU_IF/FrameData[0] Tile_X5Y15_S_CPU_IF/FrameData[10]
+ Tile_X5Y15_S_CPU_IF/FrameData[11] Tile_X5Y15_S_CPU_IF/FrameData[12] Tile_X5Y15_S_CPU_IF/FrameData[13]
+ Tile_X5Y15_S_CPU_IF/FrameData[14] Tile_X5Y15_S_CPU_IF/FrameData[15] Tile_X5Y15_S_CPU_IF/FrameData[16]
+ Tile_X5Y15_S_CPU_IF/FrameData[17] Tile_X5Y15_S_CPU_IF/FrameData[18] Tile_X5Y15_S_CPU_IF/FrameData[19]
+ Tile_X5Y15_S_CPU_IF/FrameData[1] Tile_X5Y15_S_CPU_IF/FrameData[20] Tile_X5Y15_S_CPU_IF/FrameData[21]
+ Tile_X5Y15_S_CPU_IF/FrameData[22] Tile_X5Y15_S_CPU_IF/FrameData[23] Tile_X5Y15_S_CPU_IF/FrameData[24]
+ Tile_X5Y15_S_CPU_IF/FrameData[25] Tile_X5Y15_S_CPU_IF/FrameData[26] Tile_X5Y15_S_CPU_IF/FrameData[27]
+ Tile_X5Y15_S_CPU_IF/FrameData[28] Tile_X5Y15_S_CPU_IF/FrameData[29] Tile_X5Y15_S_CPU_IF/FrameData[2]
+ Tile_X5Y15_S_CPU_IF/FrameData[30] Tile_X5Y15_S_CPU_IF/FrameData[31] Tile_X5Y15_S_CPU_IF/FrameData[3]
+ Tile_X5Y15_S_CPU_IF/FrameData[4] Tile_X5Y15_S_CPU_IF/FrameData[5] Tile_X5Y15_S_CPU_IF/FrameData[6]
+ Tile_X5Y15_S_CPU_IF/FrameData[7] Tile_X5Y15_S_CPU_IF/FrameData[8] Tile_X5Y15_S_CPU_IF/FrameData[9]
+ Tile_X6Y15_S_CPU_IF/FrameData[0] Tile_X6Y15_S_CPU_IF/FrameData[10] Tile_X6Y15_S_CPU_IF/FrameData[11]
+ Tile_X6Y15_S_CPU_IF/FrameData[12] Tile_X6Y15_S_CPU_IF/FrameData[13] Tile_X6Y15_S_CPU_IF/FrameData[14]
+ Tile_X6Y15_S_CPU_IF/FrameData[15] Tile_X6Y15_S_CPU_IF/FrameData[16] Tile_X6Y15_S_CPU_IF/FrameData[17]
+ Tile_X6Y15_S_CPU_IF/FrameData[18] Tile_X6Y15_S_CPU_IF/FrameData[19] Tile_X6Y15_S_CPU_IF/FrameData[1]
+ Tile_X6Y15_S_CPU_IF/FrameData[20] Tile_X6Y15_S_CPU_IF/FrameData[21] Tile_X6Y15_S_CPU_IF/FrameData[22]
+ Tile_X6Y15_S_CPU_IF/FrameData[23] Tile_X6Y15_S_CPU_IF/FrameData[24] Tile_X6Y15_S_CPU_IF/FrameData[25]
+ Tile_X6Y15_S_CPU_IF/FrameData[26] Tile_X6Y15_S_CPU_IF/FrameData[27] Tile_X6Y15_S_CPU_IF/FrameData[28]
+ Tile_X6Y15_S_CPU_IF/FrameData[29] Tile_X6Y15_S_CPU_IF/FrameData[2] Tile_X6Y15_S_CPU_IF/FrameData[30]
+ Tile_X6Y15_S_CPU_IF/FrameData[31] Tile_X6Y15_S_CPU_IF/FrameData[3] Tile_X6Y15_S_CPU_IF/FrameData[4]
+ Tile_X6Y15_S_CPU_IF/FrameData[5] Tile_X6Y15_S_CPU_IF/FrameData[6] Tile_X6Y15_S_CPU_IF/FrameData[7]
+ Tile_X6Y15_S_CPU_IF/FrameData[8] Tile_X6Y15_S_CPU_IF/FrameData[9] FrameStrobe[100]
+ FrameStrobe[110] FrameStrobe[111] FrameStrobe[112] FrameStrobe[113] FrameStrobe[114]
+ FrameStrobe[115] FrameStrobe[116] FrameStrobe[117] FrameStrobe[118] FrameStrobe[119]
+ FrameStrobe[101] FrameStrobe[102] FrameStrobe[103] FrameStrobe[104] FrameStrobe[105]
+ FrameStrobe[106] FrameStrobe[107] FrameStrobe[108] FrameStrobe[109] Tile_X5Y14_LUT4AB/FrameStrobe[0]
+ Tile_X5Y14_LUT4AB/FrameStrobe[10] Tile_X5Y14_LUT4AB/FrameStrobe[11] Tile_X5Y14_LUT4AB/FrameStrobe[12]
+ Tile_X5Y14_LUT4AB/FrameStrobe[13] Tile_X5Y14_LUT4AB/FrameStrobe[14] Tile_X5Y14_LUT4AB/FrameStrobe[15]
+ Tile_X5Y14_LUT4AB/FrameStrobe[16] Tile_X5Y14_LUT4AB/FrameStrobe[17] Tile_X5Y14_LUT4AB/FrameStrobe[18]
+ Tile_X5Y14_LUT4AB/FrameStrobe[19] Tile_X5Y14_LUT4AB/FrameStrobe[1] Tile_X5Y14_LUT4AB/FrameStrobe[2]
+ Tile_X5Y14_LUT4AB/FrameStrobe[3] Tile_X5Y14_LUT4AB/FrameStrobe[4] Tile_X5Y14_LUT4AB/FrameStrobe[5]
+ Tile_X5Y14_LUT4AB/FrameStrobe[6] Tile_X5Y14_LUT4AB/FrameStrobe[7] Tile_X5Y14_LUT4AB/FrameStrobe[8]
+ Tile_X5Y14_LUT4AB/FrameStrobe[9] Tile_X5Y15_I_top0 Tile_X5Y15_I_top1 Tile_X5Y15_I_top10
+ Tile_X5Y15_I_top11 Tile_X5Y15_I_top12 Tile_X5Y15_I_top13 Tile_X5Y15_I_top14 Tile_X5Y15_I_top15
+ Tile_X5Y15_I_top2 Tile_X5Y15_I_top3 Tile_X5Y15_I_top4 Tile_X5Y15_I_top5 Tile_X5Y15_I_top6
+ Tile_X5Y15_I_top7 Tile_X5Y15_I_top8 Tile_X5Y15_I_top9 Tile_X5Y14_LUT4AB/N1END[0]
+ Tile_X5Y14_LUT4AB/N1END[1] Tile_X5Y14_LUT4AB/N1END[2] Tile_X5Y14_LUT4AB/N1END[3]
+ Tile_X5Y14_LUT4AB/N2MID[0] Tile_X5Y14_LUT4AB/N2MID[1] Tile_X5Y14_LUT4AB/N2MID[2]
+ Tile_X5Y14_LUT4AB/N2MID[3] Tile_X5Y14_LUT4AB/N2MID[4] Tile_X5Y14_LUT4AB/N2MID[5]
+ Tile_X5Y14_LUT4AB/N2MID[6] Tile_X5Y14_LUT4AB/N2MID[7] Tile_X5Y14_LUT4AB/N2END[0]
+ Tile_X5Y14_LUT4AB/N2END[1] Tile_X5Y14_LUT4AB/N2END[2] Tile_X5Y14_LUT4AB/N2END[3]
+ Tile_X5Y14_LUT4AB/N2END[4] Tile_X5Y14_LUT4AB/N2END[5] Tile_X5Y14_LUT4AB/N2END[6]
+ Tile_X5Y14_LUT4AB/N2END[7] Tile_X5Y14_LUT4AB/N4END[0] Tile_X5Y14_LUT4AB/N4END[10]
+ Tile_X5Y14_LUT4AB/N4END[11] Tile_X5Y14_LUT4AB/N4END[12] Tile_X5Y14_LUT4AB/N4END[13]
+ Tile_X5Y14_LUT4AB/N4END[14] Tile_X5Y14_LUT4AB/N4END[15] Tile_X5Y14_LUT4AB/N4END[1]
+ Tile_X5Y14_LUT4AB/N4END[2] Tile_X5Y14_LUT4AB/N4END[3] Tile_X5Y14_LUT4AB/N4END[4]
+ Tile_X5Y14_LUT4AB/N4END[5] Tile_X5Y14_LUT4AB/N4END[6] Tile_X5Y14_LUT4AB/N4END[7]
+ Tile_X5Y14_LUT4AB/N4END[8] Tile_X5Y14_LUT4AB/N4END[9] Tile_X5Y14_LUT4AB/NN4END[0]
+ Tile_X5Y14_LUT4AB/NN4END[10] Tile_X5Y14_LUT4AB/NN4END[11] Tile_X5Y14_LUT4AB/NN4END[12]
+ Tile_X5Y14_LUT4AB/NN4END[13] Tile_X5Y14_LUT4AB/NN4END[14] Tile_X5Y14_LUT4AB/NN4END[15]
+ Tile_X5Y14_LUT4AB/NN4END[1] Tile_X5Y14_LUT4AB/NN4END[2] Tile_X5Y14_LUT4AB/NN4END[3]
+ Tile_X5Y14_LUT4AB/NN4END[4] Tile_X5Y14_LUT4AB/NN4END[5] Tile_X5Y14_LUT4AB/NN4END[6]
+ Tile_X5Y14_LUT4AB/NN4END[7] Tile_X5Y14_LUT4AB/NN4END[8] Tile_X5Y14_LUT4AB/NN4END[9]
+ Tile_X5Y15_O_top0 Tile_X5Y15_O_top1 Tile_X5Y15_O_top10 Tile_X5Y15_O_top11 Tile_X5Y15_O_top12
+ Tile_X5Y15_O_top13 Tile_X5Y15_O_top14 Tile_X5Y15_O_top15 Tile_X5Y15_O_top2 Tile_X5Y15_O_top3
+ Tile_X5Y15_O_top4 Tile_X5Y15_O_top5 Tile_X5Y15_O_top6 Tile_X5Y15_O_top7 Tile_X5Y15_O_top8
+ Tile_X5Y15_O_top9 Tile_X5Y14_LUT4AB/S1BEG[0] Tile_X5Y14_LUT4AB/S1BEG[1] Tile_X5Y14_LUT4AB/S1BEG[2]
+ Tile_X5Y14_LUT4AB/S1BEG[3] Tile_X5Y14_LUT4AB/S2BEGb[0] Tile_X5Y14_LUT4AB/S2BEGb[1]
+ Tile_X5Y14_LUT4AB/S2BEGb[2] Tile_X5Y14_LUT4AB/S2BEGb[3] Tile_X5Y14_LUT4AB/S2BEGb[4]
+ Tile_X5Y14_LUT4AB/S2BEGb[5] Tile_X5Y14_LUT4AB/S2BEGb[6] Tile_X5Y14_LUT4AB/S2BEGb[7]
+ Tile_X5Y14_LUT4AB/S2BEG[0] Tile_X5Y14_LUT4AB/S2BEG[1] Tile_X5Y14_LUT4AB/S2BEG[2]
+ Tile_X5Y14_LUT4AB/S2BEG[3] Tile_X5Y14_LUT4AB/S2BEG[4] Tile_X5Y14_LUT4AB/S2BEG[5]
+ Tile_X5Y14_LUT4AB/S2BEG[6] Tile_X5Y14_LUT4AB/S2BEG[7] Tile_X5Y14_LUT4AB/S4BEG[0]
+ Tile_X5Y14_LUT4AB/S4BEG[10] Tile_X5Y14_LUT4AB/S4BEG[11] Tile_X5Y14_LUT4AB/S4BEG[12]
+ Tile_X5Y14_LUT4AB/S4BEG[13] Tile_X5Y14_LUT4AB/S4BEG[14] Tile_X5Y14_LUT4AB/S4BEG[15]
+ Tile_X5Y14_LUT4AB/S4BEG[1] Tile_X5Y14_LUT4AB/S4BEG[2] Tile_X5Y14_LUT4AB/S4BEG[3]
+ Tile_X5Y14_LUT4AB/S4BEG[4] Tile_X5Y14_LUT4AB/S4BEG[5] Tile_X5Y14_LUT4AB/S4BEG[6]
+ Tile_X5Y14_LUT4AB/S4BEG[7] Tile_X5Y14_LUT4AB/S4BEG[8] Tile_X5Y14_LUT4AB/S4BEG[9]
+ Tile_X5Y14_LUT4AB/SS4BEG[0] Tile_X5Y14_LUT4AB/SS4BEG[10] Tile_X5Y14_LUT4AB/SS4BEG[11]
+ Tile_X5Y14_LUT4AB/SS4BEG[12] Tile_X5Y14_LUT4AB/SS4BEG[13] Tile_X5Y14_LUT4AB/SS4BEG[14]
+ Tile_X5Y14_LUT4AB/SS4BEG[15] Tile_X5Y14_LUT4AB/SS4BEG[1] Tile_X5Y14_LUT4AB/SS4BEG[2]
+ Tile_X5Y14_LUT4AB/SS4BEG[3] Tile_X5Y14_LUT4AB/SS4BEG[4] Tile_X5Y14_LUT4AB/SS4BEG[5]
+ Tile_X5Y14_LUT4AB/SS4BEG[6] Tile_X5Y14_LUT4AB/SS4BEG[7] Tile_X5Y14_LUT4AB/SS4BEG[8]
+ Tile_X5Y14_LUT4AB/SS4BEG[9] UserCLK Tile_X5Y14_LUT4AB/UserCLK VGND VPWR S_CPU_IF
XTile_X2Y6_LUT4AB Tile_X2Y7_LUT4AB/Co Tile_X2Y6_LUT4AB/Co Tile_X3Y6_LUT4AB/E1END[0]
+ Tile_X3Y6_LUT4AB/E1END[1] Tile_X3Y6_LUT4AB/E1END[2] Tile_X3Y6_LUT4AB/E1END[3] Tile_X2Y6_LUT4AB/E1END[0]
+ Tile_X2Y6_LUT4AB/E1END[1] Tile_X2Y6_LUT4AB/E1END[2] Tile_X2Y6_LUT4AB/E1END[3] Tile_X3Y6_LUT4AB/E2MID[0]
+ Tile_X3Y6_LUT4AB/E2MID[1] Tile_X3Y6_LUT4AB/E2MID[2] Tile_X3Y6_LUT4AB/E2MID[3] Tile_X3Y6_LUT4AB/E2MID[4]
+ Tile_X3Y6_LUT4AB/E2MID[5] Tile_X3Y6_LUT4AB/E2MID[6] Tile_X3Y6_LUT4AB/E2MID[7] Tile_X3Y6_LUT4AB/E2END[0]
+ Tile_X3Y6_LUT4AB/E2END[1] Tile_X3Y6_LUT4AB/E2END[2] Tile_X3Y6_LUT4AB/E2END[3] Tile_X3Y6_LUT4AB/E2END[4]
+ Tile_X3Y6_LUT4AB/E2END[5] Tile_X3Y6_LUT4AB/E2END[6] Tile_X3Y6_LUT4AB/E2END[7] Tile_X2Y6_LUT4AB/E2END[0]
+ Tile_X2Y6_LUT4AB/E2END[1] Tile_X2Y6_LUT4AB/E2END[2] Tile_X2Y6_LUT4AB/E2END[3] Tile_X2Y6_LUT4AB/E2END[4]
+ Tile_X2Y6_LUT4AB/E2END[5] Tile_X2Y6_LUT4AB/E2END[6] Tile_X2Y6_LUT4AB/E2END[7] Tile_X2Y6_LUT4AB/E2MID[0]
+ Tile_X2Y6_LUT4AB/E2MID[1] Tile_X2Y6_LUT4AB/E2MID[2] Tile_X2Y6_LUT4AB/E2MID[3] Tile_X2Y6_LUT4AB/E2MID[4]
+ Tile_X2Y6_LUT4AB/E2MID[5] Tile_X2Y6_LUT4AB/E2MID[6] Tile_X2Y6_LUT4AB/E2MID[7] Tile_X3Y6_LUT4AB/E6END[0]
+ Tile_X3Y6_LUT4AB/E6END[10] Tile_X3Y6_LUT4AB/E6END[11] Tile_X3Y6_LUT4AB/E6END[1]
+ Tile_X3Y6_LUT4AB/E6END[2] Tile_X3Y6_LUT4AB/E6END[3] Tile_X3Y6_LUT4AB/E6END[4] Tile_X3Y6_LUT4AB/E6END[5]
+ Tile_X3Y6_LUT4AB/E6END[6] Tile_X3Y6_LUT4AB/E6END[7] Tile_X3Y6_LUT4AB/E6END[8] Tile_X3Y6_LUT4AB/E6END[9]
+ Tile_X2Y6_LUT4AB/E6END[0] Tile_X2Y6_LUT4AB/E6END[10] Tile_X2Y6_LUT4AB/E6END[11]
+ Tile_X2Y6_LUT4AB/E6END[1] Tile_X2Y6_LUT4AB/E6END[2] Tile_X2Y6_LUT4AB/E6END[3] Tile_X2Y6_LUT4AB/E6END[4]
+ Tile_X2Y6_LUT4AB/E6END[5] Tile_X2Y6_LUT4AB/E6END[6] Tile_X2Y6_LUT4AB/E6END[7] Tile_X2Y6_LUT4AB/E6END[8]
+ Tile_X2Y6_LUT4AB/E6END[9] Tile_X3Y6_LUT4AB/EE4END[0] Tile_X3Y6_LUT4AB/EE4END[10]
+ Tile_X3Y6_LUT4AB/EE4END[11] Tile_X3Y6_LUT4AB/EE4END[12] Tile_X3Y6_LUT4AB/EE4END[13]
+ Tile_X3Y6_LUT4AB/EE4END[14] Tile_X3Y6_LUT4AB/EE4END[15] Tile_X3Y6_LUT4AB/EE4END[1]
+ Tile_X3Y6_LUT4AB/EE4END[2] Tile_X3Y6_LUT4AB/EE4END[3] Tile_X3Y6_LUT4AB/EE4END[4]
+ Tile_X3Y6_LUT4AB/EE4END[5] Tile_X3Y6_LUT4AB/EE4END[6] Tile_X3Y6_LUT4AB/EE4END[7]
+ Tile_X3Y6_LUT4AB/EE4END[8] Tile_X3Y6_LUT4AB/EE4END[9] Tile_X2Y6_LUT4AB/EE4END[0]
+ Tile_X2Y6_LUT4AB/EE4END[10] Tile_X2Y6_LUT4AB/EE4END[11] Tile_X2Y6_LUT4AB/EE4END[12]
+ Tile_X2Y6_LUT4AB/EE4END[13] Tile_X2Y6_LUT4AB/EE4END[14] Tile_X2Y6_LUT4AB/EE4END[15]
+ Tile_X2Y6_LUT4AB/EE4END[1] Tile_X2Y6_LUT4AB/EE4END[2] Tile_X2Y6_LUT4AB/EE4END[3]
+ Tile_X2Y6_LUT4AB/EE4END[4] Tile_X2Y6_LUT4AB/EE4END[5] Tile_X2Y6_LUT4AB/EE4END[6]
+ Tile_X2Y6_LUT4AB/EE4END[7] Tile_X2Y6_LUT4AB/EE4END[8] Tile_X2Y6_LUT4AB/EE4END[9]
+ Tile_X2Y6_LUT4AB/FrameData[0] Tile_X2Y6_LUT4AB/FrameData[10] Tile_X2Y6_LUT4AB/FrameData[11]
+ Tile_X2Y6_LUT4AB/FrameData[12] Tile_X2Y6_LUT4AB/FrameData[13] Tile_X2Y6_LUT4AB/FrameData[14]
+ Tile_X2Y6_LUT4AB/FrameData[15] Tile_X2Y6_LUT4AB/FrameData[16] Tile_X2Y6_LUT4AB/FrameData[17]
+ Tile_X2Y6_LUT4AB/FrameData[18] Tile_X2Y6_LUT4AB/FrameData[19] Tile_X2Y6_LUT4AB/FrameData[1]
+ Tile_X2Y6_LUT4AB/FrameData[20] Tile_X2Y6_LUT4AB/FrameData[21] Tile_X2Y6_LUT4AB/FrameData[22]
+ Tile_X2Y6_LUT4AB/FrameData[23] Tile_X2Y6_LUT4AB/FrameData[24] Tile_X2Y6_LUT4AB/FrameData[25]
+ Tile_X2Y6_LUT4AB/FrameData[26] Tile_X2Y6_LUT4AB/FrameData[27] Tile_X2Y6_LUT4AB/FrameData[28]
+ Tile_X2Y6_LUT4AB/FrameData[29] Tile_X2Y6_LUT4AB/FrameData[2] Tile_X2Y6_LUT4AB/FrameData[30]
+ Tile_X2Y6_LUT4AB/FrameData[31] Tile_X2Y6_LUT4AB/FrameData[3] Tile_X2Y6_LUT4AB/FrameData[4]
+ Tile_X2Y6_LUT4AB/FrameData[5] Tile_X2Y6_LUT4AB/FrameData[6] Tile_X2Y6_LUT4AB/FrameData[7]
+ Tile_X2Y6_LUT4AB/FrameData[8] Tile_X2Y6_LUT4AB/FrameData[9] Tile_X3Y6_LUT4AB/FrameData[0]
+ Tile_X3Y6_LUT4AB/FrameData[10] Tile_X3Y6_LUT4AB/FrameData[11] Tile_X3Y6_LUT4AB/FrameData[12]
+ Tile_X3Y6_LUT4AB/FrameData[13] Tile_X3Y6_LUT4AB/FrameData[14] Tile_X3Y6_LUT4AB/FrameData[15]
+ Tile_X3Y6_LUT4AB/FrameData[16] Tile_X3Y6_LUT4AB/FrameData[17] Tile_X3Y6_LUT4AB/FrameData[18]
+ Tile_X3Y6_LUT4AB/FrameData[19] Tile_X3Y6_LUT4AB/FrameData[1] Tile_X3Y6_LUT4AB/FrameData[20]
+ Tile_X3Y6_LUT4AB/FrameData[21] Tile_X3Y6_LUT4AB/FrameData[22] Tile_X3Y6_LUT4AB/FrameData[23]
+ Tile_X3Y6_LUT4AB/FrameData[24] Tile_X3Y6_LUT4AB/FrameData[25] Tile_X3Y6_LUT4AB/FrameData[26]
+ Tile_X3Y6_LUT4AB/FrameData[27] Tile_X3Y6_LUT4AB/FrameData[28] Tile_X3Y6_LUT4AB/FrameData[29]
+ Tile_X3Y6_LUT4AB/FrameData[2] Tile_X3Y6_LUT4AB/FrameData[30] Tile_X3Y6_LUT4AB/FrameData[31]
+ Tile_X3Y6_LUT4AB/FrameData[3] Tile_X3Y6_LUT4AB/FrameData[4] Tile_X3Y6_LUT4AB/FrameData[5]
+ Tile_X3Y6_LUT4AB/FrameData[6] Tile_X3Y6_LUT4AB/FrameData[7] Tile_X3Y6_LUT4AB/FrameData[8]
+ Tile_X3Y6_LUT4AB/FrameData[9] Tile_X2Y6_LUT4AB/FrameStrobe[0] Tile_X2Y6_LUT4AB/FrameStrobe[10]
+ Tile_X2Y6_LUT4AB/FrameStrobe[11] Tile_X2Y6_LUT4AB/FrameStrobe[12] Tile_X2Y6_LUT4AB/FrameStrobe[13]
+ Tile_X2Y6_LUT4AB/FrameStrobe[14] Tile_X2Y6_LUT4AB/FrameStrobe[15] Tile_X2Y6_LUT4AB/FrameStrobe[16]
+ Tile_X2Y6_LUT4AB/FrameStrobe[17] Tile_X2Y6_LUT4AB/FrameStrobe[18] Tile_X2Y6_LUT4AB/FrameStrobe[19]
+ Tile_X2Y6_LUT4AB/FrameStrobe[1] Tile_X2Y6_LUT4AB/FrameStrobe[2] Tile_X2Y6_LUT4AB/FrameStrobe[3]
+ Tile_X2Y6_LUT4AB/FrameStrobe[4] Tile_X2Y6_LUT4AB/FrameStrobe[5] Tile_X2Y6_LUT4AB/FrameStrobe[6]
+ Tile_X2Y6_LUT4AB/FrameStrobe[7] Tile_X2Y6_LUT4AB/FrameStrobe[8] Tile_X2Y6_LUT4AB/FrameStrobe[9]
+ Tile_X2Y5_LUT4AB/FrameStrobe[0] Tile_X2Y5_LUT4AB/FrameStrobe[10] Tile_X2Y5_LUT4AB/FrameStrobe[11]
+ Tile_X2Y5_LUT4AB/FrameStrobe[12] Tile_X2Y5_LUT4AB/FrameStrobe[13] Tile_X2Y5_LUT4AB/FrameStrobe[14]
+ Tile_X2Y5_LUT4AB/FrameStrobe[15] Tile_X2Y5_LUT4AB/FrameStrobe[16] Tile_X2Y5_LUT4AB/FrameStrobe[17]
+ Tile_X2Y5_LUT4AB/FrameStrobe[18] Tile_X2Y5_LUT4AB/FrameStrobe[19] Tile_X2Y5_LUT4AB/FrameStrobe[1]
+ Tile_X2Y5_LUT4AB/FrameStrobe[2] Tile_X2Y5_LUT4AB/FrameStrobe[3] Tile_X2Y5_LUT4AB/FrameStrobe[4]
+ Tile_X2Y5_LUT4AB/FrameStrobe[5] Tile_X2Y5_LUT4AB/FrameStrobe[6] Tile_X2Y5_LUT4AB/FrameStrobe[7]
+ Tile_X2Y5_LUT4AB/FrameStrobe[8] Tile_X2Y5_LUT4AB/FrameStrobe[9] Tile_X2Y6_LUT4AB/N1BEG[0]
+ Tile_X2Y6_LUT4AB/N1BEG[1] Tile_X2Y6_LUT4AB/N1BEG[2] Tile_X2Y6_LUT4AB/N1BEG[3] Tile_X2Y7_LUT4AB/N1BEG[0]
+ Tile_X2Y7_LUT4AB/N1BEG[1] Tile_X2Y7_LUT4AB/N1BEG[2] Tile_X2Y7_LUT4AB/N1BEG[3] Tile_X2Y6_LUT4AB/N2BEG[0]
+ Tile_X2Y6_LUT4AB/N2BEG[1] Tile_X2Y6_LUT4AB/N2BEG[2] Tile_X2Y6_LUT4AB/N2BEG[3] Tile_X2Y6_LUT4AB/N2BEG[4]
+ Tile_X2Y6_LUT4AB/N2BEG[5] Tile_X2Y6_LUT4AB/N2BEG[6] Tile_X2Y6_LUT4AB/N2BEG[7] Tile_X2Y5_LUT4AB/N2END[0]
+ Tile_X2Y5_LUT4AB/N2END[1] Tile_X2Y5_LUT4AB/N2END[2] Tile_X2Y5_LUT4AB/N2END[3] Tile_X2Y5_LUT4AB/N2END[4]
+ Tile_X2Y5_LUT4AB/N2END[5] Tile_X2Y5_LUT4AB/N2END[6] Tile_X2Y5_LUT4AB/N2END[7] Tile_X2Y6_LUT4AB/N2END[0]
+ Tile_X2Y6_LUT4AB/N2END[1] Tile_X2Y6_LUT4AB/N2END[2] Tile_X2Y6_LUT4AB/N2END[3] Tile_X2Y6_LUT4AB/N2END[4]
+ Tile_X2Y6_LUT4AB/N2END[5] Tile_X2Y6_LUT4AB/N2END[6] Tile_X2Y6_LUT4AB/N2END[7] Tile_X2Y7_LUT4AB/N2BEG[0]
+ Tile_X2Y7_LUT4AB/N2BEG[1] Tile_X2Y7_LUT4AB/N2BEG[2] Tile_X2Y7_LUT4AB/N2BEG[3] Tile_X2Y7_LUT4AB/N2BEG[4]
+ Tile_X2Y7_LUT4AB/N2BEG[5] Tile_X2Y7_LUT4AB/N2BEG[6] Tile_X2Y7_LUT4AB/N2BEG[7] Tile_X2Y6_LUT4AB/N4BEG[0]
+ Tile_X2Y6_LUT4AB/N4BEG[10] Tile_X2Y6_LUT4AB/N4BEG[11] Tile_X2Y6_LUT4AB/N4BEG[12]
+ Tile_X2Y6_LUT4AB/N4BEG[13] Tile_X2Y6_LUT4AB/N4BEG[14] Tile_X2Y6_LUT4AB/N4BEG[15]
+ Tile_X2Y6_LUT4AB/N4BEG[1] Tile_X2Y6_LUT4AB/N4BEG[2] Tile_X2Y6_LUT4AB/N4BEG[3] Tile_X2Y6_LUT4AB/N4BEG[4]
+ Tile_X2Y6_LUT4AB/N4BEG[5] Tile_X2Y6_LUT4AB/N4BEG[6] Tile_X2Y6_LUT4AB/N4BEG[7] Tile_X2Y6_LUT4AB/N4BEG[8]
+ Tile_X2Y6_LUT4AB/N4BEG[9] Tile_X2Y7_LUT4AB/N4BEG[0] Tile_X2Y7_LUT4AB/N4BEG[10] Tile_X2Y7_LUT4AB/N4BEG[11]
+ Tile_X2Y7_LUT4AB/N4BEG[12] Tile_X2Y7_LUT4AB/N4BEG[13] Tile_X2Y7_LUT4AB/N4BEG[14]
+ Tile_X2Y7_LUT4AB/N4BEG[15] Tile_X2Y7_LUT4AB/N4BEG[1] Tile_X2Y7_LUT4AB/N4BEG[2] Tile_X2Y7_LUT4AB/N4BEG[3]
+ Tile_X2Y7_LUT4AB/N4BEG[4] Tile_X2Y7_LUT4AB/N4BEG[5] Tile_X2Y7_LUT4AB/N4BEG[6] Tile_X2Y7_LUT4AB/N4BEG[7]
+ Tile_X2Y7_LUT4AB/N4BEG[8] Tile_X2Y7_LUT4AB/N4BEG[9] Tile_X2Y6_LUT4AB/NN4BEG[0] Tile_X2Y6_LUT4AB/NN4BEG[10]
+ Tile_X2Y6_LUT4AB/NN4BEG[11] Tile_X2Y6_LUT4AB/NN4BEG[12] Tile_X2Y6_LUT4AB/NN4BEG[13]
+ Tile_X2Y6_LUT4AB/NN4BEG[14] Tile_X2Y6_LUT4AB/NN4BEG[15] Tile_X2Y6_LUT4AB/NN4BEG[1]
+ Tile_X2Y6_LUT4AB/NN4BEG[2] Tile_X2Y6_LUT4AB/NN4BEG[3] Tile_X2Y6_LUT4AB/NN4BEG[4]
+ Tile_X2Y6_LUT4AB/NN4BEG[5] Tile_X2Y6_LUT4AB/NN4BEG[6] Tile_X2Y6_LUT4AB/NN4BEG[7]
+ Tile_X2Y6_LUT4AB/NN4BEG[8] Tile_X2Y6_LUT4AB/NN4BEG[9] Tile_X2Y7_LUT4AB/NN4BEG[0]
+ Tile_X2Y7_LUT4AB/NN4BEG[10] Tile_X2Y7_LUT4AB/NN4BEG[11] Tile_X2Y7_LUT4AB/NN4BEG[12]
+ Tile_X2Y7_LUT4AB/NN4BEG[13] Tile_X2Y7_LUT4AB/NN4BEG[14] Tile_X2Y7_LUT4AB/NN4BEG[15]
+ Tile_X2Y7_LUT4AB/NN4BEG[1] Tile_X2Y7_LUT4AB/NN4BEG[2] Tile_X2Y7_LUT4AB/NN4BEG[3]
+ Tile_X2Y7_LUT4AB/NN4BEG[4] Tile_X2Y7_LUT4AB/NN4BEG[5] Tile_X2Y7_LUT4AB/NN4BEG[6]
+ Tile_X2Y7_LUT4AB/NN4BEG[7] Tile_X2Y7_LUT4AB/NN4BEG[8] Tile_X2Y7_LUT4AB/NN4BEG[9]
+ Tile_X2Y7_LUT4AB/S1END[0] Tile_X2Y7_LUT4AB/S1END[1] Tile_X2Y7_LUT4AB/S1END[2] Tile_X2Y7_LUT4AB/S1END[3]
+ Tile_X2Y6_LUT4AB/S1END[0] Tile_X2Y6_LUT4AB/S1END[1] Tile_X2Y6_LUT4AB/S1END[2] Tile_X2Y6_LUT4AB/S1END[3]
+ Tile_X2Y7_LUT4AB/S2MID[0] Tile_X2Y7_LUT4AB/S2MID[1] Tile_X2Y7_LUT4AB/S2MID[2] Tile_X2Y7_LUT4AB/S2MID[3]
+ Tile_X2Y7_LUT4AB/S2MID[4] Tile_X2Y7_LUT4AB/S2MID[5] Tile_X2Y7_LUT4AB/S2MID[6] Tile_X2Y7_LUT4AB/S2MID[7]
+ Tile_X2Y7_LUT4AB/S2END[0] Tile_X2Y7_LUT4AB/S2END[1] Tile_X2Y7_LUT4AB/S2END[2] Tile_X2Y7_LUT4AB/S2END[3]
+ Tile_X2Y7_LUT4AB/S2END[4] Tile_X2Y7_LUT4AB/S2END[5] Tile_X2Y7_LUT4AB/S2END[6] Tile_X2Y7_LUT4AB/S2END[7]
+ Tile_X2Y6_LUT4AB/S2END[0] Tile_X2Y6_LUT4AB/S2END[1] Tile_X2Y6_LUT4AB/S2END[2] Tile_X2Y6_LUT4AB/S2END[3]
+ Tile_X2Y6_LUT4AB/S2END[4] Tile_X2Y6_LUT4AB/S2END[5] Tile_X2Y6_LUT4AB/S2END[6] Tile_X2Y6_LUT4AB/S2END[7]
+ Tile_X2Y6_LUT4AB/S2MID[0] Tile_X2Y6_LUT4AB/S2MID[1] Tile_X2Y6_LUT4AB/S2MID[2] Tile_X2Y6_LUT4AB/S2MID[3]
+ Tile_X2Y6_LUT4AB/S2MID[4] Tile_X2Y6_LUT4AB/S2MID[5] Tile_X2Y6_LUT4AB/S2MID[6] Tile_X2Y6_LUT4AB/S2MID[7]
+ Tile_X2Y7_LUT4AB/S4END[0] Tile_X2Y7_LUT4AB/S4END[10] Tile_X2Y7_LUT4AB/S4END[11]
+ Tile_X2Y7_LUT4AB/S4END[12] Tile_X2Y7_LUT4AB/S4END[13] Tile_X2Y7_LUT4AB/S4END[14]
+ Tile_X2Y7_LUT4AB/S4END[15] Tile_X2Y7_LUT4AB/S4END[1] Tile_X2Y7_LUT4AB/S4END[2] Tile_X2Y7_LUT4AB/S4END[3]
+ Tile_X2Y7_LUT4AB/S4END[4] Tile_X2Y7_LUT4AB/S4END[5] Tile_X2Y7_LUT4AB/S4END[6] Tile_X2Y7_LUT4AB/S4END[7]
+ Tile_X2Y7_LUT4AB/S4END[8] Tile_X2Y7_LUT4AB/S4END[9] Tile_X2Y6_LUT4AB/S4END[0] Tile_X2Y6_LUT4AB/S4END[10]
+ Tile_X2Y6_LUT4AB/S4END[11] Tile_X2Y6_LUT4AB/S4END[12] Tile_X2Y6_LUT4AB/S4END[13]
+ Tile_X2Y6_LUT4AB/S4END[14] Tile_X2Y6_LUT4AB/S4END[15] Tile_X2Y6_LUT4AB/S4END[1]
+ Tile_X2Y6_LUT4AB/S4END[2] Tile_X2Y6_LUT4AB/S4END[3] Tile_X2Y6_LUT4AB/S4END[4] Tile_X2Y6_LUT4AB/S4END[5]
+ Tile_X2Y6_LUT4AB/S4END[6] Tile_X2Y6_LUT4AB/S4END[7] Tile_X2Y6_LUT4AB/S4END[8] Tile_X2Y6_LUT4AB/S4END[9]
+ Tile_X2Y7_LUT4AB/SS4END[0] Tile_X2Y7_LUT4AB/SS4END[10] Tile_X2Y7_LUT4AB/SS4END[11]
+ Tile_X2Y7_LUT4AB/SS4END[12] Tile_X2Y7_LUT4AB/SS4END[13] Tile_X2Y7_LUT4AB/SS4END[14]
+ Tile_X2Y7_LUT4AB/SS4END[15] Tile_X2Y7_LUT4AB/SS4END[1] Tile_X2Y7_LUT4AB/SS4END[2]
+ Tile_X2Y7_LUT4AB/SS4END[3] Tile_X2Y7_LUT4AB/SS4END[4] Tile_X2Y7_LUT4AB/SS4END[5]
+ Tile_X2Y7_LUT4AB/SS4END[6] Tile_X2Y7_LUT4AB/SS4END[7] Tile_X2Y7_LUT4AB/SS4END[8]
+ Tile_X2Y7_LUT4AB/SS4END[9] Tile_X2Y6_LUT4AB/SS4END[0] Tile_X2Y6_LUT4AB/SS4END[10]
+ Tile_X2Y6_LUT4AB/SS4END[11] Tile_X2Y6_LUT4AB/SS4END[12] Tile_X2Y6_LUT4AB/SS4END[13]
+ Tile_X2Y6_LUT4AB/SS4END[14] Tile_X2Y6_LUT4AB/SS4END[15] Tile_X2Y6_LUT4AB/SS4END[1]
+ Tile_X2Y6_LUT4AB/SS4END[2] Tile_X2Y6_LUT4AB/SS4END[3] Tile_X2Y6_LUT4AB/SS4END[4]
+ Tile_X2Y6_LUT4AB/SS4END[5] Tile_X2Y6_LUT4AB/SS4END[6] Tile_X2Y6_LUT4AB/SS4END[7]
+ Tile_X2Y6_LUT4AB/SS4END[8] Tile_X2Y6_LUT4AB/SS4END[9] Tile_X2Y6_LUT4AB/UserCLK Tile_X2Y5_LUT4AB/UserCLK
+ VGND VPWR Tile_X2Y6_LUT4AB/W1BEG[0] Tile_X2Y6_LUT4AB/W1BEG[1] Tile_X2Y6_LUT4AB/W1BEG[2]
+ Tile_X2Y6_LUT4AB/W1BEG[3] Tile_X3Y6_LUT4AB/W1BEG[0] Tile_X3Y6_LUT4AB/W1BEG[1] Tile_X3Y6_LUT4AB/W1BEG[2]
+ Tile_X3Y6_LUT4AB/W1BEG[3] Tile_X2Y6_LUT4AB/W2BEG[0] Tile_X2Y6_LUT4AB/W2BEG[1] Tile_X2Y6_LUT4AB/W2BEG[2]
+ Tile_X2Y6_LUT4AB/W2BEG[3] Tile_X2Y6_LUT4AB/W2BEG[4] Tile_X2Y6_LUT4AB/W2BEG[5] Tile_X2Y6_LUT4AB/W2BEG[6]
+ Tile_X2Y6_LUT4AB/W2BEG[7] Tile_X1Y6_LUT4AB/W2END[0] Tile_X1Y6_LUT4AB/W2END[1] Tile_X1Y6_LUT4AB/W2END[2]
+ Tile_X1Y6_LUT4AB/W2END[3] Tile_X1Y6_LUT4AB/W2END[4] Tile_X1Y6_LUT4AB/W2END[5] Tile_X1Y6_LUT4AB/W2END[6]
+ Tile_X1Y6_LUT4AB/W2END[7] Tile_X2Y6_LUT4AB/W2END[0] Tile_X2Y6_LUT4AB/W2END[1] Tile_X2Y6_LUT4AB/W2END[2]
+ Tile_X2Y6_LUT4AB/W2END[3] Tile_X2Y6_LUT4AB/W2END[4] Tile_X2Y6_LUT4AB/W2END[5] Tile_X2Y6_LUT4AB/W2END[6]
+ Tile_X2Y6_LUT4AB/W2END[7] Tile_X3Y6_LUT4AB/W2BEG[0] Tile_X3Y6_LUT4AB/W2BEG[1] Tile_X3Y6_LUT4AB/W2BEG[2]
+ Tile_X3Y6_LUT4AB/W2BEG[3] Tile_X3Y6_LUT4AB/W2BEG[4] Tile_X3Y6_LUT4AB/W2BEG[5] Tile_X3Y6_LUT4AB/W2BEG[6]
+ Tile_X3Y6_LUT4AB/W2BEG[7] Tile_X2Y6_LUT4AB/W6BEG[0] Tile_X2Y6_LUT4AB/W6BEG[10] Tile_X2Y6_LUT4AB/W6BEG[11]
+ Tile_X2Y6_LUT4AB/W6BEG[1] Tile_X2Y6_LUT4AB/W6BEG[2] Tile_X2Y6_LUT4AB/W6BEG[3] Tile_X2Y6_LUT4AB/W6BEG[4]
+ Tile_X2Y6_LUT4AB/W6BEG[5] Tile_X2Y6_LUT4AB/W6BEG[6] Tile_X2Y6_LUT4AB/W6BEG[7] Tile_X2Y6_LUT4AB/W6BEG[8]
+ Tile_X2Y6_LUT4AB/W6BEG[9] Tile_X3Y6_LUT4AB/W6BEG[0] Tile_X3Y6_LUT4AB/W6BEG[10] Tile_X3Y6_LUT4AB/W6BEG[11]
+ Tile_X3Y6_LUT4AB/W6BEG[1] Tile_X3Y6_LUT4AB/W6BEG[2] Tile_X3Y6_LUT4AB/W6BEG[3] Tile_X3Y6_LUT4AB/W6BEG[4]
+ Tile_X3Y6_LUT4AB/W6BEG[5] Tile_X3Y6_LUT4AB/W6BEG[6] Tile_X3Y6_LUT4AB/W6BEG[7] Tile_X3Y6_LUT4AB/W6BEG[8]
+ Tile_X3Y6_LUT4AB/W6BEG[9] Tile_X2Y6_LUT4AB/WW4BEG[0] Tile_X2Y6_LUT4AB/WW4BEG[10]
+ Tile_X2Y6_LUT4AB/WW4BEG[11] Tile_X2Y6_LUT4AB/WW4BEG[12] Tile_X2Y6_LUT4AB/WW4BEG[13]
+ Tile_X2Y6_LUT4AB/WW4BEG[14] Tile_X2Y6_LUT4AB/WW4BEG[15] Tile_X2Y6_LUT4AB/WW4BEG[1]
+ Tile_X2Y6_LUT4AB/WW4BEG[2] Tile_X2Y6_LUT4AB/WW4BEG[3] Tile_X2Y6_LUT4AB/WW4BEG[4]
+ Tile_X2Y6_LUT4AB/WW4BEG[5] Tile_X2Y6_LUT4AB/WW4BEG[6] Tile_X2Y6_LUT4AB/WW4BEG[7]
+ Tile_X2Y6_LUT4AB/WW4BEG[8] Tile_X2Y6_LUT4AB/WW4BEG[9] Tile_X3Y6_LUT4AB/WW4BEG[0]
+ Tile_X3Y6_LUT4AB/WW4BEG[10] Tile_X3Y6_LUT4AB/WW4BEG[11] Tile_X3Y6_LUT4AB/WW4BEG[12]
+ Tile_X3Y6_LUT4AB/WW4BEG[13] Tile_X3Y6_LUT4AB/WW4BEG[14] Tile_X3Y6_LUT4AB/WW4BEG[15]
+ Tile_X3Y6_LUT4AB/WW4BEG[1] Tile_X3Y6_LUT4AB/WW4BEG[2] Tile_X3Y6_LUT4AB/WW4BEG[3]
+ Tile_X3Y6_LUT4AB/WW4BEG[4] Tile_X3Y6_LUT4AB/WW4BEG[5] Tile_X3Y6_LUT4AB/WW4BEG[6]
+ Tile_X3Y6_LUT4AB/WW4BEG[7] Tile_X3Y6_LUT4AB/WW4BEG[8] Tile_X3Y6_LUT4AB/WW4BEG[9]
+ LUT4AB
XTile_X5Y12_LUT4AB Tile_X5Y13_LUT4AB/Co Tile_X5Y12_LUT4AB/Co Tile_X6Y12_LUT4AB/E1END[0]
+ Tile_X6Y12_LUT4AB/E1END[1] Tile_X6Y12_LUT4AB/E1END[2] Tile_X6Y12_LUT4AB/E1END[3]
+ Tile_X5Y12_LUT4AB/E1END[0] Tile_X5Y12_LUT4AB/E1END[1] Tile_X5Y12_LUT4AB/E1END[2]
+ Tile_X5Y12_LUT4AB/E1END[3] Tile_X6Y12_LUT4AB/E2MID[0] Tile_X6Y12_LUT4AB/E2MID[1]
+ Tile_X6Y12_LUT4AB/E2MID[2] Tile_X6Y12_LUT4AB/E2MID[3] Tile_X6Y12_LUT4AB/E2MID[4]
+ Tile_X6Y12_LUT4AB/E2MID[5] Tile_X6Y12_LUT4AB/E2MID[6] Tile_X6Y12_LUT4AB/E2MID[7]
+ Tile_X6Y12_LUT4AB/E2END[0] Tile_X6Y12_LUT4AB/E2END[1] Tile_X6Y12_LUT4AB/E2END[2]
+ Tile_X6Y12_LUT4AB/E2END[3] Tile_X6Y12_LUT4AB/E2END[4] Tile_X6Y12_LUT4AB/E2END[5]
+ Tile_X6Y12_LUT4AB/E2END[6] Tile_X6Y12_LUT4AB/E2END[7] Tile_X5Y12_LUT4AB/E2END[0]
+ Tile_X5Y12_LUT4AB/E2END[1] Tile_X5Y12_LUT4AB/E2END[2] Tile_X5Y12_LUT4AB/E2END[3]
+ Tile_X5Y12_LUT4AB/E2END[4] Tile_X5Y12_LUT4AB/E2END[5] Tile_X5Y12_LUT4AB/E2END[6]
+ Tile_X5Y12_LUT4AB/E2END[7] Tile_X5Y12_LUT4AB/E2MID[0] Tile_X5Y12_LUT4AB/E2MID[1]
+ Tile_X5Y12_LUT4AB/E2MID[2] Tile_X5Y12_LUT4AB/E2MID[3] Tile_X5Y12_LUT4AB/E2MID[4]
+ Tile_X5Y12_LUT4AB/E2MID[5] Tile_X5Y12_LUT4AB/E2MID[6] Tile_X5Y12_LUT4AB/E2MID[7]
+ Tile_X6Y12_LUT4AB/E6END[0] Tile_X6Y12_LUT4AB/E6END[10] Tile_X6Y12_LUT4AB/E6END[11]
+ Tile_X6Y12_LUT4AB/E6END[1] Tile_X6Y12_LUT4AB/E6END[2] Tile_X6Y12_LUT4AB/E6END[3]
+ Tile_X6Y12_LUT4AB/E6END[4] Tile_X6Y12_LUT4AB/E6END[5] Tile_X6Y12_LUT4AB/E6END[6]
+ Tile_X6Y12_LUT4AB/E6END[7] Tile_X6Y12_LUT4AB/E6END[8] Tile_X6Y12_LUT4AB/E6END[9]
+ Tile_X5Y12_LUT4AB/E6END[0] Tile_X5Y12_LUT4AB/E6END[10] Tile_X5Y12_LUT4AB/E6END[11]
+ Tile_X5Y12_LUT4AB/E6END[1] Tile_X5Y12_LUT4AB/E6END[2] Tile_X5Y12_LUT4AB/E6END[3]
+ Tile_X5Y12_LUT4AB/E6END[4] Tile_X5Y12_LUT4AB/E6END[5] Tile_X5Y12_LUT4AB/E6END[6]
+ Tile_X5Y12_LUT4AB/E6END[7] Tile_X5Y12_LUT4AB/E6END[8] Tile_X5Y12_LUT4AB/E6END[9]
+ Tile_X6Y12_LUT4AB/EE4END[0] Tile_X6Y12_LUT4AB/EE4END[10] Tile_X6Y12_LUT4AB/EE4END[11]
+ Tile_X6Y12_LUT4AB/EE4END[12] Tile_X6Y12_LUT4AB/EE4END[13] Tile_X6Y12_LUT4AB/EE4END[14]
+ Tile_X6Y12_LUT4AB/EE4END[15] Tile_X6Y12_LUT4AB/EE4END[1] Tile_X6Y12_LUT4AB/EE4END[2]
+ Tile_X6Y12_LUT4AB/EE4END[3] Tile_X6Y12_LUT4AB/EE4END[4] Tile_X6Y12_LUT4AB/EE4END[5]
+ Tile_X6Y12_LUT4AB/EE4END[6] Tile_X6Y12_LUT4AB/EE4END[7] Tile_X6Y12_LUT4AB/EE4END[8]
+ Tile_X6Y12_LUT4AB/EE4END[9] Tile_X5Y12_LUT4AB/EE4END[0] Tile_X5Y12_LUT4AB/EE4END[10]
+ Tile_X5Y12_LUT4AB/EE4END[11] Tile_X5Y12_LUT4AB/EE4END[12] Tile_X5Y12_LUT4AB/EE4END[13]
+ Tile_X5Y12_LUT4AB/EE4END[14] Tile_X5Y12_LUT4AB/EE4END[15] Tile_X5Y12_LUT4AB/EE4END[1]
+ Tile_X5Y12_LUT4AB/EE4END[2] Tile_X5Y12_LUT4AB/EE4END[3] Tile_X5Y12_LUT4AB/EE4END[4]
+ Tile_X5Y12_LUT4AB/EE4END[5] Tile_X5Y12_LUT4AB/EE4END[6] Tile_X5Y12_LUT4AB/EE4END[7]
+ Tile_X5Y12_LUT4AB/EE4END[8] Tile_X5Y12_LUT4AB/EE4END[9] Tile_X5Y12_LUT4AB/FrameData[0]
+ Tile_X5Y12_LUT4AB/FrameData[10] Tile_X5Y12_LUT4AB/FrameData[11] Tile_X5Y12_LUT4AB/FrameData[12]
+ Tile_X5Y12_LUT4AB/FrameData[13] Tile_X5Y12_LUT4AB/FrameData[14] Tile_X5Y12_LUT4AB/FrameData[15]
+ Tile_X5Y12_LUT4AB/FrameData[16] Tile_X5Y12_LUT4AB/FrameData[17] Tile_X5Y12_LUT4AB/FrameData[18]
+ Tile_X5Y12_LUT4AB/FrameData[19] Tile_X5Y12_LUT4AB/FrameData[1] Tile_X5Y12_LUT4AB/FrameData[20]
+ Tile_X5Y12_LUT4AB/FrameData[21] Tile_X5Y12_LUT4AB/FrameData[22] Tile_X5Y12_LUT4AB/FrameData[23]
+ Tile_X5Y12_LUT4AB/FrameData[24] Tile_X5Y12_LUT4AB/FrameData[25] Tile_X5Y12_LUT4AB/FrameData[26]
+ Tile_X5Y12_LUT4AB/FrameData[27] Tile_X5Y12_LUT4AB/FrameData[28] Tile_X5Y12_LUT4AB/FrameData[29]
+ Tile_X5Y12_LUT4AB/FrameData[2] Tile_X5Y12_LUT4AB/FrameData[30] Tile_X5Y12_LUT4AB/FrameData[31]
+ Tile_X5Y12_LUT4AB/FrameData[3] Tile_X5Y12_LUT4AB/FrameData[4] Tile_X5Y12_LUT4AB/FrameData[5]
+ Tile_X5Y12_LUT4AB/FrameData[6] Tile_X5Y12_LUT4AB/FrameData[7] Tile_X5Y12_LUT4AB/FrameData[8]
+ Tile_X5Y12_LUT4AB/FrameData[9] Tile_X6Y12_LUT4AB/FrameData[0] Tile_X6Y12_LUT4AB/FrameData[10]
+ Tile_X6Y12_LUT4AB/FrameData[11] Tile_X6Y12_LUT4AB/FrameData[12] Tile_X6Y12_LUT4AB/FrameData[13]
+ Tile_X6Y12_LUT4AB/FrameData[14] Tile_X6Y12_LUT4AB/FrameData[15] Tile_X6Y12_LUT4AB/FrameData[16]
+ Tile_X6Y12_LUT4AB/FrameData[17] Tile_X6Y12_LUT4AB/FrameData[18] Tile_X6Y12_LUT4AB/FrameData[19]
+ Tile_X6Y12_LUT4AB/FrameData[1] Tile_X6Y12_LUT4AB/FrameData[20] Tile_X6Y12_LUT4AB/FrameData[21]
+ Tile_X6Y12_LUT4AB/FrameData[22] Tile_X6Y12_LUT4AB/FrameData[23] Tile_X6Y12_LUT4AB/FrameData[24]
+ Tile_X6Y12_LUT4AB/FrameData[25] Tile_X6Y12_LUT4AB/FrameData[26] Tile_X6Y12_LUT4AB/FrameData[27]
+ Tile_X6Y12_LUT4AB/FrameData[28] Tile_X6Y12_LUT4AB/FrameData[29] Tile_X6Y12_LUT4AB/FrameData[2]
+ Tile_X6Y12_LUT4AB/FrameData[30] Tile_X6Y12_LUT4AB/FrameData[31] Tile_X6Y12_LUT4AB/FrameData[3]
+ Tile_X6Y12_LUT4AB/FrameData[4] Tile_X6Y12_LUT4AB/FrameData[5] Tile_X6Y12_LUT4AB/FrameData[6]
+ Tile_X6Y12_LUT4AB/FrameData[7] Tile_X6Y12_LUT4AB/FrameData[8] Tile_X6Y12_LUT4AB/FrameData[9]
+ Tile_X5Y12_LUT4AB/FrameStrobe[0] Tile_X5Y12_LUT4AB/FrameStrobe[10] Tile_X5Y12_LUT4AB/FrameStrobe[11]
+ Tile_X5Y12_LUT4AB/FrameStrobe[12] Tile_X5Y12_LUT4AB/FrameStrobe[13] Tile_X5Y12_LUT4AB/FrameStrobe[14]
+ Tile_X5Y12_LUT4AB/FrameStrobe[15] Tile_X5Y12_LUT4AB/FrameStrobe[16] Tile_X5Y12_LUT4AB/FrameStrobe[17]
+ Tile_X5Y12_LUT4AB/FrameStrobe[18] Tile_X5Y12_LUT4AB/FrameStrobe[19] Tile_X5Y12_LUT4AB/FrameStrobe[1]
+ Tile_X5Y12_LUT4AB/FrameStrobe[2] Tile_X5Y12_LUT4AB/FrameStrobe[3] Tile_X5Y12_LUT4AB/FrameStrobe[4]
+ Tile_X5Y12_LUT4AB/FrameStrobe[5] Tile_X5Y12_LUT4AB/FrameStrobe[6] Tile_X5Y12_LUT4AB/FrameStrobe[7]
+ Tile_X5Y12_LUT4AB/FrameStrobe[8] Tile_X5Y12_LUT4AB/FrameStrobe[9] Tile_X5Y11_LUT4AB/FrameStrobe[0]
+ Tile_X5Y11_LUT4AB/FrameStrobe[10] Tile_X5Y11_LUT4AB/FrameStrobe[11] Tile_X5Y11_LUT4AB/FrameStrobe[12]
+ Tile_X5Y11_LUT4AB/FrameStrobe[13] Tile_X5Y11_LUT4AB/FrameStrobe[14] Tile_X5Y11_LUT4AB/FrameStrobe[15]
+ Tile_X5Y11_LUT4AB/FrameStrobe[16] Tile_X5Y11_LUT4AB/FrameStrobe[17] Tile_X5Y11_LUT4AB/FrameStrobe[18]
+ Tile_X5Y11_LUT4AB/FrameStrobe[19] Tile_X5Y11_LUT4AB/FrameStrobe[1] Tile_X5Y11_LUT4AB/FrameStrobe[2]
+ Tile_X5Y11_LUT4AB/FrameStrobe[3] Tile_X5Y11_LUT4AB/FrameStrobe[4] Tile_X5Y11_LUT4AB/FrameStrobe[5]
+ Tile_X5Y11_LUT4AB/FrameStrobe[6] Tile_X5Y11_LUT4AB/FrameStrobe[7] Tile_X5Y11_LUT4AB/FrameStrobe[8]
+ Tile_X5Y11_LUT4AB/FrameStrobe[9] Tile_X5Y12_LUT4AB/N1BEG[0] Tile_X5Y12_LUT4AB/N1BEG[1]
+ Tile_X5Y12_LUT4AB/N1BEG[2] Tile_X5Y12_LUT4AB/N1BEG[3] Tile_X5Y13_LUT4AB/N1BEG[0]
+ Tile_X5Y13_LUT4AB/N1BEG[1] Tile_X5Y13_LUT4AB/N1BEG[2] Tile_X5Y13_LUT4AB/N1BEG[3]
+ Tile_X5Y12_LUT4AB/N2BEG[0] Tile_X5Y12_LUT4AB/N2BEG[1] Tile_X5Y12_LUT4AB/N2BEG[2]
+ Tile_X5Y12_LUT4AB/N2BEG[3] Tile_X5Y12_LUT4AB/N2BEG[4] Tile_X5Y12_LUT4AB/N2BEG[5]
+ Tile_X5Y12_LUT4AB/N2BEG[6] Tile_X5Y12_LUT4AB/N2BEG[7] Tile_X5Y11_LUT4AB/N2END[0]
+ Tile_X5Y11_LUT4AB/N2END[1] Tile_X5Y11_LUT4AB/N2END[2] Tile_X5Y11_LUT4AB/N2END[3]
+ Tile_X5Y11_LUT4AB/N2END[4] Tile_X5Y11_LUT4AB/N2END[5] Tile_X5Y11_LUT4AB/N2END[6]
+ Tile_X5Y11_LUT4AB/N2END[7] Tile_X5Y12_LUT4AB/N2END[0] Tile_X5Y12_LUT4AB/N2END[1]
+ Tile_X5Y12_LUT4AB/N2END[2] Tile_X5Y12_LUT4AB/N2END[3] Tile_X5Y12_LUT4AB/N2END[4]
+ Tile_X5Y12_LUT4AB/N2END[5] Tile_X5Y12_LUT4AB/N2END[6] Tile_X5Y12_LUT4AB/N2END[7]
+ Tile_X5Y13_LUT4AB/N2BEG[0] Tile_X5Y13_LUT4AB/N2BEG[1] Tile_X5Y13_LUT4AB/N2BEG[2]
+ Tile_X5Y13_LUT4AB/N2BEG[3] Tile_X5Y13_LUT4AB/N2BEG[4] Tile_X5Y13_LUT4AB/N2BEG[5]
+ Tile_X5Y13_LUT4AB/N2BEG[6] Tile_X5Y13_LUT4AB/N2BEG[7] Tile_X5Y12_LUT4AB/N4BEG[0]
+ Tile_X5Y12_LUT4AB/N4BEG[10] Tile_X5Y12_LUT4AB/N4BEG[11] Tile_X5Y12_LUT4AB/N4BEG[12]
+ Tile_X5Y12_LUT4AB/N4BEG[13] Tile_X5Y12_LUT4AB/N4BEG[14] Tile_X5Y12_LUT4AB/N4BEG[15]
+ Tile_X5Y12_LUT4AB/N4BEG[1] Tile_X5Y12_LUT4AB/N4BEG[2] Tile_X5Y12_LUT4AB/N4BEG[3]
+ Tile_X5Y12_LUT4AB/N4BEG[4] Tile_X5Y12_LUT4AB/N4BEG[5] Tile_X5Y12_LUT4AB/N4BEG[6]
+ Tile_X5Y12_LUT4AB/N4BEG[7] Tile_X5Y12_LUT4AB/N4BEG[8] Tile_X5Y12_LUT4AB/N4BEG[9]
+ Tile_X5Y13_LUT4AB/N4BEG[0] Tile_X5Y13_LUT4AB/N4BEG[10] Tile_X5Y13_LUT4AB/N4BEG[11]
+ Tile_X5Y13_LUT4AB/N4BEG[12] Tile_X5Y13_LUT4AB/N4BEG[13] Tile_X5Y13_LUT4AB/N4BEG[14]
+ Tile_X5Y13_LUT4AB/N4BEG[15] Tile_X5Y13_LUT4AB/N4BEG[1] Tile_X5Y13_LUT4AB/N4BEG[2]
+ Tile_X5Y13_LUT4AB/N4BEG[3] Tile_X5Y13_LUT4AB/N4BEG[4] Tile_X5Y13_LUT4AB/N4BEG[5]
+ Tile_X5Y13_LUT4AB/N4BEG[6] Tile_X5Y13_LUT4AB/N4BEG[7] Tile_X5Y13_LUT4AB/N4BEG[8]
+ Tile_X5Y13_LUT4AB/N4BEG[9] Tile_X5Y12_LUT4AB/NN4BEG[0] Tile_X5Y12_LUT4AB/NN4BEG[10]
+ Tile_X5Y12_LUT4AB/NN4BEG[11] Tile_X5Y12_LUT4AB/NN4BEG[12] Tile_X5Y12_LUT4AB/NN4BEG[13]
+ Tile_X5Y12_LUT4AB/NN4BEG[14] Tile_X5Y12_LUT4AB/NN4BEG[15] Tile_X5Y12_LUT4AB/NN4BEG[1]
+ Tile_X5Y12_LUT4AB/NN4BEG[2] Tile_X5Y12_LUT4AB/NN4BEG[3] Tile_X5Y12_LUT4AB/NN4BEG[4]
+ Tile_X5Y12_LUT4AB/NN4BEG[5] Tile_X5Y12_LUT4AB/NN4BEG[6] Tile_X5Y12_LUT4AB/NN4BEG[7]
+ Tile_X5Y12_LUT4AB/NN4BEG[8] Tile_X5Y12_LUT4AB/NN4BEG[9] Tile_X5Y13_LUT4AB/NN4BEG[0]
+ Tile_X5Y13_LUT4AB/NN4BEG[10] Tile_X5Y13_LUT4AB/NN4BEG[11] Tile_X5Y13_LUT4AB/NN4BEG[12]
+ Tile_X5Y13_LUT4AB/NN4BEG[13] Tile_X5Y13_LUT4AB/NN4BEG[14] Tile_X5Y13_LUT4AB/NN4BEG[15]
+ Tile_X5Y13_LUT4AB/NN4BEG[1] Tile_X5Y13_LUT4AB/NN4BEG[2] Tile_X5Y13_LUT4AB/NN4BEG[3]
+ Tile_X5Y13_LUT4AB/NN4BEG[4] Tile_X5Y13_LUT4AB/NN4BEG[5] Tile_X5Y13_LUT4AB/NN4BEG[6]
+ Tile_X5Y13_LUT4AB/NN4BEG[7] Tile_X5Y13_LUT4AB/NN4BEG[8] Tile_X5Y13_LUT4AB/NN4BEG[9]
+ Tile_X5Y13_LUT4AB/S1END[0] Tile_X5Y13_LUT4AB/S1END[1] Tile_X5Y13_LUT4AB/S1END[2]
+ Tile_X5Y13_LUT4AB/S1END[3] Tile_X5Y12_LUT4AB/S1END[0] Tile_X5Y12_LUT4AB/S1END[1]
+ Tile_X5Y12_LUT4AB/S1END[2] Tile_X5Y12_LUT4AB/S1END[3] Tile_X5Y13_LUT4AB/S2MID[0]
+ Tile_X5Y13_LUT4AB/S2MID[1] Tile_X5Y13_LUT4AB/S2MID[2] Tile_X5Y13_LUT4AB/S2MID[3]
+ Tile_X5Y13_LUT4AB/S2MID[4] Tile_X5Y13_LUT4AB/S2MID[5] Tile_X5Y13_LUT4AB/S2MID[6]
+ Tile_X5Y13_LUT4AB/S2MID[7] Tile_X5Y13_LUT4AB/S2END[0] Tile_X5Y13_LUT4AB/S2END[1]
+ Tile_X5Y13_LUT4AB/S2END[2] Tile_X5Y13_LUT4AB/S2END[3] Tile_X5Y13_LUT4AB/S2END[4]
+ Tile_X5Y13_LUT4AB/S2END[5] Tile_X5Y13_LUT4AB/S2END[6] Tile_X5Y13_LUT4AB/S2END[7]
+ Tile_X5Y12_LUT4AB/S2END[0] Tile_X5Y12_LUT4AB/S2END[1] Tile_X5Y12_LUT4AB/S2END[2]
+ Tile_X5Y12_LUT4AB/S2END[3] Tile_X5Y12_LUT4AB/S2END[4] Tile_X5Y12_LUT4AB/S2END[5]
+ Tile_X5Y12_LUT4AB/S2END[6] Tile_X5Y12_LUT4AB/S2END[7] Tile_X5Y12_LUT4AB/S2MID[0]
+ Tile_X5Y12_LUT4AB/S2MID[1] Tile_X5Y12_LUT4AB/S2MID[2] Tile_X5Y12_LUT4AB/S2MID[3]
+ Tile_X5Y12_LUT4AB/S2MID[4] Tile_X5Y12_LUT4AB/S2MID[5] Tile_X5Y12_LUT4AB/S2MID[6]
+ Tile_X5Y12_LUT4AB/S2MID[7] Tile_X5Y13_LUT4AB/S4END[0] Tile_X5Y13_LUT4AB/S4END[10]
+ Tile_X5Y13_LUT4AB/S4END[11] Tile_X5Y13_LUT4AB/S4END[12] Tile_X5Y13_LUT4AB/S4END[13]
+ Tile_X5Y13_LUT4AB/S4END[14] Tile_X5Y13_LUT4AB/S4END[15] Tile_X5Y13_LUT4AB/S4END[1]
+ Tile_X5Y13_LUT4AB/S4END[2] Tile_X5Y13_LUT4AB/S4END[3] Tile_X5Y13_LUT4AB/S4END[4]
+ Tile_X5Y13_LUT4AB/S4END[5] Tile_X5Y13_LUT4AB/S4END[6] Tile_X5Y13_LUT4AB/S4END[7]
+ Tile_X5Y13_LUT4AB/S4END[8] Tile_X5Y13_LUT4AB/S4END[9] Tile_X5Y12_LUT4AB/S4END[0]
+ Tile_X5Y12_LUT4AB/S4END[10] Tile_X5Y12_LUT4AB/S4END[11] Tile_X5Y12_LUT4AB/S4END[12]
+ Tile_X5Y12_LUT4AB/S4END[13] Tile_X5Y12_LUT4AB/S4END[14] Tile_X5Y12_LUT4AB/S4END[15]
+ Tile_X5Y12_LUT4AB/S4END[1] Tile_X5Y12_LUT4AB/S4END[2] Tile_X5Y12_LUT4AB/S4END[3]
+ Tile_X5Y12_LUT4AB/S4END[4] Tile_X5Y12_LUT4AB/S4END[5] Tile_X5Y12_LUT4AB/S4END[6]
+ Tile_X5Y12_LUT4AB/S4END[7] Tile_X5Y12_LUT4AB/S4END[8] Tile_X5Y12_LUT4AB/S4END[9]
+ Tile_X5Y13_LUT4AB/SS4END[0] Tile_X5Y13_LUT4AB/SS4END[10] Tile_X5Y13_LUT4AB/SS4END[11]
+ Tile_X5Y13_LUT4AB/SS4END[12] Tile_X5Y13_LUT4AB/SS4END[13] Tile_X5Y13_LUT4AB/SS4END[14]
+ Tile_X5Y13_LUT4AB/SS4END[15] Tile_X5Y13_LUT4AB/SS4END[1] Tile_X5Y13_LUT4AB/SS4END[2]
+ Tile_X5Y13_LUT4AB/SS4END[3] Tile_X5Y13_LUT4AB/SS4END[4] Tile_X5Y13_LUT4AB/SS4END[5]
+ Tile_X5Y13_LUT4AB/SS4END[6] Tile_X5Y13_LUT4AB/SS4END[7] Tile_X5Y13_LUT4AB/SS4END[8]
+ Tile_X5Y13_LUT4AB/SS4END[9] Tile_X5Y12_LUT4AB/SS4END[0] Tile_X5Y12_LUT4AB/SS4END[10]
+ Tile_X5Y12_LUT4AB/SS4END[11] Tile_X5Y12_LUT4AB/SS4END[12] Tile_X5Y12_LUT4AB/SS4END[13]
+ Tile_X5Y12_LUT4AB/SS4END[14] Tile_X5Y12_LUT4AB/SS4END[15] Tile_X5Y12_LUT4AB/SS4END[1]
+ Tile_X5Y12_LUT4AB/SS4END[2] Tile_X5Y12_LUT4AB/SS4END[3] Tile_X5Y12_LUT4AB/SS4END[4]
+ Tile_X5Y12_LUT4AB/SS4END[5] Tile_X5Y12_LUT4AB/SS4END[6] Tile_X5Y12_LUT4AB/SS4END[7]
+ Tile_X5Y12_LUT4AB/SS4END[8] Tile_X5Y12_LUT4AB/SS4END[9] Tile_X5Y12_LUT4AB/UserCLK
+ Tile_X5Y11_LUT4AB/UserCLK VGND VPWR Tile_X5Y12_LUT4AB/W1BEG[0] Tile_X5Y12_LUT4AB/W1BEG[1]
+ Tile_X5Y12_LUT4AB/W1BEG[2] Tile_X5Y12_LUT4AB/W1BEG[3] Tile_X6Y12_LUT4AB/W1BEG[0]
+ Tile_X6Y12_LUT4AB/W1BEG[1] Tile_X6Y12_LUT4AB/W1BEG[2] Tile_X6Y12_LUT4AB/W1BEG[3]
+ Tile_X5Y12_LUT4AB/W2BEG[0] Tile_X5Y12_LUT4AB/W2BEG[1] Tile_X5Y12_LUT4AB/W2BEG[2]
+ Tile_X5Y12_LUT4AB/W2BEG[3] Tile_X5Y12_LUT4AB/W2BEG[4] Tile_X5Y12_LUT4AB/W2BEG[5]
+ Tile_X5Y12_LUT4AB/W2BEG[6] Tile_X5Y12_LUT4AB/W2BEG[7] Tile_X5Y12_LUT4AB/W2BEGb[0]
+ Tile_X5Y12_LUT4AB/W2BEGb[1] Tile_X5Y12_LUT4AB/W2BEGb[2] Tile_X5Y12_LUT4AB/W2BEGb[3]
+ Tile_X5Y12_LUT4AB/W2BEGb[4] Tile_X5Y12_LUT4AB/W2BEGb[5] Tile_X5Y12_LUT4AB/W2BEGb[6]
+ Tile_X5Y12_LUT4AB/W2BEGb[7] Tile_X5Y12_LUT4AB/W2END[0] Tile_X5Y12_LUT4AB/W2END[1]
+ Tile_X5Y12_LUT4AB/W2END[2] Tile_X5Y12_LUT4AB/W2END[3] Tile_X5Y12_LUT4AB/W2END[4]
+ Tile_X5Y12_LUT4AB/W2END[5] Tile_X5Y12_LUT4AB/W2END[6] Tile_X5Y12_LUT4AB/W2END[7]
+ Tile_X6Y12_LUT4AB/W2BEG[0] Tile_X6Y12_LUT4AB/W2BEG[1] Tile_X6Y12_LUT4AB/W2BEG[2]
+ Tile_X6Y12_LUT4AB/W2BEG[3] Tile_X6Y12_LUT4AB/W2BEG[4] Tile_X6Y12_LUT4AB/W2BEG[5]
+ Tile_X6Y12_LUT4AB/W2BEG[6] Tile_X6Y12_LUT4AB/W2BEG[7] Tile_X5Y12_LUT4AB/W6BEG[0]
+ Tile_X5Y12_LUT4AB/W6BEG[10] Tile_X5Y12_LUT4AB/W6BEG[11] Tile_X5Y12_LUT4AB/W6BEG[1]
+ Tile_X5Y12_LUT4AB/W6BEG[2] Tile_X5Y12_LUT4AB/W6BEG[3] Tile_X5Y12_LUT4AB/W6BEG[4]
+ Tile_X5Y12_LUT4AB/W6BEG[5] Tile_X5Y12_LUT4AB/W6BEG[6] Tile_X5Y12_LUT4AB/W6BEG[7]
+ Tile_X5Y12_LUT4AB/W6BEG[8] Tile_X5Y12_LUT4AB/W6BEG[9] Tile_X6Y12_LUT4AB/W6BEG[0]
+ Tile_X6Y12_LUT4AB/W6BEG[10] Tile_X6Y12_LUT4AB/W6BEG[11] Tile_X6Y12_LUT4AB/W6BEG[1]
+ Tile_X6Y12_LUT4AB/W6BEG[2] Tile_X6Y12_LUT4AB/W6BEG[3] Tile_X6Y12_LUT4AB/W6BEG[4]
+ Tile_X6Y12_LUT4AB/W6BEG[5] Tile_X6Y12_LUT4AB/W6BEG[6] Tile_X6Y12_LUT4AB/W6BEG[7]
+ Tile_X6Y12_LUT4AB/W6BEG[8] Tile_X6Y12_LUT4AB/W6BEG[9] Tile_X5Y12_LUT4AB/WW4BEG[0]
+ Tile_X5Y12_LUT4AB/WW4BEG[10] Tile_X5Y12_LUT4AB/WW4BEG[11] Tile_X5Y12_LUT4AB/WW4BEG[12]
+ Tile_X5Y12_LUT4AB/WW4BEG[13] Tile_X5Y12_LUT4AB/WW4BEG[14] Tile_X5Y12_LUT4AB/WW4BEG[15]
+ Tile_X5Y12_LUT4AB/WW4BEG[1] Tile_X5Y12_LUT4AB/WW4BEG[2] Tile_X5Y12_LUT4AB/WW4BEG[3]
+ Tile_X5Y12_LUT4AB/WW4BEG[4] Tile_X5Y12_LUT4AB/WW4BEG[5] Tile_X5Y12_LUT4AB/WW4BEG[6]
+ Tile_X5Y12_LUT4AB/WW4BEG[7] Tile_X5Y12_LUT4AB/WW4BEG[8] Tile_X5Y12_LUT4AB/WW4BEG[9]
+ Tile_X6Y12_LUT4AB/WW4BEG[0] Tile_X6Y12_LUT4AB/WW4BEG[10] Tile_X6Y12_LUT4AB/WW4BEG[11]
+ Tile_X6Y12_LUT4AB/WW4BEG[12] Tile_X6Y12_LUT4AB/WW4BEG[13] Tile_X6Y12_LUT4AB/WW4BEG[14]
+ Tile_X6Y12_LUT4AB/WW4BEG[15] Tile_X6Y12_LUT4AB/WW4BEG[1] Tile_X6Y12_LUT4AB/WW4BEG[2]
+ Tile_X6Y12_LUT4AB/WW4BEG[3] Tile_X6Y12_LUT4AB/WW4BEG[4] Tile_X6Y12_LUT4AB/WW4BEG[5]
+ Tile_X6Y12_LUT4AB/WW4BEG[6] Tile_X6Y12_LUT4AB/WW4BEG[7] Tile_X6Y12_LUT4AB/WW4BEG[8]
+ Tile_X6Y12_LUT4AB/WW4BEG[9] LUT4AB
XTile_X9Y1_LUT4AB Tile_X9Y2_LUT4AB/Co Tile_X9Y1_LUT4AB/Co Tile_X9Y1_LUT4AB/E1BEG[0]
+ Tile_X9Y1_LUT4AB/E1BEG[1] Tile_X9Y1_LUT4AB/E1BEG[2] Tile_X9Y1_LUT4AB/E1BEG[3] Tile_X9Y1_LUT4AB/E1END[0]
+ Tile_X9Y1_LUT4AB/E1END[1] Tile_X9Y1_LUT4AB/E1END[2] Tile_X9Y1_LUT4AB/E1END[3] Tile_X9Y1_LUT4AB/E2BEG[0]
+ Tile_X9Y1_LUT4AB/E2BEG[1] Tile_X9Y1_LUT4AB/E2BEG[2] Tile_X9Y1_LUT4AB/E2BEG[3] Tile_X9Y1_LUT4AB/E2BEG[4]
+ Tile_X9Y1_LUT4AB/E2BEG[5] Tile_X9Y1_LUT4AB/E2BEG[6] Tile_X9Y1_LUT4AB/E2BEG[7] Tile_X9Y1_LUT4AB/E2BEGb[0]
+ Tile_X9Y1_LUT4AB/E2BEGb[1] Tile_X9Y1_LUT4AB/E2BEGb[2] Tile_X9Y1_LUT4AB/E2BEGb[3]
+ Tile_X9Y1_LUT4AB/E2BEGb[4] Tile_X9Y1_LUT4AB/E2BEGb[5] Tile_X9Y1_LUT4AB/E2BEGb[6]
+ Tile_X9Y1_LUT4AB/E2BEGb[7] Tile_X9Y1_LUT4AB/E2END[0] Tile_X9Y1_LUT4AB/E2END[1] Tile_X9Y1_LUT4AB/E2END[2]
+ Tile_X9Y1_LUT4AB/E2END[3] Tile_X9Y1_LUT4AB/E2END[4] Tile_X9Y1_LUT4AB/E2END[5] Tile_X9Y1_LUT4AB/E2END[6]
+ Tile_X9Y1_LUT4AB/E2END[7] Tile_X9Y1_LUT4AB/E2MID[0] Tile_X9Y1_LUT4AB/E2MID[1] Tile_X9Y1_LUT4AB/E2MID[2]
+ Tile_X9Y1_LUT4AB/E2MID[3] Tile_X9Y1_LUT4AB/E2MID[4] Tile_X9Y1_LUT4AB/E2MID[5] Tile_X9Y1_LUT4AB/E2MID[6]
+ Tile_X9Y1_LUT4AB/E2MID[7] Tile_X9Y1_LUT4AB/E6BEG[0] Tile_X9Y1_LUT4AB/E6BEG[10] Tile_X9Y1_LUT4AB/E6BEG[11]
+ Tile_X9Y1_LUT4AB/E6BEG[1] Tile_X9Y1_LUT4AB/E6BEG[2] Tile_X9Y1_LUT4AB/E6BEG[3] Tile_X9Y1_LUT4AB/E6BEG[4]
+ Tile_X9Y1_LUT4AB/E6BEG[5] Tile_X9Y1_LUT4AB/E6BEG[6] Tile_X9Y1_LUT4AB/E6BEG[7] Tile_X9Y1_LUT4AB/E6BEG[8]
+ Tile_X9Y1_LUT4AB/E6BEG[9] Tile_X9Y1_LUT4AB/E6END[0] Tile_X9Y1_LUT4AB/E6END[10] Tile_X9Y1_LUT4AB/E6END[11]
+ Tile_X9Y1_LUT4AB/E6END[1] Tile_X9Y1_LUT4AB/E6END[2] Tile_X9Y1_LUT4AB/E6END[3] Tile_X9Y1_LUT4AB/E6END[4]
+ Tile_X9Y1_LUT4AB/E6END[5] Tile_X9Y1_LUT4AB/E6END[6] Tile_X9Y1_LUT4AB/E6END[7] Tile_X9Y1_LUT4AB/E6END[8]
+ Tile_X9Y1_LUT4AB/E6END[9] Tile_X9Y1_LUT4AB/EE4BEG[0] Tile_X9Y1_LUT4AB/EE4BEG[10]
+ Tile_X9Y1_LUT4AB/EE4BEG[11] Tile_X9Y1_LUT4AB/EE4BEG[12] Tile_X9Y1_LUT4AB/EE4BEG[13]
+ Tile_X9Y1_LUT4AB/EE4BEG[14] Tile_X9Y1_LUT4AB/EE4BEG[15] Tile_X9Y1_LUT4AB/EE4BEG[1]
+ Tile_X9Y1_LUT4AB/EE4BEG[2] Tile_X9Y1_LUT4AB/EE4BEG[3] Tile_X9Y1_LUT4AB/EE4BEG[4]
+ Tile_X9Y1_LUT4AB/EE4BEG[5] Tile_X9Y1_LUT4AB/EE4BEG[6] Tile_X9Y1_LUT4AB/EE4BEG[7]
+ Tile_X9Y1_LUT4AB/EE4BEG[8] Tile_X9Y1_LUT4AB/EE4BEG[9] Tile_X9Y1_LUT4AB/EE4END[0]
+ Tile_X9Y1_LUT4AB/EE4END[10] Tile_X9Y1_LUT4AB/EE4END[11] Tile_X9Y1_LUT4AB/EE4END[12]
+ Tile_X9Y1_LUT4AB/EE4END[13] Tile_X9Y1_LUT4AB/EE4END[14] Tile_X9Y1_LUT4AB/EE4END[15]
+ Tile_X9Y1_LUT4AB/EE4END[1] Tile_X9Y1_LUT4AB/EE4END[2] Tile_X9Y1_LUT4AB/EE4END[3]
+ Tile_X9Y1_LUT4AB/EE4END[4] Tile_X9Y1_LUT4AB/EE4END[5] Tile_X9Y1_LUT4AB/EE4END[6]
+ Tile_X9Y1_LUT4AB/EE4END[7] Tile_X9Y1_LUT4AB/EE4END[8] Tile_X9Y1_LUT4AB/EE4END[9]
+ Tile_X9Y1_LUT4AB/FrameData[0] Tile_X9Y1_LUT4AB/FrameData[10] Tile_X9Y1_LUT4AB/FrameData[11]
+ Tile_X9Y1_LUT4AB/FrameData[12] Tile_X9Y1_LUT4AB/FrameData[13] Tile_X9Y1_LUT4AB/FrameData[14]
+ Tile_X9Y1_LUT4AB/FrameData[15] Tile_X9Y1_LUT4AB/FrameData[16] Tile_X9Y1_LUT4AB/FrameData[17]
+ Tile_X9Y1_LUT4AB/FrameData[18] Tile_X9Y1_LUT4AB/FrameData[19] Tile_X9Y1_LUT4AB/FrameData[1]
+ Tile_X9Y1_LUT4AB/FrameData[20] Tile_X9Y1_LUT4AB/FrameData[21] Tile_X9Y1_LUT4AB/FrameData[22]
+ Tile_X9Y1_LUT4AB/FrameData[23] Tile_X9Y1_LUT4AB/FrameData[24] Tile_X9Y1_LUT4AB/FrameData[25]
+ Tile_X9Y1_LUT4AB/FrameData[26] Tile_X9Y1_LUT4AB/FrameData[27] Tile_X9Y1_LUT4AB/FrameData[28]
+ Tile_X9Y1_LUT4AB/FrameData[29] Tile_X9Y1_LUT4AB/FrameData[2] Tile_X9Y1_LUT4AB/FrameData[30]
+ Tile_X9Y1_LUT4AB/FrameData[31] Tile_X9Y1_LUT4AB/FrameData[3] Tile_X9Y1_LUT4AB/FrameData[4]
+ Tile_X9Y1_LUT4AB/FrameData[5] Tile_X9Y1_LUT4AB/FrameData[6] Tile_X9Y1_LUT4AB/FrameData[7]
+ Tile_X9Y1_LUT4AB/FrameData[8] Tile_X9Y1_LUT4AB/FrameData[9] Tile_X9Y1_LUT4AB/FrameData_O[0]
+ Tile_X9Y1_LUT4AB/FrameData_O[10] Tile_X9Y1_LUT4AB/FrameData_O[11] Tile_X9Y1_LUT4AB/FrameData_O[12]
+ Tile_X9Y1_LUT4AB/FrameData_O[13] Tile_X9Y1_LUT4AB/FrameData_O[14] Tile_X9Y1_LUT4AB/FrameData_O[15]
+ Tile_X9Y1_LUT4AB/FrameData_O[16] Tile_X9Y1_LUT4AB/FrameData_O[17] Tile_X9Y1_LUT4AB/FrameData_O[18]
+ Tile_X9Y1_LUT4AB/FrameData_O[19] Tile_X9Y1_LUT4AB/FrameData_O[1] Tile_X9Y1_LUT4AB/FrameData_O[20]
+ Tile_X9Y1_LUT4AB/FrameData_O[21] Tile_X9Y1_LUT4AB/FrameData_O[22] Tile_X9Y1_LUT4AB/FrameData_O[23]
+ Tile_X9Y1_LUT4AB/FrameData_O[24] Tile_X9Y1_LUT4AB/FrameData_O[25] Tile_X9Y1_LUT4AB/FrameData_O[26]
+ Tile_X9Y1_LUT4AB/FrameData_O[27] Tile_X9Y1_LUT4AB/FrameData_O[28] Tile_X9Y1_LUT4AB/FrameData_O[29]
+ Tile_X9Y1_LUT4AB/FrameData_O[2] Tile_X9Y1_LUT4AB/FrameData_O[30] Tile_X9Y1_LUT4AB/FrameData_O[31]
+ Tile_X9Y1_LUT4AB/FrameData_O[3] Tile_X9Y1_LUT4AB/FrameData_O[4] Tile_X9Y1_LUT4AB/FrameData_O[5]
+ Tile_X9Y1_LUT4AB/FrameData_O[6] Tile_X9Y1_LUT4AB/FrameData_O[7] Tile_X9Y1_LUT4AB/FrameData_O[8]
+ Tile_X9Y1_LUT4AB/FrameData_O[9] Tile_X9Y1_LUT4AB/FrameStrobe[0] Tile_X9Y1_LUT4AB/FrameStrobe[10]
+ Tile_X9Y1_LUT4AB/FrameStrobe[11] Tile_X9Y1_LUT4AB/FrameStrobe[12] Tile_X9Y1_LUT4AB/FrameStrobe[13]
+ Tile_X9Y1_LUT4AB/FrameStrobe[14] Tile_X9Y1_LUT4AB/FrameStrobe[15] Tile_X9Y1_LUT4AB/FrameStrobe[16]
+ Tile_X9Y1_LUT4AB/FrameStrobe[17] Tile_X9Y1_LUT4AB/FrameStrobe[18] Tile_X9Y1_LUT4AB/FrameStrobe[19]
+ Tile_X9Y1_LUT4AB/FrameStrobe[1] Tile_X9Y1_LUT4AB/FrameStrobe[2] Tile_X9Y1_LUT4AB/FrameStrobe[3]
+ Tile_X9Y1_LUT4AB/FrameStrobe[4] Tile_X9Y1_LUT4AB/FrameStrobe[5] Tile_X9Y1_LUT4AB/FrameStrobe[6]
+ Tile_X9Y1_LUT4AB/FrameStrobe[7] Tile_X9Y1_LUT4AB/FrameStrobe[8] Tile_X9Y1_LUT4AB/FrameStrobe[9]
+ Tile_X9Y1_LUT4AB/FrameStrobe_O[0] Tile_X9Y1_LUT4AB/FrameStrobe_O[10] Tile_X9Y1_LUT4AB/FrameStrobe_O[11]
+ Tile_X9Y1_LUT4AB/FrameStrobe_O[12] Tile_X9Y1_LUT4AB/FrameStrobe_O[13] Tile_X9Y1_LUT4AB/FrameStrobe_O[14]
+ Tile_X9Y1_LUT4AB/FrameStrobe_O[15] Tile_X9Y1_LUT4AB/FrameStrobe_O[16] Tile_X9Y1_LUT4AB/FrameStrobe_O[17]
+ Tile_X9Y1_LUT4AB/FrameStrobe_O[18] Tile_X9Y1_LUT4AB/FrameStrobe_O[19] Tile_X9Y1_LUT4AB/FrameStrobe_O[1]
+ Tile_X9Y1_LUT4AB/FrameStrobe_O[2] Tile_X9Y1_LUT4AB/FrameStrobe_O[3] Tile_X9Y1_LUT4AB/FrameStrobe_O[4]
+ Tile_X9Y1_LUT4AB/FrameStrobe_O[5] Tile_X9Y1_LUT4AB/FrameStrobe_O[6] Tile_X9Y1_LUT4AB/FrameStrobe_O[7]
+ Tile_X9Y1_LUT4AB/FrameStrobe_O[8] Tile_X9Y1_LUT4AB/FrameStrobe_O[9] Tile_X9Y1_LUT4AB/N1BEG[0]
+ Tile_X9Y1_LUT4AB/N1BEG[1] Tile_X9Y1_LUT4AB/N1BEG[2] Tile_X9Y1_LUT4AB/N1BEG[3] Tile_X9Y2_LUT4AB/N1BEG[0]
+ Tile_X9Y2_LUT4AB/N1BEG[1] Tile_X9Y2_LUT4AB/N1BEG[2] Tile_X9Y2_LUT4AB/N1BEG[3] Tile_X9Y1_LUT4AB/N2BEG[0]
+ Tile_X9Y1_LUT4AB/N2BEG[1] Tile_X9Y1_LUT4AB/N2BEG[2] Tile_X9Y1_LUT4AB/N2BEG[3] Tile_X9Y1_LUT4AB/N2BEG[4]
+ Tile_X9Y1_LUT4AB/N2BEG[5] Tile_X9Y1_LUT4AB/N2BEG[6] Tile_X9Y1_LUT4AB/N2BEG[7] Tile_X9Y1_LUT4AB/N2BEGb[0]
+ Tile_X9Y1_LUT4AB/N2BEGb[1] Tile_X9Y1_LUT4AB/N2BEGb[2] Tile_X9Y1_LUT4AB/N2BEGb[3]
+ Tile_X9Y1_LUT4AB/N2BEGb[4] Tile_X9Y1_LUT4AB/N2BEGb[5] Tile_X9Y1_LUT4AB/N2BEGb[6]
+ Tile_X9Y1_LUT4AB/N2BEGb[7] Tile_X9Y1_LUT4AB/N2END[0] Tile_X9Y1_LUT4AB/N2END[1] Tile_X9Y1_LUT4AB/N2END[2]
+ Tile_X9Y1_LUT4AB/N2END[3] Tile_X9Y1_LUT4AB/N2END[4] Tile_X9Y1_LUT4AB/N2END[5] Tile_X9Y1_LUT4AB/N2END[6]
+ Tile_X9Y1_LUT4AB/N2END[7] Tile_X9Y2_LUT4AB/N2BEG[0] Tile_X9Y2_LUT4AB/N2BEG[1] Tile_X9Y2_LUT4AB/N2BEG[2]
+ Tile_X9Y2_LUT4AB/N2BEG[3] Tile_X9Y2_LUT4AB/N2BEG[4] Tile_X9Y2_LUT4AB/N2BEG[5] Tile_X9Y2_LUT4AB/N2BEG[6]
+ Tile_X9Y2_LUT4AB/N2BEG[7] Tile_X9Y1_LUT4AB/N4BEG[0] Tile_X9Y1_LUT4AB/N4BEG[10] Tile_X9Y1_LUT4AB/N4BEG[11]
+ Tile_X9Y1_LUT4AB/N4BEG[12] Tile_X9Y1_LUT4AB/N4BEG[13] Tile_X9Y1_LUT4AB/N4BEG[14]
+ Tile_X9Y1_LUT4AB/N4BEG[15] Tile_X9Y1_LUT4AB/N4BEG[1] Tile_X9Y1_LUT4AB/N4BEG[2] Tile_X9Y1_LUT4AB/N4BEG[3]
+ Tile_X9Y1_LUT4AB/N4BEG[4] Tile_X9Y1_LUT4AB/N4BEG[5] Tile_X9Y1_LUT4AB/N4BEG[6] Tile_X9Y1_LUT4AB/N4BEG[7]
+ Tile_X9Y1_LUT4AB/N4BEG[8] Tile_X9Y1_LUT4AB/N4BEG[9] Tile_X9Y2_LUT4AB/N4BEG[0] Tile_X9Y2_LUT4AB/N4BEG[10]
+ Tile_X9Y2_LUT4AB/N4BEG[11] Tile_X9Y2_LUT4AB/N4BEG[12] Tile_X9Y2_LUT4AB/N4BEG[13]
+ Tile_X9Y2_LUT4AB/N4BEG[14] Tile_X9Y2_LUT4AB/N4BEG[15] Tile_X9Y2_LUT4AB/N4BEG[1]
+ Tile_X9Y2_LUT4AB/N4BEG[2] Tile_X9Y2_LUT4AB/N4BEG[3] Tile_X9Y2_LUT4AB/N4BEG[4] Tile_X9Y2_LUT4AB/N4BEG[5]
+ Tile_X9Y2_LUT4AB/N4BEG[6] Tile_X9Y2_LUT4AB/N4BEG[7] Tile_X9Y2_LUT4AB/N4BEG[8] Tile_X9Y2_LUT4AB/N4BEG[9]
+ Tile_X9Y1_LUT4AB/NN4BEG[0] Tile_X9Y1_LUT4AB/NN4BEG[10] Tile_X9Y1_LUT4AB/NN4BEG[11]
+ Tile_X9Y1_LUT4AB/NN4BEG[12] Tile_X9Y1_LUT4AB/NN4BEG[13] Tile_X9Y1_LUT4AB/NN4BEG[14]
+ Tile_X9Y1_LUT4AB/NN4BEG[15] Tile_X9Y1_LUT4AB/NN4BEG[1] Tile_X9Y1_LUT4AB/NN4BEG[2]
+ Tile_X9Y1_LUT4AB/NN4BEG[3] Tile_X9Y1_LUT4AB/NN4BEG[4] Tile_X9Y1_LUT4AB/NN4BEG[5]
+ Tile_X9Y1_LUT4AB/NN4BEG[6] Tile_X9Y1_LUT4AB/NN4BEG[7] Tile_X9Y1_LUT4AB/NN4BEG[8]
+ Tile_X9Y1_LUT4AB/NN4BEG[9] Tile_X9Y2_LUT4AB/NN4BEG[0] Tile_X9Y2_LUT4AB/NN4BEG[10]
+ Tile_X9Y2_LUT4AB/NN4BEG[11] Tile_X9Y2_LUT4AB/NN4BEG[12] Tile_X9Y2_LUT4AB/NN4BEG[13]
+ Tile_X9Y2_LUT4AB/NN4BEG[14] Tile_X9Y2_LUT4AB/NN4BEG[15] Tile_X9Y2_LUT4AB/NN4BEG[1]
+ Tile_X9Y2_LUT4AB/NN4BEG[2] Tile_X9Y2_LUT4AB/NN4BEG[3] Tile_X9Y2_LUT4AB/NN4BEG[4]
+ Tile_X9Y2_LUT4AB/NN4BEG[5] Tile_X9Y2_LUT4AB/NN4BEG[6] Tile_X9Y2_LUT4AB/NN4BEG[7]
+ Tile_X9Y2_LUT4AB/NN4BEG[8] Tile_X9Y2_LUT4AB/NN4BEG[9] Tile_X9Y2_LUT4AB/S1END[0]
+ Tile_X9Y2_LUT4AB/S1END[1] Tile_X9Y2_LUT4AB/S1END[2] Tile_X9Y2_LUT4AB/S1END[3] Tile_X9Y1_LUT4AB/S1END[0]
+ Tile_X9Y1_LUT4AB/S1END[1] Tile_X9Y1_LUT4AB/S1END[2] Tile_X9Y1_LUT4AB/S1END[3] Tile_X9Y2_LUT4AB/S2MID[0]
+ Tile_X9Y2_LUT4AB/S2MID[1] Tile_X9Y2_LUT4AB/S2MID[2] Tile_X9Y2_LUT4AB/S2MID[3] Tile_X9Y2_LUT4AB/S2MID[4]
+ Tile_X9Y2_LUT4AB/S2MID[5] Tile_X9Y2_LUT4AB/S2MID[6] Tile_X9Y2_LUT4AB/S2MID[7] Tile_X9Y2_LUT4AB/S2END[0]
+ Tile_X9Y2_LUT4AB/S2END[1] Tile_X9Y2_LUT4AB/S2END[2] Tile_X9Y2_LUT4AB/S2END[3] Tile_X9Y2_LUT4AB/S2END[4]
+ Tile_X9Y2_LUT4AB/S2END[5] Tile_X9Y2_LUT4AB/S2END[6] Tile_X9Y2_LUT4AB/S2END[7] Tile_X9Y1_LUT4AB/S2END[0]
+ Tile_X9Y1_LUT4AB/S2END[1] Tile_X9Y1_LUT4AB/S2END[2] Tile_X9Y1_LUT4AB/S2END[3] Tile_X9Y1_LUT4AB/S2END[4]
+ Tile_X9Y1_LUT4AB/S2END[5] Tile_X9Y1_LUT4AB/S2END[6] Tile_X9Y1_LUT4AB/S2END[7] Tile_X9Y1_LUT4AB/S2MID[0]
+ Tile_X9Y1_LUT4AB/S2MID[1] Tile_X9Y1_LUT4AB/S2MID[2] Tile_X9Y1_LUT4AB/S2MID[3] Tile_X9Y1_LUT4AB/S2MID[4]
+ Tile_X9Y1_LUT4AB/S2MID[5] Tile_X9Y1_LUT4AB/S2MID[6] Tile_X9Y1_LUT4AB/S2MID[7] Tile_X9Y2_LUT4AB/S4END[0]
+ Tile_X9Y2_LUT4AB/S4END[10] Tile_X9Y2_LUT4AB/S4END[11] Tile_X9Y2_LUT4AB/S4END[12]
+ Tile_X9Y2_LUT4AB/S4END[13] Tile_X9Y2_LUT4AB/S4END[14] Tile_X9Y2_LUT4AB/S4END[15]
+ Tile_X9Y2_LUT4AB/S4END[1] Tile_X9Y2_LUT4AB/S4END[2] Tile_X9Y2_LUT4AB/S4END[3] Tile_X9Y2_LUT4AB/S4END[4]
+ Tile_X9Y2_LUT4AB/S4END[5] Tile_X9Y2_LUT4AB/S4END[6] Tile_X9Y2_LUT4AB/S4END[7] Tile_X9Y2_LUT4AB/S4END[8]
+ Tile_X9Y2_LUT4AB/S4END[9] Tile_X9Y1_LUT4AB/S4END[0] Tile_X9Y1_LUT4AB/S4END[10] Tile_X9Y1_LUT4AB/S4END[11]
+ Tile_X9Y1_LUT4AB/S4END[12] Tile_X9Y1_LUT4AB/S4END[13] Tile_X9Y1_LUT4AB/S4END[14]
+ Tile_X9Y1_LUT4AB/S4END[15] Tile_X9Y1_LUT4AB/S4END[1] Tile_X9Y1_LUT4AB/S4END[2] Tile_X9Y1_LUT4AB/S4END[3]
+ Tile_X9Y1_LUT4AB/S4END[4] Tile_X9Y1_LUT4AB/S4END[5] Tile_X9Y1_LUT4AB/S4END[6] Tile_X9Y1_LUT4AB/S4END[7]
+ Tile_X9Y1_LUT4AB/S4END[8] Tile_X9Y1_LUT4AB/S4END[9] Tile_X9Y2_LUT4AB/SS4END[0] Tile_X9Y2_LUT4AB/SS4END[10]
+ Tile_X9Y2_LUT4AB/SS4END[11] Tile_X9Y2_LUT4AB/SS4END[12] Tile_X9Y2_LUT4AB/SS4END[13]
+ Tile_X9Y2_LUT4AB/SS4END[14] Tile_X9Y2_LUT4AB/SS4END[15] Tile_X9Y2_LUT4AB/SS4END[1]
+ Tile_X9Y2_LUT4AB/SS4END[2] Tile_X9Y2_LUT4AB/SS4END[3] Tile_X9Y2_LUT4AB/SS4END[4]
+ Tile_X9Y2_LUT4AB/SS4END[5] Tile_X9Y2_LUT4AB/SS4END[6] Tile_X9Y2_LUT4AB/SS4END[7]
+ Tile_X9Y2_LUT4AB/SS4END[8] Tile_X9Y2_LUT4AB/SS4END[9] Tile_X9Y1_LUT4AB/SS4END[0]
+ Tile_X9Y1_LUT4AB/SS4END[10] Tile_X9Y1_LUT4AB/SS4END[11] Tile_X9Y1_LUT4AB/SS4END[12]
+ Tile_X9Y1_LUT4AB/SS4END[13] Tile_X9Y1_LUT4AB/SS4END[14] Tile_X9Y1_LUT4AB/SS4END[15]
+ Tile_X9Y1_LUT4AB/SS4END[1] Tile_X9Y1_LUT4AB/SS4END[2] Tile_X9Y1_LUT4AB/SS4END[3]
+ Tile_X9Y1_LUT4AB/SS4END[4] Tile_X9Y1_LUT4AB/SS4END[5] Tile_X9Y1_LUT4AB/SS4END[6]
+ Tile_X9Y1_LUT4AB/SS4END[7] Tile_X9Y1_LUT4AB/SS4END[8] Tile_X9Y1_LUT4AB/SS4END[9]
+ Tile_X9Y1_LUT4AB/UserCLK Tile_X9Y1_LUT4AB/UserCLKo VGND VPWR Tile_X9Y1_LUT4AB/W1BEG[0]
+ Tile_X9Y1_LUT4AB/W1BEG[1] Tile_X9Y1_LUT4AB/W1BEG[2] Tile_X9Y1_LUT4AB/W1BEG[3] Tile_X9Y1_LUT4AB/W1END[0]
+ Tile_X9Y1_LUT4AB/W1END[1] Tile_X9Y1_LUT4AB/W1END[2] Tile_X9Y1_LUT4AB/W1END[3] Tile_X9Y1_LUT4AB/W2BEG[0]
+ Tile_X9Y1_LUT4AB/W2BEG[1] Tile_X9Y1_LUT4AB/W2BEG[2] Tile_X9Y1_LUT4AB/W2BEG[3] Tile_X9Y1_LUT4AB/W2BEG[4]
+ Tile_X9Y1_LUT4AB/W2BEG[5] Tile_X9Y1_LUT4AB/W2BEG[6] Tile_X9Y1_LUT4AB/W2BEG[7] Tile_X8Y1_LUT4AB/W2END[0]
+ Tile_X8Y1_LUT4AB/W2END[1] Tile_X8Y1_LUT4AB/W2END[2] Tile_X8Y1_LUT4AB/W2END[3] Tile_X8Y1_LUT4AB/W2END[4]
+ Tile_X8Y1_LUT4AB/W2END[5] Tile_X8Y1_LUT4AB/W2END[6] Tile_X8Y1_LUT4AB/W2END[7] Tile_X9Y1_LUT4AB/W2END[0]
+ Tile_X9Y1_LUT4AB/W2END[1] Tile_X9Y1_LUT4AB/W2END[2] Tile_X9Y1_LUT4AB/W2END[3] Tile_X9Y1_LUT4AB/W2END[4]
+ Tile_X9Y1_LUT4AB/W2END[5] Tile_X9Y1_LUT4AB/W2END[6] Tile_X9Y1_LUT4AB/W2END[7] Tile_X9Y1_LUT4AB/W2MID[0]
+ Tile_X9Y1_LUT4AB/W2MID[1] Tile_X9Y1_LUT4AB/W2MID[2] Tile_X9Y1_LUT4AB/W2MID[3] Tile_X9Y1_LUT4AB/W2MID[4]
+ Tile_X9Y1_LUT4AB/W2MID[5] Tile_X9Y1_LUT4AB/W2MID[6] Tile_X9Y1_LUT4AB/W2MID[7] Tile_X9Y1_LUT4AB/W6BEG[0]
+ Tile_X9Y1_LUT4AB/W6BEG[10] Tile_X9Y1_LUT4AB/W6BEG[11] Tile_X9Y1_LUT4AB/W6BEG[1]
+ Tile_X9Y1_LUT4AB/W6BEG[2] Tile_X9Y1_LUT4AB/W6BEG[3] Tile_X9Y1_LUT4AB/W6BEG[4] Tile_X9Y1_LUT4AB/W6BEG[5]
+ Tile_X9Y1_LUT4AB/W6BEG[6] Tile_X9Y1_LUT4AB/W6BEG[7] Tile_X9Y1_LUT4AB/W6BEG[8] Tile_X9Y1_LUT4AB/W6BEG[9]
+ Tile_X9Y1_LUT4AB/W6END[0] Tile_X9Y1_LUT4AB/W6END[10] Tile_X9Y1_LUT4AB/W6END[11]
+ Tile_X9Y1_LUT4AB/W6END[1] Tile_X9Y1_LUT4AB/W6END[2] Tile_X9Y1_LUT4AB/W6END[3] Tile_X9Y1_LUT4AB/W6END[4]
+ Tile_X9Y1_LUT4AB/W6END[5] Tile_X9Y1_LUT4AB/W6END[6] Tile_X9Y1_LUT4AB/W6END[7] Tile_X9Y1_LUT4AB/W6END[8]
+ Tile_X9Y1_LUT4AB/W6END[9] Tile_X9Y1_LUT4AB/WW4BEG[0] Tile_X9Y1_LUT4AB/WW4BEG[10]
+ Tile_X9Y1_LUT4AB/WW4BEG[11] Tile_X9Y1_LUT4AB/WW4BEG[12] Tile_X9Y1_LUT4AB/WW4BEG[13]
+ Tile_X9Y1_LUT4AB/WW4BEG[14] Tile_X9Y1_LUT4AB/WW4BEG[15] Tile_X9Y1_LUT4AB/WW4BEG[1]
+ Tile_X9Y1_LUT4AB/WW4BEG[2] Tile_X9Y1_LUT4AB/WW4BEG[3] Tile_X9Y1_LUT4AB/WW4BEG[4]
+ Tile_X9Y1_LUT4AB/WW4BEG[5] Tile_X9Y1_LUT4AB/WW4BEG[6] Tile_X9Y1_LUT4AB/WW4BEG[7]
+ Tile_X9Y1_LUT4AB/WW4BEG[8] Tile_X9Y1_LUT4AB/WW4BEG[9] Tile_X9Y1_LUT4AB/WW4END[0]
+ Tile_X9Y1_LUT4AB/WW4END[10] Tile_X9Y1_LUT4AB/WW4END[11] Tile_X9Y1_LUT4AB/WW4END[12]
+ Tile_X9Y1_LUT4AB/WW4END[13] Tile_X9Y1_LUT4AB/WW4END[14] Tile_X9Y1_LUT4AB/WW4END[15]
+ Tile_X9Y1_LUT4AB/WW4END[1] Tile_X9Y1_LUT4AB/WW4END[2] Tile_X9Y1_LUT4AB/WW4END[3]
+ Tile_X9Y1_LUT4AB/WW4END[4] Tile_X9Y1_LUT4AB/WW4END[5] Tile_X9Y1_LUT4AB/WW4END[6]
+ Tile_X9Y1_LUT4AB/WW4END[7] Tile_X9Y1_LUT4AB/WW4END[8] Tile_X9Y1_LUT4AB/WW4END[9]
+ LUT4AB
XTile_X8Y5_LUT4AB Tile_X8Y6_LUT4AB/Co Tile_X8Y5_LUT4AB/Co Tile_X9Y5_LUT4AB/E1END[0]
+ Tile_X9Y5_LUT4AB/E1END[1] Tile_X9Y5_LUT4AB/E1END[2] Tile_X9Y5_LUT4AB/E1END[3] Tile_X8Y5_LUT4AB/E1END[0]
+ Tile_X8Y5_LUT4AB/E1END[1] Tile_X8Y5_LUT4AB/E1END[2] Tile_X8Y5_LUT4AB/E1END[3] Tile_X9Y5_LUT4AB/E2MID[0]
+ Tile_X9Y5_LUT4AB/E2MID[1] Tile_X9Y5_LUT4AB/E2MID[2] Tile_X9Y5_LUT4AB/E2MID[3] Tile_X9Y5_LUT4AB/E2MID[4]
+ Tile_X9Y5_LUT4AB/E2MID[5] Tile_X9Y5_LUT4AB/E2MID[6] Tile_X9Y5_LUT4AB/E2MID[7] Tile_X9Y5_LUT4AB/E2END[0]
+ Tile_X9Y5_LUT4AB/E2END[1] Tile_X9Y5_LUT4AB/E2END[2] Tile_X9Y5_LUT4AB/E2END[3] Tile_X9Y5_LUT4AB/E2END[4]
+ Tile_X9Y5_LUT4AB/E2END[5] Tile_X9Y5_LUT4AB/E2END[6] Tile_X9Y5_LUT4AB/E2END[7] Tile_X8Y5_LUT4AB/E2END[0]
+ Tile_X8Y5_LUT4AB/E2END[1] Tile_X8Y5_LUT4AB/E2END[2] Tile_X8Y5_LUT4AB/E2END[3] Tile_X8Y5_LUT4AB/E2END[4]
+ Tile_X8Y5_LUT4AB/E2END[5] Tile_X8Y5_LUT4AB/E2END[6] Tile_X8Y5_LUT4AB/E2END[7] Tile_X8Y5_LUT4AB/E2MID[0]
+ Tile_X8Y5_LUT4AB/E2MID[1] Tile_X8Y5_LUT4AB/E2MID[2] Tile_X8Y5_LUT4AB/E2MID[3] Tile_X8Y5_LUT4AB/E2MID[4]
+ Tile_X8Y5_LUT4AB/E2MID[5] Tile_X8Y5_LUT4AB/E2MID[6] Tile_X8Y5_LUT4AB/E2MID[7] Tile_X9Y5_LUT4AB/E6END[0]
+ Tile_X9Y5_LUT4AB/E6END[10] Tile_X9Y5_LUT4AB/E6END[11] Tile_X9Y5_LUT4AB/E6END[1]
+ Tile_X9Y5_LUT4AB/E6END[2] Tile_X9Y5_LUT4AB/E6END[3] Tile_X9Y5_LUT4AB/E6END[4] Tile_X9Y5_LUT4AB/E6END[5]
+ Tile_X9Y5_LUT4AB/E6END[6] Tile_X9Y5_LUT4AB/E6END[7] Tile_X9Y5_LUT4AB/E6END[8] Tile_X9Y5_LUT4AB/E6END[9]
+ Tile_X8Y5_LUT4AB/E6END[0] Tile_X8Y5_LUT4AB/E6END[10] Tile_X8Y5_LUT4AB/E6END[11]
+ Tile_X8Y5_LUT4AB/E6END[1] Tile_X8Y5_LUT4AB/E6END[2] Tile_X8Y5_LUT4AB/E6END[3] Tile_X8Y5_LUT4AB/E6END[4]
+ Tile_X8Y5_LUT4AB/E6END[5] Tile_X8Y5_LUT4AB/E6END[6] Tile_X8Y5_LUT4AB/E6END[7] Tile_X8Y5_LUT4AB/E6END[8]
+ Tile_X8Y5_LUT4AB/E6END[9] Tile_X9Y5_LUT4AB/EE4END[0] Tile_X9Y5_LUT4AB/EE4END[10]
+ Tile_X9Y5_LUT4AB/EE4END[11] Tile_X9Y5_LUT4AB/EE4END[12] Tile_X9Y5_LUT4AB/EE4END[13]
+ Tile_X9Y5_LUT4AB/EE4END[14] Tile_X9Y5_LUT4AB/EE4END[15] Tile_X9Y5_LUT4AB/EE4END[1]
+ Tile_X9Y5_LUT4AB/EE4END[2] Tile_X9Y5_LUT4AB/EE4END[3] Tile_X9Y5_LUT4AB/EE4END[4]
+ Tile_X9Y5_LUT4AB/EE4END[5] Tile_X9Y5_LUT4AB/EE4END[6] Tile_X9Y5_LUT4AB/EE4END[7]
+ Tile_X9Y5_LUT4AB/EE4END[8] Tile_X9Y5_LUT4AB/EE4END[9] Tile_X8Y5_LUT4AB/EE4END[0]
+ Tile_X8Y5_LUT4AB/EE4END[10] Tile_X8Y5_LUT4AB/EE4END[11] Tile_X8Y5_LUT4AB/EE4END[12]
+ Tile_X8Y5_LUT4AB/EE4END[13] Tile_X8Y5_LUT4AB/EE4END[14] Tile_X8Y5_LUT4AB/EE4END[15]
+ Tile_X8Y5_LUT4AB/EE4END[1] Tile_X8Y5_LUT4AB/EE4END[2] Tile_X8Y5_LUT4AB/EE4END[3]
+ Tile_X8Y5_LUT4AB/EE4END[4] Tile_X8Y5_LUT4AB/EE4END[5] Tile_X8Y5_LUT4AB/EE4END[6]
+ Tile_X8Y5_LUT4AB/EE4END[7] Tile_X8Y5_LUT4AB/EE4END[8] Tile_X8Y5_LUT4AB/EE4END[9]
+ Tile_X8Y5_LUT4AB/FrameData[0] Tile_X8Y5_LUT4AB/FrameData[10] Tile_X8Y5_LUT4AB/FrameData[11]
+ Tile_X8Y5_LUT4AB/FrameData[12] Tile_X8Y5_LUT4AB/FrameData[13] Tile_X8Y5_LUT4AB/FrameData[14]
+ Tile_X8Y5_LUT4AB/FrameData[15] Tile_X8Y5_LUT4AB/FrameData[16] Tile_X8Y5_LUT4AB/FrameData[17]
+ Tile_X8Y5_LUT4AB/FrameData[18] Tile_X8Y5_LUT4AB/FrameData[19] Tile_X8Y5_LUT4AB/FrameData[1]
+ Tile_X8Y5_LUT4AB/FrameData[20] Tile_X8Y5_LUT4AB/FrameData[21] Tile_X8Y5_LUT4AB/FrameData[22]
+ Tile_X8Y5_LUT4AB/FrameData[23] Tile_X8Y5_LUT4AB/FrameData[24] Tile_X8Y5_LUT4AB/FrameData[25]
+ Tile_X8Y5_LUT4AB/FrameData[26] Tile_X8Y5_LUT4AB/FrameData[27] Tile_X8Y5_LUT4AB/FrameData[28]
+ Tile_X8Y5_LUT4AB/FrameData[29] Tile_X8Y5_LUT4AB/FrameData[2] Tile_X8Y5_LUT4AB/FrameData[30]
+ Tile_X8Y5_LUT4AB/FrameData[31] Tile_X8Y5_LUT4AB/FrameData[3] Tile_X8Y5_LUT4AB/FrameData[4]
+ Tile_X8Y5_LUT4AB/FrameData[5] Tile_X8Y5_LUT4AB/FrameData[6] Tile_X8Y5_LUT4AB/FrameData[7]
+ Tile_X8Y5_LUT4AB/FrameData[8] Tile_X8Y5_LUT4AB/FrameData[9] Tile_X9Y5_LUT4AB/FrameData[0]
+ Tile_X9Y5_LUT4AB/FrameData[10] Tile_X9Y5_LUT4AB/FrameData[11] Tile_X9Y5_LUT4AB/FrameData[12]
+ Tile_X9Y5_LUT4AB/FrameData[13] Tile_X9Y5_LUT4AB/FrameData[14] Tile_X9Y5_LUT4AB/FrameData[15]
+ Tile_X9Y5_LUT4AB/FrameData[16] Tile_X9Y5_LUT4AB/FrameData[17] Tile_X9Y5_LUT4AB/FrameData[18]
+ Tile_X9Y5_LUT4AB/FrameData[19] Tile_X9Y5_LUT4AB/FrameData[1] Tile_X9Y5_LUT4AB/FrameData[20]
+ Tile_X9Y5_LUT4AB/FrameData[21] Tile_X9Y5_LUT4AB/FrameData[22] Tile_X9Y5_LUT4AB/FrameData[23]
+ Tile_X9Y5_LUT4AB/FrameData[24] Tile_X9Y5_LUT4AB/FrameData[25] Tile_X9Y5_LUT4AB/FrameData[26]
+ Tile_X9Y5_LUT4AB/FrameData[27] Tile_X9Y5_LUT4AB/FrameData[28] Tile_X9Y5_LUT4AB/FrameData[29]
+ Tile_X9Y5_LUT4AB/FrameData[2] Tile_X9Y5_LUT4AB/FrameData[30] Tile_X9Y5_LUT4AB/FrameData[31]
+ Tile_X9Y5_LUT4AB/FrameData[3] Tile_X9Y5_LUT4AB/FrameData[4] Tile_X9Y5_LUT4AB/FrameData[5]
+ Tile_X9Y5_LUT4AB/FrameData[6] Tile_X9Y5_LUT4AB/FrameData[7] Tile_X9Y5_LUT4AB/FrameData[8]
+ Tile_X9Y5_LUT4AB/FrameData[9] Tile_X8Y5_LUT4AB/FrameStrobe[0] Tile_X8Y5_LUT4AB/FrameStrobe[10]
+ Tile_X8Y5_LUT4AB/FrameStrobe[11] Tile_X8Y5_LUT4AB/FrameStrobe[12] Tile_X8Y5_LUT4AB/FrameStrobe[13]
+ Tile_X8Y5_LUT4AB/FrameStrobe[14] Tile_X8Y5_LUT4AB/FrameStrobe[15] Tile_X8Y5_LUT4AB/FrameStrobe[16]
+ Tile_X8Y5_LUT4AB/FrameStrobe[17] Tile_X8Y5_LUT4AB/FrameStrobe[18] Tile_X8Y5_LUT4AB/FrameStrobe[19]
+ Tile_X8Y5_LUT4AB/FrameStrobe[1] Tile_X8Y5_LUT4AB/FrameStrobe[2] Tile_X8Y5_LUT4AB/FrameStrobe[3]
+ Tile_X8Y5_LUT4AB/FrameStrobe[4] Tile_X8Y5_LUT4AB/FrameStrobe[5] Tile_X8Y5_LUT4AB/FrameStrobe[6]
+ Tile_X8Y5_LUT4AB/FrameStrobe[7] Tile_X8Y5_LUT4AB/FrameStrobe[8] Tile_X8Y5_LUT4AB/FrameStrobe[9]
+ Tile_X8Y4_LUT4AB/FrameStrobe[0] Tile_X8Y4_LUT4AB/FrameStrobe[10] Tile_X8Y4_LUT4AB/FrameStrobe[11]
+ Tile_X8Y4_LUT4AB/FrameStrobe[12] Tile_X8Y4_LUT4AB/FrameStrobe[13] Tile_X8Y4_LUT4AB/FrameStrobe[14]
+ Tile_X8Y4_LUT4AB/FrameStrobe[15] Tile_X8Y4_LUT4AB/FrameStrobe[16] Tile_X8Y4_LUT4AB/FrameStrobe[17]
+ Tile_X8Y4_LUT4AB/FrameStrobe[18] Tile_X8Y4_LUT4AB/FrameStrobe[19] Tile_X8Y4_LUT4AB/FrameStrobe[1]
+ Tile_X8Y4_LUT4AB/FrameStrobe[2] Tile_X8Y4_LUT4AB/FrameStrobe[3] Tile_X8Y4_LUT4AB/FrameStrobe[4]
+ Tile_X8Y4_LUT4AB/FrameStrobe[5] Tile_X8Y4_LUT4AB/FrameStrobe[6] Tile_X8Y4_LUT4AB/FrameStrobe[7]
+ Tile_X8Y4_LUT4AB/FrameStrobe[8] Tile_X8Y4_LUT4AB/FrameStrobe[9] Tile_X8Y5_LUT4AB/N1BEG[0]
+ Tile_X8Y5_LUT4AB/N1BEG[1] Tile_X8Y5_LUT4AB/N1BEG[2] Tile_X8Y5_LUT4AB/N1BEG[3] Tile_X8Y6_LUT4AB/N1BEG[0]
+ Tile_X8Y6_LUT4AB/N1BEG[1] Tile_X8Y6_LUT4AB/N1BEG[2] Tile_X8Y6_LUT4AB/N1BEG[3] Tile_X8Y5_LUT4AB/N2BEG[0]
+ Tile_X8Y5_LUT4AB/N2BEG[1] Tile_X8Y5_LUT4AB/N2BEG[2] Tile_X8Y5_LUT4AB/N2BEG[3] Tile_X8Y5_LUT4AB/N2BEG[4]
+ Tile_X8Y5_LUT4AB/N2BEG[5] Tile_X8Y5_LUT4AB/N2BEG[6] Tile_X8Y5_LUT4AB/N2BEG[7] Tile_X8Y4_LUT4AB/N2END[0]
+ Tile_X8Y4_LUT4AB/N2END[1] Tile_X8Y4_LUT4AB/N2END[2] Tile_X8Y4_LUT4AB/N2END[3] Tile_X8Y4_LUT4AB/N2END[4]
+ Tile_X8Y4_LUT4AB/N2END[5] Tile_X8Y4_LUT4AB/N2END[6] Tile_X8Y4_LUT4AB/N2END[7] Tile_X8Y5_LUT4AB/N2END[0]
+ Tile_X8Y5_LUT4AB/N2END[1] Tile_X8Y5_LUT4AB/N2END[2] Tile_X8Y5_LUT4AB/N2END[3] Tile_X8Y5_LUT4AB/N2END[4]
+ Tile_X8Y5_LUT4AB/N2END[5] Tile_X8Y5_LUT4AB/N2END[6] Tile_X8Y5_LUT4AB/N2END[7] Tile_X8Y6_LUT4AB/N2BEG[0]
+ Tile_X8Y6_LUT4AB/N2BEG[1] Tile_X8Y6_LUT4AB/N2BEG[2] Tile_X8Y6_LUT4AB/N2BEG[3] Tile_X8Y6_LUT4AB/N2BEG[4]
+ Tile_X8Y6_LUT4AB/N2BEG[5] Tile_X8Y6_LUT4AB/N2BEG[6] Tile_X8Y6_LUT4AB/N2BEG[7] Tile_X8Y5_LUT4AB/N4BEG[0]
+ Tile_X8Y5_LUT4AB/N4BEG[10] Tile_X8Y5_LUT4AB/N4BEG[11] Tile_X8Y5_LUT4AB/N4BEG[12]
+ Tile_X8Y5_LUT4AB/N4BEG[13] Tile_X8Y5_LUT4AB/N4BEG[14] Tile_X8Y5_LUT4AB/N4BEG[15]
+ Tile_X8Y5_LUT4AB/N4BEG[1] Tile_X8Y5_LUT4AB/N4BEG[2] Tile_X8Y5_LUT4AB/N4BEG[3] Tile_X8Y5_LUT4AB/N4BEG[4]
+ Tile_X8Y5_LUT4AB/N4BEG[5] Tile_X8Y5_LUT4AB/N4BEG[6] Tile_X8Y5_LUT4AB/N4BEG[7] Tile_X8Y5_LUT4AB/N4BEG[8]
+ Tile_X8Y5_LUT4AB/N4BEG[9] Tile_X8Y6_LUT4AB/N4BEG[0] Tile_X8Y6_LUT4AB/N4BEG[10] Tile_X8Y6_LUT4AB/N4BEG[11]
+ Tile_X8Y6_LUT4AB/N4BEG[12] Tile_X8Y6_LUT4AB/N4BEG[13] Tile_X8Y6_LUT4AB/N4BEG[14]
+ Tile_X8Y6_LUT4AB/N4BEG[15] Tile_X8Y6_LUT4AB/N4BEG[1] Tile_X8Y6_LUT4AB/N4BEG[2] Tile_X8Y6_LUT4AB/N4BEG[3]
+ Tile_X8Y6_LUT4AB/N4BEG[4] Tile_X8Y6_LUT4AB/N4BEG[5] Tile_X8Y6_LUT4AB/N4BEG[6] Tile_X8Y6_LUT4AB/N4BEG[7]
+ Tile_X8Y6_LUT4AB/N4BEG[8] Tile_X8Y6_LUT4AB/N4BEG[9] Tile_X8Y5_LUT4AB/NN4BEG[0] Tile_X8Y5_LUT4AB/NN4BEG[10]
+ Tile_X8Y5_LUT4AB/NN4BEG[11] Tile_X8Y5_LUT4AB/NN4BEG[12] Tile_X8Y5_LUT4AB/NN4BEG[13]
+ Tile_X8Y5_LUT4AB/NN4BEG[14] Tile_X8Y5_LUT4AB/NN4BEG[15] Tile_X8Y5_LUT4AB/NN4BEG[1]
+ Tile_X8Y5_LUT4AB/NN4BEG[2] Tile_X8Y5_LUT4AB/NN4BEG[3] Tile_X8Y5_LUT4AB/NN4BEG[4]
+ Tile_X8Y5_LUT4AB/NN4BEG[5] Tile_X8Y5_LUT4AB/NN4BEG[6] Tile_X8Y5_LUT4AB/NN4BEG[7]
+ Tile_X8Y5_LUT4AB/NN4BEG[8] Tile_X8Y5_LUT4AB/NN4BEG[9] Tile_X8Y6_LUT4AB/NN4BEG[0]
+ Tile_X8Y6_LUT4AB/NN4BEG[10] Tile_X8Y6_LUT4AB/NN4BEG[11] Tile_X8Y6_LUT4AB/NN4BEG[12]
+ Tile_X8Y6_LUT4AB/NN4BEG[13] Tile_X8Y6_LUT4AB/NN4BEG[14] Tile_X8Y6_LUT4AB/NN4BEG[15]
+ Tile_X8Y6_LUT4AB/NN4BEG[1] Tile_X8Y6_LUT4AB/NN4BEG[2] Tile_X8Y6_LUT4AB/NN4BEG[3]
+ Tile_X8Y6_LUT4AB/NN4BEG[4] Tile_X8Y6_LUT4AB/NN4BEG[5] Tile_X8Y6_LUT4AB/NN4BEG[6]
+ Tile_X8Y6_LUT4AB/NN4BEG[7] Tile_X8Y6_LUT4AB/NN4BEG[8] Tile_X8Y6_LUT4AB/NN4BEG[9]
+ Tile_X8Y6_LUT4AB/S1END[0] Tile_X8Y6_LUT4AB/S1END[1] Tile_X8Y6_LUT4AB/S1END[2] Tile_X8Y6_LUT4AB/S1END[3]
+ Tile_X8Y5_LUT4AB/S1END[0] Tile_X8Y5_LUT4AB/S1END[1] Tile_X8Y5_LUT4AB/S1END[2] Tile_X8Y5_LUT4AB/S1END[3]
+ Tile_X8Y6_LUT4AB/S2MID[0] Tile_X8Y6_LUT4AB/S2MID[1] Tile_X8Y6_LUT4AB/S2MID[2] Tile_X8Y6_LUT4AB/S2MID[3]
+ Tile_X8Y6_LUT4AB/S2MID[4] Tile_X8Y6_LUT4AB/S2MID[5] Tile_X8Y6_LUT4AB/S2MID[6] Tile_X8Y6_LUT4AB/S2MID[7]
+ Tile_X8Y6_LUT4AB/S2END[0] Tile_X8Y6_LUT4AB/S2END[1] Tile_X8Y6_LUT4AB/S2END[2] Tile_X8Y6_LUT4AB/S2END[3]
+ Tile_X8Y6_LUT4AB/S2END[4] Tile_X8Y6_LUT4AB/S2END[5] Tile_X8Y6_LUT4AB/S2END[6] Tile_X8Y6_LUT4AB/S2END[7]
+ Tile_X8Y5_LUT4AB/S2END[0] Tile_X8Y5_LUT4AB/S2END[1] Tile_X8Y5_LUT4AB/S2END[2] Tile_X8Y5_LUT4AB/S2END[3]
+ Tile_X8Y5_LUT4AB/S2END[4] Tile_X8Y5_LUT4AB/S2END[5] Tile_X8Y5_LUT4AB/S2END[6] Tile_X8Y5_LUT4AB/S2END[7]
+ Tile_X8Y5_LUT4AB/S2MID[0] Tile_X8Y5_LUT4AB/S2MID[1] Tile_X8Y5_LUT4AB/S2MID[2] Tile_X8Y5_LUT4AB/S2MID[3]
+ Tile_X8Y5_LUT4AB/S2MID[4] Tile_X8Y5_LUT4AB/S2MID[5] Tile_X8Y5_LUT4AB/S2MID[6] Tile_X8Y5_LUT4AB/S2MID[7]
+ Tile_X8Y6_LUT4AB/S4END[0] Tile_X8Y6_LUT4AB/S4END[10] Tile_X8Y6_LUT4AB/S4END[11]
+ Tile_X8Y6_LUT4AB/S4END[12] Tile_X8Y6_LUT4AB/S4END[13] Tile_X8Y6_LUT4AB/S4END[14]
+ Tile_X8Y6_LUT4AB/S4END[15] Tile_X8Y6_LUT4AB/S4END[1] Tile_X8Y6_LUT4AB/S4END[2] Tile_X8Y6_LUT4AB/S4END[3]
+ Tile_X8Y6_LUT4AB/S4END[4] Tile_X8Y6_LUT4AB/S4END[5] Tile_X8Y6_LUT4AB/S4END[6] Tile_X8Y6_LUT4AB/S4END[7]
+ Tile_X8Y6_LUT4AB/S4END[8] Tile_X8Y6_LUT4AB/S4END[9] Tile_X8Y5_LUT4AB/S4END[0] Tile_X8Y5_LUT4AB/S4END[10]
+ Tile_X8Y5_LUT4AB/S4END[11] Tile_X8Y5_LUT4AB/S4END[12] Tile_X8Y5_LUT4AB/S4END[13]
+ Tile_X8Y5_LUT4AB/S4END[14] Tile_X8Y5_LUT4AB/S4END[15] Tile_X8Y5_LUT4AB/S4END[1]
+ Tile_X8Y5_LUT4AB/S4END[2] Tile_X8Y5_LUT4AB/S4END[3] Tile_X8Y5_LUT4AB/S4END[4] Tile_X8Y5_LUT4AB/S4END[5]
+ Tile_X8Y5_LUT4AB/S4END[6] Tile_X8Y5_LUT4AB/S4END[7] Tile_X8Y5_LUT4AB/S4END[8] Tile_X8Y5_LUT4AB/S4END[9]
+ Tile_X8Y6_LUT4AB/SS4END[0] Tile_X8Y6_LUT4AB/SS4END[10] Tile_X8Y6_LUT4AB/SS4END[11]
+ Tile_X8Y6_LUT4AB/SS4END[12] Tile_X8Y6_LUT4AB/SS4END[13] Tile_X8Y6_LUT4AB/SS4END[14]
+ Tile_X8Y6_LUT4AB/SS4END[15] Tile_X8Y6_LUT4AB/SS4END[1] Tile_X8Y6_LUT4AB/SS4END[2]
+ Tile_X8Y6_LUT4AB/SS4END[3] Tile_X8Y6_LUT4AB/SS4END[4] Tile_X8Y6_LUT4AB/SS4END[5]
+ Tile_X8Y6_LUT4AB/SS4END[6] Tile_X8Y6_LUT4AB/SS4END[7] Tile_X8Y6_LUT4AB/SS4END[8]
+ Tile_X8Y6_LUT4AB/SS4END[9] Tile_X8Y5_LUT4AB/SS4END[0] Tile_X8Y5_LUT4AB/SS4END[10]
+ Tile_X8Y5_LUT4AB/SS4END[11] Tile_X8Y5_LUT4AB/SS4END[12] Tile_X8Y5_LUT4AB/SS4END[13]
+ Tile_X8Y5_LUT4AB/SS4END[14] Tile_X8Y5_LUT4AB/SS4END[15] Tile_X8Y5_LUT4AB/SS4END[1]
+ Tile_X8Y5_LUT4AB/SS4END[2] Tile_X8Y5_LUT4AB/SS4END[3] Tile_X8Y5_LUT4AB/SS4END[4]
+ Tile_X8Y5_LUT4AB/SS4END[5] Tile_X8Y5_LUT4AB/SS4END[6] Tile_X8Y5_LUT4AB/SS4END[7]
+ Tile_X8Y5_LUT4AB/SS4END[8] Tile_X8Y5_LUT4AB/SS4END[9] Tile_X8Y5_LUT4AB/UserCLK Tile_X8Y4_LUT4AB/UserCLK
+ VGND VPWR Tile_X8Y5_LUT4AB/W1BEG[0] Tile_X8Y5_LUT4AB/W1BEG[1] Tile_X8Y5_LUT4AB/W1BEG[2]
+ Tile_X8Y5_LUT4AB/W1BEG[3] Tile_X9Y5_LUT4AB/W1BEG[0] Tile_X9Y5_LUT4AB/W1BEG[1] Tile_X9Y5_LUT4AB/W1BEG[2]
+ Tile_X9Y5_LUT4AB/W1BEG[3] Tile_X8Y5_LUT4AB/W2BEG[0] Tile_X8Y5_LUT4AB/W2BEG[1] Tile_X8Y5_LUT4AB/W2BEG[2]
+ Tile_X8Y5_LUT4AB/W2BEG[3] Tile_X8Y5_LUT4AB/W2BEG[4] Tile_X8Y5_LUT4AB/W2BEG[5] Tile_X8Y5_LUT4AB/W2BEG[6]
+ Tile_X8Y5_LUT4AB/W2BEG[7] Tile_X8Y5_LUT4AB/W2BEGb[0] Tile_X8Y5_LUT4AB/W2BEGb[1]
+ Tile_X8Y5_LUT4AB/W2BEGb[2] Tile_X8Y5_LUT4AB/W2BEGb[3] Tile_X8Y5_LUT4AB/W2BEGb[4]
+ Tile_X8Y5_LUT4AB/W2BEGb[5] Tile_X8Y5_LUT4AB/W2BEGb[6] Tile_X8Y5_LUT4AB/W2BEGb[7]
+ Tile_X8Y5_LUT4AB/W2END[0] Tile_X8Y5_LUT4AB/W2END[1] Tile_X8Y5_LUT4AB/W2END[2] Tile_X8Y5_LUT4AB/W2END[3]
+ Tile_X8Y5_LUT4AB/W2END[4] Tile_X8Y5_LUT4AB/W2END[5] Tile_X8Y5_LUT4AB/W2END[6] Tile_X8Y5_LUT4AB/W2END[7]
+ Tile_X9Y5_LUT4AB/W2BEG[0] Tile_X9Y5_LUT4AB/W2BEG[1] Tile_X9Y5_LUT4AB/W2BEG[2] Tile_X9Y5_LUT4AB/W2BEG[3]
+ Tile_X9Y5_LUT4AB/W2BEG[4] Tile_X9Y5_LUT4AB/W2BEG[5] Tile_X9Y5_LUT4AB/W2BEG[6] Tile_X9Y5_LUT4AB/W2BEG[7]
+ Tile_X8Y5_LUT4AB/W6BEG[0] Tile_X8Y5_LUT4AB/W6BEG[10] Tile_X8Y5_LUT4AB/W6BEG[11]
+ Tile_X8Y5_LUT4AB/W6BEG[1] Tile_X8Y5_LUT4AB/W6BEG[2] Tile_X8Y5_LUT4AB/W6BEG[3] Tile_X8Y5_LUT4AB/W6BEG[4]
+ Tile_X8Y5_LUT4AB/W6BEG[5] Tile_X8Y5_LUT4AB/W6BEG[6] Tile_X8Y5_LUT4AB/W6BEG[7] Tile_X8Y5_LUT4AB/W6BEG[8]
+ Tile_X8Y5_LUT4AB/W6BEG[9] Tile_X9Y5_LUT4AB/W6BEG[0] Tile_X9Y5_LUT4AB/W6BEG[10] Tile_X9Y5_LUT4AB/W6BEG[11]
+ Tile_X9Y5_LUT4AB/W6BEG[1] Tile_X9Y5_LUT4AB/W6BEG[2] Tile_X9Y5_LUT4AB/W6BEG[3] Tile_X9Y5_LUT4AB/W6BEG[4]
+ Tile_X9Y5_LUT4AB/W6BEG[5] Tile_X9Y5_LUT4AB/W6BEG[6] Tile_X9Y5_LUT4AB/W6BEG[7] Tile_X9Y5_LUT4AB/W6BEG[8]
+ Tile_X9Y5_LUT4AB/W6BEG[9] Tile_X8Y5_LUT4AB/WW4BEG[0] Tile_X8Y5_LUT4AB/WW4BEG[10]
+ Tile_X8Y5_LUT4AB/WW4BEG[11] Tile_X8Y5_LUT4AB/WW4BEG[12] Tile_X8Y5_LUT4AB/WW4BEG[13]
+ Tile_X8Y5_LUT4AB/WW4BEG[14] Tile_X8Y5_LUT4AB/WW4BEG[15] Tile_X8Y5_LUT4AB/WW4BEG[1]
+ Tile_X8Y5_LUT4AB/WW4BEG[2] Tile_X8Y5_LUT4AB/WW4BEG[3] Tile_X8Y5_LUT4AB/WW4BEG[4]
+ Tile_X8Y5_LUT4AB/WW4BEG[5] Tile_X8Y5_LUT4AB/WW4BEG[6] Tile_X8Y5_LUT4AB/WW4BEG[7]
+ Tile_X8Y5_LUT4AB/WW4BEG[8] Tile_X8Y5_LUT4AB/WW4BEG[9] Tile_X9Y5_LUT4AB/WW4BEG[0]
+ Tile_X9Y5_LUT4AB/WW4BEG[10] Tile_X9Y5_LUT4AB/WW4BEG[11] Tile_X9Y5_LUT4AB/WW4BEG[12]
+ Tile_X9Y5_LUT4AB/WW4BEG[13] Tile_X9Y5_LUT4AB/WW4BEG[14] Tile_X9Y5_LUT4AB/WW4BEG[15]
+ Tile_X9Y5_LUT4AB/WW4BEG[1] Tile_X9Y5_LUT4AB/WW4BEG[2] Tile_X9Y5_LUT4AB/WW4BEG[3]
+ Tile_X9Y5_LUT4AB/WW4BEG[4] Tile_X9Y5_LUT4AB/WW4BEG[5] Tile_X9Y5_LUT4AB/WW4BEG[6]
+ Tile_X9Y5_LUT4AB/WW4BEG[7] Tile_X9Y5_LUT4AB/WW4BEG[8] Tile_X9Y5_LUT4AB/WW4BEG[9]
+ LUT4AB
XTile_X9Y12_LUT4AB Tile_X9Y13_LUT4AB/Co Tile_X9Y12_LUT4AB/Co Tile_X9Y12_LUT4AB/E1BEG[0]
+ Tile_X9Y12_LUT4AB/E1BEG[1] Tile_X9Y12_LUT4AB/E1BEG[2] Tile_X9Y12_LUT4AB/E1BEG[3]
+ Tile_X9Y12_LUT4AB/E1END[0] Tile_X9Y12_LUT4AB/E1END[1] Tile_X9Y12_LUT4AB/E1END[2]
+ Tile_X9Y12_LUT4AB/E1END[3] Tile_X9Y12_LUT4AB/E2BEG[0] Tile_X9Y12_LUT4AB/E2BEG[1]
+ Tile_X9Y12_LUT4AB/E2BEG[2] Tile_X9Y12_LUT4AB/E2BEG[3] Tile_X9Y12_LUT4AB/E2BEG[4]
+ Tile_X9Y12_LUT4AB/E2BEG[5] Tile_X9Y12_LUT4AB/E2BEG[6] Tile_X9Y12_LUT4AB/E2BEG[7]
+ Tile_X9Y12_LUT4AB/E2BEGb[0] Tile_X9Y12_LUT4AB/E2BEGb[1] Tile_X9Y12_LUT4AB/E2BEGb[2]
+ Tile_X9Y12_LUT4AB/E2BEGb[3] Tile_X9Y12_LUT4AB/E2BEGb[4] Tile_X9Y12_LUT4AB/E2BEGb[5]
+ Tile_X9Y12_LUT4AB/E2BEGb[6] Tile_X9Y12_LUT4AB/E2BEGb[7] Tile_X9Y12_LUT4AB/E2END[0]
+ Tile_X9Y12_LUT4AB/E2END[1] Tile_X9Y12_LUT4AB/E2END[2] Tile_X9Y12_LUT4AB/E2END[3]
+ Tile_X9Y12_LUT4AB/E2END[4] Tile_X9Y12_LUT4AB/E2END[5] Tile_X9Y12_LUT4AB/E2END[6]
+ Tile_X9Y12_LUT4AB/E2END[7] Tile_X9Y12_LUT4AB/E2MID[0] Tile_X9Y12_LUT4AB/E2MID[1]
+ Tile_X9Y12_LUT4AB/E2MID[2] Tile_X9Y12_LUT4AB/E2MID[3] Tile_X9Y12_LUT4AB/E2MID[4]
+ Tile_X9Y12_LUT4AB/E2MID[5] Tile_X9Y12_LUT4AB/E2MID[6] Tile_X9Y12_LUT4AB/E2MID[7]
+ Tile_X9Y12_LUT4AB/E6BEG[0] Tile_X9Y12_LUT4AB/E6BEG[10] Tile_X9Y12_LUT4AB/E6BEG[11]
+ Tile_X9Y12_LUT4AB/E6BEG[1] Tile_X9Y12_LUT4AB/E6BEG[2] Tile_X9Y12_LUT4AB/E6BEG[3]
+ Tile_X9Y12_LUT4AB/E6BEG[4] Tile_X9Y12_LUT4AB/E6BEG[5] Tile_X9Y12_LUT4AB/E6BEG[6]
+ Tile_X9Y12_LUT4AB/E6BEG[7] Tile_X9Y12_LUT4AB/E6BEG[8] Tile_X9Y12_LUT4AB/E6BEG[9]
+ Tile_X9Y12_LUT4AB/E6END[0] Tile_X9Y12_LUT4AB/E6END[10] Tile_X9Y12_LUT4AB/E6END[11]
+ Tile_X9Y12_LUT4AB/E6END[1] Tile_X9Y12_LUT4AB/E6END[2] Tile_X9Y12_LUT4AB/E6END[3]
+ Tile_X9Y12_LUT4AB/E6END[4] Tile_X9Y12_LUT4AB/E6END[5] Tile_X9Y12_LUT4AB/E6END[6]
+ Tile_X9Y12_LUT4AB/E6END[7] Tile_X9Y12_LUT4AB/E6END[8] Tile_X9Y12_LUT4AB/E6END[9]
+ Tile_X9Y12_LUT4AB/EE4BEG[0] Tile_X9Y12_LUT4AB/EE4BEG[10] Tile_X9Y12_LUT4AB/EE4BEG[11]
+ Tile_X9Y12_LUT4AB/EE4BEG[12] Tile_X9Y12_LUT4AB/EE4BEG[13] Tile_X9Y12_LUT4AB/EE4BEG[14]
+ Tile_X9Y12_LUT4AB/EE4BEG[15] Tile_X9Y12_LUT4AB/EE4BEG[1] Tile_X9Y12_LUT4AB/EE4BEG[2]
+ Tile_X9Y12_LUT4AB/EE4BEG[3] Tile_X9Y12_LUT4AB/EE4BEG[4] Tile_X9Y12_LUT4AB/EE4BEG[5]
+ Tile_X9Y12_LUT4AB/EE4BEG[6] Tile_X9Y12_LUT4AB/EE4BEG[7] Tile_X9Y12_LUT4AB/EE4BEG[8]
+ Tile_X9Y12_LUT4AB/EE4BEG[9] Tile_X9Y12_LUT4AB/EE4END[0] Tile_X9Y12_LUT4AB/EE4END[10]
+ Tile_X9Y12_LUT4AB/EE4END[11] Tile_X9Y12_LUT4AB/EE4END[12] Tile_X9Y12_LUT4AB/EE4END[13]
+ Tile_X9Y12_LUT4AB/EE4END[14] Tile_X9Y12_LUT4AB/EE4END[15] Tile_X9Y12_LUT4AB/EE4END[1]
+ Tile_X9Y12_LUT4AB/EE4END[2] Tile_X9Y12_LUT4AB/EE4END[3] Tile_X9Y12_LUT4AB/EE4END[4]
+ Tile_X9Y12_LUT4AB/EE4END[5] Tile_X9Y12_LUT4AB/EE4END[6] Tile_X9Y12_LUT4AB/EE4END[7]
+ Tile_X9Y12_LUT4AB/EE4END[8] Tile_X9Y12_LUT4AB/EE4END[9] Tile_X9Y12_LUT4AB/FrameData[0]
+ Tile_X9Y12_LUT4AB/FrameData[10] Tile_X9Y12_LUT4AB/FrameData[11] Tile_X9Y12_LUT4AB/FrameData[12]
+ Tile_X9Y12_LUT4AB/FrameData[13] Tile_X9Y12_LUT4AB/FrameData[14] Tile_X9Y12_LUT4AB/FrameData[15]
+ Tile_X9Y12_LUT4AB/FrameData[16] Tile_X9Y12_LUT4AB/FrameData[17] Tile_X9Y12_LUT4AB/FrameData[18]
+ Tile_X9Y12_LUT4AB/FrameData[19] Tile_X9Y12_LUT4AB/FrameData[1] Tile_X9Y12_LUT4AB/FrameData[20]
+ Tile_X9Y12_LUT4AB/FrameData[21] Tile_X9Y12_LUT4AB/FrameData[22] Tile_X9Y12_LUT4AB/FrameData[23]
+ Tile_X9Y12_LUT4AB/FrameData[24] Tile_X9Y12_LUT4AB/FrameData[25] Tile_X9Y12_LUT4AB/FrameData[26]
+ Tile_X9Y12_LUT4AB/FrameData[27] Tile_X9Y12_LUT4AB/FrameData[28] Tile_X9Y12_LUT4AB/FrameData[29]
+ Tile_X9Y12_LUT4AB/FrameData[2] Tile_X9Y12_LUT4AB/FrameData[30] Tile_X9Y12_LUT4AB/FrameData[31]
+ Tile_X9Y12_LUT4AB/FrameData[3] Tile_X9Y12_LUT4AB/FrameData[4] Tile_X9Y12_LUT4AB/FrameData[5]
+ Tile_X9Y12_LUT4AB/FrameData[6] Tile_X9Y12_LUT4AB/FrameData[7] Tile_X9Y12_LUT4AB/FrameData[8]
+ Tile_X9Y12_LUT4AB/FrameData[9] Tile_X9Y12_LUT4AB/FrameData_O[0] Tile_X9Y12_LUT4AB/FrameData_O[10]
+ Tile_X9Y12_LUT4AB/FrameData_O[11] Tile_X9Y12_LUT4AB/FrameData_O[12] Tile_X9Y12_LUT4AB/FrameData_O[13]
+ Tile_X9Y12_LUT4AB/FrameData_O[14] Tile_X9Y12_LUT4AB/FrameData_O[15] Tile_X9Y12_LUT4AB/FrameData_O[16]
+ Tile_X9Y12_LUT4AB/FrameData_O[17] Tile_X9Y12_LUT4AB/FrameData_O[18] Tile_X9Y12_LUT4AB/FrameData_O[19]
+ Tile_X9Y12_LUT4AB/FrameData_O[1] Tile_X9Y12_LUT4AB/FrameData_O[20] Tile_X9Y12_LUT4AB/FrameData_O[21]
+ Tile_X9Y12_LUT4AB/FrameData_O[22] Tile_X9Y12_LUT4AB/FrameData_O[23] Tile_X9Y12_LUT4AB/FrameData_O[24]
+ Tile_X9Y12_LUT4AB/FrameData_O[25] Tile_X9Y12_LUT4AB/FrameData_O[26] Tile_X9Y12_LUT4AB/FrameData_O[27]
+ Tile_X9Y12_LUT4AB/FrameData_O[28] Tile_X9Y12_LUT4AB/FrameData_O[29] Tile_X9Y12_LUT4AB/FrameData_O[2]
+ Tile_X9Y12_LUT4AB/FrameData_O[30] Tile_X9Y12_LUT4AB/FrameData_O[31] Tile_X9Y12_LUT4AB/FrameData_O[3]
+ Tile_X9Y12_LUT4AB/FrameData_O[4] Tile_X9Y12_LUT4AB/FrameData_O[5] Tile_X9Y12_LUT4AB/FrameData_O[6]
+ Tile_X9Y12_LUT4AB/FrameData_O[7] Tile_X9Y12_LUT4AB/FrameData_O[8] Tile_X9Y12_LUT4AB/FrameData_O[9]
+ Tile_X9Y12_LUT4AB/FrameStrobe[0] Tile_X9Y12_LUT4AB/FrameStrobe[10] Tile_X9Y12_LUT4AB/FrameStrobe[11]
+ Tile_X9Y12_LUT4AB/FrameStrobe[12] Tile_X9Y12_LUT4AB/FrameStrobe[13] Tile_X9Y12_LUT4AB/FrameStrobe[14]
+ Tile_X9Y12_LUT4AB/FrameStrobe[15] Tile_X9Y12_LUT4AB/FrameStrobe[16] Tile_X9Y12_LUT4AB/FrameStrobe[17]
+ Tile_X9Y12_LUT4AB/FrameStrobe[18] Tile_X9Y12_LUT4AB/FrameStrobe[19] Tile_X9Y12_LUT4AB/FrameStrobe[1]
+ Tile_X9Y12_LUT4AB/FrameStrobe[2] Tile_X9Y12_LUT4AB/FrameStrobe[3] Tile_X9Y12_LUT4AB/FrameStrobe[4]
+ Tile_X9Y12_LUT4AB/FrameStrobe[5] Tile_X9Y12_LUT4AB/FrameStrobe[6] Tile_X9Y12_LUT4AB/FrameStrobe[7]
+ Tile_X9Y12_LUT4AB/FrameStrobe[8] Tile_X9Y12_LUT4AB/FrameStrobe[9] Tile_X9Y11_LUT4AB/FrameStrobe[0]
+ Tile_X9Y11_LUT4AB/FrameStrobe[10] Tile_X9Y11_LUT4AB/FrameStrobe[11] Tile_X9Y11_LUT4AB/FrameStrobe[12]
+ Tile_X9Y11_LUT4AB/FrameStrobe[13] Tile_X9Y11_LUT4AB/FrameStrobe[14] Tile_X9Y11_LUT4AB/FrameStrobe[15]
+ Tile_X9Y11_LUT4AB/FrameStrobe[16] Tile_X9Y11_LUT4AB/FrameStrobe[17] Tile_X9Y11_LUT4AB/FrameStrobe[18]
+ Tile_X9Y11_LUT4AB/FrameStrobe[19] Tile_X9Y11_LUT4AB/FrameStrobe[1] Tile_X9Y11_LUT4AB/FrameStrobe[2]
+ Tile_X9Y11_LUT4AB/FrameStrobe[3] Tile_X9Y11_LUT4AB/FrameStrobe[4] Tile_X9Y11_LUT4AB/FrameStrobe[5]
+ Tile_X9Y11_LUT4AB/FrameStrobe[6] Tile_X9Y11_LUT4AB/FrameStrobe[7] Tile_X9Y11_LUT4AB/FrameStrobe[8]
+ Tile_X9Y11_LUT4AB/FrameStrobe[9] Tile_X9Y12_LUT4AB/N1BEG[0] Tile_X9Y12_LUT4AB/N1BEG[1]
+ Tile_X9Y12_LUT4AB/N1BEG[2] Tile_X9Y12_LUT4AB/N1BEG[3] Tile_X9Y13_LUT4AB/N1BEG[0]
+ Tile_X9Y13_LUT4AB/N1BEG[1] Tile_X9Y13_LUT4AB/N1BEG[2] Tile_X9Y13_LUT4AB/N1BEG[3]
+ Tile_X9Y12_LUT4AB/N2BEG[0] Tile_X9Y12_LUT4AB/N2BEG[1] Tile_X9Y12_LUT4AB/N2BEG[2]
+ Tile_X9Y12_LUT4AB/N2BEG[3] Tile_X9Y12_LUT4AB/N2BEG[4] Tile_X9Y12_LUT4AB/N2BEG[5]
+ Tile_X9Y12_LUT4AB/N2BEG[6] Tile_X9Y12_LUT4AB/N2BEG[7] Tile_X9Y11_LUT4AB/N2END[0]
+ Tile_X9Y11_LUT4AB/N2END[1] Tile_X9Y11_LUT4AB/N2END[2] Tile_X9Y11_LUT4AB/N2END[3]
+ Tile_X9Y11_LUT4AB/N2END[4] Tile_X9Y11_LUT4AB/N2END[5] Tile_X9Y11_LUT4AB/N2END[6]
+ Tile_X9Y11_LUT4AB/N2END[7] Tile_X9Y12_LUT4AB/N2END[0] Tile_X9Y12_LUT4AB/N2END[1]
+ Tile_X9Y12_LUT4AB/N2END[2] Tile_X9Y12_LUT4AB/N2END[3] Tile_X9Y12_LUT4AB/N2END[4]
+ Tile_X9Y12_LUT4AB/N2END[5] Tile_X9Y12_LUT4AB/N2END[6] Tile_X9Y12_LUT4AB/N2END[7]
+ Tile_X9Y13_LUT4AB/N2BEG[0] Tile_X9Y13_LUT4AB/N2BEG[1] Tile_X9Y13_LUT4AB/N2BEG[2]
+ Tile_X9Y13_LUT4AB/N2BEG[3] Tile_X9Y13_LUT4AB/N2BEG[4] Tile_X9Y13_LUT4AB/N2BEG[5]
+ Tile_X9Y13_LUT4AB/N2BEG[6] Tile_X9Y13_LUT4AB/N2BEG[7] Tile_X9Y12_LUT4AB/N4BEG[0]
+ Tile_X9Y12_LUT4AB/N4BEG[10] Tile_X9Y12_LUT4AB/N4BEG[11] Tile_X9Y12_LUT4AB/N4BEG[12]
+ Tile_X9Y12_LUT4AB/N4BEG[13] Tile_X9Y12_LUT4AB/N4BEG[14] Tile_X9Y12_LUT4AB/N4BEG[15]
+ Tile_X9Y12_LUT4AB/N4BEG[1] Tile_X9Y12_LUT4AB/N4BEG[2] Tile_X9Y12_LUT4AB/N4BEG[3]
+ Tile_X9Y12_LUT4AB/N4BEG[4] Tile_X9Y12_LUT4AB/N4BEG[5] Tile_X9Y12_LUT4AB/N4BEG[6]
+ Tile_X9Y12_LUT4AB/N4BEG[7] Tile_X9Y12_LUT4AB/N4BEG[8] Tile_X9Y12_LUT4AB/N4BEG[9]
+ Tile_X9Y13_LUT4AB/N4BEG[0] Tile_X9Y13_LUT4AB/N4BEG[10] Tile_X9Y13_LUT4AB/N4BEG[11]
+ Tile_X9Y13_LUT4AB/N4BEG[12] Tile_X9Y13_LUT4AB/N4BEG[13] Tile_X9Y13_LUT4AB/N4BEG[14]
+ Tile_X9Y13_LUT4AB/N4BEG[15] Tile_X9Y13_LUT4AB/N4BEG[1] Tile_X9Y13_LUT4AB/N4BEG[2]
+ Tile_X9Y13_LUT4AB/N4BEG[3] Tile_X9Y13_LUT4AB/N4BEG[4] Tile_X9Y13_LUT4AB/N4BEG[5]
+ Tile_X9Y13_LUT4AB/N4BEG[6] Tile_X9Y13_LUT4AB/N4BEG[7] Tile_X9Y13_LUT4AB/N4BEG[8]
+ Tile_X9Y13_LUT4AB/N4BEG[9] Tile_X9Y12_LUT4AB/NN4BEG[0] Tile_X9Y12_LUT4AB/NN4BEG[10]
+ Tile_X9Y12_LUT4AB/NN4BEG[11] Tile_X9Y12_LUT4AB/NN4BEG[12] Tile_X9Y12_LUT4AB/NN4BEG[13]
+ Tile_X9Y12_LUT4AB/NN4BEG[14] Tile_X9Y12_LUT4AB/NN4BEG[15] Tile_X9Y12_LUT4AB/NN4BEG[1]
+ Tile_X9Y12_LUT4AB/NN4BEG[2] Tile_X9Y12_LUT4AB/NN4BEG[3] Tile_X9Y12_LUT4AB/NN4BEG[4]
+ Tile_X9Y12_LUT4AB/NN4BEG[5] Tile_X9Y12_LUT4AB/NN4BEG[6] Tile_X9Y12_LUT4AB/NN4BEG[7]
+ Tile_X9Y12_LUT4AB/NN4BEG[8] Tile_X9Y12_LUT4AB/NN4BEG[9] Tile_X9Y13_LUT4AB/NN4BEG[0]
+ Tile_X9Y13_LUT4AB/NN4BEG[10] Tile_X9Y13_LUT4AB/NN4BEG[11] Tile_X9Y13_LUT4AB/NN4BEG[12]
+ Tile_X9Y13_LUT4AB/NN4BEG[13] Tile_X9Y13_LUT4AB/NN4BEG[14] Tile_X9Y13_LUT4AB/NN4BEG[15]
+ Tile_X9Y13_LUT4AB/NN4BEG[1] Tile_X9Y13_LUT4AB/NN4BEG[2] Tile_X9Y13_LUT4AB/NN4BEG[3]
+ Tile_X9Y13_LUT4AB/NN4BEG[4] Tile_X9Y13_LUT4AB/NN4BEG[5] Tile_X9Y13_LUT4AB/NN4BEG[6]
+ Tile_X9Y13_LUT4AB/NN4BEG[7] Tile_X9Y13_LUT4AB/NN4BEG[8] Tile_X9Y13_LUT4AB/NN4BEG[9]
+ Tile_X9Y13_LUT4AB/S1END[0] Tile_X9Y13_LUT4AB/S1END[1] Tile_X9Y13_LUT4AB/S1END[2]
+ Tile_X9Y13_LUT4AB/S1END[3] Tile_X9Y12_LUT4AB/S1END[0] Tile_X9Y12_LUT4AB/S1END[1]
+ Tile_X9Y12_LUT4AB/S1END[2] Tile_X9Y12_LUT4AB/S1END[3] Tile_X9Y13_LUT4AB/S2MID[0]
+ Tile_X9Y13_LUT4AB/S2MID[1] Tile_X9Y13_LUT4AB/S2MID[2] Tile_X9Y13_LUT4AB/S2MID[3]
+ Tile_X9Y13_LUT4AB/S2MID[4] Tile_X9Y13_LUT4AB/S2MID[5] Tile_X9Y13_LUT4AB/S2MID[6]
+ Tile_X9Y13_LUT4AB/S2MID[7] Tile_X9Y13_LUT4AB/S2END[0] Tile_X9Y13_LUT4AB/S2END[1]
+ Tile_X9Y13_LUT4AB/S2END[2] Tile_X9Y13_LUT4AB/S2END[3] Tile_X9Y13_LUT4AB/S2END[4]
+ Tile_X9Y13_LUT4AB/S2END[5] Tile_X9Y13_LUT4AB/S2END[6] Tile_X9Y13_LUT4AB/S2END[7]
+ Tile_X9Y12_LUT4AB/S2END[0] Tile_X9Y12_LUT4AB/S2END[1] Tile_X9Y12_LUT4AB/S2END[2]
+ Tile_X9Y12_LUT4AB/S2END[3] Tile_X9Y12_LUT4AB/S2END[4] Tile_X9Y12_LUT4AB/S2END[5]
+ Tile_X9Y12_LUT4AB/S2END[6] Tile_X9Y12_LUT4AB/S2END[7] Tile_X9Y12_LUT4AB/S2MID[0]
+ Tile_X9Y12_LUT4AB/S2MID[1] Tile_X9Y12_LUT4AB/S2MID[2] Tile_X9Y12_LUT4AB/S2MID[3]
+ Tile_X9Y12_LUT4AB/S2MID[4] Tile_X9Y12_LUT4AB/S2MID[5] Tile_X9Y12_LUT4AB/S2MID[6]
+ Tile_X9Y12_LUT4AB/S2MID[7] Tile_X9Y13_LUT4AB/S4END[0] Tile_X9Y13_LUT4AB/S4END[10]
+ Tile_X9Y13_LUT4AB/S4END[11] Tile_X9Y13_LUT4AB/S4END[12] Tile_X9Y13_LUT4AB/S4END[13]
+ Tile_X9Y13_LUT4AB/S4END[14] Tile_X9Y13_LUT4AB/S4END[15] Tile_X9Y13_LUT4AB/S4END[1]
+ Tile_X9Y13_LUT4AB/S4END[2] Tile_X9Y13_LUT4AB/S4END[3] Tile_X9Y13_LUT4AB/S4END[4]
+ Tile_X9Y13_LUT4AB/S4END[5] Tile_X9Y13_LUT4AB/S4END[6] Tile_X9Y13_LUT4AB/S4END[7]
+ Tile_X9Y13_LUT4AB/S4END[8] Tile_X9Y13_LUT4AB/S4END[9] Tile_X9Y12_LUT4AB/S4END[0]
+ Tile_X9Y12_LUT4AB/S4END[10] Tile_X9Y12_LUT4AB/S4END[11] Tile_X9Y12_LUT4AB/S4END[12]
+ Tile_X9Y12_LUT4AB/S4END[13] Tile_X9Y12_LUT4AB/S4END[14] Tile_X9Y12_LUT4AB/S4END[15]
+ Tile_X9Y12_LUT4AB/S4END[1] Tile_X9Y12_LUT4AB/S4END[2] Tile_X9Y12_LUT4AB/S4END[3]
+ Tile_X9Y12_LUT4AB/S4END[4] Tile_X9Y12_LUT4AB/S4END[5] Tile_X9Y12_LUT4AB/S4END[6]
+ Tile_X9Y12_LUT4AB/S4END[7] Tile_X9Y12_LUT4AB/S4END[8] Tile_X9Y12_LUT4AB/S4END[9]
+ Tile_X9Y13_LUT4AB/SS4END[0] Tile_X9Y13_LUT4AB/SS4END[10] Tile_X9Y13_LUT4AB/SS4END[11]
+ Tile_X9Y13_LUT4AB/SS4END[12] Tile_X9Y13_LUT4AB/SS4END[13] Tile_X9Y13_LUT4AB/SS4END[14]
+ Tile_X9Y13_LUT4AB/SS4END[15] Tile_X9Y13_LUT4AB/SS4END[1] Tile_X9Y13_LUT4AB/SS4END[2]
+ Tile_X9Y13_LUT4AB/SS4END[3] Tile_X9Y13_LUT4AB/SS4END[4] Tile_X9Y13_LUT4AB/SS4END[5]
+ Tile_X9Y13_LUT4AB/SS4END[6] Tile_X9Y13_LUT4AB/SS4END[7] Tile_X9Y13_LUT4AB/SS4END[8]
+ Tile_X9Y13_LUT4AB/SS4END[9] Tile_X9Y12_LUT4AB/SS4END[0] Tile_X9Y12_LUT4AB/SS4END[10]
+ Tile_X9Y12_LUT4AB/SS4END[11] Tile_X9Y12_LUT4AB/SS4END[12] Tile_X9Y12_LUT4AB/SS4END[13]
+ Tile_X9Y12_LUT4AB/SS4END[14] Tile_X9Y12_LUT4AB/SS4END[15] Tile_X9Y12_LUT4AB/SS4END[1]
+ Tile_X9Y12_LUT4AB/SS4END[2] Tile_X9Y12_LUT4AB/SS4END[3] Tile_X9Y12_LUT4AB/SS4END[4]
+ Tile_X9Y12_LUT4AB/SS4END[5] Tile_X9Y12_LUT4AB/SS4END[6] Tile_X9Y12_LUT4AB/SS4END[7]
+ Tile_X9Y12_LUT4AB/SS4END[8] Tile_X9Y12_LUT4AB/SS4END[9] Tile_X9Y12_LUT4AB/UserCLK
+ Tile_X9Y11_LUT4AB/UserCLK VGND VPWR Tile_X9Y12_LUT4AB/W1BEG[0] Tile_X9Y12_LUT4AB/W1BEG[1]
+ Tile_X9Y12_LUT4AB/W1BEG[2] Tile_X9Y12_LUT4AB/W1BEG[3] Tile_X9Y12_LUT4AB/W1END[0]
+ Tile_X9Y12_LUT4AB/W1END[1] Tile_X9Y12_LUT4AB/W1END[2] Tile_X9Y12_LUT4AB/W1END[3]
+ Tile_X9Y12_LUT4AB/W2BEG[0] Tile_X9Y12_LUT4AB/W2BEG[1] Tile_X9Y12_LUT4AB/W2BEG[2]
+ Tile_X9Y12_LUT4AB/W2BEG[3] Tile_X9Y12_LUT4AB/W2BEG[4] Tile_X9Y12_LUT4AB/W2BEG[5]
+ Tile_X9Y12_LUT4AB/W2BEG[6] Tile_X9Y12_LUT4AB/W2BEG[7] Tile_X8Y12_LUT4AB/W2END[0]
+ Tile_X8Y12_LUT4AB/W2END[1] Tile_X8Y12_LUT4AB/W2END[2] Tile_X8Y12_LUT4AB/W2END[3]
+ Tile_X8Y12_LUT4AB/W2END[4] Tile_X8Y12_LUT4AB/W2END[5] Tile_X8Y12_LUT4AB/W2END[6]
+ Tile_X8Y12_LUT4AB/W2END[7] Tile_X9Y12_LUT4AB/W2END[0] Tile_X9Y12_LUT4AB/W2END[1]
+ Tile_X9Y12_LUT4AB/W2END[2] Tile_X9Y12_LUT4AB/W2END[3] Tile_X9Y12_LUT4AB/W2END[4]
+ Tile_X9Y12_LUT4AB/W2END[5] Tile_X9Y12_LUT4AB/W2END[6] Tile_X9Y12_LUT4AB/W2END[7]
+ Tile_X9Y12_LUT4AB/W2MID[0] Tile_X9Y12_LUT4AB/W2MID[1] Tile_X9Y12_LUT4AB/W2MID[2]
+ Tile_X9Y12_LUT4AB/W2MID[3] Tile_X9Y12_LUT4AB/W2MID[4] Tile_X9Y12_LUT4AB/W2MID[5]
+ Tile_X9Y12_LUT4AB/W2MID[6] Tile_X9Y12_LUT4AB/W2MID[7] Tile_X9Y12_LUT4AB/W6BEG[0]
+ Tile_X9Y12_LUT4AB/W6BEG[10] Tile_X9Y12_LUT4AB/W6BEG[11] Tile_X9Y12_LUT4AB/W6BEG[1]
+ Tile_X9Y12_LUT4AB/W6BEG[2] Tile_X9Y12_LUT4AB/W6BEG[3] Tile_X9Y12_LUT4AB/W6BEG[4]
+ Tile_X9Y12_LUT4AB/W6BEG[5] Tile_X9Y12_LUT4AB/W6BEG[6] Tile_X9Y12_LUT4AB/W6BEG[7]
+ Tile_X9Y12_LUT4AB/W6BEG[8] Tile_X9Y12_LUT4AB/W6BEG[9] Tile_X9Y12_LUT4AB/W6END[0]
+ Tile_X9Y12_LUT4AB/W6END[10] Tile_X9Y12_LUT4AB/W6END[11] Tile_X9Y12_LUT4AB/W6END[1]
+ Tile_X9Y12_LUT4AB/W6END[2] Tile_X9Y12_LUT4AB/W6END[3] Tile_X9Y12_LUT4AB/W6END[4]
+ Tile_X9Y12_LUT4AB/W6END[5] Tile_X9Y12_LUT4AB/W6END[6] Tile_X9Y12_LUT4AB/W6END[7]
+ Tile_X9Y12_LUT4AB/W6END[8] Tile_X9Y12_LUT4AB/W6END[9] Tile_X9Y12_LUT4AB/WW4BEG[0]
+ Tile_X9Y12_LUT4AB/WW4BEG[10] Tile_X9Y12_LUT4AB/WW4BEG[11] Tile_X9Y12_LUT4AB/WW4BEG[12]
+ Tile_X9Y12_LUT4AB/WW4BEG[13] Tile_X9Y12_LUT4AB/WW4BEG[14] Tile_X9Y12_LUT4AB/WW4BEG[15]
+ Tile_X9Y12_LUT4AB/WW4BEG[1] Tile_X9Y12_LUT4AB/WW4BEG[2] Tile_X9Y12_LUT4AB/WW4BEG[3]
+ Tile_X9Y12_LUT4AB/WW4BEG[4] Tile_X9Y12_LUT4AB/WW4BEG[5] Tile_X9Y12_LUT4AB/WW4BEG[6]
+ Tile_X9Y12_LUT4AB/WW4BEG[7] Tile_X9Y12_LUT4AB/WW4BEG[8] Tile_X9Y12_LUT4AB/WW4BEG[9]
+ Tile_X9Y12_LUT4AB/WW4END[0] Tile_X9Y12_LUT4AB/WW4END[10] Tile_X9Y12_LUT4AB/WW4END[11]
+ Tile_X9Y12_LUT4AB/WW4END[12] Tile_X9Y12_LUT4AB/WW4END[13] Tile_X9Y12_LUT4AB/WW4END[14]
+ Tile_X9Y12_LUT4AB/WW4END[15] Tile_X9Y12_LUT4AB/WW4END[1] Tile_X9Y12_LUT4AB/WW4END[2]
+ Tile_X9Y12_LUT4AB/WW4END[3] Tile_X9Y12_LUT4AB/WW4END[4] Tile_X9Y12_LUT4AB/WW4END[5]
+ Tile_X9Y12_LUT4AB/WW4END[6] Tile_X9Y12_LUT4AB/WW4END[7] Tile_X9Y12_LUT4AB/WW4END[8]
+ Tile_X9Y12_LUT4AB/WW4END[9] LUT4AB
XTile_X7Y0_N_term_DSP Tile_X7Y0_N_term_DSP/FrameData[0] Tile_X7Y0_N_term_DSP/FrameData[10]
+ Tile_X7Y0_N_term_DSP/FrameData[11] Tile_X7Y0_N_term_DSP/FrameData[12] Tile_X7Y0_N_term_DSP/FrameData[13]
+ Tile_X7Y0_N_term_DSP/FrameData[14] Tile_X7Y0_N_term_DSP/FrameData[15] Tile_X7Y0_N_term_DSP/FrameData[16]
+ Tile_X7Y0_N_term_DSP/FrameData[17] Tile_X7Y0_N_term_DSP/FrameData[18] Tile_X7Y0_N_term_DSP/FrameData[19]
+ Tile_X7Y0_N_term_DSP/FrameData[1] Tile_X7Y0_N_term_DSP/FrameData[20] Tile_X7Y0_N_term_DSP/FrameData[21]
+ Tile_X7Y0_N_term_DSP/FrameData[22] Tile_X7Y0_N_term_DSP/FrameData[23] Tile_X7Y0_N_term_DSP/FrameData[24]
+ Tile_X7Y0_N_term_DSP/FrameData[25] Tile_X7Y0_N_term_DSP/FrameData[26] Tile_X7Y0_N_term_DSP/FrameData[27]
+ Tile_X7Y0_N_term_DSP/FrameData[28] Tile_X7Y0_N_term_DSP/FrameData[29] Tile_X7Y0_N_term_DSP/FrameData[2]
+ Tile_X7Y0_N_term_DSP/FrameData[30] Tile_X7Y0_N_term_DSP/FrameData[31] Tile_X7Y0_N_term_DSP/FrameData[3]
+ Tile_X7Y0_N_term_DSP/FrameData[4] Tile_X7Y0_N_term_DSP/FrameData[5] Tile_X7Y0_N_term_DSP/FrameData[6]
+ Tile_X7Y0_N_term_DSP/FrameData[7] Tile_X7Y0_N_term_DSP/FrameData[8] Tile_X7Y0_N_term_DSP/FrameData[9]
+ Tile_X7Y0_N_term_DSP/FrameData_O[0] Tile_X7Y0_N_term_DSP/FrameData_O[10] Tile_X7Y0_N_term_DSP/FrameData_O[11]
+ Tile_X7Y0_N_term_DSP/FrameData_O[12] Tile_X7Y0_N_term_DSP/FrameData_O[13] Tile_X7Y0_N_term_DSP/FrameData_O[14]
+ Tile_X7Y0_N_term_DSP/FrameData_O[15] Tile_X7Y0_N_term_DSP/FrameData_O[16] Tile_X7Y0_N_term_DSP/FrameData_O[17]
+ Tile_X7Y0_N_term_DSP/FrameData_O[18] Tile_X7Y0_N_term_DSP/FrameData_O[19] Tile_X7Y0_N_term_DSP/FrameData_O[1]
+ Tile_X7Y0_N_term_DSP/FrameData_O[20] Tile_X7Y0_N_term_DSP/FrameData_O[21] Tile_X7Y0_N_term_DSP/FrameData_O[22]
+ Tile_X7Y0_N_term_DSP/FrameData_O[23] Tile_X7Y0_N_term_DSP/FrameData_O[24] Tile_X7Y0_N_term_DSP/FrameData_O[25]
+ Tile_X7Y0_N_term_DSP/FrameData_O[26] Tile_X7Y0_N_term_DSP/FrameData_O[27] Tile_X7Y0_N_term_DSP/FrameData_O[28]
+ Tile_X7Y0_N_term_DSP/FrameData_O[29] Tile_X7Y0_N_term_DSP/FrameData_O[2] Tile_X7Y0_N_term_DSP/FrameData_O[30]
+ Tile_X7Y0_N_term_DSP/FrameData_O[31] Tile_X7Y0_N_term_DSP/FrameData_O[3] Tile_X7Y0_N_term_DSP/FrameData_O[4]
+ Tile_X7Y0_N_term_DSP/FrameData_O[5] Tile_X7Y0_N_term_DSP/FrameData_O[6] Tile_X7Y0_N_term_DSP/FrameData_O[7]
+ Tile_X7Y0_N_term_DSP/FrameData_O[8] Tile_X7Y0_N_term_DSP/FrameData_O[9] Tile_X7Y0_N_term_DSP/FrameStrobe[0]
+ Tile_X7Y0_N_term_DSP/FrameStrobe[10] Tile_X7Y0_N_term_DSP/FrameStrobe[11] Tile_X7Y0_N_term_DSP/FrameStrobe[12]
+ Tile_X7Y0_N_term_DSP/FrameStrobe[13] Tile_X7Y0_N_term_DSP/FrameStrobe[14] Tile_X7Y0_N_term_DSP/FrameStrobe[15]
+ Tile_X7Y0_N_term_DSP/FrameStrobe[16] Tile_X7Y0_N_term_DSP/FrameStrobe[17] Tile_X7Y0_N_term_DSP/FrameStrobe[18]
+ Tile_X7Y0_N_term_DSP/FrameStrobe[19] Tile_X7Y0_N_term_DSP/FrameStrobe[1] Tile_X7Y0_N_term_DSP/FrameStrobe[2]
+ Tile_X7Y0_N_term_DSP/FrameStrobe[3] Tile_X7Y0_N_term_DSP/FrameStrobe[4] Tile_X7Y0_N_term_DSP/FrameStrobe[5]
+ Tile_X7Y0_N_term_DSP/FrameStrobe[6] Tile_X7Y0_N_term_DSP/FrameStrobe[7] Tile_X7Y0_N_term_DSP/FrameStrobe[8]
+ Tile_X7Y0_N_term_DSP/FrameStrobe[9] Tile_X7Y0_N_term_DSP/FrameStrobe_O[0] Tile_X7Y0_N_term_DSP/FrameStrobe_O[10]
+ Tile_X7Y0_N_term_DSP/FrameStrobe_O[11] Tile_X7Y0_N_term_DSP/FrameStrobe_O[12] Tile_X7Y0_N_term_DSP/FrameStrobe_O[13]
+ Tile_X7Y0_N_term_DSP/FrameStrobe_O[14] Tile_X7Y0_N_term_DSP/FrameStrobe_O[15] Tile_X7Y0_N_term_DSP/FrameStrobe_O[16]
+ Tile_X7Y0_N_term_DSP/FrameStrobe_O[17] Tile_X7Y0_N_term_DSP/FrameStrobe_O[18] Tile_X7Y0_N_term_DSP/FrameStrobe_O[19]
+ Tile_X7Y0_N_term_DSP/FrameStrobe_O[1] Tile_X7Y0_N_term_DSP/FrameStrobe_O[2] Tile_X7Y0_N_term_DSP/FrameStrobe_O[3]
+ Tile_X7Y0_N_term_DSP/FrameStrobe_O[4] Tile_X7Y0_N_term_DSP/FrameStrobe_O[5] Tile_X7Y0_N_term_DSP/FrameStrobe_O[6]
+ Tile_X7Y0_N_term_DSP/FrameStrobe_O[7] Tile_X7Y0_N_term_DSP/FrameStrobe_O[8] Tile_X7Y0_N_term_DSP/FrameStrobe_O[9]
+ Tile_X7Y0_N_term_DSP/N1END[0] Tile_X7Y0_N_term_DSP/N1END[1] Tile_X7Y0_N_term_DSP/N1END[2]
+ Tile_X7Y0_N_term_DSP/N1END[3] Tile_X7Y0_N_term_DSP/N2END[0] Tile_X7Y0_N_term_DSP/N2END[1]
+ Tile_X7Y0_N_term_DSP/N2END[2] Tile_X7Y0_N_term_DSP/N2END[3] Tile_X7Y0_N_term_DSP/N2END[4]
+ Tile_X7Y0_N_term_DSP/N2END[5] Tile_X7Y0_N_term_DSP/N2END[6] Tile_X7Y0_N_term_DSP/N2END[7]
+ Tile_X7Y0_N_term_DSP/N2MID[0] Tile_X7Y0_N_term_DSP/N2MID[1] Tile_X7Y0_N_term_DSP/N2MID[2]
+ Tile_X7Y0_N_term_DSP/N2MID[3] Tile_X7Y0_N_term_DSP/N2MID[4] Tile_X7Y0_N_term_DSP/N2MID[5]
+ Tile_X7Y0_N_term_DSP/N2MID[6] Tile_X7Y0_N_term_DSP/N2MID[7] Tile_X7Y0_N_term_DSP/N4END[0]
+ Tile_X7Y0_N_term_DSP/N4END[10] Tile_X7Y0_N_term_DSP/N4END[11] Tile_X7Y0_N_term_DSP/N4END[12]
+ Tile_X7Y0_N_term_DSP/N4END[13] Tile_X7Y0_N_term_DSP/N4END[14] Tile_X7Y0_N_term_DSP/N4END[15]
+ Tile_X7Y0_N_term_DSP/N4END[1] Tile_X7Y0_N_term_DSP/N4END[2] Tile_X7Y0_N_term_DSP/N4END[3]
+ Tile_X7Y0_N_term_DSP/N4END[4] Tile_X7Y0_N_term_DSP/N4END[5] Tile_X7Y0_N_term_DSP/N4END[6]
+ Tile_X7Y0_N_term_DSP/N4END[7] Tile_X7Y0_N_term_DSP/N4END[8] Tile_X7Y0_N_term_DSP/N4END[9]
+ Tile_X7Y0_N_term_DSP/NN4END[0] Tile_X7Y0_N_term_DSP/NN4END[10] Tile_X7Y0_N_term_DSP/NN4END[11]
+ Tile_X7Y0_N_term_DSP/NN4END[12] Tile_X7Y0_N_term_DSP/NN4END[13] Tile_X7Y0_N_term_DSP/NN4END[14]
+ Tile_X7Y0_N_term_DSP/NN4END[15] Tile_X7Y0_N_term_DSP/NN4END[1] Tile_X7Y0_N_term_DSP/NN4END[2]
+ Tile_X7Y0_N_term_DSP/NN4END[3] Tile_X7Y0_N_term_DSP/NN4END[4] Tile_X7Y0_N_term_DSP/NN4END[5]
+ Tile_X7Y0_N_term_DSP/NN4END[6] Tile_X7Y0_N_term_DSP/NN4END[7] Tile_X7Y0_N_term_DSP/NN4END[8]
+ Tile_X7Y0_N_term_DSP/NN4END[9] Tile_X7Y0_N_term_DSP/S1BEG[0] Tile_X7Y0_N_term_DSP/S1BEG[1]
+ Tile_X7Y0_N_term_DSP/S1BEG[2] Tile_X7Y0_N_term_DSP/S1BEG[3] Tile_X7Y0_N_term_DSP/S2BEG[0]
+ Tile_X7Y0_N_term_DSP/S2BEG[1] Tile_X7Y0_N_term_DSP/S2BEG[2] Tile_X7Y0_N_term_DSP/S2BEG[3]
+ Tile_X7Y0_N_term_DSP/S2BEG[4] Tile_X7Y0_N_term_DSP/S2BEG[5] Tile_X7Y0_N_term_DSP/S2BEG[6]
+ Tile_X7Y0_N_term_DSP/S2BEG[7] Tile_X7Y0_N_term_DSP/S2BEGb[0] Tile_X7Y0_N_term_DSP/S2BEGb[1]
+ Tile_X7Y0_N_term_DSP/S2BEGb[2] Tile_X7Y0_N_term_DSP/S2BEGb[3] Tile_X7Y0_N_term_DSP/S2BEGb[4]
+ Tile_X7Y0_N_term_DSP/S2BEGb[5] Tile_X7Y0_N_term_DSP/S2BEGb[6] Tile_X7Y0_N_term_DSP/S2BEGb[7]
+ Tile_X7Y0_N_term_DSP/S4BEG[0] Tile_X7Y0_N_term_DSP/S4BEG[10] Tile_X7Y0_N_term_DSP/S4BEG[11]
+ Tile_X7Y0_N_term_DSP/S4BEG[12] Tile_X7Y0_N_term_DSP/S4BEG[13] Tile_X7Y0_N_term_DSP/S4BEG[14]
+ Tile_X7Y0_N_term_DSP/S4BEG[15] Tile_X7Y0_N_term_DSP/S4BEG[1] Tile_X7Y0_N_term_DSP/S4BEG[2]
+ Tile_X7Y0_N_term_DSP/S4BEG[3] Tile_X7Y0_N_term_DSP/S4BEG[4] Tile_X7Y0_N_term_DSP/S4BEG[5]
+ Tile_X7Y0_N_term_DSP/S4BEG[6] Tile_X7Y0_N_term_DSP/S4BEG[7] Tile_X7Y0_N_term_DSP/S4BEG[8]
+ Tile_X7Y0_N_term_DSP/S4BEG[9] Tile_X7Y0_N_term_DSP/SS4BEG[0] Tile_X7Y0_N_term_DSP/SS4BEG[10]
+ Tile_X7Y0_N_term_DSP/SS4BEG[11] Tile_X7Y0_N_term_DSP/SS4BEG[12] Tile_X7Y0_N_term_DSP/SS4BEG[13]
+ Tile_X7Y0_N_term_DSP/SS4BEG[14] Tile_X7Y0_N_term_DSP/SS4BEG[15] Tile_X7Y0_N_term_DSP/SS4BEG[1]
+ Tile_X7Y0_N_term_DSP/SS4BEG[2] Tile_X7Y0_N_term_DSP/SS4BEG[3] Tile_X7Y0_N_term_DSP/SS4BEG[4]
+ Tile_X7Y0_N_term_DSP/SS4BEG[5] Tile_X7Y0_N_term_DSP/SS4BEG[6] Tile_X7Y0_N_term_DSP/SS4BEG[7]
+ Tile_X7Y0_N_term_DSP/SS4BEG[8] Tile_X7Y0_N_term_DSP/SS4BEG[9] Tile_X7Y0_N_term_DSP/UserCLK
+ Tile_X7Y0_N_term_DSP/UserCLKo VGND VPWR N_term_DSP
XTile_X3Y8_LUT4AB Tile_X3Y9_LUT4AB/Co Tile_X3Y8_LUT4AB/Co Tile_X3Y8_LUT4AB/E1BEG[0]
+ Tile_X3Y8_LUT4AB/E1BEG[1] Tile_X3Y8_LUT4AB/E1BEG[2] Tile_X3Y8_LUT4AB/E1BEG[3] Tile_X3Y8_LUT4AB/E1END[0]
+ Tile_X3Y8_LUT4AB/E1END[1] Tile_X3Y8_LUT4AB/E1END[2] Tile_X3Y8_LUT4AB/E1END[3] Tile_X3Y8_LUT4AB/E2BEG[0]
+ Tile_X3Y8_LUT4AB/E2BEG[1] Tile_X3Y8_LUT4AB/E2BEG[2] Tile_X3Y8_LUT4AB/E2BEG[3] Tile_X3Y8_LUT4AB/E2BEG[4]
+ Tile_X3Y8_LUT4AB/E2BEG[5] Tile_X3Y8_LUT4AB/E2BEG[6] Tile_X3Y8_LUT4AB/E2BEG[7] Tile_X4Y8_RegFile/E2END[0]
+ Tile_X4Y8_RegFile/E2END[1] Tile_X4Y8_RegFile/E2END[2] Tile_X4Y8_RegFile/E2END[3]
+ Tile_X4Y8_RegFile/E2END[4] Tile_X4Y8_RegFile/E2END[5] Tile_X4Y8_RegFile/E2END[6]
+ Tile_X4Y8_RegFile/E2END[7] Tile_X3Y8_LUT4AB/E2END[0] Tile_X3Y8_LUT4AB/E2END[1] Tile_X3Y8_LUT4AB/E2END[2]
+ Tile_X3Y8_LUT4AB/E2END[3] Tile_X3Y8_LUT4AB/E2END[4] Tile_X3Y8_LUT4AB/E2END[5] Tile_X3Y8_LUT4AB/E2END[6]
+ Tile_X3Y8_LUT4AB/E2END[7] Tile_X3Y8_LUT4AB/E2MID[0] Tile_X3Y8_LUT4AB/E2MID[1] Tile_X3Y8_LUT4AB/E2MID[2]
+ Tile_X3Y8_LUT4AB/E2MID[3] Tile_X3Y8_LUT4AB/E2MID[4] Tile_X3Y8_LUT4AB/E2MID[5] Tile_X3Y8_LUT4AB/E2MID[6]
+ Tile_X3Y8_LUT4AB/E2MID[7] Tile_X3Y8_LUT4AB/E6BEG[0] Tile_X3Y8_LUT4AB/E6BEG[10] Tile_X3Y8_LUT4AB/E6BEG[11]
+ Tile_X3Y8_LUT4AB/E6BEG[1] Tile_X3Y8_LUT4AB/E6BEG[2] Tile_X3Y8_LUT4AB/E6BEG[3] Tile_X3Y8_LUT4AB/E6BEG[4]
+ Tile_X3Y8_LUT4AB/E6BEG[5] Tile_X3Y8_LUT4AB/E6BEG[6] Tile_X3Y8_LUT4AB/E6BEG[7] Tile_X3Y8_LUT4AB/E6BEG[8]
+ Tile_X3Y8_LUT4AB/E6BEG[9] Tile_X3Y8_LUT4AB/E6END[0] Tile_X3Y8_LUT4AB/E6END[10] Tile_X3Y8_LUT4AB/E6END[11]
+ Tile_X3Y8_LUT4AB/E6END[1] Tile_X3Y8_LUT4AB/E6END[2] Tile_X3Y8_LUT4AB/E6END[3] Tile_X3Y8_LUT4AB/E6END[4]
+ Tile_X3Y8_LUT4AB/E6END[5] Tile_X3Y8_LUT4AB/E6END[6] Tile_X3Y8_LUT4AB/E6END[7] Tile_X3Y8_LUT4AB/E6END[8]
+ Tile_X3Y8_LUT4AB/E6END[9] Tile_X3Y8_LUT4AB/EE4BEG[0] Tile_X3Y8_LUT4AB/EE4BEG[10]
+ Tile_X3Y8_LUT4AB/EE4BEG[11] Tile_X3Y8_LUT4AB/EE4BEG[12] Tile_X3Y8_LUT4AB/EE4BEG[13]
+ Tile_X3Y8_LUT4AB/EE4BEG[14] Tile_X3Y8_LUT4AB/EE4BEG[15] Tile_X3Y8_LUT4AB/EE4BEG[1]
+ Tile_X3Y8_LUT4AB/EE4BEG[2] Tile_X3Y8_LUT4AB/EE4BEG[3] Tile_X3Y8_LUT4AB/EE4BEG[4]
+ Tile_X3Y8_LUT4AB/EE4BEG[5] Tile_X3Y8_LUT4AB/EE4BEG[6] Tile_X3Y8_LUT4AB/EE4BEG[7]
+ Tile_X3Y8_LUT4AB/EE4BEG[8] Tile_X3Y8_LUT4AB/EE4BEG[9] Tile_X3Y8_LUT4AB/EE4END[0]
+ Tile_X3Y8_LUT4AB/EE4END[10] Tile_X3Y8_LUT4AB/EE4END[11] Tile_X3Y8_LUT4AB/EE4END[12]
+ Tile_X3Y8_LUT4AB/EE4END[13] Tile_X3Y8_LUT4AB/EE4END[14] Tile_X3Y8_LUT4AB/EE4END[15]
+ Tile_X3Y8_LUT4AB/EE4END[1] Tile_X3Y8_LUT4AB/EE4END[2] Tile_X3Y8_LUT4AB/EE4END[3]
+ Tile_X3Y8_LUT4AB/EE4END[4] Tile_X3Y8_LUT4AB/EE4END[5] Tile_X3Y8_LUT4AB/EE4END[6]
+ Tile_X3Y8_LUT4AB/EE4END[7] Tile_X3Y8_LUT4AB/EE4END[8] Tile_X3Y8_LUT4AB/EE4END[9]
+ Tile_X3Y8_LUT4AB/FrameData[0] Tile_X3Y8_LUT4AB/FrameData[10] Tile_X3Y8_LUT4AB/FrameData[11]
+ Tile_X3Y8_LUT4AB/FrameData[12] Tile_X3Y8_LUT4AB/FrameData[13] Tile_X3Y8_LUT4AB/FrameData[14]
+ Tile_X3Y8_LUT4AB/FrameData[15] Tile_X3Y8_LUT4AB/FrameData[16] Tile_X3Y8_LUT4AB/FrameData[17]
+ Tile_X3Y8_LUT4AB/FrameData[18] Tile_X3Y8_LUT4AB/FrameData[19] Tile_X3Y8_LUT4AB/FrameData[1]
+ Tile_X3Y8_LUT4AB/FrameData[20] Tile_X3Y8_LUT4AB/FrameData[21] Tile_X3Y8_LUT4AB/FrameData[22]
+ Tile_X3Y8_LUT4AB/FrameData[23] Tile_X3Y8_LUT4AB/FrameData[24] Tile_X3Y8_LUT4AB/FrameData[25]
+ Tile_X3Y8_LUT4AB/FrameData[26] Tile_X3Y8_LUT4AB/FrameData[27] Tile_X3Y8_LUT4AB/FrameData[28]
+ Tile_X3Y8_LUT4AB/FrameData[29] Tile_X3Y8_LUT4AB/FrameData[2] Tile_X3Y8_LUT4AB/FrameData[30]
+ Tile_X3Y8_LUT4AB/FrameData[31] Tile_X3Y8_LUT4AB/FrameData[3] Tile_X3Y8_LUT4AB/FrameData[4]
+ Tile_X3Y8_LUT4AB/FrameData[5] Tile_X3Y8_LUT4AB/FrameData[6] Tile_X3Y8_LUT4AB/FrameData[7]
+ Tile_X3Y8_LUT4AB/FrameData[8] Tile_X3Y8_LUT4AB/FrameData[9] Tile_X4Y8_RegFile/FrameData[0]
+ Tile_X4Y8_RegFile/FrameData[10] Tile_X4Y8_RegFile/FrameData[11] Tile_X4Y8_RegFile/FrameData[12]
+ Tile_X4Y8_RegFile/FrameData[13] Tile_X4Y8_RegFile/FrameData[14] Tile_X4Y8_RegFile/FrameData[15]
+ Tile_X4Y8_RegFile/FrameData[16] Tile_X4Y8_RegFile/FrameData[17] Tile_X4Y8_RegFile/FrameData[18]
+ Tile_X4Y8_RegFile/FrameData[19] Tile_X4Y8_RegFile/FrameData[1] Tile_X4Y8_RegFile/FrameData[20]
+ Tile_X4Y8_RegFile/FrameData[21] Tile_X4Y8_RegFile/FrameData[22] Tile_X4Y8_RegFile/FrameData[23]
+ Tile_X4Y8_RegFile/FrameData[24] Tile_X4Y8_RegFile/FrameData[25] Tile_X4Y8_RegFile/FrameData[26]
+ Tile_X4Y8_RegFile/FrameData[27] Tile_X4Y8_RegFile/FrameData[28] Tile_X4Y8_RegFile/FrameData[29]
+ Tile_X4Y8_RegFile/FrameData[2] Tile_X4Y8_RegFile/FrameData[30] Tile_X4Y8_RegFile/FrameData[31]
+ Tile_X4Y8_RegFile/FrameData[3] Tile_X4Y8_RegFile/FrameData[4] Tile_X4Y8_RegFile/FrameData[5]
+ Tile_X4Y8_RegFile/FrameData[6] Tile_X4Y8_RegFile/FrameData[7] Tile_X4Y8_RegFile/FrameData[8]
+ Tile_X4Y8_RegFile/FrameData[9] Tile_X3Y8_LUT4AB/FrameStrobe[0] Tile_X3Y8_LUT4AB/FrameStrobe[10]
+ Tile_X3Y8_LUT4AB/FrameStrobe[11] Tile_X3Y8_LUT4AB/FrameStrobe[12] Tile_X3Y8_LUT4AB/FrameStrobe[13]
+ Tile_X3Y8_LUT4AB/FrameStrobe[14] Tile_X3Y8_LUT4AB/FrameStrobe[15] Tile_X3Y8_LUT4AB/FrameStrobe[16]
+ Tile_X3Y8_LUT4AB/FrameStrobe[17] Tile_X3Y8_LUT4AB/FrameStrobe[18] Tile_X3Y8_LUT4AB/FrameStrobe[19]
+ Tile_X3Y8_LUT4AB/FrameStrobe[1] Tile_X3Y8_LUT4AB/FrameStrobe[2] Tile_X3Y8_LUT4AB/FrameStrobe[3]
+ Tile_X3Y8_LUT4AB/FrameStrobe[4] Tile_X3Y8_LUT4AB/FrameStrobe[5] Tile_X3Y8_LUT4AB/FrameStrobe[6]
+ Tile_X3Y8_LUT4AB/FrameStrobe[7] Tile_X3Y8_LUT4AB/FrameStrobe[8] Tile_X3Y8_LUT4AB/FrameStrobe[9]
+ Tile_X3Y7_LUT4AB/FrameStrobe[0] Tile_X3Y7_LUT4AB/FrameStrobe[10] Tile_X3Y7_LUT4AB/FrameStrobe[11]
+ Tile_X3Y7_LUT4AB/FrameStrobe[12] Tile_X3Y7_LUT4AB/FrameStrobe[13] Tile_X3Y7_LUT4AB/FrameStrobe[14]
+ Tile_X3Y7_LUT4AB/FrameStrobe[15] Tile_X3Y7_LUT4AB/FrameStrobe[16] Tile_X3Y7_LUT4AB/FrameStrobe[17]
+ Tile_X3Y7_LUT4AB/FrameStrobe[18] Tile_X3Y7_LUT4AB/FrameStrobe[19] Tile_X3Y7_LUT4AB/FrameStrobe[1]
+ Tile_X3Y7_LUT4AB/FrameStrobe[2] Tile_X3Y7_LUT4AB/FrameStrobe[3] Tile_X3Y7_LUT4AB/FrameStrobe[4]
+ Tile_X3Y7_LUT4AB/FrameStrobe[5] Tile_X3Y7_LUT4AB/FrameStrobe[6] Tile_X3Y7_LUT4AB/FrameStrobe[7]
+ Tile_X3Y7_LUT4AB/FrameStrobe[8] Tile_X3Y7_LUT4AB/FrameStrobe[9] Tile_X3Y8_LUT4AB/N1BEG[0]
+ Tile_X3Y8_LUT4AB/N1BEG[1] Tile_X3Y8_LUT4AB/N1BEG[2] Tile_X3Y8_LUT4AB/N1BEG[3] Tile_X3Y9_LUT4AB/N1BEG[0]
+ Tile_X3Y9_LUT4AB/N1BEG[1] Tile_X3Y9_LUT4AB/N1BEG[2] Tile_X3Y9_LUT4AB/N1BEG[3] Tile_X3Y8_LUT4AB/N2BEG[0]
+ Tile_X3Y8_LUT4AB/N2BEG[1] Tile_X3Y8_LUT4AB/N2BEG[2] Tile_X3Y8_LUT4AB/N2BEG[3] Tile_X3Y8_LUT4AB/N2BEG[4]
+ Tile_X3Y8_LUT4AB/N2BEG[5] Tile_X3Y8_LUT4AB/N2BEG[6] Tile_X3Y8_LUT4AB/N2BEG[7] Tile_X3Y7_LUT4AB/N2END[0]
+ Tile_X3Y7_LUT4AB/N2END[1] Tile_X3Y7_LUT4AB/N2END[2] Tile_X3Y7_LUT4AB/N2END[3] Tile_X3Y7_LUT4AB/N2END[4]
+ Tile_X3Y7_LUT4AB/N2END[5] Tile_X3Y7_LUT4AB/N2END[6] Tile_X3Y7_LUT4AB/N2END[7] Tile_X3Y8_LUT4AB/N2END[0]
+ Tile_X3Y8_LUT4AB/N2END[1] Tile_X3Y8_LUT4AB/N2END[2] Tile_X3Y8_LUT4AB/N2END[3] Tile_X3Y8_LUT4AB/N2END[4]
+ Tile_X3Y8_LUT4AB/N2END[5] Tile_X3Y8_LUT4AB/N2END[6] Tile_X3Y8_LUT4AB/N2END[7] Tile_X3Y9_LUT4AB/N2BEG[0]
+ Tile_X3Y9_LUT4AB/N2BEG[1] Tile_X3Y9_LUT4AB/N2BEG[2] Tile_X3Y9_LUT4AB/N2BEG[3] Tile_X3Y9_LUT4AB/N2BEG[4]
+ Tile_X3Y9_LUT4AB/N2BEG[5] Tile_X3Y9_LUT4AB/N2BEG[6] Tile_X3Y9_LUT4AB/N2BEG[7] Tile_X3Y8_LUT4AB/N4BEG[0]
+ Tile_X3Y8_LUT4AB/N4BEG[10] Tile_X3Y8_LUT4AB/N4BEG[11] Tile_X3Y8_LUT4AB/N4BEG[12]
+ Tile_X3Y8_LUT4AB/N4BEG[13] Tile_X3Y8_LUT4AB/N4BEG[14] Tile_X3Y8_LUT4AB/N4BEG[15]
+ Tile_X3Y8_LUT4AB/N4BEG[1] Tile_X3Y8_LUT4AB/N4BEG[2] Tile_X3Y8_LUT4AB/N4BEG[3] Tile_X3Y8_LUT4AB/N4BEG[4]
+ Tile_X3Y8_LUT4AB/N4BEG[5] Tile_X3Y8_LUT4AB/N4BEG[6] Tile_X3Y8_LUT4AB/N4BEG[7] Tile_X3Y8_LUT4AB/N4BEG[8]
+ Tile_X3Y8_LUT4AB/N4BEG[9] Tile_X3Y9_LUT4AB/N4BEG[0] Tile_X3Y9_LUT4AB/N4BEG[10] Tile_X3Y9_LUT4AB/N4BEG[11]
+ Tile_X3Y9_LUT4AB/N4BEG[12] Tile_X3Y9_LUT4AB/N4BEG[13] Tile_X3Y9_LUT4AB/N4BEG[14]
+ Tile_X3Y9_LUT4AB/N4BEG[15] Tile_X3Y9_LUT4AB/N4BEG[1] Tile_X3Y9_LUT4AB/N4BEG[2] Tile_X3Y9_LUT4AB/N4BEG[3]
+ Tile_X3Y9_LUT4AB/N4BEG[4] Tile_X3Y9_LUT4AB/N4BEG[5] Tile_X3Y9_LUT4AB/N4BEG[6] Tile_X3Y9_LUT4AB/N4BEG[7]
+ Tile_X3Y9_LUT4AB/N4BEG[8] Tile_X3Y9_LUT4AB/N4BEG[9] Tile_X3Y8_LUT4AB/NN4BEG[0] Tile_X3Y8_LUT4AB/NN4BEG[10]
+ Tile_X3Y8_LUT4AB/NN4BEG[11] Tile_X3Y8_LUT4AB/NN4BEG[12] Tile_X3Y8_LUT4AB/NN4BEG[13]
+ Tile_X3Y8_LUT4AB/NN4BEG[14] Tile_X3Y8_LUT4AB/NN4BEG[15] Tile_X3Y8_LUT4AB/NN4BEG[1]
+ Tile_X3Y8_LUT4AB/NN4BEG[2] Tile_X3Y8_LUT4AB/NN4BEG[3] Tile_X3Y8_LUT4AB/NN4BEG[4]
+ Tile_X3Y8_LUT4AB/NN4BEG[5] Tile_X3Y8_LUT4AB/NN4BEG[6] Tile_X3Y8_LUT4AB/NN4BEG[7]
+ Tile_X3Y8_LUT4AB/NN4BEG[8] Tile_X3Y8_LUT4AB/NN4BEG[9] Tile_X3Y9_LUT4AB/NN4BEG[0]
+ Tile_X3Y9_LUT4AB/NN4BEG[10] Tile_X3Y9_LUT4AB/NN4BEG[11] Tile_X3Y9_LUT4AB/NN4BEG[12]
+ Tile_X3Y9_LUT4AB/NN4BEG[13] Tile_X3Y9_LUT4AB/NN4BEG[14] Tile_X3Y9_LUT4AB/NN4BEG[15]
+ Tile_X3Y9_LUT4AB/NN4BEG[1] Tile_X3Y9_LUT4AB/NN4BEG[2] Tile_X3Y9_LUT4AB/NN4BEG[3]
+ Tile_X3Y9_LUT4AB/NN4BEG[4] Tile_X3Y9_LUT4AB/NN4BEG[5] Tile_X3Y9_LUT4AB/NN4BEG[6]
+ Tile_X3Y9_LUT4AB/NN4BEG[7] Tile_X3Y9_LUT4AB/NN4BEG[8] Tile_X3Y9_LUT4AB/NN4BEG[9]
+ Tile_X3Y9_LUT4AB/S1END[0] Tile_X3Y9_LUT4AB/S1END[1] Tile_X3Y9_LUT4AB/S1END[2] Tile_X3Y9_LUT4AB/S1END[3]
+ Tile_X3Y8_LUT4AB/S1END[0] Tile_X3Y8_LUT4AB/S1END[1] Tile_X3Y8_LUT4AB/S1END[2] Tile_X3Y8_LUT4AB/S1END[3]
+ Tile_X3Y9_LUT4AB/S2MID[0] Tile_X3Y9_LUT4AB/S2MID[1] Tile_X3Y9_LUT4AB/S2MID[2] Tile_X3Y9_LUT4AB/S2MID[3]
+ Tile_X3Y9_LUT4AB/S2MID[4] Tile_X3Y9_LUT4AB/S2MID[5] Tile_X3Y9_LUT4AB/S2MID[6] Tile_X3Y9_LUT4AB/S2MID[7]
+ Tile_X3Y9_LUT4AB/S2END[0] Tile_X3Y9_LUT4AB/S2END[1] Tile_X3Y9_LUT4AB/S2END[2] Tile_X3Y9_LUT4AB/S2END[3]
+ Tile_X3Y9_LUT4AB/S2END[4] Tile_X3Y9_LUT4AB/S2END[5] Tile_X3Y9_LUT4AB/S2END[6] Tile_X3Y9_LUT4AB/S2END[7]
+ Tile_X3Y8_LUT4AB/S2END[0] Tile_X3Y8_LUT4AB/S2END[1] Tile_X3Y8_LUT4AB/S2END[2] Tile_X3Y8_LUT4AB/S2END[3]
+ Tile_X3Y8_LUT4AB/S2END[4] Tile_X3Y8_LUT4AB/S2END[5] Tile_X3Y8_LUT4AB/S2END[6] Tile_X3Y8_LUT4AB/S2END[7]
+ Tile_X3Y8_LUT4AB/S2MID[0] Tile_X3Y8_LUT4AB/S2MID[1] Tile_X3Y8_LUT4AB/S2MID[2] Tile_X3Y8_LUT4AB/S2MID[3]
+ Tile_X3Y8_LUT4AB/S2MID[4] Tile_X3Y8_LUT4AB/S2MID[5] Tile_X3Y8_LUT4AB/S2MID[6] Tile_X3Y8_LUT4AB/S2MID[7]
+ Tile_X3Y9_LUT4AB/S4END[0] Tile_X3Y9_LUT4AB/S4END[10] Tile_X3Y9_LUT4AB/S4END[11]
+ Tile_X3Y9_LUT4AB/S4END[12] Tile_X3Y9_LUT4AB/S4END[13] Tile_X3Y9_LUT4AB/S4END[14]
+ Tile_X3Y9_LUT4AB/S4END[15] Tile_X3Y9_LUT4AB/S4END[1] Tile_X3Y9_LUT4AB/S4END[2] Tile_X3Y9_LUT4AB/S4END[3]
+ Tile_X3Y9_LUT4AB/S4END[4] Tile_X3Y9_LUT4AB/S4END[5] Tile_X3Y9_LUT4AB/S4END[6] Tile_X3Y9_LUT4AB/S4END[7]
+ Tile_X3Y9_LUT4AB/S4END[8] Tile_X3Y9_LUT4AB/S4END[9] Tile_X3Y8_LUT4AB/S4END[0] Tile_X3Y8_LUT4AB/S4END[10]
+ Tile_X3Y8_LUT4AB/S4END[11] Tile_X3Y8_LUT4AB/S4END[12] Tile_X3Y8_LUT4AB/S4END[13]
+ Tile_X3Y8_LUT4AB/S4END[14] Tile_X3Y8_LUT4AB/S4END[15] Tile_X3Y8_LUT4AB/S4END[1]
+ Tile_X3Y8_LUT4AB/S4END[2] Tile_X3Y8_LUT4AB/S4END[3] Tile_X3Y8_LUT4AB/S4END[4] Tile_X3Y8_LUT4AB/S4END[5]
+ Tile_X3Y8_LUT4AB/S4END[6] Tile_X3Y8_LUT4AB/S4END[7] Tile_X3Y8_LUT4AB/S4END[8] Tile_X3Y8_LUT4AB/S4END[9]
+ Tile_X3Y9_LUT4AB/SS4END[0] Tile_X3Y9_LUT4AB/SS4END[10] Tile_X3Y9_LUT4AB/SS4END[11]
+ Tile_X3Y9_LUT4AB/SS4END[12] Tile_X3Y9_LUT4AB/SS4END[13] Tile_X3Y9_LUT4AB/SS4END[14]
+ Tile_X3Y9_LUT4AB/SS4END[15] Tile_X3Y9_LUT4AB/SS4END[1] Tile_X3Y9_LUT4AB/SS4END[2]
+ Tile_X3Y9_LUT4AB/SS4END[3] Tile_X3Y9_LUT4AB/SS4END[4] Tile_X3Y9_LUT4AB/SS4END[5]
+ Tile_X3Y9_LUT4AB/SS4END[6] Tile_X3Y9_LUT4AB/SS4END[7] Tile_X3Y9_LUT4AB/SS4END[8]
+ Tile_X3Y9_LUT4AB/SS4END[9] Tile_X3Y8_LUT4AB/SS4END[0] Tile_X3Y8_LUT4AB/SS4END[10]
+ Tile_X3Y8_LUT4AB/SS4END[11] Tile_X3Y8_LUT4AB/SS4END[12] Tile_X3Y8_LUT4AB/SS4END[13]
+ Tile_X3Y8_LUT4AB/SS4END[14] Tile_X3Y8_LUT4AB/SS4END[15] Tile_X3Y8_LUT4AB/SS4END[1]
+ Tile_X3Y8_LUT4AB/SS4END[2] Tile_X3Y8_LUT4AB/SS4END[3] Tile_X3Y8_LUT4AB/SS4END[4]
+ Tile_X3Y8_LUT4AB/SS4END[5] Tile_X3Y8_LUT4AB/SS4END[6] Tile_X3Y8_LUT4AB/SS4END[7]
+ Tile_X3Y8_LUT4AB/SS4END[8] Tile_X3Y8_LUT4AB/SS4END[9] Tile_X3Y8_LUT4AB/UserCLK Tile_X3Y7_LUT4AB/UserCLK
+ VGND VPWR Tile_X3Y8_LUT4AB/W1BEG[0] Tile_X3Y8_LUT4AB/W1BEG[1] Tile_X3Y8_LUT4AB/W1BEG[2]
+ Tile_X3Y8_LUT4AB/W1BEG[3] Tile_X3Y8_LUT4AB/W1END[0] Tile_X3Y8_LUT4AB/W1END[1] Tile_X3Y8_LUT4AB/W1END[2]
+ Tile_X3Y8_LUT4AB/W1END[3] Tile_X3Y8_LUT4AB/W2BEG[0] Tile_X3Y8_LUT4AB/W2BEG[1] Tile_X3Y8_LUT4AB/W2BEG[2]
+ Tile_X3Y8_LUT4AB/W2BEG[3] Tile_X3Y8_LUT4AB/W2BEG[4] Tile_X3Y8_LUT4AB/W2BEG[5] Tile_X3Y8_LUT4AB/W2BEG[6]
+ Tile_X3Y8_LUT4AB/W2BEG[7] Tile_X2Y8_LUT4AB/W2END[0] Tile_X2Y8_LUT4AB/W2END[1] Tile_X2Y8_LUT4AB/W2END[2]
+ Tile_X2Y8_LUT4AB/W2END[3] Tile_X2Y8_LUT4AB/W2END[4] Tile_X2Y8_LUT4AB/W2END[5] Tile_X2Y8_LUT4AB/W2END[6]
+ Tile_X2Y8_LUT4AB/W2END[7] Tile_X3Y8_LUT4AB/W2END[0] Tile_X3Y8_LUT4AB/W2END[1] Tile_X3Y8_LUT4AB/W2END[2]
+ Tile_X3Y8_LUT4AB/W2END[3] Tile_X3Y8_LUT4AB/W2END[4] Tile_X3Y8_LUT4AB/W2END[5] Tile_X3Y8_LUT4AB/W2END[6]
+ Tile_X3Y8_LUT4AB/W2END[7] Tile_X3Y8_LUT4AB/W2MID[0] Tile_X3Y8_LUT4AB/W2MID[1] Tile_X3Y8_LUT4AB/W2MID[2]
+ Tile_X3Y8_LUT4AB/W2MID[3] Tile_X3Y8_LUT4AB/W2MID[4] Tile_X3Y8_LUT4AB/W2MID[5] Tile_X3Y8_LUT4AB/W2MID[6]
+ Tile_X3Y8_LUT4AB/W2MID[7] Tile_X3Y8_LUT4AB/W6BEG[0] Tile_X3Y8_LUT4AB/W6BEG[10] Tile_X3Y8_LUT4AB/W6BEG[11]
+ Tile_X3Y8_LUT4AB/W6BEG[1] Tile_X3Y8_LUT4AB/W6BEG[2] Tile_X3Y8_LUT4AB/W6BEG[3] Tile_X3Y8_LUT4AB/W6BEG[4]
+ Tile_X3Y8_LUT4AB/W6BEG[5] Tile_X3Y8_LUT4AB/W6BEG[6] Tile_X3Y8_LUT4AB/W6BEG[7] Tile_X3Y8_LUT4AB/W6BEG[8]
+ Tile_X3Y8_LUT4AB/W6BEG[9] Tile_X3Y8_LUT4AB/W6END[0] Tile_X3Y8_LUT4AB/W6END[10] Tile_X3Y8_LUT4AB/W6END[11]
+ Tile_X3Y8_LUT4AB/W6END[1] Tile_X3Y8_LUT4AB/W6END[2] Tile_X3Y8_LUT4AB/W6END[3] Tile_X3Y8_LUT4AB/W6END[4]
+ Tile_X3Y8_LUT4AB/W6END[5] Tile_X3Y8_LUT4AB/W6END[6] Tile_X3Y8_LUT4AB/W6END[7] Tile_X3Y8_LUT4AB/W6END[8]
+ Tile_X3Y8_LUT4AB/W6END[9] Tile_X3Y8_LUT4AB/WW4BEG[0] Tile_X3Y8_LUT4AB/WW4BEG[10]
+ Tile_X3Y8_LUT4AB/WW4BEG[11] Tile_X3Y8_LUT4AB/WW4BEG[12] Tile_X3Y8_LUT4AB/WW4BEG[13]
+ Tile_X3Y8_LUT4AB/WW4BEG[14] Tile_X3Y8_LUT4AB/WW4BEG[15] Tile_X3Y8_LUT4AB/WW4BEG[1]
+ Tile_X3Y8_LUT4AB/WW4BEG[2] Tile_X3Y8_LUT4AB/WW4BEG[3] Tile_X3Y8_LUT4AB/WW4BEG[4]
+ Tile_X3Y8_LUT4AB/WW4BEG[5] Tile_X3Y8_LUT4AB/WW4BEG[6] Tile_X3Y8_LUT4AB/WW4BEG[7]
+ Tile_X3Y8_LUT4AB/WW4BEG[8] Tile_X3Y8_LUT4AB/WW4BEG[9] Tile_X3Y8_LUT4AB/WW4END[0]
+ Tile_X3Y8_LUT4AB/WW4END[10] Tile_X3Y8_LUT4AB/WW4END[11] Tile_X3Y8_LUT4AB/WW4END[12]
+ Tile_X3Y8_LUT4AB/WW4END[13] Tile_X3Y8_LUT4AB/WW4END[14] Tile_X3Y8_LUT4AB/WW4END[15]
+ Tile_X3Y8_LUT4AB/WW4END[1] Tile_X3Y8_LUT4AB/WW4END[2] Tile_X3Y8_LUT4AB/WW4END[3]
+ Tile_X3Y8_LUT4AB/WW4END[4] Tile_X3Y8_LUT4AB/WW4END[5] Tile_X3Y8_LUT4AB/WW4END[6]
+ Tile_X3Y8_LUT4AB/WW4END[7] Tile_X3Y8_LUT4AB/WW4END[8] Tile_X3Y8_LUT4AB/WW4END[9]
+ LUT4AB
XTile_X0Y11_W_IO Tile_X0Y11_A_I_top Tile_X0Y11_A_O_top Tile_X0Y11_A_T_top Tile_X0Y11_A_config_C_bit0
+ Tile_X0Y11_A_config_C_bit1 Tile_X0Y11_A_config_C_bit2 Tile_X0Y11_A_config_C_bit3
+ Tile_X0Y11_B_I_top Tile_X0Y11_B_O_top Tile_X0Y11_B_T_top Tile_X0Y11_B_config_C_bit0
+ Tile_X0Y11_B_config_C_bit1 Tile_X0Y11_B_config_C_bit2 Tile_X0Y11_B_config_C_bit3
+ Tile_X0Y11_W_IO/E1BEG[0] Tile_X0Y11_W_IO/E1BEG[1] Tile_X0Y11_W_IO/E1BEG[2] Tile_X0Y11_W_IO/E1BEG[3]
+ Tile_X0Y11_W_IO/E2BEG[0] Tile_X0Y11_W_IO/E2BEG[1] Tile_X0Y11_W_IO/E2BEG[2] Tile_X0Y11_W_IO/E2BEG[3]
+ Tile_X0Y11_W_IO/E2BEG[4] Tile_X0Y11_W_IO/E2BEG[5] Tile_X0Y11_W_IO/E2BEG[6] Tile_X0Y11_W_IO/E2BEG[7]
+ Tile_X0Y11_W_IO/E2BEGb[0] Tile_X0Y11_W_IO/E2BEGb[1] Tile_X0Y11_W_IO/E2BEGb[2] Tile_X0Y11_W_IO/E2BEGb[3]
+ Tile_X0Y11_W_IO/E2BEGb[4] Tile_X0Y11_W_IO/E2BEGb[5] Tile_X0Y11_W_IO/E2BEGb[6] Tile_X0Y11_W_IO/E2BEGb[7]
+ Tile_X0Y11_W_IO/E6BEG[0] Tile_X0Y11_W_IO/E6BEG[10] Tile_X0Y11_W_IO/E6BEG[11] Tile_X0Y11_W_IO/E6BEG[1]
+ Tile_X0Y11_W_IO/E6BEG[2] Tile_X0Y11_W_IO/E6BEG[3] Tile_X0Y11_W_IO/E6BEG[4] Tile_X0Y11_W_IO/E6BEG[5]
+ Tile_X0Y11_W_IO/E6BEG[6] Tile_X0Y11_W_IO/E6BEG[7] Tile_X0Y11_W_IO/E6BEG[8] Tile_X0Y11_W_IO/E6BEG[9]
+ Tile_X0Y11_W_IO/EE4BEG[0] Tile_X0Y11_W_IO/EE4BEG[10] Tile_X0Y11_W_IO/EE4BEG[11]
+ Tile_X0Y11_W_IO/EE4BEG[12] Tile_X0Y11_W_IO/EE4BEG[13] Tile_X0Y11_W_IO/EE4BEG[14]
+ Tile_X0Y11_W_IO/EE4BEG[15] Tile_X0Y11_W_IO/EE4BEG[1] Tile_X0Y11_W_IO/EE4BEG[2] Tile_X0Y11_W_IO/EE4BEG[3]
+ Tile_X0Y11_W_IO/EE4BEG[4] Tile_X0Y11_W_IO/EE4BEG[5] Tile_X0Y11_W_IO/EE4BEG[6] Tile_X0Y11_W_IO/EE4BEG[7]
+ Tile_X0Y11_W_IO/EE4BEG[8] Tile_X0Y11_W_IO/EE4BEG[9] FrameData[352] FrameData[362]
+ FrameData[363] FrameData[364] FrameData[365] FrameData[366] FrameData[367] FrameData[368]
+ FrameData[369] FrameData[370] FrameData[371] FrameData[353] FrameData[372] FrameData[373]
+ FrameData[374] FrameData[375] FrameData[376] FrameData[377] FrameData[378] FrameData[379]
+ FrameData[380] FrameData[381] FrameData[354] FrameData[382] FrameData[383] FrameData[355]
+ FrameData[356] FrameData[357] FrameData[358] FrameData[359] FrameData[360] FrameData[361]
+ Tile_X1Y11_LUT4AB/FrameData[0] Tile_X1Y11_LUT4AB/FrameData[10] Tile_X1Y11_LUT4AB/FrameData[11]
+ Tile_X1Y11_LUT4AB/FrameData[12] Tile_X1Y11_LUT4AB/FrameData[13] Tile_X1Y11_LUT4AB/FrameData[14]
+ Tile_X1Y11_LUT4AB/FrameData[15] Tile_X1Y11_LUT4AB/FrameData[16] Tile_X1Y11_LUT4AB/FrameData[17]
+ Tile_X1Y11_LUT4AB/FrameData[18] Tile_X1Y11_LUT4AB/FrameData[19] Tile_X1Y11_LUT4AB/FrameData[1]
+ Tile_X1Y11_LUT4AB/FrameData[20] Tile_X1Y11_LUT4AB/FrameData[21] Tile_X1Y11_LUT4AB/FrameData[22]
+ Tile_X1Y11_LUT4AB/FrameData[23] Tile_X1Y11_LUT4AB/FrameData[24] Tile_X1Y11_LUT4AB/FrameData[25]
+ Tile_X1Y11_LUT4AB/FrameData[26] Tile_X1Y11_LUT4AB/FrameData[27] Tile_X1Y11_LUT4AB/FrameData[28]
+ Tile_X1Y11_LUT4AB/FrameData[29] Tile_X1Y11_LUT4AB/FrameData[2] Tile_X1Y11_LUT4AB/FrameData[30]
+ Tile_X1Y11_LUT4AB/FrameData[31] Tile_X1Y11_LUT4AB/FrameData[3] Tile_X1Y11_LUT4AB/FrameData[4]
+ Tile_X1Y11_LUT4AB/FrameData[5] Tile_X1Y11_LUT4AB/FrameData[6] Tile_X1Y11_LUT4AB/FrameData[7]
+ Tile_X1Y11_LUT4AB/FrameData[8] Tile_X1Y11_LUT4AB/FrameData[9] Tile_X0Y11_W_IO/FrameStrobe[0]
+ Tile_X0Y11_W_IO/FrameStrobe[10] Tile_X0Y11_W_IO/FrameStrobe[11] Tile_X0Y11_W_IO/FrameStrobe[12]
+ Tile_X0Y11_W_IO/FrameStrobe[13] Tile_X0Y11_W_IO/FrameStrobe[14] Tile_X0Y11_W_IO/FrameStrobe[15]
+ Tile_X0Y11_W_IO/FrameStrobe[16] Tile_X0Y11_W_IO/FrameStrobe[17] Tile_X0Y11_W_IO/FrameStrobe[18]
+ Tile_X0Y11_W_IO/FrameStrobe[19] Tile_X0Y11_W_IO/FrameStrobe[1] Tile_X0Y11_W_IO/FrameStrobe[2]
+ Tile_X0Y11_W_IO/FrameStrobe[3] Tile_X0Y11_W_IO/FrameStrobe[4] Tile_X0Y11_W_IO/FrameStrobe[5]
+ Tile_X0Y11_W_IO/FrameStrobe[6] Tile_X0Y11_W_IO/FrameStrobe[7] Tile_X0Y11_W_IO/FrameStrobe[8]
+ Tile_X0Y11_W_IO/FrameStrobe[9] Tile_X0Y10_W_IO/FrameStrobe[0] Tile_X0Y10_W_IO/FrameStrobe[10]
+ Tile_X0Y10_W_IO/FrameStrobe[11] Tile_X0Y10_W_IO/FrameStrobe[12] Tile_X0Y10_W_IO/FrameStrobe[13]
+ Tile_X0Y10_W_IO/FrameStrobe[14] Tile_X0Y10_W_IO/FrameStrobe[15] Tile_X0Y10_W_IO/FrameStrobe[16]
+ Tile_X0Y10_W_IO/FrameStrobe[17] Tile_X0Y10_W_IO/FrameStrobe[18] Tile_X0Y10_W_IO/FrameStrobe[19]
+ Tile_X0Y10_W_IO/FrameStrobe[1] Tile_X0Y10_W_IO/FrameStrobe[2] Tile_X0Y10_W_IO/FrameStrobe[3]
+ Tile_X0Y10_W_IO/FrameStrobe[4] Tile_X0Y10_W_IO/FrameStrobe[5] Tile_X0Y10_W_IO/FrameStrobe[6]
+ Tile_X0Y10_W_IO/FrameStrobe[7] Tile_X0Y10_W_IO/FrameStrobe[8] Tile_X0Y10_W_IO/FrameStrobe[9]
+ Tile_X0Y11_W_IO/UserCLK Tile_X0Y10_W_IO/UserCLK VGND VPWR Tile_X0Y11_W_IO/W1END[0]
+ Tile_X0Y11_W_IO/W1END[1] Tile_X0Y11_W_IO/W1END[2] Tile_X0Y11_W_IO/W1END[3] Tile_X0Y11_W_IO/W2END[0]
+ Tile_X0Y11_W_IO/W2END[1] Tile_X0Y11_W_IO/W2END[2] Tile_X0Y11_W_IO/W2END[3] Tile_X0Y11_W_IO/W2END[4]
+ Tile_X0Y11_W_IO/W2END[5] Tile_X0Y11_W_IO/W2END[6] Tile_X0Y11_W_IO/W2END[7] Tile_X0Y11_W_IO/W2MID[0]
+ Tile_X0Y11_W_IO/W2MID[1] Tile_X0Y11_W_IO/W2MID[2] Tile_X0Y11_W_IO/W2MID[3] Tile_X0Y11_W_IO/W2MID[4]
+ Tile_X0Y11_W_IO/W2MID[5] Tile_X0Y11_W_IO/W2MID[6] Tile_X0Y11_W_IO/W2MID[7] Tile_X0Y11_W_IO/W6END[0]
+ Tile_X0Y11_W_IO/W6END[10] Tile_X0Y11_W_IO/W6END[11] Tile_X0Y11_W_IO/W6END[1] Tile_X0Y11_W_IO/W6END[2]
+ Tile_X0Y11_W_IO/W6END[3] Tile_X0Y11_W_IO/W6END[4] Tile_X0Y11_W_IO/W6END[5] Tile_X0Y11_W_IO/W6END[6]
+ Tile_X0Y11_W_IO/W6END[7] Tile_X0Y11_W_IO/W6END[8] Tile_X0Y11_W_IO/W6END[9] Tile_X0Y11_W_IO/WW4END[0]
+ Tile_X0Y11_W_IO/WW4END[10] Tile_X0Y11_W_IO/WW4END[11] Tile_X0Y11_W_IO/WW4END[12]
+ Tile_X0Y11_W_IO/WW4END[13] Tile_X0Y11_W_IO/WW4END[14] Tile_X0Y11_W_IO/WW4END[15]
+ Tile_X0Y11_W_IO/WW4END[1] Tile_X0Y11_W_IO/WW4END[2] Tile_X0Y11_W_IO/WW4END[3] Tile_X0Y11_W_IO/WW4END[4]
+ Tile_X0Y11_W_IO/WW4END[5] Tile_X0Y11_W_IO/WW4END[6] Tile_X0Y11_W_IO/WW4END[7] Tile_X0Y11_W_IO/WW4END[8]
+ Tile_X0Y11_W_IO/WW4END[9] W_IO
XTile_X4Y0_N_term_single2 Tile_X4Y0_N_term_single2/FrameData[0] Tile_X4Y0_N_term_single2/FrameData[10]
+ Tile_X4Y0_N_term_single2/FrameData[11] Tile_X4Y0_N_term_single2/FrameData[12] Tile_X4Y0_N_term_single2/FrameData[13]
+ Tile_X4Y0_N_term_single2/FrameData[14] Tile_X4Y0_N_term_single2/FrameData[15] Tile_X4Y0_N_term_single2/FrameData[16]
+ Tile_X4Y0_N_term_single2/FrameData[17] Tile_X4Y0_N_term_single2/FrameData[18] Tile_X4Y0_N_term_single2/FrameData[19]
+ Tile_X4Y0_N_term_single2/FrameData[1] Tile_X4Y0_N_term_single2/FrameData[20] Tile_X4Y0_N_term_single2/FrameData[21]
+ Tile_X4Y0_N_term_single2/FrameData[22] Tile_X4Y0_N_term_single2/FrameData[23] Tile_X4Y0_N_term_single2/FrameData[24]
+ Tile_X4Y0_N_term_single2/FrameData[25] Tile_X4Y0_N_term_single2/FrameData[26] Tile_X4Y0_N_term_single2/FrameData[27]
+ Tile_X4Y0_N_term_single2/FrameData[28] Tile_X4Y0_N_term_single2/FrameData[29] Tile_X4Y0_N_term_single2/FrameData[2]
+ Tile_X4Y0_N_term_single2/FrameData[30] Tile_X4Y0_N_term_single2/FrameData[31] Tile_X4Y0_N_term_single2/FrameData[3]
+ Tile_X4Y0_N_term_single2/FrameData[4] Tile_X4Y0_N_term_single2/FrameData[5] Tile_X4Y0_N_term_single2/FrameData[6]
+ Tile_X4Y0_N_term_single2/FrameData[7] Tile_X4Y0_N_term_single2/FrameData[8] Tile_X4Y0_N_term_single2/FrameData[9]
+ Tile_X5Y0_N_term_single/FrameData[0] Tile_X5Y0_N_term_single/FrameData[10] Tile_X5Y0_N_term_single/FrameData[11]
+ Tile_X5Y0_N_term_single/FrameData[12] Tile_X5Y0_N_term_single/FrameData[13] Tile_X5Y0_N_term_single/FrameData[14]
+ Tile_X5Y0_N_term_single/FrameData[15] Tile_X5Y0_N_term_single/FrameData[16] Tile_X5Y0_N_term_single/FrameData[17]
+ Tile_X5Y0_N_term_single/FrameData[18] Tile_X5Y0_N_term_single/FrameData[19] Tile_X5Y0_N_term_single/FrameData[1]
+ Tile_X5Y0_N_term_single/FrameData[20] Tile_X5Y0_N_term_single/FrameData[21] Tile_X5Y0_N_term_single/FrameData[22]
+ Tile_X5Y0_N_term_single/FrameData[23] Tile_X5Y0_N_term_single/FrameData[24] Tile_X5Y0_N_term_single/FrameData[25]
+ Tile_X5Y0_N_term_single/FrameData[26] Tile_X5Y0_N_term_single/FrameData[27] Tile_X5Y0_N_term_single/FrameData[28]
+ Tile_X5Y0_N_term_single/FrameData[29] Tile_X5Y0_N_term_single/FrameData[2] Tile_X5Y0_N_term_single/FrameData[30]
+ Tile_X5Y0_N_term_single/FrameData[31] Tile_X5Y0_N_term_single/FrameData[3] Tile_X5Y0_N_term_single/FrameData[4]
+ Tile_X5Y0_N_term_single/FrameData[5] Tile_X5Y0_N_term_single/FrameData[6] Tile_X5Y0_N_term_single/FrameData[7]
+ Tile_X5Y0_N_term_single/FrameData[8] Tile_X5Y0_N_term_single/FrameData[9] Tile_X4Y1_RegFile/FrameStrobe_O[0]
+ Tile_X4Y1_RegFile/FrameStrobe_O[10] Tile_X4Y1_RegFile/FrameStrobe_O[11] Tile_X4Y1_RegFile/FrameStrobe_O[12]
+ Tile_X4Y1_RegFile/FrameStrobe_O[13] Tile_X4Y1_RegFile/FrameStrobe_O[14] Tile_X4Y1_RegFile/FrameStrobe_O[15]
+ Tile_X4Y1_RegFile/FrameStrobe_O[16] Tile_X4Y1_RegFile/FrameStrobe_O[17] Tile_X4Y1_RegFile/FrameStrobe_O[18]
+ Tile_X4Y1_RegFile/FrameStrobe_O[19] Tile_X4Y1_RegFile/FrameStrobe_O[1] Tile_X4Y1_RegFile/FrameStrobe_O[2]
+ Tile_X4Y1_RegFile/FrameStrobe_O[3] Tile_X4Y1_RegFile/FrameStrobe_O[4] Tile_X4Y1_RegFile/FrameStrobe_O[5]
+ Tile_X4Y1_RegFile/FrameStrobe_O[6] Tile_X4Y1_RegFile/FrameStrobe_O[7] Tile_X4Y1_RegFile/FrameStrobe_O[8]
+ Tile_X4Y1_RegFile/FrameStrobe_O[9] Tile_X4Y0_N_term_single2/FrameStrobe_O[0] Tile_X4Y0_N_term_single2/FrameStrobe_O[10]
+ Tile_X4Y0_N_term_single2/FrameStrobe_O[11] Tile_X4Y0_N_term_single2/FrameStrobe_O[12]
+ Tile_X4Y0_N_term_single2/FrameStrobe_O[13] Tile_X4Y0_N_term_single2/FrameStrobe_O[14]
+ Tile_X4Y0_N_term_single2/FrameStrobe_O[15] Tile_X4Y0_N_term_single2/FrameStrobe_O[16]
+ Tile_X4Y0_N_term_single2/FrameStrobe_O[17] Tile_X4Y0_N_term_single2/FrameStrobe_O[18]
+ Tile_X4Y0_N_term_single2/FrameStrobe_O[19] Tile_X4Y0_N_term_single2/FrameStrobe_O[1]
+ Tile_X4Y0_N_term_single2/FrameStrobe_O[2] Tile_X4Y0_N_term_single2/FrameStrobe_O[3]
+ Tile_X4Y0_N_term_single2/FrameStrobe_O[4] Tile_X4Y0_N_term_single2/FrameStrobe_O[5]
+ Tile_X4Y0_N_term_single2/FrameStrobe_O[6] Tile_X4Y0_N_term_single2/FrameStrobe_O[7]
+ Tile_X4Y0_N_term_single2/FrameStrobe_O[8] Tile_X4Y0_N_term_single2/FrameStrobe_O[9]
+ Tile_X4Y1_RegFile/N1BEG[0] Tile_X4Y1_RegFile/N1BEG[1] Tile_X4Y1_RegFile/N1BEG[2]
+ Tile_X4Y1_RegFile/N1BEG[3] Tile_X4Y1_RegFile/N2BEGb[0] Tile_X4Y1_RegFile/N2BEGb[1]
+ Tile_X4Y1_RegFile/N2BEGb[2] Tile_X4Y1_RegFile/N2BEGb[3] Tile_X4Y1_RegFile/N2BEGb[4]
+ Tile_X4Y1_RegFile/N2BEGb[5] Tile_X4Y1_RegFile/N2BEGb[6] Tile_X4Y1_RegFile/N2BEGb[7]
+ Tile_X4Y1_RegFile/N2BEG[0] Tile_X4Y1_RegFile/N2BEG[1] Tile_X4Y1_RegFile/N2BEG[2]
+ Tile_X4Y1_RegFile/N2BEG[3] Tile_X4Y1_RegFile/N2BEG[4] Tile_X4Y1_RegFile/N2BEG[5]
+ Tile_X4Y1_RegFile/N2BEG[6] Tile_X4Y1_RegFile/N2BEG[7] Tile_X4Y1_RegFile/N4BEG[0]
+ Tile_X4Y1_RegFile/N4BEG[10] Tile_X4Y1_RegFile/N4BEG[11] Tile_X4Y1_RegFile/N4BEG[12]
+ Tile_X4Y1_RegFile/N4BEG[13] Tile_X4Y1_RegFile/N4BEG[14] Tile_X4Y1_RegFile/N4BEG[15]
+ Tile_X4Y1_RegFile/N4BEG[1] Tile_X4Y1_RegFile/N4BEG[2] Tile_X4Y1_RegFile/N4BEG[3]
+ Tile_X4Y1_RegFile/N4BEG[4] Tile_X4Y1_RegFile/N4BEG[5] Tile_X4Y1_RegFile/N4BEG[6]
+ Tile_X4Y1_RegFile/N4BEG[7] Tile_X4Y1_RegFile/N4BEG[8] Tile_X4Y1_RegFile/N4BEG[9]
+ Tile_X4Y1_RegFile/NN4BEG[0] Tile_X4Y1_RegFile/NN4BEG[10] Tile_X4Y1_RegFile/NN4BEG[11]
+ Tile_X4Y1_RegFile/NN4BEG[12] Tile_X4Y1_RegFile/NN4BEG[13] Tile_X4Y1_RegFile/NN4BEG[14]
+ Tile_X4Y1_RegFile/NN4BEG[15] Tile_X4Y1_RegFile/NN4BEG[1] Tile_X4Y1_RegFile/NN4BEG[2]
+ Tile_X4Y1_RegFile/NN4BEG[3] Tile_X4Y1_RegFile/NN4BEG[4] Tile_X4Y1_RegFile/NN4BEG[5]
+ Tile_X4Y1_RegFile/NN4BEG[6] Tile_X4Y1_RegFile/NN4BEG[7] Tile_X4Y1_RegFile/NN4BEG[8]
+ Tile_X4Y1_RegFile/NN4BEG[9] Tile_X4Y1_RegFile/S1END[0] Tile_X4Y1_RegFile/S1END[1]
+ Tile_X4Y1_RegFile/S1END[2] Tile_X4Y1_RegFile/S1END[3] Tile_X4Y1_RegFile/S2MID[0]
+ Tile_X4Y1_RegFile/S2MID[1] Tile_X4Y1_RegFile/S2MID[2] Tile_X4Y1_RegFile/S2MID[3]
+ Tile_X4Y1_RegFile/S2MID[4] Tile_X4Y1_RegFile/S2MID[5] Tile_X4Y1_RegFile/S2MID[6]
+ Tile_X4Y1_RegFile/S2MID[7] Tile_X4Y1_RegFile/S2END[0] Tile_X4Y1_RegFile/S2END[1]
+ Tile_X4Y1_RegFile/S2END[2] Tile_X4Y1_RegFile/S2END[3] Tile_X4Y1_RegFile/S2END[4]
+ Tile_X4Y1_RegFile/S2END[5] Tile_X4Y1_RegFile/S2END[6] Tile_X4Y1_RegFile/S2END[7]
+ Tile_X4Y1_RegFile/S4END[0] Tile_X4Y1_RegFile/S4END[10] Tile_X4Y1_RegFile/S4END[11]
+ Tile_X4Y1_RegFile/S4END[12] Tile_X4Y1_RegFile/S4END[13] Tile_X4Y1_RegFile/S4END[14]
+ Tile_X4Y1_RegFile/S4END[15] Tile_X4Y1_RegFile/S4END[1] Tile_X4Y1_RegFile/S4END[2]
+ Tile_X4Y1_RegFile/S4END[3] Tile_X4Y1_RegFile/S4END[4] Tile_X4Y1_RegFile/S4END[5]
+ Tile_X4Y1_RegFile/S4END[6] Tile_X4Y1_RegFile/S4END[7] Tile_X4Y1_RegFile/S4END[8]
+ Tile_X4Y1_RegFile/S4END[9] Tile_X4Y1_RegFile/SS4END[0] Tile_X4Y1_RegFile/SS4END[10]
+ Tile_X4Y1_RegFile/SS4END[11] Tile_X4Y1_RegFile/SS4END[12] Tile_X4Y1_RegFile/SS4END[13]
+ Tile_X4Y1_RegFile/SS4END[14] Tile_X4Y1_RegFile/SS4END[15] Tile_X4Y1_RegFile/SS4END[1]
+ Tile_X4Y1_RegFile/SS4END[2] Tile_X4Y1_RegFile/SS4END[3] Tile_X4Y1_RegFile/SS4END[4]
+ Tile_X4Y1_RegFile/SS4END[5] Tile_X4Y1_RegFile/SS4END[6] Tile_X4Y1_RegFile/SS4END[7]
+ Tile_X4Y1_RegFile/SS4END[8] Tile_X4Y1_RegFile/SS4END[9] Tile_X4Y1_RegFile/UserCLKo
+ Tile_X4Y0_N_term_single2/UserCLKo VGND VPWR N_term_single2
XTile_X6Y2_LUT4AB Tile_X6Y3_LUT4AB/Co Tile_X6Y2_LUT4AB/Co Tile_X6Y2_LUT4AB/E1BEG[0]
+ Tile_X6Y2_LUT4AB/E1BEG[1] Tile_X6Y2_LUT4AB/E1BEG[2] Tile_X6Y2_LUT4AB/E1BEG[3] Tile_X6Y2_LUT4AB/E1END[0]
+ Tile_X6Y2_LUT4AB/E1END[1] Tile_X6Y2_LUT4AB/E1END[2] Tile_X6Y2_LUT4AB/E1END[3] Tile_X6Y2_LUT4AB/E2BEG[0]
+ Tile_X6Y2_LUT4AB/E2BEG[1] Tile_X6Y2_LUT4AB/E2BEG[2] Tile_X6Y2_LUT4AB/E2BEG[3] Tile_X6Y2_LUT4AB/E2BEG[4]
+ Tile_X6Y2_LUT4AB/E2BEG[5] Tile_X6Y2_LUT4AB/E2BEG[6] Tile_X6Y2_LUT4AB/E2BEG[7] Tile_X6Y2_LUT4AB/E2BEGb[0]
+ Tile_X6Y2_LUT4AB/E2BEGb[1] Tile_X6Y2_LUT4AB/E2BEGb[2] Tile_X6Y2_LUT4AB/E2BEGb[3]
+ Tile_X6Y2_LUT4AB/E2BEGb[4] Tile_X6Y2_LUT4AB/E2BEGb[5] Tile_X6Y2_LUT4AB/E2BEGb[6]
+ Tile_X6Y2_LUT4AB/E2BEGb[7] Tile_X6Y2_LUT4AB/E2END[0] Tile_X6Y2_LUT4AB/E2END[1] Tile_X6Y2_LUT4AB/E2END[2]
+ Tile_X6Y2_LUT4AB/E2END[3] Tile_X6Y2_LUT4AB/E2END[4] Tile_X6Y2_LUT4AB/E2END[5] Tile_X6Y2_LUT4AB/E2END[6]
+ Tile_X6Y2_LUT4AB/E2END[7] Tile_X6Y2_LUT4AB/E2MID[0] Tile_X6Y2_LUT4AB/E2MID[1] Tile_X6Y2_LUT4AB/E2MID[2]
+ Tile_X6Y2_LUT4AB/E2MID[3] Tile_X6Y2_LUT4AB/E2MID[4] Tile_X6Y2_LUT4AB/E2MID[5] Tile_X6Y2_LUT4AB/E2MID[6]
+ Tile_X6Y2_LUT4AB/E2MID[7] Tile_X6Y2_LUT4AB/E6BEG[0] Tile_X6Y2_LUT4AB/E6BEG[10] Tile_X6Y2_LUT4AB/E6BEG[11]
+ Tile_X6Y2_LUT4AB/E6BEG[1] Tile_X6Y2_LUT4AB/E6BEG[2] Tile_X6Y2_LUT4AB/E6BEG[3] Tile_X6Y2_LUT4AB/E6BEG[4]
+ Tile_X6Y2_LUT4AB/E6BEG[5] Tile_X6Y2_LUT4AB/E6BEG[6] Tile_X6Y2_LUT4AB/E6BEG[7] Tile_X6Y2_LUT4AB/E6BEG[8]
+ Tile_X6Y2_LUT4AB/E6BEG[9] Tile_X6Y2_LUT4AB/E6END[0] Tile_X6Y2_LUT4AB/E6END[10] Tile_X6Y2_LUT4AB/E6END[11]
+ Tile_X6Y2_LUT4AB/E6END[1] Tile_X6Y2_LUT4AB/E6END[2] Tile_X6Y2_LUT4AB/E6END[3] Tile_X6Y2_LUT4AB/E6END[4]
+ Tile_X6Y2_LUT4AB/E6END[5] Tile_X6Y2_LUT4AB/E6END[6] Tile_X6Y2_LUT4AB/E6END[7] Tile_X6Y2_LUT4AB/E6END[8]
+ Tile_X6Y2_LUT4AB/E6END[9] Tile_X6Y2_LUT4AB/EE4BEG[0] Tile_X6Y2_LUT4AB/EE4BEG[10]
+ Tile_X6Y2_LUT4AB/EE4BEG[11] Tile_X6Y2_LUT4AB/EE4BEG[12] Tile_X6Y2_LUT4AB/EE4BEG[13]
+ Tile_X6Y2_LUT4AB/EE4BEG[14] Tile_X6Y2_LUT4AB/EE4BEG[15] Tile_X6Y2_LUT4AB/EE4BEG[1]
+ Tile_X6Y2_LUT4AB/EE4BEG[2] Tile_X6Y2_LUT4AB/EE4BEG[3] Tile_X6Y2_LUT4AB/EE4BEG[4]
+ Tile_X6Y2_LUT4AB/EE4BEG[5] Tile_X6Y2_LUT4AB/EE4BEG[6] Tile_X6Y2_LUT4AB/EE4BEG[7]
+ Tile_X6Y2_LUT4AB/EE4BEG[8] Tile_X6Y2_LUT4AB/EE4BEG[9] Tile_X6Y2_LUT4AB/EE4END[0]
+ Tile_X6Y2_LUT4AB/EE4END[10] Tile_X6Y2_LUT4AB/EE4END[11] Tile_X6Y2_LUT4AB/EE4END[12]
+ Tile_X6Y2_LUT4AB/EE4END[13] Tile_X6Y2_LUT4AB/EE4END[14] Tile_X6Y2_LUT4AB/EE4END[15]
+ Tile_X6Y2_LUT4AB/EE4END[1] Tile_X6Y2_LUT4AB/EE4END[2] Tile_X6Y2_LUT4AB/EE4END[3]
+ Tile_X6Y2_LUT4AB/EE4END[4] Tile_X6Y2_LUT4AB/EE4END[5] Tile_X6Y2_LUT4AB/EE4END[6]
+ Tile_X6Y2_LUT4AB/EE4END[7] Tile_X6Y2_LUT4AB/EE4END[8] Tile_X6Y2_LUT4AB/EE4END[9]
+ Tile_X6Y2_LUT4AB/FrameData[0] Tile_X6Y2_LUT4AB/FrameData[10] Tile_X6Y2_LUT4AB/FrameData[11]
+ Tile_X6Y2_LUT4AB/FrameData[12] Tile_X6Y2_LUT4AB/FrameData[13] Tile_X6Y2_LUT4AB/FrameData[14]
+ Tile_X6Y2_LUT4AB/FrameData[15] Tile_X6Y2_LUT4AB/FrameData[16] Tile_X6Y2_LUT4AB/FrameData[17]
+ Tile_X6Y2_LUT4AB/FrameData[18] Tile_X6Y2_LUT4AB/FrameData[19] Tile_X6Y2_LUT4AB/FrameData[1]
+ Tile_X6Y2_LUT4AB/FrameData[20] Tile_X6Y2_LUT4AB/FrameData[21] Tile_X6Y2_LUT4AB/FrameData[22]
+ Tile_X6Y2_LUT4AB/FrameData[23] Tile_X6Y2_LUT4AB/FrameData[24] Tile_X6Y2_LUT4AB/FrameData[25]
+ Tile_X6Y2_LUT4AB/FrameData[26] Tile_X6Y2_LUT4AB/FrameData[27] Tile_X6Y2_LUT4AB/FrameData[28]
+ Tile_X6Y2_LUT4AB/FrameData[29] Tile_X6Y2_LUT4AB/FrameData[2] Tile_X6Y2_LUT4AB/FrameData[30]
+ Tile_X6Y2_LUT4AB/FrameData[31] Tile_X6Y2_LUT4AB/FrameData[3] Tile_X6Y2_LUT4AB/FrameData[4]
+ Tile_X6Y2_LUT4AB/FrameData[5] Tile_X6Y2_LUT4AB/FrameData[6] Tile_X6Y2_LUT4AB/FrameData[7]
+ Tile_X6Y2_LUT4AB/FrameData[8] Tile_X6Y2_LUT4AB/FrameData[9] Tile_X6Y2_LUT4AB/FrameData_O[0]
+ Tile_X6Y2_LUT4AB/FrameData_O[10] Tile_X6Y2_LUT4AB/FrameData_O[11] Tile_X6Y2_LUT4AB/FrameData_O[12]
+ Tile_X6Y2_LUT4AB/FrameData_O[13] Tile_X6Y2_LUT4AB/FrameData_O[14] Tile_X6Y2_LUT4AB/FrameData_O[15]
+ Tile_X6Y2_LUT4AB/FrameData_O[16] Tile_X6Y2_LUT4AB/FrameData_O[17] Tile_X6Y2_LUT4AB/FrameData_O[18]
+ Tile_X6Y2_LUT4AB/FrameData_O[19] Tile_X6Y2_LUT4AB/FrameData_O[1] Tile_X6Y2_LUT4AB/FrameData_O[20]
+ Tile_X6Y2_LUT4AB/FrameData_O[21] Tile_X6Y2_LUT4AB/FrameData_O[22] Tile_X6Y2_LUT4AB/FrameData_O[23]
+ Tile_X6Y2_LUT4AB/FrameData_O[24] Tile_X6Y2_LUT4AB/FrameData_O[25] Tile_X6Y2_LUT4AB/FrameData_O[26]
+ Tile_X6Y2_LUT4AB/FrameData_O[27] Tile_X6Y2_LUT4AB/FrameData_O[28] Tile_X6Y2_LUT4AB/FrameData_O[29]
+ Tile_X6Y2_LUT4AB/FrameData_O[2] Tile_X6Y2_LUT4AB/FrameData_O[30] Tile_X6Y2_LUT4AB/FrameData_O[31]
+ Tile_X6Y2_LUT4AB/FrameData_O[3] Tile_X6Y2_LUT4AB/FrameData_O[4] Tile_X6Y2_LUT4AB/FrameData_O[5]
+ Tile_X6Y2_LUT4AB/FrameData_O[6] Tile_X6Y2_LUT4AB/FrameData_O[7] Tile_X6Y2_LUT4AB/FrameData_O[8]
+ Tile_X6Y2_LUT4AB/FrameData_O[9] Tile_X6Y2_LUT4AB/FrameStrobe[0] Tile_X6Y2_LUT4AB/FrameStrobe[10]
+ Tile_X6Y2_LUT4AB/FrameStrobe[11] Tile_X6Y2_LUT4AB/FrameStrobe[12] Tile_X6Y2_LUT4AB/FrameStrobe[13]
+ Tile_X6Y2_LUT4AB/FrameStrobe[14] Tile_X6Y2_LUT4AB/FrameStrobe[15] Tile_X6Y2_LUT4AB/FrameStrobe[16]
+ Tile_X6Y2_LUT4AB/FrameStrobe[17] Tile_X6Y2_LUT4AB/FrameStrobe[18] Tile_X6Y2_LUT4AB/FrameStrobe[19]
+ Tile_X6Y2_LUT4AB/FrameStrobe[1] Tile_X6Y2_LUT4AB/FrameStrobe[2] Tile_X6Y2_LUT4AB/FrameStrobe[3]
+ Tile_X6Y2_LUT4AB/FrameStrobe[4] Tile_X6Y2_LUT4AB/FrameStrobe[5] Tile_X6Y2_LUT4AB/FrameStrobe[6]
+ Tile_X6Y2_LUT4AB/FrameStrobe[7] Tile_X6Y2_LUT4AB/FrameStrobe[8] Tile_X6Y2_LUT4AB/FrameStrobe[9]
+ Tile_X6Y1_LUT4AB/FrameStrobe[0] Tile_X6Y1_LUT4AB/FrameStrobe[10] Tile_X6Y1_LUT4AB/FrameStrobe[11]
+ Tile_X6Y1_LUT4AB/FrameStrobe[12] Tile_X6Y1_LUT4AB/FrameStrobe[13] Tile_X6Y1_LUT4AB/FrameStrobe[14]
+ Tile_X6Y1_LUT4AB/FrameStrobe[15] Tile_X6Y1_LUT4AB/FrameStrobe[16] Tile_X6Y1_LUT4AB/FrameStrobe[17]
+ Tile_X6Y1_LUT4AB/FrameStrobe[18] Tile_X6Y1_LUT4AB/FrameStrobe[19] Tile_X6Y1_LUT4AB/FrameStrobe[1]
+ Tile_X6Y1_LUT4AB/FrameStrobe[2] Tile_X6Y1_LUT4AB/FrameStrobe[3] Tile_X6Y1_LUT4AB/FrameStrobe[4]
+ Tile_X6Y1_LUT4AB/FrameStrobe[5] Tile_X6Y1_LUT4AB/FrameStrobe[6] Tile_X6Y1_LUT4AB/FrameStrobe[7]
+ Tile_X6Y1_LUT4AB/FrameStrobe[8] Tile_X6Y1_LUT4AB/FrameStrobe[9] Tile_X6Y2_LUT4AB/N1BEG[0]
+ Tile_X6Y2_LUT4AB/N1BEG[1] Tile_X6Y2_LUT4AB/N1BEG[2] Tile_X6Y2_LUT4AB/N1BEG[3] Tile_X6Y3_LUT4AB/N1BEG[0]
+ Tile_X6Y3_LUT4AB/N1BEG[1] Tile_X6Y3_LUT4AB/N1BEG[2] Tile_X6Y3_LUT4AB/N1BEG[3] Tile_X6Y2_LUT4AB/N2BEG[0]
+ Tile_X6Y2_LUT4AB/N2BEG[1] Tile_X6Y2_LUT4AB/N2BEG[2] Tile_X6Y2_LUT4AB/N2BEG[3] Tile_X6Y2_LUT4AB/N2BEG[4]
+ Tile_X6Y2_LUT4AB/N2BEG[5] Tile_X6Y2_LUT4AB/N2BEG[6] Tile_X6Y2_LUT4AB/N2BEG[7] Tile_X6Y1_LUT4AB/N2END[0]
+ Tile_X6Y1_LUT4AB/N2END[1] Tile_X6Y1_LUT4AB/N2END[2] Tile_X6Y1_LUT4AB/N2END[3] Tile_X6Y1_LUT4AB/N2END[4]
+ Tile_X6Y1_LUT4AB/N2END[5] Tile_X6Y1_LUT4AB/N2END[6] Tile_X6Y1_LUT4AB/N2END[7] Tile_X6Y2_LUT4AB/N2END[0]
+ Tile_X6Y2_LUT4AB/N2END[1] Tile_X6Y2_LUT4AB/N2END[2] Tile_X6Y2_LUT4AB/N2END[3] Tile_X6Y2_LUT4AB/N2END[4]
+ Tile_X6Y2_LUT4AB/N2END[5] Tile_X6Y2_LUT4AB/N2END[6] Tile_X6Y2_LUT4AB/N2END[7] Tile_X6Y3_LUT4AB/N2BEG[0]
+ Tile_X6Y3_LUT4AB/N2BEG[1] Tile_X6Y3_LUT4AB/N2BEG[2] Tile_X6Y3_LUT4AB/N2BEG[3] Tile_X6Y3_LUT4AB/N2BEG[4]
+ Tile_X6Y3_LUT4AB/N2BEG[5] Tile_X6Y3_LUT4AB/N2BEG[6] Tile_X6Y3_LUT4AB/N2BEG[7] Tile_X6Y2_LUT4AB/N4BEG[0]
+ Tile_X6Y2_LUT4AB/N4BEG[10] Tile_X6Y2_LUT4AB/N4BEG[11] Tile_X6Y2_LUT4AB/N4BEG[12]
+ Tile_X6Y2_LUT4AB/N4BEG[13] Tile_X6Y2_LUT4AB/N4BEG[14] Tile_X6Y2_LUT4AB/N4BEG[15]
+ Tile_X6Y2_LUT4AB/N4BEG[1] Tile_X6Y2_LUT4AB/N4BEG[2] Tile_X6Y2_LUT4AB/N4BEG[3] Tile_X6Y2_LUT4AB/N4BEG[4]
+ Tile_X6Y2_LUT4AB/N4BEG[5] Tile_X6Y2_LUT4AB/N4BEG[6] Tile_X6Y2_LUT4AB/N4BEG[7] Tile_X6Y2_LUT4AB/N4BEG[8]
+ Tile_X6Y2_LUT4AB/N4BEG[9] Tile_X6Y3_LUT4AB/N4BEG[0] Tile_X6Y3_LUT4AB/N4BEG[10] Tile_X6Y3_LUT4AB/N4BEG[11]
+ Tile_X6Y3_LUT4AB/N4BEG[12] Tile_X6Y3_LUT4AB/N4BEG[13] Tile_X6Y3_LUT4AB/N4BEG[14]
+ Tile_X6Y3_LUT4AB/N4BEG[15] Tile_X6Y3_LUT4AB/N4BEG[1] Tile_X6Y3_LUT4AB/N4BEG[2] Tile_X6Y3_LUT4AB/N4BEG[3]
+ Tile_X6Y3_LUT4AB/N4BEG[4] Tile_X6Y3_LUT4AB/N4BEG[5] Tile_X6Y3_LUT4AB/N4BEG[6] Tile_X6Y3_LUT4AB/N4BEG[7]
+ Tile_X6Y3_LUT4AB/N4BEG[8] Tile_X6Y3_LUT4AB/N4BEG[9] Tile_X6Y2_LUT4AB/NN4BEG[0] Tile_X6Y2_LUT4AB/NN4BEG[10]
+ Tile_X6Y2_LUT4AB/NN4BEG[11] Tile_X6Y2_LUT4AB/NN4BEG[12] Tile_X6Y2_LUT4AB/NN4BEG[13]
+ Tile_X6Y2_LUT4AB/NN4BEG[14] Tile_X6Y2_LUT4AB/NN4BEG[15] Tile_X6Y2_LUT4AB/NN4BEG[1]
+ Tile_X6Y2_LUT4AB/NN4BEG[2] Tile_X6Y2_LUT4AB/NN4BEG[3] Tile_X6Y2_LUT4AB/NN4BEG[4]
+ Tile_X6Y2_LUT4AB/NN4BEG[5] Tile_X6Y2_LUT4AB/NN4BEG[6] Tile_X6Y2_LUT4AB/NN4BEG[7]
+ Tile_X6Y2_LUT4AB/NN4BEG[8] Tile_X6Y2_LUT4AB/NN4BEG[9] Tile_X6Y3_LUT4AB/NN4BEG[0]
+ Tile_X6Y3_LUT4AB/NN4BEG[10] Tile_X6Y3_LUT4AB/NN4BEG[11] Tile_X6Y3_LUT4AB/NN4BEG[12]
+ Tile_X6Y3_LUT4AB/NN4BEG[13] Tile_X6Y3_LUT4AB/NN4BEG[14] Tile_X6Y3_LUT4AB/NN4BEG[15]
+ Tile_X6Y3_LUT4AB/NN4BEG[1] Tile_X6Y3_LUT4AB/NN4BEG[2] Tile_X6Y3_LUT4AB/NN4BEG[3]
+ Tile_X6Y3_LUT4AB/NN4BEG[4] Tile_X6Y3_LUT4AB/NN4BEG[5] Tile_X6Y3_LUT4AB/NN4BEG[6]
+ Tile_X6Y3_LUT4AB/NN4BEG[7] Tile_X6Y3_LUT4AB/NN4BEG[8] Tile_X6Y3_LUT4AB/NN4BEG[9]
+ Tile_X6Y3_LUT4AB/S1END[0] Tile_X6Y3_LUT4AB/S1END[1] Tile_X6Y3_LUT4AB/S1END[2] Tile_X6Y3_LUT4AB/S1END[3]
+ Tile_X6Y2_LUT4AB/S1END[0] Tile_X6Y2_LUT4AB/S1END[1] Tile_X6Y2_LUT4AB/S1END[2] Tile_X6Y2_LUT4AB/S1END[3]
+ Tile_X6Y3_LUT4AB/S2MID[0] Tile_X6Y3_LUT4AB/S2MID[1] Tile_X6Y3_LUT4AB/S2MID[2] Tile_X6Y3_LUT4AB/S2MID[3]
+ Tile_X6Y3_LUT4AB/S2MID[4] Tile_X6Y3_LUT4AB/S2MID[5] Tile_X6Y3_LUT4AB/S2MID[6] Tile_X6Y3_LUT4AB/S2MID[7]
+ Tile_X6Y3_LUT4AB/S2END[0] Tile_X6Y3_LUT4AB/S2END[1] Tile_X6Y3_LUT4AB/S2END[2] Tile_X6Y3_LUT4AB/S2END[3]
+ Tile_X6Y3_LUT4AB/S2END[4] Tile_X6Y3_LUT4AB/S2END[5] Tile_X6Y3_LUT4AB/S2END[6] Tile_X6Y3_LUT4AB/S2END[7]
+ Tile_X6Y2_LUT4AB/S2END[0] Tile_X6Y2_LUT4AB/S2END[1] Tile_X6Y2_LUT4AB/S2END[2] Tile_X6Y2_LUT4AB/S2END[3]
+ Tile_X6Y2_LUT4AB/S2END[4] Tile_X6Y2_LUT4AB/S2END[5] Tile_X6Y2_LUT4AB/S2END[6] Tile_X6Y2_LUT4AB/S2END[7]
+ Tile_X6Y2_LUT4AB/S2MID[0] Tile_X6Y2_LUT4AB/S2MID[1] Tile_X6Y2_LUT4AB/S2MID[2] Tile_X6Y2_LUT4AB/S2MID[3]
+ Tile_X6Y2_LUT4AB/S2MID[4] Tile_X6Y2_LUT4AB/S2MID[5] Tile_X6Y2_LUT4AB/S2MID[6] Tile_X6Y2_LUT4AB/S2MID[7]
+ Tile_X6Y3_LUT4AB/S4END[0] Tile_X6Y3_LUT4AB/S4END[10] Tile_X6Y3_LUT4AB/S4END[11]
+ Tile_X6Y3_LUT4AB/S4END[12] Tile_X6Y3_LUT4AB/S4END[13] Tile_X6Y3_LUT4AB/S4END[14]
+ Tile_X6Y3_LUT4AB/S4END[15] Tile_X6Y3_LUT4AB/S4END[1] Tile_X6Y3_LUT4AB/S4END[2] Tile_X6Y3_LUT4AB/S4END[3]
+ Tile_X6Y3_LUT4AB/S4END[4] Tile_X6Y3_LUT4AB/S4END[5] Tile_X6Y3_LUT4AB/S4END[6] Tile_X6Y3_LUT4AB/S4END[7]
+ Tile_X6Y3_LUT4AB/S4END[8] Tile_X6Y3_LUT4AB/S4END[9] Tile_X6Y2_LUT4AB/S4END[0] Tile_X6Y2_LUT4AB/S4END[10]
+ Tile_X6Y2_LUT4AB/S4END[11] Tile_X6Y2_LUT4AB/S4END[12] Tile_X6Y2_LUT4AB/S4END[13]
+ Tile_X6Y2_LUT4AB/S4END[14] Tile_X6Y2_LUT4AB/S4END[15] Tile_X6Y2_LUT4AB/S4END[1]
+ Tile_X6Y2_LUT4AB/S4END[2] Tile_X6Y2_LUT4AB/S4END[3] Tile_X6Y2_LUT4AB/S4END[4] Tile_X6Y2_LUT4AB/S4END[5]
+ Tile_X6Y2_LUT4AB/S4END[6] Tile_X6Y2_LUT4AB/S4END[7] Tile_X6Y2_LUT4AB/S4END[8] Tile_X6Y2_LUT4AB/S4END[9]
+ Tile_X6Y3_LUT4AB/SS4END[0] Tile_X6Y3_LUT4AB/SS4END[10] Tile_X6Y3_LUT4AB/SS4END[11]
+ Tile_X6Y3_LUT4AB/SS4END[12] Tile_X6Y3_LUT4AB/SS4END[13] Tile_X6Y3_LUT4AB/SS4END[14]
+ Tile_X6Y3_LUT4AB/SS4END[15] Tile_X6Y3_LUT4AB/SS4END[1] Tile_X6Y3_LUT4AB/SS4END[2]
+ Tile_X6Y3_LUT4AB/SS4END[3] Tile_X6Y3_LUT4AB/SS4END[4] Tile_X6Y3_LUT4AB/SS4END[5]
+ Tile_X6Y3_LUT4AB/SS4END[6] Tile_X6Y3_LUT4AB/SS4END[7] Tile_X6Y3_LUT4AB/SS4END[8]
+ Tile_X6Y3_LUT4AB/SS4END[9] Tile_X6Y2_LUT4AB/SS4END[0] Tile_X6Y2_LUT4AB/SS4END[10]
+ Tile_X6Y2_LUT4AB/SS4END[11] Tile_X6Y2_LUT4AB/SS4END[12] Tile_X6Y2_LUT4AB/SS4END[13]
+ Tile_X6Y2_LUT4AB/SS4END[14] Tile_X6Y2_LUT4AB/SS4END[15] Tile_X6Y2_LUT4AB/SS4END[1]
+ Tile_X6Y2_LUT4AB/SS4END[2] Tile_X6Y2_LUT4AB/SS4END[3] Tile_X6Y2_LUT4AB/SS4END[4]
+ Tile_X6Y2_LUT4AB/SS4END[5] Tile_X6Y2_LUT4AB/SS4END[6] Tile_X6Y2_LUT4AB/SS4END[7]
+ Tile_X6Y2_LUT4AB/SS4END[8] Tile_X6Y2_LUT4AB/SS4END[9] Tile_X6Y2_LUT4AB/UserCLK Tile_X6Y1_LUT4AB/UserCLK
+ VGND VPWR Tile_X6Y2_LUT4AB/W1BEG[0] Tile_X6Y2_LUT4AB/W1BEG[1] Tile_X6Y2_LUT4AB/W1BEG[2]
+ Tile_X6Y2_LUT4AB/W1BEG[3] Tile_X6Y2_LUT4AB/W1END[0] Tile_X6Y2_LUT4AB/W1END[1] Tile_X6Y2_LUT4AB/W1END[2]
+ Tile_X6Y2_LUT4AB/W1END[3] Tile_X6Y2_LUT4AB/W2BEG[0] Tile_X6Y2_LUT4AB/W2BEG[1] Tile_X6Y2_LUT4AB/W2BEG[2]
+ Tile_X6Y2_LUT4AB/W2BEG[3] Tile_X6Y2_LUT4AB/W2BEG[4] Tile_X6Y2_LUT4AB/W2BEG[5] Tile_X6Y2_LUT4AB/W2BEG[6]
+ Tile_X6Y2_LUT4AB/W2BEG[7] Tile_X5Y2_LUT4AB/W2END[0] Tile_X5Y2_LUT4AB/W2END[1] Tile_X5Y2_LUT4AB/W2END[2]
+ Tile_X5Y2_LUT4AB/W2END[3] Tile_X5Y2_LUT4AB/W2END[4] Tile_X5Y2_LUT4AB/W2END[5] Tile_X5Y2_LUT4AB/W2END[6]
+ Tile_X5Y2_LUT4AB/W2END[7] Tile_X6Y2_LUT4AB/W2END[0] Tile_X6Y2_LUT4AB/W2END[1] Tile_X6Y2_LUT4AB/W2END[2]
+ Tile_X6Y2_LUT4AB/W2END[3] Tile_X6Y2_LUT4AB/W2END[4] Tile_X6Y2_LUT4AB/W2END[5] Tile_X6Y2_LUT4AB/W2END[6]
+ Tile_X6Y2_LUT4AB/W2END[7] Tile_X6Y2_LUT4AB/W2MID[0] Tile_X6Y2_LUT4AB/W2MID[1] Tile_X6Y2_LUT4AB/W2MID[2]
+ Tile_X6Y2_LUT4AB/W2MID[3] Tile_X6Y2_LUT4AB/W2MID[4] Tile_X6Y2_LUT4AB/W2MID[5] Tile_X6Y2_LUT4AB/W2MID[6]
+ Tile_X6Y2_LUT4AB/W2MID[7] Tile_X6Y2_LUT4AB/W6BEG[0] Tile_X6Y2_LUT4AB/W6BEG[10] Tile_X6Y2_LUT4AB/W6BEG[11]
+ Tile_X6Y2_LUT4AB/W6BEG[1] Tile_X6Y2_LUT4AB/W6BEG[2] Tile_X6Y2_LUT4AB/W6BEG[3] Tile_X6Y2_LUT4AB/W6BEG[4]
+ Tile_X6Y2_LUT4AB/W6BEG[5] Tile_X6Y2_LUT4AB/W6BEG[6] Tile_X6Y2_LUT4AB/W6BEG[7] Tile_X6Y2_LUT4AB/W6BEG[8]
+ Tile_X6Y2_LUT4AB/W6BEG[9] Tile_X6Y2_LUT4AB/W6END[0] Tile_X6Y2_LUT4AB/W6END[10] Tile_X6Y2_LUT4AB/W6END[11]
+ Tile_X6Y2_LUT4AB/W6END[1] Tile_X6Y2_LUT4AB/W6END[2] Tile_X6Y2_LUT4AB/W6END[3] Tile_X6Y2_LUT4AB/W6END[4]
+ Tile_X6Y2_LUT4AB/W6END[5] Tile_X6Y2_LUT4AB/W6END[6] Tile_X6Y2_LUT4AB/W6END[7] Tile_X6Y2_LUT4AB/W6END[8]
+ Tile_X6Y2_LUT4AB/W6END[9] Tile_X6Y2_LUT4AB/WW4BEG[0] Tile_X6Y2_LUT4AB/WW4BEG[10]
+ Tile_X6Y2_LUT4AB/WW4BEG[11] Tile_X6Y2_LUT4AB/WW4BEG[12] Tile_X6Y2_LUT4AB/WW4BEG[13]
+ Tile_X6Y2_LUT4AB/WW4BEG[14] Tile_X6Y2_LUT4AB/WW4BEG[15] Tile_X6Y2_LUT4AB/WW4BEG[1]
+ Tile_X6Y2_LUT4AB/WW4BEG[2] Tile_X6Y2_LUT4AB/WW4BEG[3] Tile_X6Y2_LUT4AB/WW4BEG[4]
+ Tile_X6Y2_LUT4AB/WW4BEG[5] Tile_X6Y2_LUT4AB/WW4BEG[6] Tile_X6Y2_LUT4AB/WW4BEG[7]
+ Tile_X6Y2_LUT4AB/WW4BEG[8] Tile_X6Y2_LUT4AB/WW4BEG[9] Tile_X6Y2_LUT4AB/WW4END[0]
+ Tile_X6Y2_LUT4AB/WW4END[10] Tile_X6Y2_LUT4AB/WW4END[11] Tile_X6Y2_LUT4AB/WW4END[12]
+ Tile_X6Y2_LUT4AB/WW4END[13] Tile_X6Y2_LUT4AB/WW4END[14] Tile_X6Y2_LUT4AB/WW4END[15]
+ Tile_X6Y2_LUT4AB/WW4END[1] Tile_X6Y2_LUT4AB/WW4END[2] Tile_X6Y2_LUT4AB/WW4END[3]
+ Tile_X6Y2_LUT4AB/WW4END[4] Tile_X6Y2_LUT4AB/WW4END[5] Tile_X6Y2_LUT4AB/WW4END[6]
+ Tile_X6Y2_LUT4AB/WW4END[7] Tile_X6Y2_LUT4AB/WW4END[8] Tile_X6Y2_LUT4AB/WW4END[9]
+ LUT4AB
XTile_X9Y7_LUT4AB Tile_X9Y8_LUT4AB/Co Tile_X9Y7_LUT4AB/Co Tile_X9Y7_LUT4AB/E1BEG[0]
+ Tile_X9Y7_LUT4AB/E1BEG[1] Tile_X9Y7_LUT4AB/E1BEG[2] Tile_X9Y7_LUT4AB/E1BEG[3] Tile_X9Y7_LUT4AB/E1END[0]
+ Tile_X9Y7_LUT4AB/E1END[1] Tile_X9Y7_LUT4AB/E1END[2] Tile_X9Y7_LUT4AB/E1END[3] Tile_X9Y7_LUT4AB/E2BEG[0]
+ Tile_X9Y7_LUT4AB/E2BEG[1] Tile_X9Y7_LUT4AB/E2BEG[2] Tile_X9Y7_LUT4AB/E2BEG[3] Tile_X9Y7_LUT4AB/E2BEG[4]
+ Tile_X9Y7_LUT4AB/E2BEG[5] Tile_X9Y7_LUT4AB/E2BEG[6] Tile_X9Y7_LUT4AB/E2BEG[7] Tile_X9Y7_LUT4AB/E2BEGb[0]
+ Tile_X9Y7_LUT4AB/E2BEGb[1] Tile_X9Y7_LUT4AB/E2BEGb[2] Tile_X9Y7_LUT4AB/E2BEGb[3]
+ Tile_X9Y7_LUT4AB/E2BEGb[4] Tile_X9Y7_LUT4AB/E2BEGb[5] Tile_X9Y7_LUT4AB/E2BEGb[6]
+ Tile_X9Y7_LUT4AB/E2BEGb[7] Tile_X9Y7_LUT4AB/E2END[0] Tile_X9Y7_LUT4AB/E2END[1] Tile_X9Y7_LUT4AB/E2END[2]
+ Tile_X9Y7_LUT4AB/E2END[3] Tile_X9Y7_LUT4AB/E2END[4] Tile_X9Y7_LUT4AB/E2END[5] Tile_X9Y7_LUT4AB/E2END[6]
+ Tile_X9Y7_LUT4AB/E2END[7] Tile_X9Y7_LUT4AB/E2MID[0] Tile_X9Y7_LUT4AB/E2MID[1] Tile_X9Y7_LUT4AB/E2MID[2]
+ Tile_X9Y7_LUT4AB/E2MID[3] Tile_X9Y7_LUT4AB/E2MID[4] Tile_X9Y7_LUT4AB/E2MID[5] Tile_X9Y7_LUT4AB/E2MID[6]
+ Tile_X9Y7_LUT4AB/E2MID[7] Tile_X9Y7_LUT4AB/E6BEG[0] Tile_X9Y7_LUT4AB/E6BEG[10] Tile_X9Y7_LUT4AB/E6BEG[11]
+ Tile_X9Y7_LUT4AB/E6BEG[1] Tile_X9Y7_LUT4AB/E6BEG[2] Tile_X9Y7_LUT4AB/E6BEG[3] Tile_X9Y7_LUT4AB/E6BEG[4]
+ Tile_X9Y7_LUT4AB/E6BEG[5] Tile_X9Y7_LUT4AB/E6BEG[6] Tile_X9Y7_LUT4AB/E6BEG[7] Tile_X9Y7_LUT4AB/E6BEG[8]
+ Tile_X9Y7_LUT4AB/E6BEG[9] Tile_X9Y7_LUT4AB/E6END[0] Tile_X9Y7_LUT4AB/E6END[10] Tile_X9Y7_LUT4AB/E6END[11]
+ Tile_X9Y7_LUT4AB/E6END[1] Tile_X9Y7_LUT4AB/E6END[2] Tile_X9Y7_LUT4AB/E6END[3] Tile_X9Y7_LUT4AB/E6END[4]
+ Tile_X9Y7_LUT4AB/E6END[5] Tile_X9Y7_LUT4AB/E6END[6] Tile_X9Y7_LUT4AB/E6END[7] Tile_X9Y7_LUT4AB/E6END[8]
+ Tile_X9Y7_LUT4AB/E6END[9] Tile_X9Y7_LUT4AB/EE4BEG[0] Tile_X9Y7_LUT4AB/EE4BEG[10]
+ Tile_X9Y7_LUT4AB/EE4BEG[11] Tile_X9Y7_LUT4AB/EE4BEG[12] Tile_X9Y7_LUT4AB/EE4BEG[13]
+ Tile_X9Y7_LUT4AB/EE4BEG[14] Tile_X9Y7_LUT4AB/EE4BEG[15] Tile_X9Y7_LUT4AB/EE4BEG[1]
+ Tile_X9Y7_LUT4AB/EE4BEG[2] Tile_X9Y7_LUT4AB/EE4BEG[3] Tile_X9Y7_LUT4AB/EE4BEG[4]
+ Tile_X9Y7_LUT4AB/EE4BEG[5] Tile_X9Y7_LUT4AB/EE4BEG[6] Tile_X9Y7_LUT4AB/EE4BEG[7]
+ Tile_X9Y7_LUT4AB/EE4BEG[8] Tile_X9Y7_LUT4AB/EE4BEG[9] Tile_X9Y7_LUT4AB/EE4END[0]
+ Tile_X9Y7_LUT4AB/EE4END[10] Tile_X9Y7_LUT4AB/EE4END[11] Tile_X9Y7_LUT4AB/EE4END[12]
+ Tile_X9Y7_LUT4AB/EE4END[13] Tile_X9Y7_LUT4AB/EE4END[14] Tile_X9Y7_LUT4AB/EE4END[15]
+ Tile_X9Y7_LUT4AB/EE4END[1] Tile_X9Y7_LUT4AB/EE4END[2] Tile_X9Y7_LUT4AB/EE4END[3]
+ Tile_X9Y7_LUT4AB/EE4END[4] Tile_X9Y7_LUT4AB/EE4END[5] Tile_X9Y7_LUT4AB/EE4END[6]
+ Tile_X9Y7_LUT4AB/EE4END[7] Tile_X9Y7_LUT4AB/EE4END[8] Tile_X9Y7_LUT4AB/EE4END[9]
+ Tile_X9Y7_LUT4AB/FrameData[0] Tile_X9Y7_LUT4AB/FrameData[10] Tile_X9Y7_LUT4AB/FrameData[11]
+ Tile_X9Y7_LUT4AB/FrameData[12] Tile_X9Y7_LUT4AB/FrameData[13] Tile_X9Y7_LUT4AB/FrameData[14]
+ Tile_X9Y7_LUT4AB/FrameData[15] Tile_X9Y7_LUT4AB/FrameData[16] Tile_X9Y7_LUT4AB/FrameData[17]
+ Tile_X9Y7_LUT4AB/FrameData[18] Tile_X9Y7_LUT4AB/FrameData[19] Tile_X9Y7_LUT4AB/FrameData[1]
+ Tile_X9Y7_LUT4AB/FrameData[20] Tile_X9Y7_LUT4AB/FrameData[21] Tile_X9Y7_LUT4AB/FrameData[22]
+ Tile_X9Y7_LUT4AB/FrameData[23] Tile_X9Y7_LUT4AB/FrameData[24] Tile_X9Y7_LUT4AB/FrameData[25]
+ Tile_X9Y7_LUT4AB/FrameData[26] Tile_X9Y7_LUT4AB/FrameData[27] Tile_X9Y7_LUT4AB/FrameData[28]
+ Tile_X9Y7_LUT4AB/FrameData[29] Tile_X9Y7_LUT4AB/FrameData[2] Tile_X9Y7_LUT4AB/FrameData[30]
+ Tile_X9Y7_LUT4AB/FrameData[31] Tile_X9Y7_LUT4AB/FrameData[3] Tile_X9Y7_LUT4AB/FrameData[4]
+ Tile_X9Y7_LUT4AB/FrameData[5] Tile_X9Y7_LUT4AB/FrameData[6] Tile_X9Y7_LUT4AB/FrameData[7]
+ Tile_X9Y7_LUT4AB/FrameData[8] Tile_X9Y7_LUT4AB/FrameData[9] Tile_X9Y7_LUT4AB/FrameData_O[0]
+ Tile_X9Y7_LUT4AB/FrameData_O[10] Tile_X9Y7_LUT4AB/FrameData_O[11] Tile_X9Y7_LUT4AB/FrameData_O[12]
+ Tile_X9Y7_LUT4AB/FrameData_O[13] Tile_X9Y7_LUT4AB/FrameData_O[14] Tile_X9Y7_LUT4AB/FrameData_O[15]
+ Tile_X9Y7_LUT4AB/FrameData_O[16] Tile_X9Y7_LUT4AB/FrameData_O[17] Tile_X9Y7_LUT4AB/FrameData_O[18]
+ Tile_X9Y7_LUT4AB/FrameData_O[19] Tile_X9Y7_LUT4AB/FrameData_O[1] Tile_X9Y7_LUT4AB/FrameData_O[20]
+ Tile_X9Y7_LUT4AB/FrameData_O[21] Tile_X9Y7_LUT4AB/FrameData_O[22] Tile_X9Y7_LUT4AB/FrameData_O[23]
+ Tile_X9Y7_LUT4AB/FrameData_O[24] Tile_X9Y7_LUT4AB/FrameData_O[25] Tile_X9Y7_LUT4AB/FrameData_O[26]
+ Tile_X9Y7_LUT4AB/FrameData_O[27] Tile_X9Y7_LUT4AB/FrameData_O[28] Tile_X9Y7_LUT4AB/FrameData_O[29]
+ Tile_X9Y7_LUT4AB/FrameData_O[2] Tile_X9Y7_LUT4AB/FrameData_O[30] Tile_X9Y7_LUT4AB/FrameData_O[31]
+ Tile_X9Y7_LUT4AB/FrameData_O[3] Tile_X9Y7_LUT4AB/FrameData_O[4] Tile_X9Y7_LUT4AB/FrameData_O[5]
+ Tile_X9Y7_LUT4AB/FrameData_O[6] Tile_X9Y7_LUT4AB/FrameData_O[7] Tile_X9Y7_LUT4AB/FrameData_O[8]
+ Tile_X9Y7_LUT4AB/FrameData_O[9] Tile_X9Y7_LUT4AB/FrameStrobe[0] Tile_X9Y7_LUT4AB/FrameStrobe[10]
+ Tile_X9Y7_LUT4AB/FrameStrobe[11] Tile_X9Y7_LUT4AB/FrameStrobe[12] Tile_X9Y7_LUT4AB/FrameStrobe[13]
+ Tile_X9Y7_LUT4AB/FrameStrobe[14] Tile_X9Y7_LUT4AB/FrameStrobe[15] Tile_X9Y7_LUT4AB/FrameStrobe[16]
+ Tile_X9Y7_LUT4AB/FrameStrobe[17] Tile_X9Y7_LUT4AB/FrameStrobe[18] Tile_X9Y7_LUT4AB/FrameStrobe[19]
+ Tile_X9Y7_LUT4AB/FrameStrobe[1] Tile_X9Y7_LUT4AB/FrameStrobe[2] Tile_X9Y7_LUT4AB/FrameStrobe[3]
+ Tile_X9Y7_LUT4AB/FrameStrobe[4] Tile_X9Y7_LUT4AB/FrameStrobe[5] Tile_X9Y7_LUT4AB/FrameStrobe[6]
+ Tile_X9Y7_LUT4AB/FrameStrobe[7] Tile_X9Y7_LUT4AB/FrameStrobe[8] Tile_X9Y7_LUT4AB/FrameStrobe[9]
+ Tile_X9Y6_LUT4AB/FrameStrobe[0] Tile_X9Y6_LUT4AB/FrameStrobe[10] Tile_X9Y6_LUT4AB/FrameStrobe[11]
+ Tile_X9Y6_LUT4AB/FrameStrobe[12] Tile_X9Y6_LUT4AB/FrameStrobe[13] Tile_X9Y6_LUT4AB/FrameStrobe[14]
+ Tile_X9Y6_LUT4AB/FrameStrobe[15] Tile_X9Y6_LUT4AB/FrameStrobe[16] Tile_X9Y6_LUT4AB/FrameStrobe[17]
+ Tile_X9Y6_LUT4AB/FrameStrobe[18] Tile_X9Y6_LUT4AB/FrameStrobe[19] Tile_X9Y6_LUT4AB/FrameStrobe[1]
+ Tile_X9Y6_LUT4AB/FrameStrobe[2] Tile_X9Y6_LUT4AB/FrameStrobe[3] Tile_X9Y6_LUT4AB/FrameStrobe[4]
+ Tile_X9Y6_LUT4AB/FrameStrobe[5] Tile_X9Y6_LUT4AB/FrameStrobe[6] Tile_X9Y6_LUT4AB/FrameStrobe[7]
+ Tile_X9Y6_LUT4AB/FrameStrobe[8] Tile_X9Y6_LUT4AB/FrameStrobe[9] Tile_X9Y7_LUT4AB/N1BEG[0]
+ Tile_X9Y7_LUT4AB/N1BEG[1] Tile_X9Y7_LUT4AB/N1BEG[2] Tile_X9Y7_LUT4AB/N1BEG[3] Tile_X9Y8_LUT4AB/N1BEG[0]
+ Tile_X9Y8_LUT4AB/N1BEG[1] Tile_X9Y8_LUT4AB/N1BEG[2] Tile_X9Y8_LUT4AB/N1BEG[3] Tile_X9Y7_LUT4AB/N2BEG[0]
+ Tile_X9Y7_LUT4AB/N2BEG[1] Tile_X9Y7_LUT4AB/N2BEG[2] Tile_X9Y7_LUT4AB/N2BEG[3] Tile_X9Y7_LUT4AB/N2BEG[4]
+ Tile_X9Y7_LUT4AB/N2BEG[5] Tile_X9Y7_LUT4AB/N2BEG[6] Tile_X9Y7_LUT4AB/N2BEG[7] Tile_X9Y6_LUT4AB/N2END[0]
+ Tile_X9Y6_LUT4AB/N2END[1] Tile_X9Y6_LUT4AB/N2END[2] Tile_X9Y6_LUT4AB/N2END[3] Tile_X9Y6_LUT4AB/N2END[4]
+ Tile_X9Y6_LUT4AB/N2END[5] Tile_X9Y6_LUT4AB/N2END[6] Tile_X9Y6_LUT4AB/N2END[7] Tile_X9Y7_LUT4AB/N2END[0]
+ Tile_X9Y7_LUT4AB/N2END[1] Tile_X9Y7_LUT4AB/N2END[2] Tile_X9Y7_LUT4AB/N2END[3] Tile_X9Y7_LUT4AB/N2END[4]
+ Tile_X9Y7_LUT4AB/N2END[5] Tile_X9Y7_LUT4AB/N2END[6] Tile_X9Y7_LUT4AB/N2END[7] Tile_X9Y8_LUT4AB/N2BEG[0]
+ Tile_X9Y8_LUT4AB/N2BEG[1] Tile_X9Y8_LUT4AB/N2BEG[2] Tile_X9Y8_LUT4AB/N2BEG[3] Tile_X9Y8_LUT4AB/N2BEG[4]
+ Tile_X9Y8_LUT4AB/N2BEG[5] Tile_X9Y8_LUT4AB/N2BEG[6] Tile_X9Y8_LUT4AB/N2BEG[7] Tile_X9Y7_LUT4AB/N4BEG[0]
+ Tile_X9Y7_LUT4AB/N4BEG[10] Tile_X9Y7_LUT4AB/N4BEG[11] Tile_X9Y7_LUT4AB/N4BEG[12]
+ Tile_X9Y7_LUT4AB/N4BEG[13] Tile_X9Y7_LUT4AB/N4BEG[14] Tile_X9Y7_LUT4AB/N4BEG[15]
+ Tile_X9Y7_LUT4AB/N4BEG[1] Tile_X9Y7_LUT4AB/N4BEG[2] Tile_X9Y7_LUT4AB/N4BEG[3] Tile_X9Y7_LUT4AB/N4BEG[4]
+ Tile_X9Y7_LUT4AB/N4BEG[5] Tile_X9Y7_LUT4AB/N4BEG[6] Tile_X9Y7_LUT4AB/N4BEG[7] Tile_X9Y7_LUT4AB/N4BEG[8]
+ Tile_X9Y7_LUT4AB/N4BEG[9] Tile_X9Y8_LUT4AB/N4BEG[0] Tile_X9Y8_LUT4AB/N4BEG[10] Tile_X9Y8_LUT4AB/N4BEG[11]
+ Tile_X9Y8_LUT4AB/N4BEG[12] Tile_X9Y8_LUT4AB/N4BEG[13] Tile_X9Y8_LUT4AB/N4BEG[14]
+ Tile_X9Y8_LUT4AB/N4BEG[15] Tile_X9Y8_LUT4AB/N4BEG[1] Tile_X9Y8_LUT4AB/N4BEG[2] Tile_X9Y8_LUT4AB/N4BEG[3]
+ Tile_X9Y8_LUT4AB/N4BEG[4] Tile_X9Y8_LUT4AB/N4BEG[5] Tile_X9Y8_LUT4AB/N4BEG[6] Tile_X9Y8_LUT4AB/N4BEG[7]
+ Tile_X9Y8_LUT4AB/N4BEG[8] Tile_X9Y8_LUT4AB/N4BEG[9] Tile_X9Y7_LUT4AB/NN4BEG[0] Tile_X9Y7_LUT4AB/NN4BEG[10]
+ Tile_X9Y7_LUT4AB/NN4BEG[11] Tile_X9Y7_LUT4AB/NN4BEG[12] Tile_X9Y7_LUT4AB/NN4BEG[13]
+ Tile_X9Y7_LUT4AB/NN4BEG[14] Tile_X9Y7_LUT4AB/NN4BEG[15] Tile_X9Y7_LUT4AB/NN4BEG[1]
+ Tile_X9Y7_LUT4AB/NN4BEG[2] Tile_X9Y7_LUT4AB/NN4BEG[3] Tile_X9Y7_LUT4AB/NN4BEG[4]
+ Tile_X9Y7_LUT4AB/NN4BEG[5] Tile_X9Y7_LUT4AB/NN4BEG[6] Tile_X9Y7_LUT4AB/NN4BEG[7]
+ Tile_X9Y7_LUT4AB/NN4BEG[8] Tile_X9Y7_LUT4AB/NN4BEG[9] Tile_X9Y8_LUT4AB/NN4BEG[0]
+ Tile_X9Y8_LUT4AB/NN4BEG[10] Tile_X9Y8_LUT4AB/NN4BEG[11] Tile_X9Y8_LUT4AB/NN4BEG[12]
+ Tile_X9Y8_LUT4AB/NN4BEG[13] Tile_X9Y8_LUT4AB/NN4BEG[14] Tile_X9Y8_LUT4AB/NN4BEG[15]
+ Tile_X9Y8_LUT4AB/NN4BEG[1] Tile_X9Y8_LUT4AB/NN4BEG[2] Tile_X9Y8_LUT4AB/NN4BEG[3]
+ Tile_X9Y8_LUT4AB/NN4BEG[4] Tile_X9Y8_LUT4AB/NN4BEG[5] Tile_X9Y8_LUT4AB/NN4BEG[6]
+ Tile_X9Y8_LUT4AB/NN4BEG[7] Tile_X9Y8_LUT4AB/NN4BEG[8] Tile_X9Y8_LUT4AB/NN4BEG[9]
+ Tile_X9Y8_LUT4AB/S1END[0] Tile_X9Y8_LUT4AB/S1END[1] Tile_X9Y8_LUT4AB/S1END[2] Tile_X9Y8_LUT4AB/S1END[3]
+ Tile_X9Y7_LUT4AB/S1END[0] Tile_X9Y7_LUT4AB/S1END[1] Tile_X9Y7_LUT4AB/S1END[2] Tile_X9Y7_LUT4AB/S1END[3]
+ Tile_X9Y8_LUT4AB/S2MID[0] Tile_X9Y8_LUT4AB/S2MID[1] Tile_X9Y8_LUT4AB/S2MID[2] Tile_X9Y8_LUT4AB/S2MID[3]
+ Tile_X9Y8_LUT4AB/S2MID[4] Tile_X9Y8_LUT4AB/S2MID[5] Tile_X9Y8_LUT4AB/S2MID[6] Tile_X9Y8_LUT4AB/S2MID[7]
+ Tile_X9Y8_LUT4AB/S2END[0] Tile_X9Y8_LUT4AB/S2END[1] Tile_X9Y8_LUT4AB/S2END[2] Tile_X9Y8_LUT4AB/S2END[3]
+ Tile_X9Y8_LUT4AB/S2END[4] Tile_X9Y8_LUT4AB/S2END[5] Tile_X9Y8_LUT4AB/S2END[6] Tile_X9Y8_LUT4AB/S2END[7]
+ Tile_X9Y7_LUT4AB/S2END[0] Tile_X9Y7_LUT4AB/S2END[1] Tile_X9Y7_LUT4AB/S2END[2] Tile_X9Y7_LUT4AB/S2END[3]
+ Tile_X9Y7_LUT4AB/S2END[4] Tile_X9Y7_LUT4AB/S2END[5] Tile_X9Y7_LUT4AB/S2END[6] Tile_X9Y7_LUT4AB/S2END[7]
+ Tile_X9Y7_LUT4AB/S2MID[0] Tile_X9Y7_LUT4AB/S2MID[1] Tile_X9Y7_LUT4AB/S2MID[2] Tile_X9Y7_LUT4AB/S2MID[3]
+ Tile_X9Y7_LUT4AB/S2MID[4] Tile_X9Y7_LUT4AB/S2MID[5] Tile_X9Y7_LUT4AB/S2MID[6] Tile_X9Y7_LUT4AB/S2MID[7]
+ Tile_X9Y8_LUT4AB/S4END[0] Tile_X9Y8_LUT4AB/S4END[10] Tile_X9Y8_LUT4AB/S4END[11]
+ Tile_X9Y8_LUT4AB/S4END[12] Tile_X9Y8_LUT4AB/S4END[13] Tile_X9Y8_LUT4AB/S4END[14]
+ Tile_X9Y8_LUT4AB/S4END[15] Tile_X9Y8_LUT4AB/S4END[1] Tile_X9Y8_LUT4AB/S4END[2] Tile_X9Y8_LUT4AB/S4END[3]
+ Tile_X9Y8_LUT4AB/S4END[4] Tile_X9Y8_LUT4AB/S4END[5] Tile_X9Y8_LUT4AB/S4END[6] Tile_X9Y8_LUT4AB/S4END[7]
+ Tile_X9Y8_LUT4AB/S4END[8] Tile_X9Y8_LUT4AB/S4END[9] Tile_X9Y7_LUT4AB/S4END[0] Tile_X9Y7_LUT4AB/S4END[10]
+ Tile_X9Y7_LUT4AB/S4END[11] Tile_X9Y7_LUT4AB/S4END[12] Tile_X9Y7_LUT4AB/S4END[13]
+ Tile_X9Y7_LUT4AB/S4END[14] Tile_X9Y7_LUT4AB/S4END[15] Tile_X9Y7_LUT4AB/S4END[1]
+ Tile_X9Y7_LUT4AB/S4END[2] Tile_X9Y7_LUT4AB/S4END[3] Tile_X9Y7_LUT4AB/S4END[4] Tile_X9Y7_LUT4AB/S4END[5]
+ Tile_X9Y7_LUT4AB/S4END[6] Tile_X9Y7_LUT4AB/S4END[7] Tile_X9Y7_LUT4AB/S4END[8] Tile_X9Y7_LUT4AB/S4END[9]
+ Tile_X9Y8_LUT4AB/SS4END[0] Tile_X9Y8_LUT4AB/SS4END[10] Tile_X9Y8_LUT4AB/SS4END[11]
+ Tile_X9Y8_LUT4AB/SS4END[12] Tile_X9Y8_LUT4AB/SS4END[13] Tile_X9Y8_LUT4AB/SS4END[14]
+ Tile_X9Y8_LUT4AB/SS4END[15] Tile_X9Y8_LUT4AB/SS4END[1] Tile_X9Y8_LUT4AB/SS4END[2]
+ Tile_X9Y8_LUT4AB/SS4END[3] Tile_X9Y8_LUT4AB/SS4END[4] Tile_X9Y8_LUT4AB/SS4END[5]
+ Tile_X9Y8_LUT4AB/SS4END[6] Tile_X9Y8_LUT4AB/SS4END[7] Tile_X9Y8_LUT4AB/SS4END[8]
+ Tile_X9Y8_LUT4AB/SS4END[9] Tile_X9Y7_LUT4AB/SS4END[0] Tile_X9Y7_LUT4AB/SS4END[10]
+ Tile_X9Y7_LUT4AB/SS4END[11] Tile_X9Y7_LUT4AB/SS4END[12] Tile_X9Y7_LUT4AB/SS4END[13]
+ Tile_X9Y7_LUT4AB/SS4END[14] Tile_X9Y7_LUT4AB/SS4END[15] Tile_X9Y7_LUT4AB/SS4END[1]
+ Tile_X9Y7_LUT4AB/SS4END[2] Tile_X9Y7_LUT4AB/SS4END[3] Tile_X9Y7_LUT4AB/SS4END[4]
+ Tile_X9Y7_LUT4AB/SS4END[5] Tile_X9Y7_LUT4AB/SS4END[6] Tile_X9Y7_LUT4AB/SS4END[7]
+ Tile_X9Y7_LUT4AB/SS4END[8] Tile_X9Y7_LUT4AB/SS4END[9] Tile_X9Y7_LUT4AB/UserCLK Tile_X9Y6_LUT4AB/UserCLK
+ VGND VPWR Tile_X9Y7_LUT4AB/W1BEG[0] Tile_X9Y7_LUT4AB/W1BEG[1] Tile_X9Y7_LUT4AB/W1BEG[2]
+ Tile_X9Y7_LUT4AB/W1BEG[3] Tile_X9Y7_LUT4AB/W1END[0] Tile_X9Y7_LUT4AB/W1END[1] Tile_X9Y7_LUT4AB/W1END[2]
+ Tile_X9Y7_LUT4AB/W1END[3] Tile_X9Y7_LUT4AB/W2BEG[0] Tile_X9Y7_LUT4AB/W2BEG[1] Tile_X9Y7_LUT4AB/W2BEG[2]
+ Tile_X9Y7_LUT4AB/W2BEG[3] Tile_X9Y7_LUT4AB/W2BEG[4] Tile_X9Y7_LUT4AB/W2BEG[5] Tile_X9Y7_LUT4AB/W2BEG[6]
+ Tile_X9Y7_LUT4AB/W2BEG[7] Tile_X8Y7_LUT4AB/W2END[0] Tile_X8Y7_LUT4AB/W2END[1] Tile_X8Y7_LUT4AB/W2END[2]
+ Tile_X8Y7_LUT4AB/W2END[3] Tile_X8Y7_LUT4AB/W2END[4] Tile_X8Y7_LUT4AB/W2END[5] Tile_X8Y7_LUT4AB/W2END[6]
+ Tile_X8Y7_LUT4AB/W2END[7] Tile_X9Y7_LUT4AB/W2END[0] Tile_X9Y7_LUT4AB/W2END[1] Tile_X9Y7_LUT4AB/W2END[2]
+ Tile_X9Y7_LUT4AB/W2END[3] Tile_X9Y7_LUT4AB/W2END[4] Tile_X9Y7_LUT4AB/W2END[5] Tile_X9Y7_LUT4AB/W2END[6]
+ Tile_X9Y7_LUT4AB/W2END[7] Tile_X9Y7_LUT4AB/W2MID[0] Tile_X9Y7_LUT4AB/W2MID[1] Tile_X9Y7_LUT4AB/W2MID[2]
+ Tile_X9Y7_LUT4AB/W2MID[3] Tile_X9Y7_LUT4AB/W2MID[4] Tile_X9Y7_LUT4AB/W2MID[5] Tile_X9Y7_LUT4AB/W2MID[6]
+ Tile_X9Y7_LUT4AB/W2MID[7] Tile_X9Y7_LUT4AB/W6BEG[0] Tile_X9Y7_LUT4AB/W6BEG[10] Tile_X9Y7_LUT4AB/W6BEG[11]
+ Tile_X9Y7_LUT4AB/W6BEG[1] Tile_X9Y7_LUT4AB/W6BEG[2] Tile_X9Y7_LUT4AB/W6BEG[3] Tile_X9Y7_LUT4AB/W6BEG[4]
+ Tile_X9Y7_LUT4AB/W6BEG[5] Tile_X9Y7_LUT4AB/W6BEG[6] Tile_X9Y7_LUT4AB/W6BEG[7] Tile_X9Y7_LUT4AB/W6BEG[8]
+ Tile_X9Y7_LUT4AB/W6BEG[9] Tile_X9Y7_LUT4AB/W6END[0] Tile_X9Y7_LUT4AB/W6END[10] Tile_X9Y7_LUT4AB/W6END[11]
+ Tile_X9Y7_LUT4AB/W6END[1] Tile_X9Y7_LUT4AB/W6END[2] Tile_X9Y7_LUT4AB/W6END[3] Tile_X9Y7_LUT4AB/W6END[4]
+ Tile_X9Y7_LUT4AB/W6END[5] Tile_X9Y7_LUT4AB/W6END[6] Tile_X9Y7_LUT4AB/W6END[7] Tile_X9Y7_LUT4AB/W6END[8]
+ Tile_X9Y7_LUT4AB/W6END[9] Tile_X9Y7_LUT4AB/WW4BEG[0] Tile_X9Y7_LUT4AB/WW4BEG[10]
+ Tile_X9Y7_LUT4AB/WW4BEG[11] Tile_X9Y7_LUT4AB/WW4BEG[12] Tile_X9Y7_LUT4AB/WW4BEG[13]
+ Tile_X9Y7_LUT4AB/WW4BEG[14] Tile_X9Y7_LUT4AB/WW4BEG[15] Tile_X9Y7_LUT4AB/WW4BEG[1]
+ Tile_X9Y7_LUT4AB/WW4BEG[2] Tile_X9Y7_LUT4AB/WW4BEG[3] Tile_X9Y7_LUT4AB/WW4BEG[4]
+ Tile_X9Y7_LUT4AB/WW4BEG[5] Tile_X9Y7_LUT4AB/WW4BEG[6] Tile_X9Y7_LUT4AB/WW4BEG[7]
+ Tile_X9Y7_LUT4AB/WW4BEG[8] Tile_X9Y7_LUT4AB/WW4BEG[9] Tile_X9Y7_LUT4AB/WW4END[0]
+ Tile_X9Y7_LUT4AB/WW4END[10] Tile_X9Y7_LUT4AB/WW4END[11] Tile_X9Y7_LUT4AB/WW4END[12]
+ Tile_X9Y7_LUT4AB/WW4END[13] Tile_X9Y7_LUT4AB/WW4END[14] Tile_X9Y7_LUT4AB/WW4END[15]
+ Tile_X9Y7_LUT4AB/WW4END[1] Tile_X9Y7_LUT4AB/WW4END[2] Tile_X9Y7_LUT4AB/WW4END[3]
+ Tile_X9Y7_LUT4AB/WW4END[4] Tile_X9Y7_LUT4AB/WW4END[5] Tile_X9Y7_LUT4AB/WW4END[6]
+ Tile_X9Y7_LUT4AB/WW4END[7] Tile_X9Y7_LUT4AB/WW4END[8] Tile_X9Y7_LUT4AB/WW4END[9]
+ LUT4AB
XTile_X2Y14_LUT4AB Tile_X2Y14_LUT4AB/Ci Tile_X2Y14_LUT4AB/Co Tile_X3Y14_LUT4AB/E1END[0]
+ Tile_X3Y14_LUT4AB/E1END[1] Tile_X3Y14_LUT4AB/E1END[2] Tile_X3Y14_LUT4AB/E1END[3]
+ Tile_X2Y14_LUT4AB/E1END[0] Tile_X2Y14_LUT4AB/E1END[1] Tile_X2Y14_LUT4AB/E1END[2]
+ Tile_X2Y14_LUT4AB/E1END[3] Tile_X3Y14_LUT4AB/E2MID[0] Tile_X3Y14_LUT4AB/E2MID[1]
+ Tile_X3Y14_LUT4AB/E2MID[2] Tile_X3Y14_LUT4AB/E2MID[3] Tile_X3Y14_LUT4AB/E2MID[4]
+ Tile_X3Y14_LUT4AB/E2MID[5] Tile_X3Y14_LUT4AB/E2MID[6] Tile_X3Y14_LUT4AB/E2MID[7]
+ Tile_X3Y14_LUT4AB/E2END[0] Tile_X3Y14_LUT4AB/E2END[1] Tile_X3Y14_LUT4AB/E2END[2]
+ Tile_X3Y14_LUT4AB/E2END[3] Tile_X3Y14_LUT4AB/E2END[4] Tile_X3Y14_LUT4AB/E2END[5]
+ Tile_X3Y14_LUT4AB/E2END[6] Tile_X3Y14_LUT4AB/E2END[7] Tile_X2Y14_LUT4AB/E2END[0]
+ Tile_X2Y14_LUT4AB/E2END[1] Tile_X2Y14_LUT4AB/E2END[2] Tile_X2Y14_LUT4AB/E2END[3]
+ Tile_X2Y14_LUT4AB/E2END[4] Tile_X2Y14_LUT4AB/E2END[5] Tile_X2Y14_LUT4AB/E2END[6]
+ Tile_X2Y14_LUT4AB/E2END[7] Tile_X2Y14_LUT4AB/E2MID[0] Tile_X2Y14_LUT4AB/E2MID[1]
+ Tile_X2Y14_LUT4AB/E2MID[2] Tile_X2Y14_LUT4AB/E2MID[3] Tile_X2Y14_LUT4AB/E2MID[4]
+ Tile_X2Y14_LUT4AB/E2MID[5] Tile_X2Y14_LUT4AB/E2MID[6] Tile_X2Y14_LUT4AB/E2MID[7]
+ Tile_X3Y14_LUT4AB/E6END[0] Tile_X3Y14_LUT4AB/E6END[10] Tile_X3Y14_LUT4AB/E6END[11]
+ Tile_X3Y14_LUT4AB/E6END[1] Tile_X3Y14_LUT4AB/E6END[2] Tile_X3Y14_LUT4AB/E6END[3]
+ Tile_X3Y14_LUT4AB/E6END[4] Tile_X3Y14_LUT4AB/E6END[5] Tile_X3Y14_LUT4AB/E6END[6]
+ Tile_X3Y14_LUT4AB/E6END[7] Tile_X3Y14_LUT4AB/E6END[8] Tile_X3Y14_LUT4AB/E6END[9]
+ Tile_X2Y14_LUT4AB/E6END[0] Tile_X2Y14_LUT4AB/E6END[10] Tile_X2Y14_LUT4AB/E6END[11]
+ Tile_X2Y14_LUT4AB/E6END[1] Tile_X2Y14_LUT4AB/E6END[2] Tile_X2Y14_LUT4AB/E6END[3]
+ Tile_X2Y14_LUT4AB/E6END[4] Tile_X2Y14_LUT4AB/E6END[5] Tile_X2Y14_LUT4AB/E6END[6]
+ Tile_X2Y14_LUT4AB/E6END[7] Tile_X2Y14_LUT4AB/E6END[8] Tile_X2Y14_LUT4AB/E6END[9]
+ Tile_X3Y14_LUT4AB/EE4END[0] Tile_X3Y14_LUT4AB/EE4END[10] Tile_X3Y14_LUT4AB/EE4END[11]
+ Tile_X3Y14_LUT4AB/EE4END[12] Tile_X3Y14_LUT4AB/EE4END[13] Tile_X3Y14_LUT4AB/EE4END[14]
+ Tile_X3Y14_LUT4AB/EE4END[15] Tile_X3Y14_LUT4AB/EE4END[1] Tile_X3Y14_LUT4AB/EE4END[2]
+ Tile_X3Y14_LUT4AB/EE4END[3] Tile_X3Y14_LUT4AB/EE4END[4] Tile_X3Y14_LUT4AB/EE4END[5]
+ Tile_X3Y14_LUT4AB/EE4END[6] Tile_X3Y14_LUT4AB/EE4END[7] Tile_X3Y14_LUT4AB/EE4END[8]
+ Tile_X3Y14_LUT4AB/EE4END[9] Tile_X2Y14_LUT4AB/EE4END[0] Tile_X2Y14_LUT4AB/EE4END[10]
+ Tile_X2Y14_LUT4AB/EE4END[11] Tile_X2Y14_LUT4AB/EE4END[12] Tile_X2Y14_LUT4AB/EE4END[13]
+ Tile_X2Y14_LUT4AB/EE4END[14] Tile_X2Y14_LUT4AB/EE4END[15] Tile_X2Y14_LUT4AB/EE4END[1]
+ Tile_X2Y14_LUT4AB/EE4END[2] Tile_X2Y14_LUT4AB/EE4END[3] Tile_X2Y14_LUT4AB/EE4END[4]
+ Tile_X2Y14_LUT4AB/EE4END[5] Tile_X2Y14_LUT4AB/EE4END[6] Tile_X2Y14_LUT4AB/EE4END[7]
+ Tile_X2Y14_LUT4AB/EE4END[8] Tile_X2Y14_LUT4AB/EE4END[9] Tile_X2Y14_LUT4AB/FrameData[0]
+ Tile_X2Y14_LUT4AB/FrameData[10] Tile_X2Y14_LUT4AB/FrameData[11] Tile_X2Y14_LUT4AB/FrameData[12]
+ Tile_X2Y14_LUT4AB/FrameData[13] Tile_X2Y14_LUT4AB/FrameData[14] Tile_X2Y14_LUT4AB/FrameData[15]
+ Tile_X2Y14_LUT4AB/FrameData[16] Tile_X2Y14_LUT4AB/FrameData[17] Tile_X2Y14_LUT4AB/FrameData[18]
+ Tile_X2Y14_LUT4AB/FrameData[19] Tile_X2Y14_LUT4AB/FrameData[1] Tile_X2Y14_LUT4AB/FrameData[20]
+ Tile_X2Y14_LUT4AB/FrameData[21] Tile_X2Y14_LUT4AB/FrameData[22] Tile_X2Y14_LUT4AB/FrameData[23]
+ Tile_X2Y14_LUT4AB/FrameData[24] Tile_X2Y14_LUT4AB/FrameData[25] Tile_X2Y14_LUT4AB/FrameData[26]
+ Tile_X2Y14_LUT4AB/FrameData[27] Tile_X2Y14_LUT4AB/FrameData[28] Tile_X2Y14_LUT4AB/FrameData[29]
+ Tile_X2Y14_LUT4AB/FrameData[2] Tile_X2Y14_LUT4AB/FrameData[30] Tile_X2Y14_LUT4AB/FrameData[31]
+ Tile_X2Y14_LUT4AB/FrameData[3] Tile_X2Y14_LUT4AB/FrameData[4] Tile_X2Y14_LUT4AB/FrameData[5]
+ Tile_X2Y14_LUT4AB/FrameData[6] Tile_X2Y14_LUT4AB/FrameData[7] Tile_X2Y14_LUT4AB/FrameData[8]
+ Tile_X2Y14_LUT4AB/FrameData[9] Tile_X3Y14_LUT4AB/FrameData[0] Tile_X3Y14_LUT4AB/FrameData[10]
+ Tile_X3Y14_LUT4AB/FrameData[11] Tile_X3Y14_LUT4AB/FrameData[12] Tile_X3Y14_LUT4AB/FrameData[13]
+ Tile_X3Y14_LUT4AB/FrameData[14] Tile_X3Y14_LUT4AB/FrameData[15] Tile_X3Y14_LUT4AB/FrameData[16]
+ Tile_X3Y14_LUT4AB/FrameData[17] Tile_X3Y14_LUT4AB/FrameData[18] Tile_X3Y14_LUT4AB/FrameData[19]
+ Tile_X3Y14_LUT4AB/FrameData[1] Tile_X3Y14_LUT4AB/FrameData[20] Tile_X3Y14_LUT4AB/FrameData[21]
+ Tile_X3Y14_LUT4AB/FrameData[22] Tile_X3Y14_LUT4AB/FrameData[23] Tile_X3Y14_LUT4AB/FrameData[24]
+ Tile_X3Y14_LUT4AB/FrameData[25] Tile_X3Y14_LUT4AB/FrameData[26] Tile_X3Y14_LUT4AB/FrameData[27]
+ Tile_X3Y14_LUT4AB/FrameData[28] Tile_X3Y14_LUT4AB/FrameData[29] Tile_X3Y14_LUT4AB/FrameData[2]
+ Tile_X3Y14_LUT4AB/FrameData[30] Tile_X3Y14_LUT4AB/FrameData[31] Tile_X3Y14_LUT4AB/FrameData[3]
+ Tile_X3Y14_LUT4AB/FrameData[4] Tile_X3Y14_LUT4AB/FrameData[5] Tile_X3Y14_LUT4AB/FrameData[6]
+ Tile_X3Y14_LUT4AB/FrameData[7] Tile_X3Y14_LUT4AB/FrameData[8] Tile_X3Y14_LUT4AB/FrameData[9]
+ Tile_X2Y14_LUT4AB/FrameStrobe[0] Tile_X2Y14_LUT4AB/FrameStrobe[10] Tile_X2Y14_LUT4AB/FrameStrobe[11]
+ Tile_X2Y14_LUT4AB/FrameStrobe[12] Tile_X2Y14_LUT4AB/FrameStrobe[13] Tile_X2Y14_LUT4AB/FrameStrobe[14]
+ Tile_X2Y14_LUT4AB/FrameStrobe[15] Tile_X2Y14_LUT4AB/FrameStrobe[16] Tile_X2Y14_LUT4AB/FrameStrobe[17]
+ Tile_X2Y14_LUT4AB/FrameStrobe[18] Tile_X2Y14_LUT4AB/FrameStrobe[19] Tile_X2Y14_LUT4AB/FrameStrobe[1]
+ Tile_X2Y14_LUT4AB/FrameStrobe[2] Tile_X2Y14_LUT4AB/FrameStrobe[3] Tile_X2Y14_LUT4AB/FrameStrobe[4]
+ Tile_X2Y14_LUT4AB/FrameStrobe[5] Tile_X2Y14_LUT4AB/FrameStrobe[6] Tile_X2Y14_LUT4AB/FrameStrobe[7]
+ Tile_X2Y14_LUT4AB/FrameStrobe[8] Tile_X2Y14_LUT4AB/FrameStrobe[9] Tile_X2Y13_LUT4AB/FrameStrobe[0]
+ Tile_X2Y13_LUT4AB/FrameStrobe[10] Tile_X2Y13_LUT4AB/FrameStrobe[11] Tile_X2Y13_LUT4AB/FrameStrobe[12]
+ Tile_X2Y13_LUT4AB/FrameStrobe[13] Tile_X2Y13_LUT4AB/FrameStrobe[14] Tile_X2Y13_LUT4AB/FrameStrobe[15]
+ Tile_X2Y13_LUT4AB/FrameStrobe[16] Tile_X2Y13_LUT4AB/FrameStrobe[17] Tile_X2Y13_LUT4AB/FrameStrobe[18]
+ Tile_X2Y13_LUT4AB/FrameStrobe[19] Tile_X2Y13_LUT4AB/FrameStrobe[1] Tile_X2Y13_LUT4AB/FrameStrobe[2]
+ Tile_X2Y13_LUT4AB/FrameStrobe[3] Tile_X2Y13_LUT4AB/FrameStrobe[4] Tile_X2Y13_LUT4AB/FrameStrobe[5]
+ Tile_X2Y13_LUT4AB/FrameStrobe[6] Tile_X2Y13_LUT4AB/FrameStrobe[7] Tile_X2Y13_LUT4AB/FrameStrobe[8]
+ Tile_X2Y13_LUT4AB/FrameStrobe[9] Tile_X2Y14_LUT4AB/N1BEG[0] Tile_X2Y14_LUT4AB/N1BEG[1]
+ Tile_X2Y14_LUT4AB/N1BEG[2] Tile_X2Y14_LUT4AB/N1BEG[3] Tile_X2Y14_LUT4AB/N1END[0]
+ Tile_X2Y14_LUT4AB/N1END[1] Tile_X2Y14_LUT4AB/N1END[2] Tile_X2Y14_LUT4AB/N1END[3]
+ Tile_X2Y14_LUT4AB/N2BEG[0] Tile_X2Y14_LUT4AB/N2BEG[1] Tile_X2Y14_LUT4AB/N2BEG[2]
+ Tile_X2Y14_LUT4AB/N2BEG[3] Tile_X2Y14_LUT4AB/N2BEG[4] Tile_X2Y14_LUT4AB/N2BEG[5]
+ Tile_X2Y14_LUT4AB/N2BEG[6] Tile_X2Y14_LUT4AB/N2BEG[7] Tile_X2Y13_LUT4AB/N2END[0]
+ Tile_X2Y13_LUT4AB/N2END[1] Tile_X2Y13_LUT4AB/N2END[2] Tile_X2Y13_LUT4AB/N2END[3]
+ Tile_X2Y13_LUT4AB/N2END[4] Tile_X2Y13_LUT4AB/N2END[5] Tile_X2Y13_LUT4AB/N2END[6]
+ Tile_X2Y13_LUT4AB/N2END[7] Tile_X2Y14_LUT4AB/N2END[0] Tile_X2Y14_LUT4AB/N2END[1]
+ Tile_X2Y14_LUT4AB/N2END[2] Tile_X2Y14_LUT4AB/N2END[3] Tile_X2Y14_LUT4AB/N2END[4]
+ Tile_X2Y14_LUT4AB/N2END[5] Tile_X2Y14_LUT4AB/N2END[6] Tile_X2Y14_LUT4AB/N2END[7]
+ Tile_X2Y14_LUT4AB/N2MID[0] Tile_X2Y14_LUT4AB/N2MID[1] Tile_X2Y14_LUT4AB/N2MID[2]
+ Tile_X2Y14_LUT4AB/N2MID[3] Tile_X2Y14_LUT4AB/N2MID[4] Tile_X2Y14_LUT4AB/N2MID[5]
+ Tile_X2Y14_LUT4AB/N2MID[6] Tile_X2Y14_LUT4AB/N2MID[7] Tile_X2Y14_LUT4AB/N4BEG[0]
+ Tile_X2Y14_LUT4AB/N4BEG[10] Tile_X2Y14_LUT4AB/N4BEG[11] Tile_X2Y14_LUT4AB/N4BEG[12]
+ Tile_X2Y14_LUT4AB/N4BEG[13] Tile_X2Y14_LUT4AB/N4BEG[14] Tile_X2Y14_LUT4AB/N4BEG[15]
+ Tile_X2Y14_LUT4AB/N4BEG[1] Tile_X2Y14_LUT4AB/N4BEG[2] Tile_X2Y14_LUT4AB/N4BEG[3]
+ Tile_X2Y14_LUT4AB/N4BEG[4] Tile_X2Y14_LUT4AB/N4BEG[5] Tile_X2Y14_LUT4AB/N4BEG[6]
+ Tile_X2Y14_LUT4AB/N4BEG[7] Tile_X2Y14_LUT4AB/N4BEG[8] Tile_X2Y14_LUT4AB/N4BEG[9]
+ Tile_X2Y14_LUT4AB/N4END[0] Tile_X2Y14_LUT4AB/N4END[10] Tile_X2Y14_LUT4AB/N4END[11]
+ Tile_X2Y14_LUT4AB/N4END[12] Tile_X2Y14_LUT4AB/N4END[13] Tile_X2Y14_LUT4AB/N4END[14]
+ Tile_X2Y14_LUT4AB/N4END[15] Tile_X2Y14_LUT4AB/N4END[1] Tile_X2Y14_LUT4AB/N4END[2]
+ Tile_X2Y14_LUT4AB/N4END[3] Tile_X2Y14_LUT4AB/N4END[4] Tile_X2Y14_LUT4AB/N4END[5]
+ Tile_X2Y14_LUT4AB/N4END[6] Tile_X2Y14_LUT4AB/N4END[7] Tile_X2Y14_LUT4AB/N4END[8]
+ Tile_X2Y14_LUT4AB/N4END[9] Tile_X2Y14_LUT4AB/NN4BEG[0] Tile_X2Y14_LUT4AB/NN4BEG[10]
+ Tile_X2Y14_LUT4AB/NN4BEG[11] Tile_X2Y14_LUT4AB/NN4BEG[12] Tile_X2Y14_LUT4AB/NN4BEG[13]
+ Tile_X2Y14_LUT4AB/NN4BEG[14] Tile_X2Y14_LUT4AB/NN4BEG[15] Tile_X2Y14_LUT4AB/NN4BEG[1]
+ Tile_X2Y14_LUT4AB/NN4BEG[2] Tile_X2Y14_LUT4AB/NN4BEG[3] Tile_X2Y14_LUT4AB/NN4BEG[4]
+ Tile_X2Y14_LUT4AB/NN4BEG[5] Tile_X2Y14_LUT4AB/NN4BEG[6] Tile_X2Y14_LUT4AB/NN4BEG[7]
+ Tile_X2Y14_LUT4AB/NN4BEG[8] Tile_X2Y14_LUT4AB/NN4BEG[9] Tile_X2Y14_LUT4AB/NN4END[0]
+ Tile_X2Y14_LUT4AB/NN4END[10] Tile_X2Y14_LUT4AB/NN4END[11] Tile_X2Y14_LUT4AB/NN4END[12]
+ Tile_X2Y14_LUT4AB/NN4END[13] Tile_X2Y14_LUT4AB/NN4END[14] Tile_X2Y14_LUT4AB/NN4END[15]
+ Tile_X2Y14_LUT4AB/NN4END[1] Tile_X2Y14_LUT4AB/NN4END[2] Tile_X2Y14_LUT4AB/NN4END[3]
+ Tile_X2Y14_LUT4AB/NN4END[4] Tile_X2Y14_LUT4AB/NN4END[5] Tile_X2Y14_LUT4AB/NN4END[6]
+ Tile_X2Y14_LUT4AB/NN4END[7] Tile_X2Y14_LUT4AB/NN4END[8] Tile_X2Y14_LUT4AB/NN4END[9]
+ Tile_X2Y14_LUT4AB/S1BEG[0] Tile_X2Y14_LUT4AB/S1BEG[1] Tile_X2Y14_LUT4AB/S1BEG[2]
+ Tile_X2Y14_LUT4AB/S1BEG[3] Tile_X2Y14_LUT4AB/S1END[0] Tile_X2Y14_LUT4AB/S1END[1]
+ Tile_X2Y14_LUT4AB/S1END[2] Tile_X2Y14_LUT4AB/S1END[3] Tile_X2Y14_LUT4AB/S2BEG[0]
+ Tile_X2Y14_LUT4AB/S2BEG[1] Tile_X2Y14_LUT4AB/S2BEG[2] Tile_X2Y14_LUT4AB/S2BEG[3]
+ Tile_X2Y14_LUT4AB/S2BEG[4] Tile_X2Y14_LUT4AB/S2BEG[5] Tile_X2Y14_LUT4AB/S2BEG[6]
+ Tile_X2Y14_LUT4AB/S2BEG[7] Tile_X2Y14_LUT4AB/S2BEGb[0] Tile_X2Y14_LUT4AB/S2BEGb[1]
+ Tile_X2Y14_LUT4AB/S2BEGb[2] Tile_X2Y14_LUT4AB/S2BEGb[3] Tile_X2Y14_LUT4AB/S2BEGb[4]
+ Tile_X2Y14_LUT4AB/S2BEGb[5] Tile_X2Y14_LUT4AB/S2BEGb[6] Tile_X2Y14_LUT4AB/S2BEGb[7]
+ Tile_X2Y14_LUT4AB/S2END[0] Tile_X2Y14_LUT4AB/S2END[1] Tile_X2Y14_LUT4AB/S2END[2]
+ Tile_X2Y14_LUT4AB/S2END[3] Tile_X2Y14_LUT4AB/S2END[4] Tile_X2Y14_LUT4AB/S2END[5]
+ Tile_X2Y14_LUT4AB/S2END[6] Tile_X2Y14_LUT4AB/S2END[7] Tile_X2Y14_LUT4AB/S2MID[0]
+ Tile_X2Y14_LUT4AB/S2MID[1] Tile_X2Y14_LUT4AB/S2MID[2] Tile_X2Y14_LUT4AB/S2MID[3]
+ Tile_X2Y14_LUT4AB/S2MID[4] Tile_X2Y14_LUT4AB/S2MID[5] Tile_X2Y14_LUT4AB/S2MID[6]
+ Tile_X2Y14_LUT4AB/S2MID[7] Tile_X2Y14_LUT4AB/S4BEG[0] Tile_X2Y14_LUT4AB/S4BEG[10]
+ Tile_X2Y14_LUT4AB/S4BEG[11] Tile_X2Y14_LUT4AB/S4BEG[12] Tile_X2Y14_LUT4AB/S4BEG[13]
+ Tile_X2Y14_LUT4AB/S4BEG[14] Tile_X2Y14_LUT4AB/S4BEG[15] Tile_X2Y14_LUT4AB/S4BEG[1]
+ Tile_X2Y14_LUT4AB/S4BEG[2] Tile_X2Y14_LUT4AB/S4BEG[3] Tile_X2Y14_LUT4AB/S4BEG[4]
+ Tile_X2Y14_LUT4AB/S4BEG[5] Tile_X2Y14_LUT4AB/S4BEG[6] Tile_X2Y14_LUT4AB/S4BEG[7]
+ Tile_X2Y14_LUT4AB/S4BEG[8] Tile_X2Y14_LUT4AB/S4BEG[9] Tile_X2Y14_LUT4AB/S4END[0]
+ Tile_X2Y14_LUT4AB/S4END[10] Tile_X2Y14_LUT4AB/S4END[11] Tile_X2Y14_LUT4AB/S4END[12]
+ Tile_X2Y14_LUT4AB/S4END[13] Tile_X2Y14_LUT4AB/S4END[14] Tile_X2Y14_LUT4AB/S4END[15]
+ Tile_X2Y14_LUT4AB/S4END[1] Tile_X2Y14_LUT4AB/S4END[2] Tile_X2Y14_LUT4AB/S4END[3]
+ Tile_X2Y14_LUT4AB/S4END[4] Tile_X2Y14_LUT4AB/S4END[5] Tile_X2Y14_LUT4AB/S4END[6]
+ Tile_X2Y14_LUT4AB/S4END[7] Tile_X2Y14_LUT4AB/S4END[8] Tile_X2Y14_LUT4AB/S4END[9]
+ Tile_X2Y14_LUT4AB/SS4BEG[0] Tile_X2Y14_LUT4AB/SS4BEG[10] Tile_X2Y14_LUT4AB/SS4BEG[11]
+ Tile_X2Y14_LUT4AB/SS4BEG[12] Tile_X2Y14_LUT4AB/SS4BEG[13] Tile_X2Y14_LUT4AB/SS4BEG[14]
+ Tile_X2Y14_LUT4AB/SS4BEG[15] Tile_X2Y14_LUT4AB/SS4BEG[1] Tile_X2Y14_LUT4AB/SS4BEG[2]
+ Tile_X2Y14_LUT4AB/SS4BEG[3] Tile_X2Y14_LUT4AB/SS4BEG[4] Tile_X2Y14_LUT4AB/SS4BEG[5]
+ Tile_X2Y14_LUT4AB/SS4BEG[6] Tile_X2Y14_LUT4AB/SS4BEG[7] Tile_X2Y14_LUT4AB/SS4BEG[8]
+ Tile_X2Y14_LUT4AB/SS4BEG[9] Tile_X2Y14_LUT4AB/SS4END[0] Tile_X2Y14_LUT4AB/SS4END[10]
+ Tile_X2Y14_LUT4AB/SS4END[11] Tile_X2Y14_LUT4AB/SS4END[12] Tile_X2Y14_LUT4AB/SS4END[13]
+ Tile_X2Y14_LUT4AB/SS4END[14] Tile_X2Y14_LUT4AB/SS4END[15] Tile_X2Y14_LUT4AB/SS4END[1]
+ Tile_X2Y14_LUT4AB/SS4END[2] Tile_X2Y14_LUT4AB/SS4END[3] Tile_X2Y14_LUT4AB/SS4END[4]
+ Tile_X2Y14_LUT4AB/SS4END[5] Tile_X2Y14_LUT4AB/SS4END[6] Tile_X2Y14_LUT4AB/SS4END[7]
+ Tile_X2Y14_LUT4AB/SS4END[8] Tile_X2Y14_LUT4AB/SS4END[9] Tile_X2Y14_LUT4AB/UserCLK
+ Tile_X2Y13_LUT4AB/UserCLK VGND VPWR Tile_X2Y14_LUT4AB/W1BEG[0] Tile_X2Y14_LUT4AB/W1BEG[1]
+ Tile_X2Y14_LUT4AB/W1BEG[2] Tile_X2Y14_LUT4AB/W1BEG[3] Tile_X3Y14_LUT4AB/W1BEG[0]
+ Tile_X3Y14_LUT4AB/W1BEG[1] Tile_X3Y14_LUT4AB/W1BEG[2] Tile_X3Y14_LUT4AB/W1BEG[3]
+ Tile_X2Y14_LUT4AB/W2BEG[0] Tile_X2Y14_LUT4AB/W2BEG[1] Tile_X2Y14_LUT4AB/W2BEG[2]
+ Tile_X2Y14_LUT4AB/W2BEG[3] Tile_X2Y14_LUT4AB/W2BEG[4] Tile_X2Y14_LUT4AB/W2BEG[5]
+ Tile_X2Y14_LUT4AB/W2BEG[6] Tile_X2Y14_LUT4AB/W2BEG[7] Tile_X1Y14_LUT4AB/W2END[0]
+ Tile_X1Y14_LUT4AB/W2END[1] Tile_X1Y14_LUT4AB/W2END[2] Tile_X1Y14_LUT4AB/W2END[3]
+ Tile_X1Y14_LUT4AB/W2END[4] Tile_X1Y14_LUT4AB/W2END[5] Tile_X1Y14_LUT4AB/W2END[6]
+ Tile_X1Y14_LUT4AB/W2END[7] Tile_X2Y14_LUT4AB/W2END[0] Tile_X2Y14_LUT4AB/W2END[1]
+ Tile_X2Y14_LUT4AB/W2END[2] Tile_X2Y14_LUT4AB/W2END[3] Tile_X2Y14_LUT4AB/W2END[4]
+ Tile_X2Y14_LUT4AB/W2END[5] Tile_X2Y14_LUT4AB/W2END[6] Tile_X2Y14_LUT4AB/W2END[7]
+ Tile_X3Y14_LUT4AB/W2BEG[0] Tile_X3Y14_LUT4AB/W2BEG[1] Tile_X3Y14_LUT4AB/W2BEG[2]
+ Tile_X3Y14_LUT4AB/W2BEG[3] Tile_X3Y14_LUT4AB/W2BEG[4] Tile_X3Y14_LUT4AB/W2BEG[5]
+ Tile_X3Y14_LUT4AB/W2BEG[6] Tile_X3Y14_LUT4AB/W2BEG[7] Tile_X2Y14_LUT4AB/W6BEG[0]
+ Tile_X2Y14_LUT4AB/W6BEG[10] Tile_X2Y14_LUT4AB/W6BEG[11] Tile_X2Y14_LUT4AB/W6BEG[1]
+ Tile_X2Y14_LUT4AB/W6BEG[2] Tile_X2Y14_LUT4AB/W6BEG[3] Tile_X2Y14_LUT4AB/W6BEG[4]
+ Tile_X2Y14_LUT4AB/W6BEG[5] Tile_X2Y14_LUT4AB/W6BEG[6] Tile_X2Y14_LUT4AB/W6BEG[7]
+ Tile_X2Y14_LUT4AB/W6BEG[8] Tile_X2Y14_LUT4AB/W6BEG[9] Tile_X3Y14_LUT4AB/W6BEG[0]
+ Tile_X3Y14_LUT4AB/W6BEG[10] Tile_X3Y14_LUT4AB/W6BEG[11] Tile_X3Y14_LUT4AB/W6BEG[1]
+ Tile_X3Y14_LUT4AB/W6BEG[2] Tile_X3Y14_LUT4AB/W6BEG[3] Tile_X3Y14_LUT4AB/W6BEG[4]
+ Tile_X3Y14_LUT4AB/W6BEG[5] Tile_X3Y14_LUT4AB/W6BEG[6] Tile_X3Y14_LUT4AB/W6BEG[7]
+ Tile_X3Y14_LUT4AB/W6BEG[8] Tile_X3Y14_LUT4AB/W6BEG[9] Tile_X2Y14_LUT4AB/WW4BEG[0]
+ Tile_X2Y14_LUT4AB/WW4BEG[10] Tile_X2Y14_LUT4AB/WW4BEG[11] Tile_X2Y14_LUT4AB/WW4BEG[12]
+ Tile_X2Y14_LUT4AB/WW4BEG[13] Tile_X2Y14_LUT4AB/WW4BEG[14] Tile_X2Y14_LUT4AB/WW4BEG[15]
+ Tile_X2Y14_LUT4AB/WW4BEG[1] Tile_X2Y14_LUT4AB/WW4BEG[2] Tile_X2Y14_LUT4AB/WW4BEG[3]
+ Tile_X2Y14_LUT4AB/WW4BEG[4] Tile_X2Y14_LUT4AB/WW4BEG[5] Tile_X2Y14_LUT4AB/WW4BEG[6]
+ Tile_X2Y14_LUT4AB/WW4BEG[7] Tile_X2Y14_LUT4AB/WW4BEG[8] Tile_X2Y14_LUT4AB/WW4BEG[9]
+ Tile_X3Y14_LUT4AB/WW4BEG[0] Tile_X3Y14_LUT4AB/WW4BEG[10] Tile_X3Y14_LUT4AB/WW4BEG[11]
+ Tile_X3Y14_LUT4AB/WW4BEG[12] Tile_X3Y14_LUT4AB/WW4BEG[13] Tile_X3Y14_LUT4AB/WW4BEG[14]
+ Tile_X3Y14_LUT4AB/WW4BEG[15] Tile_X3Y14_LUT4AB/WW4BEG[1] Tile_X3Y14_LUT4AB/WW4BEG[2]
+ Tile_X3Y14_LUT4AB/WW4BEG[3] Tile_X3Y14_LUT4AB/WW4BEG[4] Tile_X3Y14_LUT4AB/WW4BEG[5]
+ Tile_X3Y14_LUT4AB/WW4BEG[6] Tile_X3Y14_LUT4AB/WW4BEG[7] Tile_X3Y14_LUT4AB/WW4BEG[8]
+ Tile_X3Y14_LUT4AB/WW4BEG[9] LUT4AB
XTile_X5Y6_LUT4AB Tile_X5Y7_LUT4AB/Co Tile_X5Y6_LUT4AB/Co Tile_X6Y6_LUT4AB/E1END[0]
+ Tile_X6Y6_LUT4AB/E1END[1] Tile_X6Y6_LUT4AB/E1END[2] Tile_X6Y6_LUT4AB/E1END[3] Tile_X5Y6_LUT4AB/E1END[0]
+ Tile_X5Y6_LUT4AB/E1END[1] Tile_X5Y6_LUT4AB/E1END[2] Tile_X5Y6_LUT4AB/E1END[3] Tile_X6Y6_LUT4AB/E2MID[0]
+ Tile_X6Y6_LUT4AB/E2MID[1] Tile_X6Y6_LUT4AB/E2MID[2] Tile_X6Y6_LUT4AB/E2MID[3] Tile_X6Y6_LUT4AB/E2MID[4]
+ Tile_X6Y6_LUT4AB/E2MID[5] Tile_X6Y6_LUT4AB/E2MID[6] Tile_X6Y6_LUT4AB/E2MID[7] Tile_X6Y6_LUT4AB/E2END[0]
+ Tile_X6Y6_LUT4AB/E2END[1] Tile_X6Y6_LUT4AB/E2END[2] Tile_X6Y6_LUT4AB/E2END[3] Tile_X6Y6_LUT4AB/E2END[4]
+ Tile_X6Y6_LUT4AB/E2END[5] Tile_X6Y6_LUT4AB/E2END[6] Tile_X6Y6_LUT4AB/E2END[7] Tile_X5Y6_LUT4AB/E2END[0]
+ Tile_X5Y6_LUT4AB/E2END[1] Tile_X5Y6_LUT4AB/E2END[2] Tile_X5Y6_LUT4AB/E2END[3] Tile_X5Y6_LUT4AB/E2END[4]
+ Tile_X5Y6_LUT4AB/E2END[5] Tile_X5Y6_LUT4AB/E2END[6] Tile_X5Y6_LUT4AB/E2END[7] Tile_X5Y6_LUT4AB/E2MID[0]
+ Tile_X5Y6_LUT4AB/E2MID[1] Tile_X5Y6_LUT4AB/E2MID[2] Tile_X5Y6_LUT4AB/E2MID[3] Tile_X5Y6_LUT4AB/E2MID[4]
+ Tile_X5Y6_LUT4AB/E2MID[5] Tile_X5Y6_LUT4AB/E2MID[6] Tile_X5Y6_LUT4AB/E2MID[7] Tile_X6Y6_LUT4AB/E6END[0]
+ Tile_X6Y6_LUT4AB/E6END[10] Tile_X6Y6_LUT4AB/E6END[11] Tile_X6Y6_LUT4AB/E6END[1]
+ Tile_X6Y6_LUT4AB/E6END[2] Tile_X6Y6_LUT4AB/E6END[3] Tile_X6Y6_LUT4AB/E6END[4] Tile_X6Y6_LUT4AB/E6END[5]
+ Tile_X6Y6_LUT4AB/E6END[6] Tile_X6Y6_LUT4AB/E6END[7] Tile_X6Y6_LUT4AB/E6END[8] Tile_X6Y6_LUT4AB/E6END[9]
+ Tile_X5Y6_LUT4AB/E6END[0] Tile_X5Y6_LUT4AB/E6END[10] Tile_X5Y6_LUT4AB/E6END[11]
+ Tile_X5Y6_LUT4AB/E6END[1] Tile_X5Y6_LUT4AB/E6END[2] Tile_X5Y6_LUT4AB/E6END[3] Tile_X5Y6_LUT4AB/E6END[4]
+ Tile_X5Y6_LUT4AB/E6END[5] Tile_X5Y6_LUT4AB/E6END[6] Tile_X5Y6_LUT4AB/E6END[7] Tile_X5Y6_LUT4AB/E6END[8]
+ Tile_X5Y6_LUT4AB/E6END[9] Tile_X6Y6_LUT4AB/EE4END[0] Tile_X6Y6_LUT4AB/EE4END[10]
+ Tile_X6Y6_LUT4AB/EE4END[11] Tile_X6Y6_LUT4AB/EE4END[12] Tile_X6Y6_LUT4AB/EE4END[13]
+ Tile_X6Y6_LUT4AB/EE4END[14] Tile_X6Y6_LUT4AB/EE4END[15] Tile_X6Y6_LUT4AB/EE4END[1]
+ Tile_X6Y6_LUT4AB/EE4END[2] Tile_X6Y6_LUT4AB/EE4END[3] Tile_X6Y6_LUT4AB/EE4END[4]
+ Tile_X6Y6_LUT4AB/EE4END[5] Tile_X6Y6_LUT4AB/EE4END[6] Tile_X6Y6_LUT4AB/EE4END[7]
+ Tile_X6Y6_LUT4AB/EE4END[8] Tile_X6Y6_LUT4AB/EE4END[9] Tile_X5Y6_LUT4AB/EE4END[0]
+ Tile_X5Y6_LUT4AB/EE4END[10] Tile_X5Y6_LUT4AB/EE4END[11] Tile_X5Y6_LUT4AB/EE4END[12]
+ Tile_X5Y6_LUT4AB/EE4END[13] Tile_X5Y6_LUT4AB/EE4END[14] Tile_X5Y6_LUT4AB/EE4END[15]
+ Tile_X5Y6_LUT4AB/EE4END[1] Tile_X5Y6_LUT4AB/EE4END[2] Tile_X5Y6_LUT4AB/EE4END[3]
+ Tile_X5Y6_LUT4AB/EE4END[4] Tile_X5Y6_LUT4AB/EE4END[5] Tile_X5Y6_LUT4AB/EE4END[6]
+ Tile_X5Y6_LUT4AB/EE4END[7] Tile_X5Y6_LUT4AB/EE4END[8] Tile_X5Y6_LUT4AB/EE4END[9]
+ Tile_X5Y6_LUT4AB/FrameData[0] Tile_X5Y6_LUT4AB/FrameData[10] Tile_X5Y6_LUT4AB/FrameData[11]
+ Tile_X5Y6_LUT4AB/FrameData[12] Tile_X5Y6_LUT4AB/FrameData[13] Tile_X5Y6_LUT4AB/FrameData[14]
+ Tile_X5Y6_LUT4AB/FrameData[15] Tile_X5Y6_LUT4AB/FrameData[16] Tile_X5Y6_LUT4AB/FrameData[17]
+ Tile_X5Y6_LUT4AB/FrameData[18] Tile_X5Y6_LUT4AB/FrameData[19] Tile_X5Y6_LUT4AB/FrameData[1]
+ Tile_X5Y6_LUT4AB/FrameData[20] Tile_X5Y6_LUT4AB/FrameData[21] Tile_X5Y6_LUT4AB/FrameData[22]
+ Tile_X5Y6_LUT4AB/FrameData[23] Tile_X5Y6_LUT4AB/FrameData[24] Tile_X5Y6_LUT4AB/FrameData[25]
+ Tile_X5Y6_LUT4AB/FrameData[26] Tile_X5Y6_LUT4AB/FrameData[27] Tile_X5Y6_LUT4AB/FrameData[28]
+ Tile_X5Y6_LUT4AB/FrameData[29] Tile_X5Y6_LUT4AB/FrameData[2] Tile_X5Y6_LUT4AB/FrameData[30]
+ Tile_X5Y6_LUT4AB/FrameData[31] Tile_X5Y6_LUT4AB/FrameData[3] Tile_X5Y6_LUT4AB/FrameData[4]
+ Tile_X5Y6_LUT4AB/FrameData[5] Tile_X5Y6_LUT4AB/FrameData[6] Tile_X5Y6_LUT4AB/FrameData[7]
+ Tile_X5Y6_LUT4AB/FrameData[8] Tile_X5Y6_LUT4AB/FrameData[9] Tile_X6Y6_LUT4AB/FrameData[0]
+ Tile_X6Y6_LUT4AB/FrameData[10] Tile_X6Y6_LUT4AB/FrameData[11] Tile_X6Y6_LUT4AB/FrameData[12]
+ Tile_X6Y6_LUT4AB/FrameData[13] Tile_X6Y6_LUT4AB/FrameData[14] Tile_X6Y6_LUT4AB/FrameData[15]
+ Tile_X6Y6_LUT4AB/FrameData[16] Tile_X6Y6_LUT4AB/FrameData[17] Tile_X6Y6_LUT4AB/FrameData[18]
+ Tile_X6Y6_LUT4AB/FrameData[19] Tile_X6Y6_LUT4AB/FrameData[1] Tile_X6Y6_LUT4AB/FrameData[20]
+ Tile_X6Y6_LUT4AB/FrameData[21] Tile_X6Y6_LUT4AB/FrameData[22] Tile_X6Y6_LUT4AB/FrameData[23]
+ Tile_X6Y6_LUT4AB/FrameData[24] Tile_X6Y6_LUT4AB/FrameData[25] Tile_X6Y6_LUT4AB/FrameData[26]
+ Tile_X6Y6_LUT4AB/FrameData[27] Tile_X6Y6_LUT4AB/FrameData[28] Tile_X6Y6_LUT4AB/FrameData[29]
+ Tile_X6Y6_LUT4AB/FrameData[2] Tile_X6Y6_LUT4AB/FrameData[30] Tile_X6Y6_LUT4AB/FrameData[31]
+ Tile_X6Y6_LUT4AB/FrameData[3] Tile_X6Y6_LUT4AB/FrameData[4] Tile_X6Y6_LUT4AB/FrameData[5]
+ Tile_X6Y6_LUT4AB/FrameData[6] Tile_X6Y6_LUT4AB/FrameData[7] Tile_X6Y6_LUT4AB/FrameData[8]
+ Tile_X6Y6_LUT4AB/FrameData[9] Tile_X5Y6_LUT4AB/FrameStrobe[0] Tile_X5Y6_LUT4AB/FrameStrobe[10]
+ Tile_X5Y6_LUT4AB/FrameStrobe[11] Tile_X5Y6_LUT4AB/FrameStrobe[12] Tile_X5Y6_LUT4AB/FrameStrobe[13]
+ Tile_X5Y6_LUT4AB/FrameStrobe[14] Tile_X5Y6_LUT4AB/FrameStrobe[15] Tile_X5Y6_LUT4AB/FrameStrobe[16]
+ Tile_X5Y6_LUT4AB/FrameStrobe[17] Tile_X5Y6_LUT4AB/FrameStrobe[18] Tile_X5Y6_LUT4AB/FrameStrobe[19]
+ Tile_X5Y6_LUT4AB/FrameStrobe[1] Tile_X5Y6_LUT4AB/FrameStrobe[2] Tile_X5Y6_LUT4AB/FrameStrobe[3]
+ Tile_X5Y6_LUT4AB/FrameStrobe[4] Tile_X5Y6_LUT4AB/FrameStrobe[5] Tile_X5Y6_LUT4AB/FrameStrobe[6]
+ Tile_X5Y6_LUT4AB/FrameStrobe[7] Tile_X5Y6_LUT4AB/FrameStrobe[8] Tile_X5Y6_LUT4AB/FrameStrobe[9]
+ Tile_X5Y5_LUT4AB/FrameStrobe[0] Tile_X5Y5_LUT4AB/FrameStrobe[10] Tile_X5Y5_LUT4AB/FrameStrobe[11]
+ Tile_X5Y5_LUT4AB/FrameStrobe[12] Tile_X5Y5_LUT4AB/FrameStrobe[13] Tile_X5Y5_LUT4AB/FrameStrobe[14]
+ Tile_X5Y5_LUT4AB/FrameStrobe[15] Tile_X5Y5_LUT4AB/FrameStrobe[16] Tile_X5Y5_LUT4AB/FrameStrobe[17]
+ Tile_X5Y5_LUT4AB/FrameStrobe[18] Tile_X5Y5_LUT4AB/FrameStrobe[19] Tile_X5Y5_LUT4AB/FrameStrobe[1]
+ Tile_X5Y5_LUT4AB/FrameStrobe[2] Tile_X5Y5_LUT4AB/FrameStrobe[3] Tile_X5Y5_LUT4AB/FrameStrobe[4]
+ Tile_X5Y5_LUT4AB/FrameStrobe[5] Tile_X5Y5_LUT4AB/FrameStrobe[6] Tile_X5Y5_LUT4AB/FrameStrobe[7]
+ Tile_X5Y5_LUT4AB/FrameStrobe[8] Tile_X5Y5_LUT4AB/FrameStrobe[9] Tile_X5Y6_LUT4AB/N1BEG[0]
+ Tile_X5Y6_LUT4AB/N1BEG[1] Tile_X5Y6_LUT4AB/N1BEG[2] Tile_X5Y6_LUT4AB/N1BEG[3] Tile_X5Y7_LUT4AB/N1BEG[0]
+ Tile_X5Y7_LUT4AB/N1BEG[1] Tile_X5Y7_LUT4AB/N1BEG[2] Tile_X5Y7_LUT4AB/N1BEG[3] Tile_X5Y6_LUT4AB/N2BEG[0]
+ Tile_X5Y6_LUT4AB/N2BEG[1] Tile_X5Y6_LUT4AB/N2BEG[2] Tile_X5Y6_LUT4AB/N2BEG[3] Tile_X5Y6_LUT4AB/N2BEG[4]
+ Tile_X5Y6_LUT4AB/N2BEG[5] Tile_X5Y6_LUT4AB/N2BEG[6] Tile_X5Y6_LUT4AB/N2BEG[7] Tile_X5Y5_LUT4AB/N2END[0]
+ Tile_X5Y5_LUT4AB/N2END[1] Tile_X5Y5_LUT4AB/N2END[2] Tile_X5Y5_LUT4AB/N2END[3] Tile_X5Y5_LUT4AB/N2END[4]
+ Tile_X5Y5_LUT4AB/N2END[5] Tile_X5Y5_LUT4AB/N2END[6] Tile_X5Y5_LUT4AB/N2END[7] Tile_X5Y6_LUT4AB/N2END[0]
+ Tile_X5Y6_LUT4AB/N2END[1] Tile_X5Y6_LUT4AB/N2END[2] Tile_X5Y6_LUT4AB/N2END[3] Tile_X5Y6_LUT4AB/N2END[4]
+ Tile_X5Y6_LUT4AB/N2END[5] Tile_X5Y6_LUT4AB/N2END[6] Tile_X5Y6_LUT4AB/N2END[7] Tile_X5Y7_LUT4AB/N2BEG[0]
+ Tile_X5Y7_LUT4AB/N2BEG[1] Tile_X5Y7_LUT4AB/N2BEG[2] Tile_X5Y7_LUT4AB/N2BEG[3] Tile_X5Y7_LUT4AB/N2BEG[4]
+ Tile_X5Y7_LUT4AB/N2BEG[5] Tile_X5Y7_LUT4AB/N2BEG[6] Tile_X5Y7_LUT4AB/N2BEG[7] Tile_X5Y6_LUT4AB/N4BEG[0]
+ Tile_X5Y6_LUT4AB/N4BEG[10] Tile_X5Y6_LUT4AB/N4BEG[11] Tile_X5Y6_LUT4AB/N4BEG[12]
+ Tile_X5Y6_LUT4AB/N4BEG[13] Tile_X5Y6_LUT4AB/N4BEG[14] Tile_X5Y6_LUT4AB/N4BEG[15]
+ Tile_X5Y6_LUT4AB/N4BEG[1] Tile_X5Y6_LUT4AB/N4BEG[2] Tile_X5Y6_LUT4AB/N4BEG[3] Tile_X5Y6_LUT4AB/N4BEG[4]
+ Tile_X5Y6_LUT4AB/N4BEG[5] Tile_X5Y6_LUT4AB/N4BEG[6] Tile_X5Y6_LUT4AB/N4BEG[7] Tile_X5Y6_LUT4AB/N4BEG[8]
+ Tile_X5Y6_LUT4AB/N4BEG[9] Tile_X5Y7_LUT4AB/N4BEG[0] Tile_X5Y7_LUT4AB/N4BEG[10] Tile_X5Y7_LUT4AB/N4BEG[11]
+ Tile_X5Y7_LUT4AB/N4BEG[12] Tile_X5Y7_LUT4AB/N4BEG[13] Tile_X5Y7_LUT4AB/N4BEG[14]
+ Tile_X5Y7_LUT4AB/N4BEG[15] Tile_X5Y7_LUT4AB/N4BEG[1] Tile_X5Y7_LUT4AB/N4BEG[2] Tile_X5Y7_LUT4AB/N4BEG[3]
+ Tile_X5Y7_LUT4AB/N4BEG[4] Tile_X5Y7_LUT4AB/N4BEG[5] Tile_X5Y7_LUT4AB/N4BEG[6] Tile_X5Y7_LUT4AB/N4BEG[7]
+ Tile_X5Y7_LUT4AB/N4BEG[8] Tile_X5Y7_LUT4AB/N4BEG[9] Tile_X5Y6_LUT4AB/NN4BEG[0] Tile_X5Y6_LUT4AB/NN4BEG[10]
+ Tile_X5Y6_LUT4AB/NN4BEG[11] Tile_X5Y6_LUT4AB/NN4BEG[12] Tile_X5Y6_LUT4AB/NN4BEG[13]
+ Tile_X5Y6_LUT4AB/NN4BEG[14] Tile_X5Y6_LUT4AB/NN4BEG[15] Tile_X5Y6_LUT4AB/NN4BEG[1]
+ Tile_X5Y6_LUT4AB/NN4BEG[2] Tile_X5Y6_LUT4AB/NN4BEG[3] Tile_X5Y6_LUT4AB/NN4BEG[4]
+ Tile_X5Y6_LUT4AB/NN4BEG[5] Tile_X5Y6_LUT4AB/NN4BEG[6] Tile_X5Y6_LUT4AB/NN4BEG[7]
+ Tile_X5Y6_LUT4AB/NN4BEG[8] Tile_X5Y6_LUT4AB/NN4BEG[9] Tile_X5Y7_LUT4AB/NN4BEG[0]
+ Tile_X5Y7_LUT4AB/NN4BEG[10] Tile_X5Y7_LUT4AB/NN4BEG[11] Tile_X5Y7_LUT4AB/NN4BEG[12]
+ Tile_X5Y7_LUT4AB/NN4BEG[13] Tile_X5Y7_LUT4AB/NN4BEG[14] Tile_X5Y7_LUT4AB/NN4BEG[15]
+ Tile_X5Y7_LUT4AB/NN4BEG[1] Tile_X5Y7_LUT4AB/NN4BEG[2] Tile_X5Y7_LUT4AB/NN4BEG[3]
+ Tile_X5Y7_LUT4AB/NN4BEG[4] Tile_X5Y7_LUT4AB/NN4BEG[5] Tile_X5Y7_LUT4AB/NN4BEG[6]
+ Tile_X5Y7_LUT4AB/NN4BEG[7] Tile_X5Y7_LUT4AB/NN4BEG[8] Tile_X5Y7_LUT4AB/NN4BEG[9]
+ Tile_X5Y7_LUT4AB/S1END[0] Tile_X5Y7_LUT4AB/S1END[1] Tile_X5Y7_LUT4AB/S1END[2] Tile_X5Y7_LUT4AB/S1END[3]
+ Tile_X5Y6_LUT4AB/S1END[0] Tile_X5Y6_LUT4AB/S1END[1] Tile_X5Y6_LUT4AB/S1END[2] Tile_X5Y6_LUT4AB/S1END[3]
+ Tile_X5Y7_LUT4AB/S2MID[0] Tile_X5Y7_LUT4AB/S2MID[1] Tile_X5Y7_LUT4AB/S2MID[2] Tile_X5Y7_LUT4AB/S2MID[3]
+ Tile_X5Y7_LUT4AB/S2MID[4] Tile_X5Y7_LUT4AB/S2MID[5] Tile_X5Y7_LUT4AB/S2MID[6] Tile_X5Y7_LUT4AB/S2MID[7]
+ Tile_X5Y7_LUT4AB/S2END[0] Tile_X5Y7_LUT4AB/S2END[1] Tile_X5Y7_LUT4AB/S2END[2] Tile_X5Y7_LUT4AB/S2END[3]
+ Tile_X5Y7_LUT4AB/S2END[4] Tile_X5Y7_LUT4AB/S2END[5] Tile_X5Y7_LUT4AB/S2END[6] Tile_X5Y7_LUT4AB/S2END[7]
+ Tile_X5Y6_LUT4AB/S2END[0] Tile_X5Y6_LUT4AB/S2END[1] Tile_X5Y6_LUT4AB/S2END[2] Tile_X5Y6_LUT4AB/S2END[3]
+ Tile_X5Y6_LUT4AB/S2END[4] Tile_X5Y6_LUT4AB/S2END[5] Tile_X5Y6_LUT4AB/S2END[6] Tile_X5Y6_LUT4AB/S2END[7]
+ Tile_X5Y6_LUT4AB/S2MID[0] Tile_X5Y6_LUT4AB/S2MID[1] Tile_X5Y6_LUT4AB/S2MID[2] Tile_X5Y6_LUT4AB/S2MID[3]
+ Tile_X5Y6_LUT4AB/S2MID[4] Tile_X5Y6_LUT4AB/S2MID[5] Tile_X5Y6_LUT4AB/S2MID[6] Tile_X5Y6_LUT4AB/S2MID[7]
+ Tile_X5Y7_LUT4AB/S4END[0] Tile_X5Y7_LUT4AB/S4END[10] Tile_X5Y7_LUT4AB/S4END[11]
+ Tile_X5Y7_LUT4AB/S4END[12] Tile_X5Y7_LUT4AB/S4END[13] Tile_X5Y7_LUT4AB/S4END[14]
+ Tile_X5Y7_LUT4AB/S4END[15] Tile_X5Y7_LUT4AB/S4END[1] Tile_X5Y7_LUT4AB/S4END[2] Tile_X5Y7_LUT4AB/S4END[3]
+ Tile_X5Y7_LUT4AB/S4END[4] Tile_X5Y7_LUT4AB/S4END[5] Tile_X5Y7_LUT4AB/S4END[6] Tile_X5Y7_LUT4AB/S4END[7]
+ Tile_X5Y7_LUT4AB/S4END[8] Tile_X5Y7_LUT4AB/S4END[9] Tile_X5Y6_LUT4AB/S4END[0] Tile_X5Y6_LUT4AB/S4END[10]
+ Tile_X5Y6_LUT4AB/S4END[11] Tile_X5Y6_LUT4AB/S4END[12] Tile_X5Y6_LUT4AB/S4END[13]
+ Tile_X5Y6_LUT4AB/S4END[14] Tile_X5Y6_LUT4AB/S4END[15] Tile_X5Y6_LUT4AB/S4END[1]
+ Tile_X5Y6_LUT4AB/S4END[2] Tile_X5Y6_LUT4AB/S4END[3] Tile_X5Y6_LUT4AB/S4END[4] Tile_X5Y6_LUT4AB/S4END[5]
+ Tile_X5Y6_LUT4AB/S4END[6] Tile_X5Y6_LUT4AB/S4END[7] Tile_X5Y6_LUT4AB/S4END[8] Tile_X5Y6_LUT4AB/S4END[9]
+ Tile_X5Y7_LUT4AB/SS4END[0] Tile_X5Y7_LUT4AB/SS4END[10] Tile_X5Y7_LUT4AB/SS4END[11]
+ Tile_X5Y7_LUT4AB/SS4END[12] Tile_X5Y7_LUT4AB/SS4END[13] Tile_X5Y7_LUT4AB/SS4END[14]
+ Tile_X5Y7_LUT4AB/SS4END[15] Tile_X5Y7_LUT4AB/SS4END[1] Tile_X5Y7_LUT4AB/SS4END[2]
+ Tile_X5Y7_LUT4AB/SS4END[3] Tile_X5Y7_LUT4AB/SS4END[4] Tile_X5Y7_LUT4AB/SS4END[5]
+ Tile_X5Y7_LUT4AB/SS4END[6] Tile_X5Y7_LUT4AB/SS4END[7] Tile_X5Y7_LUT4AB/SS4END[8]
+ Tile_X5Y7_LUT4AB/SS4END[9] Tile_X5Y6_LUT4AB/SS4END[0] Tile_X5Y6_LUT4AB/SS4END[10]
+ Tile_X5Y6_LUT4AB/SS4END[11] Tile_X5Y6_LUT4AB/SS4END[12] Tile_X5Y6_LUT4AB/SS4END[13]
+ Tile_X5Y6_LUT4AB/SS4END[14] Tile_X5Y6_LUT4AB/SS4END[15] Tile_X5Y6_LUT4AB/SS4END[1]
+ Tile_X5Y6_LUT4AB/SS4END[2] Tile_X5Y6_LUT4AB/SS4END[3] Tile_X5Y6_LUT4AB/SS4END[4]
+ Tile_X5Y6_LUT4AB/SS4END[5] Tile_X5Y6_LUT4AB/SS4END[6] Tile_X5Y6_LUT4AB/SS4END[7]
+ Tile_X5Y6_LUT4AB/SS4END[8] Tile_X5Y6_LUT4AB/SS4END[9] Tile_X5Y6_LUT4AB/UserCLK Tile_X5Y5_LUT4AB/UserCLK
+ VGND VPWR Tile_X5Y6_LUT4AB/W1BEG[0] Tile_X5Y6_LUT4AB/W1BEG[1] Tile_X5Y6_LUT4AB/W1BEG[2]
+ Tile_X5Y6_LUT4AB/W1BEG[3] Tile_X6Y6_LUT4AB/W1BEG[0] Tile_X6Y6_LUT4AB/W1BEG[1] Tile_X6Y6_LUT4AB/W1BEG[2]
+ Tile_X6Y6_LUT4AB/W1BEG[3] Tile_X5Y6_LUT4AB/W2BEG[0] Tile_X5Y6_LUT4AB/W2BEG[1] Tile_X5Y6_LUT4AB/W2BEG[2]
+ Tile_X5Y6_LUT4AB/W2BEG[3] Tile_X5Y6_LUT4AB/W2BEG[4] Tile_X5Y6_LUT4AB/W2BEG[5] Tile_X5Y6_LUT4AB/W2BEG[6]
+ Tile_X5Y6_LUT4AB/W2BEG[7] Tile_X5Y6_LUT4AB/W2BEGb[0] Tile_X5Y6_LUT4AB/W2BEGb[1]
+ Tile_X5Y6_LUT4AB/W2BEGb[2] Tile_X5Y6_LUT4AB/W2BEGb[3] Tile_X5Y6_LUT4AB/W2BEGb[4]
+ Tile_X5Y6_LUT4AB/W2BEGb[5] Tile_X5Y6_LUT4AB/W2BEGb[6] Tile_X5Y6_LUT4AB/W2BEGb[7]
+ Tile_X5Y6_LUT4AB/W2END[0] Tile_X5Y6_LUT4AB/W2END[1] Tile_X5Y6_LUT4AB/W2END[2] Tile_X5Y6_LUT4AB/W2END[3]
+ Tile_X5Y6_LUT4AB/W2END[4] Tile_X5Y6_LUT4AB/W2END[5] Tile_X5Y6_LUT4AB/W2END[6] Tile_X5Y6_LUT4AB/W2END[7]
+ Tile_X6Y6_LUT4AB/W2BEG[0] Tile_X6Y6_LUT4AB/W2BEG[1] Tile_X6Y6_LUT4AB/W2BEG[2] Tile_X6Y6_LUT4AB/W2BEG[3]
+ Tile_X6Y6_LUT4AB/W2BEG[4] Tile_X6Y6_LUT4AB/W2BEG[5] Tile_X6Y6_LUT4AB/W2BEG[6] Tile_X6Y6_LUT4AB/W2BEG[7]
+ Tile_X5Y6_LUT4AB/W6BEG[0] Tile_X5Y6_LUT4AB/W6BEG[10] Tile_X5Y6_LUT4AB/W6BEG[11]
+ Tile_X5Y6_LUT4AB/W6BEG[1] Tile_X5Y6_LUT4AB/W6BEG[2] Tile_X5Y6_LUT4AB/W6BEG[3] Tile_X5Y6_LUT4AB/W6BEG[4]
+ Tile_X5Y6_LUT4AB/W6BEG[5] Tile_X5Y6_LUT4AB/W6BEG[6] Tile_X5Y6_LUT4AB/W6BEG[7] Tile_X5Y6_LUT4AB/W6BEG[8]
+ Tile_X5Y6_LUT4AB/W6BEG[9] Tile_X6Y6_LUT4AB/W6BEG[0] Tile_X6Y6_LUT4AB/W6BEG[10] Tile_X6Y6_LUT4AB/W6BEG[11]
+ Tile_X6Y6_LUT4AB/W6BEG[1] Tile_X6Y6_LUT4AB/W6BEG[2] Tile_X6Y6_LUT4AB/W6BEG[3] Tile_X6Y6_LUT4AB/W6BEG[4]
+ Tile_X6Y6_LUT4AB/W6BEG[5] Tile_X6Y6_LUT4AB/W6BEG[6] Tile_X6Y6_LUT4AB/W6BEG[7] Tile_X6Y6_LUT4AB/W6BEG[8]
+ Tile_X6Y6_LUT4AB/W6BEG[9] Tile_X5Y6_LUT4AB/WW4BEG[0] Tile_X5Y6_LUT4AB/WW4BEG[10]
+ Tile_X5Y6_LUT4AB/WW4BEG[11] Tile_X5Y6_LUT4AB/WW4BEG[12] Tile_X5Y6_LUT4AB/WW4BEG[13]
+ Tile_X5Y6_LUT4AB/WW4BEG[14] Tile_X5Y6_LUT4AB/WW4BEG[15] Tile_X5Y6_LUT4AB/WW4BEG[1]
+ Tile_X5Y6_LUT4AB/WW4BEG[2] Tile_X5Y6_LUT4AB/WW4BEG[3] Tile_X5Y6_LUT4AB/WW4BEG[4]
+ Tile_X5Y6_LUT4AB/WW4BEG[5] Tile_X5Y6_LUT4AB/WW4BEG[6] Tile_X5Y6_LUT4AB/WW4BEG[7]
+ Tile_X5Y6_LUT4AB/WW4BEG[8] Tile_X5Y6_LUT4AB/WW4BEG[9] Tile_X6Y6_LUT4AB/WW4BEG[0]
+ Tile_X6Y6_LUT4AB/WW4BEG[10] Tile_X6Y6_LUT4AB/WW4BEG[11] Tile_X6Y6_LUT4AB/WW4BEG[12]
+ Tile_X6Y6_LUT4AB/WW4BEG[13] Tile_X6Y6_LUT4AB/WW4BEG[14] Tile_X6Y6_LUT4AB/WW4BEG[15]
+ Tile_X6Y6_LUT4AB/WW4BEG[1] Tile_X6Y6_LUT4AB/WW4BEG[2] Tile_X6Y6_LUT4AB/WW4BEG[3]
+ Tile_X6Y6_LUT4AB/WW4BEG[4] Tile_X6Y6_LUT4AB/WW4BEG[5] Tile_X6Y6_LUT4AB/WW4BEG[6]
+ Tile_X6Y6_LUT4AB/WW4BEG[7] Tile_X6Y6_LUT4AB/WW4BEG[8] Tile_X6Y6_LUT4AB/WW4BEG[9]
+ LUT4AB
XTile_X8Y11_LUT4AB Tile_X8Y12_LUT4AB/Co Tile_X8Y11_LUT4AB/Co Tile_X9Y11_LUT4AB/E1END[0]
+ Tile_X9Y11_LUT4AB/E1END[1] Tile_X9Y11_LUT4AB/E1END[2] Tile_X9Y11_LUT4AB/E1END[3]
+ Tile_X8Y11_LUT4AB/E1END[0] Tile_X8Y11_LUT4AB/E1END[1] Tile_X8Y11_LUT4AB/E1END[2]
+ Tile_X8Y11_LUT4AB/E1END[3] Tile_X9Y11_LUT4AB/E2MID[0] Tile_X9Y11_LUT4AB/E2MID[1]
+ Tile_X9Y11_LUT4AB/E2MID[2] Tile_X9Y11_LUT4AB/E2MID[3] Tile_X9Y11_LUT4AB/E2MID[4]
+ Tile_X9Y11_LUT4AB/E2MID[5] Tile_X9Y11_LUT4AB/E2MID[6] Tile_X9Y11_LUT4AB/E2MID[7]
+ Tile_X9Y11_LUT4AB/E2END[0] Tile_X9Y11_LUT4AB/E2END[1] Tile_X9Y11_LUT4AB/E2END[2]
+ Tile_X9Y11_LUT4AB/E2END[3] Tile_X9Y11_LUT4AB/E2END[4] Tile_X9Y11_LUT4AB/E2END[5]
+ Tile_X9Y11_LUT4AB/E2END[6] Tile_X9Y11_LUT4AB/E2END[7] Tile_X8Y11_LUT4AB/E2END[0]
+ Tile_X8Y11_LUT4AB/E2END[1] Tile_X8Y11_LUT4AB/E2END[2] Tile_X8Y11_LUT4AB/E2END[3]
+ Tile_X8Y11_LUT4AB/E2END[4] Tile_X8Y11_LUT4AB/E2END[5] Tile_X8Y11_LUT4AB/E2END[6]
+ Tile_X8Y11_LUT4AB/E2END[7] Tile_X8Y11_LUT4AB/E2MID[0] Tile_X8Y11_LUT4AB/E2MID[1]
+ Tile_X8Y11_LUT4AB/E2MID[2] Tile_X8Y11_LUT4AB/E2MID[3] Tile_X8Y11_LUT4AB/E2MID[4]
+ Tile_X8Y11_LUT4AB/E2MID[5] Tile_X8Y11_LUT4AB/E2MID[6] Tile_X8Y11_LUT4AB/E2MID[7]
+ Tile_X9Y11_LUT4AB/E6END[0] Tile_X9Y11_LUT4AB/E6END[10] Tile_X9Y11_LUT4AB/E6END[11]
+ Tile_X9Y11_LUT4AB/E6END[1] Tile_X9Y11_LUT4AB/E6END[2] Tile_X9Y11_LUT4AB/E6END[3]
+ Tile_X9Y11_LUT4AB/E6END[4] Tile_X9Y11_LUT4AB/E6END[5] Tile_X9Y11_LUT4AB/E6END[6]
+ Tile_X9Y11_LUT4AB/E6END[7] Tile_X9Y11_LUT4AB/E6END[8] Tile_X9Y11_LUT4AB/E6END[9]
+ Tile_X8Y11_LUT4AB/E6END[0] Tile_X8Y11_LUT4AB/E6END[10] Tile_X8Y11_LUT4AB/E6END[11]
+ Tile_X8Y11_LUT4AB/E6END[1] Tile_X8Y11_LUT4AB/E6END[2] Tile_X8Y11_LUT4AB/E6END[3]
+ Tile_X8Y11_LUT4AB/E6END[4] Tile_X8Y11_LUT4AB/E6END[5] Tile_X8Y11_LUT4AB/E6END[6]
+ Tile_X8Y11_LUT4AB/E6END[7] Tile_X8Y11_LUT4AB/E6END[8] Tile_X8Y11_LUT4AB/E6END[9]
+ Tile_X9Y11_LUT4AB/EE4END[0] Tile_X9Y11_LUT4AB/EE4END[10] Tile_X9Y11_LUT4AB/EE4END[11]
+ Tile_X9Y11_LUT4AB/EE4END[12] Tile_X9Y11_LUT4AB/EE4END[13] Tile_X9Y11_LUT4AB/EE4END[14]
+ Tile_X9Y11_LUT4AB/EE4END[15] Tile_X9Y11_LUT4AB/EE4END[1] Tile_X9Y11_LUT4AB/EE4END[2]
+ Tile_X9Y11_LUT4AB/EE4END[3] Tile_X9Y11_LUT4AB/EE4END[4] Tile_X9Y11_LUT4AB/EE4END[5]
+ Tile_X9Y11_LUT4AB/EE4END[6] Tile_X9Y11_LUT4AB/EE4END[7] Tile_X9Y11_LUT4AB/EE4END[8]
+ Tile_X9Y11_LUT4AB/EE4END[9] Tile_X8Y11_LUT4AB/EE4END[0] Tile_X8Y11_LUT4AB/EE4END[10]
+ Tile_X8Y11_LUT4AB/EE4END[11] Tile_X8Y11_LUT4AB/EE4END[12] Tile_X8Y11_LUT4AB/EE4END[13]
+ Tile_X8Y11_LUT4AB/EE4END[14] Tile_X8Y11_LUT4AB/EE4END[15] Tile_X8Y11_LUT4AB/EE4END[1]
+ Tile_X8Y11_LUT4AB/EE4END[2] Tile_X8Y11_LUT4AB/EE4END[3] Tile_X8Y11_LUT4AB/EE4END[4]
+ Tile_X8Y11_LUT4AB/EE4END[5] Tile_X8Y11_LUT4AB/EE4END[6] Tile_X8Y11_LUT4AB/EE4END[7]
+ Tile_X8Y11_LUT4AB/EE4END[8] Tile_X8Y11_LUT4AB/EE4END[9] Tile_X8Y11_LUT4AB/FrameData[0]
+ Tile_X8Y11_LUT4AB/FrameData[10] Tile_X8Y11_LUT4AB/FrameData[11] Tile_X8Y11_LUT4AB/FrameData[12]
+ Tile_X8Y11_LUT4AB/FrameData[13] Tile_X8Y11_LUT4AB/FrameData[14] Tile_X8Y11_LUT4AB/FrameData[15]
+ Tile_X8Y11_LUT4AB/FrameData[16] Tile_X8Y11_LUT4AB/FrameData[17] Tile_X8Y11_LUT4AB/FrameData[18]
+ Tile_X8Y11_LUT4AB/FrameData[19] Tile_X8Y11_LUT4AB/FrameData[1] Tile_X8Y11_LUT4AB/FrameData[20]
+ Tile_X8Y11_LUT4AB/FrameData[21] Tile_X8Y11_LUT4AB/FrameData[22] Tile_X8Y11_LUT4AB/FrameData[23]
+ Tile_X8Y11_LUT4AB/FrameData[24] Tile_X8Y11_LUT4AB/FrameData[25] Tile_X8Y11_LUT4AB/FrameData[26]
+ Tile_X8Y11_LUT4AB/FrameData[27] Tile_X8Y11_LUT4AB/FrameData[28] Tile_X8Y11_LUT4AB/FrameData[29]
+ Tile_X8Y11_LUT4AB/FrameData[2] Tile_X8Y11_LUT4AB/FrameData[30] Tile_X8Y11_LUT4AB/FrameData[31]
+ Tile_X8Y11_LUT4AB/FrameData[3] Tile_X8Y11_LUT4AB/FrameData[4] Tile_X8Y11_LUT4AB/FrameData[5]
+ Tile_X8Y11_LUT4AB/FrameData[6] Tile_X8Y11_LUT4AB/FrameData[7] Tile_X8Y11_LUT4AB/FrameData[8]
+ Tile_X8Y11_LUT4AB/FrameData[9] Tile_X9Y11_LUT4AB/FrameData[0] Tile_X9Y11_LUT4AB/FrameData[10]
+ Tile_X9Y11_LUT4AB/FrameData[11] Tile_X9Y11_LUT4AB/FrameData[12] Tile_X9Y11_LUT4AB/FrameData[13]
+ Tile_X9Y11_LUT4AB/FrameData[14] Tile_X9Y11_LUT4AB/FrameData[15] Tile_X9Y11_LUT4AB/FrameData[16]
+ Tile_X9Y11_LUT4AB/FrameData[17] Tile_X9Y11_LUT4AB/FrameData[18] Tile_X9Y11_LUT4AB/FrameData[19]
+ Tile_X9Y11_LUT4AB/FrameData[1] Tile_X9Y11_LUT4AB/FrameData[20] Tile_X9Y11_LUT4AB/FrameData[21]
+ Tile_X9Y11_LUT4AB/FrameData[22] Tile_X9Y11_LUT4AB/FrameData[23] Tile_X9Y11_LUT4AB/FrameData[24]
+ Tile_X9Y11_LUT4AB/FrameData[25] Tile_X9Y11_LUT4AB/FrameData[26] Tile_X9Y11_LUT4AB/FrameData[27]
+ Tile_X9Y11_LUT4AB/FrameData[28] Tile_X9Y11_LUT4AB/FrameData[29] Tile_X9Y11_LUT4AB/FrameData[2]
+ Tile_X9Y11_LUT4AB/FrameData[30] Tile_X9Y11_LUT4AB/FrameData[31] Tile_X9Y11_LUT4AB/FrameData[3]
+ Tile_X9Y11_LUT4AB/FrameData[4] Tile_X9Y11_LUT4AB/FrameData[5] Tile_X9Y11_LUT4AB/FrameData[6]
+ Tile_X9Y11_LUT4AB/FrameData[7] Tile_X9Y11_LUT4AB/FrameData[8] Tile_X9Y11_LUT4AB/FrameData[9]
+ Tile_X8Y11_LUT4AB/FrameStrobe[0] Tile_X8Y11_LUT4AB/FrameStrobe[10] Tile_X8Y11_LUT4AB/FrameStrobe[11]
+ Tile_X8Y11_LUT4AB/FrameStrobe[12] Tile_X8Y11_LUT4AB/FrameStrobe[13] Tile_X8Y11_LUT4AB/FrameStrobe[14]
+ Tile_X8Y11_LUT4AB/FrameStrobe[15] Tile_X8Y11_LUT4AB/FrameStrobe[16] Tile_X8Y11_LUT4AB/FrameStrobe[17]
+ Tile_X8Y11_LUT4AB/FrameStrobe[18] Tile_X8Y11_LUT4AB/FrameStrobe[19] Tile_X8Y11_LUT4AB/FrameStrobe[1]
+ Tile_X8Y11_LUT4AB/FrameStrobe[2] Tile_X8Y11_LUT4AB/FrameStrobe[3] Tile_X8Y11_LUT4AB/FrameStrobe[4]
+ Tile_X8Y11_LUT4AB/FrameStrobe[5] Tile_X8Y11_LUT4AB/FrameStrobe[6] Tile_X8Y11_LUT4AB/FrameStrobe[7]
+ Tile_X8Y11_LUT4AB/FrameStrobe[8] Tile_X8Y11_LUT4AB/FrameStrobe[9] Tile_X8Y10_LUT4AB/FrameStrobe[0]
+ Tile_X8Y10_LUT4AB/FrameStrobe[10] Tile_X8Y10_LUT4AB/FrameStrobe[11] Tile_X8Y10_LUT4AB/FrameStrobe[12]
+ Tile_X8Y10_LUT4AB/FrameStrobe[13] Tile_X8Y10_LUT4AB/FrameStrobe[14] Tile_X8Y10_LUT4AB/FrameStrobe[15]
+ Tile_X8Y10_LUT4AB/FrameStrobe[16] Tile_X8Y10_LUT4AB/FrameStrobe[17] Tile_X8Y10_LUT4AB/FrameStrobe[18]
+ Tile_X8Y10_LUT4AB/FrameStrobe[19] Tile_X8Y10_LUT4AB/FrameStrobe[1] Tile_X8Y10_LUT4AB/FrameStrobe[2]
+ Tile_X8Y10_LUT4AB/FrameStrobe[3] Tile_X8Y10_LUT4AB/FrameStrobe[4] Tile_X8Y10_LUT4AB/FrameStrobe[5]
+ Tile_X8Y10_LUT4AB/FrameStrobe[6] Tile_X8Y10_LUT4AB/FrameStrobe[7] Tile_X8Y10_LUT4AB/FrameStrobe[8]
+ Tile_X8Y10_LUT4AB/FrameStrobe[9] Tile_X8Y11_LUT4AB/N1BEG[0] Tile_X8Y11_LUT4AB/N1BEG[1]
+ Tile_X8Y11_LUT4AB/N1BEG[2] Tile_X8Y11_LUT4AB/N1BEG[3] Tile_X8Y12_LUT4AB/N1BEG[0]
+ Tile_X8Y12_LUT4AB/N1BEG[1] Tile_X8Y12_LUT4AB/N1BEG[2] Tile_X8Y12_LUT4AB/N1BEG[3]
+ Tile_X8Y11_LUT4AB/N2BEG[0] Tile_X8Y11_LUT4AB/N2BEG[1] Tile_X8Y11_LUT4AB/N2BEG[2]
+ Tile_X8Y11_LUT4AB/N2BEG[3] Tile_X8Y11_LUT4AB/N2BEG[4] Tile_X8Y11_LUT4AB/N2BEG[5]
+ Tile_X8Y11_LUT4AB/N2BEG[6] Tile_X8Y11_LUT4AB/N2BEG[7] Tile_X8Y10_LUT4AB/N2END[0]
+ Tile_X8Y10_LUT4AB/N2END[1] Tile_X8Y10_LUT4AB/N2END[2] Tile_X8Y10_LUT4AB/N2END[3]
+ Tile_X8Y10_LUT4AB/N2END[4] Tile_X8Y10_LUT4AB/N2END[5] Tile_X8Y10_LUT4AB/N2END[6]
+ Tile_X8Y10_LUT4AB/N2END[7] Tile_X8Y11_LUT4AB/N2END[0] Tile_X8Y11_LUT4AB/N2END[1]
+ Tile_X8Y11_LUT4AB/N2END[2] Tile_X8Y11_LUT4AB/N2END[3] Tile_X8Y11_LUT4AB/N2END[4]
+ Tile_X8Y11_LUT4AB/N2END[5] Tile_X8Y11_LUT4AB/N2END[6] Tile_X8Y11_LUT4AB/N2END[7]
+ Tile_X8Y12_LUT4AB/N2BEG[0] Tile_X8Y12_LUT4AB/N2BEG[1] Tile_X8Y12_LUT4AB/N2BEG[2]
+ Tile_X8Y12_LUT4AB/N2BEG[3] Tile_X8Y12_LUT4AB/N2BEG[4] Tile_X8Y12_LUT4AB/N2BEG[5]
+ Tile_X8Y12_LUT4AB/N2BEG[6] Tile_X8Y12_LUT4AB/N2BEG[7] Tile_X8Y11_LUT4AB/N4BEG[0]
+ Tile_X8Y11_LUT4AB/N4BEG[10] Tile_X8Y11_LUT4AB/N4BEG[11] Tile_X8Y11_LUT4AB/N4BEG[12]
+ Tile_X8Y11_LUT4AB/N4BEG[13] Tile_X8Y11_LUT4AB/N4BEG[14] Tile_X8Y11_LUT4AB/N4BEG[15]
+ Tile_X8Y11_LUT4AB/N4BEG[1] Tile_X8Y11_LUT4AB/N4BEG[2] Tile_X8Y11_LUT4AB/N4BEG[3]
+ Tile_X8Y11_LUT4AB/N4BEG[4] Tile_X8Y11_LUT4AB/N4BEG[5] Tile_X8Y11_LUT4AB/N4BEG[6]
+ Tile_X8Y11_LUT4AB/N4BEG[7] Tile_X8Y11_LUT4AB/N4BEG[8] Tile_X8Y11_LUT4AB/N4BEG[9]
+ Tile_X8Y12_LUT4AB/N4BEG[0] Tile_X8Y12_LUT4AB/N4BEG[10] Tile_X8Y12_LUT4AB/N4BEG[11]
+ Tile_X8Y12_LUT4AB/N4BEG[12] Tile_X8Y12_LUT4AB/N4BEG[13] Tile_X8Y12_LUT4AB/N4BEG[14]
+ Tile_X8Y12_LUT4AB/N4BEG[15] Tile_X8Y12_LUT4AB/N4BEG[1] Tile_X8Y12_LUT4AB/N4BEG[2]
+ Tile_X8Y12_LUT4AB/N4BEG[3] Tile_X8Y12_LUT4AB/N4BEG[4] Tile_X8Y12_LUT4AB/N4BEG[5]
+ Tile_X8Y12_LUT4AB/N4BEG[6] Tile_X8Y12_LUT4AB/N4BEG[7] Tile_X8Y12_LUT4AB/N4BEG[8]
+ Tile_X8Y12_LUT4AB/N4BEG[9] Tile_X8Y11_LUT4AB/NN4BEG[0] Tile_X8Y11_LUT4AB/NN4BEG[10]
+ Tile_X8Y11_LUT4AB/NN4BEG[11] Tile_X8Y11_LUT4AB/NN4BEG[12] Tile_X8Y11_LUT4AB/NN4BEG[13]
+ Tile_X8Y11_LUT4AB/NN4BEG[14] Tile_X8Y11_LUT4AB/NN4BEG[15] Tile_X8Y11_LUT4AB/NN4BEG[1]
+ Tile_X8Y11_LUT4AB/NN4BEG[2] Tile_X8Y11_LUT4AB/NN4BEG[3] Tile_X8Y11_LUT4AB/NN4BEG[4]
+ Tile_X8Y11_LUT4AB/NN4BEG[5] Tile_X8Y11_LUT4AB/NN4BEG[6] Tile_X8Y11_LUT4AB/NN4BEG[7]
+ Tile_X8Y11_LUT4AB/NN4BEG[8] Tile_X8Y11_LUT4AB/NN4BEG[9] Tile_X8Y12_LUT4AB/NN4BEG[0]
+ Tile_X8Y12_LUT4AB/NN4BEG[10] Tile_X8Y12_LUT4AB/NN4BEG[11] Tile_X8Y12_LUT4AB/NN4BEG[12]
+ Tile_X8Y12_LUT4AB/NN4BEG[13] Tile_X8Y12_LUT4AB/NN4BEG[14] Tile_X8Y12_LUT4AB/NN4BEG[15]
+ Tile_X8Y12_LUT4AB/NN4BEG[1] Tile_X8Y12_LUT4AB/NN4BEG[2] Tile_X8Y12_LUT4AB/NN4BEG[3]
+ Tile_X8Y12_LUT4AB/NN4BEG[4] Tile_X8Y12_LUT4AB/NN4BEG[5] Tile_X8Y12_LUT4AB/NN4BEG[6]
+ Tile_X8Y12_LUT4AB/NN4BEG[7] Tile_X8Y12_LUT4AB/NN4BEG[8] Tile_X8Y12_LUT4AB/NN4BEG[9]
+ Tile_X8Y12_LUT4AB/S1END[0] Tile_X8Y12_LUT4AB/S1END[1] Tile_X8Y12_LUT4AB/S1END[2]
+ Tile_X8Y12_LUT4AB/S1END[3] Tile_X8Y11_LUT4AB/S1END[0] Tile_X8Y11_LUT4AB/S1END[1]
+ Tile_X8Y11_LUT4AB/S1END[2] Tile_X8Y11_LUT4AB/S1END[3] Tile_X8Y12_LUT4AB/S2MID[0]
+ Tile_X8Y12_LUT4AB/S2MID[1] Tile_X8Y12_LUT4AB/S2MID[2] Tile_X8Y12_LUT4AB/S2MID[3]
+ Tile_X8Y12_LUT4AB/S2MID[4] Tile_X8Y12_LUT4AB/S2MID[5] Tile_X8Y12_LUT4AB/S2MID[6]
+ Tile_X8Y12_LUT4AB/S2MID[7] Tile_X8Y12_LUT4AB/S2END[0] Tile_X8Y12_LUT4AB/S2END[1]
+ Tile_X8Y12_LUT4AB/S2END[2] Tile_X8Y12_LUT4AB/S2END[3] Tile_X8Y12_LUT4AB/S2END[4]
+ Tile_X8Y12_LUT4AB/S2END[5] Tile_X8Y12_LUT4AB/S2END[6] Tile_X8Y12_LUT4AB/S2END[7]
+ Tile_X8Y11_LUT4AB/S2END[0] Tile_X8Y11_LUT4AB/S2END[1] Tile_X8Y11_LUT4AB/S2END[2]
+ Tile_X8Y11_LUT4AB/S2END[3] Tile_X8Y11_LUT4AB/S2END[4] Tile_X8Y11_LUT4AB/S2END[5]
+ Tile_X8Y11_LUT4AB/S2END[6] Tile_X8Y11_LUT4AB/S2END[7] Tile_X8Y11_LUT4AB/S2MID[0]
+ Tile_X8Y11_LUT4AB/S2MID[1] Tile_X8Y11_LUT4AB/S2MID[2] Tile_X8Y11_LUT4AB/S2MID[3]
+ Tile_X8Y11_LUT4AB/S2MID[4] Tile_X8Y11_LUT4AB/S2MID[5] Tile_X8Y11_LUT4AB/S2MID[6]
+ Tile_X8Y11_LUT4AB/S2MID[7] Tile_X8Y12_LUT4AB/S4END[0] Tile_X8Y12_LUT4AB/S4END[10]
+ Tile_X8Y12_LUT4AB/S4END[11] Tile_X8Y12_LUT4AB/S4END[12] Tile_X8Y12_LUT4AB/S4END[13]
+ Tile_X8Y12_LUT4AB/S4END[14] Tile_X8Y12_LUT4AB/S4END[15] Tile_X8Y12_LUT4AB/S4END[1]
+ Tile_X8Y12_LUT4AB/S4END[2] Tile_X8Y12_LUT4AB/S4END[3] Tile_X8Y12_LUT4AB/S4END[4]
+ Tile_X8Y12_LUT4AB/S4END[5] Tile_X8Y12_LUT4AB/S4END[6] Tile_X8Y12_LUT4AB/S4END[7]
+ Tile_X8Y12_LUT4AB/S4END[8] Tile_X8Y12_LUT4AB/S4END[9] Tile_X8Y11_LUT4AB/S4END[0]
+ Tile_X8Y11_LUT4AB/S4END[10] Tile_X8Y11_LUT4AB/S4END[11] Tile_X8Y11_LUT4AB/S4END[12]
+ Tile_X8Y11_LUT4AB/S4END[13] Tile_X8Y11_LUT4AB/S4END[14] Tile_X8Y11_LUT4AB/S4END[15]
+ Tile_X8Y11_LUT4AB/S4END[1] Tile_X8Y11_LUT4AB/S4END[2] Tile_X8Y11_LUT4AB/S4END[3]
+ Tile_X8Y11_LUT4AB/S4END[4] Tile_X8Y11_LUT4AB/S4END[5] Tile_X8Y11_LUT4AB/S4END[6]
+ Tile_X8Y11_LUT4AB/S4END[7] Tile_X8Y11_LUT4AB/S4END[8] Tile_X8Y11_LUT4AB/S4END[9]
+ Tile_X8Y12_LUT4AB/SS4END[0] Tile_X8Y12_LUT4AB/SS4END[10] Tile_X8Y12_LUT4AB/SS4END[11]
+ Tile_X8Y12_LUT4AB/SS4END[12] Tile_X8Y12_LUT4AB/SS4END[13] Tile_X8Y12_LUT4AB/SS4END[14]
+ Tile_X8Y12_LUT4AB/SS4END[15] Tile_X8Y12_LUT4AB/SS4END[1] Tile_X8Y12_LUT4AB/SS4END[2]
+ Tile_X8Y12_LUT4AB/SS4END[3] Tile_X8Y12_LUT4AB/SS4END[4] Tile_X8Y12_LUT4AB/SS4END[5]
+ Tile_X8Y12_LUT4AB/SS4END[6] Tile_X8Y12_LUT4AB/SS4END[7] Tile_X8Y12_LUT4AB/SS4END[8]
+ Tile_X8Y12_LUT4AB/SS4END[9] Tile_X8Y11_LUT4AB/SS4END[0] Tile_X8Y11_LUT4AB/SS4END[10]
+ Tile_X8Y11_LUT4AB/SS4END[11] Tile_X8Y11_LUT4AB/SS4END[12] Tile_X8Y11_LUT4AB/SS4END[13]
+ Tile_X8Y11_LUT4AB/SS4END[14] Tile_X8Y11_LUT4AB/SS4END[15] Tile_X8Y11_LUT4AB/SS4END[1]
+ Tile_X8Y11_LUT4AB/SS4END[2] Tile_X8Y11_LUT4AB/SS4END[3] Tile_X8Y11_LUT4AB/SS4END[4]
+ Tile_X8Y11_LUT4AB/SS4END[5] Tile_X8Y11_LUT4AB/SS4END[6] Tile_X8Y11_LUT4AB/SS4END[7]
+ Tile_X8Y11_LUT4AB/SS4END[8] Tile_X8Y11_LUT4AB/SS4END[9] Tile_X8Y11_LUT4AB/UserCLK
+ Tile_X8Y10_LUT4AB/UserCLK VGND VPWR Tile_X8Y11_LUT4AB/W1BEG[0] Tile_X8Y11_LUT4AB/W1BEG[1]
+ Tile_X8Y11_LUT4AB/W1BEG[2] Tile_X8Y11_LUT4AB/W1BEG[3] Tile_X9Y11_LUT4AB/W1BEG[0]
+ Tile_X9Y11_LUT4AB/W1BEG[1] Tile_X9Y11_LUT4AB/W1BEG[2] Tile_X9Y11_LUT4AB/W1BEG[3]
+ Tile_X8Y11_LUT4AB/W2BEG[0] Tile_X8Y11_LUT4AB/W2BEG[1] Tile_X8Y11_LUT4AB/W2BEG[2]
+ Tile_X8Y11_LUT4AB/W2BEG[3] Tile_X8Y11_LUT4AB/W2BEG[4] Tile_X8Y11_LUT4AB/W2BEG[5]
+ Tile_X8Y11_LUT4AB/W2BEG[6] Tile_X8Y11_LUT4AB/W2BEG[7] Tile_X8Y11_LUT4AB/W2BEGb[0]
+ Tile_X8Y11_LUT4AB/W2BEGb[1] Tile_X8Y11_LUT4AB/W2BEGb[2] Tile_X8Y11_LUT4AB/W2BEGb[3]
+ Tile_X8Y11_LUT4AB/W2BEGb[4] Tile_X8Y11_LUT4AB/W2BEGb[5] Tile_X8Y11_LUT4AB/W2BEGb[6]
+ Tile_X8Y11_LUT4AB/W2BEGb[7] Tile_X8Y11_LUT4AB/W2END[0] Tile_X8Y11_LUT4AB/W2END[1]
+ Tile_X8Y11_LUT4AB/W2END[2] Tile_X8Y11_LUT4AB/W2END[3] Tile_X8Y11_LUT4AB/W2END[4]
+ Tile_X8Y11_LUT4AB/W2END[5] Tile_X8Y11_LUT4AB/W2END[6] Tile_X8Y11_LUT4AB/W2END[7]
+ Tile_X9Y11_LUT4AB/W2BEG[0] Tile_X9Y11_LUT4AB/W2BEG[1] Tile_X9Y11_LUT4AB/W2BEG[2]
+ Tile_X9Y11_LUT4AB/W2BEG[3] Tile_X9Y11_LUT4AB/W2BEG[4] Tile_X9Y11_LUT4AB/W2BEG[5]
+ Tile_X9Y11_LUT4AB/W2BEG[6] Tile_X9Y11_LUT4AB/W2BEG[7] Tile_X8Y11_LUT4AB/W6BEG[0]
+ Tile_X8Y11_LUT4AB/W6BEG[10] Tile_X8Y11_LUT4AB/W6BEG[11] Tile_X8Y11_LUT4AB/W6BEG[1]
+ Tile_X8Y11_LUT4AB/W6BEG[2] Tile_X8Y11_LUT4AB/W6BEG[3] Tile_X8Y11_LUT4AB/W6BEG[4]
+ Tile_X8Y11_LUT4AB/W6BEG[5] Tile_X8Y11_LUT4AB/W6BEG[6] Tile_X8Y11_LUT4AB/W6BEG[7]
+ Tile_X8Y11_LUT4AB/W6BEG[8] Tile_X8Y11_LUT4AB/W6BEG[9] Tile_X9Y11_LUT4AB/W6BEG[0]
+ Tile_X9Y11_LUT4AB/W6BEG[10] Tile_X9Y11_LUT4AB/W6BEG[11] Tile_X9Y11_LUT4AB/W6BEG[1]
+ Tile_X9Y11_LUT4AB/W6BEG[2] Tile_X9Y11_LUT4AB/W6BEG[3] Tile_X9Y11_LUT4AB/W6BEG[4]
+ Tile_X9Y11_LUT4AB/W6BEG[5] Tile_X9Y11_LUT4AB/W6BEG[6] Tile_X9Y11_LUT4AB/W6BEG[7]
+ Tile_X9Y11_LUT4AB/W6BEG[8] Tile_X9Y11_LUT4AB/W6BEG[9] Tile_X8Y11_LUT4AB/WW4BEG[0]
+ Tile_X8Y11_LUT4AB/WW4BEG[10] Tile_X8Y11_LUT4AB/WW4BEG[11] Tile_X8Y11_LUT4AB/WW4BEG[12]
+ Tile_X8Y11_LUT4AB/WW4BEG[13] Tile_X8Y11_LUT4AB/WW4BEG[14] Tile_X8Y11_LUT4AB/WW4BEG[15]
+ Tile_X8Y11_LUT4AB/WW4BEG[1] Tile_X8Y11_LUT4AB/WW4BEG[2] Tile_X8Y11_LUT4AB/WW4BEG[3]
+ Tile_X8Y11_LUT4AB/WW4BEG[4] Tile_X8Y11_LUT4AB/WW4BEG[5] Tile_X8Y11_LUT4AB/WW4BEG[6]
+ Tile_X8Y11_LUT4AB/WW4BEG[7] Tile_X8Y11_LUT4AB/WW4BEG[8] Tile_X8Y11_LUT4AB/WW4BEG[9]
+ Tile_X9Y11_LUT4AB/WW4BEG[0] Tile_X9Y11_LUT4AB/WW4BEG[10] Tile_X9Y11_LUT4AB/WW4BEG[11]
+ Tile_X9Y11_LUT4AB/WW4BEG[12] Tile_X9Y11_LUT4AB/WW4BEG[13] Tile_X9Y11_LUT4AB/WW4BEG[14]
+ Tile_X9Y11_LUT4AB/WW4BEG[15] Tile_X9Y11_LUT4AB/WW4BEG[1] Tile_X9Y11_LUT4AB/WW4BEG[2]
+ Tile_X9Y11_LUT4AB/WW4BEG[3] Tile_X9Y11_LUT4AB/WW4BEG[4] Tile_X9Y11_LUT4AB/WW4BEG[5]
+ Tile_X9Y11_LUT4AB/WW4BEG[6] Tile_X9Y11_LUT4AB/WW4BEG[7] Tile_X9Y11_LUT4AB/WW4BEG[8]
+ Tile_X9Y11_LUT4AB/WW4BEG[9] LUT4AB
XTile_X2Y1_LUT4AB Tile_X2Y2_LUT4AB/Co Tile_X2Y0_N_IO/Ci Tile_X3Y1_LUT4AB/E1END[0]
+ Tile_X3Y1_LUT4AB/E1END[1] Tile_X3Y1_LUT4AB/E1END[2] Tile_X3Y1_LUT4AB/E1END[3] Tile_X2Y1_LUT4AB/E1END[0]
+ Tile_X2Y1_LUT4AB/E1END[1] Tile_X2Y1_LUT4AB/E1END[2] Tile_X2Y1_LUT4AB/E1END[3] Tile_X3Y1_LUT4AB/E2MID[0]
+ Tile_X3Y1_LUT4AB/E2MID[1] Tile_X3Y1_LUT4AB/E2MID[2] Tile_X3Y1_LUT4AB/E2MID[3] Tile_X3Y1_LUT4AB/E2MID[4]
+ Tile_X3Y1_LUT4AB/E2MID[5] Tile_X3Y1_LUT4AB/E2MID[6] Tile_X3Y1_LUT4AB/E2MID[7] Tile_X3Y1_LUT4AB/E2END[0]
+ Tile_X3Y1_LUT4AB/E2END[1] Tile_X3Y1_LUT4AB/E2END[2] Tile_X3Y1_LUT4AB/E2END[3] Tile_X3Y1_LUT4AB/E2END[4]
+ Tile_X3Y1_LUT4AB/E2END[5] Tile_X3Y1_LUT4AB/E2END[6] Tile_X3Y1_LUT4AB/E2END[7] Tile_X2Y1_LUT4AB/E2END[0]
+ Tile_X2Y1_LUT4AB/E2END[1] Tile_X2Y1_LUT4AB/E2END[2] Tile_X2Y1_LUT4AB/E2END[3] Tile_X2Y1_LUT4AB/E2END[4]
+ Tile_X2Y1_LUT4AB/E2END[5] Tile_X2Y1_LUT4AB/E2END[6] Tile_X2Y1_LUT4AB/E2END[7] Tile_X2Y1_LUT4AB/E2MID[0]
+ Tile_X2Y1_LUT4AB/E2MID[1] Tile_X2Y1_LUT4AB/E2MID[2] Tile_X2Y1_LUT4AB/E2MID[3] Tile_X2Y1_LUT4AB/E2MID[4]
+ Tile_X2Y1_LUT4AB/E2MID[5] Tile_X2Y1_LUT4AB/E2MID[6] Tile_X2Y1_LUT4AB/E2MID[7] Tile_X3Y1_LUT4AB/E6END[0]
+ Tile_X3Y1_LUT4AB/E6END[10] Tile_X3Y1_LUT4AB/E6END[11] Tile_X3Y1_LUT4AB/E6END[1]
+ Tile_X3Y1_LUT4AB/E6END[2] Tile_X3Y1_LUT4AB/E6END[3] Tile_X3Y1_LUT4AB/E6END[4] Tile_X3Y1_LUT4AB/E6END[5]
+ Tile_X3Y1_LUT4AB/E6END[6] Tile_X3Y1_LUT4AB/E6END[7] Tile_X3Y1_LUT4AB/E6END[8] Tile_X3Y1_LUT4AB/E6END[9]
+ Tile_X2Y1_LUT4AB/E6END[0] Tile_X2Y1_LUT4AB/E6END[10] Tile_X2Y1_LUT4AB/E6END[11]
+ Tile_X2Y1_LUT4AB/E6END[1] Tile_X2Y1_LUT4AB/E6END[2] Tile_X2Y1_LUT4AB/E6END[3] Tile_X2Y1_LUT4AB/E6END[4]
+ Tile_X2Y1_LUT4AB/E6END[5] Tile_X2Y1_LUT4AB/E6END[6] Tile_X2Y1_LUT4AB/E6END[7] Tile_X2Y1_LUT4AB/E6END[8]
+ Tile_X2Y1_LUT4AB/E6END[9] Tile_X3Y1_LUT4AB/EE4END[0] Tile_X3Y1_LUT4AB/EE4END[10]
+ Tile_X3Y1_LUT4AB/EE4END[11] Tile_X3Y1_LUT4AB/EE4END[12] Tile_X3Y1_LUT4AB/EE4END[13]
+ Tile_X3Y1_LUT4AB/EE4END[14] Tile_X3Y1_LUT4AB/EE4END[15] Tile_X3Y1_LUT4AB/EE4END[1]
+ Tile_X3Y1_LUT4AB/EE4END[2] Tile_X3Y1_LUT4AB/EE4END[3] Tile_X3Y1_LUT4AB/EE4END[4]
+ Tile_X3Y1_LUT4AB/EE4END[5] Tile_X3Y1_LUT4AB/EE4END[6] Tile_X3Y1_LUT4AB/EE4END[7]
+ Tile_X3Y1_LUT4AB/EE4END[8] Tile_X3Y1_LUT4AB/EE4END[9] Tile_X2Y1_LUT4AB/EE4END[0]
+ Tile_X2Y1_LUT4AB/EE4END[10] Tile_X2Y1_LUT4AB/EE4END[11] Tile_X2Y1_LUT4AB/EE4END[12]
+ Tile_X2Y1_LUT4AB/EE4END[13] Tile_X2Y1_LUT4AB/EE4END[14] Tile_X2Y1_LUT4AB/EE4END[15]
+ Tile_X2Y1_LUT4AB/EE4END[1] Tile_X2Y1_LUT4AB/EE4END[2] Tile_X2Y1_LUT4AB/EE4END[3]
+ Tile_X2Y1_LUT4AB/EE4END[4] Tile_X2Y1_LUT4AB/EE4END[5] Tile_X2Y1_LUT4AB/EE4END[6]
+ Tile_X2Y1_LUT4AB/EE4END[7] Tile_X2Y1_LUT4AB/EE4END[8] Tile_X2Y1_LUT4AB/EE4END[9]
+ Tile_X2Y1_LUT4AB/FrameData[0] Tile_X2Y1_LUT4AB/FrameData[10] Tile_X2Y1_LUT4AB/FrameData[11]
+ Tile_X2Y1_LUT4AB/FrameData[12] Tile_X2Y1_LUT4AB/FrameData[13] Tile_X2Y1_LUT4AB/FrameData[14]
+ Tile_X2Y1_LUT4AB/FrameData[15] Tile_X2Y1_LUT4AB/FrameData[16] Tile_X2Y1_LUT4AB/FrameData[17]
+ Tile_X2Y1_LUT4AB/FrameData[18] Tile_X2Y1_LUT4AB/FrameData[19] Tile_X2Y1_LUT4AB/FrameData[1]
+ Tile_X2Y1_LUT4AB/FrameData[20] Tile_X2Y1_LUT4AB/FrameData[21] Tile_X2Y1_LUT4AB/FrameData[22]
+ Tile_X2Y1_LUT4AB/FrameData[23] Tile_X2Y1_LUT4AB/FrameData[24] Tile_X2Y1_LUT4AB/FrameData[25]
+ Tile_X2Y1_LUT4AB/FrameData[26] Tile_X2Y1_LUT4AB/FrameData[27] Tile_X2Y1_LUT4AB/FrameData[28]
+ Tile_X2Y1_LUT4AB/FrameData[29] Tile_X2Y1_LUT4AB/FrameData[2] Tile_X2Y1_LUT4AB/FrameData[30]
+ Tile_X2Y1_LUT4AB/FrameData[31] Tile_X2Y1_LUT4AB/FrameData[3] Tile_X2Y1_LUT4AB/FrameData[4]
+ Tile_X2Y1_LUT4AB/FrameData[5] Tile_X2Y1_LUT4AB/FrameData[6] Tile_X2Y1_LUT4AB/FrameData[7]
+ Tile_X2Y1_LUT4AB/FrameData[8] Tile_X2Y1_LUT4AB/FrameData[9] Tile_X3Y1_LUT4AB/FrameData[0]
+ Tile_X3Y1_LUT4AB/FrameData[10] Tile_X3Y1_LUT4AB/FrameData[11] Tile_X3Y1_LUT4AB/FrameData[12]
+ Tile_X3Y1_LUT4AB/FrameData[13] Tile_X3Y1_LUT4AB/FrameData[14] Tile_X3Y1_LUT4AB/FrameData[15]
+ Tile_X3Y1_LUT4AB/FrameData[16] Tile_X3Y1_LUT4AB/FrameData[17] Tile_X3Y1_LUT4AB/FrameData[18]
+ Tile_X3Y1_LUT4AB/FrameData[19] Tile_X3Y1_LUT4AB/FrameData[1] Tile_X3Y1_LUT4AB/FrameData[20]
+ Tile_X3Y1_LUT4AB/FrameData[21] Tile_X3Y1_LUT4AB/FrameData[22] Tile_X3Y1_LUT4AB/FrameData[23]
+ Tile_X3Y1_LUT4AB/FrameData[24] Tile_X3Y1_LUT4AB/FrameData[25] Tile_X3Y1_LUT4AB/FrameData[26]
+ Tile_X3Y1_LUT4AB/FrameData[27] Tile_X3Y1_LUT4AB/FrameData[28] Tile_X3Y1_LUT4AB/FrameData[29]
+ Tile_X3Y1_LUT4AB/FrameData[2] Tile_X3Y1_LUT4AB/FrameData[30] Tile_X3Y1_LUT4AB/FrameData[31]
+ Tile_X3Y1_LUT4AB/FrameData[3] Tile_X3Y1_LUT4AB/FrameData[4] Tile_X3Y1_LUT4AB/FrameData[5]
+ Tile_X3Y1_LUT4AB/FrameData[6] Tile_X3Y1_LUT4AB/FrameData[7] Tile_X3Y1_LUT4AB/FrameData[8]
+ Tile_X3Y1_LUT4AB/FrameData[9] Tile_X2Y1_LUT4AB/FrameStrobe[0] Tile_X2Y1_LUT4AB/FrameStrobe[10]
+ Tile_X2Y1_LUT4AB/FrameStrobe[11] Tile_X2Y1_LUT4AB/FrameStrobe[12] Tile_X2Y1_LUT4AB/FrameStrobe[13]
+ Tile_X2Y1_LUT4AB/FrameStrobe[14] Tile_X2Y1_LUT4AB/FrameStrobe[15] Tile_X2Y1_LUT4AB/FrameStrobe[16]
+ Tile_X2Y1_LUT4AB/FrameStrobe[17] Tile_X2Y1_LUT4AB/FrameStrobe[18] Tile_X2Y1_LUT4AB/FrameStrobe[19]
+ Tile_X2Y1_LUT4AB/FrameStrobe[1] Tile_X2Y1_LUT4AB/FrameStrobe[2] Tile_X2Y1_LUT4AB/FrameStrobe[3]
+ Tile_X2Y1_LUT4AB/FrameStrobe[4] Tile_X2Y1_LUT4AB/FrameStrobe[5] Tile_X2Y1_LUT4AB/FrameStrobe[6]
+ Tile_X2Y1_LUT4AB/FrameStrobe[7] Tile_X2Y1_LUT4AB/FrameStrobe[8] Tile_X2Y1_LUT4AB/FrameStrobe[9]
+ Tile_X2Y0_N_IO/FrameStrobe[0] Tile_X2Y0_N_IO/FrameStrobe[10] Tile_X2Y0_N_IO/FrameStrobe[11]
+ Tile_X2Y0_N_IO/FrameStrobe[12] Tile_X2Y0_N_IO/FrameStrobe[13] Tile_X2Y0_N_IO/FrameStrobe[14]
+ Tile_X2Y0_N_IO/FrameStrobe[15] Tile_X2Y0_N_IO/FrameStrobe[16] Tile_X2Y0_N_IO/FrameStrobe[17]
+ Tile_X2Y0_N_IO/FrameStrobe[18] Tile_X2Y0_N_IO/FrameStrobe[19] Tile_X2Y0_N_IO/FrameStrobe[1]
+ Tile_X2Y0_N_IO/FrameStrobe[2] Tile_X2Y0_N_IO/FrameStrobe[3] Tile_X2Y0_N_IO/FrameStrobe[4]
+ Tile_X2Y0_N_IO/FrameStrobe[5] Tile_X2Y0_N_IO/FrameStrobe[6] Tile_X2Y0_N_IO/FrameStrobe[7]
+ Tile_X2Y0_N_IO/FrameStrobe[8] Tile_X2Y0_N_IO/FrameStrobe[9] Tile_X2Y0_N_IO/N1END[0]
+ Tile_X2Y0_N_IO/N1END[1] Tile_X2Y0_N_IO/N1END[2] Tile_X2Y0_N_IO/N1END[3] Tile_X2Y2_LUT4AB/N1BEG[0]
+ Tile_X2Y2_LUT4AB/N1BEG[1] Tile_X2Y2_LUT4AB/N1BEG[2] Tile_X2Y2_LUT4AB/N1BEG[3] Tile_X2Y0_N_IO/N2MID[0]
+ Tile_X2Y0_N_IO/N2MID[1] Tile_X2Y0_N_IO/N2MID[2] Tile_X2Y0_N_IO/N2MID[3] Tile_X2Y0_N_IO/N2MID[4]
+ Tile_X2Y0_N_IO/N2MID[5] Tile_X2Y0_N_IO/N2MID[6] Tile_X2Y0_N_IO/N2MID[7] Tile_X2Y0_N_IO/N2END[0]
+ Tile_X2Y0_N_IO/N2END[1] Tile_X2Y0_N_IO/N2END[2] Tile_X2Y0_N_IO/N2END[3] Tile_X2Y0_N_IO/N2END[4]
+ Tile_X2Y0_N_IO/N2END[5] Tile_X2Y0_N_IO/N2END[6] Tile_X2Y0_N_IO/N2END[7] Tile_X2Y1_LUT4AB/N2END[0]
+ Tile_X2Y1_LUT4AB/N2END[1] Tile_X2Y1_LUT4AB/N2END[2] Tile_X2Y1_LUT4AB/N2END[3] Tile_X2Y1_LUT4AB/N2END[4]
+ Tile_X2Y1_LUT4AB/N2END[5] Tile_X2Y1_LUT4AB/N2END[6] Tile_X2Y1_LUT4AB/N2END[7] Tile_X2Y2_LUT4AB/N2BEG[0]
+ Tile_X2Y2_LUT4AB/N2BEG[1] Tile_X2Y2_LUT4AB/N2BEG[2] Tile_X2Y2_LUT4AB/N2BEG[3] Tile_X2Y2_LUT4AB/N2BEG[4]
+ Tile_X2Y2_LUT4AB/N2BEG[5] Tile_X2Y2_LUT4AB/N2BEG[6] Tile_X2Y2_LUT4AB/N2BEG[7] Tile_X2Y0_N_IO/N4END[0]
+ Tile_X2Y0_N_IO/N4END[10] Tile_X2Y0_N_IO/N4END[11] Tile_X2Y0_N_IO/N4END[12] Tile_X2Y0_N_IO/N4END[13]
+ Tile_X2Y0_N_IO/N4END[14] Tile_X2Y0_N_IO/N4END[15] Tile_X2Y0_N_IO/N4END[1] Tile_X2Y0_N_IO/N4END[2]
+ Tile_X2Y0_N_IO/N4END[3] Tile_X2Y0_N_IO/N4END[4] Tile_X2Y0_N_IO/N4END[5] Tile_X2Y0_N_IO/N4END[6]
+ Tile_X2Y0_N_IO/N4END[7] Tile_X2Y0_N_IO/N4END[8] Tile_X2Y0_N_IO/N4END[9] Tile_X2Y2_LUT4AB/N4BEG[0]
+ Tile_X2Y2_LUT4AB/N4BEG[10] Tile_X2Y2_LUT4AB/N4BEG[11] Tile_X2Y2_LUT4AB/N4BEG[12]
+ Tile_X2Y2_LUT4AB/N4BEG[13] Tile_X2Y2_LUT4AB/N4BEG[14] Tile_X2Y2_LUT4AB/N4BEG[15]
+ Tile_X2Y2_LUT4AB/N4BEG[1] Tile_X2Y2_LUT4AB/N4BEG[2] Tile_X2Y2_LUT4AB/N4BEG[3] Tile_X2Y2_LUT4AB/N4BEG[4]
+ Tile_X2Y2_LUT4AB/N4BEG[5] Tile_X2Y2_LUT4AB/N4BEG[6] Tile_X2Y2_LUT4AB/N4BEG[7] Tile_X2Y2_LUT4AB/N4BEG[8]
+ Tile_X2Y2_LUT4AB/N4BEG[9] Tile_X2Y0_N_IO/NN4END[0] Tile_X2Y0_N_IO/NN4END[10] Tile_X2Y0_N_IO/NN4END[11]
+ Tile_X2Y0_N_IO/NN4END[12] Tile_X2Y0_N_IO/NN4END[13] Tile_X2Y0_N_IO/NN4END[14] Tile_X2Y0_N_IO/NN4END[15]
+ Tile_X2Y0_N_IO/NN4END[1] Tile_X2Y0_N_IO/NN4END[2] Tile_X2Y0_N_IO/NN4END[3] Tile_X2Y0_N_IO/NN4END[4]
+ Tile_X2Y0_N_IO/NN4END[5] Tile_X2Y0_N_IO/NN4END[6] Tile_X2Y0_N_IO/NN4END[7] Tile_X2Y0_N_IO/NN4END[8]
+ Tile_X2Y0_N_IO/NN4END[9] Tile_X2Y2_LUT4AB/NN4BEG[0] Tile_X2Y2_LUT4AB/NN4BEG[10]
+ Tile_X2Y2_LUT4AB/NN4BEG[11] Tile_X2Y2_LUT4AB/NN4BEG[12] Tile_X2Y2_LUT4AB/NN4BEG[13]
+ Tile_X2Y2_LUT4AB/NN4BEG[14] Tile_X2Y2_LUT4AB/NN4BEG[15] Tile_X2Y2_LUT4AB/NN4BEG[1]
+ Tile_X2Y2_LUT4AB/NN4BEG[2] Tile_X2Y2_LUT4AB/NN4BEG[3] Tile_X2Y2_LUT4AB/NN4BEG[4]
+ Tile_X2Y2_LUT4AB/NN4BEG[5] Tile_X2Y2_LUT4AB/NN4BEG[6] Tile_X2Y2_LUT4AB/NN4BEG[7]
+ Tile_X2Y2_LUT4AB/NN4BEG[8] Tile_X2Y2_LUT4AB/NN4BEG[9] Tile_X2Y2_LUT4AB/S1END[0]
+ Tile_X2Y2_LUT4AB/S1END[1] Tile_X2Y2_LUT4AB/S1END[2] Tile_X2Y2_LUT4AB/S1END[3] Tile_X2Y0_N_IO/S1BEG[0]
+ Tile_X2Y0_N_IO/S1BEG[1] Tile_X2Y0_N_IO/S1BEG[2] Tile_X2Y0_N_IO/S1BEG[3] Tile_X2Y2_LUT4AB/S2MID[0]
+ Tile_X2Y2_LUT4AB/S2MID[1] Tile_X2Y2_LUT4AB/S2MID[2] Tile_X2Y2_LUT4AB/S2MID[3] Tile_X2Y2_LUT4AB/S2MID[4]
+ Tile_X2Y2_LUT4AB/S2MID[5] Tile_X2Y2_LUT4AB/S2MID[6] Tile_X2Y2_LUT4AB/S2MID[7] Tile_X2Y2_LUT4AB/S2END[0]
+ Tile_X2Y2_LUT4AB/S2END[1] Tile_X2Y2_LUT4AB/S2END[2] Tile_X2Y2_LUT4AB/S2END[3] Tile_X2Y2_LUT4AB/S2END[4]
+ Tile_X2Y2_LUT4AB/S2END[5] Tile_X2Y2_LUT4AB/S2END[6] Tile_X2Y2_LUT4AB/S2END[7] Tile_X2Y0_N_IO/S2BEGb[0]
+ Tile_X2Y0_N_IO/S2BEGb[1] Tile_X2Y0_N_IO/S2BEGb[2] Tile_X2Y0_N_IO/S2BEGb[3] Tile_X2Y0_N_IO/S2BEGb[4]
+ Tile_X2Y0_N_IO/S2BEGb[5] Tile_X2Y0_N_IO/S2BEGb[6] Tile_X2Y0_N_IO/S2BEGb[7] Tile_X2Y0_N_IO/S2BEG[0]
+ Tile_X2Y0_N_IO/S2BEG[1] Tile_X2Y0_N_IO/S2BEG[2] Tile_X2Y0_N_IO/S2BEG[3] Tile_X2Y0_N_IO/S2BEG[4]
+ Tile_X2Y0_N_IO/S2BEG[5] Tile_X2Y0_N_IO/S2BEG[6] Tile_X2Y0_N_IO/S2BEG[7] Tile_X2Y2_LUT4AB/S4END[0]
+ Tile_X2Y2_LUT4AB/S4END[10] Tile_X2Y2_LUT4AB/S4END[11] Tile_X2Y2_LUT4AB/S4END[12]
+ Tile_X2Y2_LUT4AB/S4END[13] Tile_X2Y2_LUT4AB/S4END[14] Tile_X2Y2_LUT4AB/S4END[15]
+ Tile_X2Y2_LUT4AB/S4END[1] Tile_X2Y2_LUT4AB/S4END[2] Tile_X2Y2_LUT4AB/S4END[3] Tile_X2Y2_LUT4AB/S4END[4]
+ Tile_X2Y2_LUT4AB/S4END[5] Tile_X2Y2_LUT4AB/S4END[6] Tile_X2Y2_LUT4AB/S4END[7] Tile_X2Y2_LUT4AB/S4END[8]
+ Tile_X2Y2_LUT4AB/S4END[9] Tile_X2Y0_N_IO/S4BEG[0] Tile_X2Y0_N_IO/S4BEG[10] Tile_X2Y0_N_IO/S4BEG[11]
+ Tile_X2Y0_N_IO/S4BEG[12] Tile_X2Y0_N_IO/S4BEG[13] Tile_X2Y0_N_IO/S4BEG[14] Tile_X2Y0_N_IO/S4BEG[15]
+ Tile_X2Y0_N_IO/S4BEG[1] Tile_X2Y0_N_IO/S4BEG[2] Tile_X2Y0_N_IO/S4BEG[3] Tile_X2Y0_N_IO/S4BEG[4]
+ Tile_X2Y0_N_IO/S4BEG[5] Tile_X2Y0_N_IO/S4BEG[6] Tile_X2Y0_N_IO/S4BEG[7] Tile_X2Y0_N_IO/S4BEG[8]
+ Tile_X2Y0_N_IO/S4BEG[9] Tile_X2Y2_LUT4AB/SS4END[0] Tile_X2Y2_LUT4AB/SS4END[10] Tile_X2Y2_LUT4AB/SS4END[11]
+ Tile_X2Y2_LUT4AB/SS4END[12] Tile_X2Y2_LUT4AB/SS4END[13] Tile_X2Y2_LUT4AB/SS4END[14]
+ Tile_X2Y2_LUT4AB/SS4END[15] Tile_X2Y2_LUT4AB/SS4END[1] Tile_X2Y2_LUT4AB/SS4END[2]
+ Tile_X2Y2_LUT4AB/SS4END[3] Tile_X2Y2_LUT4AB/SS4END[4] Tile_X2Y2_LUT4AB/SS4END[5]
+ Tile_X2Y2_LUT4AB/SS4END[6] Tile_X2Y2_LUT4AB/SS4END[7] Tile_X2Y2_LUT4AB/SS4END[8]
+ Tile_X2Y2_LUT4AB/SS4END[9] Tile_X2Y0_N_IO/SS4BEG[0] Tile_X2Y0_N_IO/SS4BEG[10] Tile_X2Y0_N_IO/SS4BEG[11]
+ Tile_X2Y0_N_IO/SS4BEG[12] Tile_X2Y0_N_IO/SS4BEG[13] Tile_X2Y0_N_IO/SS4BEG[14] Tile_X2Y0_N_IO/SS4BEG[15]
+ Tile_X2Y0_N_IO/SS4BEG[1] Tile_X2Y0_N_IO/SS4BEG[2] Tile_X2Y0_N_IO/SS4BEG[3] Tile_X2Y0_N_IO/SS4BEG[4]
+ Tile_X2Y0_N_IO/SS4BEG[5] Tile_X2Y0_N_IO/SS4BEG[6] Tile_X2Y0_N_IO/SS4BEG[7] Tile_X2Y0_N_IO/SS4BEG[8]
+ Tile_X2Y0_N_IO/SS4BEG[9] Tile_X2Y1_LUT4AB/UserCLK Tile_X2Y0_N_IO/UserCLK VGND VPWR
+ Tile_X2Y1_LUT4AB/W1BEG[0] Tile_X2Y1_LUT4AB/W1BEG[1] Tile_X2Y1_LUT4AB/W1BEG[2] Tile_X2Y1_LUT4AB/W1BEG[3]
+ Tile_X3Y1_LUT4AB/W1BEG[0] Tile_X3Y1_LUT4AB/W1BEG[1] Tile_X3Y1_LUT4AB/W1BEG[2] Tile_X3Y1_LUT4AB/W1BEG[3]
+ Tile_X2Y1_LUT4AB/W2BEG[0] Tile_X2Y1_LUT4AB/W2BEG[1] Tile_X2Y1_LUT4AB/W2BEG[2] Tile_X2Y1_LUT4AB/W2BEG[3]
+ Tile_X2Y1_LUT4AB/W2BEG[4] Tile_X2Y1_LUT4AB/W2BEG[5] Tile_X2Y1_LUT4AB/W2BEG[6] Tile_X2Y1_LUT4AB/W2BEG[7]
+ Tile_X1Y1_LUT4AB/W2END[0] Tile_X1Y1_LUT4AB/W2END[1] Tile_X1Y1_LUT4AB/W2END[2] Tile_X1Y1_LUT4AB/W2END[3]
+ Tile_X1Y1_LUT4AB/W2END[4] Tile_X1Y1_LUT4AB/W2END[5] Tile_X1Y1_LUT4AB/W2END[6] Tile_X1Y1_LUT4AB/W2END[7]
+ Tile_X2Y1_LUT4AB/W2END[0] Tile_X2Y1_LUT4AB/W2END[1] Tile_X2Y1_LUT4AB/W2END[2] Tile_X2Y1_LUT4AB/W2END[3]
+ Tile_X2Y1_LUT4AB/W2END[4] Tile_X2Y1_LUT4AB/W2END[5] Tile_X2Y1_LUT4AB/W2END[6] Tile_X2Y1_LUT4AB/W2END[7]
+ Tile_X3Y1_LUT4AB/W2BEG[0] Tile_X3Y1_LUT4AB/W2BEG[1] Tile_X3Y1_LUT4AB/W2BEG[2] Tile_X3Y1_LUT4AB/W2BEG[3]
+ Tile_X3Y1_LUT4AB/W2BEG[4] Tile_X3Y1_LUT4AB/W2BEG[5] Tile_X3Y1_LUT4AB/W2BEG[6] Tile_X3Y1_LUT4AB/W2BEG[7]
+ Tile_X2Y1_LUT4AB/W6BEG[0] Tile_X2Y1_LUT4AB/W6BEG[10] Tile_X2Y1_LUT4AB/W6BEG[11]
+ Tile_X2Y1_LUT4AB/W6BEG[1] Tile_X2Y1_LUT4AB/W6BEG[2] Tile_X2Y1_LUT4AB/W6BEG[3] Tile_X2Y1_LUT4AB/W6BEG[4]
+ Tile_X2Y1_LUT4AB/W6BEG[5] Tile_X2Y1_LUT4AB/W6BEG[6] Tile_X2Y1_LUT4AB/W6BEG[7] Tile_X2Y1_LUT4AB/W6BEG[8]
+ Tile_X2Y1_LUT4AB/W6BEG[9] Tile_X3Y1_LUT4AB/W6BEG[0] Tile_X3Y1_LUT4AB/W6BEG[10] Tile_X3Y1_LUT4AB/W6BEG[11]
+ Tile_X3Y1_LUT4AB/W6BEG[1] Tile_X3Y1_LUT4AB/W6BEG[2] Tile_X3Y1_LUT4AB/W6BEG[3] Tile_X3Y1_LUT4AB/W6BEG[4]
+ Tile_X3Y1_LUT4AB/W6BEG[5] Tile_X3Y1_LUT4AB/W6BEG[6] Tile_X3Y1_LUT4AB/W6BEG[7] Tile_X3Y1_LUT4AB/W6BEG[8]
+ Tile_X3Y1_LUT4AB/W6BEG[9] Tile_X2Y1_LUT4AB/WW4BEG[0] Tile_X2Y1_LUT4AB/WW4BEG[10]
+ Tile_X2Y1_LUT4AB/WW4BEG[11] Tile_X2Y1_LUT4AB/WW4BEG[12] Tile_X2Y1_LUT4AB/WW4BEG[13]
+ Tile_X2Y1_LUT4AB/WW4BEG[14] Tile_X2Y1_LUT4AB/WW4BEG[15] Tile_X2Y1_LUT4AB/WW4BEG[1]
+ Tile_X2Y1_LUT4AB/WW4BEG[2] Tile_X2Y1_LUT4AB/WW4BEG[3] Tile_X2Y1_LUT4AB/WW4BEG[4]
+ Tile_X2Y1_LUT4AB/WW4BEG[5] Tile_X2Y1_LUT4AB/WW4BEG[6] Tile_X2Y1_LUT4AB/WW4BEG[7]
+ Tile_X2Y1_LUT4AB/WW4BEG[8] Tile_X2Y1_LUT4AB/WW4BEG[9] Tile_X3Y1_LUT4AB/WW4BEG[0]
+ Tile_X3Y1_LUT4AB/WW4BEG[10] Tile_X3Y1_LUT4AB/WW4BEG[11] Tile_X3Y1_LUT4AB/WW4BEG[12]
+ Tile_X3Y1_LUT4AB/WW4BEG[13] Tile_X3Y1_LUT4AB/WW4BEG[14] Tile_X3Y1_LUT4AB/WW4BEG[15]
+ Tile_X3Y1_LUT4AB/WW4BEG[1] Tile_X3Y1_LUT4AB/WW4BEG[2] Tile_X3Y1_LUT4AB/WW4BEG[3]
+ Tile_X3Y1_LUT4AB/WW4BEG[4] Tile_X3Y1_LUT4AB/WW4BEG[5] Tile_X3Y1_LUT4AB/WW4BEG[6]
+ Tile_X3Y1_LUT4AB/WW4BEG[7] Tile_X3Y1_LUT4AB/WW4BEG[8] Tile_X3Y1_LUT4AB/WW4BEG[9]
+ LUT4AB
XTile_X0Y3_W_IO Tile_X0Y3_A_I_top Tile_X0Y3_A_O_top Tile_X0Y3_A_T_top Tile_X0Y3_A_config_C_bit0
+ Tile_X0Y3_A_config_C_bit1 Tile_X0Y3_A_config_C_bit2 Tile_X0Y3_A_config_C_bit3 Tile_X0Y3_B_I_top
+ Tile_X0Y3_B_O_top Tile_X0Y3_B_T_top Tile_X0Y3_B_config_C_bit0 Tile_X0Y3_B_config_C_bit1
+ Tile_X0Y3_B_config_C_bit2 Tile_X0Y3_B_config_C_bit3 Tile_X0Y3_W_IO/E1BEG[0] Tile_X0Y3_W_IO/E1BEG[1]
+ Tile_X0Y3_W_IO/E1BEG[2] Tile_X0Y3_W_IO/E1BEG[3] Tile_X0Y3_W_IO/E2BEG[0] Tile_X0Y3_W_IO/E2BEG[1]
+ Tile_X0Y3_W_IO/E2BEG[2] Tile_X0Y3_W_IO/E2BEG[3] Tile_X0Y3_W_IO/E2BEG[4] Tile_X0Y3_W_IO/E2BEG[5]
+ Tile_X0Y3_W_IO/E2BEG[6] Tile_X0Y3_W_IO/E2BEG[7] Tile_X0Y3_W_IO/E2BEGb[0] Tile_X0Y3_W_IO/E2BEGb[1]
+ Tile_X0Y3_W_IO/E2BEGb[2] Tile_X0Y3_W_IO/E2BEGb[3] Tile_X0Y3_W_IO/E2BEGb[4] Tile_X0Y3_W_IO/E2BEGb[5]
+ Tile_X0Y3_W_IO/E2BEGb[6] Tile_X0Y3_W_IO/E2BEGb[7] Tile_X0Y3_W_IO/E6BEG[0] Tile_X0Y3_W_IO/E6BEG[10]
+ Tile_X0Y3_W_IO/E6BEG[11] Tile_X0Y3_W_IO/E6BEG[1] Tile_X0Y3_W_IO/E6BEG[2] Tile_X0Y3_W_IO/E6BEG[3]
+ Tile_X0Y3_W_IO/E6BEG[4] Tile_X0Y3_W_IO/E6BEG[5] Tile_X0Y3_W_IO/E6BEG[6] Tile_X0Y3_W_IO/E6BEG[7]
+ Tile_X0Y3_W_IO/E6BEG[8] Tile_X0Y3_W_IO/E6BEG[9] Tile_X0Y3_W_IO/EE4BEG[0] Tile_X0Y3_W_IO/EE4BEG[10]
+ Tile_X0Y3_W_IO/EE4BEG[11] Tile_X0Y3_W_IO/EE4BEG[12] Tile_X0Y3_W_IO/EE4BEG[13] Tile_X0Y3_W_IO/EE4BEG[14]
+ Tile_X0Y3_W_IO/EE4BEG[15] Tile_X0Y3_W_IO/EE4BEG[1] Tile_X0Y3_W_IO/EE4BEG[2] Tile_X0Y3_W_IO/EE4BEG[3]
+ Tile_X0Y3_W_IO/EE4BEG[4] Tile_X0Y3_W_IO/EE4BEG[5] Tile_X0Y3_W_IO/EE4BEG[6] Tile_X0Y3_W_IO/EE4BEG[7]
+ Tile_X0Y3_W_IO/EE4BEG[8] Tile_X0Y3_W_IO/EE4BEG[9] FrameData[96] FrameData[106] FrameData[107]
+ FrameData[108] FrameData[109] FrameData[110] FrameData[111] FrameData[112] FrameData[113]
+ FrameData[114] FrameData[115] FrameData[97] FrameData[116] FrameData[117] FrameData[118]
+ FrameData[119] FrameData[120] FrameData[121] FrameData[122] FrameData[123] FrameData[124]
+ FrameData[125] FrameData[98] FrameData[126] FrameData[127] FrameData[99] FrameData[100]
+ FrameData[101] FrameData[102] FrameData[103] FrameData[104] FrameData[105] Tile_X1Y3_LUT4AB/FrameData[0]
+ Tile_X1Y3_LUT4AB/FrameData[10] Tile_X1Y3_LUT4AB/FrameData[11] Tile_X1Y3_LUT4AB/FrameData[12]
+ Tile_X1Y3_LUT4AB/FrameData[13] Tile_X1Y3_LUT4AB/FrameData[14] Tile_X1Y3_LUT4AB/FrameData[15]
+ Tile_X1Y3_LUT4AB/FrameData[16] Tile_X1Y3_LUT4AB/FrameData[17] Tile_X1Y3_LUT4AB/FrameData[18]
+ Tile_X1Y3_LUT4AB/FrameData[19] Tile_X1Y3_LUT4AB/FrameData[1] Tile_X1Y3_LUT4AB/FrameData[20]
+ Tile_X1Y3_LUT4AB/FrameData[21] Tile_X1Y3_LUT4AB/FrameData[22] Tile_X1Y3_LUT4AB/FrameData[23]
+ Tile_X1Y3_LUT4AB/FrameData[24] Tile_X1Y3_LUT4AB/FrameData[25] Tile_X1Y3_LUT4AB/FrameData[26]
+ Tile_X1Y3_LUT4AB/FrameData[27] Tile_X1Y3_LUT4AB/FrameData[28] Tile_X1Y3_LUT4AB/FrameData[29]
+ Tile_X1Y3_LUT4AB/FrameData[2] Tile_X1Y3_LUT4AB/FrameData[30] Tile_X1Y3_LUT4AB/FrameData[31]
+ Tile_X1Y3_LUT4AB/FrameData[3] Tile_X1Y3_LUT4AB/FrameData[4] Tile_X1Y3_LUT4AB/FrameData[5]
+ Tile_X1Y3_LUT4AB/FrameData[6] Tile_X1Y3_LUT4AB/FrameData[7] Tile_X1Y3_LUT4AB/FrameData[8]
+ Tile_X1Y3_LUT4AB/FrameData[9] Tile_X0Y3_W_IO/FrameStrobe[0] Tile_X0Y3_W_IO/FrameStrobe[10]
+ Tile_X0Y3_W_IO/FrameStrobe[11] Tile_X0Y3_W_IO/FrameStrobe[12] Tile_X0Y3_W_IO/FrameStrobe[13]
+ Tile_X0Y3_W_IO/FrameStrobe[14] Tile_X0Y3_W_IO/FrameStrobe[15] Tile_X0Y3_W_IO/FrameStrobe[16]
+ Tile_X0Y3_W_IO/FrameStrobe[17] Tile_X0Y3_W_IO/FrameStrobe[18] Tile_X0Y3_W_IO/FrameStrobe[19]
+ Tile_X0Y3_W_IO/FrameStrobe[1] Tile_X0Y3_W_IO/FrameStrobe[2] Tile_X0Y3_W_IO/FrameStrobe[3]
+ Tile_X0Y3_W_IO/FrameStrobe[4] Tile_X0Y3_W_IO/FrameStrobe[5] Tile_X0Y3_W_IO/FrameStrobe[6]
+ Tile_X0Y3_W_IO/FrameStrobe[7] Tile_X0Y3_W_IO/FrameStrobe[8] Tile_X0Y3_W_IO/FrameStrobe[9]
+ Tile_X0Y2_W_IO/FrameStrobe[0] Tile_X0Y2_W_IO/FrameStrobe[10] Tile_X0Y2_W_IO/FrameStrobe[11]
+ Tile_X0Y2_W_IO/FrameStrobe[12] Tile_X0Y2_W_IO/FrameStrobe[13] Tile_X0Y2_W_IO/FrameStrobe[14]
+ Tile_X0Y2_W_IO/FrameStrobe[15] Tile_X0Y2_W_IO/FrameStrobe[16] Tile_X0Y2_W_IO/FrameStrobe[17]
+ Tile_X0Y2_W_IO/FrameStrobe[18] Tile_X0Y2_W_IO/FrameStrobe[19] Tile_X0Y2_W_IO/FrameStrobe[1]
+ Tile_X0Y2_W_IO/FrameStrobe[2] Tile_X0Y2_W_IO/FrameStrobe[3] Tile_X0Y2_W_IO/FrameStrobe[4]
+ Tile_X0Y2_W_IO/FrameStrobe[5] Tile_X0Y2_W_IO/FrameStrobe[6] Tile_X0Y2_W_IO/FrameStrobe[7]
+ Tile_X0Y2_W_IO/FrameStrobe[8] Tile_X0Y2_W_IO/FrameStrobe[9] Tile_X0Y3_W_IO/UserCLK
+ Tile_X0Y2_W_IO/UserCLK VGND VPWR Tile_X0Y3_W_IO/W1END[0] Tile_X0Y3_W_IO/W1END[1]
+ Tile_X0Y3_W_IO/W1END[2] Tile_X0Y3_W_IO/W1END[3] Tile_X0Y3_W_IO/W2END[0] Tile_X0Y3_W_IO/W2END[1]
+ Tile_X0Y3_W_IO/W2END[2] Tile_X0Y3_W_IO/W2END[3] Tile_X0Y3_W_IO/W2END[4] Tile_X0Y3_W_IO/W2END[5]
+ Tile_X0Y3_W_IO/W2END[6] Tile_X0Y3_W_IO/W2END[7] Tile_X0Y3_W_IO/W2MID[0] Tile_X0Y3_W_IO/W2MID[1]
+ Tile_X0Y3_W_IO/W2MID[2] Tile_X0Y3_W_IO/W2MID[3] Tile_X0Y3_W_IO/W2MID[4] Tile_X0Y3_W_IO/W2MID[5]
+ Tile_X0Y3_W_IO/W2MID[6] Tile_X0Y3_W_IO/W2MID[7] Tile_X0Y3_W_IO/W6END[0] Tile_X0Y3_W_IO/W6END[10]
+ Tile_X0Y3_W_IO/W6END[11] Tile_X0Y3_W_IO/W6END[1] Tile_X0Y3_W_IO/W6END[2] Tile_X0Y3_W_IO/W6END[3]
+ Tile_X0Y3_W_IO/W6END[4] Tile_X0Y3_W_IO/W6END[5] Tile_X0Y3_W_IO/W6END[6] Tile_X0Y3_W_IO/W6END[7]
+ Tile_X0Y3_W_IO/W6END[8] Tile_X0Y3_W_IO/W6END[9] Tile_X0Y3_W_IO/WW4END[0] Tile_X0Y3_W_IO/WW4END[10]
+ Tile_X0Y3_W_IO/WW4END[11] Tile_X0Y3_W_IO/WW4END[12] Tile_X0Y3_W_IO/WW4END[13] Tile_X0Y3_W_IO/WW4END[14]
+ Tile_X0Y3_W_IO/WW4END[15] Tile_X0Y3_W_IO/WW4END[1] Tile_X0Y3_W_IO/WW4END[2] Tile_X0Y3_W_IO/WW4END[3]
+ Tile_X0Y3_W_IO/WW4END[4] Tile_X0Y3_W_IO/WW4END[5] Tile_X0Y3_W_IO/WW4END[6] Tile_X0Y3_W_IO/WW4END[7]
+ Tile_X0Y3_W_IO/WW4END[8] Tile_X0Y3_W_IO/WW4END[9] W_IO
XTile_X6Y14_LUT4AB Tile_X6Y14_LUT4AB/Ci Tile_X6Y14_LUT4AB/Co Tile_X6Y14_LUT4AB/E1BEG[0]
+ Tile_X6Y14_LUT4AB/E1BEG[1] Tile_X6Y14_LUT4AB/E1BEG[2] Tile_X6Y14_LUT4AB/E1BEG[3]
+ Tile_X6Y14_LUT4AB/E1END[0] Tile_X6Y14_LUT4AB/E1END[1] Tile_X6Y14_LUT4AB/E1END[2]
+ Tile_X6Y14_LUT4AB/E1END[3] Tile_X6Y14_LUT4AB/E2BEG[0] Tile_X6Y14_LUT4AB/E2BEG[1]
+ Tile_X6Y14_LUT4AB/E2BEG[2] Tile_X6Y14_LUT4AB/E2BEG[3] Tile_X6Y14_LUT4AB/E2BEG[4]
+ Tile_X6Y14_LUT4AB/E2BEG[5] Tile_X6Y14_LUT4AB/E2BEG[6] Tile_X6Y14_LUT4AB/E2BEG[7]
+ Tile_X6Y14_LUT4AB/E2BEGb[0] Tile_X6Y14_LUT4AB/E2BEGb[1] Tile_X6Y14_LUT4AB/E2BEGb[2]
+ Tile_X6Y14_LUT4AB/E2BEGb[3] Tile_X6Y14_LUT4AB/E2BEGb[4] Tile_X6Y14_LUT4AB/E2BEGb[5]
+ Tile_X6Y14_LUT4AB/E2BEGb[6] Tile_X6Y14_LUT4AB/E2BEGb[7] Tile_X6Y14_LUT4AB/E2END[0]
+ Tile_X6Y14_LUT4AB/E2END[1] Tile_X6Y14_LUT4AB/E2END[2] Tile_X6Y14_LUT4AB/E2END[3]
+ Tile_X6Y14_LUT4AB/E2END[4] Tile_X6Y14_LUT4AB/E2END[5] Tile_X6Y14_LUT4AB/E2END[6]
+ Tile_X6Y14_LUT4AB/E2END[7] Tile_X6Y14_LUT4AB/E2MID[0] Tile_X6Y14_LUT4AB/E2MID[1]
+ Tile_X6Y14_LUT4AB/E2MID[2] Tile_X6Y14_LUT4AB/E2MID[3] Tile_X6Y14_LUT4AB/E2MID[4]
+ Tile_X6Y14_LUT4AB/E2MID[5] Tile_X6Y14_LUT4AB/E2MID[6] Tile_X6Y14_LUT4AB/E2MID[7]
+ Tile_X6Y14_LUT4AB/E6BEG[0] Tile_X6Y14_LUT4AB/E6BEG[10] Tile_X6Y14_LUT4AB/E6BEG[11]
+ Tile_X6Y14_LUT4AB/E6BEG[1] Tile_X6Y14_LUT4AB/E6BEG[2] Tile_X6Y14_LUT4AB/E6BEG[3]
+ Tile_X6Y14_LUT4AB/E6BEG[4] Tile_X6Y14_LUT4AB/E6BEG[5] Tile_X6Y14_LUT4AB/E6BEG[6]
+ Tile_X6Y14_LUT4AB/E6BEG[7] Tile_X6Y14_LUT4AB/E6BEG[8] Tile_X6Y14_LUT4AB/E6BEG[9]
+ Tile_X6Y14_LUT4AB/E6END[0] Tile_X6Y14_LUT4AB/E6END[10] Tile_X6Y14_LUT4AB/E6END[11]
+ Tile_X6Y14_LUT4AB/E6END[1] Tile_X6Y14_LUT4AB/E6END[2] Tile_X6Y14_LUT4AB/E6END[3]
+ Tile_X6Y14_LUT4AB/E6END[4] Tile_X6Y14_LUT4AB/E6END[5] Tile_X6Y14_LUT4AB/E6END[6]
+ Tile_X6Y14_LUT4AB/E6END[7] Tile_X6Y14_LUT4AB/E6END[8] Tile_X6Y14_LUT4AB/E6END[9]
+ Tile_X6Y14_LUT4AB/EE4BEG[0] Tile_X6Y14_LUT4AB/EE4BEG[10] Tile_X6Y14_LUT4AB/EE4BEG[11]
+ Tile_X6Y14_LUT4AB/EE4BEG[12] Tile_X6Y14_LUT4AB/EE4BEG[13] Tile_X6Y14_LUT4AB/EE4BEG[14]
+ Tile_X6Y14_LUT4AB/EE4BEG[15] Tile_X6Y14_LUT4AB/EE4BEG[1] Tile_X6Y14_LUT4AB/EE4BEG[2]
+ Tile_X6Y14_LUT4AB/EE4BEG[3] Tile_X6Y14_LUT4AB/EE4BEG[4] Tile_X6Y14_LUT4AB/EE4BEG[5]
+ Tile_X6Y14_LUT4AB/EE4BEG[6] Tile_X6Y14_LUT4AB/EE4BEG[7] Tile_X6Y14_LUT4AB/EE4BEG[8]
+ Tile_X6Y14_LUT4AB/EE4BEG[9] Tile_X6Y14_LUT4AB/EE4END[0] Tile_X6Y14_LUT4AB/EE4END[10]
+ Tile_X6Y14_LUT4AB/EE4END[11] Tile_X6Y14_LUT4AB/EE4END[12] Tile_X6Y14_LUT4AB/EE4END[13]
+ Tile_X6Y14_LUT4AB/EE4END[14] Tile_X6Y14_LUT4AB/EE4END[15] Tile_X6Y14_LUT4AB/EE4END[1]
+ Tile_X6Y14_LUT4AB/EE4END[2] Tile_X6Y14_LUT4AB/EE4END[3] Tile_X6Y14_LUT4AB/EE4END[4]
+ Tile_X6Y14_LUT4AB/EE4END[5] Tile_X6Y14_LUT4AB/EE4END[6] Tile_X6Y14_LUT4AB/EE4END[7]
+ Tile_X6Y14_LUT4AB/EE4END[8] Tile_X6Y14_LUT4AB/EE4END[9] Tile_X6Y14_LUT4AB/FrameData[0]
+ Tile_X6Y14_LUT4AB/FrameData[10] Tile_X6Y14_LUT4AB/FrameData[11] Tile_X6Y14_LUT4AB/FrameData[12]
+ Tile_X6Y14_LUT4AB/FrameData[13] Tile_X6Y14_LUT4AB/FrameData[14] Tile_X6Y14_LUT4AB/FrameData[15]
+ Tile_X6Y14_LUT4AB/FrameData[16] Tile_X6Y14_LUT4AB/FrameData[17] Tile_X6Y14_LUT4AB/FrameData[18]
+ Tile_X6Y14_LUT4AB/FrameData[19] Tile_X6Y14_LUT4AB/FrameData[1] Tile_X6Y14_LUT4AB/FrameData[20]
+ Tile_X6Y14_LUT4AB/FrameData[21] Tile_X6Y14_LUT4AB/FrameData[22] Tile_X6Y14_LUT4AB/FrameData[23]
+ Tile_X6Y14_LUT4AB/FrameData[24] Tile_X6Y14_LUT4AB/FrameData[25] Tile_X6Y14_LUT4AB/FrameData[26]
+ Tile_X6Y14_LUT4AB/FrameData[27] Tile_X6Y14_LUT4AB/FrameData[28] Tile_X6Y14_LUT4AB/FrameData[29]
+ Tile_X6Y14_LUT4AB/FrameData[2] Tile_X6Y14_LUT4AB/FrameData[30] Tile_X6Y14_LUT4AB/FrameData[31]
+ Tile_X6Y14_LUT4AB/FrameData[3] Tile_X6Y14_LUT4AB/FrameData[4] Tile_X6Y14_LUT4AB/FrameData[5]
+ Tile_X6Y14_LUT4AB/FrameData[6] Tile_X6Y14_LUT4AB/FrameData[7] Tile_X6Y14_LUT4AB/FrameData[8]
+ Tile_X6Y14_LUT4AB/FrameData[9] Tile_X6Y14_LUT4AB/FrameData_O[0] Tile_X6Y14_LUT4AB/FrameData_O[10]
+ Tile_X6Y14_LUT4AB/FrameData_O[11] Tile_X6Y14_LUT4AB/FrameData_O[12] Tile_X6Y14_LUT4AB/FrameData_O[13]
+ Tile_X6Y14_LUT4AB/FrameData_O[14] Tile_X6Y14_LUT4AB/FrameData_O[15] Tile_X6Y14_LUT4AB/FrameData_O[16]
+ Tile_X6Y14_LUT4AB/FrameData_O[17] Tile_X6Y14_LUT4AB/FrameData_O[18] Tile_X6Y14_LUT4AB/FrameData_O[19]
+ Tile_X6Y14_LUT4AB/FrameData_O[1] Tile_X6Y14_LUT4AB/FrameData_O[20] Tile_X6Y14_LUT4AB/FrameData_O[21]
+ Tile_X6Y14_LUT4AB/FrameData_O[22] Tile_X6Y14_LUT4AB/FrameData_O[23] Tile_X6Y14_LUT4AB/FrameData_O[24]
+ Tile_X6Y14_LUT4AB/FrameData_O[25] Tile_X6Y14_LUT4AB/FrameData_O[26] Tile_X6Y14_LUT4AB/FrameData_O[27]
+ Tile_X6Y14_LUT4AB/FrameData_O[28] Tile_X6Y14_LUT4AB/FrameData_O[29] Tile_X6Y14_LUT4AB/FrameData_O[2]
+ Tile_X6Y14_LUT4AB/FrameData_O[30] Tile_X6Y14_LUT4AB/FrameData_O[31] Tile_X6Y14_LUT4AB/FrameData_O[3]
+ Tile_X6Y14_LUT4AB/FrameData_O[4] Tile_X6Y14_LUT4AB/FrameData_O[5] Tile_X6Y14_LUT4AB/FrameData_O[6]
+ Tile_X6Y14_LUT4AB/FrameData_O[7] Tile_X6Y14_LUT4AB/FrameData_O[8] Tile_X6Y14_LUT4AB/FrameData_O[9]
+ Tile_X6Y14_LUT4AB/FrameStrobe[0] Tile_X6Y14_LUT4AB/FrameStrobe[10] Tile_X6Y14_LUT4AB/FrameStrobe[11]
+ Tile_X6Y14_LUT4AB/FrameStrobe[12] Tile_X6Y14_LUT4AB/FrameStrobe[13] Tile_X6Y14_LUT4AB/FrameStrobe[14]
+ Tile_X6Y14_LUT4AB/FrameStrobe[15] Tile_X6Y14_LUT4AB/FrameStrobe[16] Tile_X6Y14_LUT4AB/FrameStrobe[17]
+ Tile_X6Y14_LUT4AB/FrameStrobe[18] Tile_X6Y14_LUT4AB/FrameStrobe[19] Tile_X6Y14_LUT4AB/FrameStrobe[1]
+ Tile_X6Y14_LUT4AB/FrameStrobe[2] Tile_X6Y14_LUT4AB/FrameStrobe[3] Tile_X6Y14_LUT4AB/FrameStrobe[4]
+ Tile_X6Y14_LUT4AB/FrameStrobe[5] Tile_X6Y14_LUT4AB/FrameStrobe[6] Tile_X6Y14_LUT4AB/FrameStrobe[7]
+ Tile_X6Y14_LUT4AB/FrameStrobe[8] Tile_X6Y14_LUT4AB/FrameStrobe[9] Tile_X6Y13_LUT4AB/FrameStrobe[0]
+ Tile_X6Y13_LUT4AB/FrameStrobe[10] Tile_X6Y13_LUT4AB/FrameStrobe[11] Tile_X6Y13_LUT4AB/FrameStrobe[12]
+ Tile_X6Y13_LUT4AB/FrameStrobe[13] Tile_X6Y13_LUT4AB/FrameStrobe[14] Tile_X6Y13_LUT4AB/FrameStrobe[15]
+ Tile_X6Y13_LUT4AB/FrameStrobe[16] Tile_X6Y13_LUT4AB/FrameStrobe[17] Tile_X6Y13_LUT4AB/FrameStrobe[18]
+ Tile_X6Y13_LUT4AB/FrameStrobe[19] Tile_X6Y13_LUT4AB/FrameStrobe[1] Tile_X6Y13_LUT4AB/FrameStrobe[2]
+ Tile_X6Y13_LUT4AB/FrameStrobe[3] Tile_X6Y13_LUT4AB/FrameStrobe[4] Tile_X6Y13_LUT4AB/FrameStrobe[5]
+ Tile_X6Y13_LUT4AB/FrameStrobe[6] Tile_X6Y13_LUT4AB/FrameStrobe[7] Tile_X6Y13_LUT4AB/FrameStrobe[8]
+ Tile_X6Y13_LUT4AB/FrameStrobe[9] Tile_X6Y14_LUT4AB/N1BEG[0] Tile_X6Y14_LUT4AB/N1BEG[1]
+ Tile_X6Y14_LUT4AB/N1BEG[2] Tile_X6Y14_LUT4AB/N1BEG[3] Tile_X6Y14_LUT4AB/N1END[0]
+ Tile_X6Y14_LUT4AB/N1END[1] Tile_X6Y14_LUT4AB/N1END[2] Tile_X6Y14_LUT4AB/N1END[3]
+ Tile_X6Y14_LUT4AB/N2BEG[0] Tile_X6Y14_LUT4AB/N2BEG[1] Tile_X6Y14_LUT4AB/N2BEG[2]
+ Tile_X6Y14_LUT4AB/N2BEG[3] Tile_X6Y14_LUT4AB/N2BEG[4] Tile_X6Y14_LUT4AB/N2BEG[5]
+ Tile_X6Y14_LUT4AB/N2BEG[6] Tile_X6Y14_LUT4AB/N2BEG[7] Tile_X6Y13_LUT4AB/N2END[0]
+ Tile_X6Y13_LUT4AB/N2END[1] Tile_X6Y13_LUT4AB/N2END[2] Tile_X6Y13_LUT4AB/N2END[3]
+ Tile_X6Y13_LUT4AB/N2END[4] Tile_X6Y13_LUT4AB/N2END[5] Tile_X6Y13_LUT4AB/N2END[6]
+ Tile_X6Y13_LUT4AB/N2END[7] Tile_X6Y14_LUT4AB/N2END[0] Tile_X6Y14_LUT4AB/N2END[1]
+ Tile_X6Y14_LUT4AB/N2END[2] Tile_X6Y14_LUT4AB/N2END[3] Tile_X6Y14_LUT4AB/N2END[4]
+ Tile_X6Y14_LUT4AB/N2END[5] Tile_X6Y14_LUT4AB/N2END[6] Tile_X6Y14_LUT4AB/N2END[7]
+ Tile_X6Y14_LUT4AB/N2MID[0] Tile_X6Y14_LUT4AB/N2MID[1] Tile_X6Y14_LUT4AB/N2MID[2]
+ Tile_X6Y14_LUT4AB/N2MID[3] Tile_X6Y14_LUT4AB/N2MID[4] Tile_X6Y14_LUT4AB/N2MID[5]
+ Tile_X6Y14_LUT4AB/N2MID[6] Tile_X6Y14_LUT4AB/N2MID[7] Tile_X6Y14_LUT4AB/N4BEG[0]
+ Tile_X6Y14_LUT4AB/N4BEG[10] Tile_X6Y14_LUT4AB/N4BEG[11] Tile_X6Y14_LUT4AB/N4BEG[12]
+ Tile_X6Y14_LUT4AB/N4BEG[13] Tile_X6Y14_LUT4AB/N4BEG[14] Tile_X6Y14_LUT4AB/N4BEG[15]
+ Tile_X6Y14_LUT4AB/N4BEG[1] Tile_X6Y14_LUT4AB/N4BEG[2] Tile_X6Y14_LUT4AB/N4BEG[3]
+ Tile_X6Y14_LUT4AB/N4BEG[4] Tile_X6Y14_LUT4AB/N4BEG[5] Tile_X6Y14_LUT4AB/N4BEG[6]
+ Tile_X6Y14_LUT4AB/N4BEG[7] Tile_X6Y14_LUT4AB/N4BEG[8] Tile_X6Y14_LUT4AB/N4BEG[9]
+ Tile_X6Y14_LUT4AB/N4END[0] Tile_X6Y14_LUT4AB/N4END[10] Tile_X6Y14_LUT4AB/N4END[11]
+ Tile_X6Y14_LUT4AB/N4END[12] Tile_X6Y14_LUT4AB/N4END[13] Tile_X6Y14_LUT4AB/N4END[14]
+ Tile_X6Y14_LUT4AB/N4END[15] Tile_X6Y14_LUT4AB/N4END[1] Tile_X6Y14_LUT4AB/N4END[2]
+ Tile_X6Y14_LUT4AB/N4END[3] Tile_X6Y14_LUT4AB/N4END[4] Tile_X6Y14_LUT4AB/N4END[5]
+ Tile_X6Y14_LUT4AB/N4END[6] Tile_X6Y14_LUT4AB/N4END[7] Tile_X6Y14_LUT4AB/N4END[8]
+ Tile_X6Y14_LUT4AB/N4END[9] Tile_X6Y14_LUT4AB/NN4BEG[0] Tile_X6Y14_LUT4AB/NN4BEG[10]
+ Tile_X6Y14_LUT4AB/NN4BEG[11] Tile_X6Y14_LUT4AB/NN4BEG[12] Tile_X6Y14_LUT4AB/NN4BEG[13]
+ Tile_X6Y14_LUT4AB/NN4BEG[14] Tile_X6Y14_LUT4AB/NN4BEG[15] Tile_X6Y14_LUT4AB/NN4BEG[1]
+ Tile_X6Y14_LUT4AB/NN4BEG[2] Tile_X6Y14_LUT4AB/NN4BEG[3] Tile_X6Y14_LUT4AB/NN4BEG[4]
+ Tile_X6Y14_LUT4AB/NN4BEG[5] Tile_X6Y14_LUT4AB/NN4BEG[6] Tile_X6Y14_LUT4AB/NN4BEG[7]
+ Tile_X6Y14_LUT4AB/NN4BEG[8] Tile_X6Y14_LUT4AB/NN4BEG[9] Tile_X6Y14_LUT4AB/NN4END[0]
+ Tile_X6Y14_LUT4AB/NN4END[10] Tile_X6Y14_LUT4AB/NN4END[11] Tile_X6Y14_LUT4AB/NN4END[12]
+ Tile_X6Y14_LUT4AB/NN4END[13] Tile_X6Y14_LUT4AB/NN4END[14] Tile_X6Y14_LUT4AB/NN4END[15]
+ Tile_X6Y14_LUT4AB/NN4END[1] Tile_X6Y14_LUT4AB/NN4END[2] Tile_X6Y14_LUT4AB/NN4END[3]
+ Tile_X6Y14_LUT4AB/NN4END[4] Tile_X6Y14_LUT4AB/NN4END[5] Tile_X6Y14_LUT4AB/NN4END[6]
+ Tile_X6Y14_LUT4AB/NN4END[7] Tile_X6Y14_LUT4AB/NN4END[8] Tile_X6Y14_LUT4AB/NN4END[9]
+ Tile_X6Y14_LUT4AB/S1BEG[0] Tile_X6Y14_LUT4AB/S1BEG[1] Tile_X6Y14_LUT4AB/S1BEG[2]
+ Tile_X6Y14_LUT4AB/S1BEG[3] Tile_X6Y14_LUT4AB/S1END[0] Tile_X6Y14_LUT4AB/S1END[1]
+ Tile_X6Y14_LUT4AB/S1END[2] Tile_X6Y14_LUT4AB/S1END[3] Tile_X6Y14_LUT4AB/S2BEG[0]
+ Tile_X6Y14_LUT4AB/S2BEG[1] Tile_X6Y14_LUT4AB/S2BEG[2] Tile_X6Y14_LUT4AB/S2BEG[3]
+ Tile_X6Y14_LUT4AB/S2BEG[4] Tile_X6Y14_LUT4AB/S2BEG[5] Tile_X6Y14_LUT4AB/S2BEG[6]
+ Tile_X6Y14_LUT4AB/S2BEG[7] Tile_X6Y14_LUT4AB/S2BEGb[0] Tile_X6Y14_LUT4AB/S2BEGb[1]
+ Tile_X6Y14_LUT4AB/S2BEGb[2] Tile_X6Y14_LUT4AB/S2BEGb[3] Tile_X6Y14_LUT4AB/S2BEGb[4]
+ Tile_X6Y14_LUT4AB/S2BEGb[5] Tile_X6Y14_LUT4AB/S2BEGb[6] Tile_X6Y14_LUT4AB/S2BEGb[7]
+ Tile_X6Y14_LUT4AB/S2END[0] Tile_X6Y14_LUT4AB/S2END[1] Tile_X6Y14_LUT4AB/S2END[2]
+ Tile_X6Y14_LUT4AB/S2END[3] Tile_X6Y14_LUT4AB/S2END[4] Tile_X6Y14_LUT4AB/S2END[5]
+ Tile_X6Y14_LUT4AB/S2END[6] Tile_X6Y14_LUT4AB/S2END[7] Tile_X6Y14_LUT4AB/S2MID[0]
+ Tile_X6Y14_LUT4AB/S2MID[1] Tile_X6Y14_LUT4AB/S2MID[2] Tile_X6Y14_LUT4AB/S2MID[3]
+ Tile_X6Y14_LUT4AB/S2MID[4] Tile_X6Y14_LUT4AB/S2MID[5] Tile_X6Y14_LUT4AB/S2MID[6]
+ Tile_X6Y14_LUT4AB/S2MID[7] Tile_X6Y14_LUT4AB/S4BEG[0] Tile_X6Y14_LUT4AB/S4BEG[10]
+ Tile_X6Y14_LUT4AB/S4BEG[11] Tile_X6Y14_LUT4AB/S4BEG[12] Tile_X6Y14_LUT4AB/S4BEG[13]
+ Tile_X6Y14_LUT4AB/S4BEG[14] Tile_X6Y14_LUT4AB/S4BEG[15] Tile_X6Y14_LUT4AB/S4BEG[1]
+ Tile_X6Y14_LUT4AB/S4BEG[2] Tile_X6Y14_LUT4AB/S4BEG[3] Tile_X6Y14_LUT4AB/S4BEG[4]
+ Tile_X6Y14_LUT4AB/S4BEG[5] Tile_X6Y14_LUT4AB/S4BEG[6] Tile_X6Y14_LUT4AB/S4BEG[7]
+ Tile_X6Y14_LUT4AB/S4BEG[8] Tile_X6Y14_LUT4AB/S4BEG[9] Tile_X6Y14_LUT4AB/S4END[0]
+ Tile_X6Y14_LUT4AB/S4END[10] Tile_X6Y14_LUT4AB/S4END[11] Tile_X6Y14_LUT4AB/S4END[12]
+ Tile_X6Y14_LUT4AB/S4END[13] Tile_X6Y14_LUT4AB/S4END[14] Tile_X6Y14_LUT4AB/S4END[15]
+ Tile_X6Y14_LUT4AB/S4END[1] Tile_X6Y14_LUT4AB/S4END[2] Tile_X6Y14_LUT4AB/S4END[3]
+ Tile_X6Y14_LUT4AB/S4END[4] Tile_X6Y14_LUT4AB/S4END[5] Tile_X6Y14_LUT4AB/S4END[6]
+ Tile_X6Y14_LUT4AB/S4END[7] Tile_X6Y14_LUT4AB/S4END[8] Tile_X6Y14_LUT4AB/S4END[9]
+ Tile_X6Y14_LUT4AB/SS4BEG[0] Tile_X6Y14_LUT4AB/SS4BEG[10] Tile_X6Y14_LUT4AB/SS4BEG[11]
+ Tile_X6Y14_LUT4AB/SS4BEG[12] Tile_X6Y14_LUT4AB/SS4BEG[13] Tile_X6Y14_LUT4AB/SS4BEG[14]
+ Tile_X6Y14_LUT4AB/SS4BEG[15] Tile_X6Y14_LUT4AB/SS4BEG[1] Tile_X6Y14_LUT4AB/SS4BEG[2]
+ Tile_X6Y14_LUT4AB/SS4BEG[3] Tile_X6Y14_LUT4AB/SS4BEG[4] Tile_X6Y14_LUT4AB/SS4BEG[5]
+ Tile_X6Y14_LUT4AB/SS4BEG[6] Tile_X6Y14_LUT4AB/SS4BEG[7] Tile_X6Y14_LUT4AB/SS4BEG[8]
+ Tile_X6Y14_LUT4AB/SS4BEG[9] Tile_X6Y14_LUT4AB/SS4END[0] Tile_X6Y14_LUT4AB/SS4END[10]
+ Tile_X6Y14_LUT4AB/SS4END[11] Tile_X6Y14_LUT4AB/SS4END[12] Tile_X6Y14_LUT4AB/SS4END[13]
+ Tile_X6Y14_LUT4AB/SS4END[14] Tile_X6Y14_LUT4AB/SS4END[15] Tile_X6Y14_LUT4AB/SS4END[1]
+ Tile_X6Y14_LUT4AB/SS4END[2] Tile_X6Y14_LUT4AB/SS4END[3] Tile_X6Y14_LUT4AB/SS4END[4]
+ Tile_X6Y14_LUT4AB/SS4END[5] Tile_X6Y14_LUT4AB/SS4END[6] Tile_X6Y14_LUT4AB/SS4END[7]
+ Tile_X6Y14_LUT4AB/SS4END[8] Tile_X6Y14_LUT4AB/SS4END[9] Tile_X6Y14_LUT4AB/UserCLK
+ Tile_X6Y13_LUT4AB/UserCLK VGND VPWR Tile_X6Y14_LUT4AB/W1BEG[0] Tile_X6Y14_LUT4AB/W1BEG[1]
+ Tile_X6Y14_LUT4AB/W1BEG[2] Tile_X6Y14_LUT4AB/W1BEG[3] Tile_X6Y14_LUT4AB/W1END[0]
+ Tile_X6Y14_LUT4AB/W1END[1] Tile_X6Y14_LUT4AB/W1END[2] Tile_X6Y14_LUT4AB/W1END[3]
+ Tile_X6Y14_LUT4AB/W2BEG[0] Tile_X6Y14_LUT4AB/W2BEG[1] Tile_X6Y14_LUT4AB/W2BEG[2]
+ Tile_X6Y14_LUT4AB/W2BEG[3] Tile_X6Y14_LUT4AB/W2BEG[4] Tile_X6Y14_LUT4AB/W2BEG[5]
+ Tile_X6Y14_LUT4AB/W2BEG[6] Tile_X6Y14_LUT4AB/W2BEG[7] Tile_X5Y14_LUT4AB/W2END[0]
+ Tile_X5Y14_LUT4AB/W2END[1] Tile_X5Y14_LUT4AB/W2END[2] Tile_X5Y14_LUT4AB/W2END[3]
+ Tile_X5Y14_LUT4AB/W2END[4] Tile_X5Y14_LUT4AB/W2END[5] Tile_X5Y14_LUT4AB/W2END[6]
+ Tile_X5Y14_LUT4AB/W2END[7] Tile_X6Y14_LUT4AB/W2END[0] Tile_X6Y14_LUT4AB/W2END[1]
+ Tile_X6Y14_LUT4AB/W2END[2] Tile_X6Y14_LUT4AB/W2END[3] Tile_X6Y14_LUT4AB/W2END[4]
+ Tile_X6Y14_LUT4AB/W2END[5] Tile_X6Y14_LUT4AB/W2END[6] Tile_X6Y14_LUT4AB/W2END[7]
+ Tile_X6Y14_LUT4AB/W2MID[0] Tile_X6Y14_LUT4AB/W2MID[1] Tile_X6Y14_LUT4AB/W2MID[2]
+ Tile_X6Y14_LUT4AB/W2MID[3] Tile_X6Y14_LUT4AB/W2MID[4] Tile_X6Y14_LUT4AB/W2MID[5]
+ Tile_X6Y14_LUT4AB/W2MID[6] Tile_X6Y14_LUT4AB/W2MID[7] Tile_X6Y14_LUT4AB/W6BEG[0]
+ Tile_X6Y14_LUT4AB/W6BEG[10] Tile_X6Y14_LUT4AB/W6BEG[11] Tile_X6Y14_LUT4AB/W6BEG[1]
+ Tile_X6Y14_LUT4AB/W6BEG[2] Tile_X6Y14_LUT4AB/W6BEG[3] Tile_X6Y14_LUT4AB/W6BEG[4]
+ Tile_X6Y14_LUT4AB/W6BEG[5] Tile_X6Y14_LUT4AB/W6BEG[6] Tile_X6Y14_LUT4AB/W6BEG[7]
+ Tile_X6Y14_LUT4AB/W6BEG[8] Tile_X6Y14_LUT4AB/W6BEG[9] Tile_X6Y14_LUT4AB/W6END[0]
+ Tile_X6Y14_LUT4AB/W6END[10] Tile_X6Y14_LUT4AB/W6END[11] Tile_X6Y14_LUT4AB/W6END[1]
+ Tile_X6Y14_LUT4AB/W6END[2] Tile_X6Y14_LUT4AB/W6END[3] Tile_X6Y14_LUT4AB/W6END[4]
+ Tile_X6Y14_LUT4AB/W6END[5] Tile_X6Y14_LUT4AB/W6END[6] Tile_X6Y14_LUT4AB/W6END[7]
+ Tile_X6Y14_LUT4AB/W6END[8] Tile_X6Y14_LUT4AB/W6END[9] Tile_X6Y14_LUT4AB/WW4BEG[0]
+ Tile_X6Y14_LUT4AB/WW4BEG[10] Tile_X6Y14_LUT4AB/WW4BEG[11] Tile_X6Y14_LUT4AB/WW4BEG[12]
+ Tile_X6Y14_LUT4AB/WW4BEG[13] Tile_X6Y14_LUT4AB/WW4BEG[14] Tile_X6Y14_LUT4AB/WW4BEG[15]
+ Tile_X6Y14_LUT4AB/WW4BEG[1] Tile_X6Y14_LUT4AB/WW4BEG[2] Tile_X6Y14_LUT4AB/WW4BEG[3]
+ Tile_X6Y14_LUT4AB/WW4BEG[4] Tile_X6Y14_LUT4AB/WW4BEG[5] Tile_X6Y14_LUT4AB/WW4BEG[6]
+ Tile_X6Y14_LUT4AB/WW4BEG[7] Tile_X6Y14_LUT4AB/WW4BEG[8] Tile_X6Y14_LUT4AB/WW4BEG[9]
+ Tile_X6Y14_LUT4AB/WW4END[0] Tile_X6Y14_LUT4AB/WW4END[10] Tile_X6Y14_LUT4AB/WW4END[11]
+ Tile_X6Y14_LUT4AB/WW4END[12] Tile_X6Y14_LUT4AB/WW4END[13] Tile_X6Y14_LUT4AB/WW4END[14]
+ Tile_X6Y14_LUT4AB/WW4END[15] Tile_X6Y14_LUT4AB/WW4END[1] Tile_X6Y14_LUT4AB/WW4END[2]
+ Tile_X6Y14_LUT4AB/WW4END[3] Tile_X6Y14_LUT4AB/WW4END[4] Tile_X6Y14_LUT4AB/WW4END[5]
+ Tile_X6Y14_LUT4AB/WW4END[6] Tile_X6Y14_LUT4AB/WW4END[7] Tile_X6Y14_LUT4AB/WW4END[8]
+ Tile_X6Y14_LUT4AB/WW4END[9] LUT4AB
XTile_X1Y5_LUT4AB Tile_X1Y6_LUT4AB/Co Tile_X1Y5_LUT4AB/Co Tile_X2Y5_LUT4AB/E1END[0]
+ Tile_X2Y5_LUT4AB/E1END[1] Tile_X2Y5_LUT4AB/E1END[2] Tile_X2Y5_LUT4AB/E1END[3] Tile_X0Y5_W_IO/E1BEG[0]
+ Tile_X0Y5_W_IO/E1BEG[1] Tile_X0Y5_W_IO/E1BEG[2] Tile_X0Y5_W_IO/E1BEG[3] Tile_X2Y5_LUT4AB/E2MID[0]
+ Tile_X2Y5_LUT4AB/E2MID[1] Tile_X2Y5_LUT4AB/E2MID[2] Tile_X2Y5_LUT4AB/E2MID[3] Tile_X2Y5_LUT4AB/E2MID[4]
+ Tile_X2Y5_LUT4AB/E2MID[5] Tile_X2Y5_LUT4AB/E2MID[6] Tile_X2Y5_LUT4AB/E2MID[7] Tile_X2Y5_LUT4AB/E2END[0]
+ Tile_X2Y5_LUT4AB/E2END[1] Tile_X2Y5_LUT4AB/E2END[2] Tile_X2Y5_LUT4AB/E2END[3] Tile_X2Y5_LUT4AB/E2END[4]
+ Tile_X2Y5_LUT4AB/E2END[5] Tile_X2Y5_LUT4AB/E2END[6] Tile_X2Y5_LUT4AB/E2END[7] Tile_X0Y5_W_IO/E2BEGb[0]
+ Tile_X0Y5_W_IO/E2BEGb[1] Tile_X0Y5_W_IO/E2BEGb[2] Tile_X0Y5_W_IO/E2BEGb[3] Tile_X0Y5_W_IO/E2BEGb[4]
+ Tile_X0Y5_W_IO/E2BEGb[5] Tile_X0Y5_W_IO/E2BEGb[6] Tile_X0Y5_W_IO/E2BEGb[7] Tile_X0Y5_W_IO/E2BEG[0]
+ Tile_X0Y5_W_IO/E2BEG[1] Tile_X0Y5_W_IO/E2BEG[2] Tile_X0Y5_W_IO/E2BEG[3] Tile_X0Y5_W_IO/E2BEG[4]
+ Tile_X0Y5_W_IO/E2BEG[5] Tile_X0Y5_W_IO/E2BEG[6] Tile_X0Y5_W_IO/E2BEG[7] Tile_X2Y5_LUT4AB/E6END[0]
+ Tile_X2Y5_LUT4AB/E6END[10] Tile_X2Y5_LUT4AB/E6END[11] Tile_X2Y5_LUT4AB/E6END[1]
+ Tile_X2Y5_LUT4AB/E6END[2] Tile_X2Y5_LUT4AB/E6END[3] Tile_X2Y5_LUT4AB/E6END[4] Tile_X2Y5_LUT4AB/E6END[5]
+ Tile_X2Y5_LUT4AB/E6END[6] Tile_X2Y5_LUT4AB/E6END[7] Tile_X2Y5_LUT4AB/E6END[8] Tile_X2Y5_LUT4AB/E6END[9]
+ Tile_X0Y5_W_IO/E6BEG[0] Tile_X0Y5_W_IO/E6BEG[10] Tile_X0Y5_W_IO/E6BEG[11] Tile_X0Y5_W_IO/E6BEG[1]
+ Tile_X0Y5_W_IO/E6BEG[2] Tile_X0Y5_W_IO/E6BEG[3] Tile_X0Y5_W_IO/E6BEG[4] Tile_X0Y5_W_IO/E6BEG[5]
+ Tile_X0Y5_W_IO/E6BEG[6] Tile_X0Y5_W_IO/E6BEG[7] Tile_X0Y5_W_IO/E6BEG[8] Tile_X0Y5_W_IO/E6BEG[9]
+ Tile_X2Y5_LUT4AB/EE4END[0] Tile_X2Y5_LUT4AB/EE4END[10] Tile_X2Y5_LUT4AB/EE4END[11]
+ Tile_X2Y5_LUT4AB/EE4END[12] Tile_X2Y5_LUT4AB/EE4END[13] Tile_X2Y5_LUT4AB/EE4END[14]
+ Tile_X2Y5_LUT4AB/EE4END[15] Tile_X2Y5_LUT4AB/EE4END[1] Tile_X2Y5_LUT4AB/EE4END[2]
+ Tile_X2Y5_LUT4AB/EE4END[3] Tile_X2Y5_LUT4AB/EE4END[4] Tile_X2Y5_LUT4AB/EE4END[5]
+ Tile_X2Y5_LUT4AB/EE4END[6] Tile_X2Y5_LUT4AB/EE4END[7] Tile_X2Y5_LUT4AB/EE4END[8]
+ Tile_X2Y5_LUT4AB/EE4END[9] Tile_X0Y5_W_IO/EE4BEG[0] Tile_X0Y5_W_IO/EE4BEG[10] Tile_X0Y5_W_IO/EE4BEG[11]
+ Tile_X0Y5_W_IO/EE4BEG[12] Tile_X0Y5_W_IO/EE4BEG[13] Tile_X0Y5_W_IO/EE4BEG[14] Tile_X0Y5_W_IO/EE4BEG[15]
+ Tile_X0Y5_W_IO/EE4BEG[1] Tile_X0Y5_W_IO/EE4BEG[2] Tile_X0Y5_W_IO/EE4BEG[3] Tile_X0Y5_W_IO/EE4BEG[4]
+ Tile_X0Y5_W_IO/EE4BEG[5] Tile_X0Y5_W_IO/EE4BEG[6] Tile_X0Y5_W_IO/EE4BEG[7] Tile_X0Y5_W_IO/EE4BEG[8]
+ Tile_X0Y5_W_IO/EE4BEG[9] Tile_X1Y5_LUT4AB/FrameData[0] Tile_X1Y5_LUT4AB/FrameData[10]
+ Tile_X1Y5_LUT4AB/FrameData[11] Tile_X1Y5_LUT4AB/FrameData[12] Tile_X1Y5_LUT4AB/FrameData[13]
+ Tile_X1Y5_LUT4AB/FrameData[14] Tile_X1Y5_LUT4AB/FrameData[15] Tile_X1Y5_LUT4AB/FrameData[16]
+ Tile_X1Y5_LUT4AB/FrameData[17] Tile_X1Y5_LUT4AB/FrameData[18] Tile_X1Y5_LUT4AB/FrameData[19]
+ Tile_X1Y5_LUT4AB/FrameData[1] Tile_X1Y5_LUT4AB/FrameData[20] Tile_X1Y5_LUT4AB/FrameData[21]
+ Tile_X1Y5_LUT4AB/FrameData[22] Tile_X1Y5_LUT4AB/FrameData[23] Tile_X1Y5_LUT4AB/FrameData[24]
+ Tile_X1Y5_LUT4AB/FrameData[25] Tile_X1Y5_LUT4AB/FrameData[26] Tile_X1Y5_LUT4AB/FrameData[27]
+ Tile_X1Y5_LUT4AB/FrameData[28] Tile_X1Y5_LUT4AB/FrameData[29] Tile_X1Y5_LUT4AB/FrameData[2]
+ Tile_X1Y5_LUT4AB/FrameData[30] Tile_X1Y5_LUT4AB/FrameData[31] Tile_X1Y5_LUT4AB/FrameData[3]
+ Tile_X1Y5_LUT4AB/FrameData[4] Tile_X1Y5_LUT4AB/FrameData[5] Tile_X1Y5_LUT4AB/FrameData[6]
+ Tile_X1Y5_LUT4AB/FrameData[7] Tile_X1Y5_LUT4AB/FrameData[8] Tile_X1Y5_LUT4AB/FrameData[9]
+ Tile_X2Y5_LUT4AB/FrameData[0] Tile_X2Y5_LUT4AB/FrameData[10] Tile_X2Y5_LUT4AB/FrameData[11]
+ Tile_X2Y5_LUT4AB/FrameData[12] Tile_X2Y5_LUT4AB/FrameData[13] Tile_X2Y5_LUT4AB/FrameData[14]
+ Tile_X2Y5_LUT4AB/FrameData[15] Tile_X2Y5_LUT4AB/FrameData[16] Tile_X2Y5_LUT4AB/FrameData[17]
+ Tile_X2Y5_LUT4AB/FrameData[18] Tile_X2Y5_LUT4AB/FrameData[19] Tile_X2Y5_LUT4AB/FrameData[1]
+ Tile_X2Y5_LUT4AB/FrameData[20] Tile_X2Y5_LUT4AB/FrameData[21] Tile_X2Y5_LUT4AB/FrameData[22]
+ Tile_X2Y5_LUT4AB/FrameData[23] Tile_X2Y5_LUT4AB/FrameData[24] Tile_X2Y5_LUT4AB/FrameData[25]
+ Tile_X2Y5_LUT4AB/FrameData[26] Tile_X2Y5_LUT4AB/FrameData[27] Tile_X2Y5_LUT4AB/FrameData[28]
+ Tile_X2Y5_LUT4AB/FrameData[29] Tile_X2Y5_LUT4AB/FrameData[2] Tile_X2Y5_LUT4AB/FrameData[30]
+ Tile_X2Y5_LUT4AB/FrameData[31] Tile_X2Y5_LUT4AB/FrameData[3] Tile_X2Y5_LUT4AB/FrameData[4]
+ Tile_X2Y5_LUT4AB/FrameData[5] Tile_X2Y5_LUT4AB/FrameData[6] Tile_X2Y5_LUT4AB/FrameData[7]
+ Tile_X2Y5_LUT4AB/FrameData[8] Tile_X2Y5_LUT4AB/FrameData[9] Tile_X1Y5_LUT4AB/FrameStrobe[0]
+ Tile_X1Y5_LUT4AB/FrameStrobe[10] Tile_X1Y5_LUT4AB/FrameStrobe[11] Tile_X1Y5_LUT4AB/FrameStrobe[12]
+ Tile_X1Y5_LUT4AB/FrameStrobe[13] Tile_X1Y5_LUT4AB/FrameStrobe[14] Tile_X1Y5_LUT4AB/FrameStrobe[15]
+ Tile_X1Y5_LUT4AB/FrameStrobe[16] Tile_X1Y5_LUT4AB/FrameStrobe[17] Tile_X1Y5_LUT4AB/FrameStrobe[18]
+ Tile_X1Y5_LUT4AB/FrameStrobe[19] Tile_X1Y5_LUT4AB/FrameStrobe[1] Tile_X1Y5_LUT4AB/FrameStrobe[2]
+ Tile_X1Y5_LUT4AB/FrameStrobe[3] Tile_X1Y5_LUT4AB/FrameStrobe[4] Tile_X1Y5_LUT4AB/FrameStrobe[5]
+ Tile_X1Y5_LUT4AB/FrameStrobe[6] Tile_X1Y5_LUT4AB/FrameStrobe[7] Tile_X1Y5_LUT4AB/FrameStrobe[8]
+ Tile_X1Y5_LUT4AB/FrameStrobe[9] Tile_X1Y4_LUT4AB/FrameStrobe[0] Tile_X1Y4_LUT4AB/FrameStrobe[10]
+ Tile_X1Y4_LUT4AB/FrameStrobe[11] Tile_X1Y4_LUT4AB/FrameStrobe[12] Tile_X1Y4_LUT4AB/FrameStrobe[13]
+ Tile_X1Y4_LUT4AB/FrameStrobe[14] Tile_X1Y4_LUT4AB/FrameStrobe[15] Tile_X1Y4_LUT4AB/FrameStrobe[16]
+ Tile_X1Y4_LUT4AB/FrameStrobe[17] Tile_X1Y4_LUT4AB/FrameStrobe[18] Tile_X1Y4_LUT4AB/FrameStrobe[19]
+ Tile_X1Y4_LUT4AB/FrameStrobe[1] Tile_X1Y4_LUT4AB/FrameStrobe[2] Tile_X1Y4_LUT4AB/FrameStrobe[3]
+ Tile_X1Y4_LUT4AB/FrameStrobe[4] Tile_X1Y4_LUT4AB/FrameStrobe[5] Tile_X1Y4_LUT4AB/FrameStrobe[6]
+ Tile_X1Y4_LUT4AB/FrameStrobe[7] Tile_X1Y4_LUT4AB/FrameStrobe[8] Tile_X1Y4_LUT4AB/FrameStrobe[9]
+ Tile_X1Y5_LUT4AB/N1BEG[0] Tile_X1Y5_LUT4AB/N1BEG[1] Tile_X1Y5_LUT4AB/N1BEG[2] Tile_X1Y5_LUT4AB/N1BEG[3]
+ Tile_X1Y6_LUT4AB/N1BEG[0] Tile_X1Y6_LUT4AB/N1BEG[1] Tile_X1Y6_LUT4AB/N1BEG[2] Tile_X1Y6_LUT4AB/N1BEG[3]
+ Tile_X1Y5_LUT4AB/N2BEG[0] Tile_X1Y5_LUT4AB/N2BEG[1] Tile_X1Y5_LUT4AB/N2BEG[2] Tile_X1Y5_LUT4AB/N2BEG[3]
+ Tile_X1Y5_LUT4AB/N2BEG[4] Tile_X1Y5_LUT4AB/N2BEG[5] Tile_X1Y5_LUT4AB/N2BEG[6] Tile_X1Y5_LUT4AB/N2BEG[7]
+ Tile_X1Y4_LUT4AB/N2END[0] Tile_X1Y4_LUT4AB/N2END[1] Tile_X1Y4_LUT4AB/N2END[2] Tile_X1Y4_LUT4AB/N2END[3]
+ Tile_X1Y4_LUT4AB/N2END[4] Tile_X1Y4_LUT4AB/N2END[5] Tile_X1Y4_LUT4AB/N2END[6] Tile_X1Y4_LUT4AB/N2END[7]
+ Tile_X1Y5_LUT4AB/N2END[0] Tile_X1Y5_LUT4AB/N2END[1] Tile_X1Y5_LUT4AB/N2END[2] Tile_X1Y5_LUT4AB/N2END[3]
+ Tile_X1Y5_LUT4AB/N2END[4] Tile_X1Y5_LUT4AB/N2END[5] Tile_X1Y5_LUT4AB/N2END[6] Tile_X1Y5_LUT4AB/N2END[7]
+ Tile_X1Y6_LUT4AB/N2BEG[0] Tile_X1Y6_LUT4AB/N2BEG[1] Tile_X1Y6_LUT4AB/N2BEG[2] Tile_X1Y6_LUT4AB/N2BEG[3]
+ Tile_X1Y6_LUT4AB/N2BEG[4] Tile_X1Y6_LUT4AB/N2BEG[5] Tile_X1Y6_LUT4AB/N2BEG[6] Tile_X1Y6_LUT4AB/N2BEG[7]
+ Tile_X1Y5_LUT4AB/N4BEG[0] Tile_X1Y5_LUT4AB/N4BEG[10] Tile_X1Y5_LUT4AB/N4BEG[11]
+ Tile_X1Y5_LUT4AB/N4BEG[12] Tile_X1Y5_LUT4AB/N4BEG[13] Tile_X1Y5_LUT4AB/N4BEG[14]
+ Tile_X1Y5_LUT4AB/N4BEG[15] Tile_X1Y5_LUT4AB/N4BEG[1] Tile_X1Y5_LUT4AB/N4BEG[2] Tile_X1Y5_LUT4AB/N4BEG[3]
+ Tile_X1Y5_LUT4AB/N4BEG[4] Tile_X1Y5_LUT4AB/N4BEG[5] Tile_X1Y5_LUT4AB/N4BEG[6] Tile_X1Y5_LUT4AB/N4BEG[7]
+ Tile_X1Y5_LUT4AB/N4BEG[8] Tile_X1Y5_LUT4AB/N4BEG[9] Tile_X1Y6_LUT4AB/N4BEG[0] Tile_X1Y6_LUT4AB/N4BEG[10]
+ Tile_X1Y6_LUT4AB/N4BEG[11] Tile_X1Y6_LUT4AB/N4BEG[12] Tile_X1Y6_LUT4AB/N4BEG[13]
+ Tile_X1Y6_LUT4AB/N4BEG[14] Tile_X1Y6_LUT4AB/N4BEG[15] Tile_X1Y6_LUT4AB/N4BEG[1]
+ Tile_X1Y6_LUT4AB/N4BEG[2] Tile_X1Y6_LUT4AB/N4BEG[3] Tile_X1Y6_LUT4AB/N4BEG[4] Tile_X1Y6_LUT4AB/N4BEG[5]
+ Tile_X1Y6_LUT4AB/N4BEG[6] Tile_X1Y6_LUT4AB/N4BEG[7] Tile_X1Y6_LUT4AB/N4BEG[8] Tile_X1Y6_LUT4AB/N4BEG[9]
+ Tile_X1Y5_LUT4AB/NN4BEG[0] Tile_X1Y5_LUT4AB/NN4BEG[10] Tile_X1Y5_LUT4AB/NN4BEG[11]
+ Tile_X1Y5_LUT4AB/NN4BEG[12] Tile_X1Y5_LUT4AB/NN4BEG[13] Tile_X1Y5_LUT4AB/NN4BEG[14]
+ Tile_X1Y5_LUT4AB/NN4BEG[15] Tile_X1Y5_LUT4AB/NN4BEG[1] Tile_X1Y5_LUT4AB/NN4BEG[2]
+ Tile_X1Y5_LUT4AB/NN4BEG[3] Tile_X1Y5_LUT4AB/NN4BEG[4] Tile_X1Y5_LUT4AB/NN4BEG[5]
+ Tile_X1Y5_LUT4AB/NN4BEG[6] Tile_X1Y5_LUT4AB/NN4BEG[7] Tile_X1Y5_LUT4AB/NN4BEG[8]
+ Tile_X1Y5_LUT4AB/NN4BEG[9] Tile_X1Y6_LUT4AB/NN4BEG[0] Tile_X1Y6_LUT4AB/NN4BEG[10]
+ Tile_X1Y6_LUT4AB/NN4BEG[11] Tile_X1Y6_LUT4AB/NN4BEG[12] Tile_X1Y6_LUT4AB/NN4BEG[13]
+ Tile_X1Y6_LUT4AB/NN4BEG[14] Tile_X1Y6_LUT4AB/NN4BEG[15] Tile_X1Y6_LUT4AB/NN4BEG[1]
+ Tile_X1Y6_LUT4AB/NN4BEG[2] Tile_X1Y6_LUT4AB/NN4BEG[3] Tile_X1Y6_LUT4AB/NN4BEG[4]
+ Tile_X1Y6_LUT4AB/NN4BEG[5] Tile_X1Y6_LUT4AB/NN4BEG[6] Tile_X1Y6_LUT4AB/NN4BEG[7]
+ Tile_X1Y6_LUT4AB/NN4BEG[8] Tile_X1Y6_LUT4AB/NN4BEG[9] Tile_X1Y6_LUT4AB/S1END[0]
+ Tile_X1Y6_LUT4AB/S1END[1] Tile_X1Y6_LUT4AB/S1END[2] Tile_X1Y6_LUT4AB/S1END[3] Tile_X1Y5_LUT4AB/S1END[0]
+ Tile_X1Y5_LUT4AB/S1END[1] Tile_X1Y5_LUT4AB/S1END[2] Tile_X1Y5_LUT4AB/S1END[3] Tile_X1Y6_LUT4AB/S2MID[0]
+ Tile_X1Y6_LUT4AB/S2MID[1] Tile_X1Y6_LUT4AB/S2MID[2] Tile_X1Y6_LUT4AB/S2MID[3] Tile_X1Y6_LUT4AB/S2MID[4]
+ Tile_X1Y6_LUT4AB/S2MID[5] Tile_X1Y6_LUT4AB/S2MID[6] Tile_X1Y6_LUT4AB/S2MID[7] Tile_X1Y6_LUT4AB/S2END[0]
+ Tile_X1Y6_LUT4AB/S2END[1] Tile_X1Y6_LUT4AB/S2END[2] Tile_X1Y6_LUT4AB/S2END[3] Tile_X1Y6_LUT4AB/S2END[4]
+ Tile_X1Y6_LUT4AB/S2END[5] Tile_X1Y6_LUT4AB/S2END[6] Tile_X1Y6_LUT4AB/S2END[7] Tile_X1Y5_LUT4AB/S2END[0]
+ Tile_X1Y5_LUT4AB/S2END[1] Tile_X1Y5_LUT4AB/S2END[2] Tile_X1Y5_LUT4AB/S2END[3] Tile_X1Y5_LUT4AB/S2END[4]
+ Tile_X1Y5_LUT4AB/S2END[5] Tile_X1Y5_LUT4AB/S2END[6] Tile_X1Y5_LUT4AB/S2END[7] Tile_X1Y5_LUT4AB/S2MID[0]
+ Tile_X1Y5_LUT4AB/S2MID[1] Tile_X1Y5_LUT4AB/S2MID[2] Tile_X1Y5_LUT4AB/S2MID[3] Tile_X1Y5_LUT4AB/S2MID[4]
+ Tile_X1Y5_LUT4AB/S2MID[5] Tile_X1Y5_LUT4AB/S2MID[6] Tile_X1Y5_LUT4AB/S2MID[7] Tile_X1Y6_LUT4AB/S4END[0]
+ Tile_X1Y6_LUT4AB/S4END[10] Tile_X1Y6_LUT4AB/S4END[11] Tile_X1Y6_LUT4AB/S4END[12]
+ Tile_X1Y6_LUT4AB/S4END[13] Tile_X1Y6_LUT4AB/S4END[14] Tile_X1Y6_LUT4AB/S4END[15]
+ Tile_X1Y6_LUT4AB/S4END[1] Tile_X1Y6_LUT4AB/S4END[2] Tile_X1Y6_LUT4AB/S4END[3] Tile_X1Y6_LUT4AB/S4END[4]
+ Tile_X1Y6_LUT4AB/S4END[5] Tile_X1Y6_LUT4AB/S4END[6] Tile_X1Y6_LUT4AB/S4END[7] Tile_X1Y6_LUT4AB/S4END[8]
+ Tile_X1Y6_LUT4AB/S4END[9] Tile_X1Y5_LUT4AB/S4END[0] Tile_X1Y5_LUT4AB/S4END[10] Tile_X1Y5_LUT4AB/S4END[11]
+ Tile_X1Y5_LUT4AB/S4END[12] Tile_X1Y5_LUT4AB/S4END[13] Tile_X1Y5_LUT4AB/S4END[14]
+ Tile_X1Y5_LUT4AB/S4END[15] Tile_X1Y5_LUT4AB/S4END[1] Tile_X1Y5_LUT4AB/S4END[2] Tile_X1Y5_LUT4AB/S4END[3]
+ Tile_X1Y5_LUT4AB/S4END[4] Tile_X1Y5_LUT4AB/S4END[5] Tile_X1Y5_LUT4AB/S4END[6] Tile_X1Y5_LUT4AB/S4END[7]
+ Tile_X1Y5_LUT4AB/S4END[8] Tile_X1Y5_LUT4AB/S4END[9] Tile_X1Y6_LUT4AB/SS4END[0] Tile_X1Y6_LUT4AB/SS4END[10]
+ Tile_X1Y6_LUT4AB/SS4END[11] Tile_X1Y6_LUT4AB/SS4END[12] Tile_X1Y6_LUT4AB/SS4END[13]
+ Tile_X1Y6_LUT4AB/SS4END[14] Tile_X1Y6_LUT4AB/SS4END[15] Tile_X1Y6_LUT4AB/SS4END[1]
+ Tile_X1Y6_LUT4AB/SS4END[2] Tile_X1Y6_LUT4AB/SS4END[3] Tile_X1Y6_LUT4AB/SS4END[4]
+ Tile_X1Y6_LUT4AB/SS4END[5] Tile_X1Y6_LUT4AB/SS4END[6] Tile_X1Y6_LUT4AB/SS4END[7]
+ Tile_X1Y6_LUT4AB/SS4END[8] Tile_X1Y6_LUT4AB/SS4END[9] Tile_X1Y5_LUT4AB/SS4END[0]
+ Tile_X1Y5_LUT4AB/SS4END[10] Tile_X1Y5_LUT4AB/SS4END[11] Tile_X1Y5_LUT4AB/SS4END[12]
+ Tile_X1Y5_LUT4AB/SS4END[13] Tile_X1Y5_LUT4AB/SS4END[14] Tile_X1Y5_LUT4AB/SS4END[15]
+ Tile_X1Y5_LUT4AB/SS4END[1] Tile_X1Y5_LUT4AB/SS4END[2] Tile_X1Y5_LUT4AB/SS4END[3]
+ Tile_X1Y5_LUT4AB/SS4END[4] Tile_X1Y5_LUT4AB/SS4END[5] Tile_X1Y5_LUT4AB/SS4END[6]
+ Tile_X1Y5_LUT4AB/SS4END[7] Tile_X1Y5_LUT4AB/SS4END[8] Tile_X1Y5_LUT4AB/SS4END[9]
+ Tile_X1Y5_LUT4AB/UserCLK Tile_X1Y4_LUT4AB/UserCLK VGND VPWR Tile_X0Y5_W_IO/W1END[0]
+ Tile_X0Y5_W_IO/W1END[1] Tile_X0Y5_W_IO/W1END[2] Tile_X0Y5_W_IO/W1END[3] Tile_X2Y5_LUT4AB/W1BEG[0]
+ Tile_X2Y5_LUT4AB/W1BEG[1] Tile_X2Y5_LUT4AB/W1BEG[2] Tile_X2Y5_LUT4AB/W1BEG[3] Tile_X0Y5_W_IO/W2MID[0]
+ Tile_X0Y5_W_IO/W2MID[1] Tile_X0Y5_W_IO/W2MID[2] Tile_X0Y5_W_IO/W2MID[3] Tile_X0Y5_W_IO/W2MID[4]
+ Tile_X0Y5_W_IO/W2MID[5] Tile_X0Y5_W_IO/W2MID[6] Tile_X0Y5_W_IO/W2MID[7] Tile_X0Y5_W_IO/W2END[0]
+ Tile_X0Y5_W_IO/W2END[1] Tile_X0Y5_W_IO/W2END[2] Tile_X0Y5_W_IO/W2END[3] Tile_X0Y5_W_IO/W2END[4]
+ Tile_X0Y5_W_IO/W2END[5] Tile_X0Y5_W_IO/W2END[6] Tile_X0Y5_W_IO/W2END[7] Tile_X1Y5_LUT4AB/W2END[0]
+ Tile_X1Y5_LUT4AB/W2END[1] Tile_X1Y5_LUT4AB/W2END[2] Tile_X1Y5_LUT4AB/W2END[3] Tile_X1Y5_LUT4AB/W2END[4]
+ Tile_X1Y5_LUT4AB/W2END[5] Tile_X1Y5_LUT4AB/W2END[6] Tile_X1Y5_LUT4AB/W2END[7] Tile_X2Y5_LUT4AB/W2BEG[0]
+ Tile_X2Y5_LUT4AB/W2BEG[1] Tile_X2Y5_LUT4AB/W2BEG[2] Tile_X2Y5_LUT4AB/W2BEG[3] Tile_X2Y5_LUT4AB/W2BEG[4]
+ Tile_X2Y5_LUT4AB/W2BEG[5] Tile_X2Y5_LUT4AB/W2BEG[6] Tile_X2Y5_LUT4AB/W2BEG[7] Tile_X0Y5_W_IO/W6END[0]
+ Tile_X0Y5_W_IO/W6END[10] Tile_X0Y5_W_IO/W6END[11] Tile_X0Y5_W_IO/W6END[1] Tile_X0Y5_W_IO/W6END[2]
+ Tile_X0Y5_W_IO/W6END[3] Tile_X0Y5_W_IO/W6END[4] Tile_X0Y5_W_IO/W6END[5] Tile_X0Y5_W_IO/W6END[6]
+ Tile_X0Y5_W_IO/W6END[7] Tile_X0Y5_W_IO/W6END[8] Tile_X0Y5_W_IO/W6END[9] Tile_X2Y5_LUT4AB/W6BEG[0]
+ Tile_X2Y5_LUT4AB/W6BEG[10] Tile_X2Y5_LUT4AB/W6BEG[11] Tile_X2Y5_LUT4AB/W6BEG[1]
+ Tile_X2Y5_LUT4AB/W6BEG[2] Tile_X2Y5_LUT4AB/W6BEG[3] Tile_X2Y5_LUT4AB/W6BEG[4] Tile_X2Y5_LUT4AB/W6BEG[5]
+ Tile_X2Y5_LUT4AB/W6BEG[6] Tile_X2Y5_LUT4AB/W6BEG[7] Tile_X2Y5_LUT4AB/W6BEG[8] Tile_X2Y5_LUT4AB/W6BEG[9]
+ Tile_X0Y5_W_IO/WW4END[0] Tile_X0Y5_W_IO/WW4END[10] Tile_X0Y5_W_IO/WW4END[11] Tile_X0Y5_W_IO/WW4END[12]
+ Tile_X0Y5_W_IO/WW4END[13] Tile_X0Y5_W_IO/WW4END[14] Tile_X0Y5_W_IO/WW4END[15] Tile_X0Y5_W_IO/WW4END[1]
+ Tile_X0Y5_W_IO/WW4END[2] Tile_X0Y5_W_IO/WW4END[3] Tile_X0Y5_W_IO/WW4END[4] Tile_X0Y5_W_IO/WW4END[5]
+ Tile_X0Y5_W_IO/WW4END[6] Tile_X0Y5_W_IO/WW4END[7] Tile_X0Y5_W_IO/WW4END[8] Tile_X0Y5_W_IO/WW4END[9]
+ Tile_X2Y5_LUT4AB/WW4BEG[0] Tile_X2Y5_LUT4AB/WW4BEG[10] Tile_X2Y5_LUT4AB/WW4BEG[11]
+ Tile_X2Y5_LUT4AB/WW4BEG[12] Tile_X2Y5_LUT4AB/WW4BEG[13] Tile_X2Y5_LUT4AB/WW4BEG[14]
+ Tile_X2Y5_LUT4AB/WW4BEG[15] Tile_X2Y5_LUT4AB/WW4BEG[1] Tile_X2Y5_LUT4AB/WW4BEG[2]
+ Tile_X2Y5_LUT4AB/WW4BEG[3] Tile_X2Y5_LUT4AB/WW4BEG[4] Tile_X2Y5_LUT4AB/WW4BEG[5]
+ Tile_X2Y5_LUT4AB/WW4BEG[6] Tile_X2Y5_LUT4AB/WW4BEG[7] Tile_X2Y5_LUT4AB/WW4BEG[8]
+ Tile_X2Y5_LUT4AB/WW4BEG[9] LUT4AB
XTile_X10Y9_IHP_SRAM Tile_X10Y10_ADDR_SRAM0 Tile_X10Y10_ADDR_SRAM1 Tile_X10Y10_ADDR_SRAM2
+ Tile_X10Y10_ADDR_SRAM3 Tile_X10Y10_ADDR_SRAM4 Tile_X10Y10_ADDR_SRAM5 Tile_X10Y10_ADDR_SRAM6
+ Tile_X10Y10_ADDR_SRAM7 Tile_X10Y10_ADDR_SRAM8 Tile_X10Y10_ADDR_SRAM9 Tile_X10Y10_BM_SRAM0
+ Tile_X10Y10_BM_SRAM1 Tile_X10Y10_BM_SRAM10 Tile_X10Y10_BM_SRAM11 Tile_X10Y10_BM_SRAM12
+ Tile_X10Y10_BM_SRAM13 Tile_X10Y10_BM_SRAM14 Tile_X10Y10_BM_SRAM15 Tile_X10Y10_BM_SRAM16
+ Tile_X10Y10_BM_SRAM17 Tile_X10Y10_BM_SRAM18 Tile_X10Y10_BM_SRAM19 Tile_X10Y10_BM_SRAM2
+ Tile_X10Y10_BM_SRAM20 Tile_X10Y10_BM_SRAM21 Tile_X10Y10_BM_SRAM22 Tile_X10Y10_BM_SRAM23
+ Tile_X10Y10_BM_SRAM24 Tile_X10Y10_BM_SRAM25 Tile_X10Y10_BM_SRAM26 Tile_X10Y10_BM_SRAM27
+ Tile_X10Y10_BM_SRAM28 Tile_X10Y10_BM_SRAM29 Tile_X10Y10_BM_SRAM3 Tile_X10Y10_BM_SRAM30
+ Tile_X10Y10_BM_SRAM31 Tile_X10Y10_BM_SRAM4 Tile_X10Y10_BM_SRAM5 Tile_X10Y10_BM_SRAM6
+ Tile_X10Y10_BM_SRAM7 Tile_X10Y10_BM_SRAM8 Tile_X10Y10_BM_SRAM9 Tile_X10Y10_CLK_SRAM
+ Tile_X10Y10_CONFIGURED_top Tile_X10Y10_DIN_SRAM0 Tile_X10Y10_DIN_SRAM1 Tile_X10Y10_DIN_SRAM10
+ Tile_X10Y10_DIN_SRAM11 Tile_X10Y10_DIN_SRAM12 Tile_X10Y10_DIN_SRAM13 Tile_X10Y10_DIN_SRAM14
+ Tile_X10Y10_DIN_SRAM15 Tile_X10Y10_DIN_SRAM16 Tile_X10Y10_DIN_SRAM17 Tile_X10Y10_DIN_SRAM18
+ Tile_X10Y10_DIN_SRAM19 Tile_X10Y10_DIN_SRAM2 Tile_X10Y10_DIN_SRAM20 Tile_X10Y10_DIN_SRAM21
+ Tile_X10Y10_DIN_SRAM22 Tile_X10Y10_DIN_SRAM23 Tile_X10Y10_DIN_SRAM24 Tile_X10Y10_DIN_SRAM25
+ Tile_X10Y10_DIN_SRAM26 Tile_X10Y10_DIN_SRAM27 Tile_X10Y10_DIN_SRAM28 Tile_X10Y10_DIN_SRAM29
+ Tile_X10Y10_DIN_SRAM3 Tile_X10Y10_DIN_SRAM30 Tile_X10Y10_DIN_SRAM31 Tile_X10Y10_DIN_SRAM4
+ Tile_X10Y10_DIN_SRAM5 Tile_X10Y10_DIN_SRAM6 Tile_X10Y10_DIN_SRAM7 Tile_X10Y10_DIN_SRAM8
+ Tile_X10Y10_DIN_SRAM9 Tile_X10Y10_DOUT_SRAM0 Tile_X10Y10_DOUT_SRAM1 Tile_X10Y10_DOUT_SRAM10
+ Tile_X10Y10_DOUT_SRAM11 Tile_X10Y10_DOUT_SRAM12 Tile_X10Y10_DOUT_SRAM13 Tile_X10Y10_DOUT_SRAM14
+ Tile_X10Y10_DOUT_SRAM15 Tile_X10Y10_DOUT_SRAM16 Tile_X10Y10_DOUT_SRAM17 Tile_X10Y10_DOUT_SRAM18
+ Tile_X10Y10_DOUT_SRAM19 Tile_X10Y10_DOUT_SRAM2 Tile_X10Y10_DOUT_SRAM20 Tile_X10Y10_DOUT_SRAM21
+ Tile_X10Y10_DOUT_SRAM22 Tile_X10Y10_DOUT_SRAM23 Tile_X10Y10_DOUT_SRAM24 Tile_X10Y10_DOUT_SRAM25
+ Tile_X10Y10_DOUT_SRAM26 Tile_X10Y10_DOUT_SRAM27 Tile_X10Y10_DOUT_SRAM28 Tile_X10Y10_DOUT_SRAM29
+ Tile_X10Y10_DOUT_SRAM3 Tile_X10Y10_DOUT_SRAM30 Tile_X10Y10_DOUT_SRAM31 Tile_X10Y10_DOUT_SRAM4
+ Tile_X10Y10_DOUT_SRAM5 Tile_X10Y10_DOUT_SRAM6 Tile_X10Y10_DOUT_SRAM7 Tile_X10Y10_DOUT_SRAM8
+ Tile_X10Y10_DOUT_SRAM9 Tile_X10Y10_MEN_SRAM Tile_X10Y10_REN_SRAM Tile_X10Y10_TIE_HIGH_SRAM
+ Tile_X10Y10_TIE_LOW_SRAM Tile_X9Y9_LUT4AB/E1BEG[0] Tile_X9Y9_LUT4AB/E1BEG[1] Tile_X9Y9_LUT4AB/E1BEG[2]
+ Tile_X9Y9_LUT4AB/E1BEG[3] Tile_X9Y9_LUT4AB/E2BEGb[0] Tile_X9Y9_LUT4AB/E2BEGb[1]
+ Tile_X9Y9_LUT4AB/E2BEGb[2] Tile_X9Y9_LUT4AB/E2BEGb[3] Tile_X9Y9_LUT4AB/E2BEGb[4]
+ Tile_X9Y9_LUT4AB/E2BEGb[5] Tile_X9Y9_LUT4AB/E2BEGb[6] Tile_X9Y9_LUT4AB/E2BEGb[7]
+ Tile_X9Y9_LUT4AB/E2BEG[0] Tile_X9Y9_LUT4AB/E2BEG[1] Tile_X9Y9_LUT4AB/E2BEG[2] Tile_X9Y9_LUT4AB/E2BEG[3]
+ Tile_X9Y9_LUT4AB/E2BEG[4] Tile_X9Y9_LUT4AB/E2BEG[5] Tile_X9Y9_LUT4AB/E2BEG[6] Tile_X9Y9_LUT4AB/E2BEG[7]
+ Tile_X9Y9_LUT4AB/E6BEG[0] Tile_X9Y9_LUT4AB/E6BEG[10] Tile_X9Y9_LUT4AB/E6BEG[11]
+ Tile_X9Y9_LUT4AB/E6BEG[1] Tile_X9Y9_LUT4AB/E6BEG[2] Tile_X9Y9_LUT4AB/E6BEG[3] Tile_X9Y9_LUT4AB/E6BEG[4]
+ Tile_X9Y9_LUT4AB/E6BEG[5] Tile_X9Y9_LUT4AB/E6BEG[6] Tile_X9Y9_LUT4AB/E6BEG[7] Tile_X9Y9_LUT4AB/E6BEG[8]
+ Tile_X9Y9_LUT4AB/E6BEG[9] Tile_X9Y9_LUT4AB/EE4BEG[0] Tile_X9Y9_LUT4AB/EE4BEG[10]
+ Tile_X9Y9_LUT4AB/EE4BEG[11] Tile_X9Y9_LUT4AB/EE4BEG[12] Tile_X9Y9_LUT4AB/EE4BEG[13]
+ Tile_X9Y9_LUT4AB/EE4BEG[14] Tile_X9Y9_LUT4AB/EE4BEG[15] Tile_X9Y9_LUT4AB/EE4BEG[1]
+ Tile_X9Y9_LUT4AB/EE4BEG[2] Tile_X9Y9_LUT4AB/EE4BEG[3] Tile_X9Y9_LUT4AB/EE4BEG[4]
+ Tile_X9Y9_LUT4AB/EE4BEG[5] Tile_X9Y9_LUT4AB/EE4BEG[6] Tile_X9Y9_LUT4AB/EE4BEG[7]
+ Tile_X9Y9_LUT4AB/EE4BEG[8] Tile_X9Y9_LUT4AB/EE4BEG[9] Tile_X9Y9_LUT4AB/FrameData_O[0]
+ Tile_X9Y9_LUT4AB/FrameData_O[10] Tile_X9Y9_LUT4AB/FrameData_O[11] Tile_X9Y9_LUT4AB/FrameData_O[12]
+ Tile_X9Y9_LUT4AB/FrameData_O[13] Tile_X9Y9_LUT4AB/FrameData_O[14] Tile_X9Y9_LUT4AB/FrameData_O[15]
+ Tile_X9Y9_LUT4AB/FrameData_O[16] Tile_X9Y9_LUT4AB/FrameData_O[17] Tile_X9Y9_LUT4AB/FrameData_O[18]
+ Tile_X9Y9_LUT4AB/FrameData_O[19] Tile_X9Y9_LUT4AB/FrameData_O[1] Tile_X9Y9_LUT4AB/FrameData_O[20]
+ Tile_X9Y9_LUT4AB/FrameData_O[21] Tile_X9Y9_LUT4AB/FrameData_O[22] Tile_X9Y9_LUT4AB/FrameData_O[23]
+ Tile_X9Y9_LUT4AB/FrameData_O[24] Tile_X9Y9_LUT4AB/FrameData_O[25] Tile_X9Y9_LUT4AB/FrameData_O[26]
+ Tile_X9Y9_LUT4AB/FrameData_O[27] Tile_X9Y9_LUT4AB/FrameData_O[28] Tile_X9Y9_LUT4AB/FrameData_O[29]
+ Tile_X9Y9_LUT4AB/FrameData_O[2] Tile_X9Y9_LUT4AB/FrameData_O[30] Tile_X9Y9_LUT4AB/FrameData_O[31]
+ Tile_X9Y9_LUT4AB/FrameData_O[3] Tile_X9Y9_LUT4AB/FrameData_O[4] Tile_X9Y9_LUT4AB/FrameData_O[5]
+ Tile_X9Y9_LUT4AB/FrameData_O[6] Tile_X9Y9_LUT4AB/FrameData_O[7] Tile_X9Y9_LUT4AB/FrameData_O[8]
+ Tile_X9Y9_LUT4AB/FrameData_O[9] Tile_X10Y9_IHP_SRAM/Tile_X0Y0_FrameData_O[0] Tile_X10Y9_IHP_SRAM/Tile_X0Y0_FrameData_O[10]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y0_FrameData_O[11] Tile_X10Y9_IHP_SRAM/Tile_X0Y0_FrameData_O[12]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y0_FrameData_O[13] Tile_X10Y9_IHP_SRAM/Tile_X0Y0_FrameData_O[14]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y0_FrameData_O[15] Tile_X10Y9_IHP_SRAM/Tile_X0Y0_FrameData_O[16]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y0_FrameData_O[17] Tile_X10Y9_IHP_SRAM/Tile_X0Y0_FrameData_O[18]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y0_FrameData_O[19] Tile_X10Y9_IHP_SRAM/Tile_X0Y0_FrameData_O[1]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y0_FrameData_O[20] Tile_X10Y9_IHP_SRAM/Tile_X0Y0_FrameData_O[21]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y0_FrameData_O[22] Tile_X10Y9_IHP_SRAM/Tile_X0Y0_FrameData_O[23]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y0_FrameData_O[24] Tile_X10Y9_IHP_SRAM/Tile_X0Y0_FrameData_O[25]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y0_FrameData_O[26] Tile_X10Y9_IHP_SRAM/Tile_X0Y0_FrameData_O[27]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y0_FrameData_O[28] Tile_X10Y9_IHP_SRAM/Tile_X0Y0_FrameData_O[29]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y0_FrameData_O[2] Tile_X10Y9_IHP_SRAM/Tile_X0Y0_FrameData_O[30]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y0_FrameData_O[31] Tile_X10Y9_IHP_SRAM/Tile_X0Y0_FrameData_O[3]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y0_FrameData_O[4] Tile_X10Y9_IHP_SRAM/Tile_X0Y0_FrameData_O[5]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y0_FrameData_O[6] Tile_X10Y9_IHP_SRAM/Tile_X0Y0_FrameData_O[7]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y0_FrameData_O[8] Tile_X10Y9_IHP_SRAM/Tile_X0Y0_FrameData_O[9]
+ Tile_X10Y7_IHP_SRAM/Tile_X0Y1_FrameStrobe[0] Tile_X10Y7_IHP_SRAM/Tile_X0Y1_FrameStrobe[10]
+ Tile_X10Y7_IHP_SRAM/Tile_X0Y1_FrameStrobe[11] Tile_X10Y7_IHP_SRAM/Tile_X0Y1_FrameStrobe[12]
+ Tile_X10Y7_IHP_SRAM/Tile_X0Y1_FrameStrobe[13] Tile_X10Y7_IHP_SRAM/Tile_X0Y1_FrameStrobe[14]
+ Tile_X10Y7_IHP_SRAM/Tile_X0Y1_FrameStrobe[15] Tile_X10Y7_IHP_SRAM/Tile_X0Y1_FrameStrobe[16]
+ Tile_X10Y7_IHP_SRAM/Tile_X0Y1_FrameStrobe[17] Tile_X10Y7_IHP_SRAM/Tile_X0Y1_FrameStrobe[18]
+ Tile_X10Y7_IHP_SRAM/Tile_X0Y1_FrameStrobe[19] Tile_X10Y7_IHP_SRAM/Tile_X0Y1_FrameStrobe[1]
+ Tile_X10Y7_IHP_SRAM/Tile_X0Y1_FrameStrobe[2] Tile_X10Y7_IHP_SRAM/Tile_X0Y1_FrameStrobe[3]
+ Tile_X10Y7_IHP_SRAM/Tile_X0Y1_FrameStrobe[4] Tile_X10Y7_IHP_SRAM/Tile_X0Y1_FrameStrobe[5]
+ Tile_X10Y7_IHP_SRAM/Tile_X0Y1_FrameStrobe[6] Tile_X10Y7_IHP_SRAM/Tile_X0Y1_FrameStrobe[7]
+ Tile_X10Y7_IHP_SRAM/Tile_X0Y1_FrameStrobe[8] Tile_X10Y7_IHP_SRAM/Tile_X0Y1_FrameStrobe[9]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y0_N1BEG[0] Tile_X10Y9_IHP_SRAM/Tile_X0Y0_N1BEG[1] Tile_X10Y9_IHP_SRAM/Tile_X0Y0_N1BEG[2]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y0_N1BEG[3] Tile_X10Y9_IHP_SRAM/Tile_X0Y0_N2BEG[0] Tile_X10Y9_IHP_SRAM/Tile_X0Y0_N2BEG[1]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y0_N2BEG[2] Tile_X10Y9_IHP_SRAM/Tile_X0Y0_N2BEG[3] Tile_X10Y9_IHP_SRAM/Tile_X0Y0_N2BEG[4]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y0_N2BEG[5] Tile_X10Y9_IHP_SRAM/Tile_X0Y0_N2BEG[6] Tile_X10Y9_IHP_SRAM/Tile_X0Y0_N2BEG[7]
+ Tile_X10Y7_IHP_SRAM/Tile_X0Y1_N2END[0] Tile_X10Y7_IHP_SRAM/Tile_X0Y1_N2END[1] Tile_X10Y7_IHP_SRAM/Tile_X0Y1_N2END[2]
+ Tile_X10Y7_IHP_SRAM/Tile_X0Y1_N2END[3] Tile_X10Y7_IHP_SRAM/Tile_X0Y1_N2END[4] Tile_X10Y7_IHP_SRAM/Tile_X0Y1_N2END[5]
+ Tile_X10Y7_IHP_SRAM/Tile_X0Y1_N2END[6] Tile_X10Y7_IHP_SRAM/Tile_X0Y1_N2END[7] Tile_X10Y9_IHP_SRAM/Tile_X0Y0_N4BEG[0]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y0_N4BEG[10] Tile_X10Y9_IHP_SRAM/Tile_X0Y0_N4BEG[11]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y0_N4BEG[12] Tile_X10Y9_IHP_SRAM/Tile_X0Y0_N4BEG[13]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y0_N4BEG[14] Tile_X10Y9_IHP_SRAM/Tile_X0Y0_N4BEG[15]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y0_N4BEG[1] Tile_X10Y9_IHP_SRAM/Tile_X0Y0_N4BEG[2] Tile_X10Y9_IHP_SRAM/Tile_X0Y0_N4BEG[3]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y0_N4BEG[4] Tile_X10Y9_IHP_SRAM/Tile_X0Y0_N4BEG[5] Tile_X10Y9_IHP_SRAM/Tile_X0Y0_N4BEG[6]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y0_N4BEG[7] Tile_X10Y9_IHP_SRAM/Tile_X0Y0_N4BEG[8] Tile_X10Y9_IHP_SRAM/Tile_X0Y0_N4BEG[9]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y0_S1END[0] Tile_X10Y9_IHP_SRAM/Tile_X0Y0_S1END[1] Tile_X10Y9_IHP_SRAM/Tile_X0Y0_S1END[2]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y0_S1END[3] Tile_X10Y9_IHP_SRAM/Tile_X0Y0_S2END[0] Tile_X10Y9_IHP_SRAM/Tile_X0Y0_S2END[1]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y0_S2END[2] Tile_X10Y9_IHP_SRAM/Tile_X0Y0_S2END[3] Tile_X10Y9_IHP_SRAM/Tile_X0Y0_S2END[4]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y0_S2END[5] Tile_X10Y9_IHP_SRAM/Tile_X0Y0_S2END[6] Tile_X10Y9_IHP_SRAM/Tile_X0Y0_S2END[7]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y0_S2MID[0] Tile_X10Y9_IHP_SRAM/Tile_X0Y0_S2MID[1] Tile_X10Y9_IHP_SRAM/Tile_X0Y0_S2MID[2]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y0_S2MID[3] Tile_X10Y9_IHP_SRAM/Tile_X0Y0_S2MID[4] Tile_X10Y9_IHP_SRAM/Tile_X0Y0_S2MID[5]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y0_S2MID[6] Tile_X10Y9_IHP_SRAM/Tile_X0Y0_S2MID[7] Tile_X10Y9_IHP_SRAM/Tile_X0Y0_S4END[0]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y0_S4END[10] Tile_X10Y9_IHP_SRAM/Tile_X0Y0_S4END[11]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y0_S4END[12] Tile_X10Y9_IHP_SRAM/Tile_X0Y0_S4END[13]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y0_S4END[14] Tile_X10Y9_IHP_SRAM/Tile_X0Y0_S4END[15]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y0_S4END[1] Tile_X10Y9_IHP_SRAM/Tile_X0Y0_S4END[2] Tile_X10Y9_IHP_SRAM/Tile_X0Y0_S4END[3]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y0_S4END[4] Tile_X10Y9_IHP_SRAM/Tile_X0Y0_S4END[5] Tile_X10Y9_IHP_SRAM/Tile_X0Y0_S4END[6]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y0_S4END[7] Tile_X10Y9_IHP_SRAM/Tile_X0Y0_S4END[8] Tile_X10Y9_IHP_SRAM/Tile_X0Y0_S4END[9]
+ Tile_X10Y7_IHP_SRAM/Tile_X0Y1_UserCLK Tile_X9Y9_LUT4AB/W1END[0] Tile_X9Y9_LUT4AB/W1END[1]
+ Tile_X9Y9_LUT4AB/W1END[2] Tile_X9Y9_LUT4AB/W1END[3] Tile_X9Y9_LUT4AB/W2MID[0] Tile_X9Y9_LUT4AB/W2MID[1]
+ Tile_X9Y9_LUT4AB/W2MID[2] Tile_X9Y9_LUT4AB/W2MID[3] Tile_X9Y9_LUT4AB/W2MID[4] Tile_X9Y9_LUT4AB/W2MID[5]
+ Tile_X9Y9_LUT4AB/W2MID[6] Tile_X9Y9_LUT4AB/W2MID[7] Tile_X9Y9_LUT4AB/W2END[0] Tile_X9Y9_LUT4AB/W2END[1]
+ Tile_X9Y9_LUT4AB/W2END[2] Tile_X9Y9_LUT4AB/W2END[3] Tile_X9Y9_LUT4AB/W2END[4] Tile_X9Y9_LUT4AB/W2END[5]
+ Tile_X9Y9_LUT4AB/W2END[6] Tile_X9Y9_LUT4AB/W2END[7] Tile_X9Y9_LUT4AB/W6END[0] Tile_X9Y9_LUT4AB/W6END[10]
+ Tile_X9Y9_LUT4AB/W6END[11] Tile_X9Y9_LUT4AB/W6END[1] Tile_X9Y9_LUT4AB/W6END[2] Tile_X9Y9_LUT4AB/W6END[3]
+ Tile_X9Y9_LUT4AB/W6END[4] Tile_X9Y9_LUT4AB/W6END[5] Tile_X9Y9_LUT4AB/W6END[6] Tile_X9Y9_LUT4AB/W6END[7]
+ Tile_X9Y9_LUT4AB/W6END[8] Tile_X9Y9_LUT4AB/W6END[9] Tile_X9Y9_LUT4AB/WW4END[0] Tile_X9Y9_LUT4AB/WW4END[10]
+ Tile_X9Y9_LUT4AB/WW4END[11] Tile_X9Y9_LUT4AB/WW4END[12] Tile_X9Y9_LUT4AB/WW4END[13]
+ Tile_X9Y9_LUT4AB/WW4END[14] Tile_X9Y9_LUT4AB/WW4END[15] Tile_X9Y9_LUT4AB/WW4END[1]
+ Tile_X9Y9_LUT4AB/WW4END[2] Tile_X9Y9_LUT4AB/WW4END[3] Tile_X9Y9_LUT4AB/WW4END[4]
+ Tile_X9Y9_LUT4AB/WW4END[5] Tile_X9Y9_LUT4AB/WW4END[6] Tile_X9Y9_LUT4AB/WW4END[7]
+ Tile_X9Y9_LUT4AB/WW4END[8] Tile_X9Y9_LUT4AB/WW4END[9] Tile_X9Y10_LUT4AB/E1BEG[0]
+ Tile_X9Y10_LUT4AB/E1BEG[1] Tile_X9Y10_LUT4AB/E1BEG[2] Tile_X9Y10_LUT4AB/E1BEG[3]
+ Tile_X9Y10_LUT4AB/E2BEGb[0] Tile_X9Y10_LUT4AB/E2BEGb[1] Tile_X9Y10_LUT4AB/E2BEGb[2]
+ Tile_X9Y10_LUT4AB/E2BEGb[3] Tile_X9Y10_LUT4AB/E2BEGb[4] Tile_X9Y10_LUT4AB/E2BEGb[5]
+ Tile_X9Y10_LUT4AB/E2BEGb[6] Tile_X9Y10_LUT4AB/E2BEGb[7] Tile_X9Y10_LUT4AB/E2BEG[0]
+ Tile_X9Y10_LUT4AB/E2BEG[1] Tile_X9Y10_LUT4AB/E2BEG[2] Tile_X9Y10_LUT4AB/E2BEG[3]
+ Tile_X9Y10_LUT4AB/E2BEG[4] Tile_X9Y10_LUT4AB/E2BEG[5] Tile_X9Y10_LUT4AB/E2BEG[6]
+ Tile_X9Y10_LUT4AB/E2BEG[7] Tile_X9Y10_LUT4AB/E6BEG[0] Tile_X9Y10_LUT4AB/E6BEG[10]
+ Tile_X9Y10_LUT4AB/E6BEG[11] Tile_X9Y10_LUT4AB/E6BEG[1] Tile_X9Y10_LUT4AB/E6BEG[2]
+ Tile_X9Y10_LUT4AB/E6BEG[3] Tile_X9Y10_LUT4AB/E6BEG[4] Tile_X9Y10_LUT4AB/E6BEG[5]
+ Tile_X9Y10_LUT4AB/E6BEG[6] Tile_X9Y10_LUT4AB/E6BEG[7] Tile_X9Y10_LUT4AB/E6BEG[8]
+ Tile_X9Y10_LUT4AB/E6BEG[9] Tile_X9Y10_LUT4AB/EE4BEG[0] Tile_X9Y10_LUT4AB/EE4BEG[10]
+ Tile_X9Y10_LUT4AB/EE4BEG[11] Tile_X9Y10_LUT4AB/EE4BEG[12] Tile_X9Y10_LUT4AB/EE4BEG[13]
+ Tile_X9Y10_LUT4AB/EE4BEG[14] Tile_X9Y10_LUT4AB/EE4BEG[15] Tile_X9Y10_LUT4AB/EE4BEG[1]
+ Tile_X9Y10_LUT4AB/EE4BEG[2] Tile_X9Y10_LUT4AB/EE4BEG[3] Tile_X9Y10_LUT4AB/EE4BEG[4]
+ Tile_X9Y10_LUT4AB/EE4BEG[5] Tile_X9Y10_LUT4AB/EE4BEG[6] Tile_X9Y10_LUT4AB/EE4BEG[7]
+ Tile_X9Y10_LUT4AB/EE4BEG[8] Tile_X9Y10_LUT4AB/EE4BEG[9] Tile_X9Y10_LUT4AB/FrameData_O[0]
+ Tile_X9Y10_LUT4AB/FrameData_O[10] Tile_X9Y10_LUT4AB/FrameData_O[11] Tile_X9Y10_LUT4AB/FrameData_O[12]
+ Tile_X9Y10_LUT4AB/FrameData_O[13] Tile_X9Y10_LUT4AB/FrameData_O[14] Tile_X9Y10_LUT4AB/FrameData_O[15]
+ Tile_X9Y10_LUT4AB/FrameData_O[16] Tile_X9Y10_LUT4AB/FrameData_O[17] Tile_X9Y10_LUT4AB/FrameData_O[18]
+ Tile_X9Y10_LUT4AB/FrameData_O[19] Tile_X9Y10_LUT4AB/FrameData_O[1] Tile_X9Y10_LUT4AB/FrameData_O[20]
+ Tile_X9Y10_LUT4AB/FrameData_O[21] Tile_X9Y10_LUT4AB/FrameData_O[22] Tile_X9Y10_LUT4AB/FrameData_O[23]
+ Tile_X9Y10_LUT4AB/FrameData_O[24] Tile_X9Y10_LUT4AB/FrameData_O[25] Tile_X9Y10_LUT4AB/FrameData_O[26]
+ Tile_X9Y10_LUT4AB/FrameData_O[27] Tile_X9Y10_LUT4AB/FrameData_O[28] Tile_X9Y10_LUT4AB/FrameData_O[29]
+ Tile_X9Y10_LUT4AB/FrameData_O[2] Tile_X9Y10_LUT4AB/FrameData_O[30] Tile_X9Y10_LUT4AB/FrameData_O[31]
+ Tile_X9Y10_LUT4AB/FrameData_O[3] Tile_X9Y10_LUT4AB/FrameData_O[4] Tile_X9Y10_LUT4AB/FrameData_O[5]
+ Tile_X9Y10_LUT4AB/FrameData_O[6] Tile_X9Y10_LUT4AB/FrameData_O[7] Tile_X9Y10_LUT4AB/FrameData_O[8]
+ Tile_X9Y10_LUT4AB/FrameData_O[9] Tile_X10Y9_IHP_SRAM/Tile_X0Y1_FrameData_O[0] Tile_X10Y9_IHP_SRAM/Tile_X0Y1_FrameData_O[10]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y1_FrameData_O[11] Tile_X10Y9_IHP_SRAM/Tile_X0Y1_FrameData_O[12]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y1_FrameData_O[13] Tile_X10Y9_IHP_SRAM/Tile_X0Y1_FrameData_O[14]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y1_FrameData_O[15] Tile_X10Y9_IHP_SRAM/Tile_X0Y1_FrameData_O[16]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y1_FrameData_O[17] Tile_X10Y9_IHP_SRAM/Tile_X0Y1_FrameData_O[18]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y1_FrameData_O[19] Tile_X10Y9_IHP_SRAM/Tile_X0Y1_FrameData_O[1]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y1_FrameData_O[20] Tile_X10Y9_IHP_SRAM/Tile_X0Y1_FrameData_O[21]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y1_FrameData_O[22] Tile_X10Y9_IHP_SRAM/Tile_X0Y1_FrameData_O[23]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y1_FrameData_O[24] Tile_X10Y9_IHP_SRAM/Tile_X0Y1_FrameData_O[25]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y1_FrameData_O[26] Tile_X10Y9_IHP_SRAM/Tile_X0Y1_FrameData_O[27]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y1_FrameData_O[28] Tile_X10Y9_IHP_SRAM/Tile_X0Y1_FrameData_O[29]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y1_FrameData_O[2] Tile_X10Y9_IHP_SRAM/Tile_X0Y1_FrameData_O[30]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y1_FrameData_O[31] Tile_X10Y9_IHP_SRAM/Tile_X0Y1_FrameData_O[3]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y1_FrameData_O[4] Tile_X10Y9_IHP_SRAM/Tile_X0Y1_FrameData_O[5]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y1_FrameData_O[6] Tile_X10Y9_IHP_SRAM/Tile_X0Y1_FrameData_O[7]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y1_FrameData_O[8] Tile_X10Y9_IHP_SRAM/Tile_X0Y1_FrameData_O[9]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y1_FrameStrobe[0] Tile_X10Y9_IHP_SRAM/Tile_X0Y1_FrameStrobe[10]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y1_FrameStrobe[11] Tile_X10Y9_IHP_SRAM/Tile_X0Y1_FrameStrobe[12]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y1_FrameStrobe[13] Tile_X10Y9_IHP_SRAM/Tile_X0Y1_FrameStrobe[14]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y1_FrameStrobe[15] Tile_X10Y9_IHP_SRAM/Tile_X0Y1_FrameStrobe[16]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y1_FrameStrobe[17] Tile_X10Y9_IHP_SRAM/Tile_X0Y1_FrameStrobe[18]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y1_FrameStrobe[19] Tile_X10Y9_IHP_SRAM/Tile_X0Y1_FrameStrobe[1]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y1_FrameStrobe[2] Tile_X10Y9_IHP_SRAM/Tile_X0Y1_FrameStrobe[3]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y1_FrameStrobe[4] Tile_X10Y9_IHP_SRAM/Tile_X0Y1_FrameStrobe[5]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y1_FrameStrobe[6] Tile_X10Y9_IHP_SRAM/Tile_X0Y1_FrameStrobe[7]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y1_FrameStrobe[8] Tile_X10Y9_IHP_SRAM/Tile_X0Y1_FrameStrobe[9]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y1_N1END[0] Tile_X10Y9_IHP_SRAM/Tile_X0Y1_N1END[1] Tile_X10Y9_IHP_SRAM/Tile_X0Y1_N1END[2]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y1_N1END[3] Tile_X10Y9_IHP_SRAM/Tile_X0Y1_N2END[0] Tile_X10Y9_IHP_SRAM/Tile_X0Y1_N2END[1]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y1_N2END[2] Tile_X10Y9_IHP_SRAM/Tile_X0Y1_N2END[3] Tile_X10Y9_IHP_SRAM/Tile_X0Y1_N2END[4]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y1_N2END[5] Tile_X10Y9_IHP_SRAM/Tile_X0Y1_N2END[6] Tile_X10Y9_IHP_SRAM/Tile_X0Y1_N2END[7]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y1_N2MID[0] Tile_X10Y9_IHP_SRAM/Tile_X0Y1_N2MID[1] Tile_X10Y9_IHP_SRAM/Tile_X0Y1_N2MID[2]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y1_N2MID[3] Tile_X10Y9_IHP_SRAM/Tile_X0Y1_N2MID[4] Tile_X10Y9_IHP_SRAM/Tile_X0Y1_N2MID[5]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y1_N2MID[6] Tile_X10Y9_IHP_SRAM/Tile_X0Y1_N2MID[7] Tile_X10Y9_IHP_SRAM/Tile_X0Y1_N4END[0]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y1_N4END[10] Tile_X10Y9_IHP_SRAM/Tile_X0Y1_N4END[11]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y1_N4END[12] Tile_X10Y9_IHP_SRAM/Tile_X0Y1_N4END[13]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y1_N4END[14] Tile_X10Y9_IHP_SRAM/Tile_X0Y1_N4END[15]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y1_N4END[1] Tile_X10Y9_IHP_SRAM/Tile_X0Y1_N4END[2] Tile_X10Y9_IHP_SRAM/Tile_X0Y1_N4END[3]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y1_N4END[4] Tile_X10Y9_IHP_SRAM/Tile_X0Y1_N4END[5] Tile_X10Y9_IHP_SRAM/Tile_X0Y1_N4END[6]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y1_N4END[7] Tile_X10Y9_IHP_SRAM/Tile_X0Y1_N4END[8] Tile_X10Y9_IHP_SRAM/Tile_X0Y1_N4END[9]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y1_S1BEG[0] Tile_X10Y9_IHP_SRAM/Tile_X0Y1_S1BEG[1] Tile_X10Y9_IHP_SRAM/Tile_X0Y1_S1BEG[2]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y1_S1BEG[3] Tile_X10Y9_IHP_SRAM/Tile_X0Y1_S2BEG[0] Tile_X10Y9_IHP_SRAM/Tile_X0Y1_S2BEG[1]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y1_S2BEG[2] Tile_X10Y9_IHP_SRAM/Tile_X0Y1_S2BEG[3] Tile_X10Y9_IHP_SRAM/Tile_X0Y1_S2BEG[4]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y1_S2BEG[5] Tile_X10Y9_IHP_SRAM/Tile_X0Y1_S2BEG[6] Tile_X10Y9_IHP_SRAM/Tile_X0Y1_S2BEG[7]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y1_S2BEGb[0] Tile_X10Y9_IHP_SRAM/Tile_X0Y1_S2BEGb[1]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y1_S2BEGb[2] Tile_X10Y9_IHP_SRAM/Tile_X0Y1_S2BEGb[3]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y1_S2BEGb[4] Tile_X10Y9_IHP_SRAM/Tile_X0Y1_S2BEGb[5]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y1_S2BEGb[6] Tile_X10Y9_IHP_SRAM/Tile_X0Y1_S2BEGb[7]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y1_S4BEG[0] Tile_X10Y9_IHP_SRAM/Tile_X0Y1_S4BEG[10] Tile_X10Y9_IHP_SRAM/Tile_X0Y1_S4BEG[11]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y1_S4BEG[12] Tile_X10Y9_IHP_SRAM/Tile_X0Y1_S4BEG[13]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y1_S4BEG[14] Tile_X10Y9_IHP_SRAM/Tile_X0Y1_S4BEG[15]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y1_S4BEG[1] Tile_X10Y9_IHP_SRAM/Tile_X0Y1_S4BEG[2] Tile_X10Y9_IHP_SRAM/Tile_X0Y1_S4BEG[3]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y1_S4BEG[4] Tile_X10Y9_IHP_SRAM/Tile_X0Y1_S4BEG[5] Tile_X10Y9_IHP_SRAM/Tile_X0Y1_S4BEG[6]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y1_S4BEG[7] Tile_X10Y9_IHP_SRAM/Tile_X0Y1_S4BEG[8] Tile_X10Y9_IHP_SRAM/Tile_X0Y1_S4BEG[9]
+ Tile_X10Y9_IHP_SRAM/Tile_X0Y1_UserCLK Tile_X9Y10_LUT4AB/W1END[0] Tile_X9Y10_LUT4AB/W1END[1]
+ Tile_X9Y10_LUT4AB/W1END[2] Tile_X9Y10_LUT4AB/W1END[3] Tile_X9Y10_LUT4AB/W2MID[0]
+ Tile_X9Y10_LUT4AB/W2MID[1] Tile_X9Y10_LUT4AB/W2MID[2] Tile_X9Y10_LUT4AB/W2MID[3]
+ Tile_X9Y10_LUT4AB/W2MID[4] Tile_X9Y10_LUT4AB/W2MID[5] Tile_X9Y10_LUT4AB/W2MID[6]
+ Tile_X9Y10_LUT4AB/W2MID[7] Tile_X9Y10_LUT4AB/W2END[0] Tile_X9Y10_LUT4AB/W2END[1]
+ Tile_X9Y10_LUT4AB/W2END[2] Tile_X9Y10_LUT4AB/W2END[3] Tile_X9Y10_LUT4AB/W2END[4]
+ Tile_X9Y10_LUT4AB/W2END[5] Tile_X9Y10_LUT4AB/W2END[6] Tile_X9Y10_LUT4AB/W2END[7]
+ Tile_X9Y10_LUT4AB/W6END[0] Tile_X9Y10_LUT4AB/W6END[10] Tile_X9Y10_LUT4AB/W6END[11]
+ Tile_X9Y10_LUT4AB/W6END[1] Tile_X9Y10_LUT4AB/W6END[2] Tile_X9Y10_LUT4AB/W6END[3]
+ Tile_X9Y10_LUT4AB/W6END[4] Tile_X9Y10_LUT4AB/W6END[5] Tile_X9Y10_LUT4AB/W6END[6]
+ Tile_X9Y10_LUT4AB/W6END[7] Tile_X9Y10_LUT4AB/W6END[8] Tile_X9Y10_LUT4AB/W6END[9]
+ Tile_X9Y10_LUT4AB/WW4END[0] Tile_X9Y10_LUT4AB/WW4END[10] Tile_X9Y10_LUT4AB/WW4END[11]
+ Tile_X9Y10_LUT4AB/WW4END[12] Tile_X9Y10_LUT4AB/WW4END[13] Tile_X9Y10_LUT4AB/WW4END[14]
+ Tile_X9Y10_LUT4AB/WW4END[15] Tile_X9Y10_LUT4AB/WW4END[1] Tile_X9Y10_LUT4AB/WW4END[2]
+ Tile_X9Y10_LUT4AB/WW4END[3] Tile_X9Y10_LUT4AB/WW4END[4] Tile_X9Y10_LUT4AB/WW4END[5]
+ Tile_X9Y10_LUT4AB/WW4END[6] Tile_X9Y10_LUT4AB/WW4END[7] Tile_X9Y10_LUT4AB/WW4END[8]
+ Tile_X9Y10_LUT4AB/WW4END[9] VGND VPWR Tile_X10Y10_WEN_SRAM IHP_SRAM
XTile_X6Y0_N_term_single Tile_X6Y1_LUT4AB/Co Tile_X6Y0_N_term_single/FrameData[0]
+ Tile_X6Y0_N_term_single/FrameData[10] Tile_X6Y0_N_term_single/FrameData[11] Tile_X6Y0_N_term_single/FrameData[12]
+ Tile_X6Y0_N_term_single/FrameData[13] Tile_X6Y0_N_term_single/FrameData[14] Tile_X6Y0_N_term_single/FrameData[15]
+ Tile_X6Y0_N_term_single/FrameData[16] Tile_X6Y0_N_term_single/FrameData[17] Tile_X6Y0_N_term_single/FrameData[18]
+ Tile_X6Y0_N_term_single/FrameData[19] Tile_X6Y0_N_term_single/FrameData[1] Tile_X6Y0_N_term_single/FrameData[20]
+ Tile_X6Y0_N_term_single/FrameData[21] Tile_X6Y0_N_term_single/FrameData[22] Tile_X6Y0_N_term_single/FrameData[23]
+ Tile_X6Y0_N_term_single/FrameData[24] Tile_X6Y0_N_term_single/FrameData[25] Tile_X6Y0_N_term_single/FrameData[26]
+ Tile_X6Y0_N_term_single/FrameData[27] Tile_X6Y0_N_term_single/FrameData[28] Tile_X6Y0_N_term_single/FrameData[29]
+ Tile_X6Y0_N_term_single/FrameData[2] Tile_X6Y0_N_term_single/FrameData[30] Tile_X6Y0_N_term_single/FrameData[31]
+ Tile_X6Y0_N_term_single/FrameData[3] Tile_X6Y0_N_term_single/FrameData[4] Tile_X6Y0_N_term_single/FrameData[5]
+ Tile_X6Y0_N_term_single/FrameData[6] Tile_X6Y0_N_term_single/FrameData[7] Tile_X6Y0_N_term_single/FrameData[8]
+ Tile_X6Y0_N_term_single/FrameData[9] Tile_X7Y0_N_term_DSP/FrameData[0] Tile_X7Y0_N_term_DSP/FrameData[10]
+ Tile_X7Y0_N_term_DSP/FrameData[11] Tile_X7Y0_N_term_DSP/FrameData[12] Tile_X7Y0_N_term_DSP/FrameData[13]
+ Tile_X7Y0_N_term_DSP/FrameData[14] Tile_X7Y0_N_term_DSP/FrameData[15] Tile_X7Y0_N_term_DSP/FrameData[16]
+ Tile_X7Y0_N_term_DSP/FrameData[17] Tile_X7Y0_N_term_DSP/FrameData[18] Tile_X7Y0_N_term_DSP/FrameData[19]
+ Tile_X7Y0_N_term_DSP/FrameData[1] Tile_X7Y0_N_term_DSP/FrameData[20] Tile_X7Y0_N_term_DSP/FrameData[21]
+ Tile_X7Y0_N_term_DSP/FrameData[22] Tile_X7Y0_N_term_DSP/FrameData[23] Tile_X7Y0_N_term_DSP/FrameData[24]
+ Tile_X7Y0_N_term_DSP/FrameData[25] Tile_X7Y0_N_term_DSP/FrameData[26] Tile_X7Y0_N_term_DSP/FrameData[27]
+ Tile_X7Y0_N_term_DSP/FrameData[28] Tile_X7Y0_N_term_DSP/FrameData[29] Tile_X7Y0_N_term_DSP/FrameData[2]
+ Tile_X7Y0_N_term_DSP/FrameData[30] Tile_X7Y0_N_term_DSP/FrameData[31] Tile_X7Y0_N_term_DSP/FrameData[3]
+ Tile_X7Y0_N_term_DSP/FrameData[4] Tile_X7Y0_N_term_DSP/FrameData[5] Tile_X7Y0_N_term_DSP/FrameData[6]
+ Tile_X7Y0_N_term_DSP/FrameData[7] Tile_X7Y0_N_term_DSP/FrameData[8] Tile_X7Y0_N_term_DSP/FrameData[9]
+ Tile_X6Y1_LUT4AB/FrameStrobe_O[0] Tile_X6Y1_LUT4AB/FrameStrobe_O[10] Tile_X6Y1_LUT4AB/FrameStrobe_O[11]
+ Tile_X6Y1_LUT4AB/FrameStrobe_O[12] Tile_X6Y1_LUT4AB/FrameStrobe_O[13] Tile_X6Y1_LUT4AB/FrameStrobe_O[14]
+ Tile_X6Y1_LUT4AB/FrameStrobe_O[15] Tile_X6Y1_LUT4AB/FrameStrobe_O[16] Tile_X6Y1_LUT4AB/FrameStrobe_O[17]
+ Tile_X6Y1_LUT4AB/FrameStrobe_O[18] Tile_X6Y1_LUT4AB/FrameStrobe_O[19] Tile_X6Y1_LUT4AB/FrameStrobe_O[1]
+ Tile_X6Y1_LUT4AB/FrameStrobe_O[2] Tile_X6Y1_LUT4AB/FrameStrobe_O[3] Tile_X6Y1_LUT4AB/FrameStrobe_O[4]
+ Tile_X6Y1_LUT4AB/FrameStrobe_O[5] Tile_X6Y1_LUT4AB/FrameStrobe_O[6] Tile_X6Y1_LUT4AB/FrameStrobe_O[7]
+ Tile_X6Y1_LUT4AB/FrameStrobe_O[8] Tile_X6Y1_LUT4AB/FrameStrobe_O[9] Tile_X6Y0_N_term_single/FrameStrobe_O[0]
+ Tile_X6Y0_N_term_single/FrameStrobe_O[10] Tile_X6Y0_N_term_single/FrameStrobe_O[11]
+ Tile_X6Y0_N_term_single/FrameStrobe_O[12] Tile_X6Y0_N_term_single/FrameStrobe_O[13]
+ Tile_X6Y0_N_term_single/FrameStrobe_O[14] Tile_X6Y0_N_term_single/FrameStrobe_O[15]
+ Tile_X6Y0_N_term_single/FrameStrobe_O[16] Tile_X6Y0_N_term_single/FrameStrobe_O[17]
+ Tile_X6Y0_N_term_single/FrameStrobe_O[18] Tile_X6Y0_N_term_single/FrameStrobe_O[19]
+ Tile_X6Y0_N_term_single/FrameStrobe_O[1] Tile_X6Y0_N_term_single/FrameStrobe_O[2]
+ Tile_X6Y0_N_term_single/FrameStrobe_O[3] Tile_X6Y0_N_term_single/FrameStrobe_O[4]
+ Tile_X6Y0_N_term_single/FrameStrobe_O[5] Tile_X6Y0_N_term_single/FrameStrobe_O[6]
+ Tile_X6Y0_N_term_single/FrameStrobe_O[7] Tile_X6Y0_N_term_single/FrameStrobe_O[8]
+ Tile_X6Y0_N_term_single/FrameStrobe_O[9] Tile_X6Y1_LUT4AB/N1BEG[0] Tile_X6Y1_LUT4AB/N1BEG[1]
+ Tile_X6Y1_LUT4AB/N1BEG[2] Tile_X6Y1_LUT4AB/N1BEG[3] Tile_X6Y1_LUT4AB/N2BEGb[0] Tile_X6Y1_LUT4AB/N2BEGb[1]
+ Tile_X6Y1_LUT4AB/N2BEGb[2] Tile_X6Y1_LUT4AB/N2BEGb[3] Tile_X6Y1_LUT4AB/N2BEGb[4]
+ Tile_X6Y1_LUT4AB/N2BEGb[5] Tile_X6Y1_LUT4AB/N2BEGb[6] Tile_X6Y1_LUT4AB/N2BEGb[7]
+ Tile_X6Y1_LUT4AB/N2BEG[0] Tile_X6Y1_LUT4AB/N2BEG[1] Tile_X6Y1_LUT4AB/N2BEG[2] Tile_X6Y1_LUT4AB/N2BEG[3]
+ Tile_X6Y1_LUT4AB/N2BEG[4] Tile_X6Y1_LUT4AB/N2BEG[5] Tile_X6Y1_LUT4AB/N2BEG[6] Tile_X6Y1_LUT4AB/N2BEG[7]
+ Tile_X6Y1_LUT4AB/N4BEG[0] Tile_X6Y1_LUT4AB/N4BEG[10] Tile_X6Y1_LUT4AB/N4BEG[11]
+ Tile_X6Y1_LUT4AB/N4BEG[12] Tile_X6Y1_LUT4AB/N4BEG[13] Tile_X6Y1_LUT4AB/N4BEG[14]
+ Tile_X6Y1_LUT4AB/N4BEG[15] Tile_X6Y1_LUT4AB/N4BEG[1] Tile_X6Y1_LUT4AB/N4BEG[2] Tile_X6Y1_LUT4AB/N4BEG[3]
+ Tile_X6Y1_LUT4AB/N4BEG[4] Tile_X6Y1_LUT4AB/N4BEG[5] Tile_X6Y1_LUT4AB/N4BEG[6] Tile_X6Y1_LUT4AB/N4BEG[7]
+ Tile_X6Y1_LUT4AB/N4BEG[8] Tile_X6Y1_LUT4AB/N4BEG[9] Tile_X6Y1_LUT4AB/NN4BEG[0] Tile_X6Y1_LUT4AB/NN4BEG[10]
+ Tile_X6Y1_LUT4AB/NN4BEG[11] Tile_X6Y1_LUT4AB/NN4BEG[12] Tile_X6Y1_LUT4AB/NN4BEG[13]
+ Tile_X6Y1_LUT4AB/NN4BEG[14] Tile_X6Y1_LUT4AB/NN4BEG[15] Tile_X6Y1_LUT4AB/NN4BEG[1]
+ Tile_X6Y1_LUT4AB/NN4BEG[2] Tile_X6Y1_LUT4AB/NN4BEG[3] Tile_X6Y1_LUT4AB/NN4BEG[4]
+ Tile_X6Y1_LUT4AB/NN4BEG[5] Tile_X6Y1_LUT4AB/NN4BEG[6] Tile_X6Y1_LUT4AB/NN4BEG[7]
+ Tile_X6Y1_LUT4AB/NN4BEG[8] Tile_X6Y1_LUT4AB/NN4BEG[9] Tile_X6Y1_LUT4AB/S1END[0]
+ Tile_X6Y1_LUT4AB/S1END[1] Tile_X6Y1_LUT4AB/S1END[2] Tile_X6Y1_LUT4AB/S1END[3] Tile_X6Y1_LUT4AB/S2MID[0]
+ Tile_X6Y1_LUT4AB/S2MID[1] Tile_X6Y1_LUT4AB/S2MID[2] Tile_X6Y1_LUT4AB/S2MID[3] Tile_X6Y1_LUT4AB/S2MID[4]
+ Tile_X6Y1_LUT4AB/S2MID[5] Tile_X6Y1_LUT4AB/S2MID[6] Tile_X6Y1_LUT4AB/S2MID[7] Tile_X6Y1_LUT4AB/S2END[0]
+ Tile_X6Y1_LUT4AB/S2END[1] Tile_X6Y1_LUT4AB/S2END[2] Tile_X6Y1_LUT4AB/S2END[3] Tile_X6Y1_LUT4AB/S2END[4]
+ Tile_X6Y1_LUT4AB/S2END[5] Tile_X6Y1_LUT4AB/S2END[6] Tile_X6Y1_LUT4AB/S2END[7] Tile_X6Y1_LUT4AB/S4END[0]
+ Tile_X6Y1_LUT4AB/S4END[10] Tile_X6Y1_LUT4AB/S4END[11] Tile_X6Y1_LUT4AB/S4END[12]
+ Tile_X6Y1_LUT4AB/S4END[13] Tile_X6Y1_LUT4AB/S4END[14] Tile_X6Y1_LUT4AB/S4END[15]
+ Tile_X6Y1_LUT4AB/S4END[1] Tile_X6Y1_LUT4AB/S4END[2] Tile_X6Y1_LUT4AB/S4END[3] Tile_X6Y1_LUT4AB/S4END[4]
+ Tile_X6Y1_LUT4AB/S4END[5] Tile_X6Y1_LUT4AB/S4END[6] Tile_X6Y1_LUT4AB/S4END[7] Tile_X6Y1_LUT4AB/S4END[8]
+ Tile_X6Y1_LUT4AB/S4END[9] Tile_X6Y1_LUT4AB/SS4END[0] Tile_X6Y1_LUT4AB/SS4END[10]
+ Tile_X6Y1_LUT4AB/SS4END[11] Tile_X6Y1_LUT4AB/SS4END[12] Tile_X6Y1_LUT4AB/SS4END[13]
+ Tile_X6Y1_LUT4AB/SS4END[14] Tile_X6Y1_LUT4AB/SS4END[15] Tile_X6Y1_LUT4AB/SS4END[1]
+ Tile_X6Y1_LUT4AB/SS4END[2] Tile_X6Y1_LUT4AB/SS4END[3] Tile_X6Y1_LUT4AB/SS4END[4]
+ Tile_X6Y1_LUT4AB/SS4END[5] Tile_X6Y1_LUT4AB/SS4END[6] Tile_X6Y1_LUT4AB/SS4END[7]
+ Tile_X6Y1_LUT4AB/SS4END[8] Tile_X6Y1_LUT4AB/SS4END[9] Tile_X6Y1_LUT4AB/UserCLKo
+ Tile_X6Y0_N_term_single/UserCLKo VGND VPWR N_term_single
XTile_X0Y14_W_IO Tile_X0Y14_A_I_top Tile_X0Y14_A_O_top Tile_X0Y14_A_T_top Tile_X0Y14_A_config_C_bit0
+ Tile_X0Y14_A_config_C_bit1 Tile_X0Y14_A_config_C_bit2 Tile_X0Y14_A_config_C_bit3
+ Tile_X0Y14_B_I_top Tile_X0Y14_B_O_top Tile_X0Y14_B_T_top Tile_X0Y14_B_config_C_bit0
+ Tile_X0Y14_B_config_C_bit1 Tile_X0Y14_B_config_C_bit2 Tile_X0Y14_B_config_C_bit3
+ Tile_X0Y14_W_IO/E1BEG[0] Tile_X0Y14_W_IO/E1BEG[1] Tile_X0Y14_W_IO/E1BEG[2] Tile_X0Y14_W_IO/E1BEG[3]
+ Tile_X0Y14_W_IO/E2BEG[0] Tile_X0Y14_W_IO/E2BEG[1] Tile_X0Y14_W_IO/E2BEG[2] Tile_X0Y14_W_IO/E2BEG[3]
+ Tile_X0Y14_W_IO/E2BEG[4] Tile_X0Y14_W_IO/E2BEG[5] Tile_X0Y14_W_IO/E2BEG[6] Tile_X0Y14_W_IO/E2BEG[7]
+ Tile_X0Y14_W_IO/E2BEGb[0] Tile_X0Y14_W_IO/E2BEGb[1] Tile_X0Y14_W_IO/E2BEGb[2] Tile_X0Y14_W_IO/E2BEGb[3]
+ Tile_X0Y14_W_IO/E2BEGb[4] Tile_X0Y14_W_IO/E2BEGb[5] Tile_X0Y14_W_IO/E2BEGb[6] Tile_X0Y14_W_IO/E2BEGb[7]
+ Tile_X0Y14_W_IO/E6BEG[0] Tile_X0Y14_W_IO/E6BEG[10] Tile_X0Y14_W_IO/E6BEG[11] Tile_X0Y14_W_IO/E6BEG[1]
+ Tile_X0Y14_W_IO/E6BEG[2] Tile_X0Y14_W_IO/E6BEG[3] Tile_X0Y14_W_IO/E6BEG[4] Tile_X0Y14_W_IO/E6BEG[5]
+ Tile_X0Y14_W_IO/E6BEG[6] Tile_X0Y14_W_IO/E6BEG[7] Tile_X0Y14_W_IO/E6BEG[8] Tile_X0Y14_W_IO/E6BEG[9]
+ Tile_X0Y14_W_IO/EE4BEG[0] Tile_X0Y14_W_IO/EE4BEG[10] Tile_X0Y14_W_IO/EE4BEG[11]
+ Tile_X0Y14_W_IO/EE4BEG[12] Tile_X0Y14_W_IO/EE4BEG[13] Tile_X0Y14_W_IO/EE4BEG[14]
+ Tile_X0Y14_W_IO/EE4BEG[15] Tile_X0Y14_W_IO/EE4BEG[1] Tile_X0Y14_W_IO/EE4BEG[2] Tile_X0Y14_W_IO/EE4BEG[3]
+ Tile_X0Y14_W_IO/EE4BEG[4] Tile_X0Y14_W_IO/EE4BEG[5] Tile_X0Y14_W_IO/EE4BEG[6] Tile_X0Y14_W_IO/EE4BEG[7]
+ Tile_X0Y14_W_IO/EE4BEG[8] Tile_X0Y14_W_IO/EE4BEG[9] FrameData[448] FrameData[458]
+ FrameData[459] FrameData[460] FrameData[461] FrameData[462] FrameData[463] FrameData[464]
+ FrameData[465] FrameData[466] FrameData[467] FrameData[449] FrameData[468] FrameData[469]
+ FrameData[470] FrameData[471] FrameData[472] FrameData[473] FrameData[474] FrameData[475]
+ FrameData[476] FrameData[477] FrameData[450] FrameData[478] FrameData[479] FrameData[451]
+ FrameData[452] FrameData[453] FrameData[454] FrameData[455] FrameData[456] FrameData[457]
+ Tile_X1Y14_LUT4AB/FrameData[0] Tile_X1Y14_LUT4AB/FrameData[10] Tile_X1Y14_LUT4AB/FrameData[11]
+ Tile_X1Y14_LUT4AB/FrameData[12] Tile_X1Y14_LUT4AB/FrameData[13] Tile_X1Y14_LUT4AB/FrameData[14]
+ Tile_X1Y14_LUT4AB/FrameData[15] Tile_X1Y14_LUT4AB/FrameData[16] Tile_X1Y14_LUT4AB/FrameData[17]
+ Tile_X1Y14_LUT4AB/FrameData[18] Tile_X1Y14_LUT4AB/FrameData[19] Tile_X1Y14_LUT4AB/FrameData[1]
+ Tile_X1Y14_LUT4AB/FrameData[20] Tile_X1Y14_LUT4AB/FrameData[21] Tile_X1Y14_LUT4AB/FrameData[22]
+ Tile_X1Y14_LUT4AB/FrameData[23] Tile_X1Y14_LUT4AB/FrameData[24] Tile_X1Y14_LUT4AB/FrameData[25]
+ Tile_X1Y14_LUT4AB/FrameData[26] Tile_X1Y14_LUT4AB/FrameData[27] Tile_X1Y14_LUT4AB/FrameData[28]
+ Tile_X1Y14_LUT4AB/FrameData[29] Tile_X1Y14_LUT4AB/FrameData[2] Tile_X1Y14_LUT4AB/FrameData[30]
+ Tile_X1Y14_LUT4AB/FrameData[31] Tile_X1Y14_LUT4AB/FrameData[3] Tile_X1Y14_LUT4AB/FrameData[4]
+ Tile_X1Y14_LUT4AB/FrameData[5] Tile_X1Y14_LUT4AB/FrameData[6] Tile_X1Y14_LUT4AB/FrameData[7]
+ Tile_X1Y14_LUT4AB/FrameData[8] Tile_X1Y14_LUT4AB/FrameData[9] FrameStrobe[0] FrameStrobe[10]
+ FrameStrobe[11] FrameStrobe[12] FrameStrobe[13] FrameStrobe[14] FrameStrobe[15]
+ FrameStrobe[16] FrameStrobe[17] FrameStrobe[18] FrameStrobe[19] FrameStrobe[1] FrameStrobe[2]
+ FrameStrobe[3] FrameStrobe[4] FrameStrobe[5] FrameStrobe[6] FrameStrobe[7] FrameStrobe[8]
+ FrameStrobe[9] Tile_X0Y13_W_IO/FrameStrobe[0] Tile_X0Y13_W_IO/FrameStrobe[10] Tile_X0Y13_W_IO/FrameStrobe[11]
+ Tile_X0Y13_W_IO/FrameStrobe[12] Tile_X0Y13_W_IO/FrameStrobe[13] Tile_X0Y13_W_IO/FrameStrobe[14]
+ Tile_X0Y13_W_IO/FrameStrobe[15] Tile_X0Y13_W_IO/FrameStrobe[16] Tile_X0Y13_W_IO/FrameStrobe[17]
+ Tile_X0Y13_W_IO/FrameStrobe[18] Tile_X0Y13_W_IO/FrameStrobe[19] Tile_X0Y13_W_IO/FrameStrobe[1]
+ Tile_X0Y13_W_IO/FrameStrobe[2] Tile_X0Y13_W_IO/FrameStrobe[3] Tile_X0Y13_W_IO/FrameStrobe[4]
+ Tile_X0Y13_W_IO/FrameStrobe[5] Tile_X0Y13_W_IO/FrameStrobe[6] Tile_X0Y13_W_IO/FrameStrobe[7]
+ Tile_X0Y13_W_IO/FrameStrobe[8] Tile_X0Y13_W_IO/FrameStrobe[9] UserCLK Tile_X0Y13_W_IO/UserCLK
+ VGND VPWR Tile_X0Y14_W_IO/W1END[0] Tile_X0Y14_W_IO/W1END[1] Tile_X0Y14_W_IO/W1END[2]
+ Tile_X0Y14_W_IO/W1END[3] Tile_X0Y14_W_IO/W2END[0] Tile_X0Y14_W_IO/W2END[1] Tile_X0Y14_W_IO/W2END[2]
+ Tile_X0Y14_W_IO/W2END[3] Tile_X0Y14_W_IO/W2END[4] Tile_X0Y14_W_IO/W2END[5] Tile_X0Y14_W_IO/W2END[6]
+ Tile_X0Y14_W_IO/W2END[7] Tile_X0Y14_W_IO/W2MID[0] Tile_X0Y14_W_IO/W2MID[1] Tile_X0Y14_W_IO/W2MID[2]
+ Tile_X0Y14_W_IO/W2MID[3] Tile_X0Y14_W_IO/W2MID[4] Tile_X0Y14_W_IO/W2MID[5] Tile_X0Y14_W_IO/W2MID[6]
+ Tile_X0Y14_W_IO/W2MID[7] Tile_X0Y14_W_IO/W6END[0] Tile_X0Y14_W_IO/W6END[10] Tile_X0Y14_W_IO/W6END[11]
+ Tile_X0Y14_W_IO/W6END[1] Tile_X0Y14_W_IO/W6END[2] Tile_X0Y14_W_IO/W6END[3] Tile_X0Y14_W_IO/W6END[4]
+ Tile_X0Y14_W_IO/W6END[5] Tile_X0Y14_W_IO/W6END[6] Tile_X0Y14_W_IO/W6END[7] Tile_X0Y14_W_IO/W6END[8]
+ Tile_X0Y14_W_IO/W6END[9] Tile_X0Y14_W_IO/WW4END[0] Tile_X0Y14_W_IO/WW4END[10] Tile_X0Y14_W_IO/WW4END[11]
+ Tile_X0Y14_W_IO/WW4END[12] Tile_X0Y14_W_IO/WW4END[13] Tile_X0Y14_W_IO/WW4END[14]
+ Tile_X0Y14_W_IO/WW4END[15] Tile_X0Y14_W_IO/WW4END[1] Tile_X0Y14_W_IO/WW4END[2] Tile_X0Y14_W_IO/WW4END[3]
+ Tile_X0Y14_W_IO/WW4END[4] Tile_X0Y14_W_IO/WW4END[5] Tile_X0Y14_W_IO/WW4END[6] Tile_X0Y14_W_IO/WW4END[7]
+ Tile_X0Y14_W_IO/WW4END[8] Tile_X0Y14_W_IO/WW4END[9] W_IO
XTile_X3Y10_LUT4AB Tile_X3Y11_LUT4AB/Co Tile_X3Y9_LUT4AB/Ci Tile_X3Y10_LUT4AB/E1BEG[0]
+ Tile_X3Y10_LUT4AB/E1BEG[1] Tile_X3Y10_LUT4AB/E1BEG[2] Tile_X3Y10_LUT4AB/E1BEG[3]
+ Tile_X3Y10_LUT4AB/E1END[0] Tile_X3Y10_LUT4AB/E1END[1] Tile_X3Y10_LUT4AB/E1END[2]
+ Tile_X3Y10_LUT4AB/E1END[3] Tile_X3Y10_LUT4AB/E2BEG[0] Tile_X3Y10_LUT4AB/E2BEG[1]
+ Tile_X3Y10_LUT4AB/E2BEG[2] Tile_X3Y10_LUT4AB/E2BEG[3] Tile_X3Y10_LUT4AB/E2BEG[4]
+ Tile_X3Y10_LUT4AB/E2BEG[5] Tile_X3Y10_LUT4AB/E2BEG[6] Tile_X3Y10_LUT4AB/E2BEG[7]
+ Tile_X4Y10_RegFile/E2END[0] Tile_X4Y10_RegFile/E2END[1] Tile_X4Y10_RegFile/E2END[2]
+ Tile_X4Y10_RegFile/E2END[3] Tile_X4Y10_RegFile/E2END[4] Tile_X4Y10_RegFile/E2END[5]
+ Tile_X4Y10_RegFile/E2END[6] Tile_X4Y10_RegFile/E2END[7] Tile_X3Y10_LUT4AB/E2END[0]
+ Tile_X3Y10_LUT4AB/E2END[1] Tile_X3Y10_LUT4AB/E2END[2] Tile_X3Y10_LUT4AB/E2END[3]
+ Tile_X3Y10_LUT4AB/E2END[4] Tile_X3Y10_LUT4AB/E2END[5] Tile_X3Y10_LUT4AB/E2END[6]
+ Tile_X3Y10_LUT4AB/E2END[7] Tile_X3Y10_LUT4AB/E2MID[0] Tile_X3Y10_LUT4AB/E2MID[1]
+ Tile_X3Y10_LUT4AB/E2MID[2] Tile_X3Y10_LUT4AB/E2MID[3] Tile_X3Y10_LUT4AB/E2MID[4]
+ Tile_X3Y10_LUT4AB/E2MID[5] Tile_X3Y10_LUT4AB/E2MID[6] Tile_X3Y10_LUT4AB/E2MID[7]
+ Tile_X3Y10_LUT4AB/E6BEG[0] Tile_X3Y10_LUT4AB/E6BEG[10] Tile_X3Y10_LUT4AB/E6BEG[11]
+ Tile_X3Y10_LUT4AB/E6BEG[1] Tile_X3Y10_LUT4AB/E6BEG[2] Tile_X3Y10_LUT4AB/E6BEG[3]
+ Tile_X3Y10_LUT4AB/E6BEG[4] Tile_X3Y10_LUT4AB/E6BEG[5] Tile_X3Y10_LUT4AB/E6BEG[6]
+ Tile_X3Y10_LUT4AB/E6BEG[7] Tile_X3Y10_LUT4AB/E6BEG[8] Tile_X3Y10_LUT4AB/E6BEG[9]
+ Tile_X3Y10_LUT4AB/E6END[0] Tile_X3Y10_LUT4AB/E6END[10] Tile_X3Y10_LUT4AB/E6END[11]
+ Tile_X3Y10_LUT4AB/E6END[1] Tile_X3Y10_LUT4AB/E6END[2] Tile_X3Y10_LUT4AB/E6END[3]
+ Tile_X3Y10_LUT4AB/E6END[4] Tile_X3Y10_LUT4AB/E6END[5] Tile_X3Y10_LUT4AB/E6END[6]
+ Tile_X3Y10_LUT4AB/E6END[7] Tile_X3Y10_LUT4AB/E6END[8] Tile_X3Y10_LUT4AB/E6END[9]
+ Tile_X3Y10_LUT4AB/EE4BEG[0] Tile_X3Y10_LUT4AB/EE4BEG[10] Tile_X3Y10_LUT4AB/EE4BEG[11]
+ Tile_X3Y10_LUT4AB/EE4BEG[12] Tile_X3Y10_LUT4AB/EE4BEG[13] Tile_X3Y10_LUT4AB/EE4BEG[14]
+ Tile_X3Y10_LUT4AB/EE4BEG[15] Tile_X3Y10_LUT4AB/EE4BEG[1] Tile_X3Y10_LUT4AB/EE4BEG[2]
+ Tile_X3Y10_LUT4AB/EE4BEG[3] Tile_X3Y10_LUT4AB/EE4BEG[4] Tile_X3Y10_LUT4AB/EE4BEG[5]
+ Tile_X3Y10_LUT4AB/EE4BEG[6] Tile_X3Y10_LUT4AB/EE4BEG[7] Tile_X3Y10_LUT4AB/EE4BEG[8]
+ Tile_X3Y10_LUT4AB/EE4BEG[9] Tile_X3Y10_LUT4AB/EE4END[0] Tile_X3Y10_LUT4AB/EE4END[10]
+ Tile_X3Y10_LUT4AB/EE4END[11] Tile_X3Y10_LUT4AB/EE4END[12] Tile_X3Y10_LUT4AB/EE4END[13]
+ Tile_X3Y10_LUT4AB/EE4END[14] Tile_X3Y10_LUT4AB/EE4END[15] Tile_X3Y10_LUT4AB/EE4END[1]
+ Tile_X3Y10_LUT4AB/EE4END[2] Tile_X3Y10_LUT4AB/EE4END[3] Tile_X3Y10_LUT4AB/EE4END[4]
+ Tile_X3Y10_LUT4AB/EE4END[5] Tile_X3Y10_LUT4AB/EE4END[6] Tile_X3Y10_LUT4AB/EE4END[7]
+ Tile_X3Y10_LUT4AB/EE4END[8] Tile_X3Y10_LUT4AB/EE4END[9] Tile_X3Y10_LUT4AB/FrameData[0]
+ Tile_X3Y10_LUT4AB/FrameData[10] Tile_X3Y10_LUT4AB/FrameData[11] Tile_X3Y10_LUT4AB/FrameData[12]
+ Tile_X3Y10_LUT4AB/FrameData[13] Tile_X3Y10_LUT4AB/FrameData[14] Tile_X3Y10_LUT4AB/FrameData[15]
+ Tile_X3Y10_LUT4AB/FrameData[16] Tile_X3Y10_LUT4AB/FrameData[17] Tile_X3Y10_LUT4AB/FrameData[18]
+ Tile_X3Y10_LUT4AB/FrameData[19] Tile_X3Y10_LUT4AB/FrameData[1] Tile_X3Y10_LUT4AB/FrameData[20]
+ Tile_X3Y10_LUT4AB/FrameData[21] Tile_X3Y10_LUT4AB/FrameData[22] Tile_X3Y10_LUT4AB/FrameData[23]
+ Tile_X3Y10_LUT4AB/FrameData[24] Tile_X3Y10_LUT4AB/FrameData[25] Tile_X3Y10_LUT4AB/FrameData[26]
+ Tile_X3Y10_LUT4AB/FrameData[27] Tile_X3Y10_LUT4AB/FrameData[28] Tile_X3Y10_LUT4AB/FrameData[29]
+ Tile_X3Y10_LUT4AB/FrameData[2] Tile_X3Y10_LUT4AB/FrameData[30] Tile_X3Y10_LUT4AB/FrameData[31]
+ Tile_X3Y10_LUT4AB/FrameData[3] Tile_X3Y10_LUT4AB/FrameData[4] Tile_X3Y10_LUT4AB/FrameData[5]
+ Tile_X3Y10_LUT4AB/FrameData[6] Tile_X3Y10_LUT4AB/FrameData[7] Tile_X3Y10_LUT4AB/FrameData[8]
+ Tile_X3Y10_LUT4AB/FrameData[9] Tile_X4Y10_RegFile/FrameData[0] Tile_X4Y10_RegFile/FrameData[10]
+ Tile_X4Y10_RegFile/FrameData[11] Tile_X4Y10_RegFile/FrameData[12] Tile_X4Y10_RegFile/FrameData[13]
+ Tile_X4Y10_RegFile/FrameData[14] Tile_X4Y10_RegFile/FrameData[15] Tile_X4Y10_RegFile/FrameData[16]
+ Tile_X4Y10_RegFile/FrameData[17] Tile_X4Y10_RegFile/FrameData[18] Tile_X4Y10_RegFile/FrameData[19]
+ Tile_X4Y10_RegFile/FrameData[1] Tile_X4Y10_RegFile/FrameData[20] Tile_X4Y10_RegFile/FrameData[21]
+ Tile_X4Y10_RegFile/FrameData[22] Tile_X4Y10_RegFile/FrameData[23] Tile_X4Y10_RegFile/FrameData[24]
+ Tile_X4Y10_RegFile/FrameData[25] Tile_X4Y10_RegFile/FrameData[26] Tile_X4Y10_RegFile/FrameData[27]
+ Tile_X4Y10_RegFile/FrameData[28] Tile_X4Y10_RegFile/FrameData[29] Tile_X4Y10_RegFile/FrameData[2]
+ Tile_X4Y10_RegFile/FrameData[30] Tile_X4Y10_RegFile/FrameData[31] Tile_X4Y10_RegFile/FrameData[3]
+ Tile_X4Y10_RegFile/FrameData[4] Tile_X4Y10_RegFile/FrameData[5] Tile_X4Y10_RegFile/FrameData[6]
+ Tile_X4Y10_RegFile/FrameData[7] Tile_X4Y10_RegFile/FrameData[8] Tile_X4Y10_RegFile/FrameData[9]
+ Tile_X3Y10_LUT4AB/FrameStrobe[0] Tile_X3Y10_LUT4AB/FrameStrobe[10] Tile_X3Y10_LUT4AB/FrameStrobe[11]
+ Tile_X3Y10_LUT4AB/FrameStrobe[12] Tile_X3Y10_LUT4AB/FrameStrobe[13] Tile_X3Y10_LUT4AB/FrameStrobe[14]
+ Tile_X3Y10_LUT4AB/FrameStrobe[15] Tile_X3Y10_LUT4AB/FrameStrobe[16] Tile_X3Y10_LUT4AB/FrameStrobe[17]
+ Tile_X3Y10_LUT4AB/FrameStrobe[18] Tile_X3Y10_LUT4AB/FrameStrobe[19] Tile_X3Y10_LUT4AB/FrameStrobe[1]
+ Tile_X3Y10_LUT4AB/FrameStrobe[2] Tile_X3Y10_LUT4AB/FrameStrobe[3] Tile_X3Y10_LUT4AB/FrameStrobe[4]
+ Tile_X3Y10_LUT4AB/FrameStrobe[5] Tile_X3Y10_LUT4AB/FrameStrobe[6] Tile_X3Y10_LUT4AB/FrameStrobe[7]
+ Tile_X3Y10_LUT4AB/FrameStrobe[8] Tile_X3Y10_LUT4AB/FrameStrobe[9] Tile_X3Y9_LUT4AB/FrameStrobe[0]
+ Tile_X3Y9_LUT4AB/FrameStrobe[10] Tile_X3Y9_LUT4AB/FrameStrobe[11] Tile_X3Y9_LUT4AB/FrameStrobe[12]
+ Tile_X3Y9_LUT4AB/FrameStrobe[13] Tile_X3Y9_LUT4AB/FrameStrobe[14] Tile_X3Y9_LUT4AB/FrameStrobe[15]
+ Tile_X3Y9_LUT4AB/FrameStrobe[16] Tile_X3Y9_LUT4AB/FrameStrobe[17] Tile_X3Y9_LUT4AB/FrameStrobe[18]
+ Tile_X3Y9_LUT4AB/FrameStrobe[19] Tile_X3Y9_LUT4AB/FrameStrobe[1] Tile_X3Y9_LUT4AB/FrameStrobe[2]
+ Tile_X3Y9_LUT4AB/FrameStrobe[3] Tile_X3Y9_LUT4AB/FrameStrobe[4] Tile_X3Y9_LUT4AB/FrameStrobe[5]
+ Tile_X3Y9_LUT4AB/FrameStrobe[6] Tile_X3Y9_LUT4AB/FrameStrobe[7] Tile_X3Y9_LUT4AB/FrameStrobe[8]
+ Tile_X3Y9_LUT4AB/FrameStrobe[9] Tile_X3Y9_LUT4AB/N1END[0] Tile_X3Y9_LUT4AB/N1END[1]
+ Tile_X3Y9_LUT4AB/N1END[2] Tile_X3Y9_LUT4AB/N1END[3] Tile_X3Y11_LUT4AB/N1BEG[0] Tile_X3Y11_LUT4AB/N1BEG[1]
+ Tile_X3Y11_LUT4AB/N1BEG[2] Tile_X3Y11_LUT4AB/N1BEG[3] Tile_X3Y9_LUT4AB/N2MID[0]
+ Tile_X3Y9_LUT4AB/N2MID[1] Tile_X3Y9_LUT4AB/N2MID[2] Tile_X3Y9_LUT4AB/N2MID[3] Tile_X3Y9_LUT4AB/N2MID[4]
+ Tile_X3Y9_LUT4AB/N2MID[5] Tile_X3Y9_LUT4AB/N2MID[6] Tile_X3Y9_LUT4AB/N2MID[7] Tile_X3Y9_LUT4AB/N2END[0]
+ Tile_X3Y9_LUT4AB/N2END[1] Tile_X3Y9_LUT4AB/N2END[2] Tile_X3Y9_LUT4AB/N2END[3] Tile_X3Y9_LUT4AB/N2END[4]
+ Tile_X3Y9_LUT4AB/N2END[5] Tile_X3Y9_LUT4AB/N2END[6] Tile_X3Y9_LUT4AB/N2END[7] Tile_X3Y10_LUT4AB/N2END[0]
+ Tile_X3Y10_LUT4AB/N2END[1] Tile_X3Y10_LUT4AB/N2END[2] Tile_X3Y10_LUT4AB/N2END[3]
+ Tile_X3Y10_LUT4AB/N2END[4] Tile_X3Y10_LUT4AB/N2END[5] Tile_X3Y10_LUT4AB/N2END[6]
+ Tile_X3Y10_LUT4AB/N2END[7] Tile_X3Y11_LUT4AB/N2BEG[0] Tile_X3Y11_LUT4AB/N2BEG[1]
+ Tile_X3Y11_LUT4AB/N2BEG[2] Tile_X3Y11_LUT4AB/N2BEG[3] Tile_X3Y11_LUT4AB/N2BEG[4]
+ Tile_X3Y11_LUT4AB/N2BEG[5] Tile_X3Y11_LUT4AB/N2BEG[6] Tile_X3Y11_LUT4AB/N2BEG[7]
+ Tile_X3Y9_LUT4AB/N4END[0] Tile_X3Y9_LUT4AB/N4END[10] Tile_X3Y9_LUT4AB/N4END[11]
+ Tile_X3Y9_LUT4AB/N4END[12] Tile_X3Y9_LUT4AB/N4END[13] Tile_X3Y9_LUT4AB/N4END[14]
+ Tile_X3Y9_LUT4AB/N4END[15] Tile_X3Y9_LUT4AB/N4END[1] Tile_X3Y9_LUT4AB/N4END[2] Tile_X3Y9_LUT4AB/N4END[3]
+ Tile_X3Y9_LUT4AB/N4END[4] Tile_X3Y9_LUT4AB/N4END[5] Tile_X3Y9_LUT4AB/N4END[6] Tile_X3Y9_LUT4AB/N4END[7]
+ Tile_X3Y9_LUT4AB/N4END[8] Tile_X3Y9_LUT4AB/N4END[9] Tile_X3Y11_LUT4AB/N4BEG[0] Tile_X3Y11_LUT4AB/N4BEG[10]
+ Tile_X3Y11_LUT4AB/N4BEG[11] Tile_X3Y11_LUT4AB/N4BEG[12] Tile_X3Y11_LUT4AB/N4BEG[13]
+ Tile_X3Y11_LUT4AB/N4BEG[14] Tile_X3Y11_LUT4AB/N4BEG[15] Tile_X3Y11_LUT4AB/N4BEG[1]
+ Tile_X3Y11_LUT4AB/N4BEG[2] Tile_X3Y11_LUT4AB/N4BEG[3] Tile_X3Y11_LUT4AB/N4BEG[4]
+ Tile_X3Y11_LUT4AB/N4BEG[5] Tile_X3Y11_LUT4AB/N4BEG[6] Tile_X3Y11_LUT4AB/N4BEG[7]
+ Tile_X3Y11_LUT4AB/N4BEG[8] Tile_X3Y11_LUT4AB/N4BEG[9] Tile_X3Y9_LUT4AB/NN4END[0]
+ Tile_X3Y9_LUT4AB/NN4END[10] Tile_X3Y9_LUT4AB/NN4END[11] Tile_X3Y9_LUT4AB/NN4END[12]
+ Tile_X3Y9_LUT4AB/NN4END[13] Tile_X3Y9_LUT4AB/NN4END[14] Tile_X3Y9_LUT4AB/NN4END[15]
+ Tile_X3Y9_LUT4AB/NN4END[1] Tile_X3Y9_LUT4AB/NN4END[2] Tile_X3Y9_LUT4AB/NN4END[3]
+ Tile_X3Y9_LUT4AB/NN4END[4] Tile_X3Y9_LUT4AB/NN4END[5] Tile_X3Y9_LUT4AB/NN4END[6]
+ Tile_X3Y9_LUT4AB/NN4END[7] Tile_X3Y9_LUT4AB/NN4END[8] Tile_X3Y9_LUT4AB/NN4END[9]
+ Tile_X3Y11_LUT4AB/NN4BEG[0] Tile_X3Y11_LUT4AB/NN4BEG[10] Tile_X3Y11_LUT4AB/NN4BEG[11]
+ Tile_X3Y11_LUT4AB/NN4BEG[12] Tile_X3Y11_LUT4AB/NN4BEG[13] Tile_X3Y11_LUT4AB/NN4BEG[14]
+ Tile_X3Y11_LUT4AB/NN4BEG[15] Tile_X3Y11_LUT4AB/NN4BEG[1] Tile_X3Y11_LUT4AB/NN4BEG[2]
+ Tile_X3Y11_LUT4AB/NN4BEG[3] Tile_X3Y11_LUT4AB/NN4BEG[4] Tile_X3Y11_LUT4AB/NN4BEG[5]
+ Tile_X3Y11_LUT4AB/NN4BEG[6] Tile_X3Y11_LUT4AB/NN4BEG[7] Tile_X3Y11_LUT4AB/NN4BEG[8]
+ Tile_X3Y11_LUT4AB/NN4BEG[9] Tile_X3Y11_LUT4AB/S1END[0] Tile_X3Y11_LUT4AB/S1END[1]
+ Tile_X3Y11_LUT4AB/S1END[2] Tile_X3Y11_LUT4AB/S1END[3] Tile_X3Y9_LUT4AB/S1BEG[0]
+ Tile_X3Y9_LUT4AB/S1BEG[1] Tile_X3Y9_LUT4AB/S1BEG[2] Tile_X3Y9_LUT4AB/S1BEG[3] Tile_X3Y11_LUT4AB/S2MID[0]
+ Tile_X3Y11_LUT4AB/S2MID[1] Tile_X3Y11_LUT4AB/S2MID[2] Tile_X3Y11_LUT4AB/S2MID[3]
+ Tile_X3Y11_LUT4AB/S2MID[4] Tile_X3Y11_LUT4AB/S2MID[5] Tile_X3Y11_LUT4AB/S2MID[6]
+ Tile_X3Y11_LUT4AB/S2MID[7] Tile_X3Y11_LUT4AB/S2END[0] Tile_X3Y11_LUT4AB/S2END[1]
+ Tile_X3Y11_LUT4AB/S2END[2] Tile_X3Y11_LUT4AB/S2END[3] Tile_X3Y11_LUT4AB/S2END[4]
+ Tile_X3Y11_LUT4AB/S2END[5] Tile_X3Y11_LUT4AB/S2END[6] Tile_X3Y11_LUT4AB/S2END[7]
+ Tile_X3Y9_LUT4AB/S2BEGb[0] Tile_X3Y9_LUT4AB/S2BEGb[1] Tile_X3Y9_LUT4AB/S2BEGb[2]
+ Tile_X3Y9_LUT4AB/S2BEGb[3] Tile_X3Y9_LUT4AB/S2BEGb[4] Tile_X3Y9_LUT4AB/S2BEGb[5]
+ Tile_X3Y9_LUT4AB/S2BEGb[6] Tile_X3Y9_LUT4AB/S2BEGb[7] Tile_X3Y9_LUT4AB/S2BEG[0]
+ Tile_X3Y9_LUT4AB/S2BEG[1] Tile_X3Y9_LUT4AB/S2BEG[2] Tile_X3Y9_LUT4AB/S2BEG[3] Tile_X3Y9_LUT4AB/S2BEG[4]
+ Tile_X3Y9_LUT4AB/S2BEG[5] Tile_X3Y9_LUT4AB/S2BEG[6] Tile_X3Y9_LUT4AB/S2BEG[7] Tile_X3Y11_LUT4AB/S4END[0]
+ Tile_X3Y11_LUT4AB/S4END[10] Tile_X3Y11_LUT4AB/S4END[11] Tile_X3Y11_LUT4AB/S4END[12]
+ Tile_X3Y11_LUT4AB/S4END[13] Tile_X3Y11_LUT4AB/S4END[14] Tile_X3Y11_LUT4AB/S4END[15]
+ Tile_X3Y11_LUT4AB/S4END[1] Tile_X3Y11_LUT4AB/S4END[2] Tile_X3Y11_LUT4AB/S4END[3]
+ Tile_X3Y11_LUT4AB/S4END[4] Tile_X3Y11_LUT4AB/S4END[5] Tile_X3Y11_LUT4AB/S4END[6]
+ Tile_X3Y11_LUT4AB/S4END[7] Tile_X3Y11_LUT4AB/S4END[8] Tile_X3Y11_LUT4AB/S4END[9]
+ Tile_X3Y9_LUT4AB/S4BEG[0] Tile_X3Y9_LUT4AB/S4BEG[10] Tile_X3Y9_LUT4AB/S4BEG[11]
+ Tile_X3Y9_LUT4AB/S4BEG[12] Tile_X3Y9_LUT4AB/S4BEG[13] Tile_X3Y9_LUT4AB/S4BEG[14]
+ Tile_X3Y9_LUT4AB/S4BEG[15] Tile_X3Y9_LUT4AB/S4BEG[1] Tile_X3Y9_LUT4AB/S4BEG[2] Tile_X3Y9_LUT4AB/S4BEG[3]
+ Tile_X3Y9_LUT4AB/S4BEG[4] Tile_X3Y9_LUT4AB/S4BEG[5] Tile_X3Y9_LUT4AB/S4BEG[6] Tile_X3Y9_LUT4AB/S4BEG[7]
+ Tile_X3Y9_LUT4AB/S4BEG[8] Tile_X3Y9_LUT4AB/S4BEG[9] Tile_X3Y11_LUT4AB/SS4END[0]
+ Tile_X3Y11_LUT4AB/SS4END[10] Tile_X3Y11_LUT4AB/SS4END[11] Tile_X3Y11_LUT4AB/SS4END[12]
+ Tile_X3Y11_LUT4AB/SS4END[13] Tile_X3Y11_LUT4AB/SS4END[14] Tile_X3Y11_LUT4AB/SS4END[15]
+ Tile_X3Y11_LUT4AB/SS4END[1] Tile_X3Y11_LUT4AB/SS4END[2] Tile_X3Y11_LUT4AB/SS4END[3]
+ Tile_X3Y11_LUT4AB/SS4END[4] Tile_X3Y11_LUT4AB/SS4END[5] Tile_X3Y11_LUT4AB/SS4END[6]
+ Tile_X3Y11_LUT4AB/SS4END[7] Tile_X3Y11_LUT4AB/SS4END[8] Tile_X3Y11_LUT4AB/SS4END[9]
+ Tile_X3Y9_LUT4AB/SS4BEG[0] Tile_X3Y9_LUT4AB/SS4BEG[10] Tile_X3Y9_LUT4AB/SS4BEG[11]
+ Tile_X3Y9_LUT4AB/SS4BEG[12] Tile_X3Y9_LUT4AB/SS4BEG[13] Tile_X3Y9_LUT4AB/SS4BEG[14]
+ Tile_X3Y9_LUT4AB/SS4BEG[15] Tile_X3Y9_LUT4AB/SS4BEG[1] Tile_X3Y9_LUT4AB/SS4BEG[2]
+ Tile_X3Y9_LUT4AB/SS4BEG[3] Tile_X3Y9_LUT4AB/SS4BEG[4] Tile_X3Y9_LUT4AB/SS4BEG[5]
+ Tile_X3Y9_LUT4AB/SS4BEG[6] Tile_X3Y9_LUT4AB/SS4BEG[7] Tile_X3Y9_LUT4AB/SS4BEG[8]
+ Tile_X3Y9_LUT4AB/SS4BEG[9] Tile_X3Y10_LUT4AB/UserCLK Tile_X3Y9_LUT4AB/UserCLK VGND
+ VPWR Tile_X3Y10_LUT4AB/W1BEG[0] Tile_X3Y10_LUT4AB/W1BEG[1] Tile_X3Y10_LUT4AB/W1BEG[2]
+ Tile_X3Y10_LUT4AB/W1BEG[3] Tile_X3Y10_LUT4AB/W1END[0] Tile_X3Y10_LUT4AB/W1END[1]
+ Tile_X3Y10_LUT4AB/W1END[2] Tile_X3Y10_LUT4AB/W1END[3] Tile_X3Y10_LUT4AB/W2BEG[0]
+ Tile_X3Y10_LUT4AB/W2BEG[1] Tile_X3Y10_LUT4AB/W2BEG[2] Tile_X3Y10_LUT4AB/W2BEG[3]
+ Tile_X3Y10_LUT4AB/W2BEG[4] Tile_X3Y10_LUT4AB/W2BEG[5] Tile_X3Y10_LUT4AB/W2BEG[6]
+ Tile_X3Y10_LUT4AB/W2BEG[7] Tile_X2Y10_LUT4AB/W2END[0] Tile_X2Y10_LUT4AB/W2END[1]
+ Tile_X2Y10_LUT4AB/W2END[2] Tile_X2Y10_LUT4AB/W2END[3] Tile_X2Y10_LUT4AB/W2END[4]
+ Tile_X2Y10_LUT4AB/W2END[5] Tile_X2Y10_LUT4AB/W2END[6] Tile_X2Y10_LUT4AB/W2END[7]
+ Tile_X3Y10_LUT4AB/W2END[0] Tile_X3Y10_LUT4AB/W2END[1] Tile_X3Y10_LUT4AB/W2END[2]
+ Tile_X3Y10_LUT4AB/W2END[3] Tile_X3Y10_LUT4AB/W2END[4] Tile_X3Y10_LUT4AB/W2END[5]
+ Tile_X3Y10_LUT4AB/W2END[6] Tile_X3Y10_LUT4AB/W2END[7] Tile_X3Y10_LUT4AB/W2MID[0]
+ Tile_X3Y10_LUT4AB/W2MID[1] Tile_X3Y10_LUT4AB/W2MID[2] Tile_X3Y10_LUT4AB/W2MID[3]
+ Tile_X3Y10_LUT4AB/W2MID[4] Tile_X3Y10_LUT4AB/W2MID[5] Tile_X3Y10_LUT4AB/W2MID[6]
+ Tile_X3Y10_LUT4AB/W2MID[7] Tile_X3Y10_LUT4AB/W6BEG[0] Tile_X3Y10_LUT4AB/W6BEG[10]
+ Tile_X3Y10_LUT4AB/W6BEG[11] Tile_X3Y10_LUT4AB/W6BEG[1] Tile_X3Y10_LUT4AB/W6BEG[2]
+ Tile_X3Y10_LUT4AB/W6BEG[3] Tile_X3Y10_LUT4AB/W6BEG[4] Tile_X3Y10_LUT4AB/W6BEG[5]
+ Tile_X3Y10_LUT4AB/W6BEG[6] Tile_X3Y10_LUT4AB/W6BEG[7] Tile_X3Y10_LUT4AB/W6BEG[8]
+ Tile_X3Y10_LUT4AB/W6BEG[9] Tile_X3Y10_LUT4AB/W6END[0] Tile_X3Y10_LUT4AB/W6END[10]
+ Tile_X3Y10_LUT4AB/W6END[11] Tile_X3Y10_LUT4AB/W6END[1] Tile_X3Y10_LUT4AB/W6END[2]
+ Tile_X3Y10_LUT4AB/W6END[3] Tile_X3Y10_LUT4AB/W6END[4] Tile_X3Y10_LUT4AB/W6END[5]
+ Tile_X3Y10_LUT4AB/W6END[6] Tile_X3Y10_LUT4AB/W6END[7] Tile_X3Y10_LUT4AB/W6END[8]
+ Tile_X3Y10_LUT4AB/W6END[9] Tile_X3Y10_LUT4AB/WW4BEG[0] Tile_X3Y10_LUT4AB/WW4BEG[10]
+ Tile_X3Y10_LUT4AB/WW4BEG[11] Tile_X3Y10_LUT4AB/WW4BEG[12] Tile_X3Y10_LUT4AB/WW4BEG[13]
+ Tile_X3Y10_LUT4AB/WW4BEG[14] Tile_X3Y10_LUT4AB/WW4BEG[15] Tile_X3Y10_LUT4AB/WW4BEG[1]
+ Tile_X3Y10_LUT4AB/WW4BEG[2] Tile_X3Y10_LUT4AB/WW4BEG[3] Tile_X3Y10_LUT4AB/WW4BEG[4]
+ Tile_X3Y10_LUT4AB/WW4BEG[5] Tile_X3Y10_LUT4AB/WW4BEG[6] Tile_X3Y10_LUT4AB/WW4BEG[7]
+ Tile_X3Y10_LUT4AB/WW4BEG[8] Tile_X3Y10_LUT4AB/WW4BEG[9] Tile_X3Y10_LUT4AB/WW4END[0]
+ Tile_X3Y10_LUT4AB/WW4END[10] Tile_X3Y10_LUT4AB/WW4END[11] Tile_X3Y10_LUT4AB/WW4END[12]
+ Tile_X3Y10_LUT4AB/WW4END[13] Tile_X3Y10_LUT4AB/WW4END[14] Tile_X3Y10_LUT4AB/WW4END[15]
+ Tile_X3Y10_LUT4AB/WW4END[1] Tile_X3Y10_LUT4AB/WW4END[2] Tile_X3Y10_LUT4AB/WW4END[3]
+ Tile_X3Y10_LUT4AB/WW4END[4] Tile_X3Y10_LUT4AB/WW4END[5] Tile_X3Y10_LUT4AB/WW4END[6]
+ Tile_X3Y10_LUT4AB/WW4END[7] Tile_X3Y10_LUT4AB/WW4END[8] Tile_X3Y10_LUT4AB/WW4END[9]
+ LUT4AB
XTile_X7Y5_DSP Tile_X8Y5_LUT4AB/E1END[0] Tile_X8Y5_LUT4AB/E1END[1] Tile_X8Y5_LUT4AB/E1END[2]
+ Tile_X8Y5_LUT4AB/E1END[3] Tile_X6Y5_LUT4AB/E1BEG[0] Tile_X6Y5_LUT4AB/E1BEG[1] Tile_X6Y5_LUT4AB/E1BEG[2]
+ Tile_X6Y5_LUT4AB/E1BEG[3] Tile_X8Y5_LUT4AB/E2MID[0] Tile_X8Y5_LUT4AB/E2MID[1] Tile_X8Y5_LUT4AB/E2MID[2]
+ Tile_X8Y5_LUT4AB/E2MID[3] Tile_X8Y5_LUT4AB/E2MID[4] Tile_X8Y5_LUT4AB/E2MID[5] Tile_X8Y5_LUT4AB/E2MID[6]
+ Tile_X8Y5_LUT4AB/E2MID[7] Tile_X8Y5_LUT4AB/E2END[0] Tile_X8Y5_LUT4AB/E2END[1] Tile_X8Y5_LUT4AB/E2END[2]
+ Tile_X8Y5_LUT4AB/E2END[3] Tile_X8Y5_LUT4AB/E2END[4] Tile_X8Y5_LUT4AB/E2END[5] Tile_X8Y5_LUT4AB/E2END[6]
+ Tile_X8Y5_LUT4AB/E2END[7] Tile_X6Y5_LUT4AB/E2BEGb[0] Tile_X6Y5_LUT4AB/E2BEGb[1]
+ Tile_X6Y5_LUT4AB/E2BEGb[2] Tile_X6Y5_LUT4AB/E2BEGb[3] Tile_X6Y5_LUT4AB/E2BEGb[4]
+ Tile_X6Y5_LUT4AB/E2BEGb[5] Tile_X6Y5_LUT4AB/E2BEGb[6] Tile_X6Y5_LUT4AB/E2BEGb[7]
+ Tile_X6Y5_LUT4AB/E2BEG[0] Tile_X6Y5_LUT4AB/E2BEG[1] Tile_X6Y5_LUT4AB/E2BEG[2] Tile_X6Y5_LUT4AB/E2BEG[3]
+ Tile_X6Y5_LUT4AB/E2BEG[4] Tile_X6Y5_LUT4AB/E2BEG[5] Tile_X6Y5_LUT4AB/E2BEG[6] Tile_X6Y5_LUT4AB/E2BEG[7]
+ Tile_X8Y5_LUT4AB/E6END[0] Tile_X8Y5_LUT4AB/E6END[10] Tile_X8Y5_LUT4AB/E6END[11]
+ Tile_X8Y5_LUT4AB/E6END[1] Tile_X8Y5_LUT4AB/E6END[2] Tile_X8Y5_LUT4AB/E6END[3] Tile_X8Y5_LUT4AB/E6END[4]
+ Tile_X8Y5_LUT4AB/E6END[5] Tile_X8Y5_LUT4AB/E6END[6] Tile_X8Y5_LUT4AB/E6END[7] Tile_X8Y5_LUT4AB/E6END[8]
+ Tile_X8Y5_LUT4AB/E6END[9] Tile_X6Y5_LUT4AB/E6BEG[0] Tile_X6Y5_LUT4AB/E6BEG[10] Tile_X6Y5_LUT4AB/E6BEG[11]
+ Tile_X6Y5_LUT4AB/E6BEG[1] Tile_X6Y5_LUT4AB/E6BEG[2] Tile_X6Y5_LUT4AB/E6BEG[3] Tile_X6Y5_LUT4AB/E6BEG[4]
+ Tile_X6Y5_LUT4AB/E6BEG[5] Tile_X6Y5_LUT4AB/E6BEG[6] Tile_X6Y5_LUT4AB/E6BEG[7] Tile_X6Y5_LUT4AB/E6BEG[8]
+ Tile_X6Y5_LUT4AB/E6BEG[9] Tile_X8Y5_LUT4AB/EE4END[0] Tile_X8Y5_LUT4AB/EE4END[10]
+ Tile_X8Y5_LUT4AB/EE4END[11] Tile_X8Y5_LUT4AB/EE4END[12] Tile_X8Y5_LUT4AB/EE4END[13]
+ Tile_X8Y5_LUT4AB/EE4END[14] Tile_X8Y5_LUT4AB/EE4END[15] Tile_X8Y5_LUT4AB/EE4END[1]
+ Tile_X8Y5_LUT4AB/EE4END[2] Tile_X8Y5_LUT4AB/EE4END[3] Tile_X8Y5_LUT4AB/EE4END[4]
+ Tile_X8Y5_LUT4AB/EE4END[5] Tile_X8Y5_LUT4AB/EE4END[6] Tile_X8Y5_LUT4AB/EE4END[7]
+ Tile_X8Y5_LUT4AB/EE4END[8] Tile_X8Y5_LUT4AB/EE4END[9] Tile_X6Y5_LUT4AB/EE4BEG[0]
+ Tile_X6Y5_LUT4AB/EE4BEG[10] Tile_X6Y5_LUT4AB/EE4BEG[11] Tile_X6Y5_LUT4AB/EE4BEG[12]
+ Tile_X6Y5_LUT4AB/EE4BEG[13] Tile_X6Y5_LUT4AB/EE4BEG[14] Tile_X6Y5_LUT4AB/EE4BEG[15]
+ Tile_X6Y5_LUT4AB/EE4BEG[1] Tile_X6Y5_LUT4AB/EE4BEG[2] Tile_X6Y5_LUT4AB/EE4BEG[3]
+ Tile_X6Y5_LUT4AB/EE4BEG[4] Tile_X6Y5_LUT4AB/EE4BEG[5] Tile_X6Y5_LUT4AB/EE4BEG[6]
+ Tile_X6Y5_LUT4AB/EE4BEG[7] Tile_X6Y5_LUT4AB/EE4BEG[8] Tile_X6Y5_LUT4AB/EE4BEG[9]
+ Tile_X6Y5_LUT4AB/FrameData_O[0] Tile_X6Y5_LUT4AB/FrameData_O[10] Tile_X6Y5_LUT4AB/FrameData_O[11]
+ Tile_X6Y5_LUT4AB/FrameData_O[12] Tile_X6Y5_LUT4AB/FrameData_O[13] Tile_X6Y5_LUT4AB/FrameData_O[14]
+ Tile_X6Y5_LUT4AB/FrameData_O[15] Tile_X6Y5_LUT4AB/FrameData_O[16] Tile_X6Y5_LUT4AB/FrameData_O[17]
+ Tile_X6Y5_LUT4AB/FrameData_O[18] Tile_X6Y5_LUT4AB/FrameData_O[19] Tile_X6Y5_LUT4AB/FrameData_O[1]
+ Tile_X6Y5_LUT4AB/FrameData_O[20] Tile_X6Y5_LUT4AB/FrameData_O[21] Tile_X6Y5_LUT4AB/FrameData_O[22]
+ Tile_X6Y5_LUT4AB/FrameData_O[23] Tile_X6Y5_LUT4AB/FrameData_O[24] Tile_X6Y5_LUT4AB/FrameData_O[25]
+ Tile_X6Y5_LUT4AB/FrameData_O[26] Tile_X6Y5_LUT4AB/FrameData_O[27] Tile_X6Y5_LUT4AB/FrameData_O[28]
+ Tile_X6Y5_LUT4AB/FrameData_O[29] Tile_X6Y5_LUT4AB/FrameData_O[2] Tile_X6Y5_LUT4AB/FrameData_O[30]
+ Tile_X6Y5_LUT4AB/FrameData_O[31] Tile_X6Y5_LUT4AB/FrameData_O[3] Tile_X6Y5_LUT4AB/FrameData_O[4]
+ Tile_X6Y5_LUT4AB/FrameData_O[5] Tile_X6Y5_LUT4AB/FrameData_O[6] Tile_X6Y5_LUT4AB/FrameData_O[7]
+ Tile_X6Y5_LUT4AB/FrameData_O[8] Tile_X6Y5_LUT4AB/FrameData_O[9] Tile_X8Y5_LUT4AB/FrameData[0]
+ Tile_X8Y5_LUT4AB/FrameData[10] Tile_X8Y5_LUT4AB/FrameData[11] Tile_X8Y5_LUT4AB/FrameData[12]
+ Tile_X8Y5_LUT4AB/FrameData[13] Tile_X8Y5_LUT4AB/FrameData[14] Tile_X8Y5_LUT4AB/FrameData[15]
+ Tile_X8Y5_LUT4AB/FrameData[16] Tile_X8Y5_LUT4AB/FrameData[17] Tile_X8Y5_LUT4AB/FrameData[18]
+ Tile_X8Y5_LUT4AB/FrameData[19] Tile_X8Y5_LUT4AB/FrameData[1] Tile_X8Y5_LUT4AB/FrameData[20]
+ Tile_X8Y5_LUT4AB/FrameData[21] Tile_X8Y5_LUT4AB/FrameData[22] Tile_X8Y5_LUT4AB/FrameData[23]
+ Tile_X8Y5_LUT4AB/FrameData[24] Tile_X8Y5_LUT4AB/FrameData[25] Tile_X8Y5_LUT4AB/FrameData[26]
+ Tile_X8Y5_LUT4AB/FrameData[27] Tile_X8Y5_LUT4AB/FrameData[28] Tile_X8Y5_LUT4AB/FrameData[29]
+ Tile_X8Y5_LUT4AB/FrameData[2] Tile_X8Y5_LUT4AB/FrameData[30] Tile_X8Y5_LUT4AB/FrameData[31]
+ Tile_X8Y5_LUT4AB/FrameData[3] Tile_X8Y5_LUT4AB/FrameData[4] Tile_X8Y5_LUT4AB/FrameData[5]
+ Tile_X8Y5_LUT4AB/FrameData[6] Tile_X8Y5_LUT4AB/FrameData[7] Tile_X8Y5_LUT4AB/FrameData[8]
+ Tile_X8Y5_LUT4AB/FrameData[9] Tile_X7Y3_DSP/Tile_X0Y1_FrameStrobe[0] Tile_X7Y3_DSP/Tile_X0Y1_FrameStrobe[10]
+ Tile_X7Y3_DSP/Tile_X0Y1_FrameStrobe[11] Tile_X7Y3_DSP/Tile_X0Y1_FrameStrobe[12]
+ Tile_X7Y3_DSP/Tile_X0Y1_FrameStrobe[13] Tile_X7Y3_DSP/Tile_X0Y1_FrameStrobe[14]
+ Tile_X7Y3_DSP/Tile_X0Y1_FrameStrobe[15] Tile_X7Y3_DSP/Tile_X0Y1_FrameStrobe[16]
+ Tile_X7Y3_DSP/Tile_X0Y1_FrameStrobe[17] Tile_X7Y3_DSP/Tile_X0Y1_FrameStrobe[18]
+ Tile_X7Y3_DSP/Tile_X0Y1_FrameStrobe[19] Tile_X7Y3_DSP/Tile_X0Y1_FrameStrobe[1] Tile_X7Y3_DSP/Tile_X0Y1_FrameStrobe[2]
+ Tile_X7Y3_DSP/Tile_X0Y1_FrameStrobe[3] Tile_X7Y3_DSP/Tile_X0Y1_FrameStrobe[4] Tile_X7Y3_DSP/Tile_X0Y1_FrameStrobe[5]
+ Tile_X7Y3_DSP/Tile_X0Y1_FrameStrobe[6] Tile_X7Y3_DSP/Tile_X0Y1_FrameStrobe[7] Tile_X7Y3_DSP/Tile_X0Y1_FrameStrobe[8]
+ Tile_X7Y3_DSP/Tile_X0Y1_FrameStrobe[9] Tile_X7Y5_DSP/Tile_X0Y0_N1BEG[0] Tile_X7Y5_DSP/Tile_X0Y0_N1BEG[1]
+ Tile_X7Y5_DSP/Tile_X0Y0_N1BEG[2] Tile_X7Y5_DSP/Tile_X0Y0_N1BEG[3] Tile_X7Y5_DSP/Tile_X0Y0_N2BEG[0]
+ Tile_X7Y5_DSP/Tile_X0Y0_N2BEG[1] Tile_X7Y5_DSP/Tile_X0Y0_N2BEG[2] Tile_X7Y5_DSP/Tile_X0Y0_N2BEG[3]
+ Tile_X7Y5_DSP/Tile_X0Y0_N2BEG[4] Tile_X7Y5_DSP/Tile_X0Y0_N2BEG[5] Tile_X7Y5_DSP/Tile_X0Y0_N2BEG[6]
+ Tile_X7Y5_DSP/Tile_X0Y0_N2BEG[7] Tile_X7Y3_DSP/Tile_X0Y1_N2END[0] Tile_X7Y3_DSP/Tile_X0Y1_N2END[1]
+ Tile_X7Y3_DSP/Tile_X0Y1_N2END[2] Tile_X7Y3_DSP/Tile_X0Y1_N2END[3] Tile_X7Y3_DSP/Tile_X0Y1_N2END[4]
+ Tile_X7Y3_DSP/Tile_X0Y1_N2END[5] Tile_X7Y3_DSP/Tile_X0Y1_N2END[6] Tile_X7Y3_DSP/Tile_X0Y1_N2END[7]
+ Tile_X7Y5_DSP/Tile_X0Y0_N4BEG[0] Tile_X7Y5_DSP/Tile_X0Y0_N4BEG[10] Tile_X7Y5_DSP/Tile_X0Y0_N4BEG[11]
+ Tile_X7Y5_DSP/Tile_X0Y0_N4BEG[12] Tile_X7Y5_DSP/Tile_X0Y0_N4BEG[13] Tile_X7Y5_DSP/Tile_X0Y0_N4BEG[14]
+ Tile_X7Y5_DSP/Tile_X0Y0_N4BEG[15] Tile_X7Y5_DSP/Tile_X0Y0_N4BEG[1] Tile_X7Y5_DSP/Tile_X0Y0_N4BEG[2]
+ Tile_X7Y5_DSP/Tile_X0Y0_N4BEG[3] Tile_X7Y5_DSP/Tile_X0Y0_N4BEG[4] Tile_X7Y5_DSP/Tile_X0Y0_N4BEG[5]
+ Tile_X7Y5_DSP/Tile_X0Y0_N4BEG[6] Tile_X7Y5_DSP/Tile_X0Y0_N4BEG[7] Tile_X7Y5_DSP/Tile_X0Y0_N4BEG[8]
+ Tile_X7Y5_DSP/Tile_X0Y0_N4BEG[9] Tile_X7Y5_DSP/Tile_X0Y0_NN4BEG[0] Tile_X7Y5_DSP/Tile_X0Y0_NN4BEG[10]
+ Tile_X7Y5_DSP/Tile_X0Y0_NN4BEG[11] Tile_X7Y5_DSP/Tile_X0Y0_NN4BEG[12] Tile_X7Y5_DSP/Tile_X0Y0_NN4BEG[13]
+ Tile_X7Y5_DSP/Tile_X0Y0_NN4BEG[14] Tile_X7Y5_DSP/Tile_X0Y0_NN4BEG[15] Tile_X7Y5_DSP/Tile_X0Y0_NN4BEG[1]
+ Tile_X7Y5_DSP/Tile_X0Y0_NN4BEG[2] Tile_X7Y5_DSP/Tile_X0Y0_NN4BEG[3] Tile_X7Y5_DSP/Tile_X0Y0_NN4BEG[4]
+ Tile_X7Y5_DSP/Tile_X0Y0_NN4BEG[5] Tile_X7Y5_DSP/Tile_X0Y0_NN4BEG[6] Tile_X7Y5_DSP/Tile_X0Y0_NN4BEG[7]
+ Tile_X7Y5_DSP/Tile_X0Y0_NN4BEG[8] Tile_X7Y5_DSP/Tile_X0Y0_NN4BEG[9] Tile_X7Y5_DSP/Tile_X0Y0_S1END[0]
+ Tile_X7Y5_DSP/Tile_X0Y0_S1END[1] Tile_X7Y5_DSP/Tile_X0Y0_S1END[2] Tile_X7Y5_DSP/Tile_X0Y0_S1END[3]
+ Tile_X7Y5_DSP/Tile_X0Y0_S2END[0] Tile_X7Y5_DSP/Tile_X0Y0_S2END[1] Tile_X7Y5_DSP/Tile_X0Y0_S2END[2]
+ Tile_X7Y5_DSP/Tile_X0Y0_S2END[3] Tile_X7Y5_DSP/Tile_X0Y0_S2END[4] Tile_X7Y5_DSP/Tile_X0Y0_S2END[5]
+ Tile_X7Y5_DSP/Tile_X0Y0_S2END[6] Tile_X7Y5_DSP/Tile_X0Y0_S2END[7] Tile_X7Y5_DSP/Tile_X0Y0_S2MID[0]
+ Tile_X7Y5_DSP/Tile_X0Y0_S2MID[1] Tile_X7Y5_DSP/Tile_X0Y0_S2MID[2] Tile_X7Y5_DSP/Tile_X0Y0_S2MID[3]
+ Tile_X7Y5_DSP/Tile_X0Y0_S2MID[4] Tile_X7Y5_DSP/Tile_X0Y0_S2MID[5] Tile_X7Y5_DSP/Tile_X0Y0_S2MID[6]
+ Tile_X7Y5_DSP/Tile_X0Y0_S2MID[7] Tile_X7Y5_DSP/Tile_X0Y0_S4END[0] Tile_X7Y5_DSP/Tile_X0Y0_S4END[10]
+ Tile_X7Y5_DSP/Tile_X0Y0_S4END[11] Tile_X7Y5_DSP/Tile_X0Y0_S4END[12] Tile_X7Y5_DSP/Tile_X0Y0_S4END[13]
+ Tile_X7Y5_DSP/Tile_X0Y0_S4END[14] Tile_X7Y5_DSP/Tile_X0Y0_S4END[15] Tile_X7Y5_DSP/Tile_X0Y0_S4END[1]
+ Tile_X7Y5_DSP/Tile_X0Y0_S4END[2] Tile_X7Y5_DSP/Tile_X0Y0_S4END[3] Tile_X7Y5_DSP/Tile_X0Y0_S4END[4]
+ Tile_X7Y5_DSP/Tile_X0Y0_S4END[5] Tile_X7Y5_DSP/Tile_X0Y0_S4END[6] Tile_X7Y5_DSP/Tile_X0Y0_S4END[7]
+ Tile_X7Y5_DSP/Tile_X0Y0_S4END[8] Tile_X7Y5_DSP/Tile_X0Y0_S4END[9] Tile_X7Y5_DSP/Tile_X0Y0_SS4END[0]
+ Tile_X7Y5_DSP/Tile_X0Y0_SS4END[10] Tile_X7Y5_DSP/Tile_X0Y0_SS4END[11] Tile_X7Y5_DSP/Tile_X0Y0_SS4END[12]
+ Tile_X7Y5_DSP/Tile_X0Y0_SS4END[13] Tile_X7Y5_DSP/Tile_X0Y0_SS4END[14] Tile_X7Y5_DSP/Tile_X0Y0_SS4END[15]
+ Tile_X7Y5_DSP/Tile_X0Y0_SS4END[1] Tile_X7Y5_DSP/Tile_X0Y0_SS4END[2] Tile_X7Y5_DSP/Tile_X0Y0_SS4END[3]
+ Tile_X7Y5_DSP/Tile_X0Y0_SS4END[4] Tile_X7Y5_DSP/Tile_X0Y0_SS4END[5] Tile_X7Y5_DSP/Tile_X0Y0_SS4END[6]
+ Tile_X7Y5_DSP/Tile_X0Y0_SS4END[7] Tile_X7Y5_DSP/Tile_X0Y0_SS4END[8] Tile_X7Y5_DSP/Tile_X0Y0_SS4END[9]
+ Tile_X7Y3_DSP/Tile_X0Y1_UserCLK Tile_X6Y5_LUT4AB/W1END[0] Tile_X6Y5_LUT4AB/W1END[1]
+ Tile_X6Y5_LUT4AB/W1END[2] Tile_X6Y5_LUT4AB/W1END[3] Tile_X8Y5_LUT4AB/W1BEG[0] Tile_X8Y5_LUT4AB/W1BEG[1]
+ Tile_X8Y5_LUT4AB/W1BEG[2] Tile_X8Y5_LUT4AB/W1BEG[3] Tile_X6Y5_LUT4AB/W2MID[0] Tile_X6Y5_LUT4AB/W2MID[1]
+ Tile_X6Y5_LUT4AB/W2MID[2] Tile_X6Y5_LUT4AB/W2MID[3] Tile_X6Y5_LUT4AB/W2MID[4] Tile_X6Y5_LUT4AB/W2MID[5]
+ Tile_X6Y5_LUT4AB/W2MID[6] Tile_X6Y5_LUT4AB/W2MID[7] Tile_X6Y5_LUT4AB/W2END[0] Tile_X6Y5_LUT4AB/W2END[1]
+ Tile_X6Y5_LUT4AB/W2END[2] Tile_X6Y5_LUT4AB/W2END[3] Tile_X6Y5_LUT4AB/W2END[4] Tile_X6Y5_LUT4AB/W2END[5]
+ Tile_X6Y5_LUT4AB/W2END[6] Tile_X6Y5_LUT4AB/W2END[7] Tile_X8Y5_LUT4AB/W2BEGb[0] Tile_X8Y5_LUT4AB/W2BEGb[1]
+ Tile_X8Y5_LUT4AB/W2BEGb[2] Tile_X8Y5_LUT4AB/W2BEGb[3] Tile_X8Y5_LUT4AB/W2BEGb[4]
+ Tile_X8Y5_LUT4AB/W2BEGb[5] Tile_X8Y5_LUT4AB/W2BEGb[6] Tile_X8Y5_LUT4AB/W2BEGb[7]
+ Tile_X8Y5_LUT4AB/W2BEG[0] Tile_X8Y5_LUT4AB/W2BEG[1] Tile_X8Y5_LUT4AB/W2BEG[2] Tile_X8Y5_LUT4AB/W2BEG[3]
+ Tile_X8Y5_LUT4AB/W2BEG[4] Tile_X8Y5_LUT4AB/W2BEG[5] Tile_X8Y5_LUT4AB/W2BEG[6] Tile_X8Y5_LUT4AB/W2BEG[7]
+ Tile_X6Y5_LUT4AB/W6END[0] Tile_X6Y5_LUT4AB/W6END[10] Tile_X6Y5_LUT4AB/W6END[11]
+ Tile_X6Y5_LUT4AB/W6END[1] Tile_X6Y5_LUT4AB/W6END[2] Tile_X6Y5_LUT4AB/W6END[3] Tile_X6Y5_LUT4AB/W6END[4]
+ Tile_X6Y5_LUT4AB/W6END[5] Tile_X6Y5_LUT4AB/W6END[6] Tile_X6Y5_LUT4AB/W6END[7] Tile_X6Y5_LUT4AB/W6END[8]
+ Tile_X6Y5_LUT4AB/W6END[9] Tile_X8Y5_LUT4AB/W6BEG[0] Tile_X8Y5_LUT4AB/W6BEG[10] Tile_X8Y5_LUT4AB/W6BEG[11]
+ Tile_X8Y5_LUT4AB/W6BEG[1] Tile_X8Y5_LUT4AB/W6BEG[2] Tile_X8Y5_LUT4AB/W6BEG[3] Tile_X8Y5_LUT4AB/W6BEG[4]
+ Tile_X8Y5_LUT4AB/W6BEG[5] Tile_X8Y5_LUT4AB/W6BEG[6] Tile_X8Y5_LUT4AB/W6BEG[7] Tile_X8Y5_LUT4AB/W6BEG[8]
+ Tile_X8Y5_LUT4AB/W6BEG[9] Tile_X6Y5_LUT4AB/WW4END[0] Tile_X6Y5_LUT4AB/WW4END[10]
+ Tile_X6Y5_LUT4AB/WW4END[11] Tile_X6Y5_LUT4AB/WW4END[12] Tile_X6Y5_LUT4AB/WW4END[13]
+ Tile_X6Y5_LUT4AB/WW4END[14] Tile_X6Y5_LUT4AB/WW4END[15] Tile_X6Y5_LUT4AB/WW4END[1]
+ Tile_X6Y5_LUT4AB/WW4END[2] Tile_X6Y5_LUT4AB/WW4END[3] Tile_X6Y5_LUT4AB/WW4END[4]
+ Tile_X6Y5_LUT4AB/WW4END[5] Tile_X6Y5_LUT4AB/WW4END[6] Tile_X6Y5_LUT4AB/WW4END[7]
+ Tile_X6Y5_LUT4AB/WW4END[8] Tile_X6Y5_LUT4AB/WW4END[9] Tile_X8Y5_LUT4AB/WW4BEG[0]
+ Tile_X8Y5_LUT4AB/WW4BEG[10] Tile_X8Y5_LUT4AB/WW4BEG[11] Tile_X8Y5_LUT4AB/WW4BEG[12]
+ Tile_X8Y5_LUT4AB/WW4BEG[13] Tile_X8Y5_LUT4AB/WW4BEG[14] Tile_X8Y5_LUT4AB/WW4BEG[15]
+ Tile_X8Y5_LUT4AB/WW4BEG[1] Tile_X8Y5_LUT4AB/WW4BEG[2] Tile_X8Y5_LUT4AB/WW4BEG[3]
+ Tile_X8Y5_LUT4AB/WW4BEG[4] Tile_X8Y5_LUT4AB/WW4BEG[5] Tile_X8Y5_LUT4AB/WW4BEG[6]
+ Tile_X8Y5_LUT4AB/WW4BEG[7] Tile_X8Y5_LUT4AB/WW4BEG[8] Tile_X8Y5_LUT4AB/WW4BEG[9]
+ Tile_X8Y6_LUT4AB/E1END[0] Tile_X8Y6_LUT4AB/E1END[1] Tile_X8Y6_LUT4AB/E1END[2] Tile_X8Y6_LUT4AB/E1END[3]
+ Tile_X6Y6_LUT4AB/E1BEG[0] Tile_X6Y6_LUT4AB/E1BEG[1] Tile_X6Y6_LUT4AB/E1BEG[2] Tile_X6Y6_LUT4AB/E1BEG[3]
+ Tile_X8Y6_LUT4AB/E2MID[0] Tile_X8Y6_LUT4AB/E2MID[1] Tile_X8Y6_LUT4AB/E2MID[2] Tile_X8Y6_LUT4AB/E2MID[3]
+ Tile_X8Y6_LUT4AB/E2MID[4] Tile_X8Y6_LUT4AB/E2MID[5] Tile_X8Y6_LUT4AB/E2MID[6] Tile_X8Y6_LUT4AB/E2MID[7]
+ Tile_X8Y6_LUT4AB/E2END[0] Tile_X8Y6_LUT4AB/E2END[1] Tile_X8Y6_LUT4AB/E2END[2] Tile_X8Y6_LUT4AB/E2END[3]
+ Tile_X8Y6_LUT4AB/E2END[4] Tile_X8Y6_LUT4AB/E2END[5] Tile_X8Y6_LUT4AB/E2END[6] Tile_X8Y6_LUT4AB/E2END[7]
+ Tile_X6Y6_LUT4AB/E2BEGb[0] Tile_X6Y6_LUT4AB/E2BEGb[1] Tile_X6Y6_LUT4AB/E2BEGb[2]
+ Tile_X6Y6_LUT4AB/E2BEGb[3] Tile_X6Y6_LUT4AB/E2BEGb[4] Tile_X6Y6_LUT4AB/E2BEGb[5]
+ Tile_X6Y6_LUT4AB/E2BEGb[6] Tile_X6Y6_LUT4AB/E2BEGb[7] Tile_X6Y6_LUT4AB/E2BEG[0]
+ Tile_X6Y6_LUT4AB/E2BEG[1] Tile_X6Y6_LUT4AB/E2BEG[2] Tile_X6Y6_LUT4AB/E2BEG[3] Tile_X6Y6_LUT4AB/E2BEG[4]
+ Tile_X6Y6_LUT4AB/E2BEG[5] Tile_X6Y6_LUT4AB/E2BEG[6] Tile_X6Y6_LUT4AB/E2BEG[7] Tile_X8Y6_LUT4AB/E6END[0]
+ Tile_X8Y6_LUT4AB/E6END[10] Tile_X8Y6_LUT4AB/E6END[11] Tile_X8Y6_LUT4AB/E6END[1]
+ Tile_X8Y6_LUT4AB/E6END[2] Tile_X8Y6_LUT4AB/E6END[3] Tile_X8Y6_LUT4AB/E6END[4] Tile_X8Y6_LUT4AB/E6END[5]
+ Tile_X8Y6_LUT4AB/E6END[6] Tile_X8Y6_LUT4AB/E6END[7] Tile_X8Y6_LUT4AB/E6END[8] Tile_X8Y6_LUT4AB/E6END[9]
+ Tile_X6Y6_LUT4AB/E6BEG[0] Tile_X6Y6_LUT4AB/E6BEG[10] Tile_X6Y6_LUT4AB/E6BEG[11]
+ Tile_X6Y6_LUT4AB/E6BEG[1] Tile_X6Y6_LUT4AB/E6BEG[2] Tile_X6Y6_LUT4AB/E6BEG[3] Tile_X6Y6_LUT4AB/E6BEG[4]
+ Tile_X6Y6_LUT4AB/E6BEG[5] Tile_X6Y6_LUT4AB/E6BEG[6] Tile_X6Y6_LUT4AB/E6BEG[7] Tile_X6Y6_LUT4AB/E6BEG[8]
+ Tile_X6Y6_LUT4AB/E6BEG[9] Tile_X8Y6_LUT4AB/EE4END[0] Tile_X8Y6_LUT4AB/EE4END[10]
+ Tile_X8Y6_LUT4AB/EE4END[11] Tile_X8Y6_LUT4AB/EE4END[12] Tile_X8Y6_LUT4AB/EE4END[13]
+ Tile_X8Y6_LUT4AB/EE4END[14] Tile_X8Y6_LUT4AB/EE4END[15] Tile_X8Y6_LUT4AB/EE4END[1]
+ Tile_X8Y6_LUT4AB/EE4END[2] Tile_X8Y6_LUT4AB/EE4END[3] Tile_X8Y6_LUT4AB/EE4END[4]
+ Tile_X8Y6_LUT4AB/EE4END[5] Tile_X8Y6_LUT4AB/EE4END[6] Tile_X8Y6_LUT4AB/EE4END[7]
+ Tile_X8Y6_LUT4AB/EE4END[8] Tile_X8Y6_LUT4AB/EE4END[9] Tile_X6Y6_LUT4AB/EE4BEG[0]
+ Tile_X6Y6_LUT4AB/EE4BEG[10] Tile_X6Y6_LUT4AB/EE4BEG[11] Tile_X6Y6_LUT4AB/EE4BEG[12]
+ Tile_X6Y6_LUT4AB/EE4BEG[13] Tile_X6Y6_LUT4AB/EE4BEG[14] Tile_X6Y6_LUT4AB/EE4BEG[15]
+ Tile_X6Y6_LUT4AB/EE4BEG[1] Tile_X6Y6_LUT4AB/EE4BEG[2] Tile_X6Y6_LUT4AB/EE4BEG[3]
+ Tile_X6Y6_LUT4AB/EE4BEG[4] Tile_X6Y6_LUT4AB/EE4BEG[5] Tile_X6Y6_LUT4AB/EE4BEG[6]
+ Tile_X6Y6_LUT4AB/EE4BEG[7] Tile_X6Y6_LUT4AB/EE4BEG[8] Tile_X6Y6_LUT4AB/EE4BEG[9]
+ Tile_X6Y6_LUT4AB/FrameData_O[0] Tile_X6Y6_LUT4AB/FrameData_O[10] Tile_X6Y6_LUT4AB/FrameData_O[11]
+ Tile_X6Y6_LUT4AB/FrameData_O[12] Tile_X6Y6_LUT4AB/FrameData_O[13] Tile_X6Y6_LUT4AB/FrameData_O[14]
+ Tile_X6Y6_LUT4AB/FrameData_O[15] Tile_X6Y6_LUT4AB/FrameData_O[16] Tile_X6Y6_LUT4AB/FrameData_O[17]
+ Tile_X6Y6_LUT4AB/FrameData_O[18] Tile_X6Y6_LUT4AB/FrameData_O[19] Tile_X6Y6_LUT4AB/FrameData_O[1]
+ Tile_X6Y6_LUT4AB/FrameData_O[20] Tile_X6Y6_LUT4AB/FrameData_O[21] Tile_X6Y6_LUT4AB/FrameData_O[22]
+ Tile_X6Y6_LUT4AB/FrameData_O[23] Tile_X6Y6_LUT4AB/FrameData_O[24] Tile_X6Y6_LUT4AB/FrameData_O[25]
+ Tile_X6Y6_LUT4AB/FrameData_O[26] Tile_X6Y6_LUT4AB/FrameData_O[27] Tile_X6Y6_LUT4AB/FrameData_O[28]
+ Tile_X6Y6_LUT4AB/FrameData_O[29] Tile_X6Y6_LUT4AB/FrameData_O[2] Tile_X6Y6_LUT4AB/FrameData_O[30]
+ Tile_X6Y6_LUT4AB/FrameData_O[31] Tile_X6Y6_LUT4AB/FrameData_O[3] Tile_X6Y6_LUT4AB/FrameData_O[4]
+ Tile_X6Y6_LUT4AB/FrameData_O[5] Tile_X6Y6_LUT4AB/FrameData_O[6] Tile_X6Y6_LUT4AB/FrameData_O[7]
+ Tile_X6Y6_LUT4AB/FrameData_O[8] Tile_X6Y6_LUT4AB/FrameData_O[9] Tile_X8Y6_LUT4AB/FrameData[0]
+ Tile_X8Y6_LUT4AB/FrameData[10] Tile_X8Y6_LUT4AB/FrameData[11] Tile_X8Y6_LUT4AB/FrameData[12]
+ Tile_X8Y6_LUT4AB/FrameData[13] Tile_X8Y6_LUT4AB/FrameData[14] Tile_X8Y6_LUT4AB/FrameData[15]
+ Tile_X8Y6_LUT4AB/FrameData[16] Tile_X8Y6_LUT4AB/FrameData[17] Tile_X8Y6_LUT4AB/FrameData[18]
+ Tile_X8Y6_LUT4AB/FrameData[19] Tile_X8Y6_LUT4AB/FrameData[1] Tile_X8Y6_LUT4AB/FrameData[20]
+ Tile_X8Y6_LUT4AB/FrameData[21] Tile_X8Y6_LUT4AB/FrameData[22] Tile_X8Y6_LUT4AB/FrameData[23]
+ Tile_X8Y6_LUT4AB/FrameData[24] Tile_X8Y6_LUT4AB/FrameData[25] Tile_X8Y6_LUT4AB/FrameData[26]
+ Tile_X8Y6_LUT4AB/FrameData[27] Tile_X8Y6_LUT4AB/FrameData[28] Tile_X8Y6_LUT4AB/FrameData[29]
+ Tile_X8Y6_LUT4AB/FrameData[2] Tile_X8Y6_LUT4AB/FrameData[30] Tile_X8Y6_LUT4AB/FrameData[31]
+ Tile_X8Y6_LUT4AB/FrameData[3] Tile_X8Y6_LUT4AB/FrameData[4] Tile_X8Y6_LUT4AB/FrameData[5]
+ Tile_X8Y6_LUT4AB/FrameData[6] Tile_X8Y6_LUT4AB/FrameData[7] Tile_X8Y6_LUT4AB/FrameData[8]
+ Tile_X8Y6_LUT4AB/FrameData[9] Tile_X7Y5_DSP/Tile_X0Y1_FrameStrobe[0] Tile_X7Y5_DSP/Tile_X0Y1_FrameStrobe[10]
+ Tile_X7Y5_DSP/Tile_X0Y1_FrameStrobe[11] Tile_X7Y5_DSP/Tile_X0Y1_FrameStrobe[12]
+ Tile_X7Y5_DSP/Tile_X0Y1_FrameStrobe[13] Tile_X7Y5_DSP/Tile_X0Y1_FrameStrobe[14]
+ Tile_X7Y5_DSP/Tile_X0Y1_FrameStrobe[15] Tile_X7Y5_DSP/Tile_X0Y1_FrameStrobe[16]
+ Tile_X7Y5_DSP/Tile_X0Y1_FrameStrobe[17] Tile_X7Y5_DSP/Tile_X0Y1_FrameStrobe[18]
+ Tile_X7Y5_DSP/Tile_X0Y1_FrameStrobe[19] Tile_X7Y5_DSP/Tile_X0Y1_FrameStrobe[1] Tile_X7Y5_DSP/Tile_X0Y1_FrameStrobe[2]
+ Tile_X7Y5_DSP/Tile_X0Y1_FrameStrobe[3] Tile_X7Y5_DSP/Tile_X0Y1_FrameStrobe[4] Tile_X7Y5_DSP/Tile_X0Y1_FrameStrobe[5]
+ Tile_X7Y5_DSP/Tile_X0Y1_FrameStrobe[6] Tile_X7Y5_DSP/Tile_X0Y1_FrameStrobe[7] Tile_X7Y5_DSP/Tile_X0Y1_FrameStrobe[8]
+ Tile_X7Y5_DSP/Tile_X0Y1_FrameStrobe[9] Tile_X7Y7_DSP/Tile_X0Y0_N1BEG[0] Tile_X7Y7_DSP/Tile_X0Y0_N1BEG[1]
+ Tile_X7Y7_DSP/Tile_X0Y0_N1BEG[2] Tile_X7Y7_DSP/Tile_X0Y0_N1BEG[3] Tile_X7Y5_DSP/Tile_X0Y1_N2END[0]
+ Tile_X7Y5_DSP/Tile_X0Y1_N2END[1] Tile_X7Y5_DSP/Tile_X0Y1_N2END[2] Tile_X7Y5_DSP/Tile_X0Y1_N2END[3]
+ Tile_X7Y5_DSP/Tile_X0Y1_N2END[4] Tile_X7Y5_DSP/Tile_X0Y1_N2END[5] Tile_X7Y5_DSP/Tile_X0Y1_N2END[6]
+ Tile_X7Y5_DSP/Tile_X0Y1_N2END[7] Tile_X7Y7_DSP/Tile_X0Y0_N2BEG[0] Tile_X7Y7_DSP/Tile_X0Y0_N2BEG[1]
+ Tile_X7Y7_DSP/Tile_X0Y0_N2BEG[2] Tile_X7Y7_DSP/Tile_X0Y0_N2BEG[3] Tile_X7Y7_DSP/Tile_X0Y0_N2BEG[4]
+ Tile_X7Y7_DSP/Tile_X0Y0_N2BEG[5] Tile_X7Y7_DSP/Tile_X0Y0_N2BEG[6] Tile_X7Y7_DSP/Tile_X0Y0_N2BEG[7]
+ Tile_X7Y7_DSP/Tile_X0Y0_N4BEG[0] Tile_X7Y7_DSP/Tile_X0Y0_N4BEG[10] Tile_X7Y7_DSP/Tile_X0Y0_N4BEG[11]
+ Tile_X7Y7_DSP/Tile_X0Y0_N4BEG[12] Tile_X7Y7_DSP/Tile_X0Y0_N4BEG[13] Tile_X7Y7_DSP/Tile_X0Y0_N4BEG[14]
+ Tile_X7Y7_DSP/Tile_X0Y0_N4BEG[15] Tile_X7Y7_DSP/Tile_X0Y0_N4BEG[1] Tile_X7Y7_DSP/Tile_X0Y0_N4BEG[2]
+ Tile_X7Y7_DSP/Tile_X0Y0_N4BEG[3] Tile_X7Y7_DSP/Tile_X0Y0_N4BEG[4] Tile_X7Y7_DSP/Tile_X0Y0_N4BEG[5]
+ Tile_X7Y7_DSP/Tile_X0Y0_N4BEG[6] Tile_X7Y7_DSP/Tile_X0Y0_N4BEG[7] Tile_X7Y7_DSP/Tile_X0Y0_N4BEG[8]
+ Tile_X7Y7_DSP/Tile_X0Y0_N4BEG[9] Tile_X7Y7_DSP/Tile_X0Y0_NN4BEG[0] Tile_X7Y7_DSP/Tile_X0Y0_NN4BEG[10]
+ Tile_X7Y7_DSP/Tile_X0Y0_NN4BEG[11] Tile_X7Y7_DSP/Tile_X0Y0_NN4BEG[12] Tile_X7Y7_DSP/Tile_X0Y0_NN4BEG[13]
+ Tile_X7Y7_DSP/Tile_X0Y0_NN4BEG[14] Tile_X7Y7_DSP/Tile_X0Y0_NN4BEG[15] Tile_X7Y7_DSP/Tile_X0Y0_NN4BEG[1]
+ Tile_X7Y7_DSP/Tile_X0Y0_NN4BEG[2] Tile_X7Y7_DSP/Tile_X0Y0_NN4BEG[3] Tile_X7Y7_DSP/Tile_X0Y0_NN4BEG[4]
+ Tile_X7Y7_DSP/Tile_X0Y0_NN4BEG[5] Tile_X7Y7_DSP/Tile_X0Y0_NN4BEG[6] Tile_X7Y7_DSP/Tile_X0Y0_NN4BEG[7]
+ Tile_X7Y7_DSP/Tile_X0Y0_NN4BEG[8] Tile_X7Y7_DSP/Tile_X0Y0_NN4BEG[9] Tile_X7Y7_DSP/Tile_X0Y0_S1END[0]
+ Tile_X7Y7_DSP/Tile_X0Y0_S1END[1] Tile_X7Y7_DSP/Tile_X0Y0_S1END[2] Tile_X7Y7_DSP/Tile_X0Y0_S1END[3]
+ Tile_X7Y7_DSP/Tile_X0Y0_S2MID[0] Tile_X7Y7_DSP/Tile_X0Y0_S2MID[1] Tile_X7Y7_DSP/Tile_X0Y0_S2MID[2]
+ Tile_X7Y7_DSP/Tile_X0Y0_S2MID[3] Tile_X7Y7_DSP/Tile_X0Y0_S2MID[4] Tile_X7Y7_DSP/Tile_X0Y0_S2MID[5]
+ Tile_X7Y7_DSP/Tile_X0Y0_S2MID[6] Tile_X7Y7_DSP/Tile_X0Y0_S2MID[7] Tile_X7Y7_DSP/Tile_X0Y0_S2END[0]
+ Tile_X7Y7_DSP/Tile_X0Y0_S2END[1] Tile_X7Y7_DSP/Tile_X0Y0_S2END[2] Tile_X7Y7_DSP/Tile_X0Y0_S2END[3]
+ Tile_X7Y7_DSP/Tile_X0Y0_S2END[4] Tile_X7Y7_DSP/Tile_X0Y0_S2END[5] Tile_X7Y7_DSP/Tile_X0Y0_S2END[6]
+ Tile_X7Y7_DSP/Tile_X0Y0_S2END[7] Tile_X7Y7_DSP/Tile_X0Y0_S4END[0] Tile_X7Y7_DSP/Tile_X0Y0_S4END[10]
+ Tile_X7Y7_DSP/Tile_X0Y0_S4END[11] Tile_X7Y7_DSP/Tile_X0Y0_S4END[12] Tile_X7Y7_DSP/Tile_X0Y0_S4END[13]
+ Tile_X7Y7_DSP/Tile_X0Y0_S4END[14] Tile_X7Y7_DSP/Tile_X0Y0_S4END[15] Tile_X7Y7_DSP/Tile_X0Y0_S4END[1]
+ Tile_X7Y7_DSP/Tile_X0Y0_S4END[2] Tile_X7Y7_DSP/Tile_X0Y0_S4END[3] Tile_X7Y7_DSP/Tile_X0Y0_S4END[4]
+ Tile_X7Y7_DSP/Tile_X0Y0_S4END[5] Tile_X7Y7_DSP/Tile_X0Y0_S4END[6] Tile_X7Y7_DSP/Tile_X0Y0_S4END[7]
+ Tile_X7Y7_DSP/Tile_X0Y0_S4END[8] Tile_X7Y7_DSP/Tile_X0Y0_S4END[9] Tile_X7Y7_DSP/Tile_X0Y0_SS4END[0]
+ Tile_X7Y7_DSP/Tile_X0Y0_SS4END[10] Tile_X7Y7_DSP/Tile_X0Y0_SS4END[11] Tile_X7Y7_DSP/Tile_X0Y0_SS4END[12]
+ Tile_X7Y7_DSP/Tile_X0Y0_SS4END[13] Tile_X7Y7_DSP/Tile_X0Y0_SS4END[14] Tile_X7Y7_DSP/Tile_X0Y0_SS4END[15]
+ Tile_X7Y7_DSP/Tile_X0Y0_SS4END[1] Tile_X7Y7_DSP/Tile_X0Y0_SS4END[2] Tile_X7Y7_DSP/Tile_X0Y0_SS4END[3]
+ Tile_X7Y7_DSP/Tile_X0Y0_SS4END[4] Tile_X7Y7_DSP/Tile_X0Y0_SS4END[5] Tile_X7Y7_DSP/Tile_X0Y0_SS4END[6]
+ Tile_X7Y7_DSP/Tile_X0Y0_SS4END[7] Tile_X7Y7_DSP/Tile_X0Y0_SS4END[8] Tile_X7Y7_DSP/Tile_X0Y0_SS4END[9]
+ Tile_X7Y5_DSP/Tile_X0Y1_UserCLK Tile_X6Y6_LUT4AB/W1END[0] Tile_X6Y6_LUT4AB/W1END[1]
+ Tile_X6Y6_LUT4AB/W1END[2] Tile_X6Y6_LUT4AB/W1END[3] Tile_X8Y6_LUT4AB/W1BEG[0] Tile_X8Y6_LUT4AB/W1BEG[1]
+ Tile_X8Y6_LUT4AB/W1BEG[2] Tile_X8Y6_LUT4AB/W1BEG[3] Tile_X6Y6_LUT4AB/W2MID[0] Tile_X6Y6_LUT4AB/W2MID[1]
+ Tile_X6Y6_LUT4AB/W2MID[2] Tile_X6Y6_LUT4AB/W2MID[3] Tile_X6Y6_LUT4AB/W2MID[4] Tile_X6Y6_LUT4AB/W2MID[5]
+ Tile_X6Y6_LUT4AB/W2MID[6] Tile_X6Y6_LUT4AB/W2MID[7] Tile_X6Y6_LUT4AB/W2END[0] Tile_X6Y6_LUT4AB/W2END[1]
+ Tile_X6Y6_LUT4AB/W2END[2] Tile_X6Y6_LUT4AB/W2END[3] Tile_X6Y6_LUT4AB/W2END[4] Tile_X6Y6_LUT4AB/W2END[5]
+ Tile_X6Y6_LUT4AB/W2END[6] Tile_X6Y6_LUT4AB/W2END[7] Tile_X8Y6_LUT4AB/W2BEGb[0] Tile_X8Y6_LUT4AB/W2BEGb[1]
+ Tile_X8Y6_LUT4AB/W2BEGb[2] Tile_X8Y6_LUT4AB/W2BEGb[3] Tile_X8Y6_LUT4AB/W2BEGb[4]
+ Tile_X8Y6_LUT4AB/W2BEGb[5] Tile_X8Y6_LUT4AB/W2BEGb[6] Tile_X8Y6_LUT4AB/W2BEGb[7]
+ Tile_X8Y6_LUT4AB/W2BEG[0] Tile_X8Y6_LUT4AB/W2BEG[1] Tile_X8Y6_LUT4AB/W2BEG[2] Tile_X8Y6_LUT4AB/W2BEG[3]
+ Tile_X8Y6_LUT4AB/W2BEG[4] Tile_X8Y6_LUT4AB/W2BEG[5] Tile_X8Y6_LUT4AB/W2BEG[6] Tile_X8Y6_LUT4AB/W2BEG[7]
+ Tile_X6Y6_LUT4AB/W6END[0] Tile_X6Y6_LUT4AB/W6END[10] Tile_X6Y6_LUT4AB/W6END[11]
+ Tile_X6Y6_LUT4AB/W6END[1] Tile_X6Y6_LUT4AB/W6END[2] Tile_X6Y6_LUT4AB/W6END[3] Tile_X6Y6_LUT4AB/W6END[4]
+ Tile_X6Y6_LUT4AB/W6END[5] Tile_X6Y6_LUT4AB/W6END[6] Tile_X6Y6_LUT4AB/W6END[7] Tile_X6Y6_LUT4AB/W6END[8]
+ Tile_X6Y6_LUT4AB/W6END[9] Tile_X8Y6_LUT4AB/W6BEG[0] Tile_X8Y6_LUT4AB/W6BEG[10] Tile_X8Y6_LUT4AB/W6BEG[11]
+ Tile_X8Y6_LUT4AB/W6BEG[1] Tile_X8Y6_LUT4AB/W6BEG[2] Tile_X8Y6_LUT4AB/W6BEG[3] Tile_X8Y6_LUT4AB/W6BEG[4]
+ Tile_X8Y6_LUT4AB/W6BEG[5] Tile_X8Y6_LUT4AB/W6BEG[6] Tile_X8Y6_LUT4AB/W6BEG[7] Tile_X8Y6_LUT4AB/W6BEG[8]
+ Tile_X8Y6_LUT4AB/W6BEG[9] Tile_X6Y6_LUT4AB/WW4END[0] Tile_X6Y6_LUT4AB/WW4END[10]
+ Tile_X6Y6_LUT4AB/WW4END[11] Tile_X6Y6_LUT4AB/WW4END[12] Tile_X6Y6_LUT4AB/WW4END[13]
+ Tile_X6Y6_LUT4AB/WW4END[14] Tile_X6Y6_LUT4AB/WW4END[15] Tile_X6Y6_LUT4AB/WW4END[1]
+ Tile_X6Y6_LUT4AB/WW4END[2] Tile_X6Y6_LUT4AB/WW4END[3] Tile_X6Y6_LUT4AB/WW4END[4]
+ Tile_X6Y6_LUT4AB/WW4END[5] Tile_X6Y6_LUT4AB/WW4END[6] Tile_X6Y6_LUT4AB/WW4END[7]
+ Tile_X6Y6_LUT4AB/WW4END[8] Tile_X6Y6_LUT4AB/WW4END[9] Tile_X8Y6_LUT4AB/WW4BEG[0]
+ Tile_X8Y6_LUT4AB/WW4BEG[10] Tile_X8Y6_LUT4AB/WW4BEG[11] Tile_X8Y6_LUT4AB/WW4BEG[12]
+ Tile_X8Y6_LUT4AB/WW4BEG[13] Tile_X8Y6_LUT4AB/WW4BEG[14] Tile_X8Y6_LUT4AB/WW4BEG[15]
+ Tile_X8Y6_LUT4AB/WW4BEG[1] Tile_X8Y6_LUT4AB/WW4BEG[2] Tile_X8Y6_LUT4AB/WW4BEG[3]
+ Tile_X8Y6_LUT4AB/WW4BEG[4] Tile_X8Y6_LUT4AB/WW4BEG[5] Tile_X8Y6_LUT4AB/WW4BEG[6]
+ Tile_X8Y6_LUT4AB/WW4BEG[7] Tile_X8Y6_LUT4AB/WW4BEG[8] Tile_X8Y6_LUT4AB/WW4BEG[9]
+ VGND VPWR DSP
XTile_X10Y13_IHP_SRAM Tile_X10Y14_ADDR_SRAM0 Tile_X10Y14_ADDR_SRAM1 Tile_X10Y14_ADDR_SRAM2
+ Tile_X10Y14_ADDR_SRAM3 Tile_X10Y14_ADDR_SRAM4 Tile_X10Y14_ADDR_SRAM5 Tile_X10Y14_ADDR_SRAM6
+ Tile_X10Y14_ADDR_SRAM7 Tile_X10Y14_ADDR_SRAM8 Tile_X10Y14_ADDR_SRAM9 Tile_X10Y14_BM_SRAM0
+ Tile_X10Y14_BM_SRAM1 Tile_X10Y14_BM_SRAM10 Tile_X10Y14_BM_SRAM11 Tile_X10Y14_BM_SRAM12
+ Tile_X10Y14_BM_SRAM13 Tile_X10Y14_BM_SRAM14 Tile_X10Y14_BM_SRAM15 Tile_X10Y14_BM_SRAM16
+ Tile_X10Y14_BM_SRAM17 Tile_X10Y14_BM_SRAM18 Tile_X10Y14_BM_SRAM19 Tile_X10Y14_BM_SRAM2
+ Tile_X10Y14_BM_SRAM20 Tile_X10Y14_BM_SRAM21 Tile_X10Y14_BM_SRAM22 Tile_X10Y14_BM_SRAM23
+ Tile_X10Y14_BM_SRAM24 Tile_X10Y14_BM_SRAM25 Tile_X10Y14_BM_SRAM26 Tile_X10Y14_BM_SRAM27
+ Tile_X10Y14_BM_SRAM28 Tile_X10Y14_BM_SRAM29 Tile_X10Y14_BM_SRAM3 Tile_X10Y14_BM_SRAM30
+ Tile_X10Y14_BM_SRAM31 Tile_X10Y14_BM_SRAM4 Tile_X10Y14_BM_SRAM5 Tile_X10Y14_BM_SRAM6
+ Tile_X10Y14_BM_SRAM7 Tile_X10Y14_BM_SRAM8 Tile_X10Y14_BM_SRAM9 Tile_X10Y14_CLK_SRAM
+ Tile_X10Y14_CONFIGURED_top Tile_X10Y14_DIN_SRAM0 Tile_X10Y14_DIN_SRAM1 Tile_X10Y14_DIN_SRAM10
+ Tile_X10Y14_DIN_SRAM11 Tile_X10Y14_DIN_SRAM12 Tile_X10Y14_DIN_SRAM13 Tile_X10Y14_DIN_SRAM14
+ Tile_X10Y14_DIN_SRAM15 Tile_X10Y14_DIN_SRAM16 Tile_X10Y14_DIN_SRAM17 Tile_X10Y14_DIN_SRAM18
+ Tile_X10Y14_DIN_SRAM19 Tile_X10Y14_DIN_SRAM2 Tile_X10Y14_DIN_SRAM20 Tile_X10Y14_DIN_SRAM21
+ Tile_X10Y14_DIN_SRAM22 Tile_X10Y14_DIN_SRAM23 Tile_X10Y14_DIN_SRAM24 Tile_X10Y14_DIN_SRAM25
+ Tile_X10Y14_DIN_SRAM26 Tile_X10Y14_DIN_SRAM27 Tile_X10Y14_DIN_SRAM28 Tile_X10Y14_DIN_SRAM29
+ Tile_X10Y14_DIN_SRAM3 Tile_X10Y14_DIN_SRAM30 Tile_X10Y14_DIN_SRAM31 Tile_X10Y14_DIN_SRAM4
+ Tile_X10Y14_DIN_SRAM5 Tile_X10Y14_DIN_SRAM6 Tile_X10Y14_DIN_SRAM7 Tile_X10Y14_DIN_SRAM8
+ Tile_X10Y14_DIN_SRAM9 Tile_X10Y14_DOUT_SRAM0 Tile_X10Y14_DOUT_SRAM1 Tile_X10Y14_DOUT_SRAM10
+ Tile_X10Y14_DOUT_SRAM11 Tile_X10Y14_DOUT_SRAM12 Tile_X10Y14_DOUT_SRAM13 Tile_X10Y14_DOUT_SRAM14
+ Tile_X10Y14_DOUT_SRAM15 Tile_X10Y14_DOUT_SRAM16 Tile_X10Y14_DOUT_SRAM17 Tile_X10Y14_DOUT_SRAM18
+ Tile_X10Y14_DOUT_SRAM19 Tile_X10Y14_DOUT_SRAM2 Tile_X10Y14_DOUT_SRAM20 Tile_X10Y14_DOUT_SRAM21
+ Tile_X10Y14_DOUT_SRAM22 Tile_X10Y14_DOUT_SRAM23 Tile_X10Y14_DOUT_SRAM24 Tile_X10Y14_DOUT_SRAM25
+ Tile_X10Y14_DOUT_SRAM26 Tile_X10Y14_DOUT_SRAM27 Tile_X10Y14_DOUT_SRAM28 Tile_X10Y14_DOUT_SRAM29
+ Tile_X10Y14_DOUT_SRAM3 Tile_X10Y14_DOUT_SRAM30 Tile_X10Y14_DOUT_SRAM31 Tile_X10Y14_DOUT_SRAM4
+ Tile_X10Y14_DOUT_SRAM5 Tile_X10Y14_DOUT_SRAM6 Tile_X10Y14_DOUT_SRAM7 Tile_X10Y14_DOUT_SRAM8
+ Tile_X10Y14_DOUT_SRAM9 Tile_X10Y14_MEN_SRAM Tile_X10Y14_REN_SRAM Tile_X10Y14_TIE_HIGH_SRAM
+ Tile_X10Y14_TIE_LOW_SRAM Tile_X9Y13_LUT4AB/E1BEG[0] Tile_X9Y13_LUT4AB/E1BEG[1] Tile_X9Y13_LUT4AB/E1BEG[2]
+ Tile_X9Y13_LUT4AB/E1BEG[3] Tile_X9Y13_LUT4AB/E2BEGb[0] Tile_X9Y13_LUT4AB/E2BEGb[1]
+ Tile_X9Y13_LUT4AB/E2BEGb[2] Tile_X9Y13_LUT4AB/E2BEGb[3] Tile_X9Y13_LUT4AB/E2BEGb[4]
+ Tile_X9Y13_LUT4AB/E2BEGb[5] Tile_X9Y13_LUT4AB/E2BEGb[6] Tile_X9Y13_LUT4AB/E2BEGb[7]
+ Tile_X9Y13_LUT4AB/E2BEG[0] Tile_X9Y13_LUT4AB/E2BEG[1] Tile_X9Y13_LUT4AB/E2BEG[2]
+ Tile_X9Y13_LUT4AB/E2BEG[3] Tile_X9Y13_LUT4AB/E2BEG[4] Tile_X9Y13_LUT4AB/E2BEG[5]
+ Tile_X9Y13_LUT4AB/E2BEG[6] Tile_X9Y13_LUT4AB/E2BEG[7] Tile_X9Y13_LUT4AB/E6BEG[0]
+ Tile_X9Y13_LUT4AB/E6BEG[10] Tile_X9Y13_LUT4AB/E6BEG[11] Tile_X9Y13_LUT4AB/E6BEG[1]
+ Tile_X9Y13_LUT4AB/E6BEG[2] Tile_X9Y13_LUT4AB/E6BEG[3] Tile_X9Y13_LUT4AB/E6BEG[4]
+ Tile_X9Y13_LUT4AB/E6BEG[5] Tile_X9Y13_LUT4AB/E6BEG[6] Tile_X9Y13_LUT4AB/E6BEG[7]
+ Tile_X9Y13_LUT4AB/E6BEG[8] Tile_X9Y13_LUT4AB/E6BEG[9] Tile_X9Y13_LUT4AB/EE4BEG[0]
+ Tile_X9Y13_LUT4AB/EE4BEG[10] Tile_X9Y13_LUT4AB/EE4BEG[11] Tile_X9Y13_LUT4AB/EE4BEG[12]
+ Tile_X9Y13_LUT4AB/EE4BEG[13] Tile_X9Y13_LUT4AB/EE4BEG[14] Tile_X9Y13_LUT4AB/EE4BEG[15]
+ Tile_X9Y13_LUT4AB/EE4BEG[1] Tile_X9Y13_LUT4AB/EE4BEG[2] Tile_X9Y13_LUT4AB/EE4BEG[3]
+ Tile_X9Y13_LUT4AB/EE4BEG[4] Tile_X9Y13_LUT4AB/EE4BEG[5] Tile_X9Y13_LUT4AB/EE4BEG[6]
+ Tile_X9Y13_LUT4AB/EE4BEG[7] Tile_X9Y13_LUT4AB/EE4BEG[8] Tile_X9Y13_LUT4AB/EE4BEG[9]
+ Tile_X9Y13_LUT4AB/FrameData_O[0] Tile_X9Y13_LUT4AB/FrameData_O[10] Tile_X9Y13_LUT4AB/FrameData_O[11]
+ Tile_X9Y13_LUT4AB/FrameData_O[12] Tile_X9Y13_LUT4AB/FrameData_O[13] Tile_X9Y13_LUT4AB/FrameData_O[14]
+ Tile_X9Y13_LUT4AB/FrameData_O[15] Tile_X9Y13_LUT4AB/FrameData_O[16] Tile_X9Y13_LUT4AB/FrameData_O[17]
+ Tile_X9Y13_LUT4AB/FrameData_O[18] Tile_X9Y13_LUT4AB/FrameData_O[19] Tile_X9Y13_LUT4AB/FrameData_O[1]
+ Tile_X9Y13_LUT4AB/FrameData_O[20] Tile_X9Y13_LUT4AB/FrameData_O[21] Tile_X9Y13_LUT4AB/FrameData_O[22]
+ Tile_X9Y13_LUT4AB/FrameData_O[23] Tile_X9Y13_LUT4AB/FrameData_O[24] Tile_X9Y13_LUT4AB/FrameData_O[25]
+ Tile_X9Y13_LUT4AB/FrameData_O[26] Tile_X9Y13_LUT4AB/FrameData_O[27] Tile_X9Y13_LUT4AB/FrameData_O[28]
+ Tile_X9Y13_LUT4AB/FrameData_O[29] Tile_X9Y13_LUT4AB/FrameData_O[2] Tile_X9Y13_LUT4AB/FrameData_O[30]
+ Tile_X9Y13_LUT4AB/FrameData_O[31] Tile_X9Y13_LUT4AB/FrameData_O[3] Tile_X9Y13_LUT4AB/FrameData_O[4]
+ Tile_X9Y13_LUT4AB/FrameData_O[5] Tile_X9Y13_LUT4AB/FrameData_O[6] Tile_X9Y13_LUT4AB/FrameData_O[7]
+ Tile_X9Y13_LUT4AB/FrameData_O[8] Tile_X9Y13_LUT4AB/FrameData_O[9] Tile_X10Y13_IHP_SRAM/Tile_X0Y0_FrameData_O[0]
+ Tile_X10Y13_IHP_SRAM/Tile_X0Y0_FrameData_O[10] Tile_X10Y13_IHP_SRAM/Tile_X0Y0_FrameData_O[11]
+ Tile_X10Y13_IHP_SRAM/Tile_X0Y0_FrameData_O[12] Tile_X10Y13_IHP_SRAM/Tile_X0Y0_FrameData_O[13]
+ Tile_X10Y13_IHP_SRAM/Tile_X0Y0_FrameData_O[14] Tile_X10Y13_IHP_SRAM/Tile_X0Y0_FrameData_O[15]
+ Tile_X10Y13_IHP_SRAM/Tile_X0Y0_FrameData_O[16] Tile_X10Y13_IHP_SRAM/Tile_X0Y0_FrameData_O[17]
+ Tile_X10Y13_IHP_SRAM/Tile_X0Y0_FrameData_O[18] Tile_X10Y13_IHP_SRAM/Tile_X0Y0_FrameData_O[19]
+ Tile_X10Y13_IHP_SRAM/Tile_X0Y0_FrameData_O[1] Tile_X10Y13_IHP_SRAM/Tile_X0Y0_FrameData_O[20]
+ Tile_X10Y13_IHP_SRAM/Tile_X0Y0_FrameData_O[21] Tile_X10Y13_IHP_SRAM/Tile_X0Y0_FrameData_O[22]
+ Tile_X10Y13_IHP_SRAM/Tile_X0Y0_FrameData_O[23] Tile_X10Y13_IHP_SRAM/Tile_X0Y0_FrameData_O[24]
+ Tile_X10Y13_IHP_SRAM/Tile_X0Y0_FrameData_O[25] Tile_X10Y13_IHP_SRAM/Tile_X0Y0_FrameData_O[26]
+ Tile_X10Y13_IHP_SRAM/Tile_X0Y0_FrameData_O[27] Tile_X10Y13_IHP_SRAM/Tile_X0Y0_FrameData_O[28]
+ Tile_X10Y13_IHP_SRAM/Tile_X0Y0_FrameData_O[29] Tile_X10Y13_IHP_SRAM/Tile_X0Y0_FrameData_O[2]
+ Tile_X10Y13_IHP_SRAM/Tile_X0Y0_FrameData_O[30] Tile_X10Y13_IHP_SRAM/Tile_X0Y0_FrameData_O[31]
+ Tile_X10Y13_IHP_SRAM/Tile_X0Y0_FrameData_O[3] Tile_X10Y13_IHP_SRAM/Tile_X0Y0_FrameData_O[4]
+ Tile_X10Y13_IHP_SRAM/Tile_X0Y0_FrameData_O[5] Tile_X10Y13_IHP_SRAM/Tile_X0Y0_FrameData_O[6]
+ Tile_X10Y13_IHP_SRAM/Tile_X0Y0_FrameData_O[7] Tile_X10Y13_IHP_SRAM/Tile_X0Y0_FrameData_O[8]
+ Tile_X10Y13_IHP_SRAM/Tile_X0Y0_FrameData_O[9] Tile_X10Y11_IHP_SRAM/Tile_X0Y1_FrameStrobe[0]
+ Tile_X10Y11_IHP_SRAM/Tile_X0Y1_FrameStrobe[10] Tile_X10Y11_IHP_SRAM/Tile_X0Y1_FrameStrobe[11]
+ Tile_X10Y11_IHP_SRAM/Tile_X0Y1_FrameStrobe[12] Tile_X10Y11_IHP_SRAM/Tile_X0Y1_FrameStrobe[13]
+ Tile_X10Y11_IHP_SRAM/Tile_X0Y1_FrameStrobe[14] Tile_X10Y11_IHP_SRAM/Tile_X0Y1_FrameStrobe[15]
+ Tile_X10Y11_IHP_SRAM/Tile_X0Y1_FrameStrobe[16] Tile_X10Y11_IHP_SRAM/Tile_X0Y1_FrameStrobe[17]
+ Tile_X10Y11_IHP_SRAM/Tile_X0Y1_FrameStrobe[18] Tile_X10Y11_IHP_SRAM/Tile_X0Y1_FrameStrobe[19]
+ Tile_X10Y11_IHP_SRAM/Tile_X0Y1_FrameStrobe[1] Tile_X10Y11_IHP_SRAM/Tile_X0Y1_FrameStrobe[2]
+ Tile_X10Y11_IHP_SRAM/Tile_X0Y1_FrameStrobe[3] Tile_X10Y11_IHP_SRAM/Tile_X0Y1_FrameStrobe[4]
+ Tile_X10Y11_IHP_SRAM/Tile_X0Y1_FrameStrobe[5] Tile_X10Y11_IHP_SRAM/Tile_X0Y1_FrameStrobe[6]
+ Tile_X10Y11_IHP_SRAM/Tile_X0Y1_FrameStrobe[7] Tile_X10Y11_IHP_SRAM/Tile_X0Y1_FrameStrobe[8]
+ Tile_X10Y11_IHP_SRAM/Tile_X0Y1_FrameStrobe[9] Tile_X10Y13_IHP_SRAM/Tile_X0Y0_N1BEG[0]
+ Tile_X10Y13_IHP_SRAM/Tile_X0Y0_N1BEG[1] Tile_X10Y13_IHP_SRAM/Tile_X0Y0_N1BEG[2]
+ Tile_X10Y13_IHP_SRAM/Tile_X0Y0_N1BEG[3] Tile_X10Y13_IHP_SRAM/Tile_X0Y0_N2BEG[0]
+ Tile_X10Y13_IHP_SRAM/Tile_X0Y0_N2BEG[1] Tile_X10Y13_IHP_SRAM/Tile_X0Y0_N2BEG[2]
+ Tile_X10Y13_IHP_SRAM/Tile_X0Y0_N2BEG[3] Tile_X10Y13_IHP_SRAM/Tile_X0Y0_N2BEG[4]
+ Tile_X10Y13_IHP_SRAM/Tile_X0Y0_N2BEG[5] Tile_X10Y13_IHP_SRAM/Tile_X0Y0_N2BEG[6]
+ Tile_X10Y13_IHP_SRAM/Tile_X0Y0_N2BEG[7] Tile_X10Y11_IHP_SRAM/Tile_X0Y1_N2END[0]
+ Tile_X10Y11_IHP_SRAM/Tile_X0Y1_N2END[1] Tile_X10Y11_IHP_SRAM/Tile_X0Y1_N2END[2]
+ Tile_X10Y11_IHP_SRAM/Tile_X0Y1_N2END[3] Tile_X10Y11_IHP_SRAM/Tile_X0Y1_N2END[4]
+ Tile_X10Y11_IHP_SRAM/Tile_X0Y1_N2END[5] Tile_X10Y11_IHP_SRAM/Tile_X0Y1_N2END[6]
+ Tile_X10Y11_IHP_SRAM/Tile_X0Y1_N2END[7] Tile_X10Y13_IHP_SRAM/Tile_X0Y0_N4BEG[0]
+ Tile_X10Y13_IHP_SRAM/Tile_X0Y0_N4BEG[10] Tile_X10Y13_IHP_SRAM/Tile_X0Y0_N4BEG[11]
+ Tile_X10Y13_IHP_SRAM/Tile_X0Y0_N4BEG[12] Tile_X10Y13_IHP_SRAM/Tile_X0Y0_N4BEG[13]
+ Tile_X10Y13_IHP_SRAM/Tile_X0Y0_N4BEG[14] Tile_X10Y13_IHP_SRAM/Tile_X0Y0_N4BEG[15]
+ Tile_X10Y13_IHP_SRAM/Tile_X0Y0_N4BEG[1] Tile_X10Y13_IHP_SRAM/Tile_X0Y0_N4BEG[2]
+ Tile_X10Y13_IHP_SRAM/Tile_X0Y0_N4BEG[3] Tile_X10Y13_IHP_SRAM/Tile_X0Y0_N4BEG[4]
+ Tile_X10Y13_IHP_SRAM/Tile_X0Y0_N4BEG[5] Tile_X10Y13_IHP_SRAM/Tile_X0Y0_N4BEG[6]
+ Tile_X10Y13_IHP_SRAM/Tile_X0Y0_N4BEG[7] Tile_X10Y13_IHP_SRAM/Tile_X0Y0_N4BEG[8]
+ Tile_X10Y13_IHP_SRAM/Tile_X0Y0_N4BEG[9] Tile_X10Y13_IHP_SRAM/Tile_X0Y0_S1END[0]
+ Tile_X10Y13_IHP_SRAM/Tile_X0Y0_S1END[1] Tile_X10Y13_IHP_SRAM/Tile_X0Y0_S1END[2]
+ Tile_X10Y13_IHP_SRAM/Tile_X0Y0_S1END[3] Tile_X10Y13_IHP_SRAM/Tile_X0Y0_S2END[0]
+ Tile_X10Y13_IHP_SRAM/Tile_X0Y0_S2END[1] Tile_X10Y13_IHP_SRAM/Tile_X0Y0_S2END[2]
+ Tile_X10Y13_IHP_SRAM/Tile_X0Y0_S2END[3] Tile_X10Y13_IHP_SRAM/Tile_X0Y0_S2END[4]
+ Tile_X10Y13_IHP_SRAM/Tile_X0Y0_S2END[5] Tile_X10Y13_IHP_SRAM/Tile_X0Y0_S2END[6]
+ Tile_X10Y13_IHP_SRAM/Tile_X0Y0_S2END[7] Tile_X10Y13_IHP_SRAM/Tile_X0Y0_S2MID[0]
+ Tile_X10Y13_IHP_SRAM/Tile_X0Y0_S2MID[1] Tile_X10Y13_IHP_SRAM/Tile_X0Y0_S2MID[2]
+ Tile_X10Y13_IHP_SRAM/Tile_X0Y0_S2MID[3] Tile_X10Y13_IHP_SRAM/Tile_X0Y0_S2MID[4]
+ Tile_X10Y13_IHP_SRAM/Tile_X0Y0_S2MID[5] Tile_X10Y13_IHP_SRAM/Tile_X0Y0_S2MID[6]
+ Tile_X10Y13_IHP_SRAM/Tile_X0Y0_S2MID[7] Tile_X10Y13_IHP_SRAM/Tile_X0Y0_S4END[0]
+ Tile_X10Y13_IHP_SRAM/Tile_X0Y0_S4END[10] Tile_X10Y13_IHP_SRAM/Tile_X0Y0_S4END[11]
+ Tile_X10Y13_IHP_SRAM/Tile_X0Y0_S4END[12] Tile_X10Y13_IHP_SRAM/Tile_X0Y0_S4END[13]
+ Tile_X10Y13_IHP_SRAM/Tile_X0Y0_S4END[14] Tile_X10Y13_IHP_SRAM/Tile_X0Y0_S4END[15]
+ Tile_X10Y13_IHP_SRAM/Tile_X0Y0_S4END[1] Tile_X10Y13_IHP_SRAM/Tile_X0Y0_S4END[2]
+ Tile_X10Y13_IHP_SRAM/Tile_X0Y0_S4END[3] Tile_X10Y13_IHP_SRAM/Tile_X0Y0_S4END[4]
+ Tile_X10Y13_IHP_SRAM/Tile_X0Y0_S4END[5] Tile_X10Y13_IHP_SRAM/Tile_X0Y0_S4END[6]
+ Tile_X10Y13_IHP_SRAM/Tile_X0Y0_S4END[7] Tile_X10Y13_IHP_SRAM/Tile_X0Y0_S4END[8]
+ Tile_X10Y13_IHP_SRAM/Tile_X0Y0_S4END[9] Tile_X10Y11_IHP_SRAM/Tile_X0Y1_UserCLK Tile_X9Y13_LUT4AB/W1END[0]
+ Tile_X9Y13_LUT4AB/W1END[1] Tile_X9Y13_LUT4AB/W1END[2] Tile_X9Y13_LUT4AB/W1END[3]
+ Tile_X9Y13_LUT4AB/W2MID[0] Tile_X9Y13_LUT4AB/W2MID[1] Tile_X9Y13_LUT4AB/W2MID[2]
+ Tile_X9Y13_LUT4AB/W2MID[3] Tile_X9Y13_LUT4AB/W2MID[4] Tile_X9Y13_LUT4AB/W2MID[5]
+ Tile_X9Y13_LUT4AB/W2MID[6] Tile_X9Y13_LUT4AB/W2MID[7] Tile_X9Y13_LUT4AB/W2END[0]
+ Tile_X9Y13_LUT4AB/W2END[1] Tile_X9Y13_LUT4AB/W2END[2] Tile_X9Y13_LUT4AB/W2END[3]
+ Tile_X9Y13_LUT4AB/W2END[4] Tile_X9Y13_LUT4AB/W2END[5] Tile_X9Y13_LUT4AB/W2END[6]
+ Tile_X9Y13_LUT4AB/W2END[7] Tile_X9Y13_LUT4AB/W6END[0] Tile_X9Y13_LUT4AB/W6END[10]
+ Tile_X9Y13_LUT4AB/W6END[11] Tile_X9Y13_LUT4AB/W6END[1] Tile_X9Y13_LUT4AB/W6END[2]
+ Tile_X9Y13_LUT4AB/W6END[3] Tile_X9Y13_LUT4AB/W6END[4] Tile_X9Y13_LUT4AB/W6END[5]
+ Tile_X9Y13_LUT4AB/W6END[6] Tile_X9Y13_LUT4AB/W6END[7] Tile_X9Y13_LUT4AB/W6END[8]
+ Tile_X9Y13_LUT4AB/W6END[9] Tile_X9Y13_LUT4AB/WW4END[0] Tile_X9Y13_LUT4AB/WW4END[10]
+ Tile_X9Y13_LUT4AB/WW4END[11] Tile_X9Y13_LUT4AB/WW4END[12] Tile_X9Y13_LUT4AB/WW4END[13]
+ Tile_X9Y13_LUT4AB/WW4END[14] Tile_X9Y13_LUT4AB/WW4END[15] Tile_X9Y13_LUT4AB/WW4END[1]
+ Tile_X9Y13_LUT4AB/WW4END[2] Tile_X9Y13_LUT4AB/WW4END[3] Tile_X9Y13_LUT4AB/WW4END[4]
+ Tile_X9Y13_LUT4AB/WW4END[5] Tile_X9Y13_LUT4AB/WW4END[6] Tile_X9Y13_LUT4AB/WW4END[7]
+ Tile_X9Y13_LUT4AB/WW4END[8] Tile_X9Y13_LUT4AB/WW4END[9] Tile_X9Y14_LUT4AB/E1BEG[0]
+ Tile_X9Y14_LUT4AB/E1BEG[1] Tile_X9Y14_LUT4AB/E1BEG[2] Tile_X9Y14_LUT4AB/E1BEG[3]
+ Tile_X9Y14_LUT4AB/E2BEGb[0] Tile_X9Y14_LUT4AB/E2BEGb[1] Tile_X9Y14_LUT4AB/E2BEGb[2]
+ Tile_X9Y14_LUT4AB/E2BEGb[3] Tile_X9Y14_LUT4AB/E2BEGb[4] Tile_X9Y14_LUT4AB/E2BEGb[5]
+ Tile_X9Y14_LUT4AB/E2BEGb[6] Tile_X9Y14_LUT4AB/E2BEGb[7] Tile_X9Y14_LUT4AB/E2BEG[0]
+ Tile_X9Y14_LUT4AB/E2BEG[1] Tile_X9Y14_LUT4AB/E2BEG[2] Tile_X9Y14_LUT4AB/E2BEG[3]
+ Tile_X9Y14_LUT4AB/E2BEG[4] Tile_X9Y14_LUT4AB/E2BEG[5] Tile_X9Y14_LUT4AB/E2BEG[6]
+ Tile_X9Y14_LUT4AB/E2BEG[7] Tile_X9Y14_LUT4AB/E6BEG[0] Tile_X9Y14_LUT4AB/E6BEG[10]
+ Tile_X9Y14_LUT4AB/E6BEG[11] Tile_X9Y14_LUT4AB/E6BEG[1] Tile_X9Y14_LUT4AB/E6BEG[2]
+ Tile_X9Y14_LUT4AB/E6BEG[3] Tile_X9Y14_LUT4AB/E6BEG[4] Tile_X9Y14_LUT4AB/E6BEG[5]
+ Tile_X9Y14_LUT4AB/E6BEG[6] Tile_X9Y14_LUT4AB/E6BEG[7] Tile_X9Y14_LUT4AB/E6BEG[8]
+ Tile_X9Y14_LUT4AB/E6BEG[9] Tile_X9Y14_LUT4AB/EE4BEG[0] Tile_X9Y14_LUT4AB/EE4BEG[10]
+ Tile_X9Y14_LUT4AB/EE4BEG[11] Tile_X9Y14_LUT4AB/EE4BEG[12] Tile_X9Y14_LUT4AB/EE4BEG[13]
+ Tile_X9Y14_LUT4AB/EE4BEG[14] Tile_X9Y14_LUT4AB/EE4BEG[15] Tile_X9Y14_LUT4AB/EE4BEG[1]
+ Tile_X9Y14_LUT4AB/EE4BEG[2] Tile_X9Y14_LUT4AB/EE4BEG[3] Tile_X9Y14_LUT4AB/EE4BEG[4]
+ Tile_X9Y14_LUT4AB/EE4BEG[5] Tile_X9Y14_LUT4AB/EE4BEG[6] Tile_X9Y14_LUT4AB/EE4BEG[7]
+ Tile_X9Y14_LUT4AB/EE4BEG[8] Tile_X9Y14_LUT4AB/EE4BEG[9] Tile_X9Y14_LUT4AB/FrameData_O[0]
+ Tile_X9Y14_LUT4AB/FrameData_O[10] Tile_X9Y14_LUT4AB/FrameData_O[11] Tile_X9Y14_LUT4AB/FrameData_O[12]
+ Tile_X9Y14_LUT4AB/FrameData_O[13] Tile_X9Y14_LUT4AB/FrameData_O[14] Tile_X9Y14_LUT4AB/FrameData_O[15]
+ Tile_X9Y14_LUT4AB/FrameData_O[16] Tile_X9Y14_LUT4AB/FrameData_O[17] Tile_X9Y14_LUT4AB/FrameData_O[18]
+ Tile_X9Y14_LUT4AB/FrameData_O[19] Tile_X9Y14_LUT4AB/FrameData_O[1] Tile_X9Y14_LUT4AB/FrameData_O[20]
+ Tile_X9Y14_LUT4AB/FrameData_O[21] Tile_X9Y14_LUT4AB/FrameData_O[22] Tile_X9Y14_LUT4AB/FrameData_O[23]
+ Tile_X9Y14_LUT4AB/FrameData_O[24] Tile_X9Y14_LUT4AB/FrameData_O[25] Tile_X9Y14_LUT4AB/FrameData_O[26]
+ Tile_X9Y14_LUT4AB/FrameData_O[27] Tile_X9Y14_LUT4AB/FrameData_O[28] Tile_X9Y14_LUT4AB/FrameData_O[29]
+ Tile_X9Y14_LUT4AB/FrameData_O[2] Tile_X9Y14_LUT4AB/FrameData_O[30] Tile_X9Y14_LUT4AB/FrameData_O[31]
+ Tile_X9Y14_LUT4AB/FrameData_O[3] Tile_X9Y14_LUT4AB/FrameData_O[4] Tile_X9Y14_LUT4AB/FrameData_O[5]
+ Tile_X9Y14_LUT4AB/FrameData_O[6] Tile_X9Y14_LUT4AB/FrameData_O[7] Tile_X9Y14_LUT4AB/FrameData_O[8]
+ Tile_X9Y14_LUT4AB/FrameData_O[9] Tile_X10Y13_IHP_SRAM/Tile_X0Y1_FrameData_O[0] Tile_X10Y13_IHP_SRAM/Tile_X0Y1_FrameData_O[10]
+ Tile_X10Y13_IHP_SRAM/Tile_X0Y1_FrameData_O[11] Tile_X10Y13_IHP_SRAM/Tile_X0Y1_FrameData_O[12]
+ Tile_X10Y13_IHP_SRAM/Tile_X0Y1_FrameData_O[13] Tile_X10Y13_IHP_SRAM/Tile_X0Y1_FrameData_O[14]
+ Tile_X10Y13_IHP_SRAM/Tile_X0Y1_FrameData_O[15] Tile_X10Y13_IHP_SRAM/Tile_X0Y1_FrameData_O[16]
+ Tile_X10Y13_IHP_SRAM/Tile_X0Y1_FrameData_O[17] Tile_X10Y13_IHP_SRAM/Tile_X0Y1_FrameData_O[18]
+ Tile_X10Y13_IHP_SRAM/Tile_X0Y1_FrameData_O[19] Tile_X10Y13_IHP_SRAM/Tile_X0Y1_FrameData_O[1]
+ Tile_X10Y13_IHP_SRAM/Tile_X0Y1_FrameData_O[20] Tile_X10Y13_IHP_SRAM/Tile_X0Y1_FrameData_O[21]
+ Tile_X10Y13_IHP_SRAM/Tile_X0Y1_FrameData_O[22] Tile_X10Y13_IHP_SRAM/Tile_X0Y1_FrameData_O[23]
+ Tile_X10Y13_IHP_SRAM/Tile_X0Y1_FrameData_O[24] Tile_X10Y13_IHP_SRAM/Tile_X0Y1_FrameData_O[25]
+ Tile_X10Y13_IHP_SRAM/Tile_X0Y1_FrameData_O[26] Tile_X10Y13_IHP_SRAM/Tile_X0Y1_FrameData_O[27]
+ Tile_X10Y13_IHP_SRAM/Tile_X0Y1_FrameData_O[28] Tile_X10Y13_IHP_SRAM/Tile_X0Y1_FrameData_O[29]
+ Tile_X10Y13_IHP_SRAM/Tile_X0Y1_FrameData_O[2] Tile_X10Y13_IHP_SRAM/Tile_X0Y1_FrameData_O[30]
+ Tile_X10Y13_IHP_SRAM/Tile_X0Y1_FrameData_O[31] Tile_X10Y13_IHP_SRAM/Tile_X0Y1_FrameData_O[3]
+ Tile_X10Y13_IHP_SRAM/Tile_X0Y1_FrameData_O[4] Tile_X10Y13_IHP_SRAM/Tile_X0Y1_FrameData_O[5]
+ Tile_X10Y13_IHP_SRAM/Tile_X0Y1_FrameData_O[6] Tile_X10Y13_IHP_SRAM/Tile_X0Y1_FrameData_O[7]
+ Tile_X10Y13_IHP_SRAM/Tile_X0Y1_FrameData_O[8] Tile_X10Y13_IHP_SRAM/Tile_X0Y1_FrameData_O[9]
+ Tile_X10Y15_S_term_IHP_SRAM/FrameStrobe_O[0] Tile_X10Y15_S_term_IHP_SRAM/FrameStrobe_O[10]
+ Tile_X10Y15_S_term_IHP_SRAM/FrameStrobe_O[11] Tile_X10Y15_S_term_IHP_SRAM/FrameStrobe_O[12]
+ Tile_X10Y15_S_term_IHP_SRAM/FrameStrobe_O[13] Tile_X10Y15_S_term_IHP_SRAM/FrameStrobe_O[14]
+ Tile_X10Y15_S_term_IHP_SRAM/FrameStrobe_O[15] Tile_X10Y15_S_term_IHP_SRAM/FrameStrobe_O[16]
+ Tile_X10Y15_S_term_IHP_SRAM/FrameStrobe_O[17] Tile_X10Y15_S_term_IHP_SRAM/FrameStrobe_O[18]
+ Tile_X10Y15_S_term_IHP_SRAM/FrameStrobe_O[19] Tile_X10Y15_S_term_IHP_SRAM/FrameStrobe_O[1]
+ Tile_X10Y15_S_term_IHP_SRAM/FrameStrobe_O[2] Tile_X10Y15_S_term_IHP_SRAM/FrameStrobe_O[3]
+ Tile_X10Y15_S_term_IHP_SRAM/FrameStrobe_O[4] Tile_X10Y15_S_term_IHP_SRAM/FrameStrobe_O[5]
+ Tile_X10Y15_S_term_IHP_SRAM/FrameStrobe_O[6] Tile_X10Y15_S_term_IHP_SRAM/FrameStrobe_O[7]
+ Tile_X10Y15_S_term_IHP_SRAM/FrameStrobe_O[8] Tile_X10Y15_S_term_IHP_SRAM/FrameStrobe_O[9]
+ Tile_X10Y15_S_term_IHP_SRAM/N1BEG[0] Tile_X10Y15_S_term_IHP_SRAM/N1BEG[1] Tile_X10Y15_S_term_IHP_SRAM/N1BEG[2]
+ Tile_X10Y15_S_term_IHP_SRAM/N1BEG[3] Tile_X10Y15_S_term_IHP_SRAM/N2BEGb[0] Tile_X10Y15_S_term_IHP_SRAM/N2BEGb[1]
+ Tile_X10Y15_S_term_IHP_SRAM/N2BEGb[2] Tile_X10Y15_S_term_IHP_SRAM/N2BEGb[3] Tile_X10Y15_S_term_IHP_SRAM/N2BEGb[4]
+ Tile_X10Y15_S_term_IHP_SRAM/N2BEGb[5] Tile_X10Y15_S_term_IHP_SRAM/N2BEGb[6] Tile_X10Y15_S_term_IHP_SRAM/N2BEGb[7]
+ Tile_X10Y15_S_term_IHP_SRAM/N2BEG[0] Tile_X10Y15_S_term_IHP_SRAM/N2BEG[1] Tile_X10Y15_S_term_IHP_SRAM/N2BEG[2]
+ Tile_X10Y15_S_term_IHP_SRAM/N2BEG[3] Tile_X10Y15_S_term_IHP_SRAM/N2BEG[4] Tile_X10Y15_S_term_IHP_SRAM/N2BEG[5]
+ Tile_X10Y15_S_term_IHP_SRAM/N2BEG[6] Tile_X10Y15_S_term_IHP_SRAM/N2BEG[7] Tile_X10Y15_S_term_IHP_SRAM/N4BEG[0]
+ Tile_X10Y15_S_term_IHP_SRAM/N4BEG[10] Tile_X10Y15_S_term_IHP_SRAM/N4BEG[11] Tile_X10Y15_S_term_IHP_SRAM/N4BEG[12]
+ Tile_X10Y15_S_term_IHP_SRAM/N4BEG[13] Tile_X10Y15_S_term_IHP_SRAM/N4BEG[14] Tile_X10Y15_S_term_IHP_SRAM/N4BEG[15]
+ Tile_X10Y15_S_term_IHP_SRAM/N4BEG[1] Tile_X10Y15_S_term_IHP_SRAM/N4BEG[2] Tile_X10Y15_S_term_IHP_SRAM/N4BEG[3]
+ Tile_X10Y15_S_term_IHP_SRAM/N4BEG[4] Tile_X10Y15_S_term_IHP_SRAM/N4BEG[5] Tile_X10Y15_S_term_IHP_SRAM/N4BEG[6]
+ Tile_X10Y15_S_term_IHP_SRAM/N4BEG[7] Tile_X10Y15_S_term_IHP_SRAM/N4BEG[8] Tile_X10Y15_S_term_IHP_SRAM/N4BEG[9]
+ Tile_X10Y15_S_term_IHP_SRAM/S1END[0] Tile_X10Y15_S_term_IHP_SRAM/S1END[1] Tile_X10Y15_S_term_IHP_SRAM/S1END[2]
+ Tile_X10Y15_S_term_IHP_SRAM/S1END[3] Tile_X10Y15_S_term_IHP_SRAM/S2MID[0] Tile_X10Y15_S_term_IHP_SRAM/S2MID[1]
+ Tile_X10Y15_S_term_IHP_SRAM/S2MID[2] Tile_X10Y15_S_term_IHP_SRAM/S2MID[3] Tile_X10Y15_S_term_IHP_SRAM/S2MID[4]
+ Tile_X10Y15_S_term_IHP_SRAM/S2MID[5] Tile_X10Y15_S_term_IHP_SRAM/S2MID[6] Tile_X10Y15_S_term_IHP_SRAM/S2MID[7]
+ Tile_X10Y15_S_term_IHP_SRAM/S2END[0] Tile_X10Y15_S_term_IHP_SRAM/S2END[1] Tile_X10Y15_S_term_IHP_SRAM/S2END[2]
+ Tile_X10Y15_S_term_IHP_SRAM/S2END[3] Tile_X10Y15_S_term_IHP_SRAM/S2END[4] Tile_X10Y15_S_term_IHP_SRAM/S2END[5]
+ Tile_X10Y15_S_term_IHP_SRAM/S2END[6] Tile_X10Y15_S_term_IHP_SRAM/S2END[7] Tile_X10Y15_S_term_IHP_SRAM/S4END[0]
+ Tile_X10Y15_S_term_IHP_SRAM/S4END[10] Tile_X10Y15_S_term_IHP_SRAM/S4END[11] Tile_X10Y15_S_term_IHP_SRAM/S4END[12]
+ Tile_X10Y15_S_term_IHP_SRAM/S4END[13] Tile_X10Y15_S_term_IHP_SRAM/S4END[14] Tile_X10Y15_S_term_IHP_SRAM/S4END[15]
+ Tile_X10Y15_S_term_IHP_SRAM/S4END[1] Tile_X10Y15_S_term_IHP_SRAM/S4END[2] Tile_X10Y15_S_term_IHP_SRAM/S4END[3]
+ Tile_X10Y15_S_term_IHP_SRAM/S4END[4] Tile_X10Y15_S_term_IHP_SRAM/S4END[5] Tile_X10Y15_S_term_IHP_SRAM/S4END[6]
+ Tile_X10Y15_S_term_IHP_SRAM/S4END[7] Tile_X10Y15_S_term_IHP_SRAM/S4END[8] Tile_X10Y15_S_term_IHP_SRAM/S4END[9]
+ Tile_X10Y15_S_term_IHP_SRAM/UserCLKo Tile_X9Y14_LUT4AB/W1END[0] Tile_X9Y14_LUT4AB/W1END[1]
+ Tile_X9Y14_LUT4AB/W1END[2] Tile_X9Y14_LUT4AB/W1END[3] Tile_X9Y14_LUT4AB/W2MID[0]
+ Tile_X9Y14_LUT4AB/W2MID[1] Tile_X9Y14_LUT4AB/W2MID[2] Tile_X9Y14_LUT4AB/W2MID[3]
+ Tile_X9Y14_LUT4AB/W2MID[4] Tile_X9Y14_LUT4AB/W2MID[5] Tile_X9Y14_LUT4AB/W2MID[6]
+ Tile_X9Y14_LUT4AB/W2MID[7] Tile_X9Y14_LUT4AB/W2END[0] Tile_X9Y14_LUT4AB/W2END[1]
+ Tile_X9Y14_LUT4AB/W2END[2] Tile_X9Y14_LUT4AB/W2END[3] Tile_X9Y14_LUT4AB/W2END[4]
+ Tile_X9Y14_LUT4AB/W2END[5] Tile_X9Y14_LUT4AB/W2END[6] Tile_X9Y14_LUT4AB/W2END[7]
+ Tile_X9Y14_LUT4AB/W6END[0] Tile_X9Y14_LUT4AB/W6END[10] Tile_X9Y14_LUT4AB/W6END[11]
+ Tile_X9Y14_LUT4AB/W6END[1] Tile_X9Y14_LUT4AB/W6END[2] Tile_X9Y14_LUT4AB/W6END[3]
+ Tile_X9Y14_LUT4AB/W6END[4] Tile_X9Y14_LUT4AB/W6END[5] Tile_X9Y14_LUT4AB/W6END[6]
+ Tile_X9Y14_LUT4AB/W6END[7] Tile_X9Y14_LUT4AB/W6END[8] Tile_X9Y14_LUT4AB/W6END[9]
+ Tile_X9Y14_LUT4AB/WW4END[0] Tile_X9Y14_LUT4AB/WW4END[10] Tile_X9Y14_LUT4AB/WW4END[11]
+ Tile_X9Y14_LUT4AB/WW4END[12] Tile_X9Y14_LUT4AB/WW4END[13] Tile_X9Y14_LUT4AB/WW4END[14]
+ Tile_X9Y14_LUT4AB/WW4END[15] Tile_X9Y14_LUT4AB/WW4END[1] Tile_X9Y14_LUT4AB/WW4END[2]
+ Tile_X9Y14_LUT4AB/WW4END[3] Tile_X9Y14_LUT4AB/WW4END[4] Tile_X9Y14_LUT4AB/WW4END[5]
+ Tile_X9Y14_LUT4AB/WW4END[6] Tile_X9Y14_LUT4AB/WW4END[7] Tile_X9Y14_LUT4AB/WW4END[8]
+ Tile_X9Y14_LUT4AB/WW4END[9] VGND VPWR Tile_X10Y14_WEN_SRAM IHP_SRAM
XTile_X4Y7_RegFile Tile_X5Y7_LUT4AB/E1END[0] Tile_X5Y7_LUT4AB/E1END[1] Tile_X5Y7_LUT4AB/E1END[2]
+ Tile_X5Y7_LUT4AB/E1END[3] Tile_X3Y7_LUT4AB/E1BEG[0] Tile_X3Y7_LUT4AB/E1BEG[1] Tile_X3Y7_LUT4AB/E1BEG[2]
+ Tile_X3Y7_LUT4AB/E1BEG[3] Tile_X5Y7_LUT4AB/E2MID[0] Tile_X5Y7_LUT4AB/E2MID[1] Tile_X5Y7_LUT4AB/E2MID[2]
+ Tile_X5Y7_LUT4AB/E2MID[3] Tile_X5Y7_LUT4AB/E2MID[4] Tile_X5Y7_LUT4AB/E2MID[5] Tile_X5Y7_LUT4AB/E2MID[6]
+ Tile_X5Y7_LUT4AB/E2MID[7] Tile_X5Y7_LUT4AB/E2END[0] Tile_X5Y7_LUT4AB/E2END[1] Tile_X5Y7_LUT4AB/E2END[2]
+ Tile_X5Y7_LUT4AB/E2END[3] Tile_X5Y7_LUT4AB/E2END[4] Tile_X5Y7_LUT4AB/E2END[5] Tile_X5Y7_LUT4AB/E2END[6]
+ Tile_X5Y7_LUT4AB/E2END[7] Tile_X4Y7_RegFile/E2END[0] Tile_X4Y7_RegFile/E2END[1]
+ Tile_X4Y7_RegFile/E2END[2] Tile_X4Y7_RegFile/E2END[3] Tile_X4Y7_RegFile/E2END[4]
+ Tile_X4Y7_RegFile/E2END[5] Tile_X4Y7_RegFile/E2END[6] Tile_X4Y7_RegFile/E2END[7]
+ Tile_X3Y7_LUT4AB/E2BEG[0] Tile_X3Y7_LUT4AB/E2BEG[1] Tile_X3Y7_LUT4AB/E2BEG[2] Tile_X3Y7_LUT4AB/E2BEG[3]
+ Tile_X3Y7_LUT4AB/E2BEG[4] Tile_X3Y7_LUT4AB/E2BEG[5] Tile_X3Y7_LUT4AB/E2BEG[6] Tile_X3Y7_LUT4AB/E2BEG[7]
+ Tile_X5Y7_LUT4AB/E6END[0] Tile_X5Y7_LUT4AB/E6END[10] Tile_X5Y7_LUT4AB/E6END[11]
+ Tile_X5Y7_LUT4AB/E6END[1] Tile_X5Y7_LUT4AB/E6END[2] Tile_X5Y7_LUT4AB/E6END[3] Tile_X5Y7_LUT4AB/E6END[4]
+ Tile_X5Y7_LUT4AB/E6END[5] Tile_X5Y7_LUT4AB/E6END[6] Tile_X5Y7_LUT4AB/E6END[7] Tile_X5Y7_LUT4AB/E6END[8]
+ Tile_X5Y7_LUT4AB/E6END[9] Tile_X3Y7_LUT4AB/E6BEG[0] Tile_X3Y7_LUT4AB/E6BEG[10] Tile_X3Y7_LUT4AB/E6BEG[11]
+ Tile_X3Y7_LUT4AB/E6BEG[1] Tile_X3Y7_LUT4AB/E6BEG[2] Tile_X3Y7_LUT4AB/E6BEG[3] Tile_X3Y7_LUT4AB/E6BEG[4]
+ Tile_X3Y7_LUT4AB/E6BEG[5] Tile_X3Y7_LUT4AB/E6BEG[6] Tile_X3Y7_LUT4AB/E6BEG[7] Tile_X3Y7_LUT4AB/E6BEG[8]
+ Tile_X3Y7_LUT4AB/E6BEG[9] Tile_X5Y7_LUT4AB/EE4END[0] Tile_X5Y7_LUT4AB/EE4END[10]
+ Tile_X5Y7_LUT4AB/EE4END[11] Tile_X5Y7_LUT4AB/EE4END[12] Tile_X5Y7_LUT4AB/EE4END[13]
+ Tile_X5Y7_LUT4AB/EE4END[14] Tile_X5Y7_LUT4AB/EE4END[15] Tile_X5Y7_LUT4AB/EE4END[1]
+ Tile_X5Y7_LUT4AB/EE4END[2] Tile_X5Y7_LUT4AB/EE4END[3] Tile_X5Y7_LUT4AB/EE4END[4]
+ Tile_X5Y7_LUT4AB/EE4END[5] Tile_X5Y7_LUT4AB/EE4END[6] Tile_X5Y7_LUT4AB/EE4END[7]
+ Tile_X5Y7_LUT4AB/EE4END[8] Tile_X5Y7_LUT4AB/EE4END[9] Tile_X3Y7_LUT4AB/EE4BEG[0]
+ Tile_X3Y7_LUT4AB/EE4BEG[10] Tile_X3Y7_LUT4AB/EE4BEG[11] Tile_X3Y7_LUT4AB/EE4BEG[12]
+ Tile_X3Y7_LUT4AB/EE4BEG[13] Tile_X3Y7_LUT4AB/EE4BEG[14] Tile_X3Y7_LUT4AB/EE4BEG[15]
+ Tile_X3Y7_LUT4AB/EE4BEG[1] Tile_X3Y7_LUT4AB/EE4BEG[2] Tile_X3Y7_LUT4AB/EE4BEG[3]
+ Tile_X3Y7_LUT4AB/EE4BEG[4] Tile_X3Y7_LUT4AB/EE4BEG[5] Tile_X3Y7_LUT4AB/EE4BEG[6]
+ Tile_X3Y7_LUT4AB/EE4BEG[7] Tile_X3Y7_LUT4AB/EE4BEG[8] Tile_X3Y7_LUT4AB/EE4BEG[9]
+ Tile_X4Y7_RegFile/FrameData[0] Tile_X4Y7_RegFile/FrameData[10] Tile_X4Y7_RegFile/FrameData[11]
+ Tile_X4Y7_RegFile/FrameData[12] Tile_X4Y7_RegFile/FrameData[13] Tile_X4Y7_RegFile/FrameData[14]
+ Tile_X4Y7_RegFile/FrameData[15] Tile_X4Y7_RegFile/FrameData[16] Tile_X4Y7_RegFile/FrameData[17]
+ Tile_X4Y7_RegFile/FrameData[18] Tile_X4Y7_RegFile/FrameData[19] Tile_X4Y7_RegFile/FrameData[1]
+ Tile_X4Y7_RegFile/FrameData[20] Tile_X4Y7_RegFile/FrameData[21] Tile_X4Y7_RegFile/FrameData[22]
+ Tile_X4Y7_RegFile/FrameData[23] Tile_X4Y7_RegFile/FrameData[24] Tile_X4Y7_RegFile/FrameData[25]
+ Tile_X4Y7_RegFile/FrameData[26] Tile_X4Y7_RegFile/FrameData[27] Tile_X4Y7_RegFile/FrameData[28]
+ Tile_X4Y7_RegFile/FrameData[29] Tile_X4Y7_RegFile/FrameData[2] Tile_X4Y7_RegFile/FrameData[30]
+ Tile_X4Y7_RegFile/FrameData[31] Tile_X4Y7_RegFile/FrameData[3] Tile_X4Y7_RegFile/FrameData[4]
+ Tile_X4Y7_RegFile/FrameData[5] Tile_X4Y7_RegFile/FrameData[6] Tile_X4Y7_RegFile/FrameData[7]
+ Tile_X4Y7_RegFile/FrameData[8] Tile_X4Y7_RegFile/FrameData[9] Tile_X5Y7_LUT4AB/FrameData[0]
+ Tile_X5Y7_LUT4AB/FrameData[10] Tile_X5Y7_LUT4AB/FrameData[11] Tile_X5Y7_LUT4AB/FrameData[12]
+ Tile_X5Y7_LUT4AB/FrameData[13] Tile_X5Y7_LUT4AB/FrameData[14] Tile_X5Y7_LUT4AB/FrameData[15]
+ Tile_X5Y7_LUT4AB/FrameData[16] Tile_X5Y7_LUT4AB/FrameData[17] Tile_X5Y7_LUT4AB/FrameData[18]
+ Tile_X5Y7_LUT4AB/FrameData[19] Tile_X5Y7_LUT4AB/FrameData[1] Tile_X5Y7_LUT4AB/FrameData[20]
+ Tile_X5Y7_LUT4AB/FrameData[21] Tile_X5Y7_LUT4AB/FrameData[22] Tile_X5Y7_LUT4AB/FrameData[23]
+ Tile_X5Y7_LUT4AB/FrameData[24] Tile_X5Y7_LUT4AB/FrameData[25] Tile_X5Y7_LUT4AB/FrameData[26]
+ Tile_X5Y7_LUT4AB/FrameData[27] Tile_X5Y7_LUT4AB/FrameData[28] Tile_X5Y7_LUT4AB/FrameData[29]
+ Tile_X5Y7_LUT4AB/FrameData[2] Tile_X5Y7_LUT4AB/FrameData[30] Tile_X5Y7_LUT4AB/FrameData[31]
+ Tile_X5Y7_LUT4AB/FrameData[3] Tile_X5Y7_LUT4AB/FrameData[4] Tile_X5Y7_LUT4AB/FrameData[5]
+ Tile_X5Y7_LUT4AB/FrameData[6] Tile_X5Y7_LUT4AB/FrameData[7] Tile_X5Y7_LUT4AB/FrameData[8]
+ Tile_X5Y7_LUT4AB/FrameData[9] Tile_X4Y7_RegFile/FrameStrobe[0] Tile_X4Y7_RegFile/FrameStrobe[10]
+ Tile_X4Y7_RegFile/FrameStrobe[11] Tile_X4Y7_RegFile/FrameStrobe[12] Tile_X4Y7_RegFile/FrameStrobe[13]
+ Tile_X4Y7_RegFile/FrameStrobe[14] Tile_X4Y7_RegFile/FrameStrobe[15] Tile_X4Y7_RegFile/FrameStrobe[16]
+ Tile_X4Y7_RegFile/FrameStrobe[17] Tile_X4Y7_RegFile/FrameStrobe[18] Tile_X4Y7_RegFile/FrameStrobe[19]
+ Tile_X4Y7_RegFile/FrameStrobe[1] Tile_X4Y7_RegFile/FrameStrobe[2] Tile_X4Y7_RegFile/FrameStrobe[3]
+ Tile_X4Y7_RegFile/FrameStrobe[4] Tile_X4Y7_RegFile/FrameStrobe[5] Tile_X4Y7_RegFile/FrameStrobe[6]
+ Tile_X4Y7_RegFile/FrameStrobe[7] Tile_X4Y7_RegFile/FrameStrobe[8] Tile_X4Y7_RegFile/FrameStrobe[9]
+ Tile_X4Y6_RegFile/FrameStrobe[0] Tile_X4Y6_RegFile/FrameStrobe[10] Tile_X4Y6_RegFile/FrameStrobe[11]
+ Tile_X4Y6_RegFile/FrameStrobe[12] Tile_X4Y6_RegFile/FrameStrobe[13] Tile_X4Y6_RegFile/FrameStrobe[14]
+ Tile_X4Y6_RegFile/FrameStrobe[15] Tile_X4Y6_RegFile/FrameStrobe[16] Tile_X4Y6_RegFile/FrameStrobe[17]
+ Tile_X4Y6_RegFile/FrameStrobe[18] Tile_X4Y6_RegFile/FrameStrobe[19] Tile_X4Y6_RegFile/FrameStrobe[1]
+ Tile_X4Y6_RegFile/FrameStrobe[2] Tile_X4Y6_RegFile/FrameStrobe[3] Tile_X4Y6_RegFile/FrameStrobe[4]
+ Tile_X4Y6_RegFile/FrameStrobe[5] Tile_X4Y6_RegFile/FrameStrobe[6] Tile_X4Y6_RegFile/FrameStrobe[7]
+ Tile_X4Y6_RegFile/FrameStrobe[8] Tile_X4Y6_RegFile/FrameStrobe[9] Tile_X4Y7_RegFile/N1BEG[0]
+ Tile_X4Y7_RegFile/N1BEG[1] Tile_X4Y7_RegFile/N1BEG[2] Tile_X4Y7_RegFile/N1BEG[3]
+ Tile_X4Y8_RegFile/N1BEG[0] Tile_X4Y8_RegFile/N1BEG[1] Tile_X4Y8_RegFile/N1BEG[2]
+ Tile_X4Y8_RegFile/N1BEG[3] Tile_X4Y7_RegFile/N2BEG[0] Tile_X4Y7_RegFile/N2BEG[1]
+ Tile_X4Y7_RegFile/N2BEG[2] Tile_X4Y7_RegFile/N2BEG[3] Tile_X4Y7_RegFile/N2BEG[4]
+ Tile_X4Y7_RegFile/N2BEG[5] Tile_X4Y7_RegFile/N2BEG[6] Tile_X4Y7_RegFile/N2BEG[7]
+ Tile_X4Y6_RegFile/N2END[0] Tile_X4Y6_RegFile/N2END[1] Tile_X4Y6_RegFile/N2END[2]
+ Tile_X4Y6_RegFile/N2END[3] Tile_X4Y6_RegFile/N2END[4] Tile_X4Y6_RegFile/N2END[5]
+ Tile_X4Y6_RegFile/N2END[6] Tile_X4Y6_RegFile/N2END[7] Tile_X4Y7_RegFile/N2END[0]
+ Tile_X4Y7_RegFile/N2END[1] Tile_X4Y7_RegFile/N2END[2] Tile_X4Y7_RegFile/N2END[3]
+ Tile_X4Y7_RegFile/N2END[4] Tile_X4Y7_RegFile/N2END[5] Tile_X4Y7_RegFile/N2END[6]
+ Tile_X4Y7_RegFile/N2END[7] Tile_X4Y8_RegFile/N2BEG[0] Tile_X4Y8_RegFile/N2BEG[1]
+ Tile_X4Y8_RegFile/N2BEG[2] Tile_X4Y8_RegFile/N2BEG[3] Tile_X4Y8_RegFile/N2BEG[4]
+ Tile_X4Y8_RegFile/N2BEG[5] Tile_X4Y8_RegFile/N2BEG[6] Tile_X4Y8_RegFile/N2BEG[7]
+ Tile_X4Y7_RegFile/N4BEG[0] Tile_X4Y7_RegFile/N4BEG[10] Tile_X4Y7_RegFile/N4BEG[11]
+ Tile_X4Y7_RegFile/N4BEG[12] Tile_X4Y7_RegFile/N4BEG[13] Tile_X4Y7_RegFile/N4BEG[14]
+ Tile_X4Y7_RegFile/N4BEG[15] Tile_X4Y7_RegFile/N4BEG[1] Tile_X4Y7_RegFile/N4BEG[2]
+ Tile_X4Y7_RegFile/N4BEG[3] Tile_X4Y7_RegFile/N4BEG[4] Tile_X4Y7_RegFile/N4BEG[5]
+ Tile_X4Y7_RegFile/N4BEG[6] Tile_X4Y7_RegFile/N4BEG[7] Tile_X4Y7_RegFile/N4BEG[8]
+ Tile_X4Y7_RegFile/N4BEG[9] Tile_X4Y8_RegFile/N4BEG[0] Tile_X4Y8_RegFile/N4BEG[10]
+ Tile_X4Y8_RegFile/N4BEG[11] Tile_X4Y8_RegFile/N4BEG[12] Tile_X4Y8_RegFile/N4BEG[13]
+ Tile_X4Y8_RegFile/N4BEG[14] Tile_X4Y8_RegFile/N4BEG[15] Tile_X4Y8_RegFile/N4BEG[1]
+ Tile_X4Y8_RegFile/N4BEG[2] Tile_X4Y8_RegFile/N4BEG[3] Tile_X4Y8_RegFile/N4BEG[4]
+ Tile_X4Y8_RegFile/N4BEG[5] Tile_X4Y8_RegFile/N4BEG[6] Tile_X4Y8_RegFile/N4BEG[7]
+ Tile_X4Y8_RegFile/N4BEG[8] Tile_X4Y8_RegFile/N4BEG[9] Tile_X4Y7_RegFile/NN4BEG[0]
+ Tile_X4Y7_RegFile/NN4BEG[10] Tile_X4Y7_RegFile/NN4BEG[11] Tile_X4Y7_RegFile/NN4BEG[12]
+ Tile_X4Y7_RegFile/NN4BEG[13] Tile_X4Y7_RegFile/NN4BEG[14] Tile_X4Y7_RegFile/NN4BEG[15]
+ Tile_X4Y7_RegFile/NN4BEG[1] Tile_X4Y7_RegFile/NN4BEG[2] Tile_X4Y7_RegFile/NN4BEG[3]
+ Tile_X4Y7_RegFile/NN4BEG[4] Tile_X4Y7_RegFile/NN4BEG[5] Tile_X4Y7_RegFile/NN4BEG[6]
+ Tile_X4Y7_RegFile/NN4BEG[7] Tile_X4Y7_RegFile/NN4BEG[8] Tile_X4Y7_RegFile/NN4BEG[9]
+ Tile_X4Y8_RegFile/NN4BEG[0] Tile_X4Y8_RegFile/NN4BEG[10] Tile_X4Y8_RegFile/NN4BEG[11]
+ Tile_X4Y8_RegFile/NN4BEG[12] Tile_X4Y8_RegFile/NN4BEG[13] Tile_X4Y8_RegFile/NN4BEG[14]
+ Tile_X4Y8_RegFile/NN4BEG[15] Tile_X4Y8_RegFile/NN4BEG[1] Tile_X4Y8_RegFile/NN4BEG[2]
+ Tile_X4Y8_RegFile/NN4BEG[3] Tile_X4Y8_RegFile/NN4BEG[4] Tile_X4Y8_RegFile/NN4BEG[5]
+ Tile_X4Y8_RegFile/NN4BEG[6] Tile_X4Y8_RegFile/NN4BEG[7] Tile_X4Y8_RegFile/NN4BEG[8]
+ Tile_X4Y8_RegFile/NN4BEG[9] Tile_X4Y8_RegFile/S1END[0] Tile_X4Y8_RegFile/S1END[1]
+ Tile_X4Y8_RegFile/S1END[2] Tile_X4Y8_RegFile/S1END[3] Tile_X4Y7_RegFile/S1END[0]
+ Tile_X4Y7_RegFile/S1END[1] Tile_X4Y7_RegFile/S1END[2] Tile_X4Y7_RegFile/S1END[3]
+ Tile_X4Y8_RegFile/S2MID[0] Tile_X4Y8_RegFile/S2MID[1] Tile_X4Y8_RegFile/S2MID[2]
+ Tile_X4Y8_RegFile/S2MID[3] Tile_X4Y8_RegFile/S2MID[4] Tile_X4Y8_RegFile/S2MID[5]
+ Tile_X4Y8_RegFile/S2MID[6] Tile_X4Y8_RegFile/S2MID[7] Tile_X4Y8_RegFile/S2END[0]
+ Tile_X4Y8_RegFile/S2END[1] Tile_X4Y8_RegFile/S2END[2] Tile_X4Y8_RegFile/S2END[3]
+ Tile_X4Y8_RegFile/S2END[4] Tile_X4Y8_RegFile/S2END[5] Tile_X4Y8_RegFile/S2END[6]
+ Tile_X4Y8_RegFile/S2END[7] Tile_X4Y7_RegFile/S2END[0] Tile_X4Y7_RegFile/S2END[1]
+ Tile_X4Y7_RegFile/S2END[2] Tile_X4Y7_RegFile/S2END[3] Tile_X4Y7_RegFile/S2END[4]
+ Tile_X4Y7_RegFile/S2END[5] Tile_X4Y7_RegFile/S2END[6] Tile_X4Y7_RegFile/S2END[7]
+ Tile_X4Y7_RegFile/S2MID[0] Tile_X4Y7_RegFile/S2MID[1] Tile_X4Y7_RegFile/S2MID[2]
+ Tile_X4Y7_RegFile/S2MID[3] Tile_X4Y7_RegFile/S2MID[4] Tile_X4Y7_RegFile/S2MID[5]
+ Tile_X4Y7_RegFile/S2MID[6] Tile_X4Y7_RegFile/S2MID[7] Tile_X4Y8_RegFile/S4END[0]
+ Tile_X4Y8_RegFile/S4END[10] Tile_X4Y8_RegFile/S4END[11] Tile_X4Y8_RegFile/S4END[12]
+ Tile_X4Y8_RegFile/S4END[13] Tile_X4Y8_RegFile/S4END[14] Tile_X4Y8_RegFile/S4END[15]
+ Tile_X4Y8_RegFile/S4END[1] Tile_X4Y8_RegFile/S4END[2] Tile_X4Y8_RegFile/S4END[3]
+ Tile_X4Y8_RegFile/S4END[4] Tile_X4Y8_RegFile/S4END[5] Tile_X4Y8_RegFile/S4END[6]
+ Tile_X4Y8_RegFile/S4END[7] Tile_X4Y8_RegFile/S4END[8] Tile_X4Y8_RegFile/S4END[9]
+ Tile_X4Y7_RegFile/S4END[0] Tile_X4Y7_RegFile/S4END[10] Tile_X4Y7_RegFile/S4END[11]
+ Tile_X4Y7_RegFile/S4END[12] Tile_X4Y7_RegFile/S4END[13] Tile_X4Y7_RegFile/S4END[14]
+ Tile_X4Y7_RegFile/S4END[15] Tile_X4Y7_RegFile/S4END[1] Tile_X4Y7_RegFile/S4END[2]
+ Tile_X4Y7_RegFile/S4END[3] Tile_X4Y7_RegFile/S4END[4] Tile_X4Y7_RegFile/S4END[5]
+ Tile_X4Y7_RegFile/S4END[6] Tile_X4Y7_RegFile/S4END[7] Tile_X4Y7_RegFile/S4END[8]
+ Tile_X4Y7_RegFile/S4END[9] Tile_X4Y8_RegFile/SS4END[0] Tile_X4Y8_RegFile/SS4END[10]
+ Tile_X4Y8_RegFile/SS4END[11] Tile_X4Y8_RegFile/SS4END[12] Tile_X4Y8_RegFile/SS4END[13]
+ Tile_X4Y8_RegFile/SS4END[14] Tile_X4Y8_RegFile/SS4END[15] Tile_X4Y8_RegFile/SS4END[1]
+ Tile_X4Y8_RegFile/SS4END[2] Tile_X4Y8_RegFile/SS4END[3] Tile_X4Y8_RegFile/SS4END[4]
+ Tile_X4Y8_RegFile/SS4END[5] Tile_X4Y8_RegFile/SS4END[6] Tile_X4Y8_RegFile/SS4END[7]
+ Tile_X4Y8_RegFile/SS4END[8] Tile_X4Y8_RegFile/SS4END[9] Tile_X4Y7_RegFile/SS4END[0]
+ Tile_X4Y7_RegFile/SS4END[10] Tile_X4Y7_RegFile/SS4END[11] Tile_X4Y7_RegFile/SS4END[12]
+ Tile_X4Y7_RegFile/SS4END[13] Tile_X4Y7_RegFile/SS4END[14] Tile_X4Y7_RegFile/SS4END[15]
+ Tile_X4Y7_RegFile/SS4END[1] Tile_X4Y7_RegFile/SS4END[2] Tile_X4Y7_RegFile/SS4END[3]
+ Tile_X4Y7_RegFile/SS4END[4] Tile_X4Y7_RegFile/SS4END[5] Tile_X4Y7_RegFile/SS4END[6]
+ Tile_X4Y7_RegFile/SS4END[7] Tile_X4Y7_RegFile/SS4END[8] Tile_X4Y7_RegFile/SS4END[9]
+ Tile_X4Y7_RegFile/UserCLK Tile_X4Y6_RegFile/UserCLK VGND VPWR Tile_X3Y7_LUT4AB/W1END[0]
+ Tile_X3Y7_LUT4AB/W1END[1] Tile_X3Y7_LUT4AB/W1END[2] Tile_X3Y7_LUT4AB/W1END[3] Tile_X5Y7_LUT4AB/W1BEG[0]
+ Tile_X5Y7_LUT4AB/W1BEG[1] Tile_X5Y7_LUT4AB/W1BEG[2] Tile_X5Y7_LUT4AB/W1BEG[3] Tile_X3Y7_LUT4AB/W2MID[0]
+ Tile_X3Y7_LUT4AB/W2MID[1] Tile_X3Y7_LUT4AB/W2MID[2] Tile_X3Y7_LUT4AB/W2MID[3] Tile_X3Y7_LUT4AB/W2MID[4]
+ Tile_X3Y7_LUT4AB/W2MID[5] Tile_X3Y7_LUT4AB/W2MID[6] Tile_X3Y7_LUT4AB/W2MID[7] Tile_X3Y7_LUT4AB/W2END[0]
+ Tile_X3Y7_LUT4AB/W2END[1] Tile_X3Y7_LUT4AB/W2END[2] Tile_X3Y7_LUT4AB/W2END[3] Tile_X3Y7_LUT4AB/W2END[4]
+ Tile_X3Y7_LUT4AB/W2END[5] Tile_X3Y7_LUT4AB/W2END[6] Tile_X3Y7_LUT4AB/W2END[7] Tile_X5Y7_LUT4AB/W2BEGb[0]
+ Tile_X5Y7_LUT4AB/W2BEGb[1] Tile_X5Y7_LUT4AB/W2BEGb[2] Tile_X5Y7_LUT4AB/W2BEGb[3]
+ Tile_X5Y7_LUT4AB/W2BEGb[4] Tile_X5Y7_LUT4AB/W2BEGb[5] Tile_X5Y7_LUT4AB/W2BEGb[6]
+ Tile_X5Y7_LUT4AB/W2BEGb[7] Tile_X5Y7_LUT4AB/W2BEG[0] Tile_X5Y7_LUT4AB/W2BEG[1] Tile_X5Y7_LUT4AB/W2BEG[2]
+ Tile_X5Y7_LUT4AB/W2BEG[3] Tile_X5Y7_LUT4AB/W2BEG[4] Tile_X5Y7_LUT4AB/W2BEG[5] Tile_X5Y7_LUT4AB/W2BEG[6]
+ Tile_X5Y7_LUT4AB/W2BEG[7] Tile_X3Y7_LUT4AB/W6END[0] Tile_X3Y7_LUT4AB/W6END[10] Tile_X3Y7_LUT4AB/W6END[11]
+ Tile_X3Y7_LUT4AB/W6END[1] Tile_X3Y7_LUT4AB/W6END[2] Tile_X3Y7_LUT4AB/W6END[3] Tile_X3Y7_LUT4AB/W6END[4]
+ Tile_X3Y7_LUT4AB/W6END[5] Tile_X3Y7_LUT4AB/W6END[6] Tile_X3Y7_LUT4AB/W6END[7] Tile_X3Y7_LUT4AB/W6END[8]
+ Tile_X3Y7_LUT4AB/W6END[9] Tile_X5Y7_LUT4AB/W6BEG[0] Tile_X5Y7_LUT4AB/W6BEG[10] Tile_X5Y7_LUT4AB/W6BEG[11]
+ Tile_X5Y7_LUT4AB/W6BEG[1] Tile_X5Y7_LUT4AB/W6BEG[2] Tile_X5Y7_LUT4AB/W6BEG[3] Tile_X5Y7_LUT4AB/W6BEG[4]
+ Tile_X5Y7_LUT4AB/W6BEG[5] Tile_X5Y7_LUT4AB/W6BEG[6] Tile_X5Y7_LUT4AB/W6BEG[7] Tile_X5Y7_LUT4AB/W6BEG[8]
+ Tile_X5Y7_LUT4AB/W6BEG[9] Tile_X3Y7_LUT4AB/WW4END[0] Tile_X3Y7_LUT4AB/WW4END[10]
+ Tile_X3Y7_LUT4AB/WW4END[11] Tile_X3Y7_LUT4AB/WW4END[12] Tile_X3Y7_LUT4AB/WW4END[13]
+ Tile_X3Y7_LUT4AB/WW4END[14] Tile_X3Y7_LUT4AB/WW4END[15] Tile_X3Y7_LUT4AB/WW4END[1]
+ Tile_X3Y7_LUT4AB/WW4END[2] Tile_X3Y7_LUT4AB/WW4END[3] Tile_X3Y7_LUT4AB/WW4END[4]
+ Tile_X3Y7_LUT4AB/WW4END[5] Tile_X3Y7_LUT4AB/WW4END[6] Tile_X3Y7_LUT4AB/WW4END[7]
+ Tile_X3Y7_LUT4AB/WW4END[8] Tile_X3Y7_LUT4AB/WW4END[9] Tile_X5Y7_LUT4AB/WW4BEG[0]
+ Tile_X5Y7_LUT4AB/WW4BEG[10] Tile_X5Y7_LUT4AB/WW4BEG[11] Tile_X5Y7_LUT4AB/WW4BEG[12]
+ Tile_X5Y7_LUT4AB/WW4BEG[13] Tile_X5Y7_LUT4AB/WW4BEG[14] Tile_X5Y7_LUT4AB/WW4BEG[15]
+ Tile_X5Y7_LUT4AB/WW4BEG[1] Tile_X5Y7_LUT4AB/WW4BEG[2] Tile_X5Y7_LUT4AB/WW4BEG[3]
+ Tile_X5Y7_LUT4AB/WW4BEG[4] Tile_X5Y7_LUT4AB/WW4BEG[5] Tile_X5Y7_LUT4AB/WW4BEG[6]
+ Tile_X5Y7_LUT4AB/WW4BEG[7] Tile_X5Y7_LUT4AB/WW4BEG[8] Tile_X5Y7_LUT4AB/WW4BEG[9]
+ RegFile
XTile_X1Y13_LUT4AB Tile_X1Y14_LUT4AB/Co Tile_X1Y13_LUT4AB/Co Tile_X2Y13_LUT4AB/E1END[0]
+ Tile_X2Y13_LUT4AB/E1END[1] Tile_X2Y13_LUT4AB/E1END[2] Tile_X2Y13_LUT4AB/E1END[3]
+ Tile_X0Y13_W_IO/E1BEG[0] Tile_X0Y13_W_IO/E1BEG[1] Tile_X0Y13_W_IO/E1BEG[2] Tile_X0Y13_W_IO/E1BEG[3]
+ Tile_X2Y13_LUT4AB/E2MID[0] Tile_X2Y13_LUT4AB/E2MID[1] Tile_X2Y13_LUT4AB/E2MID[2]
+ Tile_X2Y13_LUT4AB/E2MID[3] Tile_X2Y13_LUT4AB/E2MID[4] Tile_X2Y13_LUT4AB/E2MID[5]
+ Tile_X2Y13_LUT4AB/E2MID[6] Tile_X2Y13_LUT4AB/E2MID[7] Tile_X2Y13_LUT4AB/E2END[0]
+ Tile_X2Y13_LUT4AB/E2END[1] Tile_X2Y13_LUT4AB/E2END[2] Tile_X2Y13_LUT4AB/E2END[3]
+ Tile_X2Y13_LUT4AB/E2END[4] Tile_X2Y13_LUT4AB/E2END[5] Tile_X2Y13_LUT4AB/E2END[6]
+ Tile_X2Y13_LUT4AB/E2END[7] Tile_X0Y13_W_IO/E2BEGb[0] Tile_X0Y13_W_IO/E2BEGb[1] Tile_X0Y13_W_IO/E2BEGb[2]
+ Tile_X0Y13_W_IO/E2BEGb[3] Tile_X0Y13_W_IO/E2BEGb[4] Tile_X0Y13_W_IO/E2BEGb[5] Tile_X0Y13_W_IO/E2BEGb[6]
+ Tile_X0Y13_W_IO/E2BEGb[7] Tile_X0Y13_W_IO/E2BEG[0] Tile_X0Y13_W_IO/E2BEG[1] Tile_X0Y13_W_IO/E2BEG[2]
+ Tile_X0Y13_W_IO/E2BEG[3] Tile_X0Y13_W_IO/E2BEG[4] Tile_X0Y13_W_IO/E2BEG[5] Tile_X0Y13_W_IO/E2BEG[6]
+ Tile_X0Y13_W_IO/E2BEG[7] Tile_X2Y13_LUT4AB/E6END[0] Tile_X2Y13_LUT4AB/E6END[10]
+ Tile_X2Y13_LUT4AB/E6END[11] Tile_X2Y13_LUT4AB/E6END[1] Tile_X2Y13_LUT4AB/E6END[2]
+ Tile_X2Y13_LUT4AB/E6END[3] Tile_X2Y13_LUT4AB/E6END[4] Tile_X2Y13_LUT4AB/E6END[5]
+ Tile_X2Y13_LUT4AB/E6END[6] Tile_X2Y13_LUT4AB/E6END[7] Tile_X2Y13_LUT4AB/E6END[8]
+ Tile_X2Y13_LUT4AB/E6END[9] Tile_X0Y13_W_IO/E6BEG[0] Tile_X0Y13_W_IO/E6BEG[10] Tile_X0Y13_W_IO/E6BEG[11]
+ Tile_X0Y13_W_IO/E6BEG[1] Tile_X0Y13_W_IO/E6BEG[2] Tile_X0Y13_W_IO/E6BEG[3] Tile_X0Y13_W_IO/E6BEG[4]
+ Tile_X0Y13_W_IO/E6BEG[5] Tile_X0Y13_W_IO/E6BEG[6] Tile_X0Y13_W_IO/E6BEG[7] Tile_X0Y13_W_IO/E6BEG[8]
+ Tile_X0Y13_W_IO/E6BEG[9] Tile_X2Y13_LUT4AB/EE4END[0] Tile_X2Y13_LUT4AB/EE4END[10]
+ Tile_X2Y13_LUT4AB/EE4END[11] Tile_X2Y13_LUT4AB/EE4END[12] Tile_X2Y13_LUT4AB/EE4END[13]
+ Tile_X2Y13_LUT4AB/EE4END[14] Tile_X2Y13_LUT4AB/EE4END[15] Tile_X2Y13_LUT4AB/EE4END[1]
+ Tile_X2Y13_LUT4AB/EE4END[2] Tile_X2Y13_LUT4AB/EE4END[3] Tile_X2Y13_LUT4AB/EE4END[4]
+ Tile_X2Y13_LUT4AB/EE4END[5] Tile_X2Y13_LUT4AB/EE4END[6] Tile_X2Y13_LUT4AB/EE4END[7]
+ Tile_X2Y13_LUT4AB/EE4END[8] Tile_X2Y13_LUT4AB/EE4END[9] Tile_X0Y13_W_IO/EE4BEG[0]
+ Tile_X0Y13_W_IO/EE4BEG[10] Tile_X0Y13_W_IO/EE4BEG[11] Tile_X0Y13_W_IO/EE4BEG[12]
+ Tile_X0Y13_W_IO/EE4BEG[13] Tile_X0Y13_W_IO/EE4BEG[14] Tile_X0Y13_W_IO/EE4BEG[15]
+ Tile_X0Y13_W_IO/EE4BEG[1] Tile_X0Y13_W_IO/EE4BEG[2] Tile_X0Y13_W_IO/EE4BEG[3] Tile_X0Y13_W_IO/EE4BEG[4]
+ Tile_X0Y13_W_IO/EE4BEG[5] Tile_X0Y13_W_IO/EE4BEG[6] Tile_X0Y13_W_IO/EE4BEG[7] Tile_X0Y13_W_IO/EE4BEG[8]
+ Tile_X0Y13_W_IO/EE4BEG[9] Tile_X1Y13_LUT4AB/FrameData[0] Tile_X1Y13_LUT4AB/FrameData[10]
+ Tile_X1Y13_LUT4AB/FrameData[11] Tile_X1Y13_LUT4AB/FrameData[12] Tile_X1Y13_LUT4AB/FrameData[13]
+ Tile_X1Y13_LUT4AB/FrameData[14] Tile_X1Y13_LUT4AB/FrameData[15] Tile_X1Y13_LUT4AB/FrameData[16]
+ Tile_X1Y13_LUT4AB/FrameData[17] Tile_X1Y13_LUT4AB/FrameData[18] Tile_X1Y13_LUT4AB/FrameData[19]
+ Tile_X1Y13_LUT4AB/FrameData[1] Tile_X1Y13_LUT4AB/FrameData[20] Tile_X1Y13_LUT4AB/FrameData[21]
+ Tile_X1Y13_LUT4AB/FrameData[22] Tile_X1Y13_LUT4AB/FrameData[23] Tile_X1Y13_LUT4AB/FrameData[24]
+ Tile_X1Y13_LUT4AB/FrameData[25] Tile_X1Y13_LUT4AB/FrameData[26] Tile_X1Y13_LUT4AB/FrameData[27]
+ Tile_X1Y13_LUT4AB/FrameData[28] Tile_X1Y13_LUT4AB/FrameData[29] Tile_X1Y13_LUT4AB/FrameData[2]
+ Tile_X1Y13_LUT4AB/FrameData[30] Tile_X1Y13_LUT4AB/FrameData[31] Tile_X1Y13_LUT4AB/FrameData[3]
+ Tile_X1Y13_LUT4AB/FrameData[4] Tile_X1Y13_LUT4AB/FrameData[5] Tile_X1Y13_LUT4AB/FrameData[6]
+ Tile_X1Y13_LUT4AB/FrameData[7] Tile_X1Y13_LUT4AB/FrameData[8] Tile_X1Y13_LUT4AB/FrameData[9]
+ Tile_X2Y13_LUT4AB/FrameData[0] Tile_X2Y13_LUT4AB/FrameData[10] Tile_X2Y13_LUT4AB/FrameData[11]
+ Tile_X2Y13_LUT4AB/FrameData[12] Tile_X2Y13_LUT4AB/FrameData[13] Tile_X2Y13_LUT4AB/FrameData[14]
+ Tile_X2Y13_LUT4AB/FrameData[15] Tile_X2Y13_LUT4AB/FrameData[16] Tile_X2Y13_LUT4AB/FrameData[17]
+ Tile_X2Y13_LUT4AB/FrameData[18] Tile_X2Y13_LUT4AB/FrameData[19] Tile_X2Y13_LUT4AB/FrameData[1]
+ Tile_X2Y13_LUT4AB/FrameData[20] Tile_X2Y13_LUT4AB/FrameData[21] Tile_X2Y13_LUT4AB/FrameData[22]
+ Tile_X2Y13_LUT4AB/FrameData[23] Tile_X2Y13_LUT4AB/FrameData[24] Tile_X2Y13_LUT4AB/FrameData[25]
+ Tile_X2Y13_LUT4AB/FrameData[26] Tile_X2Y13_LUT4AB/FrameData[27] Tile_X2Y13_LUT4AB/FrameData[28]
+ Tile_X2Y13_LUT4AB/FrameData[29] Tile_X2Y13_LUT4AB/FrameData[2] Tile_X2Y13_LUT4AB/FrameData[30]
+ Tile_X2Y13_LUT4AB/FrameData[31] Tile_X2Y13_LUT4AB/FrameData[3] Tile_X2Y13_LUT4AB/FrameData[4]
+ Tile_X2Y13_LUT4AB/FrameData[5] Tile_X2Y13_LUT4AB/FrameData[6] Tile_X2Y13_LUT4AB/FrameData[7]
+ Tile_X2Y13_LUT4AB/FrameData[8] Tile_X2Y13_LUT4AB/FrameData[9] Tile_X1Y13_LUT4AB/FrameStrobe[0]
+ Tile_X1Y13_LUT4AB/FrameStrobe[10] Tile_X1Y13_LUT4AB/FrameStrobe[11] Tile_X1Y13_LUT4AB/FrameStrobe[12]
+ Tile_X1Y13_LUT4AB/FrameStrobe[13] Tile_X1Y13_LUT4AB/FrameStrobe[14] Tile_X1Y13_LUT4AB/FrameStrobe[15]
+ Tile_X1Y13_LUT4AB/FrameStrobe[16] Tile_X1Y13_LUT4AB/FrameStrobe[17] Tile_X1Y13_LUT4AB/FrameStrobe[18]
+ Tile_X1Y13_LUT4AB/FrameStrobe[19] Tile_X1Y13_LUT4AB/FrameStrobe[1] Tile_X1Y13_LUT4AB/FrameStrobe[2]
+ Tile_X1Y13_LUT4AB/FrameStrobe[3] Tile_X1Y13_LUT4AB/FrameStrobe[4] Tile_X1Y13_LUT4AB/FrameStrobe[5]
+ Tile_X1Y13_LUT4AB/FrameStrobe[6] Tile_X1Y13_LUT4AB/FrameStrobe[7] Tile_X1Y13_LUT4AB/FrameStrobe[8]
+ Tile_X1Y13_LUT4AB/FrameStrobe[9] Tile_X1Y12_LUT4AB/FrameStrobe[0] Tile_X1Y12_LUT4AB/FrameStrobe[10]
+ Tile_X1Y12_LUT4AB/FrameStrobe[11] Tile_X1Y12_LUT4AB/FrameStrobe[12] Tile_X1Y12_LUT4AB/FrameStrobe[13]
+ Tile_X1Y12_LUT4AB/FrameStrobe[14] Tile_X1Y12_LUT4AB/FrameStrobe[15] Tile_X1Y12_LUT4AB/FrameStrobe[16]
+ Tile_X1Y12_LUT4AB/FrameStrobe[17] Tile_X1Y12_LUT4AB/FrameStrobe[18] Tile_X1Y12_LUT4AB/FrameStrobe[19]
+ Tile_X1Y12_LUT4AB/FrameStrobe[1] Tile_X1Y12_LUT4AB/FrameStrobe[2] Tile_X1Y12_LUT4AB/FrameStrobe[3]
+ Tile_X1Y12_LUT4AB/FrameStrobe[4] Tile_X1Y12_LUT4AB/FrameStrobe[5] Tile_X1Y12_LUT4AB/FrameStrobe[6]
+ Tile_X1Y12_LUT4AB/FrameStrobe[7] Tile_X1Y12_LUT4AB/FrameStrobe[8] Tile_X1Y12_LUT4AB/FrameStrobe[9]
+ Tile_X1Y13_LUT4AB/N1BEG[0] Tile_X1Y13_LUT4AB/N1BEG[1] Tile_X1Y13_LUT4AB/N1BEG[2]
+ Tile_X1Y13_LUT4AB/N1BEG[3] Tile_X1Y14_LUT4AB/N1BEG[0] Tile_X1Y14_LUT4AB/N1BEG[1]
+ Tile_X1Y14_LUT4AB/N1BEG[2] Tile_X1Y14_LUT4AB/N1BEG[3] Tile_X1Y13_LUT4AB/N2BEG[0]
+ Tile_X1Y13_LUT4AB/N2BEG[1] Tile_X1Y13_LUT4AB/N2BEG[2] Tile_X1Y13_LUT4AB/N2BEG[3]
+ Tile_X1Y13_LUT4AB/N2BEG[4] Tile_X1Y13_LUT4AB/N2BEG[5] Tile_X1Y13_LUT4AB/N2BEG[6]
+ Tile_X1Y13_LUT4AB/N2BEG[7] Tile_X1Y12_LUT4AB/N2END[0] Tile_X1Y12_LUT4AB/N2END[1]
+ Tile_X1Y12_LUT4AB/N2END[2] Tile_X1Y12_LUT4AB/N2END[3] Tile_X1Y12_LUT4AB/N2END[4]
+ Tile_X1Y12_LUT4AB/N2END[5] Tile_X1Y12_LUT4AB/N2END[6] Tile_X1Y12_LUT4AB/N2END[7]
+ Tile_X1Y13_LUT4AB/N2END[0] Tile_X1Y13_LUT4AB/N2END[1] Tile_X1Y13_LUT4AB/N2END[2]
+ Tile_X1Y13_LUT4AB/N2END[3] Tile_X1Y13_LUT4AB/N2END[4] Tile_X1Y13_LUT4AB/N2END[5]
+ Tile_X1Y13_LUT4AB/N2END[6] Tile_X1Y13_LUT4AB/N2END[7] Tile_X1Y14_LUT4AB/N2BEG[0]
+ Tile_X1Y14_LUT4AB/N2BEG[1] Tile_X1Y14_LUT4AB/N2BEG[2] Tile_X1Y14_LUT4AB/N2BEG[3]
+ Tile_X1Y14_LUT4AB/N2BEG[4] Tile_X1Y14_LUT4AB/N2BEG[5] Tile_X1Y14_LUT4AB/N2BEG[6]
+ Tile_X1Y14_LUT4AB/N2BEG[7] Tile_X1Y13_LUT4AB/N4BEG[0] Tile_X1Y13_LUT4AB/N4BEG[10]
+ Tile_X1Y13_LUT4AB/N4BEG[11] Tile_X1Y13_LUT4AB/N4BEG[12] Tile_X1Y13_LUT4AB/N4BEG[13]
+ Tile_X1Y13_LUT4AB/N4BEG[14] Tile_X1Y13_LUT4AB/N4BEG[15] Tile_X1Y13_LUT4AB/N4BEG[1]
+ Tile_X1Y13_LUT4AB/N4BEG[2] Tile_X1Y13_LUT4AB/N4BEG[3] Tile_X1Y13_LUT4AB/N4BEG[4]
+ Tile_X1Y13_LUT4AB/N4BEG[5] Tile_X1Y13_LUT4AB/N4BEG[6] Tile_X1Y13_LUT4AB/N4BEG[7]
+ Tile_X1Y13_LUT4AB/N4BEG[8] Tile_X1Y13_LUT4AB/N4BEG[9] Tile_X1Y14_LUT4AB/N4BEG[0]
+ Tile_X1Y14_LUT4AB/N4BEG[10] Tile_X1Y14_LUT4AB/N4BEG[11] Tile_X1Y14_LUT4AB/N4BEG[12]
+ Tile_X1Y14_LUT4AB/N4BEG[13] Tile_X1Y14_LUT4AB/N4BEG[14] Tile_X1Y14_LUT4AB/N4BEG[15]
+ Tile_X1Y14_LUT4AB/N4BEG[1] Tile_X1Y14_LUT4AB/N4BEG[2] Tile_X1Y14_LUT4AB/N4BEG[3]
+ Tile_X1Y14_LUT4AB/N4BEG[4] Tile_X1Y14_LUT4AB/N4BEG[5] Tile_X1Y14_LUT4AB/N4BEG[6]
+ Tile_X1Y14_LUT4AB/N4BEG[7] Tile_X1Y14_LUT4AB/N4BEG[8] Tile_X1Y14_LUT4AB/N4BEG[9]
+ Tile_X1Y13_LUT4AB/NN4BEG[0] Tile_X1Y13_LUT4AB/NN4BEG[10] Tile_X1Y13_LUT4AB/NN4BEG[11]
+ Tile_X1Y13_LUT4AB/NN4BEG[12] Tile_X1Y13_LUT4AB/NN4BEG[13] Tile_X1Y13_LUT4AB/NN4BEG[14]
+ Tile_X1Y13_LUT4AB/NN4BEG[15] Tile_X1Y13_LUT4AB/NN4BEG[1] Tile_X1Y13_LUT4AB/NN4BEG[2]
+ Tile_X1Y13_LUT4AB/NN4BEG[3] Tile_X1Y13_LUT4AB/NN4BEG[4] Tile_X1Y13_LUT4AB/NN4BEG[5]
+ Tile_X1Y13_LUT4AB/NN4BEG[6] Tile_X1Y13_LUT4AB/NN4BEG[7] Tile_X1Y13_LUT4AB/NN4BEG[8]
+ Tile_X1Y13_LUT4AB/NN4BEG[9] Tile_X1Y14_LUT4AB/NN4BEG[0] Tile_X1Y14_LUT4AB/NN4BEG[10]
+ Tile_X1Y14_LUT4AB/NN4BEG[11] Tile_X1Y14_LUT4AB/NN4BEG[12] Tile_X1Y14_LUT4AB/NN4BEG[13]
+ Tile_X1Y14_LUT4AB/NN4BEG[14] Tile_X1Y14_LUT4AB/NN4BEG[15] Tile_X1Y14_LUT4AB/NN4BEG[1]
+ Tile_X1Y14_LUT4AB/NN4BEG[2] Tile_X1Y14_LUT4AB/NN4BEG[3] Tile_X1Y14_LUT4AB/NN4BEG[4]
+ Tile_X1Y14_LUT4AB/NN4BEG[5] Tile_X1Y14_LUT4AB/NN4BEG[6] Tile_X1Y14_LUT4AB/NN4BEG[7]
+ Tile_X1Y14_LUT4AB/NN4BEG[8] Tile_X1Y14_LUT4AB/NN4BEG[9] Tile_X1Y14_LUT4AB/S1END[0]
+ Tile_X1Y14_LUT4AB/S1END[1] Tile_X1Y14_LUT4AB/S1END[2] Tile_X1Y14_LUT4AB/S1END[3]
+ Tile_X1Y13_LUT4AB/S1END[0] Tile_X1Y13_LUT4AB/S1END[1] Tile_X1Y13_LUT4AB/S1END[2]
+ Tile_X1Y13_LUT4AB/S1END[3] Tile_X1Y14_LUT4AB/S2MID[0] Tile_X1Y14_LUT4AB/S2MID[1]
+ Tile_X1Y14_LUT4AB/S2MID[2] Tile_X1Y14_LUT4AB/S2MID[3] Tile_X1Y14_LUT4AB/S2MID[4]
+ Tile_X1Y14_LUT4AB/S2MID[5] Tile_X1Y14_LUT4AB/S2MID[6] Tile_X1Y14_LUT4AB/S2MID[7]
+ Tile_X1Y14_LUT4AB/S2END[0] Tile_X1Y14_LUT4AB/S2END[1] Tile_X1Y14_LUT4AB/S2END[2]
+ Tile_X1Y14_LUT4AB/S2END[3] Tile_X1Y14_LUT4AB/S2END[4] Tile_X1Y14_LUT4AB/S2END[5]
+ Tile_X1Y14_LUT4AB/S2END[6] Tile_X1Y14_LUT4AB/S2END[7] Tile_X1Y13_LUT4AB/S2END[0]
+ Tile_X1Y13_LUT4AB/S2END[1] Tile_X1Y13_LUT4AB/S2END[2] Tile_X1Y13_LUT4AB/S2END[3]
+ Tile_X1Y13_LUT4AB/S2END[4] Tile_X1Y13_LUT4AB/S2END[5] Tile_X1Y13_LUT4AB/S2END[6]
+ Tile_X1Y13_LUT4AB/S2END[7] Tile_X1Y13_LUT4AB/S2MID[0] Tile_X1Y13_LUT4AB/S2MID[1]
+ Tile_X1Y13_LUT4AB/S2MID[2] Tile_X1Y13_LUT4AB/S2MID[3] Tile_X1Y13_LUT4AB/S2MID[4]
+ Tile_X1Y13_LUT4AB/S2MID[5] Tile_X1Y13_LUT4AB/S2MID[6] Tile_X1Y13_LUT4AB/S2MID[7]
+ Tile_X1Y14_LUT4AB/S4END[0] Tile_X1Y14_LUT4AB/S4END[10] Tile_X1Y14_LUT4AB/S4END[11]
+ Tile_X1Y14_LUT4AB/S4END[12] Tile_X1Y14_LUT4AB/S4END[13] Tile_X1Y14_LUT4AB/S4END[14]
+ Tile_X1Y14_LUT4AB/S4END[15] Tile_X1Y14_LUT4AB/S4END[1] Tile_X1Y14_LUT4AB/S4END[2]
+ Tile_X1Y14_LUT4AB/S4END[3] Tile_X1Y14_LUT4AB/S4END[4] Tile_X1Y14_LUT4AB/S4END[5]
+ Tile_X1Y14_LUT4AB/S4END[6] Tile_X1Y14_LUT4AB/S4END[7] Tile_X1Y14_LUT4AB/S4END[8]
+ Tile_X1Y14_LUT4AB/S4END[9] Tile_X1Y13_LUT4AB/S4END[0] Tile_X1Y13_LUT4AB/S4END[10]
+ Tile_X1Y13_LUT4AB/S4END[11] Tile_X1Y13_LUT4AB/S4END[12] Tile_X1Y13_LUT4AB/S4END[13]
+ Tile_X1Y13_LUT4AB/S4END[14] Tile_X1Y13_LUT4AB/S4END[15] Tile_X1Y13_LUT4AB/S4END[1]
+ Tile_X1Y13_LUT4AB/S4END[2] Tile_X1Y13_LUT4AB/S4END[3] Tile_X1Y13_LUT4AB/S4END[4]
+ Tile_X1Y13_LUT4AB/S4END[5] Tile_X1Y13_LUT4AB/S4END[6] Tile_X1Y13_LUT4AB/S4END[7]
+ Tile_X1Y13_LUT4AB/S4END[8] Tile_X1Y13_LUT4AB/S4END[9] Tile_X1Y14_LUT4AB/SS4END[0]
+ Tile_X1Y14_LUT4AB/SS4END[10] Tile_X1Y14_LUT4AB/SS4END[11] Tile_X1Y14_LUT4AB/SS4END[12]
+ Tile_X1Y14_LUT4AB/SS4END[13] Tile_X1Y14_LUT4AB/SS4END[14] Tile_X1Y14_LUT4AB/SS4END[15]
+ Tile_X1Y14_LUT4AB/SS4END[1] Tile_X1Y14_LUT4AB/SS4END[2] Tile_X1Y14_LUT4AB/SS4END[3]
+ Tile_X1Y14_LUT4AB/SS4END[4] Tile_X1Y14_LUT4AB/SS4END[5] Tile_X1Y14_LUT4AB/SS4END[6]
+ Tile_X1Y14_LUT4AB/SS4END[7] Tile_X1Y14_LUT4AB/SS4END[8] Tile_X1Y14_LUT4AB/SS4END[9]
+ Tile_X1Y13_LUT4AB/SS4END[0] Tile_X1Y13_LUT4AB/SS4END[10] Tile_X1Y13_LUT4AB/SS4END[11]
+ Tile_X1Y13_LUT4AB/SS4END[12] Tile_X1Y13_LUT4AB/SS4END[13] Tile_X1Y13_LUT4AB/SS4END[14]
+ Tile_X1Y13_LUT4AB/SS4END[15] Tile_X1Y13_LUT4AB/SS4END[1] Tile_X1Y13_LUT4AB/SS4END[2]
+ Tile_X1Y13_LUT4AB/SS4END[3] Tile_X1Y13_LUT4AB/SS4END[4] Tile_X1Y13_LUT4AB/SS4END[5]
+ Tile_X1Y13_LUT4AB/SS4END[6] Tile_X1Y13_LUT4AB/SS4END[7] Tile_X1Y13_LUT4AB/SS4END[8]
+ Tile_X1Y13_LUT4AB/SS4END[9] Tile_X1Y13_LUT4AB/UserCLK Tile_X1Y12_LUT4AB/UserCLK
+ VGND VPWR Tile_X0Y13_W_IO/W1END[0] Tile_X0Y13_W_IO/W1END[1] Tile_X0Y13_W_IO/W1END[2]
+ Tile_X0Y13_W_IO/W1END[3] Tile_X2Y13_LUT4AB/W1BEG[0] Tile_X2Y13_LUT4AB/W1BEG[1] Tile_X2Y13_LUT4AB/W1BEG[2]
+ Tile_X2Y13_LUT4AB/W1BEG[3] Tile_X0Y13_W_IO/W2MID[0] Tile_X0Y13_W_IO/W2MID[1] Tile_X0Y13_W_IO/W2MID[2]
+ Tile_X0Y13_W_IO/W2MID[3] Tile_X0Y13_W_IO/W2MID[4] Tile_X0Y13_W_IO/W2MID[5] Tile_X0Y13_W_IO/W2MID[6]
+ Tile_X0Y13_W_IO/W2MID[7] Tile_X0Y13_W_IO/W2END[0] Tile_X0Y13_W_IO/W2END[1] Tile_X0Y13_W_IO/W2END[2]
+ Tile_X0Y13_W_IO/W2END[3] Tile_X0Y13_W_IO/W2END[4] Tile_X0Y13_W_IO/W2END[5] Tile_X0Y13_W_IO/W2END[6]
+ Tile_X0Y13_W_IO/W2END[7] Tile_X1Y13_LUT4AB/W2END[0] Tile_X1Y13_LUT4AB/W2END[1] Tile_X1Y13_LUT4AB/W2END[2]
+ Tile_X1Y13_LUT4AB/W2END[3] Tile_X1Y13_LUT4AB/W2END[4] Tile_X1Y13_LUT4AB/W2END[5]
+ Tile_X1Y13_LUT4AB/W2END[6] Tile_X1Y13_LUT4AB/W2END[7] Tile_X2Y13_LUT4AB/W2BEG[0]
+ Tile_X2Y13_LUT4AB/W2BEG[1] Tile_X2Y13_LUT4AB/W2BEG[2] Tile_X2Y13_LUT4AB/W2BEG[3]
+ Tile_X2Y13_LUT4AB/W2BEG[4] Tile_X2Y13_LUT4AB/W2BEG[5] Tile_X2Y13_LUT4AB/W2BEG[6]
+ Tile_X2Y13_LUT4AB/W2BEG[7] Tile_X0Y13_W_IO/W6END[0] Tile_X0Y13_W_IO/W6END[10] Tile_X0Y13_W_IO/W6END[11]
+ Tile_X0Y13_W_IO/W6END[1] Tile_X0Y13_W_IO/W6END[2] Tile_X0Y13_W_IO/W6END[3] Tile_X0Y13_W_IO/W6END[4]
+ Tile_X0Y13_W_IO/W6END[5] Tile_X0Y13_W_IO/W6END[6] Tile_X0Y13_W_IO/W6END[7] Tile_X0Y13_W_IO/W6END[8]
+ Tile_X0Y13_W_IO/W6END[9] Tile_X2Y13_LUT4AB/W6BEG[0] Tile_X2Y13_LUT4AB/W6BEG[10]
+ Tile_X2Y13_LUT4AB/W6BEG[11] Tile_X2Y13_LUT4AB/W6BEG[1] Tile_X2Y13_LUT4AB/W6BEG[2]
+ Tile_X2Y13_LUT4AB/W6BEG[3] Tile_X2Y13_LUT4AB/W6BEG[4] Tile_X2Y13_LUT4AB/W6BEG[5]
+ Tile_X2Y13_LUT4AB/W6BEG[6] Tile_X2Y13_LUT4AB/W6BEG[7] Tile_X2Y13_LUT4AB/W6BEG[8]
+ Tile_X2Y13_LUT4AB/W6BEG[9] Tile_X0Y13_W_IO/WW4END[0] Tile_X0Y13_W_IO/WW4END[10]
+ Tile_X0Y13_W_IO/WW4END[11] Tile_X0Y13_W_IO/WW4END[12] Tile_X0Y13_W_IO/WW4END[13]
+ Tile_X0Y13_W_IO/WW4END[14] Tile_X0Y13_W_IO/WW4END[15] Tile_X0Y13_W_IO/WW4END[1]
+ Tile_X0Y13_W_IO/WW4END[2] Tile_X0Y13_W_IO/WW4END[3] Tile_X0Y13_W_IO/WW4END[4] Tile_X0Y13_W_IO/WW4END[5]
+ Tile_X0Y13_W_IO/WW4END[6] Tile_X0Y13_W_IO/WW4END[7] Tile_X0Y13_W_IO/WW4END[8] Tile_X0Y13_W_IO/WW4END[9]
+ Tile_X2Y13_LUT4AB/WW4BEG[0] Tile_X2Y13_LUT4AB/WW4BEG[10] Tile_X2Y13_LUT4AB/WW4BEG[11]
+ Tile_X2Y13_LUT4AB/WW4BEG[12] Tile_X2Y13_LUT4AB/WW4BEG[13] Tile_X2Y13_LUT4AB/WW4BEG[14]
+ Tile_X2Y13_LUT4AB/WW4BEG[15] Tile_X2Y13_LUT4AB/WW4BEG[1] Tile_X2Y13_LUT4AB/WW4BEG[2]
+ Tile_X2Y13_LUT4AB/WW4BEG[3] Tile_X2Y13_LUT4AB/WW4BEG[4] Tile_X2Y13_LUT4AB/WW4BEG[5]
+ Tile_X2Y13_LUT4AB/WW4BEG[6] Tile_X2Y13_LUT4AB/WW4BEG[7] Tile_X2Y13_LUT4AB/WW4BEG[8]
+ Tile_X2Y13_LUT4AB/WW4BEG[9] LUT4AB
XTile_X6Y8_LUT4AB Tile_X6Y9_LUT4AB/Co Tile_X6Y8_LUT4AB/Co Tile_X6Y8_LUT4AB/E1BEG[0]
+ Tile_X6Y8_LUT4AB/E1BEG[1] Tile_X6Y8_LUT4AB/E1BEG[2] Tile_X6Y8_LUT4AB/E1BEG[3] Tile_X6Y8_LUT4AB/E1END[0]
+ Tile_X6Y8_LUT4AB/E1END[1] Tile_X6Y8_LUT4AB/E1END[2] Tile_X6Y8_LUT4AB/E1END[3] Tile_X6Y8_LUT4AB/E2BEG[0]
+ Tile_X6Y8_LUT4AB/E2BEG[1] Tile_X6Y8_LUT4AB/E2BEG[2] Tile_X6Y8_LUT4AB/E2BEG[3] Tile_X6Y8_LUT4AB/E2BEG[4]
+ Tile_X6Y8_LUT4AB/E2BEG[5] Tile_X6Y8_LUT4AB/E2BEG[6] Tile_X6Y8_LUT4AB/E2BEG[7] Tile_X6Y8_LUT4AB/E2BEGb[0]
+ Tile_X6Y8_LUT4AB/E2BEGb[1] Tile_X6Y8_LUT4AB/E2BEGb[2] Tile_X6Y8_LUT4AB/E2BEGb[3]
+ Tile_X6Y8_LUT4AB/E2BEGb[4] Tile_X6Y8_LUT4AB/E2BEGb[5] Tile_X6Y8_LUT4AB/E2BEGb[6]
+ Tile_X6Y8_LUT4AB/E2BEGb[7] Tile_X6Y8_LUT4AB/E2END[0] Tile_X6Y8_LUT4AB/E2END[1] Tile_X6Y8_LUT4AB/E2END[2]
+ Tile_X6Y8_LUT4AB/E2END[3] Tile_X6Y8_LUT4AB/E2END[4] Tile_X6Y8_LUT4AB/E2END[5] Tile_X6Y8_LUT4AB/E2END[6]
+ Tile_X6Y8_LUT4AB/E2END[7] Tile_X6Y8_LUT4AB/E2MID[0] Tile_X6Y8_LUT4AB/E2MID[1] Tile_X6Y8_LUT4AB/E2MID[2]
+ Tile_X6Y8_LUT4AB/E2MID[3] Tile_X6Y8_LUT4AB/E2MID[4] Tile_X6Y8_LUT4AB/E2MID[5] Tile_X6Y8_LUT4AB/E2MID[6]
+ Tile_X6Y8_LUT4AB/E2MID[7] Tile_X6Y8_LUT4AB/E6BEG[0] Tile_X6Y8_LUT4AB/E6BEG[10] Tile_X6Y8_LUT4AB/E6BEG[11]
+ Tile_X6Y8_LUT4AB/E6BEG[1] Tile_X6Y8_LUT4AB/E6BEG[2] Tile_X6Y8_LUT4AB/E6BEG[3] Tile_X6Y8_LUT4AB/E6BEG[4]
+ Tile_X6Y8_LUT4AB/E6BEG[5] Tile_X6Y8_LUT4AB/E6BEG[6] Tile_X6Y8_LUT4AB/E6BEG[7] Tile_X6Y8_LUT4AB/E6BEG[8]
+ Tile_X6Y8_LUT4AB/E6BEG[9] Tile_X6Y8_LUT4AB/E6END[0] Tile_X6Y8_LUT4AB/E6END[10] Tile_X6Y8_LUT4AB/E6END[11]
+ Tile_X6Y8_LUT4AB/E6END[1] Tile_X6Y8_LUT4AB/E6END[2] Tile_X6Y8_LUT4AB/E6END[3] Tile_X6Y8_LUT4AB/E6END[4]
+ Tile_X6Y8_LUT4AB/E6END[5] Tile_X6Y8_LUT4AB/E6END[6] Tile_X6Y8_LUT4AB/E6END[7] Tile_X6Y8_LUT4AB/E6END[8]
+ Tile_X6Y8_LUT4AB/E6END[9] Tile_X6Y8_LUT4AB/EE4BEG[0] Tile_X6Y8_LUT4AB/EE4BEG[10]
+ Tile_X6Y8_LUT4AB/EE4BEG[11] Tile_X6Y8_LUT4AB/EE4BEG[12] Tile_X6Y8_LUT4AB/EE4BEG[13]
+ Tile_X6Y8_LUT4AB/EE4BEG[14] Tile_X6Y8_LUT4AB/EE4BEG[15] Tile_X6Y8_LUT4AB/EE4BEG[1]
+ Tile_X6Y8_LUT4AB/EE4BEG[2] Tile_X6Y8_LUT4AB/EE4BEG[3] Tile_X6Y8_LUT4AB/EE4BEG[4]
+ Tile_X6Y8_LUT4AB/EE4BEG[5] Tile_X6Y8_LUT4AB/EE4BEG[6] Tile_X6Y8_LUT4AB/EE4BEG[7]
+ Tile_X6Y8_LUT4AB/EE4BEG[8] Tile_X6Y8_LUT4AB/EE4BEG[9] Tile_X6Y8_LUT4AB/EE4END[0]
+ Tile_X6Y8_LUT4AB/EE4END[10] Tile_X6Y8_LUT4AB/EE4END[11] Tile_X6Y8_LUT4AB/EE4END[12]
+ Tile_X6Y8_LUT4AB/EE4END[13] Tile_X6Y8_LUT4AB/EE4END[14] Tile_X6Y8_LUT4AB/EE4END[15]
+ Tile_X6Y8_LUT4AB/EE4END[1] Tile_X6Y8_LUT4AB/EE4END[2] Tile_X6Y8_LUT4AB/EE4END[3]
+ Tile_X6Y8_LUT4AB/EE4END[4] Tile_X6Y8_LUT4AB/EE4END[5] Tile_X6Y8_LUT4AB/EE4END[6]
+ Tile_X6Y8_LUT4AB/EE4END[7] Tile_X6Y8_LUT4AB/EE4END[8] Tile_X6Y8_LUT4AB/EE4END[9]
+ Tile_X6Y8_LUT4AB/FrameData[0] Tile_X6Y8_LUT4AB/FrameData[10] Tile_X6Y8_LUT4AB/FrameData[11]
+ Tile_X6Y8_LUT4AB/FrameData[12] Tile_X6Y8_LUT4AB/FrameData[13] Tile_X6Y8_LUT4AB/FrameData[14]
+ Tile_X6Y8_LUT4AB/FrameData[15] Tile_X6Y8_LUT4AB/FrameData[16] Tile_X6Y8_LUT4AB/FrameData[17]
+ Tile_X6Y8_LUT4AB/FrameData[18] Tile_X6Y8_LUT4AB/FrameData[19] Tile_X6Y8_LUT4AB/FrameData[1]
+ Tile_X6Y8_LUT4AB/FrameData[20] Tile_X6Y8_LUT4AB/FrameData[21] Tile_X6Y8_LUT4AB/FrameData[22]
+ Tile_X6Y8_LUT4AB/FrameData[23] Tile_X6Y8_LUT4AB/FrameData[24] Tile_X6Y8_LUT4AB/FrameData[25]
+ Tile_X6Y8_LUT4AB/FrameData[26] Tile_X6Y8_LUT4AB/FrameData[27] Tile_X6Y8_LUT4AB/FrameData[28]
+ Tile_X6Y8_LUT4AB/FrameData[29] Tile_X6Y8_LUT4AB/FrameData[2] Tile_X6Y8_LUT4AB/FrameData[30]
+ Tile_X6Y8_LUT4AB/FrameData[31] Tile_X6Y8_LUT4AB/FrameData[3] Tile_X6Y8_LUT4AB/FrameData[4]
+ Tile_X6Y8_LUT4AB/FrameData[5] Tile_X6Y8_LUT4AB/FrameData[6] Tile_X6Y8_LUT4AB/FrameData[7]
+ Tile_X6Y8_LUT4AB/FrameData[8] Tile_X6Y8_LUT4AB/FrameData[9] Tile_X6Y8_LUT4AB/FrameData_O[0]
+ Tile_X6Y8_LUT4AB/FrameData_O[10] Tile_X6Y8_LUT4AB/FrameData_O[11] Tile_X6Y8_LUT4AB/FrameData_O[12]
+ Tile_X6Y8_LUT4AB/FrameData_O[13] Tile_X6Y8_LUT4AB/FrameData_O[14] Tile_X6Y8_LUT4AB/FrameData_O[15]
+ Tile_X6Y8_LUT4AB/FrameData_O[16] Tile_X6Y8_LUT4AB/FrameData_O[17] Tile_X6Y8_LUT4AB/FrameData_O[18]
+ Tile_X6Y8_LUT4AB/FrameData_O[19] Tile_X6Y8_LUT4AB/FrameData_O[1] Tile_X6Y8_LUT4AB/FrameData_O[20]
+ Tile_X6Y8_LUT4AB/FrameData_O[21] Tile_X6Y8_LUT4AB/FrameData_O[22] Tile_X6Y8_LUT4AB/FrameData_O[23]
+ Tile_X6Y8_LUT4AB/FrameData_O[24] Tile_X6Y8_LUT4AB/FrameData_O[25] Tile_X6Y8_LUT4AB/FrameData_O[26]
+ Tile_X6Y8_LUT4AB/FrameData_O[27] Tile_X6Y8_LUT4AB/FrameData_O[28] Tile_X6Y8_LUT4AB/FrameData_O[29]
+ Tile_X6Y8_LUT4AB/FrameData_O[2] Tile_X6Y8_LUT4AB/FrameData_O[30] Tile_X6Y8_LUT4AB/FrameData_O[31]
+ Tile_X6Y8_LUT4AB/FrameData_O[3] Tile_X6Y8_LUT4AB/FrameData_O[4] Tile_X6Y8_LUT4AB/FrameData_O[5]
+ Tile_X6Y8_LUT4AB/FrameData_O[6] Tile_X6Y8_LUT4AB/FrameData_O[7] Tile_X6Y8_LUT4AB/FrameData_O[8]
+ Tile_X6Y8_LUT4AB/FrameData_O[9] Tile_X6Y8_LUT4AB/FrameStrobe[0] Tile_X6Y8_LUT4AB/FrameStrobe[10]
+ Tile_X6Y8_LUT4AB/FrameStrobe[11] Tile_X6Y8_LUT4AB/FrameStrobe[12] Tile_X6Y8_LUT4AB/FrameStrobe[13]
+ Tile_X6Y8_LUT4AB/FrameStrobe[14] Tile_X6Y8_LUT4AB/FrameStrobe[15] Tile_X6Y8_LUT4AB/FrameStrobe[16]
+ Tile_X6Y8_LUT4AB/FrameStrobe[17] Tile_X6Y8_LUT4AB/FrameStrobe[18] Tile_X6Y8_LUT4AB/FrameStrobe[19]
+ Tile_X6Y8_LUT4AB/FrameStrobe[1] Tile_X6Y8_LUT4AB/FrameStrobe[2] Tile_X6Y8_LUT4AB/FrameStrobe[3]
+ Tile_X6Y8_LUT4AB/FrameStrobe[4] Tile_X6Y8_LUT4AB/FrameStrobe[5] Tile_X6Y8_LUT4AB/FrameStrobe[6]
+ Tile_X6Y8_LUT4AB/FrameStrobe[7] Tile_X6Y8_LUT4AB/FrameStrobe[8] Tile_X6Y8_LUT4AB/FrameStrobe[9]
+ Tile_X6Y7_LUT4AB/FrameStrobe[0] Tile_X6Y7_LUT4AB/FrameStrobe[10] Tile_X6Y7_LUT4AB/FrameStrobe[11]
+ Tile_X6Y7_LUT4AB/FrameStrobe[12] Tile_X6Y7_LUT4AB/FrameStrobe[13] Tile_X6Y7_LUT4AB/FrameStrobe[14]
+ Tile_X6Y7_LUT4AB/FrameStrobe[15] Tile_X6Y7_LUT4AB/FrameStrobe[16] Tile_X6Y7_LUT4AB/FrameStrobe[17]
+ Tile_X6Y7_LUT4AB/FrameStrobe[18] Tile_X6Y7_LUT4AB/FrameStrobe[19] Tile_X6Y7_LUT4AB/FrameStrobe[1]
+ Tile_X6Y7_LUT4AB/FrameStrobe[2] Tile_X6Y7_LUT4AB/FrameStrobe[3] Tile_X6Y7_LUT4AB/FrameStrobe[4]
+ Tile_X6Y7_LUT4AB/FrameStrobe[5] Tile_X6Y7_LUT4AB/FrameStrobe[6] Tile_X6Y7_LUT4AB/FrameStrobe[7]
+ Tile_X6Y7_LUT4AB/FrameStrobe[8] Tile_X6Y7_LUT4AB/FrameStrobe[9] Tile_X6Y8_LUT4AB/N1BEG[0]
+ Tile_X6Y8_LUT4AB/N1BEG[1] Tile_X6Y8_LUT4AB/N1BEG[2] Tile_X6Y8_LUT4AB/N1BEG[3] Tile_X6Y9_LUT4AB/N1BEG[0]
+ Tile_X6Y9_LUT4AB/N1BEG[1] Tile_X6Y9_LUT4AB/N1BEG[2] Tile_X6Y9_LUT4AB/N1BEG[3] Tile_X6Y8_LUT4AB/N2BEG[0]
+ Tile_X6Y8_LUT4AB/N2BEG[1] Tile_X6Y8_LUT4AB/N2BEG[2] Tile_X6Y8_LUT4AB/N2BEG[3] Tile_X6Y8_LUT4AB/N2BEG[4]
+ Tile_X6Y8_LUT4AB/N2BEG[5] Tile_X6Y8_LUT4AB/N2BEG[6] Tile_X6Y8_LUT4AB/N2BEG[7] Tile_X6Y7_LUT4AB/N2END[0]
+ Tile_X6Y7_LUT4AB/N2END[1] Tile_X6Y7_LUT4AB/N2END[2] Tile_X6Y7_LUT4AB/N2END[3] Tile_X6Y7_LUT4AB/N2END[4]
+ Tile_X6Y7_LUT4AB/N2END[5] Tile_X6Y7_LUT4AB/N2END[6] Tile_X6Y7_LUT4AB/N2END[7] Tile_X6Y8_LUT4AB/N2END[0]
+ Tile_X6Y8_LUT4AB/N2END[1] Tile_X6Y8_LUT4AB/N2END[2] Tile_X6Y8_LUT4AB/N2END[3] Tile_X6Y8_LUT4AB/N2END[4]
+ Tile_X6Y8_LUT4AB/N2END[5] Tile_X6Y8_LUT4AB/N2END[6] Tile_X6Y8_LUT4AB/N2END[7] Tile_X6Y9_LUT4AB/N2BEG[0]
+ Tile_X6Y9_LUT4AB/N2BEG[1] Tile_X6Y9_LUT4AB/N2BEG[2] Tile_X6Y9_LUT4AB/N2BEG[3] Tile_X6Y9_LUT4AB/N2BEG[4]
+ Tile_X6Y9_LUT4AB/N2BEG[5] Tile_X6Y9_LUT4AB/N2BEG[6] Tile_X6Y9_LUT4AB/N2BEG[7] Tile_X6Y8_LUT4AB/N4BEG[0]
+ Tile_X6Y8_LUT4AB/N4BEG[10] Tile_X6Y8_LUT4AB/N4BEG[11] Tile_X6Y8_LUT4AB/N4BEG[12]
+ Tile_X6Y8_LUT4AB/N4BEG[13] Tile_X6Y8_LUT4AB/N4BEG[14] Tile_X6Y8_LUT4AB/N4BEG[15]
+ Tile_X6Y8_LUT4AB/N4BEG[1] Tile_X6Y8_LUT4AB/N4BEG[2] Tile_X6Y8_LUT4AB/N4BEG[3] Tile_X6Y8_LUT4AB/N4BEG[4]
+ Tile_X6Y8_LUT4AB/N4BEG[5] Tile_X6Y8_LUT4AB/N4BEG[6] Tile_X6Y8_LUT4AB/N4BEG[7] Tile_X6Y8_LUT4AB/N4BEG[8]
+ Tile_X6Y8_LUT4AB/N4BEG[9] Tile_X6Y9_LUT4AB/N4BEG[0] Tile_X6Y9_LUT4AB/N4BEG[10] Tile_X6Y9_LUT4AB/N4BEG[11]
+ Tile_X6Y9_LUT4AB/N4BEG[12] Tile_X6Y9_LUT4AB/N4BEG[13] Tile_X6Y9_LUT4AB/N4BEG[14]
+ Tile_X6Y9_LUT4AB/N4BEG[15] Tile_X6Y9_LUT4AB/N4BEG[1] Tile_X6Y9_LUT4AB/N4BEG[2] Tile_X6Y9_LUT4AB/N4BEG[3]
+ Tile_X6Y9_LUT4AB/N4BEG[4] Tile_X6Y9_LUT4AB/N4BEG[5] Tile_X6Y9_LUT4AB/N4BEG[6] Tile_X6Y9_LUT4AB/N4BEG[7]
+ Tile_X6Y9_LUT4AB/N4BEG[8] Tile_X6Y9_LUT4AB/N4BEG[9] Tile_X6Y8_LUT4AB/NN4BEG[0] Tile_X6Y8_LUT4AB/NN4BEG[10]
+ Tile_X6Y8_LUT4AB/NN4BEG[11] Tile_X6Y8_LUT4AB/NN4BEG[12] Tile_X6Y8_LUT4AB/NN4BEG[13]
+ Tile_X6Y8_LUT4AB/NN4BEG[14] Tile_X6Y8_LUT4AB/NN4BEG[15] Tile_X6Y8_LUT4AB/NN4BEG[1]
+ Tile_X6Y8_LUT4AB/NN4BEG[2] Tile_X6Y8_LUT4AB/NN4BEG[3] Tile_X6Y8_LUT4AB/NN4BEG[4]
+ Tile_X6Y8_LUT4AB/NN4BEG[5] Tile_X6Y8_LUT4AB/NN4BEG[6] Tile_X6Y8_LUT4AB/NN4BEG[7]
+ Tile_X6Y8_LUT4AB/NN4BEG[8] Tile_X6Y8_LUT4AB/NN4BEG[9] Tile_X6Y9_LUT4AB/NN4BEG[0]
+ Tile_X6Y9_LUT4AB/NN4BEG[10] Tile_X6Y9_LUT4AB/NN4BEG[11] Tile_X6Y9_LUT4AB/NN4BEG[12]
+ Tile_X6Y9_LUT4AB/NN4BEG[13] Tile_X6Y9_LUT4AB/NN4BEG[14] Tile_X6Y9_LUT4AB/NN4BEG[15]
+ Tile_X6Y9_LUT4AB/NN4BEG[1] Tile_X6Y9_LUT4AB/NN4BEG[2] Tile_X6Y9_LUT4AB/NN4BEG[3]
+ Tile_X6Y9_LUT4AB/NN4BEG[4] Tile_X6Y9_LUT4AB/NN4BEG[5] Tile_X6Y9_LUT4AB/NN4BEG[6]
+ Tile_X6Y9_LUT4AB/NN4BEG[7] Tile_X6Y9_LUT4AB/NN4BEG[8] Tile_X6Y9_LUT4AB/NN4BEG[9]
+ Tile_X6Y9_LUT4AB/S1END[0] Tile_X6Y9_LUT4AB/S1END[1] Tile_X6Y9_LUT4AB/S1END[2] Tile_X6Y9_LUT4AB/S1END[3]
+ Tile_X6Y8_LUT4AB/S1END[0] Tile_X6Y8_LUT4AB/S1END[1] Tile_X6Y8_LUT4AB/S1END[2] Tile_X6Y8_LUT4AB/S1END[3]
+ Tile_X6Y9_LUT4AB/S2MID[0] Tile_X6Y9_LUT4AB/S2MID[1] Tile_X6Y9_LUT4AB/S2MID[2] Tile_X6Y9_LUT4AB/S2MID[3]
+ Tile_X6Y9_LUT4AB/S2MID[4] Tile_X6Y9_LUT4AB/S2MID[5] Tile_X6Y9_LUT4AB/S2MID[6] Tile_X6Y9_LUT4AB/S2MID[7]
+ Tile_X6Y9_LUT4AB/S2END[0] Tile_X6Y9_LUT4AB/S2END[1] Tile_X6Y9_LUT4AB/S2END[2] Tile_X6Y9_LUT4AB/S2END[3]
+ Tile_X6Y9_LUT4AB/S2END[4] Tile_X6Y9_LUT4AB/S2END[5] Tile_X6Y9_LUT4AB/S2END[6] Tile_X6Y9_LUT4AB/S2END[7]
+ Tile_X6Y8_LUT4AB/S2END[0] Tile_X6Y8_LUT4AB/S2END[1] Tile_X6Y8_LUT4AB/S2END[2] Tile_X6Y8_LUT4AB/S2END[3]
+ Tile_X6Y8_LUT4AB/S2END[4] Tile_X6Y8_LUT4AB/S2END[5] Tile_X6Y8_LUT4AB/S2END[6] Tile_X6Y8_LUT4AB/S2END[7]
+ Tile_X6Y8_LUT4AB/S2MID[0] Tile_X6Y8_LUT4AB/S2MID[1] Tile_X6Y8_LUT4AB/S2MID[2] Tile_X6Y8_LUT4AB/S2MID[3]
+ Tile_X6Y8_LUT4AB/S2MID[4] Tile_X6Y8_LUT4AB/S2MID[5] Tile_X6Y8_LUT4AB/S2MID[6] Tile_X6Y8_LUT4AB/S2MID[7]
+ Tile_X6Y9_LUT4AB/S4END[0] Tile_X6Y9_LUT4AB/S4END[10] Tile_X6Y9_LUT4AB/S4END[11]
+ Tile_X6Y9_LUT4AB/S4END[12] Tile_X6Y9_LUT4AB/S4END[13] Tile_X6Y9_LUT4AB/S4END[14]
+ Tile_X6Y9_LUT4AB/S4END[15] Tile_X6Y9_LUT4AB/S4END[1] Tile_X6Y9_LUT4AB/S4END[2] Tile_X6Y9_LUT4AB/S4END[3]
+ Tile_X6Y9_LUT4AB/S4END[4] Tile_X6Y9_LUT4AB/S4END[5] Tile_X6Y9_LUT4AB/S4END[6] Tile_X6Y9_LUT4AB/S4END[7]
+ Tile_X6Y9_LUT4AB/S4END[8] Tile_X6Y9_LUT4AB/S4END[9] Tile_X6Y8_LUT4AB/S4END[0] Tile_X6Y8_LUT4AB/S4END[10]
+ Tile_X6Y8_LUT4AB/S4END[11] Tile_X6Y8_LUT4AB/S4END[12] Tile_X6Y8_LUT4AB/S4END[13]
+ Tile_X6Y8_LUT4AB/S4END[14] Tile_X6Y8_LUT4AB/S4END[15] Tile_X6Y8_LUT4AB/S4END[1]
+ Tile_X6Y8_LUT4AB/S4END[2] Tile_X6Y8_LUT4AB/S4END[3] Tile_X6Y8_LUT4AB/S4END[4] Tile_X6Y8_LUT4AB/S4END[5]
+ Tile_X6Y8_LUT4AB/S4END[6] Tile_X6Y8_LUT4AB/S4END[7] Tile_X6Y8_LUT4AB/S4END[8] Tile_X6Y8_LUT4AB/S4END[9]
+ Tile_X6Y9_LUT4AB/SS4END[0] Tile_X6Y9_LUT4AB/SS4END[10] Tile_X6Y9_LUT4AB/SS4END[11]
+ Tile_X6Y9_LUT4AB/SS4END[12] Tile_X6Y9_LUT4AB/SS4END[13] Tile_X6Y9_LUT4AB/SS4END[14]
+ Tile_X6Y9_LUT4AB/SS4END[15] Tile_X6Y9_LUT4AB/SS4END[1] Tile_X6Y9_LUT4AB/SS4END[2]
+ Tile_X6Y9_LUT4AB/SS4END[3] Tile_X6Y9_LUT4AB/SS4END[4] Tile_X6Y9_LUT4AB/SS4END[5]
+ Tile_X6Y9_LUT4AB/SS4END[6] Tile_X6Y9_LUT4AB/SS4END[7] Tile_X6Y9_LUT4AB/SS4END[8]
+ Tile_X6Y9_LUT4AB/SS4END[9] Tile_X6Y8_LUT4AB/SS4END[0] Tile_X6Y8_LUT4AB/SS4END[10]
+ Tile_X6Y8_LUT4AB/SS4END[11] Tile_X6Y8_LUT4AB/SS4END[12] Tile_X6Y8_LUT4AB/SS4END[13]
+ Tile_X6Y8_LUT4AB/SS4END[14] Tile_X6Y8_LUT4AB/SS4END[15] Tile_X6Y8_LUT4AB/SS4END[1]
+ Tile_X6Y8_LUT4AB/SS4END[2] Tile_X6Y8_LUT4AB/SS4END[3] Tile_X6Y8_LUT4AB/SS4END[4]
+ Tile_X6Y8_LUT4AB/SS4END[5] Tile_X6Y8_LUT4AB/SS4END[6] Tile_X6Y8_LUT4AB/SS4END[7]
+ Tile_X6Y8_LUT4AB/SS4END[8] Tile_X6Y8_LUT4AB/SS4END[9] Tile_X6Y8_LUT4AB/UserCLK Tile_X6Y7_LUT4AB/UserCLK
+ VGND VPWR Tile_X6Y8_LUT4AB/W1BEG[0] Tile_X6Y8_LUT4AB/W1BEG[1] Tile_X6Y8_LUT4AB/W1BEG[2]
+ Tile_X6Y8_LUT4AB/W1BEG[3] Tile_X6Y8_LUT4AB/W1END[0] Tile_X6Y8_LUT4AB/W1END[1] Tile_X6Y8_LUT4AB/W1END[2]
+ Tile_X6Y8_LUT4AB/W1END[3] Tile_X6Y8_LUT4AB/W2BEG[0] Tile_X6Y8_LUT4AB/W2BEG[1] Tile_X6Y8_LUT4AB/W2BEG[2]
+ Tile_X6Y8_LUT4AB/W2BEG[3] Tile_X6Y8_LUT4AB/W2BEG[4] Tile_X6Y8_LUT4AB/W2BEG[5] Tile_X6Y8_LUT4AB/W2BEG[6]
+ Tile_X6Y8_LUT4AB/W2BEG[7] Tile_X5Y8_LUT4AB/W2END[0] Tile_X5Y8_LUT4AB/W2END[1] Tile_X5Y8_LUT4AB/W2END[2]
+ Tile_X5Y8_LUT4AB/W2END[3] Tile_X5Y8_LUT4AB/W2END[4] Tile_X5Y8_LUT4AB/W2END[5] Tile_X5Y8_LUT4AB/W2END[6]
+ Tile_X5Y8_LUT4AB/W2END[7] Tile_X6Y8_LUT4AB/W2END[0] Tile_X6Y8_LUT4AB/W2END[1] Tile_X6Y8_LUT4AB/W2END[2]
+ Tile_X6Y8_LUT4AB/W2END[3] Tile_X6Y8_LUT4AB/W2END[4] Tile_X6Y8_LUT4AB/W2END[5] Tile_X6Y8_LUT4AB/W2END[6]
+ Tile_X6Y8_LUT4AB/W2END[7] Tile_X6Y8_LUT4AB/W2MID[0] Tile_X6Y8_LUT4AB/W2MID[1] Tile_X6Y8_LUT4AB/W2MID[2]
+ Tile_X6Y8_LUT4AB/W2MID[3] Tile_X6Y8_LUT4AB/W2MID[4] Tile_X6Y8_LUT4AB/W2MID[5] Tile_X6Y8_LUT4AB/W2MID[6]
+ Tile_X6Y8_LUT4AB/W2MID[7] Tile_X6Y8_LUT4AB/W6BEG[0] Tile_X6Y8_LUT4AB/W6BEG[10] Tile_X6Y8_LUT4AB/W6BEG[11]
+ Tile_X6Y8_LUT4AB/W6BEG[1] Tile_X6Y8_LUT4AB/W6BEG[2] Tile_X6Y8_LUT4AB/W6BEG[3] Tile_X6Y8_LUT4AB/W6BEG[4]
+ Tile_X6Y8_LUT4AB/W6BEG[5] Tile_X6Y8_LUT4AB/W6BEG[6] Tile_X6Y8_LUT4AB/W6BEG[7] Tile_X6Y8_LUT4AB/W6BEG[8]
+ Tile_X6Y8_LUT4AB/W6BEG[9] Tile_X6Y8_LUT4AB/W6END[0] Tile_X6Y8_LUT4AB/W6END[10] Tile_X6Y8_LUT4AB/W6END[11]
+ Tile_X6Y8_LUT4AB/W6END[1] Tile_X6Y8_LUT4AB/W6END[2] Tile_X6Y8_LUT4AB/W6END[3] Tile_X6Y8_LUT4AB/W6END[4]
+ Tile_X6Y8_LUT4AB/W6END[5] Tile_X6Y8_LUT4AB/W6END[6] Tile_X6Y8_LUT4AB/W6END[7] Tile_X6Y8_LUT4AB/W6END[8]
+ Tile_X6Y8_LUT4AB/W6END[9] Tile_X6Y8_LUT4AB/WW4BEG[0] Tile_X6Y8_LUT4AB/WW4BEG[10]
+ Tile_X6Y8_LUT4AB/WW4BEG[11] Tile_X6Y8_LUT4AB/WW4BEG[12] Tile_X6Y8_LUT4AB/WW4BEG[13]
+ Tile_X6Y8_LUT4AB/WW4BEG[14] Tile_X6Y8_LUT4AB/WW4BEG[15] Tile_X6Y8_LUT4AB/WW4BEG[1]
+ Tile_X6Y8_LUT4AB/WW4BEG[2] Tile_X6Y8_LUT4AB/WW4BEG[3] Tile_X6Y8_LUT4AB/WW4BEG[4]
+ Tile_X6Y8_LUT4AB/WW4BEG[5] Tile_X6Y8_LUT4AB/WW4BEG[6] Tile_X6Y8_LUT4AB/WW4BEG[7]
+ Tile_X6Y8_LUT4AB/WW4BEG[8] Tile_X6Y8_LUT4AB/WW4BEG[9] Tile_X6Y8_LUT4AB/WW4END[0]
+ Tile_X6Y8_LUT4AB/WW4END[10] Tile_X6Y8_LUT4AB/WW4END[11] Tile_X6Y8_LUT4AB/WW4END[12]
+ Tile_X6Y8_LUT4AB/WW4END[13] Tile_X6Y8_LUT4AB/WW4END[14] Tile_X6Y8_LUT4AB/WW4END[15]
+ Tile_X6Y8_LUT4AB/WW4END[1] Tile_X6Y8_LUT4AB/WW4END[2] Tile_X6Y8_LUT4AB/WW4END[3]
+ Tile_X6Y8_LUT4AB/WW4END[4] Tile_X6Y8_LUT4AB/WW4END[5] Tile_X6Y8_LUT4AB/WW4END[6]
+ Tile_X6Y8_LUT4AB/WW4END[7] Tile_X6Y8_LUT4AB/WW4END[8] Tile_X6Y8_LUT4AB/WW4END[9]
+ LUT4AB
.ends

