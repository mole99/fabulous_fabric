module eFPGA
    #(
        parameter MaxFramesPerCol=20,
        parameter FrameBitsPerRow=32
    )
    (
        input Tile_X1Y0_A_O_top, //EXTERNAL
        output Tile_X1Y0_A_I_top, //EXTERNAL
        output Tile_X1Y0_A_T_top, //EXTERNAL
        input Tile_X1Y0_B_O_top, //EXTERNAL
        output Tile_X1Y0_B_I_top, //EXTERNAL
        output Tile_X1Y0_B_T_top, //EXTERNAL
        output Tile_X1Y0_A_config_C_bit0, //EXTERNAL
        output Tile_X1Y0_A_config_C_bit1, //EXTERNAL
        output Tile_X1Y0_A_config_C_bit2, //EXTERNAL
        output Tile_X1Y0_A_config_C_bit3, //EXTERNAL
        output Tile_X1Y0_B_config_C_bit0, //EXTERNAL
        output Tile_X1Y0_B_config_C_bit1, //EXTERNAL
        output Tile_X1Y0_B_config_C_bit2, //EXTERNAL
        output Tile_X1Y0_B_config_C_bit3, //EXTERNAL
        input Tile_X2Y0_A_O_top, //EXTERNAL
        output Tile_X2Y0_A_I_top, //EXTERNAL
        output Tile_X2Y0_A_T_top, //EXTERNAL
        input Tile_X2Y0_B_O_top, //EXTERNAL
        output Tile_X2Y0_B_I_top, //EXTERNAL
        output Tile_X2Y0_B_T_top, //EXTERNAL
        output Tile_X2Y0_A_config_C_bit0, //EXTERNAL
        output Tile_X2Y0_A_config_C_bit1, //EXTERNAL
        output Tile_X2Y0_A_config_C_bit2, //EXTERNAL
        output Tile_X2Y0_A_config_C_bit3, //EXTERNAL
        output Tile_X2Y0_B_config_C_bit0, //EXTERNAL
        output Tile_X2Y0_B_config_C_bit1, //EXTERNAL
        output Tile_X2Y0_B_config_C_bit2, //EXTERNAL
        output Tile_X2Y0_B_config_C_bit3, //EXTERNAL
        input Tile_X0Y1_A_O_top, //EXTERNAL
        output Tile_X0Y1_A_I_top, //EXTERNAL
        output Tile_X0Y1_A_T_top, //EXTERNAL
        input Tile_X0Y1_B_O_top, //EXTERNAL
        output Tile_X0Y1_B_I_top, //EXTERNAL
        output Tile_X0Y1_B_T_top, //EXTERNAL
        output Tile_X0Y1_A_config_C_bit0, //EXTERNAL
        output Tile_X0Y1_A_config_C_bit1, //EXTERNAL
        output Tile_X0Y1_A_config_C_bit2, //EXTERNAL
        output Tile_X0Y1_A_config_C_bit3, //EXTERNAL
        output Tile_X0Y1_B_config_C_bit0, //EXTERNAL
        output Tile_X0Y1_B_config_C_bit1, //EXTERNAL
        output Tile_X0Y1_B_config_C_bit2, //EXTERNAL
        output Tile_X0Y1_B_config_C_bit3, //EXTERNAL
        input Tile_X0Y2_A_O_top, //EXTERNAL
        output Tile_X0Y2_A_I_top, //EXTERNAL
        output Tile_X0Y2_A_T_top, //EXTERNAL
        input Tile_X0Y2_B_O_top, //EXTERNAL
        output Tile_X0Y2_B_I_top, //EXTERNAL
        output Tile_X0Y2_B_T_top, //EXTERNAL
        output Tile_X0Y2_A_config_C_bit0, //EXTERNAL
        output Tile_X0Y2_A_config_C_bit1, //EXTERNAL
        output Tile_X0Y2_A_config_C_bit2, //EXTERNAL
        output Tile_X0Y2_A_config_C_bit3, //EXTERNAL
        output Tile_X0Y2_B_config_C_bit0, //EXTERNAL
        output Tile_X0Y2_B_config_C_bit1, //EXTERNAL
        output Tile_X0Y2_B_config_C_bit2, //EXTERNAL
        output Tile_X0Y2_B_config_C_bit3, //EXTERNAL
        input Tile_X10Y2_CONFIGURED_top, //EXTERNAL
        input Tile_X10Y2_DOUT_SRAM0, //EXTERNAL
        input Tile_X10Y2_DOUT_SRAM1, //EXTERNAL
        input Tile_X10Y2_DOUT_SRAM2, //EXTERNAL
        input Tile_X10Y2_DOUT_SRAM3, //EXTERNAL
        input Tile_X10Y2_DOUT_SRAM4, //EXTERNAL
        input Tile_X10Y2_DOUT_SRAM5, //EXTERNAL
        input Tile_X10Y2_DOUT_SRAM6, //EXTERNAL
        input Tile_X10Y2_DOUT_SRAM7, //EXTERNAL
        input Tile_X10Y2_DOUT_SRAM8, //EXTERNAL
        input Tile_X10Y2_DOUT_SRAM9, //EXTERNAL
        input Tile_X10Y2_DOUT_SRAM10, //EXTERNAL
        input Tile_X10Y2_DOUT_SRAM11, //EXTERNAL
        input Tile_X10Y2_DOUT_SRAM12, //EXTERNAL
        input Tile_X10Y2_DOUT_SRAM13, //EXTERNAL
        input Tile_X10Y2_DOUT_SRAM14, //EXTERNAL
        input Tile_X10Y2_DOUT_SRAM15, //EXTERNAL
        input Tile_X10Y2_DOUT_SRAM16, //EXTERNAL
        input Tile_X10Y2_DOUT_SRAM17, //EXTERNAL
        input Tile_X10Y2_DOUT_SRAM18, //EXTERNAL
        input Tile_X10Y2_DOUT_SRAM19, //EXTERNAL
        input Tile_X10Y2_DOUT_SRAM20, //EXTERNAL
        input Tile_X10Y2_DOUT_SRAM21, //EXTERNAL
        input Tile_X10Y2_DOUT_SRAM22, //EXTERNAL
        input Tile_X10Y2_DOUT_SRAM23, //EXTERNAL
        input Tile_X10Y2_DOUT_SRAM24, //EXTERNAL
        input Tile_X10Y2_DOUT_SRAM25, //EXTERNAL
        input Tile_X10Y2_DOUT_SRAM26, //EXTERNAL
        input Tile_X10Y2_DOUT_SRAM27, //EXTERNAL
        input Tile_X10Y2_DOUT_SRAM28, //EXTERNAL
        input Tile_X10Y2_DOUT_SRAM29, //EXTERNAL
        input Tile_X10Y2_DOUT_SRAM30, //EXTERNAL
        input Tile_X10Y2_DOUT_SRAM31, //EXTERNAL
        output Tile_X10Y2_ADDR_SRAM0, //EXTERNAL
        output Tile_X10Y2_ADDR_SRAM1, //EXTERNAL
        output Tile_X10Y2_ADDR_SRAM2, //EXTERNAL
        output Tile_X10Y2_ADDR_SRAM3, //EXTERNAL
        output Tile_X10Y2_ADDR_SRAM4, //EXTERNAL
        output Tile_X10Y2_ADDR_SRAM5, //EXTERNAL
        output Tile_X10Y2_ADDR_SRAM6, //EXTERNAL
        output Tile_X10Y2_ADDR_SRAM7, //EXTERNAL
        output Tile_X10Y2_ADDR_SRAM8, //EXTERNAL
        output Tile_X10Y2_ADDR_SRAM9, //EXTERNAL
        output Tile_X10Y2_BM_SRAM0, //EXTERNAL
        output Tile_X10Y2_BM_SRAM1, //EXTERNAL
        output Tile_X10Y2_BM_SRAM2, //EXTERNAL
        output Tile_X10Y2_BM_SRAM3, //EXTERNAL
        output Tile_X10Y2_BM_SRAM4, //EXTERNAL
        output Tile_X10Y2_BM_SRAM5, //EXTERNAL
        output Tile_X10Y2_BM_SRAM6, //EXTERNAL
        output Tile_X10Y2_BM_SRAM7, //EXTERNAL
        output Tile_X10Y2_BM_SRAM8, //EXTERNAL
        output Tile_X10Y2_BM_SRAM9, //EXTERNAL
        output Tile_X10Y2_BM_SRAM10, //EXTERNAL
        output Tile_X10Y2_BM_SRAM11, //EXTERNAL
        output Tile_X10Y2_BM_SRAM12, //EXTERNAL
        output Tile_X10Y2_BM_SRAM13, //EXTERNAL
        output Tile_X10Y2_BM_SRAM14, //EXTERNAL
        output Tile_X10Y2_BM_SRAM15, //EXTERNAL
        output Tile_X10Y2_BM_SRAM16, //EXTERNAL
        output Tile_X10Y2_BM_SRAM17, //EXTERNAL
        output Tile_X10Y2_BM_SRAM18, //EXTERNAL
        output Tile_X10Y2_BM_SRAM19, //EXTERNAL
        output Tile_X10Y2_BM_SRAM20, //EXTERNAL
        output Tile_X10Y2_BM_SRAM21, //EXTERNAL
        output Tile_X10Y2_BM_SRAM22, //EXTERNAL
        output Tile_X10Y2_BM_SRAM23, //EXTERNAL
        output Tile_X10Y2_BM_SRAM24, //EXTERNAL
        output Tile_X10Y2_BM_SRAM25, //EXTERNAL
        output Tile_X10Y2_BM_SRAM26, //EXTERNAL
        output Tile_X10Y2_BM_SRAM27, //EXTERNAL
        output Tile_X10Y2_BM_SRAM28, //EXTERNAL
        output Tile_X10Y2_BM_SRAM29, //EXTERNAL
        output Tile_X10Y2_BM_SRAM30, //EXTERNAL
        output Tile_X10Y2_BM_SRAM31, //EXTERNAL
        output Tile_X10Y2_CLK_SRAM, //EXTERNAL
        output Tile_X10Y2_DIN_SRAM0, //EXTERNAL
        output Tile_X10Y2_DIN_SRAM1, //EXTERNAL
        output Tile_X10Y2_DIN_SRAM2, //EXTERNAL
        output Tile_X10Y2_DIN_SRAM3, //EXTERNAL
        output Tile_X10Y2_DIN_SRAM4, //EXTERNAL
        output Tile_X10Y2_DIN_SRAM5, //EXTERNAL
        output Tile_X10Y2_DIN_SRAM6, //EXTERNAL
        output Tile_X10Y2_DIN_SRAM7, //EXTERNAL
        output Tile_X10Y2_DIN_SRAM8, //EXTERNAL
        output Tile_X10Y2_DIN_SRAM9, //EXTERNAL
        output Tile_X10Y2_DIN_SRAM10, //EXTERNAL
        output Tile_X10Y2_DIN_SRAM11, //EXTERNAL
        output Tile_X10Y2_DIN_SRAM12, //EXTERNAL
        output Tile_X10Y2_DIN_SRAM13, //EXTERNAL
        output Tile_X10Y2_DIN_SRAM14, //EXTERNAL
        output Tile_X10Y2_DIN_SRAM15, //EXTERNAL
        output Tile_X10Y2_DIN_SRAM16, //EXTERNAL
        output Tile_X10Y2_DIN_SRAM17, //EXTERNAL
        output Tile_X10Y2_DIN_SRAM18, //EXTERNAL
        output Tile_X10Y2_DIN_SRAM19, //EXTERNAL
        output Tile_X10Y2_DIN_SRAM20, //EXTERNAL
        output Tile_X10Y2_DIN_SRAM21, //EXTERNAL
        output Tile_X10Y2_DIN_SRAM22, //EXTERNAL
        output Tile_X10Y2_DIN_SRAM23, //EXTERNAL
        output Tile_X10Y2_DIN_SRAM24, //EXTERNAL
        output Tile_X10Y2_DIN_SRAM25, //EXTERNAL
        output Tile_X10Y2_DIN_SRAM26, //EXTERNAL
        output Tile_X10Y2_DIN_SRAM27, //EXTERNAL
        output Tile_X10Y2_DIN_SRAM28, //EXTERNAL
        output Tile_X10Y2_DIN_SRAM29, //EXTERNAL
        output Tile_X10Y2_DIN_SRAM30, //EXTERNAL
        output Tile_X10Y2_DIN_SRAM31, //EXTERNAL
        output Tile_X10Y2_MEN_SRAM, //EXTERNAL
        output Tile_X10Y2_REN_SRAM, //EXTERNAL
        output Tile_X10Y2_TIE_HIGH_SRAM, //EXTERNAL
        output Tile_X10Y2_TIE_LOW_SRAM, //EXTERNAL
        output Tile_X10Y2_WEN_SRAM, //EXTERNAL
        input Tile_X0Y3_A_O_top, //EXTERNAL
        output Tile_X0Y3_A_I_top, //EXTERNAL
        output Tile_X0Y3_A_T_top, //EXTERNAL
        input Tile_X0Y3_B_O_top, //EXTERNAL
        output Tile_X0Y3_B_I_top, //EXTERNAL
        output Tile_X0Y3_B_T_top, //EXTERNAL
        output Tile_X0Y3_A_config_C_bit0, //EXTERNAL
        output Tile_X0Y3_A_config_C_bit1, //EXTERNAL
        output Tile_X0Y3_A_config_C_bit2, //EXTERNAL
        output Tile_X0Y3_A_config_C_bit3, //EXTERNAL
        output Tile_X0Y3_B_config_C_bit0, //EXTERNAL
        output Tile_X0Y3_B_config_C_bit1, //EXTERNAL
        output Tile_X0Y3_B_config_C_bit2, //EXTERNAL
        output Tile_X0Y3_B_config_C_bit3, //EXTERNAL
        input Tile_X0Y4_A_O_top, //EXTERNAL
        output Tile_X0Y4_A_I_top, //EXTERNAL
        output Tile_X0Y4_A_T_top, //EXTERNAL
        input Tile_X0Y4_B_O_top, //EXTERNAL
        output Tile_X0Y4_B_I_top, //EXTERNAL
        output Tile_X0Y4_B_T_top, //EXTERNAL
        output Tile_X0Y4_A_config_C_bit0, //EXTERNAL
        output Tile_X0Y4_A_config_C_bit1, //EXTERNAL
        output Tile_X0Y4_A_config_C_bit2, //EXTERNAL
        output Tile_X0Y4_A_config_C_bit3, //EXTERNAL
        output Tile_X0Y4_B_config_C_bit0, //EXTERNAL
        output Tile_X0Y4_B_config_C_bit1, //EXTERNAL
        output Tile_X0Y4_B_config_C_bit2, //EXTERNAL
        output Tile_X0Y4_B_config_C_bit3, //EXTERNAL
        input Tile_X10Y4_CONFIGURED_top, //EXTERNAL
        input Tile_X10Y4_DOUT_SRAM0, //EXTERNAL
        input Tile_X10Y4_DOUT_SRAM1, //EXTERNAL
        input Tile_X10Y4_DOUT_SRAM2, //EXTERNAL
        input Tile_X10Y4_DOUT_SRAM3, //EXTERNAL
        input Tile_X10Y4_DOUT_SRAM4, //EXTERNAL
        input Tile_X10Y4_DOUT_SRAM5, //EXTERNAL
        input Tile_X10Y4_DOUT_SRAM6, //EXTERNAL
        input Tile_X10Y4_DOUT_SRAM7, //EXTERNAL
        input Tile_X10Y4_DOUT_SRAM8, //EXTERNAL
        input Tile_X10Y4_DOUT_SRAM9, //EXTERNAL
        input Tile_X10Y4_DOUT_SRAM10, //EXTERNAL
        input Tile_X10Y4_DOUT_SRAM11, //EXTERNAL
        input Tile_X10Y4_DOUT_SRAM12, //EXTERNAL
        input Tile_X10Y4_DOUT_SRAM13, //EXTERNAL
        input Tile_X10Y4_DOUT_SRAM14, //EXTERNAL
        input Tile_X10Y4_DOUT_SRAM15, //EXTERNAL
        input Tile_X10Y4_DOUT_SRAM16, //EXTERNAL
        input Tile_X10Y4_DOUT_SRAM17, //EXTERNAL
        input Tile_X10Y4_DOUT_SRAM18, //EXTERNAL
        input Tile_X10Y4_DOUT_SRAM19, //EXTERNAL
        input Tile_X10Y4_DOUT_SRAM20, //EXTERNAL
        input Tile_X10Y4_DOUT_SRAM21, //EXTERNAL
        input Tile_X10Y4_DOUT_SRAM22, //EXTERNAL
        input Tile_X10Y4_DOUT_SRAM23, //EXTERNAL
        input Tile_X10Y4_DOUT_SRAM24, //EXTERNAL
        input Tile_X10Y4_DOUT_SRAM25, //EXTERNAL
        input Tile_X10Y4_DOUT_SRAM26, //EXTERNAL
        input Tile_X10Y4_DOUT_SRAM27, //EXTERNAL
        input Tile_X10Y4_DOUT_SRAM28, //EXTERNAL
        input Tile_X10Y4_DOUT_SRAM29, //EXTERNAL
        input Tile_X10Y4_DOUT_SRAM30, //EXTERNAL
        input Tile_X10Y4_DOUT_SRAM31, //EXTERNAL
        output Tile_X10Y4_ADDR_SRAM0, //EXTERNAL
        output Tile_X10Y4_ADDR_SRAM1, //EXTERNAL
        output Tile_X10Y4_ADDR_SRAM2, //EXTERNAL
        output Tile_X10Y4_ADDR_SRAM3, //EXTERNAL
        output Tile_X10Y4_ADDR_SRAM4, //EXTERNAL
        output Tile_X10Y4_ADDR_SRAM5, //EXTERNAL
        output Tile_X10Y4_ADDR_SRAM6, //EXTERNAL
        output Tile_X10Y4_ADDR_SRAM7, //EXTERNAL
        output Tile_X10Y4_ADDR_SRAM8, //EXTERNAL
        output Tile_X10Y4_ADDR_SRAM9, //EXTERNAL
        output Tile_X10Y4_BM_SRAM0, //EXTERNAL
        output Tile_X10Y4_BM_SRAM1, //EXTERNAL
        output Tile_X10Y4_BM_SRAM2, //EXTERNAL
        output Tile_X10Y4_BM_SRAM3, //EXTERNAL
        output Tile_X10Y4_BM_SRAM4, //EXTERNAL
        output Tile_X10Y4_BM_SRAM5, //EXTERNAL
        output Tile_X10Y4_BM_SRAM6, //EXTERNAL
        output Tile_X10Y4_BM_SRAM7, //EXTERNAL
        output Tile_X10Y4_BM_SRAM8, //EXTERNAL
        output Tile_X10Y4_BM_SRAM9, //EXTERNAL
        output Tile_X10Y4_BM_SRAM10, //EXTERNAL
        output Tile_X10Y4_BM_SRAM11, //EXTERNAL
        output Tile_X10Y4_BM_SRAM12, //EXTERNAL
        output Tile_X10Y4_BM_SRAM13, //EXTERNAL
        output Tile_X10Y4_BM_SRAM14, //EXTERNAL
        output Tile_X10Y4_BM_SRAM15, //EXTERNAL
        output Tile_X10Y4_BM_SRAM16, //EXTERNAL
        output Tile_X10Y4_BM_SRAM17, //EXTERNAL
        output Tile_X10Y4_BM_SRAM18, //EXTERNAL
        output Tile_X10Y4_BM_SRAM19, //EXTERNAL
        output Tile_X10Y4_BM_SRAM20, //EXTERNAL
        output Tile_X10Y4_BM_SRAM21, //EXTERNAL
        output Tile_X10Y4_BM_SRAM22, //EXTERNAL
        output Tile_X10Y4_BM_SRAM23, //EXTERNAL
        output Tile_X10Y4_BM_SRAM24, //EXTERNAL
        output Tile_X10Y4_BM_SRAM25, //EXTERNAL
        output Tile_X10Y4_BM_SRAM26, //EXTERNAL
        output Tile_X10Y4_BM_SRAM27, //EXTERNAL
        output Tile_X10Y4_BM_SRAM28, //EXTERNAL
        output Tile_X10Y4_BM_SRAM29, //EXTERNAL
        output Tile_X10Y4_BM_SRAM30, //EXTERNAL
        output Tile_X10Y4_BM_SRAM31, //EXTERNAL
        output Tile_X10Y4_CLK_SRAM, //EXTERNAL
        output Tile_X10Y4_DIN_SRAM0, //EXTERNAL
        output Tile_X10Y4_DIN_SRAM1, //EXTERNAL
        output Tile_X10Y4_DIN_SRAM2, //EXTERNAL
        output Tile_X10Y4_DIN_SRAM3, //EXTERNAL
        output Tile_X10Y4_DIN_SRAM4, //EXTERNAL
        output Tile_X10Y4_DIN_SRAM5, //EXTERNAL
        output Tile_X10Y4_DIN_SRAM6, //EXTERNAL
        output Tile_X10Y4_DIN_SRAM7, //EXTERNAL
        output Tile_X10Y4_DIN_SRAM8, //EXTERNAL
        output Tile_X10Y4_DIN_SRAM9, //EXTERNAL
        output Tile_X10Y4_DIN_SRAM10, //EXTERNAL
        output Tile_X10Y4_DIN_SRAM11, //EXTERNAL
        output Tile_X10Y4_DIN_SRAM12, //EXTERNAL
        output Tile_X10Y4_DIN_SRAM13, //EXTERNAL
        output Tile_X10Y4_DIN_SRAM14, //EXTERNAL
        output Tile_X10Y4_DIN_SRAM15, //EXTERNAL
        output Tile_X10Y4_DIN_SRAM16, //EXTERNAL
        output Tile_X10Y4_DIN_SRAM17, //EXTERNAL
        output Tile_X10Y4_DIN_SRAM18, //EXTERNAL
        output Tile_X10Y4_DIN_SRAM19, //EXTERNAL
        output Tile_X10Y4_DIN_SRAM20, //EXTERNAL
        output Tile_X10Y4_DIN_SRAM21, //EXTERNAL
        output Tile_X10Y4_DIN_SRAM22, //EXTERNAL
        output Tile_X10Y4_DIN_SRAM23, //EXTERNAL
        output Tile_X10Y4_DIN_SRAM24, //EXTERNAL
        output Tile_X10Y4_DIN_SRAM25, //EXTERNAL
        output Tile_X10Y4_DIN_SRAM26, //EXTERNAL
        output Tile_X10Y4_DIN_SRAM27, //EXTERNAL
        output Tile_X10Y4_DIN_SRAM28, //EXTERNAL
        output Tile_X10Y4_DIN_SRAM29, //EXTERNAL
        output Tile_X10Y4_DIN_SRAM30, //EXTERNAL
        output Tile_X10Y4_DIN_SRAM31, //EXTERNAL
        output Tile_X10Y4_MEN_SRAM, //EXTERNAL
        output Tile_X10Y4_REN_SRAM, //EXTERNAL
        output Tile_X10Y4_TIE_HIGH_SRAM, //EXTERNAL
        output Tile_X10Y4_TIE_LOW_SRAM, //EXTERNAL
        output Tile_X10Y4_WEN_SRAM, //EXTERNAL
        input Tile_X0Y5_A_O_top, //EXTERNAL
        output Tile_X0Y5_A_I_top, //EXTERNAL
        output Tile_X0Y5_A_T_top, //EXTERNAL
        input Tile_X0Y5_B_O_top, //EXTERNAL
        output Tile_X0Y5_B_I_top, //EXTERNAL
        output Tile_X0Y5_B_T_top, //EXTERNAL
        output Tile_X0Y5_A_config_C_bit0, //EXTERNAL
        output Tile_X0Y5_A_config_C_bit1, //EXTERNAL
        output Tile_X0Y5_A_config_C_bit2, //EXTERNAL
        output Tile_X0Y5_A_config_C_bit3, //EXTERNAL
        output Tile_X0Y5_B_config_C_bit0, //EXTERNAL
        output Tile_X0Y5_B_config_C_bit1, //EXTERNAL
        output Tile_X0Y5_B_config_C_bit2, //EXTERNAL
        output Tile_X0Y5_B_config_C_bit3, //EXTERNAL
        input Tile_X0Y6_A_O_top, //EXTERNAL
        output Tile_X0Y6_A_I_top, //EXTERNAL
        output Tile_X0Y6_A_T_top, //EXTERNAL
        input Tile_X0Y6_B_O_top, //EXTERNAL
        output Tile_X0Y6_B_I_top, //EXTERNAL
        output Tile_X0Y6_B_T_top, //EXTERNAL
        output Tile_X0Y6_A_config_C_bit0, //EXTERNAL
        output Tile_X0Y6_A_config_C_bit1, //EXTERNAL
        output Tile_X0Y6_A_config_C_bit2, //EXTERNAL
        output Tile_X0Y6_A_config_C_bit3, //EXTERNAL
        output Tile_X0Y6_B_config_C_bit0, //EXTERNAL
        output Tile_X0Y6_B_config_C_bit1, //EXTERNAL
        output Tile_X0Y6_B_config_C_bit2, //EXTERNAL
        output Tile_X0Y6_B_config_C_bit3, //EXTERNAL
        input Tile_X10Y6_CONFIGURED_top, //EXTERNAL
        input Tile_X10Y6_DOUT_SRAM0, //EXTERNAL
        input Tile_X10Y6_DOUT_SRAM1, //EXTERNAL
        input Tile_X10Y6_DOUT_SRAM2, //EXTERNAL
        input Tile_X10Y6_DOUT_SRAM3, //EXTERNAL
        input Tile_X10Y6_DOUT_SRAM4, //EXTERNAL
        input Tile_X10Y6_DOUT_SRAM5, //EXTERNAL
        input Tile_X10Y6_DOUT_SRAM6, //EXTERNAL
        input Tile_X10Y6_DOUT_SRAM7, //EXTERNAL
        input Tile_X10Y6_DOUT_SRAM8, //EXTERNAL
        input Tile_X10Y6_DOUT_SRAM9, //EXTERNAL
        input Tile_X10Y6_DOUT_SRAM10, //EXTERNAL
        input Tile_X10Y6_DOUT_SRAM11, //EXTERNAL
        input Tile_X10Y6_DOUT_SRAM12, //EXTERNAL
        input Tile_X10Y6_DOUT_SRAM13, //EXTERNAL
        input Tile_X10Y6_DOUT_SRAM14, //EXTERNAL
        input Tile_X10Y6_DOUT_SRAM15, //EXTERNAL
        input Tile_X10Y6_DOUT_SRAM16, //EXTERNAL
        input Tile_X10Y6_DOUT_SRAM17, //EXTERNAL
        input Tile_X10Y6_DOUT_SRAM18, //EXTERNAL
        input Tile_X10Y6_DOUT_SRAM19, //EXTERNAL
        input Tile_X10Y6_DOUT_SRAM20, //EXTERNAL
        input Tile_X10Y6_DOUT_SRAM21, //EXTERNAL
        input Tile_X10Y6_DOUT_SRAM22, //EXTERNAL
        input Tile_X10Y6_DOUT_SRAM23, //EXTERNAL
        input Tile_X10Y6_DOUT_SRAM24, //EXTERNAL
        input Tile_X10Y6_DOUT_SRAM25, //EXTERNAL
        input Tile_X10Y6_DOUT_SRAM26, //EXTERNAL
        input Tile_X10Y6_DOUT_SRAM27, //EXTERNAL
        input Tile_X10Y6_DOUT_SRAM28, //EXTERNAL
        input Tile_X10Y6_DOUT_SRAM29, //EXTERNAL
        input Tile_X10Y6_DOUT_SRAM30, //EXTERNAL
        input Tile_X10Y6_DOUT_SRAM31, //EXTERNAL
        output Tile_X10Y6_ADDR_SRAM0, //EXTERNAL
        output Tile_X10Y6_ADDR_SRAM1, //EXTERNAL
        output Tile_X10Y6_ADDR_SRAM2, //EXTERNAL
        output Tile_X10Y6_ADDR_SRAM3, //EXTERNAL
        output Tile_X10Y6_ADDR_SRAM4, //EXTERNAL
        output Tile_X10Y6_ADDR_SRAM5, //EXTERNAL
        output Tile_X10Y6_ADDR_SRAM6, //EXTERNAL
        output Tile_X10Y6_ADDR_SRAM7, //EXTERNAL
        output Tile_X10Y6_ADDR_SRAM8, //EXTERNAL
        output Tile_X10Y6_ADDR_SRAM9, //EXTERNAL
        output Tile_X10Y6_BM_SRAM0, //EXTERNAL
        output Tile_X10Y6_BM_SRAM1, //EXTERNAL
        output Tile_X10Y6_BM_SRAM2, //EXTERNAL
        output Tile_X10Y6_BM_SRAM3, //EXTERNAL
        output Tile_X10Y6_BM_SRAM4, //EXTERNAL
        output Tile_X10Y6_BM_SRAM5, //EXTERNAL
        output Tile_X10Y6_BM_SRAM6, //EXTERNAL
        output Tile_X10Y6_BM_SRAM7, //EXTERNAL
        output Tile_X10Y6_BM_SRAM8, //EXTERNAL
        output Tile_X10Y6_BM_SRAM9, //EXTERNAL
        output Tile_X10Y6_BM_SRAM10, //EXTERNAL
        output Tile_X10Y6_BM_SRAM11, //EXTERNAL
        output Tile_X10Y6_BM_SRAM12, //EXTERNAL
        output Tile_X10Y6_BM_SRAM13, //EXTERNAL
        output Tile_X10Y6_BM_SRAM14, //EXTERNAL
        output Tile_X10Y6_BM_SRAM15, //EXTERNAL
        output Tile_X10Y6_BM_SRAM16, //EXTERNAL
        output Tile_X10Y6_BM_SRAM17, //EXTERNAL
        output Tile_X10Y6_BM_SRAM18, //EXTERNAL
        output Tile_X10Y6_BM_SRAM19, //EXTERNAL
        output Tile_X10Y6_BM_SRAM20, //EXTERNAL
        output Tile_X10Y6_BM_SRAM21, //EXTERNAL
        output Tile_X10Y6_BM_SRAM22, //EXTERNAL
        output Tile_X10Y6_BM_SRAM23, //EXTERNAL
        output Tile_X10Y6_BM_SRAM24, //EXTERNAL
        output Tile_X10Y6_BM_SRAM25, //EXTERNAL
        output Tile_X10Y6_BM_SRAM26, //EXTERNAL
        output Tile_X10Y6_BM_SRAM27, //EXTERNAL
        output Tile_X10Y6_BM_SRAM28, //EXTERNAL
        output Tile_X10Y6_BM_SRAM29, //EXTERNAL
        output Tile_X10Y6_BM_SRAM30, //EXTERNAL
        output Tile_X10Y6_BM_SRAM31, //EXTERNAL
        output Tile_X10Y6_CLK_SRAM, //EXTERNAL
        output Tile_X10Y6_DIN_SRAM0, //EXTERNAL
        output Tile_X10Y6_DIN_SRAM1, //EXTERNAL
        output Tile_X10Y6_DIN_SRAM2, //EXTERNAL
        output Tile_X10Y6_DIN_SRAM3, //EXTERNAL
        output Tile_X10Y6_DIN_SRAM4, //EXTERNAL
        output Tile_X10Y6_DIN_SRAM5, //EXTERNAL
        output Tile_X10Y6_DIN_SRAM6, //EXTERNAL
        output Tile_X10Y6_DIN_SRAM7, //EXTERNAL
        output Tile_X10Y6_DIN_SRAM8, //EXTERNAL
        output Tile_X10Y6_DIN_SRAM9, //EXTERNAL
        output Tile_X10Y6_DIN_SRAM10, //EXTERNAL
        output Tile_X10Y6_DIN_SRAM11, //EXTERNAL
        output Tile_X10Y6_DIN_SRAM12, //EXTERNAL
        output Tile_X10Y6_DIN_SRAM13, //EXTERNAL
        output Tile_X10Y6_DIN_SRAM14, //EXTERNAL
        output Tile_X10Y6_DIN_SRAM15, //EXTERNAL
        output Tile_X10Y6_DIN_SRAM16, //EXTERNAL
        output Tile_X10Y6_DIN_SRAM17, //EXTERNAL
        output Tile_X10Y6_DIN_SRAM18, //EXTERNAL
        output Tile_X10Y6_DIN_SRAM19, //EXTERNAL
        output Tile_X10Y6_DIN_SRAM20, //EXTERNAL
        output Tile_X10Y6_DIN_SRAM21, //EXTERNAL
        output Tile_X10Y6_DIN_SRAM22, //EXTERNAL
        output Tile_X10Y6_DIN_SRAM23, //EXTERNAL
        output Tile_X10Y6_DIN_SRAM24, //EXTERNAL
        output Tile_X10Y6_DIN_SRAM25, //EXTERNAL
        output Tile_X10Y6_DIN_SRAM26, //EXTERNAL
        output Tile_X10Y6_DIN_SRAM27, //EXTERNAL
        output Tile_X10Y6_DIN_SRAM28, //EXTERNAL
        output Tile_X10Y6_DIN_SRAM29, //EXTERNAL
        output Tile_X10Y6_DIN_SRAM30, //EXTERNAL
        output Tile_X10Y6_DIN_SRAM31, //EXTERNAL
        output Tile_X10Y6_MEN_SRAM, //EXTERNAL
        output Tile_X10Y6_REN_SRAM, //EXTERNAL
        output Tile_X10Y6_TIE_HIGH_SRAM, //EXTERNAL
        output Tile_X10Y6_TIE_LOW_SRAM, //EXTERNAL
        output Tile_X10Y6_WEN_SRAM, //EXTERNAL
        input Tile_X0Y7_A_O_top, //EXTERNAL
        output Tile_X0Y7_A_I_top, //EXTERNAL
        output Tile_X0Y7_A_T_top, //EXTERNAL
        input Tile_X0Y7_B_O_top, //EXTERNAL
        output Tile_X0Y7_B_I_top, //EXTERNAL
        output Tile_X0Y7_B_T_top, //EXTERNAL
        output Tile_X0Y7_A_config_C_bit0, //EXTERNAL
        output Tile_X0Y7_A_config_C_bit1, //EXTERNAL
        output Tile_X0Y7_A_config_C_bit2, //EXTERNAL
        output Tile_X0Y7_A_config_C_bit3, //EXTERNAL
        output Tile_X0Y7_B_config_C_bit0, //EXTERNAL
        output Tile_X0Y7_B_config_C_bit1, //EXTERNAL
        output Tile_X0Y7_B_config_C_bit2, //EXTERNAL
        output Tile_X0Y7_B_config_C_bit3, //EXTERNAL
        input Tile_X0Y8_A_O_top, //EXTERNAL
        output Tile_X0Y8_A_I_top, //EXTERNAL
        output Tile_X0Y8_A_T_top, //EXTERNAL
        input Tile_X0Y8_B_O_top, //EXTERNAL
        output Tile_X0Y8_B_I_top, //EXTERNAL
        output Tile_X0Y8_B_T_top, //EXTERNAL
        output Tile_X0Y8_A_config_C_bit0, //EXTERNAL
        output Tile_X0Y8_A_config_C_bit1, //EXTERNAL
        output Tile_X0Y8_A_config_C_bit2, //EXTERNAL
        output Tile_X0Y8_A_config_C_bit3, //EXTERNAL
        output Tile_X0Y8_B_config_C_bit0, //EXTERNAL
        output Tile_X0Y8_B_config_C_bit1, //EXTERNAL
        output Tile_X0Y8_B_config_C_bit2, //EXTERNAL
        output Tile_X0Y8_B_config_C_bit3, //EXTERNAL
        input Tile_X10Y8_CONFIGURED_top, //EXTERNAL
        input Tile_X10Y8_DOUT_SRAM0, //EXTERNAL
        input Tile_X10Y8_DOUT_SRAM1, //EXTERNAL
        input Tile_X10Y8_DOUT_SRAM2, //EXTERNAL
        input Tile_X10Y8_DOUT_SRAM3, //EXTERNAL
        input Tile_X10Y8_DOUT_SRAM4, //EXTERNAL
        input Tile_X10Y8_DOUT_SRAM5, //EXTERNAL
        input Tile_X10Y8_DOUT_SRAM6, //EXTERNAL
        input Tile_X10Y8_DOUT_SRAM7, //EXTERNAL
        input Tile_X10Y8_DOUT_SRAM8, //EXTERNAL
        input Tile_X10Y8_DOUT_SRAM9, //EXTERNAL
        input Tile_X10Y8_DOUT_SRAM10, //EXTERNAL
        input Tile_X10Y8_DOUT_SRAM11, //EXTERNAL
        input Tile_X10Y8_DOUT_SRAM12, //EXTERNAL
        input Tile_X10Y8_DOUT_SRAM13, //EXTERNAL
        input Tile_X10Y8_DOUT_SRAM14, //EXTERNAL
        input Tile_X10Y8_DOUT_SRAM15, //EXTERNAL
        input Tile_X10Y8_DOUT_SRAM16, //EXTERNAL
        input Tile_X10Y8_DOUT_SRAM17, //EXTERNAL
        input Tile_X10Y8_DOUT_SRAM18, //EXTERNAL
        input Tile_X10Y8_DOUT_SRAM19, //EXTERNAL
        input Tile_X10Y8_DOUT_SRAM20, //EXTERNAL
        input Tile_X10Y8_DOUT_SRAM21, //EXTERNAL
        input Tile_X10Y8_DOUT_SRAM22, //EXTERNAL
        input Tile_X10Y8_DOUT_SRAM23, //EXTERNAL
        input Tile_X10Y8_DOUT_SRAM24, //EXTERNAL
        input Tile_X10Y8_DOUT_SRAM25, //EXTERNAL
        input Tile_X10Y8_DOUT_SRAM26, //EXTERNAL
        input Tile_X10Y8_DOUT_SRAM27, //EXTERNAL
        input Tile_X10Y8_DOUT_SRAM28, //EXTERNAL
        input Tile_X10Y8_DOUT_SRAM29, //EXTERNAL
        input Tile_X10Y8_DOUT_SRAM30, //EXTERNAL
        input Tile_X10Y8_DOUT_SRAM31, //EXTERNAL
        output Tile_X10Y8_ADDR_SRAM0, //EXTERNAL
        output Tile_X10Y8_ADDR_SRAM1, //EXTERNAL
        output Tile_X10Y8_ADDR_SRAM2, //EXTERNAL
        output Tile_X10Y8_ADDR_SRAM3, //EXTERNAL
        output Tile_X10Y8_ADDR_SRAM4, //EXTERNAL
        output Tile_X10Y8_ADDR_SRAM5, //EXTERNAL
        output Tile_X10Y8_ADDR_SRAM6, //EXTERNAL
        output Tile_X10Y8_ADDR_SRAM7, //EXTERNAL
        output Tile_X10Y8_ADDR_SRAM8, //EXTERNAL
        output Tile_X10Y8_ADDR_SRAM9, //EXTERNAL
        output Tile_X10Y8_BM_SRAM0, //EXTERNAL
        output Tile_X10Y8_BM_SRAM1, //EXTERNAL
        output Tile_X10Y8_BM_SRAM2, //EXTERNAL
        output Tile_X10Y8_BM_SRAM3, //EXTERNAL
        output Tile_X10Y8_BM_SRAM4, //EXTERNAL
        output Tile_X10Y8_BM_SRAM5, //EXTERNAL
        output Tile_X10Y8_BM_SRAM6, //EXTERNAL
        output Tile_X10Y8_BM_SRAM7, //EXTERNAL
        output Tile_X10Y8_BM_SRAM8, //EXTERNAL
        output Tile_X10Y8_BM_SRAM9, //EXTERNAL
        output Tile_X10Y8_BM_SRAM10, //EXTERNAL
        output Tile_X10Y8_BM_SRAM11, //EXTERNAL
        output Tile_X10Y8_BM_SRAM12, //EXTERNAL
        output Tile_X10Y8_BM_SRAM13, //EXTERNAL
        output Tile_X10Y8_BM_SRAM14, //EXTERNAL
        output Tile_X10Y8_BM_SRAM15, //EXTERNAL
        output Tile_X10Y8_BM_SRAM16, //EXTERNAL
        output Tile_X10Y8_BM_SRAM17, //EXTERNAL
        output Tile_X10Y8_BM_SRAM18, //EXTERNAL
        output Tile_X10Y8_BM_SRAM19, //EXTERNAL
        output Tile_X10Y8_BM_SRAM20, //EXTERNAL
        output Tile_X10Y8_BM_SRAM21, //EXTERNAL
        output Tile_X10Y8_BM_SRAM22, //EXTERNAL
        output Tile_X10Y8_BM_SRAM23, //EXTERNAL
        output Tile_X10Y8_BM_SRAM24, //EXTERNAL
        output Tile_X10Y8_BM_SRAM25, //EXTERNAL
        output Tile_X10Y8_BM_SRAM26, //EXTERNAL
        output Tile_X10Y8_BM_SRAM27, //EXTERNAL
        output Tile_X10Y8_BM_SRAM28, //EXTERNAL
        output Tile_X10Y8_BM_SRAM29, //EXTERNAL
        output Tile_X10Y8_BM_SRAM30, //EXTERNAL
        output Tile_X10Y8_BM_SRAM31, //EXTERNAL
        output Tile_X10Y8_CLK_SRAM, //EXTERNAL
        output Tile_X10Y8_DIN_SRAM0, //EXTERNAL
        output Tile_X10Y8_DIN_SRAM1, //EXTERNAL
        output Tile_X10Y8_DIN_SRAM2, //EXTERNAL
        output Tile_X10Y8_DIN_SRAM3, //EXTERNAL
        output Tile_X10Y8_DIN_SRAM4, //EXTERNAL
        output Tile_X10Y8_DIN_SRAM5, //EXTERNAL
        output Tile_X10Y8_DIN_SRAM6, //EXTERNAL
        output Tile_X10Y8_DIN_SRAM7, //EXTERNAL
        output Tile_X10Y8_DIN_SRAM8, //EXTERNAL
        output Tile_X10Y8_DIN_SRAM9, //EXTERNAL
        output Tile_X10Y8_DIN_SRAM10, //EXTERNAL
        output Tile_X10Y8_DIN_SRAM11, //EXTERNAL
        output Tile_X10Y8_DIN_SRAM12, //EXTERNAL
        output Tile_X10Y8_DIN_SRAM13, //EXTERNAL
        output Tile_X10Y8_DIN_SRAM14, //EXTERNAL
        output Tile_X10Y8_DIN_SRAM15, //EXTERNAL
        output Tile_X10Y8_DIN_SRAM16, //EXTERNAL
        output Tile_X10Y8_DIN_SRAM17, //EXTERNAL
        output Tile_X10Y8_DIN_SRAM18, //EXTERNAL
        output Tile_X10Y8_DIN_SRAM19, //EXTERNAL
        output Tile_X10Y8_DIN_SRAM20, //EXTERNAL
        output Tile_X10Y8_DIN_SRAM21, //EXTERNAL
        output Tile_X10Y8_DIN_SRAM22, //EXTERNAL
        output Tile_X10Y8_DIN_SRAM23, //EXTERNAL
        output Tile_X10Y8_DIN_SRAM24, //EXTERNAL
        output Tile_X10Y8_DIN_SRAM25, //EXTERNAL
        output Tile_X10Y8_DIN_SRAM26, //EXTERNAL
        output Tile_X10Y8_DIN_SRAM27, //EXTERNAL
        output Tile_X10Y8_DIN_SRAM28, //EXTERNAL
        output Tile_X10Y8_DIN_SRAM29, //EXTERNAL
        output Tile_X10Y8_DIN_SRAM30, //EXTERNAL
        output Tile_X10Y8_DIN_SRAM31, //EXTERNAL
        output Tile_X10Y8_MEN_SRAM, //EXTERNAL
        output Tile_X10Y8_REN_SRAM, //EXTERNAL
        output Tile_X10Y8_TIE_HIGH_SRAM, //EXTERNAL
        output Tile_X10Y8_TIE_LOW_SRAM, //EXTERNAL
        output Tile_X10Y8_WEN_SRAM, //EXTERNAL
        input Tile_X0Y9_A_O_top, //EXTERNAL
        output Tile_X0Y9_A_I_top, //EXTERNAL
        output Tile_X0Y9_A_T_top, //EXTERNAL
        input Tile_X0Y9_B_O_top, //EXTERNAL
        output Tile_X0Y9_B_I_top, //EXTERNAL
        output Tile_X0Y9_B_T_top, //EXTERNAL
        output Tile_X0Y9_A_config_C_bit0, //EXTERNAL
        output Tile_X0Y9_A_config_C_bit1, //EXTERNAL
        output Tile_X0Y9_A_config_C_bit2, //EXTERNAL
        output Tile_X0Y9_A_config_C_bit3, //EXTERNAL
        output Tile_X0Y9_B_config_C_bit0, //EXTERNAL
        output Tile_X0Y9_B_config_C_bit1, //EXTERNAL
        output Tile_X0Y9_B_config_C_bit2, //EXTERNAL
        output Tile_X0Y9_B_config_C_bit3, //EXTERNAL
        input Tile_X0Y10_A_O_top, //EXTERNAL
        output Tile_X0Y10_A_I_top, //EXTERNAL
        output Tile_X0Y10_A_T_top, //EXTERNAL
        input Tile_X0Y10_B_O_top, //EXTERNAL
        output Tile_X0Y10_B_I_top, //EXTERNAL
        output Tile_X0Y10_B_T_top, //EXTERNAL
        output Tile_X0Y10_A_config_C_bit0, //EXTERNAL
        output Tile_X0Y10_A_config_C_bit1, //EXTERNAL
        output Tile_X0Y10_A_config_C_bit2, //EXTERNAL
        output Tile_X0Y10_A_config_C_bit3, //EXTERNAL
        output Tile_X0Y10_B_config_C_bit0, //EXTERNAL
        output Tile_X0Y10_B_config_C_bit1, //EXTERNAL
        output Tile_X0Y10_B_config_C_bit2, //EXTERNAL
        output Tile_X0Y10_B_config_C_bit3, //EXTERNAL
        input Tile_X10Y10_CONFIGURED_top, //EXTERNAL
        input Tile_X10Y10_DOUT_SRAM0, //EXTERNAL
        input Tile_X10Y10_DOUT_SRAM1, //EXTERNAL
        input Tile_X10Y10_DOUT_SRAM2, //EXTERNAL
        input Tile_X10Y10_DOUT_SRAM3, //EXTERNAL
        input Tile_X10Y10_DOUT_SRAM4, //EXTERNAL
        input Tile_X10Y10_DOUT_SRAM5, //EXTERNAL
        input Tile_X10Y10_DOUT_SRAM6, //EXTERNAL
        input Tile_X10Y10_DOUT_SRAM7, //EXTERNAL
        input Tile_X10Y10_DOUT_SRAM8, //EXTERNAL
        input Tile_X10Y10_DOUT_SRAM9, //EXTERNAL
        input Tile_X10Y10_DOUT_SRAM10, //EXTERNAL
        input Tile_X10Y10_DOUT_SRAM11, //EXTERNAL
        input Tile_X10Y10_DOUT_SRAM12, //EXTERNAL
        input Tile_X10Y10_DOUT_SRAM13, //EXTERNAL
        input Tile_X10Y10_DOUT_SRAM14, //EXTERNAL
        input Tile_X10Y10_DOUT_SRAM15, //EXTERNAL
        input Tile_X10Y10_DOUT_SRAM16, //EXTERNAL
        input Tile_X10Y10_DOUT_SRAM17, //EXTERNAL
        input Tile_X10Y10_DOUT_SRAM18, //EXTERNAL
        input Tile_X10Y10_DOUT_SRAM19, //EXTERNAL
        input Tile_X10Y10_DOUT_SRAM20, //EXTERNAL
        input Tile_X10Y10_DOUT_SRAM21, //EXTERNAL
        input Tile_X10Y10_DOUT_SRAM22, //EXTERNAL
        input Tile_X10Y10_DOUT_SRAM23, //EXTERNAL
        input Tile_X10Y10_DOUT_SRAM24, //EXTERNAL
        input Tile_X10Y10_DOUT_SRAM25, //EXTERNAL
        input Tile_X10Y10_DOUT_SRAM26, //EXTERNAL
        input Tile_X10Y10_DOUT_SRAM27, //EXTERNAL
        input Tile_X10Y10_DOUT_SRAM28, //EXTERNAL
        input Tile_X10Y10_DOUT_SRAM29, //EXTERNAL
        input Tile_X10Y10_DOUT_SRAM30, //EXTERNAL
        input Tile_X10Y10_DOUT_SRAM31, //EXTERNAL
        output Tile_X10Y10_ADDR_SRAM0, //EXTERNAL
        output Tile_X10Y10_ADDR_SRAM1, //EXTERNAL
        output Tile_X10Y10_ADDR_SRAM2, //EXTERNAL
        output Tile_X10Y10_ADDR_SRAM3, //EXTERNAL
        output Tile_X10Y10_ADDR_SRAM4, //EXTERNAL
        output Tile_X10Y10_ADDR_SRAM5, //EXTERNAL
        output Tile_X10Y10_ADDR_SRAM6, //EXTERNAL
        output Tile_X10Y10_ADDR_SRAM7, //EXTERNAL
        output Tile_X10Y10_ADDR_SRAM8, //EXTERNAL
        output Tile_X10Y10_ADDR_SRAM9, //EXTERNAL
        output Tile_X10Y10_BM_SRAM0, //EXTERNAL
        output Tile_X10Y10_BM_SRAM1, //EXTERNAL
        output Tile_X10Y10_BM_SRAM2, //EXTERNAL
        output Tile_X10Y10_BM_SRAM3, //EXTERNAL
        output Tile_X10Y10_BM_SRAM4, //EXTERNAL
        output Tile_X10Y10_BM_SRAM5, //EXTERNAL
        output Tile_X10Y10_BM_SRAM6, //EXTERNAL
        output Tile_X10Y10_BM_SRAM7, //EXTERNAL
        output Tile_X10Y10_BM_SRAM8, //EXTERNAL
        output Tile_X10Y10_BM_SRAM9, //EXTERNAL
        output Tile_X10Y10_BM_SRAM10, //EXTERNAL
        output Tile_X10Y10_BM_SRAM11, //EXTERNAL
        output Tile_X10Y10_BM_SRAM12, //EXTERNAL
        output Tile_X10Y10_BM_SRAM13, //EXTERNAL
        output Tile_X10Y10_BM_SRAM14, //EXTERNAL
        output Tile_X10Y10_BM_SRAM15, //EXTERNAL
        output Tile_X10Y10_BM_SRAM16, //EXTERNAL
        output Tile_X10Y10_BM_SRAM17, //EXTERNAL
        output Tile_X10Y10_BM_SRAM18, //EXTERNAL
        output Tile_X10Y10_BM_SRAM19, //EXTERNAL
        output Tile_X10Y10_BM_SRAM20, //EXTERNAL
        output Tile_X10Y10_BM_SRAM21, //EXTERNAL
        output Tile_X10Y10_BM_SRAM22, //EXTERNAL
        output Tile_X10Y10_BM_SRAM23, //EXTERNAL
        output Tile_X10Y10_BM_SRAM24, //EXTERNAL
        output Tile_X10Y10_BM_SRAM25, //EXTERNAL
        output Tile_X10Y10_BM_SRAM26, //EXTERNAL
        output Tile_X10Y10_BM_SRAM27, //EXTERNAL
        output Tile_X10Y10_BM_SRAM28, //EXTERNAL
        output Tile_X10Y10_BM_SRAM29, //EXTERNAL
        output Tile_X10Y10_BM_SRAM30, //EXTERNAL
        output Tile_X10Y10_BM_SRAM31, //EXTERNAL
        output Tile_X10Y10_CLK_SRAM, //EXTERNAL
        output Tile_X10Y10_DIN_SRAM0, //EXTERNAL
        output Tile_X10Y10_DIN_SRAM1, //EXTERNAL
        output Tile_X10Y10_DIN_SRAM2, //EXTERNAL
        output Tile_X10Y10_DIN_SRAM3, //EXTERNAL
        output Tile_X10Y10_DIN_SRAM4, //EXTERNAL
        output Tile_X10Y10_DIN_SRAM5, //EXTERNAL
        output Tile_X10Y10_DIN_SRAM6, //EXTERNAL
        output Tile_X10Y10_DIN_SRAM7, //EXTERNAL
        output Tile_X10Y10_DIN_SRAM8, //EXTERNAL
        output Tile_X10Y10_DIN_SRAM9, //EXTERNAL
        output Tile_X10Y10_DIN_SRAM10, //EXTERNAL
        output Tile_X10Y10_DIN_SRAM11, //EXTERNAL
        output Tile_X10Y10_DIN_SRAM12, //EXTERNAL
        output Tile_X10Y10_DIN_SRAM13, //EXTERNAL
        output Tile_X10Y10_DIN_SRAM14, //EXTERNAL
        output Tile_X10Y10_DIN_SRAM15, //EXTERNAL
        output Tile_X10Y10_DIN_SRAM16, //EXTERNAL
        output Tile_X10Y10_DIN_SRAM17, //EXTERNAL
        output Tile_X10Y10_DIN_SRAM18, //EXTERNAL
        output Tile_X10Y10_DIN_SRAM19, //EXTERNAL
        output Tile_X10Y10_DIN_SRAM20, //EXTERNAL
        output Tile_X10Y10_DIN_SRAM21, //EXTERNAL
        output Tile_X10Y10_DIN_SRAM22, //EXTERNAL
        output Tile_X10Y10_DIN_SRAM23, //EXTERNAL
        output Tile_X10Y10_DIN_SRAM24, //EXTERNAL
        output Tile_X10Y10_DIN_SRAM25, //EXTERNAL
        output Tile_X10Y10_DIN_SRAM26, //EXTERNAL
        output Tile_X10Y10_DIN_SRAM27, //EXTERNAL
        output Tile_X10Y10_DIN_SRAM28, //EXTERNAL
        output Tile_X10Y10_DIN_SRAM29, //EXTERNAL
        output Tile_X10Y10_DIN_SRAM30, //EXTERNAL
        output Tile_X10Y10_DIN_SRAM31, //EXTERNAL
        output Tile_X10Y10_MEN_SRAM, //EXTERNAL
        output Tile_X10Y10_REN_SRAM, //EXTERNAL
        output Tile_X10Y10_TIE_HIGH_SRAM, //EXTERNAL
        output Tile_X10Y10_TIE_LOW_SRAM, //EXTERNAL
        output Tile_X10Y10_WEN_SRAM, //EXTERNAL
        input Tile_X0Y11_A_O_top, //EXTERNAL
        output Tile_X0Y11_A_I_top, //EXTERNAL
        output Tile_X0Y11_A_T_top, //EXTERNAL
        input Tile_X0Y11_B_O_top, //EXTERNAL
        output Tile_X0Y11_B_I_top, //EXTERNAL
        output Tile_X0Y11_B_T_top, //EXTERNAL
        output Tile_X0Y11_A_config_C_bit0, //EXTERNAL
        output Tile_X0Y11_A_config_C_bit1, //EXTERNAL
        output Tile_X0Y11_A_config_C_bit2, //EXTERNAL
        output Tile_X0Y11_A_config_C_bit3, //EXTERNAL
        output Tile_X0Y11_B_config_C_bit0, //EXTERNAL
        output Tile_X0Y11_B_config_C_bit1, //EXTERNAL
        output Tile_X0Y11_B_config_C_bit2, //EXTERNAL
        output Tile_X0Y11_B_config_C_bit3, //EXTERNAL
        input Tile_X0Y12_A_O_top, //EXTERNAL
        output Tile_X0Y12_A_I_top, //EXTERNAL
        output Tile_X0Y12_A_T_top, //EXTERNAL
        input Tile_X0Y12_B_O_top, //EXTERNAL
        output Tile_X0Y12_B_I_top, //EXTERNAL
        output Tile_X0Y12_B_T_top, //EXTERNAL
        output Tile_X0Y12_A_config_C_bit0, //EXTERNAL
        output Tile_X0Y12_A_config_C_bit1, //EXTERNAL
        output Tile_X0Y12_A_config_C_bit2, //EXTERNAL
        output Tile_X0Y12_A_config_C_bit3, //EXTERNAL
        output Tile_X0Y12_B_config_C_bit0, //EXTERNAL
        output Tile_X0Y12_B_config_C_bit1, //EXTERNAL
        output Tile_X0Y12_B_config_C_bit2, //EXTERNAL
        output Tile_X0Y12_B_config_C_bit3, //EXTERNAL
        input Tile_X10Y12_CONFIGURED_top, //EXTERNAL
        input Tile_X10Y12_DOUT_SRAM0, //EXTERNAL
        input Tile_X10Y12_DOUT_SRAM1, //EXTERNAL
        input Tile_X10Y12_DOUT_SRAM2, //EXTERNAL
        input Tile_X10Y12_DOUT_SRAM3, //EXTERNAL
        input Tile_X10Y12_DOUT_SRAM4, //EXTERNAL
        input Tile_X10Y12_DOUT_SRAM5, //EXTERNAL
        input Tile_X10Y12_DOUT_SRAM6, //EXTERNAL
        input Tile_X10Y12_DOUT_SRAM7, //EXTERNAL
        input Tile_X10Y12_DOUT_SRAM8, //EXTERNAL
        input Tile_X10Y12_DOUT_SRAM9, //EXTERNAL
        input Tile_X10Y12_DOUT_SRAM10, //EXTERNAL
        input Tile_X10Y12_DOUT_SRAM11, //EXTERNAL
        input Tile_X10Y12_DOUT_SRAM12, //EXTERNAL
        input Tile_X10Y12_DOUT_SRAM13, //EXTERNAL
        input Tile_X10Y12_DOUT_SRAM14, //EXTERNAL
        input Tile_X10Y12_DOUT_SRAM15, //EXTERNAL
        input Tile_X10Y12_DOUT_SRAM16, //EXTERNAL
        input Tile_X10Y12_DOUT_SRAM17, //EXTERNAL
        input Tile_X10Y12_DOUT_SRAM18, //EXTERNAL
        input Tile_X10Y12_DOUT_SRAM19, //EXTERNAL
        input Tile_X10Y12_DOUT_SRAM20, //EXTERNAL
        input Tile_X10Y12_DOUT_SRAM21, //EXTERNAL
        input Tile_X10Y12_DOUT_SRAM22, //EXTERNAL
        input Tile_X10Y12_DOUT_SRAM23, //EXTERNAL
        input Tile_X10Y12_DOUT_SRAM24, //EXTERNAL
        input Tile_X10Y12_DOUT_SRAM25, //EXTERNAL
        input Tile_X10Y12_DOUT_SRAM26, //EXTERNAL
        input Tile_X10Y12_DOUT_SRAM27, //EXTERNAL
        input Tile_X10Y12_DOUT_SRAM28, //EXTERNAL
        input Tile_X10Y12_DOUT_SRAM29, //EXTERNAL
        input Tile_X10Y12_DOUT_SRAM30, //EXTERNAL
        input Tile_X10Y12_DOUT_SRAM31, //EXTERNAL
        output Tile_X10Y12_ADDR_SRAM0, //EXTERNAL
        output Tile_X10Y12_ADDR_SRAM1, //EXTERNAL
        output Tile_X10Y12_ADDR_SRAM2, //EXTERNAL
        output Tile_X10Y12_ADDR_SRAM3, //EXTERNAL
        output Tile_X10Y12_ADDR_SRAM4, //EXTERNAL
        output Tile_X10Y12_ADDR_SRAM5, //EXTERNAL
        output Tile_X10Y12_ADDR_SRAM6, //EXTERNAL
        output Tile_X10Y12_ADDR_SRAM7, //EXTERNAL
        output Tile_X10Y12_ADDR_SRAM8, //EXTERNAL
        output Tile_X10Y12_ADDR_SRAM9, //EXTERNAL
        output Tile_X10Y12_BM_SRAM0, //EXTERNAL
        output Tile_X10Y12_BM_SRAM1, //EXTERNAL
        output Tile_X10Y12_BM_SRAM2, //EXTERNAL
        output Tile_X10Y12_BM_SRAM3, //EXTERNAL
        output Tile_X10Y12_BM_SRAM4, //EXTERNAL
        output Tile_X10Y12_BM_SRAM5, //EXTERNAL
        output Tile_X10Y12_BM_SRAM6, //EXTERNAL
        output Tile_X10Y12_BM_SRAM7, //EXTERNAL
        output Tile_X10Y12_BM_SRAM8, //EXTERNAL
        output Tile_X10Y12_BM_SRAM9, //EXTERNAL
        output Tile_X10Y12_BM_SRAM10, //EXTERNAL
        output Tile_X10Y12_BM_SRAM11, //EXTERNAL
        output Tile_X10Y12_BM_SRAM12, //EXTERNAL
        output Tile_X10Y12_BM_SRAM13, //EXTERNAL
        output Tile_X10Y12_BM_SRAM14, //EXTERNAL
        output Tile_X10Y12_BM_SRAM15, //EXTERNAL
        output Tile_X10Y12_BM_SRAM16, //EXTERNAL
        output Tile_X10Y12_BM_SRAM17, //EXTERNAL
        output Tile_X10Y12_BM_SRAM18, //EXTERNAL
        output Tile_X10Y12_BM_SRAM19, //EXTERNAL
        output Tile_X10Y12_BM_SRAM20, //EXTERNAL
        output Tile_X10Y12_BM_SRAM21, //EXTERNAL
        output Tile_X10Y12_BM_SRAM22, //EXTERNAL
        output Tile_X10Y12_BM_SRAM23, //EXTERNAL
        output Tile_X10Y12_BM_SRAM24, //EXTERNAL
        output Tile_X10Y12_BM_SRAM25, //EXTERNAL
        output Tile_X10Y12_BM_SRAM26, //EXTERNAL
        output Tile_X10Y12_BM_SRAM27, //EXTERNAL
        output Tile_X10Y12_BM_SRAM28, //EXTERNAL
        output Tile_X10Y12_BM_SRAM29, //EXTERNAL
        output Tile_X10Y12_BM_SRAM30, //EXTERNAL
        output Tile_X10Y12_BM_SRAM31, //EXTERNAL
        output Tile_X10Y12_CLK_SRAM, //EXTERNAL
        output Tile_X10Y12_DIN_SRAM0, //EXTERNAL
        output Tile_X10Y12_DIN_SRAM1, //EXTERNAL
        output Tile_X10Y12_DIN_SRAM2, //EXTERNAL
        output Tile_X10Y12_DIN_SRAM3, //EXTERNAL
        output Tile_X10Y12_DIN_SRAM4, //EXTERNAL
        output Tile_X10Y12_DIN_SRAM5, //EXTERNAL
        output Tile_X10Y12_DIN_SRAM6, //EXTERNAL
        output Tile_X10Y12_DIN_SRAM7, //EXTERNAL
        output Tile_X10Y12_DIN_SRAM8, //EXTERNAL
        output Tile_X10Y12_DIN_SRAM9, //EXTERNAL
        output Tile_X10Y12_DIN_SRAM10, //EXTERNAL
        output Tile_X10Y12_DIN_SRAM11, //EXTERNAL
        output Tile_X10Y12_DIN_SRAM12, //EXTERNAL
        output Tile_X10Y12_DIN_SRAM13, //EXTERNAL
        output Tile_X10Y12_DIN_SRAM14, //EXTERNAL
        output Tile_X10Y12_DIN_SRAM15, //EXTERNAL
        output Tile_X10Y12_DIN_SRAM16, //EXTERNAL
        output Tile_X10Y12_DIN_SRAM17, //EXTERNAL
        output Tile_X10Y12_DIN_SRAM18, //EXTERNAL
        output Tile_X10Y12_DIN_SRAM19, //EXTERNAL
        output Tile_X10Y12_DIN_SRAM20, //EXTERNAL
        output Tile_X10Y12_DIN_SRAM21, //EXTERNAL
        output Tile_X10Y12_DIN_SRAM22, //EXTERNAL
        output Tile_X10Y12_DIN_SRAM23, //EXTERNAL
        output Tile_X10Y12_DIN_SRAM24, //EXTERNAL
        output Tile_X10Y12_DIN_SRAM25, //EXTERNAL
        output Tile_X10Y12_DIN_SRAM26, //EXTERNAL
        output Tile_X10Y12_DIN_SRAM27, //EXTERNAL
        output Tile_X10Y12_DIN_SRAM28, //EXTERNAL
        output Tile_X10Y12_DIN_SRAM29, //EXTERNAL
        output Tile_X10Y12_DIN_SRAM30, //EXTERNAL
        output Tile_X10Y12_DIN_SRAM31, //EXTERNAL
        output Tile_X10Y12_MEN_SRAM, //EXTERNAL
        output Tile_X10Y12_REN_SRAM, //EXTERNAL
        output Tile_X10Y12_TIE_HIGH_SRAM, //EXTERNAL
        output Tile_X10Y12_TIE_LOW_SRAM, //EXTERNAL
        output Tile_X10Y12_WEN_SRAM, //EXTERNAL
        input Tile_X0Y13_A_O_top, //EXTERNAL
        output Tile_X0Y13_A_I_top, //EXTERNAL
        output Tile_X0Y13_A_T_top, //EXTERNAL
        input Tile_X0Y13_B_O_top, //EXTERNAL
        output Tile_X0Y13_B_I_top, //EXTERNAL
        output Tile_X0Y13_B_T_top, //EXTERNAL
        output Tile_X0Y13_A_config_C_bit0, //EXTERNAL
        output Tile_X0Y13_A_config_C_bit1, //EXTERNAL
        output Tile_X0Y13_A_config_C_bit2, //EXTERNAL
        output Tile_X0Y13_A_config_C_bit3, //EXTERNAL
        output Tile_X0Y13_B_config_C_bit0, //EXTERNAL
        output Tile_X0Y13_B_config_C_bit1, //EXTERNAL
        output Tile_X0Y13_B_config_C_bit2, //EXTERNAL
        output Tile_X0Y13_B_config_C_bit3, //EXTERNAL
        input Tile_X0Y14_A_O_top, //EXTERNAL
        output Tile_X0Y14_A_I_top, //EXTERNAL
        output Tile_X0Y14_A_T_top, //EXTERNAL
        input Tile_X0Y14_B_O_top, //EXTERNAL
        output Tile_X0Y14_B_I_top, //EXTERNAL
        output Tile_X0Y14_B_T_top, //EXTERNAL
        output Tile_X0Y14_A_config_C_bit0, //EXTERNAL
        output Tile_X0Y14_A_config_C_bit1, //EXTERNAL
        output Tile_X0Y14_A_config_C_bit2, //EXTERNAL
        output Tile_X0Y14_A_config_C_bit3, //EXTERNAL
        output Tile_X0Y14_B_config_C_bit0, //EXTERNAL
        output Tile_X0Y14_B_config_C_bit1, //EXTERNAL
        output Tile_X0Y14_B_config_C_bit2, //EXTERNAL
        output Tile_X0Y14_B_config_C_bit3, //EXTERNAL
        input Tile_X10Y14_CONFIGURED_top, //EXTERNAL
        input Tile_X10Y14_DOUT_SRAM0, //EXTERNAL
        input Tile_X10Y14_DOUT_SRAM1, //EXTERNAL
        input Tile_X10Y14_DOUT_SRAM2, //EXTERNAL
        input Tile_X10Y14_DOUT_SRAM3, //EXTERNAL
        input Tile_X10Y14_DOUT_SRAM4, //EXTERNAL
        input Tile_X10Y14_DOUT_SRAM5, //EXTERNAL
        input Tile_X10Y14_DOUT_SRAM6, //EXTERNAL
        input Tile_X10Y14_DOUT_SRAM7, //EXTERNAL
        input Tile_X10Y14_DOUT_SRAM8, //EXTERNAL
        input Tile_X10Y14_DOUT_SRAM9, //EXTERNAL
        input Tile_X10Y14_DOUT_SRAM10, //EXTERNAL
        input Tile_X10Y14_DOUT_SRAM11, //EXTERNAL
        input Tile_X10Y14_DOUT_SRAM12, //EXTERNAL
        input Tile_X10Y14_DOUT_SRAM13, //EXTERNAL
        input Tile_X10Y14_DOUT_SRAM14, //EXTERNAL
        input Tile_X10Y14_DOUT_SRAM15, //EXTERNAL
        input Tile_X10Y14_DOUT_SRAM16, //EXTERNAL
        input Tile_X10Y14_DOUT_SRAM17, //EXTERNAL
        input Tile_X10Y14_DOUT_SRAM18, //EXTERNAL
        input Tile_X10Y14_DOUT_SRAM19, //EXTERNAL
        input Tile_X10Y14_DOUT_SRAM20, //EXTERNAL
        input Tile_X10Y14_DOUT_SRAM21, //EXTERNAL
        input Tile_X10Y14_DOUT_SRAM22, //EXTERNAL
        input Tile_X10Y14_DOUT_SRAM23, //EXTERNAL
        input Tile_X10Y14_DOUT_SRAM24, //EXTERNAL
        input Tile_X10Y14_DOUT_SRAM25, //EXTERNAL
        input Tile_X10Y14_DOUT_SRAM26, //EXTERNAL
        input Tile_X10Y14_DOUT_SRAM27, //EXTERNAL
        input Tile_X10Y14_DOUT_SRAM28, //EXTERNAL
        input Tile_X10Y14_DOUT_SRAM29, //EXTERNAL
        input Tile_X10Y14_DOUT_SRAM30, //EXTERNAL
        input Tile_X10Y14_DOUT_SRAM31, //EXTERNAL
        output Tile_X10Y14_ADDR_SRAM0, //EXTERNAL
        output Tile_X10Y14_ADDR_SRAM1, //EXTERNAL
        output Tile_X10Y14_ADDR_SRAM2, //EXTERNAL
        output Tile_X10Y14_ADDR_SRAM3, //EXTERNAL
        output Tile_X10Y14_ADDR_SRAM4, //EXTERNAL
        output Tile_X10Y14_ADDR_SRAM5, //EXTERNAL
        output Tile_X10Y14_ADDR_SRAM6, //EXTERNAL
        output Tile_X10Y14_ADDR_SRAM7, //EXTERNAL
        output Tile_X10Y14_ADDR_SRAM8, //EXTERNAL
        output Tile_X10Y14_ADDR_SRAM9, //EXTERNAL
        output Tile_X10Y14_BM_SRAM0, //EXTERNAL
        output Tile_X10Y14_BM_SRAM1, //EXTERNAL
        output Tile_X10Y14_BM_SRAM2, //EXTERNAL
        output Tile_X10Y14_BM_SRAM3, //EXTERNAL
        output Tile_X10Y14_BM_SRAM4, //EXTERNAL
        output Tile_X10Y14_BM_SRAM5, //EXTERNAL
        output Tile_X10Y14_BM_SRAM6, //EXTERNAL
        output Tile_X10Y14_BM_SRAM7, //EXTERNAL
        output Tile_X10Y14_BM_SRAM8, //EXTERNAL
        output Tile_X10Y14_BM_SRAM9, //EXTERNAL
        output Tile_X10Y14_BM_SRAM10, //EXTERNAL
        output Tile_X10Y14_BM_SRAM11, //EXTERNAL
        output Tile_X10Y14_BM_SRAM12, //EXTERNAL
        output Tile_X10Y14_BM_SRAM13, //EXTERNAL
        output Tile_X10Y14_BM_SRAM14, //EXTERNAL
        output Tile_X10Y14_BM_SRAM15, //EXTERNAL
        output Tile_X10Y14_BM_SRAM16, //EXTERNAL
        output Tile_X10Y14_BM_SRAM17, //EXTERNAL
        output Tile_X10Y14_BM_SRAM18, //EXTERNAL
        output Tile_X10Y14_BM_SRAM19, //EXTERNAL
        output Tile_X10Y14_BM_SRAM20, //EXTERNAL
        output Tile_X10Y14_BM_SRAM21, //EXTERNAL
        output Tile_X10Y14_BM_SRAM22, //EXTERNAL
        output Tile_X10Y14_BM_SRAM23, //EXTERNAL
        output Tile_X10Y14_BM_SRAM24, //EXTERNAL
        output Tile_X10Y14_BM_SRAM25, //EXTERNAL
        output Tile_X10Y14_BM_SRAM26, //EXTERNAL
        output Tile_X10Y14_BM_SRAM27, //EXTERNAL
        output Tile_X10Y14_BM_SRAM28, //EXTERNAL
        output Tile_X10Y14_BM_SRAM29, //EXTERNAL
        output Tile_X10Y14_BM_SRAM30, //EXTERNAL
        output Tile_X10Y14_BM_SRAM31, //EXTERNAL
        output Tile_X10Y14_CLK_SRAM, //EXTERNAL
        output Tile_X10Y14_DIN_SRAM0, //EXTERNAL
        output Tile_X10Y14_DIN_SRAM1, //EXTERNAL
        output Tile_X10Y14_DIN_SRAM2, //EXTERNAL
        output Tile_X10Y14_DIN_SRAM3, //EXTERNAL
        output Tile_X10Y14_DIN_SRAM4, //EXTERNAL
        output Tile_X10Y14_DIN_SRAM5, //EXTERNAL
        output Tile_X10Y14_DIN_SRAM6, //EXTERNAL
        output Tile_X10Y14_DIN_SRAM7, //EXTERNAL
        output Tile_X10Y14_DIN_SRAM8, //EXTERNAL
        output Tile_X10Y14_DIN_SRAM9, //EXTERNAL
        output Tile_X10Y14_DIN_SRAM10, //EXTERNAL
        output Tile_X10Y14_DIN_SRAM11, //EXTERNAL
        output Tile_X10Y14_DIN_SRAM12, //EXTERNAL
        output Tile_X10Y14_DIN_SRAM13, //EXTERNAL
        output Tile_X10Y14_DIN_SRAM14, //EXTERNAL
        output Tile_X10Y14_DIN_SRAM15, //EXTERNAL
        output Tile_X10Y14_DIN_SRAM16, //EXTERNAL
        output Tile_X10Y14_DIN_SRAM17, //EXTERNAL
        output Tile_X10Y14_DIN_SRAM18, //EXTERNAL
        output Tile_X10Y14_DIN_SRAM19, //EXTERNAL
        output Tile_X10Y14_DIN_SRAM20, //EXTERNAL
        output Tile_X10Y14_DIN_SRAM21, //EXTERNAL
        output Tile_X10Y14_DIN_SRAM22, //EXTERNAL
        output Tile_X10Y14_DIN_SRAM23, //EXTERNAL
        output Tile_X10Y14_DIN_SRAM24, //EXTERNAL
        output Tile_X10Y14_DIN_SRAM25, //EXTERNAL
        output Tile_X10Y14_DIN_SRAM26, //EXTERNAL
        output Tile_X10Y14_DIN_SRAM27, //EXTERNAL
        output Tile_X10Y14_DIN_SRAM28, //EXTERNAL
        output Tile_X10Y14_DIN_SRAM29, //EXTERNAL
        output Tile_X10Y14_DIN_SRAM30, //EXTERNAL
        output Tile_X10Y14_DIN_SRAM31, //EXTERNAL
        output Tile_X10Y14_MEN_SRAM, //EXTERNAL
        output Tile_X10Y14_REN_SRAM, //EXTERNAL
        output Tile_X10Y14_TIE_HIGH_SRAM, //EXTERNAL
        output Tile_X10Y14_TIE_LOW_SRAM, //EXTERNAL
        output Tile_X10Y14_WEN_SRAM, //EXTERNAL
        input Tile_X2Y15_CONFIGURED_top, //EXTERNAL
        input Tile_X2Y15_RESET_top, //EXTERNAL
        output Tile_X2Y15_BOOT_top, //EXTERNAL
        output Tile_X2Y15_SLOT_top0, //EXTERNAL
        output Tile_X2Y15_SLOT_top1, //EXTERNAL
        output Tile_X2Y15_SLOT_top2, //EXTERNAL
        output Tile_X2Y15_SLOT_top3, //EXTERNAL
        input Tile_X3Y15_CONFIGURED_top, //EXTERNAL
        output Tile_X3Y15_IRQ_top0, //EXTERNAL
        output Tile_X3Y15_IRQ_top1, //EXTERNAL
        output Tile_X3Y15_IRQ_top2, //EXTERNAL
        output Tile_X3Y15_IRQ_top3, //EXTERNAL
        input Tile_X5Y15_O_top0, //EXTERNAL
        input Tile_X5Y15_O_top1, //EXTERNAL
        input Tile_X5Y15_O_top2, //EXTERNAL
        input Tile_X5Y15_O_top3, //EXTERNAL
        input Tile_X5Y15_O_top4, //EXTERNAL
        input Tile_X5Y15_O_top5, //EXTERNAL
        input Tile_X5Y15_O_top6, //EXTERNAL
        input Tile_X5Y15_O_top7, //EXTERNAL
        input Tile_X5Y15_O_top8, //EXTERNAL
        input Tile_X5Y15_O_top9, //EXTERNAL
        input Tile_X5Y15_O_top10, //EXTERNAL
        input Tile_X5Y15_O_top11, //EXTERNAL
        input Tile_X5Y15_O_top12, //EXTERNAL
        input Tile_X5Y15_O_top13, //EXTERNAL
        input Tile_X5Y15_O_top14, //EXTERNAL
        input Tile_X5Y15_O_top15, //EXTERNAL
        output Tile_X5Y15_I_top0, //EXTERNAL
        output Tile_X5Y15_I_top1, //EXTERNAL
        output Tile_X5Y15_I_top2, //EXTERNAL
        output Tile_X5Y15_I_top3, //EXTERNAL
        output Tile_X5Y15_I_top4, //EXTERNAL
        output Tile_X5Y15_I_top5, //EXTERNAL
        output Tile_X5Y15_I_top6, //EXTERNAL
        output Tile_X5Y15_I_top7, //EXTERNAL
        output Tile_X5Y15_I_top8, //EXTERNAL
        output Tile_X5Y15_I_top9, //EXTERNAL
        output Tile_X5Y15_I_top10, //EXTERNAL
        output Tile_X5Y15_I_top11, //EXTERNAL
        output Tile_X5Y15_I_top12, //EXTERNAL
        output Tile_X5Y15_I_top13, //EXTERNAL
        output Tile_X5Y15_I_top14, //EXTERNAL
        output Tile_X5Y15_I_top15, //EXTERNAL
        input Tile_X6Y15_O_top0, //EXTERNAL
        input Tile_X6Y15_O_top1, //EXTERNAL
        input Tile_X6Y15_O_top2, //EXTERNAL
        input Tile_X6Y15_O_top3, //EXTERNAL
        input Tile_X6Y15_O_top4, //EXTERNAL
        input Tile_X6Y15_O_top5, //EXTERNAL
        input Tile_X6Y15_O_top6, //EXTERNAL
        input Tile_X6Y15_O_top7, //EXTERNAL
        input Tile_X6Y15_O_top8, //EXTERNAL
        input Tile_X6Y15_O_top9, //EXTERNAL
        input Tile_X6Y15_O_top10, //EXTERNAL
        input Tile_X6Y15_O_top11, //EXTERNAL
        input Tile_X6Y15_O_top12, //EXTERNAL
        input Tile_X6Y15_O_top13, //EXTERNAL
        input Tile_X6Y15_O_top14, //EXTERNAL
        input Tile_X6Y15_O_top15, //EXTERNAL
        output Tile_X6Y15_I_top0, //EXTERNAL
        output Tile_X6Y15_I_top1, //EXTERNAL
        output Tile_X6Y15_I_top2, //EXTERNAL
        output Tile_X6Y15_I_top3, //EXTERNAL
        output Tile_X6Y15_I_top4, //EXTERNAL
        output Tile_X6Y15_I_top5, //EXTERNAL
        output Tile_X6Y15_I_top6, //EXTERNAL
        output Tile_X6Y15_I_top7, //EXTERNAL
        output Tile_X6Y15_I_top8, //EXTERNAL
        output Tile_X6Y15_I_top9, //EXTERNAL
        output Tile_X6Y15_I_top10, //EXTERNAL
        output Tile_X6Y15_I_top11, //EXTERNAL
        output Tile_X6Y15_I_top12, //EXTERNAL
        output Tile_X6Y15_I_top13, //EXTERNAL
        output Tile_X6Y15_I_top14, //EXTERNAL
        output Tile_X6Y15_I_top15, //EXTERNAL
        input Tile_X8Y15_O_top0, //EXTERNAL
        input Tile_X8Y15_O_top1, //EXTERNAL
        input Tile_X8Y15_O_top2, //EXTERNAL
        input Tile_X8Y15_O_top3, //EXTERNAL
        input Tile_X8Y15_O_top4, //EXTERNAL
        input Tile_X8Y15_O_top5, //EXTERNAL
        input Tile_X8Y15_O_top6, //EXTERNAL
        input Tile_X8Y15_O_top7, //EXTERNAL
        input Tile_X8Y15_O_top8, //EXTERNAL
        input Tile_X8Y15_O_top9, //EXTERNAL
        input Tile_X8Y15_O_top10, //EXTERNAL
        input Tile_X8Y15_O_top11, //EXTERNAL
        input Tile_X8Y15_O_top12, //EXTERNAL
        input Tile_X8Y15_O_top13, //EXTERNAL
        input Tile_X8Y15_O_top14, //EXTERNAL
        input Tile_X8Y15_O_top15, //EXTERNAL
        output Tile_X8Y15_I_top0, //EXTERNAL
        output Tile_X8Y15_I_top1, //EXTERNAL
        output Tile_X8Y15_I_top2, //EXTERNAL
        output Tile_X8Y15_I_top3, //EXTERNAL
        output Tile_X8Y15_I_top4, //EXTERNAL
        output Tile_X8Y15_I_top5, //EXTERNAL
        output Tile_X8Y15_I_top6, //EXTERNAL
        output Tile_X8Y15_I_top7, //EXTERNAL
        output Tile_X8Y15_I_top8, //EXTERNAL
        output Tile_X8Y15_I_top9, //EXTERNAL
        output Tile_X8Y15_I_top10, //EXTERNAL
        output Tile_X8Y15_I_top11, //EXTERNAL
        output Tile_X8Y15_I_top12, //EXTERNAL
        output Tile_X8Y15_I_top13, //EXTERNAL
        output Tile_X8Y15_I_top14, //EXTERNAL
        output Tile_X8Y15_I_top15, //EXTERNAL
        input Tile_X9Y15_O_top0, //EXTERNAL
        input Tile_X9Y15_O_top1, //EXTERNAL
        input Tile_X9Y15_O_top2, //EXTERNAL
        input Tile_X9Y15_O_top3, //EXTERNAL
        input Tile_X9Y15_O_top4, //EXTERNAL
        input Tile_X9Y15_O_top5, //EXTERNAL
        input Tile_X9Y15_O_top6, //EXTERNAL
        input Tile_X9Y15_O_top7, //EXTERNAL
        input Tile_X9Y15_O_top8, //EXTERNAL
        input Tile_X9Y15_O_top9, //EXTERNAL
        input Tile_X9Y15_O_top10, //EXTERNAL
        input Tile_X9Y15_O_top11, //EXTERNAL
        input Tile_X9Y15_O_top12, //EXTERNAL
        input Tile_X9Y15_O_top13, //EXTERNAL
        input Tile_X9Y15_O_top14, //EXTERNAL
        input Tile_X9Y15_O_top15, //EXTERNAL
        output Tile_X9Y15_I_top0, //EXTERNAL
        output Tile_X9Y15_I_top1, //EXTERNAL
        output Tile_X9Y15_I_top2, //EXTERNAL
        output Tile_X9Y15_I_top3, //EXTERNAL
        output Tile_X9Y15_I_top4, //EXTERNAL
        output Tile_X9Y15_I_top5, //EXTERNAL
        output Tile_X9Y15_I_top6, //EXTERNAL
        output Tile_X9Y15_I_top7, //EXTERNAL
        output Tile_X9Y15_I_top8, //EXTERNAL
        output Tile_X9Y15_I_top9, //EXTERNAL
        output Tile_X9Y15_I_top10, //EXTERNAL
        output Tile_X9Y15_I_top11, //EXTERNAL
        output Tile_X9Y15_I_top12, //EXTERNAL
        output Tile_X9Y15_I_top13, //EXTERNAL
        output Tile_X9Y15_I_top14, //EXTERNAL
        output Tile_X9Y15_I_top15, //EXTERNAL
        input [(FrameBitsPerRow*16)-1:0] FrameData, //CONFIG_PORT
        input [(MaxFramesPerCol*11)-1:0] FrameStrobe, //CONFIG_PORT
        input UserCLK
);

 //signal declarations

wire Tile_X0Y0_UserCLKo;
wire Tile_X1Y0_UserCLKo;
wire Tile_X2Y0_UserCLKo;
wire Tile_X3Y0_UserCLKo;
wire Tile_X4Y0_UserCLKo;
wire Tile_X5Y0_UserCLKo;
wire Tile_X6Y0_UserCLKo;
wire Tile_X7Y0_UserCLKo;
wire Tile_X8Y0_UserCLKo;
wire Tile_X9Y0_UserCLKo;
wire Tile_X10Y0_UserCLKo;
wire Tile_X0Y1_UserCLKo;
wire Tile_X1Y1_UserCLKo;
wire Tile_X2Y1_UserCLKo;
wire Tile_X3Y1_UserCLKo;
wire Tile_X4Y1_UserCLKo;
wire Tile_X5Y1_UserCLKo;
wire Tile_X6Y1_UserCLKo;
wire Tile_X7Y1_UserCLKo;
wire Tile_X8Y1_UserCLKo;
wire Tile_X9Y1_UserCLKo;
wire Tile_X10Y1_UserCLKo;
wire Tile_X0Y2_UserCLKo;
wire Tile_X1Y2_UserCLKo;
wire Tile_X2Y2_UserCLKo;
wire Tile_X3Y2_UserCLKo;
wire Tile_X4Y2_UserCLKo;
wire Tile_X5Y2_UserCLKo;
wire Tile_X6Y2_UserCLKo;
wire Tile_X7Y2_UserCLKo;
wire Tile_X8Y2_UserCLKo;
wire Tile_X9Y2_UserCLKo;
wire Tile_X10Y2_UserCLKo;
wire Tile_X0Y3_UserCLKo;
wire Tile_X1Y3_UserCLKo;
wire Tile_X2Y3_UserCLKo;
wire Tile_X3Y3_UserCLKo;
wire Tile_X4Y3_UserCLKo;
wire Tile_X5Y3_UserCLKo;
wire Tile_X6Y3_UserCLKo;
wire Tile_X7Y3_UserCLKo;
wire Tile_X8Y3_UserCLKo;
wire Tile_X9Y3_UserCLKo;
wire Tile_X10Y3_UserCLKo;
wire Tile_X0Y4_UserCLKo;
wire Tile_X1Y4_UserCLKo;
wire Tile_X2Y4_UserCLKo;
wire Tile_X3Y4_UserCLKo;
wire Tile_X4Y4_UserCLKo;
wire Tile_X5Y4_UserCLKo;
wire Tile_X6Y4_UserCLKo;
wire Tile_X7Y4_UserCLKo;
wire Tile_X8Y4_UserCLKo;
wire Tile_X9Y4_UserCLKo;
wire Tile_X10Y4_UserCLKo;
wire Tile_X0Y5_UserCLKo;
wire Tile_X1Y5_UserCLKo;
wire Tile_X2Y5_UserCLKo;
wire Tile_X3Y5_UserCLKo;
wire Tile_X4Y5_UserCLKo;
wire Tile_X5Y5_UserCLKo;
wire Tile_X6Y5_UserCLKo;
wire Tile_X7Y5_UserCLKo;
wire Tile_X8Y5_UserCLKo;
wire Tile_X9Y5_UserCLKo;
wire Tile_X10Y5_UserCLKo;
wire Tile_X0Y6_UserCLKo;
wire Tile_X1Y6_UserCLKo;
wire Tile_X2Y6_UserCLKo;
wire Tile_X3Y6_UserCLKo;
wire Tile_X4Y6_UserCLKo;
wire Tile_X5Y6_UserCLKo;
wire Tile_X6Y6_UserCLKo;
wire Tile_X7Y6_UserCLKo;
wire Tile_X8Y6_UserCLKo;
wire Tile_X9Y6_UserCLKo;
wire Tile_X10Y6_UserCLKo;
wire Tile_X0Y7_UserCLKo;
wire Tile_X1Y7_UserCLKo;
wire Tile_X2Y7_UserCLKo;
wire Tile_X3Y7_UserCLKo;
wire Tile_X4Y7_UserCLKo;
wire Tile_X5Y7_UserCLKo;
wire Tile_X6Y7_UserCLKo;
wire Tile_X7Y7_UserCLKo;
wire Tile_X8Y7_UserCLKo;
wire Tile_X9Y7_UserCLKo;
wire Tile_X10Y7_UserCLKo;
wire Tile_X0Y8_UserCLKo;
wire Tile_X1Y8_UserCLKo;
wire Tile_X2Y8_UserCLKo;
wire Tile_X3Y8_UserCLKo;
wire Tile_X4Y8_UserCLKo;
wire Tile_X5Y8_UserCLKo;
wire Tile_X6Y8_UserCLKo;
wire Tile_X7Y8_UserCLKo;
wire Tile_X8Y8_UserCLKo;
wire Tile_X9Y8_UserCLKo;
wire Tile_X10Y8_UserCLKo;
wire Tile_X0Y9_UserCLKo;
wire Tile_X1Y9_UserCLKo;
wire Tile_X2Y9_UserCLKo;
wire Tile_X3Y9_UserCLKo;
wire Tile_X4Y9_UserCLKo;
wire Tile_X5Y9_UserCLKo;
wire Tile_X6Y9_UserCLKo;
wire Tile_X7Y9_UserCLKo;
wire Tile_X8Y9_UserCLKo;
wire Tile_X9Y9_UserCLKo;
wire Tile_X10Y9_UserCLKo;
wire Tile_X0Y10_UserCLKo;
wire Tile_X1Y10_UserCLKo;
wire Tile_X2Y10_UserCLKo;
wire Tile_X3Y10_UserCLKo;
wire Tile_X4Y10_UserCLKo;
wire Tile_X5Y10_UserCLKo;
wire Tile_X6Y10_UserCLKo;
wire Tile_X7Y10_UserCLKo;
wire Tile_X8Y10_UserCLKo;
wire Tile_X9Y10_UserCLKo;
wire Tile_X10Y10_UserCLKo;
wire Tile_X0Y11_UserCLKo;
wire Tile_X1Y11_UserCLKo;
wire Tile_X2Y11_UserCLKo;
wire Tile_X3Y11_UserCLKo;
wire Tile_X4Y11_UserCLKo;
wire Tile_X5Y11_UserCLKo;
wire Tile_X6Y11_UserCLKo;
wire Tile_X7Y11_UserCLKo;
wire Tile_X8Y11_UserCLKo;
wire Tile_X9Y11_UserCLKo;
wire Tile_X10Y11_UserCLKo;
wire Tile_X0Y12_UserCLKo;
wire Tile_X1Y12_UserCLKo;
wire Tile_X2Y12_UserCLKo;
wire Tile_X3Y12_UserCLKo;
wire Tile_X4Y12_UserCLKo;
wire Tile_X5Y12_UserCLKo;
wire Tile_X6Y12_UserCLKo;
wire Tile_X7Y12_UserCLKo;
wire Tile_X8Y12_UserCLKo;
wire Tile_X9Y12_UserCLKo;
wire Tile_X10Y12_UserCLKo;
wire Tile_X0Y13_UserCLKo;
wire Tile_X1Y13_UserCLKo;
wire Tile_X2Y13_UserCLKo;
wire Tile_X3Y13_UserCLKo;
wire Tile_X4Y13_UserCLKo;
wire Tile_X5Y13_UserCLKo;
wire Tile_X6Y13_UserCLKo;
wire Tile_X7Y13_UserCLKo;
wire Tile_X8Y13_UserCLKo;
wire Tile_X9Y13_UserCLKo;
wire Tile_X10Y13_UserCLKo;
wire Tile_X0Y14_UserCLKo;
wire Tile_X1Y14_UserCLKo;
wire Tile_X2Y14_UserCLKo;
wire Tile_X3Y14_UserCLKo;
wire Tile_X4Y14_UserCLKo;
wire Tile_X5Y14_UserCLKo;
wire Tile_X6Y14_UserCLKo;
wire Tile_X7Y14_UserCLKo;
wire Tile_X8Y14_UserCLKo;
wire Tile_X9Y14_UserCLKo;
wire Tile_X10Y14_UserCLKo;
wire Tile_X0Y15_UserCLKo;
wire Tile_X1Y15_UserCLKo;
wire Tile_X2Y15_UserCLKo;
wire Tile_X3Y15_UserCLKo;
wire Tile_X4Y15_UserCLKo;
wire Tile_X5Y15_UserCLKo;
wire Tile_X6Y15_UserCLKo;
wire Tile_X7Y15_UserCLKo;
wire Tile_X8Y15_UserCLKo;
wire Tile_X9Y15_UserCLKo;
wire Tile_X10Y15_UserCLKo;
 //configuration signal declarations

wire[FrameBitsPerRow -1:0] Row_Y0_FrameData;
wire[FrameBitsPerRow -1:0] Row_Y1_FrameData;
wire[FrameBitsPerRow -1:0] Row_Y2_FrameData;
wire[FrameBitsPerRow -1:0] Row_Y3_FrameData;
wire[FrameBitsPerRow -1:0] Row_Y4_FrameData;
wire[FrameBitsPerRow -1:0] Row_Y5_FrameData;
wire[FrameBitsPerRow -1:0] Row_Y6_FrameData;
wire[FrameBitsPerRow -1:0] Row_Y7_FrameData;
wire[FrameBitsPerRow -1:0] Row_Y8_FrameData;
wire[FrameBitsPerRow -1:0] Row_Y9_FrameData;
wire[FrameBitsPerRow -1:0] Row_Y10_FrameData;
wire[FrameBitsPerRow -1:0] Row_Y11_FrameData;
wire[FrameBitsPerRow -1:0] Row_Y12_FrameData;
wire[FrameBitsPerRow -1:0] Row_Y13_FrameData;
wire[FrameBitsPerRow -1:0] Row_Y14_FrameData;
wire[FrameBitsPerRow -1:0] Row_Y15_FrameData;
wire[MaxFramesPerCol - 1:0] Column_X0_FrameStrobe;
wire[MaxFramesPerCol - 1:0] Column_X1_FrameStrobe;
wire[MaxFramesPerCol - 1:0] Column_X2_FrameStrobe;
wire[MaxFramesPerCol - 1:0] Column_X3_FrameStrobe;
wire[MaxFramesPerCol - 1:0] Column_X4_FrameStrobe;
wire[MaxFramesPerCol - 1:0] Column_X5_FrameStrobe;
wire[MaxFramesPerCol - 1:0] Column_X6_FrameStrobe;
wire[MaxFramesPerCol - 1:0] Column_X7_FrameStrobe;
wire[MaxFramesPerCol - 1:0] Column_X8_FrameStrobe;
wire[MaxFramesPerCol - 1:0] Column_X9_FrameStrobe;
wire[MaxFramesPerCol - 1:0] Column_X10_FrameStrobe;
wire[FrameBitsPerRow - 1:0] Tile_X0Y0_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X1Y0_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X2Y0_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X3Y0_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X4Y0_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X5Y0_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X6Y0_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X7Y0_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X8Y0_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X9Y0_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X10Y0_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X0Y1_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X1Y1_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X2Y1_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X3Y1_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X4Y1_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X5Y1_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X6Y1_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X7Y1_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X8Y1_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X9Y1_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X10Y1_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X0Y2_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X1Y2_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X2Y2_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X3Y2_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X4Y2_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X5Y2_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X6Y2_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X7Y2_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X8Y2_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X9Y2_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X10Y2_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X0Y3_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X1Y3_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X2Y3_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X3Y3_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X4Y3_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X5Y3_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X6Y3_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X7Y3_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X8Y3_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X9Y3_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X10Y3_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X0Y4_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X1Y4_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X2Y4_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X3Y4_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X4Y4_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X5Y4_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X6Y4_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X7Y4_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X8Y4_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X9Y4_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X10Y4_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X0Y5_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X1Y5_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X2Y5_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X3Y5_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X4Y5_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X5Y5_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X6Y5_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X7Y5_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X8Y5_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X9Y5_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X10Y5_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X0Y6_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X1Y6_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X2Y6_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X3Y6_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X4Y6_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X5Y6_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X6Y6_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X7Y6_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X8Y6_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X9Y6_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X10Y6_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X0Y7_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X1Y7_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X2Y7_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X3Y7_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X4Y7_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X5Y7_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X6Y7_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X7Y7_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X8Y7_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X9Y7_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X10Y7_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X0Y8_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X1Y8_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X2Y8_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X3Y8_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X4Y8_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X5Y8_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X6Y8_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X7Y8_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X8Y8_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X9Y8_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X10Y8_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X0Y9_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X1Y9_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X2Y9_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X3Y9_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X4Y9_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X5Y9_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X6Y9_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X7Y9_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X8Y9_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X9Y9_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X10Y9_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X0Y10_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X1Y10_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X2Y10_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X3Y10_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X4Y10_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X5Y10_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X6Y10_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X7Y10_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X8Y10_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X9Y10_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X10Y10_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X0Y11_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X1Y11_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X2Y11_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X3Y11_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X4Y11_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X5Y11_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X6Y11_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X7Y11_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X8Y11_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X9Y11_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X10Y11_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X0Y12_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X1Y12_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X2Y12_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X3Y12_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X4Y12_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X5Y12_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X6Y12_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X7Y12_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X8Y12_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X9Y12_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X10Y12_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X0Y13_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X1Y13_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X2Y13_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X3Y13_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X4Y13_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X5Y13_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X6Y13_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X7Y13_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X8Y13_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X9Y13_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X10Y13_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X0Y14_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X1Y14_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X2Y14_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X3Y14_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X4Y14_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X5Y14_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X6Y14_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X7Y14_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X8Y14_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X9Y14_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X10Y14_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X0Y15_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X1Y15_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X2Y15_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X3Y15_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X4Y15_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X5Y15_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X6Y15_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X7Y15_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X8Y15_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X9Y15_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X10Y15_FrameData_O;
wire[MaxFramesPerCol - 1:0] Tile_X0Y0_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X1Y0_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X2Y0_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X3Y0_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X4Y0_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X5Y0_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X6Y0_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X7Y0_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X8Y0_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X9Y0_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X10Y0_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X0Y1_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X1Y1_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X2Y1_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X3Y1_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X4Y1_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X5Y1_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X6Y1_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X7Y1_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X8Y1_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X9Y1_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X10Y1_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X0Y2_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X1Y2_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X2Y2_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X3Y2_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X4Y2_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X5Y2_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X6Y2_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X7Y2_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X8Y2_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X9Y2_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X10Y2_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X0Y3_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X1Y3_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X2Y3_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X3Y3_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X4Y3_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X5Y3_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X6Y3_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X7Y3_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X8Y3_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X9Y3_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X10Y3_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X0Y4_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X1Y4_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X2Y4_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X3Y4_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X4Y4_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X5Y4_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X6Y4_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X7Y4_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X8Y4_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X9Y4_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X10Y4_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X0Y5_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X1Y5_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X2Y5_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X3Y5_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X4Y5_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X5Y5_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X6Y5_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X7Y5_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X8Y5_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X9Y5_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X10Y5_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X0Y6_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X1Y6_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X2Y6_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X3Y6_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X4Y6_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X5Y6_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X6Y6_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X7Y6_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X8Y6_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X9Y6_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X10Y6_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X0Y7_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X1Y7_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X2Y7_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X3Y7_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X4Y7_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X5Y7_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X6Y7_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X7Y7_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X8Y7_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X9Y7_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X10Y7_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X0Y8_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X1Y8_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X2Y8_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X3Y8_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X4Y8_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X5Y8_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X6Y8_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X7Y8_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X8Y8_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X9Y8_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X10Y8_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X0Y9_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X1Y9_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X2Y9_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X3Y9_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X4Y9_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X5Y9_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X6Y9_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X7Y9_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X8Y9_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X9Y9_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X10Y9_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X0Y10_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X1Y10_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X2Y10_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X3Y10_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X4Y10_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X5Y10_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X6Y10_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X7Y10_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X8Y10_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X9Y10_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X10Y10_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X0Y11_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X1Y11_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X2Y11_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X3Y11_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X4Y11_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X5Y11_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X6Y11_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X7Y11_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X8Y11_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X9Y11_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X10Y11_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X0Y12_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X1Y12_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X2Y12_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X3Y12_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X4Y12_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X5Y12_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X6Y12_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X7Y12_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X8Y12_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X9Y12_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X10Y12_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X0Y13_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X1Y13_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X2Y13_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X3Y13_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X4Y13_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X5Y13_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X6Y13_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X7Y13_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X8Y13_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X9Y13_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X10Y13_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X0Y14_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X1Y14_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X2Y14_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X3Y14_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X4Y14_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X5Y14_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X6Y14_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X7Y14_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X8Y14_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X9Y14_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X10Y14_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X0Y15_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X1Y15_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X2Y15_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X3Y15_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X4Y15_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X5Y15_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X6Y15_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X7Y15_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X8Y15_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X9Y15_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X10Y15_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X0Y16_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X1Y16_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X2Y16_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X3Y16_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X4Y16_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X5Y16_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X6Y16_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X7Y16_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X8Y16_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X9Y16_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X10Y16_FrameStrobe_O;
 //tile-to-tile signal declarations
wire[3:0] Tile_X1Y0_S1BEG;
wire[7:0] Tile_X1Y0_S2BEG;
wire[7:0] Tile_X1Y0_S2BEGb;
wire[15:0] Tile_X1Y0_S4BEG;
wire[15:0] Tile_X1Y0_SS4BEG;
wire[3:0] Tile_X2Y0_S1BEG;
wire[7:0] Tile_X2Y0_S2BEG;
wire[7:0] Tile_X2Y0_S2BEGb;
wire[15:0] Tile_X2Y0_S4BEG;
wire[15:0] Tile_X2Y0_SS4BEG;
wire[3:0] Tile_X3Y0_S1BEG;
wire[7:0] Tile_X3Y0_S2BEG;
wire[7:0] Tile_X3Y0_S2BEGb;
wire[15:0] Tile_X3Y0_S4BEG;
wire[15:0] Tile_X3Y0_SS4BEG;
wire[3:0] Tile_X4Y0_S1BEG;
wire[7:0] Tile_X4Y0_S2BEG;
wire[7:0] Tile_X4Y0_S2BEGb;
wire[15:0] Tile_X4Y0_S4BEG;
wire[15:0] Tile_X4Y0_SS4BEG;
wire[3:0] Tile_X5Y0_S1BEG;
wire[7:0] Tile_X5Y0_S2BEG;
wire[7:0] Tile_X5Y0_S2BEGb;
wire[15:0] Tile_X5Y0_S4BEG;
wire[15:0] Tile_X5Y0_SS4BEG;
wire[3:0] Tile_X6Y0_S1BEG;
wire[7:0] Tile_X6Y0_S2BEG;
wire[7:0] Tile_X6Y0_S2BEGb;
wire[15:0] Tile_X6Y0_S4BEG;
wire[15:0] Tile_X6Y0_SS4BEG;
wire[3:0] Tile_X7Y0_S1BEG;
wire[7:0] Tile_X7Y0_S2BEG;
wire[7:0] Tile_X7Y0_S2BEGb;
wire[15:0] Tile_X7Y0_S4BEG;
wire[15:0] Tile_X7Y0_SS4BEG;
wire[3:0] Tile_X8Y0_S1BEG;
wire[7:0] Tile_X8Y0_S2BEG;
wire[7:0] Tile_X8Y0_S2BEGb;
wire[15:0] Tile_X8Y0_S4BEG;
wire[15:0] Tile_X8Y0_SS4BEG;
wire[3:0] Tile_X9Y0_S1BEG;
wire[7:0] Tile_X9Y0_S2BEG;
wire[7:0] Tile_X9Y0_S2BEGb;
wire[15:0] Tile_X9Y0_S4BEG;
wire[15:0] Tile_X9Y0_SS4BEG;
wire[3:0] Tile_X10Y0_S1BEG;
wire[7:0] Tile_X10Y0_S2BEG;
wire[7:0] Tile_X10Y0_S2BEGb;
wire[15:0] Tile_X10Y0_S4BEG;
wire[3:0] Tile_X0Y1_E1BEG;
wire[7:0] Tile_X0Y1_E2BEG;
wire[7:0] Tile_X0Y1_E2BEGb;
wire[15:0] Tile_X0Y1_EE4BEG;
wire[11:0] Tile_X0Y1_E6BEG;
wire[3:0] Tile_X1Y1_N1BEG;
wire[7:0] Tile_X1Y1_N2BEG;
wire[7:0] Tile_X1Y1_N2BEGb;
wire[15:0] Tile_X1Y1_N4BEG;
wire[15:0] Tile_X1Y1_NN4BEG;
wire[3:0] Tile_X1Y1_E1BEG;
wire[7:0] Tile_X1Y1_E2BEG;
wire[7:0] Tile_X1Y1_E2BEGb;
wire[15:0] Tile_X1Y1_EE4BEG;
wire[11:0] Tile_X1Y1_E6BEG;
wire[3:0] Tile_X1Y1_S1BEG;
wire[7:0] Tile_X1Y1_S2BEG;
wire[7:0] Tile_X1Y1_S2BEGb;
wire[15:0] Tile_X1Y1_S4BEG;
wire[15:0] Tile_X1Y1_SS4BEG;
wire[3:0] Tile_X1Y1_W1BEG;
wire[7:0] Tile_X1Y1_W2BEG;
wire[7:0] Tile_X1Y1_W2BEGb;
wire[15:0] Tile_X1Y1_WW4BEG;
wire[11:0] Tile_X1Y1_W6BEG;
wire[0:0] Tile_X1Y1_Co;
wire[3:0] Tile_X2Y1_N1BEG;
wire[7:0] Tile_X2Y1_N2BEG;
wire[7:0] Tile_X2Y1_N2BEGb;
wire[15:0] Tile_X2Y1_N4BEG;
wire[15:0] Tile_X2Y1_NN4BEG;
wire[3:0] Tile_X2Y1_E1BEG;
wire[7:0] Tile_X2Y1_E2BEG;
wire[7:0] Tile_X2Y1_E2BEGb;
wire[15:0] Tile_X2Y1_EE4BEG;
wire[11:0] Tile_X2Y1_E6BEG;
wire[3:0] Tile_X2Y1_S1BEG;
wire[7:0] Tile_X2Y1_S2BEG;
wire[7:0] Tile_X2Y1_S2BEGb;
wire[15:0] Tile_X2Y1_S4BEG;
wire[15:0] Tile_X2Y1_SS4BEG;
wire[3:0] Tile_X2Y1_W1BEG;
wire[7:0] Tile_X2Y1_W2BEG;
wire[7:0] Tile_X2Y1_W2BEGb;
wire[15:0] Tile_X2Y1_WW4BEG;
wire[11:0] Tile_X2Y1_W6BEG;
wire[0:0] Tile_X2Y1_Co;
wire[3:0] Tile_X3Y1_N1BEG;
wire[7:0] Tile_X3Y1_N2BEG;
wire[7:0] Tile_X3Y1_N2BEGb;
wire[15:0] Tile_X3Y1_N4BEG;
wire[15:0] Tile_X3Y1_NN4BEG;
wire[3:0] Tile_X3Y1_E1BEG;
wire[7:0] Tile_X3Y1_E2BEG;
wire[7:0] Tile_X3Y1_E2BEGb;
wire[15:0] Tile_X3Y1_EE4BEG;
wire[11:0] Tile_X3Y1_E6BEG;
wire[3:0] Tile_X3Y1_S1BEG;
wire[7:0] Tile_X3Y1_S2BEG;
wire[7:0] Tile_X3Y1_S2BEGb;
wire[15:0] Tile_X3Y1_S4BEG;
wire[15:0] Tile_X3Y1_SS4BEG;
wire[3:0] Tile_X3Y1_W1BEG;
wire[7:0] Tile_X3Y1_W2BEG;
wire[7:0] Tile_X3Y1_W2BEGb;
wire[15:0] Tile_X3Y1_WW4BEG;
wire[11:0] Tile_X3Y1_W6BEG;
wire[0:0] Tile_X3Y1_Co;
wire[3:0] Tile_X4Y1_N1BEG;
wire[7:0] Tile_X4Y1_N2BEG;
wire[7:0] Tile_X4Y1_N2BEGb;
wire[15:0] Tile_X4Y1_N4BEG;
wire[15:0] Tile_X4Y1_NN4BEG;
wire[3:0] Tile_X4Y1_E1BEG;
wire[7:0] Tile_X4Y1_E2BEG;
wire[7:0] Tile_X4Y1_E2BEGb;
wire[15:0] Tile_X4Y1_EE4BEG;
wire[11:0] Tile_X4Y1_E6BEG;
wire[3:0] Tile_X4Y1_S1BEG;
wire[7:0] Tile_X4Y1_S2BEG;
wire[7:0] Tile_X4Y1_S2BEGb;
wire[15:0] Tile_X4Y1_S4BEG;
wire[15:0] Tile_X4Y1_SS4BEG;
wire[3:0] Tile_X4Y1_W1BEG;
wire[7:0] Tile_X4Y1_W2BEG;
wire[7:0] Tile_X4Y1_W2BEGb;
wire[15:0] Tile_X4Y1_WW4BEG;
wire[11:0] Tile_X4Y1_W6BEG;
wire[3:0] Tile_X5Y1_N1BEG;
wire[7:0] Tile_X5Y1_N2BEG;
wire[7:0] Tile_X5Y1_N2BEGb;
wire[15:0] Tile_X5Y1_N4BEG;
wire[15:0] Tile_X5Y1_NN4BEG;
wire[3:0] Tile_X5Y1_E1BEG;
wire[7:0] Tile_X5Y1_E2BEG;
wire[7:0] Tile_X5Y1_E2BEGb;
wire[15:0] Tile_X5Y1_EE4BEG;
wire[11:0] Tile_X5Y1_E6BEG;
wire[3:0] Tile_X5Y1_S1BEG;
wire[7:0] Tile_X5Y1_S2BEG;
wire[7:0] Tile_X5Y1_S2BEGb;
wire[15:0] Tile_X5Y1_S4BEG;
wire[15:0] Tile_X5Y1_SS4BEG;
wire[3:0] Tile_X5Y1_W1BEG;
wire[7:0] Tile_X5Y1_W2BEG;
wire[7:0] Tile_X5Y1_W2BEGb;
wire[15:0] Tile_X5Y1_WW4BEG;
wire[11:0] Tile_X5Y1_W6BEG;
wire[0:0] Tile_X5Y1_Co;
wire[3:0] Tile_X6Y1_N1BEG;
wire[7:0] Tile_X6Y1_N2BEG;
wire[7:0] Tile_X6Y1_N2BEGb;
wire[15:0] Tile_X6Y1_N4BEG;
wire[15:0] Tile_X6Y1_NN4BEG;
wire[3:0] Tile_X6Y1_E1BEG;
wire[7:0] Tile_X6Y1_E2BEG;
wire[7:0] Tile_X6Y1_E2BEGb;
wire[15:0] Tile_X6Y1_EE4BEG;
wire[11:0] Tile_X6Y1_E6BEG;
wire[3:0] Tile_X6Y1_S1BEG;
wire[7:0] Tile_X6Y1_S2BEG;
wire[7:0] Tile_X6Y1_S2BEGb;
wire[15:0] Tile_X6Y1_S4BEG;
wire[15:0] Tile_X6Y1_SS4BEG;
wire[3:0] Tile_X6Y1_W1BEG;
wire[7:0] Tile_X6Y1_W2BEG;
wire[7:0] Tile_X6Y1_W2BEGb;
wire[15:0] Tile_X6Y1_WW4BEG;
wire[11:0] Tile_X6Y1_W6BEG;
wire[0:0] Tile_X6Y1_Co;
wire[3:0] Tile_X7Y1_N1BEG;
wire[7:0] Tile_X7Y1_N2BEG;
wire[7:0] Tile_X7Y1_N2BEGb;
wire[15:0] Tile_X7Y1_N4BEG;
wire[15:0] Tile_X7Y1_NN4BEG;
wire[3:0] Tile_X7Y1_E1BEG;
wire[7:0] Tile_X7Y1_E2BEG;
wire[7:0] Tile_X7Y1_E2BEGb;
wire[15:0] Tile_X7Y1_EE4BEG;
wire[11:0] Tile_X7Y1_E6BEG;
wire[3:0] Tile_X7Y1_S1BEG;
wire[7:0] Tile_X7Y1_S2BEG;
wire[7:0] Tile_X7Y1_S2BEGb;
wire[15:0] Tile_X7Y1_S4BEG;
wire[15:0] Tile_X7Y1_SS4BEG;
wire[3:0] Tile_X7Y1_W1BEG;
wire[7:0] Tile_X7Y1_W2BEG;
wire[7:0] Tile_X7Y1_W2BEGb;
wire[15:0] Tile_X7Y1_WW4BEG;
wire[11:0] Tile_X7Y1_W6BEG;
wire[17:0] Tile_X7Y1_top2bot;
wire[3:0] Tile_X8Y1_N1BEG;
wire[7:0] Tile_X8Y1_N2BEG;
wire[7:0] Tile_X8Y1_N2BEGb;
wire[15:0] Tile_X8Y1_N4BEG;
wire[15:0] Tile_X8Y1_NN4BEG;
wire[3:0] Tile_X8Y1_E1BEG;
wire[7:0] Tile_X8Y1_E2BEG;
wire[7:0] Tile_X8Y1_E2BEGb;
wire[15:0] Tile_X8Y1_EE4BEG;
wire[11:0] Tile_X8Y1_E6BEG;
wire[3:0] Tile_X8Y1_S1BEG;
wire[7:0] Tile_X8Y1_S2BEG;
wire[7:0] Tile_X8Y1_S2BEGb;
wire[15:0] Tile_X8Y1_S4BEG;
wire[15:0] Tile_X8Y1_SS4BEG;
wire[3:0] Tile_X8Y1_W1BEG;
wire[7:0] Tile_X8Y1_W2BEG;
wire[7:0] Tile_X8Y1_W2BEGb;
wire[15:0] Tile_X8Y1_WW4BEG;
wire[11:0] Tile_X8Y1_W6BEG;
wire[0:0] Tile_X8Y1_Co;
wire[3:0] Tile_X9Y1_N1BEG;
wire[7:0] Tile_X9Y1_N2BEG;
wire[7:0] Tile_X9Y1_N2BEGb;
wire[15:0] Tile_X9Y1_N4BEG;
wire[15:0] Tile_X9Y1_NN4BEG;
wire[3:0] Tile_X9Y1_E1BEG;
wire[7:0] Tile_X9Y1_E2BEG;
wire[7:0] Tile_X9Y1_E2BEGb;
wire[15:0] Tile_X9Y1_EE4BEG;
wire[11:0] Tile_X9Y1_E6BEG;
wire[3:0] Tile_X9Y1_S1BEG;
wire[7:0] Tile_X9Y1_S2BEG;
wire[7:0] Tile_X9Y1_S2BEGb;
wire[15:0] Tile_X9Y1_S4BEG;
wire[15:0] Tile_X9Y1_SS4BEG;
wire[3:0] Tile_X9Y1_W1BEG;
wire[7:0] Tile_X9Y1_W2BEG;
wire[7:0] Tile_X9Y1_W2BEGb;
wire[15:0] Tile_X9Y1_WW4BEG;
wire[11:0] Tile_X9Y1_W6BEG;
wire[0:0] Tile_X9Y1_Co;
wire[3:0] Tile_X10Y1_N1BEG;
wire[7:0] Tile_X10Y1_N2BEG;
wire[7:0] Tile_X10Y1_N2BEGb;
wire[15:0] Tile_X10Y1_N4BEG;
wire[3:0] Tile_X10Y1_S1BEG;
wire[7:0] Tile_X10Y1_S2BEG;
wire[7:0] Tile_X10Y1_S2BEGb;
wire[15:0] Tile_X10Y1_S4BEG;
wire[3:0] Tile_X10Y1_W1BEG;
wire[7:0] Tile_X10Y1_W2BEG;
wire[7:0] Tile_X10Y1_W2BEGb;
wire[15:0] Tile_X10Y1_WW4BEG;
wire[11:0] Tile_X10Y1_W6BEG;
wire[15:0] Tile_X10Y1_top2bot_DIN;
wire[15:0] Tile_X10Y1_top2bot_BM;
wire[4:0] Tile_X10Y1_top2bot_ADDR;
wire[3:0] Tile_X0Y2_E1BEG;
wire[7:0] Tile_X0Y2_E2BEG;
wire[7:0] Tile_X0Y2_E2BEGb;
wire[15:0] Tile_X0Y2_EE4BEG;
wire[11:0] Tile_X0Y2_E6BEG;
wire[3:0] Tile_X1Y2_N1BEG;
wire[7:0] Tile_X1Y2_N2BEG;
wire[7:0] Tile_X1Y2_N2BEGb;
wire[15:0] Tile_X1Y2_N4BEG;
wire[15:0] Tile_X1Y2_NN4BEG;
wire[3:0] Tile_X1Y2_E1BEG;
wire[7:0] Tile_X1Y2_E2BEG;
wire[7:0] Tile_X1Y2_E2BEGb;
wire[15:0] Tile_X1Y2_EE4BEG;
wire[11:0] Tile_X1Y2_E6BEG;
wire[3:0] Tile_X1Y2_S1BEG;
wire[7:0] Tile_X1Y2_S2BEG;
wire[7:0] Tile_X1Y2_S2BEGb;
wire[15:0] Tile_X1Y2_S4BEG;
wire[15:0] Tile_X1Y2_SS4BEG;
wire[3:0] Tile_X1Y2_W1BEG;
wire[7:0] Tile_X1Y2_W2BEG;
wire[7:0] Tile_X1Y2_W2BEGb;
wire[15:0] Tile_X1Y2_WW4BEG;
wire[11:0] Tile_X1Y2_W6BEG;
wire[0:0] Tile_X1Y2_Co;
wire[3:0] Tile_X2Y2_N1BEG;
wire[7:0] Tile_X2Y2_N2BEG;
wire[7:0] Tile_X2Y2_N2BEGb;
wire[15:0] Tile_X2Y2_N4BEG;
wire[15:0] Tile_X2Y2_NN4BEG;
wire[3:0] Tile_X2Y2_E1BEG;
wire[7:0] Tile_X2Y2_E2BEG;
wire[7:0] Tile_X2Y2_E2BEGb;
wire[15:0] Tile_X2Y2_EE4BEG;
wire[11:0] Tile_X2Y2_E6BEG;
wire[3:0] Tile_X2Y2_S1BEG;
wire[7:0] Tile_X2Y2_S2BEG;
wire[7:0] Tile_X2Y2_S2BEGb;
wire[15:0] Tile_X2Y2_S4BEG;
wire[15:0] Tile_X2Y2_SS4BEG;
wire[3:0] Tile_X2Y2_W1BEG;
wire[7:0] Tile_X2Y2_W2BEG;
wire[7:0] Tile_X2Y2_W2BEGb;
wire[15:0] Tile_X2Y2_WW4BEG;
wire[11:0] Tile_X2Y2_W6BEG;
wire[0:0] Tile_X2Y2_Co;
wire[3:0] Tile_X3Y2_N1BEG;
wire[7:0] Tile_X3Y2_N2BEG;
wire[7:0] Tile_X3Y2_N2BEGb;
wire[15:0] Tile_X3Y2_N4BEG;
wire[15:0] Tile_X3Y2_NN4BEG;
wire[3:0] Tile_X3Y2_E1BEG;
wire[7:0] Tile_X3Y2_E2BEG;
wire[7:0] Tile_X3Y2_E2BEGb;
wire[15:0] Tile_X3Y2_EE4BEG;
wire[11:0] Tile_X3Y2_E6BEG;
wire[3:0] Tile_X3Y2_S1BEG;
wire[7:0] Tile_X3Y2_S2BEG;
wire[7:0] Tile_X3Y2_S2BEGb;
wire[15:0] Tile_X3Y2_S4BEG;
wire[15:0] Tile_X3Y2_SS4BEG;
wire[3:0] Tile_X3Y2_W1BEG;
wire[7:0] Tile_X3Y2_W2BEG;
wire[7:0] Tile_X3Y2_W2BEGb;
wire[15:0] Tile_X3Y2_WW4BEG;
wire[11:0] Tile_X3Y2_W6BEG;
wire[0:0] Tile_X3Y2_Co;
wire[3:0] Tile_X4Y2_N1BEG;
wire[7:0] Tile_X4Y2_N2BEG;
wire[7:0] Tile_X4Y2_N2BEGb;
wire[15:0] Tile_X4Y2_N4BEG;
wire[15:0] Tile_X4Y2_NN4BEG;
wire[3:0] Tile_X4Y2_E1BEG;
wire[7:0] Tile_X4Y2_E2BEG;
wire[7:0] Tile_X4Y2_E2BEGb;
wire[15:0] Tile_X4Y2_EE4BEG;
wire[11:0] Tile_X4Y2_E6BEG;
wire[3:0] Tile_X4Y2_S1BEG;
wire[7:0] Tile_X4Y2_S2BEG;
wire[7:0] Tile_X4Y2_S2BEGb;
wire[15:0] Tile_X4Y2_S4BEG;
wire[15:0] Tile_X4Y2_SS4BEG;
wire[3:0] Tile_X4Y2_W1BEG;
wire[7:0] Tile_X4Y2_W2BEG;
wire[7:0] Tile_X4Y2_W2BEGb;
wire[15:0] Tile_X4Y2_WW4BEG;
wire[11:0] Tile_X4Y2_W6BEG;
wire[3:0] Tile_X5Y2_N1BEG;
wire[7:0] Tile_X5Y2_N2BEG;
wire[7:0] Tile_X5Y2_N2BEGb;
wire[15:0] Tile_X5Y2_N4BEG;
wire[15:0] Tile_X5Y2_NN4BEG;
wire[3:0] Tile_X5Y2_E1BEG;
wire[7:0] Tile_X5Y2_E2BEG;
wire[7:0] Tile_X5Y2_E2BEGb;
wire[15:0] Tile_X5Y2_EE4BEG;
wire[11:0] Tile_X5Y2_E6BEG;
wire[3:0] Tile_X5Y2_S1BEG;
wire[7:0] Tile_X5Y2_S2BEG;
wire[7:0] Tile_X5Y2_S2BEGb;
wire[15:0] Tile_X5Y2_S4BEG;
wire[15:0] Tile_X5Y2_SS4BEG;
wire[3:0] Tile_X5Y2_W1BEG;
wire[7:0] Tile_X5Y2_W2BEG;
wire[7:0] Tile_X5Y2_W2BEGb;
wire[15:0] Tile_X5Y2_WW4BEG;
wire[11:0] Tile_X5Y2_W6BEG;
wire[0:0] Tile_X5Y2_Co;
wire[3:0] Tile_X6Y2_N1BEG;
wire[7:0] Tile_X6Y2_N2BEG;
wire[7:0] Tile_X6Y2_N2BEGb;
wire[15:0] Tile_X6Y2_N4BEG;
wire[15:0] Tile_X6Y2_NN4BEG;
wire[3:0] Tile_X6Y2_E1BEG;
wire[7:0] Tile_X6Y2_E2BEG;
wire[7:0] Tile_X6Y2_E2BEGb;
wire[15:0] Tile_X6Y2_EE4BEG;
wire[11:0] Tile_X6Y2_E6BEG;
wire[3:0] Tile_X6Y2_S1BEG;
wire[7:0] Tile_X6Y2_S2BEG;
wire[7:0] Tile_X6Y2_S2BEGb;
wire[15:0] Tile_X6Y2_S4BEG;
wire[15:0] Tile_X6Y2_SS4BEG;
wire[3:0] Tile_X6Y2_W1BEG;
wire[7:0] Tile_X6Y2_W2BEG;
wire[7:0] Tile_X6Y2_W2BEGb;
wire[15:0] Tile_X6Y2_WW4BEG;
wire[11:0] Tile_X6Y2_W6BEG;
wire[0:0] Tile_X6Y2_Co;
wire[3:0] Tile_X7Y2_N1BEG;
wire[7:0] Tile_X7Y2_N2BEG;
wire[7:0] Tile_X7Y2_N2BEGb;
wire[15:0] Tile_X7Y2_N4BEG;
wire[15:0] Tile_X7Y2_NN4BEG;
wire[3:0] Tile_X7Y2_E1BEG;
wire[7:0] Tile_X7Y2_E2BEG;
wire[7:0] Tile_X7Y2_E2BEGb;
wire[15:0] Tile_X7Y2_EE4BEG;
wire[11:0] Tile_X7Y2_E6BEG;
wire[3:0] Tile_X7Y2_S1BEG;
wire[7:0] Tile_X7Y2_S2BEG;
wire[7:0] Tile_X7Y2_S2BEGb;
wire[15:0] Tile_X7Y2_S4BEG;
wire[15:0] Tile_X7Y2_SS4BEG;
wire[3:0] Tile_X7Y2_W1BEG;
wire[7:0] Tile_X7Y2_W2BEG;
wire[7:0] Tile_X7Y2_W2BEGb;
wire[15:0] Tile_X7Y2_WW4BEG;
wire[11:0] Tile_X7Y2_W6BEG;
wire[9:0] Tile_X7Y2_bot2top;
wire[3:0] Tile_X8Y2_N1BEG;
wire[7:0] Tile_X8Y2_N2BEG;
wire[7:0] Tile_X8Y2_N2BEGb;
wire[15:0] Tile_X8Y2_N4BEG;
wire[15:0] Tile_X8Y2_NN4BEG;
wire[3:0] Tile_X8Y2_E1BEG;
wire[7:0] Tile_X8Y2_E2BEG;
wire[7:0] Tile_X8Y2_E2BEGb;
wire[15:0] Tile_X8Y2_EE4BEG;
wire[11:0] Tile_X8Y2_E6BEG;
wire[3:0] Tile_X8Y2_S1BEG;
wire[7:0] Tile_X8Y2_S2BEG;
wire[7:0] Tile_X8Y2_S2BEGb;
wire[15:0] Tile_X8Y2_S4BEG;
wire[15:0] Tile_X8Y2_SS4BEG;
wire[3:0] Tile_X8Y2_W1BEG;
wire[7:0] Tile_X8Y2_W2BEG;
wire[7:0] Tile_X8Y2_W2BEGb;
wire[15:0] Tile_X8Y2_WW4BEG;
wire[11:0] Tile_X8Y2_W6BEG;
wire[0:0] Tile_X8Y2_Co;
wire[3:0] Tile_X9Y2_N1BEG;
wire[7:0] Tile_X9Y2_N2BEG;
wire[7:0] Tile_X9Y2_N2BEGb;
wire[15:0] Tile_X9Y2_N4BEG;
wire[15:0] Tile_X9Y2_NN4BEG;
wire[3:0] Tile_X9Y2_E1BEG;
wire[7:0] Tile_X9Y2_E2BEG;
wire[7:0] Tile_X9Y2_E2BEGb;
wire[15:0] Tile_X9Y2_EE4BEG;
wire[11:0] Tile_X9Y2_E6BEG;
wire[3:0] Tile_X9Y2_S1BEG;
wire[7:0] Tile_X9Y2_S2BEG;
wire[7:0] Tile_X9Y2_S2BEGb;
wire[15:0] Tile_X9Y2_S4BEG;
wire[15:0] Tile_X9Y2_SS4BEG;
wire[3:0] Tile_X9Y2_W1BEG;
wire[7:0] Tile_X9Y2_W2BEG;
wire[7:0] Tile_X9Y2_W2BEGb;
wire[15:0] Tile_X9Y2_WW4BEG;
wire[11:0] Tile_X9Y2_W6BEG;
wire[0:0] Tile_X9Y2_Co;
wire[3:0] Tile_X10Y2_N1BEG;
wire[7:0] Tile_X10Y2_N2BEG;
wire[7:0] Tile_X10Y2_N2BEGb;
wire[15:0] Tile_X10Y2_N4BEG;
wire[3:0] Tile_X10Y2_S1BEG;
wire[7:0] Tile_X10Y2_S2BEG;
wire[7:0] Tile_X10Y2_S2BEGb;
wire[15:0] Tile_X10Y2_S4BEG;
wire[3:0] Tile_X10Y2_W1BEG;
wire[7:0] Tile_X10Y2_W2BEG;
wire[7:0] Tile_X10Y2_W2BEGb;
wire[15:0] Tile_X10Y2_WW4BEG;
wire[11:0] Tile_X10Y2_W6BEG;
wire[15:0] Tile_X10Y2_bot2top_DOUT;
wire[3:0] Tile_X0Y3_E1BEG;
wire[7:0] Tile_X0Y3_E2BEG;
wire[7:0] Tile_X0Y3_E2BEGb;
wire[15:0] Tile_X0Y3_EE4BEG;
wire[11:0] Tile_X0Y3_E6BEG;
wire[3:0] Tile_X1Y3_N1BEG;
wire[7:0] Tile_X1Y3_N2BEG;
wire[7:0] Tile_X1Y3_N2BEGb;
wire[15:0] Tile_X1Y3_N4BEG;
wire[15:0] Tile_X1Y3_NN4BEG;
wire[3:0] Tile_X1Y3_E1BEG;
wire[7:0] Tile_X1Y3_E2BEG;
wire[7:0] Tile_X1Y3_E2BEGb;
wire[15:0] Tile_X1Y3_EE4BEG;
wire[11:0] Tile_X1Y3_E6BEG;
wire[3:0] Tile_X1Y3_S1BEG;
wire[7:0] Tile_X1Y3_S2BEG;
wire[7:0] Tile_X1Y3_S2BEGb;
wire[15:0] Tile_X1Y3_S4BEG;
wire[15:0] Tile_X1Y3_SS4BEG;
wire[3:0] Tile_X1Y3_W1BEG;
wire[7:0] Tile_X1Y3_W2BEG;
wire[7:0] Tile_X1Y3_W2BEGb;
wire[15:0] Tile_X1Y3_WW4BEG;
wire[11:0] Tile_X1Y3_W6BEG;
wire[0:0] Tile_X1Y3_Co;
wire[3:0] Tile_X2Y3_N1BEG;
wire[7:0] Tile_X2Y3_N2BEG;
wire[7:0] Tile_X2Y3_N2BEGb;
wire[15:0] Tile_X2Y3_N4BEG;
wire[15:0] Tile_X2Y3_NN4BEG;
wire[3:0] Tile_X2Y3_E1BEG;
wire[7:0] Tile_X2Y3_E2BEG;
wire[7:0] Tile_X2Y3_E2BEGb;
wire[15:0] Tile_X2Y3_EE4BEG;
wire[11:0] Tile_X2Y3_E6BEG;
wire[3:0] Tile_X2Y3_S1BEG;
wire[7:0] Tile_X2Y3_S2BEG;
wire[7:0] Tile_X2Y3_S2BEGb;
wire[15:0] Tile_X2Y3_S4BEG;
wire[15:0] Tile_X2Y3_SS4BEG;
wire[3:0] Tile_X2Y3_W1BEG;
wire[7:0] Tile_X2Y3_W2BEG;
wire[7:0] Tile_X2Y3_W2BEGb;
wire[15:0] Tile_X2Y3_WW4BEG;
wire[11:0] Tile_X2Y3_W6BEG;
wire[0:0] Tile_X2Y3_Co;
wire[3:0] Tile_X3Y3_N1BEG;
wire[7:0] Tile_X3Y3_N2BEG;
wire[7:0] Tile_X3Y3_N2BEGb;
wire[15:0] Tile_X3Y3_N4BEG;
wire[15:0] Tile_X3Y3_NN4BEG;
wire[3:0] Tile_X3Y3_E1BEG;
wire[7:0] Tile_X3Y3_E2BEG;
wire[7:0] Tile_X3Y3_E2BEGb;
wire[15:0] Tile_X3Y3_EE4BEG;
wire[11:0] Tile_X3Y3_E6BEG;
wire[3:0] Tile_X3Y3_S1BEG;
wire[7:0] Tile_X3Y3_S2BEG;
wire[7:0] Tile_X3Y3_S2BEGb;
wire[15:0] Tile_X3Y3_S4BEG;
wire[15:0] Tile_X3Y3_SS4BEG;
wire[3:0] Tile_X3Y3_W1BEG;
wire[7:0] Tile_X3Y3_W2BEG;
wire[7:0] Tile_X3Y3_W2BEGb;
wire[15:0] Tile_X3Y3_WW4BEG;
wire[11:0] Tile_X3Y3_W6BEG;
wire[0:0] Tile_X3Y3_Co;
wire[3:0] Tile_X4Y3_N1BEG;
wire[7:0] Tile_X4Y3_N2BEG;
wire[7:0] Tile_X4Y3_N2BEGb;
wire[15:0] Tile_X4Y3_N4BEG;
wire[15:0] Tile_X4Y3_NN4BEG;
wire[3:0] Tile_X4Y3_E1BEG;
wire[7:0] Tile_X4Y3_E2BEG;
wire[7:0] Tile_X4Y3_E2BEGb;
wire[15:0] Tile_X4Y3_EE4BEG;
wire[11:0] Tile_X4Y3_E6BEG;
wire[3:0] Tile_X4Y3_S1BEG;
wire[7:0] Tile_X4Y3_S2BEG;
wire[7:0] Tile_X4Y3_S2BEGb;
wire[15:0] Tile_X4Y3_S4BEG;
wire[15:0] Tile_X4Y3_SS4BEG;
wire[3:0] Tile_X4Y3_W1BEG;
wire[7:0] Tile_X4Y3_W2BEG;
wire[7:0] Tile_X4Y3_W2BEGb;
wire[15:0] Tile_X4Y3_WW4BEG;
wire[11:0] Tile_X4Y3_W6BEG;
wire[3:0] Tile_X5Y3_N1BEG;
wire[7:0] Tile_X5Y3_N2BEG;
wire[7:0] Tile_X5Y3_N2BEGb;
wire[15:0] Tile_X5Y3_N4BEG;
wire[15:0] Tile_X5Y3_NN4BEG;
wire[3:0] Tile_X5Y3_E1BEG;
wire[7:0] Tile_X5Y3_E2BEG;
wire[7:0] Tile_X5Y3_E2BEGb;
wire[15:0] Tile_X5Y3_EE4BEG;
wire[11:0] Tile_X5Y3_E6BEG;
wire[3:0] Tile_X5Y3_S1BEG;
wire[7:0] Tile_X5Y3_S2BEG;
wire[7:0] Tile_X5Y3_S2BEGb;
wire[15:0] Tile_X5Y3_S4BEG;
wire[15:0] Tile_X5Y3_SS4BEG;
wire[3:0] Tile_X5Y3_W1BEG;
wire[7:0] Tile_X5Y3_W2BEG;
wire[7:0] Tile_X5Y3_W2BEGb;
wire[15:0] Tile_X5Y3_WW4BEG;
wire[11:0] Tile_X5Y3_W6BEG;
wire[0:0] Tile_X5Y3_Co;
wire[3:0] Tile_X6Y3_N1BEG;
wire[7:0] Tile_X6Y3_N2BEG;
wire[7:0] Tile_X6Y3_N2BEGb;
wire[15:0] Tile_X6Y3_N4BEG;
wire[15:0] Tile_X6Y3_NN4BEG;
wire[3:0] Tile_X6Y3_E1BEG;
wire[7:0] Tile_X6Y3_E2BEG;
wire[7:0] Tile_X6Y3_E2BEGb;
wire[15:0] Tile_X6Y3_EE4BEG;
wire[11:0] Tile_X6Y3_E6BEG;
wire[3:0] Tile_X6Y3_S1BEG;
wire[7:0] Tile_X6Y3_S2BEG;
wire[7:0] Tile_X6Y3_S2BEGb;
wire[15:0] Tile_X6Y3_S4BEG;
wire[15:0] Tile_X6Y3_SS4BEG;
wire[3:0] Tile_X6Y3_W1BEG;
wire[7:0] Tile_X6Y3_W2BEG;
wire[7:0] Tile_X6Y3_W2BEGb;
wire[15:0] Tile_X6Y3_WW4BEG;
wire[11:0] Tile_X6Y3_W6BEG;
wire[0:0] Tile_X6Y3_Co;
wire[3:0] Tile_X7Y3_N1BEG;
wire[7:0] Tile_X7Y3_N2BEG;
wire[7:0] Tile_X7Y3_N2BEGb;
wire[15:0] Tile_X7Y3_N4BEG;
wire[15:0] Tile_X7Y3_NN4BEG;
wire[3:0] Tile_X7Y3_E1BEG;
wire[7:0] Tile_X7Y3_E2BEG;
wire[7:0] Tile_X7Y3_E2BEGb;
wire[15:0] Tile_X7Y3_EE4BEG;
wire[11:0] Tile_X7Y3_E6BEG;
wire[3:0] Tile_X7Y3_S1BEG;
wire[7:0] Tile_X7Y3_S2BEG;
wire[7:0] Tile_X7Y3_S2BEGb;
wire[15:0] Tile_X7Y3_S4BEG;
wire[15:0] Tile_X7Y3_SS4BEG;
wire[3:0] Tile_X7Y3_W1BEG;
wire[7:0] Tile_X7Y3_W2BEG;
wire[7:0] Tile_X7Y3_W2BEGb;
wire[15:0] Tile_X7Y3_WW4BEG;
wire[11:0] Tile_X7Y3_W6BEG;
wire[17:0] Tile_X7Y3_top2bot;
wire[3:0] Tile_X8Y3_N1BEG;
wire[7:0] Tile_X8Y3_N2BEG;
wire[7:0] Tile_X8Y3_N2BEGb;
wire[15:0] Tile_X8Y3_N4BEG;
wire[15:0] Tile_X8Y3_NN4BEG;
wire[3:0] Tile_X8Y3_E1BEG;
wire[7:0] Tile_X8Y3_E2BEG;
wire[7:0] Tile_X8Y3_E2BEGb;
wire[15:0] Tile_X8Y3_EE4BEG;
wire[11:0] Tile_X8Y3_E6BEG;
wire[3:0] Tile_X8Y3_S1BEG;
wire[7:0] Tile_X8Y3_S2BEG;
wire[7:0] Tile_X8Y3_S2BEGb;
wire[15:0] Tile_X8Y3_S4BEG;
wire[15:0] Tile_X8Y3_SS4BEG;
wire[3:0] Tile_X8Y3_W1BEG;
wire[7:0] Tile_X8Y3_W2BEG;
wire[7:0] Tile_X8Y3_W2BEGb;
wire[15:0] Tile_X8Y3_WW4BEG;
wire[11:0] Tile_X8Y3_W6BEG;
wire[0:0] Tile_X8Y3_Co;
wire[3:0] Tile_X9Y3_N1BEG;
wire[7:0] Tile_X9Y3_N2BEG;
wire[7:0] Tile_X9Y3_N2BEGb;
wire[15:0] Tile_X9Y3_N4BEG;
wire[15:0] Tile_X9Y3_NN4BEG;
wire[3:0] Tile_X9Y3_E1BEG;
wire[7:0] Tile_X9Y3_E2BEG;
wire[7:0] Tile_X9Y3_E2BEGb;
wire[15:0] Tile_X9Y3_EE4BEG;
wire[11:0] Tile_X9Y3_E6BEG;
wire[3:0] Tile_X9Y3_S1BEG;
wire[7:0] Tile_X9Y3_S2BEG;
wire[7:0] Tile_X9Y3_S2BEGb;
wire[15:0] Tile_X9Y3_S4BEG;
wire[15:0] Tile_X9Y3_SS4BEG;
wire[3:0] Tile_X9Y3_W1BEG;
wire[7:0] Tile_X9Y3_W2BEG;
wire[7:0] Tile_X9Y3_W2BEGb;
wire[15:0] Tile_X9Y3_WW4BEG;
wire[11:0] Tile_X9Y3_W6BEG;
wire[0:0] Tile_X9Y3_Co;
wire[3:0] Tile_X10Y3_N1BEG;
wire[7:0] Tile_X10Y3_N2BEG;
wire[7:0] Tile_X10Y3_N2BEGb;
wire[15:0] Tile_X10Y3_N4BEG;
wire[3:0] Tile_X10Y3_S1BEG;
wire[7:0] Tile_X10Y3_S2BEG;
wire[7:0] Tile_X10Y3_S2BEGb;
wire[15:0] Tile_X10Y3_S4BEG;
wire[3:0] Tile_X10Y3_W1BEG;
wire[7:0] Tile_X10Y3_W2BEG;
wire[7:0] Tile_X10Y3_W2BEGb;
wire[15:0] Tile_X10Y3_WW4BEG;
wire[11:0] Tile_X10Y3_W6BEG;
wire[15:0] Tile_X10Y3_top2bot_DIN;
wire[15:0] Tile_X10Y3_top2bot_BM;
wire[4:0] Tile_X10Y3_top2bot_ADDR;
wire[3:0] Tile_X0Y4_E1BEG;
wire[7:0] Tile_X0Y4_E2BEG;
wire[7:0] Tile_X0Y4_E2BEGb;
wire[15:0] Tile_X0Y4_EE4BEG;
wire[11:0] Tile_X0Y4_E6BEG;
wire[3:0] Tile_X1Y4_N1BEG;
wire[7:0] Tile_X1Y4_N2BEG;
wire[7:0] Tile_X1Y4_N2BEGb;
wire[15:0] Tile_X1Y4_N4BEG;
wire[15:0] Tile_X1Y4_NN4BEG;
wire[3:0] Tile_X1Y4_E1BEG;
wire[7:0] Tile_X1Y4_E2BEG;
wire[7:0] Tile_X1Y4_E2BEGb;
wire[15:0] Tile_X1Y4_EE4BEG;
wire[11:0] Tile_X1Y4_E6BEG;
wire[3:0] Tile_X1Y4_S1BEG;
wire[7:0] Tile_X1Y4_S2BEG;
wire[7:0] Tile_X1Y4_S2BEGb;
wire[15:0] Tile_X1Y4_S4BEG;
wire[15:0] Tile_X1Y4_SS4BEG;
wire[3:0] Tile_X1Y4_W1BEG;
wire[7:0] Tile_X1Y4_W2BEG;
wire[7:0] Tile_X1Y4_W2BEGb;
wire[15:0] Tile_X1Y4_WW4BEG;
wire[11:0] Tile_X1Y4_W6BEG;
wire[0:0] Tile_X1Y4_Co;
wire[3:0] Tile_X2Y4_N1BEG;
wire[7:0] Tile_X2Y4_N2BEG;
wire[7:0] Tile_X2Y4_N2BEGb;
wire[15:0] Tile_X2Y4_N4BEG;
wire[15:0] Tile_X2Y4_NN4BEG;
wire[3:0] Tile_X2Y4_E1BEG;
wire[7:0] Tile_X2Y4_E2BEG;
wire[7:0] Tile_X2Y4_E2BEGb;
wire[15:0] Tile_X2Y4_EE4BEG;
wire[11:0] Tile_X2Y4_E6BEG;
wire[3:0] Tile_X2Y4_S1BEG;
wire[7:0] Tile_X2Y4_S2BEG;
wire[7:0] Tile_X2Y4_S2BEGb;
wire[15:0] Tile_X2Y4_S4BEG;
wire[15:0] Tile_X2Y4_SS4BEG;
wire[3:0] Tile_X2Y4_W1BEG;
wire[7:0] Tile_X2Y4_W2BEG;
wire[7:0] Tile_X2Y4_W2BEGb;
wire[15:0] Tile_X2Y4_WW4BEG;
wire[11:0] Tile_X2Y4_W6BEG;
wire[0:0] Tile_X2Y4_Co;
wire[3:0] Tile_X3Y4_N1BEG;
wire[7:0] Tile_X3Y4_N2BEG;
wire[7:0] Tile_X3Y4_N2BEGb;
wire[15:0] Tile_X3Y4_N4BEG;
wire[15:0] Tile_X3Y4_NN4BEG;
wire[3:0] Tile_X3Y4_E1BEG;
wire[7:0] Tile_X3Y4_E2BEG;
wire[7:0] Tile_X3Y4_E2BEGb;
wire[15:0] Tile_X3Y4_EE4BEG;
wire[11:0] Tile_X3Y4_E6BEG;
wire[3:0] Tile_X3Y4_S1BEG;
wire[7:0] Tile_X3Y4_S2BEG;
wire[7:0] Tile_X3Y4_S2BEGb;
wire[15:0] Tile_X3Y4_S4BEG;
wire[15:0] Tile_X3Y4_SS4BEG;
wire[3:0] Tile_X3Y4_W1BEG;
wire[7:0] Tile_X3Y4_W2BEG;
wire[7:0] Tile_X3Y4_W2BEGb;
wire[15:0] Tile_X3Y4_WW4BEG;
wire[11:0] Tile_X3Y4_W6BEG;
wire[0:0] Tile_X3Y4_Co;
wire[3:0] Tile_X4Y4_N1BEG;
wire[7:0] Tile_X4Y4_N2BEG;
wire[7:0] Tile_X4Y4_N2BEGb;
wire[15:0] Tile_X4Y4_N4BEG;
wire[15:0] Tile_X4Y4_NN4BEG;
wire[3:0] Tile_X4Y4_E1BEG;
wire[7:0] Tile_X4Y4_E2BEG;
wire[7:0] Tile_X4Y4_E2BEGb;
wire[15:0] Tile_X4Y4_EE4BEG;
wire[11:0] Tile_X4Y4_E6BEG;
wire[3:0] Tile_X4Y4_S1BEG;
wire[7:0] Tile_X4Y4_S2BEG;
wire[7:0] Tile_X4Y4_S2BEGb;
wire[15:0] Tile_X4Y4_S4BEG;
wire[15:0] Tile_X4Y4_SS4BEG;
wire[3:0] Tile_X4Y4_W1BEG;
wire[7:0] Tile_X4Y4_W2BEG;
wire[7:0] Tile_X4Y4_W2BEGb;
wire[15:0] Tile_X4Y4_WW4BEG;
wire[11:0] Tile_X4Y4_W6BEG;
wire[3:0] Tile_X5Y4_N1BEG;
wire[7:0] Tile_X5Y4_N2BEG;
wire[7:0] Tile_X5Y4_N2BEGb;
wire[15:0] Tile_X5Y4_N4BEG;
wire[15:0] Tile_X5Y4_NN4BEG;
wire[3:0] Tile_X5Y4_E1BEG;
wire[7:0] Tile_X5Y4_E2BEG;
wire[7:0] Tile_X5Y4_E2BEGb;
wire[15:0] Tile_X5Y4_EE4BEG;
wire[11:0] Tile_X5Y4_E6BEG;
wire[3:0] Tile_X5Y4_S1BEG;
wire[7:0] Tile_X5Y4_S2BEG;
wire[7:0] Tile_X5Y4_S2BEGb;
wire[15:0] Tile_X5Y4_S4BEG;
wire[15:0] Tile_X5Y4_SS4BEG;
wire[3:0] Tile_X5Y4_W1BEG;
wire[7:0] Tile_X5Y4_W2BEG;
wire[7:0] Tile_X5Y4_W2BEGb;
wire[15:0] Tile_X5Y4_WW4BEG;
wire[11:0] Tile_X5Y4_W6BEG;
wire[0:0] Tile_X5Y4_Co;
wire[3:0] Tile_X6Y4_N1BEG;
wire[7:0] Tile_X6Y4_N2BEG;
wire[7:0] Tile_X6Y4_N2BEGb;
wire[15:0] Tile_X6Y4_N4BEG;
wire[15:0] Tile_X6Y4_NN4BEG;
wire[3:0] Tile_X6Y4_E1BEG;
wire[7:0] Tile_X6Y4_E2BEG;
wire[7:0] Tile_X6Y4_E2BEGb;
wire[15:0] Tile_X6Y4_EE4BEG;
wire[11:0] Tile_X6Y4_E6BEG;
wire[3:0] Tile_X6Y4_S1BEG;
wire[7:0] Tile_X6Y4_S2BEG;
wire[7:0] Tile_X6Y4_S2BEGb;
wire[15:0] Tile_X6Y4_S4BEG;
wire[15:0] Tile_X6Y4_SS4BEG;
wire[3:0] Tile_X6Y4_W1BEG;
wire[7:0] Tile_X6Y4_W2BEG;
wire[7:0] Tile_X6Y4_W2BEGb;
wire[15:0] Tile_X6Y4_WW4BEG;
wire[11:0] Tile_X6Y4_W6BEG;
wire[0:0] Tile_X6Y4_Co;
wire[3:0] Tile_X7Y4_N1BEG;
wire[7:0] Tile_X7Y4_N2BEG;
wire[7:0] Tile_X7Y4_N2BEGb;
wire[15:0] Tile_X7Y4_N4BEG;
wire[15:0] Tile_X7Y4_NN4BEG;
wire[3:0] Tile_X7Y4_E1BEG;
wire[7:0] Tile_X7Y4_E2BEG;
wire[7:0] Tile_X7Y4_E2BEGb;
wire[15:0] Tile_X7Y4_EE4BEG;
wire[11:0] Tile_X7Y4_E6BEG;
wire[3:0] Tile_X7Y4_S1BEG;
wire[7:0] Tile_X7Y4_S2BEG;
wire[7:0] Tile_X7Y4_S2BEGb;
wire[15:0] Tile_X7Y4_S4BEG;
wire[15:0] Tile_X7Y4_SS4BEG;
wire[3:0] Tile_X7Y4_W1BEG;
wire[7:0] Tile_X7Y4_W2BEG;
wire[7:0] Tile_X7Y4_W2BEGb;
wire[15:0] Tile_X7Y4_WW4BEG;
wire[11:0] Tile_X7Y4_W6BEG;
wire[9:0] Tile_X7Y4_bot2top;
wire[3:0] Tile_X8Y4_N1BEG;
wire[7:0] Tile_X8Y4_N2BEG;
wire[7:0] Tile_X8Y4_N2BEGb;
wire[15:0] Tile_X8Y4_N4BEG;
wire[15:0] Tile_X8Y4_NN4BEG;
wire[3:0] Tile_X8Y4_E1BEG;
wire[7:0] Tile_X8Y4_E2BEG;
wire[7:0] Tile_X8Y4_E2BEGb;
wire[15:0] Tile_X8Y4_EE4BEG;
wire[11:0] Tile_X8Y4_E6BEG;
wire[3:0] Tile_X8Y4_S1BEG;
wire[7:0] Tile_X8Y4_S2BEG;
wire[7:0] Tile_X8Y4_S2BEGb;
wire[15:0] Tile_X8Y4_S4BEG;
wire[15:0] Tile_X8Y4_SS4BEG;
wire[3:0] Tile_X8Y4_W1BEG;
wire[7:0] Tile_X8Y4_W2BEG;
wire[7:0] Tile_X8Y4_W2BEGb;
wire[15:0] Tile_X8Y4_WW4BEG;
wire[11:0] Tile_X8Y4_W6BEG;
wire[0:0] Tile_X8Y4_Co;
wire[3:0] Tile_X9Y4_N1BEG;
wire[7:0] Tile_X9Y4_N2BEG;
wire[7:0] Tile_X9Y4_N2BEGb;
wire[15:0] Tile_X9Y4_N4BEG;
wire[15:0] Tile_X9Y4_NN4BEG;
wire[3:0] Tile_X9Y4_E1BEG;
wire[7:0] Tile_X9Y4_E2BEG;
wire[7:0] Tile_X9Y4_E2BEGb;
wire[15:0] Tile_X9Y4_EE4BEG;
wire[11:0] Tile_X9Y4_E6BEG;
wire[3:0] Tile_X9Y4_S1BEG;
wire[7:0] Tile_X9Y4_S2BEG;
wire[7:0] Tile_X9Y4_S2BEGb;
wire[15:0] Tile_X9Y4_S4BEG;
wire[15:0] Tile_X9Y4_SS4BEG;
wire[3:0] Tile_X9Y4_W1BEG;
wire[7:0] Tile_X9Y4_W2BEG;
wire[7:0] Tile_X9Y4_W2BEGb;
wire[15:0] Tile_X9Y4_WW4BEG;
wire[11:0] Tile_X9Y4_W6BEG;
wire[0:0] Tile_X9Y4_Co;
wire[3:0] Tile_X10Y4_N1BEG;
wire[7:0] Tile_X10Y4_N2BEG;
wire[7:0] Tile_X10Y4_N2BEGb;
wire[15:0] Tile_X10Y4_N4BEG;
wire[3:0] Tile_X10Y4_S1BEG;
wire[7:0] Tile_X10Y4_S2BEG;
wire[7:0] Tile_X10Y4_S2BEGb;
wire[15:0] Tile_X10Y4_S4BEG;
wire[3:0] Tile_X10Y4_W1BEG;
wire[7:0] Tile_X10Y4_W2BEG;
wire[7:0] Tile_X10Y4_W2BEGb;
wire[15:0] Tile_X10Y4_WW4BEG;
wire[11:0] Tile_X10Y4_W6BEG;
wire[15:0] Tile_X10Y4_bot2top_DOUT;
wire[3:0] Tile_X0Y5_E1BEG;
wire[7:0] Tile_X0Y5_E2BEG;
wire[7:0] Tile_X0Y5_E2BEGb;
wire[15:0] Tile_X0Y5_EE4BEG;
wire[11:0] Tile_X0Y5_E6BEG;
wire[3:0] Tile_X1Y5_N1BEG;
wire[7:0] Tile_X1Y5_N2BEG;
wire[7:0] Tile_X1Y5_N2BEGb;
wire[15:0] Tile_X1Y5_N4BEG;
wire[15:0] Tile_X1Y5_NN4BEG;
wire[3:0] Tile_X1Y5_E1BEG;
wire[7:0] Tile_X1Y5_E2BEG;
wire[7:0] Tile_X1Y5_E2BEGb;
wire[15:0] Tile_X1Y5_EE4BEG;
wire[11:0] Tile_X1Y5_E6BEG;
wire[3:0] Tile_X1Y5_S1BEG;
wire[7:0] Tile_X1Y5_S2BEG;
wire[7:0] Tile_X1Y5_S2BEGb;
wire[15:0] Tile_X1Y5_S4BEG;
wire[15:0] Tile_X1Y5_SS4BEG;
wire[3:0] Tile_X1Y5_W1BEG;
wire[7:0] Tile_X1Y5_W2BEG;
wire[7:0] Tile_X1Y5_W2BEGb;
wire[15:0] Tile_X1Y5_WW4BEG;
wire[11:0] Tile_X1Y5_W6BEG;
wire[0:0] Tile_X1Y5_Co;
wire[3:0] Tile_X2Y5_N1BEG;
wire[7:0] Tile_X2Y5_N2BEG;
wire[7:0] Tile_X2Y5_N2BEGb;
wire[15:0] Tile_X2Y5_N4BEG;
wire[15:0] Tile_X2Y5_NN4BEG;
wire[3:0] Tile_X2Y5_E1BEG;
wire[7:0] Tile_X2Y5_E2BEG;
wire[7:0] Tile_X2Y5_E2BEGb;
wire[15:0] Tile_X2Y5_EE4BEG;
wire[11:0] Tile_X2Y5_E6BEG;
wire[3:0] Tile_X2Y5_S1BEG;
wire[7:0] Tile_X2Y5_S2BEG;
wire[7:0] Tile_X2Y5_S2BEGb;
wire[15:0] Tile_X2Y5_S4BEG;
wire[15:0] Tile_X2Y5_SS4BEG;
wire[3:0] Tile_X2Y5_W1BEG;
wire[7:0] Tile_X2Y5_W2BEG;
wire[7:0] Tile_X2Y5_W2BEGb;
wire[15:0] Tile_X2Y5_WW4BEG;
wire[11:0] Tile_X2Y5_W6BEG;
wire[0:0] Tile_X2Y5_Co;
wire[3:0] Tile_X3Y5_N1BEG;
wire[7:0] Tile_X3Y5_N2BEG;
wire[7:0] Tile_X3Y5_N2BEGb;
wire[15:0] Tile_X3Y5_N4BEG;
wire[15:0] Tile_X3Y5_NN4BEG;
wire[3:0] Tile_X3Y5_E1BEG;
wire[7:0] Tile_X3Y5_E2BEG;
wire[7:0] Tile_X3Y5_E2BEGb;
wire[15:0] Tile_X3Y5_EE4BEG;
wire[11:0] Tile_X3Y5_E6BEG;
wire[3:0] Tile_X3Y5_S1BEG;
wire[7:0] Tile_X3Y5_S2BEG;
wire[7:0] Tile_X3Y5_S2BEGb;
wire[15:0] Tile_X3Y5_S4BEG;
wire[15:0] Tile_X3Y5_SS4BEG;
wire[3:0] Tile_X3Y5_W1BEG;
wire[7:0] Tile_X3Y5_W2BEG;
wire[7:0] Tile_X3Y5_W2BEGb;
wire[15:0] Tile_X3Y5_WW4BEG;
wire[11:0] Tile_X3Y5_W6BEG;
wire[0:0] Tile_X3Y5_Co;
wire[3:0] Tile_X4Y5_N1BEG;
wire[7:0] Tile_X4Y5_N2BEG;
wire[7:0] Tile_X4Y5_N2BEGb;
wire[15:0] Tile_X4Y5_N4BEG;
wire[15:0] Tile_X4Y5_NN4BEG;
wire[3:0] Tile_X4Y5_E1BEG;
wire[7:0] Tile_X4Y5_E2BEG;
wire[7:0] Tile_X4Y5_E2BEGb;
wire[15:0] Tile_X4Y5_EE4BEG;
wire[11:0] Tile_X4Y5_E6BEG;
wire[3:0] Tile_X4Y5_S1BEG;
wire[7:0] Tile_X4Y5_S2BEG;
wire[7:0] Tile_X4Y5_S2BEGb;
wire[15:0] Tile_X4Y5_S4BEG;
wire[15:0] Tile_X4Y5_SS4BEG;
wire[3:0] Tile_X4Y5_W1BEG;
wire[7:0] Tile_X4Y5_W2BEG;
wire[7:0] Tile_X4Y5_W2BEGb;
wire[15:0] Tile_X4Y5_WW4BEG;
wire[11:0] Tile_X4Y5_W6BEG;
wire[3:0] Tile_X5Y5_N1BEG;
wire[7:0] Tile_X5Y5_N2BEG;
wire[7:0] Tile_X5Y5_N2BEGb;
wire[15:0] Tile_X5Y5_N4BEG;
wire[15:0] Tile_X5Y5_NN4BEG;
wire[3:0] Tile_X5Y5_E1BEG;
wire[7:0] Tile_X5Y5_E2BEG;
wire[7:0] Tile_X5Y5_E2BEGb;
wire[15:0] Tile_X5Y5_EE4BEG;
wire[11:0] Tile_X5Y5_E6BEG;
wire[3:0] Tile_X5Y5_S1BEG;
wire[7:0] Tile_X5Y5_S2BEG;
wire[7:0] Tile_X5Y5_S2BEGb;
wire[15:0] Tile_X5Y5_S4BEG;
wire[15:0] Tile_X5Y5_SS4BEG;
wire[3:0] Tile_X5Y5_W1BEG;
wire[7:0] Tile_X5Y5_W2BEG;
wire[7:0] Tile_X5Y5_W2BEGb;
wire[15:0] Tile_X5Y5_WW4BEG;
wire[11:0] Tile_X5Y5_W6BEG;
wire[0:0] Tile_X5Y5_Co;
wire[3:0] Tile_X6Y5_N1BEG;
wire[7:0] Tile_X6Y5_N2BEG;
wire[7:0] Tile_X6Y5_N2BEGb;
wire[15:0] Tile_X6Y5_N4BEG;
wire[15:0] Tile_X6Y5_NN4BEG;
wire[3:0] Tile_X6Y5_E1BEG;
wire[7:0] Tile_X6Y5_E2BEG;
wire[7:0] Tile_X6Y5_E2BEGb;
wire[15:0] Tile_X6Y5_EE4BEG;
wire[11:0] Tile_X6Y5_E6BEG;
wire[3:0] Tile_X6Y5_S1BEG;
wire[7:0] Tile_X6Y5_S2BEG;
wire[7:0] Tile_X6Y5_S2BEGb;
wire[15:0] Tile_X6Y5_S4BEG;
wire[15:0] Tile_X6Y5_SS4BEG;
wire[3:0] Tile_X6Y5_W1BEG;
wire[7:0] Tile_X6Y5_W2BEG;
wire[7:0] Tile_X6Y5_W2BEGb;
wire[15:0] Tile_X6Y5_WW4BEG;
wire[11:0] Tile_X6Y5_W6BEG;
wire[0:0] Tile_X6Y5_Co;
wire[3:0] Tile_X7Y5_N1BEG;
wire[7:0] Tile_X7Y5_N2BEG;
wire[7:0] Tile_X7Y5_N2BEGb;
wire[15:0] Tile_X7Y5_N4BEG;
wire[15:0] Tile_X7Y5_NN4BEG;
wire[3:0] Tile_X7Y5_E1BEG;
wire[7:0] Tile_X7Y5_E2BEG;
wire[7:0] Tile_X7Y5_E2BEGb;
wire[15:0] Tile_X7Y5_EE4BEG;
wire[11:0] Tile_X7Y5_E6BEG;
wire[3:0] Tile_X7Y5_S1BEG;
wire[7:0] Tile_X7Y5_S2BEG;
wire[7:0] Tile_X7Y5_S2BEGb;
wire[15:0] Tile_X7Y5_S4BEG;
wire[15:0] Tile_X7Y5_SS4BEG;
wire[3:0] Tile_X7Y5_W1BEG;
wire[7:0] Tile_X7Y5_W2BEG;
wire[7:0] Tile_X7Y5_W2BEGb;
wire[15:0] Tile_X7Y5_WW4BEG;
wire[11:0] Tile_X7Y5_W6BEG;
wire[17:0] Tile_X7Y5_top2bot;
wire[3:0] Tile_X8Y5_N1BEG;
wire[7:0] Tile_X8Y5_N2BEG;
wire[7:0] Tile_X8Y5_N2BEGb;
wire[15:0] Tile_X8Y5_N4BEG;
wire[15:0] Tile_X8Y5_NN4BEG;
wire[3:0] Tile_X8Y5_E1BEG;
wire[7:0] Tile_X8Y5_E2BEG;
wire[7:0] Tile_X8Y5_E2BEGb;
wire[15:0] Tile_X8Y5_EE4BEG;
wire[11:0] Tile_X8Y5_E6BEG;
wire[3:0] Tile_X8Y5_S1BEG;
wire[7:0] Tile_X8Y5_S2BEG;
wire[7:0] Tile_X8Y5_S2BEGb;
wire[15:0] Tile_X8Y5_S4BEG;
wire[15:0] Tile_X8Y5_SS4BEG;
wire[3:0] Tile_X8Y5_W1BEG;
wire[7:0] Tile_X8Y5_W2BEG;
wire[7:0] Tile_X8Y5_W2BEGb;
wire[15:0] Tile_X8Y5_WW4BEG;
wire[11:0] Tile_X8Y5_W6BEG;
wire[0:0] Tile_X8Y5_Co;
wire[3:0] Tile_X9Y5_N1BEG;
wire[7:0] Tile_X9Y5_N2BEG;
wire[7:0] Tile_X9Y5_N2BEGb;
wire[15:0] Tile_X9Y5_N4BEG;
wire[15:0] Tile_X9Y5_NN4BEG;
wire[3:0] Tile_X9Y5_E1BEG;
wire[7:0] Tile_X9Y5_E2BEG;
wire[7:0] Tile_X9Y5_E2BEGb;
wire[15:0] Tile_X9Y5_EE4BEG;
wire[11:0] Tile_X9Y5_E6BEG;
wire[3:0] Tile_X9Y5_S1BEG;
wire[7:0] Tile_X9Y5_S2BEG;
wire[7:0] Tile_X9Y5_S2BEGb;
wire[15:0] Tile_X9Y5_S4BEG;
wire[15:0] Tile_X9Y5_SS4BEG;
wire[3:0] Tile_X9Y5_W1BEG;
wire[7:0] Tile_X9Y5_W2BEG;
wire[7:0] Tile_X9Y5_W2BEGb;
wire[15:0] Tile_X9Y5_WW4BEG;
wire[11:0] Tile_X9Y5_W6BEG;
wire[0:0] Tile_X9Y5_Co;
wire[3:0] Tile_X10Y5_N1BEG;
wire[7:0] Tile_X10Y5_N2BEG;
wire[7:0] Tile_X10Y5_N2BEGb;
wire[15:0] Tile_X10Y5_N4BEG;
wire[3:0] Tile_X10Y5_S1BEG;
wire[7:0] Tile_X10Y5_S2BEG;
wire[7:0] Tile_X10Y5_S2BEGb;
wire[15:0] Tile_X10Y5_S4BEG;
wire[3:0] Tile_X10Y5_W1BEG;
wire[7:0] Tile_X10Y5_W2BEG;
wire[7:0] Tile_X10Y5_W2BEGb;
wire[15:0] Tile_X10Y5_WW4BEG;
wire[11:0] Tile_X10Y5_W6BEG;
wire[15:0] Tile_X10Y5_top2bot_DIN;
wire[15:0] Tile_X10Y5_top2bot_BM;
wire[4:0] Tile_X10Y5_top2bot_ADDR;
wire[3:0] Tile_X0Y6_E1BEG;
wire[7:0] Tile_X0Y6_E2BEG;
wire[7:0] Tile_X0Y6_E2BEGb;
wire[15:0] Tile_X0Y6_EE4BEG;
wire[11:0] Tile_X0Y6_E6BEG;
wire[3:0] Tile_X1Y6_N1BEG;
wire[7:0] Tile_X1Y6_N2BEG;
wire[7:0] Tile_X1Y6_N2BEGb;
wire[15:0] Tile_X1Y6_N4BEG;
wire[15:0] Tile_X1Y6_NN4BEG;
wire[3:0] Tile_X1Y6_E1BEG;
wire[7:0] Tile_X1Y6_E2BEG;
wire[7:0] Tile_X1Y6_E2BEGb;
wire[15:0] Tile_X1Y6_EE4BEG;
wire[11:0] Tile_X1Y6_E6BEG;
wire[3:0] Tile_X1Y6_S1BEG;
wire[7:0] Tile_X1Y6_S2BEG;
wire[7:0] Tile_X1Y6_S2BEGb;
wire[15:0] Tile_X1Y6_S4BEG;
wire[15:0] Tile_X1Y6_SS4BEG;
wire[3:0] Tile_X1Y6_W1BEG;
wire[7:0] Tile_X1Y6_W2BEG;
wire[7:0] Tile_X1Y6_W2BEGb;
wire[15:0] Tile_X1Y6_WW4BEG;
wire[11:0] Tile_X1Y6_W6BEG;
wire[0:0] Tile_X1Y6_Co;
wire[3:0] Tile_X2Y6_N1BEG;
wire[7:0] Tile_X2Y6_N2BEG;
wire[7:0] Tile_X2Y6_N2BEGb;
wire[15:0] Tile_X2Y6_N4BEG;
wire[15:0] Tile_X2Y6_NN4BEG;
wire[3:0] Tile_X2Y6_E1BEG;
wire[7:0] Tile_X2Y6_E2BEG;
wire[7:0] Tile_X2Y6_E2BEGb;
wire[15:0] Tile_X2Y6_EE4BEG;
wire[11:0] Tile_X2Y6_E6BEG;
wire[3:0] Tile_X2Y6_S1BEG;
wire[7:0] Tile_X2Y6_S2BEG;
wire[7:0] Tile_X2Y6_S2BEGb;
wire[15:0] Tile_X2Y6_S4BEG;
wire[15:0] Tile_X2Y6_SS4BEG;
wire[3:0] Tile_X2Y6_W1BEG;
wire[7:0] Tile_X2Y6_W2BEG;
wire[7:0] Tile_X2Y6_W2BEGb;
wire[15:0] Tile_X2Y6_WW4BEG;
wire[11:0] Tile_X2Y6_W6BEG;
wire[0:0] Tile_X2Y6_Co;
wire[3:0] Tile_X3Y6_N1BEG;
wire[7:0] Tile_X3Y6_N2BEG;
wire[7:0] Tile_X3Y6_N2BEGb;
wire[15:0] Tile_X3Y6_N4BEG;
wire[15:0] Tile_X3Y6_NN4BEG;
wire[3:0] Tile_X3Y6_E1BEG;
wire[7:0] Tile_X3Y6_E2BEG;
wire[7:0] Tile_X3Y6_E2BEGb;
wire[15:0] Tile_X3Y6_EE4BEG;
wire[11:0] Tile_X3Y6_E6BEG;
wire[3:0] Tile_X3Y6_S1BEG;
wire[7:0] Tile_X3Y6_S2BEG;
wire[7:0] Tile_X3Y6_S2BEGb;
wire[15:0] Tile_X3Y6_S4BEG;
wire[15:0] Tile_X3Y6_SS4BEG;
wire[3:0] Tile_X3Y6_W1BEG;
wire[7:0] Tile_X3Y6_W2BEG;
wire[7:0] Tile_X3Y6_W2BEGb;
wire[15:0] Tile_X3Y6_WW4BEG;
wire[11:0] Tile_X3Y6_W6BEG;
wire[0:0] Tile_X3Y6_Co;
wire[3:0] Tile_X4Y6_N1BEG;
wire[7:0] Tile_X4Y6_N2BEG;
wire[7:0] Tile_X4Y6_N2BEGb;
wire[15:0] Tile_X4Y6_N4BEG;
wire[15:0] Tile_X4Y6_NN4BEG;
wire[3:0] Tile_X4Y6_E1BEG;
wire[7:0] Tile_X4Y6_E2BEG;
wire[7:0] Tile_X4Y6_E2BEGb;
wire[15:0] Tile_X4Y6_EE4BEG;
wire[11:0] Tile_X4Y6_E6BEG;
wire[3:0] Tile_X4Y6_S1BEG;
wire[7:0] Tile_X4Y6_S2BEG;
wire[7:0] Tile_X4Y6_S2BEGb;
wire[15:0] Tile_X4Y6_S4BEG;
wire[15:0] Tile_X4Y6_SS4BEG;
wire[3:0] Tile_X4Y6_W1BEG;
wire[7:0] Tile_X4Y6_W2BEG;
wire[7:0] Tile_X4Y6_W2BEGb;
wire[15:0] Tile_X4Y6_WW4BEG;
wire[11:0] Tile_X4Y6_W6BEG;
wire[3:0] Tile_X5Y6_N1BEG;
wire[7:0] Tile_X5Y6_N2BEG;
wire[7:0] Tile_X5Y6_N2BEGb;
wire[15:0] Tile_X5Y6_N4BEG;
wire[15:0] Tile_X5Y6_NN4BEG;
wire[3:0] Tile_X5Y6_E1BEG;
wire[7:0] Tile_X5Y6_E2BEG;
wire[7:0] Tile_X5Y6_E2BEGb;
wire[15:0] Tile_X5Y6_EE4BEG;
wire[11:0] Tile_X5Y6_E6BEG;
wire[3:0] Tile_X5Y6_S1BEG;
wire[7:0] Tile_X5Y6_S2BEG;
wire[7:0] Tile_X5Y6_S2BEGb;
wire[15:0] Tile_X5Y6_S4BEG;
wire[15:0] Tile_X5Y6_SS4BEG;
wire[3:0] Tile_X5Y6_W1BEG;
wire[7:0] Tile_X5Y6_W2BEG;
wire[7:0] Tile_X5Y6_W2BEGb;
wire[15:0] Tile_X5Y6_WW4BEG;
wire[11:0] Tile_X5Y6_W6BEG;
wire[0:0] Tile_X5Y6_Co;
wire[3:0] Tile_X6Y6_N1BEG;
wire[7:0] Tile_X6Y6_N2BEG;
wire[7:0] Tile_X6Y6_N2BEGb;
wire[15:0] Tile_X6Y6_N4BEG;
wire[15:0] Tile_X6Y6_NN4BEG;
wire[3:0] Tile_X6Y6_E1BEG;
wire[7:0] Tile_X6Y6_E2BEG;
wire[7:0] Tile_X6Y6_E2BEGb;
wire[15:0] Tile_X6Y6_EE4BEG;
wire[11:0] Tile_X6Y6_E6BEG;
wire[3:0] Tile_X6Y6_S1BEG;
wire[7:0] Tile_X6Y6_S2BEG;
wire[7:0] Tile_X6Y6_S2BEGb;
wire[15:0] Tile_X6Y6_S4BEG;
wire[15:0] Tile_X6Y6_SS4BEG;
wire[3:0] Tile_X6Y6_W1BEG;
wire[7:0] Tile_X6Y6_W2BEG;
wire[7:0] Tile_X6Y6_W2BEGb;
wire[15:0] Tile_X6Y6_WW4BEG;
wire[11:0] Tile_X6Y6_W6BEG;
wire[0:0] Tile_X6Y6_Co;
wire[3:0] Tile_X7Y6_N1BEG;
wire[7:0] Tile_X7Y6_N2BEG;
wire[7:0] Tile_X7Y6_N2BEGb;
wire[15:0] Tile_X7Y6_N4BEG;
wire[15:0] Tile_X7Y6_NN4BEG;
wire[3:0] Tile_X7Y6_E1BEG;
wire[7:0] Tile_X7Y6_E2BEG;
wire[7:0] Tile_X7Y6_E2BEGb;
wire[15:0] Tile_X7Y6_EE4BEG;
wire[11:0] Tile_X7Y6_E6BEG;
wire[3:0] Tile_X7Y6_S1BEG;
wire[7:0] Tile_X7Y6_S2BEG;
wire[7:0] Tile_X7Y6_S2BEGb;
wire[15:0] Tile_X7Y6_S4BEG;
wire[15:0] Tile_X7Y6_SS4BEG;
wire[3:0] Tile_X7Y6_W1BEG;
wire[7:0] Tile_X7Y6_W2BEG;
wire[7:0] Tile_X7Y6_W2BEGb;
wire[15:0] Tile_X7Y6_WW4BEG;
wire[11:0] Tile_X7Y6_W6BEG;
wire[9:0] Tile_X7Y6_bot2top;
wire[3:0] Tile_X8Y6_N1BEG;
wire[7:0] Tile_X8Y6_N2BEG;
wire[7:0] Tile_X8Y6_N2BEGb;
wire[15:0] Tile_X8Y6_N4BEG;
wire[15:0] Tile_X8Y6_NN4BEG;
wire[3:0] Tile_X8Y6_E1BEG;
wire[7:0] Tile_X8Y6_E2BEG;
wire[7:0] Tile_X8Y6_E2BEGb;
wire[15:0] Tile_X8Y6_EE4BEG;
wire[11:0] Tile_X8Y6_E6BEG;
wire[3:0] Tile_X8Y6_S1BEG;
wire[7:0] Tile_X8Y6_S2BEG;
wire[7:0] Tile_X8Y6_S2BEGb;
wire[15:0] Tile_X8Y6_S4BEG;
wire[15:0] Tile_X8Y6_SS4BEG;
wire[3:0] Tile_X8Y6_W1BEG;
wire[7:0] Tile_X8Y6_W2BEG;
wire[7:0] Tile_X8Y6_W2BEGb;
wire[15:0] Tile_X8Y6_WW4BEG;
wire[11:0] Tile_X8Y6_W6BEG;
wire[0:0] Tile_X8Y6_Co;
wire[3:0] Tile_X9Y6_N1BEG;
wire[7:0] Tile_X9Y6_N2BEG;
wire[7:0] Tile_X9Y6_N2BEGb;
wire[15:0] Tile_X9Y6_N4BEG;
wire[15:0] Tile_X9Y6_NN4BEG;
wire[3:0] Tile_X9Y6_E1BEG;
wire[7:0] Tile_X9Y6_E2BEG;
wire[7:0] Tile_X9Y6_E2BEGb;
wire[15:0] Tile_X9Y6_EE4BEG;
wire[11:0] Tile_X9Y6_E6BEG;
wire[3:0] Tile_X9Y6_S1BEG;
wire[7:0] Tile_X9Y6_S2BEG;
wire[7:0] Tile_X9Y6_S2BEGb;
wire[15:0] Tile_X9Y6_S4BEG;
wire[15:0] Tile_X9Y6_SS4BEG;
wire[3:0] Tile_X9Y6_W1BEG;
wire[7:0] Tile_X9Y6_W2BEG;
wire[7:0] Tile_X9Y6_W2BEGb;
wire[15:0] Tile_X9Y6_WW4BEG;
wire[11:0] Tile_X9Y6_W6BEG;
wire[0:0] Tile_X9Y6_Co;
wire[3:0] Tile_X10Y6_N1BEG;
wire[7:0] Tile_X10Y6_N2BEG;
wire[7:0] Tile_X10Y6_N2BEGb;
wire[15:0] Tile_X10Y6_N4BEG;
wire[3:0] Tile_X10Y6_S1BEG;
wire[7:0] Tile_X10Y6_S2BEG;
wire[7:0] Tile_X10Y6_S2BEGb;
wire[15:0] Tile_X10Y6_S4BEG;
wire[3:0] Tile_X10Y6_W1BEG;
wire[7:0] Tile_X10Y6_W2BEG;
wire[7:0] Tile_X10Y6_W2BEGb;
wire[15:0] Tile_X10Y6_WW4BEG;
wire[11:0] Tile_X10Y6_W6BEG;
wire[15:0] Tile_X10Y6_bot2top_DOUT;
wire[3:0] Tile_X0Y7_E1BEG;
wire[7:0] Tile_X0Y7_E2BEG;
wire[7:0] Tile_X0Y7_E2BEGb;
wire[15:0] Tile_X0Y7_EE4BEG;
wire[11:0] Tile_X0Y7_E6BEG;
wire[3:0] Tile_X1Y7_N1BEG;
wire[7:0] Tile_X1Y7_N2BEG;
wire[7:0] Tile_X1Y7_N2BEGb;
wire[15:0] Tile_X1Y7_N4BEG;
wire[15:0] Tile_X1Y7_NN4BEG;
wire[3:0] Tile_X1Y7_E1BEG;
wire[7:0] Tile_X1Y7_E2BEG;
wire[7:0] Tile_X1Y7_E2BEGb;
wire[15:0] Tile_X1Y7_EE4BEG;
wire[11:0] Tile_X1Y7_E6BEG;
wire[3:0] Tile_X1Y7_S1BEG;
wire[7:0] Tile_X1Y7_S2BEG;
wire[7:0] Tile_X1Y7_S2BEGb;
wire[15:0] Tile_X1Y7_S4BEG;
wire[15:0] Tile_X1Y7_SS4BEG;
wire[3:0] Tile_X1Y7_W1BEG;
wire[7:0] Tile_X1Y7_W2BEG;
wire[7:0] Tile_X1Y7_W2BEGb;
wire[15:0] Tile_X1Y7_WW4BEG;
wire[11:0] Tile_X1Y7_W6BEG;
wire[0:0] Tile_X1Y7_Co;
wire[3:0] Tile_X2Y7_N1BEG;
wire[7:0] Tile_X2Y7_N2BEG;
wire[7:0] Tile_X2Y7_N2BEGb;
wire[15:0] Tile_X2Y7_N4BEG;
wire[15:0] Tile_X2Y7_NN4BEG;
wire[3:0] Tile_X2Y7_E1BEG;
wire[7:0] Tile_X2Y7_E2BEG;
wire[7:0] Tile_X2Y7_E2BEGb;
wire[15:0] Tile_X2Y7_EE4BEG;
wire[11:0] Tile_X2Y7_E6BEG;
wire[3:0] Tile_X2Y7_S1BEG;
wire[7:0] Tile_X2Y7_S2BEG;
wire[7:0] Tile_X2Y7_S2BEGb;
wire[15:0] Tile_X2Y7_S4BEG;
wire[15:0] Tile_X2Y7_SS4BEG;
wire[3:0] Tile_X2Y7_W1BEG;
wire[7:0] Tile_X2Y7_W2BEG;
wire[7:0] Tile_X2Y7_W2BEGb;
wire[15:0] Tile_X2Y7_WW4BEG;
wire[11:0] Tile_X2Y7_W6BEG;
wire[0:0] Tile_X2Y7_Co;
wire[3:0] Tile_X3Y7_N1BEG;
wire[7:0] Tile_X3Y7_N2BEG;
wire[7:0] Tile_X3Y7_N2BEGb;
wire[15:0] Tile_X3Y7_N4BEG;
wire[15:0] Tile_X3Y7_NN4BEG;
wire[3:0] Tile_X3Y7_E1BEG;
wire[7:0] Tile_X3Y7_E2BEG;
wire[7:0] Tile_X3Y7_E2BEGb;
wire[15:0] Tile_X3Y7_EE4BEG;
wire[11:0] Tile_X3Y7_E6BEG;
wire[3:0] Tile_X3Y7_S1BEG;
wire[7:0] Tile_X3Y7_S2BEG;
wire[7:0] Tile_X3Y7_S2BEGb;
wire[15:0] Tile_X3Y7_S4BEG;
wire[15:0] Tile_X3Y7_SS4BEG;
wire[3:0] Tile_X3Y7_W1BEG;
wire[7:0] Tile_X3Y7_W2BEG;
wire[7:0] Tile_X3Y7_W2BEGb;
wire[15:0] Tile_X3Y7_WW4BEG;
wire[11:0] Tile_X3Y7_W6BEG;
wire[0:0] Tile_X3Y7_Co;
wire[3:0] Tile_X4Y7_N1BEG;
wire[7:0] Tile_X4Y7_N2BEG;
wire[7:0] Tile_X4Y7_N2BEGb;
wire[15:0] Tile_X4Y7_N4BEG;
wire[15:0] Tile_X4Y7_NN4BEG;
wire[3:0] Tile_X4Y7_E1BEG;
wire[7:0] Tile_X4Y7_E2BEG;
wire[7:0] Tile_X4Y7_E2BEGb;
wire[15:0] Tile_X4Y7_EE4BEG;
wire[11:0] Tile_X4Y7_E6BEG;
wire[3:0] Tile_X4Y7_S1BEG;
wire[7:0] Tile_X4Y7_S2BEG;
wire[7:0] Tile_X4Y7_S2BEGb;
wire[15:0] Tile_X4Y7_S4BEG;
wire[15:0] Tile_X4Y7_SS4BEG;
wire[3:0] Tile_X4Y7_W1BEG;
wire[7:0] Tile_X4Y7_W2BEG;
wire[7:0] Tile_X4Y7_W2BEGb;
wire[15:0] Tile_X4Y7_WW4BEG;
wire[11:0] Tile_X4Y7_W6BEG;
wire[3:0] Tile_X5Y7_N1BEG;
wire[7:0] Tile_X5Y7_N2BEG;
wire[7:0] Tile_X5Y7_N2BEGb;
wire[15:0] Tile_X5Y7_N4BEG;
wire[15:0] Tile_X5Y7_NN4BEG;
wire[3:0] Tile_X5Y7_E1BEG;
wire[7:0] Tile_X5Y7_E2BEG;
wire[7:0] Tile_X5Y7_E2BEGb;
wire[15:0] Tile_X5Y7_EE4BEG;
wire[11:0] Tile_X5Y7_E6BEG;
wire[3:0] Tile_X5Y7_S1BEG;
wire[7:0] Tile_X5Y7_S2BEG;
wire[7:0] Tile_X5Y7_S2BEGb;
wire[15:0] Tile_X5Y7_S4BEG;
wire[15:0] Tile_X5Y7_SS4BEG;
wire[3:0] Tile_X5Y7_W1BEG;
wire[7:0] Tile_X5Y7_W2BEG;
wire[7:0] Tile_X5Y7_W2BEGb;
wire[15:0] Tile_X5Y7_WW4BEG;
wire[11:0] Tile_X5Y7_W6BEG;
wire[0:0] Tile_X5Y7_Co;
wire[3:0] Tile_X6Y7_N1BEG;
wire[7:0] Tile_X6Y7_N2BEG;
wire[7:0] Tile_X6Y7_N2BEGb;
wire[15:0] Tile_X6Y7_N4BEG;
wire[15:0] Tile_X6Y7_NN4BEG;
wire[3:0] Tile_X6Y7_E1BEG;
wire[7:0] Tile_X6Y7_E2BEG;
wire[7:0] Tile_X6Y7_E2BEGb;
wire[15:0] Tile_X6Y7_EE4BEG;
wire[11:0] Tile_X6Y7_E6BEG;
wire[3:0] Tile_X6Y7_S1BEG;
wire[7:0] Tile_X6Y7_S2BEG;
wire[7:0] Tile_X6Y7_S2BEGb;
wire[15:0] Tile_X6Y7_S4BEG;
wire[15:0] Tile_X6Y7_SS4BEG;
wire[3:0] Tile_X6Y7_W1BEG;
wire[7:0] Tile_X6Y7_W2BEG;
wire[7:0] Tile_X6Y7_W2BEGb;
wire[15:0] Tile_X6Y7_WW4BEG;
wire[11:0] Tile_X6Y7_W6BEG;
wire[0:0] Tile_X6Y7_Co;
wire[3:0] Tile_X7Y7_N1BEG;
wire[7:0] Tile_X7Y7_N2BEG;
wire[7:0] Tile_X7Y7_N2BEGb;
wire[15:0] Tile_X7Y7_N4BEG;
wire[15:0] Tile_X7Y7_NN4BEG;
wire[3:0] Tile_X7Y7_E1BEG;
wire[7:0] Tile_X7Y7_E2BEG;
wire[7:0] Tile_X7Y7_E2BEGb;
wire[15:0] Tile_X7Y7_EE4BEG;
wire[11:0] Tile_X7Y7_E6BEG;
wire[3:0] Tile_X7Y7_S1BEG;
wire[7:0] Tile_X7Y7_S2BEG;
wire[7:0] Tile_X7Y7_S2BEGb;
wire[15:0] Tile_X7Y7_S4BEG;
wire[15:0] Tile_X7Y7_SS4BEG;
wire[3:0] Tile_X7Y7_W1BEG;
wire[7:0] Tile_X7Y7_W2BEG;
wire[7:0] Tile_X7Y7_W2BEGb;
wire[15:0] Tile_X7Y7_WW4BEG;
wire[11:0] Tile_X7Y7_W6BEG;
wire[17:0] Tile_X7Y7_top2bot;
wire[3:0] Tile_X8Y7_N1BEG;
wire[7:0] Tile_X8Y7_N2BEG;
wire[7:0] Tile_X8Y7_N2BEGb;
wire[15:0] Tile_X8Y7_N4BEG;
wire[15:0] Tile_X8Y7_NN4BEG;
wire[3:0] Tile_X8Y7_E1BEG;
wire[7:0] Tile_X8Y7_E2BEG;
wire[7:0] Tile_X8Y7_E2BEGb;
wire[15:0] Tile_X8Y7_EE4BEG;
wire[11:0] Tile_X8Y7_E6BEG;
wire[3:0] Tile_X8Y7_S1BEG;
wire[7:0] Tile_X8Y7_S2BEG;
wire[7:0] Tile_X8Y7_S2BEGb;
wire[15:0] Tile_X8Y7_S4BEG;
wire[15:0] Tile_X8Y7_SS4BEG;
wire[3:0] Tile_X8Y7_W1BEG;
wire[7:0] Tile_X8Y7_W2BEG;
wire[7:0] Tile_X8Y7_W2BEGb;
wire[15:0] Tile_X8Y7_WW4BEG;
wire[11:0] Tile_X8Y7_W6BEG;
wire[0:0] Tile_X8Y7_Co;
wire[3:0] Tile_X9Y7_N1BEG;
wire[7:0] Tile_X9Y7_N2BEG;
wire[7:0] Tile_X9Y7_N2BEGb;
wire[15:0] Tile_X9Y7_N4BEG;
wire[15:0] Tile_X9Y7_NN4BEG;
wire[3:0] Tile_X9Y7_E1BEG;
wire[7:0] Tile_X9Y7_E2BEG;
wire[7:0] Tile_X9Y7_E2BEGb;
wire[15:0] Tile_X9Y7_EE4BEG;
wire[11:0] Tile_X9Y7_E6BEG;
wire[3:0] Tile_X9Y7_S1BEG;
wire[7:0] Tile_X9Y7_S2BEG;
wire[7:0] Tile_X9Y7_S2BEGb;
wire[15:0] Tile_X9Y7_S4BEG;
wire[15:0] Tile_X9Y7_SS4BEG;
wire[3:0] Tile_X9Y7_W1BEG;
wire[7:0] Tile_X9Y7_W2BEG;
wire[7:0] Tile_X9Y7_W2BEGb;
wire[15:0] Tile_X9Y7_WW4BEG;
wire[11:0] Tile_X9Y7_W6BEG;
wire[0:0] Tile_X9Y7_Co;
wire[3:0] Tile_X10Y7_N1BEG;
wire[7:0] Tile_X10Y7_N2BEG;
wire[7:0] Tile_X10Y7_N2BEGb;
wire[15:0] Tile_X10Y7_N4BEG;
wire[3:0] Tile_X10Y7_S1BEG;
wire[7:0] Tile_X10Y7_S2BEG;
wire[7:0] Tile_X10Y7_S2BEGb;
wire[15:0] Tile_X10Y7_S4BEG;
wire[3:0] Tile_X10Y7_W1BEG;
wire[7:0] Tile_X10Y7_W2BEG;
wire[7:0] Tile_X10Y7_W2BEGb;
wire[15:0] Tile_X10Y7_WW4BEG;
wire[11:0] Tile_X10Y7_W6BEG;
wire[15:0] Tile_X10Y7_top2bot_DIN;
wire[15:0] Tile_X10Y7_top2bot_BM;
wire[4:0] Tile_X10Y7_top2bot_ADDR;
wire[3:0] Tile_X0Y8_E1BEG;
wire[7:0] Tile_X0Y8_E2BEG;
wire[7:0] Tile_X0Y8_E2BEGb;
wire[15:0] Tile_X0Y8_EE4BEG;
wire[11:0] Tile_X0Y8_E6BEG;
wire[3:0] Tile_X1Y8_N1BEG;
wire[7:0] Tile_X1Y8_N2BEG;
wire[7:0] Tile_X1Y8_N2BEGb;
wire[15:0] Tile_X1Y8_N4BEG;
wire[15:0] Tile_X1Y8_NN4BEG;
wire[3:0] Tile_X1Y8_E1BEG;
wire[7:0] Tile_X1Y8_E2BEG;
wire[7:0] Tile_X1Y8_E2BEGb;
wire[15:0] Tile_X1Y8_EE4BEG;
wire[11:0] Tile_X1Y8_E6BEG;
wire[3:0] Tile_X1Y8_S1BEG;
wire[7:0] Tile_X1Y8_S2BEG;
wire[7:0] Tile_X1Y8_S2BEGb;
wire[15:0] Tile_X1Y8_S4BEG;
wire[15:0] Tile_X1Y8_SS4BEG;
wire[3:0] Tile_X1Y8_W1BEG;
wire[7:0] Tile_X1Y8_W2BEG;
wire[7:0] Tile_X1Y8_W2BEGb;
wire[15:0] Tile_X1Y8_WW4BEG;
wire[11:0] Tile_X1Y8_W6BEG;
wire[0:0] Tile_X1Y8_Co;
wire[3:0] Tile_X2Y8_N1BEG;
wire[7:0] Tile_X2Y8_N2BEG;
wire[7:0] Tile_X2Y8_N2BEGb;
wire[15:0] Tile_X2Y8_N4BEG;
wire[15:0] Tile_X2Y8_NN4BEG;
wire[3:0] Tile_X2Y8_E1BEG;
wire[7:0] Tile_X2Y8_E2BEG;
wire[7:0] Tile_X2Y8_E2BEGb;
wire[15:0] Tile_X2Y8_EE4BEG;
wire[11:0] Tile_X2Y8_E6BEG;
wire[3:0] Tile_X2Y8_S1BEG;
wire[7:0] Tile_X2Y8_S2BEG;
wire[7:0] Tile_X2Y8_S2BEGb;
wire[15:0] Tile_X2Y8_S4BEG;
wire[15:0] Tile_X2Y8_SS4BEG;
wire[3:0] Tile_X2Y8_W1BEG;
wire[7:0] Tile_X2Y8_W2BEG;
wire[7:0] Tile_X2Y8_W2BEGb;
wire[15:0] Tile_X2Y8_WW4BEG;
wire[11:0] Tile_X2Y8_W6BEG;
wire[0:0] Tile_X2Y8_Co;
wire[3:0] Tile_X3Y8_N1BEG;
wire[7:0] Tile_X3Y8_N2BEG;
wire[7:0] Tile_X3Y8_N2BEGb;
wire[15:0] Tile_X3Y8_N4BEG;
wire[15:0] Tile_X3Y8_NN4BEG;
wire[3:0] Tile_X3Y8_E1BEG;
wire[7:0] Tile_X3Y8_E2BEG;
wire[7:0] Tile_X3Y8_E2BEGb;
wire[15:0] Tile_X3Y8_EE4BEG;
wire[11:0] Tile_X3Y8_E6BEG;
wire[3:0] Tile_X3Y8_S1BEG;
wire[7:0] Tile_X3Y8_S2BEG;
wire[7:0] Tile_X3Y8_S2BEGb;
wire[15:0] Tile_X3Y8_S4BEG;
wire[15:0] Tile_X3Y8_SS4BEG;
wire[3:0] Tile_X3Y8_W1BEG;
wire[7:0] Tile_X3Y8_W2BEG;
wire[7:0] Tile_X3Y8_W2BEGb;
wire[15:0] Tile_X3Y8_WW4BEG;
wire[11:0] Tile_X3Y8_W6BEG;
wire[0:0] Tile_X3Y8_Co;
wire[3:0] Tile_X4Y8_N1BEG;
wire[7:0] Tile_X4Y8_N2BEG;
wire[7:0] Tile_X4Y8_N2BEGb;
wire[15:0] Tile_X4Y8_N4BEG;
wire[15:0] Tile_X4Y8_NN4BEG;
wire[3:0] Tile_X4Y8_E1BEG;
wire[7:0] Tile_X4Y8_E2BEG;
wire[7:0] Tile_X4Y8_E2BEGb;
wire[15:0] Tile_X4Y8_EE4BEG;
wire[11:0] Tile_X4Y8_E6BEG;
wire[3:0] Tile_X4Y8_S1BEG;
wire[7:0] Tile_X4Y8_S2BEG;
wire[7:0] Tile_X4Y8_S2BEGb;
wire[15:0] Tile_X4Y8_S4BEG;
wire[15:0] Tile_X4Y8_SS4BEG;
wire[3:0] Tile_X4Y8_W1BEG;
wire[7:0] Tile_X4Y8_W2BEG;
wire[7:0] Tile_X4Y8_W2BEGb;
wire[15:0] Tile_X4Y8_WW4BEG;
wire[11:0] Tile_X4Y8_W6BEG;
wire[3:0] Tile_X5Y8_N1BEG;
wire[7:0] Tile_X5Y8_N2BEG;
wire[7:0] Tile_X5Y8_N2BEGb;
wire[15:0] Tile_X5Y8_N4BEG;
wire[15:0] Tile_X5Y8_NN4BEG;
wire[3:0] Tile_X5Y8_E1BEG;
wire[7:0] Tile_X5Y8_E2BEG;
wire[7:0] Tile_X5Y8_E2BEGb;
wire[15:0] Tile_X5Y8_EE4BEG;
wire[11:0] Tile_X5Y8_E6BEG;
wire[3:0] Tile_X5Y8_S1BEG;
wire[7:0] Tile_X5Y8_S2BEG;
wire[7:0] Tile_X5Y8_S2BEGb;
wire[15:0] Tile_X5Y8_S4BEG;
wire[15:0] Tile_X5Y8_SS4BEG;
wire[3:0] Tile_X5Y8_W1BEG;
wire[7:0] Tile_X5Y8_W2BEG;
wire[7:0] Tile_X5Y8_W2BEGb;
wire[15:0] Tile_X5Y8_WW4BEG;
wire[11:0] Tile_X5Y8_W6BEG;
wire[0:0] Tile_X5Y8_Co;
wire[3:0] Tile_X6Y8_N1BEG;
wire[7:0] Tile_X6Y8_N2BEG;
wire[7:0] Tile_X6Y8_N2BEGb;
wire[15:0] Tile_X6Y8_N4BEG;
wire[15:0] Tile_X6Y8_NN4BEG;
wire[3:0] Tile_X6Y8_E1BEG;
wire[7:0] Tile_X6Y8_E2BEG;
wire[7:0] Tile_X6Y8_E2BEGb;
wire[15:0] Tile_X6Y8_EE4BEG;
wire[11:0] Tile_X6Y8_E6BEG;
wire[3:0] Tile_X6Y8_S1BEG;
wire[7:0] Tile_X6Y8_S2BEG;
wire[7:0] Tile_X6Y8_S2BEGb;
wire[15:0] Tile_X6Y8_S4BEG;
wire[15:0] Tile_X6Y8_SS4BEG;
wire[3:0] Tile_X6Y8_W1BEG;
wire[7:0] Tile_X6Y8_W2BEG;
wire[7:0] Tile_X6Y8_W2BEGb;
wire[15:0] Tile_X6Y8_WW4BEG;
wire[11:0] Tile_X6Y8_W6BEG;
wire[0:0] Tile_X6Y8_Co;
wire[3:0] Tile_X7Y8_N1BEG;
wire[7:0] Tile_X7Y8_N2BEG;
wire[7:0] Tile_X7Y8_N2BEGb;
wire[15:0] Tile_X7Y8_N4BEG;
wire[15:0] Tile_X7Y8_NN4BEG;
wire[3:0] Tile_X7Y8_E1BEG;
wire[7:0] Tile_X7Y8_E2BEG;
wire[7:0] Tile_X7Y8_E2BEGb;
wire[15:0] Tile_X7Y8_EE4BEG;
wire[11:0] Tile_X7Y8_E6BEG;
wire[3:0] Tile_X7Y8_S1BEG;
wire[7:0] Tile_X7Y8_S2BEG;
wire[7:0] Tile_X7Y8_S2BEGb;
wire[15:0] Tile_X7Y8_S4BEG;
wire[15:0] Tile_X7Y8_SS4BEG;
wire[3:0] Tile_X7Y8_W1BEG;
wire[7:0] Tile_X7Y8_W2BEG;
wire[7:0] Tile_X7Y8_W2BEGb;
wire[15:0] Tile_X7Y8_WW4BEG;
wire[11:0] Tile_X7Y8_W6BEG;
wire[9:0] Tile_X7Y8_bot2top;
wire[3:0] Tile_X8Y8_N1BEG;
wire[7:0] Tile_X8Y8_N2BEG;
wire[7:0] Tile_X8Y8_N2BEGb;
wire[15:0] Tile_X8Y8_N4BEG;
wire[15:0] Tile_X8Y8_NN4BEG;
wire[3:0] Tile_X8Y8_E1BEG;
wire[7:0] Tile_X8Y8_E2BEG;
wire[7:0] Tile_X8Y8_E2BEGb;
wire[15:0] Tile_X8Y8_EE4BEG;
wire[11:0] Tile_X8Y8_E6BEG;
wire[3:0] Tile_X8Y8_S1BEG;
wire[7:0] Tile_X8Y8_S2BEG;
wire[7:0] Tile_X8Y8_S2BEGb;
wire[15:0] Tile_X8Y8_S4BEG;
wire[15:0] Tile_X8Y8_SS4BEG;
wire[3:0] Tile_X8Y8_W1BEG;
wire[7:0] Tile_X8Y8_W2BEG;
wire[7:0] Tile_X8Y8_W2BEGb;
wire[15:0] Tile_X8Y8_WW4BEG;
wire[11:0] Tile_X8Y8_W6BEG;
wire[0:0] Tile_X8Y8_Co;
wire[3:0] Tile_X9Y8_N1BEG;
wire[7:0] Tile_X9Y8_N2BEG;
wire[7:0] Tile_X9Y8_N2BEGb;
wire[15:0] Tile_X9Y8_N4BEG;
wire[15:0] Tile_X9Y8_NN4BEG;
wire[3:0] Tile_X9Y8_E1BEG;
wire[7:0] Tile_X9Y8_E2BEG;
wire[7:0] Tile_X9Y8_E2BEGb;
wire[15:0] Tile_X9Y8_EE4BEG;
wire[11:0] Tile_X9Y8_E6BEG;
wire[3:0] Tile_X9Y8_S1BEG;
wire[7:0] Tile_X9Y8_S2BEG;
wire[7:0] Tile_X9Y8_S2BEGb;
wire[15:0] Tile_X9Y8_S4BEG;
wire[15:0] Tile_X9Y8_SS4BEG;
wire[3:0] Tile_X9Y8_W1BEG;
wire[7:0] Tile_X9Y8_W2BEG;
wire[7:0] Tile_X9Y8_W2BEGb;
wire[15:0] Tile_X9Y8_WW4BEG;
wire[11:0] Tile_X9Y8_W6BEG;
wire[0:0] Tile_X9Y8_Co;
wire[3:0] Tile_X10Y8_N1BEG;
wire[7:0] Tile_X10Y8_N2BEG;
wire[7:0] Tile_X10Y8_N2BEGb;
wire[15:0] Tile_X10Y8_N4BEG;
wire[3:0] Tile_X10Y8_S1BEG;
wire[7:0] Tile_X10Y8_S2BEG;
wire[7:0] Tile_X10Y8_S2BEGb;
wire[15:0] Tile_X10Y8_S4BEG;
wire[3:0] Tile_X10Y8_W1BEG;
wire[7:0] Tile_X10Y8_W2BEG;
wire[7:0] Tile_X10Y8_W2BEGb;
wire[15:0] Tile_X10Y8_WW4BEG;
wire[11:0] Tile_X10Y8_W6BEG;
wire[15:0] Tile_X10Y8_bot2top_DOUT;
wire[3:0] Tile_X0Y9_E1BEG;
wire[7:0] Tile_X0Y9_E2BEG;
wire[7:0] Tile_X0Y9_E2BEGb;
wire[15:0] Tile_X0Y9_EE4BEG;
wire[11:0] Tile_X0Y9_E6BEG;
wire[3:0] Tile_X1Y9_N1BEG;
wire[7:0] Tile_X1Y9_N2BEG;
wire[7:0] Tile_X1Y9_N2BEGb;
wire[15:0] Tile_X1Y9_N4BEG;
wire[15:0] Tile_X1Y9_NN4BEG;
wire[3:0] Tile_X1Y9_E1BEG;
wire[7:0] Tile_X1Y9_E2BEG;
wire[7:0] Tile_X1Y9_E2BEGb;
wire[15:0] Tile_X1Y9_EE4BEG;
wire[11:0] Tile_X1Y9_E6BEG;
wire[3:0] Tile_X1Y9_S1BEG;
wire[7:0] Tile_X1Y9_S2BEG;
wire[7:0] Tile_X1Y9_S2BEGb;
wire[15:0] Tile_X1Y9_S4BEG;
wire[15:0] Tile_X1Y9_SS4BEG;
wire[3:0] Tile_X1Y9_W1BEG;
wire[7:0] Tile_X1Y9_W2BEG;
wire[7:0] Tile_X1Y9_W2BEGb;
wire[15:0] Tile_X1Y9_WW4BEG;
wire[11:0] Tile_X1Y9_W6BEG;
wire[0:0] Tile_X1Y9_Co;
wire[3:0] Tile_X2Y9_N1BEG;
wire[7:0] Tile_X2Y9_N2BEG;
wire[7:0] Tile_X2Y9_N2BEGb;
wire[15:0] Tile_X2Y9_N4BEG;
wire[15:0] Tile_X2Y9_NN4BEG;
wire[3:0] Tile_X2Y9_E1BEG;
wire[7:0] Tile_X2Y9_E2BEG;
wire[7:0] Tile_X2Y9_E2BEGb;
wire[15:0] Tile_X2Y9_EE4BEG;
wire[11:0] Tile_X2Y9_E6BEG;
wire[3:0] Tile_X2Y9_S1BEG;
wire[7:0] Tile_X2Y9_S2BEG;
wire[7:0] Tile_X2Y9_S2BEGb;
wire[15:0] Tile_X2Y9_S4BEG;
wire[15:0] Tile_X2Y9_SS4BEG;
wire[3:0] Tile_X2Y9_W1BEG;
wire[7:0] Tile_X2Y9_W2BEG;
wire[7:0] Tile_X2Y9_W2BEGb;
wire[15:0] Tile_X2Y9_WW4BEG;
wire[11:0] Tile_X2Y9_W6BEG;
wire[0:0] Tile_X2Y9_Co;
wire[3:0] Tile_X3Y9_N1BEG;
wire[7:0] Tile_X3Y9_N2BEG;
wire[7:0] Tile_X3Y9_N2BEGb;
wire[15:0] Tile_X3Y9_N4BEG;
wire[15:0] Tile_X3Y9_NN4BEG;
wire[3:0] Tile_X3Y9_E1BEG;
wire[7:0] Tile_X3Y9_E2BEG;
wire[7:0] Tile_X3Y9_E2BEGb;
wire[15:0] Tile_X3Y9_EE4BEG;
wire[11:0] Tile_X3Y9_E6BEG;
wire[3:0] Tile_X3Y9_S1BEG;
wire[7:0] Tile_X3Y9_S2BEG;
wire[7:0] Tile_X3Y9_S2BEGb;
wire[15:0] Tile_X3Y9_S4BEG;
wire[15:0] Tile_X3Y9_SS4BEG;
wire[3:0] Tile_X3Y9_W1BEG;
wire[7:0] Tile_X3Y9_W2BEG;
wire[7:0] Tile_X3Y9_W2BEGb;
wire[15:0] Tile_X3Y9_WW4BEG;
wire[11:0] Tile_X3Y9_W6BEG;
wire[0:0] Tile_X3Y9_Co;
wire[3:0] Tile_X4Y9_N1BEG;
wire[7:0] Tile_X4Y9_N2BEG;
wire[7:0] Tile_X4Y9_N2BEGb;
wire[15:0] Tile_X4Y9_N4BEG;
wire[15:0] Tile_X4Y9_NN4BEG;
wire[3:0] Tile_X4Y9_E1BEG;
wire[7:0] Tile_X4Y9_E2BEG;
wire[7:0] Tile_X4Y9_E2BEGb;
wire[15:0] Tile_X4Y9_EE4BEG;
wire[11:0] Tile_X4Y9_E6BEG;
wire[3:0] Tile_X4Y9_S1BEG;
wire[7:0] Tile_X4Y9_S2BEG;
wire[7:0] Tile_X4Y9_S2BEGb;
wire[15:0] Tile_X4Y9_S4BEG;
wire[15:0] Tile_X4Y9_SS4BEG;
wire[3:0] Tile_X4Y9_W1BEG;
wire[7:0] Tile_X4Y9_W2BEG;
wire[7:0] Tile_X4Y9_W2BEGb;
wire[15:0] Tile_X4Y9_WW4BEG;
wire[11:0] Tile_X4Y9_W6BEG;
wire[3:0] Tile_X5Y9_N1BEG;
wire[7:0] Tile_X5Y9_N2BEG;
wire[7:0] Tile_X5Y9_N2BEGb;
wire[15:0] Tile_X5Y9_N4BEG;
wire[15:0] Tile_X5Y9_NN4BEG;
wire[3:0] Tile_X5Y9_E1BEG;
wire[7:0] Tile_X5Y9_E2BEG;
wire[7:0] Tile_X5Y9_E2BEGb;
wire[15:0] Tile_X5Y9_EE4BEG;
wire[11:0] Tile_X5Y9_E6BEG;
wire[3:0] Tile_X5Y9_S1BEG;
wire[7:0] Tile_X5Y9_S2BEG;
wire[7:0] Tile_X5Y9_S2BEGb;
wire[15:0] Tile_X5Y9_S4BEG;
wire[15:0] Tile_X5Y9_SS4BEG;
wire[3:0] Tile_X5Y9_W1BEG;
wire[7:0] Tile_X5Y9_W2BEG;
wire[7:0] Tile_X5Y9_W2BEGb;
wire[15:0] Tile_X5Y9_WW4BEG;
wire[11:0] Tile_X5Y9_W6BEG;
wire[0:0] Tile_X5Y9_Co;
wire[3:0] Tile_X6Y9_N1BEG;
wire[7:0] Tile_X6Y9_N2BEG;
wire[7:0] Tile_X6Y9_N2BEGb;
wire[15:0] Tile_X6Y9_N4BEG;
wire[15:0] Tile_X6Y9_NN4BEG;
wire[3:0] Tile_X6Y9_E1BEG;
wire[7:0] Tile_X6Y9_E2BEG;
wire[7:0] Tile_X6Y9_E2BEGb;
wire[15:0] Tile_X6Y9_EE4BEG;
wire[11:0] Tile_X6Y9_E6BEG;
wire[3:0] Tile_X6Y9_S1BEG;
wire[7:0] Tile_X6Y9_S2BEG;
wire[7:0] Tile_X6Y9_S2BEGb;
wire[15:0] Tile_X6Y9_S4BEG;
wire[15:0] Tile_X6Y9_SS4BEG;
wire[3:0] Tile_X6Y9_W1BEG;
wire[7:0] Tile_X6Y9_W2BEG;
wire[7:0] Tile_X6Y9_W2BEGb;
wire[15:0] Tile_X6Y9_WW4BEG;
wire[11:0] Tile_X6Y9_W6BEG;
wire[0:0] Tile_X6Y9_Co;
wire[3:0] Tile_X7Y9_N1BEG;
wire[7:0] Tile_X7Y9_N2BEG;
wire[7:0] Tile_X7Y9_N2BEGb;
wire[15:0] Tile_X7Y9_N4BEG;
wire[15:0] Tile_X7Y9_NN4BEG;
wire[3:0] Tile_X7Y9_E1BEG;
wire[7:0] Tile_X7Y9_E2BEG;
wire[7:0] Tile_X7Y9_E2BEGb;
wire[15:0] Tile_X7Y9_EE4BEG;
wire[11:0] Tile_X7Y9_E6BEG;
wire[3:0] Tile_X7Y9_S1BEG;
wire[7:0] Tile_X7Y9_S2BEG;
wire[7:0] Tile_X7Y9_S2BEGb;
wire[15:0] Tile_X7Y9_S4BEG;
wire[15:0] Tile_X7Y9_SS4BEG;
wire[3:0] Tile_X7Y9_W1BEG;
wire[7:0] Tile_X7Y9_W2BEG;
wire[7:0] Tile_X7Y9_W2BEGb;
wire[15:0] Tile_X7Y9_WW4BEG;
wire[11:0] Tile_X7Y9_W6BEG;
wire[17:0] Tile_X7Y9_top2bot;
wire[3:0] Tile_X8Y9_N1BEG;
wire[7:0] Tile_X8Y9_N2BEG;
wire[7:0] Tile_X8Y9_N2BEGb;
wire[15:0] Tile_X8Y9_N4BEG;
wire[15:0] Tile_X8Y9_NN4BEG;
wire[3:0] Tile_X8Y9_E1BEG;
wire[7:0] Tile_X8Y9_E2BEG;
wire[7:0] Tile_X8Y9_E2BEGb;
wire[15:0] Tile_X8Y9_EE4BEG;
wire[11:0] Tile_X8Y9_E6BEG;
wire[3:0] Tile_X8Y9_S1BEG;
wire[7:0] Tile_X8Y9_S2BEG;
wire[7:0] Tile_X8Y9_S2BEGb;
wire[15:0] Tile_X8Y9_S4BEG;
wire[15:0] Tile_X8Y9_SS4BEG;
wire[3:0] Tile_X8Y9_W1BEG;
wire[7:0] Tile_X8Y9_W2BEG;
wire[7:0] Tile_X8Y9_W2BEGb;
wire[15:0] Tile_X8Y9_WW4BEG;
wire[11:0] Tile_X8Y9_W6BEG;
wire[0:0] Tile_X8Y9_Co;
wire[3:0] Tile_X9Y9_N1BEG;
wire[7:0] Tile_X9Y9_N2BEG;
wire[7:0] Tile_X9Y9_N2BEGb;
wire[15:0] Tile_X9Y9_N4BEG;
wire[15:0] Tile_X9Y9_NN4BEG;
wire[3:0] Tile_X9Y9_E1BEG;
wire[7:0] Tile_X9Y9_E2BEG;
wire[7:0] Tile_X9Y9_E2BEGb;
wire[15:0] Tile_X9Y9_EE4BEG;
wire[11:0] Tile_X9Y9_E6BEG;
wire[3:0] Tile_X9Y9_S1BEG;
wire[7:0] Tile_X9Y9_S2BEG;
wire[7:0] Tile_X9Y9_S2BEGb;
wire[15:0] Tile_X9Y9_S4BEG;
wire[15:0] Tile_X9Y9_SS4BEG;
wire[3:0] Tile_X9Y9_W1BEG;
wire[7:0] Tile_X9Y9_W2BEG;
wire[7:0] Tile_X9Y9_W2BEGb;
wire[15:0] Tile_X9Y9_WW4BEG;
wire[11:0] Tile_X9Y9_W6BEG;
wire[0:0] Tile_X9Y9_Co;
wire[3:0] Tile_X10Y9_N1BEG;
wire[7:0] Tile_X10Y9_N2BEG;
wire[7:0] Tile_X10Y9_N2BEGb;
wire[15:0] Tile_X10Y9_N4BEG;
wire[3:0] Tile_X10Y9_S1BEG;
wire[7:0] Tile_X10Y9_S2BEG;
wire[7:0] Tile_X10Y9_S2BEGb;
wire[15:0] Tile_X10Y9_S4BEG;
wire[3:0] Tile_X10Y9_W1BEG;
wire[7:0] Tile_X10Y9_W2BEG;
wire[7:0] Tile_X10Y9_W2BEGb;
wire[15:0] Tile_X10Y9_WW4BEG;
wire[11:0] Tile_X10Y9_W6BEG;
wire[15:0] Tile_X10Y9_top2bot_DIN;
wire[15:0] Tile_X10Y9_top2bot_BM;
wire[4:0] Tile_X10Y9_top2bot_ADDR;
wire[3:0] Tile_X0Y10_E1BEG;
wire[7:0] Tile_X0Y10_E2BEG;
wire[7:0] Tile_X0Y10_E2BEGb;
wire[15:0] Tile_X0Y10_EE4BEG;
wire[11:0] Tile_X0Y10_E6BEG;
wire[3:0] Tile_X1Y10_N1BEG;
wire[7:0] Tile_X1Y10_N2BEG;
wire[7:0] Tile_X1Y10_N2BEGb;
wire[15:0] Tile_X1Y10_N4BEG;
wire[15:0] Tile_X1Y10_NN4BEG;
wire[3:0] Tile_X1Y10_E1BEG;
wire[7:0] Tile_X1Y10_E2BEG;
wire[7:0] Tile_X1Y10_E2BEGb;
wire[15:0] Tile_X1Y10_EE4BEG;
wire[11:0] Tile_X1Y10_E6BEG;
wire[3:0] Tile_X1Y10_S1BEG;
wire[7:0] Tile_X1Y10_S2BEG;
wire[7:0] Tile_X1Y10_S2BEGb;
wire[15:0] Tile_X1Y10_S4BEG;
wire[15:0] Tile_X1Y10_SS4BEG;
wire[3:0] Tile_X1Y10_W1BEG;
wire[7:0] Tile_X1Y10_W2BEG;
wire[7:0] Tile_X1Y10_W2BEGb;
wire[15:0] Tile_X1Y10_WW4BEG;
wire[11:0] Tile_X1Y10_W6BEG;
wire[0:0] Tile_X1Y10_Co;
wire[3:0] Tile_X2Y10_N1BEG;
wire[7:0] Tile_X2Y10_N2BEG;
wire[7:0] Tile_X2Y10_N2BEGb;
wire[15:0] Tile_X2Y10_N4BEG;
wire[15:0] Tile_X2Y10_NN4BEG;
wire[3:0] Tile_X2Y10_E1BEG;
wire[7:0] Tile_X2Y10_E2BEG;
wire[7:0] Tile_X2Y10_E2BEGb;
wire[15:0] Tile_X2Y10_EE4BEG;
wire[11:0] Tile_X2Y10_E6BEG;
wire[3:0] Tile_X2Y10_S1BEG;
wire[7:0] Tile_X2Y10_S2BEG;
wire[7:0] Tile_X2Y10_S2BEGb;
wire[15:0] Tile_X2Y10_S4BEG;
wire[15:0] Tile_X2Y10_SS4BEG;
wire[3:0] Tile_X2Y10_W1BEG;
wire[7:0] Tile_X2Y10_W2BEG;
wire[7:0] Tile_X2Y10_W2BEGb;
wire[15:0] Tile_X2Y10_WW4BEG;
wire[11:0] Tile_X2Y10_W6BEG;
wire[0:0] Tile_X2Y10_Co;
wire[3:0] Tile_X3Y10_N1BEG;
wire[7:0] Tile_X3Y10_N2BEG;
wire[7:0] Tile_X3Y10_N2BEGb;
wire[15:0] Tile_X3Y10_N4BEG;
wire[15:0] Tile_X3Y10_NN4BEG;
wire[3:0] Tile_X3Y10_E1BEG;
wire[7:0] Tile_X3Y10_E2BEG;
wire[7:0] Tile_X3Y10_E2BEGb;
wire[15:0] Tile_X3Y10_EE4BEG;
wire[11:0] Tile_X3Y10_E6BEG;
wire[3:0] Tile_X3Y10_S1BEG;
wire[7:0] Tile_X3Y10_S2BEG;
wire[7:0] Tile_X3Y10_S2BEGb;
wire[15:0] Tile_X3Y10_S4BEG;
wire[15:0] Tile_X3Y10_SS4BEG;
wire[3:0] Tile_X3Y10_W1BEG;
wire[7:0] Tile_X3Y10_W2BEG;
wire[7:0] Tile_X3Y10_W2BEGb;
wire[15:0] Tile_X3Y10_WW4BEG;
wire[11:0] Tile_X3Y10_W6BEG;
wire[0:0] Tile_X3Y10_Co;
wire[3:0] Tile_X4Y10_N1BEG;
wire[7:0] Tile_X4Y10_N2BEG;
wire[7:0] Tile_X4Y10_N2BEGb;
wire[15:0] Tile_X4Y10_N4BEG;
wire[15:0] Tile_X4Y10_NN4BEG;
wire[3:0] Tile_X4Y10_E1BEG;
wire[7:0] Tile_X4Y10_E2BEG;
wire[7:0] Tile_X4Y10_E2BEGb;
wire[15:0] Tile_X4Y10_EE4BEG;
wire[11:0] Tile_X4Y10_E6BEG;
wire[3:0] Tile_X4Y10_S1BEG;
wire[7:0] Tile_X4Y10_S2BEG;
wire[7:0] Tile_X4Y10_S2BEGb;
wire[15:0] Tile_X4Y10_S4BEG;
wire[15:0] Tile_X4Y10_SS4BEG;
wire[3:0] Tile_X4Y10_W1BEG;
wire[7:0] Tile_X4Y10_W2BEG;
wire[7:0] Tile_X4Y10_W2BEGb;
wire[15:0] Tile_X4Y10_WW4BEG;
wire[11:0] Tile_X4Y10_W6BEG;
wire[3:0] Tile_X5Y10_N1BEG;
wire[7:0] Tile_X5Y10_N2BEG;
wire[7:0] Tile_X5Y10_N2BEGb;
wire[15:0] Tile_X5Y10_N4BEG;
wire[15:0] Tile_X5Y10_NN4BEG;
wire[3:0] Tile_X5Y10_E1BEG;
wire[7:0] Tile_X5Y10_E2BEG;
wire[7:0] Tile_X5Y10_E2BEGb;
wire[15:0] Tile_X5Y10_EE4BEG;
wire[11:0] Tile_X5Y10_E6BEG;
wire[3:0] Tile_X5Y10_S1BEG;
wire[7:0] Tile_X5Y10_S2BEG;
wire[7:0] Tile_X5Y10_S2BEGb;
wire[15:0] Tile_X5Y10_S4BEG;
wire[15:0] Tile_X5Y10_SS4BEG;
wire[3:0] Tile_X5Y10_W1BEG;
wire[7:0] Tile_X5Y10_W2BEG;
wire[7:0] Tile_X5Y10_W2BEGb;
wire[15:0] Tile_X5Y10_WW4BEG;
wire[11:0] Tile_X5Y10_W6BEG;
wire[0:0] Tile_X5Y10_Co;
wire[3:0] Tile_X6Y10_N1BEG;
wire[7:0] Tile_X6Y10_N2BEG;
wire[7:0] Tile_X6Y10_N2BEGb;
wire[15:0] Tile_X6Y10_N4BEG;
wire[15:0] Tile_X6Y10_NN4BEG;
wire[3:0] Tile_X6Y10_E1BEG;
wire[7:0] Tile_X6Y10_E2BEG;
wire[7:0] Tile_X6Y10_E2BEGb;
wire[15:0] Tile_X6Y10_EE4BEG;
wire[11:0] Tile_X6Y10_E6BEG;
wire[3:0] Tile_X6Y10_S1BEG;
wire[7:0] Tile_X6Y10_S2BEG;
wire[7:0] Tile_X6Y10_S2BEGb;
wire[15:0] Tile_X6Y10_S4BEG;
wire[15:0] Tile_X6Y10_SS4BEG;
wire[3:0] Tile_X6Y10_W1BEG;
wire[7:0] Tile_X6Y10_W2BEG;
wire[7:0] Tile_X6Y10_W2BEGb;
wire[15:0] Tile_X6Y10_WW4BEG;
wire[11:0] Tile_X6Y10_W6BEG;
wire[0:0] Tile_X6Y10_Co;
wire[3:0] Tile_X7Y10_N1BEG;
wire[7:0] Tile_X7Y10_N2BEG;
wire[7:0] Tile_X7Y10_N2BEGb;
wire[15:0] Tile_X7Y10_N4BEG;
wire[15:0] Tile_X7Y10_NN4BEG;
wire[3:0] Tile_X7Y10_E1BEG;
wire[7:0] Tile_X7Y10_E2BEG;
wire[7:0] Tile_X7Y10_E2BEGb;
wire[15:0] Tile_X7Y10_EE4BEG;
wire[11:0] Tile_X7Y10_E6BEG;
wire[3:0] Tile_X7Y10_S1BEG;
wire[7:0] Tile_X7Y10_S2BEG;
wire[7:0] Tile_X7Y10_S2BEGb;
wire[15:0] Tile_X7Y10_S4BEG;
wire[15:0] Tile_X7Y10_SS4BEG;
wire[3:0] Tile_X7Y10_W1BEG;
wire[7:0] Tile_X7Y10_W2BEG;
wire[7:0] Tile_X7Y10_W2BEGb;
wire[15:0] Tile_X7Y10_WW4BEG;
wire[11:0] Tile_X7Y10_W6BEG;
wire[9:0] Tile_X7Y10_bot2top;
wire[3:0] Tile_X8Y10_N1BEG;
wire[7:0] Tile_X8Y10_N2BEG;
wire[7:0] Tile_X8Y10_N2BEGb;
wire[15:0] Tile_X8Y10_N4BEG;
wire[15:0] Tile_X8Y10_NN4BEG;
wire[3:0] Tile_X8Y10_E1BEG;
wire[7:0] Tile_X8Y10_E2BEG;
wire[7:0] Tile_X8Y10_E2BEGb;
wire[15:0] Tile_X8Y10_EE4BEG;
wire[11:0] Tile_X8Y10_E6BEG;
wire[3:0] Tile_X8Y10_S1BEG;
wire[7:0] Tile_X8Y10_S2BEG;
wire[7:0] Tile_X8Y10_S2BEGb;
wire[15:0] Tile_X8Y10_S4BEG;
wire[15:0] Tile_X8Y10_SS4BEG;
wire[3:0] Tile_X8Y10_W1BEG;
wire[7:0] Tile_X8Y10_W2BEG;
wire[7:0] Tile_X8Y10_W2BEGb;
wire[15:0] Tile_X8Y10_WW4BEG;
wire[11:0] Tile_X8Y10_W6BEG;
wire[0:0] Tile_X8Y10_Co;
wire[3:0] Tile_X9Y10_N1BEG;
wire[7:0] Tile_X9Y10_N2BEG;
wire[7:0] Tile_X9Y10_N2BEGb;
wire[15:0] Tile_X9Y10_N4BEG;
wire[15:0] Tile_X9Y10_NN4BEG;
wire[3:0] Tile_X9Y10_E1BEG;
wire[7:0] Tile_X9Y10_E2BEG;
wire[7:0] Tile_X9Y10_E2BEGb;
wire[15:0] Tile_X9Y10_EE4BEG;
wire[11:0] Tile_X9Y10_E6BEG;
wire[3:0] Tile_X9Y10_S1BEG;
wire[7:0] Tile_X9Y10_S2BEG;
wire[7:0] Tile_X9Y10_S2BEGb;
wire[15:0] Tile_X9Y10_S4BEG;
wire[15:0] Tile_X9Y10_SS4BEG;
wire[3:0] Tile_X9Y10_W1BEG;
wire[7:0] Tile_X9Y10_W2BEG;
wire[7:0] Tile_X9Y10_W2BEGb;
wire[15:0] Tile_X9Y10_WW4BEG;
wire[11:0] Tile_X9Y10_W6BEG;
wire[0:0] Tile_X9Y10_Co;
wire[3:0] Tile_X10Y10_N1BEG;
wire[7:0] Tile_X10Y10_N2BEG;
wire[7:0] Tile_X10Y10_N2BEGb;
wire[15:0] Tile_X10Y10_N4BEG;
wire[3:0] Tile_X10Y10_S1BEG;
wire[7:0] Tile_X10Y10_S2BEG;
wire[7:0] Tile_X10Y10_S2BEGb;
wire[15:0] Tile_X10Y10_S4BEG;
wire[3:0] Tile_X10Y10_W1BEG;
wire[7:0] Tile_X10Y10_W2BEG;
wire[7:0] Tile_X10Y10_W2BEGb;
wire[15:0] Tile_X10Y10_WW4BEG;
wire[11:0] Tile_X10Y10_W6BEG;
wire[15:0] Tile_X10Y10_bot2top_DOUT;
wire[3:0] Tile_X0Y11_E1BEG;
wire[7:0] Tile_X0Y11_E2BEG;
wire[7:0] Tile_X0Y11_E2BEGb;
wire[15:0] Tile_X0Y11_EE4BEG;
wire[11:0] Tile_X0Y11_E6BEG;
wire[3:0] Tile_X1Y11_N1BEG;
wire[7:0] Tile_X1Y11_N2BEG;
wire[7:0] Tile_X1Y11_N2BEGb;
wire[15:0] Tile_X1Y11_N4BEG;
wire[15:0] Tile_X1Y11_NN4BEG;
wire[3:0] Tile_X1Y11_E1BEG;
wire[7:0] Tile_X1Y11_E2BEG;
wire[7:0] Tile_X1Y11_E2BEGb;
wire[15:0] Tile_X1Y11_EE4BEG;
wire[11:0] Tile_X1Y11_E6BEG;
wire[3:0] Tile_X1Y11_S1BEG;
wire[7:0] Tile_X1Y11_S2BEG;
wire[7:0] Tile_X1Y11_S2BEGb;
wire[15:0] Tile_X1Y11_S4BEG;
wire[15:0] Tile_X1Y11_SS4BEG;
wire[3:0] Tile_X1Y11_W1BEG;
wire[7:0] Tile_X1Y11_W2BEG;
wire[7:0] Tile_X1Y11_W2BEGb;
wire[15:0] Tile_X1Y11_WW4BEG;
wire[11:0] Tile_X1Y11_W6BEG;
wire[0:0] Tile_X1Y11_Co;
wire[3:0] Tile_X2Y11_N1BEG;
wire[7:0] Tile_X2Y11_N2BEG;
wire[7:0] Tile_X2Y11_N2BEGb;
wire[15:0] Tile_X2Y11_N4BEG;
wire[15:0] Tile_X2Y11_NN4BEG;
wire[3:0] Tile_X2Y11_E1BEG;
wire[7:0] Tile_X2Y11_E2BEG;
wire[7:0] Tile_X2Y11_E2BEGb;
wire[15:0] Tile_X2Y11_EE4BEG;
wire[11:0] Tile_X2Y11_E6BEG;
wire[3:0] Tile_X2Y11_S1BEG;
wire[7:0] Tile_X2Y11_S2BEG;
wire[7:0] Tile_X2Y11_S2BEGb;
wire[15:0] Tile_X2Y11_S4BEG;
wire[15:0] Tile_X2Y11_SS4BEG;
wire[3:0] Tile_X2Y11_W1BEG;
wire[7:0] Tile_X2Y11_W2BEG;
wire[7:0] Tile_X2Y11_W2BEGb;
wire[15:0] Tile_X2Y11_WW4BEG;
wire[11:0] Tile_X2Y11_W6BEG;
wire[0:0] Tile_X2Y11_Co;
wire[3:0] Tile_X3Y11_N1BEG;
wire[7:0] Tile_X3Y11_N2BEG;
wire[7:0] Tile_X3Y11_N2BEGb;
wire[15:0] Tile_X3Y11_N4BEG;
wire[15:0] Tile_X3Y11_NN4BEG;
wire[3:0] Tile_X3Y11_E1BEG;
wire[7:0] Tile_X3Y11_E2BEG;
wire[7:0] Tile_X3Y11_E2BEGb;
wire[15:0] Tile_X3Y11_EE4BEG;
wire[11:0] Tile_X3Y11_E6BEG;
wire[3:0] Tile_X3Y11_S1BEG;
wire[7:0] Tile_X3Y11_S2BEG;
wire[7:0] Tile_X3Y11_S2BEGb;
wire[15:0] Tile_X3Y11_S4BEG;
wire[15:0] Tile_X3Y11_SS4BEG;
wire[3:0] Tile_X3Y11_W1BEG;
wire[7:0] Tile_X3Y11_W2BEG;
wire[7:0] Tile_X3Y11_W2BEGb;
wire[15:0] Tile_X3Y11_WW4BEG;
wire[11:0] Tile_X3Y11_W6BEG;
wire[0:0] Tile_X3Y11_Co;
wire[3:0] Tile_X4Y11_N1BEG;
wire[7:0] Tile_X4Y11_N2BEG;
wire[7:0] Tile_X4Y11_N2BEGb;
wire[15:0] Tile_X4Y11_N4BEG;
wire[15:0] Tile_X4Y11_NN4BEG;
wire[3:0] Tile_X4Y11_E1BEG;
wire[7:0] Tile_X4Y11_E2BEG;
wire[7:0] Tile_X4Y11_E2BEGb;
wire[15:0] Tile_X4Y11_EE4BEG;
wire[11:0] Tile_X4Y11_E6BEG;
wire[3:0] Tile_X4Y11_S1BEG;
wire[7:0] Tile_X4Y11_S2BEG;
wire[7:0] Tile_X4Y11_S2BEGb;
wire[15:0] Tile_X4Y11_S4BEG;
wire[15:0] Tile_X4Y11_SS4BEG;
wire[3:0] Tile_X4Y11_W1BEG;
wire[7:0] Tile_X4Y11_W2BEG;
wire[7:0] Tile_X4Y11_W2BEGb;
wire[15:0] Tile_X4Y11_WW4BEG;
wire[11:0] Tile_X4Y11_W6BEG;
wire[3:0] Tile_X5Y11_N1BEG;
wire[7:0] Tile_X5Y11_N2BEG;
wire[7:0] Tile_X5Y11_N2BEGb;
wire[15:0] Tile_X5Y11_N4BEG;
wire[15:0] Tile_X5Y11_NN4BEG;
wire[3:0] Tile_X5Y11_E1BEG;
wire[7:0] Tile_X5Y11_E2BEG;
wire[7:0] Tile_X5Y11_E2BEGb;
wire[15:0] Tile_X5Y11_EE4BEG;
wire[11:0] Tile_X5Y11_E6BEG;
wire[3:0] Tile_X5Y11_S1BEG;
wire[7:0] Tile_X5Y11_S2BEG;
wire[7:0] Tile_X5Y11_S2BEGb;
wire[15:0] Tile_X5Y11_S4BEG;
wire[15:0] Tile_X5Y11_SS4BEG;
wire[3:0] Tile_X5Y11_W1BEG;
wire[7:0] Tile_X5Y11_W2BEG;
wire[7:0] Tile_X5Y11_W2BEGb;
wire[15:0] Tile_X5Y11_WW4BEG;
wire[11:0] Tile_X5Y11_W6BEG;
wire[0:0] Tile_X5Y11_Co;
wire[3:0] Tile_X6Y11_N1BEG;
wire[7:0] Tile_X6Y11_N2BEG;
wire[7:0] Tile_X6Y11_N2BEGb;
wire[15:0] Tile_X6Y11_N4BEG;
wire[15:0] Tile_X6Y11_NN4BEG;
wire[3:0] Tile_X6Y11_E1BEG;
wire[7:0] Tile_X6Y11_E2BEG;
wire[7:0] Tile_X6Y11_E2BEGb;
wire[15:0] Tile_X6Y11_EE4BEG;
wire[11:0] Tile_X6Y11_E6BEG;
wire[3:0] Tile_X6Y11_S1BEG;
wire[7:0] Tile_X6Y11_S2BEG;
wire[7:0] Tile_X6Y11_S2BEGb;
wire[15:0] Tile_X6Y11_S4BEG;
wire[15:0] Tile_X6Y11_SS4BEG;
wire[3:0] Tile_X6Y11_W1BEG;
wire[7:0] Tile_X6Y11_W2BEG;
wire[7:0] Tile_X6Y11_W2BEGb;
wire[15:0] Tile_X6Y11_WW4BEG;
wire[11:0] Tile_X6Y11_W6BEG;
wire[0:0] Tile_X6Y11_Co;
wire[3:0] Tile_X7Y11_N1BEG;
wire[7:0] Tile_X7Y11_N2BEG;
wire[7:0] Tile_X7Y11_N2BEGb;
wire[15:0] Tile_X7Y11_N4BEG;
wire[15:0] Tile_X7Y11_NN4BEG;
wire[3:0] Tile_X7Y11_E1BEG;
wire[7:0] Tile_X7Y11_E2BEG;
wire[7:0] Tile_X7Y11_E2BEGb;
wire[15:0] Tile_X7Y11_EE4BEG;
wire[11:0] Tile_X7Y11_E6BEG;
wire[3:0] Tile_X7Y11_S1BEG;
wire[7:0] Tile_X7Y11_S2BEG;
wire[7:0] Tile_X7Y11_S2BEGb;
wire[15:0] Tile_X7Y11_S4BEG;
wire[15:0] Tile_X7Y11_SS4BEG;
wire[3:0] Tile_X7Y11_W1BEG;
wire[7:0] Tile_X7Y11_W2BEG;
wire[7:0] Tile_X7Y11_W2BEGb;
wire[15:0] Tile_X7Y11_WW4BEG;
wire[11:0] Tile_X7Y11_W6BEG;
wire[17:0] Tile_X7Y11_top2bot;
wire[3:0] Tile_X8Y11_N1BEG;
wire[7:0] Tile_X8Y11_N2BEG;
wire[7:0] Tile_X8Y11_N2BEGb;
wire[15:0] Tile_X8Y11_N4BEG;
wire[15:0] Tile_X8Y11_NN4BEG;
wire[3:0] Tile_X8Y11_E1BEG;
wire[7:0] Tile_X8Y11_E2BEG;
wire[7:0] Tile_X8Y11_E2BEGb;
wire[15:0] Tile_X8Y11_EE4BEG;
wire[11:0] Tile_X8Y11_E6BEG;
wire[3:0] Tile_X8Y11_S1BEG;
wire[7:0] Tile_X8Y11_S2BEG;
wire[7:0] Tile_X8Y11_S2BEGb;
wire[15:0] Tile_X8Y11_S4BEG;
wire[15:0] Tile_X8Y11_SS4BEG;
wire[3:0] Tile_X8Y11_W1BEG;
wire[7:0] Tile_X8Y11_W2BEG;
wire[7:0] Tile_X8Y11_W2BEGb;
wire[15:0] Tile_X8Y11_WW4BEG;
wire[11:0] Tile_X8Y11_W6BEG;
wire[0:0] Tile_X8Y11_Co;
wire[3:0] Tile_X9Y11_N1BEG;
wire[7:0] Tile_X9Y11_N2BEG;
wire[7:0] Tile_X9Y11_N2BEGb;
wire[15:0] Tile_X9Y11_N4BEG;
wire[15:0] Tile_X9Y11_NN4BEG;
wire[3:0] Tile_X9Y11_E1BEG;
wire[7:0] Tile_X9Y11_E2BEG;
wire[7:0] Tile_X9Y11_E2BEGb;
wire[15:0] Tile_X9Y11_EE4BEG;
wire[11:0] Tile_X9Y11_E6BEG;
wire[3:0] Tile_X9Y11_S1BEG;
wire[7:0] Tile_X9Y11_S2BEG;
wire[7:0] Tile_X9Y11_S2BEGb;
wire[15:0] Tile_X9Y11_S4BEG;
wire[15:0] Tile_X9Y11_SS4BEG;
wire[3:0] Tile_X9Y11_W1BEG;
wire[7:0] Tile_X9Y11_W2BEG;
wire[7:0] Tile_X9Y11_W2BEGb;
wire[15:0] Tile_X9Y11_WW4BEG;
wire[11:0] Tile_X9Y11_W6BEG;
wire[0:0] Tile_X9Y11_Co;
wire[3:0] Tile_X10Y11_N1BEG;
wire[7:0] Tile_X10Y11_N2BEG;
wire[7:0] Tile_X10Y11_N2BEGb;
wire[15:0] Tile_X10Y11_N4BEG;
wire[3:0] Tile_X10Y11_S1BEG;
wire[7:0] Tile_X10Y11_S2BEG;
wire[7:0] Tile_X10Y11_S2BEGb;
wire[15:0] Tile_X10Y11_S4BEG;
wire[3:0] Tile_X10Y11_W1BEG;
wire[7:0] Tile_X10Y11_W2BEG;
wire[7:0] Tile_X10Y11_W2BEGb;
wire[15:0] Tile_X10Y11_WW4BEG;
wire[11:0] Tile_X10Y11_W6BEG;
wire[15:0] Tile_X10Y11_top2bot_DIN;
wire[15:0] Tile_X10Y11_top2bot_BM;
wire[4:0] Tile_X10Y11_top2bot_ADDR;
wire[3:0] Tile_X0Y12_E1BEG;
wire[7:0] Tile_X0Y12_E2BEG;
wire[7:0] Tile_X0Y12_E2BEGb;
wire[15:0] Tile_X0Y12_EE4BEG;
wire[11:0] Tile_X0Y12_E6BEG;
wire[3:0] Tile_X1Y12_N1BEG;
wire[7:0] Tile_X1Y12_N2BEG;
wire[7:0] Tile_X1Y12_N2BEGb;
wire[15:0] Tile_X1Y12_N4BEG;
wire[15:0] Tile_X1Y12_NN4BEG;
wire[3:0] Tile_X1Y12_E1BEG;
wire[7:0] Tile_X1Y12_E2BEG;
wire[7:0] Tile_X1Y12_E2BEGb;
wire[15:0] Tile_X1Y12_EE4BEG;
wire[11:0] Tile_X1Y12_E6BEG;
wire[3:0] Tile_X1Y12_S1BEG;
wire[7:0] Tile_X1Y12_S2BEG;
wire[7:0] Tile_X1Y12_S2BEGb;
wire[15:0] Tile_X1Y12_S4BEG;
wire[15:0] Tile_X1Y12_SS4BEG;
wire[3:0] Tile_X1Y12_W1BEG;
wire[7:0] Tile_X1Y12_W2BEG;
wire[7:0] Tile_X1Y12_W2BEGb;
wire[15:0] Tile_X1Y12_WW4BEG;
wire[11:0] Tile_X1Y12_W6BEG;
wire[0:0] Tile_X1Y12_Co;
wire[3:0] Tile_X2Y12_N1BEG;
wire[7:0] Tile_X2Y12_N2BEG;
wire[7:0] Tile_X2Y12_N2BEGb;
wire[15:0] Tile_X2Y12_N4BEG;
wire[15:0] Tile_X2Y12_NN4BEG;
wire[3:0] Tile_X2Y12_E1BEG;
wire[7:0] Tile_X2Y12_E2BEG;
wire[7:0] Tile_X2Y12_E2BEGb;
wire[15:0] Tile_X2Y12_EE4BEG;
wire[11:0] Tile_X2Y12_E6BEG;
wire[3:0] Tile_X2Y12_S1BEG;
wire[7:0] Tile_X2Y12_S2BEG;
wire[7:0] Tile_X2Y12_S2BEGb;
wire[15:0] Tile_X2Y12_S4BEG;
wire[15:0] Tile_X2Y12_SS4BEG;
wire[3:0] Tile_X2Y12_W1BEG;
wire[7:0] Tile_X2Y12_W2BEG;
wire[7:0] Tile_X2Y12_W2BEGb;
wire[15:0] Tile_X2Y12_WW4BEG;
wire[11:0] Tile_X2Y12_W6BEG;
wire[0:0] Tile_X2Y12_Co;
wire[3:0] Tile_X3Y12_N1BEG;
wire[7:0] Tile_X3Y12_N2BEG;
wire[7:0] Tile_X3Y12_N2BEGb;
wire[15:0] Tile_X3Y12_N4BEG;
wire[15:0] Tile_X3Y12_NN4BEG;
wire[3:0] Tile_X3Y12_E1BEG;
wire[7:0] Tile_X3Y12_E2BEG;
wire[7:0] Tile_X3Y12_E2BEGb;
wire[15:0] Tile_X3Y12_EE4BEG;
wire[11:0] Tile_X3Y12_E6BEG;
wire[3:0] Tile_X3Y12_S1BEG;
wire[7:0] Tile_X3Y12_S2BEG;
wire[7:0] Tile_X3Y12_S2BEGb;
wire[15:0] Tile_X3Y12_S4BEG;
wire[15:0] Tile_X3Y12_SS4BEG;
wire[3:0] Tile_X3Y12_W1BEG;
wire[7:0] Tile_X3Y12_W2BEG;
wire[7:0] Tile_X3Y12_W2BEGb;
wire[15:0] Tile_X3Y12_WW4BEG;
wire[11:0] Tile_X3Y12_W6BEG;
wire[0:0] Tile_X3Y12_Co;
wire[3:0] Tile_X4Y12_N1BEG;
wire[7:0] Tile_X4Y12_N2BEG;
wire[7:0] Tile_X4Y12_N2BEGb;
wire[15:0] Tile_X4Y12_N4BEG;
wire[15:0] Tile_X4Y12_NN4BEG;
wire[3:0] Tile_X4Y12_E1BEG;
wire[7:0] Tile_X4Y12_E2BEG;
wire[7:0] Tile_X4Y12_E2BEGb;
wire[15:0] Tile_X4Y12_EE4BEG;
wire[11:0] Tile_X4Y12_E6BEG;
wire[3:0] Tile_X4Y12_S1BEG;
wire[7:0] Tile_X4Y12_S2BEG;
wire[7:0] Tile_X4Y12_S2BEGb;
wire[15:0] Tile_X4Y12_S4BEG;
wire[15:0] Tile_X4Y12_SS4BEG;
wire[3:0] Tile_X4Y12_W1BEG;
wire[7:0] Tile_X4Y12_W2BEG;
wire[7:0] Tile_X4Y12_W2BEGb;
wire[15:0] Tile_X4Y12_WW4BEG;
wire[11:0] Tile_X4Y12_W6BEG;
wire[3:0] Tile_X5Y12_N1BEG;
wire[7:0] Tile_X5Y12_N2BEG;
wire[7:0] Tile_X5Y12_N2BEGb;
wire[15:0] Tile_X5Y12_N4BEG;
wire[15:0] Tile_X5Y12_NN4BEG;
wire[3:0] Tile_X5Y12_E1BEG;
wire[7:0] Tile_X5Y12_E2BEG;
wire[7:0] Tile_X5Y12_E2BEGb;
wire[15:0] Tile_X5Y12_EE4BEG;
wire[11:0] Tile_X5Y12_E6BEG;
wire[3:0] Tile_X5Y12_S1BEG;
wire[7:0] Tile_X5Y12_S2BEG;
wire[7:0] Tile_X5Y12_S2BEGb;
wire[15:0] Tile_X5Y12_S4BEG;
wire[15:0] Tile_X5Y12_SS4BEG;
wire[3:0] Tile_X5Y12_W1BEG;
wire[7:0] Tile_X5Y12_W2BEG;
wire[7:0] Tile_X5Y12_W2BEGb;
wire[15:0] Tile_X5Y12_WW4BEG;
wire[11:0] Tile_X5Y12_W6BEG;
wire[0:0] Tile_X5Y12_Co;
wire[3:0] Tile_X6Y12_N1BEG;
wire[7:0] Tile_X6Y12_N2BEG;
wire[7:0] Tile_X6Y12_N2BEGb;
wire[15:0] Tile_X6Y12_N4BEG;
wire[15:0] Tile_X6Y12_NN4BEG;
wire[3:0] Tile_X6Y12_E1BEG;
wire[7:0] Tile_X6Y12_E2BEG;
wire[7:0] Tile_X6Y12_E2BEGb;
wire[15:0] Tile_X6Y12_EE4BEG;
wire[11:0] Tile_X6Y12_E6BEG;
wire[3:0] Tile_X6Y12_S1BEG;
wire[7:0] Tile_X6Y12_S2BEG;
wire[7:0] Tile_X6Y12_S2BEGb;
wire[15:0] Tile_X6Y12_S4BEG;
wire[15:0] Tile_X6Y12_SS4BEG;
wire[3:0] Tile_X6Y12_W1BEG;
wire[7:0] Tile_X6Y12_W2BEG;
wire[7:0] Tile_X6Y12_W2BEGb;
wire[15:0] Tile_X6Y12_WW4BEG;
wire[11:0] Tile_X6Y12_W6BEG;
wire[0:0] Tile_X6Y12_Co;
wire[3:0] Tile_X7Y12_N1BEG;
wire[7:0] Tile_X7Y12_N2BEG;
wire[7:0] Tile_X7Y12_N2BEGb;
wire[15:0] Tile_X7Y12_N4BEG;
wire[15:0] Tile_X7Y12_NN4BEG;
wire[3:0] Tile_X7Y12_E1BEG;
wire[7:0] Tile_X7Y12_E2BEG;
wire[7:0] Tile_X7Y12_E2BEGb;
wire[15:0] Tile_X7Y12_EE4BEG;
wire[11:0] Tile_X7Y12_E6BEG;
wire[3:0] Tile_X7Y12_S1BEG;
wire[7:0] Tile_X7Y12_S2BEG;
wire[7:0] Tile_X7Y12_S2BEGb;
wire[15:0] Tile_X7Y12_S4BEG;
wire[15:0] Tile_X7Y12_SS4BEG;
wire[3:0] Tile_X7Y12_W1BEG;
wire[7:0] Tile_X7Y12_W2BEG;
wire[7:0] Tile_X7Y12_W2BEGb;
wire[15:0] Tile_X7Y12_WW4BEG;
wire[11:0] Tile_X7Y12_W6BEG;
wire[9:0] Tile_X7Y12_bot2top;
wire[3:0] Tile_X8Y12_N1BEG;
wire[7:0] Tile_X8Y12_N2BEG;
wire[7:0] Tile_X8Y12_N2BEGb;
wire[15:0] Tile_X8Y12_N4BEG;
wire[15:0] Tile_X8Y12_NN4BEG;
wire[3:0] Tile_X8Y12_E1BEG;
wire[7:0] Tile_X8Y12_E2BEG;
wire[7:0] Tile_X8Y12_E2BEGb;
wire[15:0] Tile_X8Y12_EE4BEG;
wire[11:0] Tile_X8Y12_E6BEG;
wire[3:0] Tile_X8Y12_S1BEG;
wire[7:0] Tile_X8Y12_S2BEG;
wire[7:0] Tile_X8Y12_S2BEGb;
wire[15:0] Tile_X8Y12_S4BEG;
wire[15:0] Tile_X8Y12_SS4BEG;
wire[3:0] Tile_X8Y12_W1BEG;
wire[7:0] Tile_X8Y12_W2BEG;
wire[7:0] Tile_X8Y12_W2BEGb;
wire[15:0] Tile_X8Y12_WW4BEG;
wire[11:0] Tile_X8Y12_W6BEG;
wire[0:0] Tile_X8Y12_Co;
wire[3:0] Tile_X9Y12_N1BEG;
wire[7:0] Tile_X9Y12_N2BEG;
wire[7:0] Tile_X9Y12_N2BEGb;
wire[15:0] Tile_X9Y12_N4BEG;
wire[15:0] Tile_X9Y12_NN4BEG;
wire[3:0] Tile_X9Y12_E1BEG;
wire[7:0] Tile_X9Y12_E2BEG;
wire[7:0] Tile_X9Y12_E2BEGb;
wire[15:0] Tile_X9Y12_EE4BEG;
wire[11:0] Tile_X9Y12_E6BEG;
wire[3:0] Tile_X9Y12_S1BEG;
wire[7:0] Tile_X9Y12_S2BEG;
wire[7:0] Tile_X9Y12_S2BEGb;
wire[15:0] Tile_X9Y12_S4BEG;
wire[15:0] Tile_X9Y12_SS4BEG;
wire[3:0] Tile_X9Y12_W1BEG;
wire[7:0] Tile_X9Y12_W2BEG;
wire[7:0] Tile_X9Y12_W2BEGb;
wire[15:0] Tile_X9Y12_WW4BEG;
wire[11:0] Tile_X9Y12_W6BEG;
wire[0:0] Tile_X9Y12_Co;
wire[3:0] Tile_X10Y12_N1BEG;
wire[7:0] Tile_X10Y12_N2BEG;
wire[7:0] Tile_X10Y12_N2BEGb;
wire[15:0] Tile_X10Y12_N4BEG;
wire[3:0] Tile_X10Y12_S1BEG;
wire[7:0] Tile_X10Y12_S2BEG;
wire[7:0] Tile_X10Y12_S2BEGb;
wire[15:0] Tile_X10Y12_S4BEG;
wire[3:0] Tile_X10Y12_W1BEG;
wire[7:0] Tile_X10Y12_W2BEG;
wire[7:0] Tile_X10Y12_W2BEGb;
wire[15:0] Tile_X10Y12_WW4BEG;
wire[11:0] Tile_X10Y12_W6BEG;
wire[15:0] Tile_X10Y12_bot2top_DOUT;
wire[3:0] Tile_X0Y13_E1BEG;
wire[7:0] Tile_X0Y13_E2BEG;
wire[7:0] Tile_X0Y13_E2BEGb;
wire[15:0] Tile_X0Y13_EE4BEG;
wire[11:0] Tile_X0Y13_E6BEG;
wire[3:0] Tile_X1Y13_N1BEG;
wire[7:0] Tile_X1Y13_N2BEG;
wire[7:0] Tile_X1Y13_N2BEGb;
wire[15:0] Tile_X1Y13_N4BEG;
wire[15:0] Tile_X1Y13_NN4BEG;
wire[3:0] Tile_X1Y13_E1BEG;
wire[7:0] Tile_X1Y13_E2BEG;
wire[7:0] Tile_X1Y13_E2BEGb;
wire[15:0] Tile_X1Y13_EE4BEG;
wire[11:0] Tile_X1Y13_E6BEG;
wire[3:0] Tile_X1Y13_S1BEG;
wire[7:0] Tile_X1Y13_S2BEG;
wire[7:0] Tile_X1Y13_S2BEGb;
wire[15:0] Tile_X1Y13_S4BEG;
wire[15:0] Tile_X1Y13_SS4BEG;
wire[3:0] Tile_X1Y13_W1BEG;
wire[7:0] Tile_X1Y13_W2BEG;
wire[7:0] Tile_X1Y13_W2BEGb;
wire[15:0] Tile_X1Y13_WW4BEG;
wire[11:0] Tile_X1Y13_W6BEG;
wire[0:0] Tile_X1Y13_Co;
wire[3:0] Tile_X2Y13_N1BEG;
wire[7:0] Tile_X2Y13_N2BEG;
wire[7:0] Tile_X2Y13_N2BEGb;
wire[15:0] Tile_X2Y13_N4BEG;
wire[15:0] Tile_X2Y13_NN4BEG;
wire[3:0] Tile_X2Y13_E1BEG;
wire[7:0] Tile_X2Y13_E2BEG;
wire[7:0] Tile_X2Y13_E2BEGb;
wire[15:0] Tile_X2Y13_EE4BEG;
wire[11:0] Tile_X2Y13_E6BEG;
wire[3:0] Tile_X2Y13_S1BEG;
wire[7:0] Tile_X2Y13_S2BEG;
wire[7:0] Tile_X2Y13_S2BEGb;
wire[15:0] Tile_X2Y13_S4BEG;
wire[15:0] Tile_X2Y13_SS4BEG;
wire[3:0] Tile_X2Y13_W1BEG;
wire[7:0] Tile_X2Y13_W2BEG;
wire[7:0] Tile_X2Y13_W2BEGb;
wire[15:0] Tile_X2Y13_WW4BEG;
wire[11:0] Tile_X2Y13_W6BEG;
wire[0:0] Tile_X2Y13_Co;
wire[3:0] Tile_X3Y13_N1BEG;
wire[7:0] Tile_X3Y13_N2BEG;
wire[7:0] Tile_X3Y13_N2BEGb;
wire[15:0] Tile_X3Y13_N4BEG;
wire[15:0] Tile_X3Y13_NN4BEG;
wire[3:0] Tile_X3Y13_E1BEG;
wire[7:0] Tile_X3Y13_E2BEG;
wire[7:0] Tile_X3Y13_E2BEGb;
wire[15:0] Tile_X3Y13_EE4BEG;
wire[11:0] Tile_X3Y13_E6BEG;
wire[3:0] Tile_X3Y13_S1BEG;
wire[7:0] Tile_X3Y13_S2BEG;
wire[7:0] Tile_X3Y13_S2BEGb;
wire[15:0] Tile_X3Y13_S4BEG;
wire[15:0] Tile_X3Y13_SS4BEG;
wire[3:0] Tile_X3Y13_W1BEG;
wire[7:0] Tile_X3Y13_W2BEG;
wire[7:0] Tile_X3Y13_W2BEGb;
wire[15:0] Tile_X3Y13_WW4BEG;
wire[11:0] Tile_X3Y13_W6BEG;
wire[0:0] Tile_X3Y13_Co;
wire[3:0] Tile_X4Y13_N1BEG;
wire[7:0] Tile_X4Y13_N2BEG;
wire[7:0] Tile_X4Y13_N2BEGb;
wire[15:0] Tile_X4Y13_N4BEG;
wire[15:0] Tile_X4Y13_NN4BEG;
wire[3:0] Tile_X4Y13_E1BEG;
wire[7:0] Tile_X4Y13_E2BEG;
wire[7:0] Tile_X4Y13_E2BEGb;
wire[15:0] Tile_X4Y13_EE4BEG;
wire[11:0] Tile_X4Y13_E6BEG;
wire[3:0] Tile_X4Y13_S1BEG;
wire[7:0] Tile_X4Y13_S2BEG;
wire[7:0] Tile_X4Y13_S2BEGb;
wire[15:0] Tile_X4Y13_S4BEG;
wire[15:0] Tile_X4Y13_SS4BEG;
wire[3:0] Tile_X4Y13_W1BEG;
wire[7:0] Tile_X4Y13_W2BEG;
wire[7:0] Tile_X4Y13_W2BEGb;
wire[15:0] Tile_X4Y13_WW4BEG;
wire[11:0] Tile_X4Y13_W6BEG;
wire[3:0] Tile_X5Y13_N1BEG;
wire[7:0] Tile_X5Y13_N2BEG;
wire[7:0] Tile_X5Y13_N2BEGb;
wire[15:0] Tile_X5Y13_N4BEG;
wire[15:0] Tile_X5Y13_NN4BEG;
wire[3:0] Tile_X5Y13_E1BEG;
wire[7:0] Tile_X5Y13_E2BEG;
wire[7:0] Tile_X5Y13_E2BEGb;
wire[15:0] Tile_X5Y13_EE4BEG;
wire[11:0] Tile_X5Y13_E6BEG;
wire[3:0] Tile_X5Y13_S1BEG;
wire[7:0] Tile_X5Y13_S2BEG;
wire[7:0] Tile_X5Y13_S2BEGb;
wire[15:0] Tile_X5Y13_S4BEG;
wire[15:0] Tile_X5Y13_SS4BEG;
wire[3:0] Tile_X5Y13_W1BEG;
wire[7:0] Tile_X5Y13_W2BEG;
wire[7:0] Tile_X5Y13_W2BEGb;
wire[15:0] Tile_X5Y13_WW4BEG;
wire[11:0] Tile_X5Y13_W6BEG;
wire[0:0] Tile_X5Y13_Co;
wire[3:0] Tile_X6Y13_N1BEG;
wire[7:0] Tile_X6Y13_N2BEG;
wire[7:0] Tile_X6Y13_N2BEGb;
wire[15:0] Tile_X6Y13_N4BEG;
wire[15:0] Tile_X6Y13_NN4BEG;
wire[3:0] Tile_X6Y13_E1BEG;
wire[7:0] Tile_X6Y13_E2BEG;
wire[7:0] Tile_X6Y13_E2BEGb;
wire[15:0] Tile_X6Y13_EE4BEG;
wire[11:0] Tile_X6Y13_E6BEG;
wire[3:0] Tile_X6Y13_S1BEG;
wire[7:0] Tile_X6Y13_S2BEG;
wire[7:0] Tile_X6Y13_S2BEGb;
wire[15:0] Tile_X6Y13_S4BEG;
wire[15:0] Tile_X6Y13_SS4BEG;
wire[3:0] Tile_X6Y13_W1BEG;
wire[7:0] Tile_X6Y13_W2BEG;
wire[7:0] Tile_X6Y13_W2BEGb;
wire[15:0] Tile_X6Y13_WW4BEG;
wire[11:0] Tile_X6Y13_W6BEG;
wire[0:0] Tile_X6Y13_Co;
wire[3:0] Tile_X7Y13_N1BEG;
wire[7:0] Tile_X7Y13_N2BEG;
wire[7:0] Tile_X7Y13_N2BEGb;
wire[15:0] Tile_X7Y13_N4BEG;
wire[15:0] Tile_X7Y13_NN4BEG;
wire[3:0] Tile_X7Y13_E1BEG;
wire[7:0] Tile_X7Y13_E2BEG;
wire[7:0] Tile_X7Y13_E2BEGb;
wire[15:0] Tile_X7Y13_EE4BEG;
wire[11:0] Tile_X7Y13_E6BEG;
wire[3:0] Tile_X7Y13_S1BEG;
wire[7:0] Tile_X7Y13_S2BEG;
wire[7:0] Tile_X7Y13_S2BEGb;
wire[15:0] Tile_X7Y13_S4BEG;
wire[15:0] Tile_X7Y13_SS4BEG;
wire[3:0] Tile_X7Y13_W1BEG;
wire[7:0] Tile_X7Y13_W2BEG;
wire[7:0] Tile_X7Y13_W2BEGb;
wire[15:0] Tile_X7Y13_WW4BEG;
wire[11:0] Tile_X7Y13_W6BEG;
wire[17:0] Tile_X7Y13_top2bot;
wire[3:0] Tile_X8Y13_N1BEG;
wire[7:0] Tile_X8Y13_N2BEG;
wire[7:0] Tile_X8Y13_N2BEGb;
wire[15:0] Tile_X8Y13_N4BEG;
wire[15:0] Tile_X8Y13_NN4BEG;
wire[3:0] Tile_X8Y13_E1BEG;
wire[7:0] Tile_X8Y13_E2BEG;
wire[7:0] Tile_X8Y13_E2BEGb;
wire[15:0] Tile_X8Y13_EE4BEG;
wire[11:0] Tile_X8Y13_E6BEG;
wire[3:0] Tile_X8Y13_S1BEG;
wire[7:0] Tile_X8Y13_S2BEG;
wire[7:0] Tile_X8Y13_S2BEGb;
wire[15:0] Tile_X8Y13_S4BEG;
wire[15:0] Tile_X8Y13_SS4BEG;
wire[3:0] Tile_X8Y13_W1BEG;
wire[7:0] Tile_X8Y13_W2BEG;
wire[7:0] Tile_X8Y13_W2BEGb;
wire[15:0] Tile_X8Y13_WW4BEG;
wire[11:0] Tile_X8Y13_W6BEG;
wire[0:0] Tile_X8Y13_Co;
wire[3:0] Tile_X9Y13_N1BEG;
wire[7:0] Tile_X9Y13_N2BEG;
wire[7:0] Tile_X9Y13_N2BEGb;
wire[15:0] Tile_X9Y13_N4BEG;
wire[15:0] Tile_X9Y13_NN4BEG;
wire[3:0] Tile_X9Y13_E1BEG;
wire[7:0] Tile_X9Y13_E2BEG;
wire[7:0] Tile_X9Y13_E2BEGb;
wire[15:0] Tile_X9Y13_EE4BEG;
wire[11:0] Tile_X9Y13_E6BEG;
wire[3:0] Tile_X9Y13_S1BEG;
wire[7:0] Tile_X9Y13_S2BEG;
wire[7:0] Tile_X9Y13_S2BEGb;
wire[15:0] Tile_X9Y13_S4BEG;
wire[15:0] Tile_X9Y13_SS4BEG;
wire[3:0] Tile_X9Y13_W1BEG;
wire[7:0] Tile_X9Y13_W2BEG;
wire[7:0] Tile_X9Y13_W2BEGb;
wire[15:0] Tile_X9Y13_WW4BEG;
wire[11:0] Tile_X9Y13_W6BEG;
wire[0:0] Tile_X9Y13_Co;
wire[3:0] Tile_X10Y13_N1BEG;
wire[7:0] Tile_X10Y13_N2BEG;
wire[7:0] Tile_X10Y13_N2BEGb;
wire[15:0] Tile_X10Y13_N4BEG;
wire[3:0] Tile_X10Y13_S1BEG;
wire[7:0] Tile_X10Y13_S2BEG;
wire[7:0] Tile_X10Y13_S2BEGb;
wire[15:0] Tile_X10Y13_S4BEG;
wire[3:0] Tile_X10Y13_W1BEG;
wire[7:0] Tile_X10Y13_W2BEG;
wire[7:0] Tile_X10Y13_W2BEGb;
wire[15:0] Tile_X10Y13_WW4BEG;
wire[11:0] Tile_X10Y13_W6BEG;
wire[15:0] Tile_X10Y13_top2bot_DIN;
wire[15:0] Tile_X10Y13_top2bot_BM;
wire[4:0] Tile_X10Y13_top2bot_ADDR;
wire[3:0] Tile_X0Y14_E1BEG;
wire[7:0] Tile_X0Y14_E2BEG;
wire[7:0] Tile_X0Y14_E2BEGb;
wire[15:0] Tile_X0Y14_EE4BEG;
wire[11:0] Tile_X0Y14_E6BEG;
wire[3:0] Tile_X1Y14_N1BEG;
wire[7:0] Tile_X1Y14_N2BEG;
wire[7:0] Tile_X1Y14_N2BEGb;
wire[15:0] Tile_X1Y14_N4BEG;
wire[15:0] Tile_X1Y14_NN4BEG;
wire[3:0] Tile_X1Y14_E1BEG;
wire[7:0] Tile_X1Y14_E2BEG;
wire[7:0] Tile_X1Y14_E2BEGb;
wire[15:0] Tile_X1Y14_EE4BEG;
wire[11:0] Tile_X1Y14_E6BEG;
wire[3:0] Tile_X1Y14_S1BEG;
wire[7:0] Tile_X1Y14_S2BEG;
wire[7:0] Tile_X1Y14_S2BEGb;
wire[15:0] Tile_X1Y14_S4BEG;
wire[15:0] Tile_X1Y14_SS4BEG;
wire[3:0] Tile_X1Y14_W1BEG;
wire[7:0] Tile_X1Y14_W2BEG;
wire[7:0] Tile_X1Y14_W2BEGb;
wire[15:0] Tile_X1Y14_WW4BEG;
wire[11:0] Tile_X1Y14_W6BEG;
wire[0:0] Tile_X1Y14_Co;
wire[3:0] Tile_X2Y14_N1BEG;
wire[7:0] Tile_X2Y14_N2BEG;
wire[7:0] Tile_X2Y14_N2BEGb;
wire[15:0] Tile_X2Y14_N4BEG;
wire[15:0] Tile_X2Y14_NN4BEG;
wire[3:0] Tile_X2Y14_E1BEG;
wire[7:0] Tile_X2Y14_E2BEG;
wire[7:0] Tile_X2Y14_E2BEGb;
wire[15:0] Tile_X2Y14_EE4BEG;
wire[11:0] Tile_X2Y14_E6BEG;
wire[3:0] Tile_X2Y14_S1BEG;
wire[7:0] Tile_X2Y14_S2BEG;
wire[7:0] Tile_X2Y14_S2BEGb;
wire[15:0] Tile_X2Y14_S4BEG;
wire[15:0] Tile_X2Y14_SS4BEG;
wire[3:0] Tile_X2Y14_W1BEG;
wire[7:0] Tile_X2Y14_W2BEG;
wire[7:0] Tile_X2Y14_W2BEGb;
wire[15:0] Tile_X2Y14_WW4BEG;
wire[11:0] Tile_X2Y14_W6BEG;
wire[0:0] Tile_X2Y14_Co;
wire[3:0] Tile_X3Y14_N1BEG;
wire[7:0] Tile_X3Y14_N2BEG;
wire[7:0] Tile_X3Y14_N2BEGb;
wire[15:0] Tile_X3Y14_N4BEG;
wire[15:0] Tile_X3Y14_NN4BEG;
wire[3:0] Tile_X3Y14_E1BEG;
wire[7:0] Tile_X3Y14_E2BEG;
wire[7:0] Tile_X3Y14_E2BEGb;
wire[15:0] Tile_X3Y14_EE4BEG;
wire[11:0] Tile_X3Y14_E6BEG;
wire[3:0] Tile_X3Y14_S1BEG;
wire[7:0] Tile_X3Y14_S2BEG;
wire[7:0] Tile_X3Y14_S2BEGb;
wire[15:0] Tile_X3Y14_S4BEG;
wire[15:0] Tile_X3Y14_SS4BEG;
wire[3:0] Tile_X3Y14_W1BEG;
wire[7:0] Tile_X3Y14_W2BEG;
wire[7:0] Tile_X3Y14_W2BEGb;
wire[15:0] Tile_X3Y14_WW4BEG;
wire[11:0] Tile_X3Y14_W6BEG;
wire[0:0] Tile_X3Y14_Co;
wire[3:0] Tile_X4Y14_N1BEG;
wire[7:0] Tile_X4Y14_N2BEG;
wire[7:0] Tile_X4Y14_N2BEGb;
wire[15:0] Tile_X4Y14_N4BEG;
wire[15:0] Tile_X4Y14_NN4BEG;
wire[3:0] Tile_X4Y14_E1BEG;
wire[7:0] Tile_X4Y14_E2BEG;
wire[7:0] Tile_X4Y14_E2BEGb;
wire[15:0] Tile_X4Y14_EE4BEG;
wire[11:0] Tile_X4Y14_E6BEG;
wire[3:0] Tile_X4Y14_S1BEG;
wire[7:0] Tile_X4Y14_S2BEG;
wire[7:0] Tile_X4Y14_S2BEGb;
wire[15:0] Tile_X4Y14_S4BEG;
wire[15:0] Tile_X4Y14_SS4BEG;
wire[3:0] Tile_X4Y14_W1BEG;
wire[7:0] Tile_X4Y14_W2BEG;
wire[7:0] Tile_X4Y14_W2BEGb;
wire[15:0] Tile_X4Y14_WW4BEG;
wire[11:0] Tile_X4Y14_W6BEG;
wire[3:0] Tile_X5Y14_N1BEG;
wire[7:0] Tile_X5Y14_N2BEG;
wire[7:0] Tile_X5Y14_N2BEGb;
wire[15:0] Tile_X5Y14_N4BEG;
wire[15:0] Tile_X5Y14_NN4BEG;
wire[3:0] Tile_X5Y14_E1BEG;
wire[7:0] Tile_X5Y14_E2BEG;
wire[7:0] Tile_X5Y14_E2BEGb;
wire[15:0] Tile_X5Y14_EE4BEG;
wire[11:0] Tile_X5Y14_E6BEG;
wire[3:0] Tile_X5Y14_S1BEG;
wire[7:0] Tile_X5Y14_S2BEG;
wire[7:0] Tile_X5Y14_S2BEGb;
wire[15:0] Tile_X5Y14_S4BEG;
wire[15:0] Tile_X5Y14_SS4BEG;
wire[3:0] Tile_X5Y14_W1BEG;
wire[7:0] Tile_X5Y14_W2BEG;
wire[7:0] Tile_X5Y14_W2BEGb;
wire[15:0] Tile_X5Y14_WW4BEG;
wire[11:0] Tile_X5Y14_W6BEG;
wire[0:0] Tile_X5Y14_Co;
wire[3:0] Tile_X6Y14_N1BEG;
wire[7:0] Tile_X6Y14_N2BEG;
wire[7:0] Tile_X6Y14_N2BEGb;
wire[15:0] Tile_X6Y14_N4BEG;
wire[15:0] Tile_X6Y14_NN4BEG;
wire[3:0] Tile_X6Y14_E1BEG;
wire[7:0] Tile_X6Y14_E2BEG;
wire[7:0] Tile_X6Y14_E2BEGb;
wire[15:0] Tile_X6Y14_EE4BEG;
wire[11:0] Tile_X6Y14_E6BEG;
wire[3:0] Tile_X6Y14_S1BEG;
wire[7:0] Tile_X6Y14_S2BEG;
wire[7:0] Tile_X6Y14_S2BEGb;
wire[15:0] Tile_X6Y14_S4BEG;
wire[15:0] Tile_X6Y14_SS4BEG;
wire[3:0] Tile_X6Y14_W1BEG;
wire[7:0] Tile_X6Y14_W2BEG;
wire[7:0] Tile_X6Y14_W2BEGb;
wire[15:0] Tile_X6Y14_WW4BEG;
wire[11:0] Tile_X6Y14_W6BEG;
wire[0:0] Tile_X6Y14_Co;
wire[3:0] Tile_X7Y14_N1BEG;
wire[7:0] Tile_X7Y14_N2BEG;
wire[7:0] Tile_X7Y14_N2BEGb;
wire[15:0] Tile_X7Y14_N4BEG;
wire[15:0] Tile_X7Y14_NN4BEG;
wire[3:0] Tile_X7Y14_E1BEG;
wire[7:0] Tile_X7Y14_E2BEG;
wire[7:0] Tile_X7Y14_E2BEGb;
wire[15:0] Tile_X7Y14_EE4BEG;
wire[11:0] Tile_X7Y14_E6BEG;
wire[3:0] Tile_X7Y14_S1BEG;
wire[7:0] Tile_X7Y14_S2BEG;
wire[7:0] Tile_X7Y14_S2BEGb;
wire[15:0] Tile_X7Y14_S4BEG;
wire[15:0] Tile_X7Y14_SS4BEG;
wire[3:0] Tile_X7Y14_W1BEG;
wire[7:0] Tile_X7Y14_W2BEG;
wire[7:0] Tile_X7Y14_W2BEGb;
wire[15:0] Tile_X7Y14_WW4BEG;
wire[11:0] Tile_X7Y14_W6BEG;
wire[9:0] Tile_X7Y14_bot2top;
wire[3:0] Tile_X8Y14_N1BEG;
wire[7:0] Tile_X8Y14_N2BEG;
wire[7:0] Tile_X8Y14_N2BEGb;
wire[15:0] Tile_X8Y14_N4BEG;
wire[15:0] Tile_X8Y14_NN4BEG;
wire[3:0] Tile_X8Y14_E1BEG;
wire[7:0] Tile_X8Y14_E2BEG;
wire[7:0] Tile_X8Y14_E2BEGb;
wire[15:0] Tile_X8Y14_EE4BEG;
wire[11:0] Tile_X8Y14_E6BEG;
wire[3:0] Tile_X8Y14_S1BEG;
wire[7:0] Tile_X8Y14_S2BEG;
wire[7:0] Tile_X8Y14_S2BEGb;
wire[15:0] Tile_X8Y14_S4BEG;
wire[15:0] Tile_X8Y14_SS4BEG;
wire[3:0] Tile_X8Y14_W1BEG;
wire[7:0] Tile_X8Y14_W2BEG;
wire[7:0] Tile_X8Y14_W2BEGb;
wire[15:0] Tile_X8Y14_WW4BEG;
wire[11:0] Tile_X8Y14_W6BEG;
wire[0:0] Tile_X8Y14_Co;
wire[3:0] Tile_X9Y14_N1BEG;
wire[7:0] Tile_X9Y14_N2BEG;
wire[7:0] Tile_X9Y14_N2BEGb;
wire[15:0] Tile_X9Y14_N4BEG;
wire[15:0] Tile_X9Y14_NN4BEG;
wire[3:0] Tile_X9Y14_E1BEG;
wire[7:0] Tile_X9Y14_E2BEG;
wire[7:0] Tile_X9Y14_E2BEGb;
wire[15:0] Tile_X9Y14_EE4BEG;
wire[11:0] Tile_X9Y14_E6BEG;
wire[3:0] Tile_X9Y14_S1BEG;
wire[7:0] Tile_X9Y14_S2BEG;
wire[7:0] Tile_X9Y14_S2BEGb;
wire[15:0] Tile_X9Y14_S4BEG;
wire[15:0] Tile_X9Y14_SS4BEG;
wire[3:0] Tile_X9Y14_W1BEG;
wire[7:0] Tile_X9Y14_W2BEG;
wire[7:0] Tile_X9Y14_W2BEGb;
wire[15:0] Tile_X9Y14_WW4BEG;
wire[11:0] Tile_X9Y14_W6BEG;
wire[0:0] Tile_X9Y14_Co;
wire[3:0] Tile_X10Y14_N1BEG;
wire[7:0] Tile_X10Y14_N2BEG;
wire[7:0] Tile_X10Y14_N2BEGb;
wire[15:0] Tile_X10Y14_N4BEG;
wire[3:0] Tile_X10Y14_S1BEG;
wire[7:0] Tile_X10Y14_S2BEG;
wire[7:0] Tile_X10Y14_S2BEGb;
wire[15:0] Tile_X10Y14_S4BEG;
wire[3:0] Tile_X10Y14_W1BEG;
wire[7:0] Tile_X10Y14_W2BEG;
wire[7:0] Tile_X10Y14_W2BEGb;
wire[15:0] Tile_X10Y14_WW4BEG;
wire[11:0] Tile_X10Y14_W6BEG;
wire[15:0] Tile_X10Y14_bot2top_DOUT;
wire[3:0] Tile_X1Y15_N1BEG;
wire[7:0] Tile_X1Y15_N2BEG;
wire[7:0] Tile_X1Y15_N2BEGb;
wire[15:0] Tile_X1Y15_N4BEG;
wire[15:0] Tile_X1Y15_NN4BEG;
wire[0:0] Tile_X1Y15_Co;
wire[3:0] Tile_X2Y15_N1BEG;
wire[7:0] Tile_X2Y15_N2BEG;
wire[7:0] Tile_X2Y15_N2BEGb;
wire[15:0] Tile_X2Y15_N4BEG;
wire[15:0] Tile_X2Y15_NN4BEG;
wire[0:0] Tile_X2Y15_Co;
wire[3:0] Tile_X3Y15_N1BEG;
wire[7:0] Tile_X3Y15_N2BEG;
wire[7:0] Tile_X3Y15_N2BEGb;
wire[15:0] Tile_X3Y15_N4BEG;
wire[15:0] Tile_X3Y15_NN4BEG;
wire[0:0] Tile_X3Y15_Co;
wire[3:0] Tile_X4Y15_N1BEG;
wire[7:0] Tile_X4Y15_N2BEG;
wire[7:0] Tile_X4Y15_N2BEGb;
wire[15:0] Tile_X4Y15_N4BEG;
wire[15:0] Tile_X4Y15_NN4BEG;
wire[3:0] Tile_X5Y15_N1BEG;
wire[7:0] Tile_X5Y15_N2BEG;
wire[7:0] Tile_X5Y15_N2BEGb;
wire[15:0] Tile_X5Y15_N4BEG;
wire[15:0] Tile_X5Y15_NN4BEG;
wire[0:0] Tile_X5Y15_Co;
wire[3:0] Tile_X6Y15_N1BEG;
wire[7:0] Tile_X6Y15_N2BEG;
wire[7:0] Tile_X6Y15_N2BEGb;
wire[15:0] Tile_X6Y15_N4BEG;
wire[15:0] Tile_X6Y15_NN4BEG;
wire[0:0] Tile_X6Y15_Co;
wire[3:0] Tile_X7Y15_N1BEG;
wire[7:0] Tile_X7Y15_N2BEG;
wire[7:0] Tile_X7Y15_N2BEGb;
wire[15:0] Tile_X7Y15_N4BEG;
wire[15:0] Tile_X7Y15_NN4BEG;
wire[3:0] Tile_X8Y15_N1BEG;
wire[7:0] Tile_X8Y15_N2BEG;
wire[7:0] Tile_X8Y15_N2BEGb;
wire[15:0] Tile_X8Y15_N4BEG;
wire[15:0] Tile_X8Y15_NN4BEG;
wire[0:0] Tile_X8Y15_Co;
wire[3:0] Tile_X9Y15_N1BEG;
wire[7:0] Tile_X9Y15_N2BEG;
wire[7:0] Tile_X9Y15_N2BEGb;
wire[15:0] Tile_X9Y15_N4BEG;
wire[15:0] Tile_X9Y15_NN4BEG;
wire[0:0] Tile_X9Y15_Co;
wire[3:0] Tile_X10Y15_N1BEG;
wire[7:0] Tile_X10Y15_N2BEG;
wire[7:0] Tile_X10Y15_N2BEGb;
wire[15:0] Tile_X10Y15_N4BEG;

assign Row_Y0_FrameData = FrameData[FrameBitsPerRow*(0+1)-1:FrameBitsPerRow*0];
assign Row_Y1_FrameData = FrameData[FrameBitsPerRow*(1+1)-1:FrameBitsPerRow*1];
assign Row_Y2_FrameData = FrameData[FrameBitsPerRow*(2+1)-1:FrameBitsPerRow*2];
assign Row_Y3_FrameData = FrameData[FrameBitsPerRow*(3+1)-1:FrameBitsPerRow*3];
assign Row_Y4_FrameData = FrameData[FrameBitsPerRow*(4+1)-1:FrameBitsPerRow*4];
assign Row_Y5_FrameData = FrameData[FrameBitsPerRow*(5+1)-1:FrameBitsPerRow*5];
assign Row_Y6_FrameData = FrameData[FrameBitsPerRow*(6+1)-1:FrameBitsPerRow*6];
assign Row_Y7_FrameData = FrameData[FrameBitsPerRow*(7+1)-1:FrameBitsPerRow*7];
assign Row_Y8_FrameData = FrameData[FrameBitsPerRow*(8+1)-1:FrameBitsPerRow*8];
assign Row_Y9_FrameData = FrameData[FrameBitsPerRow*(9+1)-1:FrameBitsPerRow*9];
assign Row_Y10_FrameData = FrameData[FrameBitsPerRow*(10+1)-1:FrameBitsPerRow*10];
assign Row_Y11_FrameData = FrameData[FrameBitsPerRow*(11+1)-1:FrameBitsPerRow*11];
assign Row_Y12_FrameData = FrameData[FrameBitsPerRow*(12+1)-1:FrameBitsPerRow*12];
assign Row_Y13_FrameData = FrameData[FrameBitsPerRow*(13+1)-1:FrameBitsPerRow*13];
assign Row_Y14_FrameData = FrameData[FrameBitsPerRow*(14+1)-1:FrameBitsPerRow*14];
assign Row_Y15_FrameData = FrameData[FrameBitsPerRow*(15+1)-1:FrameBitsPerRow*15];
assign Column_X0_FrameStrobe = FrameStrobe[MaxFramesPerCol*(0+1)-1:MaxFramesPerCol*0];
assign Column_X1_FrameStrobe = FrameStrobe[MaxFramesPerCol*(1+1)-1:MaxFramesPerCol*1];
assign Column_X2_FrameStrobe = FrameStrobe[MaxFramesPerCol*(2+1)-1:MaxFramesPerCol*2];
assign Column_X3_FrameStrobe = FrameStrobe[MaxFramesPerCol*(3+1)-1:MaxFramesPerCol*3];
assign Column_X4_FrameStrobe = FrameStrobe[MaxFramesPerCol*(4+1)-1:MaxFramesPerCol*4];
assign Column_X5_FrameStrobe = FrameStrobe[MaxFramesPerCol*(5+1)-1:MaxFramesPerCol*5];
assign Column_X6_FrameStrobe = FrameStrobe[MaxFramesPerCol*(6+1)-1:MaxFramesPerCol*6];
assign Column_X7_FrameStrobe = FrameStrobe[MaxFramesPerCol*(7+1)-1:MaxFramesPerCol*7];
assign Column_X8_FrameStrobe = FrameStrobe[MaxFramesPerCol*(8+1)-1:MaxFramesPerCol*8];
assign Column_X9_FrameStrobe = FrameStrobe[MaxFramesPerCol*(9+1)-1:MaxFramesPerCol*9];
assign Column_X10_FrameStrobe = FrameStrobe[MaxFramesPerCol*(10+1)-1:MaxFramesPerCol*10];

 //tile IO port will get directly connected to top-level tile module
N_IO Tile_X1Y0_N_IO (
    .N1END(Tile_X1Y1_N1BEG),
    .N2MID(Tile_X1Y1_N2BEG),
    .N2END(Tile_X1Y1_N2BEGb),
    .N4END(Tile_X1Y1_N4BEG),
    .NN4END(Tile_X1Y1_NN4BEG),
    .Ci(Tile_X1Y1_Co),
    .S1BEG(Tile_X1Y0_S1BEG),
    .S2BEG(Tile_X1Y0_S2BEG),
    .S2BEGb(Tile_X1Y0_S2BEGb),
    .S4BEG(Tile_X1Y0_S4BEG),
    .SS4BEG(Tile_X1Y0_SS4BEG),
    .A_O_top(Tile_X1Y0_A_O_top),
    .A_I_top(Tile_X1Y0_A_I_top),
    .A_T_top(Tile_X1Y0_A_T_top),
    .B_O_top(Tile_X1Y0_B_O_top),
    .B_I_top(Tile_X1Y0_B_I_top),
    .B_T_top(Tile_X1Y0_B_T_top),
    .A_config_C_bit0(Tile_X1Y0_A_config_C_bit0),
    .A_config_C_bit1(Tile_X1Y0_A_config_C_bit1),
    .A_config_C_bit2(Tile_X1Y0_A_config_C_bit2),
    .A_config_C_bit3(Tile_X1Y0_A_config_C_bit3),
    .B_config_C_bit0(Tile_X1Y0_B_config_C_bit0),
    .B_config_C_bit1(Tile_X1Y0_B_config_C_bit1),
    .B_config_C_bit2(Tile_X1Y0_B_config_C_bit2),
    .B_config_C_bit3(Tile_X1Y0_B_config_C_bit3),
    .UserCLK(Tile_X1Y1_UserCLKo),
    .UserCLKo(Tile_X1Y0_UserCLKo),
    .FrameData(Row_Y0_FrameData),
    .FrameData_O(Tile_X1Y0_FrameData_O),
    .FrameStrobe(Tile_X1Y1_FrameStrobe_O),
    .FrameStrobe_O(Tile_X1Y0_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
N_IO Tile_X2Y0_N_IO (
    .N1END(Tile_X2Y1_N1BEG),
    .N2MID(Tile_X2Y1_N2BEG),
    .N2END(Tile_X2Y1_N2BEGb),
    .N4END(Tile_X2Y1_N4BEG),
    .NN4END(Tile_X2Y1_NN4BEG),
    .Ci(Tile_X2Y1_Co),
    .S1BEG(Tile_X2Y0_S1BEG),
    .S2BEG(Tile_X2Y0_S2BEG),
    .S2BEGb(Tile_X2Y0_S2BEGb),
    .S4BEG(Tile_X2Y0_S4BEG),
    .SS4BEG(Tile_X2Y0_SS4BEG),
    .A_O_top(Tile_X2Y0_A_O_top),
    .A_I_top(Tile_X2Y0_A_I_top),
    .A_T_top(Tile_X2Y0_A_T_top),
    .B_O_top(Tile_X2Y0_B_O_top),
    .B_I_top(Tile_X2Y0_B_I_top),
    .B_T_top(Tile_X2Y0_B_T_top),
    .A_config_C_bit0(Tile_X2Y0_A_config_C_bit0),
    .A_config_C_bit1(Tile_X2Y0_A_config_C_bit1),
    .A_config_C_bit2(Tile_X2Y0_A_config_C_bit2),
    .A_config_C_bit3(Tile_X2Y0_A_config_C_bit3),
    .B_config_C_bit0(Tile_X2Y0_B_config_C_bit0),
    .B_config_C_bit1(Tile_X2Y0_B_config_C_bit1),
    .B_config_C_bit2(Tile_X2Y0_B_config_C_bit2),
    .B_config_C_bit3(Tile_X2Y0_B_config_C_bit3),
    .UserCLK(Tile_X2Y1_UserCLKo),
    .UserCLKo(Tile_X2Y0_UserCLKo),
    .FrameData(Tile_X1Y0_FrameData_O),
    .FrameData_O(Tile_X2Y0_FrameData_O),
    .FrameStrobe(Tile_X2Y1_FrameStrobe_O),
    .FrameStrobe_O(Tile_X2Y0_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
N_term_single Tile_X3Y0_N_term_single (
    .N1END(Tile_X3Y1_N1BEG),
    .N2MID(Tile_X3Y1_N2BEG),
    .N2END(Tile_X3Y1_N2BEGb),
    .N4END(Tile_X3Y1_N4BEG),
    .NN4END(Tile_X3Y1_NN4BEG),
    .Ci(Tile_X3Y1_Co),
    .S1BEG(Tile_X3Y0_S1BEG),
    .S2BEG(Tile_X3Y0_S2BEG),
    .S2BEGb(Tile_X3Y0_S2BEGb),
    .S4BEG(Tile_X3Y0_S4BEG),
    .SS4BEG(Tile_X3Y0_SS4BEG),
    .UserCLK(Tile_X3Y1_UserCLKo),
    .UserCLKo(Tile_X3Y0_UserCLKo),
    .FrameData(Tile_X2Y0_FrameData_O),
    .FrameData_O(Tile_X3Y0_FrameData_O),
    .FrameStrobe(Tile_X3Y1_FrameStrobe_O),
    .FrameStrobe_O(Tile_X3Y0_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
N_term_single2 Tile_X4Y0_N_term_single2 (
    .N1END(Tile_X4Y1_N1BEG),
    .N2MID(Tile_X4Y1_N2BEG),
    .N2END(Tile_X4Y1_N2BEGb),
    .N4END(Tile_X4Y1_N4BEG),
    .NN4END(Tile_X4Y1_NN4BEG),
    .S1BEG(Tile_X4Y0_S1BEG),
    .S2BEG(Tile_X4Y0_S2BEG),
    .S2BEGb(Tile_X4Y0_S2BEGb),
    .S4BEG(Tile_X4Y0_S4BEG),
    .SS4BEG(Tile_X4Y0_SS4BEG),
    .UserCLK(Tile_X4Y1_UserCLKo),
    .UserCLKo(Tile_X4Y0_UserCLKo),
    .FrameData(Tile_X3Y0_FrameData_O),
    .FrameData_O(Tile_X4Y0_FrameData_O),
    .FrameStrobe(Tile_X4Y1_FrameStrobe_O),
    .FrameStrobe_O(Tile_X4Y0_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
N_term_single Tile_X5Y0_N_term_single (
    .N1END(Tile_X5Y1_N1BEG),
    .N2MID(Tile_X5Y1_N2BEG),
    .N2END(Tile_X5Y1_N2BEGb),
    .N4END(Tile_X5Y1_N4BEG),
    .NN4END(Tile_X5Y1_NN4BEG),
    .Ci(Tile_X5Y1_Co),
    .S1BEG(Tile_X5Y0_S1BEG),
    .S2BEG(Tile_X5Y0_S2BEG),
    .S2BEGb(Tile_X5Y0_S2BEGb),
    .S4BEG(Tile_X5Y0_S4BEG),
    .SS4BEG(Tile_X5Y0_SS4BEG),
    .UserCLK(Tile_X5Y1_UserCLKo),
    .UserCLKo(Tile_X5Y0_UserCLKo),
    .FrameData(Tile_X4Y0_FrameData_O),
    .FrameData_O(Tile_X5Y0_FrameData_O),
    .FrameStrobe(Tile_X5Y1_FrameStrobe_O),
    .FrameStrobe_O(Tile_X5Y0_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
N_term_single Tile_X6Y0_N_term_single (
    .N1END(Tile_X6Y1_N1BEG),
    .N2MID(Tile_X6Y1_N2BEG),
    .N2END(Tile_X6Y1_N2BEGb),
    .N4END(Tile_X6Y1_N4BEG),
    .NN4END(Tile_X6Y1_NN4BEG),
    .Ci(Tile_X6Y1_Co),
    .S1BEG(Tile_X6Y0_S1BEG),
    .S2BEG(Tile_X6Y0_S2BEG),
    .S2BEGb(Tile_X6Y0_S2BEGb),
    .S4BEG(Tile_X6Y0_S4BEG),
    .SS4BEG(Tile_X6Y0_SS4BEG),
    .UserCLK(Tile_X6Y1_UserCLKo),
    .UserCLKo(Tile_X6Y0_UserCLKo),
    .FrameData(Tile_X5Y0_FrameData_O),
    .FrameData_O(Tile_X6Y0_FrameData_O),
    .FrameStrobe(Tile_X6Y1_FrameStrobe_O),
    .FrameStrobe_O(Tile_X6Y0_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
N_term_DSP Tile_X7Y0_N_term_DSP (
    .N1END(Tile_X7Y1_N1BEG),
    .N2MID(Tile_X7Y1_N2BEG),
    .N2END(Tile_X7Y1_N2BEGb),
    .N4END(Tile_X7Y1_N4BEG),
    .NN4END(Tile_X7Y1_NN4BEG),
    .S1BEG(Tile_X7Y0_S1BEG),
    .S2BEG(Tile_X7Y0_S2BEG),
    .S2BEGb(Tile_X7Y0_S2BEGb),
    .S4BEG(Tile_X7Y0_S4BEG),
    .SS4BEG(Tile_X7Y0_SS4BEG),
    .UserCLK(Tile_X7Y1_UserCLKo),
    .UserCLKo(Tile_X7Y0_UserCLKo),
    .FrameData(Tile_X6Y0_FrameData_O),
    .FrameData_O(Tile_X7Y0_FrameData_O),
    .FrameStrobe(Tile_X7Y1_FrameStrobe_O),
    .FrameStrobe_O(Tile_X7Y0_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
N_term_single Tile_X8Y0_N_term_single (
    .N1END(Tile_X8Y1_N1BEG),
    .N2MID(Tile_X8Y1_N2BEG),
    .N2END(Tile_X8Y1_N2BEGb),
    .N4END(Tile_X8Y1_N4BEG),
    .NN4END(Tile_X8Y1_NN4BEG),
    .Ci(Tile_X8Y1_Co),
    .S1BEG(Tile_X8Y0_S1BEG),
    .S2BEG(Tile_X8Y0_S2BEG),
    .S2BEGb(Tile_X8Y0_S2BEGb),
    .S4BEG(Tile_X8Y0_S4BEG),
    .SS4BEG(Tile_X8Y0_SS4BEG),
    .UserCLK(Tile_X8Y1_UserCLKo),
    .UserCLKo(Tile_X8Y0_UserCLKo),
    .FrameData(Tile_X7Y0_FrameData_O),
    .FrameData_O(Tile_X8Y0_FrameData_O),
    .FrameStrobe(Tile_X8Y1_FrameStrobe_O),
    .FrameStrobe_O(Tile_X8Y0_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
N_term_single Tile_X9Y0_N_term_single (
    .N1END(Tile_X9Y1_N1BEG),
    .N2MID(Tile_X9Y1_N2BEG),
    .N2END(Tile_X9Y1_N2BEGb),
    .N4END(Tile_X9Y1_N4BEG),
    .NN4END(Tile_X9Y1_NN4BEG),
    .Ci(Tile_X9Y1_Co),
    .S1BEG(Tile_X9Y0_S1BEG),
    .S2BEG(Tile_X9Y0_S2BEG),
    .S2BEGb(Tile_X9Y0_S2BEGb),
    .S4BEG(Tile_X9Y0_S4BEG),
    .SS4BEG(Tile_X9Y0_SS4BEG),
    .UserCLK(Tile_X9Y1_UserCLKo),
    .UserCLKo(Tile_X9Y0_UserCLKo),
    .FrameData(Tile_X8Y0_FrameData_O),
    .FrameData_O(Tile_X9Y0_FrameData_O),
    .FrameStrobe(Tile_X9Y1_FrameStrobe_O),
    .FrameStrobe_O(Tile_X9Y0_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
N_term_IHP_SRAM Tile_X10Y0_N_term_IHP_SRAM (
    .N1END(Tile_X10Y1_N1BEG),
    .N2MID(Tile_X10Y1_N2BEG),
    .N2END(Tile_X10Y1_N2BEGb),
    .N4END(Tile_X10Y1_N4BEG),
    .S1BEG(Tile_X10Y0_S1BEG),
    .S2BEG(Tile_X10Y0_S2BEG),
    .S2BEGb(Tile_X10Y0_S2BEGb),
    .S4BEG(Tile_X10Y0_S4BEG),
    .UserCLK(Tile_X10Y1_UserCLKo),
    .UserCLKo(Tile_X10Y0_UserCLKo),
    .FrameData(Tile_X9Y0_FrameData_O),
    .FrameData_O(Tile_X10Y0_FrameData_O),
    .FrameStrobe(Tile_X10Y1_FrameStrobe_O),
    .FrameStrobe_O(Tile_X10Y0_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
W_IO
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X0Y1_Emulate_Bitstream)
    )
`endif
    Tile_X0Y1_W_IO
    (
    .W1END(Tile_X1Y1_W1BEG),
    .W2MID(Tile_X1Y1_W2BEG),
    .W2END(Tile_X1Y1_W2BEGb),
    .WW4END(Tile_X1Y1_WW4BEG),
    .W6END(Tile_X1Y1_W6BEG),
    .E1BEG(Tile_X0Y1_E1BEG),
    .E2BEG(Tile_X0Y1_E2BEG),
    .E2BEGb(Tile_X0Y1_E2BEGb),
    .EE4BEG(Tile_X0Y1_EE4BEG),
    .E6BEG(Tile_X0Y1_E6BEG),
    .A_O_top(Tile_X0Y1_A_O_top),
    .A_I_top(Tile_X0Y1_A_I_top),
    .A_T_top(Tile_X0Y1_A_T_top),
    .B_O_top(Tile_X0Y1_B_O_top),
    .B_I_top(Tile_X0Y1_B_I_top),
    .B_T_top(Tile_X0Y1_B_T_top),
    .A_config_C_bit0(Tile_X0Y1_A_config_C_bit0),
    .A_config_C_bit1(Tile_X0Y1_A_config_C_bit1),
    .A_config_C_bit2(Tile_X0Y1_A_config_C_bit2),
    .A_config_C_bit3(Tile_X0Y1_A_config_C_bit3),
    .B_config_C_bit0(Tile_X0Y1_B_config_C_bit0),
    .B_config_C_bit1(Tile_X0Y1_B_config_C_bit1),
    .B_config_C_bit2(Tile_X0Y1_B_config_C_bit2),
    .B_config_C_bit3(Tile_X0Y1_B_config_C_bit3),
    .UserCLK(Tile_X0Y2_UserCLKo),
    .UserCLKo(Tile_X0Y1_UserCLKo),
    .FrameData(Row_Y1_FrameData),
    .FrameData_O(Tile_X0Y1_FrameData_O),
    .FrameStrobe(Tile_X0Y2_FrameStrobe_O),
    .FrameStrobe_O(Tile_X0Y1_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X1Y1_Emulate_Bitstream)
    )
`endif
    Tile_X1Y1_LUT4AB
    (
    .N1END(Tile_X1Y2_N1BEG),
    .N2MID(Tile_X1Y2_N2BEG),
    .N2END(Tile_X1Y2_N2BEGb),
    .N4END(Tile_X1Y2_N4BEG),
    .NN4END(Tile_X1Y2_NN4BEG),
    .Ci(Tile_X1Y2_Co),
    .E1END(Tile_X0Y1_E1BEG),
    .E2MID(Tile_X0Y1_E2BEG),
    .E2END(Tile_X0Y1_E2BEGb),
    .EE4END(Tile_X0Y1_EE4BEG),
    .E6END(Tile_X0Y1_E6BEG),
    .S1END(Tile_X1Y0_S1BEG),
    .S2MID(Tile_X1Y0_S2BEG),
    .S2END(Tile_X1Y0_S2BEGb),
    .S4END(Tile_X1Y0_S4BEG),
    .SS4END(Tile_X1Y0_SS4BEG),
    .W1END(Tile_X2Y1_W1BEG),
    .W2MID(Tile_X2Y1_W2BEG),
    .W2END(Tile_X2Y1_W2BEGb),
    .WW4END(Tile_X2Y1_WW4BEG),
    .W6END(Tile_X2Y1_W6BEG),
    .N1BEG(Tile_X1Y1_N1BEG),
    .N2BEG(Tile_X1Y1_N2BEG),
    .N2BEGb(Tile_X1Y1_N2BEGb),
    .N4BEG(Tile_X1Y1_N4BEG),
    .NN4BEG(Tile_X1Y1_NN4BEG),
    .E1BEG(Tile_X1Y1_E1BEG),
    .E2BEG(Tile_X1Y1_E2BEG),
    .E2BEGb(Tile_X1Y1_E2BEGb),
    .EE4BEG(Tile_X1Y1_EE4BEG),
    .E6BEG(Tile_X1Y1_E6BEG),
    .S1BEG(Tile_X1Y1_S1BEG),
    .S2BEG(Tile_X1Y1_S2BEG),
    .S2BEGb(Tile_X1Y1_S2BEGb),
    .S4BEG(Tile_X1Y1_S4BEG),
    .SS4BEG(Tile_X1Y1_SS4BEG),
    .W1BEG(Tile_X1Y1_W1BEG),
    .W2BEG(Tile_X1Y1_W2BEG),
    .W2BEGb(Tile_X1Y1_W2BEGb),
    .WW4BEG(Tile_X1Y1_WW4BEG),
    .W6BEG(Tile_X1Y1_W6BEG),
    .Co(Tile_X1Y1_Co),
    .UserCLK(Tile_X1Y2_UserCLKo),
    .UserCLKo(Tile_X1Y1_UserCLKo),
    .FrameData(Tile_X0Y1_FrameData_O),
    .FrameData_O(Tile_X1Y1_FrameData_O),
    .FrameStrobe(Tile_X1Y2_FrameStrobe_O),
    .FrameStrobe_O(Tile_X1Y1_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X2Y1_Emulate_Bitstream)
    )
`endif
    Tile_X2Y1_LUT4AB
    (
    .N1END(Tile_X2Y2_N1BEG),
    .N2MID(Tile_X2Y2_N2BEG),
    .N2END(Tile_X2Y2_N2BEGb),
    .N4END(Tile_X2Y2_N4BEG),
    .NN4END(Tile_X2Y2_NN4BEG),
    .Ci(Tile_X2Y2_Co),
    .E1END(Tile_X1Y1_E1BEG),
    .E2MID(Tile_X1Y1_E2BEG),
    .E2END(Tile_X1Y1_E2BEGb),
    .EE4END(Tile_X1Y1_EE4BEG),
    .E6END(Tile_X1Y1_E6BEG),
    .S1END(Tile_X2Y0_S1BEG),
    .S2MID(Tile_X2Y0_S2BEG),
    .S2END(Tile_X2Y0_S2BEGb),
    .S4END(Tile_X2Y0_S4BEG),
    .SS4END(Tile_X2Y0_SS4BEG),
    .W1END(Tile_X3Y1_W1BEG),
    .W2MID(Tile_X3Y1_W2BEG),
    .W2END(Tile_X3Y1_W2BEGb),
    .WW4END(Tile_X3Y1_WW4BEG),
    .W6END(Tile_X3Y1_W6BEG),
    .N1BEG(Tile_X2Y1_N1BEG),
    .N2BEG(Tile_X2Y1_N2BEG),
    .N2BEGb(Tile_X2Y1_N2BEGb),
    .N4BEG(Tile_X2Y1_N4BEG),
    .NN4BEG(Tile_X2Y1_NN4BEG),
    .E1BEG(Tile_X2Y1_E1BEG),
    .E2BEG(Tile_X2Y1_E2BEG),
    .E2BEGb(Tile_X2Y1_E2BEGb),
    .EE4BEG(Tile_X2Y1_EE4BEG),
    .E6BEG(Tile_X2Y1_E6BEG),
    .S1BEG(Tile_X2Y1_S1BEG),
    .S2BEG(Tile_X2Y1_S2BEG),
    .S2BEGb(Tile_X2Y1_S2BEGb),
    .S4BEG(Tile_X2Y1_S4BEG),
    .SS4BEG(Tile_X2Y1_SS4BEG),
    .W1BEG(Tile_X2Y1_W1BEG),
    .W2BEG(Tile_X2Y1_W2BEG),
    .W2BEGb(Tile_X2Y1_W2BEGb),
    .WW4BEG(Tile_X2Y1_WW4BEG),
    .W6BEG(Tile_X2Y1_W6BEG),
    .Co(Tile_X2Y1_Co),
    .UserCLK(Tile_X2Y2_UserCLKo),
    .UserCLKo(Tile_X2Y1_UserCLKo),
    .FrameData(Tile_X1Y1_FrameData_O),
    .FrameData_O(Tile_X2Y1_FrameData_O),
    .FrameStrobe(Tile_X2Y2_FrameStrobe_O),
    .FrameStrobe_O(Tile_X2Y1_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X3Y1_Emulate_Bitstream)
    )
`endif
    Tile_X3Y1_LUT4AB
    (
    .N1END(Tile_X3Y2_N1BEG),
    .N2MID(Tile_X3Y2_N2BEG),
    .N2END(Tile_X3Y2_N2BEGb),
    .N4END(Tile_X3Y2_N4BEG),
    .NN4END(Tile_X3Y2_NN4BEG),
    .Ci(Tile_X3Y2_Co),
    .E1END(Tile_X2Y1_E1BEG),
    .E2MID(Tile_X2Y1_E2BEG),
    .E2END(Tile_X2Y1_E2BEGb),
    .EE4END(Tile_X2Y1_EE4BEG),
    .E6END(Tile_X2Y1_E6BEG),
    .S1END(Tile_X3Y0_S1BEG),
    .S2MID(Tile_X3Y0_S2BEG),
    .S2END(Tile_X3Y0_S2BEGb),
    .S4END(Tile_X3Y0_S4BEG),
    .SS4END(Tile_X3Y0_SS4BEG),
    .W1END(Tile_X4Y1_W1BEG),
    .W2MID(Tile_X4Y1_W2BEG),
    .W2END(Tile_X4Y1_W2BEGb),
    .WW4END(Tile_X4Y1_WW4BEG),
    .W6END(Tile_X4Y1_W6BEG),
    .N1BEG(Tile_X3Y1_N1BEG),
    .N2BEG(Tile_X3Y1_N2BEG),
    .N2BEGb(Tile_X3Y1_N2BEGb),
    .N4BEG(Tile_X3Y1_N4BEG),
    .NN4BEG(Tile_X3Y1_NN4BEG),
    .E1BEG(Tile_X3Y1_E1BEG),
    .E2BEG(Tile_X3Y1_E2BEG),
    .E2BEGb(Tile_X3Y1_E2BEGb),
    .EE4BEG(Tile_X3Y1_EE4BEG),
    .E6BEG(Tile_X3Y1_E6BEG),
    .S1BEG(Tile_X3Y1_S1BEG),
    .S2BEG(Tile_X3Y1_S2BEG),
    .S2BEGb(Tile_X3Y1_S2BEGb),
    .S4BEG(Tile_X3Y1_S4BEG),
    .SS4BEG(Tile_X3Y1_SS4BEG),
    .W1BEG(Tile_X3Y1_W1BEG),
    .W2BEG(Tile_X3Y1_W2BEG),
    .W2BEGb(Tile_X3Y1_W2BEGb),
    .WW4BEG(Tile_X3Y1_WW4BEG),
    .W6BEG(Tile_X3Y1_W6BEG),
    .Co(Tile_X3Y1_Co),
    .UserCLK(Tile_X3Y2_UserCLKo),
    .UserCLKo(Tile_X3Y1_UserCLKo),
    .FrameData(Tile_X2Y1_FrameData_O),
    .FrameData_O(Tile_X3Y1_FrameData_O),
    .FrameStrobe(Tile_X3Y2_FrameStrobe_O),
    .FrameStrobe_O(Tile_X3Y1_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
RegFile
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X4Y1_Emulate_Bitstream)
    )
`endif
    Tile_X4Y1_RegFile
    (
    .N1END(Tile_X4Y2_N1BEG),
    .N2MID(Tile_X4Y2_N2BEG),
    .N2END(Tile_X4Y2_N2BEGb),
    .N4END(Tile_X4Y2_N4BEG),
    .NN4END(Tile_X4Y2_NN4BEG),
    .E1END(Tile_X3Y1_E1BEG),
    .E2MID(Tile_X3Y1_E2BEG),
    .E2END(Tile_X3Y1_E2BEGb),
    .EE4END(Tile_X3Y1_EE4BEG),
    .E6END(Tile_X3Y1_E6BEG),
    .S1END(Tile_X4Y0_S1BEG),
    .S2MID(Tile_X4Y0_S2BEG),
    .S2END(Tile_X4Y0_S2BEGb),
    .S4END(Tile_X4Y0_S4BEG),
    .SS4END(Tile_X4Y0_SS4BEG),
    .W1END(Tile_X5Y1_W1BEG),
    .W2MID(Tile_X5Y1_W2BEG),
    .W2END(Tile_X5Y1_W2BEGb),
    .WW4END(Tile_X5Y1_WW4BEG),
    .W6END(Tile_X5Y1_W6BEG),
    .N1BEG(Tile_X4Y1_N1BEG),
    .N2BEG(Tile_X4Y1_N2BEG),
    .N2BEGb(Tile_X4Y1_N2BEGb),
    .N4BEG(Tile_X4Y1_N4BEG),
    .NN4BEG(Tile_X4Y1_NN4BEG),
    .E1BEG(Tile_X4Y1_E1BEG),
    .E2BEG(Tile_X4Y1_E2BEG),
    .E2BEGb(Tile_X4Y1_E2BEGb),
    .EE4BEG(Tile_X4Y1_EE4BEG),
    .E6BEG(Tile_X4Y1_E6BEG),
    .S1BEG(Tile_X4Y1_S1BEG),
    .S2BEG(Tile_X4Y1_S2BEG),
    .S2BEGb(Tile_X4Y1_S2BEGb),
    .S4BEG(Tile_X4Y1_S4BEG),
    .SS4BEG(Tile_X4Y1_SS4BEG),
    .W1BEG(Tile_X4Y1_W1BEG),
    .W2BEG(Tile_X4Y1_W2BEG),
    .W2BEGb(Tile_X4Y1_W2BEGb),
    .WW4BEG(Tile_X4Y1_WW4BEG),
    .W6BEG(Tile_X4Y1_W6BEG),
    .UserCLK(Tile_X4Y2_UserCLKo),
    .UserCLKo(Tile_X4Y1_UserCLKo),
    .FrameData(Tile_X3Y1_FrameData_O),
    .FrameData_O(Tile_X4Y1_FrameData_O),
    .FrameStrobe(Tile_X4Y2_FrameStrobe_O),
    .FrameStrobe_O(Tile_X4Y1_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X5Y1_Emulate_Bitstream)
    )
`endif
    Tile_X5Y1_LUT4AB
    (
    .N1END(Tile_X5Y2_N1BEG),
    .N2MID(Tile_X5Y2_N2BEG),
    .N2END(Tile_X5Y2_N2BEGb),
    .N4END(Tile_X5Y2_N4BEG),
    .NN4END(Tile_X5Y2_NN4BEG),
    .Ci(Tile_X5Y2_Co),
    .E1END(Tile_X4Y1_E1BEG),
    .E2MID(Tile_X4Y1_E2BEG),
    .E2END(Tile_X4Y1_E2BEGb),
    .EE4END(Tile_X4Y1_EE4BEG),
    .E6END(Tile_X4Y1_E6BEG),
    .S1END(Tile_X5Y0_S1BEG),
    .S2MID(Tile_X5Y0_S2BEG),
    .S2END(Tile_X5Y0_S2BEGb),
    .S4END(Tile_X5Y0_S4BEG),
    .SS4END(Tile_X5Y0_SS4BEG),
    .W1END(Tile_X6Y1_W1BEG),
    .W2MID(Tile_X6Y1_W2BEG),
    .W2END(Tile_X6Y1_W2BEGb),
    .WW4END(Tile_X6Y1_WW4BEG),
    .W6END(Tile_X6Y1_W6BEG),
    .N1BEG(Tile_X5Y1_N1BEG),
    .N2BEG(Tile_X5Y1_N2BEG),
    .N2BEGb(Tile_X5Y1_N2BEGb),
    .N4BEG(Tile_X5Y1_N4BEG),
    .NN4BEG(Tile_X5Y1_NN4BEG),
    .E1BEG(Tile_X5Y1_E1BEG),
    .E2BEG(Tile_X5Y1_E2BEG),
    .E2BEGb(Tile_X5Y1_E2BEGb),
    .EE4BEG(Tile_X5Y1_EE4BEG),
    .E6BEG(Tile_X5Y1_E6BEG),
    .S1BEG(Tile_X5Y1_S1BEG),
    .S2BEG(Tile_X5Y1_S2BEG),
    .S2BEGb(Tile_X5Y1_S2BEGb),
    .S4BEG(Tile_X5Y1_S4BEG),
    .SS4BEG(Tile_X5Y1_SS4BEG),
    .W1BEG(Tile_X5Y1_W1BEG),
    .W2BEG(Tile_X5Y1_W2BEG),
    .W2BEGb(Tile_X5Y1_W2BEGb),
    .WW4BEG(Tile_X5Y1_WW4BEG),
    .W6BEG(Tile_X5Y1_W6BEG),
    .Co(Tile_X5Y1_Co),
    .UserCLK(Tile_X5Y2_UserCLKo),
    .UserCLKo(Tile_X5Y1_UserCLKo),
    .FrameData(Tile_X4Y1_FrameData_O),
    .FrameData_O(Tile_X5Y1_FrameData_O),
    .FrameStrobe(Tile_X5Y2_FrameStrobe_O),
    .FrameStrobe_O(Tile_X5Y1_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X6Y1_Emulate_Bitstream)
    )
`endif
    Tile_X6Y1_LUT4AB
    (
    .N1END(Tile_X6Y2_N1BEG),
    .N2MID(Tile_X6Y2_N2BEG),
    .N2END(Tile_X6Y2_N2BEGb),
    .N4END(Tile_X6Y2_N4BEG),
    .NN4END(Tile_X6Y2_NN4BEG),
    .Ci(Tile_X6Y2_Co),
    .E1END(Tile_X5Y1_E1BEG),
    .E2MID(Tile_X5Y1_E2BEG),
    .E2END(Tile_X5Y1_E2BEGb),
    .EE4END(Tile_X5Y1_EE4BEG),
    .E6END(Tile_X5Y1_E6BEG),
    .S1END(Tile_X6Y0_S1BEG),
    .S2MID(Tile_X6Y0_S2BEG),
    .S2END(Tile_X6Y0_S2BEGb),
    .S4END(Tile_X6Y0_S4BEG),
    .SS4END(Tile_X6Y0_SS4BEG),
    .W1END(Tile_X7Y1_W1BEG),
    .W2MID(Tile_X7Y1_W2BEG),
    .W2END(Tile_X7Y1_W2BEGb),
    .WW4END(Tile_X7Y1_WW4BEG),
    .W6END(Tile_X7Y1_W6BEG),
    .N1BEG(Tile_X6Y1_N1BEG),
    .N2BEG(Tile_X6Y1_N2BEG),
    .N2BEGb(Tile_X6Y1_N2BEGb),
    .N4BEG(Tile_X6Y1_N4BEG),
    .NN4BEG(Tile_X6Y1_NN4BEG),
    .E1BEG(Tile_X6Y1_E1BEG),
    .E2BEG(Tile_X6Y1_E2BEG),
    .E2BEGb(Tile_X6Y1_E2BEGb),
    .EE4BEG(Tile_X6Y1_EE4BEG),
    .E6BEG(Tile_X6Y1_E6BEG),
    .S1BEG(Tile_X6Y1_S1BEG),
    .S2BEG(Tile_X6Y1_S2BEG),
    .S2BEGb(Tile_X6Y1_S2BEGb),
    .S4BEG(Tile_X6Y1_S4BEG),
    .SS4BEG(Tile_X6Y1_SS4BEG),
    .W1BEG(Tile_X6Y1_W1BEG),
    .W2BEG(Tile_X6Y1_W2BEG),
    .W2BEGb(Tile_X6Y1_W2BEGb),
    .WW4BEG(Tile_X6Y1_WW4BEG),
    .W6BEG(Tile_X6Y1_W6BEG),
    .Co(Tile_X6Y1_Co),
    .UserCLK(Tile_X6Y2_UserCLKo),
    .UserCLKo(Tile_X6Y1_UserCLKo),
    .FrameData(Tile_X5Y1_FrameData_O),
    .FrameData_O(Tile_X6Y1_FrameData_O),
    .FrameStrobe(Tile_X6Y2_FrameStrobe_O),
    .FrameStrobe_O(Tile_X6Y1_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
DSP
`ifdef EMULATION
    #(
    .Tile_X0Y0_Emulate_Bitstream(`Tile_X7Y1_Emulate_Bitstream),
    .Tile_X0Y1_Emulate_Bitstream(`Tile_X7Y2_Emulate_Bitstream)
    )
`endif
    Tile_X7Y1_DSP
    (
    .Tile_X0Y0_E1END(Tile_X6Y1_E1BEG),
    .Tile_X0Y0_E2MID(Tile_X6Y1_E2BEG),
    .Tile_X0Y0_E2END(Tile_X6Y1_E2BEGb),
    .Tile_X0Y0_EE4END(Tile_X6Y1_EE4BEG),
    .Tile_X0Y0_E6END(Tile_X6Y1_E6BEG),
    .Tile_X0Y0_S1END(Tile_X7Y0_S1BEG),
    .Tile_X0Y0_S2MID(Tile_X7Y0_S2BEG),
    .Tile_X0Y0_S2END(Tile_X7Y0_S2BEGb),
    .Tile_X0Y0_S4END(Tile_X7Y0_S4BEG),
    .Tile_X0Y0_SS4END(Tile_X7Y0_SS4BEG),
    .Tile_X0Y0_W1END(Tile_X8Y1_W1BEG),
    .Tile_X0Y0_W2MID(Tile_X8Y1_W2BEG),
    .Tile_X0Y0_W2END(Tile_X8Y1_W2BEGb),
    .Tile_X0Y0_WW4END(Tile_X8Y1_WW4BEG),
    .Tile_X0Y0_W6END(Tile_X8Y1_W6BEG),
    .Tile_X0Y1_N1END(Tile_X7Y3_N1BEG),
    .Tile_X0Y1_N2MID(Tile_X7Y3_N2BEG),
    .Tile_X0Y1_N2END(Tile_X7Y3_N2BEGb),
    .Tile_X0Y1_N4END(Tile_X7Y3_N4BEG),
    .Tile_X0Y1_NN4END(Tile_X7Y3_NN4BEG),
    .Tile_X0Y1_E1END(Tile_X6Y2_E1BEG),
    .Tile_X0Y1_E2MID(Tile_X6Y2_E2BEG),
    .Tile_X0Y1_E2END(Tile_X6Y2_E2BEGb),
    .Tile_X0Y1_EE4END(Tile_X6Y2_EE4BEG),
    .Tile_X0Y1_E6END(Tile_X6Y2_E6BEG),
    .Tile_X0Y1_W1END(Tile_X8Y2_W1BEG),
    .Tile_X0Y1_W2MID(Tile_X8Y2_W2BEG),
    .Tile_X0Y1_W2END(Tile_X8Y2_W2BEGb),
    .Tile_X0Y1_WW4END(Tile_X8Y2_WW4BEG),
    .Tile_X0Y1_W6END(Tile_X8Y2_W6BEG),
    .Tile_X0Y0_N1BEG(Tile_X7Y1_N1BEG),
    .Tile_X0Y0_N2BEG(Tile_X7Y1_N2BEG),
    .Tile_X0Y0_N2BEGb(Tile_X7Y1_N2BEGb),
    .Tile_X0Y0_N4BEG(Tile_X7Y1_N4BEG),
    .Tile_X0Y0_NN4BEG(Tile_X7Y1_NN4BEG),
    .Tile_X0Y0_E1BEG(Tile_X7Y1_E1BEG),
    .Tile_X0Y0_E2BEG(Tile_X7Y1_E2BEG),
    .Tile_X0Y0_E2BEGb(Tile_X7Y1_E2BEGb),
    .Tile_X0Y0_EE4BEG(Tile_X7Y1_EE4BEG),
    .Tile_X0Y0_E6BEG(Tile_X7Y1_E6BEG),
    .Tile_X0Y0_W1BEG(Tile_X7Y1_W1BEG),
    .Tile_X0Y0_W2BEG(Tile_X7Y1_W2BEG),
    .Tile_X0Y0_W2BEGb(Tile_X7Y1_W2BEGb),
    .Tile_X0Y0_WW4BEG(Tile_X7Y1_WW4BEG),
    .Tile_X0Y0_W6BEG(Tile_X7Y1_W6BEG),
    .Tile_X0Y1_E1BEG(Tile_X7Y2_E1BEG),
    .Tile_X0Y1_E2BEG(Tile_X7Y2_E2BEG),
    .Tile_X0Y1_E2BEGb(Tile_X7Y2_E2BEGb),
    .Tile_X0Y1_EE4BEG(Tile_X7Y2_EE4BEG),
    .Tile_X0Y1_E6BEG(Tile_X7Y2_E6BEG),
    .Tile_X0Y1_S1BEG(Tile_X7Y2_S1BEG),
    .Tile_X0Y1_S2BEG(Tile_X7Y2_S2BEG),
    .Tile_X0Y1_S2BEGb(Tile_X7Y2_S2BEGb),
    .Tile_X0Y1_S4BEG(Tile_X7Y2_S4BEG),
    .Tile_X0Y1_SS4BEG(Tile_X7Y2_SS4BEG),
    .Tile_X0Y1_W1BEG(Tile_X7Y2_W1BEG),
    .Tile_X0Y1_W2BEG(Tile_X7Y2_W2BEG),
    .Tile_X0Y1_W2BEGb(Tile_X7Y2_W2BEGb),
    .Tile_X0Y1_WW4BEG(Tile_X7Y2_WW4BEG),
    .Tile_X0Y1_W6BEG(Tile_X7Y2_W6BEG),
    .Tile_X0Y0_UserCLKo(Tile_X7Y1_UserCLKo),
    .Tile_X0Y1_UserCLK(Tile_X7Y3_UserCLKo),
    .Tile_X0Y0_FrameData(Tile_X6Y1_FrameData_O),
    .Tile_X0Y0_FrameData_O(Tile_X7Y1_FrameData_O),
    .Tile_X0Y0_FrameStrobe_O(Tile_X7Y1_FrameStrobe_O),
    .Tile_X0Y1_FrameData(Tile_X6Y2_FrameData_O),
    .Tile_X0Y1_FrameData_O(Tile_X7Y2_FrameData_O),
    .Tile_X0Y1_FrameStrobe(Tile_X7Y3_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X8Y1_Emulate_Bitstream)
    )
`endif
    Tile_X8Y1_LUT4AB
    (
    .N1END(Tile_X8Y2_N1BEG),
    .N2MID(Tile_X8Y2_N2BEG),
    .N2END(Tile_X8Y2_N2BEGb),
    .N4END(Tile_X8Y2_N4BEG),
    .NN4END(Tile_X8Y2_NN4BEG),
    .Ci(Tile_X8Y2_Co),
    .E1END(Tile_X7Y1_E1BEG),
    .E2MID(Tile_X7Y1_E2BEG),
    .E2END(Tile_X7Y1_E2BEGb),
    .EE4END(Tile_X7Y1_EE4BEG),
    .E6END(Tile_X7Y1_E6BEG),
    .S1END(Tile_X8Y0_S1BEG),
    .S2MID(Tile_X8Y0_S2BEG),
    .S2END(Tile_X8Y0_S2BEGb),
    .S4END(Tile_X8Y0_S4BEG),
    .SS4END(Tile_X8Y0_SS4BEG),
    .W1END(Tile_X9Y1_W1BEG),
    .W2MID(Tile_X9Y1_W2BEG),
    .W2END(Tile_X9Y1_W2BEGb),
    .WW4END(Tile_X9Y1_WW4BEG),
    .W6END(Tile_X9Y1_W6BEG),
    .N1BEG(Tile_X8Y1_N1BEG),
    .N2BEG(Tile_X8Y1_N2BEG),
    .N2BEGb(Tile_X8Y1_N2BEGb),
    .N4BEG(Tile_X8Y1_N4BEG),
    .NN4BEG(Tile_X8Y1_NN4BEG),
    .E1BEG(Tile_X8Y1_E1BEG),
    .E2BEG(Tile_X8Y1_E2BEG),
    .E2BEGb(Tile_X8Y1_E2BEGb),
    .EE4BEG(Tile_X8Y1_EE4BEG),
    .E6BEG(Tile_X8Y1_E6BEG),
    .S1BEG(Tile_X8Y1_S1BEG),
    .S2BEG(Tile_X8Y1_S2BEG),
    .S2BEGb(Tile_X8Y1_S2BEGb),
    .S4BEG(Tile_X8Y1_S4BEG),
    .SS4BEG(Tile_X8Y1_SS4BEG),
    .W1BEG(Tile_X8Y1_W1BEG),
    .W2BEG(Tile_X8Y1_W2BEG),
    .W2BEGb(Tile_X8Y1_W2BEGb),
    .WW4BEG(Tile_X8Y1_WW4BEG),
    .W6BEG(Tile_X8Y1_W6BEG),
    .Co(Tile_X8Y1_Co),
    .UserCLK(Tile_X8Y2_UserCLKo),
    .UserCLKo(Tile_X8Y1_UserCLKo),
    .FrameData(Tile_X7Y1_FrameData_O),
    .FrameData_O(Tile_X8Y1_FrameData_O),
    .FrameStrobe(Tile_X8Y2_FrameStrobe_O),
    .FrameStrobe_O(Tile_X8Y1_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X9Y1_Emulate_Bitstream)
    )
`endif
    Tile_X9Y1_LUT4AB
    (
    .N1END(Tile_X9Y2_N1BEG),
    .N2MID(Tile_X9Y2_N2BEG),
    .N2END(Tile_X9Y2_N2BEGb),
    .N4END(Tile_X9Y2_N4BEG),
    .NN4END(Tile_X9Y2_NN4BEG),
    .Ci(Tile_X9Y2_Co),
    .E1END(Tile_X8Y1_E1BEG),
    .E2MID(Tile_X8Y1_E2BEG),
    .E2END(Tile_X8Y1_E2BEGb),
    .EE4END(Tile_X8Y1_EE4BEG),
    .E6END(Tile_X8Y1_E6BEG),
    .S1END(Tile_X9Y0_S1BEG),
    .S2MID(Tile_X9Y0_S2BEG),
    .S2END(Tile_X9Y0_S2BEGb),
    .S4END(Tile_X9Y0_S4BEG),
    .SS4END(Tile_X9Y0_SS4BEG),
    .W1END(Tile_X10Y1_W1BEG),
    .W2MID(Tile_X10Y1_W2BEG),
    .W2END(Tile_X10Y1_W2BEGb),
    .WW4END(Tile_X10Y1_WW4BEG),
    .W6END(Tile_X10Y1_W6BEG),
    .N1BEG(Tile_X9Y1_N1BEG),
    .N2BEG(Tile_X9Y1_N2BEG),
    .N2BEGb(Tile_X9Y1_N2BEGb),
    .N4BEG(Tile_X9Y1_N4BEG),
    .NN4BEG(Tile_X9Y1_NN4BEG),
    .E1BEG(Tile_X9Y1_E1BEG),
    .E2BEG(Tile_X9Y1_E2BEG),
    .E2BEGb(Tile_X9Y1_E2BEGb),
    .EE4BEG(Tile_X9Y1_EE4BEG),
    .E6BEG(Tile_X9Y1_E6BEG),
    .S1BEG(Tile_X9Y1_S1BEG),
    .S2BEG(Tile_X9Y1_S2BEG),
    .S2BEGb(Tile_X9Y1_S2BEGb),
    .S4BEG(Tile_X9Y1_S4BEG),
    .SS4BEG(Tile_X9Y1_SS4BEG),
    .W1BEG(Tile_X9Y1_W1BEG),
    .W2BEG(Tile_X9Y1_W2BEG),
    .W2BEGb(Tile_X9Y1_W2BEGb),
    .WW4BEG(Tile_X9Y1_WW4BEG),
    .W6BEG(Tile_X9Y1_W6BEG),
    .Co(Tile_X9Y1_Co),
    .UserCLK(Tile_X9Y2_UserCLKo),
    .UserCLKo(Tile_X9Y1_UserCLKo),
    .FrameData(Tile_X8Y1_FrameData_O),
    .FrameData_O(Tile_X9Y1_FrameData_O),
    .FrameStrobe(Tile_X9Y2_FrameStrobe_O),
    .FrameStrobe_O(Tile_X9Y1_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
IHP_SRAM
`ifdef EMULATION
    #(
    .Tile_X0Y0_Emulate_Bitstream(`Tile_X10Y1_Emulate_Bitstream),
    .Tile_X0Y1_Emulate_Bitstream(`Tile_X10Y2_Emulate_Bitstream)
    )
`endif
    Tile_X10Y1_IHP_SRAM
    (
    .Tile_X0Y0_E1END(Tile_X9Y1_E1BEG),
    .Tile_X0Y0_E2MID(Tile_X9Y1_E2BEG),
    .Tile_X0Y0_E2END(Tile_X9Y1_E2BEGb),
    .Tile_X0Y0_EE4END(Tile_X9Y1_EE4BEG),
    .Tile_X0Y0_E6END(Tile_X9Y1_E6BEG),
    .Tile_X0Y0_S1END(Tile_X10Y0_S1BEG),
    .Tile_X0Y0_S2MID(Tile_X10Y0_S2BEG),
    .Tile_X0Y0_S2END(Tile_X10Y0_S2BEGb),
    .Tile_X0Y0_S4END(Tile_X10Y0_S4BEG),
    .Tile_X0Y1_N1END(Tile_X10Y3_N1BEG),
    .Tile_X0Y1_N2MID(Tile_X10Y3_N2BEG),
    .Tile_X0Y1_N2END(Tile_X10Y3_N2BEGb),
    .Tile_X0Y1_N4END(Tile_X10Y3_N4BEG),
    .Tile_X0Y1_E1END(Tile_X9Y2_E1BEG),
    .Tile_X0Y1_E2MID(Tile_X9Y2_E2BEG),
    .Tile_X0Y1_E2END(Tile_X9Y2_E2BEGb),
    .Tile_X0Y1_EE4END(Tile_X9Y2_EE4BEG),
    .Tile_X0Y1_E6END(Tile_X9Y2_E6BEG),
    .Tile_X0Y0_N1BEG(Tile_X10Y1_N1BEG),
    .Tile_X0Y0_N2BEG(Tile_X10Y1_N2BEG),
    .Tile_X0Y0_N2BEGb(Tile_X10Y1_N2BEGb),
    .Tile_X0Y0_N4BEG(Tile_X10Y1_N4BEG),
    .Tile_X0Y0_W1BEG(Tile_X10Y1_W1BEG),
    .Tile_X0Y0_W2BEG(Tile_X10Y1_W2BEG),
    .Tile_X0Y0_W2BEGb(Tile_X10Y1_W2BEGb),
    .Tile_X0Y0_WW4BEG(Tile_X10Y1_WW4BEG),
    .Tile_X0Y0_W6BEG(Tile_X10Y1_W6BEG),
    .Tile_X0Y1_S1BEG(Tile_X10Y2_S1BEG),
    .Tile_X0Y1_S2BEG(Tile_X10Y2_S2BEG),
    .Tile_X0Y1_S2BEGb(Tile_X10Y2_S2BEGb),
    .Tile_X0Y1_S4BEG(Tile_X10Y2_S4BEG),
    .Tile_X0Y1_W1BEG(Tile_X10Y2_W1BEG),
    .Tile_X0Y1_W2BEG(Tile_X10Y2_W2BEG),
    .Tile_X0Y1_W2BEGb(Tile_X10Y2_W2BEGb),
    .Tile_X0Y1_WW4BEG(Tile_X10Y2_WW4BEG),
    .Tile_X0Y1_W6BEG(Tile_X10Y2_W6BEG),
    .CONFIGURED_top(Tile_X10Y2_CONFIGURED_top),
    .DOUT_SRAM0(Tile_X10Y2_DOUT_SRAM0),
    .DOUT_SRAM1(Tile_X10Y2_DOUT_SRAM1),
    .DOUT_SRAM2(Tile_X10Y2_DOUT_SRAM2),
    .DOUT_SRAM3(Tile_X10Y2_DOUT_SRAM3),
    .DOUT_SRAM4(Tile_X10Y2_DOUT_SRAM4),
    .DOUT_SRAM5(Tile_X10Y2_DOUT_SRAM5),
    .DOUT_SRAM6(Tile_X10Y2_DOUT_SRAM6),
    .DOUT_SRAM7(Tile_X10Y2_DOUT_SRAM7),
    .DOUT_SRAM8(Tile_X10Y2_DOUT_SRAM8),
    .DOUT_SRAM9(Tile_X10Y2_DOUT_SRAM9),
    .DOUT_SRAM10(Tile_X10Y2_DOUT_SRAM10),
    .DOUT_SRAM11(Tile_X10Y2_DOUT_SRAM11),
    .DOUT_SRAM12(Tile_X10Y2_DOUT_SRAM12),
    .DOUT_SRAM13(Tile_X10Y2_DOUT_SRAM13),
    .DOUT_SRAM14(Tile_X10Y2_DOUT_SRAM14),
    .DOUT_SRAM15(Tile_X10Y2_DOUT_SRAM15),
    .DOUT_SRAM16(Tile_X10Y2_DOUT_SRAM16),
    .DOUT_SRAM17(Tile_X10Y2_DOUT_SRAM17),
    .DOUT_SRAM18(Tile_X10Y2_DOUT_SRAM18),
    .DOUT_SRAM19(Tile_X10Y2_DOUT_SRAM19),
    .DOUT_SRAM20(Tile_X10Y2_DOUT_SRAM20),
    .DOUT_SRAM21(Tile_X10Y2_DOUT_SRAM21),
    .DOUT_SRAM22(Tile_X10Y2_DOUT_SRAM22),
    .DOUT_SRAM23(Tile_X10Y2_DOUT_SRAM23),
    .DOUT_SRAM24(Tile_X10Y2_DOUT_SRAM24),
    .DOUT_SRAM25(Tile_X10Y2_DOUT_SRAM25),
    .DOUT_SRAM26(Tile_X10Y2_DOUT_SRAM26),
    .DOUT_SRAM27(Tile_X10Y2_DOUT_SRAM27),
    .DOUT_SRAM28(Tile_X10Y2_DOUT_SRAM28),
    .DOUT_SRAM29(Tile_X10Y2_DOUT_SRAM29),
    .DOUT_SRAM30(Tile_X10Y2_DOUT_SRAM30),
    .DOUT_SRAM31(Tile_X10Y2_DOUT_SRAM31),
    .ADDR_SRAM0(Tile_X10Y2_ADDR_SRAM0),
    .ADDR_SRAM1(Tile_X10Y2_ADDR_SRAM1),
    .ADDR_SRAM2(Tile_X10Y2_ADDR_SRAM2),
    .ADDR_SRAM3(Tile_X10Y2_ADDR_SRAM3),
    .ADDR_SRAM4(Tile_X10Y2_ADDR_SRAM4),
    .ADDR_SRAM5(Tile_X10Y2_ADDR_SRAM5),
    .ADDR_SRAM6(Tile_X10Y2_ADDR_SRAM6),
    .ADDR_SRAM7(Tile_X10Y2_ADDR_SRAM7),
    .ADDR_SRAM8(Tile_X10Y2_ADDR_SRAM8),
    .ADDR_SRAM9(Tile_X10Y2_ADDR_SRAM9),
    .BM_SRAM0(Tile_X10Y2_BM_SRAM0),
    .BM_SRAM1(Tile_X10Y2_BM_SRAM1),
    .BM_SRAM2(Tile_X10Y2_BM_SRAM2),
    .BM_SRAM3(Tile_X10Y2_BM_SRAM3),
    .BM_SRAM4(Tile_X10Y2_BM_SRAM4),
    .BM_SRAM5(Tile_X10Y2_BM_SRAM5),
    .BM_SRAM6(Tile_X10Y2_BM_SRAM6),
    .BM_SRAM7(Tile_X10Y2_BM_SRAM7),
    .BM_SRAM8(Tile_X10Y2_BM_SRAM8),
    .BM_SRAM9(Tile_X10Y2_BM_SRAM9),
    .BM_SRAM10(Tile_X10Y2_BM_SRAM10),
    .BM_SRAM11(Tile_X10Y2_BM_SRAM11),
    .BM_SRAM12(Tile_X10Y2_BM_SRAM12),
    .BM_SRAM13(Tile_X10Y2_BM_SRAM13),
    .BM_SRAM14(Tile_X10Y2_BM_SRAM14),
    .BM_SRAM15(Tile_X10Y2_BM_SRAM15),
    .BM_SRAM16(Tile_X10Y2_BM_SRAM16),
    .BM_SRAM17(Tile_X10Y2_BM_SRAM17),
    .BM_SRAM18(Tile_X10Y2_BM_SRAM18),
    .BM_SRAM19(Tile_X10Y2_BM_SRAM19),
    .BM_SRAM20(Tile_X10Y2_BM_SRAM20),
    .BM_SRAM21(Tile_X10Y2_BM_SRAM21),
    .BM_SRAM22(Tile_X10Y2_BM_SRAM22),
    .BM_SRAM23(Tile_X10Y2_BM_SRAM23),
    .BM_SRAM24(Tile_X10Y2_BM_SRAM24),
    .BM_SRAM25(Tile_X10Y2_BM_SRAM25),
    .BM_SRAM26(Tile_X10Y2_BM_SRAM26),
    .BM_SRAM27(Tile_X10Y2_BM_SRAM27),
    .BM_SRAM28(Tile_X10Y2_BM_SRAM28),
    .BM_SRAM29(Tile_X10Y2_BM_SRAM29),
    .BM_SRAM30(Tile_X10Y2_BM_SRAM30),
    .BM_SRAM31(Tile_X10Y2_BM_SRAM31),
    .CLK_SRAM(Tile_X10Y2_CLK_SRAM),
    .DIN_SRAM0(Tile_X10Y2_DIN_SRAM0),
    .DIN_SRAM1(Tile_X10Y2_DIN_SRAM1),
    .DIN_SRAM2(Tile_X10Y2_DIN_SRAM2),
    .DIN_SRAM3(Tile_X10Y2_DIN_SRAM3),
    .DIN_SRAM4(Tile_X10Y2_DIN_SRAM4),
    .DIN_SRAM5(Tile_X10Y2_DIN_SRAM5),
    .DIN_SRAM6(Tile_X10Y2_DIN_SRAM6),
    .DIN_SRAM7(Tile_X10Y2_DIN_SRAM7),
    .DIN_SRAM8(Tile_X10Y2_DIN_SRAM8),
    .DIN_SRAM9(Tile_X10Y2_DIN_SRAM9),
    .DIN_SRAM10(Tile_X10Y2_DIN_SRAM10),
    .DIN_SRAM11(Tile_X10Y2_DIN_SRAM11),
    .DIN_SRAM12(Tile_X10Y2_DIN_SRAM12),
    .DIN_SRAM13(Tile_X10Y2_DIN_SRAM13),
    .DIN_SRAM14(Tile_X10Y2_DIN_SRAM14),
    .DIN_SRAM15(Tile_X10Y2_DIN_SRAM15),
    .DIN_SRAM16(Tile_X10Y2_DIN_SRAM16),
    .DIN_SRAM17(Tile_X10Y2_DIN_SRAM17),
    .DIN_SRAM18(Tile_X10Y2_DIN_SRAM18),
    .DIN_SRAM19(Tile_X10Y2_DIN_SRAM19),
    .DIN_SRAM20(Tile_X10Y2_DIN_SRAM20),
    .DIN_SRAM21(Tile_X10Y2_DIN_SRAM21),
    .DIN_SRAM22(Tile_X10Y2_DIN_SRAM22),
    .DIN_SRAM23(Tile_X10Y2_DIN_SRAM23),
    .DIN_SRAM24(Tile_X10Y2_DIN_SRAM24),
    .DIN_SRAM25(Tile_X10Y2_DIN_SRAM25),
    .DIN_SRAM26(Tile_X10Y2_DIN_SRAM26),
    .DIN_SRAM27(Tile_X10Y2_DIN_SRAM27),
    .DIN_SRAM28(Tile_X10Y2_DIN_SRAM28),
    .DIN_SRAM29(Tile_X10Y2_DIN_SRAM29),
    .DIN_SRAM30(Tile_X10Y2_DIN_SRAM30),
    .DIN_SRAM31(Tile_X10Y2_DIN_SRAM31),
    .MEN_SRAM(Tile_X10Y2_MEN_SRAM),
    .REN_SRAM(Tile_X10Y2_REN_SRAM),
    .TIE_HIGH_SRAM(Tile_X10Y2_TIE_HIGH_SRAM),
    .TIE_LOW_SRAM(Tile_X10Y2_TIE_LOW_SRAM),
    .WEN_SRAM(Tile_X10Y2_WEN_SRAM),
    .Tile_X0Y0_UserCLKo(Tile_X10Y1_UserCLKo),
    .Tile_X0Y1_UserCLK(Tile_X10Y3_UserCLKo),
    .Tile_X0Y0_FrameData(Tile_X9Y1_FrameData_O),
    .Tile_X0Y0_FrameData_O(Tile_X10Y1_FrameData_O),
    .Tile_X0Y0_FrameStrobe_O(Tile_X10Y1_FrameStrobe_O),
    .Tile_X0Y1_FrameData(Tile_X9Y2_FrameData_O),
    .Tile_X0Y1_FrameData_O(Tile_X10Y2_FrameData_O),
    .Tile_X0Y1_FrameStrobe(Tile_X10Y3_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
W_IO
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X0Y2_Emulate_Bitstream)
    )
`endif
    Tile_X0Y2_W_IO
    (
    .W1END(Tile_X1Y2_W1BEG),
    .W2MID(Tile_X1Y2_W2BEG),
    .W2END(Tile_X1Y2_W2BEGb),
    .WW4END(Tile_X1Y2_WW4BEG),
    .W6END(Tile_X1Y2_W6BEG),
    .E1BEG(Tile_X0Y2_E1BEG),
    .E2BEG(Tile_X0Y2_E2BEG),
    .E2BEGb(Tile_X0Y2_E2BEGb),
    .EE4BEG(Tile_X0Y2_EE4BEG),
    .E6BEG(Tile_X0Y2_E6BEG),
    .A_O_top(Tile_X0Y2_A_O_top),
    .A_I_top(Tile_X0Y2_A_I_top),
    .A_T_top(Tile_X0Y2_A_T_top),
    .B_O_top(Tile_X0Y2_B_O_top),
    .B_I_top(Tile_X0Y2_B_I_top),
    .B_T_top(Tile_X0Y2_B_T_top),
    .A_config_C_bit0(Tile_X0Y2_A_config_C_bit0),
    .A_config_C_bit1(Tile_X0Y2_A_config_C_bit1),
    .A_config_C_bit2(Tile_X0Y2_A_config_C_bit2),
    .A_config_C_bit3(Tile_X0Y2_A_config_C_bit3),
    .B_config_C_bit0(Tile_X0Y2_B_config_C_bit0),
    .B_config_C_bit1(Tile_X0Y2_B_config_C_bit1),
    .B_config_C_bit2(Tile_X0Y2_B_config_C_bit2),
    .B_config_C_bit3(Tile_X0Y2_B_config_C_bit3),
    .UserCLK(Tile_X0Y3_UserCLKo),
    .UserCLKo(Tile_X0Y2_UserCLKo),
    .FrameData(Row_Y2_FrameData),
    .FrameData_O(Tile_X0Y2_FrameData_O),
    .FrameStrobe(Tile_X0Y3_FrameStrobe_O),
    .FrameStrobe_O(Tile_X0Y2_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X1Y2_Emulate_Bitstream)
    )
`endif
    Tile_X1Y2_LUT4AB
    (
    .N1END(Tile_X1Y3_N1BEG),
    .N2MID(Tile_X1Y3_N2BEG),
    .N2END(Tile_X1Y3_N2BEGb),
    .N4END(Tile_X1Y3_N4BEG),
    .NN4END(Tile_X1Y3_NN4BEG),
    .Ci(Tile_X1Y3_Co),
    .E1END(Tile_X0Y2_E1BEG),
    .E2MID(Tile_X0Y2_E2BEG),
    .E2END(Tile_X0Y2_E2BEGb),
    .EE4END(Tile_X0Y2_EE4BEG),
    .E6END(Tile_X0Y2_E6BEG),
    .S1END(Tile_X1Y1_S1BEG),
    .S2MID(Tile_X1Y1_S2BEG),
    .S2END(Tile_X1Y1_S2BEGb),
    .S4END(Tile_X1Y1_S4BEG),
    .SS4END(Tile_X1Y1_SS4BEG),
    .W1END(Tile_X2Y2_W1BEG),
    .W2MID(Tile_X2Y2_W2BEG),
    .W2END(Tile_X2Y2_W2BEGb),
    .WW4END(Tile_X2Y2_WW4BEG),
    .W6END(Tile_X2Y2_W6BEG),
    .N1BEG(Tile_X1Y2_N1BEG),
    .N2BEG(Tile_X1Y2_N2BEG),
    .N2BEGb(Tile_X1Y2_N2BEGb),
    .N4BEG(Tile_X1Y2_N4BEG),
    .NN4BEG(Tile_X1Y2_NN4BEG),
    .E1BEG(Tile_X1Y2_E1BEG),
    .E2BEG(Tile_X1Y2_E2BEG),
    .E2BEGb(Tile_X1Y2_E2BEGb),
    .EE4BEG(Tile_X1Y2_EE4BEG),
    .E6BEG(Tile_X1Y2_E6BEG),
    .S1BEG(Tile_X1Y2_S1BEG),
    .S2BEG(Tile_X1Y2_S2BEG),
    .S2BEGb(Tile_X1Y2_S2BEGb),
    .S4BEG(Tile_X1Y2_S4BEG),
    .SS4BEG(Tile_X1Y2_SS4BEG),
    .W1BEG(Tile_X1Y2_W1BEG),
    .W2BEG(Tile_X1Y2_W2BEG),
    .W2BEGb(Tile_X1Y2_W2BEGb),
    .WW4BEG(Tile_X1Y2_WW4BEG),
    .W6BEG(Tile_X1Y2_W6BEG),
    .Co(Tile_X1Y2_Co),
    .UserCLK(Tile_X1Y3_UserCLKo),
    .UserCLKo(Tile_X1Y2_UserCLKo),
    .FrameData(Tile_X0Y2_FrameData_O),
    .FrameData_O(Tile_X1Y2_FrameData_O),
    .FrameStrobe(Tile_X1Y3_FrameStrobe_O),
    .FrameStrobe_O(Tile_X1Y2_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X2Y2_Emulate_Bitstream)
    )
`endif
    Tile_X2Y2_LUT4AB
    (
    .N1END(Tile_X2Y3_N1BEG),
    .N2MID(Tile_X2Y3_N2BEG),
    .N2END(Tile_X2Y3_N2BEGb),
    .N4END(Tile_X2Y3_N4BEG),
    .NN4END(Tile_X2Y3_NN4BEG),
    .Ci(Tile_X2Y3_Co),
    .E1END(Tile_X1Y2_E1BEG),
    .E2MID(Tile_X1Y2_E2BEG),
    .E2END(Tile_X1Y2_E2BEGb),
    .EE4END(Tile_X1Y2_EE4BEG),
    .E6END(Tile_X1Y2_E6BEG),
    .S1END(Tile_X2Y1_S1BEG),
    .S2MID(Tile_X2Y1_S2BEG),
    .S2END(Tile_X2Y1_S2BEGb),
    .S4END(Tile_X2Y1_S4BEG),
    .SS4END(Tile_X2Y1_SS4BEG),
    .W1END(Tile_X3Y2_W1BEG),
    .W2MID(Tile_X3Y2_W2BEG),
    .W2END(Tile_X3Y2_W2BEGb),
    .WW4END(Tile_X3Y2_WW4BEG),
    .W6END(Tile_X3Y2_W6BEG),
    .N1BEG(Tile_X2Y2_N1BEG),
    .N2BEG(Tile_X2Y2_N2BEG),
    .N2BEGb(Tile_X2Y2_N2BEGb),
    .N4BEG(Tile_X2Y2_N4BEG),
    .NN4BEG(Tile_X2Y2_NN4BEG),
    .E1BEG(Tile_X2Y2_E1BEG),
    .E2BEG(Tile_X2Y2_E2BEG),
    .E2BEGb(Tile_X2Y2_E2BEGb),
    .EE4BEG(Tile_X2Y2_EE4BEG),
    .E6BEG(Tile_X2Y2_E6BEG),
    .S1BEG(Tile_X2Y2_S1BEG),
    .S2BEG(Tile_X2Y2_S2BEG),
    .S2BEGb(Tile_X2Y2_S2BEGb),
    .S4BEG(Tile_X2Y2_S4BEG),
    .SS4BEG(Tile_X2Y2_SS4BEG),
    .W1BEG(Tile_X2Y2_W1BEG),
    .W2BEG(Tile_X2Y2_W2BEG),
    .W2BEGb(Tile_X2Y2_W2BEGb),
    .WW4BEG(Tile_X2Y2_WW4BEG),
    .W6BEG(Tile_X2Y2_W6BEG),
    .Co(Tile_X2Y2_Co),
    .UserCLK(Tile_X2Y3_UserCLKo),
    .UserCLKo(Tile_X2Y2_UserCLKo),
    .FrameData(Tile_X1Y2_FrameData_O),
    .FrameData_O(Tile_X2Y2_FrameData_O),
    .FrameStrobe(Tile_X2Y3_FrameStrobe_O),
    .FrameStrobe_O(Tile_X2Y2_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X3Y2_Emulate_Bitstream)
    )
`endif
    Tile_X3Y2_LUT4AB
    (
    .N1END(Tile_X3Y3_N1BEG),
    .N2MID(Tile_X3Y3_N2BEG),
    .N2END(Tile_X3Y3_N2BEGb),
    .N4END(Tile_X3Y3_N4BEG),
    .NN4END(Tile_X3Y3_NN4BEG),
    .Ci(Tile_X3Y3_Co),
    .E1END(Tile_X2Y2_E1BEG),
    .E2MID(Tile_X2Y2_E2BEG),
    .E2END(Tile_X2Y2_E2BEGb),
    .EE4END(Tile_X2Y2_EE4BEG),
    .E6END(Tile_X2Y2_E6BEG),
    .S1END(Tile_X3Y1_S1BEG),
    .S2MID(Tile_X3Y1_S2BEG),
    .S2END(Tile_X3Y1_S2BEGb),
    .S4END(Tile_X3Y1_S4BEG),
    .SS4END(Tile_X3Y1_SS4BEG),
    .W1END(Tile_X4Y2_W1BEG),
    .W2MID(Tile_X4Y2_W2BEG),
    .W2END(Tile_X4Y2_W2BEGb),
    .WW4END(Tile_X4Y2_WW4BEG),
    .W6END(Tile_X4Y2_W6BEG),
    .N1BEG(Tile_X3Y2_N1BEG),
    .N2BEG(Tile_X3Y2_N2BEG),
    .N2BEGb(Tile_X3Y2_N2BEGb),
    .N4BEG(Tile_X3Y2_N4BEG),
    .NN4BEG(Tile_X3Y2_NN4BEG),
    .E1BEG(Tile_X3Y2_E1BEG),
    .E2BEG(Tile_X3Y2_E2BEG),
    .E2BEGb(Tile_X3Y2_E2BEGb),
    .EE4BEG(Tile_X3Y2_EE4BEG),
    .E6BEG(Tile_X3Y2_E6BEG),
    .S1BEG(Tile_X3Y2_S1BEG),
    .S2BEG(Tile_X3Y2_S2BEG),
    .S2BEGb(Tile_X3Y2_S2BEGb),
    .S4BEG(Tile_X3Y2_S4BEG),
    .SS4BEG(Tile_X3Y2_SS4BEG),
    .W1BEG(Tile_X3Y2_W1BEG),
    .W2BEG(Tile_X3Y2_W2BEG),
    .W2BEGb(Tile_X3Y2_W2BEGb),
    .WW4BEG(Tile_X3Y2_WW4BEG),
    .W6BEG(Tile_X3Y2_W6BEG),
    .Co(Tile_X3Y2_Co),
    .UserCLK(Tile_X3Y3_UserCLKo),
    .UserCLKo(Tile_X3Y2_UserCLKo),
    .FrameData(Tile_X2Y2_FrameData_O),
    .FrameData_O(Tile_X3Y2_FrameData_O),
    .FrameStrobe(Tile_X3Y3_FrameStrobe_O),
    .FrameStrobe_O(Tile_X3Y2_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
RegFile
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X4Y2_Emulate_Bitstream)
    )
`endif
    Tile_X4Y2_RegFile
    (
    .N1END(Tile_X4Y3_N1BEG),
    .N2MID(Tile_X4Y3_N2BEG),
    .N2END(Tile_X4Y3_N2BEGb),
    .N4END(Tile_X4Y3_N4BEG),
    .NN4END(Tile_X4Y3_NN4BEG),
    .E1END(Tile_X3Y2_E1BEG),
    .E2MID(Tile_X3Y2_E2BEG),
    .E2END(Tile_X3Y2_E2BEGb),
    .EE4END(Tile_X3Y2_EE4BEG),
    .E6END(Tile_X3Y2_E6BEG),
    .S1END(Tile_X4Y1_S1BEG),
    .S2MID(Tile_X4Y1_S2BEG),
    .S2END(Tile_X4Y1_S2BEGb),
    .S4END(Tile_X4Y1_S4BEG),
    .SS4END(Tile_X4Y1_SS4BEG),
    .W1END(Tile_X5Y2_W1BEG),
    .W2MID(Tile_X5Y2_W2BEG),
    .W2END(Tile_X5Y2_W2BEGb),
    .WW4END(Tile_X5Y2_WW4BEG),
    .W6END(Tile_X5Y2_W6BEG),
    .N1BEG(Tile_X4Y2_N1BEG),
    .N2BEG(Tile_X4Y2_N2BEG),
    .N2BEGb(Tile_X4Y2_N2BEGb),
    .N4BEG(Tile_X4Y2_N4BEG),
    .NN4BEG(Tile_X4Y2_NN4BEG),
    .E1BEG(Tile_X4Y2_E1BEG),
    .E2BEG(Tile_X4Y2_E2BEG),
    .E2BEGb(Tile_X4Y2_E2BEGb),
    .EE4BEG(Tile_X4Y2_EE4BEG),
    .E6BEG(Tile_X4Y2_E6BEG),
    .S1BEG(Tile_X4Y2_S1BEG),
    .S2BEG(Tile_X4Y2_S2BEG),
    .S2BEGb(Tile_X4Y2_S2BEGb),
    .S4BEG(Tile_X4Y2_S4BEG),
    .SS4BEG(Tile_X4Y2_SS4BEG),
    .W1BEG(Tile_X4Y2_W1BEG),
    .W2BEG(Tile_X4Y2_W2BEG),
    .W2BEGb(Tile_X4Y2_W2BEGb),
    .WW4BEG(Tile_X4Y2_WW4BEG),
    .W6BEG(Tile_X4Y2_W6BEG),
    .UserCLK(Tile_X4Y3_UserCLKo),
    .UserCLKo(Tile_X4Y2_UserCLKo),
    .FrameData(Tile_X3Y2_FrameData_O),
    .FrameData_O(Tile_X4Y2_FrameData_O),
    .FrameStrobe(Tile_X4Y3_FrameStrobe_O),
    .FrameStrobe_O(Tile_X4Y2_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X5Y2_Emulate_Bitstream)
    )
`endif
    Tile_X5Y2_LUT4AB
    (
    .N1END(Tile_X5Y3_N1BEG),
    .N2MID(Tile_X5Y3_N2BEG),
    .N2END(Tile_X5Y3_N2BEGb),
    .N4END(Tile_X5Y3_N4BEG),
    .NN4END(Tile_X5Y3_NN4BEG),
    .Ci(Tile_X5Y3_Co),
    .E1END(Tile_X4Y2_E1BEG),
    .E2MID(Tile_X4Y2_E2BEG),
    .E2END(Tile_X4Y2_E2BEGb),
    .EE4END(Tile_X4Y2_EE4BEG),
    .E6END(Tile_X4Y2_E6BEG),
    .S1END(Tile_X5Y1_S1BEG),
    .S2MID(Tile_X5Y1_S2BEG),
    .S2END(Tile_X5Y1_S2BEGb),
    .S4END(Tile_X5Y1_S4BEG),
    .SS4END(Tile_X5Y1_SS4BEG),
    .W1END(Tile_X6Y2_W1BEG),
    .W2MID(Tile_X6Y2_W2BEG),
    .W2END(Tile_X6Y2_W2BEGb),
    .WW4END(Tile_X6Y2_WW4BEG),
    .W6END(Tile_X6Y2_W6BEG),
    .N1BEG(Tile_X5Y2_N1BEG),
    .N2BEG(Tile_X5Y2_N2BEG),
    .N2BEGb(Tile_X5Y2_N2BEGb),
    .N4BEG(Tile_X5Y2_N4BEG),
    .NN4BEG(Tile_X5Y2_NN4BEG),
    .E1BEG(Tile_X5Y2_E1BEG),
    .E2BEG(Tile_X5Y2_E2BEG),
    .E2BEGb(Tile_X5Y2_E2BEGb),
    .EE4BEG(Tile_X5Y2_EE4BEG),
    .E6BEG(Tile_X5Y2_E6BEG),
    .S1BEG(Tile_X5Y2_S1BEG),
    .S2BEG(Tile_X5Y2_S2BEG),
    .S2BEGb(Tile_X5Y2_S2BEGb),
    .S4BEG(Tile_X5Y2_S4BEG),
    .SS4BEG(Tile_X5Y2_SS4BEG),
    .W1BEG(Tile_X5Y2_W1BEG),
    .W2BEG(Tile_X5Y2_W2BEG),
    .W2BEGb(Tile_X5Y2_W2BEGb),
    .WW4BEG(Tile_X5Y2_WW4BEG),
    .W6BEG(Tile_X5Y2_W6BEG),
    .Co(Tile_X5Y2_Co),
    .UserCLK(Tile_X5Y3_UserCLKo),
    .UserCLKo(Tile_X5Y2_UserCLKo),
    .FrameData(Tile_X4Y2_FrameData_O),
    .FrameData_O(Tile_X5Y2_FrameData_O),
    .FrameStrobe(Tile_X5Y3_FrameStrobe_O),
    .FrameStrobe_O(Tile_X5Y2_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X6Y2_Emulate_Bitstream)
    )
`endif
    Tile_X6Y2_LUT4AB
    (
    .N1END(Tile_X6Y3_N1BEG),
    .N2MID(Tile_X6Y3_N2BEG),
    .N2END(Tile_X6Y3_N2BEGb),
    .N4END(Tile_X6Y3_N4BEG),
    .NN4END(Tile_X6Y3_NN4BEG),
    .Ci(Tile_X6Y3_Co),
    .E1END(Tile_X5Y2_E1BEG),
    .E2MID(Tile_X5Y2_E2BEG),
    .E2END(Tile_X5Y2_E2BEGb),
    .EE4END(Tile_X5Y2_EE4BEG),
    .E6END(Tile_X5Y2_E6BEG),
    .S1END(Tile_X6Y1_S1BEG),
    .S2MID(Tile_X6Y1_S2BEG),
    .S2END(Tile_X6Y1_S2BEGb),
    .S4END(Tile_X6Y1_S4BEG),
    .SS4END(Tile_X6Y1_SS4BEG),
    .W1END(Tile_X7Y2_W1BEG),
    .W2MID(Tile_X7Y2_W2BEG),
    .W2END(Tile_X7Y2_W2BEGb),
    .WW4END(Tile_X7Y2_WW4BEG),
    .W6END(Tile_X7Y2_W6BEG),
    .N1BEG(Tile_X6Y2_N1BEG),
    .N2BEG(Tile_X6Y2_N2BEG),
    .N2BEGb(Tile_X6Y2_N2BEGb),
    .N4BEG(Tile_X6Y2_N4BEG),
    .NN4BEG(Tile_X6Y2_NN4BEG),
    .E1BEG(Tile_X6Y2_E1BEG),
    .E2BEG(Tile_X6Y2_E2BEG),
    .E2BEGb(Tile_X6Y2_E2BEGb),
    .EE4BEG(Tile_X6Y2_EE4BEG),
    .E6BEG(Tile_X6Y2_E6BEG),
    .S1BEG(Tile_X6Y2_S1BEG),
    .S2BEG(Tile_X6Y2_S2BEG),
    .S2BEGb(Tile_X6Y2_S2BEGb),
    .S4BEG(Tile_X6Y2_S4BEG),
    .SS4BEG(Tile_X6Y2_SS4BEG),
    .W1BEG(Tile_X6Y2_W1BEG),
    .W2BEG(Tile_X6Y2_W2BEG),
    .W2BEGb(Tile_X6Y2_W2BEGb),
    .WW4BEG(Tile_X6Y2_WW4BEG),
    .W6BEG(Tile_X6Y2_W6BEG),
    .Co(Tile_X6Y2_Co),
    .UserCLK(Tile_X6Y3_UserCLKo),
    .UserCLKo(Tile_X6Y2_UserCLKo),
    .FrameData(Tile_X5Y2_FrameData_O),
    .FrameData_O(Tile_X6Y2_FrameData_O),
    .FrameStrobe(Tile_X6Y3_FrameStrobe_O),
    .FrameStrobe_O(Tile_X6Y2_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X8Y2_Emulate_Bitstream)
    )
`endif
    Tile_X8Y2_LUT4AB
    (
    .N1END(Tile_X8Y3_N1BEG),
    .N2MID(Tile_X8Y3_N2BEG),
    .N2END(Tile_X8Y3_N2BEGb),
    .N4END(Tile_X8Y3_N4BEG),
    .NN4END(Tile_X8Y3_NN4BEG),
    .Ci(Tile_X8Y3_Co),
    .E1END(Tile_X7Y2_E1BEG),
    .E2MID(Tile_X7Y2_E2BEG),
    .E2END(Tile_X7Y2_E2BEGb),
    .EE4END(Tile_X7Y2_EE4BEG),
    .E6END(Tile_X7Y2_E6BEG),
    .S1END(Tile_X8Y1_S1BEG),
    .S2MID(Tile_X8Y1_S2BEG),
    .S2END(Tile_X8Y1_S2BEGb),
    .S4END(Tile_X8Y1_S4BEG),
    .SS4END(Tile_X8Y1_SS4BEG),
    .W1END(Tile_X9Y2_W1BEG),
    .W2MID(Tile_X9Y2_W2BEG),
    .W2END(Tile_X9Y2_W2BEGb),
    .WW4END(Tile_X9Y2_WW4BEG),
    .W6END(Tile_X9Y2_W6BEG),
    .N1BEG(Tile_X8Y2_N1BEG),
    .N2BEG(Tile_X8Y2_N2BEG),
    .N2BEGb(Tile_X8Y2_N2BEGb),
    .N4BEG(Tile_X8Y2_N4BEG),
    .NN4BEG(Tile_X8Y2_NN4BEG),
    .E1BEG(Tile_X8Y2_E1BEG),
    .E2BEG(Tile_X8Y2_E2BEG),
    .E2BEGb(Tile_X8Y2_E2BEGb),
    .EE4BEG(Tile_X8Y2_EE4BEG),
    .E6BEG(Tile_X8Y2_E6BEG),
    .S1BEG(Tile_X8Y2_S1BEG),
    .S2BEG(Tile_X8Y2_S2BEG),
    .S2BEGb(Tile_X8Y2_S2BEGb),
    .S4BEG(Tile_X8Y2_S4BEG),
    .SS4BEG(Tile_X8Y2_SS4BEG),
    .W1BEG(Tile_X8Y2_W1BEG),
    .W2BEG(Tile_X8Y2_W2BEG),
    .W2BEGb(Tile_X8Y2_W2BEGb),
    .WW4BEG(Tile_X8Y2_WW4BEG),
    .W6BEG(Tile_X8Y2_W6BEG),
    .Co(Tile_X8Y2_Co),
    .UserCLK(Tile_X8Y3_UserCLKo),
    .UserCLKo(Tile_X8Y2_UserCLKo),
    .FrameData(Tile_X7Y2_FrameData_O),
    .FrameData_O(Tile_X8Y2_FrameData_O),
    .FrameStrobe(Tile_X8Y3_FrameStrobe_O),
    .FrameStrobe_O(Tile_X8Y2_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X9Y2_Emulate_Bitstream)
    )
`endif
    Tile_X9Y2_LUT4AB
    (
    .N1END(Tile_X9Y3_N1BEG),
    .N2MID(Tile_X9Y3_N2BEG),
    .N2END(Tile_X9Y3_N2BEGb),
    .N4END(Tile_X9Y3_N4BEG),
    .NN4END(Tile_X9Y3_NN4BEG),
    .Ci(Tile_X9Y3_Co),
    .E1END(Tile_X8Y2_E1BEG),
    .E2MID(Tile_X8Y2_E2BEG),
    .E2END(Tile_X8Y2_E2BEGb),
    .EE4END(Tile_X8Y2_EE4BEG),
    .E6END(Tile_X8Y2_E6BEG),
    .S1END(Tile_X9Y1_S1BEG),
    .S2MID(Tile_X9Y1_S2BEG),
    .S2END(Tile_X9Y1_S2BEGb),
    .S4END(Tile_X9Y1_S4BEG),
    .SS4END(Tile_X9Y1_SS4BEG),
    .W1END(Tile_X10Y2_W1BEG),
    .W2MID(Tile_X10Y2_W2BEG),
    .W2END(Tile_X10Y2_W2BEGb),
    .WW4END(Tile_X10Y2_WW4BEG),
    .W6END(Tile_X10Y2_W6BEG),
    .N1BEG(Tile_X9Y2_N1BEG),
    .N2BEG(Tile_X9Y2_N2BEG),
    .N2BEGb(Tile_X9Y2_N2BEGb),
    .N4BEG(Tile_X9Y2_N4BEG),
    .NN4BEG(Tile_X9Y2_NN4BEG),
    .E1BEG(Tile_X9Y2_E1BEG),
    .E2BEG(Tile_X9Y2_E2BEG),
    .E2BEGb(Tile_X9Y2_E2BEGb),
    .EE4BEG(Tile_X9Y2_EE4BEG),
    .E6BEG(Tile_X9Y2_E6BEG),
    .S1BEG(Tile_X9Y2_S1BEG),
    .S2BEG(Tile_X9Y2_S2BEG),
    .S2BEGb(Tile_X9Y2_S2BEGb),
    .S4BEG(Tile_X9Y2_S4BEG),
    .SS4BEG(Tile_X9Y2_SS4BEG),
    .W1BEG(Tile_X9Y2_W1BEG),
    .W2BEG(Tile_X9Y2_W2BEG),
    .W2BEGb(Tile_X9Y2_W2BEGb),
    .WW4BEG(Tile_X9Y2_WW4BEG),
    .W6BEG(Tile_X9Y2_W6BEG),
    .Co(Tile_X9Y2_Co),
    .UserCLK(Tile_X9Y3_UserCLKo),
    .UserCLKo(Tile_X9Y2_UserCLKo),
    .FrameData(Tile_X8Y2_FrameData_O),
    .FrameData_O(Tile_X9Y2_FrameData_O),
    .FrameStrobe(Tile_X9Y3_FrameStrobe_O),
    .FrameStrobe_O(Tile_X9Y2_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
W_IO
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X0Y3_Emulate_Bitstream)
    )
`endif
    Tile_X0Y3_W_IO
    (
    .W1END(Tile_X1Y3_W1BEG),
    .W2MID(Tile_X1Y3_W2BEG),
    .W2END(Tile_X1Y3_W2BEGb),
    .WW4END(Tile_X1Y3_WW4BEG),
    .W6END(Tile_X1Y3_W6BEG),
    .E1BEG(Tile_X0Y3_E1BEG),
    .E2BEG(Tile_X0Y3_E2BEG),
    .E2BEGb(Tile_X0Y3_E2BEGb),
    .EE4BEG(Tile_X0Y3_EE4BEG),
    .E6BEG(Tile_X0Y3_E6BEG),
    .A_O_top(Tile_X0Y3_A_O_top),
    .A_I_top(Tile_X0Y3_A_I_top),
    .A_T_top(Tile_X0Y3_A_T_top),
    .B_O_top(Tile_X0Y3_B_O_top),
    .B_I_top(Tile_X0Y3_B_I_top),
    .B_T_top(Tile_X0Y3_B_T_top),
    .A_config_C_bit0(Tile_X0Y3_A_config_C_bit0),
    .A_config_C_bit1(Tile_X0Y3_A_config_C_bit1),
    .A_config_C_bit2(Tile_X0Y3_A_config_C_bit2),
    .A_config_C_bit3(Tile_X0Y3_A_config_C_bit3),
    .B_config_C_bit0(Tile_X0Y3_B_config_C_bit0),
    .B_config_C_bit1(Tile_X0Y3_B_config_C_bit1),
    .B_config_C_bit2(Tile_X0Y3_B_config_C_bit2),
    .B_config_C_bit3(Tile_X0Y3_B_config_C_bit3),
    .UserCLK(Tile_X0Y4_UserCLKo),
    .UserCLKo(Tile_X0Y3_UserCLKo),
    .FrameData(Row_Y3_FrameData),
    .FrameData_O(Tile_X0Y3_FrameData_O),
    .FrameStrobe(Tile_X0Y4_FrameStrobe_O),
    .FrameStrobe_O(Tile_X0Y3_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X1Y3_Emulate_Bitstream)
    )
`endif
    Tile_X1Y3_LUT4AB
    (
    .N1END(Tile_X1Y4_N1BEG),
    .N2MID(Tile_X1Y4_N2BEG),
    .N2END(Tile_X1Y4_N2BEGb),
    .N4END(Tile_X1Y4_N4BEG),
    .NN4END(Tile_X1Y4_NN4BEG),
    .Ci(Tile_X1Y4_Co),
    .E1END(Tile_X0Y3_E1BEG),
    .E2MID(Tile_X0Y3_E2BEG),
    .E2END(Tile_X0Y3_E2BEGb),
    .EE4END(Tile_X0Y3_EE4BEG),
    .E6END(Tile_X0Y3_E6BEG),
    .S1END(Tile_X1Y2_S1BEG),
    .S2MID(Tile_X1Y2_S2BEG),
    .S2END(Tile_X1Y2_S2BEGb),
    .S4END(Tile_X1Y2_S4BEG),
    .SS4END(Tile_X1Y2_SS4BEG),
    .W1END(Tile_X2Y3_W1BEG),
    .W2MID(Tile_X2Y3_W2BEG),
    .W2END(Tile_X2Y3_W2BEGb),
    .WW4END(Tile_X2Y3_WW4BEG),
    .W6END(Tile_X2Y3_W6BEG),
    .N1BEG(Tile_X1Y3_N1BEG),
    .N2BEG(Tile_X1Y3_N2BEG),
    .N2BEGb(Tile_X1Y3_N2BEGb),
    .N4BEG(Tile_X1Y3_N4BEG),
    .NN4BEG(Tile_X1Y3_NN4BEG),
    .E1BEG(Tile_X1Y3_E1BEG),
    .E2BEG(Tile_X1Y3_E2BEG),
    .E2BEGb(Tile_X1Y3_E2BEGb),
    .EE4BEG(Tile_X1Y3_EE4BEG),
    .E6BEG(Tile_X1Y3_E6BEG),
    .S1BEG(Tile_X1Y3_S1BEG),
    .S2BEG(Tile_X1Y3_S2BEG),
    .S2BEGb(Tile_X1Y3_S2BEGb),
    .S4BEG(Tile_X1Y3_S4BEG),
    .SS4BEG(Tile_X1Y3_SS4BEG),
    .W1BEG(Tile_X1Y3_W1BEG),
    .W2BEG(Tile_X1Y3_W2BEG),
    .W2BEGb(Tile_X1Y3_W2BEGb),
    .WW4BEG(Tile_X1Y3_WW4BEG),
    .W6BEG(Tile_X1Y3_W6BEG),
    .Co(Tile_X1Y3_Co),
    .UserCLK(Tile_X1Y4_UserCLKo),
    .UserCLKo(Tile_X1Y3_UserCLKo),
    .FrameData(Tile_X0Y3_FrameData_O),
    .FrameData_O(Tile_X1Y3_FrameData_O),
    .FrameStrobe(Tile_X1Y4_FrameStrobe_O),
    .FrameStrobe_O(Tile_X1Y3_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X2Y3_Emulate_Bitstream)
    )
`endif
    Tile_X2Y3_LUT4AB
    (
    .N1END(Tile_X2Y4_N1BEG),
    .N2MID(Tile_X2Y4_N2BEG),
    .N2END(Tile_X2Y4_N2BEGb),
    .N4END(Tile_X2Y4_N4BEG),
    .NN4END(Tile_X2Y4_NN4BEG),
    .Ci(Tile_X2Y4_Co),
    .E1END(Tile_X1Y3_E1BEG),
    .E2MID(Tile_X1Y3_E2BEG),
    .E2END(Tile_X1Y3_E2BEGb),
    .EE4END(Tile_X1Y3_EE4BEG),
    .E6END(Tile_X1Y3_E6BEG),
    .S1END(Tile_X2Y2_S1BEG),
    .S2MID(Tile_X2Y2_S2BEG),
    .S2END(Tile_X2Y2_S2BEGb),
    .S4END(Tile_X2Y2_S4BEG),
    .SS4END(Tile_X2Y2_SS4BEG),
    .W1END(Tile_X3Y3_W1BEG),
    .W2MID(Tile_X3Y3_W2BEG),
    .W2END(Tile_X3Y3_W2BEGb),
    .WW4END(Tile_X3Y3_WW4BEG),
    .W6END(Tile_X3Y3_W6BEG),
    .N1BEG(Tile_X2Y3_N1BEG),
    .N2BEG(Tile_X2Y3_N2BEG),
    .N2BEGb(Tile_X2Y3_N2BEGb),
    .N4BEG(Tile_X2Y3_N4BEG),
    .NN4BEG(Tile_X2Y3_NN4BEG),
    .E1BEG(Tile_X2Y3_E1BEG),
    .E2BEG(Tile_X2Y3_E2BEG),
    .E2BEGb(Tile_X2Y3_E2BEGb),
    .EE4BEG(Tile_X2Y3_EE4BEG),
    .E6BEG(Tile_X2Y3_E6BEG),
    .S1BEG(Tile_X2Y3_S1BEG),
    .S2BEG(Tile_X2Y3_S2BEG),
    .S2BEGb(Tile_X2Y3_S2BEGb),
    .S4BEG(Tile_X2Y3_S4BEG),
    .SS4BEG(Tile_X2Y3_SS4BEG),
    .W1BEG(Tile_X2Y3_W1BEG),
    .W2BEG(Tile_X2Y3_W2BEG),
    .W2BEGb(Tile_X2Y3_W2BEGb),
    .WW4BEG(Tile_X2Y3_WW4BEG),
    .W6BEG(Tile_X2Y3_W6BEG),
    .Co(Tile_X2Y3_Co),
    .UserCLK(Tile_X2Y4_UserCLKo),
    .UserCLKo(Tile_X2Y3_UserCLKo),
    .FrameData(Tile_X1Y3_FrameData_O),
    .FrameData_O(Tile_X2Y3_FrameData_O),
    .FrameStrobe(Tile_X2Y4_FrameStrobe_O),
    .FrameStrobe_O(Tile_X2Y3_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X3Y3_Emulate_Bitstream)
    )
`endif
    Tile_X3Y3_LUT4AB
    (
    .N1END(Tile_X3Y4_N1BEG),
    .N2MID(Tile_X3Y4_N2BEG),
    .N2END(Tile_X3Y4_N2BEGb),
    .N4END(Tile_X3Y4_N4BEG),
    .NN4END(Tile_X3Y4_NN4BEG),
    .Ci(Tile_X3Y4_Co),
    .E1END(Tile_X2Y3_E1BEG),
    .E2MID(Tile_X2Y3_E2BEG),
    .E2END(Tile_X2Y3_E2BEGb),
    .EE4END(Tile_X2Y3_EE4BEG),
    .E6END(Tile_X2Y3_E6BEG),
    .S1END(Tile_X3Y2_S1BEG),
    .S2MID(Tile_X3Y2_S2BEG),
    .S2END(Tile_X3Y2_S2BEGb),
    .S4END(Tile_X3Y2_S4BEG),
    .SS4END(Tile_X3Y2_SS4BEG),
    .W1END(Tile_X4Y3_W1BEG),
    .W2MID(Tile_X4Y3_W2BEG),
    .W2END(Tile_X4Y3_W2BEGb),
    .WW4END(Tile_X4Y3_WW4BEG),
    .W6END(Tile_X4Y3_W6BEG),
    .N1BEG(Tile_X3Y3_N1BEG),
    .N2BEG(Tile_X3Y3_N2BEG),
    .N2BEGb(Tile_X3Y3_N2BEGb),
    .N4BEG(Tile_X3Y3_N4BEG),
    .NN4BEG(Tile_X3Y3_NN4BEG),
    .E1BEG(Tile_X3Y3_E1BEG),
    .E2BEG(Tile_X3Y3_E2BEG),
    .E2BEGb(Tile_X3Y3_E2BEGb),
    .EE4BEG(Tile_X3Y3_EE4BEG),
    .E6BEG(Tile_X3Y3_E6BEG),
    .S1BEG(Tile_X3Y3_S1BEG),
    .S2BEG(Tile_X3Y3_S2BEG),
    .S2BEGb(Tile_X3Y3_S2BEGb),
    .S4BEG(Tile_X3Y3_S4BEG),
    .SS4BEG(Tile_X3Y3_SS4BEG),
    .W1BEG(Tile_X3Y3_W1BEG),
    .W2BEG(Tile_X3Y3_W2BEG),
    .W2BEGb(Tile_X3Y3_W2BEGb),
    .WW4BEG(Tile_X3Y3_WW4BEG),
    .W6BEG(Tile_X3Y3_W6BEG),
    .Co(Tile_X3Y3_Co),
    .UserCLK(Tile_X3Y4_UserCLKo),
    .UserCLKo(Tile_X3Y3_UserCLKo),
    .FrameData(Tile_X2Y3_FrameData_O),
    .FrameData_O(Tile_X3Y3_FrameData_O),
    .FrameStrobe(Tile_X3Y4_FrameStrobe_O),
    .FrameStrobe_O(Tile_X3Y3_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
RegFile
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X4Y3_Emulate_Bitstream)
    )
`endif
    Tile_X4Y3_RegFile
    (
    .N1END(Tile_X4Y4_N1BEG),
    .N2MID(Tile_X4Y4_N2BEG),
    .N2END(Tile_X4Y4_N2BEGb),
    .N4END(Tile_X4Y4_N4BEG),
    .NN4END(Tile_X4Y4_NN4BEG),
    .E1END(Tile_X3Y3_E1BEG),
    .E2MID(Tile_X3Y3_E2BEG),
    .E2END(Tile_X3Y3_E2BEGb),
    .EE4END(Tile_X3Y3_EE4BEG),
    .E6END(Tile_X3Y3_E6BEG),
    .S1END(Tile_X4Y2_S1BEG),
    .S2MID(Tile_X4Y2_S2BEG),
    .S2END(Tile_X4Y2_S2BEGb),
    .S4END(Tile_X4Y2_S4BEG),
    .SS4END(Tile_X4Y2_SS4BEG),
    .W1END(Tile_X5Y3_W1BEG),
    .W2MID(Tile_X5Y3_W2BEG),
    .W2END(Tile_X5Y3_W2BEGb),
    .WW4END(Tile_X5Y3_WW4BEG),
    .W6END(Tile_X5Y3_W6BEG),
    .N1BEG(Tile_X4Y3_N1BEG),
    .N2BEG(Tile_X4Y3_N2BEG),
    .N2BEGb(Tile_X4Y3_N2BEGb),
    .N4BEG(Tile_X4Y3_N4BEG),
    .NN4BEG(Tile_X4Y3_NN4BEG),
    .E1BEG(Tile_X4Y3_E1BEG),
    .E2BEG(Tile_X4Y3_E2BEG),
    .E2BEGb(Tile_X4Y3_E2BEGb),
    .EE4BEG(Tile_X4Y3_EE4BEG),
    .E6BEG(Tile_X4Y3_E6BEG),
    .S1BEG(Tile_X4Y3_S1BEG),
    .S2BEG(Tile_X4Y3_S2BEG),
    .S2BEGb(Tile_X4Y3_S2BEGb),
    .S4BEG(Tile_X4Y3_S4BEG),
    .SS4BEG(Tile_X4Y3_SS4BEG),
    .W1BEG(Tile_X4Y3_W1BEG),
    .W2BEG(Tile_X4Y3_W2BEG),
    .W2BEGb(Tile_X4Y3_W2BEGb),
    .WW4BEG(Tile_X4Y3_WW4BEG),
    .W6BEG(Tile_X4Y3_W6BEG),
    .UserCLK(Tile_X4Y4_UserCLKo),
    .UserCLKo(Tile_X4Y3_UserCLKo),
    .FrameData(Tile_X3Y3_FrameData_O),
    .FrameData_O(Tile_X4Y3_FrameData_O),
    .FrameStrobe(Tile_X4Y4_FrameStrobe_O),
    .FrameStrobe_O(Tile_X4Y3_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X5Y3_Emulate_Bitstream)
    )
`endif
    Tile_X5Y3_LUT4AB
    (
    .N1END(Tile_X5Y4_N1BEG),
    .N2MID(Tile_X5Y4_N2BEG),
    .N2END(Tile_X5Y4_N2BEGb),
    .N4END(Tile_X5Y4_N4BEG),
    .NN4END(Tile_X5Y4_NN4BEG),
    .Ci(Tile_X5Y4_Co),
    .E1END(Tile_X4Y3_E1BEG),
    .E2MID(Tile_X4Y3_E2BEG),
    .E2END(Tile_X4Y3_E2BEGb),
    .EE4END(Tile_X4Y3_EE4BEG),
    .E6END(Tile_X4Y3_E6BEG),
    .S1END(Tile_X5Y2_S1BEG),
    .S2MID(Tile_X5Y2_S2BEG),
    .S2END(Tile_X5Y2_S2BEGb),
    .S4END(Tile_X5Y2_S4BEG),
    .SS4END(Tile_X5Y2_SS4BEG),
    .W1END(Tile_X6Y3_W1BEG),
    .W2MID(Tile_X6Y3_W2BEG),
    .W2END(Tile_X6Y3_W2BEGb),
    .WW4END(Tile_X6Y3_WW4BEG),
    .W6END(Tile_X6Y3_W6BEG),
    .N1BEG(Tile_X5Y3_N1BEG),
    .N2BEG(Tile_X5Y3_N2BEG),
    .N2BEGb(Tile_X5Y3_N2BEGb),
    .N4BEG(Tile_X5Y3_N4BEG),
    .NN4BEG(Tile_X5Y3_NN4BEG),
    .E1BEG(Tile_X5Y3_E1BEG),
    .E2BEG(Tile_X5Y3_E2BEG),
    .E2BEGb(Tile_X5Y3_E2BEGb),
    .EE4BEG(Tile_X5Y3_EE4BEG),
    .E6BEG(Tile_X5Y3_E6BEG),
    .S1BEG(Tile_X5Y3_S1BEG),
    .S2BEG(Tile_X5Y3_S2BEG),
    .S2BEGb(Tile_X5Y3_S2BEGb),
    .S4BEG(Tile_X5Y3_S4BEG),
    .SS4BEG(Tile_X5Y3_SS4BEG),
    .W1BEG(Tile_X5Y3_W1BEG),
    .W2BEG(Tile_X5Y3_W2BEG),
    .W2BEGb(Tile_X5Y3_W2BEGb),
    .WW4BEG(Tile_X5Y3_WW4BEG),
    .W6BEG(Tile_X5Y3_W6BEG),
    .Co(Tile_X5Y3_Co),
    .UserCLK(Tile_X5Y4_UserCLKo),
    .UserCLKo(Tile_X5Y3_UserCLKo),
    .FrameData(Tile_X4Y3_FrameData_O),
    .FrameData_O(Tile_X5Y3_FrameData_O),
    .FrameStrobe(Tile_X5Y4_FrameStrobe_O),
    .FrameStrobe_O(Tile_X5Y3_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X6Y3_Emulate_Bitstream)
    )
`endif
    Tile_X6Y3_LUT4AB
    (
    .N1END(Tile_X6Y4_N1BEG),
    .N2MID(Tile_X6Y4_N2BEG),
    .N2END(Tile_X6Y4_N2BEGb),
    .N4END(Tile_X6Y4_N4BEG),
    .NN4END(Tile_X6Y4_NN4BEG),
    .Ci(Tile_X6Y4_Co),
    .E1END(Tile_X5Y3_E1BEG),
    .E2MID(Tile_X5Y3_E2BEG),
    .E2END(Tile_X5Y3_E2BEGb),
    .EE4END(Tile_X5Y3_EE4BEG),
    .E6END(Tile_X5Y3_E6BEG),
    .S1END(Tile_X6Y2_S1BEG),
    .S2MID(Tile_X6Y2_S2BEG),
    .S2END(Tile_X6Y2_S2BEGb),
    .S4END(Tile_X6Y2_S4BEG),
    .SS4END(Tile_X6Y2_SS4BEG),
    .W1END(Tile_X7Y3_W1BEG),
    .W2MID(Tile_X7Y3_W2BEG),
    .W2END(Tile_X7Y3_W2BEGb),
    .WW4END(Tile_X7Y3_WW4BEG),
    .W6END(Tile_X7Y3_W6BEG),
    .N1BEG(Tile_X6Y3_N1BEG),
    .N2BEG(Tile_X6Y3_N2BEG),
    .N2BEGb(Tile_X6Y3_N2BEGb),
    .N4BEG(Tile_X6Y3_N4BEG),
    .NN4BEG(Tile_X6Y3_NN4BEG),
    .E1BEG(Tile_X6Y3_E1BEG),
    .E2BEG(Tile_X6Y3_E2BEG),
    .E2BEGb(Tile_X6Y3_E2BEGb),
    .EE4BEG(Tile_X6Y3_EE4BEG),
    .E6BEG(Tile_X6Y3_E6BEG),
    .S1BEG(Tile_X6Y3_S1BEG),
    .S2BEG(Tile_X6Y3_S2BEG),
    .S2BEGb(Tile_X6Y3_S2BEGb),
    .S4BEG(Tile_X6Y3_S4BEG),
    .SS4BEG(Tile_X6Y3_SS4BEG),
    .W1BEG(Tile_X6Y3_W1BEG),
    .W2BEG(Tile_X6Y3_W2BEG),
    .W2BEGb(Tile_X6Y3_W2BEGb),
    .WW4BEG(Tile_X6Y3_WW4BEG),
    .W6BEG(Tile_X6Y3_W6BEG),
    .Co(Tile_X6Y3_Co),
    .UserCLK(Tile_X6Y4_UserCLKo),
    .UserCLKo(Tile_X6Y3_UserCLKo),
    .FrameData(Tile_X5Y3_FrameData_O),
    .FrameData_O(Tile_X6Y3_FrameData_O),
    .FrameStrobe(Tile_X6Y4_FrameStrobe_O),
    .FrameStrobe_O(Tile_X6Y3_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
DSP
`ifdef EMULATION
    #(
    .Tile_X0Y0_Emulate_Bitstream(`Tile_X7Y3_Emulate_Bitstream),
    .Tile_X0Y1_Emulate_Bitstream(`Tile_X7Y4_Emulate_Bitstream)
    )
`endif
    Tile_X7Y3_DSP
    (
    .Tile_X0Y0_E1END(Tile_X6Y3_E1BEG),
    .Tile_X0Y0_E2MID(Tile_X6Y3_E2BEG),
    .Tile_X0Y0_E2END(Tile_X6Y3_E2BEGb),
    .Tile_X0Y0_EE4END(Tile_X6Y3_EE4BEG),
    .Tile_X0Y0_E6END(Tile_X6Y3_E6BEG),
    .Tile_X0Y0_S1END(Tile_X7Y2_S1BEG),
    .Tile_X0Y0_S2MID(Tile_X7Y2_S2BEG),
    .Tile_X0Y0_S2END(Tile_X7Y2_S2BEGb),
    .Tile_X0Y0_S4END(Tile_X7Y2_S4BEG),
    .Tile_X0Y0_SS4END(Tile_X7Y2_SS4BEG),
    .Tile_X0Y0_W1END(Tile_X8Y3_W1BEG),
    .Tile_X0Y0_W2MID(Tile_X8Y3_W2BEG),
    .Tile_X0Y0_W2END(Tile_X8Y3_W2BEGb),
    .Tile_X0Y0_WW4END(Tile_X8Y3_WW4BEG),
    .Tile_X0Y0_W6END(Tile_X8Y3_W6BEG),
    .Tile_X0Y1_N1END(Tile_X7Y5_N1BEG),
    .Tile_X0Y1_N2MID(Tile_X7Y5_N2BEG),
    .Tile_X0Y1_N2END(Tile_X7Y5_N2BEGb),
    .Tile_X0Y1_N4END(Tile_X7Y5_N4BEG),
    .Tile_X0Y1_NN4END(Tile_X7Y5_NN4BEG),
    .Tile_X0Y1_E1END(Tile_X6Y4_E1BEG),
    .Tile_X0Y1_E2MID(Tile_X6Y4_E2BEG),
    .Tile_X0Y1_E2END(Tile_X6Y4_E2BEGb),
    .Tile_X0Y1_EE4END(Tile_X6Y4_EE4BEG),
    .Tile_X0Y1_E6END(Tile_X6Y4_E6BEG),
    .Tile_X0Y1_W1END(Tile_X8Y4_W1BEG),
    .Tile_X0Y1_W2MID(Tile_X8Y4_W2BEG),
    .Tile_X0Y1_W2END(Tile_X8Y4_W2BEGb),
    .Tile_X0Y1_WW4END(Tile_X8Y4_WW4BEG),
    .Tile_X0Y1_W6END(Tile_X8Y4_W6BEG),
    .Tile_X0Y0_N1BEG(Tile_X7Y3_N1BEG),
    .Tile_X0Y0_N2BEG(Tile_X7Y3_N2BEG),
    .Tile_X0Y0_N2BEGb(Tile_X7Y3_N2BEGb),
    .Tile_X0Y0_N4BEG(Tile_X7Y3_N4BEG),
    .Tile_X0Y0_NN4BEG(Tile_X7Y3_NN4BEG),
    .Tile_X0Y0_E1BEG(Tile_X7Y3_E1BEG),
    .Tile_X0Y0_E2BEG(Tile_X7Y3_E2BEG),
    .Tile_X0Y0_E2BEGb(Tile_X7Y3_E2BEGb),
    .Tile_X0Y0_EE4BEG(Tile_X7Y3_EE4BEG),
    .Tile_X0Y0_E6BEG(Tile_X7Y3_E6BEG),
    .Tile_X0Y0_W1BEG(Tile_X7Y3_W1BEG),
    .Tile_X0Y0_W2BEG(Tile_X7Y3_W2BEG),
    .Tile_X0Y0_W2BEGb(Tile_X7Y3_W2BEGb),
    .Tile_X0Y0_WW4BEG(Tile_X7Y3_WW4BEG),
    .Tile_X0Y0_W6BEG(Tile_X7Y3_W6BEG),
    .Tile_X0Y1_E1BEG(Tile_X7Y4_E1BEG),
    .Tile_X0Y1_E2BEG(Tile_X7Y4_E2BEG),
    .Tile_X0Y1_E2BEGb(Tile_X7Y4_E2BEGb),
    .Tile_X0Y1_EE4BEG(Tile_X7Y4_EE4BEG),
    .Tile_X0Y1_E6BEG(Tile_X7Y4_E6BEG),
    .Tile_X0Y1_S1BEG(Tile_X7Y4_S1BEG),
    .Tile_X0Y1_S2BEG(Tile_X7Y4_S2BEG),
    .Tile_X0Y1_S2BEGb(Tile_X7Y4_S2BEGb),
    .Tile_X0Y1_S4BEG(Tile_X7Y4_S4BEG),
    .Tile_X0Y1_SS4BEG(Tile_X7Y4_SS4BEG),
    .Tile_X0Y1_W1BEG(Tile_X7Y4_W1BEG),
    .Tile_X0Y1_W2BEG(Tile_X7Y4_W2BEG),
    .Tile_X0Y1_W2BEGb(Tile_X7Y4_W2BEGb),
    .Tile_X0Y1_WW4BEG(Tile_X7Y4_WW4BEG),
    .Tile_X0Y1_W6BEG(Tile_X7Y4_W6BEG),
    .Tile_X0Y0_UserCLKo(Tile_X7Y3_UserCLKo),
    .Tile_X0Y1_UserCLK(Tile_X7Y5_UserCLKo),
    .Tile_X0Y0_FrameData(Tile_X6Y3_FrameData_O),
    .Tile_X0Y0_FrameData_O(Tile_X7Y3_FrameData_O),
    .Tile_X0Y0_FrameStrobe_O(Tile_X7Y3_FrameStrobe_O),
    .Tile_X0Y1_FrameData(Tile_X6Y4_FrameData_O),
    .Tile_X0Y1_FrameData_O(Tile_X7Y4_FrameData_O),
    .Tile_X0Y1_FrameStrobe(Tile_X7Y5_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X8Y3_Emulate_Bitstream)
    )
`endif
    Tile_X8Y3_LUT4AB
    (
    .N1END(Tile_X8Y4_N1BEG),
    .N2MID(Tile_X8Y4_N2BEG),
    .N2END(Tile_X8Y4_N2BEGb),
    .N4END(Tile_X8Y4_N4BEG),
    .NN4END(Tile_X8Y4_NN4BEG),
    .Ci(Tile_X8Y4_Co),
    .E1END(Tile_X7Y3_E1BEG),
    .E2MID(Tile_X7Y3_E2BEG),
    .E2END(Tile_X7Y3_E2BEGb),
    .EE4END(Tile_X7Y3_EE4BEG),
    .E6END(Tile_X7Y3_E6BEG),
    .S1END(Tile_X8Y2_S1BEG),
    .S2MID(Tile_X8Y2_S2BEG),
    .S2END(Tile_X8Y2_S2BEGb),
    .S4END(Tile_X8Y2_S4BEG),
    .SS4END(Tile_X8Y2_SS4BEG),
    .W1END(Tile_X9Y3_W1BEG),
    .W2MID(Tile_X9Y3_W2BEG),
    .W2END(Tile_X9Y3_W2BEGb),
    .WW4END(Tile_X9Y3_WW4BEG),
    .W6END(Tile_X9Y3_W6BEG),
    .N1BEG(Tile_X8Y3_N1BEG),
    .N2BEG(Tile_X8Y3_N2BEG),
    .N2BEGb(Tile_X8Y3_N2BEGb),
    .N4BEG(Tile_X8Y3_N4BEG),
    .NN4BEG(Tile_X8Y3_NN4BEG),
    .E1BEG(Tile_X8Y3_E1BEG),
    .E2BEG(Tile_X8Y3_E2BEG),
    .E2BEGb(Tile_X8Y3_E2BEGb),
    .EE4BEG(Tile_X8Y3_EE4BEG),
    .E6BEG(Tile_X8Y3_E6BEG),
    .S1BEG(Tile_X8Y3_S1BEG),
    .S2BEG(Tile_X8Y3_S2BEG),
    .S2BEGb(Tile_X8Y3_S2BEGb),
    .S4BEG(Tile_X8Y3_S4BEG),
    .SS4BEG(Tile_X8Y3_SS4BEG),
    .W1BEG(Tile_X8Y3_W1BEG),
    .W2BEG(Tile_X8Y3_W2BEG),
    .W2BEGb(Tile_X8Y3_W2BEGb),
    .WW4BEG(Tile_X8Y3_WW4BEG),
    .W6BEG(Tile_X8Y3_W6BEG),
    .Co(Tile_X8Y3_Co),
    .UserCLK(Tile_X8Y4_UserCLKo),
    .UserCLKo(Tile_X8Y3_UserCLKo),
    .FrameData(Tile_X7Y3_FrameData_O),
    .FrameData_O(Tile_X8Y3_FrameData_O),
    .FrameStrobe(Tile_X8Y4_FrameStrobe_O),
    .FrameStrobe_O(Tile_X8Y3_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X9Y3_Emulate_Bitstream)
    )
`endif
    Tile_X9Y3_LUT4AB
    (
    .N1END(Tile_X9Y4_N1BEG),
    .N2MID(Tile_X9Y4_N2BEG),
    .N2END(Tile_X9Y4_N2BEGb),
    .N4END(Tile_X9Y4_N4BEG),
    .NN4END(Tile_X9Y4_NN4BEG),
    .Ci(Tile_X9Y4_Co),
    .E1END(Tile_X8Y3_E1BEG),
    .E2MID(Tile_X8Y3_E2BEG),
    .E2END(Tile_X8Y3_E2BEGb),
    .EE4END(Tile_X8Y3_EE4BEG),
    .E6END(Tile_X8Y3_E6BEG),
    .S1END(Tile_X9Y2_S1BEG),
    .S2MID(Tile_X9Y2_S2BEG),
    .S2END(Tile_X9Y2_S2BEGb),
    .S4END(Tile_X9Y2_S4BEG),
    .SS4END(Tile_X9Y2_SS4BEG),
    .W1END(Tile_X10Y3_W1BEG),
    .W2MID(Tile_X10Y3_W2BEG),
    .W2END(Tile_X10Y3_W2BEGb),
    .WW4END(Tile_X10Y3_WW4BEG),
    .W6END(Tile_X10Y3_W6BEG),
    .N1BEG(Tile_X9Y3_N1BEG),
    .N2BEG(Tile_X9Y3_N2BEG),
    .N2BEGb(Tile_X9Y3_N2BEGb),
    .N4BEG(Tile_X9Y3_N4BEG),
    .NN4BEG(Tile_X9Y3_NN4BEG),
    .E1BEG(Tile_X9Y3_E1BEG),
    .E2BEG(Tile_X9Y3_E2BEG),
    .E2BEGb(Tile_X9Y3_E2BEGb),
    .EE4BEG(Tile_X9Y3_EE4BEG),
    .E6BEG(Tile_X9Y3_E6BEG),
    .S1BEG(Tile_X9Y3_S1BEG),
    .S2BEG(Tile_X9Y3_S2BEG),
    .S2BEGb(Tile_X9Y3_S2BEGb),
    .S4BEG(Tile_X9Y3_S4BEG),
    .SS4BEG(Tile_X9Y3_SS4BEG),
    .W1BEG(Tile_X9Y3_W1BEG),
    .W2BEG(Tile_X9Y3_W2BEG),
    .W2BEGb(Tile_X9Y3_W2BEGb),
    .WW4BEG(Tile_X9Y3_WW4BEG),
    .W6BEG(Tile_X9Y3_W6BEG),
    .Co(Tile_X9Y3_Co),
    .UserCLK(Tile_X9Y4_UserCLKo),
    .UserCLKo(Tile_X9Y3_UserCLKo),
    .FrameData(Tile_X8Y3_FrameData_O),
    .FrameData_O(Tile_X9Y3_FrameData_O),
    .FrameStrobe(Tile_X9Y4_FrameStrobe_O),
    .FrameStrobe_O(Tile_X9Y3_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
IHP_SRAM
`ifdef EMULATION
    #(
    .Tile_X0Y0_Emulate_Bitstream(`Tile_X10Y3_Emulate_Bitstream),
    .Tile_X0Y1_Emulate_Bitstream(`Tile_X10Y4_Emulate_Bitstream)
    )
`endif
    Tile_X10Y3_IHP_SRAM
    (
    .Tile_X0Y0_E1END(Tile_X9Y3_E1BEG),
    .Tile_X0Y0_E2MID(Tile_X9Y3_E2BEG),
    .Tile_X0Y0_E2END(Tile_X9Y3_E2BEGb),
    .Tile_X0Y0_EE4END(Tile_X9Y3_EE4BEG),
    .Tile_X0Y0_E6END(Tile_X9Y3_E6BEG),
    .Tile_X0Y0_S1END(Tile_X10Y2_S1BEG),
    .Tile_X0Y0_S2MID(Tile_X10Y2_S2BEG),
    .Tile_X0Y0_S2END(Tile_X10Y2_S2BEGb),
    .Tile_X0Y0_S4END(Tile_X10Y2_S4BEG),
    .Tile_X0Y1_N1END(Tile_X10Y5_N1BEG),
    .Tile_X0Y1_N2MID(Tile_X10Y5_N2BEG),
    .Tile_X0Y1_N2END(Tile_X10Y5_N2BEGb),
    .Tile_X0Y1_N4END(Tile_X10Y5_N4BEG),
    .Tile_X0Y1_E1END(Tile_X9Y4_E1BEG),
    .Tile_X0Y1_E2MID(Tile_X9Y4_E2BEG),
    .Tile_X0Y1_E2END(Tile_X9Y4_E2BEGb),
    .Tile_X0Y1_EE4END(Tile_X9Y4_EE4BEG),
    .Tile_X0Y1_E6END(Tile_X9Y4_E6BEG),
    .Tile_X0Y0_N1BEG(Tile_X10Y3_N1BEG),
    .Tile_X0Y0_N2BEG(Tile_X10Y3_N2BEG),
    .Tile_X0Y0_N2BEGb(Tile_X10Y3_N2BEGb),
    .Tile_X0Y0_N4BEG(Tile_X10Y3_N4BEG),
    .Tile_X0Y0_W1BEG(Tile_X10Y3_W1BEG),
    .Tile_X0Y0_W2BEG(Tile_X10Y3_W2BEG),
    .Tile_X0Y0_W2BEGb(Tile_X10Y3_W2BEGb),
    .Tile_X0Y0_WW4BEG(Tile_X10Y3_WW4BEG),
    .Tile_X0Y0_W6BEG(Tile_X10Y3_W6BEG),
    .Tile_X0Y1_S1BEG(Tile_X10Y4_S1BEG),
    .Tile_X0Y1_S2BEG(Tile_X10Y4_S2BEG),
    .Tile_X0Y1_S2BEGb(Tile_X10Y4_S2BEGb),
    .Tile_X0Y1_S4BEG(Tile_X10Y4_S4BEG),
    .Tile_X0Y1_W1BEG(Tile_X10Y4_W1BEG),
    .Tile_X0Y1_W2BEG(Tile_X10Y4_W2BEG),
    .Tile_X0Y1_W2BEGb(Tile_X10Y4_W2BEGb),
    .Tile_X0Y1_WW4BEG(Tile_X10Y4_WW4BEG),
    .Tile_X0Y1_W6BEG(Tile_X10Y4_W6BEG),
    .CONFIGURED_top(Tile_X10Y4_CONFIGURED_top),
    .DOUT_SRAM0(Tile_X10Y4_DOUT_SRAM0),
    .DOUT_SRAM1(Tile_X10Y4_DOUT_SRAM1),
    .DOUT_SRAM2(Tile_X10Y4_DOUT_SRAM2),
    .DOUT_SRAM3(Tile_X10Y4_DOUT_SRAM3),
    .DOUT_SRAM4(Tile_X10Y4_DOUT_SRAM4),
    .DOUT_SRAM5(Tile_X10Y4_DOUT_SRAM5),
    .DOUT_SRAM6(Tile_X10Y4_DOUT_SRAM6),
    .DOUT_SRAM7(Tile_X10Y4_DOUT_SRAM7),
    .DOUT_SRAM8(Tile_X10Y4_DOUT_SRAM8),
    .DOUT_SRAM9(Tile_X10Y4_DOUT_SRAM9),
    .DOUT_SRAM10(Tile_X10Y4_DOUT_SRAM10),
    .DOUT_SRAM11(Tile_X10Y4_DOUT_SRAM11),
    .DOUT_SRAM12(Tile_X10Y4_DOUT_SRAM12),
    .DOUT_SRAM13(Tile_X10Y4_DOUT_SRAM13),
    .DOUT_SRAM14(Tile_X10Y4_DOUT_SRAM14),
    .DOUT_SRAM15(Tile_X10Y4_DOUT_SRAM15),
    .DOUT_SRAM16(Tile_X10Y4_DOUT_SRAM16),
    .DOUT_SRAM17(Tile_X10Y4_DOUT_SRAM17),
    .DOUT_SRAM18(Tile_X10Y4_DOUT_SRAM18),
    .DOUT_SRAM19(Tile_X10Y4_DOUT_SRAM19),
    .DOUT_SRAM20(Tile_X10Y4_DOUT_SRAM20),
    .DOUT_SRAM21(Tile_X10Y4_DOUT_SRAM21),
    .DOUT_SRAM22(Tile_X10Y4_DOUT_SRAM22),
    .DOUT_SRAM23(Tile_X10Y4_DOUT_SRAM23),
    .DOUT_SRAM24(Tile_X10Y4_DOUT_SRAM24),
    .DOUT_SRAM25(Tile_X10Y4_DOUT_SRAM25),
    .DOUT_SRAM26(Tile_X10Y4_DOUT_SRAM26),
    .DOUT_SRAM27(Tile_X10Y4_DOUT_SRAM27),
    .DOUT_SRAM28(Tile_X10Y4_DOUT_SRAM28),
    .DOUT_SRAM29(Tile_X10Y4_DOUT_SRAM29),
    .DOUT_SRAM30(Tile_X10Y4_DOUT_SRAM30),
    .DOUT_SRAM31(Tile_X10Y4_DOUT_SRAM31),
    .ADDR_SRAM0(Tile_X10Y4_ADDR_SRAM0),
    .ADDR_SRAM1(Tile_X10Y4_ADDR_SRAM1),
    .ADDR_SRAM2(Tile_X10Y4_ADDR_SRAM2),
    .ADDR_SRAM3(Tile_X10Y4_ADDR_SRAM3),
    .ADDR_SRAM4(Tile_X10Y4_ADDR_SRAM4),
    .ADDR_SRAM5(Tile_X10Y4_ADDR_SRAM5),
    .ADDR_SRAM6(Tile_X10Y4_ADDR_SRAM6),
    .ADDR_SRAM7(Tile_X10Y4_ADDR_SRAM7),
    .ADDR_SRAM8(Tile_X10Y4_ADDR_SRAM8),
    .ADDR_SRAM9(Tile_X10Y4_ADDR_SRAM9),
    .BM_SRAM0(Tile_X10Y4_BM_SRAM0),
    .BM_SRAM1(Tile_X10Y4_BM_SRAM1),
    .BM_SRAM2(Tile_X10Y4_BM_SRAM2),
    .BM_SRAM3(Tile_X10Y4_BM_SRAM3),
    .BM_SRAM4(Tile_X10Y4_BM_SRAM4),
    .BM_SRAM5(Tile_X10Y4_BM_SRAM5),
    .BM_SRAM6(Tile_X10Y4_BM_SRAM6),
    .BM_SRAM7(Tile_X10Y4_BM_SRAM7),
    .BM_SRAM8(Tile_X10Y4_BM_SRAM8),
    .BM_SRAM9(Tile_X10Y4_BM_SRAM9),
    .BM_SRAM10(Tile_X10Y4_BM_SRAM10),
    .BM_SRAM11(Tile_X10Y4_BM_SRAM11),
    .BM_SRAM12(Tile_X10Y4_BM_SRAM12),
    .BM_SRAM13(Tile_X10Y4_BM_SRAM13),
    .BM_SRAM14(Tile_X10Y4_BM_SRAM14),
    .BM_SRAM15(Tile_X10Y4_BM_SRAM15),
    .BM_SRAM16(Tile_X10Y4_BM_SRAM16),
    .BM_SRAM17(Tile_X10Y4_BM_SRAM17),
    .BM_SRAM18(Tile_X10Y4_BM_SRAM18),
    .BM_SRAM19(Tile_X10Y4_BM_SRAM19),
    .BM_SRAM20(Tile_X10Y4_BM_SRAM20),
    .BM_SRAM21(Tile_X10Y4_BM_SRAM21),
    .BM_SRAM22(Tile_X10Y4_BM_SRAM22),
    .BM_SRAM23(Tile_X10Y4_BM_SRAM23),
    .BM_SRAM24(Tile_X10Y4_BM_SRAM24),
    .BM_SRAM25(Tile_X10Y4_BM_SRAM25),
    .BM_SRAM26(Tile_X10Y4_BM_SRAM26),
    .BM_SRAM27(Tile_X10Y4_BM_SRAM27),
    .BM_SRAM28(Tile_X10Y4_BM_SRAM28),
    .BM_SRAM29(Tile_X10Y4_BM_SRAM29),
    .BM_SRAM30(Tile_X10Y4_BM_SRAM30),
    .BM_SRAM31(Tile_X10Y4_BM_SRAM31),
    .CLK_SRAM(Tile_X10Y4_CLK_SRAM),
    .DIN_SRAM0(Tile_X10Y4_DIN_SRAM0),
    .DIN_SRAM1(Tile_X10Y4_DIN_SRAM1),
    .DIN_SRAM2(Tile_X10Y4_DIN_SRAM2),
    .DIN_SRAM3(Tile_X10Y4_DIN_SRAM3),
    .DIN_SRAM4(Tile_X10Y4_DIN_SRAM4),
    .DIN_SRAM5(Tile_X10Y4_DIN_SRAM5),
    .DIN_SRAM6(Tile_X10Y4_DIN_SRAM6),
    .DIN_SRAM7(Tile_X10Y4_DIN_SRAM7),
    .DIN_SRAM8(Tile_X10Y4_DIN_SRAM8),
    .DIN_SRAM9(Tile_X10Y4_DIN_SRAM9),
    .DIN_SRAM10(Tile_X10Y4_DIN_SRAM10),
    .DIN_SRAM11(Tile_X10Y4_DIN_SRAM11),
    .DIN_SRAM12(Tile_X10Y4_DIN_SRAM12),
    .DIN_SRAM13(Tile_X10Y4_DIN_SRAM13),
    .DIN_SRAM14(Tile_X10Y4_DIN_SRAM14),
    .DIN_SRAM15(Tile_X10Y4_DIN_SRAM15),
    .DIN_SRAM16(Tile_X10Y4_DIN_SRAM16),
    .DIN_SRAM17(Tile_X10Y4_DIN_SRAM17),
    .DIN_SRAM18(Tile_X10Y4_DIN_SRAM18),
    .DIN_SRAM19(Tile_X10Y4_DIN_SRAM19),
    .DIN_SRAM20(Tile_X10Y4_DIN_SRAM20),
    .DIN_SRAM21(Tile_X10Y4_DIN_SRAM21),
    .DIN_SRAM22(Tile_X10Y4_DIN_SRAM22),
    .DIN_SRAM23(Tile_X10Y4_DIN_SRAM23),
    .DIN_SRAM24(Tile_X10Y4_DIN_SRAM24),
    .DIN_SRAM25(Tile_X10Y4_DIN_SRAM25),
    .DIN_SRAM26(Tile_X10Y4_DIN_SRAM26),
    .DIN_SRAM27(Tile_X10Y4_DIN_SRAM27),
    .DIN_SRAM28(Tile_X10Y4_DIN_SRAM28),
    .DIN_SRAM29(Tile_X10Y4_DIN_SRAM29),
    .DIN_SRAM30(Tile_X10Y4_DIN_SRAM30),
    .DIN_SRAM31(Tile_X10Y4_DIN_SRAM31),
    .MEN_SRAM(Tile_X10Y4_MEN_SRAM),
    .REN_SRAM(Tile_X10Y4_REN_SRAM),
    .TIE_HIGH_SRAM(Tile_X10Y4_TIE_HIGH_SRAM),
    .TIE_LOW_SRAM(Tile_X10Y4_TIE_LOW_SRAM),
    .WEN_SRAM(Tile_X10Y4_WEN_SRAM),
    .Tile_X0Y0_UserCLKo(Tile_X10Y3_UserCLKo),
    .Tile_X0Y1_UserCLK(Tile_X10Y5_UserCLKo),
    .Tile_X0Y0_FrameData(Tile_X9Y3_FrameData_O),
    .Tile_X0Y0_FrameData_O(Tile_X10Y3_FrameData_O),
    .Tile_X0Y0_FrameStrobe_O(Tile_X10Y3_FrameStrobe_O),
    .Tile_X0Y1_FrameData(Tile_X9Y4_FrameData_O),
    .Tile_X0Y1_FrameData_O(Tile_X10Y4_FrameData_O),
    .Tile_X0Y1_FrameStrobe(Tile_X10Y5_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
W_IO
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X0Y4_Emulate_Bitstream)
    )
`endif
    Tile_X0Y4_W_IO
    (
    .W1END(Tile_X1Y4_W1BEG),
    .W2MID(Tile_X1Y4_W2BEG),
    .W2END(Tile_X1Y4_W2BEGb),
    .WW4END(Tile_X1Y4_WW4BEG),
    .W6END(Tile_X1Y4_W6BEG),
    .E1BEG(Tile_X0Y4_E1BEG),
    .E2BEG(Tile_X0Y4_E2BEG),
    .E2BEGb(Tile_X0Y4_E2BEGb),
    .EE4BEG(Tile_X0Y4_EE4BEG),
    .E6BEG(Tile_X0Y4_E6BEG),
    .A_O_top(Tile_X0Y4_A_O_top),
    .A_I_top(Tile_X0Y4_A_I_top),
    .A_T_top(Tile_X0Y4_A_T_top),
    .B_O_top(Tile_X0Y4_B_O_top),
    .B_I_top(Tile_X0Y4_B_I_top),
    .B_T_top(Tile_X0Y4_B_T_top),
    .A_config_C_bit0(Tile_X0Y4_A_config_C_bit0),
    .A_config_C_bit1(Tile_X0Y4_A_config_C_bit1),
    .A_config_C_bit2(Tile_X0Y4_A_config_C_bit2),
    .A_config_C_bit3(Tile_X0Y4_A_config_C_bit3),
    .B_config_C_bit0(Tile_X0Y4_B_config_C_bit0),
    .B_config_C_bit1(Tile_X0Y4_B_config_C_bit1),
    .B_config_C_bit2(Tile_X0Y4_B_config_C_bit2),
    .B_config_C_bit3(Tile_X0Y4_B_config_C_bit3),
    .UserCLK(Tile_X0Y5_UserCLKo),
    .UserCLKo(Tile_X0Y4_UserCLKo),
    .FrameData(Row_Y4_FrameData),
    .FrameData_O(Tile_X0Y4_FrameData_O),
    .FrameStrobe(Tile_X0Y5_FrameStrobe_O),
    .FrameStrobe_O(Tile_X0Y4_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X1Y4_Emulate_Bitstream)
    )
`endif
    Tile_X1Y4_LUT4AB
    (
    .N1END(Tile_X1Y5_N1BEG),
    .N2MID(Tile_X1Y5_N2BEG),
    .N2END(Tile_X1Y5_N2BEGb),
    .N4END(Tile_X1Y5_N4BEG),
    .NN4END(Tile_X1Y5_NN4BEG),
    .Ci(Tile_X1Y5_Co),
    .E1END(Tile_X0Y4_E1BEG),
    .E2MID(Tile_X0Y4_E2BEG),
    .E2END(Tile_X0Y4_E2BEGb),
    .EE4END(Tile_X0Y4_EE4BEG),
    .E6END(Tile_X0Y4_E6BEG),
    .S1END(Tile_X1Y3_S1BEG),
    .S2MID(Tile_X1Y3_S2BEG),
    .S2END(Tile_X1Y3_S2BEGb),
    .S4END(Tile_X1Y3_S4BEG),
    .SS4END(Tile_X1Y3_SS4BEG),
    .W1END(Tile_X2Y4_W1BEG),
    .W2MID(Tile_X2Y4_W2BEG),
    .W2END(Tile_X2Y4_W2BEGb),
    .WW4END(Tile_X2Y4_WW4BEG),
    .W6END(Tile_X2Y4_W6BEG),
    .N1BEG(Tile_X1Y4_N1BEG),
    .N2BEG(Tile_X1Y4_N2BEG),
    .N2BEGb(Tile_X1Y4_N2BEGb),
    .N4BEG(Tile_X1Y4_N4BEG),
    .NN4BEG(Tile_X1Y4_NN4BEG),
    .E1BEG(Tile_X1Y4_E1BEG),
    .E2BEG(Tile_X1Y4_E2BEG),
    .E2BEGb(Tile_X1Y4_E2BEGb),
    .EE4BEG(Tile_X1Y4_EE4BEG),
    .E6BEG(Tile_X1Y4_E6BEG),
    .S1BEG(Tile_X1Y4_S1BEG),
    .S2BEG(Tile_X1Y4_S2BEG),
    .S2BEGb(Tile_X1Y4_S2BEGb),
    .S4BEG(Tile_X1Y4_S4BEG),
    .SS4BEG(Tile_X1Y4_SS4BEG),
    .W1BEG(Tile_X1Y4_W1BEG),
    .W2BEG(Tile_X1Y4_W2BEG),
    .W2BEGb(Tile_X1Y4_W2BEGb),
    .WW4BEG(Tile_X1Y4_WW4BEG),
    .W6BEG(Tile_X1Y4_W6BEG),
    .Co(Tile_X1Y4_Co),
    .UserCLK(Tile_X1Y5_UserCLKo),
    .UserCLKo(Tile_X1Y4_UserCLKo),
    .FrameData(Tile_X0Y4_FrameData_O),
    .FrameData_O(Tile_X1Y4_FrameData_O),
    .FrameStrobe(Tile_X1Y5_FrameStrobe_O),
    .FrameStrobe_O(Tile_X1Y4_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X2Y4_Emulate_Bitstream)
    )
`endif
    Tile_X2Y4_LUT4AB
    (
    .N1END(Tile_X2Y5_N1BEG),
    .N2MID(Tile_X2Y5_N2BEG),
    .N2END(Tile_X2Y5_N2BEGb),
    .N4END(Tile_X2Y5_N4BEG),
    .NN4END(Tile_X2Y5_NN4BEG),
    .Ci(Tile_X2Y5_Co),
    .E1END(Tile_X1Y4_E1BEG),
    .E2MID(Tile_X1Y4_E2BEG),
    .E2END(Tile_X1Y4_E2BEGb),
    .EE4END(Tile_X1Y4_EE4BEG),
    .E6END(Tile_X1Y4_E6BEG),
    .S1END(Tile_X2Y3_S1BEG),
    .S2MID(Tile_X2Y3_S2BEG),
    .S2END(Tile_X2Y3_S2BEGb),
    .S4END(Tile_X2Y3_S4BEG),
    .SS4END(Tile_X2Y3_SS4BEG),
    .W1END(Tile_X3Y4_W1BEG),
    .W2MID(Tile_X3Y4_W2BEG),
    .W2END(Tile_X3Y4_W2BEGb),
    .WW4END(Tile_X3Y4_WW4BEG),
    .W6END(Tile_X3Y4_W6BEG),
    .N1BEG(Tile_X2Y4_N1BEG),
    .N2BEG(Tile_X2Y4_N2BEG),
    .N2BEGb(Tile_X2Y4_N2BEGb),
    .N4BEG(Tile_X2Y4_N4BEG),
    .NN4BEG(Tile_X2Y4_NN4BEG),
    .E1BEG(Tile_X2Y4_E1BEG),
    .E2BEG(Tile_X2Y4_E2BEG),
    .E2BEGb(Tile_X2Y4_E2BEGb),
    .EE4BEG(Tile_X2Y4_EE4BEG),
    .E6BEG(Tile_X2Y4_E6BEG),
    .S1BEG(Tile_X2Y4_S1BEG),
    .S2BEG(Tile_X2Y4_S2BEG),
    .S2BEGb(Tile_X2Y4_S2BEGb),
    .S4BEG(Tile_X2Y4_S4BEG),
    .SS4BEG(Tile_X2Y4_SS4BEG),
    .W1BEG(Tile_X2Y4_W1BEG),
    .W2BEG(Tile_X2Y4_W2BEG),
    .W2BEGb(Tile_X2Y4_W2BEGb),
    .WW4BEG(Tile_X2Y4_WW4BEG),
    .W6BEG(Tile_X2Y4_W6BEG),
    .Co(Tile_X2Y4_Co),
    .UserCLK(Tile_X2Y5_UserCLKo),
    .UserCLKo(Tile_X2Y4_UserCLKo),
    .FrameData(Tile_X1Y4_FrameData_O),
    .FrameData_O(Tile_X2Y4_FrameData_O),
    .FrameStrobe(Tile_X2Y5_FrameStrobe_O),
    .FrameStrobe_O(Tile_X2Y4_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X3Y4_Emulate_Bitstream)
    )
`endif
    Tile_X3Y4_LUT4AB
    (
    .N1END(Tile_X3Y5_N1BEG),
    .N2MID(Tile_X3Y5_N2BEG),
    .N2END(Tile_X3Y5_N2BEGb),
    .N4END(Tile_X3Y5_N4BEG),
    .NN4END(Tile_X3Y5_NN4BEG),
    .Ci(Tile_X3Y5_Co),
    .E1END(Tile_X2Y4_E1BEG),
    .E2MID(Tile_X2Y4_E2BEG),
    .E2END(Tile_X2Y4_E2BEGb),
    .EE4END(Tile_X2Y4_EE4BEG),
    .E6END(Tile_X2Y4_E6BEG),
    .S1END(Tile_X3Y3_S1BEG),
    .S2MID(Tile_X3Y3_S2BEG),
    .S2END(Tile_X3Y3_S2BEGb),
    .S4END(Tile_X3Y3_S4BEG),
    .SS4END(Tile_X3Y3_SS4BEG),
    .W1END(Tile_X4Y4_W1BEG),
    .W2MID(Tile_X4Y4_W2BEG),
    .W2END(Tile_X4Y4_W2BEGb),
    .WW4END(Tile_X4Y4_WW4BEG),
    .W6END(Tile_X4Y4_W6BEG),
    .N1BEG(Tile_X3Y4_N1BEG),
    .N2BEG(Tile_X3Y4_N2BEG),
    .N2BEGb(Tile_X3Y4_N2BEGb),
    .N4BEG(Tile_X3Y4_N4BEG),
    .NN4BEG(Tile_X3Y4_NN4BEG),
    .E1BEG(Tile_X3Y4_E1BEG),
    .E2BEG(Tile_X3Y4_E2BEG),
    .E2BEGb(Tile_X3Y4_E2BEGb),
    .EE4BEG(Tile_X3Y4_EE4BEG),
    .E6BEG(Tile_X3Y4_E6BEG),
    .S1BEG(Tile_X3Y4_S1BEG),
    .S2BEG(Tile_X3Y4_S2BEG),
    .S2BEGb(Tile_X3Y4_S2BEGb),
    .S4BEG(Tile_X3Y4_S4BEG),
    .SS4BEG(Tile_X3Y4_SS4BEG),
    .W1BEG(Tile_X3Y4_W1BEG),
    .W2BEG(Tile_X3Y4_W2BEG),
    .W2BEGb(Tile_X3Y4_W2BEGb),
    .WW4BEG(Tile_X3Y4_WW4BEG),
    .W6BEG(Tile_X3Y4_W6BEG),
    .Co(Tile_X3Y4_Co),
    .UserCLK(Tile_X3Y5_UserCLKo),
    .UserCLKo(Tile_X3Y4_UserCLKo),
    .FrameData(Tile_X2Y4_FrameData_O),
    .FrameData_O(Tile_X3Y4_FrameData_O),
    .FrameStrobe(Tile_X3Y5_FrameStrobe_O),
    .FrameStrobe_O(Tile_X3Y4_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
RegFile
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X4Y4_Emulate_Bitstream)
    )
`endif
    Tile_X4Y4_RegFile
    (
    .N1END(Tile_X4Y5_N1BEG),
    .N2MID(Tile_X4Y5_N2BEG),
    .N2END(Tile_X4Y5_N2BEGb),
    .N4END(Tile_X4Y5_N4BEG),
    .NN4END(Tile_X4Y5_NN4BEG),
    .E1END(Tile_X3Y4_E1BEG),
    .E2MID(Tile_X3Y4_E2BEG),
    .E2END(Tile_X3Y4_E2BEGb),
    .EE4END(Tile_X3Y4_EE4BEG),
    .E6END(Tile_X3Y4_E6BEG),
    .S1END(Tile_X4Y3_S1BEG),
    .S2MID(Tile_X4Y3_S2BEG),
    .S2END(Tile_X4Y3_S2BEGb),
    .S4END(Tile_X4Y3_S4BEG),
    .SS4END(Tile_X4Y3_SS4BEG),
    .W1END(Tile_X5Y4_W1BEG),
    .W2MID(Tile_X5Y4_W2BEG),
    .W2END(Tile_X5Y4_W2BEGb),
    .WW4END(Tile_X5Y4_WW4BEG),
    .W6END(Tile_X5Y4_W6BEG),
    .N1BEG(Tile_X4Y4_N1BEG),
    .N2BEG(Tile_X4Y4_N2BEG),
    .N2BEGb(Tile_X4Y4_N2BEGb),
    .N4BEG(Tile_X4Y4_N4BEG),
    .NN4BEG(Tile_X4Y4_NN4BEG),
    .E1BEG(Tile_X4Y4_E1BEG),
    .E2BEG(Tile_X4Y4_E2BEG),
    .E2BEGb(Tile_X4Y4_E2BEGb),
    .EE4BEG(Tile_X4Y4_EE4BEG),
    .E6BEG(Tile_X4Y4_E6BEG),
    .S1BEG(Tile_X4Y4_S1BEG),
    .S2BEG(Tile_X4Y4_S2BEG),
    .S2BEGb(Tile_X4Y4_S2BEGb),
    .S4BEG(Tile_X4Y4_S4BEG),
    .SS4BEG(Tile_X4Y4_SS4BEG),
    .W1BEG(Tile_X4Y4_W1BEG),
    .W2BEG(Tile_X4Y4_W2BEG),
    .W2BEGb(Tile_X4Y4_W2BEGb),
    .WW4BEG(Tile_X4Y4_WW4BEG),
    .W6BEG(Tile_X4Y4_W6BEG),
    .UserCLK(Tile_X4Y5_UserCLKo),
    .UserCLKo(Tile_X4Y4_UserCLKo),
    .FrameData(Tile_X3Y4_FrameData_O),
    .FrameData_O(Tile_X4Y4_FrameData_O),
    .FrameStrobe(Tile_X4Y5_FrameStrobe_O),
    .FrameStrobe_O(Tile_X4Y4_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X5Y4_Emulate_Bitstream)
    )
`endif
    Tile_X5Y4_LUT4AB
    (
    .N1END(Tile_X5Y5_N1BEG),
    .N2MID(Tile_X5Y5_N2BEG),
    .N2END(Tile_X5Y5_N2BEGb),
    .N4END(Tile_X5Y5_N4BEG),
    .NN4END(Tile_X5Y5_NN4BEG),
    .Ci(Tile_X5Y5_Co),
    .E1END(Tile_X4Y4_E1BEG),
    .E2MID(Tile_X4Y4_E2BEG),
    .E2END(Tile_X4Y4_E2BEGb),
    .EE4END(Tile_X4Y4_EE4BEG),
    .E6END(Tile_X4Y4_E6BEG),
    .S1END(Tile_X5Y3_S1BEG),
    .S2MID(Tile_X5Y3_S2BEG),
    .S2END(Tile_X5Y3_S2BEGb),
    .S4END(Tile_X5Y3_S4BEG),
    .SS4END(Tile_X5Y3_SS4BEG),
    .W1END(Tile_X6Y4_W1BEG),
    .W2MID(Tile_X6Y4_W2BEG),
    .W2END(Tile_X6Y4_W2BEGb),
    .WW4END(Tile_X6Y4_WW4BEG),
    .W6END(Tile_X6Y4_W6BEG),
    .N1BEG(Tile_X5Y4_N1BEG),
    .N2BEG(Tile_X5Y4_N2BEG),
    .N2BEGb(Tile_X5Y4_N2BEGb),
    .N4BEG(Tile_X5Y4_N4BEG),
    .NN4BEG(Tile_X5Y4_NN4BEG),
    .E1BEG(Tile_X5Y4_E1BEG),
    .E2BEG(Tile_X5Y4_E2BEG),
    .E2BEGb(Tile_X5Y4_E2BEGb),
    .EE4BEG(Tile_X5Y4_EE4BEG),
    .E6BEG(Tile_X5Y4_E6BEG),
    .S1BEG(Tile_X5Y4_S1BEG),
    .S2BEG(Tile_X5Y4_S2BEG),
    .S2BEGb(Tile_X5Y4_S2BEGb),
    .S4BEG(Tile_X5Y4_S4BEG),
    .SS4BEG(Tile_X5Y4_SS4BEG),
    .W1BEG(Tile_X5Y4_W1BEG),
    .W2BEG(Tile_X5Y4_W2BEG),
    .W2BEGb(Tile_X5Y4_W2BEGb),
    .WW4BEG(Tile_X5Y4_WW4BEG),
    .W6BEG(Tile_X5Y4_W6BEG),
    .Co(Tile_X5Y4_Co),
    .UserCLK(Tile_X5Y5_UserCLKo),
    .UserCLKo(Tile_X5Y4_UserCLKo),
    .FrameData(Tile_X4Y4_FrameData_O),
    .FrameData_O(Tile_X5Y4_FrameData_O),
    .FrameStrobe(Tile_X5Y5_FrameStrobe_O),
    .FrameStrobe_O(Tile_X5Y4_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X6Y4_Emulate_Bitstream)
    )
`endif
    Tile_X6Y4_LUT4AB
    (
    .N1END(Tile_X6Y5_N1BEG),
    .N2MID(Tile_X6Y5_N2BEG),
    .N2END(Tile_X6Y5_N2BEGb),
    .N4END(Tile_X6Y5_N4BEG),
    .NN4END(Tile_X6Y5_NN4BEG),
    .Ci(Tile_X6Y5_Co),
    .E1END(Tile_X5Y4_E1BEG),
    .E2MID(Tile_X5Y4_E2BEG),
    .E2END(Tile_X5Y4_E2BEGb),
    .EE4END(Tile_X5Y4_EE4BEG),
    .E6END(Tile_X5Y4_E6BEG),
    .S1END(Tile_X6Y3_S1BEG),
    .S2MID(Tile_X6Y3_S2BEG),
    .S2END(Tile_X6Y3_S2BEGb),
    .S4END(Tile_X6Y3_S4BEG),
    .SS4END(Tile_X6Y3_SS4BEG),
    .W1END(Tile_X7Y4_W1BEG),
    .W2MID(Tile_X7Y4_W2BEG),
    .W2END(Tile_X7Y4_W2BEGb),
    .WW4END(Tile_X7Y4_WW4BEG),
    .W6END(Tile_X7Y4_W6BEG),
    .N1BEG(Tile_X6Y4_N1BEG),
    .N2BEG(Tile_X6Y4_N2BEG),
    .N2BEGb(Tile_X6Y4_N2BEGb),
    .N4BEG(Tile_X6Y4_N4BEG),
    .NN4BEG(Tile_X6Y4_NN4BEG),
    .E1BEG(Tile_X6Y4_E1BEG),
    .E2BEG(Tile_X6Y4_E2BEG),
    .E2BEGb(Tile_X6Y4_E2BEGb),
    .EE4BEG(Tile_X6Y4_EE4BEG),
    .E6BEG(Tile_X6Y4_E6BEG),
    .S1BEG(Tile_X6Y4_S1BEG),
    .S2BEG(Tile_X6Y4_S2BEG),
    .S2BEGb(Tile_X6Y4_S2BEGb),
    .S4BEG(Tile_X6Y4_S4BEG),
    .SS4BEG(Tile_X6Y4_SS4BEG),
    .W1BEG(Tile_X6Y4_W1BEG),
    .W2BEG(Tile_X6Y4_W2BEG),
    .W2BEGb(Tile_X6Y4_W2BEGb),
    .WW4BEG(Tile_X6Y4_WW4BEG),
    .W6BEG(Tile_X6Y4_W6BEG),
    .Co(Tile_X6Y4_Co),
    .UserCLK(Tile_X6Y5_UserCLKo),
    .UserCLKo(Tile_X6Y4_UserCLKo),
    .FrameData(Tile_X5Y4_FrameData_O),
    .FrameData_O(Tile_X6Y4_FrameData_O),
    .FrameStrobe(Tile_X6Y5_FrameStrobe_O),
    .FrameStrobe_O(Tile_X6Y4_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X8Y4_Emulate_Bitstream)
    )
`endif
    Tile_X8Y4_LUT4AB
    (
    .N1END(Tile_X8Y5_N1BEG),
    .N2MID(Tile_X8Y5_N2BEG),
    .N2END(Tile_X8Y5_N2BEGb),
    .N4END(Tile_X8Y5_N4BEG),
    .NN4END(Tile_X8Y5_NN4BEG),
    .Ci(Tile_X8Y5_Co),
    .E1END(Tile_X7Y4_E1BEG),
    .E2MID(Tile_X7Y4_E2BEG),
    .E2END(Tile_X7Y4_E2BEGb),
    .EE4END(Tile_X7Y4_EE4BEG),
    .E6END(Tile_X7Y4_E6BEG),
    .S1END(Tile_X8Y3_S1BEG),
    .S2MID(Tile_X8Y3_S2BEG),
    .S2END(Tile_X8Y3_S2BEGb),
    .S4END(Tile_X8Y3_S4BEG),
    .SS4END(Tile_X8Y3_SS4BEG),
    .W1END(Tile_X9Y4_W1BEG),
    .W2MID(Tile_X9Y4_W2BEG),
    .W2END(Tile_X9Y4_W2BEGb),
    .WW4END(Tile_X9Y4_WW4BEG),
    .W6END(Tile_X9Y4_W6BEG),
    .N1BEG(Tile_X8Y4_N1BEG),
    .N2BEG(Tile_X8Y4_N2BEG),
    .N2BEGb(Tile_X8Y4_N2BEGb),
    .N4BEG(Tile_X8Y4_N4BEG),
    .NN4BEG(Tile_X8Y4_NN4BEG),
    .E1BEG(Tile_X8Y4_E1BEG),
    .E2BEG(Tile_X8Y4_E2BEG),
    .E2BEGb(Tile_X8Y4_E2BEGb),
    .EE4BEG(Tile_X8Y4_EE4BEG),
    .E6BEG(Tile_X8Y4_E6BEG),
    .S1BEG(Tile_X8Y4_S1BEG),
    .S2BEG(Tile_X8Y4_S2BEG),
    .S2BEGb(Tile_X8Y4_S2BEGb),
    .S4BEG(Tile_X8Y4_S4BEG),
    .SS4BEG(Tile_X8Y4_SS4BEG),
    .W1BEG(Tile_X8Y4_W1BEG),
    .W2BEG(Tile_X8Y4_W2BEG),
    .W2BEGb(Tile_X8Y4_W2BEGb),
    .WW4BEG(Tile_X8Y4_WW4BEG),
    .W6BEG(Tile_X8Y4_W6BEG),
    .Co(Tile_X8Y4_Co),
    .UserCLK(Tile_X8Y5_UserCLKo),
    .UserCLKo(Tile_X8Y4_UserCLKo),
    .FrameData(Tile_X7Y4_FrameData_O),
    .FrameData_O(Tile_X8Y4_FrameData_O),
    .FrameStrobe(Tile_X8Y5_FrameStrobe_O),
    .FrameStrobe_O(Tile_X8Y4_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X9Y4_Emulate_Bitstream)
    )
`endif
    Tile_X9Y4_LUT4AB
    (
    .N1END(Tile_X9Y5_N1BEG),
    .N2MID(Tile_X9Y5_N2BEG),
    .N2END(Tile_X9Y5_N2BEGb),
    .N4END(Tile_X9Y5_N4BEG),
    .NN4END(Tile_X9Y5_NN4BEG),
    .Ci(Tile_X9Y5_Co),
    .E1END(Tile_X8Y4_E1BEG),
    .E2MID(Tile_X8Y4_E2BEG),
    .E2END(Tile_X8Y4_E2BEGb),
    .EE4END(Tile_X8Y4_EE4BEG),
    .E6END(Tile_X8Y4_E6BEG),
    .S1END(Tile_X9Y3_S1BEG),
    .S2MID(Tile_X9Y3_S2BEG),
    .S2END(Tile_X9Y3_S2BEGb),
    .S4END(Tile_X9Y3_S4BEG),
    .SS4END(Tile_X9Y3_SS4BEG),
    .W1END(Tile_X10Y4_W1BEG),
    .W2MID(Tile_X10Y4_W2BEG),
    .W2END(Tile_X10Y4_W2BEGb),
    .WW4END(Tile_X10Y4_WW4BEG),
    .W6END(Tile_X10Y4_W6BEG),
    .N1BEG(Tile_X9Y4_N1BEG),
    .N2BEG(Tile_X9Y4_N2BEG),
    .N2BEGb(Tile_X9Y4_N2BEGb),
    .N4BEG(Tile_X9Y4_N4BEG),
    .NN4BEG(Tile_X9Y4_NN4BEG),
    .E1BEG(Tile_X9Y4_E1BEG),
    .E2BEG(Tile_X9Y4_E2BEG),
    .E2BEGb(Tile_X9Y4_E2BEGb),
    .EE4BEG(Tile_X9Y4_EE4BEG),
    .E6BEG(Tile_X9Y4_E6BEG),
    .S1BEG(Tile_X9Y4_S1BEG),
    .S2BEG(Tile_X9Y4_S2BEG),
    .S2BEGb(Tile_X9Y4_S2BEGb),
    .S4BEG(Tile_X9Y4_S4BEG),
    .SS4BEG(Tile_X9Y4_SS4BEG),
    .W1BEG(Tile_X9Y4_W1BEG),
    .W2BEG(Tile_X9Y4_W2BEG),
    .W2BEGb(Tile_X9Y4_W2BEGb),
    .WW4BEG(Tile_X9Y4_WW4BEG),
    .W6BEG(Tile_X9Y4_W6BEG),
    .Co(Tile_X9Y4_Co),
    .UserCLK(Tile_X9Y5_UserCLKo),
    .UserCLKo(Tile_X9Y4_UserCLKo),
    .FrameData(Tile_X8Y4_FrameData_O),
    .FrameData_O(Tile_X9Y4_FrameData_O),
    .FrameStrobe(Tile_X9Y5_FrameStrobe_O),
    .FrameStrobe_O(Tile_X9Y4_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
W_IO
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X0Y5_Emulate_Bitstream)
    )
`endif
    Tile_X0Y5_W_IO
    (
    .W1END(Tile_X1Y5_W1BEG),
    .W2MID(Tile_X1Y5_W2BEG),
    .W2END(Tile_X1Y5_W2BEGb),
    .WW4END(Tile_X1Y5_WW4BEG),
    .W6END(Tile_X1Y5_W6BEG),
    .E1BEG(Tile_X0Y5_E1BEG),
    .E2BEG(Tile_X0Y5_E2BEG),
    .E2BEGb(Tile_X0Y5_E2BEGb),
    .EE4BEG(Tile_X0Y5_EE4BEG),
    .E6BEG(Tile_X0Y5_E6BEG),
    .A_O_top(Tile_X0Y5_A_O_top),
    .A_I_top(Tile_X0Y5_A_I_top),
    .A_T_top(Tile_X0Y5_A_T_top),
    .B_O_top(Tile_X0Y5_B_O_top),
    .B_I_top(Tile_X0Y5_B_I_top),
    .B_T_top(Tile_X0Y5_B_T_top),
    .A_config_C_bit0(Tile_X0Y5_A_config_C_bit0),
    .A_config_C_bit1(Tile_X0Y5_A_config_C_bit1),
    .A_config_C_bit2(Tile_X0Y5_A_config_C_bit2),
    .A_config_C_bit3(Tile_X0Y5_A_config_C_bit3),
    .B_config_C_bit0(Tile_X0Y5_B_config_C_bit0),
    .B_config_C_bit1(Tile_X0Y5_B_config_C_bit1),
    .B_config_C_bit2(Tile_X0Y5_B_config_C_bit2),
    .B_config_C_bit3(Tile_X0Y5_B_config_C_bit3),
    .UserCLK(Tile_X0Y6_UserCLKo),
    .UserCLKo(Tile_X0Y5_UserCLKo),
    .FrameData(Row_Y5_FrameData),
    .FrameData_O(Tile_X0Y5_FrameData_O),
    .FrameStrobe(Tile_X0Y6_FrameStrobe_O),
    .FrameStrobe_O(Tile_X0Y5_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X1Y5_Emulate_Bitstream)
    )
`endif
    Tile_X1Y5_LUT4AB
    (
    .N1END(Tile_X1Y6_N1BEG),
    .N2MID(Tile_X1Y6_N2BEG),
    .N2END(Tile_X1Y6_N2BEGb),
    .N4END(Tile_X1Y6_N4BEG),
    .NN4END(Tile_X1Y6_NN4BEG),
    .Ci(Tile_X1Y6_Co),
    .E1END(Tile_X0Y5_E1BEG),
    .E2MID(Tile_X0Y5_E2BEG),
    .E2END(Tile_X0Y5_E2BEGb),
    .EE4END(Tile_X0Y5_EE4BEG),
    .E6END(Tile_X0Y5_E6BEG),
    .S1END(Tile_X1Y4_S1BEG),
    .S2MID(Tile_X1Y4_S2BEG),
    .S2END(Tile_X1Y4_S2BEGb),
    .S4END(Tile_X1Y4_S4BEG),
    .SS4END(Tile_X1Y4_SS4BEG),
    .W1END(Tile_X2Y5_W1BEG),
    .W2MID(Tile_X2Y5_W2BEG),
    .W2END(Tile_X2Y5_W2BEGb),
    .WW4END(Tile_X2Y5_WW4BEG),
    .W6END(Tile_X2Y5_W6BEG),
    .N1BEG(Tile_X1Y5_N1BEG),
    .N2BEG(Tile_X1Y5_N2BEG),
    .N2BEGb(Tile_X1Y5_N2BEGb),
    .N4BEG(Tile_X1Y5_N4BEG),
    .NN4BEG(Tile_X1Y5_NN4BEG),
    .E1BEG(Tile_X1Y5_E1BEG),
    .E2BEG(Tile_X1Y5_E2BEG),
    .E2BEGb(Tile_X1Y5_E2BEGb),
    .EE4BEG(Tile_X1Y5_EE4BEG),
    .E6BEG(Tile_X1Y5_E6BEG),
    .S1BEG(Tile_X1Y5_S1BEG),
    .S2BEG(Tile_X1Y5_S2BEG),
    .S2BEGb(Tile_X1Y5_S2BEGb),
    .S4BEG(Tile_X1Y5_S4BEG),
    .SS4BEG(Tile_X1Y5_SS4BEG),
    .W1BEG(Tile_X1Y5_W1BEG),
    .W2BEG(Tile_X1Y5_W2BEG),
    .W2BEGb(Tile_X1Y5_W2BEGb),
    .WW4BEG(Tile_X1Y5_WW4BEG),
    .W6BEG(Tile_X1Y5_W6BEG),
    .Co(Tile_X1Y5_Co),
    .UserCLK(Tile_X1Y6_UserCLKo),
    .UserCLKo(Tile_X1Y5_UserCLKo),
    .FrameData(Tile_X0Y5_FrameData_O),
    .FrameData_O(Tile_X1Y5_FrameData_O),
    .FrameStrobe(Tile_X1Y6_FrameStrobe_O),
    .FrameStrobe_O(Tile_X1Y5_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X2Y5_Emulate_Bitstream)
    )
`endif
    Tile_X2Y5_LUT4AB
    (
    .N1END(Tile_X2Y6_N1BEG),
    .N2MID(Tile_X2Y6_N2BEG),
    .N2END(Tile_X2Y6_N2BEGb),
    .N4END(Tile_X2Y6_N4BEG),
    .NN4END(Tile_X2Y6_NN4BEG),
    .Ci(Tile_X2Y6_Co),
    .E1END(Tile_X1Y5_E1BEG),
    .E2MID(Tile_X1Y5_E2BEG),
    .E2END(Tile_X1Y5_E2BEGb),
    .EE4END(Tile_X1Y5_EE4BEG),
    .E6END(Tile_X1Y5_E6BEG),
    .S1END(Tile_X2Y4_S1BEG),
    .S2MID(Tile_X2Y4_S2BEG),
    .S2END(Tile_X2Y4_S2BEGb),
    .S4END(Tile_X2Y4_S4BEG),
    .SS4END(Tile_X2Y4_SS4BEG),
    .W1END(Tile_X3Y5_W1BEG),
    .W2MID(Tile_X3Y5_W2BEG),
    .W2END(Tile_X3Y5_W2BEGb),
    .WW4END(Tile_X3Y5_WW4BEG),
    .W6END(Tile_X3Y5_W6BEG),
    .N1BEG(Tile_X2Y5_N1BEG),
    .N2BEG(Tile_X2Y5_N2BEG),
    .N2BEGb(Tile_X2Y5_N2BEGb),
    .N4BEG(Tile_X2Y5_N4BEG),
    .NN4BEG(Tile_X2Y5_NN4BEG),
    .E1BEG(Tile_X2Y5_E1BEG),
    .E2BEG(Tile_X2Y5_E2BEG),
    .E2BEGb(Tile_X2Y5_E2BEGb),
    .EE4BEG(Tile_X2Y5_EE4BEG),
    .E6BEG(Tile_X2Y5_E6BEG),
    .S1BEG(Tile_X2Y5_S1BEG),
    .S2BEG(Tile_X2Y5_S2BEG),
    .S2BEGb(Tile_X2Y5_S2BEGb),
    .S4BEG(Tile_X2Y5_S4BEG),
    .SS4BEG(Tile_X2Y5_SS4BEG),
    .W1BEG(Tile_X2Y5_W1BEG),
    .W2BEG(Tile_X2Y5_W2BEG),
    .W2BEGb(Tile_X2Y5_W2BEGb),
    .WW4BEG(Tile_X2Y5_WW4BEG),
    .W6BEG(Tile_X2Y5_W6BEG),
    .Co(Tile_X2Y5_Co),
    .UserCLK(Tile_X2Y6_UserCLKo),
    .UserCLKo(Tile_X2Y5_UserCLKo),
    .FrameData(Tile_X1Y5_FrameData_O),
    .FrameData_O(Tile_X2Y5_FrameData_O),
    .FrameStrobe(Tile_X2Y6_FrameStrobe_O),
    .FrameStrobe_O(Tile_X2Y5_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X3Y5_Emulate_Bitstream)
    )
`endif
    Tile_X3Y5_LUT4AB
    (
    .N1END(Tile_X3Y6_N1BEG),
    .N2MID(Tile_X3Y6_N2BEG),
    .N2END(Tile_X3Y6_N2BEGb),
    .N4END(Tile_X3Y6_N4BEG),
    .NN4END(Tile_X3Y6_NN4BEG),
    .Ci(Tile_X3Y6_Co),
    .E1END(Tile_X2Y5_E1BEG),
    .E2MID(Tile_X2Y5_E2BEG),
    .E2END(Tile_X2Y5_E2BEGb),
    .EE4END(Tile_X2Y5_EE4BEG),
    .E6END(Tile_X2Y5_E6BEG),
    .S1END(Tile_X3Y4_S1BEG),
    .S2MID(Tile_X3Y4_S2BEG),
    .S2END(Tile_X3Y4_S2BEGb),
    .S4END(Tile_X3Y4_S4BEG),
    .SS4END(Tile_X3Y4_SS4BEG),
    .W1END(Tile_X4Y5_W1BEG),
    .W2MID(Tile_X4Y5_W2BEG),
    .W2END(Tile_X4Y5_W2BEGb),
    .WW4END(Tile_X4Y5_WW4BEG),
    .W6END(Tile_X4Y5_W6BEG),
    .N1BEG(Tile_X3Y5_N1BEG),
    .N2BEG(Tile_X3Y5_N2BEG),
    .N2BEGb(Tile_X3Y5_N2BEGb),
    .N4BEG(Tile_X3Y5_N4BEG),
    .NN4BEG(Tile_X3Y5_NN4BEG),
    .E1BEG(Tile_X3Y5_E1BEG),
    .E2BEG(Tile_X3Y5_E2BEG),
    .E2BEGb(Tile_X3Y5_E2BEGb),
    .EE4BEG(Tile_X3Y5_EE4BEG),
    .E6BEG(Tile_X3Y5_E6BEG),
    .S1BEG(Tile_X3Y5_S1BEG),
    .S2BEG(Tile_X3Y5_S2BEG),
    .S2BEGb(Tile_X3Y5_S2BEGb),
    .S4BEG(Tile_X3Y5_S4BEG),
    .SS4BEG(Tile_X3Y5_SS4BEG),
    .W1BEG(Tile_X3Y5_W1BEG),
    .W2BEG(Tile_X3Y5_W2BEG),
    .W2BEGb(Tile_X3Y5_W2BEGb),
    .WW4BEG(Tile_X3Y5_WW4BEG),
    .W6BEG(Tile_X3Y5_W6BEG),
    .Co(Tile_X3Y5_Co),
    .UserCLK(Tile_X3Y6_UserCLKo),
    .UserCLKo(Tile_X3Y5_UserCLKo),
    .FrameData(Tile_X2Y5_FrameData_O),
    .FrameData_O(Tile_X3Y5_FrameData_O),
    .FrameStrobe(Tile_X3Y6_FrameStrobe_O),
    .FrameStrobe_O(Tile_X3Y5_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
RegFile
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X4Y5_Emulate_Bitstream)
    )
`endif
    Tile_X4Y5_RegFile
    (
    .N1END(Tile_X4Y6_N1BEG),
    .N2MID(Tile_X4Y6_N2BEG),
    .N2END(Tile_X4Y6_N2BEGb),
    .N4END(Tile_X4Y6_N4BEG),
    .NN4END(Tile_X4Y6_NN4BEG),
    .E1END(Tile_X3Y5_E1BEG),
    .E2MID(Tile_X3Y5_E2BEG),
    .E2END(Tile_X3Y5_E2BEGb),
    .EE4END(Tile_X3Y5_EE4BEG),
    .E6END(Tile_X3Y5_E6BEG),
    .S1END(Tile_X4Y4_S1BEG),
    .S2MID(Tile_X4Y4_S2BEG),
    .S2END(Tile_X4Y4_S2BEGb),
    .S4END(Tile_X4Y4_S4BEG),
    .SS4END(Tile_X4Y4_SS4BEG),
    .W1END(Tile_X5Y5_W1BEG),
    .W2MID(Tile_X5Y5_W2BEG),
    .W2END(Tile_X5Y5_W2BEGb),
    .WW4END(Tile_X5Y5_WW4BEG),
    .W6END(Tile_X5Y5_W6BEG),
    .N1BEG(Tile_X4Y5_N1BEG),
    .N2BEG(Tile_X4Y5_N2BEG),
    .N2BEGb(Tile_X4Y5_N2BEGb),
    .N4BEG(Tile_X4Y5_N4BEG),
    .NN4BEG(Tile_X4Y5_NN4BEG),
    .E1BEG(Tile_X4Y5_E1BEG),
    .E2BEG(Tile_X4Y5_E2BEG),
    .E2BEGb(Tile_X4Y5_E2BEGb),
    .EE4BEG(Tile_X4Y5_EE4BEG),
    .E6BEG(Tile_X4Y5_E6BEG),
    .S1BEG(Tile_X4Y5_S1BEG),
    .S2BEG(Tile_X4Y5_S2BEG),
    .S2BEGb(Tile_X4Y5_S2BEGb),
    .S4BEG(Tile_X4Y5_S4BEG),
    .SS4BEG(Tile_X4Y5_SS4BEG),
    .W1BEG(Tile_X4Y5_W1BEG),
    .W2BEG(Tile_X4Y5_W2BEG),
    .W2BEGb(Tile_X4Y5_W2BEGb),
    .WW4BEG(Tile_X4Y5_WW4BEG),
    .W6BEG(Tile_X4Y5_W6BEG),
    .UserCLK(Tile_X4Y6_UserCLKo),
    .UserCLKo(Tile_X4Y5_UserCLKo),
    .FrameData(Tile_X3Y5_FrameData_O),
    .FrameData_O(Tile_X4Y5_FrameData_O),
    .FrameStrobe(Tile_X4Y6_FrameStrobe_O),
    .FrameStrobe_O(Tile_X4Y5_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X5Y5_Emulate_Bitstream)
    )
`endif
    Tile_X5Y5_LUT4AB
    (
    .N1END(Tile_X5Y6_N1BEG),
    .N2MID(Tile_X5Y6_N2BEG),
    .N2END(Tile_X5Y6_N2BEGb),
    .N4END(Tile_X5Y6_N4BEG),
    .NN4END(Tile_X5Y6_NN4BEG),
    .Ci(Tile_X5Y6_Co),
    .E1END(Tile_X4Y5_E1BEG),
    .E2MID(Tile_X4Y5_E2BEG),
    .E2END(Tile_X4Y5_E2BEGb),
    .EE4END(Tile_X4Y5_EE4BEG),
    .E6END(Tile_X4Y5_E6BEG),
    .S1END(Tile_X5Y4_S1BEG),
    .S2MID(Tile_X5Y4_S2BEG),
    .S2END(Tile_X5Y4_S2BEGb),
    .S4END(Tile_X5Y4_S4BEG),
    .SS4END(Tile_X5Y4_SS4BEG),
    .W1END(Tile_X6Y5_W1BEG),
    .W2MID(Tile_X6Y5_W2BEG),
    .W2END(Tile_X6Y5_W2BEGb),
    .WW4END(Tile_X6Y5_WW4BEG),
    .W6END(Tile_X6Y5_W6BEG),
    .N1BEG(Tile_X5Y5_N1BEG),
    .N2BEG(Tile_X5Y5_N2BEG),
    .N2BEGb(Tile_X5Y5_N2BEGb),
    .N4BEG(Tile_X5Y5_N4BEG),
    .NN4BEG(Tile_X5Y5_NN4BEG),
    .E1BEG(Tile_X5Y5_E1BEG),
    .E2BEG(Tile_X5Y5_E2BEG),
    .E2BEGb(Tile_X5Y5_E2BEGb),
    .EE4BEG(Tile_X5Y5_EE4BEG),
    .E6BEG(Tile_X5Y5_E6BEG),
    .S1BEG(Tile_X5Y5_S1BEG),
    .S2BEG(Tile_X5Y5_S2BEG),
    .S2BEGb(Tile_X5Y5_S2BEGb),
    .S4BEG(Tile_X5Y5_S4BEG),
    .SS4BEG(Tile_X5Y5_SS4BEG),
    .W1BEG(Tile_X5Y5_W1BEG),
    .W2BEG(Tile_X5Y5_W2BEG),
    .W2BEGb(Tile_X5Y5_W2BEGb),
    .WW4BEG(Tile_X5Y5_WW4BEG),
    .W6BEG(Tile_X5Y5_W6BEG),
    .Co(Tile_X5Y5_Co),
    .UserCLK(Tile_X5Y6_UserCLKo),
    .UserCLKo(Tile_X5Y5_UserCLKo),
    .FrameData(Tile_X4Y5_FrameData_O),
    .FrameData_O(Tile_X5Y5_FrameData_O),
    .FrameStrobe(Tile_X5Y6_FrameStrobe_O),
    .FrameStrobe_O(Tile_X5Y5_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X6Y5_Emulate_Bitstream)
    )
`endif
    Tile_X6Y5_LUT4AB
    (
    .N1END(Tile_X6Y6_N1BEG),
    .N2MID(Tile_X6Y6_N2BEG),
    .N2END(Tile_X6Y6_N2BEGb),
    .N4END(Tile_X6Y6_N4BEG),
    .NN4END(Tile_X6Y6_NN4BEG),
    .Ci(Tile_X6Y6_Co),
    .E1END(Tile_X5Y5_E1BEG),
    .E2MID(Tile_X5Y5_E2BEG),
    .E2END(Tile_X5Y5_E2BEGb),
    .EE4END(Tile_X5Y5_EE4BEG),
    .E6END(Tile_X5Y5_E6BEG),
    .S1END(Tile_X6Y4_S1BEG),
    .S2MID(Tile_X6Y4_S2BEG),
    .S2END(Tile_X6Y4_S2BEGb),
    .S4END(Tile_X6Y4_S4BEG),
    .SS4END(Tile_X6Y4_SS4BEG),
    .W1END(Tile_X7Y5_W1BEG),
    .W2MID(Tile_X7Y5_W2BEG),
    .W2END(Tile_X7Y5_W2BEGb),
    .WW4END(Tile_X7Y5_WW4BEG),
    .W6END(Tile_X7Y5_W6BEG),
    .N1BEG(Tile_X6Y5_N1BEG),
    .N2BEG(Tile_X6Y5_N2BEG),
    .N2BEGb(Tile_X6Y5_N2BEGb),
    .N4BEG(Tile_X6Y5_N4BEG),
    .NN4BEG(Tile_X6Y5_NN4BEG),
    .E1BEG(Tile_X6Y5_E1BEG),
    .E2BEG(Tile_X6Y5_E2BEG),
    .E2BEGb(Tile_X6Y5_E2BEGb),
    .EE4BEG(Tile_X6Y5_EE4BEG),
    .E6BEG(Tile_X6Y5_E6BEG),
    .S1BEG(Tile_X6Y5_S1BEG),
    .S2BEG(Tile_X6Y5_S2BEG),
    .S2BEGb(Tile_X6Y5_S2BEGb),
    .S4BEG(Tile_X6Y5_S4BEG),
    .SS4BEG(Tile_X6Y5_SS4BEG),
    .W1BEG(Tile_X6Y5_W1BEG),
    .W2BEG(Tile_X6Y5_W2BEG),
    .W2BEGb(Tile_X6Y5_W2BEGb),
    .WW4BEG(Tile_X6Y5_WW4BEG),
    .W6BEG(Tile_X6Y5_W6BEG),
    .Co(Tile_X6Y5_Co),
    .UserCLK(Tile_X6Y6_UserCLKo),
    .UserCLKo(Tile_X6Y5_UserCLKo),
    .FrameData(Tile_X5Y5_FrameData_O),
    .FrameData_O(Tile_X6Y5_FrameData_O),
    .FrameStrobe(Tile_X6Y6_FrameStrobe_O),
    .FrameStrobe_O(Tile_X6Y5_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
DSP
`ifdef EMULATION
    #(
    .Tile_X0Y0_Emulate_Bitstream(`Tile_X7Y5_Emulate_Bitstream),
    .Tile_X0Y1_Emulate_Bitstream(`Tile_X7Y6_Emulate_Bitstream)
    )
`endif
    Tile_X7Y5_DSP
    (
    .Tile_X0Y0_E1END(Tile_X6Y5_E1BEG),
    .Tile_X0Y0_E2MID(Tile_X6Y5_E2BEG),
    .Tile_X0Y0_E2END(Tile_X6Y5_E2BEGb),
    .Tile_X0Y0_EE4END(Tile_X6Y5_EE4BEG),
    .Tile_X0Y0_E6END(Tile_X6Y5_E6BEG),
    .Tile_X0Y0_S1END(Tile_X7Y4_S1BEG),
    .Tile_X0Y0_S2MID(Tile_X7Y4_S2BEG),
    .Tile_X0Y0_S2END(Tile_X7Y4_S2BEGb),
    .Tile_X0Y0_S4END(Tile_X7Y4_S4BEG),
    .Tile_X0Y0_SS4END(Tile_X7Y4_SS4BEG),
    .Tile_X0Y0_W1END(Tile_X8Y5_W1BEG),
    .Tile_X0Y0_W2MID(Tile_X8Y5_W2BEG),
    .Tile_X0Y0_W2END(Tile_X8Y5_W2BEGb),
    .Tile_X0Y0_WW4END(Tile_X8Y5_WW4BEG),
    .Tile_X0Y0_W6END(Tile_X8Y5_W6BEG),
    .Tile_X0Y1_N1END(Tile_X7Y7_N1BEG),
    .Tile_X0Y1_N2MID(Tile_X7Y7_N2BEG),
    .Tile_X0Y1_N2END(Tile_X7Y7_N2BEGb),
    .Tile_X0Y1_N4END(Tile_X7Y7_N4BEG),
    .Tile_X0Y1_NN4END(Tile_X7Y7_NN4BEG),
    .Tile_X0Y1_E1END(Tile_X6Y6_E1BEG),
    .Tile_X0Y1_E2MID(Tile_X6Y6_E2BEG),
    .Tile_X0Y1_E2END(Tile_X6Y6_E2BEGb),
    .Tile_X0Y1_EE4END(Tile_X6Y6_EE4BEG),
    .Tile_X0Y1_E6END(Tile_X6Y6_E6BEG),
    .Tile_X0Y1_W1END(Tile_X8Y6_W1BEG),
    .Tile_X0Y1_W2MID(Tile_X8Y6_W2BEG),
    .Tile_X0Y1_W2END(Tile_X8Y6_W2BEGb),
    .Tile_X0Y1_WW4END(Tile_X8Y6_WW4BEG),
    .Tile_X0Y1_W6END(Tile_X8Y6_W6BEG),
    .Tile_X0Y0_N1BEG(Tile_X7Y5_N1BEG),
    .Tile_X0Y0_N2BEG(Tile_X7Y5_N2BEG),
    .Tile_X0Y0_N2BEGb(Tile_X7Y5_N2BEGb),
    .Tile_X0Y0_N4BEG(Tile_X7Y5_N4BEG),
    .Tile_X0Y0_NN4BEG(Tile_X7Y5_NN4BEG),
    .Tile_X0Y0_E1BEG(Tile_X7Y5_E1BEG),
    .Tile_X0Y0_E2BEG(Tile_X7Y5_E2BEG),
    .Tile_X0Y0_E2BEGb(Tile_X7Y5_E2BEGb),
    .Tile_X0Y0_EE4BEG(Tile_X7Y5_EE4BEG),
    .Tile_X0Y0_E6BEG(Tile_X7Y5_E6BEG),
    .Tile_X0Y0_W1BEG(Tile_X7Y5_W1BEG),
    .Tile_X0Y0_W2BEG(Tile_X7Y5_W2BEG),
    .Tile_X0Y0_W2BEGb(Tile_X7Y5_W2BEGb),
    .Tile_X0Y0_WW4BEG(Tile_X7Y5_WW4BEG),
    .Tile_X0Y0_W6BEG(Tile_X7Y5_W6BEG),
    .Tile_X0Y1_E1BEG(Tile_X7Y6_E1BEG),
    .Tile_X0Y1_E2BEG(Tile_X7Y6_E2BEG),
    .Tile_X0Y1_E2BEGb(Tile_X7Y6_E2BEGb),
    .Tile_X0Y1_EE4BEG(Tile_X7Y6_EE4BEG),
    .Tile_X0Y1_E6BEG(Tile_X7Y6_E6BEG),
    .Tile_X0Y1_S1BEG(Tile_X7Y6_S1BEG),
    .Tile_X0Y1_S2BEG(Tile_X7Y6_S2BEG),
    .Tile_X0Y1_S2BEGb(Tile_X7Y6_S2BEGb),
    .Tile_X0Y1_S4BEG(Tile_X7Y6_S4BEG),
    .Tile_X0Y1_SS4BEG(Tile_X7Y6_SS4BEG),
    .Tile_X0Y1_W1BEG(Tile_X7Y6_W1BEG),
    .Tile_X0Y1_W2BEG(Tile_X7Y6_W2BEG),
    .Tile_X0Y1_W2BEGb(Tile_X7Y6_W2BEGb),
    .Tile_X0Y1_WW4BEG(Tile_X7Y6_WW4BEG),
    .Tile_X0Y1_W6BEG(Tile_X7Y6_W6BEG),
    .Tile_X0Y0_UserCLKo(Tile_X7Y5_UserCLKo),
    .Tile_X0Y1_UserCLK(Tile_X7Y7_UserCLKo),
    .Tile_X0Y0_FrameData(Tile_X6Y5_FrameData_O),
    .Tile_X0Y0_FrameData_O(Tile_X7Y5_FrameData_O),
    .Tile_X0Y0_FrameStrobe_O(Tile_X7Y5_FrameStrobe_O),
    .Tile_X0Y1_FrameData(Tile_X6Y6_FrameData_O),
    .Tile_X0Y1_FrameData_O(Tile_X7Y6_FrameData_O),
    .Tile_X0Y1_FrameStrobe(Tile_X7Y7_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X8Y5_Emulate_Bitstream)
    )
`endif
    Tile_X8Y5_LUT4AB
    (
    .N1END(Tile_X8Y6_N1BEG),
    .N2MID(Tile_X8Y6_N2BEG),
    .N2END(Tile_X8Y6_N2BEGb),
    .N4END(Tile_X8Y6_N4BEG),
    .NN4END(Tile_X8Y6_NN4BEG),
    .Ci(Tile_X8Y6_Co),
    .E1END(Tile_X7Y5_E1BEG),
    .E2MID(Tile_X7Y5_E2BEG),
    .E2END(Tile_X7Y5_E2BEGb),
    .EE4END(Tile_X7Y5_EE4BEG),
    .E6END(Tile_X7Y5_E6BEG),
    .S1END(Tile_X8Y4_S1BEG),
    .S2MID(Tile_X8Y4_S2BEG),
    .S2END(Tile_X8Y4_S2BEGb),
    .S4END(Tile_X8Y4_S4BEG),
    .SS4END(Tile_X8Y4_SS4BEG),
    .W1END(Tile_X9Y5_W1BEG),
    .W2MID(Tile_X9Y5_W2BEG),
    .W2END(Tile_X9Y5_W2BEGb),
    .WW4END(Tile_X9Y5_WW4BEG),
    .W6END(Tile_X9Y5_W6BEG),
    .N1BEG(Tile_X8Y5_N1BEG),
    .N2BEG(Tile_X8Y5_N2BEG),
    .N2BEGb(Tile_X8Y5_N2BEGb),
    .N4BEG(Tile_X8Y5_N4BEG),
    .NN4BEG(Tile_X8Y5_NN4BEG),
    .E1BEG(Tile_X8Y5_E1BEG),
    .E2BEG(Tile_X8Y5_E2BEG),
    .E2BEGb(Tile_X8Y5_E2BEGb),
    .EE4BEG(Tile_X8Y5_EE4BEG),
    .E6BEG(Tile_X8Y5_E6BEG),
    .S1BEG(Tile_X8Y5_S1BEG),
    .S2BEG(Tile_X8Y5_S2BEG),
    .S2BEGb(Tile_X8Y5_S2BEGb),
    .S4BEG(Tile_X8Y5_S4BEG),
    .SS4BEG(Tile_X8Y5_SS4BEG),
    .W1BEG(Tile_X8Y5_W1BEG),
    .W2BEG(Tile_X8Y5_W2BEG),
    .W2BEGb(Tile_X8Y5_W2BEGb),
    .WW4BEG(Tile_X8Y5_WW4BEG),
    .W6BEG(Tile_X8Y5_W6BEG),
    .Co(Tile_X8Y5_Co),
    .UserCLK(Tile_X8Y6_UserCLKo),
    .UserCLKo(Tile_X8Y5_UserCLKo),
    .FrameData(Tile_X7Y5_FrameData_O),
    .FrameData_O(Tile_X8Y5_FrameData_O),
    .FrameStrobe(Tile_X8Y6_FrameStrobe_O),
    .FrameStrobe_O(Tile_X8Y5_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X9Y5_Emulate_Bitstream)
    )
`endif
    Tile_X9Y5_LUT4AB
    (
    .N1END(Tile_X9Y6_N1BEG),
    .N2MID(Tile_X9Y6_N2BEG),
    .N2END(Tile_X9Y6_N2BEGb),
    .N4END(Tile_X9Y6_N4BEG),
    .NN4END(Tile_X9Y6_NN4BEG),
    .Ci(Tile_X9Y6_Co),
    .E1END(Tile_X8Y5_E1BEG),
    .E2MID(Tile_X8Y5_E2BEG),
    .E2END(Tile_X8Y5_E2BEGb),
    .EE4END(Tile_X8Y5_EE4BEG),
    .E6END(Tile_X8Y5_E6BEG),
    .S1END(Tile_X9Y4_S1BEG),
    .S2MID(Tile_X9Y4_S2BEG),
    .S2END(Tile_X9Y4_S2BEGb),
    .S4END(Tile_X9Y4_S4BEG),
    .SS4END(Tile_X9Y4_SS4BEG),
    .W1END(Tile_X10Y5_W1BEG),
    .W2MID(Tile_X10Y5_W2BEG),
    .W2END(Tile_X10Y5_W2BEGb),
    .WW4END(Tile_X10Y5_WW4BEG),
    .W6END(Tile_X10Y5_W6BEG),
    .N1BEG(Tile_X9Y5_N1BEG),
    .N2BEG(Tile_X9Y5_N2BEG),
    .N2BEGb(Tile_X9Y5_N2BEGb),
    .N4BEG(Tile_X9Y5_N4BEG),
    .NN4BEG(Tile_X9Y5_NN4BEG),
    .E1BEG(Tile_X9Y5_E1BEG),
    .E2BEG(Tile_X9Y5_E2BEG),
    .E2BEGb(Tile_X9Y5_E2BEGb),
    .EE4BEG(Tile_X9Y5_EE4BEG),
    .E6BEG(Tile_X9Y5_E6BEG),
    .S1BEG(Tile_X9Y5_S1BEG),
    .S2BEG(Tile_X9Y5_S2BEG),
    .S2BEGb(Tile_X9Y5_S2BEGb),
    .S4BEG(Tile_X9Y5_S4BEG),
    .SS4BEG(Tile_X9Y5_SS4BEG),
    .W1BEG(Tile_X9Y5_W1BEG),
    .W2BEG(Tile_X9Y5_W2BEG),
    .W2BEGb(Tile_X9Y5_W2BEGb),
    .WW4BEG(Tile_X9Y5_WW4BEG),
    .W6BEG(Tile_X9Y5_W6BEG),
    .Co(Tile_X9Y5_Co),
    .UserCLK(Tile_X9Y6_UserCLKo),
    .UserCLKo(Tile_X9Y5_UserCLKo),
    .FrameData(Tile_X8Y5_FrameData_O),
    .FrameData_O(Tile_X9Y5_FrameData_O),
    .FrameStrobe(Tile_X9Y6_FrameStrobe_O),
    .FrameStrobe_O(Tile_X9Y5_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
IHP_SRAM
`ifdef EMULATION
    #(
    .Tile_X0Y0_Emulate_Bitstream(`Tile_X10Y5_Emulate_Bitstream),
    .Tile_X0Y1_Emulate_Bitstream(`Tile_X10Y6_Emulate_Bitstream)
    )
`endif
    Tile_X10Y5_IHP_SRAM
    (
    .Tile_X0Y0_E1END(Tile_X9Y5_E1BEG),
    .Tile_X0Y0_E2MID(Tile_X9Y5_E2BEG),
    .Tile_X0Y0_E2END(Tile_X9Y5_E2BEGb),
    .Tile_X0Y0_EE4END(Tile_X9Y5_EE4BEG),
    .Tile_X0Y0_E6END(Tile_X9Y5_E6BEG),
    .Tile_X0Y0_S1END(Tile_X10Y4_S1BEG),
    .Tile_X0Y0_S2MID(Tile_X10Y4_S2BEG),
    .Tile_X0Y0_S2END(Tile_X10Y4_S2BEGb),
    .Tile_X0Y0_S4END(Tile_X10Y4_S4BEG),
    .Tile_X0Y1_N1END(Tile_X10Y7_N1BEG),
    .Tile_X0Y1_N2MID(Tile_X10Y7_N2BEG),
    .Tile_X0Y1_N2END(Tile_X10Y7_N2BEGb),
    .Tile_X0Y1_N4END(Tile_X10Y7_N4BEG),
    .Tile_X0Y1_E1END(Tile_X9Y6_E1BEG),
    .Tile_X0Y1_E2MID(Tile_X9Y6_E2BEG),
    .Tile_X0Y1_E2END(Tile_X9Y6_E2BEGb),
    .Tile_X0Y1_EE4END(Tile_X9Y6_EE4BEG),
    .Tile_X0Y1_E6END(Tile_X9Y6_E6BEG),
    .Tile_X0Y0_N1BEG(Tile_X10Y5_N1BEG),
    .Tile_X0Y0_N2BEG(Tile_X10Y5_N2BEG),
    .Tile_X0Y0_N2BEGb(Tile_X10Y5_N2BEGb),
    .Tile_X0Y0_N4BEG(Tile_X10Y5_N4BEG),
    .Tile_X0Y0_W1BEG(Tile_X10Y5_W1BEG),
    .Tile_X0Y0_W2BEG(Tile_X10Y5_W2BEG),
    .Tile_X0Y0_W2BEGb(Tile_X10Y5_W2BEGb),
    .Tile_X0Y0_WW4BEG(Tile_X10Y5_WW4BEG),
    .Tile_X0Y0_W6BEG(Tile_X10Y5_W6BEG),
    .Tile_X0Y1_S1BEG(Tile_X10Y6_S1BEG),
    .Tile_X0Y1_S2BEG(Tile_X10Y6_S2BEG),
    .Tile_X0Y1_S2BEGb(Tile_X10Y6_S2BEGb),
    .Tile_X0Y1_S4BEG(Tile_X10Y6_S4BEG),
    .Tile_X0Y1_W1BEG(Tile_X10Y6_W1BEG),
    .Tile_X0Y1_W2BEG(Tile_X10Y6_W2BEG),
    .Tile_X0Y1_W2BEGb(Tile_X10Y6_W2BEGb),
    .Tile_X0Y1_WW4BEG(Tile_X10Y6_WW4BEG),
    .Tile_X0Y1_W6BEG(Tile_X10Y6_W6BEG),
    .CONFIGURED_top(Tile_X10Y6_CONFIGURED_top),
    .DOUT_SRAM0(Tile_X10Y6_DOUT_SRAM0),
    .DOUT_SRAM1(Tile_X10Y6_DOUT_SRAM1),
    .DOUT_SRAM2(Tile_X10Y6_DOUT_SRAM2),
    .DOUT_SRAM3(Tile_X10Y6_DOUT_SRAM3),
    .DOUT_SRAM4(Tile_X10Y6_DOUT_SRAM4),
    .DOUT_SRAM5(Tile_X10Y6_DOUT_SRAM5),
    .DOUT_SRAM6(Tile_X10Y6_DOUT_SRAM6),
    .DOUT_SRAM7(Tile_X10Y6_DOUT_SRAM7),
    .DOUT_SRAM8(Tile_X10Y6_DOUT_SRAM8),
    .DOUT_SRAM9(Tile_X10Y6_DOUT_SRAM9),
    .DOUT_SRAM10(Tile_X10Y6_DOUT_SRAM10),
    .DOUT_SRAM11(Tile_X10Y6_DOUT_SRAM11),
    .DOUT_SRAM12(Tile_X10Y6_DOUT_SRAM12),
    .DOUT_SRAM13(Tile_X10Y6_DOUT_SRAM13),
    .DOUT_SRAM14(Tile_X10Y6_DOUT_SRAM14),
    .DOUT_SRAM15(Tile_X10Y6_DOUT_SRAM15),
    .DOUT_SRAM16(Tile_X10Y6_DOUT_SRAM16),
    .DOUT_SRAM17(Tile_X10Y6_DOUT_SRAM17),
    .DOUT_SRAM18(Tile_X10Y6_DOUT_SRAM18),
    .DOUT_SRAM19(Tile_X10Y6_DOUT_SRAM19),
    .DOUT_SRAM20(Tile_X10Y6_DOUT_SRAM20),
    .DOUT_SRAM21(Tile_X10Y6_DOUT_SRAM21),
    .DOUT_SRAM22(Tile_X10Y6_DOUT_SRAM22),
    .DOUT_SRAM23(Tile_X10Y6_DOUT_SRAM23),
    .DOUT_SRAM24(Tile_X10Y6_DOUT_SRAM24),
    .DOUT_SRAM25(Tile_X10Y6_DOUT_SRAM25),
    .DOUT_SRAM26(Tile_X10Y6_DOUT_SRAM26),
    .DOUT_SRAM27(Tile_X10Y6_DOUT_SRAM27),
    .DOUT_SRAM28(Tile_X10Y6_DOUT_SRAM28),
    .DOUT_SRAM29(Tile_X10Y6_DOUT_SRAM29),
    .DOUT_SRAM30(Tile_X10Y6_DOUT_SRAM30),
    .DOUT_SRAM31(Tile_X10Y6_DOUT_SRAM31),
    .ADDR_SRAM0(Tile_X10Y6_ADDR_SRAM0),
    .ADDR_SRAM1(Tile_X10Y6_ADDR_SRAM1),
    .ADDR_SRAM2(Tile_X10Y6_ADDR_SRAM2),
    .ADDR_SRAM3(Tile_X10Y6_ADDR_SRAM3),
    .ADDR_SRAM4(Tile_X10Y6_ADDR_SRAM4),
    .ADDR_SRAM5(Tile_X10Y6_ADDR_SRAM5),
    .ADDR_SRAM6(Tile_X10Y6_ADDR_SRAM6),
    .ADDR_SRAM7(Tile_X10Y6_ADDR_SRAM7),
    .ADDR_SRAM8(Tile_X10Y6_ADDR_SRAM8),
    .ADDR_SRAM9(Tile_X10Y6_ADDR_SRAM9),
    .BM_SRAM0(Tile_X10Y6_BM_SRAM0),
    .BM_SRAM1(Tile_X10Y6_BM_SRAM1),
    .BM_SRAM2(Tile_X10Y6_BM_SRAM2),
    .BM_SRAM3(Tile_X10Y6_BM_SRAM3),
    .BM_SRAM4(Tile_X10Y6_BM_SRAM4),
    .BM_SRAM5(Tile_X10Y6_BM_SRAM5),
    .BM_SRAM6(Tile_X10Y6_BM_SRAM6),
    .BM_SRAM7(Tile_X10Y6_BM_SRAM7),
    .BM_SRAM8(Tile_X10Y6_BM_SRAM8),
    .BM_SRAM9(Tile_X10Y6_BM_SRAM9),
    .BM_SRAM10(Tile_X10Y6_BM_SRAM10),
    .BM_SRAM11(Tile_X10Y6_BM_SRAM11),
    .BM_SRAM12(Tile_X10Y6_BM_SRAM12),
    .BM_SRAM13(Tile_X10Y6_BM_SRAM13),
    .BM_SRAM14(Tile_X10Y6_BM_SRAM14),
    .BM_SRAM15(Tile_X10Y6_BM_SRAM15),
    .BM_SRAM16(Tile_X10Y6_BM_SRAM16),
    .BM_SRAM17(Tile_X10Y6_BM_SRAM17),
    .BM_SRAM18(Tile_X10Y6_BM_SRAM18),
    .BM_SRAM19(Tile_X10Y6_BM_SRAM19),
    .BM_SRAM20(Tile_X10Y6_BM_SRAM20),
    .BM_SRAM21(Tile_X10Y6_BM_SRAM21),
    .BM_SRAM22(Tile_X10Y6_BM_SRAM22),
    .BM_SRAM23(Tile_X10Y6_BM_SRAM23),
    .BM_SRAM24(Tile_X10Y6_BM_SRAM24),
    .BM_SRAM25(Tile_X10Y6_BM_SRAM25),
    .BM_SRAM26(Tile_X10Y6_BM_SRAM26),
    .BM_SRAM27(Tile_X10Y6_BM_SRAM27),
    .BM_SRAM28(Tile_X10Y6_BM_SRAM28),
    .BM_SRAM29(Tile_X10Y6_BM_SRAM29),
    .BM_SRAM30(Tile_X10Y6_BM_SRAM30),
    .BM_SRAM31(Tile_X10Y6_BM_SRAM31),
    .CLK_SRAM(Tile_X10Y6_CLK_SRAM),
    .DIN_SRAM0(Tile_X10Y6_DIN_SRAM0),
    .DIN_SRAM1(Tile_X10Y6_DIN_SRAM1),
    .DIN_SRAM2(Tile_X10Y6_DIN_SRAM2),
    .DIN_SRAM3(Tile_X10Y6_DIN_SRAM3),
    .DIN_SRAM4(Tile_X10Y6_DIN_SRAM4),
    .DIN_SRAM5(Tile_X10Y6_DIN_SRAM5),
    .DIN_SRAM6(Tile_X10Y6_DIN_SRAM6),
    .DIN_SRAM7(Tile_X10Y6_DIN_SRAM7),
    .DIN_SRAM8(Tile_X10Y6_DIN_SRAM8),
    .DIN_SRAM9(Tile_X10Y6_DIN_SRAM9),
    .DIN_SRAM10(Tile_X10Y6_DIN_SRAM10),
    .DIN_SRAM11(Tile_X10Y6_DIN_SRAM11),
    .DIN_SRAM12(Tile_X10Y6_DIN_SRAM12),
    .DIN_SRAM13(Tile_X10Y6_DIN_SRAM13),
    .DIN_SRAM14(Tile_X10Y6_DIN_SRAM14),
    .DIN_SRAM15(Tile_X10Y6_DIN_SRAM15),
    .DIN_SRAM16(Tile_X10Y6_DIN_SRAM16),
    .DIN_SRAM17(Tile_X10Y6_DIN_SRAM17),
    .DIN_SRAM18(Tile_X10Y6_DIN_SRAM18),
    .DIN_SRAM19(Tile_X10Y6_DIN_SRAM19),
    .DIN_SRAM20(Tile_X10Y6_DIN_SRAM20),
    .DIN_SRAM21(Tile_X10Y6_DIN_SRAM21),
    .DIN_SRAM22(Tile_X10Y6_DIN_SRAM22),
    .DIN_SRAM23(Tile_X10Y6_DIN_SRAM23),
    .DIN_SRAM24(Tile_X10Y6_DIN_SRAM24),
    .DIN_SRAM25(Tile_X10Y6_DIN_SRAM25),
    .DIN_SRAM26(Tile_X10Y6_DIN_SRAM26),
    .DIN_SRAM27(Tile_X10Y6_DIN_SRAM27),
    .DIN_SRAM28(Tile_X10Y6_DIN_SRAM28),
    .DIN_SRAM29(Tile_X10Y6_DIN_SRAM29),
    .DIN_SRAM30(Tile_X10Y6_DIN_SRAM30),
    .DIN_SRAM31(Tile_X10Y6_DIN_SRAM31),
    .MEN_SRAM(Tile_X10Y6_MEN_SRAM),
    .REN_SRAM(Tile_X10Y6_REN_SRAM),
    .TIE_HIGH_SRAM(Tile_X10Y6_TIE_HIGH_SRAM),
    .TIE_LOW_SRAM(Tile_X10Y6_TIE_LOW_SRAM),
    .WEN_SRAM(Tile_X10Y6_WEN_SRAM),
    .Tile_X0Y0_UserCLKo(Tile_X10Y5_UserCLKo),
    .Tile_X0Y1_UserCLK(Tile_X10Y7_UserCLKo),
    .Tile_X0Y0_FrameData(Tile_X9Y5_FrameData_O),
    .Tile_X0Y0_FrameData_O(Tile_X10Y5_FrameData_O),
    .Tile_X0Y0_FrameStrobe_O(Tile_X10Y5_FrameStrobe_O),
    .Tile_X0Y1_FrameData(Tile_X9Y6_FrameData_O),
    .Tile_X0Y1_FrameData_O(Tile_X10Y6_FrameData_O),
    .Tile_X0Y1_FrameStrobe(Tile_X10Y7_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
W_IO
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X0Y6_Emulate_Bitstream)
    )
`endif
    Tile_X0Y6_W_IO
    (
    .W1END(Tile_X1Y6_W1BEG),
    .W2MID(Tile_X1Y6_W2BEG),
    .W2END(Tile_X1Y6_W2BEGb),
    .WW4END(Tile_X1Y6_WW4BEG),
    .W6END(Tile_X1Y6_W6BEG),
    .E1BEG(Tile_X0Y6_E1BEG),
    .E2BEG(Tile_X0Y6_E2BEG),
    .E2BEGb(Tile_X0Y6_E2BEGb),
    .EE4BEG(Tile_X0Y6_EE4BEG),
    .E6BEG(Tile_X0Y6_E6BEG),
    .A_O_top(Tile_X0Y6_A_O_top),
    .A_I_top(Tile_X0Y6_A_I_top),
    .A_T_top(Tile_X0Y6_A_T_top),
    .B_O_top(Tile_X0Y6_B_O_top),
    .B_I_top(Tile_X0Y6_B_I_top),
    .B_T_top(Tile_X0Y6_B_T_top),
    .A_config_C_bit0(Tile_X0Y6_A_config_C_bit0),
    .A_config_C_bit1(Tile_X0Y6_A_config_C_bit1),
    .A_config_C_bit2(Tile_X0Y6_A_config_C_bit2),
    .A_config_C_bit3(Tile_X0Y6_A_config_C_bit3),
    .B_config_C_bit0(Tile_X0Y6_B_config_C_bit0),
    .B_config_C_bit1(Tile_X0Y6_B_config_C_bit1),
    .B_config_C_bit2(Tile_X0Y6_B_config_C_bit2),
    .B_config_C_bit3(Tile_X0Y6_B_config_C_bit3),
    .UserCLK(Tile_X0Y7_UserCLKo),
    .UserCLKo(Tile_X0Y6_UserCLKo),
    .FrameData(Row_Y6_FrameData),
    .FrameData_O(Tile_X0Y6_FrameData_O),
    .FrameStrobe(Tile_X0Y7_FrameStrobe_O),
    .FrameStrobe_O(Tile_X0Y6_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X1Y6_Emulate_Bitstream)
    )
`endif
    Tile_X1Y6_LUT4AB
    (
    .N1END(Tile_X1Y7_N1BEG),
    .N2MID(Tile_X1Y7_N2BEG),
    .N2END(Tile_X1Y7_N2BEGb),
    .N4END(Tile_X1Y7_N4BEG),
    .NN4END(Tile_X1Y7_NN4BEG),
    .Ci(Tile_X1Y7_Co),
    .E1END(Tile_X0Y6_E1BEG),
    .E2MID(Tile_X0Y6_E2BEG),
    .E2END(Tile_X0Y6_E2BEGb),
    .EE4END(Tile_X0Y6_EE4BEG),
    .E6END(Tile_X0Y6_E6BEG),
    .S1END(Tile_X1Y5_S1BEG),
    .S2MID(Tile_X1Y5_S2BEG),
    .S2END(Tile_X1Y5_S2BEGb),
    .S4END(Tile_X1Y5_S4BEG),
    .SS4END(Tile_X1Y5_SS4BEG),
    .W1END(Tile_X2Y6_W1BEG),
    .W2MID(Tile_X2Y6_W2BEG),
    .W2END(Tile_X2Y6_W2BEGb),
    .WW4END(Tile_X2Y6_WW4BEG),
    .W6END(Tile_X2Y6_W6BEG),
    .N1BEG(Tile_X1Y6_N1BEG),
    .N2BEG(Tile_X1Y6_N2BEG),
    .N2BEGb(Tile_X1Y6_N2BEGb),
    .N4BEG(Tile_X1Y6_N4BEG),
    .NN4BEG(Tile_X1Y6_NN4BEG),
    .E1BEG(Tile_X1Y6_E1BEG),
    .E2BEG(Tile_X1Y6_E2BEG),
    .E2BEGb(Tile_X1Y6_E2BEGb),
    .EE4BEG(Tile_X1Y6_EE4BEG),
    .E6BEG(Tile_X1Y6_E6BEG),
    .S1BEG(Tile_X1Y6_S1BEG),
    .S2BEG(Tile_X1Y6_S2BEG),
    .S2BEGb(Tile_X1Y6_S2BEGb),
    .S4BEG(Tile_X1Y6_S4BEG),
    .SS4BEG(Tile_X1Y6_SS4BEG),
    .W1BEG(Tile_X1Y6_W1BEG),
    .W2BEG(Tile_X1Y6_W2BEG),
    .W2BEGb(Tile_X1Y6_W2BEGb),
    .WW4BEG(Tile_X1Y6_WW4BEG),
    .W6BEG(Tile_X1Y6_W6BEG),
    .Co(Tile_X1Y6_Co),
    .UserCLK(Tile_X1Y7_UserCLKo),
    .UserCLKo(Tile_X1Y6_UserCLKo),
    .FrameData(Tile_X0Y6_FrameData_O),
    .FrameData_O(Tile_X1Y6_FrameData_O),
    .FrameStrobe(Tile_X1Y7_FrameStrobe_O),
    .FrameStrobe_O(Tile_X1Y6_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X2Y6_Emulate_Bitstream)
    )
`endif
    Tile_X2Y6_LUT4AB
    (
    .N1END(Tile_X2Y7_N1BEG),
    .N2MID(Tile_X2Y7_N2BEG),
    .N2END(Tile_X2Y7_N2BEGb),
    .N4END(Tile_X2Y7_N4BEG),
    .NN4END(Tile_X2Y7_NN4BEG),
    .Ci(Tile_X2Y7_Co),
    .E1END(Tile_X1Y6_E1BEG),
    .E2MID(Tile_X1Y6_E2BEG),
    .E2END(Tile_X1Y6_E2BEGb),
    .EE4END(Tile_X1Y6_EE4BEG),
    .E6END(Tile_X1Y6_E6BEG),
    .S1END(Tile_X2Y5_S1BEG),
    .S2MID(Tile_X2Y5_S2BEG),
    .S2END(Tile_X2Y5_S2BEGb),
    .S4END(Tile_X2Y5_S4BEG),
    .SS4END(Tile_X2Y5_SS4BEG),
    .W1END(Tile_X3Y6_W1BEG),
    .W2MID(Tile_X3Y6_W2BEG),
    .W2END(Tile_X3Y6_W2BEGb),
    .WW4END(Tile_X3Y6_WW4BEG),
    .W6END(Tile_X3Y6_W6BEG),
    .N1BEG(Tile_X2Y6_N1BEG),
    .N2BEG(Tile_X2Y6_N2BEG),
    .N2BEGb(Tile_X2Y6_N2BEGb),
    .N4BEG(Tile_X2Y6_N4BEG),
    .NN4BEG(Tile_X2Y6_NN4BEG),
    .E1BEG(Tile_X2Y6_E1BEG),
    .E2BEG(Tile_X2Y6_E2BEG),
    .E2BEGb(Tile_X2Y6_E2BEGb),
    .EE4BEG(Tile_X2Y6_EE4BEG),
    .E6BEG(Tile_X2Y6_E6BEG),
    .S1BEG(Tile_X2Y6_S1BEG),
    .S2BEG(Tile_X2Y6_S2BEG),
    .S2BEGb(Tile_X2Y6_S2BEGb),
    .S4BEG(Tile_X2Y6_S4BEG),
    .SS4BEG(Tile_X2Y6_SS4BEG),
    .W1BEG(Tile_X2Y6_W1BEG),
    .W2BEG(Tile_X2Y6_W2BEG),
    .W2BEGb(Tile_X2Y6_W2BEGb),
    .WW4BEG(Tile_X2Y6_WW4BEG),
    .W6BEG(Tile_X2Y6_W6BEG),
    .Co(Tile_X2Y6_Co),
    .UserCLK(Tile_X2Y7_UserCLKo),
    .UserCLKo(Tile_X2Y6_UserCLKo),
    .FrameData(Tile_X1Y6_FrameData_O),
    .FrameData_O(Tile_X2Y6_FrameData_O),
    .FrameStrobe(Tile_X2Y7_FrameStrobe_O),
    .FrameStrobe_O(Tile_X2Y6_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X3Y6_Emulate_Bitstream)
    )
`endif
    Tile_X3Y6_LUT4AB
    (
    .N1END(Tile_X3Y7_N1BEG),
    .N2MID(Tile_X3Y7_N2BEG),
    .N2END(Tile_X3Y7_N2BEGb),
    .N4END(Tile_X3Y7_N4BEG),
    .NN4END(Tile_X3Y7_NN4BEG),
    .Ci(Tile_X3Y7_Co),
    .E1END(Tile_X2Y6_E1BEG),
    .E2MID(Tile_X2Y6_E2BEG),
    .E2END(Tile_X2Y6_E2BEGb),
    .EE4END(Tile_X2Y6_EE4BEG),
    .E6END(Tile_X2Y6_E6BEG),
    .S1END(Tile_X3Y5_S1BEG),
    .S2MID(Tile_X3Y5_S2BEG),
    .S2END(Tile_X3Y5_S2BEGb),
    .S4END(Tile_X3Y5_S4BEG),
    .SS4END(Tile_X3Y5_SS4BEG),
    .W1END(Tile_X4Y6_W1BEG),
    .W2MID(Tile_X4Y6_W2BEG),
    .W2END(Tile_X4Y6_W2BEGb),
    .WW4END(Tile_X4Y6_WW4BEG),
    .W6END(Tile_X4Y6_W6BEG),
    .N1BEG(Tile_X3Y6_N1BEG),
    .N2BEG(Tile_X3Y6_N2BEG),
    .N2BEGb(Tile_X3Y6_N2BEGb),
    .N4BEG(Tile_X3Y6_N4BEG),
    .NN4BEG(Tile_X3Y6_NN4BEG),
    .E1BEG(Tile_X3Y6_E1BEG),
    .E2BEG(Tile_X3Y6_E2BEG),
    .E2BEGb(Tile_X3Y6_E2BEGb),
    .EE4BEG(Tile_X3Y6_EE4BEG),
    .E6BEG(Tile_X3Y6_E6BEG),
    .S1BEG(Tile_X3Y6_S1BEG),
    .S2BEG(Tile_X3Y6_S2BEG),
    .S2BEGb(Tile_X3Y6_S2BEGb),
    .S4BEG(Tile_X3Y6_S4BEG),
    .SS4BEG(Tile_X3Y6_SS4BEG),
    .W1BEG(Tile_X3Y6_W1BEG),
    .W2BEG(Tile_X3Y6_W2BEG),
    .W2BEGb(Tile_X3Y6_W2BEGb),
    .WW4BEG(Tile_X3Y6_WW4BEG),
    .W6BEG(Tile_X3Y6_W6BEG),
    .Co(Tile_X3Y6_Co),
    .UserCLK(Tile_X3Y7_UserCLKo),
    .UserCLKo(Tile_X3Y6_UserCLKo),
    .FrameData(Tile_X2Y6_FrameData_O),
    .FrameData_O(Tile_X3Y6_FrameData_O),
    .FrameStrobe(Tile_X3Y7_FrameStrobe_O),
    .FrameStrobe_O(Tile_X3Y6_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
RegFile
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X4Y6_Emulate_Bitstream)
    )
`endif
    Tile_X4Y6_RegFile
    (
    .N1END(Tile_X4Y7_N1BEG),
    .N2MID(Tile_X4Y7_N2BEG),
    .N2END(Tile_X4Y7_N2BEGb),
    .N4END(Tile_X4Y7_N4BEG),
    .NN4END(Tile_X4Y7_NN4BEG),
    .E1END(Tile_X3Y6_E1BEG),
    .E2MID(Tile_X3Y6_E2BEG),
    .E2END(Tile_X3Y6_E2BEGb),
    .EE4END(Tile_X3Y6_EE4BEG),
    .E6END(Tile_X3Y6_E6BEG),
    .S1END(Tile_X4Y5_S1BEG),
    .S2MID(Tile_X4Y5_S2BEG),
    .S2END(Tile_X4Y5_S2BEGb),
    .S4END(Tile_X4Y5_S4BEG),
    .SS4END(Tile_X4Y5_SS4BEG),
    .W1END(Tile_X5Y6_W1BEG),
    .W2MID(Tile_X5Y6_W2BEG),
    .W2END(Tile_X5Y6_W2BEGb),
    .WW4END(Tile_X5Y6_WW4BEG),
    .W6END(Tile_X5Y6_W6BEG),
    .N1BEG(Tile_X4Y6_N1BEG),
    .N2BEG(Tile_X4Y6_N2BEG),
    .N2BEGb(Tile_X4Y6_N2BEGb),
    .N4BEG(Tile_X4Y6_N4BEG),
    .NN4BEG(Tile_X4Y6_NN4BEG),
    .E1BEG(Tile_X4Y6_E1BEG),
    .E2BEG(Tile_X4Y6_E2BEG),
    .E2BEGb(Tile_X4Y6_E2BEGb),
    .EE4BEG(Tile_X4Y6_EE4BEG),
    .E6BEG(Tile_X4Y6_E6BEG),
    .S1BEG(Tile_X4Y6_S1BEG),
    .S2BEG(Tile_X4Y6_S2BEG),
    .S2BEGb(Tile_X4Y6_S2BEGb),
    .S4BEG(Tile_X4Y6_S4BEG),
    .SS4BEG(Tile_X4Y6_SS4BEG),
    .W1BEG(Tile_X4Y6_W1BEG),
    .W2BEG(Tile_X4Y6_W2BEG),
    .W2BEGb(Tile_X4Y6_W2BEGb),
    .WW4BEG(Tile_X4Y6_WW4BEG),
    .W6BEG(Tile_X4Y6_W6BEG),
    .UserCLK(Tile_X4Y7_UserCLKo),
    .UserCLKo(Tile_X4Y6_UserCLKo),
    .FrameData(Tile_X3Y6_FrameData_O),
    .FrameData_O(Tile_X4Y6_FrameData_O),
    .FrameStrobe(Tile_X4Y7_FrameStrobe_O),
    .FrameStrobe_O(Tile_X4Y6_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X5Y6_Emulate_Bitstream)
    )
`endif
    Tile_X5Y6_LUT4AB
    (
    .N1END(Tile_X5Y7_N1BEG),
    .N2MID(Tile_X5Y7_N2BEG),
    .N2END(Tile_X5Y7_N2BEGb),
    .N4END(Tile_X5Y7_N4BEG),
    .NN4END(Tile_X5Y7_NN4BEG),
    .Ci(Tile_X5Y7_Co),
    .E1END(Tile_X4Y6_E1BEG),
    .E2MID(Tile_X4Y6_E2BEG),
    .E2END(Tile_X4Y6_E2BEGb),
    .EE4END(Tile_X4Y6_EE4BEG),
    .E6END(Tile_X4Y6_E6BEG),
    .S1END(Tile_X5Y5_S1BEG),
    .S2MID(Tile_X5Y5_S2BEG),
    .S2END(Tile_X5Y5_S2BEGb),
    .S4END(Tile_X5Y5_S4BEG),
    .SS4END(Tile_X5Y5_SS4BEG),
    .W1END(Tile_X6Y6_W1BEG),
    .W2MID(Tile_X6Y6_W2BEG),
    .W2END(Tile_X6Y6_W2BEGb),
    .WW4END(Tile_X6Y6_WW4BEG),
    .W6END(Tile_X6Y6_W6BEG),
    .N1BEG(Tile_X5Y6_N1BEG),
    .N2BEG(Tile_X5Y6_N2BEG),
    .N2BEGb(Tile_X5Y6_N2BEGb),
    .N4BEG(Tile_X5Y6_N4BEG),
    .NN4BEG(Tile_X5Y6_NN4BEG),
    .E1BEG(Tile_X5Y6_E1BEG),
    .E2BEG(Tile_X5Y6_E2BEG),
    .E2BEGb(Tile_X5Y6_E2BEGb),
    .EE4BEG(Tile_X5Y6_EE4BEG),
    .E6BEG(Tile_X5Y6_E6BEG),
    .S1BEG(Tile_X5Y6_S1BEG),
    .S2BEG(Tile_X5Y6_S2BEG),
    .S2BEGb(Tile_X5Y6_S2BEGb),
    .S4BEG(Tile_X5Y6_S4BEG),
    .SS4BEG(Tile_X5Y6_SS4BEG),
    .W1BEG(Tile_X5Y6_W1BEG),
    .W2BEG(Tile_X5Y6_W2BEG),
    .W2BEGb(Tile_X5Y6_W2BEGb),
    .WW4BEG(Tile_X5Y6_WW4BEG),
    .W6BEG(Tile_X5Y6_W6BEG),
    .Co(Tile_X5Y6_Co),
    .UserCLK(Tile_X5Y7_UserCLKo),
    .UserCLKo(Tile_X5Y6_UserCLKo),
    .FrameData(Tile_X4Y6_FrameData_O),
    .FrameData_O(Tile_X5Y6_FrameData_O),
    .FrameStrobe(Tile_X5Y7_FrameStrobe_O),
    .FrameStrobe_O(Tile_X5Y6_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X6Y6_Emulate_Bitstream)
    )
`endif
    Tile_X6Y6_LUT4AB
    (
    .N1END(Tile_X6Y7_N1BEG),
    .N2MID(Tile_X6Y7_N2BEG),
    .N2END(Tile_X6Y7_N2BEGb),
    .N4END(Tile_X6Y7_N4BEG),
    .NN4END(Tile_X6Y7_NN4BEG),
    .Ci(Tile_X6Y7_Co),
    .E1END(Tile_X5Y6_E1BEG),
    .E2MID(Tile_X5Y6_E2BEG),
    .E2END(Tile_X5Y6_E2BEGb),
    .EE4END(Tile_X5Y6_EE4BEG),
    .E6END(Tile_X5Y6_E6BEG),
    .S1END(Tile_X6Y5_S1BEG),
    .S2MID(Tile_X6Y5_S2BEG),
    .S2END(Tile_X6Y5_S2BEGb),
    .S4END(Tile_X6Y5_S4BEG),
    .SS4END(Tile_X6Y5_SS4BEG),
    .W1END(Tile_X7Y6_W1BEG),
    .W2MID(Tile_X7Y6_W2BEG),
    .W2END(Tile_X7Y6_W2BEGb),
    .WW4END(Tile_X7Y6_WW4BEG),
    .W6END(Tile_X7Y6_W6BEG),
    .N1BEG(Tile_X6Y6_N1BEG),
    .N2BEG(Tile_X6Y6_N2BEG),
    .N2BEGb(Tile_X6Y6_N2BEGb),
    .N4BEG(Tile_X6Y6_N4BEG),
    .NN4BEG(Tile_X6Y6_NN4BEG),
    .E1BEG(Tile_X6Y6_E1BEG),
    .E2BEG(Tile_X6Y6_E2BEG),
    .E2BEGb(Tile_X6Y6_E2BEGb),
    .EE4BEG(Tile_X6Y6_EE4BEG),
    .E6BEG(Tile_X6Y6_E6BEG),
    .S1BEG(Tile_X6Y6_S1BEG),
    .S2BEG(Tile_X6Y6_S2BEG),
    .S2BEGb(Tile_X6Y6_S2BEGb),
    .S4BEG(Tile_X6Y6_S4BEG),
    .SS4BEG(Tile_X6Y6_SS4BEG),
    .W1BEG(Tile_X6Y6_W1BEG),
    .W2BEG(Tile_X6Y6_W2BEG),
    .W2BEGb(Tile_X6Y6_W2BEGb),
    .WW4BEG(Tile_X6Y6_WW4BEG),
    .W6BEG(Tile_X6Y6_W6BEG),
    .Co(Tile_X6Y6_Co),
    .UserCLK(Tile_X6Y7_UserCLKo),
    .UserCLKo(Tile_X6Y6_UserCLKo),
    .FrameData(Tile_X5Y6_FrameData_O),
    .FrameData_O(Tile_X6Y6_FrameData_O),
    .FrameStrobe(Tile_X6Y7_FrameStrobe_O),
    .FrameStrobe_O(Tile_X6Y6_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X8Y6_Emulate_Bitstream)
    )
`endif
    Tile_X8Y6_LUT4AB
    (
    .N1END(Tile_X8Y7_N1BEG),
    .N2MID(Tile_X8Y7_N2BEG),
    .N2END(Tile_X8Y7_N2BEGb),
    .N4END(Tile_X8Y7_N4BEG),
    .NN4END(Tile_X8Y7_NN4BEG),
    .Ci(Tile_X8Y7_Co),
    .E1END(Tile_X7Y6_E1BEG),
    .E2MID(Tile_X7Y6_E2BEG),
    .E2END(Tile_X7Y6_E2BEGb),
    .EE4END(Tile_X7Y6_EE4BEG),
    .E6END(Tile_X7Y6_E6BEG),
    .S1END(Tile_X8Y5_S1BEG),
    .S2MID(Tile_X8Y5_S2BEG),
    .S2END(Tile_X8Y5_S2BEGb),
    .S4END(Tile_X8Y5_S4BEG),
    .SS4END(Tile_X8Y5_SS4BEG),
    .W1END(Tile_X9Y6_W1BEG),
    .W2MID(Tile_X9Y6_W2BEG),
    .W2END(Tile_X9Y6_W2BEGb),
    .WW4END(Tile_X9Y6_WW4BEG),
    .W6END(Tile_X9Y6_W6BEG),
    .N1BEG(Tile_X8Y6_N1BEG),
    .N2BEG(Tile_X8Y6_N2BEG),
    .N2BEGb(Tile_X8Y6_N2BEGb),
    .N4BEG(Tile_X8Y6_N4BEG),
    .NN4BEG(Tile_X8Y6_NN4BEG),
    .E1BEG(Tile_X8Y6_E1BEG),
    .E2BEG(Tile_X8Y6_E2BEG),
    .E2BEGb(Tile_X8Y6_E2BEGb),
    .EE4BEG(Tile_X8Y6_EE4BEG),
    .E6BEG(Tile_X8Y6_E6BEG),
    .S1BEG(Tile_X8Y6_S1BEG),
    .S2BEG(Tile_X8Y6_S2BEG),
    .S2BEGb(Tile_X8Y6_S2BEGb),
    .S4BEG(Tile_X8Y6_S4BEG),
    .SS4BEG(Tile_X8Y6_SS4BEG),
    .W1BEG(Tile_X8Y6_W1BEG),
    .W2BEG(Tile_X8Y6_W2BEG),
    .W2BEGb(Tile_X8Y6_W2BEGb),
    .WW4BEG(Tile_X8Y6_WW4BEG),
    .W6BEG(Tile_X8Y6_W6BEG),
    .Co(Tile_X8Y6_Co),
    .UserCLK(Tile_X8Y7_UserCLKo),
    .UserCLKo(Tile_X8Y6_UserCLKo),
    .FrameData(Tile_X7Y6_FrameData_O),
    .FrameData_O(Tile_X8Y6_FrameData_O),
    .FrameStrobe(Tile_X8Y7_FrameStrobe_O),
    .FrameStrobe_O(Tile_X8Y6_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X9Y6_Emulate_Bitstream)
    )
`endif
    Tile_X9Y6_LUT4AB
    (
    .N1END(Tile_X9Y7_N1BEG),
    .N2MID(Tile_X9Y7_N2BEG),
    .N2END(Tile_X9Y7_N2BEGb),
    .N4END(Tile_X9Y7_N4BEG),
    .NN4END(Tile_X9Y7_NN4BEG),
    .Ci(Tile_X9Y7_Co),
    .E1END(Tile_X8Y6_E1BEG),
    .E2MID(Tile_X8Y6_E2BEG),
    .E2END(Tile_X8Y6_E2BEGb),
    .EE4END(Tile_X8Y6_EE4BEG),
    .E6END(Tile_X8Y6_E6BEG),
    .S1END(Tile_X9Y5_S1BEG),
    .S2MID(Tile_X9Y5_S2BEG),
    .S2END(Tile_X9Y5_S2BEGb),
    .S4END(Tile_X9Y5_S4BEG),
    .SS4END(Tile_X9Y5_SS4BEG),
    .W1END(Tile_X10Y6_W1BEG),
    .W2MID(Tile_X10Y6_W2BEG),
    .W2END(Tile_X10Y6_W2BEGb),
    .WW4END(Tile_X10Y6_WW4BEG),
    .W6END(Tile_X10Y6_W6BEG),
    .N1BEG(Tile_X9Y6_N1BEG),
    .N2BEG(Tile_X9Y6_N2BEG),
    .N2BEGb(Tile_X9Y6_N2BEGb),
    .N4BEG(Tile_X9Y6_N4BEG),
    .NN4BEG(Tile_X9Y6_NN4BEG),
    .E1BEG(Tile_X9Y6_E1BEG),
    .E2BEG(Tile_X9Y6_E2BEG),
    .E2BEGb(Tile_X9Y6_E2BEGb),
    .EE4BEG(Tile_X9Y6_EE4BEG),
    .E6BEG(Tile_X9Y6_E6BEG),
    .S1BEG(Tile_X9Y6_S1BEG),
    .S2BEG(Tile_X9Y6_S2BEG),
    .S2BEGb(Tile_X9Y6_S2BEGb),
    .S4BEG(Tile_X9Y6_S4BEG),
    .SS4BEG(Tile_X9Y6_SS4BEG),
    .W1BEG(Tile_X9Y6_W1BEG),
    .W2BEG(Tile_X9Y6_W2BEG),
    .W2BEGb(Tile_X9Y6_W2BEGb),
    .WW4BEG(Tile_X9Y6_WW4BEG),
    .W6BEG(Tile_X9Y6_W6BEG),
    .Co(Tile_X9Y6_Co),
    .UserCLK(Tile_X9Y7_UserCLKo),
    .UserCLKo(Tile_X9Y6_UserCLKo),
    .FrameData(Tile_X8Y6_FrameData_O),
    .FrameData_O(Tile_X9Y6_FrameData_O),
    .FrameStrobe(Tile_X9Y7_FrameStrobe_O),
    .FrameStrobe_O(Tile_X9Y6_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
W_IO
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X0Y7_Emulate_Bitstream)
    )
`endif
    Tile_X0Y7_W_IO
    (
    .W1END(Tile_X1Y7_W1BEG),
    .W2MID(Tile_X1Y7_W2BEG),
    .W2END(Tile_X1Y7_W2BEGb),
    .WW4END(Tile_X1Y7_WW4BEG),
    .W6END(Tile_X1Y7_W6BEG),
    .E1BEG(Tile_X0Y7_E1BEG),
    .E2BEG(Tile_X0Y7_E2BEG),
    .E2BEGb(Tile_X0Y7_E2BEGb),
    .EE4BEG(Tile_X0Y7_EE4BEG),
    .E6BEG(Tile_X0Y7_E6BEG),
    .A_O_top(Tile_X0Y7_A_O_top),
    .A_I_top(Tile_X0Y7_A_I_top),
    .A_T_top(Tile_X0Y7_A_T_top),
    .B_O_top(Tile_X0Y7_B_O_top),
    .B_I_top(Tile_X0Y7_B_I_top),
    .B_T_top(Tile_X0Y7_B_T_top),
    .A_config_C_bit0(Tile_X0Y7_A_config_C_bit0),
    .A_config_C_bit1(Tile_X0Y7_A_config_C_bit1),
    .A_config_C_bit2(Tile_X0Y7_A_config_C_bit2),
    .A_config_C_bit3(Tile_X0Y7_A_config_C_bit3),
    .B_config_C_bit0(Tile_X0Y7_B_config_C_bit0),
    .B_config_C_bit1(Tile_X0Y7_B_config_C_bit1),
    .B_config_C_bit2(Tile_X0Y7_B_config_C_bit2),
    .B_config_C_bit3(Tile_X0Y7_B_config_C_bit3),
    .UserCLK(Tile_X0Y8_UserCLKo),
    .UserCLKo(Tile_X0Y7_UserCLKo),
    .FrameData(Row_Y7_FrameData),
    .FrameData_O(Tile_X0Y7_FrameData_O),
    .FrameStrobe(Tile_X0Y8_FrameStrobe_O),
    .FrameStrobe_O(Tile_X0Y7_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X1Y7_Emulate_Bitstream)
    )
`endif
    Tile_X1Y7_LUT4AB
    (
    .N1END(Tile_X1Y8_N1BEG),
    .N2MID(Tile_X1Y8_N2BEG),
    .N2END(Tile_X1Y8_N2BEGb),
    .N4END(Tile_X1Y8_N4BEG),
    .NN4END(Tile_X1Y8_NN4BEG),
    .Ci(Tile_X1Y8_Co),
    .E1END(Tile_X0Y7_E1BEG),
    .E2MID(Tile_X0Y7_E2BEG),
    .E2END(Tile_X0Y7_E2BEGb),
    .EE4END(Tile_X0Y7_EE4BEG),
    .E6END(Tile_X0Y7_E6BEG),
    .S1END(Tile_X1Y6_S1BEG),
    .S2MID(Tile_X1Y6_S2BEG),
    .S2END(Tile_X1Y6_S2BEGb),
    .S4END(Tile_X1Y6_S4BEG),
    .SS4END(Tile_X1Y6_SS4BEG),
    .W1END(Tile_X2Y7_W1BEG),
    .W2MID(Tile_X2Y7_W2BEG),
    .W2END(Tile_X2Y7_W2BEGb),
    .WW4END(Tile_X2Y7_WW4BEG),
    .W6END(Tile_X2Y7_W6BEG),
    .N1BEG(Tile_X1Y7_N1BEG),
    .N2BEG(Tile_X1Y7_N2BEG),
    .N2BEGb(Tile_X1Y7_N2BEGb),
    .N4BEG(Tile_X1Y7_N4BEG),
    .NN4BEG(Tile_X1Y7_NN4BEG),
    .E1BEG(Tile_X1Y7_E1BEG),
    .E2BEG(Tile_X1Y7_E2BEG),
    .E2BEGb(Tile_X1Y7_E2BEGb),
    .EE4BEG(Tile_X1Y7_EE4BEG),
    .E6BEG(Tile_X1Y7_E6BEG),
    .S1BEG(Tile_X1Y7_S1BEG),
    .S2BEG(Tile_X1Y7_S2BEG),
    .S2BEGb(Tile_X1Y7_S2BEGb),
    .S4BEG(Tile_X1Y7_S4BEG),
    .SS4BEG(Tile_X1Y7_SS4BEG),
    .W1BEG(Tile_X1Y7_W1BEG),
    .W2BEG(Tile_X1Y7_W2BEG),
    .W2BEGb(Tile_X1Y7_W2BEGb),
    .WW4BEG(Tile_X1Y7_WW4BEG),
    .W6BEG(Tile_X1Y7_W6BEG),
    .Co(Tile_X1Y7_Co),
    .UserCLK(Tile_X1Y8_UserCLKo),
    .UserCLKo(Tile_X1Y7_UserCLKo),
    .FrameData(Tile_X0Y7_FrameData_O),
    .FrameData_O(Tile_X1Y7_FrameData_O),
    .FrameStrobe(Tile_X1Y8_FrameStrobe_O),
    .FrameStrobe_O(Tile_X1Y7_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X2Y7_Emulate_Bitstream)
    )
`endif
    Tile_X2Y7_LUT4AB
    (
    .N1END(Tile_X2Y8_N1BEG),
    .N2MID(Tile_X2Y8_N2BEG),
    .N2END(Tile_X2Y8_N2BEGb),
    .N4END(Tile_X2Y8_N4BEG),
    .NN4END(Tile_X2Y8_NN4BEG),
    .Ci(Tile_X2Y8_Co),
    .E1END(Tile_X1Y7_E1BEG),
    .E2MID(Tile_X1Y7_E2BEG),
    .E2END(Tile_X1Y7_E2BEGb),
    .EE4END(Tile_X1Y7_EE4BEG),
    .E6END(Tile_X1Y7_E6BEG),
    .S1END(Tile_X2Y6_S1BEG),
    .S2MID(Tile_X2Y6_S2BEG),
    .S2END(Tile_X2Y6_S2BEGb),
    .S4END(Tile_X2Y6_S4BEG),
    .SS4END(Tile_X2Y6_SS4BEG),
    .W1END(Tile_X3Y7_W1BEG),
    .W2MID(Tile_X3Y7_W2BEG),
    .W2END(Tile_X3Y7_W2BEGb),
    .WW4END(Tile_X3Y7_WW4BEG),
    .W6END(Tile_X3Y7_W6BEG),
    .N1BEG(Tile_X2Y7_N1BEG),
    .N2BEG(Tile_X2Y7_N2BEG),
    .N2BEGb(Tile_X2Y7_N2BEGb),
    .N4BEG(Tile_X2Y7_N4BEG),
    .NN4BEG(Tile_X2Y7_NN4BEG),
    .E1BEG(Tile_X2Y7_E1BEG),
    .E2BEG(Tile_X2Y7_E2BEG),
    .E2BEGb(Tile_X2Y7_E2BEGb),
    .EE4BEG(Tile_X2Y7_EE4BEG),
    .E6BEG(Tile_X2Y7_E6BEG),
    .S1BEG(Tile_X2Y7_S1BEG),
    .S2BEG(Tile_X2Y7_S2BEG),
    .S2BEGb(Tile_X2Y7_S2BEGb),
    .S4BEG(Tile_X2Y7_S4BEG),
    .SS4BEG(Tile_X2Y7_SS4BEG),
    .W1BEG(Tile_X2Y7_W1BEG),
    .W2BEG(Tile_X2Y7_W2BEG),
    .W2BEGb(Tile_X2Y7_W2BEGb),
    .WW4BEG(Tile_X2Y7_WW4BEG),
    .W6BEG(Tile_X2Y7_W6BEG),
    .Co(Tile_X2Y7_Co),
    .UserCLK(Tile_X2Y8_UserCLKo),
    .UserCLKo(Tile_X2Y7_UserCLKo),
    .FrameData(Tile_X1Y7_FrameData_O),
    .FrameData_O(Tile_X2Y7_FrameData_O),
    .FrameStrobe(Tile_X2Y8_FrameStrobe_O),
    .FrameStrobe_O(Tile_X2Y7_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X3Y7_Emulate_Bitstream)
    )
`endif
    Tile_X3Y7_LUT4AB
    (
    .N1END(Tile_X3Y8_N1BEG),
    .N2MID(Tile_X3Y8_N2BEG),
    .N2END(Tile_X3Y8_N2BEGb),
    .N4END(Tile_X3Y8_N4BEG),
    .NN4END(Tile_X3Y8_NN4BEG),
    .Ci(Tile_X3Y8_Co),
    .E1END(Tile_X2Y7_E1BEG),
    .E2MID(Tile_X2Y7_E2BEG),
    .E2END(Tile_X2Y7_E2BEGb),
    .EE4END(Tile_X2Y7_EE4BEG),
    .E6END(Tile_X2Y7_E6BEG),
    .S1END(Tile_X3Y6_S1BEG),
    .S2MID(Tile_X3Y6_S2BEG),
    .S2END(Tile_X3Y6_S2BEGb),
    .S4END(Tile_X3Y6_S4BEG),
    .SS4END(Tile_X3Y6_SS4BEG),
    .W1END(Tile_X4Y7_W1BEG),
    .W2MID(Tile_X4Y7_W2BEG),
    .W2END(Tile_X4Y7_W2BEGb),
    .WW4END(Tile_X4Y7_WW4BEG),
    .W6END(Tile_X4Y7_W6BEG),
    .N1BEG(Tile_X3Y7_N1BEG),
    .N2BEG(Tile_X3Y7_N2BEG),
    .N2BEGb(Tile_X3Y7_N2BEGb),
    .N4BEG(Tile_X3Y7_N4BEG),
    .NN4BEG(Tile_X3Y7_NN4BEG),
    .E1BEG(Tile_X3Y7_E1BEG),
    .E2BEG(Tile_X3Y7_E2BEG),
    .E2BEGb(Tile_X3Y7_E2BEGb),
    .EE4BEG(Tile_X3Y7_EE4BEG),
    .E6BEG(Tile_X3Y7_E6BEG),
    .S1BEG(Tile_X3Y7_S1BEG),
    .S2BEG(Tile_X3Y7_S2BEG),
    .S2BEGb(Tile_X3Y7_S2BEGb),
    .S4BEG(Tile_X3Y7_S4BEG),
    .SS4BEG(Tile_X3Y7_SS4BEG),
    .W1BEG(Tile_X3Y7_W1BEG),
    .W2BEG(Tile_X3Y7_W2BEG),
    .W2BEGb(Tile_X3Y7_W2BEGb),
    .WW4BEG(Tile_X3Y7_WW4BEG),
    .W6BEG(Tile_X3Y7_W6BEG),
    .Co(Tile_X3Y7_Co),
    .UserCLK(Tile_X3Y8_UserCLKo),
    .UserCLKo(Tile_X3Y7_UserCLKo),
    .FrameData(Tile_X2Y7_FrameData_O),
    .FrameData_O(Tile_X3Y7_FrameData_O),
    .FrameStrobe(Tile_X3Y8_FrameStrobe_O),
    .FrameStrobe_O(Tile_X3Y7_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
RegFile
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X4Y7_Emulate_Bitstream)
    )
`endif
    Tile_X4Y7_RegFile
    (
    .N1END(Tile_X4Y8_N1BEG),
    .N2MID(Tile_X4Y8_N2BEG),
    .N2END(Tile_X4Y8_N2BEGb),
    .N4END(Tile_X4Y8_N4BEG),
    .NN4END(Tile_X4Y8_NN4BEG),
    .E1END(Tile_X3Y7_E1BEG),
    .E2MID(Tile_X3Y7_E2BEG),
    .E2END(Tile_X3Y7_E2BEGb),
    .EE4END(Tile_X3Y7_EE4BEG),
    .E6END(Tile_X3Y7_E6BEG),
    .S1END(Tile_X4Y6_S1BEG),
    .S2MID(Tile_X4Y6_S2BEG),
    .S2END(Tile_X4Y6_S2BEGb),
    .S4END(Tile_X4Y6_S4BEG),
    .SS4END(Tile_X4Y6_SS4BEG),
    .W1END(Tile_X5Y7_W1BEG),
    .W2MID(Tile_X5Y7_W2BEG),
    .W2END(Tile_X5Y7_W2BEGb),
    .WW4END(Tile_X5Y7_WW4BEG),
    .W6END(Tile_X5Y7_W6BEG),
    .N1BEG(Tile_X4Y7_N1BEG),
    .N2BEG(Tile_X4Y7_N2BEG),
    .N2BEGb(Tile_X4Y7_N2BEGb),
    .N4BEG(Tile_X4Y7_N4BEG),
    .NN4BEG(Tile_X4Y7_NN4BEG),
    .E1BEG(Tile_X4Y7_E1BEG),
    .E2BEG(Tile_X4Y7_E2BEG),
    .E2BEGb(Tile_X4Y7_E2BEGb),
    .EE4BEG(Tile_X4Y7_EE4BEG),
    .E6BEG(Tile_X4Y7_E6BEG),
    .S1BEG(Tile_X4Y7_S1BEG),
    .S2BEG(Tile_X4Y7_S2BEG),
    .S2BEGb(Tile_X4Y7_S2BEGb),
    .S4BEG(Tile_X4Y7_S4BEG),
    .SS4BEG(Tile_X4Y7_SS4BEG),
    .W1BEG(Tile_X4Y7_W1BEG),
    .W2BEG(Tile_X4Y7_W2BEG),
    .W2BEGb(Tile_X4Y7_W2BEGb),
    .WW4BEG(Tile_X4Y7_WW4BEG),
    .W6BEG(Tile_X4Y7_W6BEG),
    .UserCLK(Tile_X4Y8_UserCLKo),
    .UserCLKo(Tile_X4Y7_UserCLKo),
    .FrameData(Tile_X3Y7_FrameData_O),
    .FrameData_O(Tile_X4Y7_FrameData_O),
    .FrameStrobe(Tile_X4Y8_FrameStrobe_O),
    .FrameStrobe_O(Tile_X4Y7_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X5Y7_Emulate_Bitstream)
    )
`endif
    Tile_X5Y7_LUT4AB
    (
    .N1END(Tile_X5Y8_N1BEG),
    .N2MID(Tile_X5Y8_N2BEG),
    .N2END(Tile_X5Y8_N2BEGb),
    .N4END(Tile_X5Y8_N4BEG),
    .NN4END(Tile_X5Y8_NN4BEG),
    .Ci(Tile_X5Y8_Co),
    .E1END(Tile_X4Y7_E1BEG),
    .E2MID(Tile_X4Y7_E2BEG),
    .E2END(Tile_X4Y7_E2BEGb),
    .EE4END(Tile_X4Y7_EE4BEG),
    .E6END(Tile_X4Y7_E6BEG),
    .S1END(Tile_X5Y6_S1BEG),
    .S2MID(Tile_X5Y6_S2BEG),
    .S2END(Tile_X5Y6_S2BEGb),
    .S4END(Tile_X5Y6_S4BEG),
    .SS4END(Tile_X5Y6_SS4BEG),
    .W1END(Tile_X6Y7_W1BEG),
    .W2MID(Tile_X6Y7_W2BEG),
    .W2END(Tile_X6Y7_W2BEGb),
    .WW4END(Tile_X6Y7_WW4BEG),
    .W6END(Tile_X6Y7_W6BEG),
    .N1BEG(Tile_X5Y7_N1BEG),
    .N2BEG(Tile_X5Y7_N2BEG),
    .N2BEGb(Tile_X5Y7_N2BEGb),
    .N4BEG(Tile_X5Y7_N4BEG),
    .NN4BEG(Tile_X5Y7_NN4BEG),
    .E1BEG(Tile_X5Y7_E1BEG),
    .E2BEG(Tile_X5Y7_E2BEG),
    .E2BEGb(Tile_X5Y7_E2BEGb),
    .EE4BEG(Tile_X5Y7_EE4BEG),
    .E6BEG(Tile_X5Y7_E6BEG),
    .S1BEG(Tile_X5Y7_S1BEG),
    .S2BEG(Tile_X5Y7_S2BEG),
    .S2BEGb(Tile_X5Y7_S2BEGb),
    .S4BEG(Tile_X5Y7_S4BEG),
    .SS4BEG(Tile_X5Y7_SS4BEG),
    .W1BEG(Tile_X5Y7_W1BEG),
    .W2BEG(Tile_X5Y7_W2BEG),
    .W2BEGb(Tile_X5Y7_W2BEGb),
    .WW4BEG(Tile_X5Y7_WW4BEG),
    .W6BEG(Tile_X5Y7_W6BEG),
    .Co(Tile_X5Y7_Co),
    .UserCLK(Tile_X5Y8_UserCLKo),
    .UserCLKo(Tile_X5Y7_UserCLKo),
    .FrameData(Tile_X4Y7_FrameData_O),
    .FrameData_O(Tile_X5Y7_FrameData_O),
    .FrameStrobe(Tile_X5Y8_FrameStrobe_O),
    .FrameStrobe_O(Tile_X5Y7_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X6Y7_Emulate_Bitstream)
    )
`endif
    Tile_X6Y7_LUT4AB
    (
    .N1END(Tile_X6Y8_N1BEG),
    .N2MID(Tile_X6Y8_N2BEG),
    .N2END(Tile_X6Y8_N2BEGb),
    .N4END(Tile_X6Y8_N4BEG),
    .NN4END(Tile_X6Y8_NN4BEG),
    .Ci(Tile_X6Y8_Co),
    .E1END(Tile_X5Y7_E1BEG),
    .E2MID(Tile_X5Y7_E2BEG),
    .E2END(Tile_X5Y7_E2BEGb),
    .EE4END(Tile_X5Y7_EE4BEG),
    .E6END(Tile_X5Y7_E6BEG),
    .S1END(Tile_X6Y6_S1BEG),
    .S2MID(Tile_X6Y6_S2BEG),
    .S2END(Tile_X6Y6_S2BEGb),
    .S4END(Tile_X6Y6_S4BEG),
    .SS4END(Tile_X6Y6_SS4BEG),
    .W1END(Tile_X7Y7_W1BEG),
    .W2MID(Tile_X7Y7_W2BEG),
    .W2END(Tile_X7Y7_W2BEGb),
    .WW4END(Tile_X7Y7_WW4BEG),
    .W6END(Tile_X7Y7_W6BEG),
    .N1BEG(Tile_X6Y7_N1BEG),
    .N2BEG(Tile_X6Y7_N2BEG),
    .N2BEGb(Tile_X6Y7_N2BEGb),
    .N4BEG(Tile_X6Y7_N4BEG),
    .NN4BEG(Tile_X6Y7_NN4BEG),
    .E1BEG(Tile_X6Y7_E1BEG),
    .E2BEG(Tile_X6Y7_E2BEG),
    .E2BEGb(Tile_X6Y7_E2BEGb),
    .EE4BEG(Tile_X6Y7_EE4BEG),
    .E6BEG(Tile_X6Y7_E6BEG),
    .S1BEG(Tile_X6Y7_S1BEG),
    .S2BEG(Tile_X6Y7_S2BEG),
    .S2BEGb(Tile_X6Y7_S2BEGb),
    .S4BEG(Tile_X6Y7_S4BEG),
    .SS4BEG(Tile_X6Y7_SS4BEG),
    .W1BEG(Tile_X6Y7_W1BEG),
    .W2BEG(Tile_X6Y7_W2BEG),
    .W2BEGb(Tile_X6Y7_W2BEGb),
    .WW4BEG(Tile_X6Y7_WW4BEG),
    .W6BEG(Tile_X6Y7_W6BEG),
    .Co(Tile_X6Y7_Co),
    .UserCLK(Tile_X6Y8_UserCLKo),
    .UserCLKo(Tile_X6Y7_UserCLKo),
    .FrameData(Tile_X5Y7_FrameData_O),
    .FrameData_O(Tile_X6Y7_FrameData_O),
    .FrameStrobe(Tile_X6Y8_FrameStrobe_O),
    .FrameStrobe_O(Tile_X6Y7_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
DSP
`ifdef EMULATION
    #(
    .Tile_X0Y0_Emulate_Bitstream(`Tile_X7Y7_Emulate_Bitstream),
    .Tile_X0Y1_Emulate_Bitstream(`Tile_X7Y8_Emulate_Bitstream)
    )
`endif
    Tile_X7Y7_DSP
    (
    .Tile_X0Y0_E1END(Tile_X6Y7_E1BEG),
    .Tile_X0Y0_E2MID(Tile_X6Y7_E2BEG),
    .Tile_X0Y0_E2END(Tile_X6Y7_E2BEGb),
    .Tile_X0Y0_EE4END(Tile_X6Y7_EE4BEG),
    .Tile_X0Y0_E6END(Tile_X6Y7_E6BEG),
    .Tile_X0Y0_S1END(Tile_X7Y6_S1BEG),
    .Tile_X0Y0_S2MID(Tile_X7Y6_S2BEG),
    .Tile_X0Y0_S2END(Tile_X7Y6_S2BEGb),
    .Tile_X0Y0_S4END(Tile_X7Y6_S4BEG),
    .Tile_X0Y0_SS4END(Tile_X7Y6_SS4BEG),
    .Tile_X0Y0_W1END(Tile_X8Y7_W1BEG),
    .Tile_X0Y0_W2MID(Tile_X8Y7_W2BEG),
    .Tile_X0Y0_W2END(Tile_X8Y7_W2BEGb),
    .Tile_X0Y0_WW4END(Tile_X8Y7_WW4BEG),
    .Tile_X0Y0_W6END(Tile_X8Y7_W6BEG),
    .Tile_X0Y1_N1END(Tile_X7Y9_N1BEG),
    .Tile_X0Y1_N2MID(Tile_X7Y9_N2BEG),
    .Tile_X0Y1_N2END(Tile_X7Y9_N2BEGb),
    .Tile_X0Y1_N4END(Tile_X7Y9_N4BEG),
    .Tile_X0Y1_NN4END(Tile_X7Y9_NN4BEG),
    .Tile_X0Y1_E1END(Tile_X6Y8_E1BEG),
    .Tile_X0Y1_E2MID(Tile_X6Y8_E2BEG),
    .Tile_X0Y1_E2END(Tile_X6Y8_E2BEGb),
    .Tile_X0Y1_EE4END(Tile_X6Y8_EE4BEG),
    .Tile_X0Y1_E6END(Tile_X6Y8_E6BEG),
    .Tile_X0Y1_W1END(Tile_X8Y8_W1BEG),
    .Tile_X0Y1_W2MID(Tile_X8Y8_W2BEG),
    .Tile_X0Y1_W2END(Tile_X8Y8_W2BEGb),
    .Tile_X0Y1_WW4END(Tile_X8Y8_WW4BEG),
    .Tile_X0Y1_W6END(Tile_X8Y8_W6BEG),
    .Tile_X0Y0_N1BEG(Tile_X7Y7_N1BEG),
    .Tile_X0Y0_N2BEG(Tile_X7Y7_N2BEG),
    .Tile_X0Y0_N2BEGb(Tile_X7Y7_N2BEGb),
    .Tile_X0Y0_N4BEG(Tile_X7Y7_N4BEG),
    .Tile_X0Y0_NN4BEG(Tile_X7Y7_NN4BEG),
    .Tile_X0Y0_E1BEG(Tile_X7Y7_E1BEG),
    .Tile_X0Y0_E2BEG(Tile_X7Y7_E2BEG),
    .Tile_X0Y0_E2BEGb(Tile_X7Y7_E2BEGb),
    .Tile_X0Y0_EE4BEG(Tile_X7Y7_EE4BEG),
    .Tile_X0Y0_E6BEG(Tile_X7Y7_E6BEG),
    .Tile_X0Y0_W1BEG(Tile_X7Y7_W1BEG),
    .Tile_X0Y0_W2BEG(Tile_X7Y7_W2BEG),
    .Tile_X0Y0_W2BEGb(Tile_X7Y7_W2BEGb),
    .Tile_X0Y0_WW4BEG(Tile_X7Y7_WW4BEG),
    .Tile_X0Y0_W6BEG(Tile_X7Y7_W6BEG),
    .Tile_X0Y1_E1BEG(Tile_X7Y8_E1BEG),
    .Tile_X0Y1_E2BEG(Tile_X7Y8_E2BEG),
    .Tile_X0Y1_E2BEGb(Tile_X7Y8_E2BEGb),
    .Tile_X0Y1_EE4BEG(Tile_X7Y8_EE4BEG),
    .Tile_X0Y1_E6BEG(Tile_X7Y8_E6BEG),
    .Tile_X0Y1_S1BEG(Tile_X7Y8_S1BEG),
    .Tile_X0Y1_S2BEG(Tile_X7Y8_S2BEG),
    .Tile_X0Y1_S2BEGb(Tile_X7Y8_S2BEGb),
    .Tile_X0Y1_S4BEG(Tile_X7Y8_S4BEG),
    .Tile_X0Y1_SS4BEG(Tile_X7Y8_SS4BEG),
    .Tile_X0Y1_W1BEG(Tile_X7Y8_W1BEG),
    .Tile_X0Y1_W2BEG(Tile_X7Y8_W2BEG),
    .Tile_X0Y1_W2BEGb(Tile_X7Y8_W2BEGb),
    .Tile_X0Y1_WW4BEG(Tile_X7Y8_WW4BEG),
    .Tile_X0Y1_W6BEG(Tile_X7Y8_W6BEG),
    .Tile_X0Y0_UserCLKo(Tile_X7Y7_UserCLKo),
    .Tile_X0Y1_UserCLK(Tile_X7Y9_UserCLKo),
    .Tile_X0Y0_FrameData(Tile_X6Y7_FrameData_O),
    .Tile_X0Y0_FrameData_O(Tile_X7Y7_FrameData_O),
    .Tile_X0Y0_FrameStrobe_O(Tile_X7Y7_FrameStrobe_O),
    .Tile_X0Y1_FrameData(Tile_X6Y8_FrameData_O),
    .Tile_X0Y1_FrameData_O(Tile_X7Y8_FrameData_O),
    .Tile_X0Y1_FrameStrobe(Tile_X7Y9_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X8Y7_Emulate_Bitstream)
    )
`endif
    Tile_X8Y7_LUT4AB
    (
    .N1END(Tile_X8Y8_N1BEG),
    .N2MID(Tile_X8Y8_N2BEG),
    .N2END(Tile_X8Y8_N2BEGb),
    .N4END(Tile_X8Y8_N4BEG),
    .NN4END(Tile_X8Y8_NN4BEG),
    .Ci(Tile_X8Y8_Co),
    .E1END(Tile_X7Y7_E1BEG),
    .E2MID(Tile_X7Y7_E2BEG),
    .E2END(Tile_X7Y7_E2BEGb),
    .EE4END(Tile_X7Y7_EE4BEG),
    .E6END(Tile_X7Y7_E6BEG),
    .S1END(Tile_X8Y6_S1BEG),
    .S2MID(Tile_X8Y6_S2BEG),
    .S2END(Tile_X8Y6_S2BEGb),
    .S4END(Tile_X8Y6_S4BEG),
    .SS4END(Tile_X8Y6_SS4BEG),
    .W1END(Tile_X9Y7_W1BEG),
    .W2MID(Tile_X9Y7_W2BEG),
    .W2END(Tile_X9Y7_W2BEGb),
    .WW4END(Tile_X9Y7_WW4BEG),
    .W6END(Tile_X9Y7_W6BEG),
    .N1BEG(Tile_X8Y7_N1BEG),
    .N2BEG(Tile_X8Y7_N2BEG),
    .N2BEGb(Tile_X8Y7_N2BEGb),
    .N4BEG(Tile_X8Y7_N4BEG),
    .NN4BEG(Tile_X8Y7_NN4BEG),
    .E1BEG(Tile_X8Y7_E1BEG),
    .E2BEG(Tile_X8Y7_E2BEG),
    .E2BEGb(Tile_X8Y7_E2BEGb),
    .EE4BEG(Tile_X8Y7_EE4BEG),
    .E6BEG(Tile_X8Y7_E6BEG),
    .S1BEG(Tile_X8Y7_S1BEG),
    .S2BEG(Tile_X8Y7_S2BEG),
    .S2BEGb(Tile_X8Y7_S2BEGb),
    .S4BEG(Tile_X8Y7_S4BEG),
    .SS4BEG(Tile_X8Y7_SS4BEG),
    .W1BEG(Tile_X8Y7_W1BEG),
    .W2BEG(Tile_X8Y7_W2BEG),
    .W2BEGb(Tile_X8Y7_W2BEGb),
    .WW4BEG(Tile_X8Y7_WW4BEG),
    .W6BEG(Tile_X8Y7_W6BEG),
    .Co(Tile_X8Y7_Co),
    .UserCLK(Tile_X8Y8_UserCLKo),
    .UserCLKo(Tile_X8Y7_UserCLKo),
    .FrameData(Tile_X7Y7_FrameData_O),
    .FrameData_O(Tile_X8Y7_FrameData_O),
    .FrameStrobe(Tile_X8Y8_FrameStrobe_O),
    .FrameStrobe_O(Tile_X8Y7_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X9Y7_Emulate_Bitstream)
    )
`endif
    Tile_X9Y7_LUT4AB
    (
    .N1END(Tile_X9Y8_N1BEG),
    .N2MID(Tile_X9Y8_N2BEG),
    .N2END(Tile_X9Y8_N2BEGb),
    .N4END(Tile_X9Y8_N4BEG),
    .NN4END(Tile_X9Y8_NN4BEG),
    .Ci(Tile_X9Y8_Co),
    .E1END(Tile_X8Y7_E1BEG),
    .E2MID(Tile_X8Y7_E2BEG),
    .E2END(Tile_X8Y7_E2BEGb),
    .EE4END(Tile_X8Y7_EE4BEG),
    .E6END(Tile_X8Y7_E6BEG),
    .S1END(Tile_X9Y6_S1BEG),
    .S2MID(Tile_X9Y6_S2BEG),
    .S2END(Tile_X9Y6_S2BEGb),
    .S4END(Tile_X9Y6_S4BEG),
    .SS4END(Tile_X9Y6_SS4BEG),
    .W1END(Tile_X10Y7_W1BEG),
    .W2MID(Tile_X10Y7_W2BEG),
    .W2END(Tile_X10Y7_W2BEGb),
    .WW4END(Tile_X10Y7_WW4BEG),
    .W6END(Tile_X10Y7_W6BEG),
    .N1BEG(Tile_X9Y7_N1BEG),
    .N2BEG(Tile_X9Y7_N2BEG),
    .N2BEGb(Tile_X9Y7_N2BEGb),
    .N4BEG(Tile_X9Y7_N4BEG),
    .NN4BEG(Tile_X9Y7_NN4BEG),
    .E1BEG(Tile_X9Y7_E1BEG),
    .E2BEG(Tile_X9Y7_E2BEG),
    .E2BEGb(Tile_X9Y7_E2BEGb),
    .EE4BEG(Tile_X9Y7_EE4BEG),
    .E6BEG(Tile_X9Y7_E6BEG),
    .S1BEG(Tile_X9Y7_S1BEG),
    .S2BEG(Tile_X9Y7_S2BEG),
    .S2BEGb(Tile_X9Y7_S2BEGb),
    .S4BEG(Tile_X9Y7_S4BEG),
    .SS4BEG(Tile_X9Y7_SS4BEG),
    .W1BEG(Tile_X9Y7_W1BEG),
    .W2BEG(Tile_X9Y7_W2BEG),
    .W2BEGb(Tile_X9Y7_W2BEGb),
    .WW4BEG(Tile_X9Y7_WW4BEG),
    .W6BEG(Tile_X9Y7_W6BEG),
    .Co(Tile_X9Y7_Co),
    .UserCLK(Tile_X9Y8_UserCLKo),
    .UserCLKo(Tile_X9Y7_UserCLKo),
    .FrameData(Tile_X8Y7_FrameData_O),
    .FrameData_O(Tile_X9Y7_FrameData_O),
    .FrameStrobe(Tile_X9Y8_FrameStrobe_O),
    .FrameStrobe_O(Tile_X9Y7_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
IHP_SRAM
`ifdef EMULATION
    #(
    .Tile_X0Y0_Emulate_Bitstream(`Tile_X10Y7_Emulate_Bitstream),
    .Tile_X0Y1_Emulate_Bitstream(`Tile_X10Y8_Emulate_Bitstream)
    )
`endif
    Tile_X10Y7_IHP_SRAM
    (
    .Tile_X0Y0_E1END(Tile_X9Y7_E1BEG),
    .Tile_X0Y0_E2MID(Tile_X9Y7_E2BEG),
    .Tile_X0Y0_E2END(Tile_X9Y7_E2BEGb),
    .Tile_X0Y0_EE4END(Tile_X9Y7_EE4BEG),
    .Tile_X0Y0_E6END(Tile_X9Y7_E6BEG),
    .Tile_X0Y0_S1END(Tile_X10Y6_S1BEG),
    .Tile_X0Y0_S2MID(Tile_X10Y6_S2BEG),
    .Tile_X0Y0_S2END(Tile_X10Y6_S2BEGb),
    .Tile_X0Y0_S4END(Tile_X10Y6_S4BEG),
    .Tile_X0Y1_N1END(Tile_X10Y9_N1BEG),
    .Tile_X0Y1_N2MID(Tile_X10Y9_N2BEG),
    .Tile_X0Y1_N2END(Tile_X10Y9_N2BEGb),
    .Tile_X0Y1_N4END(Tile_X10Y9_N4BEG),
    .Tile_X0Y1_E1END(Tile_X9Y8_E1BEG),
    .Tile_X0Y1_E2MID(Tile_X9Y8_E2BEG),
    .Tile_X0Y1_E2END(Tile_X9Y8_E2BEGb),
    .Tile_X0Y1_EE4END(Tile_X9Y8_EE4BEG),
    .Tile_X0Y1_E6END(Tile_X9Y8_E6BEG),
    .Tile_X0Y0_N1BEG(Tile_X10Y7_N1BEG),
    .Tile_X0Y0_N2BEG(Tile_X10Y7_N2BEG),
    .Tile_X0Y0_N2BEGb(Tile_X10Y7_N2BEGb),
    .Tile_X0Y0_N4BEG(Tile_X10Y7_N4BEG),
    .Tile_X0Y0_W1BEG(Tile_X10Y7_W1BEG),
    .Tile_X0Y0_W2BEG(Tile_X10Y7_W2BEG),
    .Tile_X0Y0_W2BEGb(Tile_X10Y7_W2BEGb),
    .Tile_X0Y0_WW4BEG(Tile_X10Y7_WW4BEG),
    .Tile_X0Y0_W6BEG(Tile_X10Y7_W6BEG),
    .Tile_X0Y1_S1BEG(Tile_X10Y8_S1BEG),
    .Tile_X0Y1_S2BEG(Tile_X10Y8_S2BEG),
    .Tile_X0Y1_S2BEGb(Tile_X10Y8_S2BEGb),
    .Tile_X0Y1_S4BEG(Tile_X10Y8_S4BEG),
    .Tile_X0Y1_W1BEG(Tile_X10Y8_W1BEG),
    .Tile_X0Y1_W2BEG(Tile_X10Y8_W2BEG),
    .Tile_X0Y1_W2BEGb(Tile_X10Y8_W2BEGb),
    .Tile_X0Y1_WW4BEG(Tile_X10Y8_WW4BEG),
    .Tile_X0Y1_W6BEG(Tile_X10Y8_W6BEG),
    .CONFIGURED_top(Tile_X10Y8_CONFIGURED_top),
    .DOUT_SRAM0(Tile_X10Y8_DOUT_SRAM0),
    .DOUT_SRAM1(Tile_X10Y8_DOUT_SRAM1),
    .DOUT_SRAM2(Tile_X10Y8_DOUT_SRAM2),
    .DOUT_SRAM3(Tile_X10Y8_DOUT_SRAM3),
    .DOUT_SRAM4(Tile_X10Y8_DOUT_SRAM4),
    .DOUT_SRAM5(Tile_X10Y8_DOUT_SRAM5),
    .DOUT_SRAM6(Tile_X10Y8_DOUT_SRAM6),
    .DOUT_SRAM7(Tile_X10Y8_DOUT_SRAM7),
    .DOUT_SRAM8(Tile_X10Y8_DOUT_SRAM8),
    .DOUT_SRAM9(Tile_X10Y8_DOUT_SRAM9),
    .DOUT_SRAM10(Tile_X10Y8_DOUT_SRAM10),
    .DOUT_SRAM11(Tile_X10Y8_DOUT_SRAM11),
    .DOUT_SRAM12(Tile_X10Y8_DOUT_SRAM12),
    .DOUT_SRAM13(Tile_X10Y8_DOUT_SRAM13),
    .DOUT_SRAM14(Tile_X10Y8_DOUT_SRAM14),
    .DOUT_SRAM15(Tile_X10Y8_DOUT_SRAM15),
    .DOUT_SRAM16(Tile_X10Y8_DOUT_SRAM16),
    .DOUT_SRAM17(Tile_X10Y8_DOUT_SRAM17),
    .DOUT_SRAM18(Tile_X10Y8_DOUT_SRAM18),
    .DOUT_SRAM19(Tile_X10Y8_DOUT_SRAM19),
    .DOUT_SRAM20(Tile_X10Y8_DOUT_SRAM20),
    .DOUT_SRAM21(Tile_X10Y8_DOUT_SRAM21),
    .DOUT_SRAM22(Tile_X10Y8_DOUT_SRAM22),
    .DOUT_SRAM23(Tile_X10Y8_DOUT_SRAM23),
    .DOUT_SRAM24(Tile_X10Y8_DOUT_SRAM24),
    .DOUT_SRAM25(Tile_X10Y8_DOUT_SRAM25),
    .DOUT_SRAM26(Tile_X10Y8_DOUT_SRAM26),
    .DOUT_SRAM27(Tile_X10Y8_DOUT_SRAM27),
    .DOUT_SRAM28(Tile_X10Y8_DOUT_SRAM28),
    .DOUT_SRAM29(Tile_X10Y8_DOUT_SRAM29),
    .DOUT_SRAM30(Tile_X10Y8_DOUT_SRAM30),
    .DOUT_SRAM31(Tile_X10Y8_DOUT_SRAM31),
    .ADDR_SRAM0(Tile_X10Y8_ADDR_SRAM0),
    .ADDR_SRAM1(Tile_X10Y8_ADDR_SRAM1),
    .ADDR_SRAM2(Tile_X10Y8_ADDR_SRAM2),
    .ADDR_SRAM3(Tile_X10Y8_ADDR_SRAM3),
    .ADDR_SRAM4(Tile_X10Y8_ADDR_SRAM4),
    .ADDR_SRAM5(Tile_X10Y8_ADDR_SRAM5),
    .ADDR_SRAM6(Tile_X10Y8_ADDR_SRAM6),
    .ADDR_SRAM7(Tile_X10Y8_ADDR_SRAM7),
    .ADDR_SRAM8(Tile_X10Y8_ADDR_SRAM8),
    .ADDR_SRAM9(Tile_X10Y8_ADDR_SRAM9),
    .BM_SRAM0(Tile_X10Y8_BM_SRAM0),
    .BM_SRAM1(Tile_X10Y8_BM_SRAM1),
    .BM_SRAM2(Tile_X10Y8_BM_SRAM2),
    .BM_SRAM3(Tile_X10Y8_BM_SRAM3),
    .BM_SRAM4(Tile_X10Y8_BM_SRAM4),
    .BM_SRAM5(Tile_X10Y8_BM_SRAM5),
    .BM_SRAM6(Tile_X10Y8_BM_SRAM6),
    .BM_SRAM7(Tile_X10Y8_BM_SRAM7),
    .BM_SRAM8(Tile_X10Y8_BM_SRAM8),
    .BM_SRAM9(Tile_X10Y8_BM_SRAM9),
    .BM_SRAM10(Tile_X10Y8_BM_SRAM10),
    .BM_SRAM11(Tile_X10Y8_BM_SRAM11),
    .BM_SRAM12(Tile_X10Y8_BM_SRAM12),
    .BM_SRAM13(Tile_X10Y8_BM_SRAM13),
    .BM_SRAM14(Tile_X10Y8_BM_SRAM14),
    .BM_SRAM15(Tile_X10Y8_BM_SRAM15),
    .BM_SRAM16(Tile_X10Y8_BM_SRAM16),
    .BM_SRAM17(Tile_X10Y8_BM_SRAM17),
    .BM_SRAM18(Tile_X10Y8_BM_SRAM18),
    .BM_SRAM19(Tile_X10Y8_BM_SRAM19),
    .BM_SRAM20(Tile_X10Y8_BM_SRAM20),
    .BM_SRAM21(Tile_X10Y8_BM_SRAM21),
    .BM_SRAM22(Tile_X10Y8_BM_SRAM22),
    .BM_SRAM23(Tile_X10Y8_BM_SRAM23),
    .BM_SRAM24(Tile_X10Y8_BM_SRAM24),
    .BM_SRAM25(Tile_X10Y8_BM_SRAM25),
    .BM_SRAM26(Tile_X10Y8_BM_SRAM26),
    .BM_SRAM27(Tile_X10Y8_BM_SRAM27),
    .BM_SRAM28(Tile_X10Y8_BM_SRAM28),
    .BM_SRAM29(Tile_X10Y8_BM_SRAM29),
    .BM_SRAM30(Tile_X10Y8_BM_SRAM30),
    .BM_SRAM31(Tile_X10Y8_BM_SRAM31),
    .CLK_SRAM(Tile_X10Y8_CLK_SRAM),
    .DIN_SRAM0(Tile_X10Y8_DIN_SRAM0),
    .DIN_SRAM1(Tile_X10Y8_DIN_SRAM1),
    .DIN_SRAM2(Tile_X10Y8_DIN_SRAM2),
    .DIN_SRAM3(Tile_X10Y8_DIN_SRAM3),
    .DIN_SRAM4(Tile_X10Y8_DIN_SRAM4),
    .DIN_SRAM5(Tile_X10Y8_DIN_SRAM5),
    .DIN_SRAM6(Tile_X10Y8_DIN_SRAM6),
    .DIN_SRAM7(Tile_X10Y8_DIN_SRAM7),
    .DIN_SRAM8(Tile_X10Y8_DIN_SRAM8),
    .DIN_SRAM9(Tile_X10Y8_DIN_SRAM9),
    .DIN_SRAM10(Tile_X10Y8_DIN_SRAM10),
    .DIN_SRAM11(Tile_X10Y8_DIN_SRAM11),
    .DIN_SRAM12(Tile_X10Y8_DIN_SRAM12),
    .DIN_SRAM13(Tile_X10Y8_DIN_SRAM13),
    .DIN_SRAM14(Tile_X10Y8_DIN_SRAM14),
    .DIN_SRAM15(Tile_X10Y8_DIN_SRAM15),
    .DIN_SRAM16(Tile_X10Y8_DIN_SRAM16),
    .DIN_SRAM17(Tile_X10Y8_DIN_SRAM17),
    .DIN_SRAM18(Tile_X10Y8_DIN_SRAM18),
    .DIN_SRAM19(Tile_X10Y8_DIN_SRAM19),
    .DIN_SRAM20(Tile_X10Y8_DIN_SRAM20),
    .DIN_SRAM21(Tile_X10Y8_DIN_SRAM21),
    .DIN_SRAM22(Tile_X10Y8_DIN_SRAM22),
    .DIN_SRAM23(Tile_X10Y8_DIN_SRAM23),
    .DIN_SRAM24(Tile_X10Y8_DIN_SRAM24),
    .DIN_SRAM25(Tile_X10Y8_DIN_SRAM25),
    .DIN_SRAM26(Tile_X10Y8_DIN_SRAM26),
    .DIN_SRAM27(Tile_X10Y8_DIN_SRAM27),
    .DIN_SRAM28(Tile_X10Y8_DIN_SRAM28),
    .DIN_SRAM29(Tile_X10Y8_DIN_SRAM29),
    .DIN_SRAM30(Tile_X10Y8_DIN_SRAM30),
    .DIN_SRAM31(Tile_X10Y8_DIN_SRAM31),
    .MEN_SRAM(Tile_X10Y8_MEN_SRAM),
    .REN_SRAM(Tile_X10Y8_REN_SRAM),
    .TIE_HIGH_SRAM(Tile_X10Y8_TIE_HIGH_SRAM),
    .TIE_LOW_SRAM(Tile_X10Y8_TIE_LOW_SRAM),
    .WEN_SRAM(Tile_X10Y8_WEN_SRAM),
    .Tile_X0Y0_UserCLKo(Tile_X10Y7_UserCLKo),
    .Tile_X0Y1_UserCLK(Tile_X10Y9_UserCLKo),
    .Tile_X0Y0_FrameData(Tile_X9Y7_FrameData_O),
    .Tile_X0Y0_FrameData_O(Tile_X10Y7_FrameData_O),
    .Tile_X0Y0_FrameStrobe_O(Tile_X10Y7_FrameStrobe_O),
    .Tile_X0Y1_FrameData(Tile_X9Y8_FrameData_O),
    .Tile_X0Y1_FrameData_O(Tile_X10Y8_FrameData_O),
    .Tile_X0Y1_FrameStrobe(Tile_X10Y9_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
W_IO
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X0Y8_Emulate_Bitstream)
    )
`endif
    Tile_X0Y8_W_IO
    (
    .W1END(Tile_X1Y8_W1BEG),
    .W2MID(Tile_X1Y8_W2BEG),
    .W2END(Tile_X1Y8_W2BEGb),
    .WW4END(Tile_X1Y8_WW4BEG),
    .W6END(Tile_X1Y8_W6BEG),
    .E1BEG(Tile_X0Y8_E1BEG),
    .E2BEG(Tile_X0Y8_E2BEG),
    .E2BEGb(Tile_X0Y8_E2BEGb),
    .EE4BEG(Tile_X0Y8_EE4BEG),
    .E6BEG(Tile_X0Y8_E6BEG),
    .A_O_top(Tile_X0Y8_A_O_top),
    .A_I_top(Tile_X0Y8_A_I_top),
    .A_T_top(Tile_X0Y8_A_T_top),
    .B_O_top(Tile_X0Y8_B_O_top),
    .B_I_top(Tile_X0Y8_B_I_top),
    .B_T_top(Tile_X0Y8_B_T_top),
    .A_config_C_bit0(Tile_X0Y8_A_config_C_bit0),
    .A_config_C_bit1(Tile_X0Y8_A_config_C_bit1),
    .A_config_C_bit2(Tile_X0Y8_A_config_C_bit2),
    .A_config_C_bit3(Tile_X0Y8_A_config_C_bit3),
    .B_config_C_bit0(Tile_X0Y8_B_config_C_bit0),
    .B_config_C_bit1(Tile_X0Y8_B_config_C_bit1),
    .B_config_C_bit2(Tile_X0Y8_B_config_C_bit2),
    .B_config_C_bit3(Tile_X0Y8_B_config_C_bit3),
    .UserCLK(Tile_X0Y9_UserCLKo),
    .UserCLKo(Tile_X0Y8_UserCLKo),
    .FrameData(Row_Y8_FrameData),
    .FrameData_O(Tile_X0Y8_FrameData_O),
    .FrameStrobe(Tile_X0Y9_FrameStrobe_O),
    .FrameStrobe_O(Tile_X0Y8_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X1Y8_Emulate_Bitstream)
    )
`endif
    Tile_X1Y8_LUT4AB
    (
    .N1END(Tile_X1Y9_N1BEG),
    .N2MID(Tile_X1Y9_N2BEG),
    .N2END(Tile_X1Y9_N2BEGb),
    .N4END(Tile_X1Y9_N4BEG),
    .NN4END(Tile_X1Y9_NN4BEG),
    .Ci(Tile_X1Y9_Co),
    .E1END(Tile_X0Y8_E1BEG),
    .E2MID(Tile_X0Y8_E2BEG),
    .E2END(Tile_X0Y8_E2BEGb),
    .EE4END(Tile_X0Y8_EE4BEG),
    .E6END(Tile_X0Y8_E6BEG),
    .S1END(Tile_X1Y7_S1BEG),
    .S2MID(Tile_X1Y7_S2BEG),
    .S2END(Tile_X1Y7_S2BEGb),
    .S4END(Tile_X1Y7_S4BEG),
    .SS4END(Tile_X1Y7_SS4BEG),
    .W1END(Tile_X2Y8_W1BEG),
    .W2MID(Tile_X2Y8_W2BEG),
    .W2END(Tile_X2Y8_W2BEGb),
    .WW4END(Tile_X2Y8_WW4BEG),
    .W6END(Tile_X2Y8_W6BEG),
    .N1BEG(Tile_X1Y8_N1BEG),
    .N2BEG(Tile_X1Y8_N2BEG),
    .N2BEGb(Tile_X1Y8_N2BEGb),
    .N4BEG(Tile_X1Y8_N4BEG),
    .NN4BEG(Tile_X1Y8_NN4BEG),
    .E1BEG(Tile_X1Y8_E1BEG),
    .E2BEG(Tile_X1Y8_E2BEG),
    .E2BEGb(Tile_X1Y8_E2BEGb),
    .EE4BEG(Tile_X1Y8_EE4BEG),
    .E6BEG(Tile_X1Y8_E6BEG),
    .S1BEG(Tile_X1Y8_S1BEG),
    .S2BEG(Tile_X1Y8_S2BEG),
    .S2BEGb(Tile_X1Y8_S2BEGb),
    .S4BEG(Tile_X1Y8_S4BEG),
    .SS4BEG(Tile_X1Y8_SS4BEG),
    .W1BEG(Tile_X1Y8_W1BEG),
    .W2BEG(Tile_X1Y8_W2BEG),
    .W2BEGb(Tile_X1Y8_W2BEGb),
    .WW4BEG(Tile_X1Y8_WW4BEG),
    .W6BEG(Tile_X1Y8_W6BEG),
    .Co(Tile_X1Y8_Co),
    .UserCLK(Tile_X1Y9_UserCLKo),
    .UserCLKo(Tile_X1Y8_UserCLKo),
    .FrameData(Tile_X0Y8_FrameData_O),
    .FrameData_O(Tile_X1Y8_FrameData_O),
    .FrameStrobe(Tile_X1Y9_FrameStrobe_O),
    .FrameStrobe_O(Tile_X1Y8_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X2Y8_Emulate_Bitstream)
    )
`endif
    Tile_X2Y8_LUT4AB
    (
    .N1END(Tile_X2Y9_N1BEG),
    .N2MID(Tile_X2Y9_N2BEG),
    .N2END(Tile_X2Y9_N2BEGb),
    .N4END(Tile_X2Y9_N4BEG),
    .NN4END(Tile_X2Y9_NN4BEG),
    .Ci(Tile_X2Y9_Co),
    .E1END(Tile_X1Y8_E1BEG),
    .E2MID(Tile_X1Y8_E2BEG),
    .E2END(Tile_X1Y8_E2BEGb),
    .EE4END(Tile_X1Y8_EE4BEG),
    .E6END(Tile_X1Y8_E6BEG),
    .S1END(Tile_X2Y7_S1BEG),
    .S2MID(Tile_X2Y7_S2BEG),
    .S2END(Tile_X2Y7_S2BEGb),
    .S4END(Tile_X2Y7_S4BEG),
    .SS4END(Tile_X2Y7_SS4BEG),
    .W1END(Tile_X3Y8_W1BEG),
    .W2MID(Tile_X3Y8_W2BEG),
    .W2END(Tile_X3Y8_W2BEGb),
    .WW4END(Tile_X3Y8_WW4BEG),
    .W6END(Tile_X3Y8_W6BEG),
    .N1BEG(Tile_X2Y8_N1BEG),
    .N2BEG(Tile_X2Y8_N2BEG),
    .N2BEGb(Tile_X2Y8_N2BEGb),
    .N4BEG(Tile_X2Y8_N4BEG),
    .NN4BEG(Tile_X2Y8_NN4BEG),
    .E1BEG(Tile_X2Y8_E1BEG),
    .E2BEG(Tile_X2Y8_E2BEG),
    .E2BEGb(Tile_X2Y8_E2BEGb),
    .EE4BEG(Tile_X2Y8_EE4BEG),
    .E6BEG(Tile_X2Y8_E6BEG),
    .S1BEG(Tile_X2Y8_S1BEG),
    .S2BEG(Tile_X2Y8_S2BEG),
    .S2BEGb(Tile_X2Y8_S2BEGb),
    .S4BEG(Tile_X2Y8_S4BEG),
    .SS4BEG(Tile_X2Y8_SS4BEG),
    .W1BEG(Tile_X2Y8_W1BEG),
    .W2BEG(Tile_X2Y8_W2BEG),
    .W2BEGb(Tile_X2Y8_W2BEGb),
    .WW4BEG(Tile_X2Y8_WW4BEG),
    .W6BEG(Tile_X2Y8_W6BEG),
    .Co(Tile_X2Y8_Co),
    .UserCLK(Tile_X2Y9_UserCLKo),
    .UserCLKo(Tile_X2Y8_UserCLKo),
    .FrameData(Tile_X1Y8_FrameData_O),
    .FrameData_O(Tile_X2Y8_FrameData_O),
    .FrameStrobe(Tile_X2Y9_FrameStrobe_O),
    .FrameStrobe_O(Tile_X2Y8_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X3Y8_Emulate_Bitstream)
    )
`endif
    Tile_X3Y8_LUT4AB
    (
    .N1END(Tile_X3Y9_N1BEG),
    .N2MID(Tile_X3Y9_N2BEG),
    .N2END(Tile_X3Y9_N2BEGb),
    .N4END(Tile_X3Y9_N4BEG),
    .NN4END(Tile_X3Y9_NN4BEG),
    .Ci(Tile_X3Y9_Co),
    .E1END(Tile_X2Y8_E1BEG),
    .E2MID(Tile_X2Y8_E2BEG),
    .E2END(Tile_X2Y8_E2BEGb),
    .EE4END(Tile_X2Y8_EE4BEG),
    .E6END(Tile_X2Y8_E6BEG),
    .S1END(Tile_X3Y7_S1BEG),
    .S2MID(Tile_X3Y7_S2BEG),
    .S2END(Tile_X3Y7_S2BEGb),
    .S4END(Tile_X3Y7_S4BEG),
    .SS4END(Tile_X3Y7_SS4BEG),
    .W1END(Tile_X4Y8_W1BEG),
    .W2MID(Tile_X4Y8_W2BEG),
    .W2END(Tile_X4Y8_W2BEGb),
    .WW4END(Tile_X4Y8_WW4BEG),
    .W6END(Tile_X4Y8_W6BEG),
    .N1BEG(Tile_X3Y8_N1BEG),
    .N2BEG(Tile_X3Y8_N2BEG),
    .N2BEGb(Tile_X3Y8_N2BEGb),
    .N4BEG(Tile_X3Y8_N4BEG),
    .NN4BEG(Tile_X3Y8_NN4BEG),
    .E1BEG(Tile_X3Y8_E1BEG),
    .E2BEG(Tile_X3Y8_E2BEG),
    .E2BEGb(Tile_X3Y8_E2BEGb),
    .EE4BEG(Tile_X3Y8_EE4BEG),
    .E6BEG(Tile_X3Y8_E6BEG),
    .S1BEG(Tile_X3Y8_S1BEG),
    .S2BEG(Tile_X3Y8_S2BEG),
    .S2BEGb(Tile_X3Y8_S2BEGb),
    .S4BEG(Tile_X3Y8_S4BEG),
    .SS4BEG(Tile_X3Y8_SS4BEG),
    .W1BEG(Tile_X3Y8_W1BEG),
    .W2BEG(Tile_X3Y8_W2BEG),
    .W2BEGb(Tile_X3Y8_W2BEGb),
    .WW4BEG(Tile_X3Y8_WW4BEG),
    .W6BEG(Tile_X3Y8_W6BEG),
    .Co(Tile_X3Y8_Co),
    .UserCLK(Tile_X3Y9_UserCLKo),
    .UserCLKo(Tile_X3Y8_UserCLKo),
    .FrameData(Tile_X2Y8_FrameData_O),
    .FrameData_O(Tile_X3Y8_FrameData_O),
    .FrameStrobe(Tile_X3Y9_FrameStrobe_O),
    .FrameStrobe_O(Tile_X3Y8_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
RegFile
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X4Y8_Emulate_Bitstream)
    )
`endif
    Tile_X4Y8_RegFile
    (
    .N1END(Tile_X4Y9_N1BEG),
    .N2MID(Tile_X4Y9_N2BEG),
    .N2END(Tile_X4Y9_N2BEGb),
    .N4END(Tile_X4Y9_N4BEG),
    .NN4END(Tile_X4Y9_NN4BEG),
    .E1END(Tile_X3Y8_E1BEG),
    .E2MID(Tile_X3Y8_E2BEG),
    .E2END(Tile_X3Y8_E2BEGb),
    .EE4END(Tile_X3Y8_EE4BEG),
    .E6END(Tile_X3Y8_E6BEG),
    .S1END(Tile_X4Y7_S1BEG),
    .S2MID(Tile_X4Y7_S2BEG),
    .S2END(Tile_X4Y7_S2BEGb),
    .S4END(Tile_X4Y7_S4BEG),
    .SS4END(Tile_X4Y7_SS4BEG),
    .W1END(Tile_X5Y8_W1BEG),
    .W2MID(Tile_X5Y8_W2BEG),
    .W2END(Tile_X5Y8_W2BEGb),
    .WW4END(Tile_X5Y8_WW4BEG),
    .W6END(Tile_X5Y8_W6BEG),
    .N1BEG(Tile_X4Y8_N1BEG),
    .N2BEG(Tile_X4Y8_N2BEG),
    .N2BEGb(Tile_X4Y8_N2BEGb),
    .N4BEG(Tile_X4Y8_N4BEG),
    .NN4BEG(Tile_X4Y8_NN4BEG),
    .E1BEG(Tile_X4Y8_E1BEG),
    .E2BEG(Tile_X4Y8_E2BEG),
    .E2BEGb(Tile_X4Y8_E2BEGb),
    .EE4BEG(Tile_X4Y8_EE4BEG),
    .E6BEG(Tile_X4Y8_E6BEG),
    .S1BEG(Tile_X4Y8_S1BEG),
    .S2BEG(Tile_X4Y8_S2BEG),
    .S2BEGb(Tile_X4Y8_S2BEGb),
    .S4BEG(Tile_X4Y8_S4BEG),
    .SS4BEG(Tile_X4Y8_SS4BEG),
    .W1BEG(Tile_X4Y8_W1BEG),
    .W2BEG(Tile_X4Y8_W2BEG),
    .W2BEGb(Tile_X4Y8_W2BEGb),
    .WW4BEG(Tile_X4Y8_WW4BEG),
    .W6BEG(Tile_X4Y8_W6BEG),
    .UserCLK(Tile_X4Y9_UserCLKo),
    .UserCLKo(Tile_X4Y8_UserCLKo),
    .FrameData(Tile_X3Y8_FrameData_O),
    .FrameData_O(Tile_X4Y8_FrameData_O),
    .FrameStrobe(Tile_X4Y9_FrameStrobe_O),
    .FrameStrobe_O(Tile_X4Y8_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X5Y8_Emulate_Bitstream)
    )
`endif
    Tile_X5Y8_LUT4AB
    (
    .N1END(Tile_X5Y9_N1BEG),
    .N2MID(Tile_X5Y9_N2BEG),
    .N2END(Tile_X5Y9_N2BEGb),
    .N4END(Tile_X5Y9_N4BEG),
    .NN4END(Tile_X5Y9_NN4BEG),
    .Ci(Tile_X5Y9_Co),
    .E1END(Tile_X4Y8_E1BEG),
    .E2MID(Tile_X4Y8_E2BEG),
    .E2END(Tile_X4Y8_E2BEGb),
    .EE4END(Tile_X4Y8_EE4BEG),
    .E6END(Tile_X4Y8_E6BEG),
    .S1END(Tile_X5Y7_S1BEG),
    .S2MID(Tile_X5Y7_S2BEG),
    .S2END(Tile_X5Y7_S2BEGb),
    .S4END(Tile_X5Y7_S4BEG),
    .SS4END(Tile_X5Y7_SS4BEG),
    .W1END(Tile_X6Y8_W1BEG),
    .W2MID(Tile_X6Y8_W2BEG),
    .W2END(Tile_X6Y8_W2BEGb),
    .WW4END(Tile_X6Y8_WW4BEG),
    .W6END(Tile_X6Y8_W6BEG),
    .N1BEG(Tile_X5Y8_N1BEG),
    .N2BEG(Tile_X5Y8_N2BEG),
    .N2BEGb(Tile_X5Y8_N2BEGb),
    .N4BEG(Tile_X5Y8_N4BEG),
    .NN4BEG(Tile_X5Y8_NN4BEG),
    .E1BEG(Tile_X5Y8_E1BEG),
    .E2BEG(Tile_X5Y8_E2BEG),
    .E2BEGb(Tile_X5Y8_E2BEGb),
    .EE4BEG(Tile_X5Y8_EE4BEG),
    .E6BEG(Tile_X5Y8_E6BEG),
    .S1BEG(Tile_X5Y8_S1BEG),
    .S2BEG(Tile_X5Y8_S2BEG),
    .S2BEGb(Tile_X5Y8_S2BEGb),
    .S4BEG(Tile_X5Y8_S4BEG),
    .SS4BEG(Tile_X5Y8_SS4BEG),
    .W1BEG(Tile_X5Y8_W1BEG),
    .W2BEG(Tile_X5Y8_W2BEG),
    .W2BEGb(Tile_X5Y8_W2BEGb),
    .WW4BEG(Tile_X5Y8_WW4BEG),
    .W6BEG(Tile_X5Y8_W6BEG),
    .Co(Tile_X5Y8_Co),
    .UserCLK(Tile_X5Y9_UserCLKo),
    .UserCLKo(Tile_X5Y8_UserCLKo),
    .FrameData(Tile_X4Y8_FrameData_O),
    .FrameData_O(Tile_X5Y8_FrameData_O),
    .FrameStrobe(Tile_X5Y9_FrameStrobe_O),
    .FrameStrobe_O(Tile_X5Y8_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X6Y8_Emulate_Bitstream)
    )
`endif
    Tile_X6Y8_LUT4AB
    (
    .N1END(Tile_X6Y9_N1BEG),
    .N2MID(Tile_X6Y9_N2BEG),
    .N2END(Tile_X6Y9_N2BEGb),
    .N4END(Tile_X6Y9_N4BEG),
    .NN4END(Tile_X6Y9_NN4BEG),
    .Ci(Tile_X6Y9_Co),
    .E1END(Tile_X5Y8_E1BEG),
    .E2MID(Tile_X5Y8_E2BEG),
    .E2END(Tile_X5Y8_E2BEGb),
    .EE4END(Tile_X5Y8_EE4BEG),
    .E6END(Tile_X5Y8_E6BEG),
    .S1END(Tile_X6Y7_S1BEG),
    .S2MID(Tile_X6Y7_S2BEG),
    .S2END(Tile_X6Y7_S2BEGb),
    .S4END(Tile_X6Y7_S4BEG),
    .SS4END(Tile_X6Y7_SS4BEG),
    .W1END(Tile_X7Y8_W1BEG),
    .W2MID(Tile_X7Y8_W2BEG),
    .W2END(Tile_X7Y8_W2BEGb),
    .WW4END(Tile_X7Y8_WW4BEG),
    .W6END(Tile_X7Y8_W6BEG),
    .N1BEG(Tile_X6Y8_N1BEG),
    .N2BEG(Tile_X6Y8_N2BEG),
    .N2BEGb(Tile_X6Y8_N2BEGb),
    .N4BEG(Tile_X6Y8_N4BEG),
    .NN4BEG(Tile_X6Y8_NN4BEG),
    .E1BEG(Tile_X6Y8_E1BEG),
    .E2BEG(Tile_X6Y8_E2BEG),
    .E2BEGb(Tile_X6Y8_E2BEGb),
    .EE4BEG(Tile_X6Y8_EE4BEG),
    .E6BEG(Tile_X6Y8_E6BEG),
    .S1BEG(Tile_X6Y8_S1BEG),
    .S2BEG(Tile_X6Y8_S2BEG),
    .S2BEGb(Tile_X6Y8_S2BEGb),
    .S4BEG(Tile_X6Y8_S4BEG),
    .SS4BEG(Tile_X6Y8_SS4BEG),
    .W1BEG(Tile_X6Y8_W1BEG),
    .W2BEG(Tile_X6Y8_W2BEG),
    .W2BEGb(Tile_X6Y8_W2BEGb),
    .WW4BEG(Tile_X6Y8_WW4BEG),
    .W6BEG(Tile_X6Y8_W6BEG),
    .Co(Tile_X6Y8_Co),
    .UserCLK(Tile_X6Y9_UserCLKo),
    .UserCLKo(Tile_X6Y8_UserCLKo),
    .FrameData(Tile_X5Y8_FrameData_O),
    .FrameData_O(Tile_X6Y8_FrameData_O),
    .FrameStrobe(Tile_X6Y9_FrameStrobe_O),
    .FrameStrobe_O(Tile_X6Y8_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X8Y8_Emulate_Bitstream)
    )
`endif
    Tile_X8Y8_LUT4AB
    (
    .N1END(Tile_X8Y9_N1BEG),
    .N2MID(Tile_X8Y9_N2BEG),
    .N2END(Tile_X8Y9_N2BEGb),
    .N4END(Tile_X8Y9_N4BEG),
    .NN4END(Tile_X8Y9_NN4BEG),
    .Ci(Tile_X8Y9_Co),
    .E1END(Tile_X7Y8_E1BEG),
    .E2MID(Tile_X7Y8_E2BEG),
    .E2END(Tile_X7Y8_E2BEGb),
    .EE4END(Tile_X7Y8_EE4BEG),
    .E6END(Tile_X7Y8_E6BEG),
    .S1END(Tile_X8Y7_S1BEG),
    .S2MID(Tile_X8Y7_S2BEG),
    .S2END(Tile_X8Y7_S2BEGb),
    .S4END(Tile_X8Y7_S4BEG),
    .SS4END(Tile_X8Y7_SS4BEG),
    .W1END(Tile_X9Y8_W1BEG),
    .W2MID(Tile_X9Y8_W2BEG),
    .W2END(Tile_X9Y8_W2BEGb),
    .WW4END(Tile_X9Y8_WW4BEG),
    .W6END(Tile_X9Y8_W6BEG),
    .N1BEG(Tile_X8Y8_N1BEG),
    .N2BEG(Tile_X8Y8_N2BEG),
    .N2BEGb(Tile_X8Y8_N2BEGb),
    .N4BEG(Tile_X8Y8_N4BEG),
    .NN4BEG(Tile_X8Y8_NN4BEG),
    .E1BEG(Tile_X8Y8_E1BEG),
    .E2BEG(Tile_X8Y8_E2BEG),
    .E2BEGb(Tile_X8Y8_E2BEGb),
    .EE4BEG(Tile_X8Y8_EE4BEG),
    .E6BEG(Tile_X8Y8_E6BEG),
    .S1BEG(Tile_X8Y8_S1BEG),
    .S2BEG(Tile_X8Y8_S2BEG),
    .S2BEGb(Tile_X8Y8_S2BEGb),
    .S4BEG(Tile_X8Y8_S4BEG),
    .SS4BEG(Tile_X8Y8_SS4BEG),
    .W1BEG(Tile_X8Y8_W1BEG),
    .W2BEG(Tile_X8Y8_W2BEG),
    .W2BEGb(Tile_X8Y8_W2BEGb),
    .WW4BEG(Tile_X8Y8_WW4BEG),
    .W6BEG(Tile_X8Y8_W6BEG),
    .Co(Tile_X8Y8_Co),
    .UserCLK(Tile_X8Y9_UserCLKo),
    .UserCLKo(Tile_X8Y8_UserCLKo),
    .FrameData(Tile_X7Y8_FrameData_O),
    .FrameData_O(Tile_X8Y8_FrameData_O),
    .FrameStrobe(Tile_X8Y9_FrameStrobe_O),
    .FrameStrobe_O(Tile_X8Y8_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X9Y8_Emulate_Bitstream)
    )
`endif
    Tile_X9Y8_LUT4AB
    (
    .N1END(Tile_X9Y9_N1BEG),
    .N2MID(Tile_X9Y9_N2BEG),
    .N2END(Tile_X9Y9_N2BEGb),
    .N4END(Tile_X9Y9_N4BEG),
    .NN4END(Tile_X9Y9_NN4BEG),
    .Ci(Tile_X9Y9_Co),
    .E1END(Tile_X8Y8_E1BEG),
    .E2MID(Tile_X8Y8_E2BEG),
    .E2END(Tile_X8Y8_E2BEGb),
    .EE4END(Tile_X8Y8_EE4BEG),
    .E6END(Tile_X8Y8_E6BEG),
    .S1END(Tile_X9Y7_S1BEG),
    .S2MID(Tile_X9Y7_S2BEG),
    .S2END(Tile_X9Y7_S2BEGb),
    .S4END(Tile_X9Y7_S4BEG),
    .SS4END(Tile_X9Y7_SS4BEG),
    .W1END(Tile_X10Y8_W1BEG),
    .W2MID(Tile_X10Y8_W2BEG),
    .W2END(Tile_X10Y8_W2BEGb),
    .WW4END(Tile_X10Y8_WW4BEG),
    .W6END(Tile_X10Y8_W6BEG),
    .N1BEG(Tile_X9Y8_N1BEG),
    .N2BEG(Tile_X9Y8_N2BEG),
    .N2BEGb(Tile_X9Y8_N2BEGb),
    .N4BEG(Tile_X9Y8_N4BEG),
    .NN4BEG(Tile_X9Y8_NN4BEG),
    .E1BEG(Tile_X9Y8_E1BEG),
    .E2BEG(Tile_X9Y8_E2BEG),
    .E2BEGb(Tile_X9Y8_E2BEGb),
    .EE4BEG(Tile_X9Y8_EE4BEG),
    .E6BEG(Tile_X9Y8_E6BEG),
    .S1BEG(Tile_X9Y8_S1BEG),
    .S2BEG(Tile_X9Y8_S2BEG),
    .S2BEGb(Tile_X9Y8_S2BEGb),
    .S4BEG(Tile_X9Y8_S4BEG),
    .SS4BEG(Tile_X9Y8_SS4BEG),
    .W1BEG(Tile_X9Y8_W1BEG),
    .W2BEG(Tile_X9Y8_W2BEG),
    .W2BEGb(Tile_X9Y8_W2BEGb),
    .WW4BEG(Tile_X9Y8_WW4BEG),
    .W6BEG(Tile_X9Y8_W6BEG),
    .Co(Tile_X9Y8_Co),
    .UserCLK(Tile_X9Y9_UserCLKo),
    .UserCLKo(Tile_X9Y8_UserCLKo),
    .FrameData(Tile_X8Y8_FrameData_O),
    .FrameData_O(Tile_X9Y8_FrameData_O),
    .FrameStrobe(Tile_X9Y9_FrameStrobe_O),
    .FrameStrobe_O(Tile_X9Y8_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
W_IO
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X0Y9_Emulate_Bitstream)
    )
`endif
    Tile_X0Y9_W_IO
    (
    .W1END(Tile_X1Y9_W1BEG),
    .W2MID(Tile_X1Y9_W2BEG),
    .W2END(Tile_X1Y9_W2BEGb),
    .WW4END(Tile_X1Y9_WW4BEG),
    .W6END(Tile_X1Y9_W6BEG),
    .E1BEG(Tile_X0Y9_E1BEG),
    .E2BEG(Tile_X0Y9_E2BEG),
    .E2BEGb(Tile_X0Y9_E2BEGb),
    .EE4BEG(Tile_X0Y9_EE4BEG),
    .E6BEG(Tile_X0Y9_E6BEG),
    .A_O_top(Tile_X0Y9_A_O_top),
    .A_I_top(Tile_X0Y9_A_I_top),
    .A_T_top(Tile_X0Y9_A_T_top),
    .B_O_top(Tile_X0Y9_B_O_top),
    .B_I_top(Tile_X0Y9_B_I_top),
    .B_T_top(Tile_X0Y9_B_T_top),
    .A_config_C_bit0(Tile_X0Y9_A_config_C_bit0),
    .A_config_C_bit1(Tile_X0Y9_A_config_C_bit1),
    .A_config_C_bit2(Tile_X0Y9_A_config_C_bit2),
    .A_config_C_bit3(Tile_X0Y9_A_config_C_bit3),
    .B_config_C_bit0(Tile_X0Y9_B_config_C_bit0),
    .B_config_C_bit1(Tile_X0Y9_B_config_C_bit1),
    .B_config_C_bit2(Tile_X0Y9_B_config_C_bit2),
    .B_config_C_bit3(Tile_X0Y9_B_config_C_bit3),
    .UserCLK(Tile_X0Y10_UserCLKo),
    .UserCLKo(Tile_X0Y9_UserCLKo),
    .FrameData(Row_Y9_FrameData),
    .FrameData_O(Tile_X0Y9_FrameData_O),
    .FrameStrobe(Tile_X0Y10_FrameStrobe_O),
    .FrameStrobe_O(Tile_X0Y9_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X1Y9_Emulate_Bitstream)
    )
`endif
    Tile_X1Y9_LUT4AB
    (
    .N1END(Tile_X1Y10_N1BEG),
    .N2MID(Tile_X1Y10_N2BEG),
    .N2END(Tile_X1Y10_N2BEGb),
    .N4END(Tile_X1Y10_N4BEG),
    .NN4END(Tile_X1Y10_NN4BEG),
    .Ci(Tile_X1Y10_Co),
    .E1END(Tile_X0Y9_E1BEG),
    .E2MID(Tile_X0Y9_E2BEG),
    .E2END(Tile_X0Y9_E2BEGb),
    .EE4END(Tile_X0Y9_EE4BEG),
    .E6END(Tile_X0Y9_E6BEG),
    .S1END(Tile_X1Y8_S1BEG),
    .S2MID(Tile_X1Y8_S2BEG),
    .S2END(Tile_X1Y8_S2BEGb),
    .S4END(Tile_X1Y8_S4BEG),
    .SS4END(Tile_X1Y8_SS4BEG),
    .W1END(Tile_X2Y9_W1BEG),
    .W2MID(Tile_X2Y9_W2BEG),
    .W2END(Tile_X2Y9_W2BEGb),
    .WW4END(Tile_X2Y9_WW4BEG),
    .W6END(Tile_X2Y9_W6BEG),
    .N1BEG(Tile_X1Y9_N1BEG),
    .N2BEG(Tile_X1Y9_N2BEG),
    .N2BEGb(Tile_X1Y9_N2BEGb),
    .N4BEG(Tile_X1Y9_N4BEG),
    .NN4BEG(Tile_X1Y9_NN4BEG),
    .E1BEG(Tile_X1Y9_E1BEG),
    .E2BEG(Tile_X1Y9_E2BEG),
    .E2BEGb(Tile_X1Y9_E2BEGb),
    .EE4BEG(Tile_X1Y9_EE4BEG),
    .E6BEG(Tile_X1Y9_E6BEG),
    .S1BEG(Tile_X1Y9_S1BEG),
    .S2BEG(Tile_X1Y9_S2BEG),
    .S2BEGb(Tile_X1Y9_S2BEGb),
    .S4BEG(Tile_X1Y9_S4BEG),
    .SS4BEG(Tile_X1Y9_SS4BEG),
    .W1BEG(Tile_X1Y9_W1BEG),
    .W2BEG(Tile_X1Y9_W2BEG),
    .W2BEGb(Tile_X1Y9_W2BEGb),
    .WW4BEG(Tile_X1Y9_WW4BEG),
    .W6BEG(Tile_X1Y9_W6BEG),
    .Co(Tile_X1Y9_Co),
    .UserCLK(Tile_X1Y10_UserCLKo),
    .UserCLKo(Tile_X1Y9_UserCLKo),
    .FrameData(Tile_X0Y9_FrameData_O),
    .FrameData_O(Tile_X1Y9_FrameData_O),
    .FrameStrobe(Tile_X1Y10_FrameStrobe_O),
    .FrameStrobe_O(Tile_X1Y9_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X2Y9_Emulate_Bitstream)
    )
`endif
    Tile_X2Y9_LUT4AB
    (
    .N1END(Tile_X2Y10_N1BEG),
    .N2MID(Tile_X2Y10_N2BEG),
    .N2END(Tile_X2Y10_N2BEGb),
    .N4END(Tile_X2Y10_N4BEG),
    .NN4END(Tile_X2Y10_NN4BEG),
    .Ci(Tile_X2Y10_Co),
    .E1END(Tile_X1Y9_E1BEG),
    .E2MID(Tile_X1Y9_E2BEG),
    .E2END(Tile_X1Y9_E2BEGb),
    .EE4END(Tile_X1Y9_EE4BEG),
    .E6END(Tile_X1Y9_E6BEG),
    .S1END(Tile_X2Y8_S1BEG),
    .S2MID(Tile_X2Y8_S2BEG),
    .S2END(Tile_X2Y8_S2BEGb),
    .S4END(Tile_X2Y8_S4BEG),
    .SS4END(Tile_X2Y8_SS4BEG),
    .W1END(Tile_X3Y9_W1BEG),
    .W2MID(Tile_X3Y9_W2BEG),
    .W2END(Tile_X3Y9_W2BEGb),
    .WW4END(Tile_X3Y9_WW4BEG),
    .W6END(Tile_X3Y9_W6BEG),
    .N1BEG(Tile_X2Y9_N1BEG),
    .N2BEG(Tile_X2Y9_N2BEG),
    .N2BEGb(Tile_X2Y9_N2BEGb),
    .N4BEG(Tile_X2Y9_N4BEG),
    .NN4BEG(Tile_X2Y9_NN4BEG),
    .E1BEG(Tile_X2Y9_E1BEG),
    .E2BEG(Tile_X2Y9_E2BEG),
    .E2BEGb(Tile_X2Y9_E2BEGb),
    .EE4BEG(Tile_X2Y9_EE4BEG),
    .E6BEG(Tile_X2Y9_E6BEG),
    .S1BEG(Tile_X2Y9_S1BEG),
    .S2BEG(Tile_X2Y9_S2BEG),
    .S2BEGb(Tile_X2Y9_S2BEGb),
    .S4BEG(Tile_X2Y9_S4BEG),
    .SS4BEG(Tile_X2Y9_SS4BEG),
    .W1BEG(Tile_X2Y9_W1BEG),
    .W2BEG(Tile_X2Y9_W2BEG),
    .W2BEGb(Tile_X2Y9_W2BEGb),
    .WW4BEG(Tile_X2Y9_WW4BEG),
    .W6BEG(Tile_X2Y9_W6BEG),
    .Co(Tile_X2Y9_Co),
    .UserCLK(Tile_X2Y10_UserCLKo),
    .UserCLKo(Tile_X2Y9_UserCLKo),
    .FrameData(Tile_X1Y9_FrameData_O),
    .FrameData_O(Tile_X2Y9_FrameData_O),
    .FrameStrobe(Tile_X2Y10_FrameStrobe_O),
    .FrameStrobe_O(Tile_X2Y9_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X3Y9_Emulate_Bitstream)
    )
`endif
    Tile_X3Y9_LUT4AB
    (
    .N1END(Tile_X3Y10_N1BEG),
    .N2MID(Tile_X3Y10_N2BEG),
    .N2END(Tile_X3Y10_N2BEGb),
    .N4END(Tile_X3Y10_N4BEG),
    .NN4END(Tile_X3Y10_NN4BEG),
    .Ci(Tile_X3Y10_Co),
    .E1END(Tile_X2Y9_E1BEG),
    .E2MID(Tile_X2Y9_E2BEG),
    .E2END(Tile_X2Y9_E2BEGb),
    .EE4END(Tile_X2Y9_EE4BEG),
    .E6END(Tile_X2Y9_E6BEG),
    .S1END(Tile_X3Y8_S1BEG),
    .S2MID(Tile_X3Y8_S2BEG),
    .S2END(Tile_X3Y8_S2BEGb),
    .S4END(Tile_X3Y8_S4BEG),
    .SS4END(Tile_X3Y8_SS4BEG),
    .W1END(Tile_X4Y9_W1BEG),
    .W2MID(Tile_X4Y9_W2BEG),
    .W2END(Tile_X4Y9_W2BEGb),
    .WW4END(Tile_X4Y9_WW4BEG),
    .W6END(Tile_X4Y9_W6BEG),
    .N1BEG(Tile_X3Y9_N1BEG),
    .N2BEG(Tile_X3Y9_N2BEG),
    .N2BEGb(Tile_X3Y9_N2BEGb),
    .N4BEG(Tile_X3Y9_N4BEG),
    .NN4BEG(Tile_X3Y9_NN4BEG),
    .E1BEG(Tile_X3Y9_E1BEG),
    .E2BEG(Tile_X3Y9_E2BEG),
    .E2BEGb(Tile_X3Y9_E2BEGb),
    .EE4BEG(Tile_X3Y9_EE4BEG),
    .E6BEG(Tile_X3Y9_E6BEG),
    .S1BEG(Tile_X3Y9_S1BEG),
    .S2BEG(Tile_X3Y9_S2BEG),
    .S2BEGb(Tile_X3Y9_S2BEGb),
    .S4BEG(Tile_X3Y9_S4BEG),
    .SS4BEG(Tile_X3Y9_SS4BEG),
    .W1BEG(Tile_X3Y9_W1BEG),
    .W2BEG(Tile_X3Y9_W2BEG),
    .W2BEGb(Tile_X3Y9_W2BEGb),
    .WW4BEG(Tile_X3Y9_WW4BEG),
    .W6BEG(Tile_X3Y9_W6BEG),
    .Co(Tile_X3Y9_Co),
    .UserCLK(Tile_X3Y10_UserCLKo),
    .UserCLKo(Tile_X3Y9_UserCLKo),
    .FrameData(Tile_X2Y9_FrameData_O),
    .FrameData_O(Tile_X3Y9_FrameData_O),
    .FrameStrobe(Tile_X3Y10_FrameStrobe_O),
    .FrameStrobe_O(Tile_X3Y9_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
RegFile
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X4Y9_Emulate_Bitstream)
    )
`endif
    Tile_X4Y9_RegFile
    (
    .N1END(Tile_X4Y10_N1BEG),
    .N2MID(Tile_X4Y10_N2BEG),
    .N2END(Tile_X4Y10_N2BEGb),
    .N4END(Tile_X4Y10_N4BEG),
    .NN4END(Tile_X4Y10_NN4BEG),
    .E1END(Tile_X3Y9_E1BEG),
    .E2MID(Tile_X3Y9_E2BEG),
    .E2END(Tile_X3Y9_E2BEGb),
    .EE4END(Tile_X3Y9_EE4BEG),
    .E6END(Tile_X3Y9_E6BEG),
    .S1END(Tile_X4Y8_S1BEG),
    .S2MID(Tile_X4Y8_S2BEG),
    .S2END(Tile_X4Y8_S2BEGb),
    .S4END(Tile_X4Y8_S4BEG),
    .SS4END(Tile_X4Y8_SS4BEG),
    .W1END(Tile_X5Y9_W1BEG),
    .W2MID(Tile_X5Y9_W2BEG),
    .W2END(Tile_X5Y9_W2BEGb),
    .WW4END(Tile_X5Y9_WW4BEG),
    .W6END(Tile_X5Y9_W6BEG),
    .N1BEG(Tile_X4Y9_N1BEG),
    .N2BEG(Tile_X4Y9_N2BEG),
    .N2BEGb(Tile_X4Y9_N2BEGb),
    .N4BEG(Tile_X4Y9_N4BEG),
    .NN4BEG(Tile_X4Y9_NN4BEG),
    .E1BEG(Tile_X4Y9_E1BEG),
    .E2BEG(Tile_X4Y9_E2BEG),
    .E2BEGb(Tile_X4Y9_E2BEGb),
    .EE4BEG(Tile_X4Y9_EE4BEG),
    .E6BEG(Tile_X4Y9_E6BEG),
    .S1BEG(Tile_X4Y9_S1BEG),
    .S2BEG(Tile_X4Y9_S2BEG),
    .S2BEGb(Tile_X4Y9_S2BEGb),
    .S4BEG(Tile_X4Y9_S4BEG),
    .SS4BEG(Tile_X4Y9_SS4BEG),
    .W1BEG(Tile_X4Y9_W1BEG),
    .W2BEG(Tile_X4Y9_W2BEG),
    .W2BEGb(Tile_X4Y9_W2BEGb),
    .WW4BEG(Tile_X4Y9_WW4BEG),
    .W6BEG(Tile_X4Y9_W6BEG),
    .UserCLK(Tile_X4Y10_UserCLKo),
    .UserCLKo(Tile_X4Y9_UserCLKo),
    .FrameData(Tile_X3Y9_FrameData_O),
    .FrameData_O(Tile_X4Y9_FrameData_O),
    .FrameStrobe(Tile_X4Y10_FrameStrobe_O),
    .FrameStrobe_O(Tile_X4Y9_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X5Y9_Emulate_Bitstream)
    )
`endif
    Tile_X5Y9_LUT4AB
    (
    .N1END(Tile_X5Y10_N1BEG),
    .N2MID(Tile_X5Y10_N2BEG),
    .N2END(Tile_X5Y10_N2BEGb),
    .N4END(Tile_X5Y10_N4BEG),
    .NN4END(Tile_X5Y10_NN4BEG),
    .Ci(Tile_X5Y10_Co),
    .E1END(Tile_X4Y9_E1BEG),
    .E2MID(Tile_X4Y9_E2BEG),
    .E2END(Tile_X4Y9_E2BEGb),
    .EE4END(Tile_X4Y9_EE4BEG),
    .E6END(Tile_X4Y9_E6BEG),
    .S1END(Tile_X5Y8_S1BEG),
    .S2MID(Tile_X5Y8_S2BEG),
    .S2END(Tile_X5Y8_S2BEGb),
    .S4END(Tile_X5Y8_S4BEG),
    .SS4END(Tile_X5Y8_SS4BEG),
    .W1END(Tile_X6Y9_W1BEG),
    .W2MID(Tile_X6Y9_W2BEG),
    .W2END(Tile_X6Y9_W2BEGb),
    .WW4END(Tile_X6Y9_WW4BEG),
    .W6END(Tile_X6Y9_W6BEG),
    .N1BEG(Tile_X5Y9_N1BEG),
    .N2BEG(Tile_X5Y9_N2BEG),
    .N2BEGb(Tile_X5Y9_N2BEGb),
    .N4BEG(Tile_X5Y9_N4BEG),
    .NN4BEG(Tile_X5Y9_NN4BEG),
    .E1BEG(Tile_X5Y9_E1BEG),
    .E2BEG(Tile_X5Y9_E2BEG),
    .E2BEGb(Tile_X5Y9_E2BEGb),
    .EE4BEG(Tile_X5Y9_EE4BEG),
    .E6BEG(Tile_X5Y9_E6BEG),
    .S1BEG(Tile_X5Y9_S1BEG),
    .S2BEG(Tile_X5Y9_S2BEG),
    .S2BEGb(Tile_X5Y9_S2BEGb),
    .S4BEG(Tile_X5Y9_S4BEG),
    .SS4BEG(Tile_X5Y9_SS4BEG),
    .W1BEG(Tile_X5Y9_W1BEG),
    .W2BEG(Tile_X5Y9_W2BEG),
    .W2BEGb(Tile_X5Y9_W2BEGb),
    .WW4BEG(Tile_X5Y9_WW4BEG),
    .W6BEG(Tile_X5Y9_W6BEG),
    .Co(Tile_X5Y9_Co),
    .UserCLK(Tile_X5Y10_UserCLKo),
    .UserCLKo(Tile_X5Y9_UserCLKo),
    .FrameData(Tile_X4Y9_FrameData_O),
    .FrameData_O(Tile_X5Y9_FrameData_O),
    .FrameStrobe(Tile_X5Y10_FrameStrobe_O),
    .FrameStrobe_O(Tile_X5Y9_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X6Y9_Emulate_Bitstream)
    )
`endif
    Tile_X6Y9_LUT4AB
    (
    .N1END(Tile_X6Y10_N1BEG),
    .N2MID(Tile_X6Y10_N2BEG),
    .N2END(Tile_X6Y10_N2BEGb),
    .N4END(Tile_X6Y10_N4BEG),
    .NN4END(Tile_X6Y10_NN4BEG),
    .Ci(Tile_X6Y10_Co),
    .E1END(Tile_X5Y9_E1BEG),
    .E2MID(Tile_X5Y9_E2BEG),
    .E2END(Tile_X5Y9_E2BEGb),
    .EE4END(Tile_X5Y9_EE4BEG),
    .E6END(Tile_X5Y9_E6BEG),
    .S1END(Tile_X6Y8_S1BEG),
    .S2MID(Tile_X6Y8_S2BEG),
    .S2END(Tile_X6Y8_S2BEGb),
    .S4END(Tile_X6Y8_S4BEG),
    .SS4END(Tile_X6Y8_SS4BEG),
    .W1END(Tile_X7Y9_W1BEG),
    .W2MID(Tile_X7Y9_W2BEG),
    .W2END(Tile_X7Y9_W2BEGb),
    .WW4END(Tile_X7Y9_WW4BEG),
    .W6END(Tile_X7Y9_W6BEG),
    .N1BEG(Tile_X6Y9_N1BEG),
    .N2BEG(Tile_X6Y9_N2BEG),
    .N2BEGb(Tile_X6Y9_N2BEGb),
    .N4BEG(Tile_X6Y9_N4BEG),
    .NN4BEG(Tile_X6Y9_NN4BEG),
    .E1BEG(Tile_X6Y9_E1BEG),
    .E2BEG(Tile_X6Y9_E2BEG),
    .E2BEGb(Tile_X6Y9_E2BEGb),
    .EE4BEG(Tile_X6Y9_EE4BEG),
    .E6BEG(Tile_X6Y9_E6BEG),
    .S1BEG(Tile_X6Y9_S1BEG),
    .S2BEG(Tile_X6Y9_S2BEG),
    .S2BEGb(Tile_X6Y9_S2BEGb),
    .S4BEG(Tile_X6Y9_S4BEG),
    .SS4BEG(Tile_X6Y9_SS4BEG),
    .W1BEG(Tile_X6Y9_W1BEG),
    .W2BEG(Tile_X6Y9_W2BEG),
    .W2BEGb(Tile_X6Y9_W2BEGb),
    .WW4BEG(Tile_X6Y9_WW4BEG),
    .W6BEG(Tile_X6Y9_W6BEG),
    .Co(Tile_X6Y9_Co),
    .UserCLK(Tile_X6Y10_UserCLKo),
    .UserCLKo(Tile_X6Y9_UserCLKo),
    .FrameData(Tile_X5Y9_FrameData_O),
    .FrameData_O(Tile_X6Y9_FrameData_O),
    .FrameStrobe(Tile_X6Y10_FrameStrobe_O),
    .FrameStrobe_O(Tile_X6Y9_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
DSP
`ifdef EMULATION
    #(
    .Tile_X0Y0_Emulate_Bitstream(`Tile_X7Y9_Emulate_Bitstream),
    .Tile_X0Y1_Emulate_Bitstream(`Tile_X7Y10_Emulate_Bitstream)
    )
`endif
    Tile_X7Y9_DSP
    (
    .Tile_X0Y0_E1END(Tile_X6Y9_E1BEG),
    .Tile_X0Y0_E2MID(Tile_X6Y9_E2BEG),
    .Tile_X0Y0_E2END(Tile_X6Y9_E2BEGb),
    .Tile_X0Y0_EE4END(Tile_X6Y9_EE4BEG),
    .Tile_X0Y0_E6END(Tile_X6Y9_E6BEG),
    .Tile_X0Y0_S1END(Tile_X7Y8_S1BEG),
    .Tile_X0Y0_S2MID(Tile_X7Y8_S2BEG),
    .Tile_X0Y0_S2END(Tile_X7Y8_S2BEGb),
    .Tile_X0Y0_S4END(Tile_X7Y8_S4BEG),
    .Tile_X0Y0_SS4END(Tile_X7Y8_SS4BEG),
    .Tile_X0Y0_W1END(Tile_X8Y9_W1BEG),
    .Tile_X0Y0_W2MID(Tile_X8Y9_W2BEG),
    .Tile_X0Y0_W2END(Tile_X8Y9_W2BEGb),
    .Tile_X0Y0_WW4END(Tile_X8Y9_WW4BEG),
    .Tile_X0Y0_W6END(Tile_X8Y9_W6BEG),
    .Tile_X0Y1_N1END(Tile_X7Y11_N1BEG),
    .Tile_X0Y1_N2MID(Tile_X7Y11_N2BEG),
    .Tile_X0Y1_N2END(Tile_X7Y11_N2BEGb),
    .Tile_X0Y1_N4END(Tile_X7Y11_N4BEG),
    .Tile_X0Y1_NN4END(Tile_X7Y11_NN4BEG),
    .Tile_X0Y1_E1END(Tile_X6Y10_E1BEG),
    .Tile_X0Y1_E2MID(Tile_X6Y10_E2BEG),
    .Tile_X0Y1_E2END(Tile_X6Y10_E2BEGb),
    .Tile_X0Y1_EE4END(Tile_X6Y10_EE4BEG),
    .Tile_X0Y1_E6END(Tile_X6Y10_E6BEG),
    .Tile_X0Y1_W1END(Tile_X8Y10_W1BEG),
    .Tile_X0Y1_W2MID(Tile_X8Y10_W2BEG),
    .Tile_X0Y1_W2END(Tile_X8Y10_W2BEGb),
    .Tile_X0Y1_WW4END(Tile_X8Y10_WW4BEG),
    .Tile_X0Y1_W6END(Tile_X8Y10_W6BEG),
    .Tile_X0Y0_N1BEG(Tile_X7Y9_N1BEG),
    .Tile_X0Y0_N2BEG(Tile_X7Y9_N2BEG),
    .Tile_X0Y0_N2BEGb(Tile_X7Y9_N2BEGb),
    .Tile_X0Y0_N4BEG(Tile_X7Y9_N4BEG),
    .Tile_X0Y0_NN4BEG(Tile_X7Y9_NN4BEG),
    .Tile_X0Y0_E1BEG(Tile_X7Y9_E1BEG),
    .Tile_X0Y0_E2BEG(Tile_X7Y9_E2BEG),
    .Tile_X0Y0_E2BEGb(Tile_X7Y9_E2BEGb),
    .Tile_X0Y0_EE4BEG(Tile_X7Y9_EE4BEG),
    .Tile_X0Y0_E6BEG(Tile_X7Y9_E6BEG),
    .Tile_X0Y0_W1BEG(Tile_X7Y9_W1BEG),
    .Tile_X0Y0_W2BEG(Tile_X7Y9_W2BEG),
    .Tile_X0Y0_W2BEGb(Tile_X7Y9_W2BEGb),
    .Tile_X0Y0_WW4BEG(Tile_X7Y9_WW4BEG),
    .Tile_X0Y0_W6BEG(Tile_X7Y9_W6BEG),
    .Tile_X0Y1_E1BEG(Tile_X7Y10_E1BEG),
    .Tile_X0Y1_E2BEG(Tile_X7Y10_E2BEG),
    .Tile_X0Y1_E2BEGb(Tile_X7Y10_E2BEGb),
    .Tile_X0Y1_EE4BEG(Tile_X7Y10_EE4BEG),
    .Tile_X0Y1_E6BEG(Tile_X7Y10_E6BEG),
    .Tile_X0Y1_S1BEG(Tile_X7Y10_S1BEG),
    .Tile_X0Y1_S2BEG(Tile_X7Y10_S2BEG),
    .Tile_X0Y1_S2BEGb(Tile_X7Y10_S2BEGb),
    .Tile_X0Y1_S4BEG(Tile_X7Y10_S4BEG),
    .Tile_X0Y1_SS4BEG(Tile_X7Y10_SS4BEG),
    .Tile_X0Y1_W1BEG(Tile_X7Y10_W1BEG),
    .Tile_X0Y1_W2BEG(Tile_X7Y10_W2BEG),
    .Tile_X0Y1_W2BEGb(Tile_X7Y10_W2BEGb),
    .Tile_X0Y1_WW4BEG(Tile_X7Y10_WW4BEG),
    .Tile_X0Y1_W6BEG(Tile_X7Y10_W6BEG),
    .Tile_X0Y0_UserCLKo(Tile_X7Y9_UserCLKo),
    .Tile_X0Y1_UserCLK(Tile_X7Y11_UserCLKo),
    .Tile_X0Y0_FrameData(Tile_X6Y9_FrameData_O),
    .Tile_X0Y0_FrameData_O(Tile_X7Y9_FrameData_O),
    .Tile_X0Y0_FrameStrobe_O(Tile_X7Y9_FrameStrobe_O),
    .Tile_X0Y1_FrameData(Tile_X6Y10_FrameData_O),
    .Tile_X0Y1_FrameData_O(Tile_X7Y10_FrameData_O),
    .Tile_X0Y1_FrameStrobe(Tile_X7Y11_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X8Y9_Emulate_Bitstream)
    )
`endif
    Tile_X8Y9_LUT4AB
    (
    .N1END(Tile_X8Y10_N1BEG),
    .N2MID(Tile_X8Y10_N2BEG),
    .N2END(Tile_X8Y10_N2BEGb),
    .N4END(Tile_X8Y10_N4BEG),
    .NN4END(Tile_X8Y10_NN4BEG),
    .Ci(Tile_X8Y10_Co),
    .E1END(Tile_X7Y9_E1BEG),
    .E2MID(Tile_X7Y9_E2BEG),
    .E2END(Tile_X7Y9_E2BEGb),
    .EE4END(Tile_X7Y9_EE4BEG),
    .E6END(Tile_X7Y9_E6BEG),
    .S1END(Tile_X8Y8_S1BEG),
    .S2MID(Tile_X8Y8_S2BEG),
    .S2END(Tile_X8Y8_S2BEGb),
    .S4END(Tile_X8Y8_S4BEG),
    .SS4END(Tile_X8Y8_SS4BEG),
    .W1END(Tile_X9Y9_W1BEG),
    .W2MID(Tile_X9Y9_W2BEG),
    .W2END(Tile_X9Y9_W2BEGb),
    .WW4END(Tile_X9Y9_WW4BEG),
    .W6END(Tile_X9Y9_W6BEG),
    .N1BEG(Tile_X8Y9_N1BEG),
    .N2BEG(Tile_X8Y9_N2BEG),
    .N2BEGb(Tile_X8Y9_N2BEGb),
    .N4BEG(Tile_X8Y9_N4BEG),
    .NN4BEG(Tile_X8Y9_NN4BEG),
    .E1BEG(Tile_X8Y9_E1BEG),
    .E2BEG(Tile_X8Y9_E2BEG),
    .E2BEGb(Tile_X8Y9_E2BEGb),
    .EE4BEG(Tile_X8Y9_EE4BEG),
    .E6BEG(Tile_X8Y9_E6BEG),
    .S1BEG(Tile_X8Y9_S1BEG),
    .S2BEG(Tile_X8Y9_S2BEG),
    .S2BEGb(Tile_X8Y9_S2BEGb),
    .S4BEG(Tile_X8Y9_S4BEG),
    .SS4BEG(Tile_X8Y9_SS4BEG),
    .W1BEG(Tile_X8Y9_W1BEG),
    .W2BEG(Tile_X8Y9_W2BEG),
    .W2BEGb(Tile_X8Y9_W2BEGb),
    .WW4BEG(Tile_X8Y9_WW4BEG),
    .W6BEG(Tile_X8Y9_W6BEG),
    .Co(Tile_X8Y9_Co),
    .UserCLK(Tile_X8Y10_UserCLKo),
    .UserCLKo(Tile_X8Y9_UserCLKo),
    .FrameData(Tile_X7Y9_FrameData_O),
    .FrameData_O(Tile_X8Y9_FrameData_O),
    .FrameStrobe(Tile_X8Y10_FrameStrobe_O),
    .FrameStrobe_O(Tile_X8Y9_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X9Y9_Emulate_Bitstream)
    )
`endif
    Tile_X9Y9_LUT4AB
    (
    .N1END(Tile_X9Y10_N1BEG),
    .N2MID(Tile_X9Y10_N2BEG),
    .N2END(Tile_X9Y10_N2BEGb),
    .N4END(Tile_X9Y10_N4BEG),
    .NN4END(Tile_X9Y10_NN4BEG),
    .Ci(Tile_X9Y10_Co),
    .E1END(Tile_X8Y9_E1BEG),
    .E2MID(Tile_X8Y9_E2BEG),
    .E2END(Tile_X8Y9_E2BEGb),
    .EE4END(Tile_X8Y9_EE4BEG),
    .E6END(Tile_X8Y9_E6BEG),
    .S1END(Tile_X9Y8_S1BEG),
    .S2MID(Tile_X9Y8_S2BEG),
    .S2END(Tile_X9Y8_S2BEGb),
    .S4END(Tile_X9Y8_S4BEG),
    .SS4END(Tile_X9Y8_SS4BEG),
    .W1END(Tile_X10Y9_W1BEG),
    .W2MID(Tile_X10Y9_W2BEG),
    .W2END(Tile_X10Y9_W2BEGb),
    .WW4END(Tile_X10Y9_WW4BEG),
    .W6END(Tile_X10Y9_W6BEG),
    .N1BEG(Tile_X9Y9_N1BEG),
    .N2BEG(Tile_X9Y9_N2BEG),
    .N2BEGb(Tile_X9Y9_N2BEGb),
    .N4BEG(Tile_X9Y9_N4BEG),
    .NN4BEG(Tile_X9Y9_NN4BEG),
    .E1BEG(Tile_X9Y9_E1BEG),
    .E2BEG(Tile_X9Y9_E2BEG),
    .E2BEGb(Tile_X9Y9_E2BEGb),
    .EE4BEG(Tile_X9Y9_EE4BEG),
    .E6BEG(Tile_X9Y9_E6BEG),
    .S1BEG(Tile_X9Y9_S1BEG),
    .S2BEG(Tile_X9Y9_S2BEG),
    .S2BEGb(Tile_X9Y9_S2BEGb),
    .S4BEG(Tile_X9Y9_S4BEG),
    .SS4BEG(Tile_X9Y9_SS4BEG),
    .W1BEG(Tile_X9Y9_W1BEG),
    .W2BEG(Tile_X9Y9_W2BEG),
    .W2BEGb(Tile_X9Y9_W2BEGb),
    .WW4BEG(Tile_X9Y9_WW4BEG),
    .W6BEG(Tile_X9Y9_W6BEG),
    .Co(Tile_X9Y9_Co),
    .UserCLK(Tile_X9Y10_UserCLKo),
    .UserCLKo(Tile_X9Y9_UserCLKo),
    .FrameData(Tile_X8Y9_FrameData_O),
    .FrameData_O(Tile_X9Y9_FrameData_O),
    .FrameStrobe(Tile_X9Y10_FrameStrobe_O),
    .FrameStrobe_O(Tile_X9Y9_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
IHP_SRAM
`ifdef EMULATION
    #(
    .Tile_X0Y0_Emulate_Bitstream(`Tile_X10Y9_Emulate_Bitstream),
    .Tile_X0Y1_Emulate_Bitstream(`Tile_X10Y10_Emulate_Bitstream)
    )
`endif
    Tile_X10Y9_IHP_SRAM
    (
    .Tile_X0Y0_E1END(Tile_X9Y9_E1BEG),
    .Tile_X0Y0_E2MID(Tile_X9Y9_E2BEG),
    .Tile_X0Y0_E2END(Tile_X9Y9_E2BEGb),
    .Tile_X0Y0_EE4END(Tile_X9Y9_EE4BEG),
    .Tile_X0Y0_E6END(Tile_X9Y9_E6BEG),
    .Tile_X0Y0_S1END(Tile_X10Y8_S1BEG),
    .Tile_X0Y0_S2MID(Tile_X10Y8_S2BEG),
    .Tile_X0Y0_S2END(Tile_X10Y8_S2BEGb),
    .Tile_X0Y0_S4END(Tile_X10Y8_S4BEG),
    .Tile_X0Y1_N1END(Tile_X10Y11_N1BEG),
    .Tile_X0Y1_N2MID(Tile_X10Y11_N2BEG),
    .Tile_X0Y1_N2END(Tile_X10Y11_N2BEGb),
    .Tile_X0Y1_N4END(Tile_X10Y11_N4BEG),
    .Tile_X0Y1_E1END(Tile_X9Y10_E1BEG),
    .Tile_X0Y1_E2MID(Tile_X9Y10_E2BEG),
    .Tile_X0Y1_E2END(Tile_X9Y10_E2BEGb),
    .Tile_X0Y1_EE4END(Tile_X9Y10_EE4BEG),
    .Tile_X0Y1_E6END(Tile_X9Y10_E6BEG),
    .Tile_X0Y0_N1BEG(Tile_X10Y9_N1BEG),
    .Tile_X0Y0_N2BEG(Tile_X10Y9_N2BEG),
    .Tile_X0Y0_N2BEGb(Tile_X10Y9_N2BEGb),
    .Tile_X0Y0_N4BEG(Tile_X10Y9_N4BEG),
    .Tile_X0Y0_W1BEG(Tile_X10Y9_W1BEG),
    .Tile_X0Y0_W2BEG(Tile_X10Y9_W2BEG),
    .Tile_X0Y0_W2BEGb(Tile_X10Y9_W2BEGb),
    .Tile_X0Y0_WW4BEG(Tile_X10Y9_WW4BEG),
    .Tile_X0Y0_W6BEG(Tile_X10Y9_W6BEG),
    .Tile_X0Y1_S1BEG(Tile_X10Y10_S1BEG),
    .Tile_X0Y1_S2BEG(Tile_X10Y10_S2BEG),
    .Tile_X0Y1_S2BEGb(Tile_X10Y10_S2BEGb),
    .Tile_X0Y1_S4BEG(Tile_X10Y10_S4BEG),
    .Tile_X0Y1_W1BEG(Tile_X10Y10_W1BEG),
    .Tile_X0Y1_W2BEG(Tile_X10Y10_W2BEG),
    .Tile_X0Y1_W2BEGb(Tile_X10Y10_W2BEGb),
    .Tile_X0Y1_WW4BEG(Tile_X10Y10_WW4BEG),
    .Tile_X0Y1_W6BEG(Tile_X10Y10_W6BEG),
    .CONFIGURED_top(Tile_X10Y10_CONFIGURED_top),
    .DOUT_SRAM0(Tile_X10Y10_DOUT_SRAM0),
    .DOUT_SRAM1(Tile_X10Y10_DOUT_SRAM1),
    .DOUT_SRAM2(Tile_X10Y10_DOUT_SRAM2),
    .DOUT_SRAM3(Tile_X10Y10_DOUT_SRAM3),
    .DOUT_SRAM4(Tile_X10Y10_DOUT_SRAM4),
    .DOUT_SRAM5(Tile_X10Y10_DOUT_SRAM5),
    .DOUT_SRAM6(Tile_X10Y10_DOUT_SRAM6),
    .DOUT_SRAM7(Tile_X10Y10_DOUT_SRAM7),
    .DOUT_SRAM8(Tile_X10Y10_DOUT_SRAM8),
    .DOUT_SRAM9(Tile_X10Y10_DOUT_SRAM9),
    .DOUT_SRAM10(Tile_X10Y10_DOUT_SRAM10),
    .DOUT_SRAM11(Tile_X10Y10_DOUT_SRAM11),
    .DOUT_SRAM12(Tile_X10Y10_DOUT_SRAM12),
    .DOUT_SRAM13(Tile_X10Y10_DOUT_SRAM13),
    .DOUT_SRAM14(Tile_X10Y10_DOUT_SRAM14),
    .DOUT_SRAM15(Tile_X10Y10_DOUT_SRAM15),
    .DOUT_SRAM16(Tile_X10Y10_DOUT_SRAM16),
    .DOUT_SRAM17(Tile_X10Y10_DOUT_SRAM17),
    .DOUT_SRAM18(Tile_X10Y10_DOUT_SRAM18),
    .DOUT_SRAM19(Tile_X10Y10_DOUT_SRAM19),
    .DOUT_SRAM20(Tile_X10Y10_DOUT_SRAM20),
    .DOUT_SRAM21(Tile_X10Y10_DOUT_SRAM21),
    .DOUT_SRAM22(Tile_X10Y10_DOUT_SRAM22),
    .DOUT_SRAM23(Tile_X10Y10_DOUT_SRAM23),
    .DOUT_SRAM24(Tile_X10Y10_DOUT_SRAM24),
    .DOUT_SRAM25(Tile_X10Y10_DOUT_SRAM25),
    .DOUT_SRAM26(Tile_X10Y10_DOUT_SRAM26),
    .DOUT_SRAM27(Tile_X10Y10_DOUT_SRAM27),
    .DOUT_SRAM28(Tile_X10Y10_DOUT_SRAM28),
    .DOUT_SRAM29(Tile_X10Y10_DOUT_SRAM29),
    .DOUT_SRAM30(Tile_X10Y10_DOUT_SRAM30),
    .DOUT_SRAM31(Tile_X10Y10_DOUT_SRAM31),
    .ADDR_SRAM0(Tile_X10Y10_ADDR_SRAM0),
    .ADDR_SRAM1(Tile_X10Y10_ADDR_SRAM1),
    .ADDR_SRAM2(Tile_X10Y10_ADDR_SRAM2),
    .ADDR_SRAM3(Tile_X10Y10_ADDR_SRAM3),
    .ADDR_SRAM4(Tile_X10Y10_ADDR_SRAM4),
    .ADDR_SRAM5(Tile_X10Y10_ADDR_SRAM5),
    .ADDR_SRAM6(Tile_X10Y10_ADDR_SRAM6),
    .ADDR_SRAM7(Tile_X10Y10_ADDR_SRAM7),
    .ADDR_SRAM8(Tile_X10Y10_ADDR_SRAM8),
    .ADDR_SRAM9(Tile_X10Y10_ADDR_SRAM9),
    .BM_SRAM0(Tile_X10Y10_BM_SRAM0),
    .BM_SRAM1(Tile_X10Y10_BM_SRAM1),
    .BM_SRAM2(Tile_X10Y10_BM_SRAM2),
    .BM_SRAM3(Tile_X10Y10_BM_SRAM3),
    .BM_SRAM4(Tile_X10Y10_BM_SRAM4),
    .BM_SRAM5(Tile_X10Y10_BM_SRAM5),
    .BM_SRAM6(Tile_X10Y10_BM_SRAM6),
    .BM_SRAM7(Tile_X10Y10_BM_SRAM7),
    .BM_SRAM8(Tile_X10Y10_BM_SRAM8),
    .BM_SRAM9(Tile_X10Y10_BM_SRAM9),
    .BM_SRAM10(Tile_X10Y10_BM_SRAM10),
    .BM_SRAM11(Tile_X10Y10_BM_SRAM11),
    .BM_SRAM12(Tile_X10Y10_BM_SRAM12),
    .BM_SRAM13(Tile_X10Y10_BM_SRAM13),
    .BM_SRAM14(Tile_X10Y10_BM_SRAM14),
    .BM_SRAM15(Tile_X10Y10_BM_SRAM15),
    .BM_SRAM16(Tile_X10Y10_BM_SRAM16),
    .BM_SRAM17(Tile_X10Y10_BM_SRAM17),
    .BM_SRAM18(Tile_X10Y10_BM_SRAM18),
    .BM_SRAM19(Tile_X10Y10_BM_SRAM19),
    .BM_SRAM20(Tile_X10Y10_BM_SRAM20),
    .BM_SRAM21(Tile_X10Y10_BM_SRAM21),
    .BM_SRAM22(Tile_X10Y10_BM_SRAM22),
    .BM_SRAM23(Tile_X10Y10_BM_SRAM23),
    .BM_SRAM24(Tile_X10Y10_BM_SRAM24),
    .BM_SRAM25(Tile_X10Y10_BM_SRAM25),
    .BM_SRAM26(Tile_X10Y10_BM_SRAM26),
    .BM_SRAM27(Tile_X10Y10_BM_SRAM27),
    .BM_SRAM28(Tile_X10Y10_BM_SRAM28),
    .BM_SRAM29(Tile_X10Y10_BM_SRAM29),
    .BM_SRAM30(Tile_X10Y10_BM_SRAM30),
    .BM_SRAM31(Tile_X10Y10_BM_SRAM31),
    .CLK_SRAM(Tile_X10Y10_CLK_SRAM),
    .DIN_SRAM0(Tile_X10Y10_DIN_SRAM0),
    .DIN_SRAM1(Tile_X10Y10_DIN_SRAM1),
    .DIN_SRAM2(Tile_X10Y10_DIN_SRAM2),
    .DIN_SRAM3(Tile_X10Y10_DIN_SRAM3),
    .DIN_SRAM4(Tile_X10Y10_DIN_SRAM4),
    .DIN_SRAM5(Tile_X10Y10_DIN_SRAM5),
    .DIN_SRAM6(Tile_X10Y10_DIN_SRAM6),
    .DIN_SRAM7(Tile_X10Y10_DIN_SRAM7),
    .DIN_SRAM8(Tile_X10Y10_DIN_SRAM8),
    .DIN_SRAM9(Tile_X10Y10_DIN_SRAM9),
    .DIN_SRAM10(Tile_X10Y10_DIN_SRAM10),
    .DIN_SRAM11(Tile_X10Y10_DIN_SRAM11),
    .DIN_SRAM12(Tile_X10Y10_DIN_SRAM12),
    .DIN_SRAM13(Tile_X10Y10_DIN_SRAM13),
    .DIN_SRAM14(Tile_X10Y10_DIN_SRAM14),
    .DIN_SRAM15(Tile_X10Y10_DIN_SRAM15),
    .DIN_SRAM16(Tile_X10Y10_DIN_SRAM16),
    .DIN_SRAM17(Tile_X10Y10_DIN_SRAM17),
    .DIN_SRAM18(Tile_X10Y10_DIN_SRAM18),
    .DIN_SRAM19(Tile_X10Y10_DIN_SRAM19),
    .DIN_SRAM20(Tile_X10Y10_DIN_SRAM20),
    .DIN_SRAM21(Tile_X10Y10_DIN_SRAM21),
    .DIN_SRAM22(Tile_X10Y10_DIN_SRAM22),
    .DIN_SRAM23(Tile_X10Y10_DIN_SRAM23),
    .DIN_SRAM24(Tile_X10Y10_DIN_SRAM24),
    .DIN_SRAM25(Tile_X10Y10_DIN_SRAM25),
    .DIN_SRAM26(Tile_X10Y10_DIN_SRAM26),
    .DIN_SRAM27(Tile_X10Y10_DIN_SRAM27),
    .DIN_SRAM28(Tile_X10Y10_DIN_SRAM28),
    .DIN_SRAM29(Tile_X10Y10_DIN_SRAM29),
    .DIN_SRAM30(Tile_X10Y10_DIN_SRAM30),
    .DIN_SRAM31(Tile_X10Y10_DIN_SRAM31),
    .MEN_SRAM(Tile_X10Y10_MEN_SRAM),
    .REN_SRAM(Tile_X10Y10_REN_SRAM),
    .TIE_HIGH_SRAM(Tile_X10Y10_TIE_HIGH_SRAM),
    .TIE_LOW_SRAM(Tile_X10Y10_TIE_LOW_SRAM),
    .WEN_SRAM(Tile_X10Y10_WEN_SRAM),
    .Tile_X0Y0_UserCLKo(Tile_X10Y9_UserCLKo),
    .Tile_X0Y1_UserCLK(Tile_X10Y11_UserCLKo),
    .Tile_X0Y0_FrameData(Tile_X9Y9_FrameData_O),
    .Tile_X0Y0_FrameData_O(Tile_X10Y9_FrameData_O),
    .Tile_X0Y0_FrameStrobe_O(Tile_X10Y9_FrameStrobe_O),
    .Tile_X0Y1_FrameData(Tile_X9Y10_FrameData_O),
    .Tile_X0Y1_FrameData_O(Tile_X10Y10_FrameData_O),
    .Tile_X0Y1_FrameStrobe(Tile_X10Y11_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
W_IO
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X0Y10_Emulate_Bitstream)
    )
`endif
    Tile_X0Y10_W_IO
    (
    .W1END(Tile_X1Y10_W1BEG),
    .W2MID(Tile_X1Y10_W2BEG),
    .W2END(Tile_X1Y10_W2BEGb),
    .WW4END(Tile_X1Y10_WW4BEG),
    .W6END(Tile_X1Y10_W6BEG),
    .E1BEG(Tile_X0Y10_E1BEG),
    .E2BEG(Tile_X0Y10_E2BEG),
    .E2BEGb(Tile_X0Y10_E2BEGb),
    .EE4BEG(Tile_X0Y10_EE4BEG),
    .E6BEG(Tile_X0Y10_E6BEG),
    .A_O_top(Tile_X0Y10_A_O_top),
    .A_I_top(Tile_X0Y10_A_I_top),
    .A_T_top(Tile_X0Y10_A_T_top),
    .B_O_top(Tile_X0Y10_B_O_top),
    .B_I_top(Tile_X0Y10_B_I_top),
    .B_T_top(Tile_X0Y10_B_T_top),
    .A_config_C_bit0(Tile_X0Y10_A_config_C_bit0),
    .A_config_C_bit1(Tile_X0Y10_A_config_C_bit1),
    .A_config_C_bit2(Tile_X0Y10_A_config_C_bit2),
    .A_config_C_bit3(Tile_X0Y10_A_config_C_bit3),
    .B_config_C_bit0(Tile_X0Y10_B_config_C_bit0),
    .B_config_C_bit1(Tile_X0Y10_B_config_C_bit1),
    .B_config_C_bit2(Tile_X0Y10_B_config_C_bit2),
    .B_config_C_bit3(Tile_X0Y10_B_config_C_bit3),
    .UserCLK(Tile_X0Y11_UserCLKo),
    .UserCLKo(Tile_X0Y10_UserCLKo),
    .FrameData(Row_Y10_FrameData),
    .FrameData_O(Tile_X0Y10_FrameData_O),
    .FrameStrobe(Tile_X0Y11_FrameStrobe_O),
    .FrameStrobe_O(Tile_X0Y10_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X1Y10_Emulate_Bitstream)
    )
`endif
    Tile_X1Y10_LUT4AB
    (
    .N1END(Tile_X1Y11_N1BEG),
    .N2MID(Tile_X1Y11_N2BEG),
    .N2END(Tile_X1Y11_N2BEGb),
    .N4END(Tile_X1Y11_N4BEG),
    .NN4END(Tile_X1Y11_NN4BEG),
    .Ci(Tile_X1Y11_Co),
    .E1END(Tile_X0Y10_E1BEG),
    .E2MID(Tile_X0Y10_E2BEG),
    .E2END(Tile_X0Y10_E2BEGb),
    .EE4END(Tile_X0Y10_EE4BEG),
    .E6END(Tile_X0Y10_E6BEG),
    .S1END(Tile_X1Y9_S1BEG),
    .S2MID(Tile_X1Y9_S2BEG),
    .S2END(Tile_X1Y9_S2BEGb),
    .S4END(Tile_X1Y9_S4BEG),
    .SS4END(Tile_X1Y9_SS4BEG),
    .W1END(Tile_X2Y10_W1BEG),
    .W2MID(Tile_X2Y10_W2BEG),
    .W2END(Tile_X2Y10_W2BEGb),
    .WW4END(Tile_X2Y10_WW4BEG),
    .W6END(Tile_X2Y10_W6BEG),
    .N1BEG(Tile_X1Y10_N1BEG),
    .N2BEG(Tile_X1Y10_N2BEG),
    .N2BEGb(Tile_X1Y10_N2BEGb),
    .N4BEG(Tile_X1Y10_N4BEG),
    .NN4BEG(Tile_X1Y10_NN4BEG),
    .E1BEG(Tile_X1Y10_E1BEG),
    .E2BEG(Tile_X1Y10_E2BEG),
    .E2BEGb(Tile_X1Y10_E2BEGb),
    .EE4BEG(Tile_X1Y10_EE4BEG),
    .E6BEG(Tile_X1Y10_E6BEG),
    .S1BEG(Tile_X1Y10_S1BEG),
    .S2BEG(Tile_X1Y10_S2BEG),
    .S2BEGb(Tile_X1Y10_S2BEGb),
    .S4BEG(Tile_X1Y10_S4BEG),
    .SS4BEG(Tile_X1Y10_SS4BEG),
    .W1BEG(Tile_X1Y10_W1BEG),
    .W2BEG(Tile_X1Y10_W2BEG),
    .W2BEGb(Tile_X1Y10_W2BEGb),
    .WW4BEG(Tile_X1Y10_WW4BEG),
    .W6BEG(Tile_X1Y10_W6BEG),
    .Co(Tile_X1Y10_Co),
    .UserCLK(Tile_X1Y11_UserCLKo),
    .UserCLKo(Tile_X1Y10_UserCLKo),
    .FrameData(Tile_X0Y10_FrameData_O),
    .FrameData_O(Tile_X1Y10_FrameData_O),
    .FrameStrobe(Tile_X1Y11_FrameStrobe_O),
    .FrameStrobe_O(Tile_X1Y10_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X2Y10_Emulate_Bitstream)
    )
`endif
    Tile_X2Y10_LUT4AB
    (
    .N1END(Tile_X2Y11_N1BEG),
    .N2MID(Tile_X2Y11_N2BEG),
    .N2END(Tile_X2Y11_N2BEGb),
    .N4END(Tile_X2Y11_N4BEG),
    .NN4END(Tile_X2Y11_NN4BEG),
    .Ci(Tile_X2Y11_Co),
    .E1END(Tile_X1Y10_E1BEG),
    .E2MID(Tile_X1Y10_E2BEG),
    .E2END(Tile_X1Y10_E2BEGb),
    .EE4END(Tile_X1Y10_EE4BEG),
    .E6END(Tile_X1Y10_E6BEG),
    .S1END(Tile_X2Y9_S1BEG),
    .S2MID(Tile_X2Y9_S2BEG),
    .S2END(Tile_X2Y9_S2BEGb),
    .S4END(Tile_X2Y9_S4BEG),
    .SS4END(Tile_X2Y9_SS4BEG),
    .W1END(Tile_X3Y10_W1BEG),
    .W2MID(Tile_X3Y10_W2BEG),
    .W2END(Tile_X3Y10_W2BEGb),
    .WW4END(Tile_X3Y10_WW4BEG),
    .W6END(Tile_X3Y10_W6BEG),
    .N1BEG(Tile_X2Y10_N1BEG),
    .N2BEG(Tile_X2Y10_N2BEG),
    .N2BEGb(Tile_X2Y10_N2BEGb),
    .N4BEG(Tile_X2Y10_N4BEG),
    .NN4BEG(Tile_X2Y10_NN4BEG),
    .E1BEG(Tile_X2Y10_E1BEG),
    .E2BEG(Tile_X2Y10_E2BEG),
    .E2BEGb(Tile_X2Y10_E2BEGb),
    .EE4BEG(Tile_X2Y10_EE4BEG),
    .E6BEG(Tile_X2Y10_E6BEG),
    .S1BEG(Tile_X2Y10_S1BEG),
    .S2BEG(Tile_X2Y10_S2BEG),
    .S2BEGb(Tile_X2Y10_S2BEGb),
    .S4BEG(Tile_X2Y10_S4BEG),
    .SS4BEG(Tile_X2Y10_SS4BEG),
    .W1BEG(Tile_X2Y10_W1BEG),
    .W2BEG(Tile_X2Y10_W2BEG),
    .W2BEGb(Tile_X2Y10_W2BEGb),
    .WW4BEG(Tile_X2Y10_WW4BEG),
    .W6BEG(Tile_X2Y10_W6BEG),
    .Co(Tile_X2Y10_Co),
    .UserCLK(Tile_X2Y11_UserCLKo),
    .UserCLKo(Tile_X2Y10_UserCLKo),
    .FrameData(Tile_X1Y10_FrameData_O),
    .FrameData_O(Tile_X2Y10_FrameData_O),
    .FrameStrobe(Tile_X2Y11_FrameStrobe_O),
    .FrameStrobe_O(Tile_X2Y10_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X3Y10_Emulate_Bitstream)
    )
`endif
    Tile_X3Y10_LUT4AB
    (
    .N1END(Tile_X3Y11_N1BEG),
    .N2MID(Tile_X3Y11_N2BEG),
    .N2END(Tile_X3Y11_N2BEGb),
    .N4END(Tile_X3Y11_N4BEG),
    .NN4END(Tile_X3Y11_NN4BEG),
    .Ci(Tile_X3Y11_Co),
    .E1END(Tile_X2Y10_E1BEG),
    .E2MID(Tile_X2Y10_E2BEG),
    .E2END(Tile_X2Y10_E2BEGb),
    .EE4END(Tile_X2Y10_EE4BEG),
    .E6END(Tile_X2Y10_E6BEG),
    .S1END(Tile_X3Y9_S1BEG),
    .S2MID(Tile_X3Y9_S2BEG),
    .S2END(Tile_X3Y9_S2BEGb),
    .S4END(Tile_X3Y9_S4BEG),
    .SS4END(Tile_X3Y9_SS4BEG),
    .W1END(Tile_X4Y10_W1BEG),
    .W2MID(Tile_X4Y10_W2BEG),
    .W2END(Tile_X4Y10_W2BEGb),
    .WW4END(Tile_X4Y10_WW4BEG),
    .W6END(Tile_X4Y10_W6BEG),
    .N1BEG(Tile_X3Y10_N1BEG),
    .N2BEG(Tile_X3Y10_N2BEG),
    .N2BEGb(Tile_X3Y10_N2BEGb),
    .N4BEG(Tile_X3Y10_N4BEG),
    .NN4BEG(Tile_X3Y10_NN4BEG),
    .E1BEG(Tile_X3Y10_E1BEG),
    .E2BEG(Tile_X3Y10_E2BEG),
    .E2BEGb(Tile_X3Y10_E2BEGb),
    .EE4BEG(Tile_X3Y10_EE4BEG),
    .E6BEG(Tile_X3Y10_E6BEG),
    .S1BEG(Tile_X3Y10_S1BEG),
    .S2BEG(Tile_X3Y10_S2BEG),
    .S2BEGb(Tile_X3Y10_S2BEGb),
    .S4BEG(Tile_X3Y10_S4BEG),
    .SS4BEG(Tile_X3Y10_SS4BEG),
    .W1BEG(Tile_X3Y10_W1BEG),
    .W2BEG(Tile_X3Y10_W2BEG),
    .W2BEGb(Tile_X3Y10_W2BEGb),
    .WW4BEG(Tile_X3Y10_WW4BEG),
    .W6BEG(Tile_X3Y10_W6BEG),
    .Co(Tile_X3Y10_Co),
    .UserCLK(Tile_X3Y11_UserCLKo),
    .UserCLKo(Tile_X3Y10_UserCLKo),
    .FrameData(Tile_X2Y10_FrameData_O),
    .FrameData_O(Tile_X3Y10_FrameData_O),
    .FrameStrobe(Tile_X3Y11_FrameStrobe_O),
    .FrameStrobe_O(Tile_X3Y10_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
RegFile
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X4Y10_Emulate_Bitstream)
    )
`endif
    Tile_X4Y10_RegFile
    (
    .N1END(Tile_X4Y11_N1BEG),
    .N2MID(Tile_X4Y11_N2BEG),
    .N2END(Tile_X4Y11_N2BEGb),
    .N4END(Tile_X4Y11_N4BEG),
    .NN4END(Tile_X4Y11_NN4BEG),
    .E1END(Tile_X3Y10_E1BEG),
    .E2MID(Tile_X3Y10_E2BEG),
    .E2END(Tile_X3Y10_E2BEGb),
    .EE4END(Tile_X3Y10_EE4BEG),
    .E6END(Tile_X3Y10_E6BEG),
    .S1END(Tile_X4Y9_S1BEG),
    .S2MID(Tile_X4Y9_S2BEG),
    .S2END(Tile_X4Y9_S2BEGb),
    .S4END(Tile_X4Y9_S4BEG),
    .SS4END(Tile_X4Y9_SS4BEG),
    .W1END(Tile_X5Y10_W1BEG),
    .W2MID(Tile_X5Y10_W2BEG),
    .W2END(Tile_X5Y10_W2BEGb),
    .WW4END(Tile_X5Y10_WW4BEG),
    .W6END(Tile_X5Y10_W6BEG),
    .N1BEG(Tile_X4Y10_N1BEG),
    .N2BEG(Tile_X4Y10_N2BEG),
    .N2BEGb(Tile_X4Y10_N2BEGb),
    .N4BEG(Tile_X4Y10_N4BEG),
    .NN4BEG(Tile_X4Y10_NN4BEG),
    .E1BEG(Tile_X4Y10_E1BEG),
    .E2BEG(Tile_X4Y10_E2BEG),
    .E2BEGb(Tile_X4Y10_E2BEGb),
    .EE4BEG(Tile_X4Y10_EE4BEG),
    .E6BEG(Tile_X4Y10_E6BEG),
    .S1BEG(Tile_X4Y10_S1BEG),
    .S2BEG(Tile_X4Y10_S2BEG),
    .S2BEGb(Tile_X4Y10_S2BEGb),
    .S4BEG(Tile_X4Y10_S4BEG),
    .SS4BEG(Tile_X4Y10_SS4BEG),
    .W1BEG(Tile_X4Y10_W1BEG),
    .W2BEG(Tile_X4Y10_W2BEG),
    .W2BEGb(Tile_X4Y10_W2BEGb),
    .WW4BEG(Tile_X4Y10_WW4BEG),
    .W6BEG(Tile_X4Y10_W6BEG),
    .UserCLK(Tile_X4Y11_UserCLKo),
    .UserCLKo(Tile_X4Y10_UserCLKo),
    .FrameData(Tile_X3Y10_FrameData_O),
    .FrameData_O(Tile_X4Y10_FrameData_O),
    .FrameStrobe(Tile_X4Y11_FrameStrobe_O),
    .FrameStrobe_O(Tile_X4Y10_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X5Y10_Emulate_Bitstream)
    )
`endif
    Tile_X5Y10_LUT4AB
    (
    .N1END(Tile_X5Y11_N1BEG),
    .N2MID(Tile_X5Y11_N2BEG),
    .N2END(Tile_X5Y11_N2BEGb),
    .N4END(Tile_X5Y11_N4BEG),
    .NN4END(Tile_X5Y11_NN4BEG),
    .Ci(Tile_X5Y11_Co),
    .E1END(Tile_X4Y10_E1BEG),
    .E2MID(Tile_X4Y10_E2BEG),
    .E2END(Tile_X4Y10_E2BEGb),
    .EE4END(Tile_X4Y10_EE4BEG),
    .E6END(Tile_X4Y10_E6BEG),
    .S1END(Tile_X5Y9_S1BEG),
    .S2MID(Tile_X5Y9_S2BEG),
    .S2END(Tile_X5Y9_S2BEGb),
    .S4END(Tile_X5Y9_S4BEG),
    .SS4END(Tile_X5Y9_SS4BEG),
    .W1END(Tile_X6Y10_W1BEG),
    .W2MID(Tile_X6Y10_W2BEG),
    .W2END(Tile_X6Y10_W2BEGb),
    .WW4END(Tile_X6Y10_WW4BEG),
    .W6END(Tile_X6Y10_W6BEG),
    .N1BEG(Tile_X5Y10_N1BEG),
    .N2BEG(Tile_X5Y10_N2BEG),
    .N2BEGb(Tile_X5Y10_N2BEGb),
    .N4BEG(Tile_X5Y10_N4BEG),
    .NN4BEG(Tile_X5Y10_NN4BEG),
    .E1BEG(Tile_X5Y10_E1BEG),
    .E2BEG(Tile_X5Y10_E2BEG),
    .E2BEGb(Tile_X5Y10_E2BEGb),
    .EE4BEG(Tile_X5Y10_EE4BEG),
    .E6BEG(Tile_X5Y10_E6BEG),
    .S1BEG(Tile_X5Y10_S1BEG),
    .S2BEG(Tile_X5Y10_S2BEG),
    .S2BEGb(Tile_X5Y10_S2BEGb),
    .S4BEG(Tile_X5Y10_S4BEG),
    .SS4BEG(Tile_X5Y10_SS4BEG),
    .W1BEG(Tile_X5Y10_W1BEG),
    .W2BEG(Tile_X5Y10_W2BEG),
    .W2BEGb(Tile_X5Y10_W2BEGb),
    .WW4BEG(Tile_X5Y10_WW4BEG),
    .W6BEG(Tile_X5Y10_W6BEG),
    .Co(Tile_X5Y10_Co),
    .UserCLK(Tile_X5Y11_UserCLKo),
    .UserCLKo(Tile_X5Y10_UserCLKo),
    .FrameData(Tile_X4Y10_FrameData_O),
    .FrameData_O(Tile_X5Y10_FrameData_O),
    .FrameStrobe(Tile_X5Y11_FrameStrobe_O),
    .FrameStrobe_O(Tile_X5Y10_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X6Y10_Emulate_Bitstream)
    )
`endif
    Tile_X6Y10_LUT4AB
    (
    .N1END(Tile_X6Y11_N1BEG),
    .N2MID(Tile_X6Y11_N2BEG),
    .N2END(Tile_X6Y11_N2BEGb),
    .N4END(Tile_X6Y11_N4BEG),
    .NN4END(Tile_X6Y11_NN4BEG),
    .Ci(Tile_X6Y11_Co),
    .E1END(Tile_X5Y10_E1BEG),
    .E2MID(Tile_X5Y10_E2BEG),
    .E2END(Tile_X5Y10_E2BEGb),
    .EE4END(Tile_X5Y10_EE4BEG),
    .E6END(Tile_X5Y10_E6BEG),
    .S1END(Tile_X6Y9_S1BEG),
    .S2MID(Tile_X6Y9_S2BEG),
    .S2END(Tile_X6Y9_S2BEGb),
    .S4END(Tile_X6Y9_S4BEG),
    .SS4END(Tile_X6Y9_SS4BEG),
    .W1END(Tile_X7Y10_W1BEG),
    .W2MID(Tile_X7Y10_W2BEG),
    .W2END(Tile_X7Y10_W2BEGb),
    .WW4END(Tile_X7Y10_WW4BEG),
    .W6END(Tile_X7Y10_W6BEG),
    .N1BEG(Tile_X6Y10_N1BEG),
    .N2BEG(Tile_X6Y10_N2BEG),
    .N2BEGb(Tile_X6Y10_N2BEGb),
    .N4BEG(Tile_X6Y10_N4BEG),
    .NN4BEG(Tile_X6Y10_NN4BEG),
    .E1BEG(Tile_X6Y10_E1BEG),
    .E2BEG(Tile_X6Y10_E2BEG),
    .E2BEGb(Tile_X6Y10_E2BEGb),
    .EE4BEG(Tile_X6Y10_EE4BEG),
    .E6BEG(Tile_X6Y10_E6BEG),
    .S1BEG(Tile_X6Y10_S1BEG),
    .S2BEG(Tile_X6Y10_S2BEG),
    .S2BEGb(Tile_X6Y10_S2BEGb),
    .S4BEG(Tile_X6Y10_S4BEG),
    .SS4BEG(Tile_X6Y10_SS4BEG),
    .W1BEG(Tile_X6Y10_W1BEG),
    .W2BEG(Tile_X6Y10_W2BEG),
    .W2BEGb(Tile_X6Y10_W2BEGb),
    .WW4BEG(Tile_X6Y10_WW4BEG),
    .W6BEG(Tile_X6Y10_W6BEG),
    .Co(Tile_X6Y10_Co),
    .UserCLK(Tile_X6Y11_UserCLKo),
    .UserCLKo(Tile_X6Y10_UserCLKo),
    .FrameData(Tile_X5Y10_FrameData_O),
    .FrameData_O(Tile_X6Y10_FrameData_O),
    .FrameStrobe(Tile_X6Y11_FrameStrobe_O),
    .FrameStrobe_O(Tile_X6Y10_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X8Y10_Emulate_Bitstream)
    )
`endif
    Tile_X8Y10_LUT4AB
    (
    .N1END(Tile_X8Y11_N1BEG),
    .N2MID(Tile_X8Y11_N2BEG),
    .N2END(Tile_X8Y11_N2BEGb),
    .N4END(Tile_X8Y11_N4BEG),
    .NN4END(Tile_X8Y11_NN4BEG),
    .Ci(Tile_X8Y11_Co),
    .E1END(Tile_X7Y10_E1BEG),
    .E2MID(Tile_X7Y10_E2BEG),
    .E2END(Tile_X7Y10_E2BEGb),
    .EE4END(Tile_X7Y10_EE4BEG),
    .E6END(Tile_X7Y10_E6BEG),
    .S1END(Tile_X8Y9_S1BEG),
    .S2MID(Tile_X8Y9_S2BEG),
    .S2END(Tile_X8Y9_S2BEGb),
    .S4END(Tile_X8Y9_S4BEG),
    .SS4END(Tile_X8Y9_SS4BEG),
    .W1END(Tile_X9Y10_W1BEG),
    .W2MID(Tile_X9Y10_W2BEG),
    .W2END(Tile_X9Y10_W2BEGb),
    .WW4END(Tile_X9Y10_WW4BEG),
    .W6END(Tile_X9Y10_W6BEG),
    .N1BEG(Tile_X8Y10_N1BEG),
    .N2BEG(Tile_X8Y10_N2BEG),
    .N2BEGb(Tile_X8Y10_N2BEGb),
    .N4BEG(Tile_X8Y10_N4BEG),
    .NN4BEG(Tile_X8Y10_NN4BEG),
    .E1BEG(Tile_X8Y10_E1BEG),
    .E2BEG(Tile_X8Y10_E2BEG),
    .E2BEGb(Tile_X8Y10_E2BEGb),
    .EE4BEG(Tile_X8Y10_EE4BEG),
    .E6BEG(Tile_X8Y10_E6BEG),
    .S1BEG(Tile_X8Y10_S1BEG),
    .S2BEG(Tile_X8Y10_S2BEG),
    .S2BEGb(Tile_X8Y10_S2BEGb),
    .S4BEG(Tile_X8Y10_S4BEG),
    .SS4BEG(Tile_X8Y10_SS4BEG),
    .W1BEG(Tile_X8Y10_W1BEG),
    .W2BEG(Tile_X8Y10_W2BEG),
    .W2BEGb(Tile_X8Y10_W2BEGb),
    .WW4BEG(Tile_X8Y10_WW4BEG),
    .W6BEG(Tile_X8Y10_W6BEG),
    .Co(Tile_X8Y10_Co),
    .UserCLK(Tile_X8Y11_UserCLKo),
    .UserCLKo(Tile_X8Y10_UserCLKo),
    .FrameData(Tile_X7Y10_FrameData_O),
    .FrameData_O(Tile_X8Y10_FrameData_O),
    .FrameStrobe(Tile_X8Y11_FrameStrobe_O),
    .FrameStrobe_O(Tile_X8Y10_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X9Y10_Emulate_Bitstream)
    )
`endif
    Tile_X9Y10_LUT4AB
    (
    .N1END(Tile_X9Y11_N1BEG),
    .N2MID(Tile_X9Y11_N2BEG),
    .N2END(Tile_X9Y11_N2BEGb),
    .N4END(Tile_X9Y11_N4BEG),
    .NN4END(Tile_X9Y11_NN4BEG),
    .Ci(Tile_X9Y11_Co),
    .E1END(Tile_X8Y10_E1BEG),
    .E2MID(Tile_X8Y10_E2BEG),
    .E2END(Tile_X8Y10_E2BEGb),
    .EE4END(Tile_X8Y10_EE4BEG),
    .E6END(Tile_X8Y10_E6BEG),
    .S1END(Tile_X9Y9_S1BEG),
    .S2MID(Tile_X9Y9_S2BEG),
    .S2END(Tile_X9Y9_S2BEGb),
    .S4END(Tile_X9Y9_S4BEG),
    .SS4END(Tile_X9Y9_SS4BEG),
    .W1END(Tile_X10Y10_W1BEG),
    .W2MID(Tile_X10Y10_W2BEG),
    .W2END(Tile_X10Y10_W2BEGb),
    .WW4END(Tile_X10Y10_WW4BEG),
    .W6END(Tile_X10Y10_W6BEG),
    .N1BEG(Tile_X9Y10_N1BEG),
    .N2BEG(Tile_X9Y10_N2BEG),
    .N2BEGb(Tile_X9Y10_N2BEGb),
    .N4BEG(Tile_X9Y10_N4BEG),
    .NN4BEG(Tile_X9Y10_NN4BEG),
    .E1BEG(Tile_X9Y10_E1BEG),
    .E2BEG(Tile_X9Y10_E2BEG),
    .E2BEGb(Tile_X9Y10_E2BEGb),
    .EE4BEG(Tile_X9Y10_EE4BEG),
    .E6BEG(Tile_X9Y10_E6BEG),
    .S1BEG(Tile_X9Y10_S1BEG),
    .S2BEG(Tile_X9Y10_S2BEG),
    .S2BEGb(Tile_X9Y10_S2BEGb),
    .S4BEG(Tile_X9Y10_S4BEG),
    .SS4BEG(Tile_X9Y10_SS4BEG),
    .W1BEG(Tile_X9Y10_W1BEG),
    .W2BEG(Tile_X9Y10_W2BEG),
    .W2BEGb(Tile_X9Y10_W2BEGb),
    .WW4BEG(Tile_X9Y10_WW4BEG),
    .W6BEG(Tile_X9Y10_W6BEG),
    .Co(Tile_X9Y10_Co),
    .UserCLK(Tile_X9Y11_UserCLKo),
    .UserCLKo(Tile_X9Y10_UserCLKo),
    .FrameData(Tile_X8Y10_FrameData_O),
    .FrameData_O(Tile_X9Y10_FrameData_O),
    .FrameStrobe(Tile_X9Y11_FrameStrobe_O),
    .FrameStrobe_O(Tile_X9Y10_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
W_IO
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X0Y11_Emulate_Bitstream)
    )
`endif
    Tile_X0Y11_W_IO
    (
    .W1END(Tile_X1Y11_W1BEG),
    .W2MID(Tile_X1Y11_W2BEG),
    .W2END(Tile_X1Y11_W2BEGb),
    .WW4END(Tile_X1Y11_WW4BEG),
    .W6END(Tile_X1Y11_W6BEG),
    .E1BEG(Tile_X0Y11_E1BEG),
    .E2BEG(Tile_X0Y11_E2BEG),
    .E2BEGb(Tile_X0Y11_E2BEGb),
    .EE4BEG(Tile_X0Y11_EE4BEG),
    .E6BEG(Tile_X0Y11_E6BEG),
    .A_O_top(Tile_X0Y11_A_O_top),
    .A_I_top(Tile_X0Y11_A_I_top),
    .A_T_top(Tile_X0Y11_A_T_top),
    .B_O_top(Tile_X0Y11_B_O_top),
    .B_I_top(Tile_X0Y11_B_I_top),
    .B_T_top(Tile_X0Y11_B_T_top),
    .A_config_C_bit0(Tile_X0Y11_A_config_C_bit0),
    .A_config_C_bit1(Tile_X0Y11_A_config_C_bit1),
    .A_config_C_bit2(Tile_X0Y11_A_config_C_bit2),
    .A_config_C_bit3(Tile_X0Y11_A_config_C_bit3),
    .B_config_C_bit0(Tile_X0Y11_B_config_C_bit0),
    .B_config_C_bit1(Tile_X0Y11_B_config_C_bit1),
    .B_config_C_bit2(Tile_X0Y11_B_config_C_bit2),
    .B_config_C_bit3(Tile_X0Y11_B_config_C_bit3),
    .UserCLK(Tile_X0Y12_UserCLKo),
    .UserCLKo(Tile_X0Y11_UserCLKo),
    .FrameData(Row_Y11_FrameData),
    .FrameData_O(Tile_X0Y11_FrameData_O),
    .FrameStrobe(Tile_X0Y12_FrameStrobe_O),
    .FrameStrobe_O(Tile_X0Y11_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X1Y11_Emulate_Bitstream)
    )
`endif
    Tile_X1Y11_LUT4AB
    (
    .N1END(Tile_X1Y12_N1BEG),
    .N2MID(Tile_X1Y12_N2BEG),
    .N2END(Tile_X1Y12_N2BEGb),
    .N4END(Tile_X1Y12_N4BEG),
    .NN4END(Tile_X1Y12_NN4BEG),
    .Ci(Tile_X1Y12_Co),
    .E1END(Tile_X0Y11_E1BEG),
    .E2MID(Tile_X0Y11_E2BEG),
    .E2END(Tile_X0Y11_E2BEGb),
    .EE4END(Tile_X0Y11_EE4BEG),
    .E6END(Tile_X0Y11_E6BEG),
    .S1END(Tile_X1Y10_S1BEG),
    .S2MID(Tile_X1Y10_S2BEG),
    .S2END(Tile_X1Y10_S2BEGb),
    .S4END(Tile_X1Y10_S4BEG),
    .SS4END(Tile_X1Y10_SS4BEG),
    .W1END(Tile_X2Y11_W1BEG),
    .W2MID(Tile_X2Y11_W2BEG),
    .W2END(Tile_X2Y11_W2BEGb),
    .WW4END(Tile_X2Y11_WW4BEG),
    .W6END(Tile_X2Y11_W6BEG),
    .N1BEG(Tile_X1Y11_N1BEG),
    .N2BEG(Tile_X1Y11_N2BEG),
    .N2BEGb(Tile_X1Y11_N2BEGb),
    .N4BEG(Tile_X1Y11_N4BEG),
    .NN4BEG(Tile_X1Y11_NN4BEG),
    .E1BEG(Tile_X1Y11_E1BEG),
    .E2BEG(Tile_X1Y11_E2BEG),
    .E2BEGb(Tile_X1Y11_E2BEGb),
    .EE4BEG(Tile_X1Y11_EE4BEG),
    .E6BEG(Tile_X1Y11_E6BEG),
    .S1BEG(Tile_X1Y11_S1BEG),
    .S2BEG(Tile_X1Y11_S2BEG),
    .S2BEGb(Tile_X1Y11_S2BEGb),
    .S4BEG(Tile_X1Y11_S4BEG),
    .SS4BEG(Tile_X1Y11_SS4BEG),
    .W1BEG(Tile_X1Y11_W1BEG),
    .W2BEG(Tile_X1Y11_W2BEG),
    .W2BEGb(Tile_X1Y11_W2BEGb),
    .WW4BEG(Tile_X1Y11_WW4BEG),
    .W6BEG(Tile_X1Y11_W6BEG),
    .Co(Tile_X1Y11_Co),
    .UserCLK(Tile_X1Y12_UserCLKo),
    .UserCLKo(Tile_X1Y11_UserCLKo),
    .FrameData(Tile_X0Y11_FrameData_O),
    .FrameData_O(Tile_X1Y11_FrameData_O),
    .FrameStrobe(Tile_X1Y12_FrameStrobe_O),
    .FrameStrobe_O(Tile_X1Y11_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X2Y11_Emulate_Bitstream)
    )
`endif
    Tile_X2Y11_LUT4AB
    (
    .N1END(Tile_X2Y12_N1BEG),
    .N2MID(Tile_X2Y12_N2BEG),
    .N2END(Tile_X2Y12_N2BEGb),
    .N4END(Tile_X2Y12_N4BEG),
    .NN4END(Tile_X2Y12_NN4BEG),
    .Ci(Tile_X2Y12_Co),
    .E1END(Tile_X1Y11_E1BEG),
    .E2MID(Tile_X1Y11_E2BEG),
    .E2END(Tile_X1Y11_E2BEGb),
    .EE4END(Tile_X1Y11_EE4BEG),
    .E6END(Tile_X1Y11_E6BEG),
    .S1END(Tile_X2Y10_S1BEG),
    .S2MID(Tile_X2Y10_S2BEG),
    .S2END(Tile_X2Y10_S2BEGb),
    .S4END(Tile_X2Y10_S4BEG),
    .SS4END(Tile_X2Y10_SS4BEG),
    .W1END(Tile_X3Y11_W1BEG),
    .W2MID(Tile_X3Y11_W2BEG),
    .W2END(Tile_X3Y11_W2BEGb),
    .WW4END(Tile_X3Y11_WW4BEG),
    .W6END(Tile_X3Y11_W6BEG),
    .N1BEG(Tile_X2Y11_N1BEG),
    .N2BEG(Tile_X2Y11_N2BEG),
    .N2BEGb(Tile_X2Y11_N2BEGb),
    .N4BEG(Tile_X2Y11_N4BEG),
    .NN4BEG(Tile_X2Y11_NN4BEG),
    .E1BEG(Tile_X2Y11_E1BEG),
    .E2BEG(Tile_X2Y11_E2BEG),
    .E2BEGb(Tile_X2Y11_E2BEGb),
    .EE4BEG(Tile_X2Y11_EE4BEG),
    .E6BEG(Tile_X2Y11_E6BEG),
    .S1BEG(Tile_X2Y11_S1BEG),
    .S2BEG(Tile_X2Y11_S2BEG),
    .S2BEGb(Tile_X2Y11_S2BEGb),
    .S4BEG(Tile_X2Y11_S4BEG),
    .SS4BEG(Tile_X2Y11_SS4BEG),
    .W1BEG(Tile_X2Y11_W1BEG),
    .W2BEG(Tile_X2Y11_W2BEG),
    .W2BEGb(Tile_X2Y11_W2BEGb),
    .WW4BEG(Tile_X2Y11_WW4BEG),
    .W6BEG(Tile_X2Y11_W6BEG),
    .Co(Tile_X2Y11_Co),
    .UserCLK(Tile_X2Y12_UserCLKo),
    .UserCLKo(Tile_X2Y11_UserCLKo),
    .FrameData(Tile_X1Y11_FrameData_O),
    .FrameData_O(Tile_X2Y11_FrameData_O),
    .FrameStrobe(Tile_X2Y12_FrameStrobe_O),
    .FrameStrobe_O(Tile_X2Y11_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X3Y11_Emulate_Bitstream)
    )
`endif
    Tile_X3Y11_LUT4AB
    (
    .N1END(Tile_X3Y12_N1BEG),
    .N2MID(Tile_X3Y12_N2BEG),
    .N2END(Tile_X3Y12_N2BEGb),
    .N4END(Tile_X3Y12_N4BEG),
    .NN4END(Tile_X3Y12_NN4BEG),
    .Ci(Tile_X3Y12_Co),
    .E1END(Tile_X2Y11_E1BEG),
    .E2MID(Tile_X2Y11_E2BEG),
    .E2END(Tile_X2Y11_E2BEGb),
    .EE4END(Tile_X2Y11_EE4BEG),
    .E6END(Tile_X2Y11_E6BEG),
    .S1END(Tile_X3Y10_S1BEG),
    .S2MID(Tile_X3Y10_S2BEG),
    .S2END(Tile_X3Y10_S2BEGb),
    .S4END(Tile_X3Y10_S4BEG),
    .SS4END(Tile_X3Y10_SS4BEG),
    .W1END(Tile_X4Y11_W1BEG),
    .W2MID(Tile_X4Y11_W2BEG),
    .W2END(Tile_X4Y11_W2BEGb),
    .WW4END(Tile_X4Y11_WW4BEG),
    .W6END(Tile_X4Y11_W6BEG),
    .N1BEG(Tile_X3Y11_N1BEG),
    .N2BEG(Tile_X3Y11_N2BEG),
    .N2BEGb(Tile_X3Y11_N2BEGb),
    .N4BEG(Tile_X3Y11_N4BEG),
    .NN4BEG(Tile_X3Y11_NN4BEG),
    .E1BEG(Tile_X3Y11_E1BEG),
    .E2BEG(Tile_X3Y11_E2BEG),
    .E2BEGb(Tile_X3Y11_E2BEGb),
    .EE4BEG(Tile_X3Y11_EE4BEG),
    .E6BEG(Tile_X3Y11_E6BEG),
    .S1BEG(Tile_X3Y11_S1BEG),
    .S2BEG(Tile_X3Y11_S2BEG),
    .S2BEGb(Tile_X3Y11_S2BEGb),
    .S4BEG(Tile_X3Y11_S4BEG),
    .SS4BEG(Tile_X3Y11_SS4BEG),
    .W1BEG(Tile_X3Y11_W1BEG),
    .W2BEG(Tile_X3Y11_W2BEG),
    .W2BEGb(Tile_X3Y11_W2BEGb),
    .WW4BEG(Tile_X3Y11_WW4BEG),
    .W6BEG(Tile_X3Y11_W6BEG),
    .Co(Tile_X3Y11_Co),
    .UserCLK(Tile_X3Y12_UserCLKo),
    .UserCLKo(Tile_X3Y11_UserCLKo),
    .FrameData(Tile_X2Y11_FrameData_O),
    .FrameData_O(Tile_X3Y11_FrameData_O),
    .FrameStrobe(Tile_X3Y12_FrameStrobe_O),
    .FrameStrobe_O(Tile_X3Y11_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
RegFile
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X4Y11_Emulate_Bitstream)
    )
`endif
    Tile_X4Y11_RegFile
    (
    .N1END(Tile_X4Y12_N1BEG),
    .N2MID(Tile_X4Y12_N2BEG),
    .N2END(Tile_X4Y12_N2BEGb),
    .N4END(Tile_X4Y12_N4BEG),
    .NN4END(Tile_X4Y12_NN4BEG),
    .E1END(Tile_X3Y11_E1BEG),
    .E2MID(Tile_X3Y11_E2BEG),
    .E2END(Tile_X3Y11_E2BEGb),
    .EE4END(Tile_X3Y11_EE4BEG),
    .E6END(Tile_X3Y11_E6BEG),
    .S1END(Tile_X4Y10_S1BEG),
    .S2MID(Tile_X4Y10_S2BEG),
    .S2END(Tile_X4Y10_S2BEGb),
    .S4END(Tile_X4Y10_S4BEG),
    .SS4END(Tile_X4Y10_SS4BEG),
    .W1END(Tile_X5Y11_W1BEG),
    .W2MID(Tile_X5Y11_W2BEG),
    .W2END(Tile_X5Y11_W2BEGb),
    .WW4END(Tile_X5Y11_WW4BEG),
    .W6END(Tile_X5Y11_W6BEG),
    .N1BEG(Tile_X4Y11_N1BEG),
    .N2BEG(Tile_X4Y11_N2BEG),
    .N2BEGb(Tile_X4Y11_N2BEGb),
    .N4BEG(Tile_X4Y11_N4BEG),
    .NN4BEG(Tile_X4Y11_NN4BEG),
    .E1BEG(Tile_X4Y11_E1BEG),
    .E2BEG(Tile_X4Y11_E2BEG),
    .E2BEGb(Tile_X4Y11_E2BEGb),
    .EE4BEG(Tile_X4Y11_EE4BEG),
    .E6BEG(Tile_X4Y11_E6BEG),
    .S1BEG(Tile_X4Y11_S1BEG),
    .S2BEG(Tile_X4Y11_S2BEG),
    .S2BEGb(Tile_X4Y11_S2BEGb),
    .S4BEG(Tile_X4Y11_S4BEG),
    .SS4BEG(Tile_X4Y11_SS4BEG),
    .W1BEG(Tile_X4Y11_W1BEG),
    .W2BEG(Tile_X4Y11_W2BEG),
    .W2BEGb(Tile_X4Y11_W2BEGb),
    .WW4BEG(Tile_X4Y11_WW4BEG),
    .W6BEG(Tile_X4Y11_W6BEG),
    .UserCLK(Tile_X4Y12_UserCLKo),
    .UserCLKo(Tile_X4Y11_UserCLKo),
    .FrameData(Tile_X3Y11_FrameData_O),
    .FrameData_O(Tile_X4Y11_FrameData_O),
    .FrameStrobe(Tile_X4Y12_FrameStrobe_O),
    .FrameStrobe_O(Tile_X4Y11_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X5Y11_Emulate_Bitstream)
    )
`endif
    Tile_X5Y11_LUT4AB
    (
    .N1END(Tile_X5Y12_N1BEG),
    .N2MID(Tile_X5Y12_N2BEG),
    .N2END(Tile_X5Y12_N2BEGb),
    .N4END(Tile_X5Y12_N4BEG),
    .NN4END(Tile_X5Y12_NN4BEG),
    .Ci(Tile_X5Y12_Co),
    .E1END(Tile_X4Y11_E1BEG),
    .E2MID(Tile_X4Y11_E2BEG),
    .E2END(Tile_X4Y11_E2BEGb),
    .EE4END(Tile_X4Y11_EE4BEG),
    .E6END(Tile_X4Y11_E6BEG),
    .S1END(Tile_X5Y10_S1BEG),
    .S2MID(Tile_X5Y10_S2BEG),
    .S2END(Tile_X5Y10_S2BEGb),
    .S4END(Tile_X5Y10_S4BEG),
    .SS4END(Tile_X5Y10_SS4BEG),
    .W1END(Tile_X6Y11_W1BEG),
    .W2MID(Tile_X6Y11_W2BEG),
    .W2END(Tile_X6Y11_W2BEGb),
    .WW4END(Tile_X6Y11_WW4BEG),
    .W6END(Tile_X6Y11_W6BEG),
    .N1BEG(Tile_X5Y11_N1BEG),
    .N2BEG(Tile_X5Y11_N2BEG),
    .N2BEGb(Tile_X5Y11_N2BEGb),
    .N4BEG(Tile_X5Y11_N4BEG),
    .NN4BEG(Tile_X5Y11_NN4BEG),
    .E1BEG(Tile_X5Y11_E1BEG),
    .E2BEG(Tile_X5Y11_E2BEG),
    .E2BEGb(Tile_X5Y11_E2BEGb),
    .EE4BEG(Tile_X5Y11_EE4BEG),
    .E6BEG(Tile_X5Y11_E6BEG),
    .S1BEG(Tile_X5Y11_S1BEG),
    .S2BEG(Tile_X5Y11_S2BEG),
    .S2BEGb(Tile_X5Y11_S2BEGb),
    .S4BEG(Tile_X5Y11_S4BEG),
    .SS4BEG(Tile_X5Y11_SS4BEG),
    .W1BEG(Tile_X5Y11_W1BEG),
    .W2BEG(Tile_X5Y11_W2BEG),
    .W2BEGb(Tile_X5Y11_W2BEGb),
    .WW4BEG(Tile_X5Y11_WW4BEG),
    .W6BEG(Tile_X5Y11_W6BEG),
    .Co(Tile_X5Y11_Co),
    .UserCLK(Tile_X5Y12_UserCLKo),
    .UserCLKo(Tile_X5Y11_UserCLKo),
    .FrameData(Tile_X4Y11_FrameData_O),
    .FrameData_O(Tile_X5Y11_FrameData_O),
    .FrameStrobe(Tile_X5Y12_FrameStrobe_O),
    .FrameStrobe_O(Tile_X5Y11_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X6Y11_Emulate_Bitstream)
    )
`endif
    Tile_X6Y11_LUT4AB
    (
    .N1END(Tile_X6Y12_N1BEG),
    .N2MID(Tile_X6Y12_N2BEG),
    .N2END(Tile_X6Y12_N2BEGb),
    .N4END(Tile_X6Y12_N4BEG),
    .NN4END(Tile_X6Y12_NN4BEG),
    .Ci(Tile_X6Y12_Co),
    .E1END(Tile_X5Y11_E1BEG),
    .E2MID(Tile_X5Y11_E2BEG),
    .E2END(Tile_X5Y11_E2BEGb),
    .EE4END(Tile_X5Y11_EE4BEG),
    .E6END(Tile_X5Y11_E6BEG),
    .S1END(Tile_X6Y10_S1BEG),
    .S2MID(Tile_X6Y10_S2BEG),
    .S2END(Tile_X6Y10_S2BEGb),
    .S4END(Tile_X6Y10_S4BEG),
    .SS4END(Tile_X6Y10_SS4BEG),
    .W1END(Tile_X7Y11_W1BEG),
    .W2MID(Tile_X7Y11_W2BEG),
    .W2END(Tile_X7Y11_W2BEGb),
    .WW4END(Tile_X7Y11_WW4BEG),
    .W6END(Tile_X7Y11_W6BEG),
    .N1BEG(Tile_X6Y11_N1BEG),
    .N2BEG(Tile_X6Y11_N2BEG),
    .N2BEGb(Tile_X6Y11_N2BEGb),
    .N4BEG(Tile_X6Y11_N4BEG),
    .NN4BEG(Tile_X6Y11_NN4BEG),
    .E1BEG(Tile_X6Y11_E1BEG),
    .E2BEG(Tile_X6Y11_E2BEG),
    .E2BEGb(Tile_X6Y11_E2BEGb),
    .EE4BEG(Tile_X6Y11_EE4BEG),
    .E6BEG(Tile_X6Y11_E6BEG),
    .S1BEG(Tile_X6Y11_S1BEG),
    .S2BEG(Tile_X6Y11_S2BEG),
    .S2BEGb(Tile_X6Y11_S2BEGb),
    .S4BEG(Tile_X6Y11_S4BEG),
    .SS4BEG(Tile_X6Y11_SS4BEG),
    .W1BEG(Tile_X6Y11_W1BEG),
    .W2BEG(Tile_X6Y11_W2BEG),
    .W2BEGb(Tile_X6Y11_W2BEGb),
    .WW4BEG(Tile_X6Y11_WW4BEG),
    .W6BEG(Tile_X6Y11_W6BEG),
    .Co(Tile_X6Y11_Co),
    .UserCLK(Tile_X6Y12_UserCLKo),
    .UserCLKo(Tile_X6Y11_UserCLKo),
    .FrameData(Tile_X5Y11_FrameData_O),
    .FrameData_O(Tile_X6Y11_FrameData_O),
    .FrameStrobe(Tile_X6Y12_FrameStrobe_O),
    .FrameStrobe_O(Tile_X6Y11_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
DSP
`ifdef EMULATION
    #(
    .Tile_X0Y0_Emulate_Bitstream(`Tile_X7Y11_Emulate_Bitstream),
    .Tile_X0Y1_Emulate_Bitstream(`Tile_X7Y12_Emulate_Bitstream)
    )
`endif
    Tile_X7Y11_DSP
    (
    .Tile_X0Y0_E1END(Tile_X6Y11_E1BEG),
    .Tile_X0Y0_E2MID(Tile_X6Y11_E2BEG),
    .Tile_X0Y0_E2END(Tile_X6Y11_E2BEGb),
    .Tile_X0Y0_EE4END(Tile_X6Y11_EE4BEG),
    .Tile_X0Y0_E6END(Tile_X6Y11_E6BEG),
    .Tile_X0Y0_S1END(Tile_X7Y10_S1BEG),
    .Tile_X0Y0_S2MID(Tile_X7Y10_S2BEG),
    .Tile_X0Y0_S2END(Tile_X7Y10_S2BEGb),
    .Tile_X0Y0_S4END(Tile_X7Y10_S4BEG),
    .Tile_X0Y0_SS4END(Tile_X7Y10_SS4BEG),
    .Tile_X0Y0_W1END(Tile_X8Y11_W1BEG),
    .Tile_X0Y0_W2MID(Tile_X8Y11_W2BEG),
    .Tile_X0Y0_W2END(Tile_X8Y11_W2BEGb),
    .Tile_X0Y0_WW4END(Tile_X8Y11_WW4BEG),
    .Tile_X0Y0_W6END(Tile_X8Y11_W6BEG),
    .Tile_X0Y1_N1END(Tile_X7Y13_N1BEG),
    .Tile_X0Y1_N2MID(Tile_X7Y13_N2BEG),
    .Tile_X0Y1_N2END(Tile_X7Y13_N2BEGb),
    .Tile_X0Y1_N4END(Tile_X7Y13_N4BEG),
    .Tile_X0Y1_NN4END(Tile_X7Y13_NN4BEG),
    .Tile_X0Y1_E1END(Tile_X6Y12_E1BEG),
    .Tile_X0Y1_E2MID(Tile_X6Y12_E2BEG),
    .Tile_X0Y1_E2END(Tile_X6Y12_E2BEGb),
    .Tile_X0Y1_EE4END(Tile_X6Y12_EE4BEG),
    .Tile_X0Y1_E6END(Tile_X6Y12_E6BEG),
    .Tile_X0Y1_W1END(Tile_X8Y12_W1BEG),
    .Tile_X0Y1_W2MID(Tile_X8Y12_W2BEG),
    .Tile_X0Y1_W2END(Tile_X8Y12_W2BEGb),
    .Tile_X0Y1_WW4END(Tile_X8Y12_WW4BEG),
    .Tile_X0Y1_W6END(Tile_X8Y12_W6BEG),
    .Tile_X0Y0_N1BEG(Tile_X7Y11_N1BEG),
    .Tile_X0Y0_N2BEG(Tile_X7Y11_N2BEG),
    .Tile_X0Y0_N2BEGb(Tile_X7Y11_N2BEGb),
    .Tile_X0Y0_N4BEG(Tile_X7Y11_N4BEG),
    .Tile_X0Y0_NN4BEG(Tile_X7Y11_NN4BEG),
    .Tile_X0Y0_E1BEG(Tile_X7Y11_E1BEG),
    .Tile_X0Y0_E2BEG(Tile_X7Y11_E2BEG),
    .Tile_X0Y0_E2BEGb(Tile_X7Y11_E2BEGb),
    .Tile_X0Y0_EE4BEG(Tile_X7Y11_EE4BEG),
    .Tile_X0Y0_E6BEG(Tile_X7Y11_E6BEG),
    .Tile_X0Y0_W1BEG(Tile_X7Y11_W1BEG),
    .Tile_X0Y0_W2BEG(Tile_X7Y11_W2BEG),
    .Tile_X0Y0_W2BEGb(Tile_X7Y11_W2BEGb),
    .Tile_X0Y0_WW4BEG(Tile_X7Y11_WW4BEG),
    .Tile_X0Y0_W6BEG(Tile_X7Y11_W6BEG),
    .Tile_X0Y1_E1BEG(Tile_X7Y12_E1BEG),
    .Tile_X0Y1_E2BEG(Tile_X7Y12_E2BEG),
    .Tile_X0Y1_E2BEGb(Tile_X7Y12_E2BEGb),
    .Tile_X0Y1_EE4BEG(Tile_X7Y12_EE4BEG),
    .Tile_X0Y1_E6BEG(Tile_X7Y12_E6BEG),
    .Tile_X0Y1_S1BEG(Tile_X7Y12_S1BEG),
    .Tile_X0Y1_S2BEG(Tile_X7Y12_S2BEG),
    .Tile_X0Y1_S2BEGb(Tile_X7Y12_S2BEGb),
    .Tile_X0Y1_S4BEG(Tile_X7Y12_S4BEG),
    .Tile_X0Y1_SS4BEG(Tile_X7Y12_SS4BEG),
    .Tile_X0Y1_W1BEG(Tile_X7Y12_W1BEG),
    .Tile_X0Y1_W2BEG(Tile_X7Y12_W2BEG),
    .Tile_X0Y1_W2BEGb(Tile_X7Y12_W2BEGb),
    .Tile_X0Y1_WW4BEG(Tile_X7Y12_WW4BEG),
    .Tile_X0Y1_W6BEG(Tile_X7Y12_W6BEG),
    .Tile_X0Y0_UserCLKo(Tile_X7Y11_UserCLKo),
    .Tile_X0Y1_UserCLK(Tile_X7Y13_UserCLKo),
    .Tile_X0Y0_FrameData(Tile_X6Y11_FrameData_O),
    .Tile_X0Y0_FrameData_O(Tile_X7Y11_FrameData_O),
    .Tile_X0Y0_FrameStrobe_O(Tile_X7Y11_FrameStrobe_O),
    .Tile_X0Y1_FrameData(Tile_X6Y12_FrameData_O),
    .Tile_X0Y1_FrameData_O(Tile_X7Y12_FrameData_O),
    .Tile_X0Y1_FrameStrobe(Tile_X7Y13_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X8Y11_Emulate_Bitstream)
    )
`endif
    Tile_X8Y11_LUT4AB
    (
    .N1END(Tile_X8Y12_N1BEG),
    .N2MID(Tile_X8Y12_N2BEG),
    .N2END(Tile_X8Y12_N2BEGb),
    .N4END(Tile_X8Y12_N4BEG),
    .NN4END(Tile_X8Y12_NN4BEG),
    .Ci(Tile_X8Y12_Co),
    .E1END(Tile_X7Y11_E1BEG),
    .E2MID(Tile_X7Y11_E2BEG),
    .E2END(Tile_X7Y11_E2BEGb),
    .EE4END(Tile_X7Y11_EE4BEG),
    .E6END(Tile_X7Y11_E6BEG),
    .S1END(Tile_X8Y10_S1BEG),
    .S2MID(Tile_X8Y10_S2BEG),
    .S2END(Tile_X8Y10_S2BEGb),
    .S4END(Tile_X8Y10_S4BEG),
    .SS4END(Tile_X8Y10_SS4BEG),
    .W1END(Tile_X9Y11_W1BEG),
    .W2MID(Tile_X9Y11_W2BEG),
    .W2END(Tile_X9Y11_W2BEGb),
    .WW4END(Tile_X9Y11_WW4BEG),
    .W6END(Tile_X9Y11_W6BEG),
    .N1BEG(Tile_X8Y11_N1BEG),
    .N2BEG(Tile_X8Y11_N2BEG),
    .N2BEGb(Tile_X8Y11_N2BEGb),
    .N4BEG(Tile_X8Y11_N4BEG),
    .NN4BEG(Tile_X8Y11_NN4BEG),
    .E1BEG(Tile_X8Y11_E1BEG),
    .E2BEG(Tile_X8Y11_E2BEG),
    .E2BEGb(Tile_X8Y11_E2BEGb),
    .EE4BEG(Tile_X8Y11_EE4BEG),
    .E6BEG(Tile_X8Y11_E6BEG),
    .S1BEG(Tile_X8Y11_S1BEG),
    .S2BEG(Tile_X8Y11_S2BEG),
    .S2BEGb(Tile_X8Y11_S2BEGb),
    .S4BEG(Tile_X8Y11_S4BEG),
    .SS4BEG(Tile_X8Y11_SS4BEG),
    .W1BEG(Tile_X8Y11_W1BEG),
    .W2BEG(Tile_X8Y11_W2BEG),
    .W2BEGb(Tile_X8Y11_W2BEGb),
    .WW4BEG(Tile_X8Y11_WW4BEG),
    .W6BEG(Tile_X8Y11_W6BEG),
    .Co(Tile_X8Y11_Co),
    .UserCLK(Tile_X8Y12_UserCLKo),
    .UserCLKo(Tile_X8Y11_UserCLKo),
    .FrameData(Tile_X7Y11_FrameData_O),
    .FrameData_O(Tile_X8Y11_FrameData_O),
    .FrameStrobe(Tile_X8Y12_FrameStrobe_O),
    .FrameStrobe_O(Tile_X8Y11_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X9Y11_Emulate_Bitstream)
    )
`endif
    Tile_X9Y11_LUT4AB
    (
    .N1END(Tile_X9Y12_N1BEG),
    .N2MID(Tile_X9Y12_N2BEG),
    .N2END(Tile_X9Y12_N2BEGb),
    .N4END(Tile_X9Y12_N4BEG),
    .NN4END(Tile_X9Y12_NN4BEG),
    .Ci(Tile_X9Y12_Co),
    .E1END(Tile_X8Y11_E1BEG),
    .E2MID(Tile_X8Y11_E2BEG),
    .E2END(Tile_X8Y11_E2BEGb),
    .EE4END(Tile_X8Y11_EE4BEG),
    .E6END(Tile_X8Y11_E6BEG),
    .S1END(Tile_X9Y10_S1BEG),
    .S2MID(Tile_X9Y10_S2BEG),
    .S2END(Tile_X9Y10_S2BEGb),
    .S4END(Tile_X9Y10_S4BEG),
    .SS4END(Tile_X9Y10_SS4BEG),
    .W1END(Tile_X10Y11_W1BEG),
    .W2MID(Tile_X10Y11_W2BEG),
    .W2END(Tile_X10Y11_W2BEGb),
    .WW4END(Tile_X10Y11_WW4BEG),
    .W6END(Tile_X10Y11_W6BEG),
    .N1BEG(Tile_X9Y11_N1BEG),
    .N2BEG(Tile_X9Y11_N2BEG),
    .N2BEGb(Tile_X9Y11_N2BEGb),
    .N4BEG(Tile_X9Y11_N4BEG),
    .NN4BEG(Tile_X9Y11_NN4BEG),
    .E1BEG(Tile_X9Y11_E1BEG),
    .E2BEG(Tile_X9Y11_E2BEG),
    .E2BEGb(Tile_X9Y11_E2BEGb),
    .EE4BEG(Tile_X9Y11_EE4BEG),
    .E6BEG(Tile_X9Y11_E6BEG),
    .S1BEG(Tile_X9Y11_S1BEG),
    .S2BEG(Tile_X9Y11_S2BEG),
    .S2BEGb(Tile_X9Y11_S2BEGb),
    .S4BEG(Tile_X9Y11_S4BEG),
    .SS4BEG(Tile_X9Y11_SS4BEG),
    .W1BEG(Tile_X9Y11_W1BEG),
    .W2BEG(Tile_X9Y11_W2BEG),
    .W2BEGb(Tile_X9Y11_W2BEGb),
    .WW4BEG(Tile_X9Y11_WW4BEG),
    .W6BEG(Tile_X9Y11_W6BEG),
    .Co(Tile_X9Y11_Co),
    .UserCLK(Tile_X9Y12_UserCLKo),
    .UserCLKo(Tile_X9Y11_UserCLKo),
    .FrameData(Tile_X8Y11_FrameData_O),
    .FrameData_O(Tile_X9Y11_FrameData_O),
    .FrameStrobe(Tile_X9Y12_FrameStrobe_O),
    .FrameStrobe_O(Tile_X9Y11_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
IHP_SRAM
`ifdef EMULATION
    #(
    .Tile_X0Y0_Emulate_Bitstream(`Tile_X10Y11_Emulate_Bitstream),
    .Tile_X0Y1_Emulate_Bitstream(`Tile_X10Y12_Emulate_Bitstream)
    )
`endif
    Tile_X10Y11_IHP_SRAM
    (
    .Tile_X0Y0_E1END(Tile_X9Y11_E1BEG),
    .Tile_X0Y0_E2MID(Tile_X9Y11_E2BEG),
    .Tile_X0Y0_E2END(Tile_X9Y11_E2BEGb),
    .Tile_X0Y0_EE4END(Tile_X9Y11_EE4BEG),
    .Tile_X0Y0_E6END(Tile_X9Y11_E6BEG),
    .Tile_X0Y0_S1END(Tile_X10Y10_S1BEG),
    .Tile_X0Y0_S2MID(Tile_X10Y10_S2BEG),
    .Tile_X0Y0_S2END(Tile_X10Y10_S2BEGb),
    .Tile_X0Y0_S4END(Tile_X10Y10_S4BEG),
    .Tile_X0Y1_N1END(Tile_X10Y13_N1BEG),
    .Tile_X0Y1_N2MID(Tile_X10Y13_N2BEG),
    .Tile_X0Y1_N2END(Tile_X10Y13_N2BEGb),
    .Tile_X0Y1_N4END(Tile_X10Y13_N4BEG),
    .Tile_X0Y1_E1END(Tile_X9Y12_E1BEG),
    .Tile_X0Y1_E2MID(Tile_X9Y12_E2BEG),
    .Tile_X0Y1_E2END(Tile_X9Y12_E2BEGb),
    .Tile_X0Y1_EE4END(Tile_X9Y12_EE4BEG),
    .Tile_X0Y1_E6END(Tile_X9Y12_E6BEG),
    .Tile_X0Y0_N1BEG(Tile_X10Y11_N1BEG),
    .Tile_X0Y0_N2BEG(Tile_X10Y11_N2BEG),
    .Tile_X0Y0_N2BEGb(Tile_X10Y11_N2BEGb),
    .Tile_X0Y0_N4BEG(Tile_X10Y11_N4BEG),
    .Tile_X0Y0_W1BEG(Tile_X10Y11_W1BEG),
    .Tile_X0Y0_W2BEG(Tile_X10Y11_W2BEG),
    .Tile_X0Y0_W2BEGb(Tile_X10Y11_W2BEGb),
    .Tile_X0Y0_WW4BEG(Tile_X10Y11_WW4BEG),
    .Tile_X0Y0_W6BEG(Tile_X10Y11_W6BEG),
    .Tile_X0Y1_S1BEG(Tile_X10Y12_S1BEG),
    .Tile_X0Y1_S2BEG(Tile_X10Y12_S2BEG),
    .Tile_X0Y1_S2BEGb(Tile_X10Y12_S2BEGb),
    .Tile_X0Y1_S4BEG(Tile_X10Y12_S4BEG),
    .Tile_X0Y1_W1BEG(Tile_X10Y12_W1BEG),
    .Tile_X0Y1_W2BEG(Tile_X10Y12_W2BEG),
    .Tile_X0Y1_W2BEGb(Tile_X10Y12_W2BEGb),
    .Tile_X0Y1_WW4BEG(Tile_X10Y12_WW4BEG),
    .Tile_X0Y1_W6BEG(Tile_X10Y12_W6BEG),
    .CONFIGURED_top(Tile_X10Y12_CONFIGURED_top),
    .DOUT_SRAM0(Tile_X10Y12_DOUT_SRAM0),
    .DOUT_SRAM1(Tile_X10Y12_DOUT_SRAM1),
    .DOUT_SRAM2(Tile_X10Y12_DOUT_SRAM2),
    .DOUT_SRAM3(Tile_X10Y12_DOUT_SRAM3),
    .DOUT_SRAM4(Tile_X10Y12_DOUT_SRAM4),
    .DOUT_SRAM5(Tile_X10Y12_DOUT_SRAM5),
    .DOUT_SRAM6(Tile_X10Y12_DOUT_SRAM6),
    .DOUT_SRAM7(Tile_X10Y12_DOUT_SRAM7),
    .DOUT_SRAM8(Tile_X10Y12_DOUT_SRAM8),
    .DOUT_SRAM9(Tile_X10Y12_DOUT_SRAM9),
    .DOUT_SRAM10(Tile_X10Y12_DOUT_SRAM10),
    .DOUT_SRAM11(Tile_X10Y12_DOUT_SRAM11),
    .DOUT_SRAM12(Tile_X10Y12_DOUT_SRAM12),
    .DOUT_SRAM13(Tile_X10Y12_DOUT_SRAM13),
    .DOUT_SRAM14(Tile_X10Y12_DOUT_SRAM14),
    .DOUT_SRAM15(Tile_X10Y12_DOUT_SRAM15),
    .DOUT_SRAM16(Tile_X10Y12_DOUT_SRAM16),
    .DOUT_SRAM17(Tile_X10Y12_DOUT_SRAM17),
    .DOUT_SRAM18(Tile_X10Y12_DOUT_SRAM18),
    .DOUT_SRAM19(Tile_X10Y12_DOUT_SRAM19),
    .DOUT_SRAM20(Tile_X10Y12_DOUT_SRAM20),
    .DOUT_SRAM21(Tile_X10Y12_DOUT_SRAM21),
    .DOUT_SRAM22(Tile_X10Y12_DOUT_SRAM22),
    .DOUT_SRAM23(Tile_X10Y12_DOUT_SRAM23),
    .DOUT_SRAM24(Tile_X10Y12_DOUT_SRAM24),
    .DOUT_SRAM25(Tile_X10Y12_DOUT_SRAM25),
    .DOUT_SRAM26(Tile_X10Y12_DOUT_SRAM26),
    .DOUT_SRAM27(Tile_X10Y12_DOUT_SRAM27),
    .DOUT_SRAM28(Tile_X10Y12_DOUT_SRAM28),
    .DOUT_SRAM29(Tile_X10Y12_DOUT_SRAM29),
    .DOUT_SRAM30(Tile_X10Y12_DOUT_SRAM30),
    .DOUT_SRAM31(Tile_X10Y12_DOUT_SRAM31),
    .ADDR_SRAM0(Tile_X10Y12_ADDR_SRAM0),
    .ADDR_SRAM1(Tile_X10Y12_ADDR_SRAM1),
    .ADDR_SRAM2(Tile_X10Y12_ADDR_SRAM2),
    .ADDR_SRAM3(Tile_X10Y12_ADDR_SRAM3),
    .ADDR_SRAM4(Tile_X10Y12_ADDR_SRAM4),
    .ADDR_SRAM5(Tile_X10Y12_ADDR_SRAM5),
    .ADDR_SRAM6(Tile_X10Y12_ADDR_SRAM6),
    .ADDR_SRAM7(Tile_X10Y12_ADDR_SRAM7),
    .ADDR_SRAM8(Tile_X10Y12_ADDR_SRAM8),
    .ADDR_SRAM9(Tile_X10Y12_ADDR_SRAM9),
    .BM_SRAM0(Tile_X10Y12_BM_SRAM0),
    .BM_SRAM1(Tile_X10Y12_BM_SRAM1),
    .BM_SRAM2(Tile_X10Y12_BM_SRAM2),
    .BM_SRAM3(Tile_X10Y12_BM_SRAM3),
    .BM_SRAM4(Tile_X10Y12_BM_SRAM4),
    .BM_SRAM5(Tile_X10Y12_BM_SRAM5),
    .BM_SRAM6(Tile_X10Y12_BM_SRAM6),
    .BM_SRAM7(Tile_X10Y12_BM_SRAM7),
    .BM_SRAM8(Tile_X10Y12_BM_SRAM8),
    .BM_SRAM9(Tile_X10Y12_BM_SRAM9),
    .BM_SRAM10(Tile_X10Y12_BM_SRAM10),
    .BM_SRAM11(Tile_X10Y12_BM_SRAM11),
    .BM_SRAM12(Tile_X10Y12_BM_SRAM12),
    .BM_SRAM13(Tile_X10Y12_BM_SRAM13),
    .BM_SRAM14(Tile_X10Y12_BM_SRAM14),
    .BM_SRAM15(Tile_X10Y12_BM_SRAM15),
    .BM_SRAM16(Tile_X10Y12_BM_SRAM16),
    .BM_SRAM17(Tile_X10Y12_BM_SRAM17),
    .BM_SRAM18(Tile_X10Y12_BM_SRAM18),
    .BM_SRAM19(Tile_X10Y12_BM_SRAM19),
    .BM_SRAM20(Tile_X10Y12_BM_SRAM20),
    .BM_SRAM21(Tile_X10Y12_BM_SRAM21),
    .BM_SRAM22(Tile_X10Y12_BM_SRAM22),
    .BM_SRAM23(Tile_X10Y12_BM_SRAM23),
    .BM_SRAM24(Tile_X10Y12_BM_SRAM24),
    .BM_SRAM25(Tile_X10Y12_BM_SRAM25),
    .BM_SRAM26(Tile_X10Y12_BM_SRAM26),
    .BM_SRAM27(Tile_X10Y12_BM_SRAM27),
    .BM_SRAM28(Tile_X10Y12_BM_SRAM28),
    .BM_SRAM29(Tile_X10Y12_BM_SRAM29),
    .BM_SRAM30(Tile_X10Y12_BM_SRAM30),
    .BM_SRAM31(Tile_X10Y12_BM_SRAM31),
    .CLK_SRAM(Tile_X10Y12_CLK_SRAM),
    .DIN_SRAM0(Tile_X10Y12_DIN_SRAM0),
    .DIN_SRAM1(Tile_X10Y12_DIN_SRAM1),
    .DIN_SRAM2(Tile_X10Y12_DIN_SRAM2),
    .DIN_SRAM3(Tile_X10Y12_DIN_SRAM3),
    .DIN_SRAM4(Tile_X10Y12_DIN_SRAM4),
    .DIN_SRAM5(Tile_X10Y12_DIN_SRAM5),
    .DIN_SRAM6(Tile_X10Y12_DIN_SRAM6),
    .DIN_SRAM7(Tile_X10Y12_DIN_SRAM7),
    .DIN_SRAM8(Tile_X10Y12_DIN_SRAM8),
    .DIN_SRAM9(Tile_X10Y12_DIN_SRAM9),
    .DIN_SRAM10(Tile_X10Y12_DIN_SRAM10),
    .DIN_SRAM11(Tile_X10Y12_DIN_SRAM11),
    .DIN_SRAM12(Tile_X10Y12_DIN_SRAM12),
    .DIN_SRAM13(Tile_X10Y12_DIN_SRAM13),
    .DIN_SRAM14(Tile_X10Y12_DIN_SRAM14),
    .DIN_SRAM15(Tile_X10Y12_DIN_SRAM15),
    .DIN_SRAM16(Tile_X10Y12_DIN_SRAM16),
    .DIN_SRAM17(Tile_X10Y12_DIN_SRAM17),
    .DIN_SRAM18(Tile_X10Y12_DIN_SRAM18),
    .DIN_SRAM19(Tile_X10Y12_DIN_SRAM19),
    .DIN_SRAM20(Tile_X10Y12_DIN_SRAM20),
    .DIN_SRAM21(Tile_X10Y12_DIN_SRAM21),
    .DIN_SRAM22(Tile_X10Y12_DIN_SRAM22),
    .DIN_SRAM23(Tile_X10Y12_DIN_SRAM23),
    .DIN_SRAM24(Tile_X10Y12_DIN_SRAM24),
    .DIN_SRAM25(Tile_X10Y12_DIN_SRAM25),
    .DIN_SRAM26(Tile_X10Y12_DIN_SRAM26),
    .DIN_SRAM27(Tile_X10Y12_DIN_SRAM27),
    .DIN_SRAM28(Tile_X10Y12_DIN_SRAM28),
    .DIN_SRAM29(Tile_X10Y12_DIN_SRAM29),
    .DIN_SRAM30(Tile_X10Y12_DIN_SRAM30),
    .DIN_SRAM31(Tile_X10Y12_DIN_SRAM31),
    .MEN_SRAM(Tile_X10Y12_MEN_SRAM),
    .REN_SRAM(Tile_X10Y12_REN_SRAM),
    .TIE_HIGH_SRAM(Tile_X10Y12_TIE_HIGH_SRAM),
    .TIE_LOW_SRAM(Tile_X10Y12_TIE_LOW_SRAM),
    .WEN_SRAM(Tile_X10Y12_WEN_SRAM),
    .Tile_X0Y0_UserCLKo(Tile_X10Y11_UserCLKo),
    .Tile_X0Y1_UserCLK(Tile_X10Y13_UserCLKo),
    .Tile_X0Y0_FrameData(Tile_X9Y11_FrameData_O),
    .Tile_X0Y0_FrameData_O(Tile_X10Y11_FrameData_O),
    .Tile_X0Y0_FrameStrobe_O(Tile_X10Y11_FrameStrobe_O),
    .Tile_X0Y1_FrameData(Tile_X9Y12_FrameData_O),
    .Tile_X0Y1_FrameData_O(Tile_X10Y12_FrameData_O),
    .Tile_X0Y1_FrameStrobe(Tile_X10Y13_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
W_IO
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X0Y12_Emulate_Bitstream)
    )
`endif
    Tile_X0Y12_W_IO
    (
    .W1END(Tile_X1Y12_W1BEG),
    .W2MID(Tile_X1Y12_W2BEG),
    .W2END(Tile_X1Y12_W2BEGb),
    .WW4END(Tile_X1Y12_WW4BEG),
    .W6END(Tile_X1Y12_W6BEG),
    .E1BEG(Tile_X0Y12_E1BEG),
    .E2BEG(Tile_X0Y12_E2BEG),
    .E2BEGb(Tile_X0Y12_E2BEGb),
    .EE4BEG(Tile_X0Y12_EE4BEG),
    .E6BEG(Tile_X0Y12_E6BEG),
    .A_O_top(Tile_X0Y12_A_O_top),
    .A_I_top(Tile_X0Y12_A_I_top),
    .A_T_top(Tile_X0Y12_A_T_top),
    .B_O_top(Tile_X0Y12_B_O_top),
    .B_I_top(Tile_X0Y12_B_I_top),
    .B_T_top(Tile_X0Y12_B_T_top),
    .A_config_C_bit0(Tile_X0Y12_A_config_C_bit0),
    .A_config_C_bit1(Tile_X0Y12_A_config_C_bit1),
    .A_config_C_bit2(Tile_X0Y12_A_config_C_bit2),
    .A_config_C_bit3(Tile_X0Y12_A_config_C_bit3),
    .B_config_C_bit0(Tile_X0Y12_B_config_C_bit0),
    .B_config_C_bit1(Tile_X0Y12_B_config_C_bit1),
    .B_config_C_bit2(Tile_X0Y12_B_config_C_bit2),
    .B_config_C_bit3(Tile_X0Y12_B_config_C_bit3),
    .UserCLK(Tile_X0Y13_UserCLKo),
    .UserCLKo(Tile_X0Y12_UserCLKo),
    .FrameData(Row_Y12_FrameData),
    .FrameData_O(Tile_X0Y12_FrameData_O),
    .FrameStrobe(Tile_X0Y13_FrameStrobe_O),
    .FrameStrobe_O(Tile_X0Y12_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X1Y12_Emulate_Bitstream)
    )
`endif
    Tile_X1Y12_LUT4AB
    (
    .N1END(Tile_X1Y13_N1BEG),
    .N2MID(Tile_X1Y13_N2BEG),
    .N2END(Tile_X1Y13_N2BEGb),
    .N4END(Tile_X1Y13_N4BEG),
    .NN4END(Tile_X1Y13_NN4BEG),
    .Ci(Tile_X1Y13_Co),
    .E1END(Tile_X0Y12_E1BEG),
    .E2MID(Tile_X0Y12_E2BEG),
    .E2END(Tile_X0Y12_E2BEGb),
    .EE4END(Tile_X0Y12_EE4BEG),
    .E6END(Tile_X0Y12_E6BEG),
    .S1END(Tile_X1Y11_S1BEG),
    .S2MID(Tile_X1Y11_S2BEG),
    .S2END(Tile_X1Y11_S2BEGb),
    .S4END(Tile_X1Y11_S4BEG),
    .SS4END(Tile_X1Y11_SS4BEG),
    .W1END(Tile_X2Y12_W1BEG),
    .W2MID(Tile_X2Y12_W2BEG),
    .W2END(Tile_X2Y12_W2BEGb),
    .WW4END(Tile_X2Y12_WW4BEG),
    .W6END(Tile_X2Y12_W6BEG),
    .N1BEG(Tile_X1Y12_N1BEG),
    .N2BEG(Tile_X1Y12_N2BEG),
    .N2BEGb(Tile_X1Y12_N2BEGb),
    .N4BEG(Tile_X1Y12_N4BEG),
    .NN4BEG(Tile_X1Y12_NN4BEG),
    .E1BEG(Tile_X1Y12_E1BEG),
    .E2BEG(Tile_X1Y12_E2BEG),
    .E2BEGb(Tile_X1Y12_E2BEGb),
    .EE4BEG(Tile_X1Y12_EE4BEG),
    .E6BEG(Tile_X1Y12_E6BEG),
    .S1BEG(Tile_X1Y12_S1BEG),
    .S2BEG(Tile_X1Y12_S2BEG),
    .S2BEGb(Tile_X1Y12_S2BEGb),
    .S4BEG(Tile_X1Y12_S4BEG),
    .SS4BEG(Tile_X1Y12_SS4BEG),
    .W1BEG(Tile_X1Y12_W1BEG),
    .W2BEG(Tile_X1Y12_W2BEG),
    .W2BEGb(Tile_X1Y12_W2BEGb),
    .WW4BEG(Tile_X1Y12_WW4BEG),
    .W6BEG(Tile_X1Y12_W6BEG),
    .Co(Tile_X1Y12_Co),
    .UserCLK(Tile_X1Y13_UserCLKo),
    .UserCLKo(Tile_X1Y12_UserCLKo),
    .FrameData(Tile_X0Y12_FrameData_O),
    .FrameData_O(Tile_X1Y12_FrameData_O),
    .FrameStrobe(Tile_X1Y13_FrameStrobe_O),
    .FrameStrobe_O(Tile_X1Y12_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X2Y12_Emulate_Bitstream)
    )
`endif
    Tile_X2Y12_LUT4AB
    (
    .N1END(Tile_X2Y13_N1BEG),
    .N2MID(Tile_X2Y13_N2BEG),
    .N2END(Tile_X2Y13_N2BEGb),
    .N4END(Tile_X2Y13_N4BEG),
    .NN4END(Tile_X2Y13_NN4BEG),
    .Ci(Tile_X2Y13_Co),
    .E1END(Tile_X1Y12_E1BEG),
    .E2MID(Tile_X1Y12_E2BEG),
    .E2END(Tile_X1Y12_E2BEGb),
    .EE4END(Tile_X1Y12_EE4BEG),
    .E6END(Tile_X1Y12_E6BEG),
    .S1END(Tile_X2Y11_S1BEG),
    .S2MID(Tile_X2Y11_S2BEG),
    .S2END(Tile_X2Y11_S2BEGb),
    .S4END(Tile_X2Y11_S4BEG),
    .SS4END(Tile_X2Y11_SS4BEG),
    .W1END(Tile_X3Y12_W1BEG),
    .W2MID(Tile_X3Y12_W2BEG),
    .W2END(Tile_X3Y12_W2BEGb),
    .WW4END(Tile_X3Y12_WW4BEG),
    .W6END(Tile_X3Y12_W6BEG),
    .N1BEG(Tile_X2Y12_N1BEG),
    .N2BEG(Tile_X2Y12_N2BEG),
    .N2BEGb(Tile_X2Y12_N2BEGb),
    .N4BEG(Tile_X2Y12_N4BEG),
    .NN4BEG(Tile_X2Y12_NN4BEG),
    .E1BEG(Tile_X2Y12_E1BEG),
    .E2BEG(Tile_X2Y12_E2BEG),
    .E2BEGb(Tile_X2Y12_E2BEGb),
    .EE4BEG(Tile_X2Y12_EE4BEG),
    .E6BEG(Tile_X2Y12_E6BEG),
    .S1BEG(Tile_X2Y12_S1BEG),
    .S2BEG(Tile_X2Y12_S2BEG),
    .S2BEGb(Tile_X2Y12_S2BEGb),
    .S4BEG(Tile_X2Y12_S4BEG),
    .SS4BEG(Tile_X2Y12_SS4BEG),
    .W1BEG(Tile_X2Y12_W1BEG),
    .W2BEG(Tile_X2Y12_W2BEG),
    .W2BEGb(Tile_X2Y12_W2BEGb),
    .WW4BEG(Tile_X2Y12_WW4BEG),
    .W6BEG(Tile_X2Y12_W6BEG),
    .Co(Tile_X2Y12_Co),
    .UserCLK(Tile_X2Y13_UserCLKo),
    .UserCLKo(Tile_X2Y12_UserCLKo),
    .FrameData(Tile_X1Y12_FrameData_O),
    .FrameData_O(Tile_X2Y12_FrameData_O),
    .FrameStrobe(Tile_X2Y13_FrameStrobe_O),
    .FrameStrobe_O(Tile_X2Y12_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X3Y12_Emulate_Bitstream)
    )
`endif
    Tile_X3Y12_LUT4AB
    (
    .N1END(Tile_X3Y13_N1BEG),
    .N2MID(Tile_X3Y13_N2BEG),
    .N2END(Tile_X3Y13_N2BEGb),
    .N4END(Tile_X3Y13_N4BEG),
    .NN4END(Tile_X3Y13_NN4BEG),
    .Ci(Tile_X3Y13_Co),
    .E1END(Tile_X2Y12_E1BEG),
    .E2MID(Tile_X2Y12_E2BEG),
    .E2END(Tile_X2Y12_E2BEGb),
    .EE4END(Tile_X2Y12_EE4BEG),
    .E6END(Tile_X2Y12_E6BEG),
    .S1END(Tile_X3Y11_S1BEG),
    .S2MID(Tile_X3Y11_S2BEG),
    .S2END(Tile_X3Y11_S2BEGb),
    .S4END(Tile_X3Y11_S4BEG),
    .SS4END(Tile_X3Y11_SS4BEG),
    .W1END(Tile_X4Y12_W1BEG),
    .W2MID(Tile_X4Y12_W2BEG),
    .W2END(Tile_X4Y12_W2BEGb),
    .WW4END(Tile_X4Y12_WW4BEG),
    .W6END(Tile_X4Y12_W6BEG),
    .N1BEG(Tile_X3Y12_N1BEG),
    .N2BEG(Tile_X3Y12_N2BEG),
    .N2BEGb(Tile_X3Y12_N2BEGb),
    .N4BEG(Tile_X3Y12_N4BEG),
    .NN4BEG(Tile_X3Y12_NN4BEG),
    .E1BEG(Tile_X3Y12_E1BEG),
    .E2BEG(Tile_X3Y12_E2BEG),
    .E2BEGb(Tile_X3Y12_E2BEGb),
    .EE4BEG(Tile_X3Y12_EE4BEG),
    .E6BEG(Tile_X3Y12_E6BEG),
    .S1BEG(Tile_X3Y12_S1BEG),
    .S2BEG(Tile_X3Y12_S2BEG),
    .S2BEGb(Tile_X3Y12_S2BEGb),
    .S4BEG(Tile_X3Y12_S4BEG),
    .SS4BEG(Tile_X3Y12_SS4BEG),
    .W1BEG(Tile_X3Y12_W1BEG),
    .W2BEG(Tile_X3Y12_W2BEG),
    .W2BEGb(Tile_X3Y12_W2BEGb),
    .WW4BEG(Tile_X3Y12_WW4BEG),
    .W6BEG(Tile_X3Y12_W6BEG),
    .Co(Tile_X3Y12_Co),
    .UserCLK(Tile_X3Y13_UserCLKo),
    .UserCLKo(Tile_X3Y12_UserCLKo),
    .FrameData(Tile_X2Y12_FrameData_O),
    .FrameData_O(Tile_X3Y12_FrameData_O),
    .FrameStrobe(Tile_X3Y13_FrameStrobe_O),
    .FrameStrobe_O(Tile_X3Y12_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
RegFile
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X4Y12_Emulate_Bitstream)
    )
`endif
    Tile_X4Y12_RegFile
    (
    .N1END(Tile_X4Y13_N1BEG),
    .N2MID(Tile_X4Y13_N2BEG),
    .N2END(Tile_X4Y13_N2BEGb),
    .N4END(Tile_X4Y13_N4BEG),
    .NN4END(Tile_X4Y13_NN4BEG),
    .E1END(Tile_X3Y12_E1BEG),
    .E2MID(Tile_X3Y12_E2BEG),
    .E2END(Tile_X3Y12_E2BEGb),
    .EE4END(Tile_X3Y12_EE4BEG),
    .E6END(Tile_X3Y12_E6BEG),
    .S1END(Tile_X4Y11_S1BEG),
    .S2MID(Tile_X4Y11_S2BEG),
    .S2END(Tile_X4Y11_S2BEGb),
    .S4END(Tile_X4Y11_S4BEG),
    .SS4END(Tile_X4Y11_SS4BEG),
    .W1END(Tile_X5Y12_W1BEG),
    .W2MID(Tile_X5Y12_W2BEG),
    .W2END(Tile_X5Y12_W2BEGb),
    .WW4END(Tile_X5Y12_WW4BEG),
    .W6END(Tile_X5Y12_W6BEG),
    .N1BEG(Tile_X4Y12_N1BEG),
    .N2BEG(Tile_X4Y12_N2BEG),
    .N2BEGb(Tile_X4Y12_N2BEGb),
    .N4BEG(Tile_X4Y12_N4BEG),
    .NN4BEG(Tile_X4Y12_NN4BEG),
    .E1BEG(Tile_X4Y12_E1BEG),
    .E2BEG(Tile_X4Y12_E2BEG),
    .E2BEGb(Tile_X4Y12_E2BEGb),
    .EE4BEG(Tile_X4Y12_EE4BEG),
    .E6BEG(Tile_X4Y12_E6BEG),
    .S1BEG(Tile_X4Y12_S1BEG),
    .S2BEG(Tile_X4Y12_S2BEG),
    .S2BEGb(Tile_X4Y12_S2BEGb),
    .S4BEG(Tile_X4Y12_S4BEG),
    .SS4BEG(Tile_X4Y12_SS4BEG),
    .W1BEG(Tile_X4Y12_W1BEG),
    .W2BEG(Tile_X4Y12_W2BEG),
    .W2BEGb(Tile_X4Y12_W2BEGb),
    .WW4BEG(Tile_X4Y12_WW4BEG),
    .W6BEG(Tile_X4Y12_W6BEG),
    .UserCLK(Tile_X4Y13_UserCLKo),
    .UserCLKo(Tile_X4Y12_UserCLKo),
    .FrameData(Tile_X3Y12_FrameData_O),
    .FrameData_O(Tile_X4Y12_FrameData_O),
    .FrameStrobe(Tile_X4Y13_FrameStrobe_O),
    .FrameStrobe_O(Tile_X4Y12_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X5Y12_Emulate_Bitstream)
    )
`endif
    Tile_X5Y12_LUT4AB
    (
    .N1END(Tile_X5Y13_N1BEG),
    .N2MID(Tile_X5Y13_N2BEG),
    .N2END(Tile_X5Y13_N2BEGb),
    .N4END(Tile_X5Y13_N4BEG),
    .NN4END(Tile_X5Y13_NN4BEG),
    .Ci(Tile_X5Y13_Co),
    .E1END(Tile_X4Y12_E1BEG),
    .E2MID(Tile_X4Y12_E2BEG),
    .E2END(Tile_X4Y12_E2BEGb),
    .EE4END(Tile_X4Y12_EE4BEG),
    .E6END(Tile_X4Y12_E6BEG),
    .S1END(Tile_X5Y11_S1BEG),
    .S2MID(Tile_X5Y11_S2BEG),
    .S2END(Tile_X5Y11_S2BEGb),
    .S4END(Tile_X5Y11_S4BEG),
    .SS4END(Tile_X5Y11_SS4BEG),
    .W1END(Tile_X6Y12_W1BEG),
    .W2MID(Tile_X6Y12_W2BEG),
    .W2END(Tile_X6Y12_W2BEGb),
    .WW4END(Tile_X6Y12_WW4BEG),
    .W6END(Tile_X6Y12_W6BEG),
    .N1BEG(Tile_X5Y12_N1BEG),
    .N2BEG(Tile_X5Y12_N2BEG),
    .N2BEGb(Tile_X5Y12_N2BEGb),
    .N4BEG(Tile_X5Y12_N4BEG),
    .NN4BEG(Tile_X5Y12_NN4BEG),
    .E1BEG(Tile_X5Y12_E1BEG),
    .E2BEG(Tile_X5Y12_E2BEG),
    .E2BEGb(Tile_X5Y12_E2BEGb),
    .EE4BEG(Tile_X5Y12_EE4BEG),
    .E6BEG(Tile_X5Y12_E6BEG),
    .S1BEG(Tile_X5Y12_S1BEG),
    .S2BEG(Tile_X5Y12_S2BEG),
    .S2BEGb(Tile_X5Y12_S2BEGb),
    .S4BEG(Tile_X5Y12_S4BEG),
    .SS4BEG(Tile_X5Y12_SS4BEG),
    .W1BEG(Tile_X5Y12_W1BEG),
    .W2BEG(Tile_X5Y12_W2BEG),
    .W2BEGb(Tile_X5Y12_W2BEGb),
    .WW4BEG(Tile_X5Y12_WW4BEG),
    .W6BEG(Tile_X5Y12_W6BEG),
    .Co(Tile_X5Y12_Co),
    .UserCLK(Tile_X5Y13_UserCLKo),
    .UserCLKo(Tile_X5Y12_UserCLKo),
    .FrameData(Tile_X4Y12_FrameData_O),
    .FrameData_O(Tile_X5Y12_FrameData_O),
    .FrameStrobe(Tile_X5Y13_FrameStrobe_O),
    .FrameStrobe_O(Tile_X5Y12_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X6Y12_Emulate_Bitstream)
    )
`endif
    Tile_X6Y12_LUT4AB
    (
    .N1END(Tile_X6Y13_N1BEG),
    .N2MID(Tile_X6Y13_N2BEG),
    .N2END(Tile_X6Y13_N2BEGb),
    .N4END(Tile_X6Y13_N4BEG),
    .NN4END(Tile_X6Y13_NN4BEG),
    .Ci(Tile_X6Y13_Co),
    .E1END(Tile_X5Y12_E1BEG),
    .E2MID(Tile_X5Y12_E2BEG),
    .E2END(Tile_X5Y12_E2BEGb),
    .EE4END(Tile_X5Y12_EE4BEG),
    .E6END(Tile_X5Y12_E6BEG),
    .S1END(Tile_X6Y11_S1BEG),
    .S2MID(Tile_X6Y11_S2BEG),
    .S2END(Tile_X6Y11_S2BEGb),
    .S4END(Tile_X6Y11_S4BEG),
    .SS4END(Tile_X6Y11_SS4BEG),
    .W1END(Tile_X7Y12_W1BEG),
    .W2MID(Tile_X7Y12_W2BEG),
    .W2END(Tile_X7Y12_W2BEGb),
    .WW4END(Tile_X7Y12_WW4BEG),
    .W6END(Tile_X7Y12_W6BEG),
    .N1BEG(Tile_X6Y12_N1BEG),
    .N2BEG(Tile_X6Y12_N2BEG),
    .N2BEGb(Tile_X6Y12_N2BEGb),
    .N4BEG(Tile_X6Y12_N4BEG),
    .NN4BEG(Tile_X6Y12_NN4BEG),
    .E1BEG(Tile_X6Y12_E1BEG),
    .E2BEG(Tile_X6Y12_E2BEG),
    .E2BEGb(Tile_X6Y12_E2BEGb),
    .EE4BEG(Tile_X6Y12_EE4BEG),
    .E6BEG(Tile_X6Y12_E6BEG),
    .S1BEG(Tile_X6Y12_S1BEG),
    .S2BEG(Tile_X6Y12_S2BEG),
    .S2BEGb(Tile_X6Y12_S2BEGb),
    .S4BEG(Tile_X6Y12_S4BEG),
    .SS4BEG(Tile_X6Y12_SS4BEG),
    .W1BEG(Tile_X6Y12_W1BEG),
    .W2BEG(Tile_X6Y12_W2BEG),
    .W2BEGb(Tile_X6Y12_W2BEGb),
    .WW4BEG(Tile_X6Y12_WW4BEG),
    .W6BEG(Tile_X6Y12_W6BEG),
    .Co(Tile_X6Y12_Co),
    .UserCLK(Tile_X6Y13_UserCLKo),
    .UserCLKo(Tile_X6Y12_UserCLKo),
    .FrameData(Tile_X5Y12_FrameData_O),
    .FrameData_O(Tile_X6Y12_FrameData_O),
    .FrameStrobe(Tile_X6Y13_FrameStrobe_O),
    .FrameStrobe_O(Tile_X6Y12_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X8Y12_Emulate_Bitstream)
    )
`endif
    Tile_X8Y12_LUT4AB
    (
    .N1END(Tile_X8Y13_N1BEG),
    .N2MID(Tile_X8Y13_N2BEG),
    .N2END(Tile_X8Y13_N2BEGb),
    .N4END(Tile_X8Y13_N4BEG),
    .NN4END(Tile_X8Y13_NN4BEG),
    .Ci(Tile_X8Y13_Co),
    .E1END(Tile_X7Y12_E1BEG),
    .E2MID(Tile_X7Y12_E2BEG),
    .E2END(Tile_X7Y12_E2BEGb),
    .EE4END(Tile_X7Y12_EE4BEG),
    .E6END(Tile_X7Y12_E6BEG),
    .S1END(Tile_X8Y11_S1BEG),
    .S2MID(Tile_X8Y11_S2BEG),
    .S2END(Tile_X8Y11_S2BEGb),
    .S4END(Tile_X8Y11_S4BEG),
    .SS4END(Tile_X8Y11_SS4BEG),
    .W1END(Tile_X9Y12_W1BEG),
    .W2MID(Tile_X9Y12_W2BEG),
    .W2END(Tile_X9Y12_W2BEGb),
    .WW4END(Tile_X9Y12_WW4BEG),
    .W6END(Tile_X9Y12_W6BEG),
    .N1BEG(Tile_X8Y12_N1BEG),
    .N2BEG(Tile_X8Y12_N2BEG),
    .N2BEGb(Tile_X8Y12_N2BEGb),
    .N4BEG(Tile_X8Y12_N4BEG),
    .NN4BEG(Tile_X8Y12_NN4BEG),
    .E1BEG(Tile_X8Y12_E1BEG),
    .E2BEG(Tile_X8Y12_E2BEG),
    .E2BEGb(Tile_X8Y12_E2BEGb),
    .EE4BEG(Tile_X8Y12_EE4BEG),
    .E6BEG(Tile_X8Y12_E6BEG),
    .S1BEG(Tile_X8Y12_S1BEG),
    .S2BEG(Tile_X8Y12_S2BEG),
    .S2BEGb(Tile_X8Y12_S2BEGb),
    .S4BEG(Tile_X8Y12_S4BEG),
    .SS4BEG(Tile_X8Y12_SS4BEG),
    .W1BEG(Tile_X8Y12_W1BEG),
    .W2BEG(Tile_X8Y12_W2BEG),
    .W2BEGb(Tile_X8Y12_W2BEGb),
    .WW4BEG(Tile_X8Y12_WW4BEG),
    .W6BEG(Tile_X8Y12_W6BEG),
    .Co(Tile_X8Y12_Co),
    .UserCLK(Tile_X8Y13_UserCLKo),
    .UserCLKo(Tile_X8Y12_UserCLKo),
    .FrameData(Tile_X7Y12_FrameData_O),
    .FrameData_O(Tile_X8Y12_FrameData_O),
    .FrameStrobe(Tile_X8Y13_FrameStrobe_O),
    .FrameStrobe_O(Tile_X8Y12_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X9Y12_Emulate_Bitstream)
    )
`endif
    Tile_X9Y12_LUT4AB
    (
    .N1END(Tile_X9Y13_N1BEG),
    .N2MID(Tile_X9Y13_N2BEG),
    .N2END(Tile_X9Y13_N2BEGb),
    .N4END(Tile_X9Y13_N4BEG),
    .NN4END(Tile_X9Y13_NN4BEG),
    .Ci(Tile_X9Y13_Co),
    .E1END(Tile_X8Y12_E1BEG),
    .E2MID(Tile_X8Y12_E2BEG),
    .E2END(Tile_X8Y12_E2BEGb),
    .EE4END(Tile_X8Y12_EE4BEG),
    .E6END(Tile_X8Y12_E6BEG),
    .S1END(Tile_X9Y11_S1BEG),
    .S2MID(Tile_X9Y11_S2BEG),
    .S2END(Tile_X9Y11_S2BEGb),
    .S4END(Tile_X9Y11_S4BEG),
    .SS4END(Tile_X9Y11_SS4BEG),
    .W1END(Tile_X10Y12_W1BEG),
    .W2MID(Tile_X10Y12_W2BEG),
    .W2END(Tile_X10Y12_W2BEGb),
    .WW4END(Tile_X10Y12_WW4BEG),
    .W6END(Tile_X10Y12_W6BEG),
    .N1BEG(Tile_X9Y12_N1BEG),
    .N2BEG(Tile_X9Y12_N2BEG),
    .N2BEGb(Tile_X9Y12_N2BEGb),
    .N4BEG(Tile_X9Y12_N4BEG),
    .NN4BEG(Tile_X9Y12_NN4BEG),
    .E1BEG(Tile_X9Y12_E1BEG),
    .E2BEG(Tile_X9Y12_E2BEG),
    .E2BEGb(Tile_X9Y12_E2BEGb),
    .EE4BEG(Tile_X9Y12_EE4BEG),
    .E6BEG(Tile_X9Y12_E6BEG),
    .S1BEG(Tile_X9Y12_S1BEG),
    .S2BEG(Tile_X9Y12_S2BEG),
    .S2BEGb(Tile_X9Y12_S2BEGb),
    .S4BEG(Tile_X9Y12_S4BEG),
    .SS4BEG(Tile_X9Y12_SS4BEG),
    .W1BEG(Tile_X9Y12_W1BEG),
    .W2BEG(Tile_X9Y12_W2BEG),
    .W2BEGb(Tile_X9Y12_W2BEGb),
    .WW4BEG(Tile_X9Y12_WW4BEG),
    .W6BEG(Tile_X9Y12_W6BEG),
    .Co(Tile_X9Y12_Co),
    .UserCLK(Tile_X9Y13_UserCLKo),
    .UserCLKo(Tile_X9Y12_UserCLKo),
    .FrameData(Tile_X8Y12_FrameData_O),
    .FrameData_O(Tile_X9Y12_FrameData_O),
    .FrameStrobe(Tile_X9Y13_FrameStrobe_O),
    .FrameStrobe_O(Tile_X9Y12_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
W_IO
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X0Y13_Emulate_Bitstream)
    )
`endif
    Tile_X0Y13_W_IO
    (
    .W1END(Tile_X1Y13_W1BEG),
    .W2MID(Tile_X1Y13_W2BEG),
    .W2END(Tile_X1Y13_W2BEGb),
    .WW4END(Tile_X1Y13_WW4BEG),
    .W6END(Tile_X1Y13_W6BEG),
    .E1BEG(Tile_X0Y13_E1BEG),
    .E2BEG(Tile_X0Y13_E2BEG),
    .E2BEGb(Tile_X0Y13_E2BEGb),
    .EE4BEG(Tile_X0Y13_EE4BEG),
    .E6BEG(Tile_X0Y13_E6BEG),
    .A_O_top(Tile_X0Y13_A_O_top),
    .A_I_top(Tile_X0Y13_A_I_top),
    .A_T_top(Tile_X0Y13_A_T_top),
    .B_O_top(Tile_X0Y13_B_O_top),
    .B_I_top(Tile_X0Y13_B_I_top),
    .B_T_top(Tile_X0Y13_B_T_top),
    .A_config_C_bit0(Tile_X0Y13_A_config_C_bit0),
    .A_config_C_bit1(Tile_X0Y13_A_config_C_bit1),
    .A_config_C_bit2(Tile_X0Y13_A_config_C_bit2),
    .A_config_C_bit3(Tile_X0Y13_A_config_C_bit3),
    .B_config_C_bit0(Tile_X0Y13_B_config_C_bit0),
    .B_config_C_bit1(Tile_X0Y13_B_config_C_bit1),
    .B_config_C_bit2(Tile_X0Y13_B_config_C_bit2),
    .B_config_C_bit3(Tile_X0Y13_B_config_C_bit3),
    .UserCLK(Tile_X0Y14_UserCLKo),
    .UserCLKo(Tile_X0Y13_UserCLKo),
    .FrameData(Row_Y13_FrameData),
    .FrameData_O(Tile_X0Y13_FrameData_O),
    .FrameStrobe(Tile_X0Y14_FrameStrobe_O),
    .FrameStrobe_O(Tile_X0Y13_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X1Y13_Emulate_Bitstream)
    )
`endif
    Tile_X1Y13_LUT4AB
    (
    .N1END(Tile_X1Y14_N1BEG),
    .N2MID(Tile_X1Y14_N2BEG),
    .N2END(Tile_X1Y14_N2BEGb),
    .N4END(Tile_X1Y14_N4BEG),
    .NN4END(Tile_X1Y14_NN4BEG),
    .Ci(Tile_X1Y14_Co),
    .E1END(Tile_X0Y13_E1BEG),
    .E2MID(Tile_X0Y13_E2BEG),
    .E2END(Tile_X0Y13_E2BEGb),
    .EE4END(Tile_X0Y13_EE4BEG),
    .E6END(Tile_X0Y13_E6BEG),
    .S1END(Tile_X1Y12_S1BEG),
    .S2MID(Tile_X1Y12_S2BEG),
    .S2END(Tile_X1Y12_S2BEGb),
    .S4END(Tile_X1Y12_S4BEG),
    .SS4END(Tile_X1Y12_SS4BEG),
    .W1END(Tile_X2Y13_W1BEG),
    .W2MID(Tile_X2Y13_W2BEG),
    .W2END(Tile_X2Y13_W2BEGb),
    .WW4END(Tile_X2Y13_WW4BEG),
    .W6END(Tile_X2Y13_W6BEG),
    .N1BEG(Tile_X1Y13_N1BEG),
    .N2BEG(Tile_X1Y13_N2BEG),
    .N2BEGb(Tile_X1Y13_N2BEGb),
    .N4BEG(Tile_X1Y13_N4BEG),
    .NN4BEG(Tile_X1Y13_NN4BEG),
    .E1BEG(Tile_X1Y13_E1BEG),
    .E2BEG(Tile_X1Y13_E2BEG),
    .E2BEGb(Tile_X1Y13_E2BEGb),
    .EE4BEG(Tile_X1Y13_EE4BEG),
    .E6BEG(Tile_X1Y13_E6BEG),
    .S1BEG(Tile_X1Y13_S1BEG),
    .S2BEG(Tile_X1Y13_S2BEG),
    .S2BEGb(Tile_X1Y13_S2BEGb),
    .S4BEG(Tile_X1Y13_S4BEG),
    .SS4BEG(Tile_X1Y13_SS4BEG),
    .W1BEG(Tile_X1Y13_W1BEG),
    .W2BEG(Tile_X1Y13_W2BEG),
    .W2BEGb(Tile_X1Y13_W2BEGb),
    .WW4BEG(Tile_X1Y13_WW4BEG),
    .W6BEG(Tile_X1Y13_W6BEG),
    .Co(Tile_X1Y13_Co),
    .UserCLK(Tile_X1Y14_UserCLKo),
    .UserCLKo(Tile_X1Y13_UserCLKo),
    .FrameData(Tile_X0Y13_FrameData_O),
    .FrameData_O(Tile_X1Y13_FrameData_O),
    .FrameStrobe(Tile_X1Y14_FrameStrobe_O),
    .FrameStrobe_O(Tile_X1Y13_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X2Y13_Emulate_Bitstream)
    )
`endif
    Tile_X2Y13_LUT4AB
    (
    .N1END(Tile_X2Y14_N1BEG),
    .N2MID(Tile_X2Y14_N2BEG),
    .N2END(Tile_X2Y14_N2BEGb),
    .N4END(Tile_X2Y14_N4BEG),
    .NN4END(Tile_X2Y14_NN4BEG),
    .Ci(Tile_X2Y14_Co),
    .E1END(Tile_X1Y13_E1BEG),
    .E2MID(Tile_X1Y13_E2BEG),
    .E2END(Tile_X1Y13_E2BEGb),
    .EE4END(Tile_X1Y13_EE4BEG),
    .E6END(Tile_X1Y13_E6BEG),
    .S1END(Tile_X2Y12_S1BEG),
    .S2MID(Tile_X2Y12_S2BEG),
    .S2END(Tile_X2Y12_S2BEGb),
    .S4END(Tile_X2Y12_S4BEG),
    .SS4END(Tile_X2Y12_SS4BEG),
    .W1END(Tile_X3Y13_W1BEG),
    .W2MID(Tile_X3Y13_W2BEG),
    .W2END(Tile_X3Y13_W2BEGb),
    .WW4END(Tile_X3Y13_WW4BEG),
    .W6END(Tile_X3Y13_W6BEG),
    .N1BEG(Tile_X2Y13_N1BEG),
    .N2BEG(Tile_X2Y13_N2BEG),
    .N2BEGb(Tile_X2Y13_N2BEGb),
    .N4BEG(Tile_X2Y13_N4BEG),
    .NN4BEG(Tile_X2Y13_NN4BEG),
    .E1BEG(Tile_X2Y13_E1BEG),
    .E2BEG(Tile_X2Y13_E2BEG),
    .E2BEGb(Tile_X2Y13_E2BEGb),
    .EE4BEG(Tile_X2Y13_EE4BEG),
    .E6BEG(Tile_X2Y13_E6BEG),
    .S1BEG(Tile_X2Y13_S1BEG),
    .S2BEG(Tile_X2Y13_S2BEG),
    .S2BEGb(Tile_X2Y13_S2BEGb),
    .S4BEG(Tile_X2Y13_S4BEG),
    .SS4BEG(Tile_X2Y13_SS4BEG),
    .W1BEG(Tile_X2Y13_W1BEG),
    .W2BEG(Tile_X2Y13_W2BEG),
    .W2BEGb(Tile_X2Y13_W2BEGb),
    .WW4BEG(Tile_X2Y13_WW4BEG),
    .W6BEG(Tile_X2Y13_W6BEG),
    .Co(Tile_X2Y13_Co),
    .UserCLK(Tile_X2Y14_UserCLKo),
    .UserCLKo(Tile_X2Y13_UserCLKo),
    .FrameData(Tile_X1Y13_FrameData_O),
    .FrameData_O(Tile_X2Y13_FrameData_O),
    .FrameStrobe(Tile_X2Y14_FrameStrobe_O),
    .FrameStrobe_O(Tile_X2Y13_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X3Y13_Emulate_Bitstream)
    )
`endif
    Tile_X3Y13_LUT4AB
    (
    .N1END(Tile_X3Y14_N1BEG),
    .N2MID(Tile_X3Y14_N2BEG),
    .N2END(Tile_X3Y14_N2BEGb),
    .N4END(Tile_X3Y14_N4BEG),
    .NN4END(Tile_X3Y14_NN4BEG),
    .Ci(Tile_X3Y14_Co),
    .E1END(Tile_X2Y13_E1BEG),
    .E2MID(Tile_X2Y13_E2BEG),
    .E2END(Tile_X2Y13_E2BEGb),
    .EE4END(Tile_X2Y13_EE4BEG),
    .E6END(Tile_X2Y13_E6BEG),
    .S1END(Tile_X3Y12_S1BEG),
    .S2MID(Tile_X3Y12_S2BEG),
    .S2END(Tile_X3Y12_S2BEGb),
    .S4END(Tile_X3Y12_S4BEG),
    .SS4END(Tile_X3Y12_SS4BEG),
    .W1END(Tile_X4Y13_W1BEG),
    .W2MID(Tile_X4Y13_W2BEG),
    .W2END(Tile_X4Y13_W2BEGb),
    .WW4END(Tile_X4Y13_WW4BEG),
    .W6END(Tile_X4Y13_W6BEG),
    .N1BEG(Tile_X3Y13_N1BEG),
    .N2BEG(Tile_X3Y13_N2BEG),
    .N2BEGb(Tile_X3Y13_N2BEGb),
    .N4BEG(Tile_X3Y13_N4BEG),
    .NN4BEG(Tile_X3Y13_NN4BEG),
    .E1BEG(Tile_X3Y13_E1BEG),
    .E2BEG(Tile_X3Y13_E2BEG),
    .E2BEGb(Tile_X3Y13_E2BEGb),
    .EE4BEG(Tile_X3Y13_EE4BEG),
    .E6BEG(Tile_X3Y13_E6BEG),
    .S1BEG(Tile_X3Y13_S1BEG),
    .S2BEG(Tile_X3Y13_S2BEG),
    .S2BEGb(Tile_X3Y13_S2BEGb),
    .S4BEG(Tile_X3Y13_S4BEG),
    .SS4BEG(Tile_X3Y13_SS4BEG),
    .W1BEG(Tile_X3Y13_W1BEG),
    .W2BEG(Tile_X3Y13_W2BEG),
    .W2BEGb(Tile_X3Y13_W2BEGb),
    .WW4BEG(Tile_X3Y13_WW4BEG),
    .W6BEG(Tile_X3Y13_W6BEG),
    .Co(Tile_X3Y13_Co),
    .UserCLK(Tile_X3Y14_UserCLKo),
    .UserCLKo(Tile_X3Y13_UserCLKo),
    .FrameData(Tile_X2Y13_FrameData_O),
    .FrameData_O(Tile_X3Y13_FrameData_O),
    .FrameStrobe(Tile_X3Y14_FrameStrobe_O),
    .FrameStrobe_O(Tile_X3Y13_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
RegFile
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X4Y13_Emulate_Bitstream)
    )
`endif
    Tile_X4Y13_RegFile
    (
    .N1END(Tile_X4Y14_N1BEG),
    .N2MID(Tile_X4Y14_N2BEG),
    .N2END(Tile_X4Y14_N2BEGb),
    .N4END(Tile_X4Y14_N4BEG),
    .NN4END(Tile_X4Y14_NN4BEG),
    .E1END(Tile_X3Y13_E1BEG),
    .E2MID(Tile_X3Y13_E2BEG),
    .E2END(Tile_X3Y13_E2BEGb),
    .EE4END(Tile_X3Y13_EE4BEG),
    .E6END(Tile_X3Y13_E6BEG),
    .S1END(Tile_X4Y12_S1BEG),
    .S2MID(Tile_X4Y12_S2BEG),
    .S2END(Tile_X4Y12_S2BEGb),
    .S4END(Tile_X4Y12_S4BEG),
    .SS4END(Tile_X4Y12_SS4BEG),
    .W1END(Tile_X5Y13_W1BEG),
    .W2MID(Tile_X5Y13_W2BEG),
    .W2END(Tile_X5Y13_W2BEGb),
    .WW4END(Tile_X5Y13_WW4BEG),
    .W6END(Tile_X5Y13_W6BEG),
    .N1BEG(Tile_X4Y13_N1BEG),
    .N2BEG(Tile_X4Y13_N2BEG),
    .N2BEGb(Tile_X4Y13_N2BEGb),
    .N4BEG(Tile_X4Y13_N4BEG),
    .NN4BEG(Tile_X4Y13_NN4BEG),
    .E1BEG(Tile_X4Y13_E1BEG),
    .E2BEG(Tile_X4Y13_E2BEG),
    .E2BEGb(Tile_X4Y13_E2BEGb),
    .EE4BEG(Tile_X4Y13_EE4BEG),
    .E6BEG(Tile_X4Y13_E6BEG),
    .S1BEG(Tile_X4Y13_S1BEG),
    .S2BEG(Tile_X4Y13_S2BEG),
    .S2BEGb(Tile_X4Y13_S2BEGb),
    .S4BEG(Tile_X4Y13_S4BEG),
    .SS4BEG(Tile_X4Y13_SS4BEG),
    .W1BEG(Tile_X4Y13_W1BEG),
    .W2BEG(Tile_X4Y13_W2BEG),
    .W2BEGb(Tile_X4Y13_W2BEGb),
    .WW4BEG(Tile_X4Y13_WW4BEG),
    .W6BEG(Tile_X4Y13_W6BEG),
    .UserCLK(Tile_X4Y14_UserCLKo),
    .UserCLKo(Tile_X4Y13_UserCLKo),
    .FrameData(Tile_X3Y13_FrameData_O),
    .FrameData_O(Tile_X4Y13_FrameData_O),
    .FrameStrobe(Tile_X4Y14_FrameStrobe_O),
    .FrameStrobe_O(Tile_X4Y13_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X5Y13_Emulate_Bitstream)
    )
`endif
    Tile_X5Y13_LUT4AB
    (
    .N1END(Tile_X5Y14_N1BEG),
    .N2MID(Tile_X5Y14_N2BEG),
    .N2END(Tile_X5Y14_N2BEGb),
    .N4END(Tile_X5Y14_N4BEG),
    .NN4END(Tile_X5Y14_NN4BEG),
    .Ci(Tile_X5Y14_Co),
    .E1END(Tile_X4Y13_E1BEG),
    .E2MID(Tile_X4Y13_E2BEG),
    .E2END(Tile_X4Y13_E2BEGb),
    .EE4END(Tile_X4Y13_EE4BEG),
    .E6END(Tile_X4Y13_E6BEG),
    .S1END(Tile_X5Y12_S1BEG),
    .S2MID(Tile_X5Y12_S2BEG),
    .S2END(Tile_X5Y12_S2BEGb),
    .S4END(Tile_X5Y12_S4BEG),
    .SS4END(Tile_X5Y12_SS4BEG),
    .W1END(Tile_X6Y13_W1BEG),
    .W2MID(Tile_X6Y13_W2BEG),
    .W2END(Tile_X6Y13_W2BEGb),
    .WW4END(Tile_X6Y13_WW4BEG),
    .W6END(Tile_X6Y13_W6BEG),
    .N1BEG(Tile_X5Y13_N1BEG),
    .N2BEG(Tile_X5Y13_N2BEG),
    .N2BEGb(Tile_X5Y13_N2BEGb),
    .N4BEG(Tile_X5Y13_N4BEG),
    .NN4BEG(Tile_X5Y13_NN4BEG),
    .E1BEG(Tile_X5Y13_E1BEG),
    .E2BEG(Tile_X5Y13_E2BEG),
    .E2BEGb(Tile_X5Y13_E2BEGb),
    .EE4BEG(Tile_X5Y13_EE4BEG),
    .E6BEG(Tile_X5Y13_E6BEG),
    .S1BEG(Tile_X5Y13_S1BEG),
    .S2BEG(Tile_X5Y13_S2BEG),
    .S2BEGb(Tile_X5Y13_S2BEGb),
    .S4BEG(Tile_X5Y13_S4BEG),
    .SS4BEG(Tile_X5Y13_SS4BEG),
    .W1BEG(Tile_X5Y13_W1BEG),
    .W2BEG(Tile_X5Y13_W2BEG),
    .W2BEGb(Tile_X5Y13_W2BEGb),
    .WW4BEG(Tile_X5Y13_WW4BEG),
    .W6BEG(Tile_X5Y13_W6BEG),
    .Co(Tile_X5Y13_Co),
    .UserCLK(Tile_X5Y14_UserCLKo),
    .UserCLKo(Tile_X5Y13_UserCLKo),
    .FrameData(Tile_X4Y13_FrameData_O),
    .FrameData_O(Tile_X5Y13_FrameData_O),
    .FrameStrobe(Tile_X5Y14_FrameStrobe_O),
    .FrameStrobe_O(Tile_X5Y13_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X6Y13_Emulate_Bitstream)
    )
`endif
    Tile_X6Y13_LUT4AB
    (
    .N1END(Tile_X6Y14_N1BEG),
    .N2MID(Tile_X6Y14_N2BEG),
    .N2END(Tile_X6Y14_N2BEGb),
    .N4END(Tile_X6Y14_N4BEG),
    .NN4END(Tile_X6Y14_NN4BEG),
    .Ci(Tile_X6Y14_Co),
    .E1END(Tile_X5Y13_E1BEG),
    .E2MID(Tile_X5Y13_E2BEG),
    .E2END(Tile_X5Y13_E2BEGb),
    .EE4END(Tile_X5Y13_EE4BEG),
    .E6END(Tile_X5Y13_E6BEG),
    .S1END(Tile_X6Y12_S1BEG),
    .S2MID(Tile_X6Y12_S2BEG),
    .S2END(Tile_X6Y12_S2BEGb),
    .S4END(Tile_X6Y12_S4BEG),
    .SS4END(Tile_X6Y12_SS4BEG),
    .W1END(Tile_X7Y13_W1BEG),
    .W2MID(Tile_X7Y13_W2BEG),
    .W2END(Tile_X7Y13_W2BEGb),
    .WW4END(Tile_X7Y13_WW4BEG),
    .W6END(Tile_X7Y13_W6BEG),
    .N1BEG(Tile_X6Y13_N1BEG),
    .N2BEG(Tile_X6Y13_N2BEG),
    .N2BEGb(Tile_X6Y13_N2BEGb),
    .N4BEG(Tile_X6Y13_N4BEG),
    .NN4BEG(Tile_X6Y13_NN4BEG),
    .E1BEG(Tile_X6Y13_E1BEG),
    .E2BEG(Tile_X6Y13_E2BEG),
    .E2BEGb(Tile_X6Y13_E2BEGb),
    .EE4BEG(Tile_X6Y13_EE4BEG),
    .E6BEG(Tile_X6Y13_E6BEG),
    .S1BEG(Tile_X6Y13_S1BEG),
    .S2BEG(Tile_X6Y13_S2BEG),
    .S2BEGb(Tile_X6Y13_S2BEGb),
    .S4BEG(Tile_X6Y13_S4BEG),
    .SS4BEG(Tile_X6Y13_SS4BEG),
    .W1BEG(Tile_X6Y13_W1BEG),
    .W2BEG(Tile_X6Y13_W2BEG),
    .W2BEGb(Tile_X6Y13_W2BEGb),
    .WW4BEG(Tile_X6Y13_WW4BEG),
    .W6BEG(Tile_X6Y13_W6BEG),
    .Co(Tile_X6Y13_Co),
    .UserCLK(Tile_X6Y14_UserCLKo),
    .UserCLKo(Tile_X6Y13_UserCLKo),
    .FrameData(Tile_X5Y13_FrameData_O),
    .FrameData_O(Tile_X6Y13_FrameData_O),
    .FrameStrobe(Tile_X6Y14_FrameStrobe_O),
    .FrameStrobe_O(Tile_X6Y13_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
DSP
`ifdef EMULATION
    #(
    .Tile_X0Y0_Emulate_Bitstream(`Tile_X7Y13_Emulate_Bitstream),
    .Tile_X0Y1_Emulate_Bitstream(`Tile_X7Y14_Emulate_Bitstream)
    )
`endif
    Tile_X7Y13_DSP
    (
    .Tile_X0Y0_E1END(Tile_X6Y13_E1BEG),
    .Tile_X0Y0_E2MID(Tile_X6Y13_E2BEG),
    .Tile_X0Y0_E2END(Tile_X6Y13_E2BEGb),
    .Tile_X0Y0_EE4END(Tile_X6Y13_EE4BEG),
    .Tile_X0Y0_E6END(Tile_X6Y13_E6BEG),
    .Tile_X0Y0_S1END(Tile_X7Y12_S1BEG),
    .Tile_X0Y0_S2MID(Tile_X7Y12_S2BEG),
    .Tile_X0Y0_S2END(Tile_X7Y12_S2BEGb),
    .Tile_X0Y0_S4END(Tile_X7Y12_S4BEG),
    .Tile_X0Y0_SS4END(Tile_X7Y12_SS4BEG),
    .Tile_X0Y0_W1END(Tile_X8Y13_W1BEG),
    .Tile_X0Y0_W2MID(Tile_X8Y13_W2BEG),
    .Tile_X0Y0_W2END(Tile_X8Y13_W2BEGb),
    .Tile_X0Y0_WW4END(Tile_X8Y13_WW4BEG),
    .Tile_X0Y0_W6END(Tile_X8Y13_W6BEG),
    .Tile_X0Y1_N1END(Tile_X7Y15_N1BEG),
    .Tile_X0Y1_N2MID(Tile_X7Y15_N2BEG),
    .Tile_X0Y1_N2END(Tile_X7Y15_N2BEGb),
    .Tile_X0Y1_N4END(Tile_X7Y15_N4BEG),
    .Tile_X0Y1_NN4END(Tile_X7Y15_NN4BEG),
    .Tile_X0Y1_E1END(Tile_X6Y14_E1BEG),
    .Tile_X0Y1_E2MID(Tile_X6Y14_E2BEG),
    .Tile_X0Y1_E2END(Tile_X6Y14_E2BEGb),
    .Tile_X0Y1_EE4END(Tile_X6Y14_EE4BEG),
    .Tile_X0Y1_E6END(Tile_X6Y14_E6BEG),
    .Tile_X0Y1_W1END(Tile_X8Y14_W1BEG),
    .Tile_X0Y1_W2MID(Tile_X8Y14_W2BEG),
    .Tile_X0Y1_W2END(Tile_X8Y14_W2BEGb),
    .Tile_X0Y1_WW4END(Tile_X8Y14_WW4BEG),
    .Tile_X0Y1_W6END(Tile_X8Y14_W6BEG),
    .Tile_X0Y0_N1BEG(Tile_X7Y13_N1BEG),
    .Tile_X0Y0_N2BEG(Tile_X7Y13_N2BEG),
    .Tile_X0Y0_N2BEGb(Tile_X7Y13_N2BEGb),
    .Tile_X0Y0_N4BEG(Tile_X7Y13_N4BEG),
    .Tile_X0Y0_NN4BEG(Tile_X7Y13_NN4BEG),
    .Tile_X0Y0_E1BEG(Tile_X7Y13_E1BEG),
    .Tile_X0Y0_E2BEG(Tile_X7Y13_E2BEG),
    .Tile_X0Y0_E2BEGb(Tile_X7Y13_E2BEGb),
    .Tile_X0Y0_EE4BEG(Tile_X7Y13_EE4BEG),
    .Tile_X0Y0_E6BEG(Tile_X7Y13_E6BEG),
    .Tile_X0Y0_W1BEG(Tile_X7Y13_W1BEG),
    .Tile_X0Y0_W2BEG(Tile_X7Y13_W2BEG),
    .Tile_X0Y0_W2BEGb(Tile_X7Y13_W2BEGb),
    .Tile_X0Y0_WW4BEG(Tile_X7Y13_WW4BEG),
    .Tile_X0Y0_W6BEG(Tile_X7Y13_W6BEG),
    .Tile_X0Y1_E1BEG(Tile_X7Y14_E1BEG),
    .Tile_X0Y1_E2BEG(Tile_X7Y14_E2BEG),
    .Tile_X0Y1_E2BEGb(Tile_X7Y14_E2BEGb),
    .Tile_X0Y1_EE4BEG(Tile_X7Y14_EE4BEG),
    .Tile_X0Y1_E6BEG(Tile_X7Y14_E6BEG),
    .Tile_X0Y1_S1BEG(Tile_X7Y14_S1BEG),
    .Tile_X0Y1_S2BEG(Tile_X7Y14_S2BEG),
    .Tile_X0Y1_S2BEGb(Tile_X7Y14_S2BEGb),
    .Tile_X0Y1_S4BEG(Tile_X7Y14_S4BEG),
    .Tile_X0Y1_SS4BEG(Tile_X7Y14_SS4BEG),
    .Tile_X0Y1_W1BEG(Tile_X7Y14_W1BEG),
    .Tile_X0Y1_W2BEG(Tile_X7Y14_W2BEG),
    .Tile_X0Y1_W2BEGb(Tile_X7Y14_W2BEGb),
    .Tile_X0Y1_WW4BEG(Tile_X7Y14_WW4BEG),
    .Tile_X0Y1_W6BEG(Tile_X7Y14_W6BEG),
    .Tile_X0Y0_UserCLKo(Tile_X7Y13_UserCLKo),
    .Tile_X0Y1_UserCLK(Tile_X7Y15_UserCLKo),
    .Tile_X0Y0_FrameData(Tile_X6Y13_FrameData_O),
    .Tile_X0Y0_FrameData_O(Tile_X7Y13_FrameData_O),
    .Tile_X0Y0_FrameStrobe_O(Tile_X7Y13_FrameStrobe_O),
    .Tile_X0Y1_FrameData(Tile_X6Y14_FrameData_O),
    .Tile_X0Y1_FrameData_O(Tile_X7Y14_FrameData_O),
    .Tile_X0Y1_FrameStrobe(Tile_X7Y15_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X8Y13_Emulate_Bitstream)
    )
`endif
    Tile_X8Y13_LUT4AB
    (
    .N1END(Tile_X8Y14_N1BEG),
    .N2MID(Tile_X8Y14_N2BEG),
    .N2END(Tile_X8Y14_N2BEGb),
    .N4END(Tile_X8Y14_N4BEG),
    .NN4END(Tile_X8Y14_NN4BEG),
    .Ci(Tile_X8Y14_Co),
    .E1END(Tile_X7Y13_E1BEG),
    .E2MID(Tile_X7Y13_E2BEG),
    .E2END(Tile_X7Y13_E2BEGb),
    .EE4END(Tile_X7Y13_EE4BEG),
    .E6END(Tile_X7Y13_E6BEG),
    .S1END(Tile_X8Y12_S1BEG),
    .S2MID(Tile_X8Y12_S2BEG),
    .S2END(Tile_X8Y12_S2BEGb),
    .S4END(Tile_X8Y12_S4BEG),
    .SS4END(Tile_X8Y12_SS4BEG),
    .W1END(Tile_X9Y13_W1BEG),
    .W2MID(Tile_X9Y13_W2BEG),
    .W2END(Tile_X9Y13_W2BEGb),
    .WW4END(Tile_X9Y13_WW4BEG),
    .W6END(Tile_X9Y13_W6BEG),
    .N1BEG(Tile_X8Y13_N1BEG),
    .N2BEG(Tile_X8Y13_N2BEG),
    .N2BEGb(Tile_X8Y13_N2BEGb),
    .N4BEG(Tile_X8Y13_N4BEG),
    .NN4BEG(Tile_X8Y13_NN4BEG),
    .E1BEG(Tile_X8Y13_E1BEG),
    .E2BEG(Tile_X8Y13_E2BEG),
    .E2BEGb(Tile_X8Y13_E2BEGb),
    .EE4BEG(Tile_X8Y13_EE4BEG),
    .E6BEG(Tile_X8Y13_E6BEG),
    .S1BEG(Tile_X8Y13_S1BEG),
    .S2BEG(Tile_X8Y13_S2BEG),
    .S2BEGb(Tile_X8Y13_S2BEGb),
    .S4BEG(Tile_X8Y13_S4BEG),
    .SS4BEG(Tile_X8Y13_SS4BEG),
    .W1BEG(Tile_X8Y13_W1BEG),
    .W2BEG(Tile_X8Y13_W2BEG),
    .W2BEGb(Tile_X8Y13_W2BEGb),
    .WW4BEG(Tile_X8Y13_WW4BEG),
    .W6BEG(Tile_X8Y13_W6BEG),
    .Co(Tile_X8Y13_Co),
    .UserCLK(Tile_X8Y14_UserCLKo),
    .UserCLKo(Tile_X8Y13_UserCLKo),
    .FrameData(Tile_X7Y13_FrameData_O),
    .FrameData_O(Tile_X8Y13_FrameData_O),
    .FrameStrobe(Tile_X8Y14_FrameStrobe_O),
    .FrameStrobe_O(Tile_X8Y13_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X9Y13_Emulate_Bitstream)
    )
`endif
    Tile_X9Y13_LUT4AB
    (
    .N1END(Tile_X9Y14_N1BEG),
    .N2MID(Tile_X9Y14_N2BEG),
    .N2END(Tile_X9Y14_N2BEGb),
    .N4END(Tile_X9Y14_N4BEG),
    .NN4END(Tile_X9Y14_NN4BEG),
    .Ci(Tile_X9Y14_Co),
    .E1END(Tile_X8Y13_E1BEG),
    .E2MID(Tile_X8Y13_E2BEG),
    .E2END(Tile_X8Y13_E2BEGb),
    .EE4END(Tile_X8Y13_EE4BEG),
    .E6END(Tile_X8Y13_E6BEG),
    .S1END(Tile_X9Y12_S1BEG),
    .S2MID(Tile_X9Y12_S2BEG),
    .S2END(Tile_X9Y12_S2BEGb),
    .S4END(Tile_X9Y12_S4BEG),
    .SS4END(Tile_X9Y12_SS4BEG),
    .W1END(Tile_X10Y13_W1BEG),
    .W2MID(Tile_X10Y13_W2BEG),
    .W2END(Tile_X10Y13_W2BEGb),
    .WW4END(Tile_X10Y13_WW4BEG),
    .W6END(Tile_X10Y13_W6BEG),
    .N1BEG(Tile_X9Y13_N1BEG),
    .N2BEG(Tile_X9Y13_N2BEG),
    .N2BEGb(Tile_X9Y13_N2BEGb),
    .N4BEG(Tile_X9Y13_N4BEG),
    .NN4BEG(Tile_X9Y13_NN4BEG),
    .E1BEG(Tile_X9Y13_E1BEG),
    .E2BEG(Tile_X9Y13_E2BEG),
    .E2BEGb(Tile_X9Y13_E2BEGb),
    .EE4BEG(Tile_X9Y13_EE4BEG),
    .E6BEG(Tile_X9Y13_E6BEG),
    .S1BEG(Tile_X9Y13_S1BEG),
    .S2BEG(Tile_X9Y13_S2BEG),
    .S2BEGb(Tile_X9Y13_S2BEGb),
    .S4BEG(Tile_X9Y13_S4BEG),
    .SS4BEG(Tile_X9Y13_SS4BEG),
    .W1BEG(Tile_X9Y13_W1BEG),
    .W2BEG(Tile_X9Y13_W2BEG),
    .W2BEGb(Tile_X9Y13_W2BEGb),
    .WW4BEG(Tile_X9Y13_WW4BEG),
    .W6BEG(Tile_X9Y13_W6BEG),
    .Co(Tile_X9Y13_Co),
    .UserCLK(Tile_X9Y14_UserCLKo),
    .UserCLKo(Tile_X9Y13_UserCLKo),
    .FrameData(Tile_X8Y13_FrameData_O),
    .FrameData_O(Tile_X9Y13_FrameData_O),
    .FrameStrobe(Tile_X9Y14_FrameStrobe_O),
    .FrameStrobe_O(Tile_X9Y13_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
IHP_SRAM
`ifdef EMULATION
    #(
    .Tile_X0Y0_Emulate_Bitstream(`Tile_X10Y13_Emulate_Bitstream),
    .Tile_X0Y1_Emulate_Bitstream(`Tile_X10Y14_Emulate_Bitstream)
    )
`endif
    Tile_X10Y13_IHP_SRAM
    (
    .Tile_X0Y0_E1END(Tile_X9Y13_E1BEG),
    .Tile_X0Y0_E2MID(Tile_X9Y13_E2BEG),
    .Tile_X0Y0_E2END(Tile_X9Y13_E2BEGb),
    .Tile_X0Y0_EE4END(Tile_X9Y13_EE4BEG),
    .Tile_X0Y0_E6END(Tile_X9Y13_E6BEG),
    .Tile_X0Y0_S1END(Tile_X10Y12_S1BEG),
    .Tile_X0Y0_S2MID(Tile_X10Y12_S2BEG),
    .Tile_X0Y0_S2END(Tile_X10Y12_S2BEGb),
    .Tile_X0Y0_S4END(Tile_X10Y12_S4BEG),
    .Tile_X0Y1_N1END(Tile_X10Y15_N1BEG),
    .Tile_X0Y1_N2MID(Tile_X10Y15_N2BEG),
    .Tile_X0Y1_N2END(Tile_X10Y15_N2BEGb),
    .Tile_X0Y1_N4END(Tile_X10Y15_N4BEG),
    .Tile_X0Y1_E1END(Tile_X9Y14_E1BEG),
    .Tile_X0Y1_E2MID(Tile_X9Y14_E2BEG),
    .Tile_X0Y1_E2END(Tile_X9Y14_E2BEGb),
    .Tile_X0Y1_EE4END(Tile_X9Y14_EE4BEG),
    .Tile_X0Y1_E6END(Tile_X9Y14_E6BEG),
    .Tile_X0Y0_N1BEG(Tile_X10Y13_N1BEG),
    .Tile_X0Y0_N2BEG(Tile_X10Y13_N2BEG),
    .Tile_X0Y0_N2BEGb(Tile_X10Y13_N2BEGb),
    .Tile_X0Y0_N4BEG(Tile_X10Y13_N4BEG),
    .Tile_X0Y0_W1BEG(Tile_X10Y13_W1BEG),
    .Tile_X0Y0_W2BEG(Tile_X10Y13_W2BEG),
    .Tile_X0Y0_W2BEGb(Tile_X10Y13_W2BEGb),
    .Tile_X0Y0_WW4BEG(Tile_X10Y13_WW4BEG),
    .Tile_X0Y0_W6BEG(Tile_X10Y13_W6BEG),
    .Tile_X0Y1_S1BEG(Tile_X10Y14_S1BEG),
    .Tile_X0Y1_S2BEG(Tile_X10Y14_S2BEG),
    .Tile_X0Y1_S2BEGb(Tile_X10Y14_S2BEGb),
    .Tile_X0Y1_S4BEG(Tile_X10Y14_S4BEG),
    .Tile_X0Y1_W1BEG(Tile_X10Y14_W1BEG),
    .Tile_X0Y1_W2BEG(Tile_X10Y14_W2BEG),
    .Tile_X0Y1_W2BEGb(Tile_X10Y14_W2BEGb),
    .Tile_X0Y1_WW4BEG(Tile_X10Y14_WW4BEG),
    .Tile_X0Y1_W6BEG(Tile_X10Y14_W6BEG),
    .CONFIGURED_top(Tile_X10Y14_CONFIGURED_top),
    .DOUT_SRAM0(Tile_X10Y14_DOUT_SRAM0),
    .DOUT_SRAM1(Tile_X10Y14_DOUT_SRAM1),
    .DOUT_SRAM2(Tile_X10Y14_DOUT_SRAM2),
    .DOUT_SRAM3(Tile_X10Y14_DOUT_SRAM3),
    .DOUT_SRAM4(Tile_X10Y14_DOUT_SRAM4),
    .DOUT_SRAM5(Tile_X10Y14_DOUT_SRAM5),
    .DOUT_SRAM6(Tile_X10Y14_DOUT_SRAM6),
    .DOUT_SRAM7(Tile_X10Y14_DOUT_SRAM7),
    .DOUT_SRAM8(Tile_X10Y14_DOUT_SRAM8),
    .DOUT_SRAM9(Tile_X10Y14_DOUT_SRAM9),
    .DOUT_SRAM10(Tile_X10Y14_DOUT_SRAM10),
    .DOUT_SRAM11(Tile_X10Y14_DOUT_SRAM11),
    .DOUT_SRAM12(Tile_X10Y14_DOUT_SRAM12),
    .DOUT_SRAM13(Tile_X10Y14_DOUT_SRAM13),
    .DOUT_SRAM14(Tile_X10Y14_DOUT_SRAM14),
    .DOUT_SRAM15(Tile_X10Y14_DOUT_SRAM15),
    .DOUT_SRAM16(Tile_X10Y14_DOUT_SRAM16),
    .DOUT_SRAM17(Tile_X10Y14_DOUT_SRAM17),
    .DOUT_SRAM18(Tile_X10Y14_DOUT_SRAM18),
    .DOUT_SRAM19(Tile_X10Y14_DOUT_SRAM19),
    .DOUT_SRAM20(Tile_X10Y14_DOUT_SRAM20),
    .DOUT_SRAM21(Tile_X10Y14_DOUT_SRAM21),
    .DOUT_SRAM22(Tile_X10Y14_DOUT_SRAM22),
    .DOUT_SRAM23(Tile_X10Y14_DOUT_SRAM23),
    .DOUT_SRAM24(Tile_X10Y14_DOUT_SRAM24),
    .DOUT_SRAM25(Tile_X10Y14_DOUT_SRAM25),
    .DOUT_SRAM26(Tile_X10Y14_DOUT_SRAM26),
    .DOUT_SRAM27(Tile_X10Y14_DOUT_SRAM27),
    .DOUT_SRAM28(Tile_X10Y14_DOUT_SRAM28),
    .DOUT_SRAM29(Tile_X10Y14_DOUT_SRAM29),
    .DOUT_SRAM30(Tile_X10Y14_DOUT_SRAM30),
    .DOUT_SRAM31(Tile_X10Y14_DOUT_SRAM31),
    .ADDR_SRAM0(Tile_X10Y14_ADDR_SRAM0),
    .ADDR_SRAM1(Tile_X10Y14_ADDR_SRAM1),
    .ADDR_SRAM2(Tile_X10Y14_ADDR_SRAM2),
    .ADDR_SRAM3(Tile_X10Y14_ADDR_SRAM3),
    .ADDR_SRAM4(Tile_X10Y14_ADDR_SRAM4),
    .ADDR_SRAM5(Tile_X10Y14_ADDR_SRAM5),
    .ADDR_SRAM6(Tile_X10Y14_ADDR_SRAM6),
    .ADDR_SRAM7(Tile_X10Y14_ADDR_SRAM7),
    .ADDR_SRAM8(Tile_X10Y14_ADDR_SRAM8),
    .ADDR_SRAM9(Tile_X10Y14_ADDR_SRAM9),
    .BM_SRAM0(Tile_X10Y14_BM_SRAM0),
    .BM_SRAM1(Tile_X10Y14_BM_SRAM1),
    .BM_SRAM2(Tile_X10Y14_BM_SRAM2),
    .BM_SRAM3(Tile_X10Y14_BM_SRAM3),
    .BM_SRAM4(Tile_X10Y14_BM_SRAM4),
    .BM_SRAM5(Tile_X10Y14_BM_SRAM5),
    .BM_SRAM6(Tile_X10Y14_BM_SRAM6),
    .BM_SRAM7(Tile_X10Y14_BM_SRAM7),
    .BM_SRAM8(Tile_X10Y14_BM_SRAM8),
    .BM_SRAM9(Tile_X10Y14_BM_SRAM9),
    .BM_SRAM10(Tile_X10Y14_BM_SRAM10),
    .BM_SRAM11(Tile_X10Y14_BM_SRAM11),
    .BM_SRAM12(Tile_X10Y14_BM_SRAM12),
    .BM_SRAM13(Tile_X10Y14_BM_SRAM13),
    .BM_SRAM14(Tile_X10Y14_BM_SRAM14),
    .BM_SRAM15(Tile_X10Y14_BM_SRAM15),
    .BM_SRAM16(Tile_X10Y14_BM_SRAM16),
    .BM_SRAM17(Tile_X10Y14_BM_SRAM17),
    .BM_SRAM18(Tile_X10Y14_BM_SRAM18),
    .BM_SRAM19(Tile_X10Y14_BM_SRAM19),
    .BM_SRAM20(Tile_X10Y14_BM_SRAM20),
    .BM_SRAM21(Tile_X10Y14_BM_SRAM21),
    .BM_SRAM22(Tile_X10Y14_BM_SRAM22),
    .BM_SRAM23(Tile_X10Y14_BM_SRAM23),
    .BM_SRAM24(Tile_X10Y14_BM_SRAM24),
    .BM_SRAM25(Tile_X10Y14_BM_SRAM25),
    .BM_SRAM26(Tile_X10Y14_BM_SRAM26),
    .BM_SRAM27(Tile_X10Y14_BM_SRAM27),
    .BM_SRAM28(Tile_X10Y14_BM_SRAM28),
    .BM_SRAM29(Tile_X10Y14_BM_SRAM29),
    .BM_SRAM30(Tile_X10Y14_BM_SRAM30),
    .BM_SRAM31(Tile_X10Y14_BM_SRAM31),
    .CLK_SRAM(Tile_X10Y14_CLK_SRAM),
    .DIN_SRAM0(Tile_X10Y14_DIN_SRAM0),
    .DIN_SRAM1(Tile_X10Y14_DIN_SRAM1),
    .DIN_SRAM2(Tile_X10Y14_DIN_SRAM2),
    .DIN_SRAM3(Tile_X10Y14_DIN_SRAM3),
    .DIN_SRAM4(Tile_X10Y14_DIN_SRAM4),
    .DIN_SRAM5(Tile_X10Y14_DIN_SRAM5),
    .DIN_SRAM6(Tile_X10Y14_DIN_SRAM6),
    .DIN_SRAM7(Tile_X10Y14_DIN_SRAM7),
    .DIN_SRAM8(Tile_X10Y14_DIN_SRAM8),
    .DIN_SRAM9(Tile_X10Y14_DIN_SRAM9),
    .DIN_SRAM10(Tile_X10Y14_DIN_SRAM10),
    .DIN_SRAM11(Tile_X10Y14_DIN_SRAM11),
    .DIN_SRAM12(Tile_X10Y14_DIN_SRAM12),
    .DIN_SRAM13(Tile_X10Y14_DIN_SRAM13),
    .DIN_SRAM14(Tile_X10Y14_DIN_SRAM14),
    .DIN_SRAM15(Tile_X10Y14_DIN_SRAM15),
    .DIN_SRAM16(Tile_X10Y14_DIN_SRAM16),
    .DIN_SRAM17(Tile_X10Y14_DIN_SRAM17),
    .DIN_SRAM18(Tile_X10Y14_DIN_SRAM18),
    .DIN_SRAM19(Tile_X10Y14_DIN_SRAM19),
    .DIN_SRAM20(Tile_X10Y14_DIN_SRAM20),
    .DIN_SRAM21(Tile_X10Y14_DIN_SRAM21),
    .DIN_SRAM22(Tile_X10Y14_DIN_SRAM22),
    .DIN_SRAM23(Tile_X10Y14_DIN_SRAM23),
    .DIN_SRAM24(Tile_X10Y14_DIN_SRAM24),
    .DIN_SRAM25(Tile_X10Y14_DIN_SRAM25),
    .DIN_SRAM26(Tile_X10Y14_DIN_SRAM26),
    .DIN_SRAM27(Tile_X10Y14_DIN_SRAM27),
    .DIN_SRAM28(Tile_X10Y14_DIN_SRAM28),
    .DIN_SRAM29(Tile_X10Y14_DIN_SRAM29),
    .DIN_SRAM30(Tile_X10Y14_DIN_SRAM30),
    .DIN_SRAM31(Tile_X10Y14_DIN_SRAM31),
    .MEN_SRAM(Tile_X10Y14_MEN_SRAM),
    .REN_SRAM(Tile_X10Y14_REN_SRAM),
    .TIE_HIGH_SRAM(Tile_X10Y14_TIE_HIGH_SRAM),
    .TIE_LOW_SRAM(Tile_X10Y14_TIE_LOW_SRAM),
    .WEN_SRAM(Tile_X10Y14_WEN_SRAM),
    .Tile_X0Y0_UserCLKo(Tile_X10Y13_UserCLKo),
    .Tile_X0Y1_UserCLK(Tile_X10Y15_UserCLKo),
    .Tile_X0Y0_FrameData(Tile_X9Y13_FrameData_O),
    .Tile_X0Y0_FrameData_O(Tile_X10Y13_FrameData_O),
    .Tile_X0Y0_FrameStrobe_O(Tile_X10Y13_FrameStrobe_O),
    .Tile_X0Y1_FrameData(Tile_X9Y14_FrameData_O),
    .Tile_X0Y1_FrameData_O(Tile_X10Y14_FrameData_O),
    .Tile_X0Y1_FrameStrobe(Tile_X10Y15_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
W_IO
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X0Y14_Emulate_Bitstream)
    )
`endif
    Tile_X0Y14_W_IO
    (
    .W1END(Tile_X1Y14_W1BEG),
    .W2MID(Tile_X1Y14_W2BEG),
    .W2END(Tile_X1Y14_W2BEGb),
    .WW4END(Tile_X1Y14_WW4BEG),
    .W6END(Tile_X1Y14_W6BEG),
    .E1BEG(Tile_X0Y14_E1BEG),
    .E2BEG(Tile_X0Y14_E2BEG),
    .E2BEGb(Tile_X0Y14_E2BEGb),
    .EE4BEG(Tile_X0Y14_EE4BEG),
    .E6BEG(Tile_X0Y14_E6BEG),
    .A_O_top(Tile_X0Y14_A_O_top),
    .A_I_top(Tile_X0Y14_A_I_top),
    .A_T_top(Tile_X0Y14_A_T_top),
    .B_O_top(Tile_X0Y14_B_O_top),
    .B_I_top(Tile_X0Y14_B_I_top),
    .B_T_top(Tile_X0Y14_B_T_top),
    .A_config_C_bit0(Tile_X0Y14_A_config_C_bit0),
    .A_config_C_bit1(Tile_X0Y14_A_config_C_bit1),
    .A_config_C_bit2(Tile_X0Y14_A_config_C_bit2),
    .A_config_C_bit3(Tile_X0Y14_A_config_C_bit3),
    .B_config_C_bit0(Tile_X0Y14_B_config_C_bit0),
    .B_config_C_bit1(Tile_X0Y14_B_config_C_bit1),
    .B_config_C_bit2(Tile_X0Y14_B_config_C_bit2),
    .B_config_C_bit3(Tile_X0Y14_B_config_C_bit3),
    .UserCLK(UserCLK),
    .UserCLKo(Tile_X0Y14_UserCLKo),
    .FrameData(Row_Y14_FrameData),
    .FrameData_O(Tile_X0Y14_FrameData_O),
    .FrameStrobe(Column_X0_FrameStrobe),
    .FrameStrobe_O(Tile_X0Y14_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X1Y14_Emulate_Bitstream)
    )
`endif
    Tile_X1Y14_LUT4AB
    (
    .N1END(Tile_X1Y15_N1BEG),
    .N2MID(Tile_X1Y15_N2BEG),
    .N2END(Tile_X1Y15_N2BEGb),
    .N4END(Tile_X1Y15_N4BEG),
    .NN4END(Tile_X1Y15_NN4BEG),
    .Ci(Tile_X1Y15_Co),
    .E1END(Tile_X0Y14_E1BEG),
    .E2MID(Tile_X0Y14_E2BEG),
    .E2END(Tile_X0Y14_E2BEGb),
    .EE4END(Tile_X0Y14_EE4BEG),
    .E6END(Tile_X0Y14_E6BEG),
    .S1END(Tile_X1Y13_S1BEG),
    .S2MID(Tile_X1Y13_S2BEG),
    .S2END(Tile_X1Y13_S2BEGb),
    .S4END(Tile_X1Y13_S4BEG),
    .SS4END(Tile_X1Y13_SS4BEG),
    .W1END(Tile_X2Y14_W1BEG),
    .W2MID(Tile_X2Y14_W2BEG),
    .W2END(Tile_X2Y14_W2BEGb),
    .WW4END(Tile_X2Y14_WW4BEG),
    .W6END(Tile_X2Y14_W6BEG),
    .N1BEG(Tile_X1Y14_N1BEG),
    .N2BEG(Tile_X1Y14_N2BEG),
    .N2BEGb(Tile_X1Y14_N2BEGb),
    .N4BEG(Tile_X1Y14_N4BEG),
    .NN4BEG(Tile_X1Y14_NN4BEG),
    .E1BEG(Tile_X1Y14_E1BEG),
    .E2BEG(Tile_X1Y14_E2BEG),
    .E2BEGb(Tile_X1Y14_E2BEGb),
    .EE4BEG(Tile_X1Y14_EE4BEG),
    .E6BEG(Tile_X1Y14_E6BEG),
    .S1BEG(Tile_X1Y14_S1BEG),
    .S2BEG(Tile_X1Y14_S2BEG),
    .S2BEGb(Tile_X1Y14_S2BEGb),
    .S4BEG(Tile_X1Y14_S4BEG),
    .SS4BEG(Tile_X1Y14_SS4BEG),
    .W1BEG(Tile_X1Y14_W1BEG),
    .W2BEG(Tile_X1Y14_W2BEG),
    .W2BEGb(Tile_X1Y14_W2BEGb),
    .WW4BEG(Tile_X1Y14_WW4BEG),
    .W6BEG(Tile_X1Y14_W6BEG),
    .Co(Tile_X1Y14_Co),
    .UserCLK(Tile_X1Y15_UserCLKo),
    .UserCLKo(Tile_X1Y14_UserCLKo),
    .FrameData(Tile_X0Y14_FrameData_O),
    .FrameData_O(Tile_X1Y14_FrameData_O),
    .FrameStrobe(Tile_X1Y15_FrameStrobe_O),
    .FrameStrobe_O(Tile_X1Y14_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X2Y14_Emulate_Bitstream)
    )
`endif
    Tile_X2Y14_LUT4AB
    (
    .N1END(Tile_X2Y15_N1BEG),
    .N2MID(Tile_X2Y15_N2BEG),
    .N2END(Tile_X2Y15_N2BEGb),
    .N4END(Tile_X2Y15_N4BEG),
    .NN4END(Tile_X2Y15_NN4BEG),
    .Ci(Tile_X2Y15_Co),
    .E1END(Tile_X1Y14_E1BEG),
    .E2MID(Tile_X1Y14_E2BEG),
    .E2END(Tile_X1Y14_E2BEGb),
    .EE4END(Tile_X1Y14_EE4BEG),
    .E6END(Tile_X1Y14_E6BEG),
    .S1END(Tile_X2Y13_S1BEG),
    .S2MID(Tile_X2Y13_S2BEG),
    .S2END(Tile_X2Y13_S2BEGb),
    .S4END(Tile_X2Y13_S4BEG),
    .SS4END(Tile_X2Y13_SS4BEG),
    .W1END(Tile_X3Y14_W1BEG),
    .W2MID(Tile_X3Y14_W2BEG),
    .W2END(Tile_X3Y14_W2BEGb),
    .WW4END(Tile_X3Y14_WW4BEG),
    .W6END(Tile_X3Y14_W6BEG),
    .N1BEG(Tile_X2Y14_N1BEG),
    .N2BEG(Tile_X2Y14_N2BEG),
    .N2BEGb(Tile_X2Y14_N2BEGb),
    .N4BEG(Tile_X2Y14_N4BEG),
    .NN4BEG(Tile_X2Y14_NN4BEG),
    .E1BEG(Tile_X2Y14_E1BEG),
    .E2BEG(Tile_X2Y14_E2BEG),
    .E2BEGb(Tile_X2Y14_E2BEGb),
    .EE4BEG(Tile_X2Y14_EE4BEG),
    .E6BEG(Tile_X2Y14_E6BEG),
    .S1BEG(Tile_X2Y14_S1BEG),
    .S2BEG(Tile_X2Y14_S2BEG),
    .S2BEGb(Tile_X2Y14_S2BEGb),
    .S4BEG(Tile_X2Y14_S4BEG),
    .SS4BEG(Tile_X2Y14_SS4BEG),
    .W1BEG(Tile_X2Y14_W1BEG),
    .W2BEG(Tile_X2Y14_W2BEG),
    .W2BEGb(Tile_X2Y14_W2BEGb),
    .WW4BEG(Tile_X2Y14_WW4BEG),
    .W6BEG(Tile_X2Y14_W6BEG),
    .Co(Tile_X2Y14_Co),
    .UserCLK(Tile_X2Y15_UserCLKo),
    .UserCLKo(Tile_X2Y14_UserCLKo),
    .FrameData(Tile_X1Y14_FrameData_O),
    .FrameData_O(Tile_X2Y14_FrameData_O),
    .FrameStrobe(Tile_X2Y15_FrameStrobe_O),
    .FrameStrobe_O(Tile_X2Y14_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X3Y14_Emulate_Bitstream)
    )
`endif
    Tile_X3Y14_LUT4AB
    (
    .N1END(Tile_X3Y15_N1BEG),
    .N2MID(Tile_X3Y15_N2BEG),
    .N2END(Tile_X3Y15_N2BEGb),
    .N4END(Tile_X3Y15_N4BEG),
    .NN4END(Tile_X3Y15_NN4BEG),
    .Ci(Tile_X3Y15_Co),
    .E1END(Tile_X2Y14_E1BEG),
    .E2MID(Tile_X2Y14_E2BEG),
    .E2END(Tile_X2Y14_E2BEGb),
    .EE4END(Tile_X2Y14_EE4BEG),
    .E6END(Tile_X2Y14_E6BEG),
    .S1END(Tile_X3Y13_S1BEG),
    .S2MID(Tile_X3Y13_S2BEG),
    .S2END(Tile_X3Y13_S2BEGb),
    .S4END(Tile_X3Y13_S4BEG),
    .SS4END(Tile_X3Y13_SS4BEG),
    .W1END(Tile_X4Y14_W1BEG),
    .W2MID(Tile_X4Y14_W2BEG),
    .W2END(Tile_X4Y14_W2BEGb),
    .WW4END(Tile_X4Y14_WW4BEG),
    .W6END(Tile_X4Y14_W6BEG),
    .N1BEG(Tile_X3Y14_N1BEG),
    .N2BEG(Tile_X3Y14_N2BEG),
    .N2BEGb(Tile_X3Y14_N2BEGb),
    .N4BEG(Tile_X3Y14_N4BEG),
    .NN4BEG(Tile_X3Y14_NN4BEG),
    .E1BEG(Tile_X3Y14_E1BEG),
    .E2BEG(Tile_X3Y14_E2BEG),
    .E2BEGb(Tile_X3Y14_E2BEGb),
    .EE4BEG(Tile_X3Y14_EE4BEG),
    .E6BEG(Tile_X3Y14_E6BEG),
    .S1BEG(Tile_X3Y14_S1BEG),
    .S2BEG(Tile_X3Y14_S2BEG),
    .S2BEGb(Tile_X3Y14_S2BEGb),
    .S4BEG(Tile_X3Y14_S4BEG),
    .SS4BEG(Tile_X3Y14_SS4BEG),
    .W1BEG(Tile_X3Y14_W1BEG),
    .W2BEG(Tile_X3Y14_W2BEG),
    .W2BEGb(Tile_X3Y14_W2BEGb),
    .WW4BEG(Tile_X3Y14_WW4BEG),
    .W6BEG(Tile_X3Y14_W6BEG),
    .Co(Tile_X3Y14_Co),
    .UserCLK(Tile_X3Y15_UserCLKo),
    .UserCLKo(Tile_X3Y14_UserCLKo),
    .FrameData(Tile_X2Y14_FrameData_O),
    .FrameData_O(Tile_X3Y14_FrameData_O),
    .FrameStrobe(Tile_X3Y15_FrameStrobe_O),
    .FrameStrobe_O(Tile_X3Y14_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
RegFile
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X4Y14_Emulate_Bitstream)
    )
`endif
    Tile_X4Y14_RegFile
    (
    .N1END(Tile_X4Y15_N1BEG),
    .N2MID(Tile_X4Y15_N2BEG),
    .N2END(Tile_X4Y15_N2BEGb),
    .N4END(Tile_X4Y15_N4BEG),
    .NN4END(Tile_X4Y15_NN4BEG),
    .E1END(Tile_X3Y14_E1BEG),
    .E2MID(Tile_X3Y14_E2BEG),
    .E2END(Tile_X3Y14_E2BEGb),
    .EE4END(Tile_X3Y14_EE4BEG),
    .E6END(Tile_X3Y14_E6BEG),
    .S1END(Tile_X4Y13_S1BEG),
    .S2MID(Tile_X4Y13_S2BEG),
    .S2END(Tile_X4Y13_S2BEGb),
    .S4END(Tile_X4Y13_S4BEG),
    .SS4END(Tile_X4Y13_SS4BEG),
    .W1END(Tile_X5Y14_W1BEG),
    .W2MID(Tile_X5Y14_W2BEG),
    .W2END(Tile_X5Y14_W2BEGb),
    .WW4END(Tile_X5Y14_WW4BEG),
    .W6END(Tile_X5Y14_W6BEG),
    .N1BEG(Tile_X4Y14_N1BEG),
    .N2BEG(Tile_X4Y14_N2BEG),
    .N2BEGb(Tile_X4Y14_N2BEGb),
    .N4BEG(Tile_X4Y14_N4BEG),
    .NN4BEG(Tile_X4Y14_NN4BEG),
    .E1BEG(Tile_X4Y14_E1BEG),
    .E2BEG(Tile_X4Y14_E2BEG),
    .E2BEGb(Tile_X4Y14_E2BEGb),
    .EE4BEG(Tile_X4Y14_EE4BEG),
    .E6BEG(Tile_X4Y14_E6BEG),
    .S1BEG(Tile_X4Y14_S1BEG),
    .S2BEG(Tile_X4Y14_S2BEG),
    .S2BEGb(Tile_X4Y14_S2BEGb),
    .S4BEG(Tile_X4Y14_S4BEG),
    .SS4BEG(Tile_X4Y14_SS4BEG),
    .W1BEG(Tile_X4Y14_W1BEG),
    .W2BEG(Tile_X4Y14_W2BEG),
    .W2BEGb(Tile_X4Y14_W2BEGb),
    .WW4BEG(Tile_X4Y14_WW4BEG),
    .W6BEG(Tile_X4Y14_W6BEG),
    .UserCLK(Tile_X4Y15_UserCLKo),
    .UserCLKo(Tile_X4Y14_UserCLKo),
    .FrameData(Tile_X3Y14_FrameData_O),
    .FrameData_O(Tile_X4Y14_FrameData_O),
    .FrameStrobe(Tile_X4Y15_FrameStrobe_O),
    .FrameStrobe_O(Tile_X4Y14_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X5Y14_Emulate_Bitstream)
    )
`endif
    Tile_X5Y14_LUT4AB
    (
    .N1END(Tile_X5Y15_N1BEG),
    .N2MID(Tile_X5Y15_N2BEG),
    .N2END(Tile_X5Y15_N2BEGb),
    .N4END(Tile_X5Y15_N4BEG),
    .NN4END(Tile_X5Y15_NN4BEG),
    .Ci(Tile_X5Y15_Co),
    .E1END(Tile_X4Y14_E1BEG),
    .E2MID(Tile_X4Y14_E2BEG),
    .E2END(Tile_X4Y14_E2BEGb),
    .EE4END(Tile_X4Y14_EE4BEG),
    .E6END(Tile_X4Y14_E6BEG),
    .S1END(Tile_X5Y13_S1BEG),
    .S2MID(Tile_X5Y13_S2BEG),
    .S2END(Tile_X5Y13_S2BEGb),
    .S4END(Tile_X5Y13_S4BEG),
    .SS4END(Tile_X5Y13_SS4BEG),
    .W1END(Tile_X6Y14_W1BEG),
    .W2MID(Tile_X6Y14_W2BEG),
    .W2END(Tile_X6Y14_W2BEGb),
    .WW4END(Tile_X6Y14_WW4BEG),
    .W6END(Tile_X6Y14_W6BEG),
    .N1BEG(Tile_X5Y14_N1BEG),
    .N2BEG(Tile_X5Y14_N2BEG),
    .N2BEGb(Tile_X5Y14_N2BEGb),
    .N4BEG(Tile_X5Y14_N4BEG),
    .NN4BEG(Tile_X5Y14_NN4BEG),
    .E1BEG(Tile_X5Y14_E1BEG),
    .E2BEG(Tile_X5Y14_E2BEG),
    .E2BEGb(Tile_X5Y14_E2BEGb),
    .EE4BEG(Tile_X5Y14_EE4BEG),
    .E6BEG(Tile_X5Y14_E6BEG),
    .S1BEG(Tile_X5Y14_S1BEG),
    .S2BEG(Tile_X5Y14_S2BEG),
    .S2BEGb(Tile_X5Y14_S2BEGb),
    .S4BEG(Tile_X5Y14_S4BEG),
    .SS4BEG(Tile_X5Y14_SS4BEG),
    .W1BEG(Tile_X5Y14_W1BEG),
    .W2BEG(Tile_X5Y14_W2BEG),
    .W2BEGb(Tile_X5Y14_W2BEGb),
    .WW4BEG(Tile_X5Y14_WW4BEG),
    .W6BEG(Tile_X5Y14_W6BEG),
    .Co(Tile_X5Y14_Co),
    .UserCLK(Tile_X5Y15_UserCLKo),
    .UserCLKo(Tile_X5Y14_UserCLKo),
    .FrameData(Tile_X4Y14_FrameData_O),
    .FrameData_O(Tile_X5Y14_FrameData_O),
    .FrameStrobe(Tile_X5Y15_FrameStrobe_O),
    .FrameStrobe_O(Tile_X5Y14_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X6Y14_Emulate_Bitstream)
    )
`endif
    Tile_X6Y14_LUT4AB
    (
    .N1END(Tile_X6Y15_N1BEG),
    .N2MID(Tile_X6Y15_N2BEG),
    .N2END(Tile_X6Y15_N2BEGb),
    .N4END(Tile_X6Y15_N4BEG),
    .NN4END(Tile_X6Y15_NN4BEG),
    .Ci(Tile_X6Y15_Co),
    .E1END(Tile_X5Y14_E1BEG),
    .E2MID(Tile_X5Y14_E2BEG),
    .E2END(Tile_X5Y14_E2BEGb),
    .EE4END(Tile_X5Y14_EE4BEG),
    .E6END(Tile_X5Y14_E6BEG),
    .S1END(Tile_X6Y13_S1BEG),
    .S2MID(Tile_X6Y13_S2BEG),
    .S2END(Tile_X6Y13_S2BEGb),
    .S4END(Tile_X6Y13_S4BEG),
    .SS4END(Tile_X6Y13_SS4BEG),
    .W1END(Tile_X7Y14_W1BEG),
    .W2MID(Tile_X7Y14_W2BEG),
    .W2END(Tile_X7Y14_W2BEGb),
    .WW4END(Tile_X7Y14_WW4BEG),
    .W6END(Tile_X7Y14_W6BEG),
    .N1BEG(Tile_X6Y14_N1BEG),
    .N2BEG(Tile_X6Y14_N2BEG),
    .N2BEGb(Tile_X6Y14_N2BEGb),
    .N4BEG(Tile_X6Y14_N4BEG),
    .NN4BEG(Tile_X6Y14_NN4BEG),
    .E1BEG(Tile_X6Y14_E1BEG),
    .E2BEG(Tile_X6Y14_E2BEG),
    .E2BEGb(Tile_X6Y14_E2BEGb),
    .EE4BEG(Tile_X6Y14_EE4BEG),
    .E6BEG(Tile_X6Y14_E6BEG),
    .S1BEG(Tile_X6Y14_S1BEG),
    .S2BEG(Tile_X6Y14_S2BEG),
    .S2BEGb(Tile_X6Y14_S2BEGb),
    .S4BEG(Tile_X6Y14_S4BEG),
    .SS4BEG(Tile_X6Y14_SS4BEG),
    .W1BEG(Tile_X6Y14_W1BEG),
    .W2BEG(Tile_X6Y14_W2BEG),
    .W2BEGb(Tile_X6Y14_W2BEGb),
    .WW4BEG(Tile_X6Y14_WW4BEG),
    .W6BEG(Tile_X6Y14_W6BEG),
    .Co(Tile_X6Y14_Co),
    .UserCLK(Tile_X6Y15_UserCLKo),
    .UserCLKo(Tile_X6Y14_UserCLKo),
    .FrameData(Tile_X5Y14_FrameData_O),
    .FrameData_O(Tile_X6Y14_FrameData_O),
    .FrameStrobe(Tile_X6Y15_FrameStrobe_O),
    .FrameStrobe_O(Tile_X6Y14_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X8Y14_Emulate_Bitstream)
    )
`endif
    Tile_X8Y14_LUT4AB
    (
    .N1END(Tile_X8Y15_N1BEG),
    .N2MID(Tile_X8Y15_N2BEG),
    .N2END(Tile_X8Y15_N2BEGb),
    .N4END(Tile_X8Y15_N4BEG),
    .NN4END(Tile_X8Y15_NN4BEG),
    .Ci(Tile_X8Y15_Co),
    .E1END(Tile_X7Y14_E1BEG),
    .E2MID(Tile_X7Y14_E2BEG),
    .E2END(Tile_X7Y14_E2BEGb),
    .EE4END(Tile_X7Y14_EE4BEG),
    .E6END(Tile_X7Y14_E6BEG),
    .S1END(Tile_X8Y13_S1BEG),
    .S2MID(Tile_X8Y13_S2BEG),
    .S2END(Tile_X8Y13_S2BEGb),
    .S4END(Tile_X8Y13_S4BEG),
    .SS4END(Tile_X8Y13_SS4BEG),
    .W1END(Tile_X9Y14_W1BEG),
    .W2MID(Tile_X9Y14_W2BEG),
    .W2END(Tile_X9Y14_W2BEGb),
    .WW4END(Tile_X9Y14_WW4BEG),
    .W6END(Tile_X9Y14_W6BEG),
    .N1BEG(Tile_X8Y14_N1BEG),
    .N2BEG(Tile_X8Y14_N2BEG),
    .N2BEGb(Tile_X8Y14_N2BEGb),
    .N4BEG(Tile_X8Y14_N4BEG),
    .NN4BEG(Tile_X8Y14_NN4BEG),
    .E1BEG(Tile_X8Y14_E1BEG),
    .E2BEG(Tile_X8Y14_E2BEG),
    .E2BEGb(Tile_X8Y14_E2BEGb),
    .EE4BEG(Tile_X8Y14_EE4BEG),
    .E6BEG(Tile_X8Y14_E6BEG),
    .S1BEG(Tile_X8Y14_S1BEG),
    .S2BEG(Tile_X8Y14_S2BEG),
    .S2BEGb(Tile_X8Y14_S2BEGb),
    .S4BEG(Tile_X8Y14_S4BEG),
    .SS4BEG(Tile_X8Y14_SS4BEG),
    .W1BEG(Tile_X8Y14_W1BEG),
    .W2BEG(Tile_X8Y14_W2BEG),
    .W2BEGb(Tile_X8Y14_W2BEGb),
    .WW4BEG(Tile_X8Y14_WW4BEG),
    .W6BEG(Tile_X8Y14_W6BEG),
    .Co(Tile_X8Y14_Co),
    .UserCLK(Tile_X8Y15_UserCLKo),
    .UserCLKo(Tile_X8Y14_UserCLKo),
    .FrameData(Tile_X7Y14_FrameData_O),
    .FrameData_O(Tile_X8Y14_FrameData_O),
    .FrameStrobe(Tile_X8Y15_FrameStrobe_O),
    .FrameStrobe_O(Tile_X8Y14_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X9Y14_Emulate_Bitstream)
    )
`endif
    Tile_X9Y14_LUT4AB
    (
    .N1END(Tile_X9Y15_N1BEG),
    .N2MID(Tile_X9Y15_N2BEG),
    .N2END(Tile_X9Y15_N2BEGb),
    .N4END(Tile_X9Y15_N4BEG),
    .NN4END(Tile_X9Y15_NN4BEG),
    .Ci(Tile_X9Y15_Co),
    .E1END(Tile_X8Y14_E1BEG),
    .E2MID(Tile_X8Y14_E2BEG),
    .E2END(Tile_X8Y14_E2BEGb),
    .EE4END(Tile_X8Y14_EE4BEG),
    .E6END(Tile_X8Y14_E6BEG),
    .S1END(Tile_X9Y13_S1BEG),
    .S2MID(Tile_X9Y13_S2BEG),
    .S2END(Tile_X9Y13_S2BEGb),
    .S4END(Tile_X9Y13_S4BEG),
    .SS4END(Tile_X9Y13_SS4BEG),
    .W1END(Tile_X10Y14_W1BEG),
    .W2MID(Tile_X10Y14_W2BEG),
    .W2END(Tile_X10Y14_W2BEGb),
    .WW4END(Tile_X10Y14_WW4BEG),
    .W6END(Tile_X10Y14_W6BEG),
    .N1BEG(Tile_X9Y14_N1BEG),
    .N2BEG(Tile_X9Y14_N2BEG),
    .N2BEGb(Tile_X9Y14_N2BEGb),
    .N4BEG(Tile_X9Y14_N4BEG),
    .NN4BEG(Tile_X9Y14_NN4BEG),
    .E1BEG(Tile_X9Y14_E1BEG),
    .E2BEG(Tile_X9Y14_E2BEG),
    .E2BEGb(Tile_X9Y14_E2BEGb),
    .EE4BEG(Tile_X9Y14_EE4BEG),
    .E6BEG(Tile_X9Y14_E6BEG),
    .S1BEG(Tile_X9Y14_S1BEG),
    .S2BEG(Tile_X9Y14_S2BEG),
    .S2BEGb(Tile_X9Y14_S2BEGb),
    .S4BEG(Tile_X9Y14_S4BEG),
    .SS4BEG(Tile_X9Y14_SS4BEG),
    .W1BEG(Tile_X9Y14_W1BEG),
    .W2BEG(Tile_X9Y14_W2BEG),
    .W2BEGb(Tile_X9Y14_W2BEGb),
    .WW4BEG(Tile_X9Y14_WW4BEG),
    .W6BEG(Tile_X9Y14_W6BEG),
    .Co(Tile_X9Y14_Co),
    .UserCLK(Tile_X9Y15_UserCLKo),
    .UserCLKo(Tile_X9Y14_UserCLKo),
    .FrameData(Tile_X8Y14_FrameData_O),
    .FrameData_O(Tile_X9Y14_FrameData_O),
    .FrameStrobe(Tile_X9Y15_FrameStrobe_O),
    .FrameStrobe_O(Tile_X9Y14_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
S_term_single Tile_X1Y15_S_term_single (
    .S1END(Tile_X1Y14_S1BEG),
    .S2MID(Tile_X1Y14_S2BEG),
    .S2END(Tile_X1Y14_S2BEGb),
    .S4END(Tile_X1Y14_S4BEG),
    .SS4END(Tile_X1Y14_SS4BEG),
    .N1BEG(Tile_X1Y15_N1BEG),
    .N2BEG(Tile_X1Y15_N2BEG),
    .N2BEGb(Tile_X1Y15_N2BEGb),
    .N4BEG(Tile_X1Y15_N4BEG),
    .NN4BEG(Tile_X1Y15_NN4BEG),
    .Co(Tile_X1Y15_Co),
    .UserCLK(UserCLK),
    .UserCLKo(Tile_X1Y15_UserCLKo),
    .FrameData(Row_Y15_FrameData),
    .FrameData_O(Tile_X1Y15_FrameData_O),
    .FrameStrobe(Column_X1_FrameStrobe),
    .FrameStrobe_O(Tile_X1Y15_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
S_WARMBOOT Tile_X2Y15_S_WARMBOOT (
    .S1END(Tile_X2Y14_S1BEG),
    .S2MID(Tile_X2Y14_S2BEG),
    .S2END(Tile_X2Y14_S2BEGb),
    .S4END(Tile_X2Y14_S4BEG),
    .SS4END(Tile_X2Y14_SS4BEG),
    .N1BEG(Tile_X2Y15_N1BEG),
    .N2BEG(Tile_X2Y15_N2BEG),
    .N2BEGb(Tile_X2Y15_N2BEGb),
    .N4BEG(Tile_X2Y15_N4BEG),
    .NN4BEG(Tile_X2Y15_NN4BEG),
    .Co(Tile_X2Y15_Co),
    .CONFIGURED_top(Tile_X2Y15_CONFIGURED_top),
    .RESET_top(Tile_X2Y15_RESET_top),
    .BOOT_top(Tile_X2Y15_BOOT_top),
    .SLOT_top0(Tile_X2Y15_SLOT_top0),
    .SLOT_top1(Tile_X2Y15_SLOT_top1),
    .SLOT_top2(Tile_X2Y15_SLOT_top2),
    .SLOT_top3(Tile_X2Y15_SLOT_top3),
    .UserCLK(UserCLK),
    .UserCLKo(Tile_X2Y15_UserCLKo),
    .FrameData(Tile_X1Y15_FrameData_O),
    .FrameData_O(Tile_X2Y15_FrameData_O),
    .FrameStrobe(Column_X2_FrameStrobe),
    .FrameStrobe_O(Tile_X2Y15_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
S_CPU_IRQ Tile_X3Y15_S_CPU_IRQ (
    .S1END(Tile_X3Y14_S1BEG),
    .S2MID(Tile_X3Y14_S2BEG),
    .S2END(Tile_X3Y14_S2BEGb),
    .S4END(Tile_X3Y14_S4BEG),
    .SS4END(Tile_X3Y14_SS4BEG),
    .N1BEG(Tile_X3Y15_N1BEG),
    .N2BEG(Tile_X3Y15_N2BEG),
    .N2BEGb(Tile_X3Y15_N2BEGb),
    .N4BEG(Tile_X3Y15_N4BEG),
    .NN4BEG(Tile_X3Y15_NN4BEG),
    .Co(Tile_X3Y15_Co),
    .CONFIGURED_top(Tile_X3Y15_CONFIGURED_top),
    .IRQ_top0(Tile_X3Y15_IRQ_top0),
    .IRQ_top1(Tile_X3Y15_IRQ_top1),
    .IRQ_top2(Tile_X3Y15_IRQ_top2),
    .IRQ_top3(Tile_X3Y15_IRQ_top3),
    .UserCLK(UserCLK),
    .UserCLKo(Tile_X3Y15_UserCLKo),
    .FrameData(Tile_X2Y15_FrameData_O),
    .FrameData_O(Tile_X3Y15_FrameData_O),
    .FrameStrobe(Column_X3_FrameStrobe),
    .FrameStrobe_O(Tile_X3Y15_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
S_term_single2 Tile_X4Y15_S_term_single2 (
    .S1END(Tile_X4Y14_S1BEG),
    .S2MID(Tile_X4Y14_S2BEG),
    .S2END(Tile_X4Y14_S2BEGb),
    .S4END(Tile_X4Y14_S4BEG),
    .SS4END(Tile_X4Y14_SS4BEG),
    .N1BEG(Tile_X4Y15_N1BEG),
    .N2BEG(Tile_X4Y15_N2BEG),
    .N2BEGb(Tile_X4Y15_N2BEGb),
    .N4BEG(Tile_X4Y15_N4BEG),
    .NN4BEG(Tile_X4Y15_NN4BEG),
    .UserCLK(UserCLK),
    .UserCLKo(Tile_X4Y15_UserCLKo),
    .FrameData(Tile_X3Y15_FrameData_O),
    .FrameData_O(Tile_X4Y15_FrameData_O),
    .FrameStrobe(Column_X4_FrameStrobe),
    .FrameStrobe_O(Tile_X4Y15_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
S_CPU_IF Tile_X5Y15_S_CPU_IF (
    .S1END(Tile_X5Y14_S1BEG),
    .S2MID(Tile_X5Y14_S2BEG),
    .S2END(Tile_X5Y14_S2BEGb),
    .S4END(Tile_X5Y14_S4BEG),
    .SS4END(Tile_X5Y14_SS4BEG),
    .N1BEG(Tile_X5Y15_N1BEG),
    .N2BEG(Tile_X5Y15_N2BEG),
    .N2BEGb(Tile_X5Y15_N2BEGb),
    .N4BEG(Tile_X5Y15_N4BEG),
    .NN4BEG(Tile_X5Y15_NN4BEG),
    .Co(Tile_X5Y15_Co),
    .O_top0(Tile_X5Y15_O_top0),
    .O_top1(Tile_X5Y15_O_top1),
    .O_top2(Tile_X5Y15_O_top2),
    .O_top3(Tile_X5Y15_O_top3),
    .O_top4(Tile_X5Y15_O_top4),
    .O_top5(Tile_X5Y15_O_top5),
    .O_top6(Tile_X5Y15_O_top6),
    .O_top7(Tile_X5Y15_O_top7),
    .O_top8(Tile_X5Y15_O_top8),
    .O_top9(Tile_X5Y15_O_top9),
    .O_top10(Tile_X5Y15_O_top10),
    .O_top11(Tile_X5Y15_O_top11),
    .O_top12(Tile_X5Y15_O_top12),
    .O_top13(Tile_X5Y15_O_top13),
    .O_top14(Tile_X5Y15_O_top14),
    .O_top15(Tile_X5Y15_O_top15),
    .I_top0(Tile_X5Y15_I_top0),
    .I_top1(Tile_X5Y15_I_top1),
    .I_top2(Tile_X5Y15_I_top2),
    .I_top3(Tile_X5Y15_I_top3),
    .I_top4(Tile_X5Y15_I_top4),
    .I_top5(Tile_X5Y15_I_top5),
    .I_top6(Tile_X5Y15_I_top6),
    .I_top7(Tile_X5Y15_I_top7),
    .I_top8(Tile_X5Y15_I_top8),
    .I_top9(Tile_X5Y15_I_top9),
    .I_top10(Tile_X5Y15_I_top10),
    .I_top11(Tile_X5Y15_I_top11),
    .I_top12(Tile_X5Y15_I_top12),
    .I_top13(Tile_X5Y15_I_top13),
    .I_top14(Tile_X5Y15_I_top14),
    .I_top15(Tile_X5Y15_I_top15),
    .UserCLK(UserCLK),
    .UserCLKo(Tile_X5Y15_UserCLKo),
    .FrameData(Tile_X4Y15_FrameData_O),
    .FrameData_O(Tile_X5Y15_FrameData_O),
    .FrameStrobe(Column_X5_FrameStrobe),
    .FrameStrobe_O(Tile_X5Y15_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
S_CPU_IF Tile_X6Y15_S_CPU_IF (
    .S1END(Tile_X6Y14_S1BEG),
    .S2MID(Tile_X6Y14_S2BEG),
    .S2END(Tile_X6Y14_S2BEGb),
    .S4END(Tile_X6Y14_S4BEG),
    .SS4END(Tile_X6Y14_SS4BEG),
    .N1BEG(Tile_X6Y15_N1BEG),
    .N2BEG(Tile_X6Y15_N2BEG),
    .N2BEGb(Tile_X6Y15_N2BEGb),
    .N4BEG(Tile_X6Y15_N4BEG),
    .NN4BEG(Tile_X6Y15_NN4BEG),
    .Co(Tile_X6Y15_Co),
    .O_top0(Tile_X6Y15_O_top0),
    .O_top1(Tile_X6Y15_O_top1),
    .O_top2(Tile_X6Y15_O_top2),
    .O_top3(Tile_X6Y15_O_top3),
    .O_top4(Tile_X6Y15_O_top4),
    .O_top5(Tile_X6Y15_O_top5),
    .O_top6(Tile_X6Y15_O_top6),
    .O_top7(Tile_X6Y15_O_top7),
    .O_top8(Tile_X6Y15_O_top8),
    .O_top9(Tile_X6Y15_O_top9),
    .O_top10(Tile_X6Y15_O_top10),
    .O_top11(Tile_X6Y15_O_top11),
    .O_top12(Tile_X6Y15_O_top12),
    .O_top13(Tile_X6Y15_O_top13),
    .O_top14(Tile_X6Y15_O_top14),
    .O_top15(Tile_X6Y15_O_top15),
    .I_top0(Tile_X6Y15_I_top0),
    .I_top1(Tile_X6Y15_I_top1),
    .I_top2(Tile_X6Y15_I_top2),
    .I_top3(Tile_X6Y15_I_top3),
    .I_top4(Tile_X6Y15_I_top4),
    .I_top5(Tile_X6Y15_I_top5),
    .I_top6(Tile_X6Y15_I_top6),
    .I_top7(Tile_X6Y15_I_top7),
    .I_top8(Tile_X6Y15_I_top8),
    .I_top9(Tile_X6Y15_I_top9),
    .I_top10(Tile_X6Y15_I_top10),
    .I_top11(Tile_X6Y15_I_top11),
    .I_top12(Tile_X6Y15_I_top12),
    .I_top13(Tile_X6Y15_I_top13),
    .I_top14(Tile_X6Y15_I_top14),
    .I_top15(Tile_X6Y15_I_top15),
    .UserCLK(UserCLK),
    .UserCLKo(Tile_X6Y15_UserCLKo),
    .FrameData(Tile_X5Y15_FrameData_O),
    .FrameData_O(Tile_X6Y15_FrameData_O),
    .FrameStrobe(Column_X6_FrameStrobe),
    .FrameStrobe_O(Tile_X6Y15_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
S_term_DSP Tile_X7Y15_S_term_DSP (
    .S1END(Tile_X7Y14_S1BEG),
    .S2MID(Tile_X7Y14_S2BEG),
    .S2END(Tile_X7Y14_S2BEGb),
    .S4END(Tile_X7Y14_S4BEG),
    .SS4END(Tile_X7Y14_SS4BEG),
    .N1BEG(Tile_X7Y15_N1BEG),
    .N2BEG(Tile_X7Y15_N2BEG),
    .N2BEGb(Tile_X7Y15_N2BEGb),
    .N4BEG(Tile_X7Y15_N4BEG),
    .NN4BEG(Tile_X7Y15_NN4BEG),
    .UserCLK(UserCLK),
    .UserCLKo(Tile_X7Y15_UserCLKo),
    .FrameData(Tile_X6Y15_FrameData_O),
    .FrameData_O(Tile_X7Y15_FrameData_O),
    .FrameStrobe(Column_X7_FrameStrobe),
    .FrameStrobe_O(Tile_X7Y15_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
S_CPU_IF Tile_X8Y15_S_CPU_IF (
    .S1END(Tile_X8Y14_S1BEG),
    .S2MID(Tile_X8Y14_S2BEG),
    .S2END(Tile_X8Y14_S2BEGb),
    .S4END(Tile_X8Y14_S4BEG),
    .SS4END(Tile_X8Y14_SS4BEG),
    .N1BEG(Tile_X8Y15_N1BEG),
    .N2BEG(Tile_X8Y15_N2BEG),
    .N2BEGb(Tile_X8Y15_N2BEGb),
    .N4BEG(Tile_X8Y15_N4BEG),
    .NN4BEG(Tile_X8Y15_NN4BEG),
    .Co(Tile_X8Y15_Co),
    .O_top0(Tile_X8Y15_O_top0),
    .O_top1(Tile_X8Y15_O_top1),
    .O_top2(Tile_X8Y15_O_top2),
    .O_top3(Tile_X8Y15_O_top3),
    .O_top4(Tile_X8Y15_O_top4),
    .O_top5(Tile_X8Y15_O_top5),
    .O_top6(Tile_X8Y15_O_top6),
    .O_top7(Tile_X8Y15_O_top7),
    .O_top8(Tile_X8Y15_O_top8),
    .O_top9(Tile_X8Y15_O_top9),
    .O_top10(Tile_X8Y15_O_top10),
    .O_top11(Tile_X8Y15_O_top11),
    .O_top12(Tile_X8Y15_O_top12),
    .O_top13(Tile_X8Y15_O_top13),
    .O_top14(Tile_X8Y15_O_top14),
    .O_top15(Tile_X8Y15_O_top15),
    .I_top0(Tile_X8Y15_I_top0),
    .I_top1(Tile_X8Y15_I_top1),
    .I_top2(Tile_X8Y15_I_top2),
    .I_top3(Tile_X8Y15_I_top3),
    .I_top4(Tile_X8Y15_I_top4),
    .I_top5(Tile_X8Y15_I_top5),
    .I_top6(Tile_X8Y15_I_top6),
    .I_top7(Tile_X8Y15_I_top7),
    .I_top8(Tile_X8Y15_I_top8),
    .I_top9(Tile_X8Y15_I_top9),
    .I_top10(Tile_X8Y15_I_top10),
    .I_top11(Tile_X8Y15_I_top11),
    .I_top12(Tile_X8Y15_I_top12),
    .I_top13(Tile_X8Y15_I_top13),
    .I_top14(Tile_X8Y15_I_top14),
    .I_top15(Tile_X8Y15_I_top15),
    .UserCLK(UserCLK),
    .UserCLKo(Tile_X8Y15_UserCLKo),
    .FrameData(Tile_X7Y15_FrameData_O),
    .FrameData_O(Tile_X8Y15_FrameData_O),
    .FrameStrobe(Column_X8_FrameStrobe),
    .FrameStrobe_O(Tile_X8Y15_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
S_CPU_IF Tile_X9Y15_S_CPU_IF (
    .S1END(Tile_X9Y14_S1BEG),
    .S2MID(Tile_X9Y14_S2BEG),
    .S2END(Tile_X9Y14_S2BEGb),
    .S4END(Tile_X9Y14_S4BEG),
    .SS4END(Tile_X9Y14_SS4BEG),
    .N1BEG(Tile_X9Y15_N1BEG),
    .N2BEG(Tile_X9Y15_N2BEG),
    .N2BEGb(Tile_X9Y15_N2BEGb),
    .N4BEG(Tile_X9Y15_N4BEG),
    .NN4BEG(Tile_X9Y15_NN4BEG),
    .Co(Tile_X9Y15_Co),
    .O_top0(Tile_X9Y15_O_top0),
    .O_top1(Tile_X9Y15_O_top1),
    .O_top2(Tile_X9Y15_O_top2),
    .O_top3(Tile_X9Y15_O_top3),
    .O_top4(Tile_X9Y15_O_top4),
    .O_top5(Tile_X9Y15_O_top5),
    .O_top6(Tile_X9Y15_O_top6),
    .O_top7(Tile_X9Y15_O_top7),
    .O_top8(Tile_X9Y15_O_top8),
    .O_top9(Tile_X9Y15_O_top9),
    .O_top10(Tile_X9Y15_O_top10),
    .O_top11(Tile_X9Y15_O_top11),
    .O_top12(Tile_X9Y15_O_top12),
    .O_top13(Tile_X9Y15_O_top13),
    .O_top14(Tile_X9Y15_O_top14),
    .O_top15(Tile_X9Y15_O_top15),
    .I_top0(Tile_X9Y15_I_top0),
    .I_top1(Tile_X9Y15_I_top1),
    .I_top2(Tile_X9Y15_I_top2),
    .I_top3(Tile_X9Y15_I_top3),
    .I_top4(Tile_X9Y15_I_top4),
    .I_top5(Tile_X9Y15_I_top5),
    .I_top6(Tile_X9Y15_I_top6),
    .I_top7(Tile_X9Y15_I_top7),
    .I_top8(Tile_X9Y15_I_top8),
    .I_top9(Tile_X9Y15_I_top9),
    .I_top10(Tile_X9Y15_I_top10),
    .I_top11(Tile_X9Y15_I_top11),
    .I_top12(Tile_X9Y15_I_top12),
    .I_top13(Tile_X9Y15_I_top13),
    .I_top14(Tile_X9Y15_I_top14),
    .I_top15(Tile_X9Y15_I_top15),
    .UserCLK(UserCLK),
    .UserCLKo(Tile_X9Y15_UserCLKo),
    .FrameData(Tile_X8Y15_FrameData_O),
    .FrameData_O(Tile_X9Y15_FrameData_O),
    .FrameStrobe(Column_X9_FrameStrobe),
    .FrameStrobe_O(Tile_X9Y15_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
S_term_IHP_SRAM Tile_X10Y15_S_term_IHP_SRAM (
    .S1END(Tile_X10Y14_S1BEG),
    .S2MID(Tile_X10Y14_S2BEG),
    .S2END(Tile_X10Y14_S2BEGb),
    .S4END(Tile_X10Y14_S4BEG),
    .N1BEG(Tile_X10Y15_N1BEG),
    .N2BEG(Tile_X10Y15_N2BEG),
    .N2BEGb(Tile_X10Y15_N2BEGb),
    .N4BEG(Tile_X10Y15_N4BEG),
    .UserCLK(UserCLK),
    .UserCLKo(Tile_X10Y15_UserCLKo),
    .FrameData(Tile_X9Y15_FrameData_O),
    .FrameData_O(Tile_X10Y15_FrameData_O),
    .FrameStrobe(Column_X10_FrameStrobe),
    .FrameStrobe_O(Tile_X10Y15_FrameStrobe_O)
);

endmodule