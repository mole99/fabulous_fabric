magic
tech sky130A
magscale 1 2
timestamp 1740405677
<< metal1 >>
rect 481910 696328 481916 696380
rect 481968 696368 481974 696380
rect 482554 696368 482560 696380
rect 481968 696340 482560 696368
rect 481968 696328 481974 696340
rect 482554 696328 482560 696340
rect 482612 696328 482618 696380
rect 482554 696192 482560 696244
rect 482612 696232 482618 696244
rect 482922 696232 482928 696244
rect 482612 696204 482928 696232
rect 482612 696192 482618 696204
rect 482922 696192 482928 696204
rect 482980 696192 482986 696244
rect 479978 685040 479984 685092
rect 480036 685080 480042 685092
rect 480254 685080 480260 685092
rect 480036 685052 480260 685080
rect 480036 685040 480042 685052
rect 480254 685040 480260 685052
rect 480312 685040 480318 685092
rect 7650 17212 7656 17264
rect 7708 17252 7714 17264
rect 7708 17224 15102 17252
rect 7708 17212 7714 17224
rect 15074 17196 15102 17224
rect 9214 17144 9220 17196
rect 9272 17184 9278 17196
rect 14596 17184 14602 17196
rect 9272 17156 14602 17184
rect 9272 17144 9278 17156
rect 14596 17144 14602 17156
rect 14654 17144 14660 17196
rect 15056 17144 15062 17196
rect 15114 17144 15120 17196
rect 6178 17076 6184 17128
rect 6236 17116 6242 17128
rect 11376 17116 11382 17128
rect 6236 17088 11382 17116
rect 6236 17076 6242 17088
rect 11376 17076 11382 17088
rect 11434 17076 11440 17128
rect 7558 17008 7564 17060
rect 7616 17048 7622 17060
rect 20116 17048 20122 17060
rect 7616 17020 20122 17048
rect 7616 17008 7622 17020
rect 20116 17008 20122 17020
rect 20174 17008 20180 17060
rect 8846 16940 8852 16992
rect 8904 16980 8910 16992
rect 18322 16980 18328 16992
rect 8904 16952 18328 16980
rect 8904 16940 8910 16952
rect 18322 16940 18328 16952
rect 18380 16940 18386 16992
rect 7374 16872 7380 16924
rect 7432 16912 7438 16924
rect 19242 16912 19248 16924
rect 7432 16884 19248 16912
rect 7432 16872 7438 16884
rect 19242 16872 19248 16884
rect 19300 16872 19306 16924
rect 8478 16804 8484 16856
rect 8536 16844 8542 16856
rect 19702 16844 19708 16856
rect 8536 16816 19708 16844
rect 8536 16804 8542 16816
rect 19702 16804 19708 16816
rect 19760 16804 19766 16856
rect 8110 16532 8116 16584
rect 8168 16572 8174 16584
rect 16482 16572 16488 16584
rect 8168 16544 16488 16572
rect 8168 16532 8174 16544
rect 16482 16532 16488 16544
rect 16540 16532 16546 16584
<< via1 >>
rect 481916 696328 481968 696380
rect 482560 696328 482612 696380
rect 482560 696192 482612 696244
rect 482928 696192 482980 696244
rect 479984 685040 480036 685092
rect 480260 685040 480312 685092
rect 7656 17212 7708 17264
rect 9220 17144 9272 17196
rect 14602 17144 14654 17196
rect 15062 17144 15114 17196
rect 6184 17076 6236 17128
rect 11382 17076 11434 17128
rect 7564 17008 7616 17060
rect 20122 17008 20174 17060
rect 8852 16940 8904 16992
rect 18328 16940 18380 16992
rect 7380 16872 7432 16924
rect 19248 16872 19300 16924
rect 8484 16804 8536 16856
rect 19708 16804 19760 16856
rect 8116 16532 8168 16584
rect 16488 16532 16540 16584
<< metal2 >>
rect 7746 755834 7802 756500
rect 8390 755834 8446 756500
rect 7746 755806 7880 755834
rect 7746 755700 7802 755806
rect 7852 741074 7880 755806
rect 8312 755806 8446 755834
rect 8312 745521 8340 755806
rect 8390 755700 8446 755806
rect 9034 755834 9090 756500
rect 9678 755834 9734 756500
rect 10322 755834 10378 756500
rect 10966 755834 11022 756500
rect 9034 755806 9168 755834
rect 9034 755700 9090 755806
rect 9140 747153 9168 755806
rect 9678 755806 9812 755834
rect 9678 755700 9734 755806
rect 9126 747144 9182 747153
rect 9126 747079 9182 747088
rect 9784 746337 9812 755806
rect 10322 755806 10456 755834
rect 10322 755700 10378 755806
rect 9770 746328 9826 746337
rect 9770 746263 9826 746272
rect 8298 745512 8354 745521
rect 8298 745447 8354 745456
rect 10428 743073 10456 755806
rect 10888 755806 11022 755834
rect 10888 750734 10916 755806
rect 10966 755700 11022 755806
rect 11610 755834 11666 756500
rect 12254 755834 12310 756500
rect 11610 755806 11744 755834
rect 11610 755700 11666 755806
rect 10888 750706 11008 750734
rect 10414 743064 10470 743073
rect 10414 742999 10470 743008
rect 7760 741046 7880 741074
rect 7760 738721 7788 741046
rect 10980 739265 11008 750706
rect 11716 743889 11744 755806
rect 12176 755806 12310 755834
rect 11702 743880 11758 743889
rect 11702 743815 11758 743824
rect 12176 741985 12204 755806
rect 12254 755700 12310 755806
rect 12898 755834 12954 756500
rect 13542 755834 13598 756500
rect 12898 755806 13032 755834
rect 12898 755700 12954 755806
rect 13004 746609 13032 755806
rect 13464 755806 13598 755834
rect 12990 746600 13046 746609
rect 12990 746535 13046 746544
rect 13464 744977 13492 755806
rect 13542 755700 13598 755806
rect 14186 755834 14242 756500
rect 14830 755834 14886 756500
rect 14186 755806 14320 755834
rect 14186 755700 14242 755806
rect 13450 744968 13506 744977
rect 13450 744903 13506 744912
rect 12162 741976 12218 741985
rect 12162 741911 12218 741920
rect 14292 741074 14320 755806
rect 14752 755806 14886 755834
rect 14752 742801 14780 755806
rect 14830 755700 14886 755806
rect 15474 755834 15530 756500
rect 16118 755834 16174 756500
rect 15474 755806 15608 755834
rect 15474 755700 15530 755806
rect 14738 742792 14794 742801
rect 14738 742727 14794 742736
rect 15580 741713 15608 755806
rect 16040 755806 16174 755834
rect 16040 750734 16068 755806
rect 16118 755700 16174 755806
rect 16762 755834 16818 756500
rect 17406 755834 17462 756500
rect 16762 755806 16896 755834
rect 16762 755700 16818 755806
rect 16040 750706 16160 750734
rect 15566 741704 15622 741713
rect 15566 741639 15622 741648
rect 14200 741046 14320 741074
rect 10966 739256 11022 739265
rect 10966 739191 11022 739200
rect 14200 738993 14228 741046
rect 16132 740625 16160 750706
rect 16868 741074 16896 755806
rect 17328 755806 17462 755834
rect 17328 743617 17356 755806
rect 17406 755700 17462 755806
rect 18050 755834 18106 756500
rect 18694 755834 18750 756500
rect 18050 755806 18184 755834
rect 18050 755700 18106 755806
rect 18156 746065 18184 755806
rect 18616 755806 18750 755834
rect 18142 746056 18198 746065
rect 18142 745991 18198 746000
rect 18616 745249 18644 755806
rect 18694 755700 18750 755806
rect 19338 755834 19394 756500
rect 19982 755834 20038 756500
rect 20626 755834 20682 756500
rect 21270 755834 21326 756500
rect 19338 755806 19472 755834
rect 19338 755700 19394 755806
rect 18602 745240 18658 745249
rect 18602 745175 18658 745184
rect 19444 744161 19472 755806
rect 19904 755806 20038 755834
rect 19430 744152 19486 744161
rect 19430 744087 19486 744096
rect 17314 743608 17370 743617
rect 17314 743543 17370 743552
rect 19904 742257 19932 755806
rect 19982 755700 20038 755806
rect 20548 755806 20682 755834
rect 20442 755712 20498 755721
rect 20442 755647 20498 755656
rect 20074 755440 20130 755449
rect 20074 755375 20130 755384
rect 19890 742248 19946 742257
rect 19890 742183 19946 742192
rect 16776 741046 16896 741074
rect 16118 740616 16174 740625
rect 16118 740551 16174 740560
rect 16776 739809 16804 741046
rect 20088 740353 20116 755375
rect 20258 754896 20314 754905
rect 20258 754831 20314 754840
rect 20166 749592 20222 749601
rect 20166 749527 20222 749536
rect 20074 740344 20130 740353
rect 20074 740279 20130 740288
rect 16762 739800 16818 739809
rect 16762 739735 16818 739744
rect 20180 739537 20208 749527
rect 20272 744705 20300 754831
rect 20350 754080 20406 754089
rect 20350 754015 20406 754024
rect 20258 744696 20314 744705
rect 20258 744631 20314 744640
rect 20364 741169 20392 754015
rect 20456 753114 20484 755647
rect 20548 753250 20576 755806
rect 20626 755700 20682 755806
rect 21192 755806 21326 755834
rect 20548 753222 20668 753250
rect 20456 753086 20576 753114
rect 20442 752720 20498 752729
rect 20442 752655 20498 752664
rect 20350 741160 20406 741169
rect 20350 741095 20406 741104
rect 20456 740897 20484 752655
rect 20548 745793 20576 753086
rect 20534 745784 20590 745793
rect 20534 745719 20590 745728
rect 20640 742529 20668 753222
rect 21192 749465 21220 755806
rect 21270 755700 21326 755806
rect 21914 755834 21970 756500
rect 22558 755834 22614 756500
rect 23202 755834 23258 756500
rect 23846 755834 23902 756500
rect 24490 755834 24546 756500
rect 25134 755834 25190 756500
rect 21914 755806 22048 755834
rect 21914 755700 21970 755806
rect 21454 753536 21510 753545
rect 21454 753471 21510 753480
rect 21178 749456 21234 749465
rect 21178 749391 21234 749400
rect 21086 744446 21142 744455
rect 21468 744432 21496 753471
rect 22020 749601 22048 755806
rect 22296 755806 22614 755834
rect 22296 753545 22324 755806
rect 22558 755700 22614 755806
rect 22940 755806 23258 755834
rect 22282 753536 22338 753545
rect 22282 753471 22338 753480
rect 22006 749592 22062 749601
rect 22006 749527 22062 749536
rect 22940 748476 22968 755806
rect 23202 755700 23258 755806
rect 23584 755806 23902 755834
rect 23584 754905 23612 755806
rect 23846 755700 23902 755806
rect 24044 755806 24546 755834
rect 23570 754896 23626 754905
rect 23570 754831 23626 754840
rect 24044 748476 24072 755806
rect 24490 755700 24546 755806
rect 25056 755806 25190 755834
rect 25056 748762 25084 755806
rect 25134 755700 25190 755806
rect 25778 755834 25834 756500
rect 26422 755834 26478 756500
rect 25778 755806 25912 755834
rect 25778 755700 25834 755806
rect 25056 748734 25174 748762
rect 25146 748476 25174 748734
rect 25884 748649 25912 755806
rect 26252 755806 26478 755834
rect 25870 748640 25926 748649
rect 25870 748575 25926 748584
rect 26252 748476 26280 755806
rect 26422 755700 26478 755806
rect 26790 755848 26846 755857
rect 27066 755834 27122 756500
rect 27710 755834 27766 756500
rect 28354 755834 28410 756500
rect 28998 755834 29054 756500
rect 29642 755834 29698 756500
rect 30286 755834 30342 756500
rect 30930 755834 30986 756500
rect 31574 755834 31630 756500
rect 32218 755834 32274 756500
rect 32862 755834 32918 756500
rect 33506 755834 33562 756500
rect 34150 755834 34206 756500
rect 34794 755834 34850 756500
rect 35438 755834 35494 756500
rect 26846 755806 27122 755834
rect 26790 755783 26846 755792
rect 27066 755700 27122 755806
rect 27356 755806 27766 755834
rect 27356 748476 27384 755806
rect 27710 755700 27766 755806
rect 28000 755806 28410 755834
rect 28000 755041 28028 755806
rect 28354 755700 28410 755806
rect 28460 755806 29054 755834
rect 27986 755032 28042 755041
rect 27986 754967 28042 754976
rect 28460 748476 28488 755806
rect 28998 755700 29054 755806
rect 29564 755806 29698 755834
rect 29564 748476 29592 755806
rect 29642 755700 29698 755806
rect 30024 755806 30342 755834
rect 30024 752729 30052 755806
rect 30286 755700 30342 755806
rect 30668 755806 30986 755834
rect 30010 752720 30066 752729
rect 30010 752655 30066 752664
rect 30668 748476 30696 755806
rect 30930 755700 30986 755806
rect 31312 755806 31630 755834
rect 31312 755721 31340 755806
rect 31298 755712 31354 755721
rect 31574 755700 31630 755806
rect 31772 755806 32274 755834
rect 31298 755647 31354 755656
rect 31772 748476 31800 755806
rect 32218 755700 32274 755806
rect 32784 755806 32918 755834
rect 32784 748762 32812 755806
rect 32862 755700 32918 755806
rect 33152 755806 33562 755834
rect 33152 754089 33180 755806
rect 33506 755700 33562 755806
rect 33980 755806 34206 755834
rect 33138 754080 33194 754089
rect 33138 754015 33194 754024
rect 32784 748734 32902 748762
rect 32874 748476 32902 748734
rect 33980 748476 34008 755806
rect 34150 755700 34206 755806
rect 34532 755806 34850 755834
rect 34532 755449 34560 755806
rect 34794 755700 34850 755806
rect 35084 755806 35494 755834
rect 34518 755440 34574 755449
rect 34518 755375 34574 755384
rect 35084 748476 35112 755806
rect 35438 755700 35494 755806
rect 36082 755834 36138 756500
rect 37370 755834 37426 756500
rect 36082 755806 36216 755834
rect 36082 755700 36138 755806
rect 36188 748476 36216 755806
rect 37292 755806 37426 755834
rect 37292 748476 37320 755806
rect 37370 755700 37426 755806
rect 63774 755834 63830 756500
rect 65062 755834 65118 756500
rect 66350 755834 66406 756500
rect 63774 755806 64000 755834
rect 63774 755700 63830 755806
rect 63972 748762 64000 755806
rect 63938 748734 64000 748762
rect 64984 755806 65118 755834
rect 64984 748762 65012 755806
rect 65062 755700 65118 755806
rect 66180 755806 66406 755834
rect 66180 748762 66208 755806
rect 66350 755700 66406 755806
rect 66994 755834 67050 756500
rect 68282 755834 68338 756500
rect 69570 755834 69626 756500
rect 70858 755834 70914 756500
rect 66994 755806 67312 755834
rect 66994 755700 67050 755806
rect 67284 748762 67312 755806
rect 68282 755806 68416 755834
rect 68282 755700 68338 755806
rect 68388 748762 68416 755806
rect 69492 755806 69626 755834
rect 69492 748762 69520 755806
rect 69570 755700 69626 755806
rect 70596 755806 70914 755834
rect 70596 748762 70624 755806
rect 70858 755700 70914 755806
rect 71502 755834 71558 756500
rect 72790 755834 72846 756500
rect 74078 755834 74134 756500
rect 71502 755806 71728 755834
rect 71502 755700 71558 755806
rect 71700 748762 71728 755806
rect 64984 748734 65058 748762
rect 63938 748476 63966 748734
rect 65030 748476 65058 748734
rect 66146 748734 66208 748762
rect 67250 748734 67312 748762
rect 68354 748734 68416 748762
rect 69458 748734 69520 748762
rect 70562 748734 70624 748762
rect 71666 748734 71728 748762
rect 72712 755806 72846 755834
rect 72712 748762 72740 755806
rect 72790 755700 72846 755806
rect 73908 755806 74134 755834
rect 73908 748762 73936 755806
rect 74078 755700 74134 755806
rect 74722 755834 74778 756500
rect 76010 755834 76066 756500
rect 77298 755834 77354 756500
rect 78586 755834 78642 756500
rect 153934 755834 153990 756500
rect 155222 755834 155278 756500
rect 155866 755834 155922 756500
rect 74722 755806 75040 755834
rect 74722 755700 74778 755806
rect 75012 748762 75040 755806
rect 76010 755806 76144 755834
rect 76010 755700 76066 755806
rect 76116 748762 76144 755806
rect 77220 755806 77354 755834
rect 77220 748762 77248 755806
rect 77298 755700 77354 755806
rect 78324 755806 78642 755834
rect 78324 748762 78352 755806
rect 78586 755700 78642 755806
rect 153856 755806 153990 755834
rect 72712 748734 72786 748762
rect 66146 748476 66174 748734
rect 67250 748476 67278 748734
rect 68354 748476 68382 748734
rect 69458 748476 69486 748734
rect 70562 748476 70590 748734
rect 71666 748476 71694 748734
rect 72758 748476 72786 748734
rect 73874 748734 73936 748762
rect 74978 748734 75040 748762
rect 76082 748734 76144 748762
rect 77186 748734 77248 748762
rect 78290 748734 78352 748762
rect 153856 748762 153884 755806
rect 153934 755700 153990 755806
rect 155052 755806 155278 755834
rect 153856 748734 153966 748762
rect 73874 748476 73902 748734
rect 74978 748476 75006 748734
rect 76082 748476 76110 748734
rect 77186 748476 77214 748734
rect 78290 748476 78318 748734
rect 153938 748476 153966 748734
rect 155052 748476 155080 755806
rect 155222 755700 155278 755806
rect 155788 755806 155922 755834
rect 155788 750734 155816 755806
rect 155866 755700 155922 755806
rect 157154 755834 157210 756500
rect 158442 755834 158498 756500
rect 159730 755834 159786 756500
rect 157154 755806 157288 755834
rect 157154 755700 157210 755806
rect 155788 750706 156092 750734
rect 156064 748762 156092 750706
rect 156064 748734 156174 748762
rect 156146 748476 156174 748734
rect 157260 748476 157288 755806
rect 158364 755806 158498 755834
rect 158364 748476 158392 755806
rect 158442 755700 158498 755806
rect 159468 755806 159786 755834
rect 159468 748476 159496 755806
rect 159730 755700 159786 755806
rect 160374 755834 160430 756500
rect 161662 755834 161718 756500
rect 162950 755834 163006 756500
rect 160374 755806 160600 755834
rect 160374 755700 160430 755806
rect 160572 748476 160600 755806
rect 161584 755806 161718 755834
rect 161584 748762 161612 755806
rect 161662 755700 161718 755806
rect 162780 755806 163006 755834
rect 161584 748734 161694 748762
rect 161666 748476 161694 748734
rect 162780 748476 162808 755806
rect 162950 755700 163006 755806
rect 163594 755834 163650 756500
rect 164882 755834 164938 756500
rect 166170 755834 166226 756500
rect 167458 755834 167514 756500
rect 163594 755806 163912 755834
rect 163594 755700 163650 755806
rect 163884 748476 163912 755806
rect 164882 755806 165016 755834
rect 164882 755700 164938 755806
rect 164988 748476 165016 755806
rect 166092 755806 166226 755834
rect 166092 748476 166120 755806
rect 166170 755700 166226 755806
rect 167196 755806 167514 755834
rect 167196 748476 167224 755806
rect 167458 755700 167514 755806
rect 168102 755834 168158 756500
rect 195150 755834 195206 756500
rect 168102 755806 168328 755834
rect 168102 755700 168158 755806
rect 168300 748476 168328 755806
rect 194980 755806 195206 755834
rect 194980 748762 195008 755806
rect 195150 755700 195206 755806
rect 195794 755834 195850 756500
rect 197082 755834 197138 756500
rect 198370 755834 198426 756500
rect 199658 755834 199714 756500
rect 195794 755806 195928 755834
rect 195794 755700 195850 755806
rect 195900 750734 195928 755806
rect 197082 755806 197216 755834
rect 197082 755700 197138 755806
rect 195900 750706 196020 750734
rect 194938 748734 195008 748762
rect 195992 748762 196020 750706
rect 197188 748762 197216 755806
rect 198292 755806 198426 755834
rect 198292 748762 198320 755806
rect 198370 755700 198426 755806
rect 199396 755806 199714 755834
rect 199396 748762 199424 755806
rect 199658 755700 199714 755806
rect 200302 755834 200358 756500
rect 201590 755834 201646 756500
rect 202878 755834 202934 756500
rect 200302 755806 200528 755834
rect 200302 755700 200358 755806
rect 200500 748762 200528 755806
rect 195992 748734 196066 748762
rect 194938 748476 194966 748734
rect 196038 748476 196066 748734
rect 197146 748734 197216 748762
rect 198250 748734 198320 748762
rect 199354 748734 199424 748762
rect 200458 748734 200528 748762
rect 201512 755806 201646 755834
rect 201512 748762 201540 755806
rect 201590 755700 201646 755806
rect 202708 755806 202934 755834
rect 202708 748762 202736 755806
rect 202878 755700 202934 755806
rect 203522 755834 203578 756500
rect 204810 755834 204866 756500
rect 206098 755834 206154 756500
rect 207386 755834 207442 756500
rect 203522 755806 203840 755834
rect 203522 755700 203578 755806
rect 203812 748762 203840 755806
rect 204810 755806 204944 755834
rect 204810 755700 204866 755806
rect 204916 748762 204944 755806
rect 206020 755806 206154 755834
rect 206020 748762 206048 755806
rect 206098 755700 206154 755806
rect 207124 755806 207442 755834
rect 207124 748762 207152 755806
rect 207386 755700 207442 755806
rect 208030 755834 208086 756500
rect 209318 755834 209374 756500
rect 208030 755806 208256 755834
rect 208030 755700 208086 755806
rect 208228 748762 208256 755806
rect 201512 748734 201586 748762
rect 197146 748476 197174 748734
rect 198250 748476 198278 748734
rect 199354 748476 199382 748734
rect 200458 748476 200486 748734
rect 201558 748476 201586 748734
rect 202666 748734 202736 748762
rect 203770 748734 203840 748762
rect 204874 748734 204944 748762
rect 205978 748734 206048 748762
rect 207082 748734 207152 748762
rect 208186 748734 208256 748762
rect 209240 755806 209374 755834
rect 209240 748762 209268 755806
rect 209318 755700 209374 755806
rect 235722 755834 235778 756500
rect 237010 755834 237066 756500
rect 238298 755834 238354 756500
rect 235722 755806 235948 755834
rect 235722 755700 235778 755806
rect 235920 748762 235948 755806
rect 237010 755806 237144 755834
rect 237010 755700 237066 755806
rect 237116 748762 237144 755806
rect 238220 755806 238354 755834
rect 238220 748762 238248 755806
rect 238298 755700 238354 755806
rect 238942 755834 238998 756500
rect 240230 755834 240286 756500
rect 241518 755834 241574 756500
rect 242806 755834 242862 756500
rect 238942 755806 239352 755834
rect 238942 755700 238998 755806
rect 239324 748762 239352 755806
rect 240230 755806 240456 755834
rect 240230 755700 240286 755806
rect 240428 748762 240456 755806
rect 209240 748734 209314 748762
rect 235920 748734 235966 748762
rect 202666 748476 202694 748734
rect 203770 748476 203798 748734
rect 204874 748476 204902 748734
rect 205978 748476 206006 748734
rect 207082 748476 207110 748734
rect 208186 748476 208214 748734
rect 209286 748476 209314 748734
rect 235938 748476 235966 748734
rect 237042 748734 237144 748762
rect 238146 748734 238248 748762
rect 239250 748734 239352 748762
rect 240354 748734 240456 748762
rect 241440 755806 241574 755834
rect 241440 748762 241468 755806
rect 241518 755700 241574 755806
rect 242636 755806 242862 755834
rect 242636 748762 242664 755806
rect 242806 755700 242862 755806
rect 243450 755834 243506 756500
rect 244738 755834 244794 756500
rect 246026 755834 246082 756500
rect 243450 755806 243768 755834
rect 243450 755700 243506 755806
rect 243740 748762 243768 755806
rect 244738 755806 244872 755834
rect 244738 755700 244794 755806
rect 244844 748762 244872 755806
rect 245948 755806 246082 755834
rect 245948 748762 245976 755806
rect 246026 755700 246082 755806
rect 246670 755834 246726 756500
rect 247958 755834 248014 756500
rect 249246 755834 249302 756500
rect 250534 755834 250590 756500
rect 322018 755834 322074 756500
rect 323306 755834 323362 756500
rect 246670 755806 246988 755834
rect 246670 755700 246726 755806
rect 241440 748734 241486 748762
rect 237042 748476 237070 748734
rect 238146 748476 238174 748734
rect 239250 748476 239278 748734
rect 240354 748476 240382 748734
rect 241458 748476 241486 748734
rect 242562 748734 242664 748762
rect 243666 748734 243768 748762
rect 244770 748734 244872 748762
rect 245874 748734 245976 748762
rect 246960 748762 246988 755806
rect 247958 755806 248184 755834
rect 247958 755700 248014 755806
rect 248156 748762 248184 755806
rect 246960 748734 247006 748762
rect 242562 748476 242590 748734
rect 243666 748476 243694 748734
rect 244770 748476 244798 748734
rect 245874 748476 245902 748734
rect 246978 748476 247006 748734
rect 248082 748734 248184 748762
rect 249168 755806 249302 755834
rect 249168 748762 249196 755806
rect 249246 755700 249302 755806
rect 250364 755806 250590 755834
rect 250364 748762 250392 755806
rect 250534 755700 250590 755806
rect 321940 755806 322074 755834
rect 249168 748734 249214 748762
rect 248082 748476 248110 748734
rect 249186 748476 249214 748734
rect 250290 748734 250392 748762
rect 250290 748476 250318 748734
rect 321940 748476 321968 755806
rect 322018 755700 322074 755806
rect 323044 755806 323362 755834
rect 323044 748476 323072 755806
rect 323306 755700 323362 755806
rect 323950 755834 324006 756500
rect 325238 755834 325294 756500
rect 326526 755834 326582 756500
rect 323950 755806 324176 755834
rect 323950 755700 324006 755806
rect 324148 748476 324176 755806
rect 325160 755806 325294 755834
rect 325160 748762 325188 755806
rect 325238 755700 325294 755806
rect 326356 755806 326582 755834
rect 325160 748734 325278 748762
rect 325250 748476 325278 748734
rect 326356 748476 326384 755806
rect 326526 755700 326582 755806
rect 327170 755834 327226 756500
rect 328458 755834 328514 756500
rect 329746 755834 329802 756500
rect 331034 755834 331090 756500
rect 327170 755806 327488 755834
rect 327170 755700 327226 755806
rect 327460 748476 327488 755806
rect 328458 755806 328592 755834
rect 328458 755700 328514 755806
rect 328564 748476 328592 755806
rect 329668 755806 329802 755834
rect 329668 748476 329696 755806
rect 329746 755700 329802 755806
rect 330772 755806 331090 755834
rect 330772 748476 330800 755806
rect 331034 755700 331090 755806
rect 331678 755834 331734 756500
rect 332966 755834 333022 756500
rect 334254 755834 334310 756500
rect 331678 755806 331904 755834
rect 331678 755700 331734 755806
rect 331876 748476 331904 755806
rect 332888 755806 333022 755834
rect 332888 748762 332916 755806
rect 332966 755700 333022 755806
rect 334084 755806 334310 755834
rect 332888 748734 333006 748762
rect 332978 748476 333006 748734
rect 334084 748476 334112 755806
rect 334254 755700 334310 755806
rect 334898 755834 334954 756500
rect 336186 755834 336242 756500
rect 363234 755834 363290 756500
rect 334898 755806 335216 755834
rect 334898 755700 334954 755806
rect 335188 748476 335216 755806
rect 336186 755806 336320 755834
rect 336186 755700 336242 755806
rect 336292 748476 336320 755806
rect 362972 755806 363290 755834
rect 362972 748762 363000 755806
rect 363234 755700 363290 755806
rect 363878 755834 363934 756500
rect 365166 755834 365222 756500
rect 366454 755834 366510 756500
rect 363878 755806 364104 755834
rect 363878 755700 363934 755806
rect 364076 748762 364104 755806
rect 362938 748734 363000 748762
rect 364042 748734 364104 748762
rect 365088 755806 365222 755834
rect 365088 748762 365116 755806
rect 365166 755700 365222 755806
rect 366284 755806 366510 755834
rect 366284 748762 366312 755806
rect 366454 755700 366510 755806
rect 367098 755834 367154 756500
rect 368386 755834 368442 756500
rect 369674 755834 369730 756500
rect 370962 755834 371018 756500
rect 367098 755806 367416 755834
rect 367098 755700 367154 755806
rect 367388 748762 367416 755806
rect 368308 755806 368442 755834
rect 368308 750734 368336 755806
rect 368386 755700 368442 755806
rect 369596 755806 369730 755834
rect 368308 750706 368520 750734
rect 368492 748762 368520 750706
rect 369596 748762 369624 755806
rect 369674 755700 369730 755806
rect 370700 755806 371018 755834
rect 370700 748762 370728 755806
rect 370962 755700 371018 755806
rect 371606 755834 371662 756500
rect 372894 755834 372950 756500
rect 374182 755834 374238 756500
rect 371606 755806 371832 755834
rect 371606 755700 371662 755806
rect 371804 748762 371832 755806
rect 365088 748734 365162 748762
rect 362938 748476 362966 748734
rect 364042 748476 364070 748734
rect 365134 748476 365162 748734
rect 366250 748734 366312 748762
rect 367354 748734 367416 748762
rect 368458 748734 368520 748762
rect 369562 748734 369624 748762
rect 370666 748734 370728 748762
rect 371770 748734 371832 748762
rect 372816 755806 372950 755834
rect 372816 748762 372844 755806
rect 372894 755700 372950 755806
rect 374012 755806 374238 755834
rect 374012 748762 374040 755806
rect 374182 755700 374238 755806
rect 374826 755834 374882 756500
rect 376114 755834 376170 756500
rect 377402 755834 377458 756500
rect 374826 755806 375144 755834
rect 374826 755700 374882 755806
rect 375116 748762 375144 755806
rect 376114 755806 376248 755834
rect 376114 755700 376170 755806
rect 376220 748762 376248 755806
rect 377324 755806 377458 755834
rect 377324 748762 377352 755806
rect 377402 755700 377458 755806
rect 403806 755834 403862 756500
rect 405094 755834 405150 756500
rect 406382 755834 406438 756500
rect 407026 755834 407082 756500
rect 403806 755806 404032 755834
rect 403806 755700 403862 755806
rect 404004 748762 404032 755806
rect 372816 748734 372890 748762
rect 366250 748476 366278 748734
rect 367354 748476 367382 748734
rect 368458 748476 368486 748734
rect 369562 748476 369590 748734
rect 370666 748476 370694 748734
rect 371770 748476 371798 748734
rect 372862 748476 372890 748734
rect 373978 748734 374040 748762
rect 375082 748734 375144 748762
rect 376186 748734 376248 748762
rect 377290 748734 377352 748762
rect 403938 748734 404032 748762
rect 405016 755806 405150 755834
rect 405016 748762 405044 755806
rect 405094 755700 405150 755806
rect 406212 755806 406438 755834
rect 406212 748762 406240 755806
rect 406382 755700 406438 755806
rect 406948 755806 407082 755834
rect 406948 750734 406976 755806
rect 407026 755700 407082 755806
rect 408314 755834 408370 756500
rect 409602 755834 409658 756500
rect 408314 755806 408448 755834
rect 408314 755700 408370 755806
rect 406948 750706 407252 750734
rect 405016 748734 405070 748762
rect 373978 748476 374006 748734
rect 375082 748476 375110 748734
rect 376186 748476 376214 748734
rect 377290 748476 377318 748734
rect 403938 748476 403966 748734
rect 405042 748476 405070 748734
rect 406146 748734 406240 748762
rect 407224 748762 407252 750706
rect 408420 748762 408448 755806
rect 409524 755806 409658 755834
rect 409524 748762 409552 755806
rect 409602 755700 409658 755806
rect 410246 755834 410302 756500
rect 411534 755834 411590 756500
rect 412822 755834 412878 756500
rect 414110 755834 414166 756500
rect 410246 755806 410656 755834
rect 410246 755700 410302 755806
rect 410628 748762 410656 755806
rect 411534 755806 411760 755834
rect 411534 755700 411590 755806
rect 411732 748762 411760 755806
rect 407224 748734 407278 748762
rect 406146 748476 406174 748734
rect 407250 748476 407278 748734
rect 408354 748734 408448 748762
rect 409458 748734 409552 748762
rect 410562 748734 410656 748762
rect 411666 748734 411760 748762
rect 412744 755806 412878 755834
rect 412744 748762 412772 755806
rect 412822 755700 412878 755806
rect 413940 755806 414166 755834
rect 413940 748762 413968 755806
rect 414110 755700 414166 755806
rect 414754 755834 414810 756500
rect 416042 755834 416098 756500
rect 417330 755834 417386 756500
rect 417974 755834 418030 756500
rect 414754 755806 415072 755834
rect 414754 755700 414810 755806
rect 415044 748762 415072 755806
rect 416042 755806 416176 755834
rect 416042 755700 416098 755806
rect 416148 748762 416176 755806
rect 417252 755806 417386 755834
rect 417252 748762 417280 755806
rect 417330 755700 417386 755806
rect 417896 755806 418030 755834
rect 417896 750734 417924 755806
rect 417974 755700 418030 755806
rect 478786 753536 478842 753545
rect 478786 753471 478842 753480
rect 478142 751496 478198 751505
rect 478142 751431 478198 751440
rect 417896 750706 418292 750734
rect 412744 748734 412798 748762
rect 408354 748476 408382 748734
rect 409458 748476 409486 748734
rect 410562 748476 410590 748734
rect 411666 748476 411694 748734
rect 412770 748476 412798 748734
rect 413874 748734 413968 748762
rect 414978 748734 415072 748762
rect 416082 748734 416176 748762
rect 417186 748734 417280 748762
rect 418264 748762 418292 750706
rect 418264 748734 418318 748762
rect 413874 748476 413902 748734
rect 414978 748476 415006 748734
rect 416082 748476 416110 748734
rect 417186 748476 417214 748734
rect 418290 748476 418318 748734
rect 21142 744404 21496 744432
rect 21086 744381 21142 744390
rect 20626 742520 20682 742529
rect 20626 742455 20682 742464
rect 20442 740888 20498 740897
rect 20442 740823 20498 740832
rect 20166 739528 20222 739537
rect 20166 739463 20222 739472
rect 14186 738984 14242 738993
rect 14186 738919 14242 738928
rect 7746 738712 7802 738721
rect 7746 738647 7802 738656
rect 478050 724976 478106 724985
rect 478050 724911 478106 724920
rect 477958 722256 478014 722265
rect 477958 722191 478014 722200
rect 477038 716952 477094 716961
rect 477038 716887 477094 716896
rect 477052 702434 477080 716887
rect 477314 713416 477370 713425
rect 477314 713351 477370 713360
rect 477130 712192 477186 712201
rect 477130 712127 477186 712136
rect 476960 702406 477080 702434
rect 476960 673454 476988 702406
rect 477144 698294 477172 712127
rect 477144 698266 477264 698294
rect 476960 673426 477172 673454
rect 477144 671333 477172 673426
rect 477130 671324 477186 671333
rect 477130 671259 477186 671268
rect 477236 670789 477264 698266
rect 477328 695813 477356 713351
rect 477406 709200 477462 709209
rect 477406 709135 477462 709144
rect 477314 695804 477370 695813
rect 477314 695739 477370 695748
rect 477420 692345 477448 709135
rect 477972 696969 478000 722191
rect 477958 696960 478014 696969
rect 477958 696895 478014 696904
rect 478064 694249 478092 724911
rect 478050 694240 478106 694249
rect 478050 694175 478106 694184
rect 477406 692336 477462 692345
rect 477406 692271 477462 692280
rect 478156 680241 478184 751431
rect 478694 748776 478750 748785
rect 478694 748711 478750 748720
rect 478602 747416 478658 747425
rect 478602 747351 478658 747360
rect 478326 739936 478382 739945
rect 478326 739871 478382 739880
rect 478234 724296 478290 724305
rect 478234 724231 478290 724240
rect 478248 691393 478276 724231
rect 478234 691384 478290 691393
rect 478234 691319 478290 691328
rect 478142 680232 478198 680241
rect 478142 680167 478198 680176
rect 478340 679833 478368 739871
rect 478510 739256 478566 739265
rect 478510 739191 478566 739200
rect 478418 727016 478474 727025
rect 478418 726951 478474 726960
rect 478432 684457 478460 726951
rect 478418 684448 478474 684457
rect 478418 684383 478474 684392
rect 478524 681873 478552 739191
rect 478510 681864 478566 681873
rect 478510 681799 478566 681808
rect 478326 679824 478382 679833
rect 478326 679759 478382 679768
rect 478616 678473 478644 747351
rect 478708 679017 478736 748711
rect 478694 679008 478750 679017
rect 478694 678943 478750 678952
rect 478602 678464 478658 678473
rect 478602 678399 478658 678408
rect 478800 677657 478828 753471
rect 486146 752856 486202 752865
rect 486146 752791 486202 752800
rect 480902 752176 480958 752185
rect 480902 752111 480958 752120
rect 479522 749456 479578 749465
rect 479522 749391 479578 749400
rect 479430 738576 479486 738585
rect 479430 738511 479486 738520
rect 479338 717496 479394 717505
rect 479338 717431 479394 717440
rect 479352 695609 479380 717431
rect 479444 716961 479472 738511
rect 479430 716952 479486 716961
rect 479430 716887 479486 716896
rect 479430 698320 479486 698329
rect 479430 698255 479486 698264
rect 479338 695600 479394 695609
rect 479338 695535 479394 695544
rect 478786 677648 478842 677657
rect 478786 677583 478842 677592
rect 479444 677521 479472 698255
rect 479536 684321 479564 749391
rect 479798 741976 479854 741985
rect 479798 741911 479854 741920
rect 479614 741296 479670 741305
rect 479614 741231 479670 741240
rect 479628 685001 479656 741231
rect 479706 726336 479762 726345
rect 479706 726271 479762 726280
rect 479720 693025 479748 726271
rect 479706 693016 479762 693025
rect 479706 692951 479762 692960
rect 479812 685953 479840 741911
rect 480166 740616 480222 740625
rect 480166 740551 480222 740560
rect 479982 729736 480038 729745
rect 479982 729671 480038 729680
rect 479890 718176 479946 718185
rect 479890 718111 479946 718120
rect 479798 685944 479854 685953
rect 479798 685879 479854 685888
rect 479904 685137 479932 718111
rect 479996 686225 480024 729671
rect 480074 720216 480130 720225
rect 480074 720151 480130 720160
rect 479982 686216 480038 686225
rect 479982 686151 480038 686160
rect 479890 685128 479946 685137
rect 479890 685063 479946 685072
rect 479984 685092 480036 685098
rect 479984 685034 480036 685040
rect 479614 684992 479670 685001
rect 479614 684927 479670 684936
rect 479522 684312 479578 684321
rect 479522 684247 479578 684256
rect 479430 677512 479486 677521
rect 479430 677447 479486 677456
rect 479996 676977 480024 685034
rect 480088 680377 480116 720151
rect 480180 685817 480208 740551
rect 480810 727696 480866 727705
rect 480810 727631 480866 727640
rect 480824 690033 480852 727631
rect 480810 690024 480866 690033
rect 480810 689959 480866 689968
rect 480916 688401 480944 752111
rect 483754 750816 483810 750825
rect 483754 750751 483810 750760
rect 482282 750136 482338 750145
rect 482282 750071 482338 750080
rect 480994 743336 481050 743345
rect 480994 743271 481050 743280
rect 480902 688392 480958 688401
rect 480902 688327 480958 688336
rect 480166 685808 480222 685817
rect 480166 685743 480222 685752
rect 480166 685264 480222 685273
rect 480166 685199 480222 685208
rect 480074 680368 480130 680377
rect 480074 680303 480130 680312
rect 479982 676968 480038 676977
rect 479982 676903 480038 676912
rect 480180 675889 480208 685199
rect 480258 685128 480314 685137
rect 480258 685063 480260 685072
rect 480312 685063 480314 685072
rect 480260 685034 480312 685040
rect 481008 682145 481036 743271
rect 481178 742656 481234 742665
rect 481178 742591 481234 742600
rect 481086 728376 481142 728385
rect 481086 728311 481142 728320
rect 480994 682136 481050 682145
rect 480994 682071 481050 682080
rect 481100 681601 481128 728311
rect 481192 687857 481220 742591
rect 481454 735856 481510 735865
rect 481454 735791 481510 735800
rect 481362 732456 481418 732465
rect 481362 732391 481418 732400
rect 481270 729056 481326 729065
rect 481270 728991 481326 729000
rect 481178 687848 481234 687857
rect 481178 687783 481234 687792
rect 481284 682417 481312 728991
rect 481376 692753 481404 732391
rect 481362 692744 481418 692753
rect 481362 692679 481418 692688
rect 481270 682408 481326 682417
rect 481270 682343 481326 682352
rect 481086 681592 481142 681601
rect 481086 681527 481142 681536
rect 480166 675880 480222 675889
rect 480166 675815 480222 675824
rect 481468 675073 481496 735791
rect 481546 734496 481602 734505
rect 481546 734431 481602 734440
rect 481560 676161 481588 734431
rect 482098 721576 482154 721585
rect 482098 721511 482154 721520
rect 482112 712201 482140 721511
rect 482190 716816 482246 716825
rect 482190 716751 482246 716760
rect 482098 712192 482154 712201
rect 482098 712127 482154 712136
rect 482098 712056 482154 712065
rect 482098 711991 482154 712000
rect 481916 696380 481968 696386
rect 481916 696322 481968 696328
rect 481928 689761 481956 696322
rect 482006 695056 482062 695065
rect 482006 694991 482062 695000
rect 481914 689752 481970 689761
rect 481914 689687 481970 689696
rect 482020 678337 482048 694991
rect 482112 689217 482140 711991
rect 482204 709209 482232 716751
rect 482190 709200 482246 709209
rect 482190 709135 482246 709144
rect 482190 703760 482246 703769
rect 482190 703695 482246 703704
rect 482098 689208 482154 689217
rect 482098 689143 482154 689152
rect 482006 678328 482062 678337
rect 482006 678263 482062 678272
rect 482204 678201 482232 703695
rect 482296 692481 482324 750071
rect 483662 746736 483718 746745
rect 483662 746671 483718 746680
rect 482374 745376 482430 745385
rect 482374 745311 482430 745320
rect 482388 696017 482416 745311
rect 482834 744696 482890 744705
rect 482834 744631 482890 744640
rect 482650 731096 482706 731105
rect 482650 731031 482706 731040
rect 482466 730416 482522 730425
rect 482466 730351 482522 730360
rect 482374 696008 482430 696017
rect 482374 695943 482430 695952
rect 482480 694657 482508 730351
rect 482558 723616 482614 723625
rect 482558 723551 482614 723560
rect 482572 696386 482600 723551
rect 482560 696380 482612 696386
rect 482560 696322 482612 696328
rect 482560 696244 482612 696250
rect 482560 696186 482612 696192
rect 482466 694648 482522 694657
rect 482466 694583 482522 694592
rect 482572 692889 482600 696186
rect 482664 695473 482692 731031
rect 482742 718856 482798 718865
rect 482742 718791 482798 718800
rect 482650 695464 482706 695473
rect 482650 695399 482706 695408
rect 482558 692880 482614 692889
rect 482558 692815 482614 692824
rect 482282 692472 482338 692481
rect 482282 692407 482338 692416
rect 482282 689888 482338 689897
rect 482282 689823 482338 689832
rect 482190 678192 482246 678201
rect 482190 678127 482246 678136
rect 481546 676152 481602 676161
rect 481546 676087 481602 676096
rect 482296 676025 482324 689823
rect 482756 679017 482784 718791
rect 482848 696130 482876 744631
rect 482926 744016 482982 744025
rect 482926 743951 482982 743960
rect 482940 696250 482968 743951
rect 483478 701856 483534 701865
rect 483478 701791 483534 701800
rect 482928 696244 482980 696250
rect 482928 696186 482980 696192
rect 482848 696102 482968 696130
rect 482834 694376 482890 694385
rect 482834 694311 482890 694320
rect 482848 685817 482876 694311
rect 482940 694249 482968 696102
rect 482926 694240 482982 694249
rect 482926 694175 482982 694184
rect 482926 692744 482982 692753
rect 482926 692679 482982 692688
rect 482834 685808 482890 685817
rect 482834 685743 482890 685752
rect 482940 680377 482968 692679
rect 483492 684457 483520 701791
rect 483570 699816 483626 699825
rect 483570 699751 483626 699760
rect 483584 690033 483612 699751
rect 483570 690024 483626 690033
rect 483570 689959 483626 689968
rect 483478 684448 483534 684457
rect 483478 684383 483534 684392
rect 482926 680368 482982 680377
rect 482926 680303 482982 680312
rect 482742 679008 482798 679017
rect 482742 678943 482798 678952
rect 482282 676016 482338 676025
rect 482282 675951 482338 675960
rect 481454 675064 481510 675073
rect 481454 674999 481510 675008
rect 483676 671945 483704 746671
rect 483768 691257 483796 750751
rect 486160 750734 486188 752791
rect 486160 750706 486464 750734
rect 486146 748096 486202 748105
rect 486146 748031 486202 748040
rect 483938 746056 483994 746065
rect 483938 745991 483994 746000
rect 483846 731776 483902 731785
rect 483846 731711 483902 731720
rect 483860 696969 483888 731711
rect 483846 696960 483902 696969
rect 483846 696895 483902 696904
rect 483754 691248 483810 691257
rect 483754 691183 483810 691192
rect 483952 690441 483980 745991
rect 486160 741074 486188 748031
rect 486160 741046 486372 741074
rect 486146 737896 486202 737905
rect 486146 737831 486202 737840
rect 484306 736536 484362 736545
rect 484306 736471 484362 736480
rect 484214 733816 484270 733825
rect 484214 733751 484270 733760
rect 484122 733136 484178 733145
rect 484122 733071 484178 733080
rect 484030 714096 484086 714105
rect 484030 714031 484086 714040
rect 483938 690432 483994 690441
rect 483938 690367 483994 690376
rect 484044 676297 484072 714031
rect 484136 694113 484164 733071
rect 484122 694104 484178 694113
rect 484122 694039 484178 694048
rect 484030 676288 484086 676297
rect 484030 676223 484086 676232
rect 484228 676161 484256 733751
rect 484214 676152 484270 676161
rect 484214 676087 484270 676096
rect 484320 674801 484348 736471
rect 486160 731414 486188 737831
rect 486160 731386 486280 731414
rect 486146 703896 486202 703905
rect 486146 703831 486202 703840
rect 486160 692753 486188 703831
rect 486146 692744 486202 692753
rect 486146 692679 486202 692688
rect 486252 685273 486280 731386
rect 486344 689897 486372 741046
rect 486330 689888 486386 689897
rect 486330 689823 486386 689832
rect 486238 685264 486294 685273
rect 486238 685199 486294 685208
rect 486436 685137 486464 750706
rect 486422 685128 486478 685137
rect 486422 685063 486478 685072
rect 484306 674792 484362 674801
rect 484306 674727 484362 674736
rect 483662 671936 483718 671945
rect 483662 671871 483718 671880
rect 477222 670780 477278 670789
rect 477222 670715 477278 670724
rect 481546 630456 481602 630465
rect 481546 630391 481602 630400
rect 481454 628416 481510 628425
rect 481454 628351 481510 628360
rect 478786 625016 478842 625025
rect 478786 624951 478842 624960
rect 478694 624336 478750 624345
rect 478694 624271 478750 624280
rect 478708 601769 478736 624271
rect 478694 601760 478750 601769
rect 478694 601695 478750 601704
rect 478800 599185 478828 624951
rect 481468 604489 481496 628351
rect 481454 604480 481510 604489
rect 481454 604415 481510 604424
rect 481560 603129 481588 630391
rect 482926 629776 482982 629785
rect 482926 629711 482982 629720
rect 482834 627736 482890 627745
rect 482834 627671 482890 627680
rect 482282 620256 482338 620265
rect 482282 620191 482338 620200
rect 482296 607073 482324 620191
rect 482848 607209 482876 627671
rect 482834 607200 482890 607209
rect 482834 607135 482890 607144
rect 482282 607064 482338 607073
rect 482282 606999 482338 607008
rect 481546 603120 481602 603129
rect 481546 603055 481602 603064
rect 482940 601769 482968 629711
rect 484306 629096 484362 629105
rect 484306 629031 484362 629040
rect 484214 627056 484270 627065
rect 484214 626991 484270 627000
rect 483662 616856 483718 616865
rect 483662 616791 483718 616800
rect 483676 602857 483704 616791
rect 484228 607209 484256 626991
rect 484214 607200 484270 607209
rect 484214 607135 484270 607144
rect 484320 607073 484348 629031
rect 484306 607064 484362 607073
rect 484306 606999 484362 607008
rect 483662 602848 483718 602857
rect 483662 602783 483718 602792
rect 482926 601760 482982 601769
rect 482926 601695 482982 601704
rect 478786 599176 478842 599185
rect 478786 599111 478842 599120
rect 481546 587888 481602 587897
rect 481546 587823 481602 587832
rect 480166 587208 480222 587217
rect 480166 587143 480222 587152
rect 477130 584760 477186 584769
rect 477130 584695 477186 584704
rect 477144 569945 477172 584695
rect 480074 581632 480130 581641
rect 480074 581567 480130 581576
rect 477130 569936 477186 569945
rect 477130 569871 477186 569880
rect 480088 567225 480116 581567
rect 480074 567216 480130 567225
rect 480074 567151 480130 567160
rect 480180 566545 480208 587143
rect 481454 580952 481510 580961
rect 481454 580887 481510 580896
rect 481362 579048 481418 579057
rect 481362 578983 481418 578992
rect 480166 566536 480222 566545
rect 480166 566471 480222 566480
rect 481376 561785 481404 578983
rect 481362 561776 481418 561785
rect 481362 561711 481418 561720
rect 481468 557025 481496 580887
rect 481560 558385 481588 587823
rect 483662 584624 483718 584633
rect 483662 584559 483718 584568
rect 482926 582448 482982 582457
rect 482926 582383 482982 582392
rect 482834 579592 482890 579601
rect 482834 579527 482890 579536
rect 482848 561105 482876 579527
rect 482834 561096 482890 561105
rect 482834 561031 482890 561040
rect 482940 559745 482968 582383
rect 483676 570625 483704 584559
rect 484306 581632 484362 581641
rect 484306 581567 484362 581576
rect 483662 570616 483718 570625
rect 483662 570551 483718 570560
rect 482926 559736 482982 559745
rect 482926 559671 482982 559680
rect 481546 558376 481602 558385
rect 481546 558311 481602 558320
rect 484320 557705 484348 581567
rect 484306 557696 484362 557705
rect 484306 557631 484362 557640
rect 481454 557016 481510 557025
rect 481454 556951 481510 556960
rect 481546 540016 481602 540025
rect 481546 539951 481602 539960
rect 481454 538656 481510 538665
rect 481454 538591 481510 538600
rect 478786 534576 478842 534585
rect 478786 534511 478842 534520
rect 478694 533216 478750 533225
rect 478694 533151 478750 533160
rect 478602 517304 478658 517313
rect 478602 517239 478658 517248
rect 478616 516905 478644 517239
rect 478602 516896 478658 516905
rect 478602 516831 478658 516840
rect 478708 513369 478736 533151
rect 478694 513360 478750 513369
rect 478694 513295 478750 513304
rect 478800 511873 478828 534511
rect 481468 514865 481496 538591
rect 481454 514856 481510 514865
rect 481454 514791 481510 514800
rect 481560 513369 481588 539951
rect 482926 539336 482982 539345
rect 482926 539271 482982 539280
rect 482834 537296 482890 537305
rect 482834 537231 482890 537240
rect 482848 516225 482876 537231
rect 482834 516216 482890 516225
rect 482834 516151 482890 516160
rect 482940 513777 482968 539271
rect 484306 537976 484362 537985
rect 484306 537911 484362 537920
rect 484214 535936 484270 535945
rect 484214 535871 484270 535880
rect 483662 530496 483718 530505
rect 483662 530431 483718 530440
rect 483676 516497 483704 530431
rect 483662 516488 483718 516497
rect 483662 516423 483718 516432
rect 484228 516361 484256 535871
rect 484214 516352 484270 516361
rect 484214 516287 484270 516296
rect 484320 515001 484348 537911
rect 484306 514992 484362 515001
rect 484306 514927 484362 514936
rect 482926 513768 482982 513777
rect 482926 513703 482982 513712
rect 481546 513360 481602 513369
rect 481546 513295 481602 513304
rect 478786 511864 478842 511873
rect 478786 511799 478842 511808
rect 481546 496904 481602 496913
rect 481546 496839 481602 496848
rect 480166 494320 480222 494329
rect 480166 494255 480222 494264
rect 478786 492688 478842 492697
rect 478786 492623 478842 492632
rect 478800 468625 478828 492623
rect 480074 491192 480130 491201
rect 480074 491127 480130 491136
rect 480088 477465 480116 491127
rect 480074 477456 480130 477465
rect 480074 477391 480130 477400
rect 480180 476785 480208 494255
rect 481454 488608 481510 488617
rect 481454 488543 481510 488552
rect 480166 476776 480222 476785
rect 480166 476711 480222 476720
rect 478786 468616 478842 468625
rect 478786 468551 478842 468560
rect 481468 466585 481496 488543
rect 481560 469305 481588 496839
rect 486422 496224 486478 496233
rect 486422 496159 486478 496168
rect 482926 494728 482982 494737
rect 482926 494663 482982 494672
rect 484306 494728 484362 494737
rect 484306 494663 484362 494672
rect 482282 493640 482338 493649
rect 482282 493575 482338 493584
rect 482296 481545 482324 493575
rect 482834 492688 482890 492697
rect 482834 492623 482890 492632
rect 482282 481536 482338 481545
rect 482282 481471 482338 481480
rect 482848 470665 482876 492623
rect 482834 470656 482890 470665
rect 482834 470591 482890 470600
rect 481546 469296 481602 469305
rect 481546 469231 481602 469240
rect 482940 467945 482968 494663
rect 484214 494048 484270 494057
rect 484214 493983 484270 493992
rect 484228 469985 484256 493983
rect 484214 469976 484270 469985
rect 484214 469911 484270 469920
rect 482926 467936 482982 467945
rect 482926 467871 482982 467880
rect 484320 467265 484348 494663
rect 486436 480254 486464 496159
rect 486160 480226 486464 480254
rect 486160 478145 486188 480226
rect 486146 478136 486202 478145
rect 486146 478071 486202 478080
rect 484306 467256 484362 467265
rect 484306 467191 484362 467200
rect 481454 466576 481510 466585
rect 481454 466511 481510 466520
rect 482926 459776 482982 459785
rect 482926 459711 482982 459720
rect 479522 459096 479578 459105
rect 479522 459031 479578 459040
rect 478786 455016 478842 455025
rect 478786 454951 478842 454960
rect 478694 454336 478750 454345
rect 478694 454271 478750 454280
rect 478510 450936 478566 450945
rect 478510 450871 478566 450880
rect 478418 449576 478474 449585
rect 478418 449511 478474 449520
rect 478432 427281 478460 449511
rect 478418 427272 478474 427281
rect 478418 427207 478474 427216
rect 477406 424824 477462 424833
rect 477406 424759 477462 424768
rect 477420 424439 477448 424759
rect 477406 424430 477462 424439
rect 477406 424365 477462 424374
rect 477406 423464 477462 423473
rect 477406 423399 477462 423408
rect 477420 423079 477448 423399
rect 477406 423070 477462 423079
rect 477406 423005 477462 423014
rect 478524 421025 478552 450871
rect 478602 450256 478658 450265
rect 478602 450191 478658 450200
rect 478510 421016 478566 421025
rect 478510 420951 478566 420960
rect 478616 418305 478644 450191
rect 478602 418296 478658 418305
rect 478602 418231 478658 418240
rect 478708 416673 478736 454271
rect 478694 416664 478750 416673
rect 478694 416599 478750 416608
rect 478800 415313 478828 454951
rect 479536 418169 479564 459031
rect 482834 457736 482890 457745
rect 482834 457671 482890 457680
rect 482742 456376 482798 456385
rect 482742 456311 482798 456320
rect 480902 453656 480958 453665
rect 480902 453591 480958 453600
rect 480166 446176 480222 446185
rect 480166 446111 480222 446120
rect 479982 445496 480038 445505
rect 479982 445431 480038 445440
rect 479890 444136 479946 444145
rect 479890 444071 479946 444080
rect 479904 427281 479932 444071
rect 479890 427272 479946 427281
rect 479890 427207 479946 427216
rect 479996 424561 480024 445431
rect 480074 444816 480130 444825
rect 480074 444751 480130 444760
rect 479982 424552 480038 424561
rect 479982 424487 480038 424496
rect 479522 418160 479578 418169
rect 479522 418095 479578 418104
rect 480088 417353 480116 444751
rect 480180 419529 480208 446111
rect 480916 424153 480944 453591
rect 481546 452296 481602 452305
rect 481546 452231 481602 452240
rect 481454 451616 481510 451625
rect 481454 451551 481510 451560
rect 480902 424144 480958 424153
rect 480902 424079 480958 424088
rect 481468 421433 481496 451551
rect 481560 423609 481588 452231
rect 482650 448896 482706 448905
rect 482650 448831 482706 448840
rect 482006 429448 482062 429457
rect 482006 429383 482062 429392
rect 482020 426193 482048 429383
rect 482664 426193 482692 448831
rect 482006 426184 482062 426193
rect 482006 426119 482062 426128
rect 482650 426184 482706 426193
rect 482650 426119 482706 426128
rect 481546 423600 481602 423609
rect 481546 423535 481602 423544
rect 481454 421424 481510 421433
rect 481454 421359 481510 421368
rect 481454 420064 481510 420073
rect 481454 419999 481510 420008
rect 481468 419801 481496 419999
rect 482756 419801 482784 456311
rect 481454 419792 481510 419801
rect 481454 419727 481510 419736
rect 482742 419792 482798 419801
rect 482742 419727 482798 419736
rect 482848 419665 482876 457671
rect 482834 419656 482890 419665
rect 482834 419591 482890 419600
rect 480166 419520 480222 419529
rect 480166 419455 480222 419464
rect 480074 417344 480130 417353
rect 480074 417279 480130 417288
rect 482940 416673 482968 459711
rect 484306 458416 484362 458425
rect 484306 458351 484362 458360
rect 484214 457056 484270 457065
rect 484214 456991 484270 457000
rect 484122 455696 484178 455705
rect 484122 455631 484178 455640
rect 484030 448216 484086 448225
rect 484030 448151 484086 448160
rect 484044 424969 484072 448151
rect 483110 424960 483166 424969
rect 483110 424895 483166 424904
rect 484030 424960 484086 424969
rect 484030 424895 484086 424904
rect 483124 424561 483152 424895
rect 483110 424552 483166 424561
rect 483110 424487 483166 424496
rect 484136 423609 484164 455631
rect 484122 423600 484178 423609
rect 484122 423535 484178 423544
rect 484228 416673 484256 456991
rect 482926 416664 482982 416673
rect 482926 416599 482982 416608
rect 484214 416664 484270 416673
rect 484214 416599 484270 416608
rect 484320 415313 484348 458351
rect 486146 446856 486202 446865
rect 486146 446791 486202 446800
rect 486160 441614 486188 446791
rect 486160 441586 486280 441614
rect 486146 438016 486202 438025
rect 486146 437951 486202 437960
rect 486054 424552 486110 424561
rect 486160 424538 486188 437951
rect 486252 429457 486280 441586
rect 486238 429448 486294 429457
rect 486238 429383 486294 429392
rect 486110 424510 486188 424538
rect 486054 424487 486110 424496
rect 478786 415304 478842 415313
rect 478786 415239 478842 415248
rect 484306 415304 484362 415313
rect 484306 415239 484362 415248
rect 478786 399528 478842 399537
rect 478786 399463 478842 399472
rect 478694 398848 478750 398857
rect 478694 398783 478750 398792
rect 478708 387705 478736 398783
rect 478694 387696 478750 387705
rect 478694 387631 478750 387640
rect 478800 387025 478828 399463
rect 479522 398848 479578 398857
rect 479522 398783 479578 398792
rect 478786 387016 478842 387025
rect 478786 386951 478842 386960
rect 479536 386345 479564 398783
rect 479522 386336 479578 386345
rect 479522 386271 479578 386280
rect 481546 360496 481602 360505
rect 481546 360431 481602 360440
rect 481454 358456 481510 358465
rect 481454 358391 481510 358400
rect 478786 355056 478842 355065
rect 478786 354991 478842 355000
rect 478694 353696 478750 353705
rect 478694 353631 478750 353640
rect 477130 349616 477186 349625
rect 477130 349551 477186 349560
rect 477144 335821 477172 349551
rect 477130 335812 477186 335821
rect 477130 335747 477186 335756
rect 478708 334121 478736 353631
rect 478694 334112 478750 334121
rect 478694 334047 478750 334056
rect 478800 329633 478828 354991
rect 481468 336705 481496 358391
rect 481454 336696 481510 336705
rect 481454 336631 481510 336640
rect 481560 334121 481588 360431
rect 484306 359816 484362 359825
rect 484306 359751 484362 359760
rect 482926 359136 482982 359145
rect 482926 359071 482982 359080
rect 482282 346896 482338 346905
rect 482282 346831 482338 346840
rect 481546 334112 481602 334121
rect 481546 334047 481602 334056
rect 482296 332761 482324 346831
rect 482940 336705 482968 359071
rect 484214 357776 484270 357785
rect 484214 357711 484270 357720
rect 484228 336705 484256 357711
rect 482926 336696 482982 336705
rect 482926 336631 482982 336640
rect 484214 336696 484270 336705
rect 484214 336631 484270 336640
rect 484320 334121 484348 359751
rect 484306 334112 484362 334121
rect 484306 334047 484362 334056
rect 482282 332752 482338 332761
rect 482282 332687 482338 332696
rect 478786 329624 478842 329633
rect 478786 329559 478842 329568
rect 481546 318744 481602 318753
rect 481546 318679 481602 318688
rect 480166 314936 480222 314945
rect 480166 314871 480222 314880
rect 480074 311264 480130 311273
rect 480074 311199 480130 311208
rect 479982 310448 480038 310457
rect 479982 310383 480038 310392
rect 479996 297945 480024 310383
rect 479982 297936 480038 297945
rect 479982 297871 480038 297880
rect 480088 297265 480116 311199
rect 480074 297256 480130 297265
rect 480074 297191 480130 297200
rect 480180 296585 480208 314871
rect 481454 310448 481510 310457
rect 481454 310383 481510 310392
rect 480166 296576 480222 296585
rect 480166 296511 480222 296520
rect 481468 287065 481496 310383
rect 481560 288425 481588 318679
rect 486054 314800 486110 314809
rect 486054 314735 486110 314744
rect 482282 314528 482338 314537
rect 482282 314463 482338 314472
rect 482296 300665 482324 314463
rect 482926 311944 482982 311953
rect 482926 311879 482982 311888
rect 482834 308952 482890 308961
rect 482834 308887 482890 308896
rect 482282 300656 482338 300665
rect 482282 300591 482338 300600
rect 482848 289785 482876 308887
rect 482834 289776 482890 289785
rect 482834 289711 482890 289720
rect 481546 288416 481602 288425
rect 481546 288351 481602 288360
rect 482940 287745 482968 311879
rect 484306 311264 484362 311273
rect 484306 311199 484362 311208
rect 484320 289105 484348 311199
rect 486068 299985 486096 314735
rect 486054 299976 486110 299985
rect 486054 299911 486110 299920
rect 484306 289096 484362 289105
rect 484306 289031 484362 289040
rect 482926 287736 482982 287745
rect 482926 287671 482982 287680
rect 481454 287056 481510 287065
rect 481454 286991 481510 287000
rect 481546 270056 481602 270065
rect 481546 269991 481602 270000
rect 481454 268016 481510 268025
rect 481454 267951 481510 267960
rect 478694 264616 478750 264625
rect 478694 264551 478750 264560
rect 478602 263256 478658 263265
rect 478602 263191 478658 263200
rect 478616 247081 478644 263191
rect 478602 247072 478658 247081
rect 478602 247007 478658 247016
rect 478708 245721 478736 264551
rect 478786 263936 478842 263945
rect 478786 263871 478842 263880
rect 478694 245712 478750 245721
rect 478694 245647 478750 245656
rect 478800 242865 478828 263871
rect 481468 247081 481496 267951
rect 481454 247072 481510 247081
rect 481454 247007 481510 247016
rect 481560 244361 481588 269991
rect 482926 269376 482982 269385
rect 482926 269311 482982 269320
rect 482834 266656 482890 266665
rect 482834 266591 482890 266600
rect 482848 247081 482876 266591
rect 482834 247072 482890 247081
rect 482834 247007 482890 247016
rect 482940 245721 482968 269311
rect 484306 268696 484362 268705
rect 484306 268631 484362 268640
rect 483662 255776 483718 255785
rect 483662 255711 483718 255720
rect 483202 248296 483258 248305
rect 483202 248231 483258 248240
rect 483216 248033 483244 248231
rect 483202 248024 483258 248033
rect 483202 247959 483258 247968
rect 482926 245712 482982 245721
rect 482926 245647 482982 245656
rect 481546 244352 481602 244361
rect 481546 244287 481602 244296
rect 478786 242856 478842 242865
rect 478786 242791 478842 242800
rect 483676 241777 483704 255711
rect 484320 243545 484348 268631
rect 484306 243536 484362 243545
rect 484306 243471 484362 243480
rect 483662 241768 483718 241777
rect 483662 241703 483718 241712
rect 482926 241496 482982 241505
rect 482926 241431 482982 241440
rect 482940 240417 482968 241431
rect 482926 240408 482982 240417
rect 482926 240343 482982 240352
rect 481546 226400 481602 226409
rect 481546 226335 481602 226344
rect 481454 224088 481510 224097
rect 481454 224023 481510 224032
rect 481468 223825 481496 224023
rect 481454 223816 481510 223825
rect 481454 223751 481510 223760
rect 480166 223680 480222 223689
rect 480166 223615 480222 223624
rect 478786 220960 478842 220969
rect 478786 220895 478842 220904
rect 477406 219350 477462 219359
rect 477406 219285 477462 219294
rect 478694 219328 478750 219337
rect 477420 218385 477448 219285
rect 478694 219263 478750 219272
rect 477406 218376 477462 218385
rect 477406 218311 477462 218320
rect 478708 198665 478736 219263
rect 478694 198656 478750 198665
rect 478694 198591 478750 198600
rect 478800 197985 478828 220895
rect 480180 206825 480208 223615
rect 481454 221368 481510 221377
rect 481454 221303 481510 221312
rect 481468 221105 481496 221303
rect 481454 221096 481510 221105
rect 481454 221031 481510 221040
rect 481454 220960 481510 220969
rect 481454 220895 481510 220904
rect 480166 206816 480222 206825
rect 480166 206751 480222 206760
rect 478786 197976 478842 197985
rect 478786 197911 478842 197920
rect 481468 196625 481496 220895
rect 481560 199345 481588 226335
rect 486422 226128 486478 226137
rect 486422 226063 486478 226072
rect 482926 223680 482982 223689
rect 482926 223615 482982 223624
rect 484306 223680 484362 223689
rect 484306 223615 484362 223624
rect 482834 220960 482890 220969
rect 482834 220895 482890 220904
rect 482848 202065 482876 220895
rect 482834 202056 482890 202065
rect 482834 201991 482890 202000
rect 482940 200705 482968 223615
rect 484214 222320 484270 222329
rect 484214 222255 484270 222264
rect 482926 200696 482982 200705
rect 482926 200631 482982 200640
rect 484228 200025 484256 222255
rect 484214 200016 484270 200025
rect 484214 199951 484270 199960
rect 481546 199336 481602 199345
rect 481546 199271 481602 199280
rect 484320 197305 484348 223615
rect 486436 209774 486464 226063
rect 486160 209746 486464 209774
rect 486160 208185 486188 209746
rect 486146 208176 486202 208185
rect 486146 208111 486202 208120
rect 484306 197296 484362 197305
rect 484306 197231 484362 197240
rect 481454 196616 481510 196625
rect 481454 196551 481510 196560
rect 482926 192536 482982 192545
rect 482926 192471 482982 192480
rect 478142 191856 478198 191865
rect 478142 191791 478198 191800
rect 478156 144673 478184 191791
rect 480166 190496 480222 190505
rect 480166 190431 480222 190440
rect 479522 189816 479578 189825
rect 479522 189751 479578 189760
rect 478694 185736 478750 185745
rect 478694 185671 478750 185680
rect 478602 184376 478658 184385
rect 478602 184311 478658 184320
rect 478510 180976 478566 180985
rect 478510 180911 478566 180920
rect 478524 152969 478552 180911
rect 478510 152960 478566 152969
rect 478510 152895 478566 152904
rect 478616 152697 478644 184311
rect 478602 152688 478658 152697
rect 478602 152623 478658 152632
rect 478708 147801 478736 185671
rect 478786 185056 478842 185065
rect 478786 184991 478842 185000
rect 478694 147792 478750 147801
rect 478694 147727 478750 147736
rect 478800 144809 478828 184991
rect 479536 147121 479564 189751
rect 479982 177576 480038 177585
rect 479982 177511 480038 177520
rect 479890 176216 479946 176225
rect 479890 176151 479946 176160
rect 479904 156777 479932 176151
rect 479890 156768 479946 156777
rect 479890 156703 479946 156712
rect 479996 148753 480024 177511
rect 480074 176896 480130 176905
rect 480074 176831 480130 176840
rect 480088 148889 480116 176831
rect 480074 148880 480130 148889
rect 480074 148815 480130 148824
rect 479982 148744 480038 148753
rect 479982 148679 480038 148688
rect 479522 147112 479578 147121
rect 479522 147047 479578 147056
rect 480180 146441 480208 190431
rect 482834 188456 482890 188465
rect 482834 188391 482890 188400
rect 482742 187096 482798 187105
rect 482742 187031 482798 187040
rect 480902 183696 480958 183705
rect 480902 183631 480958 183640
rect 480916 154193 480944 183631
rect 480994 183016 481050 183025
rect 480994 182951 481050 182960
rect 481008 154737 481036 182951
rect 481546 182336 481602 182345
rect 481546 182271 481602 182280
rect 481454 175536 481510 175545
rect 481454 175471 481510 175480
rect 480994 154728 481050 154737
rect 480994 154663 481050 154672
rect 480902 154184 480958 154193
rect 480902 154119 480958 154128
rect 481468 147121 481496 175471
rect 481560 153105 481588 182271
rect 482650 179616 482706 179625
rect 482650 179551 482706 179560
rect 481638 162752 481694 162761
rect 481638 162687 481694 162696
rect 481652 155961 481680 162687
rect 481638 155952 481694 155961
rect 481638 155887 481694 155896
rect 481546 153096 481602 153105
rect 481546 153031 481602 153040
rect 482664 150521 482692 179551
rect 482650 150512 482706 150521
rect 482650 150447 482706 150456
rect 482756 149161 482784 187031
rect 482848 149297 482876 188391
rect 482834 149288 482890 149297
rect 482834 149223 482890 149232
rect 482742 149152 482798 149161
rect 482742 149087 482798 149096
rect 481454 147112 481510 147121
rect 481454 147047 481510 147056
rect 480166 146432 480222 146441
rect 480166 146367 480222 146376
rect 482940 146305 482968 192471
rect 484030 191176 484086 191185
rect 484030 191111 484086 191120
rect 483938 178936 483994 178945
rect 483938 178871 483994 178880
rect 483662 166696 483718 166705
rect 483662 166631 483718 166640
rect 483676 152833 483704 166631
rect 483952 157457 483980 178871
rect 483938 157448 483994 157457
rect 483938 157383 483994 157392
rect 484044 155961 484072 191111
rect 484306 189136 484362 189145
rect 484306 189071 484362 189080
rect 484214 187776 484270 187785
rect 484214 187711 484270 187720
rect 484122 186416 484178 186425
rect 484122 186351 484178 186360
rect 484030 155952 484086 155961
rect 484030 155887 484086 155896
rect 483662 152824 483718 152833
rect 483662 152759 483718 152768
rect 483110 151736 483166 151745
rect 483110 151671 483166 151680
rect 483124 150929 483152 151671
rect 483110 150920 483166 150929
rect 483110 150855 483166 150864
rect 484136 150521 484164 186351
rect 484122 150512 484178 150521
rect 484122 150447 484178 150456
rect 484228 147801 484256 187711
rect 484214 147792 484270 147801
rect 484214 147727 484270 147736
rect 484320 146305 484348 189071
rect 486146 178256 486202 178265
rect 486146 178191 486202 178200
rect 486160 171134 486188 178191
rect 486068 171106 486188 171134
rect 486068 162761 486096 171106
rect 486146 168056 486202 168065
rect 486146 167991 486202 168000
rect 486054 162752 486110 162761
rect 486054 162687 486110 162696
rect 486160 161474 486188 167991
rect 486160 161446 486280 161474
rect 486252 154873 486280 161446
rect 486238 154864 486294 154873
rect 486238 154799 486294 154808
rect 482926 146296 482982 146305
rect 482926 146231 482982 146240
rect 484306 146296 484362 146305
rect 484306 146231 484362 146240
rect 478786 144800 478842 144809
rect 478786 144735 478842 144744
rect 478142 144664 478198 144673
rect 478142 144599 478198 144608
rect 483662 135144 483718 135153
rect 483662 135079 483718 135088
rect 483676 119785 483704 135079
rect 483662 119776 483718 119785
rect 483662 119711 483718 119720
rect 481546 90536 481602 90545
rect 481546 90471 481602 90480
rect 481454 88496 481510 88505
rect 481454 88431 481510 88440
rect 478694 85096 478750 85105
rect 478694 85031 478750 85040
rect 478708 63753 478736 85031
rect 478786 84416 478842 84425
rect 478786 84351 478842 84360
rect 478694 63744 478750 63753
rect 478694 63679 478750 63688
rect 478800 60625 478828 84351
rect 480166 81016 480222 81025
rect 480166 80951 480222 80960
rect 480180 66201 480208 80951
rect 481468 67561 481496 88431
rect 481454 67552 481510 67561
rect 481454 67487 481510 67496
rect 480166 66192 480222 66201
rect 480166 66127 480222 66136
rect 481560 62257 481588 90471
rect 484306 89856 484362 89865
rect 484306 89791 484362 89800
rect 482926 89176 482982 89185
rect 482926 89111 482982 89120
rect 482834 87136 482890 87145
rect 482834 87071 482890 87080
rect 482282 79656 482338 79665
rect 482282 79591 482338 79600
rect 482296 64161 482324 79591
rect 482848 67561 482876 87071
rect 482834 67552 482890 67561
rect 482834 67487 482890 67496
rect 482282 64152 482338 64161
rect 482282 64087 482338 64096
rect 482940 62257 482968 89111
rect 484214 87816 484270 87825
rect 484214 87751 484270 87760
rect 484228 67561 484256 87751
rect 484214 67552 484270 67561
rect 484214 67487 484270 67496
rect 484320 65929 484348 89791
rect 484306 65920 484362 65929
rect 484306 65855 484362 65864
rect 481546 62248 481602 62257
rect 481546 62183 481602 62192
rect 482926 62248 482982 62257
rect 482926 62183 482982 62192
rect 478786 60616 478842 60625
rect 478786 60551 478842 60560
rect 481546 48240 481602 48249
rect 481546 48175 481602 48184
rect 477222 47424 477278 47433
rect 477222 47359 477278 47368
rect 477236 47025 477264 47359
rect 477222 47016 477278 47025
rect 477222 46951 477278 46960
rect 480166 44432 480222 44441
rect 480166 44367 480222 44376
rect 480074 39944 480130 39953
rect 480074 39879 480130 39888
rect 6182 32056 6238 32065
rect 6182 31991 6238 32000
rect 4802 31376 4858 31385
rect 4802 31311 4858 31320
rect 1122 30696 1178 30705
rect 1122 30631 1178 30640
rect 1136 28937 1164 30631
rect 1122 28928 1178 28937
rect 1122 28863 1178 28872
rect 202 28384 258 28393
rect 202 28319 258 28328
rect 216 18057 244 28319
rect 1306 27976 1362 27985
rect 1306 27911 1362 27920
rect 1214 26616 1270 26625
rect 1214 26551 1270 26560
rect 1228 22001 1256 26551
rect 1320 23769 1348 27911
rect 3422 23896 3478 23905
rect 3422 23831 3478 23840
rect 1306 23760 1362 23769
rect 1306 23695 1362 23704
rect 1214 21992 1270 22001
rect 1214 21927 1270 21936
rect 202 18048 258 18057
rect 202 17983 258 17992
rect 3436 16153 3464 23831
rect 4816 16561 4844 31311
rect 4894 29336 4950 29345
rect 4894 29271 4950 29280
rect 4908 16833 4936 29271
rect 5078 28928 5134 28937
rect 5078 28863 5134 28872
rect 5092 17921 5120 28863
rect 5538 23216 5594 23225
rect 5538 23151 5594 23160
rect 5078 17912 5134 17921
rect 5078 17847 5134 17856
rect 4894 16824 4950 16833
rect 4894 16759 4950 16768
rect 5552 16697 5580 23151
rect 6196 17134 6224 31991
rect 7102 31240 7158 31249
rect 7102 31175 7158 31184
rect 6458 23080 6514 23089
rect 6458 23015 6514 23024
rect 6184 17128 6236 17134
rect 6184 17070 6236 17076
rect 5538 16688 5594 16697
rect 5538 16623 5594 16632
rect 4802 16552 4858 16561
rect 4802 16487 4858 16496
rect 3422 16144 3478 16153
rect 3422 16079 3478 16088
rect 6472 800 6500 23015
rect 7116 800 7144 31175
rect 9310 30424 9366 30433
rect 9310 30359 9366 30368
rect 7562 30016 7618 30025
rect 7562 29951 7618 29960
rect 7378 23760 7434 23769
rect 7378 23695 7434 23704
rect 7392 16930 7420 23695
rect 7576 17066 7604 29951
rect 8666 28792 8722 28801
rect 8666 28727 8722 28736
rect 8206 27976 8262 27985
rect 8206 27911 8262 27920
rect 7654 27296 7710 27305
rect 7654 27231 7710 27240
rect 7668 17270 7696 27231
rect 8022 27160 8078 27169
rect 8022 27095 8078 27104
rect 7746 23896 7802 23905
rect 7746 23831 7802 23840
rect 7656 17264 7708 17270
rect 7656 17206 7708 17212
rect 7564 17060 7616 17066
rect 7564 17002 7616 17008
rect 7380 16924 7432 16930
rect 7380 16866 7432 16872
rect 7760 800 7788 23831
rect 8036 1057 8064 27095
rect 8116 16584 8168 16590
rect 8114 16552 8116 16561
rect 8168 16552 8170 16561
rect 8114 16487 8170 16496
rect 8220 6914 8248 27911
rect 8482 18048 8538 18057
rect 8482 17983 8538 17992
rect 8496 16862 8524 17983
rect 8484 16856 8536 16862
rect 8484 16798 8536 16804
rect 8128 6886 8248 6914
rect 8022 1048 8078 1057
rect 8022 983 8078 992
rect 8128 921 8156 6886
rect 8390 1320 8446 1329
rect 8390 1255 8446 1264
rect 8114 912 8170 921
rect 8114 847 8170 856
rect 8404 800 8432 1255
rect 8680 1193 8708 28727
rect 8942 25256 8998 25265
rect 8942 25191 8998 25200
rect 8850 21992 8906 22001
rect 8850 21927 8906 21936
rect 8864 16998 8892 21927
rect 8852 16992 8904 16998
rect 8852 16934 8904 16940
rect 8956 16289 8984 25191
rect 9034 24712 9090 24721
rect 9034 24647 9090 24656
rect 8942 16280 8998 16289
rect 8942 16215 8998 16224
rect 8666 1184 8722 1193
rect 8666 1119 8722 1128
rect 9048 800 9076 24647
rect 9126 20496 9182 20505
rect 9126 20431 9182 20440
rect 9140 17513 9168 20431
rect 9218 17912 9274 17921
rect 9218 17847 9274 17856
rect 9126 17504 9182 17513
rect 9126 17439 9182 17448
rect 9232 17202 9260 17847
rect 9220 17196 9272 17202
rect 9220 17138 9272 17144
rect 9324 4185 9352 30359
rect 9586 29540 9642 29549
rect 9586 29475 9642 29484
rect 9402 26344 9458 26353
rect 9402 26279 9458 26288
rect 9310 4176 9366 4185
rect 9310 4111 9366 4120
rect 9416 1329 9444 26279
rect 9494 19816 9550 19825
rect 9494 19751 9550 19760
rect 9508 16969 9536 19751
rect 9494 16960 9550 16969
rect 9494 16895 9550 16904
rect 9402 1320 9458 1329
rect 9600 1306 9628 29475
rect 480088 27305 480116 39879
rect 480074 27296 480130 27305
rect 480074 27231 480130 27240
rect 480180 26625 480208 44367
rect 480166 26616 480222 26625
rect 480166 26551 480222 26560
rect 481560 18465 481588 48175
rect 486422 44704 486478 44713
rect 486422 44639 486478 44648
rect 483110 44296 483166 44305
rect 483110 44231 483166 44240
rect 482926 41440 482982 41449
rect 482926 41375 482982 41384
rect 482834 39944 482890 39953
rect 482834 39879 482890 39888
rect 482848 21185 482876 39879
rect 482834 21176 482890 21185
rect 482834 21111 482890 21120
rect 482940 19825 482968 41375
rect 483124 30705 483152 44231
rect 484306 43344 484362 43353
rect 484306 43279 484362 43288
rect 483294 43208 483350 43217
rect 483294 43143 483350 43152
rect 483308 42945 483336 43143
rect 483294 42936 483350 42945
rect 483294 42871 483350 42880
rect 484214 41440 484270 41449
rect 484214 41375 484270 41384
rect 483110 30696 483166 30705
rect 483110 30631 483166 30640
rect 482926 19816 482982 19825
rect 482926 19751 482982 19760
rect 484228 19145 484256 41375
rect 484214 19136 484270 19145
rect 484214 19071 484270 19080
rect 481546 18456 481602 18465
rect 481546 18391 481602 18400
rect 484320 17785 484348 43279
rect 486436 35894 486464 44639
rect 486160 35866 486464 35894
rect 486160 30025 486188 35866
rect 486146 30016 486202 30025
rect 486146 29951 486202 29960
rect 484306 17776 484362 17785
rect 484306 17711 484362 17720
rect 10980 8265 11008 17278
rect 11394 17134 11422 17272
rect 11382 17128 11434 17134
rect 11382 17070 11434 17076
rect 11900 16833 11928 17278
rect 12360 16969 12388 17278
rect 12346 16960 12402 16969
rect 12346 16895 12402 16904
rect 11886 16824 11942 16833
rect 11886 16759 11942 16768
rect 12820 16017 12848 17278
rect 13234 17105 13262 17272
rect 13694 17105 13722 17272
rect 13220 17096 13276 17105
rect 13220 17031 13276 17040
rect 13680 17096 13736 17105
rect 13680 17031 13736 17040
rect 14200 16697 14228 17278
rect 14614 17202 14642 17272
rect 15074 17202 15102 17272
rect 14602 17196 14654 17202
rect 14602 17138 14654 17144
rect 15062 17196 15114 17202
rect 15062 17138 15114 17144
rect 14186 16688 14242 16697
rect 14186 16623 14242 16632
rect 15580 16153 15608 17278
rect 16040 16289 16068 17278
rect 16500 16590 16528 17278
rect 16488 16584 16540 16590
rect 16960 16561 16988 17278
rect 17420 16969 17448 17278
rect 17834 17105 17862 17272
rect 17820 17096 17876 17105
rect 17820 17031 17876 17040
rect 18340 16998 18368 17278
rect 18754 17105 18782 17272
rect 18740 17096 18796 17105
rect 18740 17031 18796 17040
rect 18328 16992 18380 16998
rect 17406 16960 17462 16969
rect 18328 16934 18380 16940
rect 19260 16930 19288 17278
rect 17406 16895 17462 16904
rect 19248 16924 19300 16930
rect 19248 16866 19300 16872
rect 19720 16862 19748 17278
rect 20134 17066 20162 17272
rect 20122 17060 20174 17066
rect 20122 17002 20174 17008
rect 19708 16856 19760 16862
rect 19708 16798 19760 16804
rect 16488 16526 16540 16532
rect 16946 16552 17002 16561
rect 16946 16487 17002 16496
rect 16026 16280 16082 16289
rect 16026 16215 16082 16224
rect 15566 16144 15622 16153
rect 15566 16079 15622 16088
rect 12806 16008 12862 16017
rect 12806 15943 12862 15952
rect 18878 13696 18934 13705
rect 18878 13631 18934 13640
rect 18892 13025 18920 13631
rect 18878 13016 18934 13025
rect 18878 12951 18934 12960
rect 11518 12336 11574 12345
rect 11518 12271 11574 12280
rect 11532 12186 11560 12271
rect 11794 12200 11850 12209
rect 11532 12158 11794 12186
rect 11794 12135 11850 12144
rect 20350 9072 20406 9081
rect 20350 9007 20406 9016
rect 10966 8256 11022 8265
rect 10966 8191 11022 8200
rect 14186 8256 14242 8265
rect 14186 8191 14242 8200
rect 14200 5953 14228 8191
rect 20364 7993 20392 9007
rect 21086 8256 21142 8265
rect 21142 8214 21496 8242
rect 21086 8191 21142 8200
rect 20350 7984 20406 7993
rect 20350 7919 20406 7928
rect 20534 7984 20590 7993
rect 20534 7919 20590 7928
rect 14186 5944 14242 5953
rect 14186 5879 14242 5888
rect 11610 5672 11666 5681
rect 11610 5607 11666 5616
rect 10322 1320 10378 1329
rect 9600 1278 9720 1306
rect 9402 1255 9458 1264
rect 9692 800 9720 1278
rect 10322 1255 10378 1264
rect 10336 800 10364 1255
rect 10966 1184 11022 1193
rect 10966 1119 11022 1128
rect 10980 800 11008 1119
rect 11624 800 11652 5607
rect 12898 4176 12954 4185
rect 12898 4111 12954 4120
rect 12254 1048 12310 1057
rect 12254 983 12310 992
rect 12268 800 12296 983
rect 12912 800 12940 4111
rect 13542 912 13598 921
rect 13542 847 13598 856
rect 13556 800 13584 847
rect 14200 800 14228 5879
rect 20548 3482 20576 7919
rect 21086 7712 21142 7721
rect 21086 7647 21142 7656
rect 20626 7440 20682 7449
rect 20626 7375 20682 7384
rect 20640 3641 20668 7375
rect 21100 6914 21128 7647
rect 21100 6886 21312 6914
rect 20626 3632 20682 3641
rect 20626 3567 20682 3576
rect 20548 3454 20668 3482
rect 20640 800 20668 3454
rect 21284 800 21312 6886
rect 6458 0 6514 800
rect 7102 0 7158 800
rect 7746 0 7802 800
rect 8390 0 8446 800
rect 9034 0 9090 800
rect 9678 0 9734 800
rect 10322 0 10378 800
rect 10966 0 11022 800
rect 11610 0 11666 800
rect 12254 0 12310 800
rect 12898 0 12954 800
rect 13542 0 13598 800
rect 14186 0 14242 800
rect 20626 0 20682 800
rect 21270 0 21326 800
rect 21468 762 21496 8214
rect 22558 3632 22614 3641
rect 22558 3567 22614 3576
rect 21836 870 21956 898
rect 21836 762 21864 870
rect 21928 800 21956 870
rect 22572 800 22600 3567
rect 21468 734 21864 762
rect 21914 0 21970 800
rect 22558 0 22614 800
rect 22940 762 22968 6028
rect 23124 870 23244 898
rect 23124 762 23152 870
rect 23216 800 23244 870
rect 24504 800 24532 6028
rect 25792 870 25912 898
rect 25792 800 25820 870
rect 22940 734 23152 762
rect 23202 0 23258 800
rect 24490 0 24546 800
rect 25778 0 25834 800
rect 25884 762 25912 870
rect 26068 762 26096 6028
rect 27632 1578 27660 6028
rect 29196 5953 29224 6028
rect 29182 5944 29238 5953
rect 29182 5879 29238 5888
rect 30760 3074 30788 6028
rect 32322 5794 32350 6028
rect 32232 5766 32350 5794
rect 30760 3046 30972 3074
rect 27632 1550 27752 1578
rect 27724 800 27752 1550
rect 30944 800 30972 3046
rect 32232 800 32260 5766
rect 25884 734 26096 762
rect 27710 0 27766 800
rect 30930 0 30986 800
rect 32218 0 32274 800
rect 33888 762 33916 6028
rect 34072 870 34192 898
rect 34072 762 34100 870
rect 34164 800 34192 870
rect 35452 800 35480 6028
rect 36740 870 36860 898
rect 36740 800 36768 870
rect 33888 734 34100 762
rect 34150 0 34206 800
rect 35438 0 35494 800
rect 36726 0 36782 800
rect 36832 762 36860 870
rect 37016 762 37044 6028
rect 38580 1306 38608 6028
rect 40142 5794 40170 6028
rect 39960 5766 40170 5794
rect 38580 1278 38700 1306
rect 38672 800 38700 1278
rect 39960 800 39988 5766
rect 41708 3074 41736 6028
rect 43270 5794 43298 6028
rect 43180 5766 43298 5794
rect 41708 3046 41920 3074
rect 41892 800 41920 3046
rect 43180 800 43208 5766
rect 36832 734 37044 762
rect 38658 0 38714 800
rect 39946 0 40002 800
rect 41878 0 41934 800
rect 43166 0 43222 800
rect 44836 762 44864 6028
rect 45020 870 45140 898
rect 45020 762 45048 870
rect 45112 800 45140 870
rect 46400 800 46428 6028
rect 47688 870 47808 898
rect 47688 800 47716 870
rect 44836 734 45048 762
rect 45098 0 45154 800
rect 46386 0 46442 800
rect 47674 0 47730 800
rect 47780 762 47808 870
rect 47964 762 47992 6028
rect 49528 3074 49556 6028
rect 51090 5794 51118 6028
rect 50908 5766 51118 5794
rect 49528 3046 49648 3074
rect 49620 800 49648 3046
rect 50908 800 50936 5766
rect 52656 3074 52684 6028
rect 54218 5794 54246 6028
rect 54128 5766 54246 5794
rect 52656 3046 52868 3074
rect 52840 800 52868 3046
rect 54128 800 54156 5766
rect 47780 734 47992 762
rect 49606 0 49662 800
rect 50894 0 50950 800
rect 52826 0 52882 800
rect 54114 0 54170 800
rect 55784 762 55812 6028
rect 55968 870 56088 898
rect 55968 762 55996 870
rect 56060 800 56088 870
rect 57348 800 57376 6028
rect 58636 870 58756 898
rect 58636 800 58664 870
rect 55784 734 55996 762
rect 56046 0 56102 800
rect 57334 0 57390 800
rect 58622 0 58678 800
rect 58728 762 58756 870
rect 58912 762 58940 6028
rect 60476 3074 60504 6028
rect 63570 5794 63598 6028
rect 65042 5794 65070 6028
rect 66502 5794 66530 6028
rect 63570 5766 63816 5794
rect 65042 5766 65104 5794
rect 60476 3046 60596 3074
rect 60568 800 60596 3046
rect 63788 800 63816 5766
rect 65076 800 65104 5766
rect 66364 5766 66530 5794
rect 67986 5794 68014 6028
rect 69458 5794 69486 6028
rect 70918 5794 70946 6028
rect 72390 5953 72418 6028
rect 72376 5944 72432 5953
rect 72376 5879 72432 5888
rect 67986 5766 68048 5794
rect 69458 5766 69612 5794
rect 66364 800 66392 5766
rect 58728 734 58940 762
rect 60554 0 60610 800
rect 63774 0 63830 800
rect 65062 0 65118 800
rect 66350 0 66406 800
rect 68020 762 68048 5766
rect 68204 870 68324 898
rect 68204 762 68232 870
rect 68296 800 68324 870
rect 69584 800 69612 5766
rect 70872 5766 70946 5794
rect 73874 5794 73902 6028
rect 75346 5794 75374 6028
rect 76806 5794 76834 6028
rect 73874 5766 74120 5794
rect 75346 5766 75408 5794
rect 70872 800 70900 5766
rect 74092 800 74120 5766
rect 75380 800 75408 5766
rect 76668 5766 76834 5794
rect 78290 5794 78318 6028
rect 79762 5794 79790 6028
rect 81222 5794 81250 6028
rect 82694 5794 82722 6028
rect 78290 5766 78352 5794
rect 79762 5766 79916 5794
rect 76668 800 76696 5766
rect 68020 734 68232 762
rect 68282 0 68338 800
rect 69570 0 69626 800
rect 70858 0 70914 800
rect 74078 0 74134 800
rect 75366 0 75422 800
rect 76654 0 76710 800
rect 78324 762 78352 5766
rect 78508 870 78628 898
rect 78508 762 78536 870
rect 78600 800 78628 870
rect 79888 800 79916 5766
rect 81176 5766 81250 5794
rect 82464 5766 82722 5794
rect 84178 5794 84206 6028
rect 85650 5794 85678 6028
rect 87110 5794 87138 6028
rect 84178 5766 84424 5794
rect 85650 5766 85712 5794
rect 81176 800 81204 5766
rect 82464 800 82492 5766
rect 84396 800 84424 5766
rect 85684 800 85712 5766
rect 86972 5766 87138 5794
rect 88594 5794 88622 6028
rect 90066 5794 90094 6028
rect 91526 5794 91554 6028
rect 92998 5794 93026 6028
rect 88594 5766 88656 5794
rect 90066 5766 90220 5794
rect 86972 800 87000 5766
rect 78324 734 78536 762
rect 78586 0 78642 800
rect 79874 0 79930 800
rect 81162 0 81218 800
rect 82450 0 82506 800
rect 84382 0 84438 800
rect 85670 0 85726 800
rect 86958 0 87014 800
rect 88628 762 88656 5766
rect 88812 870 88932 898
rect 88812 762 88840 870
rect 88904 800 88932 870
rect 90192 800 90220 5766
rect 91480 5766 91554 5794
rect 92768 5766 93026 5794
rect 94482 5794 94510 6028
rect 95954 5794 95982 6028
rect 97414 5794 97442 6028
rect 94482 5766 94728 5794
rect 95954 5766 96016 5794
rect 91480 800 91508 5766
rect 92768 800 92796 5766
rect 94700 800 94728 5766
rect 95988 800 96016 5766
rect 97276 5766 97442 5794
rect 98898 5794 98926 6028
rect 100370 5794 100398 6028
rect 101830 5794 101858 6028
rect 104662 5953 104690 6028
rect 104648 5944 104704 5953
rect 104648 5879 104704 5888
rect 106962 5794 106990 6028
rect 98898 5766 98960 5794
rect 100370 5766 100524 5794
rect 97276 800 97304 5766
rect 88628 734 88840 762
rect 88890 0 88946 800
rect 90178 0 90234 800
rect 91466 0 91522 800
rect 92754 0 92810 800
rect 94686 0 94742 800
rect 95974 0 96030 800
rect 97262 0 97318 800
rect 98932 762 98960 5766
rect 99116 870 99236 898
rect 99116 762 99144 870
rect 99208 800 99236 870
rect 100496 800 100524 5766
rect 101784 5766 101858 5794
rect 106936 5766 106990 5794
rect 109262 5794 109290 6028
rect 111562 5794 111590 6028
rect 109262 5766 109540 5794
rect 101784 800 101812 5766
rect 106936 800 106964 5766
rect 109512 800 109540 5766
rect 111444 5766 111590 5794
rect 113862 5794 113890 6028
rect 116162 5794 116190 6028
rect 113862 5766 114048 5794
rect 111444 800 111472 5766
rect 114020 800 114048 5766
rect 115952 5766 116190 5794
rect 118462 5794 118490 6028
rect 120762 5794 120790 6028
rect 123062 5794 123090 6028
rect 118462 5766 118556 5794
rect 115952 800 115980 5766
rect 118528 800 118556 5766
rect 120736 5766 120790 5794
rect 123036 5766 123090 5794
rect 125362 5794 125390 6028
rect 127662 5794 127690 6028
rect 125362 5766 125456 5794
rect 120460 870 120580 898
rect 120460 800 120488 870
rect 98932 734 99144 762
rect 99194 0 99250 800
rect 100482 0 100538 800
rect 101770 0 101826 800
rect 106922 0 106978 800
rect 109498 0 109554 800
rect 111430 0 111486 800
rect 114006 0 114062 800
rect 115938 0 115994 800
rect 118514 0 118570 800
rect 120446 0 120502 800
rect 120552 762 120580 870
rect 120736 762 120764 5766
rect 123036 800 123064 5766
rect 125428 1306 125456 5766
rect 127544 5766 127690 5794
rect 129962 5794 129990 6028
rect 132262 5794 132290 6028
rect 129962 5766 130148 5794
rect 125428 1278 125640 1306
rect 125612 800 125640 1278
rect 127544 800 127572 5766
rect 130120 800 130148 5766
rect 132236 5766 132290 5794
rect 134562 5794 134590 6028
rect 136862 5794 136890 6028
rect 139162 5794 139190 6028
rect 134562 5766 134656 5794
rect 132236 4706 132264 5766
rect 132052 4678 132264 4706
rect 132052 800 132080 4678
rect 134628 800 134656 5766
rect 136560 5766 136890 5794
rect 139136 5766 139190 5794
rect 141462 5794 141490 6028
rect 143762 5794 143790 6028
rect 141462 5766 141740 5794
rect 136560 800 136588 5766
rect 139136 800 139164 5766
rect 141712 800 141740 5766
rect 143644 5766 143790 5794
rect 146062 5794 146090 6028
rect 148362 5794 148390 6028
rect 146062 5766 146248 5794
rect 143644 800 143672 5766
rect 146220 800 146248 5766
rect 148336 5766 148390 5794
rect 150682 5794 150710 6028
rect 150682 5766 150756 5794
rect 148336 4570 148364 5766
rect 148152 4542 148364 4570
rect 148152 800 148180 4542
rect 150728 800 150756 5766
rect 153304 870 153424 898
rect 153304 800 153332 870
rect 120552 734 120764 762
rect 123022 0 123078 800
rect 125598 0 125654 800
rect 127530 0 127586 800
rect 130106 0 130162 800
rect 132038 0 132094 800
rect 134614 0 134670 800
rect 136546 0 136602 800
rect 139122 0 139178 800
rect 141698 0 141754 800
rect 143630 0 143686 800
rect 146206 0 146262 800
rect 148138 0 148194 800
rect 150714 0 150770 800
rect 153290 0 153346 800
rect 153396 762 153424 870
rect 153580 762 153608 6028
rect 153396 734 153608 762
rect 154316 762 154344 6028
rect 155052 3074 155080 6028
rect 155788 3074 155816 6028
rect 155052 3046 155264 3074
rect 155788 3046 155908 3074
rect 154500 870 154620 898
rect 154500 762 154528 870
rect 154592 800 154620 870
rect 155236 800 155264 3046
rect 155880 800 155908 3046
rect 156524 800 156552 6028
rect 157250 5794 157278 6028
rect 157986 5794 158014 6028
rect 158722 5794 158750 6028
rect 157168 5766 157278 5794
rect 157812 5766 158014 5794
rect 158456 5766 158750 5794
rect 157168 800 157196 5766
rect 157812 800 157840 5766
rect 158456 800 158484 5766
rect 154316 734 154528 762
rect 154578 0 154634 800
rect 155222 0 155278 800
rect 155866 0 155922 800
rect 156510 0 156566 800
rect 157154 0 157210 800
rect 157798 0 157854 800
rect 158442 0 158498 800
rect 159468 762 159496 6028
rect 160204 3074 160232 6028
rect 160940 3074 160968 6028
rect 160204 3046 160416 3074
rect 160940 3046 161060 3074
rect 159652 870 159772 898
rect 159652 762 159680 870
rect 159744 800 159772 870
rect 160388 800 160416 3046
rect 161032 800 161060 3046
rect 161676 800 161704 6028
rect 162402 5794 162430 6028
rect 163138 5794 163166 6028
rect 162320 5766 162430 5794
rect 162964 5766 163166 5794
rect 162320 800 162348 5766
rect 162964 800 162992 5766
rect 163608 870 163728 898
rect 163608 800 163636 870
rect 159468 734 159680 762
rect 159730 0 159786 800
rect 160374 0 160430 800
rect 161018 0 161074 800
rect 161662 0 161718 800
rect 162306 0 162362 800
rect 162950 0 163006 800
rect 163594 0 163650 800
rect 163700 762 163728 870
rect 163884 762 163912 6028
rect 163700 734 163912 762
rect 164620 762 164648 6028
rect 165356 3074 165384 6028
rect 166092 3074 166120 6028
rect 165356 3046 165568 3074
rect 166092 3046 166212 3074
rect 164804 870 164924 898
rect 164804 762 164832 870
rect 164896 800 164924 870
rect 165540 800 165568 3046
rect 166184 800 166212 3046
rect 166828 800 166856 6028
rect 167554 5794 167582 6028
rect 168290 5794 168318 6028
rect 167472 5766 167582 5794
rect 168116 5766 168318 5794
rect 167472 800 167500 5766
rect 168116 800 168144 5766
rect 168760 870 168880 898
rect 168760 800 168788 870
rect 164620 734 164832 762
rect 164882 0 164938 800
rect 165526 0 165582 800
rect 166170 0 166226 800
rect 166814 0 166870 800
rect 167458 0 167514 800
rect 168102 0 168158 800
rect 168746 0 168802 800
rect 168852 762 168880 870
rect 169036 762 169064 6028
rect 168852 734 169064 762
rect 169772 762 169800 6028
rect 170508 3074 170536 6028
rect 171244 3074 171272 6028
rect 170508 3046 170720 3074
rect 171244 3046 171364 3074
rect 169956 870 170076 898
rect 169956 762 169984 870
rect 170048 800 170076 870
rect 170692 800 170720 3046
rect 171336 800 171364 3046
rect 171980 800 172008 6028
rect 172706 5794 172734 6028
rect 173442 5794 173470 6028
rect 172624 5766 172734 5794
rect 173268 5766 173470 5794
rect 172624 800 172652 5766
rect 173268 800 173296 5766
rect 173912 870 174032 898
rect 173912 800 173940 870
rect 169772 734 169984 762
rect 170034 0 170090 800
rect 170678 0 170734 800
rect 171322 0 171378 800
rect 171966 0 172022 800
rect 172610 0 172666 800
rect 173254 0 173310 800
rect 173898 0 173954 800
rect 174004 762 174032 870
rect 174188 762 174216 6028
rect 174004 734 174216 762
rect 174924 762 174952 6028
rect 175660 3074 175688 6028
rect 176396 3074 176424 6028
rect 177122 5953 177150 6028
rect 177108 5944 177164 5953
rect 177108 5879 177164 5888
rect 177858 5794 177886 6028
rect 178594 5794 178622 6028
rect 177776 5766 177886 5794
rect 178420 5766 178622 5794
rect 175660 3046 175872 3074
rect 176396 3046 176516 3074
rect 175108 870 175228 898
rect 175108 762 175136 870
rect 175200 800 175228 870
rect 175844 800 175872 3046
rect 176488 800 176516 3046
rect 177776 800 177804 5766
rect 178420 800 178448 5766
rect 179064 870 179184 898
rect 179064 800 179092 870
rect 174924 734 175136 762
rect 175186 0 175242 800
rect 175830 0 175886 800
rect 176474 0 176530 800
rect 177762 0 177818 800
rect 178406 0 178462 800
rect 179050 0 179106 800
rect 179156 762 179184 870
rect 179340 762 179368 6028
rect 179156 734 179368 762
rect 180076 762 180104 6028
rect 180812 3074 180840 6028
rect 181548 3074 181576 6028
rect 180812 3046 181024 3074
rect 181548 3046 181668 3074
rect 180260 870 180380 898
rect 180260 762 180288 870
rect 180352 800 180380 870
rect 180996 800 181024 3046
rect 181640 800 181668 3046
rect 182284 800 182312 6028
rect 183010 5794 183038 6028
rect 183746 5794 183774 6028
rect 182928 5766 183038 5794
rect 183572 5766 183774 5794
rect 182928 800 182956 5766
rect 183572 800 183600 5766
rect 184216 870 184336 898
rect 184216 800 184244 870
rect 180076 734 180288 762
rect 180338 0 180394 800
rect 180982 0 181038 800
rect 181626 0 181682 800
rect 182270 0 182326 800
rect 182914 0 182970 800
rect 183558 0 183614 800
rect 184202 0 184258 800
rect 184308 762 184336 870
rect 184492 762 184520 6028
rect 184308 734 184520 762
rect 185228 762 185256 6028
rect 185964 3074 185992 6028
rect 186700 3074 186728 6028
rect 185964 3046 186176 3074
rect 186700 3046 186820 3074
rect 185412 870 185532 898
rect 185412 762 185440 870
rect 185504 800 185532 870
rect 186148 800 186176 3046
rect 186792 800 186820 3046
rect 187436 800 187464 6028
rect 188162 5794 188190 6028
rect 188898 5794 188926 6028
rect 188080 5766 188190 5794
rect 188724 5766 188926 5794
rect 188080 800 188108 5766
rect 188724 800 188752 5766
rect 189368 870 189488 898
rect 189368 800 189396 870
rect 185228 734 185440 762
rect 185490 0 185546 800
rect 186134 0 186190 800
rect 186778 0 186834 800
rect 187422 0 187478 800
rect 188066 0 188122 800
rect 188710 0 188766 800
rect 189354 0 189410 800
rect 189460 762 189488 870
rect 189644 762 189672 6028
rect 189460 734 189672 762
rect 190380 762 190408 6028
rect 191116 3074 191144 6028
rect 191116 3046 191328 3074
rect 190564 870 190684 898
rect 190564 762 190592 870
rect 190656 800 190684 870
rect 191300 800 191328 3046
rect 191852 1442 191880 6028
rect 194566 5794 194594 6028
rect 195302 5794 195330 6028
rect 196038 5794 196066 6028
rect 194520 5766 194594 5794
rect 195164 5766 195330 5794
rect 195808 5766 196066 5794
rect 196778 5794 196806 6028
rect 197514 5794 197542 6028
rect 198250 5794 198278 6028
rect 198986 5794 199014 6028
rect 199718 5794 199746 6028
rect 200454 5794 200482 6028
rect 201190 5794 201218 6028
rect 196778 5766 196848 5794
rect 197514 5766 197768 5794
rect 198250 5766 198412 5794
rect 198986 5766 199056 5794
rect 191852 1414 191972 1442
rect 191944 800 191972 1414
rect 194520 800 194548 5766
rect 195164 800 195192 5766
rect 195808 800 195836 5766
rect 190380 734 190592 762
rect 190642 0 190698 800
rect 191286 0 191342 800
rect 191930 0 191986 800
rect 194506 0 194562 800
rect 195150 0 195206 800
rect 195794 0 195850 800
rect 196820 762 196848 5766
rect 197004 870 197124 898
rect 197004 762 197032 870
rect 197096 800 197124 870
rect 197740 800 197768 5766
rect 198384 800 198412 5766
rect 199028 800 199056 5766
rect 199672 5766 199746 5794
rect 200316 5766 200482 5794
rect 200960 5766 201218 5794
rect 201930 5794 201958 6028
rect 202666 5794 202694 6028
rect 203402 5794 203430 6028
rect 204138 5794 204166 6028
rect 204870 5794 204898 6028
rect 205606 5794 205634 6028
rect 206342 5794 206370 6028
rect 201930 5766 202000 5794
rect 202666 5766 202736 5794
rect 203402 5766 203564 5794
rect 204138 5766 204208 5794
rect 199672 800 199700 5766
rect 200316 800 200344 5766
rect 200960 800 200988 5766
rect 196820 734 197032 762
rect 197082 0 197138 800
rect 197726 0 197782 800
rect 198370 0 198426 800
rect 199014 0 199070 800
rect 199658 0 199714 800
rect 200302 0 200358 800
rect 200946 0 201002 800
rect 201972 762 202000 5766
rect 202708 1306 202736 5766
rect 202708 1278 202920 1306
rect 202156 870 202276 898
rect 202156 762 202184 870
rect 202248 800 202276 870
rect 202892 800 202920 1278
rect 203536 800 203564 5766
rect 204180 800 204208 5766
rect 204824 5766 204898 5794
rect 205468 5766 205634 5794
rect 206112 5766 206370 5794
rect 207082 5794 207110 6028
rect 207818 5794 207846 6028
rect 208554 5794 208582 6028
rect 209290 5794 209318 6028
rect 210022 5794 210050 6028
rect 210758 5794 210786 6028
rect 211494 5794 211522 6028
rect 207082 5766 207152 5794
rect 207818 5766 208072 5794
rect 208554 5766 208716 5794
rect 209290 5766 209360 5794
rect 204824 800 204852 5766
rect 205468 800 205496 5766
rect 206112 800 206140 5766
rect 201972 734 202184 762
rect 202234 0 202290 800
rect 202878 0 202934 800
rect 203522 0 203578 800
rect 204166 0 204222 800
rect 204810 0 204866 800
rect 205454 0 205510 800
rect 206098 0 206154 800
rect 207124 762 207152 5766
rect 207308 870 207428 898
rect 207308 762 207336 870
rect 207400 800 207428 870
rect 208044 800 208072 5766
rect 208688 800 208716 5766
rect 209332 800 209360 5766
rect 209976 5766 210050 5794
rect 210620 5766 210786 5794
rect 211264 5766 211522 5794
rect 212234 5794 212262 6028
rect 212970 5794 212998 6028
rect 213706 5794 213734 6028
rect 214442 5794 214470 6028
rect 215174 5794 215202 6028
rect 215910 5794 215938 6028
rect 216646 5794 216674 6028
rect 212234 5766 212304 5794
rect 212970 5766 213224 5794
rect 213706 5766 213868 5794
rect 214442 5766 214512 5794
rect 209976 800 210004 5766
rect 210620 800 210648 5766
rect 211264 800 211292 5766
rect 207124 734 207336 762
rect 207386 0 207442 800
rect 208030 0 208086 800
rect 208674 0 208730 800
rect 209318 0 209374 800
rect 209962 0 210018 800
rect 210606 0 210662 800
rect 211250 0 211306 800
rect 212276 762 212304 5766
rect 212460 870 212580 898
rect 212460 762 212488 870
rect 212552 800 212580 870
rect 213196 800 213224 5766
rect 213840 800 213868 5766
rect 214484 800 214512 5766
rect 215128 5766 215202 5794
rect 215772 5766 215938 5794
rect 216416 5766 216674 5794
rect 217386 5794 217414 6028
rect 218118 5953 218146 6028
rect 218104 5944 218160 5953
rect 218104 5879 218160 5888
rect 218858 5794 218886 6028
rect 219594 5794 219622 6028
rect 220326 5794 220354 6028
rect 221062 5794 221090 6028
rect 221798 5794 221826 6028
rect 217386 5766 217456 5794
rect 218858 5766 219020 5794
rect 219594 5766 219664 5794
rect 215128 800 215156 5766
rect 215772 800 215800 5766
rect 216416 800 216444 5766
rect 212276 734 212488 762
rect 212538 0 212594 800
rect 213182 0 213238 800
rect 213826 0 213882 800
rect 214470 0 214526 800
rect 215114 0 215170 800
rect 215758 0 215814 800
rect 216402 0 216458 800
rect 217428 762 217456 5766
rect 217612 870 217732 898
rect 217612 762 217640 870
rect 217704 800 217732 870
rect 218992 800 219020 5766
rect 219636 800 219664 5766
rect 220280 5766 220354 5794
rect 220924 5766 221090 5794
rect 221568 5766 221826 5794
rect 222538 5794 222566 6028
rect 223274 5794 223302 6028
rect 224010 5794 224038 6028
rect 224746 5794 224774 6028
rect 225478 5794 225506 6028
rect 226214 5794 226242 6028
rect 226950 5794 226978 6028
rect 222538 5766 222608 5794
rect 223274 5766 223528 5794
rect 224010 5766 224172 5794
rect 224746 5766 224816 5794
rect 220280 800 220308 5766
rect 220924 800 220952 5766
rect 221568 800 221596 5766
rect 217428 734 217640 762
rect 217690 0 217746 800
rect 218978 0 219034 800
rect 219622 0 219678 800
rect 220266 0 220322 800
rect 220910 0 220966 800
rect 221554 0 221610 800
rect 222580 762 222608 5766
rect 222764 870 222884 898
rect 222764 762 222792 870
rect 222856 800 222884 870
rect 223500 800 223528 5766
rect 224144 800 224172 5766
rect 224788 800 224816 5766
rect 225432 5766 225506 5794
rect 226076 5766 226242 5794
rect 226720 5766 226978 5794
rect 227690 5794 227718 6028
rect 228426 5794 228454 6028
rect 229162 5794 229190 6028
rect 229898 5794 229926 6028
rect 230630 5794 230658 6028
rect 231366 5794 231394 6028
rect 232102 5794 232130 6028
rect 227690 5766 227760 5794
rect 228426 5766 228680 5794
rect 229162 5766 229324 5794
rect 229898 5766 229968 5794
rect 225432 800 225460 5766
rect 226076 800 226104 5766
rect 226720 800 226748 5766
rect 222580 734 222792 762
rect 222842 0 222898 800
rect 223486 0 223542 800
rect 224130 0 224186 800
rect 224774 0 224830 800
rect 225418 0 225474 800
rect 226062 0 226118 800
rect 226706 0 226762 800
rect 227732 762 227760 5766
rect 227916 870 228036 898
rect 227916 762 227944 870
rect 228008 800 228036 870
rect 228652 800 228680 5766
rect 229296 800 229324 5766
rect 229940 800 229968 5766
rect 230584 5766 230658 5794
rect 231228 5766 231394 5794
rect 231872 5766 232130 5794
rect 232842 5794 232870 6028
rect 235598 5794 235626 6028
rect 236334 5794 236362 6028
rect 232842 5766 232912 5794
rect 235598 5766 235764 5794
rect 236334 5766 236408 5794
rect 230584 800 230612 5766
rect 231228 800 231256 5766
rect 231872 800 231900 5766
rect 227732 734 227944 762
rect 227994 0 228050 800
rect 228638 0 228694 800
rect 229282 0 229338 800
rect 229926 0 229982 800
rect 230570 0 230626 800
rect 231214 0 231270 800
rect 231858 0 231914 800
rect 232884 762 232912 5766
rect 233068 870 233188 898
rect 233068 762 233096 870
rect 233160 800 233188 870
rect 235736 800 235764 5766
rect 236380 800 236408 5766
rect 237024 800 237052 6028
rect 237760 3074 237788 6028
rect 237668 3046 237788 3074
rect 237668 800 237696 3046
rect 238496 1714 238524 6028
rect 238312 1686 238524 1714
rect 238312 800 238340 1686
rect 238956 870 239076 898
rect 238956 800 238984 870
rect 232884 734 233096 762
rect 233146 0 233202 800
rect 235722 0 235778 800
rect 236366 0 236422 800
rect 237010 0 237066 800
rect 237654 0 237710 800
rect 238298 0 238354 800
rect 238942 0 238998 800
rect 239048 762 239076 870
rect 239232 762 239260 6028
rect 240014 5794 240042 6028
rect 240750 5794 240778 6028
rect 240014 5766 240088 5794
rect 240750 5766 240916 5794
rect 240060 1306 240088 5766
rect 240060 1278 240272 1306
rect 240244 800 240272 1278
rect 240888 800 240916 5766
rect 241440 1306 241468 6028
rect 241440 1278 241560 1306
rect 241532 800 241560 1278
rect 242176 800 242204 6028
rect 242912 5658 242940 6028
rect 242820 5630 242940 5658
rect 242820 800 242848 5630
rect 243648 1714 243676 6028
rect 244384 5658 244412 6028
rect 245166 5794 245194 6028
rect 245902 5794 245930 6028
rect 246638 5794 246666 6028
rect 245166 5766 245424 5794
rect 245902 5766 246068 5794
rect 246638 5766 246712 5794
rect 243464 1686 243676 1714
rect 244108 5630 244412 5658
rect 243464 800 243492 1686
rect 244108 800 244136 5630
rect 245396 800 245424 5766
rect 246040 800 246068 5766
rect 246684 800 246712 5766
rect 247328 800 247356 6028
rect 248064 3074 248092 6028
rect 247972 3046 248092 3074
rect 247972 800 248000 3046
rect 248800 1714 248828 6028
rect 248616 1686 248828 1714
rect 248616 800 248644 1686
rect 249260 870 249380 898
rect 249260 800 249288 870
rect 239048 734 239260 762
rect 240230 0 240286 800
rect 240874 0 240930 800
rect 241518 0 241574 800
rect 242162 0 242218 800
rect 242806 0 242862 800
rect 243450 0 243506 800
rect 244094 0 244150 800
rect 245382 0 245438 800
rect 246026 0 246082 800
rect 246670 0 246726 800
rect 247314 0 247370 800
rect 247958 0 248014 800
rect 248602 0 248658 800
rect 249246 0 249302 800
rect 249352 762 249380 870
rect 249536 762 249564 6028
rect 250318 5794 250346 6028
rect 251054 5794 251082 6028
rect 251790 5794 251818 6028
rect 250318 5766 250576 5794
rect 251054 5766 251128 5794
rect 251790 5766 251864 5794
rect 250548 800 250576 5766
rect 251100 1306 251128 5766
rect 251100 1278 251220 1306
rect 251192 800 251220 1278
rect 251836 800 251864 5766
rect 252480 800 252508 6028
rect 253216 3074 253244 6028
rect 253952 5658 253980 6028
rect 253124 3046 253244 3074
rect 253768 5630 253980 5658
rect 253124 800 253152 3046
rect 253768 800 253796 5630
rect 254412 870 254532 898
rect 254412 800 254440 870
rect 249352 734 249564 762
rect 250534 0 250590 800
rect 251178 0 251234 800
rect 251822 0 251878 800
rect 252466 0 252522 800
rect 253110 0 253166 800
rect 253754 0 253810 800
rect 254398 0 254454 800
rect 254504 762 254532 870
rect 254688 762 254716 6028
rect 255470 5794 255498 6028
rect 256206 5794 256234 6028
rect 256942 5794 256970 6028
rect 255470 5766 255728 5794
rect 256206 5766 256372 5794
rect 256942 5766 257016 5794
rect 255700 800 255728 5766
rect 256344 800 256372 5766
rect 256988 800 257016 5766
rect 257632 800 257660 6028
rect 258368 3074 258396 6028
rect 259150 5953 259178 6028
rect 259136 5944 259192 5953
rect 259136 5879 259192 5888
rect 258276 3046 258396 3074
rect 258276 800 258304 3046
rect 259564 870 259684 898
rect 259564 800 259592 870
rect 254504 734 254716 762
rect 255686 0 255742 800
rect 256330 0 256386 800
rect 256974 0 257030 800
rect 257618 0 257674 800
rect 258262 0 258318 800
rect 259550 0 259606 800
rect 259656 762 259684 870
rect 259840 762 259868 6028
rect 260622 5794 260650 6028
rect 261358 5794 261386 6028
rect 262094 5794 262122 6028
rect 260622 5766 260696 5794
rect 261358 5766 261524 5794
rect 262094 5766 262168 5794
rect 260668 1306 260696 5766
rect 260668 1278 260880 1306
rect 260852 800 260880 1278
rect 261496 800 261524 5766
rect 262140 800 262168 5766
rect 262784 800 262812 6028
rect 263520 3074 263548 6028
rect 263428 3046 263548 3074
rect 263428 800 263456 3046
rect 264256 1714 264284 6028
rect 264992 5658 265020 6028
rect 265774 5794 265802 6028
rect 266510 5794 266538 6028
rect 267246 5794 267274 6028
rect 265774 5766 266032 5794
rect 266510 5766 266676 5794
rect 267246 5766 267320 5794
rect 264072 1686 264284 1714
rect 264716 5630 265020 5658
rect 264072 800 264100 1686
rect 264716 800 264744 5630
rect 266004 800 266032 5766
rect 266648 800 266676 5766
rect 267292 800 267320 5766
rect 267936 800 267964 6028
rect 268672 3074 268700 6028
rect 268580 3046 268700 3074
rect 268580 800 268608 3046
rect 269408 1714 269436 6028
rect 269224 1686 269436 1714
rect 269224 800 269252 1686
rect 269868 870 269988 898
rect 269868 800 269896 870
rect 259656 734 259868 762
rect 260838 0 260894 800
rect 261482 0 261538 800
rect 262126 0 262182 800
rect 262770 0 262826 800
rect 263414 0 263470 800
rect 264058 0 264114 800
rect 264702 0 264758 800
rect 265990 0 266046 800
rect 266634 0 266690 800
rect 267278 0 267334 800
rect 267922 0 267978 800
rect 268566 0 268622 800
rect 269210 0 269266 800
rect 269854 0 269910 800
rect 269960 762 269988 870
rect 270144 762 270172 6028
rect 270926 5794 270954 6028
rect 271662 5794 271690 6028
rect 272398 5794 272426 6028
rect 270926 5766 271184 5794
rect 271662 5766 271828 5794
rect 272398 5766 272472 5794
rect 271156 800 271184 5766
rect 271800 800 271828 5766
rect 272444 800 272472 5766
rect 273088 800 273116 6028
rect 273824 3074 273852 6028
rect 276570 5953 276598 6028
rect 276556 5944 276612 5953
rect 276556 5879 276612 5888
rect 273732 3046 273852 3074
rect 273732 800 273760 3046
rect 278700 1306 278728 6028
rect 278700 1278 278912 1306
rect 278884 800 278912 1278
rect 280816 800 280844 6028
rect 282918 5794 282946 6028
rect 282748 5766 282946 5794
rect 282748 800 282776 5766
rect 269960 734 270172 762
rect 271142 0 271198 800
rect 271786 0 271842 800
rect 272430 0 272486 800
rect 273074 0 273130 800
rect 273718 0 273774 800
rect 278870 0 278926 800
rect 280802 0 280858 800
rect 282734 0 282790 800
rect 285048 762 285076 6028
rect 287164 3074 287192 6028
rect 289266 5794 289294 6028
rect 291382 5794 291410 6028
rect 289188 5766 289294 5794
rect 291120 5766 291410 5794
rect 287164 3046 287284 3074
rect 285232 870 285352 898
rect 285232 762 285260 870
rect 285324 800 285352 870
rect 287256 800 287284 3046
rect 289188 800 289216 5766
rect 291120 800 291148 5766
rect 293512 3074 293540 6028
rect 293512 3046 293724 3074
rect 293696 800 293724 3046
rect 295628 800 295656 6028
rect 297730 5794 297758 6028
rect 297560 5766 297758 5794
rect 297560 800 297588 5766
rect 285048 734 285260 762
rect 285310 0 285366 800
rect 287242 0 287298 800
rect 289174 0 289230 800
rect 291106 0 291162 800
rect 293682 0 293738 800
rect 295614 0 295670 800
rect 297546 0 297602 800
rect 299860 762 299888 6028
rect 301976 1170 302004 6028
rect 304078 5794 304106 6028
rect 304000 5766 304106 5794
rect 301976 1142 302096 1170
rect 300044 870 300164 898
rect 300044 762 300072 870
rect 300136 800 300164 870
rect 302068 800 302096 1142
rect 304000 800 304028 5766
rect 305932 870 306052 898
rect 305932 800 305960 870
rect 299860 734 300072 762
rect 300122 0 300178 800
rect 302054 0 302110 800
rect 303986 0 304042 800
rect 305918 0 305974 800
rect 306024 762 306052 870
rect 306208 762 306236 6028
rect 308324 3074 308352 6028
rect 308324 3046 308536 3074
rect 308508 800 308536 3046
rect 310440 800 310468 6028
rect 312542 5794 312570 6028
rect 312372 5766 312570 5794
rect 312372 800 312400 5766
rect 306024 734 306236 762
rect 308494 0 308550 800
rect 310426 0 310482 800
rect 312358 0 312414 800
rect 314672 762 314700 6028
rect 316788 3074 316816 6028
rect 318890 5794 318918 6028
rect 321570 5794 321598 6028
rect 318812 5766 318918 5794
rect 321388 5766 321598 5794
rect 316788 3046 316908 3074
rect 314856 870 314976 898
rect 314856 762 314884 870
rect 314948 800 314976 870
rect 316880 800 316908 3046
rect 318812 800 318840 5766
rect 321388 800 321416 5766
rect 322032 870 322152 898
rect 322032 800 322060 870
rect 314672 734 314884 762
rect 314934 0 314990 800
rect 316866 0 316922 800
rect 318798 0 318854 800
rect 321374 0 321430 800
rect 322018 0 322074 800
rect 322124 762 322152 870
rect 322308 762 322336 6028
rect 322124 734 322336 762
rect 323044 762 323072 6028
rect 323780 3074 323808 6028
rect 324516 3074 324544 6028
rect 323780 3046 323992 3074
rect 324516 3046 324636 3074
rect 323228 870 323348 898
rect 323228 762 323256 870
rect 323320 800 323348 870
rect 323964 800 323992 3046
rect 324608 800 324636 3046
rect 325252 800 325280 6028
rect 325986 5794 326014 6028
rect 326722 5794 326750 6028
rect 325896 5766 326014 5794
rect 326540 5766 326750 5794
rect 325896 800 325924 5766
rect 326540 800 326568 5766
rect 327184 870 327304 898
rect 327184 800 327212 870
rect 323044 734 323256 762
rect 323306 0 323362 800
rect 323950 0 324006 800
rect 324594 0 324650 800
rect 325238 0 325294 800
rect 325882 0 325938 800
rect 326526 0 326582 800
rect 327170 0 327226 800
rect 327276 762 327304 870
rect 327460 762 327488 6028
rect 327276 734 327488 762
rect 328196 762 328224 6028
rect 328932 3074 328960 6028
rect 329668 3074 329696 6028
rect 328932 3046 329144 3074
rect 329668 3046 329788 3074
rect 328380 870 328500 898
rect 328380 762 328408 870
rect 328472 800 328500 870
rect 329116 800 329144 3046
rect 329760 800 329788 3046
rect 330404 800 330432 6028
rect 331138 5794 331166 6028
rect 331874 5794 331902 6028
rect 332610 5794 332638 6028
rect 331048 5766 331166 5794
rect 331692 5766 331902 5794
rect 332336 5766 332638 5794
rect 331048 800 331076 5766
rect 331692 800 331720 5766
rect 332336 800 332364 5766
rect 328196 734 328408 762
rect 328458 0 328514 800
rect 329102 0 329158 800
rect 329746 0 329802 800
rect 330390 0 330446 800
rect 331034 0 331090 800
rect 331678 0 331734 800
rect 332322 0 332378 800
rect 333348 762 333376 6028
rect 334084 3074 334112 6028
rect 334820 3074 334848 6028
rect 334084 3046 334296 3074
rect 334820 3046 334940 3074
rect 333532 870 333652 898
rect 333532 762 333560 870
rect 333624 800 333652 870
rect 334268 800 334296 3046
rect 334912 800 334940 3046
rect 335556 800 335584 6028
rect 336290 5794 336318 6028
rect 337026 5794 337054 6028
rect 336200 5766 336318 5794
rect 336844 5766 337054 5794
rect 336200 800 336228 5766
rect 336844 800 336872 5766
rect 337488 870 337608 898
rect 337488 800 337516 870
rect 333348 734 333560 762
rect 333610 0 333666 800
rect 334254 0 334310 800
rect 334898 0 334954 800
rect 335542 0 335598 800
rect 336186 0 336242 800
rect 336830 0 336886 800
rect 337474 0 337530 800
rect 337580 762 337608 870
rect 337764 762 337792 6028
rect 337580 734 337792 762
rect 338500 762 338528 6028
rect 339236 3074 339264 6028
rect 339972 3074 340000 6028
rect 339236 3046 339448 3074
rect 339972 3046 340092 3074
rect 338684 870 338804 898
rect 338684 762 338712 870
rect 338776 800 338804 870
rect 339420 800 339448 3046
rect 340064 800 340092 3046
rect 340708 800 340736 6028
rect 341442 5794 341470 6028
rect 342178 5794 342206 6028
rect 341352 5766 341470 5794
rect 341996 5766 342206 5794
rect 341352 800 341380 5766
rect 341996 800 342024 5766
rect 342640 870 342760 898
rect 342640 800 342668 870
rect 338500 734 338712 762
rect 338762 0 338818 800
rect 339406 0 339462 800
rect 340050 0 340106 800
rect 340694 0 340750 800
rect 341338 0 341394 800
rect 341982 0 342038 800
rect 342626 0 342682 800
rect 342732 762 342760 870
rect 342916 762 342944 6028
rect 342732 734 342944 762
rect 343652 762 343680 6028
rect 344388 3074 344416 6028
rect 345124 5953 345152 6028
rect 345110 5944 345166 5953
rect 345110 5879 345166 5888
rect 344388 3046 344600 3074
rect 343836 870 343956 898
rect 343836 762 343864 870
rect 343928 800 343956 870
rect 344572 800 344600 3046
rect 345860 800 345888 6028
rect 346594 5794 346622 6028
rect 347330 5794 347358 6028
rect 346504 5766 346622 5794
rect 347148 5766 347358 5794
rect 346504 800 346532 5766
rect 347148 800 347176 5766
rect 347792 870 347912 898
rect 347792 800 347820 870
rect 343652 734 343864 762
rect 343914 0 343970 800
rect 344558 0 344614 800
rect 345846 0 345902 800
rect 346490 0 346546 800
rect 347134 0 347190 800
rect 347778 0 347834 800
rect 347884 762 347912 870
rect 348068 762 348096 6028
rect 347884 734 348096 762
rect 348804 762 348832 6028
rect 349540 3074 349568 6028
rect 350276 3074 350304 6028
rect 349540 3046 349752 3074
rect 350276 3046 350396 3074
rect 348988 870 349108 898
rect 348988 762 349016 870
rect 349080 800 349108 870
rect 349724 800 349752 3046
rect 350368 800 350396 3046
rect 351012 800 351040 6028
rect 351746 5794 351774 6028
rect 352482 5794 352510 6028
rect 351656 5766 351774 5794
rect 352300 5766 352510 5794
rect 351656 800 351684 5766
rect 352300 800 352328 5766
rect 352944 870 353064 898
rect 352944 800 352972 870
rect 348804 734 349016 762
rect 349066 0 349122 800
rect 349710 0 349766 800
rect 350354 0 350410 800
rect 350998 0 351054 800
rect 351642 0 351698 800
rect 352286 0 352342 800
rect 352930 0 352986 800
rect 353036 762 353064 870
rect 353220 762 353248 6028
rect 353036 734 353248 762
rect 353956 762 353984 6028
rect 354692 3074 354720 6028
rect 355428 3074 355456 6028
rect 354692 3046 354904 3074
rect 355428 3046 355548 3074
rect 354140 870 354260 898
rect 354140 762 354168 870
rect 354232 800 354260 870
rect 354876 800 354904 3046
rect 355520 800 355548 3046
rect 356164 800 356192 6028
rect 356898 5794 356926 6028
rect 357634 5794 357662 6028
rect 356808 5766 356926 5794
rect 357452 5766 357662 5794
rect 356808 800 356836 5766
rect 357452 800 357480 5766
rect 358096 870 358216 898
rect 358096 800 358124 870
rect 353956 734 354168 762
rect 354218 0 354274 800
rect 354862 0 354918 800
rect 355506 0 355562 800
rect 356150 0 356206 800
rect 356794 0 356850 800
rect 357438 0 357494 800
rect 358082 0 358138 800
rect 358188 762 358216 870
rect 358372 762 358400 6028
rect 358188 734 358400 762
rect 359108 762 359136 6028
rect 359844 3074 359872 6028
rect 362386 5794 362414 6028
rect 363478 5794 363506 6028
rect 364582 5794 364610 6028
rect 362386 5766 362632 5794
rect 359844 3046 360056 3074
rect 359292 870 359412 898
rect 359292 762 359320 870
rect 359384 800 359412 870
rect 360028 800 360056 3046
rect 362604 800 362632 5766
rect 363248 5766 363506 5794
rect 364536 5766 364610 5794
rect 365698 5794 365726 6028
rect 366802 5794 366830 6028
rect 367894 5794 367922 6028
rect 365698 5766 365852 5794
rect 366802 5766 366864 5794
rect 363248 800 363276 5766
rect 364536 800 364564 5766
rect 365824 800 365852 5766
rect 359108 734 359320 762
rect 359370 0 359426 800
rect 360014 0 360070 800
rect 362590 0 362646 800
rect 363234 0 363290 800
rect 364522 0 364578 800
rect 365810 0 365866 800
rect 366836 762 366864 5766
rect 367756 5766 367922 5794
rect 369010 5794 369038 6028
rect 370114 5794 370142 6028
rect 371206 5794 371234 6028
rect 372310 5794 372338 6028
rect 369010 5766 369072 5794
rect 370114 5766 370360 5794
rect 367020 870 367140 898
rect 367020 762 367048 870
rect 367112 800 367140 870
rect 367756 800 367784 5766
rect 369044 800 369072 5766
rect 370332 800 370360 5766
rect 370976 5766 371234 5794
rect 372264 5766 372338 5794
rect 373426 5794 373454 6028
rect 374530 5794 374558 6028
rect 375622 5794 375650 6028
rect 373426 5766 373580 5794
rect 374530 5766 374592 5794
rect 370976 800 371004 5766
rect 372264 800 372292 5766
rect 373552 800 373580 5766
rect 366836 734 367048 762
rect 367098 0 367154 800
rect 367742 0 367798 800
rect 369030 0 369086 800
rect 370318 0 370374 800
rect 370962 0 371018 800
rect 372250 0 372306 800
rect 373538 0 373594 800
rect 374564 762 374592 5766
rect 375484 5766 375650 5794
rect 376738 5794 376766 6028
rect 377842 5794 377870 6028
rect 378934 5953 378962 6028
rect 378920 5944 378976 5953
rect 378920 5879 378976 5888
rect 380050 5794 380078 6028
rect 381154 5794 381182 6028
rect 382258 5794 382286 6028
rect 383362 5817 383390 6028
rect 383348 5808 383404 5817
rect 376738 5766 376800 5794
rect 377842 5766 378088 5794
rect 380050 5766 380112 5794
rect 381154 5766 381216 5794
rect 382258 5766 382320 5794
rect 374748 870 374868 898
rect 374748 762 374776 870
rect 374840 800 374868 870
rect 375484 800 375512 5766
rect 376772 800 376800 5766
rect 378060 800 378088 5766
rect 374564 734 374776 762
rect 374826 0 374882 800
rect 375470 0 375526 800
rect 376758 0 376814 800
rect 378046 0 378102 800
rect 380084 377 380112 5766
rect 380070 368 380126 377
rect 380070 303 380126 312
rect 381188 241 381216 5766
rect 382292 513 382320 5766
rect 384466 5794 384494 6028
rect 385570 5794 385598 6028
rect 386674 5794 386702 6028
rect 387778 5794 387806 6028
rect 388882 5794 388910 6028
rect 389986 5794 390014 6028
rect 391090 5794 391118 6028
rect 392194 5794 392222 6028
rect 392858 5808 392914 5817
rect 384466 5766 384528 5794
rect 385570 5766 385632 5794
rect 386674 5766 386736 5794
rect 387778 5766 388484 5794
rect 388882 5766 388944 5794
rect 389986 5766 390048 5794
rect 391090 5766 391152 5794
rect 392194 5766 392256 5794
rect 383348 5743 383404 5752
rect 384500 1193 384528 5766
rect 385604 1329 385632 5766
rect 385590 1320 385646 1329
rect 385590 1255 385646 1264
rect 386418 1320 386474 1329
rect 386418 1255 386474 1264
rect 384486 1184 384542 1193
rect 384486 1119 384542 1128
rect 386432 800 386460 1255
rect 386708 1057 386736 5766
rect 387706 1184 387762 1193
rect 387706 1119 387762 1128
rect 386694 1048 386750 1057
rect 386694 983 386750 992
rect 386984 870 387104 898
rect 382278 504 382334 513
rect 382278 439 382334 448
rect 381174 232 381230 241
rect 381174 167 381230 176
rect 386418 0 386474 800
rect 386984 241 387012 870
rect 387076 800 387104 870
rect 387720 800 387748 1119
rect 388272 870 388392 898
rect 386970 232 387026 241
rect 386970 167 387026 176
rect 387062 0 387118 800
rect 387706 0 387762 800
rect 388272 513 388300 870
rect 388364 800 388392 870
rect 388258 504 388314 513
rect 388258 439 388314 448
rect 388350 0 388406 800
rect 388456 762 388484 5766
rect 388916 1329 388944 5766
rect 388902 1320 388958 1329
rect 388902 1255 388958 1264
rect 389638 1320 389694 1329
rect 389638 1255 389694 1264
rect 388916 870 389036 898
rect 388916 762 388944 870
rect 389008 800 389036 870
rect 389652 800 389680 1255
rect 388456 734 388944 762
rect 388994 0 389050 800
rect 389638 0 389694 800
rect 390020 762 390048 5766
rect 390926 1048 390982 1057
rect 390926 983 390982 992
rect 390204 870 390324 898
rect 390204 762 390232 870
rect 390296 800 390324 870
rect 390940 800 390968 983
rect 390020 734 390232 762
rect 390282 0 390338 800
rect 390926 0 390982 800
rect 391124 762 391152 5766
rect 391492 870 391612 898
rect 391492 762 391520 870
rect 391584 800 391612 870
rect 392228 800 392256 5766
rect 393298 5794 393326 6028
rect 394402 5794 394430 6028
rect 395494 5794 395522 6028
rect 393298 5766 393544 5794
rect 394402 5766 394464 5794
rect 392858 5743 392914 5752
rect 392872 800 392900 5743
rect 393516 800 393544 5766
rect 394068 870 394188 898
rect 391124 734 391520 762
rect 391570 0 391626 800
rect 392214 0 392270 800
rect 392858 0 392914 800
rect 393502 0 393558 800
rect 394068 377 394096 870
rect 394160 800 394188 870
rect 394054 368 394110 377
rect 394054 303 394110 312
rect 394146 0 394202 800
rect 394436 762 394464 5766
rect 395448 5766 395522 5794
rect 396610 5794 396638 6028
rect 397714 5794 397742 6028
rect 398806 5794 398834 6028
rect 396610 5766 396764 5794
rect 397714 5766 397776 5794
rect 394712 870 394832 898
rect 394712 762 394740 870
rect 394804 800 394832 870
rect 395448 800 395476 5766
rect 396736 800 396764 5766
rect 394436 734 394740 762
rect 394790 0 394846 800
rect 395434 0 395490 800
rect 396722 0 396778 800
rect 397748 762 397776 5766
rect 398668 5766 398834 5794
rect 399922 5794 399950 6028
rect 401026 5794 401054 6028
rect 403386 5794 403414 6028
rect 404766 5794 404794 6028
rect 399922 5766 399984 5794
rect 401026 5766 401272 5794
rect 397932 870 398052 898
rect 397932 762 397960 870
rect 398024 800 398052 870
rect 398668 800 398696 5766
rect 399956 800 399984 5766
rect 401244 800 401272 5766
rect 403360 5766 403414 5794
rect 404740 5766 404794 5794
rect 406146 5794 406174 6028
rect 407526 5794 407554 6028
rect 408906 5794 408934 6028
rect 410286 5794 410314 6028
rect 411666 5794 411694 6028
rect 413046 5794 413074 6028
rect 414426 5953 414454 6028
rect 414412 5944 414468 5953
rect 414412 5879 414468 5888
rect 406146 5766 406424 5794
rect 407526 5766 407712 5794
rect 408906 5766 409000 5794
rect 403360 4570 403388 5766
rect 403176 4542 403388 4570
rect 403176 800 403204 4542
rect 404464 870 404584 898
rect 404464 800 404492 870
rect 397748 734 397960 762
rect 398010 0 398066 800
rect 398654 0 398710 800
rect 399942 0 399998 800
rect 401230 0 401286 800
rect 403162 0 403218 800
rect 404450 0 404506 800
rect 404556 762 404584 870
rect 404740 762 404768 5766
rect 406396 800 406424 5766
rect 407684 800 407712 5766
rect 408972 800 409000 5766
rect 410260 5766 410314 5794
rect 411548 5766 411694 5794
rect 413020 5766 413074 5794
rect 415806 5794 415834 6028
rect 417186 5794 417214 6028
rect 418566 5794 418594 6028
rect 419946 5794 419974 6028
rect 421326 5794 421354 6028
rect 422706 5794 422734 6028
rect 424086 5794 424114 6028
rect 415806 5766 416084 5794
rect 417186 5766 417372 5794
rect 418566 5766 418660 5794
rect 410260 800 410288 5766
rect 411548 800 411576 5766
rect 413020 4706 413048 5766
rect 412836 4678 413048 4706
rect 412836 800 412864 4678
rect 416056 800 416084 5766
rect 417344 800 417372 5766
rect 418632 800 418660 5766
rect 419920 5766 419974 5794
rect 421208 5766 421354 5794
rect 422680 5766 422734 5794
rect 424060 5766 424114 5794
rect 425466 5794 425494 6028
rect 426846 5794 426874 6028
rect 428226 5794 428254 6028
rect 429606 5794 429634 6028
rect 430986 5794 431014 6028
rect 432366 5794 432394 6028
rect 433746 5794 433774 6028
rect 425466 5766 425744 5794
rect 426846 5766 427032 5794
rect 428226 5766 428320 5794
rect 419920 800 419948 5766
rect 421208 800 421236 5766
rect 422680 4570 422708 5766
rect 422496 4542 422708 4570
rect 422496 800 422524 4542
rect 423784 870 423904 898
rect 423784 800 423812 870
rect 404556 734 404768 762
rect 406382 0 406438 800
rect 407670 0 407726 800
rect 408958 0 409014 800
rect 410246 0 410302 800
rect 411534 0 411590 800
rect 412822 0 412878 800
rect 416042 0 416098 800
rect 417330 0 417386 800
rect 418618 0 418674 800
rect 419906 0 419962 800
rect 421194 0 421250 800
rect 422482 0 422538 800
rect 423770 0 423826 800
rect 423876 762 423904 870
rect 424060 762 424088 5766
rect 425716 800 425744 5766
rect 427004 800 427032 5766
rect 428292 800 428320 5766
rect 429580 5766 429634 5794
rect 430868 5766 431014 5794
rect 432340 5766 432394 5794
rect 433720 5766 433774 5794
rect 435126 5794 435154 6028
rect 436506 5794 436534 6028
rect 437886 5794 437914 6028
rect 439266 5794 439294 6028
rect 440646 5794 440674 6028
rect 442026 5794 442054 6028
rect 444478 5953 444506 6028
rect 444464 5944 444520 5953
rect 444464 5879 444520 5888
rect 435126 5766 435404 5794
rect 436506 5766 436692 5794
rect 437886 5766 437980 5794
rect 429580 800 429608 5766
rect 430868 800 430896 5766
rect 432340 4706 432368 5766
rect 432156 4678 432368 4706
rect 432156 800 432184 4678
rect 433444 870 433564 898
rect 433444 800 433472 870
rect 423876 734 424088 762
rect 425702 0 425758 800
rect 426990 0 427046 800
rect 428278 0 428334 800
rect 429566 0 429622 800
rect 430854 0 430910 800
rect 432142 0 432198 800
rect 433430 0 433486 800
rect 433536 762 433564 870
rect 433720 762 433748 5766
rect 435376 800 435404 5766
rect 436664 800 436692 5766
rect 437952 800 437980 5766
rect 439240 5766 439294 5794
rect 440528 5766 440674 5794
rect 441816 5766 442054 5794
rect 439240 800 439268 5766
rect 440528 800 440556 5766
rect 441816 800 441844 5766
rect 433536 734 433748 762
rect 435362 0 435418 800
rect 436650 0 436706 800
rect 437938 0 437994 800
rect 439226 0 439282 800
rect 440514 0 440570 800
rect 441802 0 441858 800
rect 446048 762 446076 6028
rect 446232 870 446352 898
rect 446232 762 446260 870
rect 446324 800 446352 870
rect 447612 800 447640 6028
rect 448900 870 449020 898
rect 448900 800 448928 870
rect 446048 734 446260 762
rect 446310 0 446366 800
rect 447598 0 447654 800
rect 448886 0 448942 800
rect 448992 762 449020 870
rect 449176 762 449204 6028
rect 450740 3074 450768 6028
rect 452298 5794 452326 6028
rect 452120 5766 452326 5794
rect 450740 3046 450860 3074
rect 450832 800 450860 3046
rect 452120 800 452148 5766
rect 453868 1306 453896 6028
rect 455426 5794 455454 6028
rect 455340 5766 455454 5794
rect 453868 1278 454080 1306
rect 454052 800 454080 1278
rect 455340 800 455368 5766
rect 448992 734 449204 762
rect 450818 0 450874 800
rect 452106 0 452162 800
rect 454038 0 454094 800
rect 455326 0 455382 800
rect 456996 762 457024 6028
rect 457180 870 457300 898
rect 457180 762 457208 870
rect 457272 800 457300 870
rect 458560 800 458588 6028
rect 459848 870 459968 898
rect 459848 800 459876 870
rect 456996 734 457208 762
rect 457258 0 457314 800
rect 458546 0 458602 800
rect 459834 0 459890 800
rect 459940 762 459968 870
rect 460124 762 460152 6028
rect 461688 3074 461716 6028
rect 463246 5794 463274 6028
rect 463068 5766 463274 5794
rect 461688 3046 461808 3074
rect 461780 800 461808 3046
rect 463068 800 463096 5766
rect 464816 3074 464844 6028
rect 466374 5794 466402 6028
rect 466288 5766 466402 5794
rect 464816 3046 465028 3074
rect 465000 800 465028 3046
rect 466288 800 466316 5766
rect 459940 734 460152 762
rect 461766 0 461822 800
rect 463054 0 463110 800
rect 464986 0 465042 800
rect 466274 0 466330 800
rect 467944 762 467972 6028
rect 468128 870 468248 898
rect 468128 762 468156 870
rect 468220 800 468248 870
rect 469508 800 469536 6028
rect 470796 870 470916 898
rect 470796 800 470824 870
rect 467944 734 468156 762
rect 468206 0 468262 800
rect 469494 0 469550 800
rect 470782 0 470838 800
rect 470888 762 470916 870
rect 471072 762 471100 6028
rect 472636 3074 472664 6028
rect 474194 5794 474222 6028
rect 474016 5766 474222 5794
rect 472636 3046 472756 3074
rect 472728 800 472756 3046
rect 474016 800 474044 5766
rect 475764 3074 475792 6028
rect 475764 3046 475976 3074
rect 475948 800 475976 3046
rect 470888 734 471100 762
rect 472714 0 472770 800
rect 474002 0 474058 800
rect 475934 0 475990 800
<< via2 >>
rect 9126 747088 9182 747144
rect 9770 746272 9826 746328
rect 8298 745456 8354 745512
rect 10414 743008 10470 743064
rect 11702 743824 11758 743880
rect 12990 746544 13046 746600
rect 13450 744912 13506 744968
rect 12162 741920 12218 741976
rect 14738 742736 14794 742792
rect 15566 741648 15622 741704
rect 10966 739200 11022 739256
rect 18142 746000 18198 746056
rect 18602 745184 18658 745240
rect 19430 744096 19486 744152
rect 17314 743552 17370 743608
rect 20442 755656 20498 755712
rect 20074 755384 20130 755440
rect 19890 742192 19946 742248
rect 16118 740560 16174 740616
rect 20258 754840 20314 754896
rect 20166 749536 20222 749592
rect 20074 740288 20130 740344
rect 16762 739744 16818 739800
rect 20350 754024 20406 754080
rect 20258 744640 20314 744696
rect 20442 752664 20498 752720
rect 20350 741104 20406 741160
rect 20534 745728 20590 745784
rect 21454 753480 21510 753536
rect 21178 749400 21234 749456
rect 21086 744390 21142 744446
rect 22282 753480 22338 753536
rect 22006 749536 22062 749592
rect 23570 754840 23626 754896
rect 25870 748584 25926 748640
rect 26790 755792 26846 755848
rect 27986 754976 28042 755032
rect 30010 752664 30066 752720
rect 31298 755656 31354 755712
rect 33138 754024 33194 754080
rect 34518 755384 34574 755440
rect 478786 753480 478842 753536
rect 478142 751440 478198 751496
rect 20626 742464 20682 742520
rect 20442 740832 20498 740888
rect 20166 739472 20222 739528
rect 14186 738928 14242 738984
rect 7746 738656 7802 738712
rect 478050 724920 478106 724976
rect 477958 722200 478014 722256
rect 477038 716896 477094 716952
rect 477314 713360 477370 713416
rect 477130 712136 477186 712192
rect 477130 671268 477186 671324
rect 477406 709144 477462 709200
rect 477314 695748 477370 695804
rect 477958 696904 478014 696960
rect 478050 694184 478106 694240
rect 477406 692280 477462 692336
rect 478694 748720 478750 748776
rect 478602 747360 478658 747416
rect 478326 739880 478382 739936
rect 478234 724240 478290 724296
rect 478234 691328 478290 691384
rect 478142 680176 478198 680232
rect 478510 739200 478566 739256
rect 478418 726960 478474 727016
rect 478418 684392 478474 684448
rect 478510 681808 478566 681864
rect 478326 679768 478382 679824
rect 478694 678952 478750 679008
rect 478602 678408 478658 678464
rect 486146 752800 486202 752856
rect 480902 752120 480958 752176
rect 479522 749400 479578 749456
rect 479430 738520 479486 738576
rect 479338 717440 479394 717496
rect 479430 716896 479486 716952
rect 479430 698264 479486 698320
rect 479338 695544 479394 695600
rect 478786 677592 478842 677648
rect 479798 741920 479854 741976
rect 479614 741240 479670 741296
rect 479706 726280 479762 726336
rect 479706 692960 479762 693016
rect 480166 740560 480222 740616
rect 479982 729680 480038 729736
rect 479890 718120 479946 718176
rect 479798 685888 479854 685944
rect 480074 720160 480130 720216
rect 479982 686160 480038 686216
rect 479890 685072 479946 685128
rect 479614 684936 479670 684992
rect 479522 684256 479578 684312
rect 479430 677456 479486 677512
rect 480810 727640 480866 727696
rect 480810 689968 480866 690024
rect 483754 750760 483810 750816
rect 482282 750080 482338 750136
rect 480994 743280 481050 743336
rect 480902 688336 480958 688392
rect 480166 685752 480222 685808
rect 480166 685208 480222 685264
rect 480074 680312 480130 680368
rect 479982 676912 480038 676968
rect 480258 685092 480314 685128
rect 480258 685072 480260 685092
rect 480260 685072 480312 685092
rect 480312 685072 480314 685092
rect 481178 742600 481234 742656
rect 481086 728320 481142 728376
rect 480994 682080 481050 682136
rect 481454 735800 481510 735856
rect 481362 732400 481418 732456
rect 481270 729000 481326 729056
rect 481178 687792 481234 687848
rect 481362 692688 481418 692744
rect 481270 682352 481326 682408
rect 481086 681536 481142 681592
rect 480166 675824 480222 675880
rect 481546 734440 481602 734496
rect 482098 721520 482154 721576
rect 482190 716760 482246 716816
rect 482098 712136 482154 712192
rect 482098 712000 482154 712056
rect 482006 695000 482062 695056
rect 481914 689696 481970 689752
rect 482190 709144 482246 709200
rect 482190 703704 482246 703760
rect 482098 689152 482154 689208
rect 482006 678272 482062 678328
rect 483662 746680 483718 746736
rect 482374 745320 482430 745376
rect 482834 744640 482890 744696
rect 482650 731040 482706 731096
rect 482466 730360 482522 730416
rect 482374 695952 482430 696008
rect 482558 723560 482614 723616
rect 482466 694592 482522 694648
rect 482742 718800 482798 718856
rect 482650 695408 482706 695464
rect 482558 692824 482614 692880
rect 482282 692416 482338 692472
rect 482282 689832 482338 689888
rect 482190 678136 482246 678192
rect 481546 676096 481602 676152
rect 482926 743960 482982 744016
rect 483478 701800 483534 701856
rect 482834 694320 482890 694376
rect 482926 694184 482982 694240
rect 482926 692688 482982 692744
rect 482834 685752 482890 685808
rect 483570 699760 483626 699816
rect 483570 689968 483626 690024
rect 483478 684392 483534 684448
rect 482926 680312 482982 680368
rect 482742 678952 482798 679008
rect 482282 675960 482338 676016
rect 481454 675008 481510 675064
rect 486146 748040 486202 748096
rect 483938 746000 483994 746056
rect 483846 731720 483902 731776
rect 483846 696904 483902 696960
rect 483754 691192 483810 691248
rect 486146 737840 486202 737896
rect 484306 736480 484362 736536
rect 484214 733760 484270 733816
rect 484122 733080 484178 733136
rect 484030 714040 484086 714096
rect 483938 690376 483994 690432
rect 484122 694048 484178 694104
rect 484030 676232 484086 676288
rect 484214 676096 484270 676152
rect 486146 703840 486202 703896
rect 486146 692688 486202 692744
rect 486330 689832 486386 689888
rect 486238 685208 486294 685264
rect 486422 685072 486478 685128
rect 484306 674736 484362 674792
rect 483662 671880 483718 671936
rect 477222 670724 477278 670780
rect 481546 630400 481602 630456
rect 481454 628360 481510 628416
rect 478786 624960 478842 625016
rect 478694 624280 478750 624336
rect 478694 601704 478750 601760
rect 481454 604424 481510 604480
rect 482926 629720 482982 629776
rect 482834 627680 482890 627736
rect 482282 620200 482338 620256
rect 482834 607144 482890 607200
rect 482282 607008 482338 607064
rect 481546 603064 481602 603120
rect 484306 629040 484362 629096
rect 484214 627000 484270 627056
rect 483662 616800 483718 616856
rect 484214 607144 484270 607200
rect 484306 607008 484362 607064
rect 483662 602792 483718 602848
rect 482926 601704 482982 601760
rect 478786 599120 478842 599176
rect 481546 587832 481602 587888
rect 480166 587152 480222 587208
rect 477130 584704 477186 584760
rect 480074 581576 480130 581632
rect 477130 569880 477186 569936
rect 480074 567160 480130 567216
rect 481454 580896 481510 580952
rect 481362 578992 481418 579048
rect 480166 566480 480222 566536
rect 481362 561720 481418 561776
rect 483662 584568 483718 584624
rect 482926 582392 482982 582448
rect 482834 579536 482890 579592
rect 482834 561040 482890 561096
rect 484306 581576 484362 581632
rect 483662 570560 483718 570616
rect 482926 559680 482982 559736
rect 481546 558320 481602 558376
rect 484306 557640 484362 557696
rect 481454 556960 481510 557016
rect 481546 539960 481602 540016
rect 481454 538600 481510 538656
rect 478786 534520 478842 534576
rect 478694 533160 478750 533216
rect 478602 517248 478658 517304
rect 478602 516840 478658 516896
rect 478694 513304 478750 513360
rect 481454 514800 481510 514856
rect 482926 539280 482982 539336
rect 482834 537240 482890 537296
rect 482834 516160 482890 516216
rect 484306 537920 484362 537976
rect 484214 535880 484270 535936
rect 483662 530440 483718 530496
rect 483662 516432 483718 516488
rect 484214 516296 484270 516352
rect 484306 514936 484362 514992
rect 482926 513712 482982 513768
rect 481546 513304 481602 513360
rect 478786 511808 478842 511864
rect 481546 496848 481602 496904
rect 480166 494264 480222 494320
rect 478786 492632 478842 492688
rect 480074 491136 480130 491192
rect 480074 477400 480130 477456
rect 481454 488552 481510 488608
rect 480166 476720 480222 476776
rect 478786 468560 478842 468616
rect 486422 496168 486478 496224
rect 482926 494672 482982 494728
rect 484306 494672 484362 494728
rect 482282 493584 482338 493640
rect 482834 492632 482890 492688
rect 482282 481480 482338 481536
rect 482834 470600 482890 470656
rect 481546 469240 481602 469296
rect 484214 493992 484270 494048
rect 484214 469920 484270 469976
rect 482926 467880 482982 467936
rect 486146 478080 486202 478136
rect 484306 467200 484362 467256
rect 481454 466520 481510 466576
rect 482926 459720 482982 459776
rect 479522 459040 479578 459096
rect 478786 454960 478842 455016
rect 478694 454280 478750 454336
rect 478510 450880 478566 450936
rect 478418 449520 478474 449576
rect 478418 427216 478474 427272
rect 477406 424768 477462 424824
rect 477406 424374 477462 424430
rect 477406 423408 477462 423464
rect 477406 423014 477462 423070
rect 478602 450200 478658 450256
rect 478510 420960 478566 421016
rect 478602 418240 478658 418296
rect 478694 416608 478750 416664
rect 482834 457680 482890 457736
rect 482742 456320 482798 456376
rect 480902 453600 480958 453656
rect 480166 446120 480222 446176
rect 479982 445440 480038 445496
rect 479890 444080 479946 444136
rect 479890 427216 479946 427272
rect 480074 444760 480130 444816
rect 479982 424496 480038 424552
rect 479522 418104 479578 418160
rect 481546 452240 481602 452296
rect 481454 451560 481510 451616
rect 480902 424088 480958 424144
rect 482650 448840 482706 448896
rect 482006 429392 482062 429448
rect 482006 426128 482062 426184
rect 482650 426128 482706 426184
rect 481546 423544 481602 423600
rect 481454 421368 481510 421424
rect 481454 420008 481510 420064
rect 481454 419736 481510 419792
rect 482742 419736 482798 419792
rect 482834 419600 482890 419656
rect 480166 419464 480222 419520
rect 480074 417288 480130 417344
rect 484306 458360 484362 458416
rect 484214 457000 484270 457056
rect 484122 455640 484178 455696
rect 484030 448160 484086 448216
rect 483110 424904 483166 424960
rect 484030 424904 484086 424960
rect 483110 424496 483166 424552
rect 484122 423544 484178 423600
rect 482926 416608 482982 416664
rect 484214 416608 484270 416664
rect 486146 446800 486202 446856
rect 486146 437960 486202 438016
rect 486054 424496 486110 424552
rect 486238 429392 486294 429448
rect 478786 415248 478842 415304
rect 484306 415248 484362 415304
rect 478786 399472 478842 399528
rect 478694 398792 478750 398848
rect 478694 387640 478750 387696
rect 479522 398792 479578 398848
rect 478786 386960 478842 387016
rect 479522 386280 479578 386336
rect 481546 360440 481602 360496
rect 481454 358400 481510 358456
rect 478786 355000 478842 355056
rect 478694 353640 478750 353696
rect 477130 349560 477186 349616
rect 477130 335756 477186 335812
rect 478694 334056 478750 334112
rect 481454 336640 481510 336696
rect 484306 359760 484362 359816
rect 482926 359080 482982 359136
rect 482282 346840 482338 346896
rect 481546 334056 481602 334112
rect 484214 357720 484270 357776
rect 482926 336640 482982 336696
rect 484214 336640 484270 336696
rect 484306 334056 484362 334112
rect 482282 332696 482338 332752
rect 478786 329568 478842 329624
rect 481546 318688 481602 318744
rect 480166 314880 480222 314936
rect 480074 311208 480130 311264
rect 479982 310392 480038 310448
rect 479982 297880 480038 297936
rect 480074 297200 480130 297256
rect 481454 310392 481510 310448
rect 480166 296520 480222 296576
rect 486054 314744 486110 314800
rect 482282 314472 482338 314528
rect 482926 311888 482982 311944
rect 482834 308896 482890 308952
rect 482282 300600 482338 300656
rect 482834 289720 482890 289776
rect 481546 288360 481602 288416
rect 484306 311208 484362 311264
rect 486054 299920 486110 299976
rect 484306 289040 484362 289096
rect 482926 287680 482982 287736
rect 481454 287000 481510 287056
rect 481546 270000 481602 270056
rect 481454 267960 481510 268016
rect 478694 264560 478750 264616
rect 478602 263200 478658 263256
rect 478602 247016 478658 247072
rect 478786 263880 478842 263936
rect 478694 245656 478750 245712
rect 481454 247016 481510 247072
rect 482926 269320 482982 269376
rect 482834 266600 482890 266656
rect 482834 247016 482890 247072
rect 484306 268640 484362 268696
rect 483662 255720 483718 255776
rect 483202 248240 483258 248296
rect 483202 247968 483258 248024
rect 482926 245656 482982 245712
rect 481546 244296 481602 244352
rect 478786 242800 478842 242856
rect 484306 243480 484362 243536
rect 483662 241712 483718 241768
rect 482926 241440 482982 241496
rect 482926 240352 482982 240408
rect 481546 226344 481602 226400
rect 481454 224032 481510 224088
rect 481454 223760 481510 223816
rect 480166 223624 480222 223680
rect 478786 220904 478842 220960
rect 477406 219294 477462 219350
rect 478694 219272 478750 219328
rect 477406 218320 477462 218376
rect 478694 198600 478750 198656
rect 481454 221312 481510 221368
rect 481454 221040 481510 221096
rect 481454 220904 481510 220960
rect 480166 206760 480222 206816
rect 478786 197920 478842 197976
rect 486422 226072 486478 226128
rect 482926 223624 482982 223680
rect 484306 223624 484362 223680
rect 482834 220904 482890 220960
rect 482834 202000 482890 202056
rect 484214 222264 484270 222320
rect 482926 200640 482982 200696
rect 484214 199960 484270 200016
rect 481546 199280 481602 199336
rect 486146 208120 486202 208176
rect 484306 197240 484362 197296
rect 481454 196560 481510 196616
rect 482926 192480 482982 192536
rect 478142 191800 478198 191856
rect 480166 190440 480222 190496
rect 479522 189760 479578 189816
rect 478694 185680 478750 185736
rect 478602 184320 478658 184376
rect 478510 180920 478566 180976
rect 478510 152904 478566 152960
rect 478602 152632 478658 152688
rect 478786 185000 478842 185056
rect 478694 147736 478750 147792
rect 479982 177520 480038 177576
rect 479890 176160 479946 176216
rect 479890 156712 479946 156768
rect 480074 176840 480130 176896
rect 480074 148824 480130 148880
rect 479982 148688 480038 148744
rect 479522 147056 479578 147112
rect 482834 188400 482890 188456
rect 482742 187040 482798 187096
rect 480902 183640 480958 183696
rect 480994 182960 481050 183016
rect 481546 182280 481602 182336
rect 481454 175480 481510 175536
rect 480994 154672 481050 154728
rect 480902 154128 480958 154184
rect 482650 179560 482706 179616
rect 481638 162696 481694 162752
rect 481638 155896 481694 155952
rect 481546 153040 481602 153096
rect 482650 150456 482706 150512
rect 482834 149232 482890 149288
rect 482742 149096 482798 149152
rect 481454 147056 481510 147112
rect 480166 146376 480222 146432
rect 484030 191120 484086 191176
rect 483938 178880 483994 178936
rect 483662 166640 483718 166696
rect 483938 157392 483994 157448
rect 484306 189080 484362 189136
rect 484214 187720 484270 187776
rect 484122 186360 484178 186416
rect 484030 155896 484086 155952
rect 483662 152768 483718 152824
rect 483110 151680 483166 151736
rect 483110 150864 483166 150920
rect 484122 150456 484178 150512
rect 484214 147736 484270 147792
rect 486146 178200 486202 178256
rect 486146 168000 486202 168056
rect 486054 162696 486110 162752
rect 486238 154808 486294 154864
rect 482926 146240 482982 146296
rect 484306 146240 484362 146296
rect 478786 144744 478842 144800
rect 478142 144608 478198 144664
rect 483662 135088 483718 135144
rect 483662 119720 483718 119776
rect 481546 90480 481602 90536
rect 481454 88440 481510 88496
rect 478694 85040 478750 85096
rect 478786 84360 478842 84416
rect 478694 63688 478750 63744
rect 480166 80960 480222 81016
rect 481454 67496 481510 67552
rect 480166 66136 480222 66192
rect 484306 89800 484362 89856
rect 482926 89120 482982 89176
rect 482834 87080 482890 87136
rect 482282 79600 482338 79656
rect 482834 67496 482890 67552
rect 482282 64096 482338 64152
rect 484214 87760 484270 87816
rect 484214 67496 484270 67552
rect 484306 65864 484362 65920
rect 481546 62192 481602 62248
rect 482926 62192 482982 62248
rect 478786 60560 478842 60616
rect 481546 48184 481602 48240
rect 477222 47368 477278 47424
rect 477222 46960 477278 47016
rect 480166 44376 480222 44432
rect 480074 39888 480130 39944
rect 6182 32000 6238 32056
rect 4802 31320 4858 31376
rect 1122 30640 1178 30696
rect 1122 28872 1178 28928
rect 202 28328 258 28384
rect 1306 27920 1362 27976
rect 1214 26560 1270 26616
rect 3422 23840 3478 23896
rect 1306 23704 1362 23760
rect 1214 21936 1270 21992
rect 202 17992 258 18048
rect 4894 29280 4950 29336
rect 5078 28872 5134 28928
rect 5538 23160 5594 23216
rect 5078 17856 5134 17912
rect 4894 16768 4950 16824
rect 7102 31184 7158 31240
rect 6458 23024 6514 23080
rect 5538 16632 5594 16688
rect 4802 16496 4858 16552
rect 3422 16088 3478 16144
rect 9310 30368 9366 30424
rect 7562 29960 7618 30016
rect 7378 23704 7434 23760
rect 8666 28736 8722 28792
rect 8206 27920 8262 27976
rect 7654 27240 7710 27296
rect 8022 27104 8078 27160
rect 7746 23840 7802 23896
rect 8114 16532 8116 16552
rect 8116 16532 8168 16552
rect 8168 16532 8170 16552
rect 8114 16496 8170 16532
rect 8482 17992 8538 18048
rect 8022 992 8078 1048
rect 8390 1264 8446 1320
rect 8114 856 8170 912
rect 8942 25200 8998 25256
rect 8850 21936 8906 21992
rect 9034 24656 9090 24712
rect 8942 16224 8998 16280
rect 8666 1128 8722 1184
rect 9126 20440 9182 20496
rect 9218 17856 9274 17912
rect 9126 17448 9182 17504
rect 9586 29484 9642 29540
rect 9402 26288 9458 26344
rect 9310 4120 9366 4176
rect 9494 19760 9550 19816
rect 9494 16904 9550 16960
rect 9402 1264 9458 1320
rect 480074 27240 480130 27296
rect 480166 26560 480222 26616
rect 486422 44648 486478 44704
rect 483110 44240 483166 44296
rect 482926 41384 482982 41440
rect 482834 39888 482890 39944
rect 482834 21120 482890 21176
rect 484306 43288 484362 43344
rect 483294 43152 483350 43208
rect 483294 42880 483350 42936
rect 484214 41384 484270 41440
rect 483110 30640 483166 30696
rect 482926 19760 482982 19816
rect 484214 19080 484270 19136
rect 481546 18400 481602 18456
rect 486146 29960 486202 30016
rect 484306 17720 484362 17776
rect 12346 16904 12402 16960
rect 11886 16768 11942 16824
rect 13220 17040 13276 17096
rect 13680 17040 13736 17096
rect 14186 16632 14242 16688
rect 17820 17040 17876 17096
rect 18740 17040 18796 17096
rect 17406 16904 17462 16960
rect 16946 16496 17002 16552
rect 16026 16224 16082 16280
rect 15566 16088 15622 16144
rect 12806 15952 12862 16008
rect 18878 13640 18934 13696
rect 18878 12960 18934 13016
rect 11518 12280 11574 12336
rect 11794 12144 11850 12200
rect 20350 9016 20406 9072
rect 10966 8200 11022 8256
rect 14186 8200 14242 8256
rect 21086 8200 21142 8256
rect 20350 7928 20406 7984
rect 20534 7928 20590 7984
rect 14186 5888 14242 5944
rect 11610 5616 11666 5672
rect 10322 1264 10378 1320
rect 10966 1128 11022 1184
rect 12898 4120 12954 4176
rect 12254 992 12310 1048
rect 13542 856 13598 912
rect 21086 7656 21142 7712
rect 20626 7384 20682 7440
rect 20626 3576 20682 3632
rect 22558 3576 22614 3632
rect 29182 5888 29238 5944
rect 72376 5888 72432 5944
rect 104648 5888 104704 5944
rect 177108 5888 177164 5944
rect 218104 5888 218160 5944
rect 259136 5888 259192 5944
rect 276556 5888 276612 5944
rect 345110 5888 345166 5944
rect 378920 5888 378976 5944
rect 380070 312 380126 368
rect 383348 5752 383404 5808
rect 385590 1264 385646 1320
rect 386418 1264 386474 1320
rect 384486 1128 384542 1184
rect 387706 1128 387762 1184
rect 386694 992 386750 1048
rect 382278 448 382334 504
rect 381174 176 381230 232
rect 386970 176 387026 232
rect 388258 448 388314 504
rect 388902 1264 388958 1320
rect 389638 1264 389694 1320
rect 390926 992 390982 1048
rect 392858 5752 392914 5808
rect 394054 312 394110 368
rect 414412 5888 414468 5944
rect 444464 5888 444520 5944
<< metal3 >>
rect 21214 755788 21220 755852
rect 21284 755850 21290 755852
rect 26785 755850 26851 755853
rect 21284 755848 26851 755850
rect 21284 755792 26790 755848
rect 26846 755792 26851 755848
rect 21284 755790 26851 755792
rect 21284 755788 21290 755790
rect 26785 755787 26851 755790
rect 20437 755714 20503 755717
rect 31293 755714 31359 755717
rect 20437 755712 31359 755714
rect 20437 755656 20442 755712
rect 20498 755656 31298 755712
rect 31354 755656 31359 755712
rect 20437 755654 31359 755656
rect 20437 755651 20503 755654
rect 31293 755651 31359 755654
rect 20069 755442 20135 755445
rect 34513 755442 34579 755445
rect 20069 755440 34579 755442
rect 20069 755384 20074 755440
rect 20130 755384 34518 755440
rect 34574 755384 34579 755440
rect 20069 755382 34579 755384
rect 20069 755379 20135 755382
rect 34513 755379 34579 755382
rect 19926 754972 19932 755036
rect 19996 755034 20002 755036
rect 27981 755034 28047 755037
rect 19996 755032 28047 755034
rect 19996 754976 27986 755032
rect 28042 754976 28047 755032
rect 19996 754974 28047 754976
rect 19996 754972 20002 754974
rect 27981 754971 28047 754974
rect 20253 754898 20319 754901
rect 23565 754898 23631 754901
rect 20253 754896 23631 754898
rect 20253 754840 20258 754896
rect 20314 754840 23570 754896
rect 23626 754840 23631 754896
rect 20253 754838 23631 754840
rect 20253 754835 20319 754838
rect 23565 754835 23631 754838
rect 20345 754082 20411 754085
rect 33133 754082 33199 754085
rect 20345 754080 33199 754082
rect 20345 754024 20350 754080
rect 20406 754024 33138 754080
rect 33194 754024 33199 754080
rect 20345 754022 33199 754024
rect 20345 754019 20411 754022
rect 33133 754019 33199 754022
rect 21449 753538 21515 753541
rect 22277 753538 22343 753541
rect 21449 753536 22343 753538
rect 21449 753480 21454 753536
rect 21510 753480 22282 753536
rect 22338 753480 22343 753536
rect 21449 753478 22343 753480
rect 21449 753475 21515 753478
rect 22277 753475 22343 753478
rect 478781 753538 478847 753541
rect 486200 753538 487000 753568
rect 478781 753536 487000 753538
rect 478781 753480 478786 753536
rect 478842 753480 487000 753536
rect 478781 753478 487000 753480
rect 478781 753475 478847 753478
rect 486200 753448 487000 753478
rect 486200 752861 487000 752888
rect 486141 752856 487000 752861
rect 486141 752800 486146 752856
rect 486202 752800 487000 752856
rect 486141 752795 487000 752800
rect 486200 752768 487000 752795
rect 20437 752722 20503 752725
rect 30005 752722 30071 752725
rect 20437 752720 30071 752722
rect 20437 752664 20442 752720
rect 20498 752664 30010 752720
rect 30066 752664 30071 752720
rect 20437 752662 30071 752664
rect 20437 752659 20503 752662
rect 30005 752659 30071 752662
rect 480897 752178 480963 752181
rect 486200 752178 487000 752208
rect 480897 752176 487000 752178
rect 480897 752120 480902 752176
rect 480958 752120 487000 752176
rect 480897 752118 487000 752120
rect 480897 752115 480963 752118
rect 486200 752088 487000 752118
rect 478137 751498 478203 751501
rect 486200 751498 487000 751528
rect 478137 751496 487000 751498
rect 478137 751440 478142 751496
rect 478198 751440 487000 751496
rect 478137 751438 487000 751440
rect 478137 751435 478203 751438
rect 486200 751408 487000 751438
rect 483749 750818 483815 750821
rect 486200 750818 487000 750848
rect 483749 750816 487000 750818
rect 483749 750760 483754 750816
rect 483810 750760 487000 750816
rect 483749 750758 487000 750760
rect 483749 750755 483815 750758
rect 486200 750728 487000 750758
rect 482277 750138 482343 750141
rect 486200 750138 487000 750168
rect 482277 750136 487000 750138
rect 482277 750080 482282 750136
rect 482338 750080 487000 750136
rect 482277 750078 487000 750080
rect 482277 750075 482343 750078
rect 486200 750048 487000 750078
rect 20161 749594 20227 749597
rect 22001 749594 22067 749597
rect 20161 749592 22067 749594
rect 20161 749536 20166 749592
rect 20222 749536 22006 749592
rect 22062 749536 22067 749592
rect 20161 749534 22067 749536
rect 20161 749531 20227 749534
rect 22001 749531 22067 749534
rect 20662 749396 20668 749460
rect 20732 749458 20738 749460
rect 21173 749458 21239 749461
rect 20732 749456 21239 749458
rect 20732 749400 21178 749456
rect 21234 749400 21239 749456
rect 20732 749398 21239 749400
rect 20732 749396 20738 749398
rect 21173 749395 21239 749398
rect 479517 749458 479583 749461
rect 486200 749458 487000 749488
rect 479517 749456 487000 749458
rect 479517 749400 479522 749456
rect 479578 749400 487000 749456
rect 479517 749398 487000 749400
rect 479517 749395 479583 749398
rect 486200 749368 487000 749398
rect 478689 748778 478755 748781
rect 486200 748778 487000 748808
rect 478689 748776 487000 748778
rect 478689 748720 478694 748776
rect 478750 748720 487000 748776
rect 478689 748718 487000 748720
rect 478689 748715 478755 748718
rect 486200 748688 487000 748718
rect 20478 748580 20484 748644
rect 20548 748642 20554 748644
rect 25865 748642 25931 748645
rect 20548 748640 25931 748642
rect 20548 748584 25870 748640
rect 25926 748584 25931 748640
rect 20548 748582 25931 748584
rect 20548 748580 20554 748582
rect 25865 748579 25931 748582
rect 486200 748101 487000 748128
rect 486141 748096 487000 748101
rect 486141 748040 486146 748096
rect 486202 748040 487000 748096
rect 486141 748035 487000 748040
rect 486200 748008 487000 748035
rect 478597 747418 478663 747421
rect 486200 747418 487000 747448
rect 478597 747416 487000 747418
rect 478597 747360 478602 747416
rect 478658 747360 487000 747416
rect 478597 747358 487000 747360
rect 478597 747355 478663 747358
rect 486200 747328 487000 747358
rect 9121 747146 9187 747149
rect 9121 747144 21282 747146
rect 9121 747088 9126 747144
rect 9182 747088 21282 747144
rect 9121 747086 21282 747088
rect 9121 747083 9187 747086
rect 21272 746834 21278 746898
rect 21342 746834 21348 746898
rect 483657 746738 483723 746741
rect 486200 746738 487000 746768
rect 483657 746736 487000 746738
rect 483657 746680 483662 746736
rect 483718 746680 487000 746736
rect 483657 746678 487000 746680
rect 483657 746675 483723 746678
rect 486200 746648 487000 746678
rect 12985 746602 13051 746605
rect 12985 746600 21282 746602
rect 12985 746544 12990 746600
rect 13046 746544 21282 746600
rect 12985 746542 21282 746544
rect 12985 746539 13051 746542
rect 9765 746330 9831 746333
rect 9765 746328 21282 746330
rect 9765 746272 9770 746328
rect 9826 746272 21282 746328
rect 9765 746270 21282 746272
rect 9765 746267 9831 746270
rect 18137 746058 18203 746061
rect 483933 746058 483999 746061
rect 486200 746058 487000 746088
rect 18137 746056 21282 746058
rect 18137 746000 18142 746056
rect 18198 746000 21282 746056
rect 18137 745998 21282 746000
rect 483933 746056 487000 746058
rect 483933 746000 483938 746056
rect 483994 746000 487000 746056
rect 483933 745998 487000 746000
rect 18137 745995 18203 745998
rect 483933 745995 483999 745998
rect 486200 745968 487000 745998
rect 20529 745786 20595 745789
rect 20529 745784 21282 745786
rect 20529 745728 20534 745784
rect 20590 745728 21282 745784
rect 20529 745726 21282 745728
rect 20529 745723 20595 745726
rect 8293 745514 8359 745517
rect 8293 745512 21282 745514
rect 8293 745456 8298 745512
rect 8354 745456 21282 745512
rect 8293 745454 21282 745456
rect 8293 745451 8359 745454
rect 482369 745378 482435 745381
rect 486200 745378 487000 745408
rect 482369 745376 487000 745378
rect 482369 745320 482374 745376
rect 482430 745320 487000 745376
rect 482369 745318 487000 745320
rect 482369 745315 482435 745318
rect 486200 745288 487000 745318
rect 18597 745242 18663 745245
rect 18597 745240 21282 745242
rect 18597 745184 18602 745240
rect 18658 745184 21282 745240
rect 18597 745182 21282 745184
rect 18597 745179 18663 745182
rect 13445 744970 13511 744973
rect 13445 744968 21282 744970
rect 13445 744912 13450 744968
rect 13506 744912 21282 744968
rect 13445 744910 21282 744912
rect 13445 744907 13511 744910
rect 20253 744698 20319 744701
rect 482829 744698 482895 744701
rect 486200 744698 487000 744728
rect 20253 744696 21282 744698
rect 20253 744640 20258 744696
rect 20314 744640 21282 744696
rect 20253 744638 21282 744640
rect 482829 744696 487000 744698
rect 482829 744640 482834 744696
rect 482890 744640 487000 744696
rect 482829 744638 487000 744640
rect 20253 744635 20319 744638
rect 482829 744635 482895 744638
rect 486200 744608 487000 744638
rect 21081 744448 21147 744451
rect 21081 744446 21282 744448
rect 21081 744390 21086 744446
rect 21142 744390 21282 744446
rect 21081 744388 21282 744390
rect 21081 744385 21147 744388
rect 19425 744154 19491 744157
rect 19425 744152 21282 744154
rect 19425 744096 19430 744152
rect 19486 744096 21282 744152
rect 19425 744094 21282 744096
rect 19425 744091 19491 744094
rect 482921 744018 482987 744021
rect 486200 744018 487000 744048
rect 482921 744016 487000 744018
rect 482921 743960 482926 744016
rect 482982 743960 487000 744016
rect 482921 743958 487000 743960
rect 482921 743955 482987 743958
rect 486200 743928 487000 743958
rect 11697 743882 11763 743885
rect 11697 743880 21282 743882
rect 11697 743824 11702 743880
rect 11758 743824 21282 743880
rect 11697 743822 21282 743824
rect 11697 743819 11763 743822
rect 17309 743610 17375 743613
rect 17309 743608 21282 743610
rect 17309 743552 17314 743608
rect 17370 743552 21282 743608
rect 17309 743550 21282 743552
rect 17309 743547 17375 743550
rect 19926 743276 19932 743340
rect 19996 743338 20002 743340
rect 480989 743338 481055 743341
rect 486200 743338 487000 743368
rect 19996 743278 21282 743338
rect 480989 743336 487000 743338
rect 480989 743280 480994 743336
rect 481050 743280 487000 743336
rect 480989 743278 487000 743280
rect 19996 743276 20002 743278
rect 480989 743275 481055 743278
rect 486200 743248 487000 743278
rect 10409 743066 10475 743069
rect 10409 743064 21282 743066
rect 10409 743008 10414 743064
rect 10470 743008 21282 743064
rect 10409 743006 21282 743008
rect 10409 743003 10475 743006
rect 14733 742794 14799 742797
rect 14733 742792 21282 742794
rect 14733 742736 14738 742792
rect 14794 742736 21282 742792
rect 14733 742734 21282 742736
rect 14733 742731 14799 742734
rect 481173 742658 481239 742661
rect 486200 742658 487000 742688
rect 481173 742656 487000 742658
rect 481173 742600 481178 742656
rect 481234 742600 487000 742656
rect 481173 742598 487000 742600
rect 481173 742595 481239 742598
rect 486200 742568 487000 742598
rect 20621 742522 20687 742525
rect 20621 742520 21282 742522
rect 20621 742464 20626 742520
rect 20682 742464 21282 742520
rect 20621 742462 21282 742464
rect 20621 742459 20687 742462
rect 19885 742250 19951 742253
rect 19885 742248 21282 742250
rect 19885 742192 19890 742248
rect 19946 742192 21282 742248
rect 19885 742190 21282 742192
rect 19885 742187 19951 742190
rect 12157 741978 12223 741981
rect 479793 741978 479859 741981
rect 486200 741978 487000 742008
rect 12157 741976 21282 741978
rect 12157 741920 12162 741976
rect 12218 741920 21282 741976
rect 12157 741918 21282 741920
rect 479793 741976 487000 741978
rect 479793 741920 479798 741976
rect 479854 741920 487000 741976
rect 479793 741918 487000 741920
rect 12157 741915 12223 741918
rect 479793 741915 479859 741918
rect 486200 741888 487000 741918
rect 15561 741706 15627 741709
rect 15561 741704 21282 741706
rect 15561 741648 15566 741704
rect 15622 741648 21282 741704
rect 15561 741646 21282 741648
rect 15561 741643 15627 741646
rect 20662 741394 20668 741458
rect 20732 741456 20738 741458
rect 20732 741396 21282 741456
rect 20732 741394 20738 741396
rect 479609 741298 479675 741301
rect 486200 741298 487000 741328
rect 479609 741296 487000 741298
rect 479609 741240 479614 741296
rect 479670 741240 487000 741296
rect 479609 741238 487000 741240
rect 479609 741235 479675 741238
rect 486200 741208 487000 741238
rect 20345 741162 20411 741165
rect 20345 741160 21282 741162
rect 20345 741104 20350 741160
rect 20406 741104 21282 741160
rect 20345 741102 21282 741104
rect 20345 741099 20411 741102
rect 20437 740890 20503 740893
rect 20437 740888 21282 740890
rect 20437 740832 20442 740888
rect 20498 740832 21282 740888
rect 20437 740830 21282 740832
rect 20437 740827 20503 740830
rect 16113 740618 16179 740621
rect 480161 740618 480227 740621
rect 486200 740618 487000 740648
rect 16113 740616 21282 740618
rect 16113 740560 16118 740616
rect 16174 740560 21282 740616
rect 16113 740558 21282 740560
rect 480161 740616 487000 740618
rect 480161 740560 480166 740616
rect 480222 740560 487000 740616
rect 480161 740558 487000 740560
rect 16113 740555 16179 740558
rect 480161 740555 480227 740558
rect 486200 740528 487000 740558
rect 20069 740346 20135 740349
rect 20069 740344 21282 740346
rect 20069 740288 20074 740344
rect 20130 740288 21282 740344
rect 20069 740286 21282 740288
rect 20069 740283 20135 740286
rect 20478 740012 20484 740076
rect 20548 740074 20554 740076
rect 20548 740014 21282 740074
rect 20548 740012 20554 740014
rect 478321 739938 478387 739941
rect 486200 739938 487000 739968
rect 478321 739936 487000 739938
rect 478321 739880 478326 739936
rect 478382 739880 487000 739936
rect 478321 739878 487000 739880
rect 478321 739875 478387 739878
rect 486200 739848 487000 739878
rect 16757 739802 16823 739805
rect 16757 739800 21282 739802
rect 16757 739744 16762 739800
rect 16818 739744 21282 739800
rect 16757 739742 21282 739744
rect 16757 739739 16823 739742
rect 20161 739530 20227 739533
rect 20161 739528 21282 739530
rect 20161 739472 20166 739528
rect 20222 739472 21282 739528
rect 20161 739470 21282 739472
rect 20161 739467 20227 739470
rect 10961 739258 11027 739261
rect 478505 739258 478571 739261
rect 486200 739258 487000 739288
rect 10961 739256 21282 739258
rect 10961 739200 10966 739256
rect 11022 739200 21282 739256
rect 10961 739198 21282 739200
rect 478505 739256 487000 739258
rect 478505 739200 478510 739256
rect 478566 739200 487000 739256
rect 478505 739198 487000 739200
rect 10961 739195 11027 739198
rect 478505 739195 478571 739198
rect 486200 739168 487000 739198
rect 14181 738986 14247 738989
rect 14181 738984 21282 738986
rect 14181 738928 14186 738984
rect 14242 738928 21282 738984
rect 14181 738926 21282 738928
rect 14181 738923 14247 738926
rect 7741 738714 7807 738717
rect 7741 738712 21282 738714
rect 7741 738656 7746 738712
rect 7802 738656 21282 738712
rect 7741 738654 21282 738656
rect 7741 738651 7807 738654
rect 479425 738578 479491 738581
rect 486200 738578 487000 738608
rect 479425 738576 487000 738578
rect 479425 738520 479430 738576
rect 479486 738520 487000 738576
rect 479425 738518 487000 738520
rect 479425 738515 479491 738518
rect 486200 738488 487000 738518
rect 486200 737901 487000 737928
rect 486141 737896 487000 737901
rect 486141 737840 486146 737896
rect 486202 737840 487000 737896
rect 486141 737835 487000 737840
rect 486200 737808 487000 737835
rect 480110 737156 480116 737220
rect 480180 737218 480186 737220
rect 486200 737218 487000 737248
rect 480180 737158 487000 737218
rect 480180 737156 480186 737158
rect 486200 737128 487000 737158
rect 484301 736538 484367 736541
rect 486200 736538 487000 736568
rect 484301 736536 487000 736538
rect 484301 736480 484306 736536
rect 484362 736480 487000 736536
rect 484301 736478 487000 736480
rect 484301 736475 484367 736478
rect 486200 736448 487000 736478
rect 481449 735858 481515 735861
rect 486200 735858 487000 735888
rect 481449 735856 487000 735858
rect 481449 735800 481454 735856
rect 481510 735800 487000 735856
rect 481449 735798 487000 735800
rect 481449 735795 481515 735798
rect 486200 735768 487000 735798
rect 482870 735116 482876 735180
rect 482940 735178 482946 735180
rect 486200 735178 487000 735208
rect 482940 735118 487000 735178
rect 482940 735116 482946 735118
rect 486200 735088 487000 735118
rect 481541 734498 481607 734501
rect 486200 734498 487000 734528
rect 481541 734496 487000 734498
rect 481541 734440 481546 734496
rect 481602 734440 487000 734496
rect 481541 734438 487000 734440
rect 481541 734435 481607 734438
rect 486200 734408 487000 734438
rect 484209 733818 484275 733821
rect 486200 733818 487000 733848
rect 484209 733816 487000 733818
rect 484209 733760 484214 733816
rect 484270 733760 487000 733816
rect 484209 733758 487000 733760
rect 484209 733755 484275 733758
rect 486200 733728 487000 733758
rect 0 733138 800 733168
rect 484117 733138 484183 733141
rect 486200 733138 487000 733168
rect 0 733078 10032 733138
rect 484117 733136 487000 733138
rect 484117 733080 484122 733136
rect 484178 733080 487000 733136
rect 484117 733078 487000 733080
rect 0 733048 800 733078
rect 484117 733075 484183 733078
rect 486200 733048 487000 733078
rect 0 732458 800 732488
rect 481357 732458 481423 732461
rect 486200 732458 487000 732488
rect 0 732398 9506 732458
rect 0 732368 800 732398
rect 9446 732360 9506 732398
rect 481357 732456 487000 732458
rect 481357 732400 481362 732456
rect 481418 732400 487000 732456
rect 481357 732398 487000 732400
rect 481357 732395 481423 732398
rect 486200 732368 487000 732398
rect 9446 732300 10060 732360
rect 0 731778 800 731808
rect 483841 731778 483907 731781
rect 486200 731778 487000 731808
rect 0 731718 9506 731778
rect 0 731688 800 731718
rect 9446 731544 9506 731718
rect 483841 731776 487000 731778
rect 483841 731720 483846 731776
rect 483902 731720 487000 731776
rect 483841 731718 487000 731720
rect 483841 731715 483907 731718
rect 486200 731688 487000 731718
rect 9446 731484 10060 731544
rect 482645 731098 482711 731101
rect 486200 731098 487000 731128
rect 482645 731096 487000 731098
rect 482645 731040 482650 731096
rect 482706 731040 487000 731096
rect 482645 731038 487000 731040
rect 482645 731035 482711 731038
rect 486200 731008 487000 731038
rect 9446 730612 10060 730672
rect 0 730418 800 730448
rect 9446 730418 9506 730612
rect 0 730358 9506 730418
rect 482461 730418 482527 730421
rect 486200 730418 487000 730448
rect 482461 730416 487000 730418
rect 482461 730360 482466 730416
rect 482522 730360 487000 730416
rect 482461 730358 487000 730360
rect 0 730328 800 730358
rect 482461 730355 482527 730358
rect 486200 730328 487000 730358
rect 9446 729796 10060 729856
rect 0 729738 800 729768
rect 9446 729738 9506 729796
rect 0 729678 9506 729738
rect 479977 729738 480043 729741
rect 486200 729738 487000 729768
rect 479977 729736 487000 729738
rect 479977 729680 479982 729736
rect 480038 729680 487000 729736
rect 479977 729678 487000 729680
rect 0 729648 800 729678
rect 479977 729675 480043 729678
rect 486200 729648 487000 729678
rect 0 729058 800 729088
rect 481265 729058 481331 729061
rect 486200 729058 487000 729088
rect 0 728998 10032 729058
rect 481265 729056 487000 729058
rect 481265 729000 481270 729056
rect 481326 729000 487000 729056
rect 481265 728998 487000 729000
rect 0 728968 800 728998
rect 481265 728995 481331 728998
rect 486200 728968 487000 728998
rect 0 728378 800 728408
rect 481081 728378 481147 728381
rect 486200 728378 487000 728408
rect 0 728318 9506 728378
rect 0 728288 800 728318
rect 9446 728280 9506 728318
rect 481081 728376 487000 728378
rect 481081 728320 481086 728376
rect 481142 728320 487000 728376
rect 481081 728318 487000 728320
rect 481081 728315 481147 728318
rect 486200 728288 487000 728318
rect 9446 728220 10060 728280
rect 0 727698 800 727728
rect 480805 727698 480871 727701
rect 486200 727698 487000 727728
rect 0 727638 9506 727698
rect 0 727608 800 727638
rect 9446 727464 9506 727638
rect 480805 727696 487000 727698
rect 480805 727640 480810 727696
rect 480866 727640 487000 727696
rect 480805 727638 487000 727640
rect 480805 727635 480871 727638
rect 486200 727608 487000 727638
rect 9446 727404 10060 727464
rect 478413 727018 478479 727021
rect 486200 727018 487000 727048
rect 478413 727016 487000 727018
rect 478413 726960 478418 727016
rect 478474 726960 487000 727016
rect 478413 726958 487000 726960
rect 478413 726955 478479 726958
rect 486200 726928 487000 726958
rect 9446 726532 10060 726592
rect 0 726338 800 726368
rect 9446 726338 9506 726532
rect 0 726278 9506 726338
rect 479701 726338 479767 726341
rect 486200 726338 487000 726368
rect 479701 726336 487000 726338
rect 479701 726280 479706 726336
rect 479762 726280 487000 726336
rect 479701 726278 487000 726280
rect 0 726248 800 726278
rect 479701 726275 479767 726278
rect 486200 726248 487000 726278
rect 9446 725716 10060 725776
rect 0 725658 800 725688
rect 9446 725658 9506 725716
rect 0 725598 9506 725658
rect 0 725568 800 725598
rect 483606 725596 483612 725660
rect 483676 725658 483682 725660
rect 486200 725658 487000 725688
rect 483676 725598 487000 725658
rect 483676 725596 483682 725598
rect 486200 725568 487000 725598
rect 0 724978 800 725008
rect 478045 724978 478111 724981
rect 486200 724978 487000 725008
rect 0 724918 10032 724978
rect 478045 724976 487000 724978
rect 478045 724920 478050 724976
rect 478106 724920 487000 724976
rect 478045 724918 487000 724920
rect 0 724888 800 724918
rect 478045 724915 478111 724918
rect 486200 724888 487000 724918
rect 0 724298 800 724328
rect 478229 724298 478295 724301
rect 486200 724298 487000 724328
rect 0 724238 9506 724298
rect 0 724208 800 724238
rect 9446 724200 9506 724238
rect 478229 724296 487000 724298
rect 478229 724240 478234 724296
rect 478290 724240 487000 724296
rect 478229 724238 487000 724240
rect 478229 724235 478295 724238
rect 486200 724208 487000 724238
rect 9446 724140 10060 724200
rect 0 723618 800 723648
rect 482553 723618 482619 723621
rect 486200 723618 487000 723648
rect 0 723558 9506 723618
rect 0 723528 800 723558
rect 9446 723384 9506 723558
rect 482553 723616 487000 723618
rect 482553 723560 482558 723616
rect 482614 723560 487000 723616
rect 482553 723558 487000 723560
rect 482553 723555 482619 723558
rect 486200 723528 487000 723558
rect 9446 723324 10060 723384
rect 483974 722876 483980 722940
rect 484044 722938 484050 722940
rect 486200 722938 487000 722968
rect 484044 722878 487000 722938
rect 484044 722876 484050 722878
rect 486200 722848 487000 722878
rect 9446 722452 10060 722512
rect 0 722258 800 722288
rect 9446 722258 9506 722452
rect 0 722198 9506 722258
rect 477953 722258 478019 722261
rect 486200 722258 487000 722288
rect 477953 722256 487000 722258
rect 477953 722200 477958 722256
rect 478014 722200 487000 722256
rect 477953 722198 487000 722200
rect 0 722168 800 722198
rect 477953 722195 478019 722198
rect 486200 722168 487000 722198
rect 9446 721636 10060 721696
rect 0 721578 800 721608
rect 9446 721578 9506 721636
rect 0 721518 9506 721578
rect 482093 721578 482159 721581
rect 486200 721578 487000 721608
rect 482093 721576 487000 721578
rect 482093 721520 482098 721576
rect 482154 721520 487000 721576
rect 482093 721518 487000 721520
rect 0 721488 800 721518
rect 482093 721515 482159 721518
rect 486200 721488 487000 721518
rect 0 720898 800 720928
rect 0 720838 10032 720898
rect 0 720808 800 720838
rect 484894 720836 484900 720900
rect 484964 720898 484970 720900
rect 486200 720898 487000 720928
rect 484964 720838 487000 720898
rect 484964 720836 484970 720838
rect 486200 720808 487000 720838
rect 0 720218 800 720248
rect 480069 720218 480135 720221
rect 486200 720218 487000 720248
rect 0 720158 9506 720218
rect 0 720128 800 720158
rect 9446 720120 9506 720158
rect 480069 720216 487000 720218
rect 480069 720160 480074 720216
rect 480130 720160 487000 720216
rect 480069 720158 487000 720160
rect 480069 720155 480135 720158
rect 486200 720128 487000 720158
rect 9446 720060 10060 720120
rect 0 719538 800 719568
rect 0 719478 9506 719538
rect 0 719448 800 719478
rect 9446 719304 9506 719478
rect 483790 719476 483796 719540
rect 483860 719538 483866 719540
rect 486200 719538 487000 719568
rect 483860 719478 487000 719538
rect 483860 719476 483866 719478
rect 486200 719448 487000 719478
rect 9446 719244 10060 719304
rect 482737 718858 482803 718861
rect 486200 718858 487000 718888
rect 482737 718856 487000 718858
rect 482737 718800 482742 718856
rect 482798 718800 487000 718856
rect 482737 718798 487000 718800
rect 482737 718795 482803 718798
rect 486200 718768 487000 718798
rect 9446 718372 10060 718432
rect 0 718178 800 718208
rect 9446 718178 9506 718372
rect 0 718118 9506 718178
rect 479885 718178 479951 718181
rect 486200 718178 487000 718208
rect 479885 718176 487000 718178
rect 479885 718120 479890 718176
rect 479946 718120 487000 718176
rect 479885 718118 487000 718120
rect 0 718088 800 718118
rect 479885 718115 479951 718118
rect 486200 718088 487000 718118
rect 6870 717574 10032 717634
rect 0 717498 800 717528
rect 6870 717498 6930 717574
rect 0 717438 6930 717498
rect 479333 717498 479399 717501
rect 486200 717498 487000 717528
rect 479333 717496 487000 717498
rect 479333 717440 479338 717496
rect 479394 717440 487000 717496
rect 479333 717438 487000 717440
rect 0 717408 800 717438
rect 479333 717435 479399 717438
rect 486200 717408 487000 717438
rect 477033 716954 477099 716957
rect 479425 716954 479491 716957
rect 477033 716952 479491 716954
rect 477033 716896 477038 716952
rect 477094 716896 479430 716952
rect 479486 716896 479491 716952
rect 477033 716894 479491 716896
rect 477033 716891 477099 716894
rect 479425 716891 479491 716894
rect 0 716818 800 716848
rect 482185 716818 482251 716821
rect 486200 716818 487000 716848
rect 0 716758 10032 716818
rect 482185 716816 487000 716818
rect 482185 716760 482190 716816
rect 482246 716760 487000 716816
rect 482185 716758 487000 716760
rect 0 716728 800 716758
rect 482185 716755 482251 716758
rect 486200 716728 487000 716758
rect 0 716138 800 716168
rect 0 716078 9506 716138
rect 0 716048 800 716078
rect 9446 716040 9506 716078
rect 479374 716076 479380 716140
rect 479444 716138 479450 716140
rect 486200 716138 487000 716168
rect 479444 716078 487000 716138
rect 479444 716076 479450 716078
rect 486200 716048 487000 716078
rect 9446 715980 10060 716040
rect 0 715458 800 715488
rect 0 715398 9506 715458
rect 0 715368 800 715398
rect 9446 715224 9506 715398
rect 480846 715396 480852 715460
rect 480916 715458 480922 715460
rect 486200 715458 487000 715488
rect 480916 715398 487000 715458
rect 480916 715396 480922 715398
rect 486200 715368 487000 715398
rect 9446 715164 10060 715224
rect 481030 714716 481036 714780
rect 481100 714778 481106 714780
rect 486200 714778 487000 714808
rect 481100 714718 487000 714778
rect 481100 714716 481106 714718
rect 486200 714688 487000 714718
rect 9446 714292 10060 714352
rect 0 714098 800 714128
rect 9446 714098 9506 714292
rect 0 714038 9506 714098
rect 484025 714098 484091 714101
rect 486200 714098 487000 714128
rect 484025 714096 487000 714098
rect 484025 714040 484030 714096
rect 484086 714040 487000 714096
rect 484025 714038 487000 714040
rect 0 714008 800 714038
rect 484025 714035 484091 714038
rect 486200 714008 487000 714038
rect 6870 713494 10032 713554
rect 0 713418 800 713448
rect 6870 713418 6930 713494
rect 0 713358 6930 713418
rect 477309 713418 477375 713421
rect 486200 713418 487000 713448
rect 477309 713416 487000 713418
rect 477309 713360 477314 713416
rect 477370 713360 487000 713416
rect 477309 713358 487000 713360
rect 0 713328 800 713358
rect 477309 713355 477375 713358
rect 486200 713328 487000 713358
rect 0 712738 800 712768
rect 486200 712740 487000 712768
rect 0 712678 10032 712738
rect 0 712648 800 712678
rect 486200 712676 486372 712740
rect 486436 712676 487000 712740
rect 486200 712648 487000 712676
rect 477125 712194 477191 712197
rect 482093 712194 482159 712197
rect 477125 712192 482159 712194
rect 477125 712136 477130 712192
rect 477186 712136 482098 712192
rect 482154 712136 482159 712192
rect 477125 712134 482159 712136
rect 477125 712131 477191 712134
rect 482093 712131 482159 712134
rect 0 712058 800 712088
rect 482093 712058 482159 712061
rect 486200 712058 487000 712088
rect 0 711998 9506 712058
rect 0 711968 800 711998
rect 9446 711960 9506 711998
rect 482093 712056 487000 712058
rect 482093 712000 482098 712056
rect 482154 712000 487000 712056
rect 482093 711998 487000 712000
rect 482093 711995 482159 711998
rect 486200 711968 487000 711998
rect 9446 711900 10060 711960
rect 0 711378 800 711408
rect 0 711318 9506 711378
rect 0 711288 800 711318
rect 9446 711144 9506 711318
rect 478086 711316 478092 711380
rect 478156 711378 478162 711380
rect 486200 711378 487000 711408
rect 478156 711318 487000 711378
rect 478156 711316 478162 711318
rect 486200 711288 487000 711318
rect 9446 711084 10060 711144
rect 484158 710636 484164 710700
rect 484228 710698 484234 710700
rect 486200 710698 487000 710728
rect 484228 710638 487000 710698
rect 484228 710636 484234 710638
rect 486200 710608 487000 710638
rect 9446 710212 10060 710272
rect 0 710018 800 710048
rect 9446 710018 9506 710212
rect 0 709958 9506 710018
rect 0 709928 800 709958
rect 477166 709956 477172 710020
rect 477236 710018 477242 710020
rect 486200 710018 487000 710048
rect 477236 709958 487000 710018
rect 477236 709956 477242 709958
rect 486200 709928 487000 709958
rect 6870 709414 10032 709474
rect 0 709338 800 709368
rect 6870 709338 6930 709414
rect 0 709278 6930 709338
rect 0 709248 800 709278
rect 478270 709276 478276 709340
rect 478340 709338 478346 709340
rect 486200 709338 487000 709368
rect 478340 709278 487000 709338
rect 478340 709276 478346 709278
rect 486200 709248 487000 709278
rect 477401 709202 477467 709205
rect 482185 709202 482251 709205
rect 477401 709200 482251 709202
rect 477401 709144 477406 709200
rect 477462 709144 482190 709200
rect 482246 709144 482251 709200
rect 477401 709142 482251 709144
rect 477401 709139 477467 709142
rect 482185 709139 482251 709142
rect 0 708658 800 708688
rect 0 708598 10032 708658
rect 0 708568 800 708598
rect 485998 708596 486004 708660
rect 486068 708658 486074 708660
rect 486200 708658 487000 708688
rect 486068 708598 487000 708658
rect 486068 708596 486074 708598
rect 486200 708568 487000 708598
rect 0 707978 800 708008
rect 0 707918 4170 707978
rect 0 707888 800 707918
rect 4110 707842 4170 707918
rect 485814 707916 485820 707980
rect 485884 707978 485890 707980
rect 486200 707978 487000 708008
rect 485884 707918 487000 707978
rect 485884 707916 485890 707918
rect 486200 707888 487000 707918
rect 4110 707782 10032 707842
rect 0 707298 800 707328
rect 0 707238 9506 707298
rect 0 707208 800 707238
rect 9446 707064 9506 707238
rect 478454 707236 478460 707300
rect 478524 707298 478530 707300
rect 486200 707298 487000 707328
rect 478524 707238 487000 707298
rect 478524 707236 478530 707238
rect 486200 707208 487000 707238
rect 9446 707004 10060 707064
rect 485078 706556 485084 706620
rect 485148 706618 485154 706620
rect 486200 706618 487000 706648
rect 485148 706558 487000 706618
rect 485148 706556 485154 706558
rect 486200 706528 487000 706558
rect 9446 706132 10060 706192
rect 0 705938 800 705968
rect 9446 705938 9506 706132
rect 0 705878 9506 705938
rect 0 705848 800 705878
rect 485262 705876 485268 705940
rect 485332 705938 485338 705940
rect 486200 705938 487000 705968
rect 485332 705878 487000 705938
rect 485332 705876 485338 705878
rect 486200 705848 487000 705878
rect 9446 705316 10060 705376
rect 0 705258 800 705288
rect 9446 705258 9506 705316
rect 0 705198 9506 705258
rect 0 705168 800 705198
rect 481398 705196 481404 705260
rect 481468 705258 481474 705260
rect 486200 705258 487000 705288
rect 481468 705198 487000 705258
rect 481468 705196 481474 705198
rect 486200 705168 487000 705198
rect 0 704578 800 704608
rect 0 704518 10032 704578
rect 0 704488 800 704518
rect 485630 704516 485636 704580
rect 485700 704578 485706 704580
rect 486200 704578 487000 704608
rect 485700 704518 487000 704578
rect 485700 704516 485706 704518
rect 486200 704488 487000 704518
rect 0 703898 800 703928
rect 486200 703901 487000 703928
rect 0 703838 4170 703898
rect 0 703808 800 703838
rect 4110 703762 4170 703838
rect 486141 703896 487000 703901
rect 486141 703840 486146 703896
rect 486202 703840 487000 703896
rect 486141 703835 487000 703840
rect 486200 703808 487000 703835
rect 482185 703762 482251 703765
rect 482870 703762 482876 703764
rect 4110 703702 10032 703762
rect 482185 703760 482876 703762
rect 482185 703704 482190 703760
rect 482246 703704 482876 703760
rect 482185 703702 482876 703704
rect 482185 703699 482251 703702
rect 482870 703700 482876 703702
rect 482940 703700 482946 703764
rect 0 703218 800 703248
rect 0 703158 9506 703218
rect 0 703128 800 703158
rect 9446 702984 9506 703158
rect 485446 703156 485452 703220
rect 485516 703218 485522 703220
rect 486200 703218 487000 703248
rect 485516 703158 487000 703218
rect 485516 703156 485522 703158
rect 486200 703128 487000 703158
rect 9446 702924 10060 702984
rect 479742 702476 479748 702540
rect 479812 702538 479818 702540
rect 486200 702538 487000 702568
rect 479812 702478 487000 702538
rect 479812 702476 479818 702478
rect 486200 702448 487000 702478
rect 9446 702052 10060 702112
rect 0 701858 800 701888
rect 9446 701858 9506 702052
rect 0 701798 9506 701858
rect 483473 701858 483539 701861
rect 486200 701858 487000 701888
rect 483473 701856 487000 701858
rect 483473 701800 483478 701856
rect 483534 701800 487000 701856
rect 483473 701798 487000 701800
rect 0 701768 800 701798
rect 483473 701795 483539 701798
rect 486200 701768 487000 701798
rect 9446 701236 10060 701296
rect 0 701178 800 701208
rect 9446 701178 9506 701236
rect 0 701118 9506 701178
rect 486200 701180 487000 701208
rect 0 701088 800 701118
rect 486200 701116 486372 701180
rect 486436 701116 487000 701180
rect 486200 701088 487000 701116
rect 0 700498 800 700528
rect 0 700438 10032 700498
rect 0 700408 800 700438
rect 479926 700436 479932 700500
rect 479996 700498 480002 700500
rect 486200 700498 487000 700528
rect 479996 700438 487000 700498
rect 479996 700436 480002 700438
rect 486200 700408 487000 700438
rect 0 699818 800 699848
rect 483565 699818 483631 699821
rect 486200 699818 487000 699848
rect 0 699758 4170 699818
rect 0 699728 800 699758
rect 4110 699682 4170 699758
rect 483565 699816 487000 699818
rect 483565 699760 483570 699816
rect 483626 699760 487000 699816
rect 483565 699758 487000 699760
rect 483565 699755 483631 699758
rect 486200 699728 487000 699758
rect 4110 699622 10032 699682
rect 478638 699348 478644 699412
rect 478708 699410 478714 699412
rect 484894 699410 484900 699412
rect 478708 699350 484900 699410
rect 478708 699348 478714 699350
rect 484894 699348 484900 699350
rect 484964 699348 484970 699412
rect 0 699138 800 699168
rect 0 699078 9506 699138
rect 0 699048 800 699078
rect 9446 698904 9506 699078
rect 482870 699076 482876 699140
rect 482940 699138 482946 699140
rect 486200 699138 487000 699168
rect 482940 699078 487000 699138
rect 482940 699076 482946 699078
rect 486200 699048 487000 699078
rect 9446 698844 10060 698904
rect 482318 698396 482324 698460
rect 482388 698458 482394 698460
rect 486200 698458 487000 698488
rect 482388 698398 487000 698458
rect 482388 698396 482394 698398
rect 486200 698368 487000 698398
rect 479425 698322 479491 698325
rect 480110 698322 480116 698324
rect 479425 698320 480116 698322
rect 479425 698264 479430 698320
rect 479486 698264 480116 698320
rect 479425 698262 480116 698264
rect 479425 698259 479491 698262
rect 480110 698260 480116 698262
rect 480180 698260 480186 698324
rect 478638 698186 478644 698188
rect 476968 698126 478644 698186
rect 478638 698124 478644 698126
rect 478708 698124 478714 698188
rect 9446 697972 10060 698032
rect 0 697778 800 697808
rect 9446 697778 9506 697972
rect 485262 697914 485268 697916
rect 476968 697854 485268 697914
rect 485262 697852 485268 697854
rect 485332 697852 485338 697916
rect 486200 697778 487000 697808
rect 0 697718 9506 697778
rect 477358 697718 487000 697778
rect 0 697688 800 697718
rect 477358 697710 477418 697718
rect 476940 697650 477418 697710
rect 486200 697688 487000 697718
rect 483606 697370 483612 697372
rect 476968 697310 483612 697370
rect 483606 697308 483612 697310
rect 483676 697308 483682 697372
rect 483974 697234 483980 697236
rect 9446 697156 10060 697216
rect 477358 697174 483980 697234
rect 477358 697166 477418 697174
rect 483974 697172 483980 697174
rect 484044 697172 484050 697236
rect 0 697098 800 697128
rect 9446 697098 9506 697156
rect 476940 697106 477418 697166
rect 0 697038 9506 697098
rect 0 697008 800 697038
rect 483422 697036 483428 697100
rect 483492 697098 483498 697100
rect 486200 697098 487000 697128
rect 483492 697038 487000 697098
rect 483492 697036 483498 697038
rect 486200 697008 487000 697038
rect 477534 696900 477540 696964
rect 477604 696962 477610 696964
rect 477953 696962 478019 696965
rect 477604 696960 478019 696962
rect 477604 696904 477958 696960
rect 478014 696904 478019 696960
rect 477604 696902 478019 696904
rect 477604 696900 477610 696902
rect 477953 696899 478019 696902
rect 483606 696900 483612 696964
rect 483676 696962 483682 696964
rect 483841 696962 483907 696965
rect 483676 696960 483907 696962
rect 483676 696904 483846 696960
rect 483902 696904 483907 696960
rect 483676 696902 483907 696904
rect 483676 696900 483682 696902
rect 483841 696899 483907 696902
rect 483790 696826 483796 696828
rect 476968 696766 483796 696826
rect 483790 696764 483796 696766
rect 483860 696764 483866 696828
rect 485814 696554 485820 696556
rect 476968 696494 485820 696554
rect 485814 696492 485820 696494
rect 485884 696492 485890 696556
rect 0 696418 800 696448
rect 0 696358 10032 696418
rect 0 696328 800 696358
rect 481582 696356 481588 696420
rect 481652 696418 481658 696420
rect 486200 696418 487000 696448
rect 481652 696358 487000 696418
rect 481652 696356 481658 696358
rect 486200 696328 487000 696358
rect 482870 696282 482876 696284
rect 476968 696222 482876 696282
rect 482870 696220 482876 696222
rect 482940 696220 482946 696284
rect 482369 696010 482435 696013
rect 476968 696008 482435 696010
rect 476968 695952 482374 696008
rect 482430 695952 482435 696008
rect 476968 695950 482435 695952
rect 482369 695947 482435 695950
rect 477309 695806 477375 695809
rect 476940 695804 477375 695806
rect 476940 695748 477314 695804
rect 477370 695748 477375 695804
rect 476940 695746 477375 695748
rect 477309 695743 477375 695746
rect 485262 695676 485268 695740
rect 485332 695738 485338 695740
rect 486200 695738 487000 695768
rect 485332 695678 487000 695738
rect 485332 695676 485338 695678
rect 486200 695648 487000 695678
rect 478822 695540 478828 695604
rect 478892 695602 478898 695604
rect 479333 695602 479399 695605
rect 478892 695600 479399 695602
rect 478892 695544 479338 695600
rect 479394 695544 479399 695600
rect 478892 695542 479399 695544
rect 478892 695540 478898 695542
rect 479333 695539 479399 695542
rect 482645 695466 482711 695469
rect 476968 695464 482711 695466
rect 476968 695408 482650 695464
rect 482706 695408 482711 695464
rect 476968 695406 482711 695408
rect 482645 695403 482711 695406
rect 485446 695194 485452 695196
rect 476968 695134 485452 695194
rect 485446 695132 485452 695134
rect 485516 695132 485522 695196
rect 482001 695058 482067 695061
rect 486200 695058 487000 695088
rect 482001 695056 487000 695058
rect 482001 695000 482006 695056
rect 482062 695000 487000 695056
rect 482001 694998 487000 695000
rect 482001 694995 482067 694998
rect 486200 694968 487000 694998
rect 478270 694922 478276 694924
rect 476968 694862 478276 694922
rect 478270 694860 478276 694862
rect 478340 694860 478346 694924
rect 482461 694650 482527 694653
rect 476968 694648 482527 694650
rect 476968 694592 482466 694648
rect 482522 694592 482527 694648
rect 476968 694590 482527 694592
rect 482461 694587 482527 694590
rect 485630 694514 485636 694516
rect 477358 694454 485636 694514
rect 477358 694446 477418 694454
rect 485630 694452 485636 694454
rect 485700 694452 485706 694516
rect 476940 694386 477418 694446
rect 482829 694378 482895 694381
rect 486200 694378 487000 694408
rect 482829 694376 487000 694378
rect 482829 694320 482834 694376
rect 482890 694320 487000 694376
rect 482829 694318 487000 694320
rect 482829 694315 482895 694318
rect 486200 694288 487000 694318
rect 477718 694180 477724 694244
rect 477788 694242 477794 694244
rect 478045 694242 478111 694245
rect 482921 694242 482987 694245
rect 477788 694240 478111 694242
rect 477788 694184 478050 694240
rect 478106 694184 478111 694240
rect 477788 694182 478111 694184
rect 477788 694180 477794 694182
rect 478045 694179 478111 694182
rect 482878 694240 482987 694242
rect 482878 694184 482926 694240
rect 482982 694184 482987 694240
rect 482878 694179 482987 694184
rect 482878 694106 482938 694179
rect 476968 694046 482938 694106
rect 483974 694044 483980 694108
rect 484044 694106 484050 694108
rect 484117 694106 484183 694109
rect 484044 694104 484183 694106
rect 484044 694048 484122 694104
rect 484178 694048 484183 694104
rect 484044 694046 484183 694048
rect 484044 694044 484050 694046
rect 484117 694043 484183 694046
rect 485998 693834 486004 693836
rect 476968 693774 486004 693834
rect 485998 693772 486004 693774
rect 486068 693772 486074 693836
rect 486200 693698 487000 693728
rect 477358 693638 487000 693698
rect 477358 693630 477418 693638
rect 476940 693570 477418 693630
rect 486200 693608 487000 693638
rect 480478 693500 480484 693564
rect 480548 693562 480554 693564
rect 481030 693562 481036 693564
rect 480548 693502 481036 693562
rect 480548 693500 480554 693502
rect 481030 693500 481036 693502
rect 481100 693500 481106 693564
rect 480846 693364 480852 693428
rect 480916 693364 480922 693428
rect 476924 693228 476930 693292
rect 476994 693228 477000 693292
rect 480854 693156 480914 693364
rect 480846 693092 480852 693156
rect 480916 693092 480922 693156
rect 479701 693018 479767 693021
rect 476968 693016 479767 693018
rect 476968 692960 479706 693016
rect 479762 692960 479767 693016
rect 476968 692958 479767 692960
rect 479701 692955 479767 692958
rect 482134 692956 482140 693020
rect 482204 693018 482210 693020
rect 486200 693018 487000 693048
rect 482204 692958 487000 693018
rect 482204 692956 482210 692958
rect 486200 692928 487000 692958
rect 482553 692882 482619 692885
rect 482510 692880 482619 692882
rect 482510 692824 482558 692880
rect 482614 692824 482619 692880
rect 482510 692819 482619 692824
rect 476968 692686 477234 692746
rect 477174 692610 477234 692686
rect 481214 692684 481220 692748
rect 481284 692746 481290 692748
rect 481357 692746 481423 692749
rect 481284 692744 481423 692746
rect 481284 692688 481362 692744
rect 481418 692688 481423 692744
rect 481284 692686 481423 692688
rect 481284 692684 481290 692686
rect 481357 692683 481423 692686
rect 482510 692610 482570 692819
rect 482921 692746 482987 692749
rect 486141 692746 486207 692749
rect 482921 692744 486207 692746
rect 482921 692688 482926 692744
rect 482982 692688 486146 692744
rect 486202 692688 486207 692744
rect 482921 692686 486207 692688
rect 482921 692683 482987 692686
rect 486141 692683 486207 692686
rect 477174 692550 482570 692610
rect 482277 692474 482343 692477
rect 476968 692472 482343 692474
rect 476968 692416 482282 692472
rect 482338 692416 482343 692472
rect 476968 692414 482343 692416
rect 482277 692411 482343 692414
rect 477166 692276 477172 692340
rect 477236 692338 477242 692340
rect 477401 692338 477467 692341
rect 477236 692336 477467 692338
rect 477236 692280 477406 692336
rect 477462 692280 477467 692336
rect 477236 692278 477467 692280
rect 477236 692276 477242 692278
rect 477401 692275 477467 692278
rect 478638 692276 478644 692340
rect 478708 692338 478714 692340
rect 486200 692338 487000 692368
rect 478708 692278 487000 692338
rect 478708 692276 478714 692278
rect 486200 692248 487000 692278
rect 485998 692202 486004 692204
rect 476968 692142 486004 692202
rect 485998 692140 486004 692142
rect 486068 692140 486074 692204
rect 478086 691930 478092 691932
rect 476968 691870 478092 691930
rect 478086 691868 478092 691870
rect 478156 691868 478162 691932
rect 481582 691658 481588 691660
rect 476968 691598 481588 691658
rect 481582 691596 481588 691598
rect 481652 691596 481658 691660
rect 485814 691596 485820 691660
rect 485884 691658 485890 691660
rect 486200 691658 487000 691688
rect 485884 691598 487000 691658
rect 485884 691596 485890 691598
rect 486200 691568 487000 691598
rect 476968 691326 477786 691386
rect 477726 691250 477786 691326
rect 477902 691324 477908 691388
rect 477972 691386 477978 691388
rect 478229 691386 478295 691389
rect 477972 691384 478295 691386
rect 477972 691328 478234 691384
rect 478290 691328 478295 691384
rect 477972 691326 478295 691328
rect 477972 691324 477978 691326
rect 478229 691323 478295 691326
rect 483749 691250 483815 691253
rect 477726 691248 483815 691250
rect 477726 691192 483754 691248
rect 483810 691192 483815 691248
rect 477726 691190 483815 691192
rect 483749 691187 483815 691190
rect 478638 691114 478644 691116
rect 476968 691054 478644 691114
rect 478638 691052 478644 691054
rect 478708 691052 478714 691116
rect 484342 690916 484348 690980
rect 484412 690978 484418 690980
rect 486200 690978 487000 691008
rect 484412 690918 487000 690978
rect 484412 690916 484418 690918
rect 486200 690888 487000 690918
rect 483974 690842 483980 690844
rect 476968 690782 483980 690842
rect 483974 690780 483980 690782
rect 484044 690780 484050 690844
rect 483606 690570 483612 690572
rect 476968 690510 483612 690570
rect 483606 690508 483612 690510
rect 483676 690508 483682 690572
rect 483933 690434 483999 690437
rect 477358 690432 483999 690434
rect 477358 690376 483938 690432
rect 483994 690376 483999 690432
rect 477358 690374 483999 690376
rect 477358 690366 477418 690374
rect 483933 690371 483999 690374
rect 476940 690306 477418 690366
rect 483606 690236 483612 690300
rect 483676 690298 483682 690300
rect 486200 690298 487000 690328
rect 483676 690238 487000 690298
rect 483676 690236 483682 690238
rect 486200 690208 487000 690238
rect 476968 689966 480178 690026
rect 480118 689890 480178 689966
rect 480294 689964 480300 690028
rect 480364 690026 480370 690028
rect 480805 690026 480871 690029
rect 480364 690024 480871 690026
rect 480364 689968 480810 690024
rect 480866 689968 480871 690024
rect 480364 689966 480871 689968
rect 480364 689964 480370 689966
rect 480805 689963 480871 689966
rect 483054 689964 483060 690028
rect 483124 690026 483130 690028
rect 483565 690026 483631 690029
rect 483124 690024 483631 690026
rect 483124 689968 483570 690024
rect 483626 689968 483631 690024
rect 483124 689966 483631 689968
rect 483124 689964 483130 689966
rect 483565 689963 483631 689966
rect 482277 689890 482343 689893
rect 486325 689890 486391 689893
rect 480118 689830 482202 689890
rect 481909 689754 481975 689757
rect 476968 689752 481975 689754
rect 476968 689696 481914 689752
rect 481970 689696 481975 689752
rect 476968 689694 481975 689696
rect 482142 689754 482202 689830
rect 482277 689888 486391 689890
rect 482277 689832 482282 689888
rect 482338 689832 486330 689888
rect 486386 689832 486391 689888
rect 482277 689830 486391 689832
rect 482277 689827 482343 689830
rect 486325 689827 486391 689830
rect 484158 689754 484164 689756
rect 482142 689694 484164 689754
rect 481909 689691 481975 689694
rect 484158 689692 484164 689694
rect 484228 689692 484234 689756
rect 486200 689618 487000 689648
rect 477358 689558 487000 689618
rect 477358 689550 477418 689558
rect 476940 689490 477418 689550
rect 486200 689528 487000 689558
rect 482093 689210 482159 689213
rect 476968 689208 482159 689210
rect 476968 689152 482098 689208
rect 482154 689152 482159 689208
rect 476968 689150 482159 689152
rect 482093 689147 482159 689150
rect 481214 689074 481220 689076
rect 477174 689014 481220 689074
rect 477174 689006 477234 689014
rect 481214 689012 481220 689014
rect 481284 689012 481290 689076
rect 476940 688946 477234 689006
rect 486200 688938 487000 688968
rect 477358 688878 487000 688938
rect 477358 688734 477418 688878
rect 486200 688848 487000 688878
rect 476940 688674 477418 688734
rect 480897 688394 480963 688397
rect 476968 688392 480963 688394
rect 476968 688336 480902 688392
rect 480958 688336 480963 688392
rect 476968 688334 480963 688336
rect 480897 688331 480963 688334
rect 0 688258 800 688288
rect 0 688198 9506 688258
rect 0 688168 800 688198
rect 9446 688176 9506 688198
rect 481030 688196 481036 688260
rect 481100 688258 481106 688260
rect 486200 688258 487000 688288
rect 481100 688198 487000 688258
rect 481100 688196 481106 688198
rect 9446 688116 10060 688176
rect 486200 688168 487000 688198
rect 485262 688122 485268 688124
rect 476968 688062 485268 688122
rect 485262 688060 485268 688062
rect 485332 688060 485338 688124
rect 481173 687850 481239 687853
rect 476968 687848 481239 687850
rect 476968 687792 481178 687848
rect 481234 687792 481239 687848
rect 476968 687790 481239 687792
rect 481173 687787 481239 687790
rect 0 687578 800 687608
rect 480478 687578 480484 687580
rect 0 687518 9506 687578
rect 476968 687518 480484 687578
rect 0 687488 800 687518
rect 9446 687374 9506 687518
rect 480478 687516 480484 687518
rect 480548 687516 480554 687580
rect 486200 687578 487000 687608
rect 483246 687518 487000 687578
rect 483246 687442 483306 687518
rect 486200 687488 487000 687518
rect 477358 687382 483306 687442
rect 477358 687374 477418 687382
rect 9446 687314 10060 687374
rect 476940 687314 477418 687374
rect 481214 687108 481220 687172
rect 481284 687170 481290 687172
rect 485630 687170 485636 687172
rect 481284 687110 485636 687170
rect 481284 687108 481290 687110
rect 485630 687108 485636 687110
rect 485700 687108 485706 687172
rect 480846 687034 480852 687036
rect 476968 686974 480852 687034
rect 480846 686972 480852 686974
rect 480916 686972 480922 687036
rect 485446 686836 485452 686900
rect 485516 686898 485522 686900
rect 486200 686898 487000 686928
rect 485516 686838 487000 686898
rect 485516 686836 485522 686838
rect 486200 686808 487000 686838
rect 482318 686762 482324 686764
rect 476968 686702 482324 686762
rect 482318 686700 482324 686702
rect 482388 686700 482394 686764
rect 479374 686490 479380 686492
rect 6870 686430 10032 686490
rect 476968 686430 479380 686490
rect 0 686218 800 686248
rect 6870 686218 6930 686430
rect 479374 686428 479380 686430
rect 479444 686428 479450 686492
rect 479977 686218 480043 686221
rect 0 686158 6930 686218
rect 476968 686216 480043 686218
rect 476968 686160 479982 686216
rect 480038 686160 480043 686216
rect 476968 686158 480043 686160
rect 0 686128 800 686158
rect 479977 686155 480043 686158
rect 483238 686156 483244 686220
rect 483308 686218 483314 686220
rect 486200 686218 487000 686248
rect 483308 686158 487000 686218
rect 483308 686156 483314 686158
rect 486200 686128 487000 686158
rect 479793 685946 479859 685949
rect 476968 685944 479859 685946
rect 476968 685888 479798 685944
rect 479854 685888 479859 685944
rect 476968 685886 479859 685888
rect 479793 685883 479859 685886
rect 479558 685748 479564 685812
rect 479628 685810 479634 685812
rect 480161 685810 480227 685813
rect 479628 685808 480227 685810
rect 479628 685752 480166 685808
rect 480222 685752 480227 685808
rect 479628 685750 480227 685752
rect 479628 685748 479634 685750
rect 480161 685747 480227 685750
rect 481582 685748 481588 685812
rect 481652 685810 481658 685812
rect 482829 685810 482895 685813
rect 481652 685808 482895 685810
rect 481652 685752 482834 685808
rect 482890 685752 482895 685808
rect 481652 685750 482895 685752
rect 481652 685748 481658 685750
rect 482829 685747 482895 685750
rect 478822 685674 478828 685676
rect 6870 685614 10032 685674
rect 476968 685614 478828 685674
rect 0 685538 800 685568
rect 6870 685538 6930 685614
rect 478822 685612 478828 685614
rect 478892 685612 478898 685676
rect 0 685478 6930 685538
rect 0 685448 800 685478
rect 480110 685476 480116 685540
rect 480180 685538 480186 685540
rect 486200 685538 487000 685568
rect 480180 685478 487000 685538
rect 480180 685476 480186 685478
rect 486200 685448 487000 685478
rect 479742 685402 479748 685404
rect 476968 685342 479748 685402
rect 479742 685340 479748 685342
rect 479812 685340 479818 685404
rect 480161 685266 480227 685269
rect 486233 685266 486299 685269
rect 480161 685264 486299 685266
rect 480161 685208 480166 685264
rect 480222 685208 486238 685264
rect 486294 685208 486299 685264
rect 480161 685206 486299 685208
rect 480161 685203 480227 685206
rect 486233 685203 486299 685206
rect 479885 685130 479951 685133
rect 476968 685128 479951 685130
rect 476968 685072 479890 685128
rect 479946 685072 479951 685128
rect 476968 685070 479951 685072
rect 479885 685067 479951 685070
rect 480253 685130 480319 685133
rect 486417 685130 486483 685133
rect 480253 685128 486483 685130
rect 480253 685072 480258 685128
rect 480314 685072 486422 685128
rect 486478 685072 486483 685128
rect 480253 685070 486483 685072
rect 480253 685067 480319 685070
rect 486417 685067 486483 685070
rect 479609 684994 479675 684997
rect 477358 684992 479675 684994
rect 477358 684936 479614 684992
rect 479670 684936 479675 684992
rect 477358 684934 479675 684936
rect 477358 684926 477418 684934
rect 479609 684931 479675 684934
rect 0 684858 800 684888
rect 476940 684866 477418 684926
rect 0 684798 10032 684858
rect 0 684768 800 684798
rect 479374 684796 479380 684860
rect 479444 684858 479450 684860
rect 486200 684858 487000 684888
rect 479444 684798 487000 684858
rect 479444 684796 479450 684798
rect 486200 684768 487000 684798
rect 483238 684722 483244 684724
rect 477358 684662 483244 684722
rect 477358 684654 477418 684662
rect 483238 684660 483244 684662
rect 483308 684660 483314 684724
rect 476940 684594 477418 684654
rect 483238 684524 483244 684588
rect 483308 684586 483314 684588
rect 483606 684586 483612 684588
rect 483308 684526 483612 684586
rect 483308 684524 483314 684526
rect 483606 684524 483612 684526
rect 483676 684524 483682 684588
rect 478270 684388 478276 684452
rect 478340 684450 478346 684452
rect 478413 684450 478479 684453
rect 478340 684448 478479 684450
rect 478340 684392 478418 684448
rect 478474 684392 478479 684448
rect 478340 684390 478479 684392
rect 478340 684388 478346 684390
rect 478413 684387 478479 684390
rect 483473 684450 483539 684453
rect 483606 684450 483612 684452
rect 483473 684448 483612 684450
rect 483473 684392 483478 684448
rect 483534 684392 483612 684448
rect 483473 684390 483612 684392
rect 483473 684387 483539 684390
rect 483606 684388 483612 684390
rect 483676 684388 483682 684452
rect 479517 684314 479583 684317
rect 476968 684312 479583 684314
rect 476968 684256 479522 684312
rect 479578 684256 479583 684312
rect 476968 684254 479583 684256
rect 479517 684251 479583 684254
rect 0 684178 800 684208
rect 0 684118 9506 684178
rect 0 684088 800 684118
rect 9446 684110 9506 684118
rect 479742 684116 479748 684180
rect 479812 684178 479818 684180
rect 486200 684178 487000 684208
rect 479812 684118 487000 684178
rect 479812 684116 479818 684118
rect 9446 684050 10060 684110
rect 486200 684088 487000 684118
rect 479926 684042 479932 684044
rect 476968 683982 479932 684042
rect 479926 683980 479932 683982
rect 479996 683980 480002 684044
rect 479558 683770 479564 683772
rect 476968 683710 479564 683770
rect 479558 683708 479564 683710
rect 479628 683708 479634 683772
rect 0 683498 800 683528
rect 477534 683498 477540 683500
rect 0 683438 9506 683498
rect 476968 683438 477540 683498
rect 0 683408 800 683438
rect 9446 683294 9506 683438
rect 477534 683436 477540 683438
rect 477604 683436 477610 683500
rect 484710 683436 484716 683500
rect 484780 683498 484786 683500
rect 486200 683498 487000 683528
rect 484780 683438 487000 683498
rect 484780 683436 484786 683438
rect 486200 683408 487000 683438
rect 9446 683234 10060 683294
rect 484342 683226 484348 683228
rect 476968 683166 484348 683226
rect 484342 683164 484348 683166
rect 484412 683164 484418 683228
rect 477718 682954 477724 682956
rect 476968 682894 477724 682954
rect 477718 682892 477724 682894
rect 477788 682892 477794 682956
rect 484526 682756 484532 682820
rect 484596 682818 484602 682820
rect 486200 682818 487000 682848
rect 484596 682758 487000 682818
rect 484596 682756 484602 682758
rect 486200 682728 487000 682758
rect 481398 682682 481404 682684
rect 476968 682622 481404 682682
rect 481398 682620 481404 682622
rect 481468 682620 481474 682684
rect 481265 682410 481331 682413
rect 6870 682350 10032 682410
rect 476968 682408 481331 682410
rect 476968 682352 481270 682408
rect 481326 682352 481331 682408
rect 476968 682350 481331 682352
rect 0 682138 800 682168
rect 6870 682138 6930 682350
rect 481265 682347 481331 682350
rect 480989 682138 481055 682141
rect 0 682078 6930 682138
rect 476968 682136 481055 682138
rect 476968 682080 480994 682136
rect 481050 682080 481055 682136
rect 476968 682078 481055 682080
rect 0 682048 800 682078
rect 480989 682075 481055 682078
rect 484342 682076 484348 682140
rect 484412 682138 484418 682140
rect 486200 682138 487000 682168
rect 484412 682078 487000 682138
rect 484412 682076 484418 682078
rect 486200 682048 487000 682078
rect 484710 682002 484716 682004
rect 477358 681942 484716 682002
rect 477358 681934 477418 681942
rect 484710 681940 484716 681942
rect 484780 681940 484786 682004
rect 476940 681874 477418 681934
rect 478086 681804 478092 681868
rect 478156 681866 478162 681868
rect 478505 681866 478571 681869
rect 478156 681864 478571 681866
rect 478156 681808 478510 681864
rect 478566 681808 478571 681864
rect 478156 681806 478571 681808
rect 478156 681804 478162 681806
rect 478505 681803 478571 681806
rect 481081 681594 481147 681597
rect 6870 681534 10032 681594
rect 476968 681592 481147 681594
rect 476968 681536 481086 681592
rect 481142 681536 481147 681592
rect 476968 681534 481147 681536
rect 0 681458 800 681488
rect 6870 681458 6930 681534
rect 481081 681531 481147 681534
rect 0 681398 6930 681458
rect 0 681368 800 681398
rect 485630 681396 485636 681460
rect 485700 681458 485706 681460
rect 486200 681458 487000 681488
rect 485700 681398 487000 681458
rect 485700 681396 485706 681398
rect 486200 681368 487000 681398
rect 484342 681322 484348 681324
rect 476968 681262 484348 681322
rect 484342 681260 484348 681262
rect 484412 681260 484418 681324
rect 480294 681186 480300 681188
rect 477358 681126 480300 681186
rect 477358 681118 477418 681126
rect 480294 681124 480300 681126
rect 480364 681124 480370 681188
rect 476940 681058 477418 681118
rect 482134 680914 482140 680916
rect 477358 680854 482140 680914
rect 477358 680846 477418 680854
rect 482134 680852 482140 680854
rect 482204 680852 482210 680916
rect 0 680778 800 680808
rect 476940 680786 477418 680846
rect 0 680718 10032 680778
rect 0 680688 800 680718
rect 481398 680716 481404 680780
rect 481468 680778 481474 680780
rect 486200 680778 487000 680808
rect 481468 680718 487000 680778
rect 481468 680716 481474 680718
rect 486200 680688 487000 680718
rect 480110 680506 480116 680508
rect 476968 680446 480116 680506
rect 480110 680444 480116 680446
rect 480180 680444 480186 680508
rect 479190 680308 479196 680372
rect 479260 680370 479266 680372
rect 480069 680370 480135 680373
rect 479260 680368 480135 680370
rect 479260 680312 480074 680368
rect 480130 680312 480135 680368
rect 479260 680310 480135 680312
rect 479260 680308 479266 680310
rect 480069 680307 480135 680310
rect 482134 680308 482140 680372
rect 482204 680370 482210 680372
rect 482921 680370 482987 680373
rect 482204 680368 482987 680370
rect 482204 680312 482926 680368
rect 482982 680312 482987 680368
rect 482204 680310 482987 680312
rect 482204 680308 482210 680310
rect 482921 680307 482987 680310
rect 478137 680234 478203 680237
rect 476968 680232 478203 680234
rect 476968 680176 478142 680232
rect 478198 680176 478203 680232
rect 476968 680174 478203 680176
rect 478137 680171 478203 680174
rect 0 680098 800 680128
rect 486200 680100 487000 680128
rect 0 680038 9506 680098
rect 0 680008 800 680038
rect 9446 680030 9506 680038
rect 486200 680036 486372 680100
rect 486436 680036 487000 680100
rect 9446 679970 10060 680030
rect 486200 680008 487000 680036
rect 478270 679962 478276 679964
rect 476968 679902 478276 679962
rect 478270 679900 478276 679902
rect 478340 679900 478346 679964
rect 478321 679826 478387 679829
rect 477358 679824 478387 679826
rect 477358 679768 478326 679824
rect 478382 679768 478387 679824
rect 477358 679766 478387 679768
rect 477358 679758 477418 679766
rect 478321 679763 478387 679766
rect 476940 679698 477418 679758
rect 477718 679628 477724 679692
rect 477788 679690 477794 679692
rect 485078 679690 485084 679692
rect 477788 679630 485084 679690
rect 477788 679628 477794 679630
rect 485078 679628 485084 679630
rect 485148 679628 485154 679692
rect 485814 679554 485820 679556
rect 477358 679494 485820 679554
rect 477358 679486 477418 679494
rect 485814 679492 485820 679494
rect 485884 679492 485890 679556
rect 0 679418 800 679448
rect 476940 679426 477418 679486
rect 0 679358 9506 679418
rect 0 679328 800 679358
rect 9446 679214 9506 679358
rect 9446 679154 10060 679214
rect 478454 679146 478460 679148
rect 476968 679086 478460 679146
rect 478454 679084 478460 679086
rect 478524 679084 478530 679148
rect 483054 679084 483060 679148
rect 483124 679146 483130 679148
rect 483790 679146 483796 679148
rect 483124 679086 483796 679146
rect 483124 679084 483130 679086
rect 483790 679084 483796 679086
rect 483860 679084 483866 679148
rect 478689 679010 478755 679013
rect 478646 679008 478755 679010
rect 478646 678952 478694 679008
rect 478750 678952 478755 679008
rect 478646 678947 478755 678952
rect 481950 678948 481956 679012
rect 482020 679010 482026 679012
rect 482737 679010 482803 679013
rect 482020 679008 482803 679010
rect 482020 678952 482742 679008
rect 482798 678952 482803 679008
rect 482020 678950 482803 678952
rect 482020 678948 482026 678950
rect 482737 678947 482803 678950
rect 477902 678874 477908 678876
rect 476968 678814 477908 678874
rect 477902 678812 477908 678814
rect 477972 678812 477978 678876
rect 478646 678738 478706 678947
rect 477358 678678 478706 678738
rect 477358 678670 477418 678678
rect 476940 678610 477418 678670
rect 478454 678404 478460 678468
rect 478524 678466 478530 678468
rect 478597 678466 478663 678469
rect 478524 678464 478663 678466
rect 478524 678408 478602 678464
rect 478658 678408 478663 678464
rect 478524 678406 478663 678408
rect 478524 678404 478530 678406
rect 478597 678403 478663 678406
rect 483054 678404 483060 678468
rect 483124 678466 483130 678468
rect 483422 678466 483428 678468
rect 483124 678406 483428 678466
rect 483124 678404 483130 678406
rect 483422 678404 483428 678406
rect 483492 678404 483498 678468
rect 482001 678330 482067 678333
rect 6870 678270 10032 678330
rect 476968 678328 482067 678330
rect 476968 678272 482006 678328
rect 482062 678272 482067 678328
rect 476968 678270 482067 678272
rect 0 678058 800 678088
rect 6870 678058 6930 678270
rect 482001 678267 482067 678270
rect 481766 678132 481772 678196
rect 481836 678194 481842 678196
rect 482185 678194 482251 678197
rect 481836 678192 482251 678194
rect 481836 678136 482190 678192
rect 482246 678136 482251 678192
rect 481836 678134 482251 678136
rect 481836 678132 481842 678134
rect 482185 678131 482251 678134
rect 478086 678058 478092 678060
rect 0 677998 6930 678058
rect 476968 677998 478092 678058
rect 0 677968 800 677998
rect 478086 677996 478092 677998
rect 478156 677996 478162 678060
rect 481398 677786 481404 677788
rect 476968 677726 481404 677786
rect 481398 677724 481404 677726
rect 481468 677724 481474 677788
rect 478781 677650 478847 677653
rect 477542 677648 478847 677650
rect 477542 677592 478786 677648
rect 478842 677592 478847 677648
rect 477542 677590 478847 677592
rect 477542 677582 477602 677590
rect 478781 677587 478847 677590
rect 476940 677522 477602 677582
rect 6870 677454 10032 677514
rect 0 677378 800 677408
rect 6870 677378 6930 677454
rect 479006 677452 479012 677516
rect 479076 677514 479082 677516
rect 479425 677514 479491 677517
rect 479076 677512 479491 677514
rect 479076 677456 479430 677512
rect 479486 677456 479491 677512
rect 479076 677454 479491 677456
rect 479076 677452 479082 677454
rect 479425 677451 479491 677454
rect 0 677318 6930 677378
rect 0 677288 800 677318
rect 481030 677242 481036 677244
rect 476968 677182 481036 677242
rect 481030 677180 481036 677182
rect 481100 677180 481106 677244
rect 479977 676970 480043 676973
rect 476968 676968 480043 676970
rect 476968 676912 479982 676968
rect 480038 676912 480043 676968
rect 476968 676910 480043 676912
rect 479977 676907 480043 676910
rect 485446 676834 485452 676836
rect 477358 676774 485452 676834
rect 477358 676766 477418 676774
rect 485446 676772 485452 676774
rect 485516 676772 485522 676836
rect 0 676698 800 676728
rect 476940 676706 477418 676766
rect 0 676638 10032 676698
rect 0 676608 800 676638
rect 483054 676562 483060 676564
rect 477358 676502 483060 676562
rect 477358 676494 477418 676502
rect 483054 676500 483060 676502
rect 483124 676500 483130 676564
rect 476940 676434 477418 676494
rect 483054 676228 483060 676292
rect 483124 676290 483130 676292
rect 484025 676290 484091 676293
rect 483124 676288 484091 676290
rect 483124 676232 484030 676288
rect 484086 676232 484091 676288
rect 483124 676230 484091 676232
rect 483124 676228 483130 676230
rect 484025 676227 484091 676230
rect 476968 676094 480270 676154
rect 0 676018 800 676048
rect 480210 676018 480270 676094
rect 480662 676092 480668 676156
rect 480732 676154 480738 676156
rect 481541 676154 481607 676157
rect 480732 676152 481607 676154
rect 480732 676096 481546 676152
rect 481602 676096 481607 676152
rect 480732 676094 481607 676096
rect 480732 676092 480738 676094
rect 481541 676091 481607 676094
rect 483606 676092 483612 676156
rect 483676 676154 483682 676156
rect 484209 676154 484275 676157
rect 483676 676152 484275 676154
rect 483676 676096 484214 676152
rect 484270 676096 484275 676152
rect 483676 676094 484275 676096
rect 483676 676092 483682 676094
rect 484209 676091 484275 676094
rect 482277 676018 482343 676021
rect 0 675958 9506 676018
rect 480210 676016 482343 676018
rect 480210 675960 482282 676016
rect 482338 675960 482343 676016
rect 480210 675958 482343 675960
rect 0 675928 800 675958
rect 9446 675950 9506 675958
rect 482277 675955 482343 675958
rect 9446 675890 10060 675950
rect 479374 675882 479380 675884
rect 476968 675822 479380 675882
rect 479374 675820 479380 675822
rect 479444 675820 479450 675884
rect 479558 675820 479564 675884
rect 479628 675882 479634 675884
rect 480161 675882 480227 675885
rect 479628 675880 480227 675882
rect 479628 675824 480166 675880
rect 480222 675824 480227 675880
rect 479628 675822 480227 675824
rect 479628 675820 479634 675822
rect 480161 675819 480227 675822
rect 482134 675610 482140 675612
rect 476968 675550 482140 675610
rect 482134 675548 482140 675550
rect 482204 675548 482210 675612
rect 483790 675474 483796 675476
rect 477358 675414 483796 675474
rect 477358 675406 477418 675414
rect 483790 675412 483796 675414
rect 483860 675412 483866 675476
rect 0 675338 800 675368
rect 476940 675346 477418 675406
rect 0 675278 9506 675338
rect 0 675248 800 675278
rect 9446 675134 9506 675278
rect 9446 675074 10060 675134
rect 481449 675066 481515 675069
rect 476968 675064 481515 675066
rect 476968 675008 481454 675064
rect 481510 675008 481515 675064
rect 476968 675006 481515 675008
rect 481449 675003 481515 675006
rect 479742 674794 479748 674796
rect 476968 674734 479748 674794
rect 479742 674732 479748 674734
rect 479812 674732 479818 674796
rect 483790 674732 483796 674796
rect 483860 674794 483866 674796
rect 484301 674794 484367 674797
rect 483860 674792 484367 674794
rect 483860 674736 484306 674792
rect 484362 674736 484367 674792
rect 483860 674734 484367 674736
rect 483860 674732 483866 674734
rect 484301 674731 484367 674734
rect 484526 674658 484532 674660
rect 477358 674598 484532 674658
rect 477358 674590 477418 674598
rect 484526 674596 484532 674598
rect 484596 674596 484602 674660
rect 476940 674530 477418 674590
rect 486366 674386 486372 674388
rect 477358 674326 486372 674386
rect 477358 674318 477418 674326
rect 486366 674324 486372 674326
rect 486436 674324 486442 674388
rect 476940 674258 477418 674318
rect 6870 674190 10032 674250
rect 0 673978 800 674008
rect 6870 673978 6930 674190
rect 483054 674114 483060 674116
rect 477358 674054 483060 674114
rect 477358 674046 477418 674054
rect 483054 674052 483060 674054
rect 483124 674052 483130 674116
rect 476940 673986 477418 674046
rect 0 673918 6930 673978
rect 0 673888 800 673918
rect 478454 673706 478460 673708
rect 476968 673646 478460 673706
rect 478454 673644 478460 673646
rect 478524 673644 478530 673708
rect 479190 673434 479196 673436
rect 6870 673374 10032 673434
rect 476968 673374 479196 673434
rect 0 673298 800 673328
rect 6870 673298 6930 673374
rect 479190 673372 479196 673374
rect 479260 673372 479266 673436
rect 0 673238 6930 673298
rect 0 673208 800 673238
rect 480662 673162 480668 673164
rect 476968 673102 480668 673162
rect 480662 673100 480668 673102
rect 480732 673100 480738 673164
rect 481950 672890 481956 672892
rect 476968 672830 481956 672890
rect 481950 672828 481956 672830
rect 482020 672828 482026 672892
rect 0 672618 800 672648
rect 480846 672618 480852 672620
rect 0 672558 10032 672618
rect 476968 672558 480852 672618
rect 0 672528 800 672558
rect 480846 672556 480852 672558
rect 480916 672556 480922 672620
rect 485630 672482 485636 672484
rect 477358 672422 485636 672482
rect 477358 672414 477418 672422
rect 485630 672420 485636 672422
rect 485700 672420 485706 672484
rect 476940 672354 477418 672414
rect 483606 672074 483612 672076
rect 476968 672014 483612 672074
rect 483606 672012 483612 672014
rect 483676 672012 483682 672076
rect 0 671938 800 671968
rect 483657 671938 483723 671941
rect 0 671878 9506 671938
rect 0 671848 800 671878
rect 9446 671870 9506 671878
rect 477358 671936 483723 671938
rect 477358 671880 483662 671936
rect 483718 671880 483723 671936
rect 477358 671878 483723 671880
rect 477358 671870 477418 671878
rect 483657 671875 483723 671878
rect 9446 671810 10060 671870
rect 476940 671810 477418 671870
rect 483238 671666 483244 671668
rect 477358 671606 483244 671666
rect 477358 671598 477418 671606
rect 483238 671604 483244 671606
rect 483308 671604 483314 671668
rect 476940 671538 477418 671598
rect 477125 671326 477191 671329
rect 476940 671324 477191 671326
rect 0 671258 800 671288
rect 476940 671268 477130 671324
rect 477186 671268 477191 671324
rect 476940 671266 477191 671268
rect 477125 671263 477191 671266
rect 0 671198 9506 671258
rect 0 671168 800 671198
rect 9446 671054 9506 671198
rect 9446 670994 10060 671054
rect 477718 670986 477724 670988
rect 476968 670926 477724 670986
rect 477718 670924 477724 670926
rect 477788 670924 477794 670988
rect 477217 670782 477283 670785
rect 476940 670780 477283 670782
rect 476940 670724 477222 670780
rect 477278 670724 477283 670780
rect 476940 670722 477283 670724
rect 477217 670719 477283 670722
rect 476902 670448 476908 670512
rect 476972 670448 476978 670512
rect 481582 670170 481588 670172
rect 6870 670110 10032 670170
rect 476968 670110 481588 670170
rect 0 669898 800 669928
rect 6870 669898 6930 670110
rect 481582 670108 481588 670110
rect 481652 670108 481658 670172
rect 479558 669898 479564 669900
rect 0 669838 6930 669898
rect 476968 669838 479564 669898
rect 0 669808 800 669838
rect 479558 669836 479564 669838
rect 479628 669836 479634 669900
rect 479006 669626 479012 669628
rect 476968 669566 479012 669626
rect 479006 669564 479012 669566
rect 479076 669564 479082 669628
rect 481766 669354 481772 669356
rect 6870 669294 10032 669354
rect 476968 669294 481772 669354
rect 0 669218 800 669248
rect 6870 669218 6930 669294
rect 481766 669292 481772 669294
rect 481836 669292 481842 669356
rect 483790 669218 483796 669220
rect 0 669158 6930 669218
rect 477358 669158 483796 669218
rect 0 669128 800 669158
rect 477358 669150 477418 669158
rect 483790 669156 483796 669158
rect 483860 669156 483866 669220
rect 476940 669090 477418 669150
rect 483422 668946 483428 668948
rect 477358 668886 483428 668946
rect 477358 668878 477418 668886
rect 483422 668884 483428 668886
rect 483492 668884 483498 668948
rect 476940 668818 477418 668878
rect 0 668538 800 668568
rect 0 668478 10032 668538
rect 0 668448 800 668478
rect 0 667858 800 667888
rect 0 667798 9506 667858
rect 0 667768 800 667798
rect 9446 667790 9506 667798
rect 9446 667730 10060 667790
rect 0 667178 800 667208
rect 0 667118 9506 667178
rect 0 667088 800 667118
rect 9446 666974 9506 667118
rect 9446 666914 10060 666974
rect 6870 666030 10032 666090
rect 0 665818 800 665848
rect 6870 665818 6930 666030
rect 0 665758 6930 665818
rect 0 665728 800 665758
rect 6870 665214 10032 665274
rect 0 665138 800 665168
rect 6870 665138 6930 665214
rect 0 665078 6930 665138
rect 0 665048 800 665078
rect 0 664458 800 664488
rect 0 664398 10032 664458
rect 0 664368 800 664398
rect 0 663778 800 663808
rect 0 663718 9506 663778
rect 0 663688 800 663718
rect 9446 663710 9506 663718
rect 9446 663650 10060 663710
rect 0 663098 800 663128
rect 0 663038 9506 663098
rect 0 663008 800 663038
rect 9446 662894 9506 663038
rect 9446 662834 10060 662894
rect 6870 661950 10032 662010
rect 0 661738 800 661768
rect 6870 661738 6930 661950
rect 0 661678 6930 661738
rect 0 661648 800 661678
rect 6870 661134 10032 661194
rect 0 661058 800 661088
rect 6870 661058 6930 661134
rect 0 660998 6930 661058
rect 0 660968 800 660998
rect 0 660378 800 660408
rect 0 660318 10032 660378
rect 0 660288 800 660318
rect 0 659698 800 659728
rect 0 659638 4170 659698
rect 0 659608 800 659638
rect 4110 659562 4170 659638
rect 4110 659502 10032 659562
rect 0 659018 800 659048
rect 0 658958 9506 659018
rect 0 658928 800 658958
rect 9446 658814 9506 658958
rect 9446 658754 10060 658814
rect 6870 657870 10032 657930
rect 0 657658 800 657688
rect 6870 657658 6930 657870
rect 0 657598 6930 657658
rect 0 657568 800 657598
rect 6870 657054 10032 657114
rect 0 656978 800 657008
rect 6870 656978 6930 657054
rect 0 656918 6930 656978
rect 0 656888 800 656918
rect 0 656298 800 656328
rect 0 656238 10032 656298
rect 0 656208 800 656238
rect 0 655618 800 655648
rect 0 655558 4170 655618
rect 0 655528 800 655558
rect 4110 655482 4170 655558
rect 4110 655422 10032 655482
rect 0 654938 800 654968
rect 0 654878 9506 654938
rect 0 654848 800 654878
rect 9446 654734 9506 654878
rect 9446 654674 10060 654734
rect 6870 653790 10032 653850
rect 0 653578 800 653608
rect 6870 653578 6930 653790
rect 0 653518 6930 653578
rect 0 653488 800 653518
rect 6870 652974 10032 653034
rect 0 652898 800 652928
rect 6870 652898 6930 652974
rect 0 652838 6930 652898
rect 0 652808 800 652838
rect 0 652218 800 652248
rect 0 652158 10032 652218
rect 0 652128 800 652158
rect 0 651538 800 651568
rect 0 651478 9506 651538
rect 0 651448 800 651478
rect 9446 651470 9506 651478
rect 9446 651410 10060 651470
rect 0 643378 800 643408
rect 0 643318 4170 643378
rect 0 643288 800 643318
rect 4110 643106 4170 643318
rect 4110 643046 10038 643106
rect 6870 642230 10038 642290
rect 0 642018 800 642048
rect 6870 642018 6930 642230
rect 0 641958 6930 642018
rect 0 641928 800 641958
rect 6870 641414 10038 641474
rect 0 641338 800 641368
rect 6870 641338 6930 641414
rect 0 641278 6930 641338
rect 0 641248 800 641278
rect 0 640658 800 640688
rect 0 640598 10038 640658
rect 0 640568 800 640598
rect 0 639978 800 640008
rect 0 639918 9506 639978
rect 0 639888 800 639918
rect 9446 639912 9506 639918
rect 9446 639852 10060 639912
rect 0 639298 800 639328
rect 0 639238 9506 639298
rect 0 639208 800 639238
rect 9446 639096 9506 639238
rect 9446 639036 10060 639096
rect 6870 638150 10038 638210
rect 0 637938 800 637968
rect 6870 637938 6930 638150
rect 0 637878 6930 637938
rect 0 637848 800 637878
rect 6870 637334 10038 637394
rect 0 637258 800 637288
rect 6870 637258 6930 637334
rect 0 637198 6930 637258
rect 0 637168 800 637198
rect 0 636578 800 636608
rect 0 636518 10038 636578
rect 0 636488 800 636518
rect 0 635898 800 635928
rect 0 635838 9506 635898
rect 0 635808 800 635838
rect 9446 635832 9506 635838
rect 9446 635772 10060 635832
rect 0 635218 800 635248
rect 0 635158 9506 635218
rect 0 635128 800 635158
rect 9446 635016 9506 635158
rect 9446 634956 10060 635016
rect 6870 634070 10038 634130
rect 0 633858 800 633888
rect 6870 633858 6930 634070
rect 0 633798 6930 633858
rect 0 633768 800 633798
rect 6870 633254 10038 633314
rect 0 633178 800 633208
rect 6870 633178 6930 633254
rect 0 633118 6930 633178
rect 0 633088 800 633118
rect 0 632498 800 632528
rect 0 632438 10038 632498
rect 0 632408 800 632438
rect 0 631818 800 631848
rect 0 631758 9506 631818
rect 0 631728 800 631758
rect 9446 631752 9506 631758
rect 9446 631692 10060 631752
rect 0 631138 800 631168
rect 0 631078 9506 631138
rect 0 631048 800 631078
rect 9446 630936 9506 631078
rect 9446 630876 10060 630936
rect 481541 630458 481607 630461
rect 486200 630458 487000 630488
rect 481541 630456 487000 630458
rect 481541 630400 481546 630456
rect 481602 630400 487000 630456
rect 481541 630398 487000 630400
rect 481541 630395 481607 630398
rect 486200 630368 487000 630398
rect 6870 629990 10038 630050
rect 0 629778 800 629808
rect 6870 629778 6930 629990
rect 0 629718 6930 629778
rect 482921 629778 482987 629781
rect 486200 629778 487000 629808
rect 482921 629776 487000 629778
rect 482921 629720 482926 629776
rect 482982 629720 487000 629776
rect 482921 629718 487000 629720
rect 0 629688 800 629718
rect 482921 629715 482987 629718
rect 486200 629688 487000 629718
rect 6870 629174 10038 629234
rect 0 629098 800 629128
rect 6870 629098 6930 629174
rect 0 629038 6930 629098
rect 484301 629098 484367 629101
rect 486200 629098 487000 629128
rect 484301 629096 487000 629098
rect 484301 629040 484306 629096
rect 484362 629040 487000 629096
rect 484301 629038 487000 629040
rect 0 629008 800 629038
rect 484301 629035 484367 629038
rect 486200 629008 487000 629038
rect 0 628418 800 628448
rect 481449 628418 481515 628421
rect 486200 628418 487000 628448
rect 0 628358 10038 628418
rect 481449 628416 487000 628418
rect 481449 628360 481454 628416
rect 481510 628360 487000 628416
rect 481449 628358 487000 628360
rect 0 628328 800 628358
rect 481449 628355 481515 628358
rect 486200 628328 487000 628358
rect 0 627738 800 627768
rect 482829 627738 482895 627741
rect 486200 627738 487000 627768
rect 0 627678 9506 627738
rect 0 627648 800 627678
rect 9446 627672 9506 627678
rect 482829 627736 487000 627738
rect 482829 627680 482834 627736
rect 482890 627680 487000 627736
rect 482829 627678 487000 627680
rect 482829 627675 482895 627678
rect 9446 627612 10060 627672
rect 486200 627648 487000 627678
rect 0 627058 800 627088
rect 484209 627058 484275 627061
rect 486200 627058 487000 627088
rect 0 626998 9506 627058
rect 0 626968 800 626998
rect 9446 626856 9506 626998
rect 484209 627056 487000 627058
rect 484209 627000 484214 627056
rect 484270 627000 487000 627056
rect 484209 626998 487000 627000
rect 484209 626995 484275 626998
rect 486200 626968 487000 626998
rect 9446 626796 10060 626856
rect 482134 626316 482140 626380
rect 482204 626378 482210 626380
rect 486200 626378 487000 626408
rect 482204 626318 487000 626378
rect 482204 626316 482210 626318
rect 486200 626288 487000 626318
rect 6870 625910 10038 625970
rect 0 625698 800 625728
rect 6870 625698 6930 625910
rect 0 625638 6930 625698
rect 0 625608 800 625638
rect 480846 625636 480852 625700
rect 480916 625698 480922 625700
rect 486200 625698 487000 625728
rect 480916 625638 487000 625698
rect 480916 625636 480922 625638
rect 486200 625608 487000 625638
rect 6870 625094 10038 625154
rect 0 625018 800 625048
rect 6870 625018 6930 625094
rect 0 624958 6930 625018
rect 478781 625018 478847 625021
rect 486200 625018 487000 625048
rect 478781 625016 487000 625018
rect 478781 624960 478786 625016
rect 478842 624960 487000 625016
rect 478781 624958 487000 624960
rect 0 624928 800 624958
rect 478781 624955 478847 624958
rect 486200 624928 487000 624958
rect 0 624338 800 624368
rect 478689 624338 478755 624341
rect 486200 624338 487000 624368
rect 0 624278 10038 624338
rect 478689 624336 487000 624338
rect 478689 624280 478694 624336
rect 478750 624280 487000 624336
rect 478689 624278 487000 624280
rect 0 624248 800 624278
rect 478689 624275 478755 624278
rect 486200 624248 487000 624278
rect 0 623658 800 623688
rect 0 623598 9506 623658
rect 0 623568 800 623598
rect 9446 623592 9506 623598
rect 478086 623596 478092 623660
rect 478156 623658 478162 623660
rect 486200 623658 487000 623688
rect 478156 623598 487000 623658
rect 478156 623596 478162 623598
rect 9446 623532 10060 623592
rect 486200 623568 487000 623598
rect 0 622978 800 623008
rect 0 622918 9506 622978
rect 0 622888 800 622918
rect 9446 622776 9506 622918
rect 478270 622916 478276 622980
rect 478340 622978 478346 622980
rect 486200 622978 487000 623008
rect 478340 622918 487000 622978
rect 478340 622916 478346 622918
rect 486200 622888 487000 622918
rect 9446 622716 10060 622776
rect 483606 622236 483612 622300
rect 483676 622298 483682 622300
rect 486200 622298 487000 622328
rect 483676 622238 487000 622298
rect 483676 622236 483682 622238
rect 486200 622208 487000 622238
rect 6870 621830 10038 621890
rect 0 621618 800 621648
rect 6870 621618 6930 621830
rect 0 621558 6930 621618
rect 0 621528 800 621558
rect 478454 621556 478460 621620
rect 478524 621618 478530 621620
rect 486200 621618 487000 621648
rect 478524 621558 487000 621618
rect 478524 621556 478530 621558
rect 486200 621528 487000 621558
rect 6870 621014 10038 621074
rect 0 620938 800 620968
rect 6870 620938 6930 621014
rect 0 620878 6930 620938
rect 0 620848 800 620878
rect 479374 620876 479380 620940
rect 479444 620938 479450 620940
rect 486200 620938 487000 620968
rect 479444 620878 487000 620938
rect 479444 620876 479450 620878
rect 486200 620848 487000 620878
rect 0 620258 800 620288
rect 482277 620258 482343 620261
rect 486200 620258 487000 620288
rect 0 620198 10038 620258
rect 482277 620256 487000 620258
rect 482277 620200 482282 620256
rect 482338 620200 487000 620256
rect 482277 620198 487000 620200
rect 0 620168 800 620198
rect 482277 620195 482343 620198
rect 486200 620168 487000 620198
rect 0 619578 800 619608
rect 0 619518 9506 619578
rect 0 619488 800 619518
rect 9446 619512 9506 619518
rect 485814 619516 485820 619580
rect 485884 619578 485890 619580
rect 486200 619578 487000 619608
rect 485884 619518 487000 619578
rect 485884 619516 485890 619518
rect 9446 619452 10060 619512
rect 486200 619488 487000 619518
rect 0 618898 800 618928
rect 0 618838 9506 618898
rect 0 618808 800 618838
rect 9446 618696 9506 618838
rect 483790 618836 483796 618900
rect 483860 618898 483866 618900
rect 486200 618898 487000 618928
rect 483860 618838 487000 618898
rect 483860 618836 483866 618838
rect 486200 618808 487000 618838
rect 9446 618636 10060 618696
rect 479558 618156 479564 618220
rect 479628 618218 479634 618220
rect 486200 618218 487000 618248
rect 479628 618158 487000 618218
rect 479628 618156 479634 618158
rect 486200 618128 487000 618158
rect 6870 617750 10038 617810
rect 0 617538 800 617568
rect 6870 617538 6930 617750
rect 0 617478 6930 617538
rect 0 617448 800 617478
rect 481030 617476 481036 617540
rect 481100 617538 481106 617540
rect 486200 617538 487000 617568
rect 481100 617478 487000 617538
rect 481100 617476 481106 617478
rect 486200 617448 487000 617478
rect 6870 616934 10038 616994
rect 0 616858 800 616888
rect 6870 616858 6930 616934
rect 0 616798 6930 616858
rect 483657 616858 483723 616861
rect 486200 616858 487000 616888
rect 483657 616856 487000 616858
rect 483657 616800 483662 616856
rect 483718 616800 487000 616856
rect 483657 616798 487000 616800
rect 0 616768 800 616798
rect 483657 616795 483723 616798
rect 486200 616768 487000 616798
rect 0 616178 800 616208
rect 0 616118 10038 616178
rect 0 616088 800 616118
rect 479926 616116 479932 616180
rect 479996 616178 480002 616180
rect 486200 616178 487000 616208
rect 479996 616118 487000 616178
rect 479996 616116 480002 616118
rect 486200 616088 487000 616118
rect 0 615498 800 615528
rect 0 615438 9506 615498
rect 0 615408 800 615438
rect 9446 615432 9506 615438
rect 485262 615436 485268 615500
rect 485332 615498 485338 615500
rect 486200 615498 487000 615528
rect 485332 615438 487000 615498
rect 485332 615436 485338 615438
rect 9446 615372 10060 615432
rect 486200 615408 487000 615438
rect 0 614818 800 614848
rect 0 614758 9506 614818
rect 0 614728 800 614758
rect 9446 614616 9506 614758
rect 485998 614756 486004 614820
rect 486068 614818 486074 614820
rect 486200 614818 487000 614848
rect 486068 614758 487000 614818
rect 486068 614756 486074 614758
rect 486200 614728 487000 614758
rect 9446 614556 10060 614616
rect 481214 614076 481220 614140
rect 481284 614138 481290 614140
rect 486200 614138 487000 614168
rect 481284 614078 487000 614138
rect 481284 614076 481290 614078
rect 486200 614048 487000 614078
rect 6870 613670 10038 613730
rect 0 613458 800 613488
rect 6870 613458 6930 613670
rect 0 613398 6930 613458
rect 0 613368 800 613398
rect 478638 613396 478644 613460
rect 478708 613458 478714 613460
rect 486200 613458 487000 613488
rect 478708 613398 487000 613458
rect 478708 613396 478714 613398
rect 486200 613368 487000 613398
rect 6870 612854 10038 612914
rect 0 612778 800 612808
rect 6870 612778 6930 612854
rect 0 612718 6930 612778
rect 0 612688 800 612718
rect 482870 612716 482876 612780
rect 482940 612778 482946 612780
rect 486200 612778 487000 612808
rect 482940 612718 487000 612778
rect 482940 612716 482946 612718
rect 486200 612688 487000 612718
rect 0 612098 800 612128
rect 0 612038 10038 612098
rect 0 612008 800 612038
rect 479742 612036 479748 612100
rect 479812 612098 479818 612100
rect 486200 612098 487000 612128
rect 479812 612038 487000 612098
rect 479812 612036 479818 612038
rect 486200 612008 487000 612038
rect 0 611418 800 611448
rect 0 611358 4170 611418
rect 0 611328 800 611358
rect 4110 611282 4170 611358
rect 482686 611356 482692 611420
rect 482756 611418 482762 611420
rect 486200 611418 487000 611448
rect 482756 611358 487000 611418
rect 482756 611356 482762 611358
rect 486200 611328 487000 611358
rect 4110 611222 10038 611282
rect 0 610738 800 610768
rect 0 610678 9506 610738
rect 0 610648 800 610678
rect 9446 610536 9506 610678
rect 483422 610676 483428 610740
rect 483492 610738 483498 610740
rect 486200 610738 487000 610768
rect 483492 610678 487000 610738
rect 483492 610676 483498 610678
rect 486200 610648 487000 610678
rect 9446 610476 10060 610536
rect 477350 609996 477356 610060
rect 477420 610058 477426 610060
rect 486200 610058 487000 610088
rect 477420 609998 487000 610058
rect 477420 609996 477426 609998
rect 486200 609968 487000 609998
rect 6870 609590 10038 609650
rect 0 609378 800 609408
rect 6870 609378 6930 609590
rect 0 609318 6930 609378
rect 486200 609380 487000 609408
rect 0 609288 800 609318
rect 486200 609316 486372 609380
rect 486436 609316 487000 609380
rect 486200 609288 487000 609316
rect 6870 608774 10038 608834
rect 0 608698 800 608728
rect 6870 608698 6930 608774
rect 0 608638 6930 608698
rect 0 608608 800 608638
rect 485630 608636 485636 608700
rect 485700 608698 485706 608700
rect 486200 608698 487000 608728
rect 485700 608638 487000 608698
rect 485700 608636 485706 608638
rect 486200 608608 487000 608638
rect 482870 608154 482876 608156
rect 476940 608094 482876 608154
rect 482870 608092 482876 608094
rect 482940 608092 482946 608156
rect 0 608018 800 608048
rect 0 607958 10038 608018
rect 0 607928 800 607958
rect 484710 607956 484716 608020
rect 484780 608018 484786 608020
rect 486200 608018 487000 608048
rect 484780 607958 487000 608018
rect 484780 607956 484786 607958
rect 486200 607928 487000 607958
rect 479926 607882 479932 607884
rect 476940 607822 479932 607882
rect 479926 607820 479932 607822
rect 479996 607820 480002 607884
rect 486366 607746 486372 607748
rect 477358 607696 486372 607746
rect 476928 607686 486372 607696
rect 476928 607636 477418 607686
rect 486366 607684 486372 607686
rect 486436 607684 486442 607748
rect 477350 607424 477356 607426
rect 0 607338 800 607368
rect 476928 607364 477356 607424
rect 477350 607362 477356 607364
rect 477420 607362 477426 607426
rect 0 607278 4170 607338
rect 0 607248 800 607278
rect 4110 607202 4170 607278
rect 481766 607276 481772 607340
rect 481836 607338 481842 607340
rect 486200 607338 487000 607368
rect 481836 607278 487000 607338
rect 481836 607276 481842 607278
rect 486200 607248 487000 607278
rect 4110 607142 10038 607202
rect 481582 607140 481588 607204
rect 481652 607202 481658 607204
rect 482829 607202 482895 607205
rect 481652 607200 482895 607202
rect 481652 607144 482834 607200
rect 482890 607144 482895 607200
rect 481652 607142 482895 607144
rect 481652 607140 481658 607142
rect 482829 607139 482895 607142
rect 483238 607140 483244 607204
rect 483308 607202 483314 607204
rect 484209 607202 484275 607205
rect 483308 607200 484275 607202
rect 483308 607144 484214 607200
rect 484270 607144 484275 607200
rect 483308 607142 484275 607144
rect 483308 607140 483314 607142
rect 484209 607139 484275 607142
rect 482277 607066 482343 607069
rect 476940 607064 482343 607066
rect 476940 607008 482282 607064
rect 482338 607008 482343 607064
rect 476940 607006 482343 607008
rect 482277 607003 482343 607006
rect 483054 607004 483060 607068
rect 483124 607066 483130 607068
rect 484301 607066 484367 607069
rect 483124 607064 484367 607066
rect 483124 607008 484306 607064
rect 484362 607008 484367 607064
rect 483124 607006 484367 607008
rect 483124 607004 483130 607006
rect 484301 607003 484367 607006
rect 483422 606930 483428 606932
rect 477358 606880 483428 606930
rect 476928 606870 483428 606880
rect 476928 606820 477418 606870
rect 483422 606868 483428 606870
rect 483492 606868 483498 606932
rect 0 606658 800 606688
rect 486200 606658 487000 606688
rect 0 606598 9506 606658
rect 477358 606608 487000 606658
rect 0 606568 800 606598
rect 9446 606454 9506 606598
rect 476928 606598 487000 606608
rect 476928 606548 477418 606598
rect 486200 606568 487000 606598
rect 9446 606394 10032 606454
rect 482686 606250 482692 606252
rect 476940 606190 482692 606250
rect 482686 606188 482692 606190
rect 482756 606188 482762 606252
rect 479558 605978 479564 605980
rect 476940 605918 479564 605978
rect 479558 605916 479564 605918
rect 479628 605916 479634 605980
rect 484894 605916 484900 605980
rect 484964 605978 484970 605980
rect 486200 605978 487000 606008
rect 484964 605918 487000 605978
rect 484964 605916 484970 605918
rect 486200 605888 487000 605918
rect 481766 605706 481772 605708
rect 476940 605646 481772 605706
rect 481766 605644 481772 605646
rect 481836 605644 481842 605708
rect 483790 605570 483796 605572
rect 477358 605520 483796 605570
rect 476928 605510 483796 605520
rect 476928 605460 477418 605510
rect 483790 605508 483796 605510
rect 483860 605508 483866 605572
rect 486200 605298 487000 605328
rect 477358 605248 487000 605298
rect 476928 605238 487000 605248
rect 476928 605188 477418 605238
rect 486200 605208 487000 605238
rect 478638 604890 478644 604892
rect 476940 604830 478644 604890
rect 478638 604828 478644 604830
rect 478708 604828 478714 604892
rect 481214 604618 481220 604620
rect 476940 604558 481220 604618
rect 481214 604556 481220 604558
rect 481284 604556 481290 604620
rect 484526 604556 484532 604620
rect 484596 604618 484602 604620
rect 486200 604618 487000 604648
rect 484596 604558 487000 604618
rect 484596 604556 484602 604558
rect 486200 604528 487000 604558
rect 480294 604420 480300 604484
rect 480364 604482 480370 604484
rect 481449 604482 481515 604485
rect 480364 604480 481515 604482
rect 480364 604424 481454 604480
rect 481510 604424 481515 604480
rect 480364 604422 481515 604424
rect 480364 604420 480370 604422
rect 481449 604419 481515 604422
rect 484710 604346 484716 604348
rect 476940 604286 484716 604346
rect 484710 604284 484716 604286
rect 484780 604284 484786 604348
rect 485998 604210 486004 604212
rect 477358 604160 486004 604210
rect 476928 604150 486004 604160
rect 476928 604100 477418 604150
rect 485998 604148 486004 604150
rect 486068 604148 486074 604212
rect 486200 603938 487000 603968
rect 477358 603888 487000 603938
rect 476928 603878 487000 603888
rect 476928 603828 477418 603878
rect 486200 603848 487000 603878
rect 485262 603666 485268 603668
rect 477358 603616 485268 603666
rect 476928 603606 485268 603616
rect 476928 603556 477418 603606
rect 485262 603604 485268 603606
rect 485332 603604 485338 603668
rect 485814 603394 485820 603396
rect 477358 603344 485820 603394
rect 476928 603334 485820 603344
rect 476928 603284 477418 603334
rect 485814 603332 485820 603334
rect 485884 603332 485890 603396
rect 484342 603196 484348 603260
rect 484412 603258 484418 603260
rect 486200 603258 487000 603288
rect 484412 603198 487000 603258
rect 484412 603196 484418 603198
rect 486200 603168 487000 603198
rect 480478 603060 480484 603124
rect 480548 603122 480554 603124
rect 481541 603122 481607 603125
rect 480548 603120 481607 603122
rect 480548 603064 481546 603120
rect 481602 603064 481607 603120
rect 480548 603062 481607 603064
rect 480548 603060 480554 603062
rect 481541 603059 481607 603062
rect 484526 602986 484532 602988
rect 476940 602926 484532 602986
rect 484526 602924 484532 602926
rect 484596 602924 484602 602988
rect 483657 602850 483723 602853
rect 477358 602848 483723 602850
rect 477358 602800 483662 602848
rect 476928 602792 483662 602800
rect 483718 602792 483723 602848
rect 476928 602790 483723 602792
rect 476928 602740 477418 602790
rect 483657 602787 483723 602790
rect 481398 602516 481404 602580
rect 481468 602578 481474 602580
rect 486200 602578 487000 602608
rect 481468 602518 487000 602578
rect 481468 602516 481474 602518
rect 486200 602488 487000 602518
rect 479742 602442 479748 602444
rect 476940 602382 479748 602442
rect 479742 602380 479748 602382
rect 479812 602380 479818 602444
rect 481030 602170 481036 602172
rect 476940 602110 481036 602170
rect 481030 602108 481036 602110
rect 481100 602108 481106 602172
rect 479374 601898 479380 601900
rect 476940 601838 479380 601898
rect 479374 601836 479380 601838
rect 479444 601836 479450 601900
rect 483422 601836 483428 601900
rect 483492 601898 483498 601900
rect 486200 601898 487000 601928
rect 483492 601838 487000 601898
rect 483492 601836 483498 601838
rect 486200 601808 487000 601838
rect 477718 601700 477724 601764
rect 477788 601762 477794 601764
rect 478689 601762 478755 601765
rect 477788 601760 478755 601762
rect 477788 601704 478694 601760
rect 478750 601704 478755 601760
rect 477788 601702 478755 601704
rect 477788 601700 477794 601702
rect 478689 601699 478755 601702
rect 481766 601700 481772 601764
rect 481836 601762 481842 601764
rect 482921 601762 482987 601765
rect 481836 601760 482987 601762
rect 481836 601704 482926 601760
rect 482982 601704 482987 601760
rect 481836 601702 482987 601704
rect 481836 601700 481842 601702
rect 482921 601699 482987 601702
rect 484894 601626 484900 601628
rect 476940 601566 484900 601626
rect 484894 601564 484900 601566
rect 484964 601564 484970 601628
rect 484342 601490 484348 601492
rect 477358 601440 484348 601490
rect 476928 601430 484348 601440
rect 476928 601380 477418 601430
rect 484342 601428 484348 601430
rect 484412 601428 484418 601492
rect 483422 601354 483428 601356
rect 483062 601294 483428 601354
rect 481398 601082 481404 601084
rect 476940 601022 481404 601082
rect 481398 601020 481404 601022
rect 481468 601020 481474 601084
rect 483062 600946 483122 601294
rect 483422 601292 483428 601294
rect 483492 601292 483498 601356
rect 486200 601218 487000 601248
rect 477358 600896 483122 600946
rect 476928 600886 483122 600896
rect 483246 601158 487000 601218
rect 476928 600836 477418 600886
rect 483246 600674 483306 601158
rect 486200 601128 487000 601158
rect 477358 600624 483306 600674
rect 476928 600614 483306 600624
rect 476928 600564 477418 600614
rect 483422 600476 483428 600540
rect 483492 600538 483498 600540
rect 486200 600538 487000 600568
rect 483492 600478 487000 600538
rect 483492 600476 483498 600478
rect 486200 600448 487000 600478
rect 485630 600266 485636 600268
rect 476940 600206 485636 600266
rect 485630 600204 485636 600206
rect 485700 600204 485706 600268
rect 483422 600130 483428 600132
rect 477358 600080 483428 600130
rect 476928 600070 483428 600080
rect 476928 600020 477418 600070
rect 483422 600068 483428 600070
rect 483492 600068 483498 600132
rect 486200 599858 487000 599888
rect 477358 599808 487000 599858
rect 476928 599798 487000 599808
rect 476928 599748 477418 599798
rect 486200 599768 487000 599798
rect 478454 599450 478460 599452
rect 476940 599390 478460 599450
rect 478454 599388 478460 599390
rect 478524 599388 478530 599452
rect 483606 599314 483612 599316
rect 477358 599264 483612 599314
rect 476928 599254 483612 599264
rect 476928 599204 477418 599254
rect 483606 599252 483612 599254
rect 483676 599252 483682 599316
rect 477902 599116 477908 599180
rect 477972 599178 477978 599180
rect 478781 599178 478847 599181
rect 486200 599178 487000 599208
rect 477972 599176 478847 599178
rect 477972 599120 478786 599176
rect 478842 599120 478847 599176
rect 477972 599118 478847 599120
rect 477972 599116 477978 599118
rect 478781 599115 478847 599118
rect 484534 599118 487000 599178
rect 484534 598906 484594 599118
rect 486200 599088 487000 599118
rect 476940 598846 484594 598906
rect 478270 598634 478276 598636
rect 476940 598574 478276 598634
rect 478270 598572 478276 598574
rect 478340 598572 478346 598636
rect 486200 598498 487000 598528
rect 477358 598448 487000 598498
rect 476928 598438 487000 598448
rect 476928 598388 477418 598438
rect 486200 598408 487000 598438
rect 9446 598060 10060 598120
rect 478086 598090 478092 598092
rect 0 597818 800 597848
rect 9446 597818 9506 598060
rect 476940 598030 478092 598090
rect 478086 598028 478092 598030
rect 478156 598028 478162 598092
rect 477718 597818 477724 597820
rect 0 597758 9506 597818
rect 476940 597758 477724 597818
rect 0 597728 800 597758
rect 477718 597756 477724 597758
rect 477788 597756 477794 597820
rect 486200 597818 487000 597848
rect 481774 597758 487000 597818
rect 481774 597546 481834 597758
rect 486200 597728 487000 597758
rect 476940 597486 481834 597546
rect 9446 597244 10060 597304
rect 477902 597274 477908 597276
rect 0 597138 800 597168
rect 9446 597138 9506 597244
rect 476940 597214 477908 597274
rect 477902 597212 477908 597214
rect 477972 597212 477978 597276
rect 486200 597138 487000 597168
rect 0 597078 9506 597138
rect 477358 597088 487000 597138
rect 476928 597078 487000 597088
rect 0 597048 800 597078
rect 476928 597028 477418 597078
rect 486200 597048 487000 597078
rect 480846 596730 480852 596732
rect 476940 596670 480852 596730
rect 480846 596668 480852 596670
rect 480916 596668 480922 596732
rect 0 596458 800 596488
rect 9446 596458 10060 596488
rect 482134 596458 482140 596460
rect 0 596428 10060 596458
rect 0 596398 9506 596428
rect 476940 596398 482140 596458
rect 0 596368 800 596398
rect 482134 596396 482140 596398
rect 482204 596396 482210 596460
rect 486200 596458 487000 596488
rect 484718 596398 487000 596458
rect 484718 596186 484778 596398
rect 486200 596368 487000 596398
rect 476940 596126 484778 596186
rect 483238 596050 483244 596052
rect 477358 596000 483244 596050
rect 476928 595990 483244 596000
rect 476928 595940 477418 595990
rect 483238 595988 483244 595990
rect 483308 595988 483314 596052
rect 0 595778 800 595808
rect 486200 595778 487000 595808
rect 0 595728 9506 595778
rect 477358 595728 487000 595778
rect 0 595718 10060 595728
rect 0 595688 800 595718
rect 9446 595668 10060 595718
rect 476928 595718 487000 595728
rect 476928 595668 477418 595718
rect 486200 595688 487000 595718
rect 481582 595370 481588 595372
rect 476940 595310 481588 595370
rect 481582 595308 481588 595310
rect 481652 595308 481658 595372
rect 0 595098 800 595128
rect 480294 595098 480300 595100
rect 0 595038 9506 595098
rect 476940 595038 480300 595098
rect 0 595008 800 595038
rect 9446 594912 9506 595038
rect 480294 595036 480300 595038
rect 480364 595036 480370 595100
rect 486200 595098 487000 595128
rect 483246 595038 487000 595098
rect 483246 594962 483306 595038
rect 486200 595008 487000 595038
rect 477358 594912 483306 594962
rect 9446 594852 10060 594912
rect 476928 594902 483306 594912
rect 476928 594852 477418 594902
rect 483054 594690 483060 594692
rect 477358 594640 483060 594690
rect 476928 594630 483060 594640
rect 476928 594580 477418 594630
rect 483054 594628 483060 594630
rect 483124 594628 483130 594692
rect 486200 594418 487000 594448
rect 477358 594368 487000 594418
rect 476928 594358 487000 594368
rect 476928 594308 477418 594358
rect 486200 594328 487000 594358
rect 9446 593980 10060 594040
rect 481766 594010 481772 594012
rect 0 593738 800 593768
rect 9446 593738 9506 593980
rect 476940 593950 481772 594010
rect 481766 593948 481772 593950
rect 481836 593948 481842 594012
rect 480478 593738 480484 593740
rect 0 593678 9506 593738
rect 476940 593678 480484 593738
rect 0 593648 800 593678
rect 480478 593676 480484 593678
rect 480548 593676 480554 593740
rect 486200 593738 487000 593768
rect 483246 593678 487000 593738
rect 483246 593602 483306 593678
rect 486200 593648 487000 593678
rect 477358 593552 483306 593602
rect 476928 593542 483306 593552
rect 476928 593492 477418 593542
rect 477358 593280 483306 593330
rect 476928 593270 483306 593280
rect 9446 593164 10060 593224
rect 476928 593220 477418 593270
rect 0 593058 800 593088
rect 9446 593058 9506 593164
rect 483054 593058 483060 593060
rect 0 592998 9506 593058
rect 477358 593008 483060 593058
rect 476928 592998 483060 593008
rect 0 592968 800 592998
rect 476928 592948 477418 592998
rect 483054 592996 483060 592998
rect 483124 592996 483130 593060
rect 483246 593058 483306 593270
rect 486200 593058 487000 593088
rect 483246 592998 487000 593058
rect 486200 592968 487000 592998
rect 480662 592650 480668 592652
rect 476940 592590 480668 592650
rect 480662 592588 480668 592590
rect 480732 592588 480738 592652
rect 0 592378 800 592408
rect 9446 592378 10060 592408
rect 486200 592378 487000 592408
rect 0 592348 10060 592378
rect 0 592318 9506 592348
rect 476940 592318 487000 592378
rect 0 592288 800 592318
rect 486200 592288 487000 592318
rect 483606 592242 483612 592244
rect 477358 592192 483612 592242
rect 476928 592182 483612 592192
rect 476928 592132 477418 592182
rect 483606 592180 483612 592182
rect 483676 592180 483682 592244
rect 476940 591774 480270 591834
rect 0 591698 800 591728
rect 480210 591698 480270 591774
rect 486200 591698 487000 591728
rect 0 591648 9506 591698
rect 0 591638 10060 591648
rect 480210 591638 487000 591698
rect 0 591608 800 591638
rect 9446 591588 10060 591638
rect 486200 591608 487000 591638
rect 481766 591562 481772 591564
rect 476940 591502 481772 591562
rect 481766 591500 481772 591502
rect 481836 591500 481842 591564
rect 483790 591426 483796 591428
rect 477358 591376 483796 591426
rect 476928 591366 483796 591376
rect 476928 591316 477418 591366
rect 483790 591364 483796 591366
rect 483860 591364 483866 591428
rect 0 591018 800 591048
rect 486200 591018 487000 591048
rect 0 590958 9506 591018
rect 476940 590958 487000 591018
rect 0 590928 800 590958
rect 9446 590832 9506 590958
rect 486200 590928 487000 590958
rect 9446 590772 10060 590832
rect 481582 590746 481588 590748
rect 476940 590686 481588 590746
rect 481582 590684 481588 590686
rect 481652 590684 481658 590748
rect 476940 590414 480270 590474
rect 480210 590338 480270 590414
rect 486200 590338 487000 590368
rect 480210 590278 487000 590338
rect 486200 590248 487000 590278
rect 480294 590202 480300 590204
rect 476940 590142 480300 590202
rect 480294 590140 480300 590142
rect 480364 590140 480370 590204
rect 9446 589900 10060 589960
rect 482134 589930 482140 589932
rect 0 589658 800 589688
rect 9446 589658 9506 589900
rect 476940 589870 482140 589930
rect 482134 589868 482140 589870
rect 482204 589868 482210 589932
rect 486200 589658 487000 589688
rect 0 589598 9506 589658
rect 476940 589598 487000 589658
rect 0 589568 800 589598
rect 486200 589568 487000 589598
rect 483974 589522 483980 589524
rect 477358 589472 483980 589522
rect 476928 589462 483980 589472
rect 476928 589412 477418 589462
rect 483974 589460 483980 589462
rect 484044 589460 484050 589524
rect 9446 589084 10060 589144
rect 0 588978 800 589008
rect 9446 588978 9506 589084
rect 476940 589054 480270 589114
rect 0 588918 9506 588978
rect 480210 588978 480270 589054
rect 486200 588978 487000 589008
rect 480210 588918 487000 588978
rect 0 588888 800 588918
rect 486200 588888 487000 588918
rect 480846 588842 480852 588844
rect 476940 588782 480852 588842
rect 480846 588780 480852 588782
rect 480916 588780 480922 588844
rect 482318 588570 482324 588572
rect 476940 588510 482324 588570
rect 482318 588508 482324 588510
rect 482388 588508 482394 588572
rect 0 588298 800 588328
rect 9446 588298 10060 588328
rect 486200 588298 487000 588328
rect 0 588268 10060 588298
rect 0 588238 9506 588268
rect 476940 588238 487000 588298
rect 0 588208 800 588238
rect 486200 588208 487000 588238
rect 481030 588026 481036 588028
rect 476940 587966 481036 588026
rect 481030 587964 481036 587966
rect 481100 587964 481106 588028
rect 480662 587828 480668 587892
rect 480732 587890 480738 587892
rect 481541 587890 481607 587893
rect 480732 587888 481607 587890
rect 480732 587832 481546 587888
rect 481602 587832 481607 587888
rect 480732 587830 481607 587832
rect 480732 587828 480738 587830
rect 481541 587827 481607 587830
rect 476940 587694 480270 587754
rect 0 587618 800 587648
rect 480210 587618 480270 587694
rect 486200 587618 487000 587648
rect 0 587568 9506 587618
rect 0 587558 10060 587568
rect 480210 587558 487000 587618
rect 0 587528 800 587558
rect 9446 587508 10060 587558
rect 486200 587528 487000 587558
rect 481214 587482 481220 587484
rect 476940 587422 481220 587482
rect 481214 587420 481220 587422
rect 481284 587420 481290 587484
rect 480161 587210 480227 587213
rect 476940 587208 480227 587210
rect 476940 587152 480166 587208
rect 480222 587152 480227 587208
rect 476940 587150 480227 587152
rect 480161 587147 480227 587150
rect 0 586938 800 586968
rect 486200 586938 487000 586968
rect 0 586878 9506 586938
rect 476940 586878 487000 586938
rect 0 586848 800 586878
rect 9446 586752 9506 586878
rect 486200 586848 487000 586878
rect 9446 586692 10060 586752
rect 479742 586666 479748 586668
rect 476940 586606 479748 586666
rect 479742 586604 479748 586606
rect 479812 586604 479818 586668
rect 476940 586334 483306 586394
rect 483246 586258 483306 586334
rect 486200 586258 487000 586288
rect 477358 586208 482938 586258
rect 476928 586198 482938 586208
rect 483246 586198 487000 586258
rect 476928 586148 477418 586198
rect 482878 585986 482938 586198
rect 486200 586168 487000 586198
rect 486182 585986 486188 585988
rect 482878 585926 486188 585986
rect 486182 585924 486188 585926
rect 486252 585924 486258 585988
rect 9446 585820 10060 585880
rect 486366 585850 486372 585852
rect 0 585578 800 585608
rect 9446 585578 9506 585820
rect 476940 585790 486372 585850
rect 486366 585788 486372 585790
rect 486436 585788 486442 585852
rect 486200 585578 487000 585608
rect 0 585518 9506 585578
rect 476940 585518 487000 585578
rect 0 585488 800 585518
rect 486200 585488 487000 585518
rect 478086 585306 478092 585308
rect 476940 585246 478092 585306
rect 478086 585244 478092 585246
rect 478156 585244 478162 585308
rect 9446 585004 10060 585064
rect 0 584898 800 584928
rect 9446 584898 9506 585004
rect 476940 584974 480270 585034
rect 0 584838 9506 584898
rect 480210 584898 480270 584974
rect 486200 584898 487000 584928
rect 480210 584838 487000 584898
rect 0 584808 800 584838
rect 486200 584808 487000 584838
rect 477125 584762 477191 584765
rect 476940 584760 477191 584762
rect 476940 584704 477130 584760
rect 477186 584704 477191 584760
rect 476940 584702 477191 584704
rect 477125 584699 477191 584702
rect 483657 584626 483723 584629
rect 477358 584624 483723 584626
rect 477358 584576 483662 584624
rect 476928 584568 483662 584576
rect 483718 584568 483723 584624
rect 476928 584566 483723 584568
rect 476928 584516 477418 584566
rect 483657 584563 483723 584566
rect 0 584218 800 584248
rect 9446 584218 10060 584248
rect 486200 584218 487000 584248
rect 0 584188 10060 584218
rect 0 584158 9506 584188
rect 476940 584158 487000 584218
rect 0 584128 800 584158
rect 486200 584128 487000 584158
rect 478270 583946 478276 583948
rect 476940 583886 478276 583946
rect 478270 583884 478276 583886
rect 478340 583884 478346 583948
rect 476940 583614 480270 583674
rect 0 583538 800 583568
rect 480210 583538 480270 583614
rect 486200 583538 487000 583568
rect 0 583488 9506 583538
rect 0 583478 10060 583488
rect 480210 583478 487000 583538
rect 0 583448 800 583478
rect 9446 583428 10060 583478
rect 486200 583448 487000 583478
rect 478638 583402 478644 583404
rect 476940 583342 478644 583402
rect 478638 583340 478644 583342
rect 478708 583340 478714 583404
rect 478454 583130 478460 583132
rect 476940 583070 478460 583130
rect 478454 583068 478460 583070
rect 478524 583068 478530 583132
rect 0 582858 800 582888
rect 486200 582858 487000 582888
rect 0 582798 9506 582858
rect 476940 582798 487000 582858
rect 0 582768 800 582798
rect 9446 582672 9506 582798
rect 486200 582768 487000 582798
rect 9446 582612 10060 582672
rect 485446 582586 485452 582588
rect 476940 582526 485452 582586
rect 485446 582524 485452 582526
rect 485516 582524 485522 582588
rect 481766 582388 481772 582452
rect 481836 582450 481842 582452
rect 482921 582450 482987 582453
rect 481836 582448 482987 582450
rect 481836 582392 482926 582448
rect 482982 582392 482987 582448
rect 481836 582390 482987 582392
rect 481836 582388 481842 582390
rect 482921 582387 482987 582390
rect 476940 582254 483306 582314
rect 483246 582178 483306 582254
rect 486200 582178 487000 582208
rect 483246 582118 487000 582178
rect 486200 582088 487000 582118
rect 485998 582042 486004 582044
rect 476940 581982 486004 582042
rect 485998 581980 486004 581982
rect 486068 581980 486074 582044
rect 485262 581906 485268 581908
rect 477358 581856 485268 581906
rect 476928 581846 485268 581856
rect 9446 581740 10060 581800
rect 476928 581796 477418 581846
rect 485262 581844 485268 581846
rect 485332 581844 485338 581908
rect 0 581498 800 581528
rect 9446 581498 9506 581740
rect 479742 581572 479748 581636
rect 479812 581634 479818 581636
rect 480069 581634 480135 581637
rect 479812 581632 480135 581634
rect 479812 581576 480074 581632
rect 480130 581576 480135 581632
rect 479812 581574 480135 581576
rect 479812 581572 479818 581574
rect 480069 581571 480135 581574
rect 483054 581572 483060 581636
rect 483124 581634 483130 581636
rect 484301 581634 484367 581637
rect 483124 581632 484367 581634
rect 483124 581576 484306 581632
rect 484362 581576 484367 581632
rect 483124 581574 484367 581576
rect 483124 581572 483130 581574
rect 484301 581571 484367 581574
rect 486200 581498 487000 581528
rect 0 581438 9506 581498
rect 476940 581438 487000 581498
rect 0 581408 800 581438
rect 486200 581408 487000 581438
rect 485814 581362 485820 581364
rect 477358 581312 485820 581362
rect 476928 581302 485820 581312
rect 476928 581252 477418 581302
rect 485814 581300 485820 581302
rect 485884 581300 485890 581364
rect 9446 580924 10060 580984
rect 0 580818 800 580848
rect 9446 580818 9506 580924
rect 476940 580894 480270 580954
rect 0 580758 9506 580818
rect 480210 580818 480270 580894
rect 481214 580892 481220 580956
rect 481284 580954 481290 580956
rect 481449 580954 481515 580957
rect 481284 580952 481515 580954
rect 481284 580896 481454 580952
rect 481510 580896 481515 580952
rect 481284 580894 481515 580896
rect 481284 580892 481290 580894
rect 481449 580891 481515 580894
rect 486200 580818 487000 580848
rect 480210 580758 487000 580818
rect 0 580728 800 580758
rect 486200 580728 487000 580758
rect 485078 580682 485084 580684
rect 476940 580622 485084 580682
rect 485078 580620 485084 580622
rect 485148 580620 485154 580684
rect 485630 580546 485636 580548
rect 477358 580496 485636 580546
rect 476928 580486 485636 580496
rect 476928 580436 477418 580486
rect 485630 580484 485636 580486
rect 485700 580484 485706 580548
rect 0 580138 800 580168
rect 9446 580138 10060 580168
rect 486200 580138 487000 580168
rect 0 580108 10060 580138
rect 0 580078 9506 580108
rect 476940 580078 487000 580138
rect 0 580048 800 580078
rect 486200 580048 487000 580078
rect 477350 579866 477356 579868
rect 476940 579806 477356 579866
rect 477350 579804 477356 579806
rect 477420 579804 477426 579868
rect 476940 579534 480270 579594
rect 0 579458 800 579488
rect 480210 579458 480270 579534
rect 481582 579532 481588 579596
rect 481652 579594 481658 579596
rect 482829 579594 482895 579597
rect 481652 579592 482895 579594
rect 481652 579536 482834 579592
rect 482890 579536 482895 579592
rect 481652 579534 482895 579536
rect 481652 579532 481658 579534
rect 482829 579531 482895 579534
rect 486200 579458 487000 579488
rect 0 579408 9506 579458
rect 0 579398 10060 579408
rect 480210 579398 487000 579458
rect 0 579368 800 579398
rect 9446 579348 10060 579398
rect 486200 579368 487000 579398
rect 482870 579322 482876 579324
rect 476940 579262 482876 579322
rect 482870 579260 482876 579262
rect 482940 579260 482946 579324
rect 477358 579136 483306 579186
rect 476928 579126 483306 579136
rect 476928 579076 477418 579126
rect 480294 578988 480300 579052
rect 480364 579050 480370 579052
rect 481357 579050 481423 579053
rect 480364 579048 481423 579050
rect 480364 578992 481362 579048
rect 481418 578992 481423 579048
rect 480364 578990 481423 578992
rect 480364 578988 480370 578990
rect 481357 578987 481423 578990
rect 0 578778 800 578808
rect 476940 578778 477418 578808
rect 482502 578778 482508 578780
rect 0 578718 9506 578778
rect 476940 578748 482508 578778
rect 477358 578718 482508 578748
rect 0 578688 800 578718
rect 9446 578592 9506 578718
rect 482502 578716 482508 578718
rect 482572 578716 482578 578780
rect 483246 578778 483306 579126
rect 486200 578778 487000 578808
rect 483246 578718 487000 578778
rect 486200 578688 487000 578718
rect 9446 578532 10060 578592
rect 482870 578036 482876 578100
rect 482940 578098 482946 578100
rect 486200 578098 487000 578128
rect 482940 578038 487000 578098
rect 482940 578036 482946 578038
rect 486200 578008 487000 578038
rect 9446 577660 10060 577720
rect 0 577418 800 577448
rect 9446 577418 9506 577660
rect 0 577358 9506 577418
rect 0 577328 800 577358
rect 477350 577356 477356 577420
rect 477420 577418 477426 577420
rect 486200 577418 487000 577448
rect 477420 577358 487000 577418
rect 477420 577356 477426 577358
rect 486200 577328 487000 577358
rect 9446 576874 10060 576904
rect 5582 576844 10060 576874
rect 5582 576814 9506 576844
rect 0 576738 800 576768
rect 5582 576738 5642 576814
rect 0 576678 5642 576738
rect 0 576648 800 576678
rect 485630 576676 485636 576740
rect 485700 576738 485706 576740
rect 486200 576738 487000 576768
rect 485700 576678 487000 576738
rect 485700 576676 485706 576678
rect 486200 576648 487000 576678
rect 0 576058 800 576088
rect 9446 576058 10060 576088
rect 0 576028 10060 576058
rect 0 575998 9506 576028
rect 0 575968 800 575998
rect 485078 575996 485084 576060
rect 485148 576058 485154 576060
rect 486200 576058 487000 576088
rect 485148 575998 487000 576058
rect 485148 575996 485154 575998
rect 486200 575968 487000 575998
rect 0 575378 800 575408
rect 0 575328 9506 575378
rect 0 575318 10060 575328
rect 0 575288 800 575318
rect 9446 575268 10060 575318
rect 485814 575316 485820 575380
rect 485884 575378 485890 575380
rect 486200 575378 487000 575408
rect 485884 575318 487000 575378
rect 485884 575316 485890 575318
rect 486200 575288 487000 575318
rect 0 574698 800 574728
rect 0 574638 9506 574698
rect 0 574608 800 574638
rect 9446 574512 9506 574638
rect 485262 574636 485268 574700
rect 485332 574698 485338 574700
rect 486200 574698 487000 574728
rect 485332 574638 487000 574698
rect 485332 574636 485338 574638
rect 486200 574608 487000 574638
rect 9446 574452 10060 574512
rect 485998 573956 486004 574020
rect 486068 574018 486074 574020
rect 486200 574018 487000 574048
rect 486068 573958 487000 574018
rect 486068 573956 486074 573958
rect 486200 573928 487000 573958
rect 9446 573580 10060 573640
rect 0 573338 800 573368
rect 9446 573338 9506 573580
rect 0 573278 9506 573338
rect 0 573248 800 573278
rect 485446 573276 485452 573340
rect 485516 573338 485522 573340
rect 486200 573338 487000 573368
rect 485516 573278 487000 573338
rect 485516 573276 485522 573278
rect 486200 573248 487000 573278
rect 9446 572794 10060 572824
rect 6870 572764 10060 572794
rect 6870 572734 9506 572764
rect 0 572658 800 572688
rect 6870 572658 6930 572734
rect 0 572598 6930 572658
rect 0 572568 800 572598
rect 478454 572596 478460 572660
rect 478524 572658 478530 572660
rect 486200 572658 487000 572688
rect 478524 572598 487000 572658
rect 478524 572596 478530 572598
rect 486200 572568 487000 572598
rect 0 571978 800 572008
rect 9446 571978 10060 572008
rect 0 571948 10060 571978
rect 0 571918 9506 571948
rect 0 571888 800 571918
rect 478638 571916 478644 571980
rect 478708 571978 478714 571980
rect 486200 571978 487000 572008
rect 478708 571918 487000 571978
rect 478708 571916 478714 571918
rect 486200 571888 487000 571918
rect 0 571298 800 571328
rect 0 571248 9506 571298
rect 0 571238 10060 571248
rect 0 571208 800 571238
rect 9446 571188 10060 571238
rect 478270 571236 478276 571300
rect 478340 571298 478346 571300
rect 486200 571298 487000 571328
rect 478340 571238 487000 571298
rect 478340 571236 478346 571238
rect 486200 571208 487000 571238
rect 0 570618 800 570648
rect 483657 570618 483723 570621
rect 486200 570618 487000 570648
rect 0 570558 9506 570618
rect 0 570528 800 570558
rect 9446 570432 9506 570558
rect 483657 570616 487000 570618
rect 483657 570560 483662 570616
rect 483718 570560 487000 570616
rect 483657 570558 487000 570560
rect 483657 570555 483723 570558
rect 486200 570528 487000 570558
rect 9446 570372 10060 570432
rect 477125 569938 477191 569941
rect 486200 569938 487000 569968
rect 477125 569936 487000 569938
rect 477125 569880 477130 569936
rect 477186 569880 487000 569936
rect 477125 569878 487000 569880
rect 477125 569875 477191 569878
rect 486200 569848 487000 569878
rect 9446 569500 10060 569560
rect 0 569258 800 569288
rect 9446 569258 9506 569500
rect 0 569198 9506 569258
rect 0 569168 800 569198
rect 478086 569196 478092 569260
rect 478156 569258 478162 569260
rect 486200 569258 487000 569288
rect 478156 569198 487000 569258
rect 478156 569196 478162 569198
rect 486200 569168 487000 569198
rect 9446 568714 10060 568744
rect 6870 568684 10060 568714
rect 6870 568654 9506 568684
rect 0 568578 800 568608
rect 6870 568578 6930 568654
rect 0 568518 6930 568578
rect 486200 568580 487000 568608
rect 0 568488 800 568518
rect 486200 568516 486372 568580
rect 486436 568516 487000 568580
rect 486200 568488 487000 568516
rect 0 567898 800 567928
rect 9446 567898 10060 567928
rect 0 567868 10060 567898
rect 486200 567900 487000 567928
rect 0 567838 9506 567868
rect 0 567808 800 567838
rect 486200 567836 486372 567900
rect 486436 567836 487000 567900
rect 486200 567808 487000 567836
rect 0 567218 800 567248
rect 480069 567218 480135 567221
rect 486200 567218 487000 567248
rect 0 567158 4906 567218
rect 0 567128 800 567158
rect 4846 567082 4906 567158
rect 480069 567216 487000 567218
rect 480069 567160 480074 567216
rect 480130 567160 487000 567216
rect 480069 567158 487000 567160
rect 480069 567155 480135 567158
rect 486200 567128 487000 567158
rect 9446 567082 10060 567112
rect 4846 567052 10060 567082
rect 4846 567022 9506 567052
rect 0 566538 800 566568
rect 480161 566538 480227 566541
rect 486200 566538 487000 566568
rect 0 566478 9506 566538
rect 0 566448 800 566478
rect 9446 566352 9506 566478
rect 480161 566536 487000 566538
rect 480161 566480 480166 566536
rect 480222 566480 487000 566536
rect 480161 566478 487000 566480
rect 480161 566475 480227 566478
rect 486200 566448 487000 566478
rect 9446 566292 10060 566352
rect 482502 565796 482508 565860
rect 482572 565858 482578 565860
rect 486200 565858 487000 565888
rect 482572 565798 487000 565858
rect 482572 565796 482578 565798
rect 486200 565768 487000 565798
rect 9446 565420 10060 565480
rect 0 565178 800 565208
rect 9446 565178 9506 565420
rect 0 565118 9506 565178
rect 0 565088 800 565118
rect 481030 565116 481036 565180
rect 481100 565178 481106 565180
rect 486200 565178 487000 565208
rect 481100 565118 487000 565178
rect 481100 565116 481106 565118
rect 486200 565088 487000 565118
rect 9446 564604 10060 564664
rect 0 564498 800 564528
rect 9446 564498 9506 564604
rect 0 564438 9506 564498
rect 0 564408 800 564438
rect 482318 564436 482324 564500
rect 482388 564498 482394 564500
rect 486200 564498 487000 564528
rect 482388 564438 487000 564498
rect 482388 564436 482394 564438
rect 486200 564408 487000 564438
rect 0 563818 800 563848
rect 9446 563818 10060 563848
rect 0 563788 10060 563818
rect 0 563758 9506 563788
rect 0 563728 800 563758
rect 480846 563756 480852 563820
rect 480916 563818 480922 563820
rect 486200 563818 487000 563848
rect 480916 563758 487000 563818
rect 480916 563756 480922 563758
rect 486200 563728 487000 563758
rect 0 563138 800 563168
rect 0 563078 4170 563138
rect 0 563048 800 563078
rect 4110 563002 4170 563078
rect 483974 563076 483980 563140
rect 484044 563138 484050 563140
rect 486200 563138 487000 563168
rect 484044 563078 487000 563138
rect 484044 563076 484050 563078
rect 486200 563048 487000 563078
rect 9446 563002 10060 563032
rect 4110 562972 10060 563002
rect 4110 562942 9506 562972
rect 0 562458 800 562488
rect 0 562398 9506 562458
rect 0 562368 800 562398
rect 9446 562272 9506 562398
rect 482134 562396 482140 562460
rect 482204 562458 482210 562460
rect 486200 562458 487000 562488
rect 482204 562398 487000 562458
rect 482204 562396 482210 562398
rect 486200 562368 487000 562398
rect 9446 562212 10060 562272
rect 481357 561778 481423 561781
rect 486200 561778 487000 561808
rect 481357 561776 487000 561778
rect 481357 561720 481362 561776
rect 481418 561720 487000 561776
rect 481357 561718 487000 561720
rect 481357 561715 481423 561718
rect 486200 561688 487000 561718
rect 9446 561340 10060 561400
rect 0 561098 800 561128
rect 9446 561098 9506 561340
rect 0 561038 9506 561098
rect 482829 561098 482895 561101
rect 486200 561098 487000 561128
rect 482829 561096 487000 561098
rect 482829 561040 482834 561096
rect 482890 561040 487000 561096
rect 482829 561038 487000 561040
rect 0 561008 800 561038
rect 482829 561035 482895 561038
rect 486200 561008 487000 561038
rect 483790 560356 483796 560420
rect 483860 560418 483866 560420
rect 486200 560418 487000 560448
rect 483860 560358 487000 560418
rect 483860 560356 483866 560358
rect 486200 560328 487000 560358
rect 482921 559738 482987 559741
rect 486200 559738 487000 559768
rect 482921 559736 487000 559738
rect 482921 559680 482926 559736
rect 482982 559680 487000 559736
rect 482921 559678 487000 559680
rect 482921 559675 482987 559678
rect 486200 559648 487000 559678
rect 483606 558996 483612 559060
rect 483676 559058 483682 559060
rect 486200 559058 487000 559088
rect 483676 558998 487000 559058
rect 483676 558996 483682 558998
rect 486200 558968 487000 558998
rect 481541 558378 481607 558381
rect 486200 558378 487000 558408
rect 481541 558376 487000 558378
rect 481541 558320 481546 558376
rect 481602 558320 487000 558376
rect 481541 558318 487000 558320
rect 481541 558315 481607 558318
rect 486200 558288 487000 558318
rect 484301 557698 484367 557701
rect 486200 557698 487000 557728
rect 484301 557696 487000 557698
rect 484301 557640 484306 557696
rect 484362 557640 487000 557696
rect 484301 557638 487000 557640
rect 484301 557635 484367 557638
rect 486200 557608 487000 557638
rect 481449 557018 481515 557021
rect 486200 557018 487000 557048
rect 481449 557016 487000 557018
rect 481449 556960 481454 557016
rect 481510 556960 487000 557016
rect 481449 556958 487000 556960
rect 481449 556955 481515 556958
rect 486200 556928 487000 556958
rect 9446 553060 10060 553120
rect 0 552938 800 552968
rect 9446 552938 9506 553060
rect 0 552878 9506 552938
rect 0 552848 800 552878
rect 0 552258 800 552288
rect 9446 552258 10060 552304
rect 0 552244 10060 552258
rect 0 552198 9506 552244
rect 0 552168 800 552198
rect 0 551578 800 551608
rect 0 551544 9506 551578
rect 0 551518 10060 551544
rect 0 551488 800 551518
rect 9446 551484 10060 551518
rect 0 550898 800 550928
rect 0 550838 9506 550898
rect 0 550808 800 550838
rect 9446 550728 9506 550838
rect 9446 550668 10060 550728
rect 0 550218 800 550248
rect 0 550158 9506 550218
rect 0 550128 800 550158
rect 9446 549912 9506 550158
rect 9446 549852 10060 549912
rect 9446 548980 10060 549040
rect 0 548858 800 548888
rect 9446 548858 9506 548980
rect 0 548798 9506 548858
rect 0 548768 800 548798
rect 0 548178 800 548208
rect 9446 548178 10060 548224
rect 0 548164 10060 548178
rect 0 548118 9506 548164
rect 0 548088 800 548118
rect 0 547498 800 547528
rect 0 547464 9506 547498
rect 0 547438 10060 547464
rect 0 547408 800 547438
rect 9446 547404 10060 547438
rect 0 546818 800 546848
rect 0 546758 9506 546818
rect 0 546728 800 546758
rect 9446 546648 9506 546758
rect 9446 546588 10060 546648
rect 0 546138 800 546168
rect 0 546078 9506 546138
rect 0 546048 800 546078
rect 9446 545832 9506 546078
rect 9446 545772 10060 545832
rect 9446 544900 10060 544960
rect 0 544778 800 544808
rect 9446 544778 9506 544900
rect 0 544718 9506 544778
rect 0 544688 800 544718
rect 0 544098 800 544128
rect 9446 544098 10060 544144
rect 0 544084 10060 544098
rect 0 544038 9506 544084
rect 0 544008 800 544038
rect 0 543418 800 543448
rect 0 543384 9506 543418
rect 0 543358 10060 543384
rect 0 543328 800 543358
rect 9446 543324 10060 543358
rect 0 542738 800 542768
rect 0 542678 9506 542738
rect 0 542648 800 542678
rect 9446 542568 9506 542678
rect 9446 542508 10060 542568
rect 0 542058 800 542088
rect 0 541998 9506 542058
rect 0 541968 800 541998
rect 9446 541752 9506 541998
rect 9446 541692 10060 541752
rect 9446 540820 10060 540880
rect 0 540698 800 540728
rect 9446 540698 9506 540820
rect 0 540638 9506 540698
rect 0 540608 800 540638
rect 0 540018 800 540048
rect 9446 540018 10060 540064
rect 0 540004 10060 540018
rect 481541 540018 481607 540021
rect 486200 540018 487000 540048
rect 481541 540016 487000 540018
rect 0 539958 9506 540004
rect 481541 539960 481546 540016
rect 481602 539960 487000 540016
rect 481541 539958 487000 539960
rect 0 539928 800 539958
rect 481541 539955 481607 539958
rect 486200 539928 487000 539958
rect 0 539338 800 539368
rect 482921 539338 482987 539341
rect 486200 539338 487000 539368
rect 0 539304 9506 539338
rect 482921 539336 487000 539338
rect 0 539278 10060 539304
rect 0 539248 800 539278
rect 9446 539244 10060 539278
rect 482921 539280 482926 539336
rect 482982 539280 487000 539336
rect 482921 539278 487000 539280
rect 482921 539275 482987 539278
rect 486200 539248 487000 539278
rect 0 538658 800 538688
rect 481449 538658 481515 538661
rect 486200 538658 487000 538688
rect 0 538598 9506 538658
rect 0 538568 800 538598
rect 9446 538488 9506 538598
rect 481449 538656 487000 538658
rect 481449 538600 481454 538656
rect 481510 538600 487000 538656
rect 481449 538598 487000 538600
rect 481449 538595 481515 538598
rect 486200 538568 487000 538598
rect 9446 538428 10060 538488
rect 0 537978 800 538008
rect 484301 537978 484367 537981
rect 486200 537978 487000 538008
rect 0 537918 9506 537978
rect 0 537888 800 537918
rect 9446 537672 9506 537918
rect 484301 537976 487000 537978
rect 484301 537920 484306 537976
rect 484362 537920 487000 537976
rect 484301 537918 487000 537920
rect 484301 537915 484367 537918
rect 486200 537888 487000 537918
rect 9446 537612 10060 537672
rect 482829 537298 482895 537301
rect 486200 537298 487000 537328
rect 482829 537296 487000 537298
rect 482829 537240 482834 537296
rect 482890 537240 487000 537296
rect 482829 537238 487000 537240
rect 482829 537235 482895 537238
rect 486200 537208 487000 537238
rect 9446 536740 10060 536800
rect 0 536618 800 536648
rect 9446 536618 9506 536740
rect 0 536558 9506 536618
rect 0 536528 800 536558
rect 480846 536556 480852 536620
rect 480916 536618 480922 536620
rect 486200 536618 487000 536648
rect 480916 536558 487000 536618
rect 480916 536556 480922 536558
rect 486200 536528 487000 536558
rect 0 535938 800 535968
rect 9446 535938 10060 535984
rect 0 535924 10060 535938
rect 484209 535938 484275 535941
rect 486200 535938 487000 535968
rect 484209 535936 487000 535938
rect 0 535878 9506 535924
rect 484209 535880 484214 535936
rect 484270 535880 487000 535936
rect 484209 535878 487000 535880
rect 0 535848 800 535878
rect 484209 535875 484275 535878
rect 486200 535848 487000 535878
rect 0 535258 800 535288
rect 0 535224 9506 535258
rect 0 535198 10060 535224
rect 0 535168 800 535198
rect 9446 535164 10060 535198
rect 482134 535196 482140 535260
rect 482204 535258 482210 535260
rect 486200 535258 487000 535288
rect 482204 535198 487000 535258
rect 482204 535196 482210 535198
rect 486200 535168 487000 535198
rect 0 534578 800 534608
rect 478781 534578 478847 534581
rect 486200 534578 487000 534608
rect 0 534518 9506 534578
rect 0 534488 800 534518
rect 9446 534408 9506 534518
rect 478781 534576 487000 534578
rect 478781 534520 478786 534576
rect 478842 534520 487000 534576
rect 478781 534518 487000 534520
rect 478781 534515 478847 534518
rect 486200 534488 487000 534518
rect 9446 534348 10060 534408
rect 0 533898 800 533928
rect 0 533838 9506 533898
rect 0 533808 800 533838
rect 9446 533592 9506 533838
rect 478086 533836 478092 533900
rect 478156 533898 478162 533900
rect 486200 533898 487000 533928
rect 478156 533838 487000 533898
rect 478156 533836 478162 533838
rect 486200 533808 487000 533838
rect 9446 533532 10060 533592
rect 478689 533218 478755 533221
rect 486200 533218 487000 533248
rect 478689 533216 487000 533218
rect 478689 533160 478694 533216
rect 478750 533160 487000 533216
rect 478689 533158 487000 533160
rect 478689 533155 478755 533158
rect 486200 533128 487000 533158
rect 6870 532776 9506 532810
rect 6870 532750 10060 532776
rect 0 532538 800 532568
rect 6870 532538 6930 532750
rect 9446 532716 10060 532750
rect 0 532478 6930 532538
rect 0 532448 800 532478
rect 478270 532476 478276 532540
rect 478340 532538 478346 532540
rect 486200 532538 487000 532568
rect 478340 532478 487000 532538
rect 478340 532476 478346 532478
rect 486200 532448 487000 532478
rect 0 531858 800 531888
rect 9446 531858 10060 531904
rect 0 531844 10060 531858
rect 0 531798 9506 531844
rect 0 531768 800 531798
rect 483606 531796 483612 531860
rect 483676 531858 483682 531860
rect 486200 531858 487000 531888
rect 483676 531798 487000 531858
rect 483676 531796 483682 531798
rect 486200 531768 487000 531798
rect 0 531178 800 531208
rect 0 531144 9506 531178
rect 0 531118 10060 531144
rect 0 531088 800 531118
rect 9446 531084 10060 531118
rect 481030 531116 481036 531180
rect 481100 531178 481106 531180
rect 486200 531178 487000 531208
rect 481100 531118 487000 531178
rect 481100 531116 481106 531118
rect 486200 531088 487000 531118
rect 0 530498 800 530528
rect 483657 530498 483723 530501
rect 486200 530498 487000 530528
rect 0 530438 9506 530498
rect 0 530408 800 530438
rect 9446 530328 9506 530438
rect 483657 530496 487000 530498
rect 483657 530440 483662 530496
rect 483718 530440 487000 530496
rect 483657 530438 487000 530440
rect 483657 530435 483723 530438
rect 486200 530408 487000 530438
rect 9446 530268 10060 530328
rect 0 529818 800 529848
rect 0 529758 9506 529818
rect 0 529728 800 529758
rect 9446 529512 9506 529758
rect 479558 529756 479564 529820
rect 479628 529818 479634 529820
rect 486200 529818 487000 529848
rect 479628 529758 487000 529818
rect 479628 529756 479634 529758
rect 486200 529728 487000 529758
rect 9446 529452 10060 529512
rect 485078 529076 485084 529140
rect 485148 529138 485154 529140
rect 486200 529138 487000 529168
rect 485148 529078 487000 529138
rect 485148 529076 485154 529078
rect 486200 529048 487000 529078
rect 9446 528594 10060 528640
rect 5582 528580 10060 528594
rect 5582 528534 9506 528580
rect 0 528458 800 528488
rect 5582 528458 5642 528534
rect 0 528398 5642 528458
rect 486200 528460 487000 528488
rect 0 528368 800 528398
rect 486200 528396 486372 528460
rect 486436 528396 487000 528460
rect 486200 528368 487000 528396
rect 0 527778 800 527808
rect 9446 527778 10060 527824
rect 0 527764 10060 527778
rect 0 527718 9506 527764
rect 0 527688 800 527718
rect 485262 527716 485268 527780
rect 485332 527778 485338 527780
rect 486200 527778 487000 527808
rect 485332 527718 487000 527778
rect 485332 527716 485338 527718
rect 486200 527688 487000 527718
rect 0 527098 800 527128
rect 0 527064 9506 527098
rect 0 527038 10060 527064
rect 0 527008 800 527038
rect 9446 527004 10060 527038
rect 481214 527036 481220 527100
rect 481284 527098 481290 527100
rect 486200 527098 487000 527128
rect 481284 527038 487000 527098
rect 481284 527036 481290 527038
rect 486200 527008 487000 527038
rect 0 526418 800 526448
rect 0 526358 9506 526418
rect 0 526328 800 526358
rect 9446 526248 9506 526358
rect 479374 526356 479380 526420
rect 479444 526418 479450 526420
rect 486200 526418 487000 526448
rect 479444 526358 487000 526418
rect 479444 526356 479450 526358
rect 486200 526328 487000 526358
rect 9446 526188 10060 526248
rect 0 525738 800 525768
rect 0 525678 9506 525738
rect 0 525648 800 525678
rect 9446 525432 9506 525678
rect 483974 525676 483980 525740
rect 484044 525738 484050 525740
rect 486200 525738 487000 525768
rect 484044 525678 487000 525738
rect 484044 525676 484050 525678
rect 486200 525648 487000 525678
rect 9446 525372 10060 525432
rect 485998 524996 486004 525060
rect 486068 525058 486074 525060
rect 486200 525058 487000 525088
rect 486068 524998 487000 525058
rect 486068 524996 486074 524998
rect 486200 524968 487000 524998
rect 9446 524514 10060 524560
rect 6870 524500 10060 524514
rect 6870 524454 9506 524500
rect 0 524378 800 524408
rect 6870 524378 6930 524454
rect 0 524318 6930 524378
rect 0 524288 800 524318
rect 479742 524316 479748 524380
rect 479812 524378 479818 524380
rect 486200 524378 487000 524408
rect 479812 524318 487000 524378
rect 479812 524316 479818 524318
rect 486200 524288 487000 524318
rect 0 523698 800 523728
rect 9446 523698 10060 523744
rect 0 523684 10060 523698
rect 0 523638 9506 523684
rect 0 523608 800 523638
rect 483790 523636 483796 523700
rect 483860 523698 483866 523700
rect 486200 523698 487000 523728
rect 483860 523638 487000 523698
rect 483860 523636 483866 523638
rect 486200 523608 487000 523638
rect 0 523018 800 523048
rect 0 522984 9506 523018
rect 0 522958 10060 522984
rect 0 522928 800 522958
rect 9446 522924 10060 522958
rect 480662 522956 480668 523020
rect 480732 523018 480738 523020
rect 486200 523018 487000 523048
rect 480732 522958 487000 523018
rect 480732 522956 480738 522958
rect 486200 522928 487000 522958
rect 0 522338 800 522368
rect 486200 522340 487000 522368
rect 0 522278 9506 522338
rect 0 522248 800 522278
rect 9446 522168 9506 522278
rect 486200 522276 486372 522340
rect 486436 522276 487000 522340
rect 486200 522248 487000 522276
rect 9446 522108 10060 522168
rect 0 521658 800 521688
rect 0 521598 9506 521658
rect 0 521568 800 521598
rect 9446 521352 9506 521598
rect 485814 521596 485820 521660
rect 485884 521658 485890 521660
rect 486200 521658 487000 521688
rect 485884 521598 487000 521658
rect 485884 521596 485890 521598
rect 486200 521568 487000 521598
rect 9446 521292 10060 521352
rect 484526 520916 484532 520980
rect 484596 520978 484602 520980
rect 486200 520978 487000 521008
rect 484596 520918 487000 520978
rect 484596 520916 484602 520918
rect 486200 520888 487000 520918
rect 9446 520420 10060 520480
rect 0 520298 800 520328
rect 9446 520298 9506 520420
rect 0 520238 9506 520298
rect 0 520208 800 520238
rect 484710 520236 484716 520300
rect 484780 520298 484786 520300
rect 486200 520298 487000 520328
rect 484780 520238 487000 520298
rect 484780 520236 484786 520238
rect 486200 520208 487000 520238
rect 0 519618 800 519648
rect 9446 519618 10060 519664
rect 0 519604 10060 519618
rect 0 519558 9506 519604
rect 0 519528 800 519558
rect 484342 519556 484348 519620
rect 484412 519618 484418 519620
rect 486200 519618 487000 519648
rect 484412 519558 487000 519618
rect 484412 519556 484418 519558
rect 486200 519528 487000 519558
rect 0 518938 800 518968
rect 0 518878 4906 518938
rect 0 518848 800 518878
rect 4846 518802 4906 518878
rect 484894 518876 484900 518940
rect 484964 518938 484970 518940
rect 486200 518938 487000 518968
rect 484964 518878 487000 518938
rect 484964 518876 484970 518878
rect 486200 518848 487000 518878
rect 9446 518802 10060 518848
rect 4846 518788 10060 518802
rect 4846 518742 9506 518788
rect 0 518258 800 518288
rect 479558 518258 479564 518260
rect 0 518198 9506 518258
rect 477358 518240 479564 518258
rect 0 518168 800 518198
rect 9446 518088 9506 518198
rect 476940 518198 479564 518240
rect 476940 518180 477418 518198
rect 479558 518196 479564 518198
rect 479628 518196 479634 518260
rect 479926 518196 479932 518260
rect 479996 518258 480002 518260
rect 486200 518258 487000 518288
rect 479996 518198 487000 518258
rect 479996 518196 480002 518198
rect 486200 518168 487000 518198
rect 9446 518028 10060 518088
rect 483974 517986 483980 517988
rect 477358 517968 483980 517986
rect 476940 517926 483980 517968
rect 476940 517908 477418 517926
rect 483974 517924 483980 517926
rect 484044 517924 484050 517988
rect 484342 517714 484348 517716
rect 477358 517696 484348 517714
rect 476940 517654 484348 517696
rect 476940 517636 477418 517654
rect 484342 517652 484348 517654
rect 484412 517652 484418 517716
rect 0 517578 800 517608
rect 486200 517578 487000 517608
rect 0 517518 4170 517578
rect 0 517488 800 517518
rect 4110 517442 4170 517518
rect 483246 517518 487000 517578
rect 483246 517442 483306 517518
rect 486200 517488 487000 517518
rect 4110 517382 9506 517442
rect 477358 517424 483306 517442
rect 9446 517272 9506 517382
rect 476940 517382 483306 517424
rect 476940 517364 477418 517382
rect 478597 517306 478663 517309
rect 486182 517306 486188 517308
rect 478597 517304 486188 517306
rect 9446 517212 10060 517272
rect 478597 517248 478602 517304
rect 478658 517248 486188 517304
rect 478597 517246 486188 517248
rect 478597 517243 478663 517246
rect 486182 517244 486188 517246
rect 486252 517244 486258 517308
rect 484710 517170 484716 517172
rect 477358 517152 484716 517170
rect 476940 517110 484716 517152
rect 476940 517092 477418 517110
rect 484710 517108 484716 517110
rect 484780 517108 484786 517172
rect 478597 516898 478663 516901
rect 486200 516898 487000 516928
rect 477358 516896 478663 516898
rect 477358 516880 478602 516896
rect 476940 516840 478602 516880
rect 478658 516840 478663 516896
rect 476940 516838 478663 516840
rect 476940 516820 477418 516838
rect 478597 516835 478663 516838
rect 480210 516838 487000 516898
rect 478454 516700 478460 516764
rect 478524 516762 478530 516764
rect 480210 516762 480270 516838
rect 486200 516808 487000 516838
rect 478524 516702 480270 516762
rect 478524 516700 478530 516702
rect 484526 516626 484532 516628
rect 477358 516608 484532 516626
rect 476940 516566 484532 516608
rect 476940 516548 477418 516566
rect 484526 516564 484532 516566
rect 484596 516564 484602 516628
rect 483657 516490 483723 516493
rect 480210 516488 483723 516490
rect 480210 516432 483662 516488
rect 483718 516432 483723 516488
rect 480210 516430 483723 516432
rect 9446 516340 10060 516400
rect 480210 516354 480270 516430
rect 483657 516427 483723 516430
rect 0 516218 800 516248
rect 9446 516218 9506 516340
rect 477358 516336 480270 516354
rect 476940 516294 480270 516336
rect 476940 516276 477418 516294
rect 483054 516292 483060 516356
rect 483124 516354 483130 516356
rect 484209 516354 484275 516357
rect 483124 516352 484275 516354
rect 483124 516296 484214 516352
rect 484270 516296 484275 516352
rect 483124 516294 484275 516296
rect 483124 516292 483130 516294
rect 484209 516291 484275 516294
rect 0 516158 9506 516218
rect 0 516128 800 516158
rect 481582 516156 481588 516220
rect 481652 516218 481658 516220
rect 482829 516218 482895 516221
rect 486200 516218 487000 516248
rect 481652 516216 482895 516218
rect 481652 516160 482834 516216
rect 482890 516160 482895 516216
rect 481652 516158 482895 516160
rect 481652 516156 481658 516158
rect 482829 516155 482895 516158
rect 483246 516158 487000 516218
rect 483246 516082 483306 516158
rect 486200 516128 487000 516158
rect 477358 516064 483306 516082
rect 476940 516022 483306 516064
rect 476940 516004 477418 516022
rect 485998 515810 486004 515812
rect 477358 515792 486004 515810
rect 476940 515750 486004 515792
rect 476940 515732 477418 515750
rect 485998 515748 486004 515750
rect 486068 515748 486074 515812
rect 484894 515674 484900 515676
rect 480210 515614 484900 515674
rect 480210 515538 480270 515614
rect 484894 515612 484900 515614
rect 484964 515612 484970 515676
rect 477358 515520 480270 515538
rect 476940 515478 480270 515520
rect 476940 515460 477418 515478
rect 483422 515476 483428 515540
rect 483492 515538 483498 515540
rect 486200 515538 487000 515568
rect 483492 515478 487000 515538
rect 483492 515476 483498 515478
rect 486200 515448 487000 515478
rect 480662 515266 480668 515268
rect 477358 515248 480668 515266
rect 476940 515206 480668 515248
rect 476940 515188 477418 515206
rect 480662 515204 480668 515206
rect 480732 515204 480738 515268
rect 483790 515130 483796 515132
rect 480210 515070 483796 515130
rect 480210 514994 480270 515070
rect 483790 515068 483796 515070
rect 483860 515068 483866 515132
rect 477358 514976 480270 514994
rect 476940 514934 480270 514976
rect 476940 514916 477418 514934
rect 483238 514932 483244 514996
rect 483308 514994 483314 514996
rect 484301 514994 484367 514997
rect 483308 514992 484367 514994
rect 483308 514936 484306 514992
rect 484362 514936 484367 514992
rect 483308 514934 484367 514936
rect 483308 514932 483314 514934
rect 484301 514931 484367 514934
rect 480478 514796 480484 514860
rect 480548 514858 480554 514860
rect 481449 514858 481515 514861
rect 486200 514858 487000 514888
rect 480548 514856 481515 514858
rect 480548 514800 481454 514856
rect 481510 514800 481515 514856
rect 480548 514798 481515 514800
rect 480548 514796 480554 514798
rect 481449 514795 481515 514798
rect 482878 514798 487000 514858
rect 482878 514722 482938 514798
rect 486200 514768 487000 514798
rect 477358 514704 482938 514722
rect 476940 514662 482938 514704
rect 476940 514644 477418 514662
rect 479742 514450 479748 514452
rect 477358 514432 479748 514450
rect 476940 514390 479748 514432
rect 476940 514372 477418 514390
rect 479742 514388 479748 514390
rect 479812 514388 479818 514452
rect 483422 514178 483428 514180
rect 477358 514160 483428 514178
rect 476940 514118 483428 514160
rect 476940 514100 477418 514118
rect 483422 514116 483428 514118
rect 483492 514116 483498 514180
rect 484342 514116 484348 514180
rect 484412 514178 484418 514180
rect 486200 514178 487000 514208
rect 484412 514118 487000 514178
rect 484412 514116 484418 514118
rect 486200 514088 487000 514118
rect 485814 513906 485820 513908
rect 477358 513888 485820 513906
rect 476940 513846 485820 513888
rect 476940 513828 477418 513846
rect 485814 513844 485820 513846
rect 485884 513844 485890 513908
rect 481766 513708 481772 513772
rect 481836 513770 481842 513772
rect 482921 513770 482987 513773
rect 481836 513768 482987 513770
rect 481836 513712 482926 513768
rect 482982 513712 482987 513768
rect 481836 513710 482987 513712
rect 481836 513708 481842 513710
rect 482921 513707 482987 513710
rect 485078 513634 485084 513636
rect 477358 513616 485084 513634
rect 476940 513574 485084 513616
rect 476940 513556 477418 513574
rect 485078 513572 485084 513574
rect 485148 513572 485154 513636
rect 484526 513436 484532 513500
rect 484596 513498 484602 513500
rect 486200 513498 487000 513528
rect 484596 513438 487000 513498
rect 484596 513436 484602 513438
rect 486200 513408 487000 513438
rect 477534 513300 477540 513364
rect 477604 513362 477610 513364
rect 478689 513362 478755 513365
rect 477604 513360 478755 513362
rect 477604 513304 478694 513360
rect 478750 513304 478755 513360
rect 477604 513302 478755 513304
rect 477604 513300 477610 513302
rect 478689 513299 478755 513302
rect 480662 513300 480668 513364
rect 480732 513362 480738 513364
rect 481541 513362 481607 513365
rect 480732 513360 481607 513362
rect 480732 513304 481546 513360
rect 481602 513304 481607 513360
rect 480732 513302 481607 513304
rect 480732 513300 480738 513302
rect 481541 513299 481607 513302
rect 476940 513228 477418 513288
rect 477358 513226 477418 513228
rect 479926 513226 479932 513228
rect 477358 513166 479932 513226
rect 479926 513164 479932 513166
rect 479996 513164 480002 513228
rect 479374 513090 479380 513092
rect 477174 513072 479380 513090
rect 476940 513030 479380 513072
rect 476940 513012 477234 513030
rect 479374 513028 479380 513030
rect 479444 513028 479450 513092
rect 484342 512954 484348 512956
rect 477358 512894 484348 512954
rect 477358 512800 477418 512894
rect 484342 512892 484348 512894
rect 484412 512892 484418 512956
rect 476940 512740 477418 512800
rect 478822 512756 478828 512820
rect 478892 512818 478898 512820
rect 486200 512818 487000 512848
rect 478892 512758 487000 512818
rect 478892 512756 478898 512758
rect 486200 512728 487000 512758
rect 481214 512546 481220 512548
rect 477358 512528 481220 512546
rect 476940 512486 481220 512528
rect 476940 512468 477418 512486
rect 481214 512484 481220 512486
rect 481284 512484 481290 512548
rect 485262 512274 485268 512276
rect 477358 512256 485268 512274
rect 476940 512214 485268 512256
rect 476940 512196 477418 512214
rect 485262 512212 485268 512214
rect 485332 512212 485338 512276
rect 484342 512076 484348 512140
rect 484412 512138 484418 512140
rect 486200 512138 487000 512168
rect 484412 512078 487000 512138
rect 484412 512076 484418 512078
rect 486200 512048 487000 512078
rect 481030 512002 481036 512004
rect 477358 511984 481036 512002
rect 476940 511942 481036 511984
rect 476940 511924 477418 511942
rect 481030 511940 481036 511942
rect 481100 511940 481106 512004
rect 478638 511804 478644 511868
rect 478708 511866 478714 511868
rect 478781 511866 478847 511869
rect 478708 511864 478847 511866
rect 478708 511808 478786 511864
rect 478842 511808 478847 511864
rect 478708 511806 478847 511808
rect 478708 511804 478714 511806
rect 478781 511803 478847 511806
rect 478454 511730 478460 511732
rect 477174 511712 478460 511730
rect 476940 511670 478460 511712
rect 476940 511652 477234 511670
rect 478454 511668 478460 511670
rect 478524 511668 478530 511732
rect 485630 511594 485636 511596
rect 477358 511534 485636 511594
rect 477358 511440 477418 511534
rect 485630 511532 485636 511534
rect 485700 511532 485706 511596
rect 476940 511380 477418 511440
rect 481398 511396 481404 511460
rect 481468 511458 481474 511460
rect 486200 511458 487000 511488
rect 481468 511398 487000 511458
rect 481468 511396 481474 511398
rect 486200 511368 487000 511398
rect 484342 511186 484348 511188
rect 477358 511168 484348 511186
rect 476940 511126 484348 511168
rect 476940 511108 477418 511126
rect 484342 511124 484348 511126
rect 484412 511124 484418 511188
rect 484526 510914 484532 510916
rect 477358 510896 484532 510914
rect 476940 510854 484532 510896
rect 476940 510836 477418 510854
rect 484526 510852 484532 510854
rect 484596 510852 484602 510916
rect 486200 510778 487000 510808
rect 483246 510718 487000 510778
rect 478822 510642 478828 510644
rect 476990 510624 478828 510642
rect 476940 510582 478828 510624
rect 476940 510564 477050 510582
rect 478822 510580 478828 510582
rect 478892 510580 478898 510644
rect 483246 510370 483306 510718
rect 486200 510688 487000 510718
rect 477358 510352 483306 510370
rect 476940 510310 483306 510352
rect 476940 510292 477418 510310
rect 481398 510098 481404 510100
rect 477358 510080 481404 510098
rect 476940 510038 481404 510080
rect 476940 510020 477418 510038
rect 481398 510036 481404 510038
rect 481468 510036 481474 510100
rect 486200 510098 487000 510128
rect 483246 510038 487000 510098
rect 483246 509826 483306 510038
rect 486200 510008 487000 510038
rect 477358 509808 483306 509826
rect 476940 509766 483306 509808
rect 476940 509748 477418 509766
rect 483606 509554 483612 509556
rect 477358 509536 483612 509554
rect 476940 509494 483612 509536
rect 476940 509476 477418 509494
rect 483606 509492 483612 509494
rect 483676 509492 483682 509556
rect 486200 509418 487000 509448
rect 480210 509358 487000 509418
rect 480210 509282 480270 509358
rect 486200 509328 487000 509358
rect 477358 509264 480270 509282
rect 476940 509222 480270 509264
rect 476940 509204 477418 509222
rect 478270 509010 478276 509012
rect 477358 508992 478276 509010
rect 476940 508950 478276 508992
rect 476940 508932 477418 508950
rect 478270 508948 478276 508950
rect 478340 508948 478346 509012
rect 486200 508738 487000 508768
rect 477358 508720 487000 508738
rect 476940 508678 487000 508720
rect 476940 508660 477418 508678
rect 486200 508648 487000 508678
rect 477534 508466 477540 508468
rect 477358 508448 477540 508466
rect 476940 508406 477540 508448
rect 476940 508388 477418 508406
rect 477534 508404 477540 508406
rect 477604 508404 477610 508468
rect 478086 508194 478092 508196
rect 477174 508176 478092 508194
rect 476940 508134 478092 508176
rect 0 508058 800 508088
rect 9446 508066 10032 508126
rect 476940 508116 477234 508134
rect 478086 508132 478092 508134
rect 478156 508132 478162 508196
rect 9446 508058 9506 508066
rect 486200 508058 487000 508088
rect 0 507998 9506 508058
rect 477358 507998 487000 508058
rect 0 507968 800 507998
rect 477358 507904 477418 507998
rect 486200 507968 487000 507998
rect 476940 507844 477418 507904
rect 478638 507650 478644 507652
rect 477358 507632 478644 507650
rect 476940 507590 478644 507632
rect 476940 507572 477418 507590
rect 478638 507588 478644 507590
rect 478708 507588 478714 507652
rect 0 507378 800 507408
rect 486200 507378 487000 507408
rect 0 507360 9506 507378
rect 477358 507360 487000 507378
rect 0 507318 10060 507360
rect 0 507288 800 507318
rect 9446 507300 10060 507318
rect 476940 507318 487000 507360
rect 476940 507300 477418 507318
rect 486200 507288 487000 507318
rect 482134 507106 482140 507108
rect 477358 507088 482140 507106
rect 476940 507046 482140 507088
rect 476940 507028 477418 507046
rect 482134 507044 482140 507046
rect 482204 507044 482210 507108
rect 483054 506834 483060 506836
rect 477358 506816 483060 506834
rect 476940 506774 483060 506816
rect 476940 506756 477418 506774
rect 483054 506772 483060 506774
rect 483124 506772 483130 506836
rect 0 506698 800 506728
rect 486200 506698 487000 506728
rect 0 506638 9506 506698
rect 0 506608 800 506638
rect 9446 506544 9506 506638
rect 480210 506638 487000 506698
rect 480210 506562 480270 506638
rect 486200 506608 487000 506638
rect 477358 506544 480270 506562
rect 9446 506484 10060 506544
rect 476940 506502 480270 506544
rect 476940 506484 477418 506502
rect 480846 506290 480852 506292
rect 477358 506272 480852 506290
rect 476940 506230 480852 506272
rect 476940 506212 477418 506230
rect 480846 506228 480852 506230
rect 480916 506228 480922 506292
rect 0 506018 800 506048
rect 486200 506018 487000 506048
rect 0 505958 9506 506018
rect 477358 506000 487000 506018
rect 0 505928 800 505958
rect 9446 505728 9506 505958
rect 476940 505958 487000 506000
rect 476940 505940 477418 505958
rect 486200 505928 487000 505958
rect 481582 505746 481588 505748
rect 477358 505728 481588 505746
rect 9446 505668 10060 505728
rect 476940 505686 481588 505728
rect 476940 505668 477418 505686
rect 481582 505684 481588 505686
rect 481652 505684 481658 505748
rect 483238 505474 483244 505476
rect 477358 505456 483244 505474
rect 476940 505414 483244 505456
rect 476940 505396 477418 505414
rect 483238 505412 483244 505414
rect 483308 505412 483314 505476
rect 486200 505338 487000 505368
rect 480210 505278 487000 505338
rect 480210 505202 480270 505278
rect 486200 505248 487000 505278
rect 477358 505184 480270 505202
rect 476940 505142 480270 505184
rect 476940 505124 477418 505142
rect 480478 504930 480484 504932
rect 477358 504912 480484 504930
rect 476940 504870 480484 504912
rect 9446 504796 10060 504856
rect 476940 504852 477418 504870
rect 480478 504868 480484 504870
rect 480548 504868 480554 504932
rect 0 504658 800 504688
rect 9446 504658 9506 504796
rect 486200 504658 487000 504688
rect 0 504598 9506 504658
rect 477358 504640 487000 504658
rect 476940 504598 487000 504640
rect 0 504568 800 504598
rect 476940 504580 477418 504598
rect 486200 504568 487000 504598
rect 481766 504386 481772 504388
rect 477358 504368 481772 504386
rect 476940 504326 481772 504368
rect 476940 504308 477418 504326
rect 481766 504324 481772 504326
rect 481836 504324 481842 504388
rect 480662 504114 480668 504116
rect 477358 504096 480668 504114
rect 476940 504054 480668 504096
rect 0 503978 800 504008
rect 9446 503980 10060 504040
rect 476940 504036 477418 504054
rect 480662 504052 480668 504054
rect 480732 504052 480738 504116
rect 9446 503978 9506 503980
rect 486200 503978 487000 504008
rect 0 503918 9506 503978
rect 480210 503918 487000 503978
rect 0 503888 800 503918
rect 480210 503842 480270 503918
rect 486200 503888 487000 503918
rect 477358 503824 480270 503842
rect 476940 503782 480270 503824
rect 476940 503764 477418 503782
rect 477358 503552 483306 503570
rect 476940 503510 483306 503552
rect 476940 503492 477418 503510
rect 0 503298 800 503328
rect 483054 503298 483060 503300
rect 0 503280 9506 503298
rect 477358 503280 483060 503298
rect 0 503238 10060 503280
rect 0 503208 800 503238
rect 9446 503220 10060 503238
rect 476940 503238 483060 503280
rect 476940 503220 477418 503238
rect 483054 503236 483060 503238
rect 483124 503236 483130 503300
rect 483246 503298 483306 503510
rect 486200 503298 487000 503328
rect 483246 503238 487000 503298
rect 486200 503208 487000 503238
rect 476940 502892 477418 502952
rect 477358 502890 477418 502892
rect 481766 502890 481772 502892
rect 477358 502830 481772 502890
rect 481766 502828 481772 502830
rect 481836 502828 481842 502892
rect 0 502618 800 502648
rect 476940 502620 477418 502680
rect 477358 502618 477418 502620
rect 486200 502618 487000 502648
rect 0 502558 9506 502618
rect 477358 502558 487000 502618
rect 0 502528 800 502558
rect 9446 502464 9506 502558
rect 486200 502528 487000 502558
rect 477534 502482 477540 502484
rect 477358 502464 477540 502482
rect 9446 502404 10060 502464
rect 476940 502422 477540 502464
rect 476940 502404 477418 502422
rect 477534 502420 477540 502422
rect 477604 502420 477610 502484
rect 476940 502076 477418 502136
rect 477358 502074 477418 502076
rect 477358 502014 480270 502074
rect 0 501938 800 501968
rect 480210 501938 480270 502014
rect 486200 501938 487000 501968
rect 0 501878 9506 501938
rect 480210 501878 487000 501938
rect 0 501848 800 501878
rect 9446 501648 9506 501878
rect 476940 501804 477418 501864
rect 486200 501848 487000 501878
rect 477358 501802 477418 501804
rect 480662 501802 480668 501804
rect 477358 501742 480668 501802
rect 480662 501740 480668 501742
rect 480732 501740 480738 501804
rect 483422 501666 483428 501668
rect 477358 501648 483428 501666
rect 9446 501588 10060 501648
rect 476940 501606 483428 501648
rect 476940 501588 477418 501606
rect 483422 501604 483428 501606
rect 483492 501604 483498 501668
rect 476940 501260 477418 501320
rect 477358 501258 477418 501260
rect 486200 501258 487000 501288
rect 477358 501198 487000 501258
rect 486200 501168 487000 501198
rect 476940 500988 477418 501048
rect 477358 500986 477418 500988
rect 481582 500986 481588 500988
rect 477358 500926 481588 500986
rect 481582 500924 481588 500926
rect 481652 500924 481658 500988
rect 9446 500716 10060 500776
rect 476940 500716 477418 500776
rect 0 500578 800 500608
rect 9446 500578 9506 500716
rect 477358 500714 477418 500716
rect 477358 500654 480270 500714
rect 0 500518 9506 500578
rect 480210 500578 480270 500654
rect 486200 500578 487000 500608
rect 480210 500518 487000 500578
rect 0 500488 800 500518
rect 476940 500444 477418 500504
rect 486200 500488 487000 500518
rect 477358 500442 477418 500444
rect 480846 500442 480852 500444
rect 477358 500382 480852 500442
rect 480846 500380 480852 500382
rect 480916 500380 480922 500444
rect 483606 500306 483612 500308
rect 477358 500288 483612 500306
rect 476940 500246 483612 500288
rect 476940 500228 477418 500246
rect 483606 500244 483612 500246
rect 483676 500244 483682 500308
rect 0 499898 800 499928
rect 9446 499900 10060 499960
rect 476940 499900 477418 499960
rect 9446 499898 9506 499900
rect 0 499838 9506 499898
rect 477358 499898 477418 499900
rect 486200 499898 487000 499928
rect 477358 499838 487000 499898
rect 0 499808 800 499838
rect 486200 499808 487000 499838
rect 476940 499628 477418 499688
rect 477358 499626 477418 499628
rect 482134 499626 482140 499628
rect 477358 499566 482140 499626
rect 482134 499564 482140 499566
rect 482204 499564 482210 499628
rect 476940 499356 477418 499416
rect 477358 499354 477418 499356
rect 477358 499294 480270 499354
rect 0 499218 800 499248
rect 480210 499218 480270 499294
rect 486200 499218 487000 499248
rect 0 499200 9506 499218
rect 0 499158 10060 499200
rect 480210 499158 487000 499218
rect 0 499128 800 499158
rect 9446 499140 10060 499158
rect 476940 499084 477418 499144
rect 486200 499128 487000 499158
rect 477358 499082 477418 499084
rect 481030 499082 481036 499084
rect 477358 499022 481036 499082
rect 481030 499020 481036 499022
rect 481100 499020 481106 499084
rect 483790 498946 483796 498948
rect 477358 498928 483796 498946
rect 476940 498886 483796 498928
rect 476940 498868 477418 498886
rect 483790 498884 483796 498886
rect 483860 498884 483866 498948
rect 0 498538 800 498568
rect 476940 498540 477418 498600
rect 477358 498538 477418 498540
rect 486200 498538 487000 498568
rect 0 498478 9506 498538
rect 477358 498478 487000 498538
rect 0 498448 800 498478
rect 9446 498384 9506 498478
rect 486200 498448 487000 498478
rect 9446 498324 10060 498384
rect 476940 498268 477418 498328
rect 477358 498266 477418 498268
rect 482318 498266 482324 498268
rect 477358 498206 482324 498266
rect 482318 498204 482324 498206
rect 482388 498204 482394 498268
rect 476940 497996 477418 498056
rect 477358 497994 477418 497996
rect 477358 497934 480270 497994
rect 0 497858 800 497888
rect 480210 497858 480270 497934
rect 486200 497858 487000 497888
rect 0 497798 9506 497858
rect 480210 497798 487000 497858
rect 0 497768 800 497798
rect 9446 497568 9506 497798
rect 476940 497724 477418 497784
rect 486200 497768 487000 497798
rect 477358 497722 477418 497724
rect 481214 497722 481220 497724
rect 477358 497662 481220 497722
rect 481214 497660 481220 497662
rect 481284 497660 481290 497724
rect 9446 497508 10060 497568
rect 476940 497452 477418 497512
rect 477358 497450 477418 497452
rect 480294 497450 480300 497452
rect 477358 497390 480300 497450
rect 480294 497388 480300 497390
rect 480364 497388 480370 497452
rect 476940 497180 477418 497240
rect 477358 497178 477418 497180
rect 486200 497178 487000 497208
rect 477358 497118 487000 497178
rect 486200 497088 487000 497118
rect 476940 496908 477418 496968
rect 477358 496906 477418 496908
rect 480110 496906 480116 496908
rect 477358 496846 480116 496906
rect 480110 496844 480116 496846
rect 480180 496844 480186 496908
rect 480662 496844 480668 496908
rect 480732 496906 480738 496908
rect 481541 496906 481607 496909
rect 480732 496904 481607 496906
rect 480732 496848 481546 496904
rect 481602 496848 481607 496904
rect 480732 496846 481607 496848
rect 480732 496844 480738 496846
rect 481541 496843 481607 496846
rect 9446 496636 10060 496696
rect 476940 496636 477418 496696
rect 0 496498 800 496528
rect 9446 496498 9506 496636
rect 0 496438 9506 496498
rect 477358 496498 477418 496636
rect 486200 496498 487000 496528
rect 477358 496438 487000 496498
rect 0 496408 800 496438
rect 476940 496364 477234 496424
rect 486200 496408 487000 496438
rect 477174 496362 477234 496364
rect 479558 496362 479564 496364
rect 477174 496302 479564 496362
rect 479558 496300 479564 496302
rect 479628 496300 479634 496364
rect 486417 496226 486483 496229
rect 477358 496224 486483 496226
rect 477358 496208 486422 496224
rect 476940 496168 486422 496208
rect 486478 496168 486483 496224
rect 476940 496166 486483 496168
rect 476940 496148 477418 496166
rect 486417 496163 486483 496166
rect 0 495818 800 495848
rect 9446 495820 10060 495880
rect 476940 495820 477418 495880
rect 9446 495818 9506 495820
rect 0 495758 9506 495818
rect 477358 495818 477418 495820
rect 486200 495818 487000 495848
rect 477358 495758 487000 495818
rect 0 495728 800 495758
rect 486200 495728 487000 495758
rect 476940 495548 477418 495608
rect 477358 495546 477418 495548
rect 478086 495546 478092 495548
rect 477358 495486 478092 495546
rect 478086 495484 478092 495486
rect 478156 495484 478162 495548
rect 476940 495276 477418 495336
rect 0 495138 800 495168
rect 477358 495138 477418 495276
rect 486200 495138 487000 495168
rect 0 495120 9506 495138
rect 0 495078 10060 495120
rect 477358 495078 487000 495138
rect 0 495048 800 495078
rect 9446 495060 10060 495078
rect 476940 495004 477234 495064
rect 486200 495048 487000 495078
rect 477174 495002 477234 495004
rect 478270 495002 478276 495004
rect 477174 494942 478276 495002
rect 478270 494940 478276 494942
rect 478340 494940 478346 495004
rect 485998 494866 486004 494868
rect 477358 494848 486004 494866
rect 476940 494806 486004 494848
rect 476940 494788 477418 494806
rect 485998 494804 486004 494806
rect 486068 494804 486074 494868
rect 481766 494668 481772 494732
rect 481836 494730 481842 494732
rect 482921 494730 482987 494733
rect 481836 494728 482987 494730
rect 481836 494672 482926 494728
rect 482982 494672 482987 494728
rect 481836 494670 482987 494672
rect 481836 494668 481842 494670
rect 482921 494667 482987 494670
rect 483054 494668 483060 494732
rect 483124 494730 483130 494732
rect 484301 494730 484367 494733
rect 483124 494728 484367 494730
rect 483124 494672 484306 494728
rect 484362 494672 484367 494728
rect 483124 494670 484367 494672
rect 483124 494668 483130 494670
rect 484301 494667 484367 494670
rect 0 494458 800 494488
rect 476940 494460 477418 494520
rect 477358 494458 477418 494460
rect 486200 494458 487000 494488
rect 0 494398 9506 494458
rect 477358 494398 487000 494458
rect 0 494368 800 494398
rect 9446 494304 9506 494398
rect 486200 494368 487000 494398
rect 480161 494324 480227 494325
rect 480110 494322 480116 494324
rect 9446 494244 10060 494304
rect 480070 494262 480116 494322
rect 480180 494320 480227 494324
rect 480222 494264 480227 494320
rect 480110 494260 480116 494262
rect 480180 494260 480227 494264
rect 480161 494259 480227 494260
rect 476940 494188 477418 494248
rect 477358 494186 477418 494188
rect 486182 494186 486188 494188
rect 477358 494126 486188 494186
rect 486182 494124 486188 494126
rect 486252 494124 486258 494188
rect 483422 493988 483428 494052
rect 483492 494050 483498 494052
rect 484209 494050 484275 494053
rect 483492 494048 484275 494050
rect 483492 493992 484214 494048
rect 484270 493992 484275 494048
rect 483492 493990 484275 493992
rect 483492 493988 483498 493990
rect 484209 493987 484275 493990
rect 476940 493916 477418 493976
rect 477358 493914 477418 493916
rect 477358 493854 480270 493914
rect 0 493778 800 493808
rect 480210 493778 480270 493854
rect 486200 493778 487000 493808
rect 0 493718 9506 493778
rect 480210 493718 487000 493778
rect 0 493688 800 493718
rect 9446 493488 9506 493718
rect 476940 493644 477418 493704
rect 486200 493688 487000 493718
rect 477358 493642 477418 493644
rect 482277 493642 482343 493645
rect 477358 493640 482343 493642
rect 477358 493584 482282 493640
rect 482338 493584 482343 493640
rect 477358 493582 482343 493584
rect 482277 493579 482343 493582
rect 483974 493506 483980 493508
rect 477358 493488 483980 493506
rect 9446 493428 10060 493488
rect 476940 493446 483980 493488
rect 476940 493428 477418 493446
rect 483974 493444 483980 493446
rect 484044 493444 484050 493508
rect 476940 493100 477418 493160
rect 477358 493098 477418 493100
rect 486200 493098 487000 493128
rect 477358 493038 487000 493098
rect 486200 493008 487000 493038
rect 476940 492828 477418 492888
rect 477358 492826 477418 492828
rect 478454 492826 478460 492828
rect 477358 492766 478460 492826
rect 478454 492764 478460 492766
rect 478524 492764 478530 492828
rect 6870 492672 10058 492690
rect 6870 492630 10060 492672
rect 0 492418 800 492448
rect 6870 492418 6930 492630
rect 9998 492612 10060 492630
rect 477534 492628 477540 492692
rect 477604 492690 477610 492692
rect 478781 492690 478847 492693
rect 477604 492688 478847 492690
rect 477604 492632 478786 492688
rect 478842 492632 478847 492688
rect 477604 492630 478847 492632
rect 477604 492628 477610 492630
rect 478781 492627 478847 492630
rect 481582 492628 481588 492692
rect 481652 492690 481658 492692
rect 482829 492690 482895 492693
rect 481652 492688 482895 492690
rect 481652 492632 482834 492688
rect 482890 492632 482895 492688
rect 481652 492630 482895 492632
rect 481652 492628 481658 492630
rect 482829 492627 482895 492630
rect 476940 492556 477418 492616
rect 0 492358 6930 492418
rect 477358 492418 477418 492556
rect 486200 492418 487000 492448
rect 477358 492358 487000 492418
rect 0 492328 800 492358
rect 476940 492284 477234 492344
rect 486200 492328 487000 492358
rect 477174 492282 477234 492284
rect 478822 492282 478828 492284
rect 477174 492222 478828 492282
rect 478822 492220 478828 492222
rect 478892 492220 478898 492284
rect 476940 492012 477418 492072
rect 477358 492010 477418 492012
rect 481950 492010 481956 492012
rect 477358 491950 481956 492010
rect 481950 491948 481956 491950
rect 482020 491948 482026 492012
rect 0 491738 800 491768
rect 9446 491740 10060 491800
rect 476940 491740 477418 491800
rect 9446 491738 9506 491740
rect 0 491678 9506 491738
rect 477358 491738 477418 491740
rect 486200 491738 487000 491768
rect 477358 491678 487000 491738
rect 0 491648 800 491678
rect 486200 491648 487000 491678
rect 481766 491602 481772 491604
rect 477358 491584 481772 491602
rect 476940 491542 481772 491584
rect 476940 491524 477418 491542
rect 481766 491540 481772 491542
rect 481836 491540 481842 491604
rect 477358 491312 483306 491330
rect 476940 491270 483306 491312
rect 476940 491252 477418 491270
rect 479558 491132 479564 491196
rect 479628 491194 479634 491196
rect 480069 491194 480135 491197
rect 479628 491192 480135 491194
rect 479628 491136 480074 491192
rect 480130 491136 480135 491192
rect 479628 491134 480135 491136
rect 479628 491132 479634 491134
rect 480069 491131 480135 491134
rect 0 491058 800 491088
rect 483246 491058 483306 491270
rect 486200 491058 487000 491088
rect 0 491040 9506 491058
rect 0 490998 10060 491040
rect 483246 490998 487000 491058
rect 0 490968 800 490998
rect 9446 490980 10060 490998
rect 476940 490924 477418 490984
rect 486200 490968 487000 490998
rect 477358 490922 477418 490924
rect 484894 490922 484900 490924
rect 477358 490862 484900 490922
rect 484894 490860 484900 490862
rect 484964 490860 484970 490924
rect 484526 490786 484532 490788
rect 477358 490768 484532 490786
rect 476940 490726 484532 490768
rect 476940 490708 477418 490726
rect 484526 490724 484532 490726
rect 484596 490724 484602 490788
rect 0 490378 800 490408
rect 476940 490380 477418 490440
rect 477358 490378 477418 490380
rect 486200 490378 487000 490408
rect 0 490318 9506 490378
rect 477358 490318 487000 490378
rect 0 490288 800 490318
rect 9446 490224 9506 490318
rect 486200 490288 487000 490318
rect 9446 490164 10060 490224
rect 477350 490168 477356 490170
rect 476940 490108 477356 490168
rect 477350 490106 477356 490108
rect 477420 490106 477426 490170
rect 477358 489952 484778 489970
rect 476940 489910 484778 489952
rect 476940 489892 477418 489910
rect 0 489698 800 489728
rect 484718 489698 484778 489910
rect 486200 489698 487000 489728
rect 0 489638 9506 489698
rect 484718 489638 487000 489698
rect 0 489608 800 489638
rect 9446 489408 9506 489638
rect 476940 489564 477418 489624
rect 486200 489608 487000 489638
rect 477358 489562 477418 489564
rect 484342 489562 484348 489564
rect 477358 489502 484348 489562
rect 484342 489500 484348 489502
rect 484412 489500 484418 489564
rect 483238 489426 483244 489428
rect 477358 489408 483244 489426
rect 9446 489348 10060 489408
rect 476940 489366 483244 489408
rect 476940 489348 477418 489366
rect 483238 489364 483244 489366
rect 483308 489364 483314 489428
rect 476940 489020 477418 489080
rect 477358 489018 477418 489020
rect 486200 489018 487000 489048
rect 477358 488958 487000 489018
rect 486200 488928 487000 488958
rect 476940 488748 477418 488808
rect 477358 488746 477418 488748
rect 485446 488746 485452 488748
rect 477358 488686 485452 488746
rect 485446 488684 485452 488686
rect 485516 488684 485522 488748
rect 6870 488592 9506 488610
rect 6870 488550 10060 488592
rect 0 488338 800 488368
rect 6870 488338 6930 488550
rect 9446 488532 10060 488550
rect 480294 488548 480300 488612
rect 480364 488610 480370 488612
rect 481449 488610 481515 488613
rect 480364 488608 481515 488610
rect 480364 488552 481454 488608
rect 481510 488552 481515 488608
rect 480364 488550 481515 488552
rect 480364 488548 480370 488550
rect 481449 488547 481515 488550
rect 0 488278 6930 488338
rect 0 488248 800 488278
rect 483238 488276 483244 488340
rect 483308 488338 483314 488340
rect 486200 488338 487000 488368
rect 483308 488278 487000 488338
rect 483308 488276 483314 488278
rect 486200 488248 487000 488278
rect 0 487658 800 487688
rect 9446 487660 10060 487720
rect 9446 487658 9506 487660
rect 0 487598 9506 487658
rect 0 487568 800 487598
rect 484342 487596 484348 487660
rect 484412 487658 484418 487660
rect 486200 487658 487000 487688
rect 484412 487598 487000 487658
rect 484412 487596 484418 487598
rect 486200 487568 487000 487598
rect 0 486978 800 487008
rect 0 486960 9506 486978
rect 0 486918 10060 486960
rect 0 486888 800 486918
rect 9446 486900 10060 486918
rect 477350 486916 477356 486980
rect 477420 486978 477426 486980
rect 486200 486978 487000 487008
rect 477420 486918 487000 486978
rect 477420 486916 477426 486918
rect 486200 486888 487000 486918
rect 0 486298 800 486328
rect 0 486238 9506 486298
rect 0 486208 800 486238
rect 9446 486144 9506 486238
rect 484526 486236 484532 486300
rect 484596 486298 484602 486300
rect 486200 486298 487000 486328
rect 484596 486238 487000 486298
rect 484596 486236 484602 486238
rect 486200 486208 487000 486238
rect 9446 486084 10060 486144
rect 0 485618 800 485648
rect 0 485558 9506 485618
rect 0 485528 800 485558
rect 9446 485328 9506 485558
rect 484894 485556 484900 485620
rect 484964 485618 484970 485620
rect 486200 485618 487000 485648
rect 484964 485558 487000 485618
rect 484964 485556 484970 485558
rect 486200 485528 487000 485558
rect 9446 485268 10060 485328
rect 481766 484876 481772 484940
rect 481836 484938 481842 484940
rect 486200 484938 487000 484968
rect 481836 484878 487000 484938
rect 481836 484876 481842 484878
rect 486200 484848 487000 484878
rect 6870 484512 9506 484530
rect 6870 484470 10060 484512
rect 0 484258 800 484288
rect 6870 484258 6930 484470
rect 9446 484452 10060 484470
rect 0 484198 6930 484258
rect 0 484168 800 484198
rect 481950 484196 481956 484260
rect 482020 484258 482026 484260
rect 486200 484258 487000 484288
rect 482020 484198 487000 484258
rect 482020 484196 482026 484198
rect 486200 484168 487000 484198
rect 0 483578 800 483608
rect 9446 483580 10060 483640
rect 9446 483578 9506 483580
rect 0 483518 9506 483578
rect 0 483488 800 483518
rect 478822 483516 478828 483580
rect 478892 483578 478898 483580
rect 486200 483578 487000 483608
rect 478892 483518 487000 483578
rect 478892 483516 478898 483518
rect 486200 483488 487000 483518
rect 0 482898 800 482928
rect 0 482880 9506 482898
rect 0 482838 10060 482880
rect 0 482808 800 482838
rect 9446 482820 10060 482838
rect 478454 482836 478460 482900
rect 478524 482898 478530 482900
rect 486200 482898 487000 482928
rect 478524 482838 487000 482898
rect 478524 482836 478530 482838
rect 486200 482808 487000 482838
rect 0 482218 800 482248
rect 0 482158 9506 482218
rect 0 482128 800 482158
rect 9446 482064 9506 482158
rect 483974 482156 483980 482220
rect 484044 482218 484050 482220
rect 486200 482218 487000 482248
rect 484044 482158 487000 482218
rect 484044 482156 484050 482158
rect 486200 482128 487000 482158
rect 9446 482004 10060 482064
rect 0 481538 800 481568
rect 482277 481538 482343 481541
rect 486200 481538 487000 481568
rect 0 481478 9506 481538
rect 0 481448 800 481478
rect 9446 481248 9506 481478
rect 482277 481536 487000 481538
rect 482277 481480 482282 481536
rect 482338 481480 487000 481536
rect 482277 481478 487000 481480
rect 482277 481475 482343 481478
rect 486200 481448 487000 481478
rect 9446 481188 10060 481248
rect 486200 480860 487000 480888
rect 486200 480796 486372 480860
rect 486436 480796 487000 480860
rect 486200 480768 487000 480796
rect 9446 480316 10060 480376
rect 9446 480314 9506 480316
rect 5582 480254 9506 480314
rect 0 480178 800 480208
rect 5582 480178 5642 480254
rect 0 480118 5642 480178
rect 0 480088 800 480118
rect 485998 480116 486004 480180
rect 486068 480178 486074 480180
rect 486200 480178 487000 480208
rect 486068 480118 487000 480178
rect 486068 480116 486074 480118
rect 486200 480088 487000 480118
rect 0 479498 800 479528
rect 9446 479500 10060 479560
rect 9446 479498 9506 479500
rect 0 479438 9506 479498
rect 0 479408 800 479438
rect 478270 479436 478276 479500
rect 478340 479498 478346 479500
rect 486200 479498 487000 479528
rect 478340 479438 487000 479498
rect 478340 479436 478346 479438
rect 486200 479408 487000 479438
rect 0 478818 800 478848
rect 0 478800 9506 478818
rect 0 478758 10060 478800
rect 0 478728 800 478758
rect 9446 478740 10060 478758
rect 478086 478756 478092 478820
rect 478156 478818 478162 478820
rect 486200 478818 487000 478848
rect 478156 478758 487000 478818
rect 478156 478756 478162 478758
rect 486200 478728 487000 478758
rect 0 478138 800 478168
rect 486200 478141 487000 478168
rect 0 478078 9506 478138
rect 0 478048 800 478078
rect 9446 477984 9506 478078
rect 486141 478136 487000 478141
rect 486141 478080 486146 478136
rect 486202 478080 487000 478136
rect 486141 478075 487000 478080
rect 486200 478048 487000 478075
rect 9446 477924 10060 477984
rect 0 477458 800 477488
rect 480069 477458 480135 477461
rect 486200 477458 487000 477488
rect 0 477398 9506 477458
rect 0 477368 800 477398
rect 9446 477168 9506 477398
rect 480069 477456 487000 477458
rect 480069 477400 480074 477456
rect 480130 477400 487000 477456
rect 480069 477398 487000 477400
rect 480069 477395 480135 477398
rect 486200 477368 487000 477398
rect 9446 477108 10060 477168
rect 480161 476778 480227 476781
rect 486200 476778 487000 476808
rect 480161 476776 487000 476778
rect 480161 476720 480166 476776
rect 480222 476720 487000 476776
rect 480161 476718 487000 476720
rect 480161 476715 480227 476718
rect 486200 476688 487000 476718
rect 9446 476236 10060 476296
rect 9446 476234 9506 476236
rect 6870 476174 9506 476234
rect 0 476098 800 476128
rect 6870 476098 6930 476174
rect 0 476038 6930 476098
rect 0 476008 800 476038
rect 485446 476036 485452 476100
rect 485516 476098 485522 476100
rect 486200 476098 487000 476128
rect 485516 476038 487000 476098
rect 485516 476036 485522 476038
rect 486200 476008 487000 476038
rect 0 475418 800 475448
rect 9446 475420 10060 475480
rect 9446 475418 9506 475420
rect 0 475358 9506 475418
rect 0 475328 800 475358
rect 481214 475356 481220 475420
rect 481284 475418 481290 475420
rect 486200 475418 487000 475448
rect 481284 475358 487000 475418
rect 481284 475356 481290 475358
rect 486200 475328 487000 475358
rect 0 474738 800 474768
rect 0 474720 9506 474738
rect 0 474678 10060 474720
rect 0 474648 800 474678
rect 9446 474660 10060 474678
rect 482318 474676 482324 474740
rect 482388 474738 482394 474740
rect 486200 474738 487000 474768
rect 482388 474678 487000 474738
rect 482388 474676 482394 474678
rect 486200 474648 487000 474678
rect 0 474058 800 474088
rect 0 473998 9506 474058
rect 0 473968 800 473998
rect 9446 473904 9506 473998
rect 483790 473996 483796 474060
rect 483860 474058 483866 474060
rect 486200 474058 487000 474088
rect 483860 473998 487000 474058
rect 483860 473996 483866 473998
rect 486200 473968 487000 473998
rect 9446 473844 10060 473904
rect 0 473378 800 473408
rect 0 473318 4170 473378
rect 0 473288 800 473318
rect 4110 473242 4170 473318
rect 481030 473316 481036 473380
rect 481100 473378 481106 473380
rect 486200 473378 487000 473408
rect 481100 473318 487000 473378
rect 481100 473316 481106 473318
rect 486200 473288 487000 473318
rect 4110 473182 9506 473242
rect 9446 473088 9506 473182
rect 9446 473028 10060 473088
rect 482134 472636 482140 472700
rect 482204 472698 482210 472700
rect 486200 472698 487000 472728
rect 482204 472638 487000 472698
rect 482204 472636 482210 472638
rect 486200 472608 487000 472638
rect 9446 472156 10060 472216
rect 0 472018 800 472048
rect 9446 472018 9506 472156
rect 0 471958 9506 472018
rect 0 471928 800 471958
rect 483606 471956 483612 472020
rect 483676 472018 483682 472020
rect 486200 472018 487000 472048
rect 483676 471958 487000 472018
rect 483676 471956 483682 471958
rect 486200 471928 487000 471958
rect 0 471338 800 471368
rect 9446 471340 10060 471400
rect 9446 471338 9506 471340
rect 0 471278 9506 471338
rect 0 471248 800 471278
rect 480846 471276 480852 471340
rect 480916 471338 480922 471340
rect 486200 471338 487000 471368
rect 480916 471278 487000 471338
rect 480916 471276 480922 471278
rect 486200 471248 487000 471278
rect 482829 470658 482895 470661
rect 486200 470658 487000 470688
rect 482829 470656 487000 470658
rect 482829 470600 482834 470656
rect 482890 470600 487000 470656
rect 482829 470598 487000 470600
rect 482829 470595 482895 470598
rect 486200 470568 487000 470598
rect 484209 469978 484275 469981
rect 486200 469978 487000 470008
rect 484209 469976 487000 469978
rect 484209 469920 484214 469976
rect 484270 469920 487000 469976
rect 484209 469918 487000 469920
rect 484209 469915 484275 469918
rect 486200 469888 487000 469918
rect 481541 469298 481607 469301
rect 486200 469298 487000 469328
rect 481541 469296 487000 469298
rect 481541 469240 481546 469296
rect 481602 469240 487000 469296
rect 481541 469238 487000 469240
rect 481541 469235 481607 469238
rect 486200 469208 487000 469238
rect 478781 468618 478847 468621
rect 486200 468618 487000 468648
rect 478781 468616 487000 468618
rect 478781 468560 478786 468616
rect 478842 468560 487000 468616
rect 478781 468558 487000 468560
rect 478781 468555 478847 468558
rect 486200 468528 487000 468558
rect 482921 467938 482987 467941
rect 486200 467938 487000 467968
rect 482921 467936 487000 467938
rect 482921 467880 482926 467936
rect 482982 467880 487000 467936
rect 482921 467878 487000 467880
rect 482921 467875 482987 467878
rect 486200 467848 487000 467878
rect 484301 467258 484367 467261
rect 486200 467258 487000 467288
rect 484301 467256 487000 467258
rect 484301 467200 484306 467256
rect 484362 467200 487000 467256
rect 484301 467198 487000 467200
rect 484301 467195 484367 467198
rect 486200 467168 487000 467198
rect 481449 466578 481515 466581
rect 486200 466578 487000 466608
rect 481449 466576 487000 466578
rect 481449 466520 481454 466576
rect 481510 466520 487000 466576
rect 481449 466518 487000 466520
rect 481449 466515 481515 466518
rect 486200 466488 487000 466518
rect 0 463178 800 463208
rect 0 463118 10032 463178
rect 0 463088 800 463118
rect 0 462498 800 462528
rect 0 462438 6930 462498
rect 0 462408 800 462438
rect 6870 462362 6930 462438
rect 6870 462302 10032 462362
rect 0 461818 800 461848
rect 0 461758 6930 461818
rect 0 461728 800 461758
rect 6870 461546 6930 461758
rect 6870 461486 10032 461546
rect 9446 460602 10060 460662
rect 0 460458 800 460488
rect 9446 460458 9506 460602
rect 0 460398 9506 460458
rect 0 460368 800 460398
rect 0 459778 800 459808
rect 9446 459786 10060 459846
rect 9446 459778 9506 459786
rect 0 459718 9506 459778
rect 482921 459778 482987 459781
rect 486200 459778 487000 459808
rect 482921 459776 487000 459778
rect 482921 459720 482926 459776
rect 482982 459720 487000 459776
rect 482921 459718 487000 459720
rect 0 459688 800 459718
rect 482921 459715 482987 459718
rect 486200 459688 487000 459718
rect 0 459098 800 459128
rect 479517 459098 479583 459101
rect 486200 459098 487000 459128
rect 0 459038 10032 459098
rect 479517 459096 487000 459098
rect 479517 459040 479522 459096
rect 479578 459040 487000 459096
rect 479517 459038 487000 459040
rect 0 459008 800 459038
rect 479517 459035 479583 459038
rect 486200 459008 487000 459038
rect 0 458418 800 458448
rect 484301 458418 484367 458421
rect 486200 458418 487000 458448
rect 0 458358 6930 458418
rect 0 458328 800 458358
rect 6870 458282 6930 458358
rect 484301 458416 487000 458418
rect 484301 458360 484306 458416
rect 484362 458360 487000 458416
rect 484301 458358 487000 458360
rect 484301 458355 484367 458358
rect 486200 458328 487000 458358
rect 6870 458222 10032 458282
rect 0 457738 800 457768
rect 482829 457738 482895 457741
rect 486200 457738 487000 457768
rect 0 457678 6930 457738
rect 0 457648 800 457678
rect 6870 457466 6930 457678
rect 482829 457736 487000 457738
rect 482829 457680 482834 457736
rect 482890 457680 487000 457736
rect 482829 457678 487000 457680
rect 482829 457675 482895 457678
rect 486200 457648 487000 457678
rect 6870 457406 10032 457466
rect 484209 457058 484275 457061
rect 486200 457058 487000 457088
rect 484209 457056 487000 457058
rect 484209 457000 484214 457056
rect 484270 457000 487000 457056
rect 484209 456998 487000 457000
rect 484209 456995 484275 456998
rect 486200 456968 487000 456998
rect 9446 456522 10060 456582
rect 0 456378 800 456408
rect 9446 456378 9506 456522
rect 0 456318 9506 456378
rect 482737 456378 482803 456381
rect 486200 456378 487000 456408
rect 482737 456376 487000 456378
rect 482737 456320 482742 456376
rect 482798 456320 487000 456376
rect 482737 456318 487000 456320
rect 0 456288 800 456318
rect 482737 456315 482803 456318
rect 486200 456288 487000 456318
rect 0 455698 800 455728
rect 9446 455706 10060 455766
rect 9446 455698 9506 455706
rect 0 455638 9506 455698
rect 484117 455698 484183 455701
rect 486200 455698 487000 455728
rect 484117 455696 487000 455698
rect 484117 455640 484122 455696
rect 484178 455640 487000 455696
rect 484117 455638 487000 455640
rect 0 455608 800 455638
rect 484117 455635 484183 455638
rect 486200 455608 487000 455638
rect 0 455018 800 455048
rect 478781 455018 478847 455021
rect 486200 455018 487000 455048
rect 0 454958 10032 455018
rect 478781 455016 487000 455018
rect 478781 454960 478786 455016
rect 478842 454960 487000 455016
rect 478781 454958 487000 454960
rect 0 454928 800 454958
rect 478781 454955 478847 454958
rect 486200 454928 487000 454958
rect 0 454338 800 454368
rect 478689 454338 478755 454341
rect 486200 454338 487000 454368
rect 0 454278 6930 454338
rect 0 454248 800 454278
rect 6870 454202 6930 454278
rect 478689 454336 487000 454338
rect 478689 454280 478694 454336
rect 478750 454280 487000 454336
rect 478689 454278 487000 454280
rect 478689 454275 478755 454278
rect 486200 454248 487000 454278
rect 6870 454142 10032 454202
rect 0 453658 800 453688
rect 480897 453658 480963 453661
rect 486200 453658 487000 453688
rect 0 453598 6930 453658
rect 0 453568 800 453598
rect 6870 453386 6930 453598
rect 480897 453656 487000 453658
rect 480897 453600 480902 453656
rect 480958 453600 487000 453656
rect 480897 453598 487000 453600
rect 480897 453595 480963 453598
rect 486200 453568 487000 453598
rect 6870 453326 10032 453386
rect 483606 452916 483612 452980
rect 483676 452978 483682 452980
rect 486200 452978 487000 453008
rect 483676 452918 487000 452978
rect 483676 452916 483682 452918
rect 486200 452888 487000 452918
rect 9446 452442 10060 452502
rect 0 452298 800 452328
rect 9446 452298 9506 452442
rect 0 452238 9506 452298
rect 481541 452298 481607 452301
rect 486200 452298 487000 452328
rect 481541 452296 487000 452298
rect 481541 452240 481546 452296
rect 481602 452240 487000 452296
rect 481541 452238 487000 452240
rect 0 452208 800 452238
rect 481541 452235 481607 452238
rect 486200 452208 487000 452238
rect 0 451618 800 451648
rect 9446 451626 10060 451686
rect 9446 451618 9506 451626
rect 0 451558 9506 451618
rect 481449 451618 481515 451621
rect 486200 451618 487000 451648
rect 481449 451616 487000 451618
rect 481449 451560 481454 451616
rect 481510 451560 487000 451616
rect 481449 451558 487000 451560
rect 0 451528 800 451558
rect 481449 451555 481515 451558
rect 486200 451528 487000 451558
rect 0 450938 800 450968
rect 478505 450938 478571 450941
rect 486200 450938 487000 450968
rect 0 450878 10032 450938
rect 478505 450936 487000 450938
rect 478505 450880 478510 450936
rect 478566 450880 487000 450936
rect 478505 450878 487000 450880
rect 0 450848 800 450878
rect 478505 450875 478571 450878
rect 486200 450848 487000 450878
rect 0 450258 800 450288
rect 478597 450258 478663 450261
rect 486200 450258 487000 450288
rect 0 450198 6930 450258
rect 0 450168 800 450198
rect 6870 450122 6930 450198
rect 478597 450256 487000 450258
rect 478597 450200 478602 450256
rect 478658 450200 487000 450256
rect 478597 450198 487000 450200
rect 478597 450195 478663 450198
rect 486200 450168 487000 450198
rect 6870 450062 10032 450122
rect 0 449578 800 449608
rect 478413 449578 478479 449581
rect 486200 449578 487000 449608
rect 0 449518 6930 449578
rect 0 449488 800 449518
rect 6870 449306 6930 449518
rect 478413 449576 487000 449578
rect 478413 449520 478418 449576
rect 478474 449520 487000 449576
rect 478413 449518 487000 449520
rect 478413 449515 478479 449518
rect 486200 449488 487000 449518
rect 6870 449246 10032 449306
rect 482645 448898 482711 448901
rect 486200 448898 487000 448928
rect 482645 448896 487000 448898
rect 482645 448840 482650 448896
rect 482706 448840 487000 448896
rect 482645 448838 487000 448840
rect 482645 448835 482711 448838
rect 486200 448808 487000 448838
rect 9446 448362 10060 448422
rect 0 448218 800 448248
rect 9446 448218 9506 448362
rect 0 448158 9506 448218
rect 484025 448218 484091 448221
rect 486200 448218 487000 448248
rect 484025 448216 487000 448218
rect 484025 448160 484030 448216
rect 484086 448160 487000 448216
rect 484025 448158 487000 448160
rect 0 448128 800 448158
rect 484025 448155 484091 448158
rect 486200 448128 487000 448158
rect 0 447538 800 447568
rect 9446 447546 10060 447606
rect 9446 447538 9506 447546
rect 0 447478 9506 447538
rect 0 447448 800 447478
rect 478086 447476 478092 447540
rect 478156 447538 478162 447540
rect 486200 447538 487000 447568
rect 478156 447478 487000 447538
rect 478156 447476 478162 447478
rect 486200 447448 487000 447478
rect 0 446858 800 446888
rect 486200 446861 487000 446888
rect 0 446798 10032 446858
rect 486141 446856 487000 446861
rect 486141 446800 486146 446856
rect 486202 446800 487000 446856
rect 0 446768 800 446798
rect 486141 446795 487000 446800
rect 486200 446768 487000 446795
rect 0 446178 800 446208
rect 480161 446178 480227 446181
rect 486200 446178 487000 446208
rect 0 446118 6930 446178
rect 0 446088 800 446118
rect 6870 446042 6930 446118
rect 480161 446176 487000 446178
rect 480161 446120 480166 446176
rect 480222 446120 487000 446176
rect 480161 446118 487000 446120
rect 480161 446115 480227 446118
rect 486200 446088 487000 446118
rect 6870 445982 10032 446042
rect 0 445498 800 445528
rect 479977 445498 480043 445501
rect 486200 445498 487000 445528
rect 0 445438 6930 445498
rect 0 445408 800 445438
rect 6870 445226 6930 445438
rect 479977 445496 487000 445498
rect 479977 445440 479982 445496
rect 480038 445440 487000 445496
rect 479977 445438 487000 445440
rect 479977 445435 480043 445438
rect 486200 445408 487000 445438
rect 6870 445166 10032 445226
rect 480069 444818 480135 444821
rect 486200 444818 487000 444848
rect 480069 444816 487000 444818
rect 480069 444760 480074 444816
rect 480130 444760 487000 444816
rect 480069 444758 487000 444760
rect 480069 444755 480135 444758
rect 486200 444728 487000 444758
rect 6870 444350 10032 444410
rect 0 444138 800 444168
rect 6870 444138 6930 444350
rect 0 444078 6930 444138
rect 479885 444138 479951 444141
rect 486200 444138 487000 444168
rect 479885 444136 487000 444138
rect 479885 444080 479890 444136
rect 479946 444080 487000 444136
rect 479885 444078 487000 444080
rect 0 444048 800 444078
rect 479885 444075 479951 444078
rect 486200 444048 487000 444078
rect 0 443458 800 443488
rect 9446 443466 10060 443526
rect 9446 443458 9506 443466
rect 0 443398 9506 443458
rect 0 443368 800 443398
rect 479374 443396 479380 443460
rect 479444 443458 479450 443460
rect 486200 443458 487000 443488
rect 479444 443398 487000 443458
rect 479444 443396 479450 443398
rect 486200 443368 487000 443398
rect 0 442778 800 442808
rect 0 442718 10032 442778
rect 0 442688 800 442718
rect 479558 442716 479564 442780
rect 479628 442778 479634 442780
rect 486200 442778 487000 442808
rect 479628 442718 487000 442778
rect 479628 442716 479634 442718
rect 486200 442688 487000 442718
rect 0 442098 800 442128
rect 0 442038 6930 442098
rect 0 442008 800 442038
rect 6870 441962 6930 442038
rect 478270 442036 478276 442100
rect 478340 442098 478346 442100
rect 486200 442098 487000 442128
rect 478340 442038 487000 442098
rect 478340 442036 478346 442038
rect 486200 442008 487000 442038
rect 6870 441902 10032 441962
rect 0 441418 800 441448
rect 0 441358 6930 441418
rect 0 441328 800 441358
rect 6870 441146 6930 441358
rect 478638 441356 478644 441420
rect 478708 441418 478714 441420
rect 486200 441418 487000 441448
rect 478708 441358 487000 441418
rect 478708 441356 478714 441358
rect 486200 441328 487000 441358
rect 6870 441086 10032 441146
rect 482134 440676 482140 440740
rect 482204 440738 482210 440740
rect 486200 440738 487000 440768
rect 482204 440678 487000 440738
rect 482204 440676 482210 440678
rect 486200 440648 487000 440678
rect 6870 440270 10032 440330
rect 0 440058 800 440088
rect 6870 440058 6930 440270
rect 0 439998 6930 440058
rect 0 439968 800 439998
rect 480846 439996 480852 440060
rect 480916 440058 480922 440060
rect 486200 440058 487000 440088
rect 480916 439998 487000 440058
rect 480916 439996 480922 439998
rect 486200 439968 487000 439998
rect 0 439378 800 439408
rect 9446 439386 10060 439446
rect 9446 439378 9506 439386
rect 0 439318 9506 439378
rect 0 439288 800 439318
rect 485630 439316 485636 439380
rect 485700 439378 485706 439380
rect 486200 439378 487000 439408
rect 485700 439318 487000 439378
rect 485700 439316 485706 439318
rect 486200 439288 487000 439318
rect 0 438698 800 438728
rect 0 438638 10032 438698
rect 0 438608 800 438638
rect 483790 438636 483796 438700
rect 483860 438698 483866 438700
rect 486200 438698 487000 438728
rect 483860 438638 487000 438698
rect 483860 438636 483866 438638
rect 486200 438608 487000 438638
rect 0 438018 800 438048
rect 486200 438021 487000 438048
rect 0 437958 6930 438018
rect 0 437928 800 437958
rect 6870 437882 6930 437958
rect 486141 438016 487000 438021
rect 486141 437960 486146 438016
rect 486202 437960 487000 438016
rect 486141 437955 487000 437960
rect 486200 437928 487000 437955
rect 6870 437822 10032 437882
rect 0 437338 800 437368
rect 0 437278 6930 437338
rect 0 437248 800 437278
rect 6870 437066 6930 437278
rect 485262 437276 485268 437340
rect 485332 437338 485338 437340
rect 486200 437338 487000 437368
rect 485332 437278 487000 437338
rect 485332 437276 485338 437278
rect 486200 437248 487000 437278
rect 6870 437006 10032 437066
rect 486200 436660 487000 436688
rect 486200 436596 486372 436660
rect 486436 436596 487000 436660
rect 486200 436568 487000 436596
rect 9446 436122 10060 436182
rect 9446 436114 9506 436122
rect 6870 436054 9506 436114
rect 0 435978 800 436008
rect 6870 435978 6930 436054
rect 0 435918 6930 435978
rect 0 435888 800 435918
rect 485078 435916 485084 435980
rect 485148 435978 485154 435980
rect 486200 435978 487000 436008
rect 485148 435918 487000 435978
rect 485148 435916 485154 435918
rect 486200 435888 487000 435918
rect 0 435298 800 435328
rect 9446 435306 10060 435366
rect 9446 435298 9506 435306
rect 0 435238 9506 435298
rect 0 435208 800 435238
rect 485814 435236 485820 435300
rect 485884 435298 485890 435300
rect 486200 435298 487000 435328
rect 485884 435238 487000 435298
rect 485884 435236 485890 435238
rect 486200 435208 487000 435238
rect 0 434618 800 434648
rect 0 434558 10032 434618
rect 0 434528 800 434558
rect 484526 434556 484532 434620
rect 484596 434618 484602 434620
rect 486200 434618 487000 434648
rect 484596 434558 487000 434618
rect 484596 434556 484602 434558
rect 486200 434528 487000 434558
rect 0 433938 800 433968
rect 0 433878 6930 433938
rect 0 433848 800 433878
rect 6870 433802 6930 433878
rect 485998 433876 486004 433940
rect 486068 433938 486074 433940
rect 486200 433938 487000 433968
rect 486068 433878 487000 433938
rect 486068 433876 486074 433878
rect 486200 433848 487000 433878
rect 6870 433742 10032 433802
rect 0 433258 800 433288
rect 0 433198 6930 433258
rect 0 433168 800 433198
rect 6870 432986 6930 433198
rect 480110 433196 480116 433260
rect 480180 433258 480186 433260
rect 486200 433258 487000 433288
rect 480180 433198 487000 433258
rect 480180 433196 480186 433198
rect 486200 433168 487000 433198
rect 6870 432926 10032 432986
rect 477350 432516 477356 432580
rect 477420 432578 477426 432580
rect 486200 432578 487000 432608
rect 477420 432518 487000 432578
rect 477420 432516 477426 432518
rect 486200 432488 487000 432518
rect 9446 432042 10060 432102
rect 9446 432034 9506 432042
rect 5582 431974 9506 432034
rect 0 431898 800 431928
rect 5582 431898 5642 431974
rect 0 431838 5642 431898
rect 0 431808 800 431838
rect 484710 431836 484716 431900
rect 484780 431898 484786 431900
rect 486200 431898 487000 431928
rect 484780 431838 487000 431898
rect 484780 431836 484786 431838
rect 486200 431808 487000 431838
rect 0 431218 800 431248
rect 9446 431226 10060 431286
rect 9446 431218 9506 431226
rect 0 431158 9506 431218
rect 0 431128 800 431158
rect 481582 431156 481588 431220
rect 481652 431218 481658 431220
rect 486200 431218 487000 431248
rect 481652 431158 487000 431218
rect 481652 431156 481658 431158
rect 486200 431128 487000 431158
rect 0 430538 800 430568
rect 0 430478 10032 430538
rect 0 430448 800 430478
rect 483238 430476 483244 430540
rect 483308 430538 483314 430540
rect 486200 430538 487000 430568
rect 483308 430478 487000 430538
rect 483308 430476 483314 430478
rect 486200 430448 487000 430478
rect 0 429858 800 429888
rect 0 429798 6930 429858
rect 0 429768 800 429798
rect 6870 429722 6930 429798
rect 484342 429796 484348 429860
rect 484412 429858 484418 429860
rect 486200 429858 487000 429888
rect 484412 429798 487000 429858
rect 484412 429796 484418 429798
rect 486200 429768 487000 429798
rect 6870 429662 10032 429722
rect 482001 429450 482067 429453
rect 486233 429450 486299 429453
rect 482001 429448 486299 429450
rect 482001 429392 482006 429448
rect 482062 429392 486238 429448
rect 486294 429392 486299 429448
rect 482001 429390 486299 429392
rect 482001 429387 482067 429390
rect 486233 429387 486299 429390
rect 0 429178 800 429208
rect 0 429118 6930 429178
rect 0 429088 800 429118
rect 6870 428906 6930 429118
rect 483054 429116 483060 429180
rect 483124 429178 483130 429180
rect 486200 429178 487000 429208
rect 483124 429118 487000 429178
rect 483124 429116 483130 429118
rect 486200 429088 487000 429118
rect 6870 428846 10032 428906
rect 484894 428436 484900 428500
rect 484964 428498 484970 428500
rect 486200 428498 487000 428528
rect 484964 428438 487000 428498
rect 484964 428436 484970 428438
rect 486200 428408 487000 428438
rect 484526 428226 484532 428228
rect 476940 428166 484532 428226
rect 484526 428164 484532 428166
rect 484596 428164 484602 428228
rect 9446 427962 10060 428022
rect 9446 427954 9506 427962
rect 485630 427954 485636 427956
rect 6870 427894 9506 427954
rect 476940 427894 485636 427954
rect 0 427818 800 427848
rect 6870 427818 6930 427894
rect 485630 427892 485636 427894
rect 485700 427892 485706 427956
rect 486200 427818 487000 427848
rect 0 427758 6930 427818
rect 477358 427758 487000 427818
rect 0 427728 800 427758
rect 477358 427696 477418 427758
rect 486200 427728 487000 427758
rect 476928 427636 477418 427696
rect 484342 427410 484348 427412
rect 476940 427350 484348 427410
rect 484342 427348 484348 427350
rect 484412 427348 484418 427412
rect 477534 427212 477540 427276
rect 477604 427274 477610 427276
rect 478413 427274 478479 427277
rect 479885 427276 479951 427277
rect 479885 427274 479932 427276
rect 477604 427272 478479 427274
rect 477604 427216 478418 427272
rect 478474 427216 478479 427272
rect 477604 427214 478479 427216
rect 479840 427272 479932 427274
rect 479840 427216 479890 427272
rect 479840 427214 479932 427216
rect 477604 427212 477610 427214
rect 478413 427211 478479 427214
rect 479885 427212 479932 427214
rect 479996 427212 480002 427276
rect 479885 427211 479951 427212
rect 0 427138 800 427168
rect 9446 427146 10060 427206
rect 9446 427138 9506 427146
rect 486200 427138 487000 427168
rect 0 427078 9506 427138
rect 476940 427078 487000 427138
rect 0 427048 800 427078
rect 486200 427048 487000 427078
rect 483238 426866 483244 426868
rect 476940 426806 483244 426866
rect 483238 426804 483244 426806
rect 483308 426804 483314 426868
rect 481582 426594 481588 426596
rect 476940 426534 481588 426594
rect 481582 426532 481588 426534
rect 481652 426532 481658 426596
rect 0 426458 800 426488
rect 486200 426458 487000 426488
rect 0 426398 10032 426458
rect 484350 426398 487000 426458
rect 0 426368 800 426398
rect 484350 426322 484410 426398
rect 486200 426368 487000 426398
rect 476940 426262 484410 426322
rect 482001 426188 482067 426189
rect 481950 426186 481956 426188
rect 481910 426126 481956 426186
rect 482020 426184 482067 426188
rect 482062 426128 482067 426184
rect 481950 426124 481956 426126
rect 482020 426124 482067 426128
rect 482502 426124 482508 426188
rect 482572 426186 482578 426188
rect 482645 426186 482711 426189
rect 482572 426184 482711 426186
rect 482572 426128 482650 426184
rect 482706 426128 482711 426184
rect 482572 426126 482711 426128
rect 482572 426124 482578 426126
rect 482001 426123 482067 426124
rect 482645 426123 482711 426126
rect 484710 426050 484716 426052
rect 476940 425990 484716 426050
rect 484710 425988 484716 425990
rect 484780 425988 484786 426052
rect 486200 425780 487000 425808
rect 480846 425778 480852 425780
rect 476940 425718 480852 425778
rect 480846 425716 480852 425718
rect 480916 425716 480922 425780
rect 486200 425716 486372 425780
rect 486436 425716 487000 425780
rect 486200 425688 487000 425716
rect 477350 425520 477356 425522
rect 476928 425460 477356 425520
rect 477350 425458 477356 425460
rect 477420 425458 477426 425522
rect 480110 425234 480116 425236
rect 476940 425174 480116 425234
rect 480110 425172 480116 425174
rect 480180 425172 480186 425236
rect 482870 425036 482876 425100
rect 482940 425098 482946 425100
rect 486200 425098 487000 425128
rect 482940 425038 487000 425098
rect 482940 425036 482946 425038
rect 486200 425008 487000 425038
rect 483105 424962 483171 424965
rect 476940 424960 483171 424962
rect 476940 424904 483110 424960
rect 483166 424904 483171 424960
rect 476940 424902 483171 424904
rect 483105 424899 483171 424902
rect 483238 424900 483244 424964
rect 483308 424962 483314 424964
rect 484025 424962 484091 424965
rect 483308 424960 484091 424962
rect 483308 424904 484030 424960
rect 484086 424904 484091 424960
rect 483308 424902 484091 424904
rect 483308 424900 483314 424902
rect 484025 424899 484091 424902
rect 477401 424826 477467 424829
rect 486366 424826 486372 424828
rect 477401 424824 486372 424826
rect 477401 424768 477406 424824
rect 477462 424768 486372 424824
rect 477401 424766 486372 424768
rect 477401 424763 477467 424766
rect 486366 424764 486372 424766
rect 486436 424764 486442 424828
rect 483606 424690 483612 424692
rect 476940 424630 483612 424690
rect 483606 424628 483612 424630
rect 483676 424628 483682 424692
rect 479742 424492 479748 424556
rect 479812 424554 479818 424556
rect 479977 424554 480043 424557
rect 479812 424552 480043 424554
rect 479812 424496 479982 424552
rect 480038 424496 480043 424552
rect 479812 424494 480043 424496
rect 479812 424492 479818 424494
rect 479977 424491 480043 424494
rect 483105 424554 483171 424557
rect 486049 424554 486115 424557
rect 483105 424552 486115 424554
rect 483105 424496 483110 424552
rect 483166 424496 486054 424552
rect 486110 424496 486115 424552
rect 483105 424494 486115 424496
rect 483105 424491 483171 424494
rect 486049 424491 486115 424494
rect 477401 424432 477467 424435
rect 476928 424430 477467 424432
rect 476928 424374 477406 424430
rect 477462 424374 477467 424430
rect 476928 424372 477467 424374
rect 477401 424369 477467 424372
rect 484342 424356 484348 424420
rect 484412 424418 484418 424420
rect 486200 424418 487000 424448
rect 484412 424358 487000 424418
rect 484412 424356 484418 424358
rect 486200 424328 487000 424358
rect 480897 424146 480963 424149
rect 476940 424144 480963 424146
rect 476940 424088 480902 424144
rect 480958 424088 480963 424144
rect 476940 424086 480963 424088
rect 480897 424083 480963 424086
rect 485814 423874 485820 423876
rect 476940 423814 485820 423874
rect 485814 423812 485820 423814
rect 485884 423812 485890 423876
rect 484526 423676 484532 423740
rect 484596 423738 484602 423740
rect 486200 423738 487000 423768
rect 484596 423678 487000 423738
rect 484596 423676 484602 423678
rect 486200 423648 487000 423678
rect 476940 423542 481098 423602
rect 477401 423466 477467 423469
rect 481038 423466 481098 423542
rect 481214 423540 481220 423604
rect 481284 423602 481290 423604
rect 481541 423602 481607 423605
rect 481284 423600 481607 423602
rect 481284 423544 481546 423600
rect 481602 423544 481607 423600
rect 481284 423542 481607 423544
rect 481284 423540 481290 423542
rect 481541 423539 481607 423542
rect 483422 423540 483428 423604
rect 483492 423602 483498 423604
rect 484117 423602 484183 423605
rect 483492 423600 484183 423602
rect 483492 423544 484122 423600
rect 484178 423544 484183 423600
rect 483492 423542 484183 423544
rect 483492 423540 483498 423542
rect 484117 423539 484183 423542
rect 482870 423466 482876 423468
rect 477401 423464 480914 423466
rect 477401 423408 477406 423464
rect 477462 423408 480914 423464
rect 477401 423406 480914 423408
rect 481038 423406 482876 423466
rect 477401 423403 477467 423406
rect 480854 423330 480914 423406
rect 482870 423404 482876 423406
rect 482940 423404 482946 423468
rect 483054 423330 483060 423332
rect 480854 423270 483060 423330
rect 483054 423268 483060 423270
rect 483124 423268 483130 423332
rect 476940 423202 477602 423262
rect 477542 423194 477602 423202
rect 485078 423194 485084 423196
rect 477542 423134 485084 423194
rect 485078 423132 485084 423134
rect 485148 423132 485154 423196
rect 477401 423072 477467 423075
rect 476928 423070 477467 423072
rect 476928 423014 477406 423070
rect 477462 423014 477467 423070
rect 476928 423012 477467 423014
rect 477401 423009 477467 423012
rect 480846 422996 480852 423060
rect 480916 423058 480922 423060
rect 486200 423058 487000 423088
rect 480916 422998 487000 423058
rect 480916 422996 480922 422998
rect 486200 422968 487000 422998
rect 486182 422786 486188 422788
rect 476940 422726 486188 422786
rect 486182 422724 486188 422726
rect 486252 422724 486258 422788
rect 485262 422514 485268 422516
rect 476940 422454 485268 422514
rect 485262 422452 485268 422454
rect 485332 422452 485338 422516
rect 484710 422316 484716 422380
rect 484780 422378 484786 422380
rect 486200 422378 487000 422408
rect 484780 422318 487000 422378
rect 484780 422316 484786 422318
rect 486200 422288 487000 422318
rect 484342 422242 484348 422244
rect 476940 422182 484348 422242
rect 484342 422180 484348 422182
rect 484412 422180 484418 422244
rect 478638 421970 478644 421972
rect 476940 421910 478644 421970
rect 478638 421908 478644 421910
rect 478708 421908 478714 421972
rect 485998 421834 486004 421836
rect 477358 421774 486004 421834
rect 477358 421712 477418 421774
rect 485998 421772 486004 421774
rect 486068 421772 486074 421836
rect 476928 421652 477418 421712
rect 486200 421698 487000 421728
rect 484902 421638 487000 421698
rect 481449 421426 481515 421429
rect 476940 421424 481515 421426
rect 476940 421368 481454 421424
rect 481510 421368 481515 421424
rect 476940 421366 481515 421368
rect 481449 421363 481515 421366
rect 484710 421290 484716 421292
rect 477358 421230 484716 421290
rect 477358 421168 477418 421230
rect 484710 421228 484716 421230
rect 484780 421228 484786 421292
rect 476928 421108 477418 421168
rect 484902 421154 484962 421638
rect 486200 421608 487000 421638
rect 482694 421094 484962 421154
rect 477902 420956 477908 421020
rect 477972 421018 477978 421020
rect 478505 421018 478571 421021
rect 477972 421016 478571 421018
rect 477972 420960 478510 421016
rect 478566 420960 478571 421016
rect 477972 420958 478571 420960
rect 477972 420956 477978 420958
rect 478505 420955 478571 420958
rect 482694 420882 482754 421094
rect 486200 421018 487000 421048
rect 476940 420822 482754 420882
rect 482878 420958 487000 421018
rect 482878 420610 482938 420958
rect 486200 420928 487000 420958
rect 476940 420550 482938 420610
rect 482134 420474 482140 420476
rect 477358 420414 482140 420474
rect 477358 420352 477418 420414
rect 482134 420412 482140 420414
rect 482204 420412 482210 420476
rect 476928 420292 477418 420352
rect 485814 420276 485820 420340
rect 485884 420338 485890 420340
rect 486200 420338 487000 420368
rect 485884 420278 487000 420338
rect 485884 420276 485890 420278
rect 486200 420248 487000 420278
rect 481214 420066 481220 420068
rect 476940 420006 481220 420066
rect 481214 420004 481220 420006
rect 481284 420004 481290 420068
rect 481449 420066 481515 420069
rect 484894 420066 484900 420068
rect 481449 420064 484900 420066
rect 481449 420008 481454 420064
rect 481510 420008 484900 420064
rect 481449 420006 484900 420008
rect 481449 420003 481515 420006
rect 484894 420004 484900 420006
rect 484964 420004 484970 420068
rect 481398 419868 481404 419932
rect 481468 419930 481474 419932
rect 481468 419870 483122 419930
rect 481468 419868 481474 419870
rect 481449 419794 481515 419797
rect 476940 419792 481515 419794
rect 476940 419736 481454 419792
rect 481510 419736 481515 419792
rect 476940 419734 481515 419736
rect 481449 419731 481515 419734
rect 481582 419732 481588 419796
rect 481652 419794 481658 419796
rect 482737 419794 482803 419797
rect 481652 419792 482803 419794
rect 481652 419736 482742 419792
rect 482798 419736 482803 419792
rect 481652 419734 482803 419736
rect 481652 419732 481658 419734
rect 482737 419731 482803 419734
rect 481950 419596 481956 419660
rect 482020 419658 482026 419660
rect 482829 419658 482895 419661
rect 482020 419656 482895 419658
rect 482020 419600 482834 419656
rect 482890 419600 482895 419656
rect 482020 419598 482895 419600
rect 483062 419658 483122 419870
rect 486200 419658 487000 419688
rect 483062 419598 487000 419658
rect 482020 419596 482026 419598
rect 482829 419595 482895 419598
rect 486200 419568 487000 419598
rect 480161 419524 480227 419525
rect 480110 419522 480116 419524
rect 480070 419462 480116 419522
rect 480180 419520 480227 419524
rect 480222 419464 480227 419520
rect 480110 419460 480116 419462
rect 480180 419460 480227 419464
rect 480161 419459 480227 419460
rect 476940 419394 477602 419454
rect 477542 419386 477602 419394
rect 484526 419386 484532 419388
rect 477542 419326 484532 419386
rect 484526 419324 484532 419326
rect 484596 419324 484602 419388
rect 478270 419250 478276 419252
rect 476940 419190 478276 419250
rect 478270 419188 478276 419190
rect 478340 419188 478346 419252
rect 486200 418978 487000 419008
rect 476940 418918 487000 418978
rect 486200 418888 487000 418918
rect 479558 418706 479564 418708
rect 476940 418646 479564 418706
rect 479558 418644 479564 418646
rect 479628 418644 479634 418708
rect 479374 418434 479380 418436
rect 476940 418374 479380 418434
rect 479374 418372 479380 418374
rect 479444 418372 479450 418436
rect 0 418298 800 418328
rect 0 418238 4170 418298
rect 0 418208 800 418238
rect 4110 418162 4170 418238
rect 478270 418236 478276 418300
rect 478340 418298 478346 418300
rect 478597 418298 478663 418301
rect 478340 418296 478663 418298
rect 478340 418240 478602 418296
rect 478658 418240 478663 418296
rect 478340 418238 478663 418240
rect 478340 418236 478346 418238
rect 478597 418235 478663 418238
rect 483238 418236 483244 418300
rect 483308 418298 483314 418300
rect 486200 418298 487000 418328
rect 483308 418238 487000 418298
rect 483308 418236 483314 418238
rect 486200 418208 487000 418238
rect 479517 418162 479583 418165
rect 4110 418102 10032 418162
rect 476940 418160 479583 418162
rect 476940 418104 479522 418160
rect 479578 418104 479583 418160
rect 476940 418102 479583 418104
rect 479517 418099 479583 418102
rect 479926 417890 479932 417892
rect 476940 417830 479932 417890
rect 479926 417828 479932 417830
rect 479996 417828 480002 417892
rect 0 417618 800 417648
rect 486200 417618 487000 417648
rect 0 417558 9506 417618
rect 476940 417558 487000 417618
rect 0 417528 800 417558
rect 9446 417360 9506 417558
rect 486200 417528 487000 417558
rect 9446 417300 10060 417360
rect 480069 417346 480135 417349
rect 476940 417344 480135 417346
rect 476940 417288 480074 417344
rect 480130 417288 480135 417344
rect 476940 417286 480135 417288
rect 480069 417283 480135 417286
rect 479742 417074 479748 417076
rect 476940 417014 479748 417074
rect 479742 417012 479748 417014
rect 479812 417012 479818 417076
rect 484342 416876 484348 416940
rect 484412 416938 484418 416940
rect 486200 416938 487000 416968
rect 484412 416878 487000 416938
rect 484412 416876 484418 416878
rect 486200 416848 487000 416878
rect 483238 416802 483244 416804
rect 476940 416742 483244 416802
rect 483238 416740 483244 416742
rect 483308 416740 483314 416804
rect 478689 416668 478755 416669
rect 478638 416604 478644 416668
rect 478708 416666 478755 416668
rect 478708 416664 478800 416666
rect 478750 416608 478800 416664
rect 478708 416606 478800 416608
rect 478708 416604 478755 416606
rect 482318 416604 482324 416668
rect 482388 416666 482394 416668
rect 482921 416666 482987 416669
rect 482388 416664 482987 416666
rect 482388 416608 482926 416664
rect 482982 416608 482987 416664
rect 482388 416606 482987 416608
rect 482388 416604 482394 416606
rect 478689 416603 478755 416604
rect 482921 416603 482987 416606
rect 483054 416604 483060 416668
rect 483124 416666 483130 416668
rect 484209 416666 484275 416669
rect 483124 416664 484275 416666
rect 483124 416608 484214 416664
rect 484270 416608 484275 416664
rect 483124 416606 484275 416608
rect 483124 416604 483130 416606
rect 484209 416603 484275 416606
rect 480110 416530 480116 416532
rect 9446 416428 10060 416488
rect 476940 416470 480116 416530
rect 480110 416468 480116 416470
rect 480180 416468 480186 416532
rect 0 416258 800 416288
rect 9446 416258 9506 416428
rect 483790 416258 483796 416260
rect 0 416198 9506 416258
rect 476940 416198 483796 416258
rect 0 416168 800 416198
rect 483790 416196 483796 416198
rect 483860 416196 483866 416260
rect 484526 416196 484532 416260
rect 484596 416258 484602 416260
rect 486200 416258 487000 416288
rect 484596 416198 487000 416258
rect 484596 416196 484602 416198
rect 486200 416168 487000 416198
rect 481766 415986 481772 415988
rect 476940 415926 481772 415986
rect 481766 415924 481772 415926
rect 481836 415924 481842 415988
rect 478086 415714 478092 415716
rect 9446 415612 10060 415672
rect 476940 415654 478092 415714
rect 478086 415652 478092 415654
rect 478156 415652 478162 415716
rect 0 415578 800 415608
rect 9446 415578 9506 415612
rect 0 415518 9506 415578
rect 0 415488 800 415518
rect 484710 415516 484716 415580
rect 484780 415578 484786 415580
rect 486200 415578 487000 415608
rect 484780 415518 487000 415578
rect 484780 415516 484786 415518
rect 486200 415488 487000 415518
rect 484342 415442 484348 415444
rect 476940 415382 484348 415442
rect 484342 415380 484348 415382
rect 484412 415380 484418 415444
rect 478454 415244 478460 415308
rect 478524 415306 478530 415308
rect 478781 415306 478847 415309
rect 478524 415304 478847 415306
rect 478524 415248 478786 415304
rect 478842 415248 478847 415304
rect 478524 415246 478847 415248
rect 478524 415244 478530 415246
rect 478781 415243 478847 415246
rect 483606 415244 483612 415308
rect 483676 415306 483682 415308
rect 484301 415306 484367 415309
rect 483676 415304 484367 415306
rect 483676 415248 484306 415304
rect 484362 415248 484367 415304
rect 483676 415246 484367 415248
rect 483676 415244 483682 415246
rect 484301 415243 484367 415246
rect 482870 415170 482876 415172
rect 476940 415110 482876 415170
rect 482870 415108 482876 415110
rect 482940 415108 482946 415172
rect 0 414898 800 414928
rect 486200 414898 487000 414928
rect 0 414838 10032 414898
rect 476940 414838 487000 414898
rect 0 414808 800 414838
rect 486200 414808 487000 414838
rect 482502 414626 482508 414628
rect 476940 414566 482508 414626
rect 482502 414564 482508 414566
rect 482572 414564 482578 414628
rect 477534 414354 477540 414356
rect 476940 414294 477540 414354
rect 477534 414292 477540 414294
rect 477604 414292 477610 414356
rect 0 414218 800 414248
rect 0 414158 9506 414218
rect 0 414128 800 414158
rect 9446 414096 9506 414158
rect 479926 414156 479932 414220
rect 479996 414218 480002 414220
rect 486200 414218 487000 414248
rect 479996 414158 487000 414218
rect 479996 414156 480002 414158
rect 486200 414128 487000 414158
rect 9446 414036 10060 414096
rect 484526 414082 484532 414084
rect 476940 414022 484532 414082
rect 484526 414020 484532 414022
rect 484596 414020 484602 414084
rect 478270 413810 478276 413812
rect 476940 413750 478276 413810
rect 478270 413748 478276 413750
rect 478340 413748 478346 413812
rect 0 413538 800 413568
rect 481398 413538 481404 413540
rect 0 413478 9506 413538
rect 476940 413478 481404 413538
rect 0 413448 800 413478
rect 9446 413280 9506 413478
rect 481398 413476 481404 413478
rect 481468 413476 481474 413540
rect 484158 413476 484164 413540
rect 484228 413538 484234 413540
rect 486200 413538 487000 413568
rect 484228 413478 487000 413538
rect 484228 413476 484234 413478
rect 486200 413448 487000 413478
rect 9446 413220 10060 413280
rect 477902 413266 477908 413268
rect 476940 413206 477908 413266
rect 477902 413204 477908 413206
rect 477972 413204 477978 413268
rect 478638 412994 478644 412996
rect 476940 412934 478644 412994
rect 478638 412932 478644 412934
rect 478708 412932 478714 412996
rect 480294 412796 480300 412860
rect 480364 412858 480370 412860
rect 486200 412858 487000 412888
rect 480364 412798 487000 412858
rect 480364 412796 480370 412798
rect 486200 412768 487000 412798
rect 484710 412722 484716 412724
rect 476940 412662 484716 412722
rect 484710 412660 484716 412662
rect 484780 412660 484786 412724
rect 485814 412450 485820 412452
rect 9446 412348 10060 412408
rect 476940 412390 485820 412450
rect 485814 412388 485820 412390
rect 485884 412388 485890 412452
rect 0 412178 800 412208
rect 9446 412178 9506 412348
rect 480846 412178 480852 412180
rect 0 412118 9506 412178
rect 476940 412118 480852 412178
rect 0 412088 800 412118
rect 480846 412116 480852 412118
rect 480916 412116 480922 412180
rect 484342 412116 484348 412180
rect 484412 412178 484418 412180
rect 486200 412178 487000 412208
rect 484412 412118 487000 412178
rect 484412 412116 484418 412118
rect 486200 412088 487000 412118
rect 480294 411906 480300 411908
rect 476940 411846 480300 411906
rect 480294 411844 480300 411846
rect 480364 411844 480370 411908
rect 479926 411634 479932 411636
rect 9446 411532 10060 411592
rect 476940 411574 479932 411634
rect 479926 411572 479932 411574
rect 479996 411572 480002 411636
rect 0 411498 800 411528
rect 9446 411498 9506 411532
rect 0 411438 9506 411498
rect 0 411408 800 411438
rect 484526 411436 484532 411500
rect 484596 411498 484602 411500
rect 486200 411498 487000 411528
rect 484596 411438 487000 411498
rect 484596 411436 484602 411438
rect 486200 411408 487000 411438
rect 484158 411362 484164 411364
rect 476940 411302 484164 411362
rect 484158 411300 484164 411302
rect 484228 411300 484234 411364
rect 484342 411090 484348 411092
rect 476940 411030 484348 411090
rect 484342 411028 484348 411030
rect 484412 411028 484418 411092
rect 0 410818 800 410848
rect 486200 410818 487000 410848
rect 0 410758 10032 410818
rect 476940 410758 487000 410818
rect 0 410728 800 410758
rect 486200 410728 487000 410758
rect 478454 410546 478460 410548
rect 476940 410486 478460 410546
rect 478454 410484 478460 410486
rect 478524 410484 478530 410548
rect 483422 410274 483428 410276
rect 476940 410214 483428 410274
rect 483422 410212 483428 410214
rect 483492 410212 483498 410276
rect 0 410138 800 410168
rect 0 410078 9506 410138
rect 0 410048 800 410078
rect 9446 410016 9506 410078
rect 482870 410076 482876 410140
rect 482940 410138 482946 410140
rect 486200 410138 487000 410168
rect 482940 410078 487000 410138
rect 482940 410076 482946 410078
rect 486200 410048 487000 410078
rect 9446 409956 10060 410016
rect 484526 410002 484532 410004
rect 476940 409942 484532 410002
rect 484526 409940 484532 409942
rect 484596 409940 484602 410004
rect 481582 409730 481588 409732
rect 476940 409670 481588 409730
rect 481582 409668 481588 409670
rect 481652 409668 481658 409732
rect 0 409458 800 409488
rect 486200 409458 487000 409488
rect 0 409398 9506 409458
rect 476940 409398 487000 409458
rect 0 409368 800 409398
rect 9446 409200 9506 409398
rect 486200 409368 487000 409398
rect 9446 409140 10060 409200
rect 483054 409186 483060 409188
rect 476940 409126 483060 409186
rect 483054 409124 483060 409126
rect 483124 409124 483130 409188
rect 481950 408914 481956 408916
rect 476940 408854 481956 408914
rect 481950 408852 481956 408854
rect 482020 408852 482026 408916
rect 484342 408716 484348 408780
rect 484412 408778 484418 408780
rect 486200 408778 487000 408808
rect 484412 408718 487000 408778
rect 484412 408716 484418 408718
rect 486200 408688 487000 408718
rect 482870 408642 482876 408644
rect 476940 408582 482876 408642
rect 482870 408580 482876 408582
rect 482940 408580 482946 408644
rect 483606 408370 483612 408372
rect 9446 408268 10060 408328
rect 476940 408310 483612 408370
rect 483606 408308 483612 408310
rect 483676 408308 483682 408372
rect 0 408098 800 408128
rect 9446 408098 9506 408268
rect 486200 408098 487000 408128
rect 0 408038 9506 408098
rect 476940 408038 487000 408098
rect 0 408008 800 408038
rect 486200 408008 487000 408038
rect 484342 407826 484348 407828
rect 476940 407766 484348 407826
rect 484342 407764 484348 407766
rect 484412 407764 484418 407828
rect 482318 407554 482324 407556
rect 9446 407452 10060 407512
rect 476940 407494 482324 407554
rect 482318 407492 482324 407494
rect 482388 407492 482394 407556
rect 0 407418 800 407448
rect 9446 407418 9506 407452
rect 486200 407418 487000 407448
rect 0 407358 9506 407418
rect 477358 407358 487000 407418
rect 0 407328 800 407358
rect 477358 407296 477418 407358
rect 486200 407328 487000 407358
rect 476928 407236 477418 407296
rect 476940 406882 477602 406942
rect 0 406738 800 406768
rect 477542 406738 477602 406882
rect 486200 406738 487000 406768
rect 0 406678 10032 406738
rect 477542 406678 487000 406738
rect 0 406648 800 406678
rect 476940 406610 477418 406670
rect 486200 406648 487000 406678
rect 477358 406602 477418 406610
rect 477534 406602 477540 406604
rect 477358 406542 477540 406602
rect 477534 406540 477540 406542
rect 477604 406540 477610 406604
rect 477718 406466 477724 406468
rect 476940 406406 477724 406466
rect 477718 406404 477724 406406
rect 477788 406404 477794 406468
rect 0 406058 800 406088
rect 476940 406066 477602 406126
rect 477542 406058 477602 406066
rect 486200 406058 487000 406088
rect 0 405998 9506 406058
rect 477542 405998 487000 406058
rect 0 405968 800 405998
rect 9446 405936 9506 405998
rect 486200 405968 487000 405998
rect 9446 405876 10060 405936
rect 476940 405794 477602 405854
rect 477542 405786 477602 405794
rect 486182 405786 486188 405788
rect 477542 405726 486188 405786
rect 486182 405724 486188 405726
rect 486252 405724 486258 405788
rect 476940 405522 477602 405582
rect 0 405378 800 405408
rect 477542 405378 477602 405522
rect 486200 405378 487000 405408
rect 0 405318 9506 405378
rect 477542 405318 487000 405378
rect 0 405288 800 405318
rect 9446 405120 9506 405318
rect 476940 405250 477418 405310
rect 486200 405288 487000 405318
rect 477358 405242 477418 405250
rect 479374 405242 479380 405244
rect 477358 405182 479380 405242
rect 479374 405180 479380 405182
rect 479444 405180 479450 405244
rect 9446 405060 10060 405120
rect 485998 405106 486004 405108
rect 476940 405046 486004 405106
rect 485998 405044 486004 405046
rect 486068 405044 486074 405108
rect 476940 404706 477602 404766
rect 477542 404698 477602 404706
rect 486200 404698 487000 404728
rect 477542 404638 487000 404698
rect 486200 404608 487000 404638
rect 476940 404434 477602 404494
rect 477542 404426 477602 404434
rect 486182 404426 486188 404428
rect 477542 404366 486188 404426
rect 486182 404364 486188 404366
rect 486252 404364 486258 404428
rect 9446 404188 10060 404248
rect 0 404018 800 404048
rect 9446 404018 9506 404188
rect 476940 404162 477602 404222
rect 0 403958 9506 404018
rect 477542 404018 477602 404162
rect 486200 404018 487000 404048
rect 477542 403958 487000 404018
rect 0 403928 800 403958
rect 476940 403890 477418 403950
rect 486200 403928 487000 403958
rect 477358 403882 477418 403890
rect 479558 403882 479564 403884
rect 477358 403822 479564 403882
rect 479558 403820 479564 403822
rect 479628 403820 479634 403884
rect 479742 403746 479748 403748
rect 476940 403686 479748 403746
rect 479742 403684 479748 403686
rect 479812 403684 479818 403748
rect 9446 403372 10060 403432
rect 0 403338 800 403368
rect 9446 403338 9506 403372
rect 476940 403346 477602 403406
rect 0 403278 9506 403338
rect 477542 403338 477602 403346
rect 486200 403338 487000 403368
rect 477542 403278 487000 403338
rect 0 403248 800 403278
rect 486200 403248 487000 403278
rect 480846 403202 480852 403204
rect 476940 403142 480852 403202
rect 480846 403140 480852 403142
rect 480916 403140 480922 403204
rect 476940 402802 477602 402862
rect 0 402658 800 402688
rect 477542 402658 477602 402802
rect 486200 402658 487000 402688
rect 0 402598 10032 402658
rect 477542 402598 487000 402658
rect 0 402568 800 402598
rect 476940 402530 477418 402590
rect 486200 402568 487000 402598
rect 477358 402522 477418 402530
rect 478086 402522 478092 402524
rect 477358 402462 478092 402522
rect 478086 402460 478092 402462
rect 478156 402460 478162 402524
rect 483238 402386 483244 402388
rect 476940 402326 483244 402386
rect 483238 402324 483244 402326
rect 483308 402324 483314 402388
rect 0 401978 800 402008
rect 476940 401986 477602 402046
rect 477542 401978 477602 401986
rect 486200 401978 487000 402008
rect 0 401918 9506 401978
rect 477542 401918 487000 401978
rect 0 401888 800 401918
rect 9446 401856 9506 401918
rect 486200 401888 487000 401918
rect 9446 401796 10060 401856
rect 477350 401774 477356 401776
rect 476940 401714 477356 401774
rect 477350 401712 477356 401714
rect 477420 401712 477426 401776
rect 476940 401442 477602 401502
rect 477542 401434 477602 401442
rect 477542 401374 480270 401434
rect 0 401298 800 401328
rect 480210 401298 480270 401374
rect 486200 401298 487000 401328
rect 0 401238 9506 401298
rect 480210 401238 487000 401298
rect 0 401208 800 401238
rect 9446 401040 9506 401238
rect 476940 401170 477602 401230
rect 486200 401208 487000 401238
rect 477542 401162 477602 401170
rect 484894 401162 484900 401164
rect 477542 401102 484900 401162
rect 484894 401100 484900 401102
rect 484964 401100 484970 401164
rect 9446 400980 10060 401040
rect 484710 401026 484716 401028
rect 476940 400966 484716 401026
rect 484710 400964 484716 400966
rect 484780 400964 484786 401028
rect 476940 400626 477602 400686
rect 477542 400618 477602 400626
rect 486200 400618 487000 400648
rect 477542 400558 487000 400618
rect 486200 400528 487000 400558
rect 476940 400354 477602 400414
rect 477542 400346 477602 400354
rect 484526 400346 484532 400348
rect 477542 400286 484532 400346
rect 484526 400284 484532 400286
rect 484596 400284 484602 400348
rect 9446 400108 10060 400168
rect 0 399938 800 399968
rect 9446 399938 9506 400108
rect 476940 400082 477602 400142
rect 477542 400074 477602 400082
rect 477542 400014 480270 400074
rect 0 399878 9506 399938
rect 480210 399938 480270 400014
rect 486200 399938 487000 399968
rect 480210 399878 487000 399938
rect 0 399848 800 399878
rect 476940 399810 477602 399870
rect 486200 399848 487000 399878
rect 477542 399802 477602 399810
rect 484342 399802 484348 399804
rect 477542 399742 484348 399802
rect 484342 399740 484348 399742
rect 484412 399740 484418 399804
rect 478638 399666 478644 399668
rect 476940 399606 478644 399666
rect 478638 399604 478644 399606
rect 478708 399604 478714 399668
rect 477534 399468 477540 399532
rect 477604 399530 477610 399532
rect 478781 399530 478847 399533
rect 477604 399528 478847 399530
rect 477604 399472 478786 399528
rect 478842 399472 478847 399528
rect 477604 399470 478847 399472
rect 477604 399468 477610 399470
rect 478781 399467 478847 399470
rect 9446 399292 10060 399352
rect 0 399258 800 399288
rect 9446 399258 9506 399292
rect 476940 399266 477602 399326
rect 0 399198 9506 399258
rect 477542 399258 477602 399266
rect 486200 399258 487000 399288
rect 477542 399198 487000 399258
rect 0 399168 800 399198
rect 486200 399168 487000 399198
rect 476940 398994 477602 399054
rect 477542 398986 477602 398994
rect 477542 398926 480270 398986
rect 476940 398790 477602 398850
rect 477542 398714 477602 398790
rect 477718 398788 477724 398852
rect 477788 398850 477794 398852
rect 478689 398850 478755 398853
rect 479517 398850 479583 398853
rect 477788 398848 478755 398850
rect 477788 398792 478694 398848
rect 478750 398792 478755 398848
rect 477788 398790 478755 398792
rect 477788 398788 477794 398790
rect 478689 398787 478755 398790
rect 478830 398848 479583 398850
rect 478830 398792 479522 398848
rect 479578 398792 479583 398848
rect 478830 398790 479583 398792
rect 478830 398714 478890 398790
rect 479517 398787 479583 398790
rect 477542 398654 478890 398714
rect 0 398578 800 398608
rect 480210 398578 480270 398926
rect 486200 398578 487000 398608
rect 0 398518 10032 398578
rect 480210 398518 487000 398578
rect 0 398488 800 398518
rect 486200 398488 487000 398518
rect 0 397898 800 397928
rect 0 397838 9506 397898
rect 0 397808 800 397838
rect 9446 397776 9506 397838
rect 478638 397836 478644 397900
rect 478708 397898 478714 397900
rect 486200 397898 487000 397928
rect 478708 397838 487000 397898
rect 478708 397836 478714 397838
rect 486200 397808 487000 397838
rect 9446 397716 10060 397776
rect 0 397218 800 397248
rect 0 397158 9506 397218
rect 0 397128 800 397158
rect 9446 396960 9506 397158
rect 484342 397156 484348 397220
rect 484412 397218 484418 397220
rect 486200 397218 487000 397248
rect 484412 397158 487000 397218
rect 484412 397156 484418 397158
rect 486200 397128 487000 397158
rect 9446 396900 10060 396960
rect 484526 396476 484532 396540
rect 484596 396538 484602 396540
rect 486200 396538 487000 396568
rect 484596 396478 487000 396538
rect 484596 396476 484602 396478
rect 486200 396448 487000 396478
rect 6870 396070 10032 396130
rect 0 395858 800 395888
rect 6870 395858 6930 396070
rect 0 395798 6930 395858
rect 0 395768 800 395798
rect 484710 395796 484716 395860
rect 484780 395858 484786 395860
rect 486200 395858 487000 395888
rect 484780 395798 487000 395858
rect 484780 395796 484786 395798
rect 486200 395768 487000 395798
rect 9446 395212 10060 395272
rect 0 395178 800 395208
rect 9446 395178 9506 395212
rect 0 395118 9506 395178
rect 0 395088 800 395118
rect 484894 395116 484900 395180
rect 484964 395178 484970 395180
rect 486200 395178 487000 395208
rect 484964 395118 487000 395178
rect 484964 395116 484970 395118
rect 486200 395088 487000 395118
rect 0 394498 800 394528
rect 0 394438 10032 394498
rect 0 394408 800 394438
rect 477350 394436 477356 394500
rect 477420 394498 477426 394500
rect 486200 394498 487000 394528
rect 477420 394438 487000 394498
rect 477420 394436 477426 394438
rect 486200 394408 487000 394438
rect 0 393818 800 393848
rect 0 393758 9506 393818
rect 0 393728 800 393758
rect 9446 393696 9506 393758
rect 483238 393756 483244 393820
rect 483308 393818 483314 393820
rect 486200 393818 487000 393848
rect 483308 393758 487000 393818
rect 483308 393756 483314 393758
rect 486200 393728 487000 393758
rect 9446 393636 10060 393696
rect 0 393138 800 393168
rect 0 393078 9506 393138
rect 0 393048 800 393078
rect 9446 392880 9506 393078
rect 478086 393076 478092 393140
rect 478156 393138 478162 393140
rect 486200 393138 487000 393168
rect 478156 393078 487000 393138
rect 478156 393076 478162 393078
rect 486200 393048 487000 393078
rect 9446 392820 10060 392880
rect 480846 392396 480852 392460
rect 480916 392458 480922 392460
rect 486200 392458 487000 392488
rect 480916 392398 487000 392458
rect 480916 392396 480922 392398
rect 486200 392368 487000 392398
rect 6870 391990 10032 392050
rect 0 391778 800 391808
rect 6870 391778 6930 391990
rect 0 391718 6930 391778
rect 0 391688 800 391718
rect 479742 391716 479748 391780
rect 479812 391778 479818 391780
rect 486200 391778 487000 391808
rect 479812 391718 487000 391778
rect 479812 391716 479818 391718
rect 486200 391688 487000 391718
rect 9446 391132 10060 391192
rect 0 391098 800 391128
rect 9446 391098 9506 391132
rect 0 391038 9506 391098
rect 0 391008 800 391038
rect 479558 391036 479564 391100
rect 479628 391098 479634 391100
rect 486200 391098 487000 391128
rect 479628 391038 487000 391098
rect 479628 391036 479634 391038
rect 486200 391008 487000 391038
rect 0 390418 800 390448
rect 486200 390420 487000 390448
rect 0 390358 10032 390418
rect 0 390328 800 390358
rect 486200 390356 486372 390420
rect 486436 390356 487000 390420
rect 486200 390328 487000 390356
rect 0 389738 800 389768
rect 0 389678 9506 389738
rect 0 389648 800 389678
rect 9446 389616 9506 389678
rect 485998 389676 486004 389740
rect 486068 389738 486074 389740
rect 486200 389738 487000 389768
rect 486068 389678 487000 389738
rect 486068 389676 486074 389678
rect 486200 389648 487000 389678
rect 9446 389556 10060 389616
rect 0 389058 800 389088
rect 0 388998 9506 389058
rect 0 388968 800 388998
rect 9446 388800 9506 388998
rect 479374 388996 479380 389060
rect 479444 389058 479450 389060
rect 486200 389058 487000 389088
rect 479444 388998 487000 389058
rect 479444 388996 479450 388998
rect 486200 388968 487000 388998
rect 9446 388740 10060 388800
rect 486200 388380 487000 388408
rect 486200 388316 486556 388380
rect 486620 388316 487000 388380
rect 486200 388288 487000 388316
rect 9446 387868 10060 387928
rect 9446 387834 9506 387868
rect 6870 387774 9506 387834
rect 0 387698 800 387728
rect 6870 387698 6930 387774
rect 0 387638 6930 387698
rect 478689 387698 478755 387701
rect 486200 387698 487000 387728
rect 478689 387696 487000 387698
rect 478689 387640 478694 387696
rect 478750 387640 487000 387696
rect 478689 387638 487000 387640
rect 0 387608 800 387638
rect 478689 387635 478755 387638
rect 486200 387608 487000 387638
rect 9446 387052 10060 387112
rect 0 387018 800 387048
rect 9446 387018 9506 387052
rect 0 386958 9506 387018
rect 478781 387018 478847 387021
rect 486200 387018 487000 387048
rect 478781 387016 487000 387018
rect 478781 386960 478786 387016
rect 478842 386960 487000 387016
rect 478781 386958 487000 386960
rect 0 386928 800 386958
rect 478781 386955 478847 386958
rect 486200 386928 487000 386958
rect 0 386338 800 386368
rect 479517 386338 479583 386341
rect 486200 386338 487000 386368
rect 0 386278 10032 386338
rect 479517 386336 487000 386338
rect 479517 386280 479522 386336
rect 479578 386280 487000 386336
rect 479517 386278 487000 386280
rect 0 386248 800 386278
rect 479517 386275 479583 386278
rect 486200 386248 487000 386278
rect 0 385658 800 385688
rect 0 385598 9506 385658
rect 0 385568 800 385598
rect 9446 385536 9506 385598
rect 9446 385476 10060 385536
rect 0 384978 800 385008
rect 0 384918 9506 384978
rect 0 384888 800 384918
rect 9446 384720 9506 384918
rect 9446 384660 10060 384720
rect 9446 383788 10060 383848
rect 9446 383754 9506 383788
rect 5582 383694 9506 383754
rect 0 383618 800 383648
rect 5582 383618 5642 383694
rect 0 383558 5642 383618
rect 0 383528 800 383558
rect 9446 382972 10060 383032
rect 0 382938 800 382968
rect 9446 382938 9506 382972
rect 0 382878 9506 382938
rect 0 382848 800 382878
rect 0 382258 800 382288
rect 0 382198 10032 382258
rect 0 382168 800 382198
rect 0 381578 800 381608
rect 0 381518 9506 381578
rect 0 381488 800 381518
rect 9446 381456 9506 381518
rect 9446 381396 10060 381456
rect 0 373418 800 373448
rect 0 373358 9506 373418
rect 0 373328 800 373358
rect 9446 373176 9506 373358
rect 9446 373116 10032 373176
rect 9446 372244 10032 372304
rect 0 372058 800 372088
rect 9446 372058 9506 372244
rect 0 371998 9506 372058
rect 0 371968 800 371998
rect 9446 371428 10032 371488
rect 0 371378 800 371408
rect 9446 371378 9506 371428
rect 0 371318 9506 371378
rect 0 371288 800 371318
rect 0 370698 800 370728
rect 0 370638 10032 370698
rect 0 370608 800 370638
rect 0 370018 800 370048
rect 0 369958 9506 370018
rect 0 369928 800 369958
rect 9446 369912 9506 369958
rect 9446 369852 10032 369912
rect 0 369338 800 369368
rect 0 369278 9506 369338
rect 0 369248 800 369278
rect 9446 369096 9506 369278
rect 9446 369036 10032 369096
rect 9446 368164 10032 368224
rect 0 367978 800 368008
rect 9446 367978 9506 368164
rect 0 367918 9506 367978
rect 0 367888 800 367918
rect 9446 367348 10032 367408
rect 0 367298 800 367328
rect 9446 367298 9506 367348
rect 0 367238 9506 367298
rect 0 367208 800 367238
rect 0 366618 800 366648
rect 0 366558 10032 366618
rect 0 366528 800 366558
rect 0 365938 800 365968
rect 0 365878 9506 365938
rect 0 365848 800 365878
rect 9446 365832 9506 365878
rect 9446 365772 10032 365832
rect 0 365258 800 365288
rect 0 365198 9506 365258
rect 0 365168 800 365198
rect 9446 365016 9506 365198
rect 9446 364956 10032 365016
rect 9446 364084 10032 364144
rect 0 363898 800 363928
rect 9446 363898 9506 364084
rect 0 363838 9506 363898
rect 0 363808 800 363838
rect 9446 363268 10032 363328
rect 0 363218 800 363248
rect 9446 363218 9506 363268
rect 0 363158 9506 363218
rect 0 363128 800 363158
rect 0 362538 800 362568
rect 0 362478 10032 362538
rect 0 362448 800 362478
rect 0 361858 800 361888
rect 0 361798 9506 361858
rect 0 361768 800 361798
rect 9446 361752 9506 361798
rect 9446 361692 10032 361752
rect 0 361178 800 361208
rect 0 361118 9506 361178
rect 0 361088 800 361118
rect 9446 360936 9506 361118
rect 9446 360876 10032 360936
rect 481541 360498 481607 360501
rect 486200 360498 487000 360528
rect 481541 360496 487000 360498
rect 481541 360440 481546 360496
rect 481602 360440 487000 360496
rect 481541 360438 487000 360440
rect 481541 360435 481607 360438
rect 486200 360408 487000 360438
rect 9446 360004 10032 360064
rect 0 359818 800 359848
rect 9446 359818 9506 360004
rect 0 359758 9506 359818
rect 484301 359818 484367 359821
rect 486200 359818 487000 359848
rect 484301 359816 487000 359818
rect 484301 359760 484306 359816
rect 484362 359760 487000 359816
rect 484301 359758 487000 359760
rect 0 359728 800 359758
rect 484301 359755 484367 359758
rect 486200 359728 487000 359758
rect 9446 359188 10032 359248
rect 0 359138 800 359168
rect 9446 359138 9506 359188
rect 0 359078 9506 359138
rect 482921 359138 482987 359141
rect 486200 359138 487000 359168
rect 482921 359136 487000 359138
rect 482921 359080 482926 359136
rect 482982 359080 487000 359136
rect 482921 359078 487000 359080
rect 0 359048 800 359078
rect 482921 359075 482987 359078
rect 486200 359048 487000 359078
rect 0 358458 800 358488
rect 481449 358458 481515 358461
rect 486200 358458 487000 358488
rect 0 358398 10032 358458
rect 481449 358456 487000 358458
rect 481449 358400 481454 358456
rect 481510 358400 487000 358456
rect 481449 358398 487000 358400
rect 0 358368 800 358398
rect 481449 358395 481515 358398
rect 486200 358368 487000 358398
rect 0 357778 800 357808
rect 484209 357778 484275 357781
rect 486200 357778 487000 357808
rect 0 357718 9506 357778
rect 0 357688 800 357718
rect 9446 357672 9506 357718
rect 484209 357776 487000 357778
rect 484209 357720 484214 357776
rect 484270 357720 487000 357776
rect 484209 357718 487000 357720
rect 484209 357715 484275 357718
rect 486200 357688 487000 357718
rect 9446 357612 10032 357672
rect 0 357098 800 357128
rect 0 357038 9506 357098
rect 0 357008 800 357038
rect 9446 356856 9506 357038
rect 482134 357036 482140 357100
rect 482204 357098 482210 357100
rect 486200 357098 487000 357128
rect 482204 357038 487000 357098
rect 482204 357036 482210 357038
rect 486200 357008 487000 357038
rect 9446 356796 10032 356856
rect 483606 356356 483612 356420
rect 483676 356418 483682 356420
rect 486200 356418 487000 356448
rect 483676 356358 487000 356418
rect 483676 356356 483682 356358
rect 486200 356328 487000 356358
rect 9446 355924 10032 355984
rect 0 355738 800 355768
rect 9446 355738 9506 355924
rect 0 355678 9506 355738
rect 0 355648 800 355678
rect 480846 355676 480852 355740
rect 480916 355738 480922 355740
rect 486200 355738 487000 355768
rect 480916 355678 487000 355738
rect 480916 355676 480922 355678
rect 486200 355648 487000 355678
rect 9446 355108 10032 355168
rect 0 355058 800 355088
rect 9446 355058 9506 355108
rect 0 354998 9506 355058
rect 478781 355058 478847 355061
rect 486200 355058 487000 355088
rect 478781 355056 487000 355058
rect 478781 355000 478786 355056
rect 478842 355000 487000 355056
rect 478781 354998 487000 355000
rect 0 354968 800 354998
rect 478781 354995 478847 354998
rect 486200 354968 487000 354998
rect 0 354378 800 354408
rect 0 354318 10032 354378
rect 0 354288 800 354318
rect 478086 354316 478092 354380
rect 478156 354378 478162 354380
rect 486200 354378 487000 354408
rect 478156 354318 487000 354378
rect 478156 354316 478162 354318
rect 486200 354288 487000 354318
rect 0 353698 800 353728
rect 478689 353698 478755 353701
rect 486200 353698 487000 353728
rect 0 353638 9506 353698
rect 0 353608 800 353638
rect 9446 353592 9506 353638
rect 478689 353696 487000 353698
rect 478689 353640 478694 353696
rect 478750 353640 487000 353696
rect 478689 353638 487000 353640
rect 478689 353635 478755 353638
rect 486200 353608 487000 353638
rect 9446 353532 10032 353592
rect 0 353018 800 353048
rect 0 352958 9506 353018
rect 0 352928 800 352958
rect 9446 352776 9506 352958
rect 478270 352956 478276 353020
rect 478340 353018 478346 353020
rect 486200 353018 487000 353048
rect 478340 352958 487000 353018
rect 478340 352956 478346 352958
rect 486200 352928 487000 352958
rect 9446 352716 10032 352776
rect 478454 352276 478460 352340
rect 478524 352338 478530 352340
rect 486200 352338 487000 352368
rect 478524 352278 487000 352338
rect 478524 352276 478530 352278
rect 486200 352248 487000 352278
rect 6870 351870 10032 351930
rect 0 351658 800 351688
rect 6870 351658 6930 351870
rect 0 351598 6930 351658
rect 0 351568 800 351598
rect 481030 351596 481036 351660
rect 481100 351658 481106 351660
rect 486200 351658 487000 351688
rect 481100 351598 487000 351658
rect 481100 351596 481106 351598
rect 486200 351568 487000 351598
rect 9446 351028 10032 351088
rect 0 350978 800 351008
rect 9446 350978 9506 351028
rect 0 350918 9506 350978
rect 0 350888 800 350918
rect 482318 350916 482324 350980
rect 482388 350978 482394 350980
rect 486200 350978 487000 351008
rect 482388 350918 487000 350978
rect 482388 350916 482394 350918
rect 486200 350888 487000 350918
rect 0 350298 800 350328
rect 0 350238 10032 350298
rect 0 350208 800 350238
rect 477902 350236 477908 350300
rect 477972 350298 477978 350300
rect 486200 350298 487000 350328
rect 477972 350238 487000 350298
rect 477972 350236 477978 350238
rect 486200 350208 487000 350238
rect 0 349618 800 349648
rect 477125 349618 477191 349621
rect 486200 349618 487000 349648
rect 0 349558 9506 349618
rect 0 349528 800 349558
rect 9446 349512 9506 349558
rect 477125 349616 487000 349618
rect 477125 349560 477130 349616
rect 477186 349560 487000 349616
rect 477125 349558 487000 349560
rect 477125 349555 477191 349558
rect 486200 349528 487000 349558
rect 9446 349452 10032 349512
rect 481214 348876 481220 348940
rect 481284 348938 481290 348940
rect 486200 348938 487000 348968
rect 481284 348878 487000 348938
rect 481284 348876 481290 348878
rect 486200 348848 487000 348878
rect 9446 348580 10032 348640
rect 0 348258 800 348288
rect 9446 348258 9506 348580
rect 0 348198 9506 348258
rect 0 348168 800 348198
rect 482686 348196 482692 348260
rect 482756 348258 482762 348260
rect 486200 348258 487000 348288
rect 482756 348198 487000 348258
rect 482756 348196 482762 348198
rect 486200 348168 487000 348198
rect 6870 347790 10032 347850
rect 0 347578 800 347608
rect 6870 347578 6930 347790
rect 0 347518 6930 347578
rect 0 347488 800 347518
rect 482502 347516 482508 347580
rect 482572 347578 482578 347580
rect 486200 347578 487000 347608
rect 482572 347518 487000 347578
rect 482572 347516 482578 347518
rect 486200 347488 487000 347518
rect 9446 346948 10032 347008
rect 0 346898 800 346928
rect 9446 346898 9506 346948
rect 0 346838 9506 346898
rect 482277 346898 482343 346901
rect 486200 346898 487000 346928
rect 482277 346896 487000 346898
rect 482277 346840 482282 346896
rect 482338 346840 487000 346896
rect 482277 346838 487000 346840
rect 0 346808 800 346838
rect 482277 346835 482343 346838
rect 486200 346808 487000 346838
rect 0 346218 800 346248
rect 0 346158 10032 346218
rect 0 346128 800 346158
rect 483790 346156 483796 346220
rect 483860 346218 483866 346220
rect 486200 346218 487000 346248
rect 483860 346158 487000 346218
rect 483860 346156 483866 346158
rect 486200 346128 487000 346158
rect 0 345538 800 345568
rect 0 345478 9506 345538
rect 0 345448 800 345478
rect 9446 345432 9506 345478
rect 479374 345476 479380 345540
rect 479444 345538 479450 345540
rect 486200 345538 487000 345568
rect 479444 345478 487000 345538
rect 479444 345476 479450 345478
rect 486200 345448 487000 345478
rect 9446 345372 10032 345432
rect 0 344858 800 344888
rect 0 344798 9506 344858
rect 0 344768 800 344798
rect 9446 344616 9506 344798
rect 485998 344796 486004 344860
rect 486068 344858 486074 344860
rect 486200 344858 487000 344888
rect 486068 344798 487000 344858
rect 486068 344796 486074 344798
rect 486200 344768 487000 344798
rect 9446 344556 10032 344616
rect 481398 344116 481404 344180
rect 481468 344178 481474 344180
rect 486200 344178 487000 344208
rect 481468 344118 487000 344178
rect 481468 344116 481474 344118
rect 486200 344088 487000 344118
rect 6870 343710 10032 343770
rect 0 343498 800 343528
rect 6870 343498 6930 343710
rect 0 343438 6930 343498
rect 0 343408 800 343438
rect 479742 343436 479748 343500
rect 479812 343498 479818 343500
rect 486200 343498 487000 343528
rect 479812 343438 487000 343498
rect 479812 343436 479818 343438
rect 486200 343408 487000 343438
rect 9446 342868 10032 342928
rect 0 342818 800 342848
rect 9446 342818 9506 342868
rect 0 342758 9506 342818
rect 0 342728 800 342758
rect 483974 342756 483980 342820
rect 484044 342818 484050 342820
rect 486200 342818 487000 342848
rect 484044 342758 487000 342818
rect 484044 342756 484050 342758
rect 486200 342728 487000 342758
rect 0 342138 800 342168
rect 0 342078 10032 342138
rect 0 342048 800 342078
rect 483422 342076 483428 342140
rect 483492 342138 483498 342140
rect 486200 342138 487000 342168
rect 483492 342078 487000 342138
rect 483492 342076 483498 342078
rect 486200 342048 487000 342078
rect 0 341458 800 341488
rect 0 341398 9506 341458
rect 0 341368 800 341398
rect 9446 341352 9506 341398
rect 484342 341396 484348 341460
rect 484412 341458 484418 341460
rect 486200 341458 487000 341488
rect 484412 341398 487000 341458
rect 484412 341396 484418 341398
rect 486200 341368 487000 341398
rect 9446 341292 10032 341352
rect 0 340778 800 340808
rect 0 340718 9506 340778
rect 0 340688 800 340718
rect 9446 340536 9506 340718
rect 477350 340716 477356 340780
rect 477420 340778 477426 340780
rect 486200 340778 487000 340808
rect 477420 340718 487000 340778
rect 477420 340716 477426 340718
rect 486200 340688 487000 340718
rect 9446 340476 10032 340536
rect 478822 340036 478828 340100
rect 478892 340098 478898 340100
rect 486200 340098 487000 340128
rect 478892 340038 487000 340098
rect 478892 340036 478898 340038
rect 486200 340008 487000 340038
rect 9446 339604 10032 339664
rect 9446 339554 9506 339604
rect 6870 339494 9506 339554
rect 0 339418 800 339448
rect 6870 339418 6930 339494
rect 0 339358 6930 339418
rect 0 339328 800 339358
rect 483238 339356 483244 339420
rect 483308 339418 483314 339420
rect 486200 339418 487000 339448
rect 483308 339358 487000 339418
rect 483308 339356 483314 339358
rect 486200 339328 487000 339358
rect 9446 338788 10032 338848
rect 0 338738 800 338768
rect 9446 338738 9506 338788
rect 0 338678 9506 338738
rect 0 338648 800 338678
rect 479558 338676 479564 338740
rect 479628 338738 479634 338740
rect 486200 338738 487000 338768
rect 479628 338678 487000 338738
rect 479628 338676 479634 338678
rect 486200 338648 487000 338678
rect 483422 338194 483428 338196
rect 476968 338134 483428 338194
rect 483422 338132 483428 338134
rect 483492 338132 483498 338196
rect 0 338058 800 338088
rect 486200 338058 487000 338088
rect 0 337998 10032 338058
rect 477358 337998 487000 338058
rect 0 337968 800 337998
rect 477358 337990 477418 337998
rect 476940 337930 477418 337990
rect 486200 337968 487000 337998
rect 483238 337650 483244 337652
rect 476968 337590 483244 337650
rect 483238 337588 483244 337590
rect 483308 337588 483314 337652
rect 478822 337514 478828 337516
rect 477174 337454 478828 337514
rect 477174 337446 477234 337454
rect 478822 337452 478828 337454
rect 478892 337452 478898 337516
rect 0 337378 800 337408
rect 476940 337386 477234 337446
rect 486200 337378 487000 337408
rect 0 337318 9506 337378
rect 0 337288 800 337318
rect 9446 337272 9506 337318
rect 477358 337318 487000 337378
rect 9446 337212 10032 337272
rect 477358 337174 477418 337318
rect 486200 337288 487000 337318
rect 476940 337114 477418 337174
rect 477350 336902 477356 336904
rect 476940 336842 477356 336902
rect 477350 336840 477356 336842
rect 477420 336840 477426 336904
rect 0 336698 800 336728
rect 0 336638 9506 336698
rect 0 336608 800 336638
rect 9446 336456 9506 336638
rect 480294 336636 480300 336700
rect 480364 336698 480370 336700
rect 481449 336698 481515 336701
rect 480364 336696 481515 336698
rect 480364 336640 481454 336696
rect 481510 336640 481515 336696
rect 480364 336638 481515 336640
rect 480364 336636 480370 336638
rect 481449 336635 481515 336638
rect 481766 336636 481772 336700
rect 481836 336698 481842 336700
rect 482921 336698 482987 336701
rect 481836 336696 482987 336698
rect 481836 336640 482926 336696
rect 482982 336640 482987 336696
rect 481836 336638 482987 336640
rect 481836 336636 481842 336638
rect 482921 336635 482987 336638
rect 483054 336636 483060 336700
rect 483124 336698 483130 336700
rect 484209 336698 484275 336701
rect 483124 336696 484275 336698
rect 483124 336640 484214 336696
rect 484270 336640 484275 336696
rect 483124 336638 484275 336640
rect 483124 336636 483130 336638
rect 484209 336635 484275 336638
rect 484710 336636 484716 336700
rect 484780 336698 484786 336700
rect 486200 336698 487000 336728
rect 484780 336638 487000 336698
rect 484780 336636 484786 336638
rect 486200 336608 487000 336638
rect 482686 336562 482692 336564
rect 476968 336502 482692 336562
rect 482686 336500 482692 336502
rect 482756 336500 482762 336564
rect 9446 336396 10032 336456
rect 484342 336290 484348 336292
rect 476968 336230 484348 336290
rect 484342 336228 484348 336230
rect 484412 336228 484418 336292
rect 481214 336018 481220 336020
rect 476968 335958 481220 336018
rect 481214 335956 481220 335958
rect 481284 335956 481290 336020
rect 486200 336018 487000 336048
rect 483246 335958 487000 336018
rect 477350 335820 477356 335884
rect 477420 335882 477426 335884
rect 483246 335882 483306 335958
rect 486200 335928 487000 335958
rect 477420 335822 483306 335882
rect 477420 335820 477426 335822
rect 477125 335814 477191 335817
rect 476940 335812 477191 335814
rect 476940 335756 477130 335812
rect 477186 335756 477191 335812
rect 476940 335754 477191 335756
rect 477125 335751 477191 335754
rect 483974 335474 483980 335476
rect 476968 335414 483980 335474
rect 483974 335412 483980 335414
rect 484044 335412 484050 335476
rect 484342 335276 484348 335340
rect 484412 335338 484418 335340
rect 486200 335338 487000 335368
rect 484412 335278 487000 335338
rect 484412 335276 484418 335278
rect 486200 335248 487000 335278
rect 477902 335202 477908 335204
rect 476968 335142 477908 335202
rect 477902 335140 477908 335142
rect 477972 335140 477978 335204
rect 479742 334930 479748 334932
rect 476968 334870 479748 334930
rect 479742 334868 479748 334870
rect 479812 334868 479818 334932
rect 481398 334794 481404 334796
rect 477358 334734 481404 334794
rect 477358 334726 477418 334734
rect 481398 334732 481404 334734
rect 481468 334732 481474 334796
rect 476940 334666 477418 334726
rect 479006 334596 479012 334660
rect 479076 334658 479082 334660
rect 486200 334658 487000 334688
rect 479076 334598 487000 334658
rect 479076 334596 479082 334598
rect 486200 334568 487000 334598
rect 484710 334386 484716 334388
rect 476968 334326 484716 334386
rect 484710 334324 484716 334326
rect 484780 334324 484786 334388
rect 485998 334250 486004 334252
rect 477358 334190 486004 334250
rect 477358 334182 477418 334190
rect 485998 334188 486004 334190
rect 486068 334188 486074 334252
rect 476940 334122 477418 334182
rect 478689 334116 478755 334117
rect 478638 334052 478644 334116
rect 478708 334114 478755 334116
rect 478708 334112 478800 334114
rect 478750 334056 478800 334112
rect 478708 334054 478800 334056
rect 478708 334052 478755 334054
rect 480478 334052 480484 334116
rect 480548 334114 480554 334116
rect 481541 334114 481607 334117
rect 480548 334112 481607 334114
rect 480548 334056 481546 334112
rect 481602 334056 481607 334112
rect 480548 334054 481607 334056
rect 480548 334052 480554 334054
rect 478689 334051 478755 334052
rect 481541 334051 481607 334054
rect 483238 334052 483244 334116
rect 483308 334114 483314 334116
rect 484301 334114 484367 334117
rect 483308 334112 484367 334114
rect 483308 334056 484306 334112
rect 484362 334056 484367 334112
rect 483308 334054 484367 334056
rect 483308 334052 483314 334054
rect 484301 334051 484367 334054
rect 478822 333916 478828 333980
rect 478892 333978 478898 333980
rect 486200 333978 487000 334008
rect 478892 333918 487000 333978
rect 478892 333916 478898 333918
rect 477350 333910 477356 333912
rect 476940 333850 477356 333910
rect 477350 333848 477356 333850
rect 477420 333848 477426 333912
rect 486200 333888 487000 333918
rect 479374 333570 479380 333572
rect 476968 333510 479380 333570
rect 479374 333508 479380 333510
rect 479444 333508 479450 333572
rect 483790 333434 483796 333436
rect 477358 333374 483796 333434
rect 477358 333366 477418 333374
rect 483790 333372 483796 333374
rect 483860 333372 483866 333436
rect 476940 333306 477418 333366
rect 483422 333236 483428 333300
rect 483492 333298 483498 333300
rect 486200 333298 487000 333328
rect 483492 333238 487000 333298
rect 483492 333236 483498 333238
rect 486200 333208 487000 333238
rect 484342 333026 484348 333028
rect 476968 332966 484348 333026
rect 484342 332964 484348 332966
rect 484412 332964 484418 333028
rect 482277 332754 482343 332757
rect 476968 332752 482343 332754
rect 476968 332696 482282 332752
rect 482338 332696 482343 332752
rect 476968 332694 482343 332696
rect 482277 332691 482343 332694
rect 477350 332556 477356 332620
rect 477420 332618 477426 332620
rect 486200 332618 487000 332648
rect 477420 332558 487000 332618
rect 477420 332556 477426 332558
rect 486200 332528 487000 332558
rect 479006 332482 479012 332484
rect 476968 332422 479012 332482
rect 479006 332420 479012 332422
rect 479076 332420 479082 332484
rect 482502 332210 482508 332212
rect 476968 332150 482508 332210
rect 482502 332148 482508 332150
rect 482572 332148 482578 332212
rect 482318 332074 482324 332076
rect 477358 332014 482324 332074
rect 477358 332006 477418 332014
rect 482318 332012 482324 332014
rect 482388 332012 482394 332076
rect 476940 331946 477418 332006
rect 482870 331876 482876 331940
rect 482940 331938 482946 331940
rect 486200 331938 487000 331968
rect 482940 331878 487000 331938
rect 482940 331876 482946 331878
rect 486200 331848 487000 331878
rect 478822 331666 478828 331668
rect 476968 331606 478828 331666
rect 478822 331604 478828 331606
rect 478892 331604 478898 331668
rect 483422 331394 483428 331396
rect 476968 331334 483428 331394
rect 483422 331332 483428 331334
rect 483492 331332 483498 331396
rect 486200 331258 487000 331288
rect 483062 331198 487000 331258
rect 477350 331190 477356 331192
rect 476940 331130 477356 331190
rect 477350 331128 477356 331130
rect 477420 331128 477426 331192
rect 479558 330850 479564 330852
rect 476968 330790 479564 330850
rect 479558 330788 479564 330790
rect 479628 330788 479634 330852
rect 482870 330578 482876 330580
rect 476968 330518 482876 330578
rect 482870 330516 482876 330518
rect 482940 330516 482946 330580
rect 483062 330306 483122 331198
rect 486200 331168 487000 331198
rect 486200 330578 487000 330608
rect 476968 330246 483122 330306
rect 483246 330518 487000 330578
rect 483246 330034 483306 330518
rect 486200 330488 487000 330518
rect 476968 329974 483306 330034
rect 486200 329898 487000 329928
rect 484350 329838 487000 329898
rect 484350 329762 484410 329838
rect 486200 329808 487000 329838
rect 476968 329702 484410 329762
rect 477902 329564 477908 329628
rect 477972 329626 477978 329628
rect 478781 329626 478847 329629
rect 477972 329624 478847 329626
rect 477972 329568 478786 329624
rect 478842 329568 478847 329624
rect 477972 329566 478847 329568
rect 477972 329564 477978 329566
rect 478781 329563 478847 329566
rect 481030 329490 481036 329492
rect 476968 329430 481036 329490
rect 481030 329428 481036 329430
rect 481100 329428 481106 329492
rect 478454 329354 478460 329356
rect 477174 329294 478460 329354
rect 477174 329286 477234 329294
rect 478454 329292 478460 329294
rect 478524 329292 478530 329356
rect 476940 329226 477234 329286
rect 486200 329218 487000 329248
rect 477358 329158 487000 329218
rect 477358 329014 477418 329158
rect 486200 329128 487000 329158
rect 476940 328954 477418 329014
rect 478270 328674 478276 328676
rect 476968 328614 478276 328674
rect 478270 328612 478276 328614
rect 478340 328612 478346 328676
rect 486200 328538 487000 328568
rect 482970 328478 487000 328538
rect 482970 328402 483030 328478
rect 486200 328448 487000 328478
rect 476968 328342 483030 328402
rect 478638 328130 478644 328132
rect 9446 328060 10060 328120
rect 476968 328070 478644 328130
rect 478638 328068 478644 328070
rect 478708 328068 478714 328132
rect 0 327858 800 327888
rect 9446 327858 9506 328060
rect 478086 327994 478092 327996
rect 477174 327934 478092 327994
rect 477174 327926 477234 327934
rect 478086 327932 478092 327934
rect 478156 327932 478162 327996
rect 476940 327866 477234 327926
rect 486200 327858 487000 327888
rect 0 327798 9506 327858
rect 477358 327798 487000 327858
rect 0 327768 800 327798
rect 477358 327654 477418 327798
rect 486200 327768 487000 327798
rect 476940 327594 477418 327654
rect 477902 327314 477908 327316
rect 9446 327244 10060 327304
rect 476968 327254 477908 327314
rect 477902 327252 477908 327254
rect 477972 327252 477978 327316
rect 0 327178 800 327208
rect 9446 327178 9506 327244
rect 486200 327178 487000 327208
rect 0 327118 9506 327178
rect 484350 327118 487000 327178
rect 0 327088 800 327118
rect 484350 327042 484410 327118
rect 486200 327088 487000 327118
rect 476968 326982 484410 327042
rect 480846 326770 480852 326772
rect 476968 326710 480852 326770
rect 480846 326708 480852 326710
rect 480916 326708 480922 326772
rect 483606 326634 483612 326636
rect 477358 326574 483612 326634
rect 477358 326566 477418 326574
rect 483606 326572 483612 326574
rect 483676 326572 483682 326636
rect 0 326498 800 326528
rect 476940 326506 477418 326566
rect 486200 326498 487000 326528
rect 0 326438 10032 326498
rect 483246 326438 487000 326498
rect 0 326408 800 326438
rect 483246 326226 483306 326438
rect 486200 326408 487000 326438
rect 476968 326166 483306 326226
rect 482134 325954 482140 325956
rect 476968 325894 482140 325954
rect 482134 325892 482140 325894
rect 482204 325892 482210 325956
rect 0 325818 800 325848
rect 486200 325818 487000 325848
rect 0 325758 4906 325818
rect 0 325728 800 325758
rect 4846 325682 4906 325758
rect 482970 325758 487000 325818
rect 482970 325682 483030 325758
rect 486200 325728 487000 325758
rect 4846 325622 10032 325682
rect 476968 325622 483030 325682
rect 483054 325410 483060 325412
rect 476968 325350 483060 325410
rect 483054 325348 483060 325350
rect 483124 325348 483130 325412
rect 0 325138 800 325168
rect 480294 325138 480300 325140
rect 0 325078 9506 325138
rect 476968 325078 480300 325138
rect 0 325048 800 325078
rect 9446 324934 9506 325078
rect 480294 325076 480300 325078
rect 480364 325076 480370 325140
rect 486200 325138 487000 325168
rect 483246 325078 487000 325138
rect 9446 324874 10060 324934
rect 483246 324866 483306 325078
rect 486200 325048 487000 325078
rect 476968 324806 483306 324866
rect 481766 324594 481772 324596
rect 476968 324534 481772 324594
rect 481766 324532 481772 324534
rect 481836 324532 481842 324596
rect 486200 324458 487000 324488
rect 482970 324398 487000 324458
rect 482970 324322 483030 324398
rect 486200 324368 487000 324398
rect 476968 324262 483030 324322
rect 483238 324050 483244 324052
rect 9446 323980 10060 324040
rect 476968 323990 483244 324050
rect 483238 323988 483244 323990
rect 483308 323988 483314 324052
rect 0 323778 800 323808
rect 9446 323778 9506 323980
rect 480478 323778 480484 323780
rect 0 323718 9506 323778
rect 476968 323718 480484 323778
rect 0 323688 800 323718
rect 480478 323716 480484 323718
rect 480548 323716 480554 323780
rect 486200 323778 487000 323808
rect 483246 323718 487000 323778
rect 483246 323506 483306 323718
rect 486200 323688 487000 323718
rect 476968 323446 483306 323506
rect 9446 323164 10060 323224
rect 476940 323164 477418 323224
rect 0 323098 800 323128
rect 9446 323098 9506 323164
rect 0 323038 9506 323098
rect 477358 323098 477418 323164
rect 486200 323098 487000 323128
rect 477358 323038 487000 323098
rect 0 323008 800 323038
rect 486200 323008 487000 323038
rect 481766 322962 481772 322964
rect 476968 322902 481772 322962
rect 481766 322900 481772 322902
rect 481836 322900 481842 322964
rect 480662 322690 480668 322692
rect 476968 322630 480668 322690
rect 480662 322628 480668 322630
rect 480732 322628 480738 322692
rect 0 322418 800 322448
rect 486200 322418 487000 322448
rect 0 322358 10032 322418
rect 476968 322358 487000 322418
rect 0 322328 800 322358
rect 486200 322328 487000 322358
rect 483054 322146 483060 322148
rect 476968 322086 483060 322146
rect 483054 322084 483060 322086
rect 483124 322084 483130 322148
rect 476940 321804 477418 321864
rect 0 321738 800 321768
rect 477358 321738 477418 321804
rect 486200 321738 487000 321768
rect 0 321678 9506 321738
rect 477358 321678 487000 321738
rect 0 321648 800 321678
rect 9446 321670 9506 321678
rect 9446 321610 10060 321670
rect 486200 321648 487000 321678
rect 481582 321602 481588 321604
rect 476968 321542 481588 321602
rect 481582 321540 481588 321542
rect 481652 321540 481658 321604
rect 480846 321330 480852 321332
rect 476968 321270 480852 321330
rect 480846 321268 480852 321270
rect 480916 321268 480922 321332
rect 0 321058 800 321088
rect 486200 321058 487000 321088
rect 0 320998 9506 321058
rect 476968 320998 487000 321058
rect 0 320968 800 320998
rect 9446 320854 9506 320998
rect 486200 320968 487000 320998
rect 9446 320794 10060 320854
rect 483606 320786 483612 320788
rect 476968 320726 483612 320786
rect 483606 320724 483612 320726
rect 483676 320724 483682 320788
rect 476940 320444 477418 320504
rect 477358 320378 477418 320444
rect 486200 320378 487000 320408
rect 477358 320318 487000 320378
rect 486200 320288 487000 320318
rect 483790 320242 483796 320244
rect 476968 320182 483796 320242
rect 483790 320180 483796 320182
rect 483860 320180 483866 320244
rect 483974 319970 483980 319972
rect 9446 319900 10060 319960
rect 476968 319910 483980 319970
rect 483974 319908 483980 319910
rect 484044 319908 484050 319972
rect 0 319698 800 319728
rect 9446 319698 9506 319900
rect 486200 319698 487000 319728
rect 0 319638 9506 319698
rect 476968 319638 487000 319698
rect 0 319608 800 319638
rect 486200 319608 487000 319638
rect 481030 319426 481036 319428
rect 476968 319366 481036 319426
rect 481030 319364 481036 319366
rect 481100 319364 481106 319428
rect 9446 319084 10060 319144
rect 476940 319084 477418 319144
rect 0 319018 800 319048
rect 9446 319018 9506 319084
rect 0 318958 9506 319018
rect 477358 319018 477418 319084
rect 486200 319018 487000 319048
rect 477358 318958 487000 319018
rect 0 318928 800 318958
rect 486200 318928 487000 318958
rect 482134 318882 482140 318884
rect 476968 318822 482140 318882
rect 482134 318820 482140 318822
rect 482204 318820 482210 318884
rect 480662 318684 480668 318748
rect 480732 318746 480738 318748
rect 481541 318746 481607 318749
rect 480732 318744 481607 318746
rect 480732 318688 481546 318744
rect 481602 318688 481607 318744
rect 480732 318686 481607 318688
rect 480732 318684 480738 318686
rect 481541 318683 481607 318686
rect 482318 318610 482324 318612
rect 476968 318550 482324 318610
rect 482318 318548 482324 318550
rect 482388 318548 482394 318612
rect 0 318338 800 318368
rect 486200 318338 487000 318368
rect 0 318278 10032 318338
rect 476968 318278 487000 318338
rect 0 318248 800 318278
rect 486200 318248 487000 318278
rect 481214 318066 481220 318068
rect 476968 318006 481220 318066
rect 481214 318004 481220 318006
rect 481284 318004 481290 318068
rect 476968 317734 483306 317794
rect 0 317658 800 317688
rect 481398 317658 481404 317660
rect 0 317598 9506 317658
rect 0 317568 800 317598
rect 9446 317590 9506 317598
rect 477358 317598 481404 317658
rect 477358 317590 477418 317598
rect 481398 317596 481404 317598
rect 481468 317596 481474 317660
rect 483246 317658 483306 317734
rect 486200 317658 487000 317688
rect 483246 317598 487000 317658
rect 9446 317530 10060 317590
rect 476940 317530 477418 317590
rect 486200 317568 487000 317598
rect 479374 317250 479380 317252
rect 476968 317190 479380 317250
rect 479374 317188 479380 317190
rect 479444 317188 479450 317252
rect 0 316978 800 317008
rect 486200 316978 487000 317008
rect 0 316918 9506 316978
rect 476968 316918 487000 316978
rect 0 316888 800 316918
rect 9446 316774 9506 316918
rect 486200 316888 487000 316918
rect 9446 316714 10060 316774
rect 479742 316706 479748 316708
rect 476968 316646 479748 316706
rect 479742 316644 479748 316646
rect 479812 316644 479818 316708
rect 476940 316364 477418 316424
rect 477358 316298 477418 316364
rect 486200 316298 487000 316328
rect 477358 316238 487000 316298
rect 486200 316208 487000 316238
rect 479926 316162 479932 316164
rect 476968 316102 479932 316162
rect 479926 316100 479932 316102
rect 479996 316100 480002 316164
rect 478086 315890 478092 315892
rect 9446 315820 10060 315880
rect 476968 315830 478092 315890
rect 478086 315828 478092 315830
rect 478156 315828 478162 315892
rect 0 315618 800 315648
rect 9446 315618 9506 315820
rect 486200 315618 487000 315648
rect 0 315558 9506 315618
rect 476968 315558 487000 315618
rect 0 315528 800 315558
rect 486200 315528 487000 315558
rect 478270 315346 478276 315348
rect 476968 315286 478276 315346
rect 478270 315284 478276 315286
rect 478340 315284 478346 315348
rect 9446 315004 10060 315064
rect 476968 315014 483306 315074
rect 0 314938 800 314968
rect 9446 314938 9506 315004
rect 0 314878 9506 314938
rect 0 314848 800 314878
rect 479374 314876 479380 314940
rect 479444 314938 479450 314940
rect 480161 314938 480227 314941
rect 479444 314936 480227 314938
rect 479444 314880 480166 314936
rect 480222 314880 480227 314936
rect 479444 314878 480227 314880
rect 483246 314938 483306 315014
rect 486200 314938 487000 314968
rect 483246 314878 487000 314938
rect 479444 314876 479450 314878
rect 480161 314875 480227 314878
rect 486200 314848 487000 314878
rect 486049 314802 486115 314805
rect 476968 314800 486115 314802
rect 476968 314744 486054 314800
rect 486110 314744 486115 314800
rect 476968 314742 486115 314744
rect 486049 314739 486115 314742
rect 482277 314530 482343 314533
rect 476968 314528 482343 314530
rect 476968 314472 482282 314528
rect 482338 314472 482343 314528
rect 476968 314470 482343 314472
rect 482277 314467 482343 314470
rect 0 314258 800 314288
rect 486200 314258 487000 314288
rect 0 314198 10032 314258
rect 476968 314198 487000 314258
rect 0 314168 800 314198
rect 486200 314168 487000 314198
rect 486182 313986 486188 313988
rect 476968 313926 486188 313986
rect 486182 313924 486188 313926
rect 486252 313924 486258 313988
rect 476940 313644 477418 313704
rect 0 313578 800 313608
rect 477358 313578 477418 313644
rect 486200 313578 487000 313608
rect 0 313518 9506 313578
rect 477358 313518 487000 313578
rect 0 313488 800 313518
rect 9446 313510 9506 313518
rect 9446 313450 10060 313510
rect 486200 313488 487000 313518
rect 485078 313442 485084 313444
rect 476968 313382 485084 313442
rect 485078 313380 485084 313382
rect 485148 313380 485154 313444
rect 485998 313170 486004 313172
rect 476968 313110 486004 313170
rect 485998 313108 486004 313110
rect 486068 313108 486074 313172
rect 0 312898 800 312928
rect 486200 312898 487000 312928
rect 0 312838 9506 312898
rect 476968 312838 487000 312898
rect 0 312808 800 312838
rect 9446 312694 9506 312838
rect 486200 312808 487000 312838
rect 9446 312634 10060 312694
rect 485814 312626 485820 312628
rect 476968 312566 485820 312626
rect 485814 312564 485820 312566
rect 485884 312564 485890 312628
rect 476940 312284 477418 312344
rect 477358 312218 477418 312284
rect 486200 312218 487000 312248
rect 477358 312158 487000 312218
rect 486200 312128 487000 312158
rect 485630 312082 485636 312084
rect 476968 312022 485636 312082
rect 485630 312020 485636 312022
rect 485700 312020 485706 312084
rect 481766 311884 481772 311948
rect 481836 311946 481842 311948
rect 482921 311946 482987 311949
rect 481836 311944 482987 311946
rect 481836 311888 482926 311944
rect 482982 311888 482987 311944
rect 481836 311886 482987 311888
rect 481836 311884 481842 311886
rect 482921 311883 482987 311886
rect 484894 311810 484900 311812
rect 9446 311740 10060 311800
rect 476968 311750 484900 311810
rect 484894 311748 484900 311750
rect 484964 311748 484970 311812
rect 0 311538 800 311568
rect 9446 311538 9506 311740
rect 486200 311538 487000 311568
rect 0 311478 9506 311538
rect 476968 311478 487000 311538
rect 0 311448 800 311478
rect 486200 311448 487000 311478
rect 476940 311196 477418 311256
rect 479742 311204 479748 311268
rect 479812 311266 479818 311268
rect 480069 311266 480135 311269
rect 479812 311264 480135 311266
rect 479812 311208 480074 311264
rect 480130 311208 480135 311264
rect 479812 311206 480135 311208
rect 479812 311204 479818 311206
rect 480069 311203 480135 311206
rect 483054 311204 483060 311268
rect 483124 311266 483130 311268
rect 484301 311266 484367 311269
rect 483124 311264 484367 311266
rect 483124 311208 484306 311264
rect 484362 311208 484367 311264
rect 483124 311206 484367 311208
rect 483124 311204 483130 311206
rect 484301 311203 484367 311206
rect 477358 311130 477418 311196
rect 485262 311130 485268 311132
rect 477358 311070 485268 311130
rect 485262 311068 485268 311070
rect 485332 311068 485338 311132
rect 9446 310924 10060 310984
rect 476940 310924 477418 310984
rect 0 310858 800 310888
rect 9446 310858 9506 310924
rect 0 310798 9506 310858
rect 477358 310858 477418 310924
rect 486200 310858 487000 310888
rect 477358 310798 487000 310858
rect 0 310768 800 310798
rect 486200 310768 487000 310798
rect 485446 310722 485452 310724
rect 476968 310662 485452 310722
rect 485446 310660 485452 310662
rect 485516 310660 485522 310724
rect 479977 310452 480043 310453
rect 481449 310452 481515 310453
rect 478638 310450 478644 310452
rect 476968 310390 478644 310450
rect 478638 310388 478644 310390
rect 478708 310388 478714 310452
rect 479926 310450 479932 310452
rect 479886 310390 479932 310450
rect 479996 310448 480043 310452
rect 481398 310450 481404 310452
rect 480038 310392 480043 310448
rect 479926 310388 479932 310390
rect 479996 310388 480043 310392
rect 481358 310390 481404 310450
rect 481468 310448 481515 310452
rect 481510 310392 481515 310448
rect 481398 310388 481404 310390
rect 481468 310388 481515 310392
rect 479977 310387 480043 310388
rect 481449 310387 481515 310388
rect 0 310178 800 310208
rect 486200 310178 487000 310208
rect 0 310118 10032 310178
rect 476968 310118 487000 310178
rect 0 310088 800 310118
rect 486200 310088 487000 310118
rect 482870 309906 482876 309908
rect 476968 309846 482876 309906
rect 482870 309844 482876 309846
rect 482940 309844 482946 309908
rect 476940 309564 477418 309624
rect 0 309498 800 309528
rect 477358 309498 477418 309564
rect 486200 309498 487000 309528
rect 0 309438 9506 309498
rect 477358 309438 487000 309498
rect 0 309408 800 309438
rect 9446 309430 9506 309438
rect 9446 309370 10060 309430
rect 486200 309408 487000 309438
rect 484342 309362 484348 309364
rect 476968 309302 484348 309362
rect 484342 309300 484348 309302
rect 484412 309300 484418 309364
rect 476968 309030 483306 309090
rect 481582 308892 481588 308956
rect 481652 308954 481658 308956
rect 482829 308954 482895 308957
rect 481652 308952 482895 308954
rect 481652 308896 482834 308952
rect 482890 308896 482895 308952
rect 481652 308894 482895 308896
rect 481652 308892 481658 308894
rect 482829 308891 482895 308894
rect 0 308818 800 308848
rect 483246 308818 483306 309030
rect 486200 308818 487000 308848
rect 0 308758 9506 308818
rect 0 308728 800 308758
rect 9446 308614 9506 308758
rect 476940 308748 477418 308808
rect 483246 308758 487000 308818
rect 9446 308554 10060 308614
rect 477358 308546 477418 308748
rect 486200 308728 487000 308758
rect 486182 308546 486188 308548
rect 477358 308486 486188 308546
rect 486182 308484 486188 308486
rect 486252 308484 486258 308548
rect 484342 308076 484348 308140
rect 484412 308138 484418 308140
rect 486200 308138 487000 308168
rect 484412 308078 487000 308138
rect 484412 308076 484418 308078
rect 486200 308048 487000 308078
rect 9446 307660 10060 307720
rect 0 307458 800 307488
rect 9446 307458 9506 307660
rect 0 307398 9506 307458
rect 0 307368 800 307398
rect 482870 307396 482876 307460
rect 482940 307458 482946 307460
rect 486200 307458 487000 307488
rect 482940 307398 487000 307458
rect 482940 307396 482946 307398
rect 486200 307368 487000 307398
rect 9446 306844 10060 306904
rect 0 306778 800 306808
rect 9446 306778 9506 306844
rect 0 306718 9506 306778
rect 0 306688 800 306718
rect 478638 306716 478644 306780
rect 478708 306778 478714 306780
rect 486200 306778 487000 306808
rect 478708 306718 487000 306778
rect 478708 306716 478714 306718
rect 486200 306688 487000 306718
rect 0 306098 800 306128
rect 0 306038 10032 306098
rect 0 306008 800 306038
rect 485446 306036 485452 306100
rect 485516 306098 485522 306100
rect 486200 306098 487000 306128
rect 485516 306038 487000 306098
rect 485516 306036 485522 306038
rect 486200 306008 487000 306038
rect 0 305418 800 305448
rect 0 305358 9506 305418
rect 0 305328 800 305358
rect 9446 305350 9506 305358
rect 485262 305356 485268 305420
rect 485332 305418 485338 305420
rect 486200 305418 487000 305448
rect 485332 305358 487000 305418
rect 485332 305356 485338 305358
rect 9446 305290 10060 305350
rect 486200 305328 487000 305358
rect 0 304738 800 304768
rect 0 304678 9506 304738
rect 0 304648 800 304678
rect 9446 304534 9506 304678
rect 484894 304676 484900 304740
rect 484964 304738 484970 304740
rect 486200 304738 487000 304768
rect 484964 304678 487000 304738
rect 484964 304676 484970 304678
rect 486200 304648 487000 304678
rect 9446 304474 10060 304534
rect 485630 303996 485636 304060
rect 485700 304058 485706 304060
rect 486200 304058 487000 304088
rect 485700 303998 487000 304058
rect 485700 303996 485706 303998
rect 486200 303968 487000 303998
rect 6870 303590 10032 303650
rect 0 303378 800 303408
rect 6870 303378 6930 303590
rect 0 303318 6930 303378
rect 0 303288 800 303318
rect 485814 303316 485820 303380
rect 485884 303378 485890 303380
rect 486200 303378 487000 303408
rect 485884 303318 487000 303378
rect 485884 303316 485890 303318
rect 486200 303288 487000 303318
rect 9446 302764 10060 302824
rect 0 302698 800 302728
rect 9446 302698 9506 302764
rect 0 302638 9506 302698
rect 0 302608 800 302638
rect 485998 302636 486004 302700
rect 486068 302698 486074 302700
rect 486200 302698 487000 302728
rect 486068 302638 487000 302698
rect 486068 302636 486074 302638
rect 486200 302608 487000 302638
rect 0 302018 800 302048
rect 0 301958 10032 302018
rect 0 301928 800 301958
rect 485078 301956 485084 302020
rect 485148 302018 485154 302020
rect 486200 302018 487000 302048
rect 485148 301958 487000 302018
rect 485148 301956 485154 301958
rect 486200 301928 487000 301958
rect 0 301338 800 301368
rect 486200 301340 487000 301368
rect 0 301278 9506 301338
rect 0 301248 800 301278
rect 9446 301270 9506 301278
rect 486200 301276 486372 301340
rect 486436 301276 487000 301340
rect 9446 301210 10060 301270
rect 486200 301248 487000 301276
rect 0 300658 800 300688
rect 482277 300658 482343 300661
rect 486200 300658 487000 300688
rect 0 300598 9506 300658
rect 0 300568 800 300598
rect 9446 300454 9506 300598
rect 482277 300656 487000 300658
rect 482277 300600 482282 300656
rect 482338 300600 487000 300656
rect 482277 300598 487000 300600
rect 482277 300595 482343 300598
rect 486200 300568 487000 300598
rect 9446 300394 10060 300454
rect 486049 299978 486115 299981
rect 486200 299978 487000 300008
rect 486049 299976 487000 299978
rect 486049 299920 486054 299976
rect 486110 299920 487000 299976
rect 486049 299918 487000 299920
rect 486049 299915 486115 299918
rect 486200 299888 487000 299918
rect 6870 299510 10032 299570
rect 0 299298 800 299328
rect 6870 299298 6930 299510
rect 0 299238 6930 299298
rect 0 299208 800 299238
rect 478270 299236 478276 299300
rect 478340 299298 478346 299300
rect 486200 299298 487000 299328
rect 478340 299238 487000 299298
rect 478340 299236 478346 299238
rect 486200 299208 487000 299238
rect 9446 298684 10060 298744
rect 0 298618 800 298648
rect 9446 298618 9506 298684
rect 0 298558 9506 298618
rect 0 298528 800 298558
rect 478086 298556 478092 298620
rect 478156 298618 478162 298620
rect 486200 298618 487000 298648
rect 478156 298558 487000 298618
rect 478156 298556 478162 298558
rect 486200 298528 487000 298558
rect 0 297938 800 297968
rect 479977 297938 480043 297941
rect 486200 297938 487000 297968
rect 0 297878 10032 297938
rect 479977 297936 487000 297938
rect 479977 297880 479982 297936
rect 480038 297880 487000 297936
rect 479977 297878 487000 297880
rect 0 297848 800 297878
rect 479977 297875 480043 297878
rect 486200 297848 487000 297878
rect 0 297258 800 297288
rect 480069 297258 480135 297261
rect 486200 297258 487000 297288
rect 0 297198 9506 297258
rect 0 297168 800 297198
rect 9446 297190 9506 297198
rect 480069 297256 487000 297258
rect 480069 297200 480074 297256
rect 480130 297200 487000 297256
rect 480069 297198 487000 297200
rect 480069 297195 480135 297198
rect 9446 297130 10060 297190
rect 486200 297168 487000 297198
rect 0 296578 800 296608
rect 480161 296578 480227 296581
rect 486200 296578 487000 296608
rect 0 296518 9506 296578
rect 0 296488 800 296518
rect 9446 296374 9506 296518
rect 480161 296576 487000 296578
rect 480161 296520 480166 296576
rect 480222 296520 487000 296576
rect 480161 296518 487000 296520
rect 480161 296515 480227 296518
rect 486200 296488 487000 296518
rect 9446 296314 10060 296374
rect 486200 295900 487000 295928
rect 486200 295836 486372 295900
rect 486436 295836 487000 295900
rect 486200 295808 487000 295836
rect 9446 295420 10060 295480
rect 9446 295354 9506 295420
rect 6870 295294 9506 295354
rect 0 295218 800 295248
rect 6870 295218 6930 295294
rect 0 295158 6930 295218
rect 0 295128 800 295158
rect 481214 295156 481220 295220
rect 481284 295218 481290 295220
rect 486200 295218 487000 295248
rect 481284 295158 487000 295218
rect 481284 295156 481290 295158
rect 486200 295128 487000 295158
rect 9446 294604 10060 294664
rect 0 294538 800 294568
rect 9446 294538 9506 294604
rect 0 294478 9506 294538
rect 0 294448 800 294478
rect 482318 294476 482324 294540
rect 482388 294538 482394 294540
rect 486200 294538 487000 294568
rect 482388 294478 487000 294538
rect 482388 294476 482394 294478
rect 486200 294448 487000 294478
rect 0 293858 800 293888
rect 0 293798 10032 293858
rect 0 293768 800 293798
rect 482134 293796 482140 293860
rect 482204 293858 482210 293860
rect 486200 293858 487000 293888
rect 482204 293798 487000 293858
rect 482204 293796 482210 293798
rect 486200 293768 487000 293798
rect 0 293178 800 293208
rect 0 293118 9506 293178
rect 0 293088 800 293118
rect 9446 293110 9506 293118
rect 481030 293116 481036 293180
rect 481100 293178 481106 293180
rect 486200 293178 487000 293208
rect 481100 293118 487000 293178
rect 481100 293116 481106 293118
rect 9446 293050 10060 293110
rect 486200 293088 487000 293118
rect 0 292498 800 292528
rect 0 292438 9506 292498
rect 0 292408 800 292438
rect 9446 292294 9506 292438
rect 483974 292436 483980 292500
rect 484044 292498 484050 292500
rect 486200 292498 487000 292528
rect 484044 292438 487000 292498
rect 484044 292436 484050 292438
rect 486200 292408 487000 292438
rect 9446 292234 10060 292294
rect 483790 291756 483796 291820
rect 483860 291818 483866 291820
rect 486200 291818 487000 291848
rect 483860 291758 487000 291818
rect 483860 291756 483866 291758
rect 486200 291728 487000 291758
rect 9446 291340 10060 291400
rect 9446 291274 9506 291340
rect 6870 291214 9506 291274
rect 0 291138 800 291168
rect 6870 291138 6930 291214
rect 0 291078 6930 291138
rect 0 291048 800 291078
rect 483606 291076 483612 291140
rect 483676 291138 483682 291140
rect 486200 291138 487000 291168
rect 483676 291078 487000 291138
rect 483676 291076 483682 291078
rect 486200 291048 487000 291078
rect 480846 290396 480852 290460
rect 480916 290458 480922 290460
rect 486200 290458 487000 290488
rect 480916 290398 487000 290458
rect 480916 290396 480922 290398
rect 486200 290368 487000 290398
rect 482829 289778 482895 289781
rect 486200 289778 487000 289808
rect 482829 289776 487000 289778
rect 482829 289720 482834 289776
rect 482890 289720 487000 289776
rect 482829 289718 487000 289720
rect 482829 289715 482895 289718
rect 486200 289688 487000 289718
rect 484301 289098 484367 289101
rect 486200 289098 487000 289128
rect 484301 289096 487000 289098
rect 484301 289040 484306 289096
rect 484362 289040 487000 289096
rect 484301 289038 487000 289040
rect 484301 289035 484367 289038
rect 486200 289008 487000 289038
rect 481541 288418 481607 288421
rect 486200 288418 487000 288448
rect 481541 288416 487000 288418
rect 481541 288360 481546 288416
rect 481602 288360 487000 288416
rect 481541 288358 487000 288360
rect 481541 288355 481607 288358
rect 486200 288328 487000 288358
rect 482921 287738 482987 287741
rect 486200 287738 487000 287768
rect 482921 287736 487000 287738
rect 482921 287680 482926 287736
rect 482982 287680 487000 287736
rect 482921 287678 487000 287680
rect 482921 287675 482987 287678
rect 486200 287648 487000 287678
rect 481449 287058 481515 287061
rect 486200 287058 487000 287088
rect 481449 287056 487000 287058
rect 481449 287000 481454 287056
rect 481510 287000 487000 287056
rect 481449 286998 487000 287000
rect 481449 286995 481515 286998
rect 486200 286968 487000 286998
rect 6870 283054 10032 283114
rect 0 282978 800 283008
rect 6870 282978 6930 283054
rect 0 282918 6930 282978
rect 0 282888 800 282918
rect 0 282298 800 282328
rect 0 282238 10060 282298
rect 0 282208 800 282238
rect 0 281618 800 281648
rect 0 281558 4170 281618
rect 0 281528 800 281558
rect 4110 281482 4170 281558
rect 4110 281422 10060 281482
rect 0 280938 800 280968
rect 0 280878 6930 280938
rect 0 280848 800 280878
rect 6870 280802 6930 280878
rect 6870 280742 9506 280802
rect 9446 280734 9506 280742
rect 9446 280674 10060 280734
rect 6870 279790 10060 279850
rect 0 279578 800 279608
rect 6870 279578 6930 279790
rect 0 279518 6930 279578
rect 0 279488 800 279518
rect 6870 278974 10060 279034
rect 0 278898 800 278928
rect 6870 278898 6930 278974
rect 0 278838 6930 278898
rect 0 278808 800 278838
rect 0 278218 800 278248
rect 0 278158 10060 278218
rect 0 278128 800 278158
rect 0 277538 800 277568
rect 0 277478 4906 277538
rect 0 277448 800 277478
rect 4846 277402 4906 277478
rect 4846 277342 10060 277402
rect 0 276858 800 276888
rect 0 276798 6930 276858
rect 0 276768 800 276798
rect 6870 276722 6930 276798
rect 6870 276662 9506 276722
rect 9446 276654 9506 276662
rect 9446 276594 10060 276654
rect 6870 275710 10060 275770
rect 0 275498 800 275528
rect 6870 275498 6930 275710
rect 0 275438 6930 275498
rect 0 275408 800 275438
rect 6870 274894 10060 274954
rect 0 274818 800 274848
rect 6870 274818 6930 274894
rect 0 274758 6930 274818
rect 0 274728 800 274758
rect 0 274138 800 274168
rect 0 274078 10060 274138
rect 0 274048 800 274078
rect 0 273458 800 273488
rect 0 273398 9506 273458
rect 0 273368 800 273398
rect 9446 273390 9506 273398
rect 9446 273330 10060 273390
rect 0 272778 800 272808
rect 0 272718 6930 272778
rect 0 272688 800 272718
rect 6870 272642 6930 272718
rect 6870 272582 9506 272642
rect 9446 272574 9506 272582
rect 9446 272514 10060 272574
rect 6870 271630 10060 271690
rect 0 271418 800 271448
rect 6870 271418 6930 271630
rect 0 271358 6930 271418
rect 0 271328 800 271358
rect 6870 270814 10060 270874
rect 0 270738 800 270768
rect 6870 270738 6930 270814
rect 0 270678 6930 270738
rect 0 270648 800 270678
rect 0 270058 800 270088
rect 481541 270058 481607 270061
rect 486200 270058 487000 270088
rect 0 269998 10060 270058
rect 481541 270056 487000 270058
rect 481541 270000 481546 270056
rect 481602 270000 487000 270056
rect 481541 269998 487000 270000
rect 0 269968 800 269998
rect 481541 269995 481607 269998
rect 486200 269968 487000 269998
rect 0 269378 800 269408
rect 482921 269378 482987 269381
rect 486200 269378 487000 269408
rect 0 269318 9506 269378
rect 0 269288 800 269318
rect 9446 269310 9506 269318
rect 482921 269376 487000 269378
rect 482921 269320 482926 269376
rect 482982 269320 487000 269376
rect 482921 269318 487000 269320
rect 482921 269315 482987 269318
rect 9446 269250 10060 269310
rect 486200 269288 487000 269318
rect 0 268698 800 268728
rect 484301 268698 484367 268701
rect 486200 268698 487000 268728
rect 0 268638 6930 268698
rect 0 268608 800 268638
rect 6870 268562 6930 268638
rect 484301 268696 487000 268698
rect 484301 268640 484306 268696
rect 484362 268640 487000 268696
rect 484301 268638 487000 268640
rect 484301 268635 484367 268638
rect 486200 268608 487000 268638
rect 6870 268502 9506 268562
rect 9446 268494 9506 268502
rect 9446 268434 10060 268494
rect 481449 268018 481515 268021
rect 486200 268018 487000 268048
rect 481449 268016 487000 268018
rect 481449 267960 481454 268016
rect 481510 267960 487000 268016
rect 481449 267958 487000 267960
rect 481449 267955 481515 267958
rect 486200 267928 487000 267958
rect 6870 267550 10060 267610
rect 0 267338 800 267368
rect 6870 267338 6930 267550
rect 0 267278 6930 267338
rect 0 267248 800 267278
rect 483606 267276 483612 267340
rect 483676 267338 483682 267340
rect 486200 267338 487000 267368
rect 483676 267278 487000 267338
rect 483676 267276 483682 267278
rect 486200 267248 487000 267278
rect 6870 266734 10060 266794
rect 0 266658 800 266688
rect 6870 266658 6930 266734
rect 0 266598 6930 266658
rect 482829 266658 482895 266661
rect 486200 266658 487000 266688
rect 482829 266656 487000 266658
rect 482829 266600 482834 266656
rect 482890 266600 487000 266656
rect 482829 266598 487000 266600
rect 0 266568 800 266598
rect 482829 266595 482895 266598
rect 486200 266568 487000 266598
rect 0 265978 800 266008
rect 0 265918 10060 265978
rect 0 265888 800 265918
rect 483790 265916 483796 265980
rect 483860 265978 483866 265980
rect 486200 265978 487000 266008
rect 483860 265918 487000 265978
rect 483860 265916 483866 265918
rect 486200 265888 487000 265918
rect 0 265298 800 265328
rect 0 265238 9506 265298
rect 0 265208 800 265238
rect 9446 265230 9506 265238
rect 480846 265236 480852 265300
rect 480916 265298 480922 265300
rect 486200 265298 487000 265328
rect 480916 265238 487000 265298
rect 480916 265236 480922 265238
rect 9446 265170 10060 265230
rect 486200 265208 487000 265238
rect 0 264618 800 264648
rect 478689 264618 478755 264621
rect 486200 264618 487000 264648
rect 0 264558 6930 264618
rect 0 264528 800 264558
rect 6870 264482 6930 264558
rect 478689 264616 487000 264618
rect 478689 264560 478694 264616
rect 478750 264560 487000 264616
rect 478689 264558 487000 264560
rect 478689 264555 478755 264558
rect 486200 264528 487000 264558
rect 6870 264422 9506 264482
rect 9446 264414 9506 264422
rect 9446 264354 10060 264414
rect 478781 263938 478847 263941
rect 486200 263938 487000 263968
rect 478781 263936 487000 263938
rect 478781 263880 478786 263936
rect 478842 263880 487000 263936
rect 478781 263878 487000 263880
rect 478781 263875 478847 263878
rect 486200 263848 487000 263878
rect 6870 263470 10060 263530
rect 0 263258 800 263288
rect 6870 263258 6930 263470
rect 0 263198 6930 263258
rect 478597 263258 478663 263261
rect 486200 263258 487000 263288
rect 478597 263256 487000 263258
rect 478597 263200 478602 263256
rect 478658 263200 487000 263256
rect 478597 263198 487000 263200
rect 0 263168 800 263198
rect 478597 263195 478663 263198
rect 486200 263168 487000 263198
rect 6870 262654 10060 262714
rect 0 262578 800 262608
rect 6870 262578 6930 262654
rect 0 262518 6930 262578
rect 0 262488 800 262518
rect 478086 262516 478092 262580
rect 478156 262578 478162 262580
rect 486200 262578 487000 262608
rect 478156 262518 487000 262578
rect 478156 262516 478162 262518
rect 486200 262488 487000 262518
rect 0 261898 800 261928
rect 0 261838 10060 261898
rect 0 261808 800 261838
rect 482134 261836 482140 261900
rect 482204 261898 482210 261900
rect 486200 261898 487000 261928
rect 482204 261838 487000 261898
rect 482204 261836 482210 261838
rect 486200 261808 487000 261838
rect 0 261218 800 261248
rect 0 261158 9506 261218
rect 0 261128 800 261158
rect 9446 261150 9506 261158
rect 478270 261156 478276 261220
rect 478340 261218 478346 261220
rect 486200 261218 487000 261248
rect 478340 261158 487000 261218
rect 478340 261156 478346 261158
rect 9446 261090 10060 261150
rect 486200 261128 487000 261158
rect 0 260538 800 260568
rect 0 260478 6930 260538
rect 0 260448 800 260478
rect 6870 260402 6930 260478
rect 482318 260476 482324 260540
rect 482388 260538 482394 260540
rect 486200 260538 487000 260568
rect 482388 260478 487000 260538
rect 482388 260476 482394 260478
rect 486200 260448 487000 260478
rect 6870 260342 9506 260402
rect 9446 260334 9506 260342
rect 9446 260274 10060 260334
rect 485630 259796 485636 259860
rect 485700 259858 485706 259860
rect 486200 259858 487000 259888
rect 485700 259798 487000 259858
rect 485700 259796 485706 259798
rect 486200 259768 487000 259798
rect 6870 259390 10060 259450
rect 0 259178 800 259208
rect 6870 259178 6930 259390
rect 0 259118 6930 259178
rect 0 259088 800 259118
rect 481030 259116 481036 259180
rect 481100 259178 481106 259180
rect 486200 259178 487000 259208
rect 481100 259118 487000 259178
rect 481100 259116 481106 259118
rect 486200 259088 487000 259118
rect 6870 258574 10060 258634
rect 0 258498 800 258528
rect 6870 258498 6930 258574
rect 0 258438 6930 258498
rect 0 258408 800 258438
rect 479558 258436 479564 258500
rect 479628 258498 479634 258500
rect 486200 258498 487000 258528
rect 479628 258438 487000 258498
rect 479628 258436 479634 258438
rect 486200 258408 487000 258438
rect 0 257818 800 257848
rect 0 257758 10060 257818
rect 0 257728 800 257758
rect 483974 257756 483980 257820
rect 484044 257818 484050 257820
rect 486200 257818 487000 257848
rect 484044 257758 487000 257818
rect 484044 257756 484050 257758
rect 486200 257728 487000 257758
rect 0 257138 800 257168
rect 0 257078 9506 257138
rect 0 257048 800 257078
rect 9446 257070 9506 257078
rect 485446 257076 485452 257140
rect 485516 257138 485522 257140
rect 486200 257138 487000 257168
rect 485516 257078 487000 257138
rect 485516 257076 485522 257078
rect 9446 257010 10060 257070
rect 486200 257048 487000 257078
rect 0 256458 800 256488
rect 0 256398 6930 256458
rect 0 256368 800 256398
rect 6870 256322 6930 256398
rect 479374 256396 479380 256460
rect 479444 256458 479450 256460
rect 486200 256458 487000 256488
rect 479444 256398 487000 256458
rect 479444 256396 479450 256398
rect 486200 256368 487000 256398
rect 6870 256262 9506 256322
rect 9446 256254 9506 256262
rect 9446 256194 10060 256254
rect 483657 255778 483723 255781
rect 486200 255778 487000 255808
rect 483657 255776 487000 255778
rect 483657 255720 483662 255776
rect 483718 255720 487000 255776
rect 483657 255718 487000 255720
rect 483657 255715 483723 255718
rect 486200 255688 487000 255718
rect 6870 255310 10060 255370
rect 0 255098 800 255128
rect 6870 255098 6930 255310
rect 0 255038 6930 255098
rect 0 255008 800 255038
rect 479742 255036 479748 255100
rect 479812 255098 479818 255100
rect 486200 255098 487000 255128
rect 479812 255038 487000 255098
rect 479812 255036 479818 255038
rect 486200 255008 487000 255038
rect 6870 254494 10060 254554
rect 0 254418 800 254448
rect 6870 254418 6930 254494
rect 0 254358 6930 254418
rect 486200 254420 487000 254448
rect 0 254328 800 254358
rect 486200 254356 486372 254420
rect 486436 254356 487000 254420
rect 486200 254328 487000 254356
rect 0 253738 800 253768
rect 0 253678 10060 253738
rect 0 253648 800 253678
rect 485814 253676 485820 253740
rect 485884 253738 485890 253740
rect 486200 253738 487000 253768
rect 485884 253678 487000 253738
rect 485884 253676 485890 253678
rect 486200 253648 487000 253678
rect 0 253058 800 253088
rect 0 252998 9506 253058
rect 0 252968 800 252998
rect 9446 252990 9506 252998
rect 479926 252996 479932 253060
rect 479996 253058 480002 253060
rect 486200 253058 487000 253088
rect 479996 252998 487000 253058
rect 479996 252996 480002 252998
rect 9446 252930 10060 252990
rect 486200 252968 487000 252998
rect 0 252378 800 252408
rect 0 252318 6930 252378
rect 0 252288 800 252318
rect 6870 252242 6930 252318
rect 481214 252316 481220 252380
rect 481284 252378 481290 252380
rect 486200 252378 487000 252408
rect 481284 252318 487000 252378
rect 481284 252316 481290 252318
rect 486200 252288 487000 252318
rect 6870 252182 9506 252242
rect 9446 252174 9506 252182
rect 9446 252114 10060 252174
rect 485998 251636 486004 251700
rect 486068 251698 486074 251700
rect 486200 251698 487000 251728
rect 486068 251638 487000 251698
rect 486068 251636 486074 251638
rect 486200 251608 487000 251638
rect 6870 251230 10060 251290
rect 0 251018 800 251048
rect 6870 251018 6930 251230
rect 0 250958 6930 251018
rect 0 250928 800 250958
rect 484526 250956 484532 251020
rect 484596 251018 484602 251020
rect 486200 251018 487000 251048
rect 484596 250958 487000 251018
rect 484596 250956 484602 250958
rect 486200 250928 487000 250958
rect 6870 250414 10060 250474
rect 0 250338 800 250368
rect 6870 250338 6930 250414
rect 0 250278 6930 250338
rect 0 250248 800 250278
rect 484710 250276 484716 250340
rect 484780 250338 484786 250340
rect 486200 250338 487000 250368
rect 484780 250278 487000 250338
rect 484780 250276 484786 250278
rect 486200 250248 487000 250278
rect 0 249658 800 249688
rect 0 249598 10060 249658
rect 0 249568 800 249598
rect 481582 249596 481588 249660
rect 481652 249658 481658 249660
rect 486200 249658 487000 249688
rect 481652 249598 487000 249658
rect 481652 249596 481658 249598
rect 486200 249568 487000 249598
rect 0 248978 800 249008
rect 0 248918 9506 248978
rect 0 248888 800 248918
rect 9446 248910 9506 248918
rect 484342 248916 484348 248980
rect 484412 248978 484418 248980
rect 486200 248978 487000 249008
rect 484412 248918 487000 248978
rect 484412 248916 484418 248918
rect 9446 248850 10060 248910
rect 486200 248888 487000 248918
rect 0 248298 800 248328
rect 483197 248298 483263 248301
rect 486200 248298 487000 248328
rect 0 248238 6930 248298
rect 0 248208 800 248238
rect 6870 248162 6930 248238
rect 483197 248296 487000 248298
rect 483197 248240 483202 248296
rect 483258 248240 487000 248296
rect 483197 248238 487000 248240
rect 483197 248235 483263 248238
rect 486200 248208 487000 248238
rect 476940 248162 477418 248184
rect 485998 248162 486004 248164
rect 6870 248102 9506 248162
rect 476940 248124 486004 248162
rect 477358 248102 486004 248124
rect 9446 248094 9506 248102
rect 485998 248100 486004 248102
rect 486068 248100 486074 248164
rect 9446 248034 10060 248094
rect 477534 247964 477540 248028
rect 477604 248026 477610 248028
rect 483197 248026 483263 248029
rect 477604 248024 483263 248026
rect 477604 247968 483202 248024
rect 483258 247968 483263 248024
rect 477604 247966 483263 247968
rect 477604 247964 477610 247966
rect 483197 247963 483263 247966
rect 476940 247890 477418 247912
rect 481214 247890 481220 247892
rect 476940 247852 481220 247890
rect 477358 247830 481220 247852
rect 481214 247828 481220 247830
rect 481284 247828 481290 247892
rect 481582 247754 481588 247756
rect 477358 247696 481588 247754
rect 476940 247694 481588 247696
rect 476940 247636 477418 247694
rect 481582 247692 481588 247694
rect 481652 247692 481658 247756
rect 482870 247556 482876 247620
rect 482940 247618 482946 247620
rect 486200 247618 487000 247648
rect 482940 247558 487000 247618
rect 482940 247556 482946 247558
rect 486200 247528 487000 247558
rect 484342 247482 484348 247484
rect 477358 247424 484348 247482
rect 476940 247422 484348 247424
rect 476940 247364 477418 247422
rect 484342 247420 484348 247422
rect 484412 247420 484418 247484
rect 484710 247210 484716 247212
rect 6870 247150 10060 247210
rect 477358 247152 484716 247210
rect 476940 247150 484716 247152
rect 0 246938 800 246968
rect 6870 246938 6930 247150
rect 476940 247092 477418 247150
rect 484710 247148 484716 247150
rect 484780 247148 484786 247212
rect 477534 247012 477540 247076
rect 477604 247074 477610 247076
rect 478597 247074 478663 247077
rect 477604 247072 478663 247074
rect 477604 247016 478602 247072
rect 478658 247016 478663 247072
rect 477604 247014 478663 247016
rect 477604 247012 477610 247014
rect 478597 247011 478663 247014
rect 480294 247012 480300 247076
rect 480364 247074 480370 247076
rect 481449 247074 481515 247077
rect 480364 247072 481515 247074
rect 480364 247016 481454 247072
rect 481510 247016 481515 247072
rect 480364 247014 481515 247016
rect 480364 247012 480370 247014
rect 481449 247011 481515 247014
rect 481766 247012 481772 247076
rect 481836 247074 481842 247076
rect 482829 247074 482895 247077
rect 481836 247072 482895 247074
rect 481836 247016 482834 247072
rect 482890 247016 482895 247072
rect 481836 247014 482895 247016
rect 481836 247012 481842 247014
rect 482829 247011 482895 247014
rect 0 246878 6930 246938
rect 477166 246880 477172 246882
rect 0 246848 800 246878
rect 476940 246820 477172 246880
rect 477166 246818 477172 246820
rect 477236 246818 477242 246882
rect 477350 246876 477356 246940
rect 477420 246938 477426 246940
rect 486200 246938 487000 246968
rect 477420 246878 487000 246938
rect 477420 246876 477426 246878
rect 486200 246848 487000 246878
rect 484526 246666 484532 246668
rect 477358 246608 484532 246666
rect 476940 246606 484532 246608
rect 476940 246548 477418 246606
rect 484526 246604 484532 246606
rect 484596 246604 484602 246668
rect 9446 246340 10060 246400
rect 479558 246394 479564 246396
rect 0 246258 800 246288
rect 9446 246258 9506 246340
rect 477358 246336 479564 246394
rect 476940 246334 479564 246336
rect 476940 246276 477418 246334
rect 479558 246332 479564 246334
rect 479628 246332 479634 246396
rect 0 246198 9506 246258
rect 0 246168 800 246198
rect 483238 246196 483244 246260
rect 483308 246258 483314 246260
rect 486200 246258 487000 246288
rect 483308 246198 487000 246258
rect 483308 246196 483314 246198
rect 486200 246168 487000 246198
rect 482870 246122 482876 246124
rect 477358 246064 482876 246122
rect 476940 246062 482876 246064
rect 476940 246004 477418 246062
rect 482870 246060 482876 246062
rect 482940 246060 482946 246124
rect 481030 245850 481036 245852
rect 477358 245792 481036 245850
rect 476940 245790 481036 245792
rect 476940 245732 477418 245790
rect 481030 245788 481036 245790
rect 481100 245788 481106 245852
rect 477718 245652 477724 245716
rect 477788 245714 477794 245716
rect 478689 245714 478755 245717
rect 477788 245712 478755 245714
rect 477788 245656 478694 245712
rect 478750 245656 478755 245712
rect 477788 245654 478755 245656
rect 477788 245652 477794 245654
rect 478689 245651 478755 245654
rect 481582 245652 481588 245716
rect 481652 245714 481658 245716
rect 482921 245714 482987 245717
rect 481652 245712 482987 245714
rect 481652 245656 482926 245712
rect 482982 245656 482987 245712
rect 481652 245654 482987 245656
rect 481652 245652 481658 245654
rect 482921 245651 482987 245654
rect 477350 245520 477356 245522
rect 476940 245460 477356 245520
rect 477350 245458 477356 245460
rect 477420 245458 477426 245522
rect 484526 245516 484532 245580
rect 484596 245578 484602 245580
rect 486200 245578 487000 245608
rect 484596 245518 487000 245578
rect 484596 245516 484602 245518
rect 486200 245488 487000 245518
rect 479926 245306 479932 245308
rect 477358 245248 479932 245306
rect 476940 245246 479932 245248
rect 476940 245188 477418 245246
rect 479926 245244 479932 245246
rect 479996 245244 480002 245308
rect 485814 245034 485820 245036
rect 477358 244976 485820 245034
rect 476940 244974 485820 244976
rect 476940 244916 477418 244974
rect 485814 244972 485820 244974
rect 485884 244972 485890 245036
rect 484342 244836 484348 244900
rect 484412 244898 484418 244900
rect 486200 244898 487000 244928
rect 484412 244838 487000 244898
rect 484412 244836 484418 244838
rect 486200 244808 487000 244838
rect 483238 244762 483244 244764
rect 477358 244704 483244 244762
rect 476940 244702 483244 244704
rect 476940 244644 477418 244702
rect 483238 244700 483244 244702
rect 483308 244700 483314 244764
rect 486182 244490 486188 244492
rect 477358 244432 486188 244490
rect 476940 244430 486188 244432
rect 476940 244372 477418 244430
rect 486182 244428 486188 244430
rect 486252 244428 486258 244492
rect 480478 244292 480484 244356
rect 480548 244354 480554 244356
rect 481541 244354 481607 244357
rect 480548 244352 481607 244354
rect 480548 244296 481546 244352
rect 481602 244296 481607 244352
rect 480548 244294 481607 244296
rect 480548 244292 480554 244294
rect 481541 244291 481607 244294
rect 484894 244156 484900 244220
rect 484964 244218 484970 244220
rect 486200 244218 487000 244248
rect 484964 244158 487000 244218
rect 484964 244156 484970 244158
rect 486200 244128 487000 244158
rect 476940 244082 477418 244104
rect 485630 244082 485636 244084
rect 476940 244044 485636 244082
rect 477358 244022 485636 244044
rect 485630 244020 485636 244022
rect 485700 244020 485706 244084
rect 479742 243946 479748 243948
rect 477358 243888 479748 243946
rect 476940 243886 479748 243888
rect 476940 243828 477418 243886
rect 479742 243884 479748 243886
rect 479812 243884 479818 243948
rect 482318 243674 482324 243676
rect 477358 243616 482324 243674
rect 476940 243614 482324 243616
rect 476940 243556 477418 243614
rect 482318 243612 482324 243614
rect 482388 243612 482394 243676
rect 483054 243476 483060 243540
rect 483124 243538 483130 243540
rect 484301 243538 484367 243541
rect 483124 243536 484367 243538
rect 483124 243480 484306 243536
rect 484362 243480 484367 243536
rect 483124 243478 484367 243480
rect 483124 243476 483130 243478
rect 484301 243475 484367 243478
rect 484710 243476 484716 243540
rect 484780 243538 484786 243540
rect 486200 243538 487000 243568
rect 484780 243478 487000 243538
rect 484780 243476 484786 243478
rect 486200 243448 487000 243478
rect 476940 243266 477418 243288
rect 484526 243266 484532 243268
rect 476940 243228 484532 243266
rect 477358 243206 484532 243228
rect 484526 243204 484532 243206
rect 484596 243204 484602 243268
rect 479374 243130 479380 243132
rect 477358 243072 479380 243130
rect 476940 243070 479380 243072
rect 476940 243012 477418 243070
rect 479374 243068 479380 243070
rect 479444 243068 479450 243132
rect 477902 242796 477908 242860
rect 477972 242858 477978 242860
rect 478781 242858 478847 242861
rect 477972 242856 478847 242858
rect 477972 242800 478786 242856
rect 478842 242800 478847 242856
rect 477972 242798 478847 242800
rect 477972 242796 477978 242798
rect 478781 242795 478847 242798
rect 483238 242796 483244 242860
rect 483308 242858 483314 242860
rect 486200 242858 487000 242888
rect 483308 242798 487000 242858
rect 483308 242796 483314 242798
rect 486200 242768 487000 242798
rect 476940 242722 477418 242744
rect 484342 242722 484348 242724
rect 476940 242684 484348 242722
rect 477358 242662 484348 242684
rect 484342 242660 484348 242662
rect 484412 242660 484418 242724
rect 485446 242586 485452 242588
rect 477358 242528 485452 242586
rect 476940 242526 485452 242528
rect 476940 242468 477418 242526
rect 485446 242524 485452 242526
rect 485516 242524 485522 242588
rect 483974 242314 483980 242316
rect 477358 242256 483980 242314
rect 476940 242254 483980 242256
rect 476940 242196 477418 242254
rect 483974 242252 483980 242254
rect 484044 242252 484050 242316
rect 484342 242116 484348 242180
rect 484412 242178 484418 242180
rect 486200 242178 487000 242208
rect 484412 242118 487000 242178
rect 484412 242116 484418 242118
rect 486200 242088 487000 242118
rect 478270 242042 478276 242044
rect 477358 241984 478276 242042
rect 476940 241982 478276 241984
rect 476940 241924 477418 241982
rect 478270 241980 478276 241982
rect 478340 241980 478346 242044
rect 483657 241770 483723 241773
rect 477358 241768 483723 241770
rect 477358 241712 483662 241768
rect 483718 241712 483723 241768
rect 476940 241710 483723 241712
rect 476940 241652 477418 241710
rect 483657 241707 483723 241710
rect 482921 241498 482987 241501
rect 486200 241498 487000 241528
rect 482921 241496 487000 241498
rect 482921 241440 482926 241496
rect 482982 241440 487000 241496
rect 482921 241438 487000 241440
rect 482921 241435 482987 241438
rect 486200 241408 487000 241438
rect 476940 241362 477418 241384
rect 484894 241362 484900 241364
rect 476940 241324 484900 241362
rect 477358 241302 484900 241324
rect 484894 241300 484900 241302
rect 484964 241300 484970 241364
rect 484710 241226 484716 241228
rect 477358 241168 484716 241226
rect 476940 241166 484716 241168
rect 476940 241108 477418 241166
rect 484710 241164 484716 241166
rect 484780 241164 484786 241228
rect 483238 241090 483244 241092
rect 480210 241030 483244 241090
rect 480210 240954 480270 241030
rect 483238 241028 483244 241030
rect 483308 241028 483314 241092
rect 484342 240954 484348 240956
rect 477358 240896 480270 240954
rect 476940 240894 480270 240896
rect 482694 240894 484348 240954
rect 476940 240836 477418 240894
rect 476940 240546 477418 240568
rect 482694 240546 482754 240894
rect 484342 240892 484348 240894
rect 484412 240892 484418 240956
rect 486200 240818 487000 240848
rect 476940 240508 482754 240546
rect 477358 240486 482754 240508
rect 483062 240758 487000 240818
rect 482921 240410 482987 240413
rect 477358 240408 482987 240410
rect 477358 240352 482926 240408
rect 482982 240352 482987 240408
rect 476940 240350 482987 240352
rect 476940 240292 477418 240350
rect 482921 240347 482987 240350
rect 483062 240138 483122 240758
rect 486200 240728 487000 240758
rect 486200 240138 487000 240168
rect 477358 240080 483122 240138
rect 476940 240078 483122 240080
rect 483246 240078 487000 240138
rect 476940 240020 477418 240078
rect 483246 239866 483306 240078
rect 486200 240048 487000 240078
rect 477358 239808 483306 239866
rect 476940 239806 483306 239808
rect 476940 239748 477418 239806
rect 482134 239594 482140 239596
rect 477358 239536 482140 239594
rect 476940 239534 482140 239536
rect 476940 239476 477418 239534
rect 482134 239532 482140 239534
rect 482204 239532 482210 239596
rect 486200 239458 487000 239488
rect 480210 239398 487000 239458
rect 480210 239322 480270 239398
rect 486200 239368 487000 239398
rect 477358 239264 480270 239322
rect 476940 239262 480270 239264
rect 476940 239204 477418 239262
rect 478086 239050 478092 239052
rect 477358 238992 478092 239050
rect 476940 238990 478092 238992
rect 476940 238932 477418 238990
rect 478086 238988 478092 238990
rect 478156 238988 478162 239052
rect 486200 238778 487000 238808
rect 484718 238718 487000 238778
rect 476940 238642 477418 238664
rect 484718 238642 484778 238718
rect 486200 238688 487000 238718
rect 476940 238604 484778 238642
rect 477358 238582 484778 238604
rect 477534 238506 477540 238508
rect 477358 238448 477540 238506
rect 476940 238446 477540 238448
rect 476940 238388 477418 238446
rect 477534 238444 477540 238446
rect 477604 238444 477610 238508
rect 477902 238234 477908 238236
rect 477174 238176 477908 238234
rect 476940 238174 477908 238176
rect 0 238098 800 238128
rect 476940 238116 477234 238174
rect 477902 238172 477908 238174
rect 477972 238172 477978 238236
rect 486200 238098 487000 238128
rect 0 238038 10060 238098
rect 477358 238038 487000 238098
rect 0 238008 800 238038
rect 477358 237904 477418 238038
rect 486200 238008 487000 238038
rect 476940 237844 477418 237904
rect 477718 237690 477724 237692
rect 477358 237632 477724 237690
rect 476940 237630 477724 237632
rect 476940 237572 477418 237630
rect 477718 237628 477724 237630
rect 477788 237628 477794 237692
rect 0 237418 800 237448
rect 486200 237418 487000 237448
rect 0 237358 4170 237418
rect 0 237328 800 237358
rect 4110 237282 4170 237358
rect 484350 237358 487000 237418
rect 476940 237282 477418 237304
rect 484350 237282 484410 237358
rect 486200 237328 487000 237358
rect 4110 237222 10060 237282
rect 476940 237244 484410 237282
rect 477358 237222 484410 237244
rect 480846 237146 480852 237148
rect 477358 237088 480852 237146
rect 476940 237086 480852 237088
rect 476940 237028 477418 237086
rect 480846 237084 480852 237086
rect 480916 237084 480922 237148
rect 483790 236874 483796 236876
rect 477358 236816 483796 236874
rect 476940 236814 483796 236816
rect 0 236738 800 236768
rect 476940 236756 477418 236814
rect 483790 236812 483796 236814
rect 483860 236812 483866 236876
rect 486200 236738 487000 236768
rect 0 236678 9506 236738
rect 0 236648 800 236678
rect 9446 236544 9506 236678
rect 480210 236678 487000 236738
rect 480210 236602 480270 236678
rect 486200 236648 487000 236678
rect 477358 236544 480270 236602
rect 9446 236484 10060 236544
rect 476940 236542 480270 236544
rect 476940 236484 477418 236542
rect 481766 236330 481772 236332
rect 477358 236272 481772 236330
rect 476940 236270 481772 236272
rect 476940 236212 477418 236270
rect 481766 236268 481772 236270
rect 481836 236268 481842 236332
rect 486200 236058 487000 236088
rect 482970 235998 487000 236058
rect 476940 235922 477418 235944
rect 482970 235922 483030 235998
rect 486200 235968 487000 235998
rect 476940 235884 483030 235922
rect 477358 235862 483030 235884
rect 483606 235786 483612 235788
rect 477358 235728 483612 235786
rect 476940 235726 483612 235728
rect 476940 235668 477418 235726
rect 483606 235724 483612 235726
rect 483676 235724 483682 235788
rect 6870 235590 10060 235650
rect 0 235378 800 235408
rect 6870 235378 6930 235590
rect 480294 235514 480300 235516
rect 477358 235456 480300 235514
rect 476940 235454 480300 235456
rect 476940 235396 477418 235454
rect 480294 235452 480300 235454
rect 480364 235452 480370 235516
rect 486200 235378 487000 235408
rect 0 235318 6930 235378
rect 480210 235318 487000 235378
rect 0 235288 800 235318
rect 480210 235242 480270 235318
rect 486200 235288 487000 235318
rect 477358 235184 480270 235242
rect 476940 235182 480270 235184
rect 476940 235124 477418 235182
rect 483054 234970 483060 234972
rect 477358 234912 483060 234970
rect 476940 234910 483060 234912
rect 476940 234852 477418 234910
rect 483054 234908 483060 234910
rect 483124 234908 483130 234972
rect 6870 234774 10060 234834
rect 0 234698 800 234728
rect 6870 234698 6930 234774
rect 486200 234698 487000 234728
rect 0 234638 6930 234698
rect 482970 234638 487000 234698
rect 0 234608 800 234638
rect 476940 234562 477418 234584
rect 482970 234562 483030 234638
rect 486200 234608 487000 234638
rect 476940 234524 483030 234562
rect 477358 234502 483030 234524
rect 481582 234426 481588 234428
rect 477358 234368 481588 234426
rect 476940 234366 481588 234368
rect 476940 234308 477418 234366
rect 481582 234364 481588 234366
rect 481652 234364 481658 234428
rect 480478 234154 480484 234156
rect 477358 234096 480484 234154
rect 476940 234094 480484 234096
rect 0 234018 800 234048
rect 476940 234036 477418 234094
rect 480478 234092 480484 234094
rect 480548 234092 480554 234156
rect 486200 234018 487000 234048
rect 0 233958 10060 234018
rect 480210 233958 487000 234018
rect 0 233928 800 233958
rect 480210 233882 480270 233958
rect 486200 233928 487000 233958
rect 477358 233824 480270 233882
rect 476940 233822 480270 233824
rect 476940 233764 477418 233822
rect 476940 233474 477418 233496
rect 476940 233436 480270 233474
rect 477358 233414 480270 233436
rect 0 233338 800 233368
rect 480210 233338 480270 233414
rect 486200 233338 487000 233368
rect 0 233278 4170 233338
rect 480210 233278 487000 233338
rect 0 233248 800 233278
rect 4110 233202 4170 233278
rect 486200 233248 487000 233278
rect 476940 233202 477418 233224
rect 483054 233202 483060 233204
rect 4110 233142 10060 233202
rect 476940 233164 483060 233202
rect 477358 233142 483060 233164
rect 483054 233140 483060 233142
rect 483124 233140 483130 233204
rect 476940 232930 477418 232952
rect 476940 232892 480270 232930
rect 477358 232870 480270 232892
rect 477718 232794 477724 232796
rect 477174 232736 477724 232794
rect 476940 232734 477724 232736
rect 0 232658 800 232688
rect 476940 232676 477234 232734
rect 477718 232732 477724 232734
rect 477788 232732 477794 232796
rect 480210 232658 480270 232870
rect 486200 232658 487000 232688
rect 0 232598 9506 232658
rect 480210 232598 487000 232658
rect 0 232568 800 232598
rect 9446 232464 9506 232598
rect 486200 232568 487000 232598
rect 9446 232404 10060 232464
rect 476940 232386 477418 232408
rect 477534 232386 477540 232388
rect 476940 232348 477540 232386
rect 477358 232326 477540 232348
rect 477534 232324 477540 232326
rect 477604 232324 477610 232388
rect 476940 232114 477418 232136
rect 476940 232076 480270 232114
rect 477358 232054 480270 232076
rect 480210 231978 480270 232054
rect 486200 231978 487000 232008
rect 480210 231918 487000 231978
rect 486200 231888 487000 231918
rect 476940 231842 477418 231864
rect 480662 231842 480668 231844
rect 476940 231804 480668 231842
rect 477358 231782 480668 231804
rect 480662 231780 480668 231782
rect 480732 231780 480738 231844
rect 483422 231706 483428 231708
rect 477358 231648 483428 231706
rect 476940 231646 483428 231648
rect 476940 231588 477418 231646
rect 483422 231644 483428 231646
rect 483492 231644 483498 231708
rect 6870 231510 10060 231570
rect 0 231298 800 231328
rect 6870 231298 6930 231510
rect 0 231238 6930 231298
rect 476940 231298 477418 231320
rect 486200 231298 487000 231328
rect 476940 231260 487000 231298
rect 477358 231238 487000 231260
rect 0 231208 800 231238
rect 486200 231208 487000 231238
rect 476940 231026 477418 231048
rect 482870 231026 482876 231028
rect 476940 230988 482876 231026
rect 477358 230966 482876 230988
rect 482870 230964 482876 230966
rect 482940 230964 482946 231028
rect 6870 230694 10060 230754
rect 476940 230716 477418 230776
rect 0 230618 800 230648
rect 6870 230618 6930 230694
rect 0 230558 6930 230618
rect 477358 230618 477418 230716
rect 486200 230618 487000 230648
rect 477358 230558 487000 230618
rect 0 230528 800 230558
rect 486200 230528 487000 230558
rect 476940 230482 477050 230504
rect 480846 230482 480852 230484
rect 476940 230444 480852 230482
rect 476990 230422 480852 230444
rect 480846 230420 480852 230422
rect 480916 230420 480922 230484
rect 476940 230210 477418 230232
rect 481582 230210 481588 230212
rect 476940 230172 481588 230210
rect 477358 230150 481588 230172
rect 481582 230148 481588 230150
rect 481652 230148 481658 230212
rect 0 229938 800 229968
rect 476940 229938 477418 229960
rect 486200 229938 487000 229968
rect 0 229878 10060 229938
rect 476940 229900 487000 229938
rect 477358 229878 487000 229900
rect 0 229848 800 229878
rect 486200 229848 487000 229878
rect 483606 229802 483612 229804
rect 477358 229744 483612 229802
rect 476940 229742 483612 229744
rect 476940 229684 477418 229742
rect 483606 229740 483612 229742
rect 483676 229740 483682 229804
rect 477358 229472 483306 229530
rect 476940 229470 483306 229472
rect 476940 229412 477418 229470
rect 0 229258 800 229288
rect 483246 229258 483306 229470
rect 486200 229258 487000 229288
rect 0 229200 9506 229258
rect 0 229198 10060 229200
rect 483246 229198 487000 229258
rect 0 229168 800 229198
rect 9446 229140 10060 229198
rect 486200 229168 487000 229198
rect 476940 229122 477418 229144
rect 483790 229122 483796 229124
rect 476940 229084 483796 229122
rect 477358 229062 483796 229084
rect 483790 229060 483796 229062
rect 483860 229060 483866 229124
rect 476940 228850 477418 228872
rect 482134 228850 482140 228852
rect 476940 228812 482140 228850
rect 477358 228790 482140 228812
rect 482134 228788 482140 228790
rect 482204 228788 482210 228852
rect 0 228578 800 228608
rect 476940 228578 477418 228600
rect 486200 228578 487000 228608
rect 0 228518 9506 228578
rect 476940 228540 487000 228578
rect 477358 228518 487000 228540
rect 0 228488 800 228518
rect 9446 228384 9506 228518
rect 486200 228488 487000 228518
rect 9446 228324 10060 228384
rect 476940 228306 477418 228328
rect 480478 228306 480484 228308
rect 476940 228268 480484 228306
rect 477358 228246 480484 228268
rect 480478 228244 480484 228246
rect 480548 228244 480554 228308
rect 476940 228034 477418 228056
rect 476940 227996 480270 228034
rect 477358 227974 480270 227996
rect 480210 227898 480270 227974
rect 486200 227898 487000 227928
rect 480210 227838 487000 227898
rect 486200 227808 487000 227838
rect 476940 227762 477418 227784
rect 482318 227762 482324 227764
rect 476940 227724 482324 227762
rect 477358 227702 482324 227724
rect 482318 227700 482324 227702
rect 482388 227700 482394 227764
rect 476940 227490 477418 227512
rect 481030 227490 481036 227492
rect 6870 227430 10060 227490
rect 476940 227452 481036 227490
rect 477358 227430 481036 227452
rect 0 227218 800 227248
rect 6870 227218 6930 227430
rect 481030 227428 481036 227430
rect 481100 227428 481106 227492
rect 0 227158 6930 227218
rect 476940 227218 477418 227240
rect 486200 227218 487000 227248
rect 476940 227180 487000 227218
rect 477358 227158 487000 227180
rect 0 227128 800 227158
rect 486200 227128 487000 227158
rect 476940 226946 477418 226968
rect 480110 226946 480116 226948
rect 476940 226908 480116 226946
rect 477358 226886 480116 226908
rect 480110 226884 480116 226886
rect 480180 226884 480186 226948
rect 476940 226674 477418 226696
rect 6870 226614 10060 226674
rect 476940 226636 480270 226674
rect 477358 226614 480270 226636
rect 0 226538 800 226568
rect 6870 226538 6930 226614
rect 0 226478 6930 226538
rect 480210 226538 480270 226614
rect 486200 226538 487000 226568
rect 480210 226478 487000 226538
rect 0 226448 800 226478
rect 486200 226448 487000 226478
rect 476940 226402 477418 226424
rect 476940 226364 480546 226402
rect 477358 226342 480546 226364
rect 480486 226266 480546 226342
rect 480662 226340 480668 226404
rect 480732 226402 480738 226404
rect 481541 226402 481607 226405
rect 480732 226400 481607 226402
rect 480732 226344 481546 226400
rect 481602 226344 481607 226400
rect 480732 226342 481607 226344
rect 480732 226340 480738 226342
rect 481541 226339 481607 226342
rect 481214 226266 481220 226268
rect 480486 226206 481220 226266
rect 481214 226204 481220 226206
rect 481284 226204 481290 226268
rect 476940 226130 477418 226152
rect 486417 226130 486483 226133
rect 476940 226128 486483 226130
rect 476940 226092 486422 226128
rect 477358 226072 486422 226092
rect 486478 226072 486483 226128
rect 477358 226070 486483 226072
rect 486417 226067 486483 226070
rect 0 225858 800 225888
rect 476940 225858 477418 225880
rect 486200 225858 487000 225888
rect 0 225798 10060 225858
rect 476940 225820 487000 225858
rect 477358 225798 487000 225820
rect 0 225768 800 225798
rect 486200 225768 487000 225798
rect 476940 225586 477418 225608
rect 479558 225586 479564 225588
rect 476940 225548 479564 225586
rect 477358 225526 479564 225548
rect 479558 225524 479564 225526
rect 479628 225524 479634 225588
rect 476940 225276 477418 225336
rect 0 225178 800 225208
rect 477358 225178 477418 225276
rect 486200 225178 487000 225208
rect 0 225120 9506 225178
rect 0 225118 10060 225120
rect 477358 225118 487000 225178
rect 0 225088 800 225118
rect 9446 225060 10060 225118
rect 486200 225088 487000 225118
rect 476940 225042 477234 225064
rect 479374 225042 479380 225044
rect 476940 225004 479380 225042
rect 477174 224982 479380 225004
rect 479374 224980 479380 224982
rect 479444 224980 479450 225044
rect 476940 224770 477418 224792
rect 486182 224770 486188 224772
rect 476940 224732 486188 224770
rect 477358 224710 486188 224732
rect 486182 224708 486188 224710
rect 486252 224708 486258 224772
rect 0 224498 800 224528
rect 476940 224498 477418 224520
rect 486200 224498 487000 224528
rect 0 224438 9506 224498
rect 476940 224460 487000 224498
rect 477358 224438 487000 224460
rect 0 224408 800 224438
rect 9446 224304 9506 224438
rect 486200 224408 487000 224438
rect 9446 224244 10060 224304
rect 476940 224226 477418 224248
rect 482502 224226 482508 224228
rect 476940 224188 482508 224226
rect 477358 224166 482508 224188
rect 482502 224164 482508 224166
rect 482572 224164 482578 224228
rect 481449 224090 481515 224093
rect 485446 224090 485452 224092
rect 481449 224088 485452 224090
rect 481449 224032 481454 224088
rect 481510 224032 485452 224088
rect 481449 224030 485452 224032
rect 481449 224027 481515 224030
rect 485446 224028 485452 224030
rect 485516 224028 485522 224092
rect 476940 223954 477418 223976
rect 476940 223916 481650 223954
rect 477358 223894 481650 223916
rect 481449 223818 481515 223821
rect 477358 223816 481515 223818
rect 477358 223760 481454 223816
rect 481510 223760 481515 223816
rect 476940 223758 481515 223760
rect 481590 223818 481650 223894
rect 486200 223818 487000 223848
rect 481590 223758 487000 223818
rect 476940 223700 477418 223758
rect 481449 223755 481515 223758
rect 486200 223728 487000 223758
rect 480161 223684 480227 223685
rect 482921 223684 482987 223685
rect 480110 223682 480116 223684
rect 480070 223622 480116 223682
rect 480180 223680 480227 223684
rect 482870 223682 482876 223684
rect 480222 223624 480227 223680
rect 480110 223620 480116 223622
rect 480180 223620 480227 223624
rect 482830 223622 482876 223682
rect 482940 223680 482987 223684
rect 482982 223624 482987 223680
rect 482870 223620 482876 223622
rect 482940 223620 482987 223624
rect 483054 223620 483060 223684
rect 483124 223682 483130 223684
rect 484301 223682 484367 223685
rect 483124 223680 484367 223682
rect 483124 223624 484306 223680
rect 484362 223624 484367 223680
rect 483124 223622 484367 223624
rect 483124 223620 483130 223622
rect 480161 223619 480227 223620
rect 482921 223619 482987 223620
rect 484301 223619 484367 223622
rect 476940 223410 477418 223432
rect 486182 223410 486188 223412
rect 6870 223350 10060 223410
rect 476940 223372 486188 223410
rect 477358 223350 486188 223372
rect 0 223138 800 223168
rect 6870 223138 6930 223350
rect 486182 223348 486188 223350
rect 486252 223348 486258 223412
rect 0 223078 6930 223138
rect 476940 223138 477418 223160
rect 486200 223138 487000 223168
rect 476940 223100 487000 223138
rect 477358 223078 487000 223100
rect 0 223048 800 223078
rect 486200 223048 487000 223078
rect 476940 222866 477418 222888
rect 483974 222866 483980 222868
rect 476940 222828 483980 222866
rect 477358 222806 483980 222828
rect 483974 222804 483980 222806
rect 484044 222804 484050 222868
rect 476940 222594 477418 222616
rect 6870 222534 10060 222594
rect 476940 222556 481650 222594
rect 477358 222534 481650 222556
rect 0 222458 800 222488
rect 6870 222458 6930 222534
rect 0 222398 6930 222458
rect 481590 222458 481650 222534
rect 486200 222458 487000 222488
rect 481590 222398 487000 222458
rect 0 222368 800 222398
rect 486200 222368 487000 222398
rect 476940 222322 477418 222344
rect 476940 222284 483306 222322
rect 477358 222262 483306 222284
rect 483246 222186 483306 222262
rect 483422 222260 483428 222324
rect 483492 222322 483498 222324
rect 484209 222322 484275 222325
rect 485998 222322 486004 222324
rect 483492 222320 484275 222322
rect 483492 222264 484214 222320
rect 484270 222264 484275 222320
rect 483492 222262 484275 222264
rect 483492 222260 483498 222262
rect 484209 222259 484275 222262
rect 484350 222262 486004 222322
rect 484350 222186 484410 222262
rect 485998 222260 486004 222262
rect 486068 222260 486074 222324
rect 483246 222126 484410 222186
rect 476940 222050 477418 222072
rect 485262 222050 485268 222052
rect 476940 222012 485268 222050
rect 477358 221990 485268 222012
rect 485262 221988 485268 221990
rect 485332 221988 485338 222052
rect 0 221778 800 221808
rect 476940 221778 477418 221800
rect 486200 221778 487000 221808
rect 0 221718 10060 221778
rect 476940 221740 487000 221778
rect 477358 221718 487000 221740
rect 0 221688 800 221718
rect 486200 221688 487000 221718
rect 476940 221506 477418 221528
rect 485078 221506 485084 221508
rect 476940 221468 485084 221506
rect 477358 221446 485084 221468
rect 485078 221444 485084 221446
rect 485148 221444 485154 221508
rect 481449 221370 481515 221373
rect 484710 221370 484716 221372
rect 481449 221368 484716 221370
rect 481449 221312 481454 221368
rect 481510 221312 484716 221368
rect 481449 221310 484716 221312
rect 481449 221307 481515 221310
rect 484710 221308 484716 221310
rect 484780 221308 484786 221372
rect 476940 221234 477418 221256
rect 476940 221196 481650 221234
rect 477358 221174 481650 221196
rect 0 221098 800 221128
rect 481449 221098 481515 221101
rect 0 221040 9506 221098
rect 477358 221096 481515 221098
rect 477358 221040 481454 221096
rect 481510 221040 481515 221096
rect 0 221038 10060 221040
rect 0 221008 800 221038
rect 9446 220980 10060 221038
rect 476940 221038 481515 221040
rect 481590 221098 481650 221174
rect 486200 221098 487000 221128
rect 481590 221038 487000 221098
rect 476940 220980 477418 221038
rect 481449 221035 481515 221038
rect 486200 221008 487000 221038
rect 477718 220900 477724 220964
rect 477788 220962 477794 220964
rect 478781 220962 478847 220965
rect 477788 220960 478847 220962
rect 477788 220904 478786 220960
rect 478842 220904 478847 220960
rect 477788 220902 478847 220904
rect 477788 220900 477794 220902
rect 478781 220899 478847 220902
rect 481030 220900 481036 220964
rect 481100 220962 481106 220964
rect 481449 220962 481515 220965
rect 481100 220960 481515 220962
rect 481100 220904 481454 220960
rect 481510 220904 481515 220960
rect 481100 220902 481515 220904
rect 481100 220900 481106 220902
rect 481449 220899 481515 220902
rect 481582 220900 481588 220964
rect 481652 220962 481658 220964
rect 482829 220962 482895 220965
rect 481652 220960 482895 220962
rect 481652 220904 482834 220960
rect 482890 220904 482895 220960
rect 481652 220902 482895 220904
rect 481652 220900 481658 220902
rect 482829 220899 482895 220902
rect 476940 220690 477418 220712
rect 484526 220690 484532 220692
rect 476940 220652 484532 220690
rect 477358 220630 484532 220652
rect 484526 220628 484532 220630
rect 484596 220628 484602 220692
rect 0 220418 800 220448
rect 476940 220418 477418 220440
rect 486200 220418 487000 220448
rect 0 220358 9506 220418
rect 476940 220380 487000 220418
rect 477358 220358 487000 220380
rect 0 220328 800 220358
rect 9446 220224 9506 220358
rect 486200 220328 487000 220358
rect 9446 220164 10060 220224
rect 476940 220146 477418 220168
rect 484342 220146 484348 220148
rect 476940 220108 484348 220146
rect 477358 220086 484348 220108
rect 484342 220084 484348 220086
rect 484412 220084 484418 220148
rect 480478 219948 480484 220012
rect 480548 220010 480554 220012
rect 481030 220010 481036 220012
rect 480548 219950 481036 220010
rect 480548 219948 480554 219950
rect 481030 219948 481036 219950
rect 481100 219948 481106 220012
rect 476940 219874 477418 219896
rect 476940 219836 481650 219874
rect 477358 219814 481650 219836
rect 481590 219738 481650 219814
rect 486200 219738 487000 219768
rect 481590 219678 487000 219738
rect 486200 219648 487000 219678
rect 476940 219602 477418 219624
rect 483054 219602 483060 219604
rect 476940 219564 483060 219602
rect 477358 219542 483060 219564
rect 483054 219540 483060 219542
rect 483124 219540 483130 219604
rect 477401 219352 477467 219355
rect 476940 219350 477467 219352
rect 6870 219270 10060 219330
rect 476940 219294 477406 219350
rect 477462 219294 477467 219350
rect 476940 219292 477467 219294
rect 477401 219289 477467 219292
rect 0 219058 800 219088
rect 6870 219058 6930 219270
rect 477534 219268 477540 219332
rect 477604 219330 477610 219332
rect 478689 219330 478755 219333
rect 477604 219328 478755 219330
rect 477604 219272 478694 219328
rect 478750 219272 478755 219328
rect 477604 219270 478755 219272
rect 477604 219268 477610 219270
rect 478689 219267 478755 219270
rect 0 218998 6930 219058
rect 476940 219058 477418 219080
rect 486200 219058 487000 219088
rect 476940 219020 487000 219058
rect 477358 218998 487000 219020
rect 0 218968 800 218998
rect 486200 218968 487000 218998
rect 481398 218786 481404 218788
rect 476940 218726 481404 218786
rect 481398 218724 481404 218726
rect 481468 218724 481474 218788
rect 6870 218454 10060 218514
rect 0 218378 800 218408
rect 6870 218378 6930 218454
rect 0 218318 6930 218378
rect 477401 218378 477467 218381
rect 486200 218378 487000 218408
rect 477401 218376 487000 218378
rect 477401 218320 477406 218376
rect 477462 218320 487000 218376
rect 477401 218318 487000 218320
rect 0 218288 800 218318
rect 477401 218315 477467 218318
rect 486200 218288 487000 218318
rect 0 217698 800 217728
rect 0 217638 10060 217698
rect 0 217608 800 217638
rect 483054 217636 483060 217700
rect 483124 217698 483130 217700
rect 486200 217698 487000 217728
rect 483124 217638 487000 217698
rect 483124 217636 483130 217638
rect 486200 217608 487000 217638
rect 0 217018 800 217048
rect 0 216960 9506 217018
rect 0 216958 10060 216960
rect 0 216928 800 216958
rect 9446 216900 10060 216958
rect 484342 216956 484348 217020
rect 484412 217018 484418 217020
rect 486200 217018 487000 217048
rect 484412 216958 487000 217018
rect 484412 216956 484418 216958
rect 486200 216928 487000 216958
rect 0 216338 800 216368
rect 0 216278 9506 216338
rect 0 216248 800 216278
rect 9446 216144 9506 216278
rect 484526 216276 484532 216340
rect 484596 216338 484602 216340
rect 486200 216338 487000 216368
rect 484596 216278 487000 216338
rect 484596 216276 484602 216278
rect 486200 216248 487000 216278
rect 9446 216084 10060 216144
rect 484710 215596 484716 215660
rect 484780 215658 484786 215660
rect 486200 215658 487000 215688
rect 484780 215598 487000 215658
rect 484780 215596 484786 215598
rect 486200 215568 487000 215598
rect 6870 215190 10060 215250
rect 0 214978 800 215008
rect 6870 214978 6930 215190
rect 0 214918 6930 214978
rect 0 214888 800 214918
rect 485078 214916 485084 214980
rect 485148 214978 485154 214980
rect 486200 214978 487000 215008
rect 485148 214918 487000 214978
rect 485148 214916 485154 214918
rect 486200 214888 487000 214918
rect 6870 214374 10060 214434
rect 0 214298 800 214328
rect 6870 214298 6930 214374
rect 0 214238 6930 214298
rect 0 214208 800 214238
rect 485262 214236 485268 214300
rect 485332 214298 485338 214300
rect 486200 214298 487000 214328
rect 485332 214238 487000 214298
rect 485332 214236 485338 214238
rect 486200 214208 487000 214238
rect 0 213618 800 213648
rect 0 213558 10060 213618
rect 0 213528 800 213558
rect 485998 213556 486004 213620
rect 486068 213618 486074 213620
rect 486200 213618 487000 213648
rect 486068 213558 487000 213618
rect 486068 213556 486074 213558
rect 486200 213528 487000 213558
rect 483974 212876 483980 212940
rect 484044 212938 484050 212940
rect 486200 212938 487000 212968
rect 484044 212878 487000 212938
rect 484044 212876 484050 212878
rect 486200 212848 487000 212878
rect 6870 212742 10060 212802
rect 0 212258 800 212288
rect 6870 212258 6930 212742
rect 0 212198 6930 212258
rect 486200 212260 487000 212288
rect 0 212168 800 212198
rect 486200 212196 486372 212260
rect 486436 212196 487000 212260
rect 486200 212168 487000 212196
rect 6870 211926 10060 211986
rect 0 211578 800 211608
rect 6870 211578 6930 211926
rect 0 211518 6930 211578
rect 0 211488 800 211518
rect 485446 211516 485452 211580
rect 485516 211578 485522 211580
rect 486200 211578 487000 211608
rect 485516 211518 487000 211578
rect 485516 211516 485522 211518
rect 486200 211488 487000 211518
rect 6870 211110 10060 211170
rect 0 210898 800 210928
rect 6870 210898 6930 211110
rect 0 210838 6930 210898
rect 0 210808 800 210838
rect 482502 210836 482508 210900
rect 482572 210898 482578 210900
rect 486200 210898 487000 210928
rect 482572 210838 487000 210898
rect 482572 210836 482578 210838
rect 486200 210808 487000 210838
rect 6870 210294 10060 210354
rect 0 210218 800 210248
rect 6870 210218 6930 210294
rect 0 210158 6930 210218
rect 486200 210220 487000 210248
rect 0 210128 800 210158
rect 486200 210156 486556 210220
rect 486620 210156 487000 210220
rect 486200 210128 487000 210156
rect 0 209538 800 209568
rect 0 209478 10060 209538
rect 0 209448 800 209478
rect 479374 209476 479380 209540
rect 479444 209538 479450 209540
rect 486200 209538 487000 209568
rect 479444 209478 487000 209538
rect 479444 209476 479450 209478
rect 486200 209448 487000 209478
rect 0 208858 800 208888
rect 0 208800 9506 208858
rect 0 208798 10060 208800
rect 0 208768 800 208798
rect 9446 208740 10060 208798
rect 479558 208796 479564 208860
rect 479628 208858 479634 208860
rect 486200 208858 487000 208888
rect 479628 208798 487000 208858
rect 479628 208796 479634 208798
rect 486200 208768 487000 208798
rect 0 208178 800 208208
rect 486200 208181 487000 208208
rect 0 208118 9506 208178
rect 0 208088 800 208118
rect 9446 207984 9506 208118
rect 486141 208176 487000 208181
rect 486141 208120 486146 208176
rect 486202 208120 487000 208176
rect 486141 208115 487000 208120
rect 486200 208088 487000 208115
rect 9446 207924 10060 207984
rect 481214 207436 481220 207500
rect 481284 207498 481290 207500
rect 486200 207498 487000 207528
rect 481284 207438 487000 207498
rect 481284 207436 481290 207438
rect 486200 207408 487000 207438
rect 6870 207030 10060 207090
rect 0 206818 800 206848
rect 6870 206818 6930 207030
rect 0 206758 6930 206818
rect 480161 206818 480227 206821
rect 486200 206818 487000 206848
rect 480161 206816 487000 206818
rect 480161 206760 480166 206816
rect 480222 206760 487000 206816
rect 480161 206758 487000 206760
rect 0 206728 800 206758
rect 480161 206755 480227 206758
rect 486200 206728 487000 206758
rect 6870 206214 10060 206274
rect 0 206138 800 206168
rect 6870 206138 6930 206214
rect 0 206078 6930 206138
rect 0 206048 800 206078
rect 481398 206076 481404 206140
rect 481468 206138 481474 206140
rect 486200 206138 487000 206168
rect 481468 206078 487000 206138
rect 481468 206076 481474 206078
rect 486200 206048 487000 206078
rect 0 205458 800 205488
rect 0 205398 10060 205458
rect 0 205368 800 205398
rect 482318 205396 482324 205460
rect 482388 205458 482394 205460
rect 486200 205458 487000 205488
rect 482388 205398 487000 205458
rect 482388 205396 482394 205398
rect 486200 205368 487000 205398
rect 0 204778 800 204808
rect 0 204720 9506 204778
rect 0 204718 10060 204720
rect 0 204688 800 204718
rect 9446 204660 10060 204718
rect 481030 204716 481036 204780
rect 481100 204778 481106 204780
rect 486200 204778 487000 204808
rect 481100 204718 487000 204778
rect 481100 204716 481106 204718
rect 486200 204688 487000 204718
rect 0 204098 800 204128
rect 0 204038 9506 204098
rect 0 204008 800 204038
rect 9446 203904 9506 204038
rect 482134 204036 482140 204100
rect 482204 204098 482210 204100
rect 486200 204098 487000 204128
rect 482204 204038 487000 204098
rect 482204 204036 482210 204038
rect 486200 204008 487000 204038
rect 9446 203844 10060 203904
rect 483790 203356 483796 203420
rect 483860 203418 483866 203420
rect 486200 203418 487000 203448
rect 483860 203358 487000 203418
rect 483860 203356 483866 203358
rect 486200 203328 487000 203358
rect 6870 202950 10060 203010
rect 0 202738 800 202768
rect 6870 202738 6930 202950
rect 0 202678 6930 202738
rect 0 202648 800 202678
rect 483606 202676 483612 202740
rect 483676 202738 483682 202740
rect 486200 202738 487000 202768
rect 483676 202678 487000 202738
rect 483676 202676 483682 202678
rect 486200 202648 487000 202678
rect 6870 202134 10060 202194
rect 0 202058 800 202088
rect 6870 202058 6930 202134
rect 0 201998 6930 202058
rect 482829 202058 482895 202061
rect 486200 202058 487000 202088
rect 482829 202056 487000 202058
rect 482829 202000 482834 202056
rect 482890 202000 487000 202056
rect 482829 201998 487000 202000
rect 0 201968 800 201998
rect 482829 201995 482895 201998
rect 486200 201968 487000 201998
rect 0 201378 800 201408
rect 9446 201378 10060 201400
rect 0 201340 10060 201378
rect 0 201318 9506 201340
rect 0 201288 800 201318
rect 480846 201316 480852 201380
rect 480916 201378 480922 201380
rect 486200 201378 487000 201408
rect 480916 201318 487000 201378
rect 480916 201316 480922 201318
rect 486200 201288 487000 201318
rect 482921 200698 482987 200701
rect 486200 200698 487000 200728
rect 482921 200696 487000 200698
rect 482921 200640 482926 200696
rect 482982 200640 487000 200696
rect 482921 200638 487000 200640
rect 482921 200635 482987 200638
rect 486200 200608 487000 200638
rect 484209 200018 484275 200021
rect 486200 200018 487000 200048
rect 484209 200016 487000 200018
rect 484209 199960 484214 200016
rect 484270 199960 487000 200016
rect 484209 199958 487000 199960
rect 484209 199955 484275 199958
rect 486200 199928 487000 199958
rect 481541 199338 481607 199341
rect 486200 199338 487000 199368
rect 481541 199336 487000 199338
rect 481541 199280 481546 199336
rect 481602 199280 487000 199336
rect 481541 199278 487000 199280
rect 481541 199275 481607 199278
rect 486200 199248 487000 199278
rect 478689 198658 478755 198661
rect 486200 198658 487000 198688
rect 478689 198656 487000 198658
rect 478689 198600 478694 198656
rect 478750 198600 487000 198656
rect 478689 198598 487000 198600
rect 478689 198595 478755 198598
rect 486200 198568 487000 198598
rect 478781 197978 478847 197981
rect 486200 197978 487000 198008
rect 478781 197976 487000 197978
rect 478781 197920 478786 197976
rect 478842 197920 487000 197976
rect 478781 197918 487000 197920
rect 478781 197915 478847 197918
rect 486200 197888 487000 197918
rect 484301 197298 484367 197301
rect 486200 197298 487000 197328
rect 484301 197296 487000 197298
rect 484301 197240 484306 197296
rect 484362 197240 487000 197296
rect 484301 197238 487000 197240
rect 484301 197235 484367 197238
rect 486200 197208 487000 197238
rect 481449 196618 481515 196621
rect 486200 196618 487000 196648
rect 481449 196616 487000 196618
rect 481449 196560 481454 196616
rect 481510 196560 487000 196616
rect 481449 196558 487000 196560
rect 481449 196555 481515 196558
rect 486200 196528 487000 196558
rect 0 193218 800 193248
rect 0 193176 9506 193218
rect 0 193158 10032 193176
rect 0 193128 800 193158
rect 9446 193116 10032 193158
rect 0 192538 800 192568
rect 482921 192538 482987 192541
rect 486200 192538 487000 192568
rect 0 192478 9506 192538
rect 0 192448 800 192478
rect 9446 192360 9506 192478
rect 482921 192536 487000 192538
rect 482921 192480 482926 192536
rect 482982 192480 487000 192536
rect 482921 192478 487000 192480
rect 482921 192475 482987 192478
rect 486200 192448 487000 192478
rect 9446 192300 10032 192360
rect 478137 191858 478203 191861
rect 486200 191858 487000 191888
rect 478137 191856 487000 191858
rect 478137 191800 478142 191856
rect 478198 191800 487000 191856
rect 478137 191798 487000 191800
rect 478137 191795 478203 191798
rect 486200 191768 487000 191798
rect 9446 191428 10032 191488
rect 0 191178 800 191208
rect 9446 191178 9506 191428
rect 0 191118 9506 191178
rect 484025 191178 484091 191181
rect 486200 191178 487000 191208
rect 484025 191176 487000 191178
rect 484025 191120 484030 191176
rect 484086 191120 487000 191176
rect 484025 191118 487000 191120
rect 0 191088 800 191118
rect 484025 191115 484091 191118
rect 486200 191088 487000 191118
rect 9446 190612 10032 190672
rect 0 190498 800 190528
rect 9446 190498 9506 190612
rect 0 190438 9506 190498
rect 480161 190498 480227 190501
rect 486200 190498 487000 190528
rect 480161 190496 487000 190498
rect 480161 190440 480166 190496
rect 480222 190440 487000 190496
rect 480161 190438 487000 190440
rect 0 190408 800 190438
rect 480161 190435 480227 190438
rect 486200 190408 487000 190438
rect 0 189818 800 189848
rect 9446 189818 10032 189856
rect 0 189796 10032 189818
rect 479517 189818 479583 189821
rect 486200 189818 487000 189848
rect 479517 189816 487000 189818
rect 0 189758 9506 189796
rect 479517 189760 479522 189816
rect 479578 189760 487000 189816
rect 479517 189758 487000 189760
rect 0 189728 800 189758
rect 479517 189755 479583 189758
rect 486200 189728 487000 189758
rect 0 189138 800 189168
rect 484301 189138 484367 189141
rect 486200 189138 487000 189168
rect 0 189078 4170 189138
rect 0 189048 800 189078
rect 4110 189002 4170 189078
rect 484301 189136 487000 189138
rect 484301 189080 484306 189136
rect 484362 189080 487000 189136
rect 484301 189078 487000 189080
rect 484301 189075 484367 189078
rect 486200 189048 487000 189078
rect 9446 189002 10032 189040
rect 4110 188980 10032 189002
rect 4110 188942 9506 188980
rect 0 188458 800 188488
rect 482829 188458 482895 188461
rect 486200 188458 487000 188488
rect 0 188398 9506 188458
rect 0 188368 800 188398
rect 9446 188280 9506 188398
rect 482829 188456 487000 188458
rect 482829 188400 482834 188456
rect 482890 188400 487000 188456
rect 482829 188398 487000 188400
rect 482829 188395 482895 188398
rect 486200 188368 487000 188398
rect 9446 188220 10032 188280
rect 484209 187778 484275 187781
rect 486200 187778 487000 187808
rect 484209 187776 487000 187778
rect 484209 187720 484214 187776
rect 484270 187720 487000 187776
rect 484209 187718 487000 187720
rect 484209 187715 484275 187718
rect 486200 187688 487000 187718
rect 9446 187348 10032 187408
rect 0 187098 800 187128
rect 9446 187098 9506 187348
rect 0 187038 9506 187098
rect 482737 187098 482803 187101
rect 486200 187098 487000 187128
rect 482737 187096 487000 187098
rect 482737 187040 482742 187096
rect 482798 187040 487000 187096
rect 482737 187038 487000 187040
rect 0 187008 800 187038
rect 482737 187035 482803 187038
rect 486200 187008 487000 187038
rect 9446 186532 10032 186592
rect 0 186418 800 186448
rect 9446 186418 9506 186532
rect 0 186358 9506 186418
rect 484117 186418 484183 186421
rect 486200 186418 487000 186448
rect 484117 186416 487000 186418
rect 484117 186360 484122 186416
rect 484178 186360 487000 186416
rect 484117 186358 487000 186360
rect 0 186328 800 186358
rect 484117 186355 484183 186358
rect 486200 186328 487000 186358
rect 0 185738 800 185768
rect 9446 185738 10032 185776
rect 0 185716 10032 185738
rect 478689 185738 478755 185741
rect 486200 185738 487000 185768
rect 478689 185736 487000 185738
rect 0 185678 9506 185716
rect 478689 185680 478694 185736
rect 478750 185680 487000 185736
rect 478689 185678 487000 185680
rect 0 185648 800 185678
rect 478689 185675 478755 185678
rect 486200 185648 487000 185678
rect 0 185058 800 185088
rect 478781 185058 478847 185061
rect 486200 185058 487000 185088
rect 0 185016 9506 185058
rect 478781 185056 487000 185058
rect 0 184998 10032 185016
rect 0 184968 800 184998
rect 9446 184956 10032 184998
rect 478781 185000 478786 185056
rect 478842 185000 487000 185056
rect 478781 184998 487000 185000
rect 478781 184995 478847 184998
rect 486200 184968 487000 184998
rect 0 184378 800 184408
rect 478597 184378 478663 184381
rect 486200 184378 487000 184408
rect 0 184318 9506 184378
rect 0 184288 800 184318
rect 9446 184200 9506 184318
rect 478597 184376 487000 184378
rect 478597 184320 478602 184376
rect 478658 184320 487000 184376
rect 478597 184318 487000 184320
rect 478597 184315 478663 184318
rect 486200 184288 487000 184318
rect 9446 184140 10032 184200
rect 480897 183698 480963 183701
rect 486200 183698 487000 183728
rect 480897 183696 487000 183698
rect 480897 183640 480902 183696
rect 480958 183640 487000 183696
rect 480897 183638 487000 183640
rect 480897 183635 480963 183638
rect 486200 183608 487000 183638
rect 9446 183268 10032 183328
rect 0 183018 800 183048
rect 9446 183018 9506 183268
rect 0 182958 9506 183018
rect 480989 183018 481055 183021
rect 486200 183018 487000 183048
rect 480989 183016 487000 183018
rect 480989 182960 480994 183016
rect 481050 182960 487000 183016
rect 480989 182958 487000 182960
rect 0 182928 800 182958
rect 480989 182955 481055 182958
rect 486200 182928 487000 182958
rect 9446 182452 10032 182512
rect 0 182338 800 182368
rect 9446 182338 9506 182452
rect 0 182278 9506 182338
rect 481541 182338 481607 182341
rect 486200 182338 487000 182368
rect 481541 182336 487000 182338
rect 481541 182280 481546 182336
rect 481602 182280 487000 182336
rect 481541 182278 487000 182280
rect 0 182248 800 182278
rect 481541 182275 481607 182278
rect 486200 182248 487000 182278
rect 0 181658 800 181688
rect 9446 181658 10032 181696
rect 0 181636 10032 181658
rect 0 181598 9506 181636
rect 0 181568 800 181598
rect 482134 181596 482140 181660
rect 482204 181658 482210 181660
rect 486200 181658 487000 181688
rect 482204 181598 487000 181658
rect 482204 181596 482210 181598
rect 486200 181568 487000 181598
rect 0 180978 800 181008
rect 478505 180978 478571 180981
rect 486200 180978 487000 181008
rect 0 180936 9506 180978
rect 478505 180976 487000 180978
rect 0 180918 10032 180936
rect 0 180888 800 180918
rect 9446 180876 10032 180918
rect 478505 180920 478510 180976
rect 478566 180920 487000 180976
rect 478505 180918 487000 180920
rect 478505 180915 478571 180918
rect 486200 180888 487000 180918
rect 0 180298 800 180328
rect 0 180238 9506 180298
rect 0 180208 800 180238
rect 9446 180120 9506 180238
rect 478270 180236 478276 180300
rect 478340 180298 478346 180300
rect 486200 180298 487000 180328
rect 478340 180238 487000 180298
rect 478340 180236 478346 180238
rect 486200 180208 487000 180238
rect 9446 180060 10032 180120
rect 482645 179618 482711 179621
rect 486200 179618 487000 179648
rect 482645 179616 487000 179618
rect 482645 179560 482650 179616
rect 482706 179560 487000 179616
rect 482645 179558 487000 179560
rect 482645 179555 482711 179558
rect 486200 179528 487000 179558
rect 9446 179188 10032 179248
rect 0 178938 800 178968
rect 9446 178938 9506 179188
rect 0 178878 9506 178938
rect 483933 178938 483999 178941
rect 486200 178938 487000 178968
rect 483933 178936 487000 178938
rect 483933 178880 483938 178936
rect 483994 178880 487000 178936
rect 483933 178878 487000 178880
rect 0 178848 800 178878
rect 483933 178875 483999 178878
rect 486200 178848 487000 178878
rect 9446 178372 10032 178432
rect 0 178258 800 178288
rect 9446 178258 9506 178372
rect 486200 178261 487000 178288
rect 0 178198 9506 178258
rect 486141 178256 487000 178261
rect 486141 178200 486146 178256
rect 486202 178200 487000 178256
rect 0 178168 800 178198
rect 486141 178195 487000 178200
rect 486200 178168 487000 178195
rect 0 177578 800 177608
rect 9446 177578 10032 177616
rect 0 177556 10032 177578
rect 479977 177578 480043 177581
rect 486200 177578 487000 177608
rect 479977 177576 487000 177578
rect 0 177518 9506 177556
rect 479977 177520 479982 177576
rect 480038 177520 487000 177576
rect 479977 177518 487000 177520
rect 0 177488 800 177518
rect 479977 177515 480043 177518
rect 486200 177488 487000 177518
rect 0 176898 800 176928
rect 480069 176898 480135 176901
rect 486200 176898 487000 176928
rect 0 176856 9506 176898
rect 480069 176896 487000 176898
rect 0 176838 10032 176856
rect 0 176808 800 176838
rect 9446 176796 10032 176838
rect 480069 176840 480074 176896
rect 480130 176840 487000 176896
rect 480069 176838 487000 176840
rect 480069 176835 480135 176838
rect 486200 176808 487000 176838
rect 0 176218 800 176248
rect 479885 176218 479951 176221
rect 486200 176218 487000 176248
rect 0 176158 9506 176218
rect 0 176128 800 176158
rect 9446 176040 9506 176158
rect 479885 176216 487000 176218
rect 479885 176160 479890 176216
rect 479946 176160 487000 176216
rect 479885 176158 487000 176160
rect 479885 176155 479951 176158
rect 486200 176128 487000 176158
rect 9446 175980 10032 176040
rect 481449 175538 481515 175541
rect 486200 175538 487000 175568
rect 481449 175536 487000 175538
rect 481449 175480 481454 175536
rect 481510 175480 487000 175536
rect 481449 175478 487000 175480
rect 481449 175475 481515 175478
rect 486200 175448 487000 175478
rect 9446 175108 10032 175168
rect 0 174858 800 174888
rect 9446 174858 9506 175108
rect 0 174798 9506 174858
rect 0 174768 800 174798
rect 479374 174796 479380 174860
rect 479444 174858 479450 174860
rect 486200 174858 487000 174888
rect 479444 174798 487000 174858
rect 479444 174796 479450 174798
rect 486200 174768 487000 174798
rect 9446 174292 10032 174352
rect 0 174178 800 174208
rect 9446 174178 9506 174292
rect 0 174118 9506 174178
rect 0 174088 800 174118
rect 478086 174116 478092 174180
rect 478156 174178 478162 174180
rect 486200 174178 487000 174208
rect 478156 174118 487000 174178
rect 478156 174116 478162 174118
rect 486200 174088 487000 174118
rect 0 173498 800 173528
rect 9446 173498 10032 173536
rect 0 173476 10032 173498
rect 0 173438 9506 173476
rect 0 173408 800 173438
rect 483606 173436 483612 173500
rect 483676 173498 483682 173500
rect 486200 173498 487000 173528
rect 483676 173438 487000 173498
rect 483676 173436 483682 173438
rect 486200 173408 487000 173438
rect 0 172818 800 172848
rect 0 172776 9506 172818
rect 0 172758 10032 172776
rect 0 172728 800 172758
rect 9446 172716 10032 172758
rect 479558 172756 479564 172820
rect 479628 172818 479634 172820
rect 486200 172818 487000 172848
rect 479628 172758 487000 172818
rect 479628 172756 479634 172758
rect 486200 172728 487000 172758
rect 0 172138 800 172168
rect 0 172078 9506 172138
rect 0 172048 800 172078
rect 9446 171960 9506 172078
rect 482318 172076 482324 172140
rect 482388 172138 482394 172140
rect 486200 172138 487000 172168
rect 482388 172078 487000 172138
rect 482388 172076 482394 172078
rect 486200 172048 487000 172078
rect 9446 171900 10032 171960
rect 477902 171396 477908 171460
rect 477972 171458 477978 171460
rect 486200 171458 487000 171488
rect 477972 171398 487000 171458
rect 477972 171396 477978 171398
rect 486200 171368 487000 171398
rect 9446 171028 10032 171088
rect 0 170778 800 170808
rect 9446 170778 9506 171028
rect 0 170718 9506 170778
rect 0 170688 800 170718
rect 482502 170716 482508 170780
rect 482572 170778 482578 170780
rect 486200 170778 487000 170808
rect 482572 170718 487000 170778
rect 482572 170716 482578 170718
rect 486200 170688 487000 170718
rect 9446 170212 10032 170272
rect 0 170098 800 170128
rect 9446 170098 9506 170212
rect 0 170038 9506 170098
rect 0 170008 800 170038
rect 485262 170036 485268 170100
rect 485332 170098 485338 170100
rect 486200 170098 487000 170128
rect 485332 170038 487000 170098
rect 485332 170036 485338 170038
rect 486200 170008 487000 170038
rect 0 169418 800 169448
rect 9446 169418 10032 169456
rect 0 169396 10032 169418
rect 0 169358 9506 169396
rect 0 169328 800 169358
rect 483790 169356 483796 169420
rect 483860 169418 483866 169420
rect 486200 169418 487000 169448
rect 483860 169358 487000 169418
rect 483860 169356 483866 169358
rect 486200 169328 487000 169358
rect 0 168738 800 168768
rect 0 168696 9506 168738
rect 0 168678 10032 168696
rect 0 168648 800 168678
rect 9446 168636 10032 168678
rect 485998 168676 486004 168740
rect 486068 168738 486074 168740
rect 486200 168738 487000 168768
rect 486068 168678 487000 168738
rect 486068 168676 486074 168678
rect 486200 168648 487000 168678
rect 0 168058 800 168088
rect 486200 168061 487000 168088
rect 0 167998 9506 168058
rect 0 167968 800 167998
rect 9446 167880 9506 167998
rect 486141 168056 487000 168061
rect 486141 168000 486146 168056
rect 486202 168000 487000 168056
rect 486141 167995 487000 168000
rect 486200 167968 487000 167995
rect 9446 167820 10032 167880
rect 485446 167316 485452 167380
rect 485516 167378 485522 167380
rect 486200 167378 487000 167408
rect 485516 167318 487000 167378
rect 485516 167316 485522 167318
rect 486200 167288 487000 167318
rect 6870 167064 9506 167106
rect 6870 167046 10032 167064
rect 0 166698 800 166728
rect 6870 166698 6930 167046
rect 9446 167004 10032 167046
rect 0 166638 6930 166698
rect 483657 166698 483723 166701
rect 486200 166698 487000 166728
rect 483657 166696 487000 166698
rect 483657 166640 483662 166696
rect 483718 166640 487000 166696
rect 483657 166638 487000 166640
rect 0 166608 800 166638
rect 483657 166635 483723 166638
rect 486200 166608 487000 166638
rect 9446 166132 10032 166192
rect 0 166018 800 166048
rect 9446 166018 9506 166132
rect 0 165958 9506 166018
rect 0 165928 800 165958
rect 479742 165956 479748 166020
rect 479812 166018 479818 166020
rect 486200 166018 487000 166048
rect 479812 165958 487000 166018
rect 479812 165956 479818 165958
rect 486200 165928 487000 165958
rect 0 165338 800 165368
rect 9446 165338 10032 165376
rect 0 165316 10032 165338
rect 0 165278 9506 165316
rect 0 165248 800 165278
rect 485814 165276 485820 165340
rect 485884 165338 485890 165340
rect 486200 165338 487000 165368
rect 485884 165278 487000 165338
rect 485884 165276 485890 165278
rect 486200 165248 487000 165278
rect 0 164658 800 164688
rect 486200 164660 487000 164688
rect 0 164616 9506 164658
rect 0 164598 10032 164616
rect 0 164568 800 164598
rect 9446 164556 10032 164598
rect 486200 164596 486372 164660
rect 486436 164596 487000 164660
rect 486200 164568 487000 164596
rect 0 163978 800 164008
rect 0 163918 9506 163978
rect 0 163888 800 163918
rect 9446 163800 9506 163918
rect 480846 163916 480852 163980
rect 480916 163978 480922 163980
rect 486200 163978 487000 164008
rect 480916 163918 487000 163978
rect 480916 163916 480922 163918
rect 486200 163888 487000 163918
rect 9446 163740 10032 163800
rect 480294 163236 480300 163300
rect 480364 163298 480370 163300
rect 486200 163298 487000 163328
rect 480364 163238 487000 163298
rect 480364 163236 480370 163238
rect 486200 163208 487000 163238
rect 9446 162890 10032 162928
rect 6870 162868 10032 162890
rect 6870 162830 9506 162868
rect 0 162618 800 162648
rect 6870 162618 6930 162830
rect 481633 162754 481699 162757
rect 486049 162754 486115 162757
rect 481633 162752 486115 162754
rect 481633 162696 481638 162752
rect 481694 162696 486054 162752
rect 486110 162696 486115 162752
rect 481633 162694 486115 162696
rect 481633 162691 481699 162694
rect 486049 162691 486115 162694
rect 0 162558 6930 162618
rect 0 162528 800 162558
rect 484158 162556 484164 162620
rect 484228 162618 484234 162620
rect 486200 162618 487000 162648
rect 484228 162558 487000 162618
rect 484228 162556 484234 162558
rect 486200 162528 487000 162558
rect 9446 162052 10032 162112
rect 0 161938 800 161968
rect 9446 161938 9506 162052
rect 0 161878 9506 161938
rect 0 161848 800 161878
rect 484710 161876 484716 161940
rect 484780 161938 484786 161940
rect 486200 161938 487000 161968
rect 484780 161878 487000 161938
rect 484780 161876 484786 161878
rect 486200 161848 487000 161878
rect 0 161258 800 161288
rect 9446 161258 10032 161296
rect 0 161236 10032 161258
rect 0 161198 9506 161236
rect 0 161168 800 161198
rect 485630 161196 485636 161260
rect 485700 161258 485706 161260
rect 486200 161258 487000 161288
rect 485700 161198 487000 161258
rect 485700 161196 485706 161198
rect 486200 161168 487000 161198
rect 0 160578 800 160608
rect 0 160536 9506 160578
rect 0 160518 10032 160536
rect 0 160488 800 160518
rect 9446 160476 10032 160518
rect 482870 160516 482876 160580
rect 482940 160578 482946 160580
rect 486200 160578 487000 160608
rect 482940 160518 487000 160578
rect 482940 160516 482946 160518
rect 486200 160488 487000 160518
rect 0 159898 800 159928
rect 0 159838 9506 159898
rect 0 159808 800 159838
rect 9446 159720 9506 159838
rect 483238 159836 483244 159900
rect 483308 159898 483314 159900
rect 486200 159898 487000 159928
rect 483308 159838 487000 159898
rect 483308 159836 483314 159838
rect 486200 159808 487000 159838
rect 9446 159660 10032 159720
rect 480478 159156 480484 159220
rect 480548 159218 480554 159220
rect 486200 159218 487000 159248
rect 480548 159158 487000 159218
rect 480548 159156 480554 159158
rect 486200 159128 487000 159158
rect 9446 158810 10032 158848
rect 6870 158788 10032 158810
rect 6870 158750 9506 158788
rect 0 158538 800 158568
rect 6870 158538 6930 158750
rect 0 158478 6930 158538
rect 0 158448 800 158478
rect 477166 158476 477172 158540
rect 477236 158538 477242 158540
rect 486200 158538 487000 158568
rect 477236 158478 487000 158538
rect 477236 158476 477242 158478
rect 486200 158448 487000 158478
rect 486182 158266 486188 158268
rect 477358 158240 486188 158266
rect 476940 158206 486188 158240
rect 476940 158180 477418 158206
rect 486182 158204 486188 158206
rect 486252 158204 486258 158268
rect 9446 157972 10032 158032
rect 483790 157994 483796 157996
rect 0 157858 800 157888
rect 9446 157858 9506 157972
rect 477358 157968 483796 157994
rect 476940 157934 483796 157968
rect 476940 157908 477418 157934
rect 483790 157932 483796 157934
rect 483860 157932 483866 157996
rect 486200 157858 487000 157888
rect 0 157798 9506 157858
rect 480210 157798 487000 157858
rect 0 157768 800 157798
rect 480210 157722 480270 157798
rect 486200 157768 487000 157798
rect 477174 157696 480270 157722
rect 476940 157662 480270 157696
rect 476940 157636 477234 157662
rect 483238 157586 483244 157588
rect 477358 157526 483244 157586
rect 477358 157424 477418 157526
rect 483238 157524 483244 157526
rect 483308 157524 483314 157588
rect 476940 157364 477418 157424
rect 483054 157388 483060 157452
rect 483124 157450 483130 157452
rect 483933 157450 483999 157453
rect 483124 157448 483999 157450
rect 483124 157392 483938 157448
rect 483994 157392 483999 157448
rect 483124 157390 483999 157392
rect 483124 157388 483130 157390
rect 483933 157387 483999 157390
rect 0 157178 800 157208
rect 9446 157178 10032 157216
rect 486200 157178 487000 157208
rect 0 157156 10032 157178
rect 0 157118 9506 157156
rect 477358 157152 487000 157178
rect 476940 157118 487000 157152
rect 0 157088 800 157118
rect 476940 157092 477418 157118
rect 486200 157088 487000 157118
rect 482870 156906 482876 156908
rect 477358 156880 482876 156906
rect 476940 156846 482876 156880
rect 476940 156820 477418 156846
rect 482870 156844 482876 156846
rect 482940 156844 482946 156908
rect 479885 156770 479951 156773
rect 480110 156770 480116 156772
rect 479885 156768 480116 156770
rect 479885 156712 479890 156768
rect 479946 156712 480116 156768
rect 479885 156710 480116 156712
rect 479885 156707 479951 156710
rect 480110 156708 480116 156710
rect 480180 156708 480186 156772
rect 485998 156634 486004 156636
rect 477358 156608 486004 156634
rect 476940 156574 486004 156608
rect 476940 156548 477418 156574
rect 485998 156572 486004 156574
rect 486068 156572 486074 156636
rect 0 156498 800 156528
rect 486200 156498 487000 156528
rect 0 156456 9506 156498
rect 0 156438 10032 156456
rect 0 156408 800 156438
rect 9446 156396 10032 156438
rect 480210 156438 487000 156498
rect 480210 156362 480270 156438
rect 486200 156408 487000 156438
rect 477358 156336 480270 156362
rect 476940 156302 480270 156336
rect 476940 156276 477418 156302
rect 484710 156090 484716 156092
rect 477358 156064 484716 156090
rect 476940 156030 484716 156064
rect 476940 156004 477418 156030
rect 484710 156028 484716 156030
rect 484780 156028 484786 156092
rect 481633 155956 481699 155957
rect 481582 155954 481588 155956
rect 481542 155894 481588 155954
rect 481652 155952 481699 155956
rect 481694 155896 481699 155952
rect 481582 155892 481588 155894
rect 481652 155892 481699 155896
rect 483238 155892 483244 155956
rect 483308 155954 483314 155956
rect 484025 155954 484091 155957
rect 485262 155954 485268 155956
rect 483308 155952 484091 155954
rect 483308 155896 484030 155952
rect 484086 155896 484091 155952
rect 483308 155894 484091 155896
rect 483308 155892 483314 155894
rect 481633 155891 481699 155892
rect 484025 155891 484091 155894
rect 484166 155894 485268 155954
rect 484166 155818 484226 155894
rect 485262 155892 485268 155894
rect 485332 155892 485338 155956
rect 477358 155792 484226 155818
rect 476940 155758 484226 155792
rect 476940 155732 477418 155758
rect 484342 155756 484348 155820
rect 484412 155818 484418 155820
rect 486200 155818 487000 155848
rect 484412 155758 487000 155818
rect 484412 155756 484418 155758
rect 486200 155728 487000 155758
rect 484158 155546 484164 155548
rect 477358 155520 484164 155546
rect 476940 155486 484164 155520
rect 476940 155460 477418 155486
rect 484158 155484 484164 155486
rect 484228 155484 484234 155548
rect 480294 155274 480300 155276
rect 477358 155248 480300 155274
rect 476940 155214 480300 155248
rect 476940 155188 477418 155214
rect 480294 155212 480300 155214
rect 480364 155212 480370 155276
rect 484526 155076 484532 155140
rect 484596 155138 484602 155140
rect 486200 155138 487000 155168
rect 484596 155078 487000 155138
rect 484596 155076 484602 155078
rect 486200 155048 487000 155078
rect 476940 154866 477418 154920
rect 486233 154866 486299 154869
rect 476940 154864 486299 154866
rect 476940 154860 486238 154864
rect 477358 154808 486238 154860
rect 486294 154808 486299 154864
rect 477358 154806 486299 154808
rect 486233 154803 486299 154806
rect 480989 154730 481055 154733
rect 477358 154728 481055 154730
rect 477358 154704 480994 154728
rect 476940 154672 480994 154704
rect 481050 154672 481055 154728
rect 476940 154670 481055 154672
rect 476940 154644 477418 154670
rect 480989 154667 481055 154670
rect 478638 154396 478644 154460
rect 478708 154458 478714 154460
rect 486200 154458 487000 154488
rect 478708 154398 487000 154458
rect 478708 154396 478714 154398
rect 476940 154322 477418 154376
rect 486200 154368 487000 154398
rect 484342 154322 484348 154324
rect 476940 154316 484348 154322
rect 477358 154262 484348 154316
rect 484342 154260 484348 154262
rect 484412 154260 484418 154324
rect 480897 154186 480963 154189
rect 477358 154184 480963 154186
rect 477358 154160 480902 154184
rect 476940 154128 480902 154160
rect 480958 154128 480963 154184
rect 476940 154126 480963 154128
rect 476940 154100 477418 154126
rect 480897 154123 480963 154126
rect 485814 153914 485820 153916
rect 477358 153888 485820 153914
rect 476940 153854 485820 153888
rect 476940 153828 477418 153854
rect 485814 153852 485820 153854
rect 485884 153852 485890 153916
rect 479926 153716 479932 153780
rect 479996 153778 480002 153780
rect 486200 153778 487000 153808
rect 479996 153718 487000 153778
rect 479996 153716 480002 153718
rect 486200 153688 487000 153718
rect 476940 153506 477418 153560
rect 484526 153506 484532 153508
rect 476940 153500 484532 153506
rect 477358 153446 484532 153500
rect 484526 153444 484532 153446
rect 484596 153444 484602 153508
rect 479742 153370 479748 153372
rect 477358 153344 479748 153370
rect 476940 153310 479748 153344
rect 476940 153284 477418 153310
rect 479742 153308 479748 153310
rect 479812 153308 479818 153372
rect 480478 153098 480484 153100
rect 477358 153072 480484 153098
rect 476940 153038 480484 153072
rect 476940 153012 477418 153038
rect 480478 153036 480484 153038
rect 480548 153036 480554 153100
rect 480662 153036 480668 153100
rect 480732 153098 480738 153100
rect 481541 153098 481607 153101
rect 480732 153096 481607 153098
rect 480732 153040 481546 153096
rect 481602 153040 481607 153096
rect 480732 153038 481607 153040
rect 480732 153036 480738 153038
rect 481541 153035 481607 153038
rect 485998 153036 486004 153100
rect 486068 153098 486074 153100
rect 486200 153098 487000 153128
rect 486068 153038 487000 153098
rect 486068 153036 486074 153038
rect 486200 153008 487000 153038
rect 477718 152900 477724 152964
rect 477788 152962 477794 152964
rect 478505 152962 478571 152965
rect 477788 152960 478571 152962
rect 477788 152904 478510 152960
rect 478566 152904 478571 152960
rect 477788 152902 478571 152904
rect 477788 152900 477794 152902
rect 478505 152899 478571 152902
rect 483657 152826 483723 152829
rect 477358 152824 483723 152826
rect 477358 152800 483662 152824
rect 476940 152768 483662 152800
rect 483718 152768 483723 152824
rect 476940 152766 483723 152768
rect 476940 152740 477418 152766
rect 483657 152763 483723 152766
rect 477534 152628 477540 152692
rect 477604 152690 477610 152692
rect 478597 152690 478663 152693
rect 477604 152688 478663 152690
rect 477604 152632 478602 152688
rect 478658 152632 478663 152688
rect 477604 152630 478663 152632
rect 477604 152628 477610 152630
rect 478597 152627 478663 152630
rect 485446 152554 485452 152556
rect 477358 152528 485452 152554
rect 476940 152494 485452 152528
rect 476940 152468 477418 152494
rect 485446 152492 485452 152494
rect 485516 152492 485522 152556
rect 484710 152356 484716 152420
rect 484780 152418 484786 152420
rect 486200 152418 487000 152448
rect 484780 152358 487000 152418
rect 484780 152356 484786 152358
rect 486200 152328 487000 152358
rect 478638 152282 478644 152284
rect 477358 152256 478644 152282
rect 476940 152222 478644 152256
rect 476940 152196 477418 152222
rect 478638 152220 478644 152222
rect 478708 152220 478714 152284
rect 477902 152010 477908 152012
rect 477358 151984 477908 152010
rect 476940 151950 477908 151984
rect 476940 151924 477418 151950
rect 477902 151948 477908 151950
rect 477972 151948 477978 152012
rect 480846 151738 480852 151740
rect 477358 151712 480852 151738
rect 476940 151678 480852 151712
rect 476940 151652 477418 151678
rect 480846 151676 480852 151678
rect 480916 151676 480922 151740
rect 483105 151738 483171 151741
rect 486200 151738 487000 151768
rect 483105 151736 487000 151738
rect 483105 151680 483110 151736
rect 483166 151680 487000 151736
rect 483105 151678 487000 151680
rect 483105 151675 483171 151678
rect 486200 151648 487000 151678
rect 482134 151466 482140 151468
rect 477358 151440 482140 151466
rect 476940 151406 482140 151440
rect 476940 151380 477418 151406
rect 482134 151404 482140 151406
rect 482204 151404 482210 151468
rect 484710 151194 484716 151196
rect 477358 151168 484716 151194
rect 476940 151134 484716 151168
rect 476940 151108 477418 151134
rect 484710 151132 484716 151134
rect 484780 151132 484786 151196
rect 486200 151058 487000 151088
rect 483246 150998 487000 151058
rect 483105 150922 483171 150925
rect 477358 150920 483171 150922
rect 477358 150896 483110 150920
rect 476940 150864 483110 150896
rect 483166 150864 483171 150920
rect 476940 150862 483171 150864
rect 476940 150836 477418 150862
rect 483105 150859 483171 150862
rect 483246 150650 483306 150998
rect 486200 150968 487000 150998
rect 477358 150624 483306 150650
rect 476940 150590 483306 150624
rect 476940 150564 477418 150590
rect 481950 150452 481956 150516
rect 482020 150514 482026 150516
rect 482645 150514 482711 150517
rect 482020 150512 482711 150514
rect 482020 150456 482650 150512
rect 482706 150456 482711 150512
rect 482020 150454 482711 150456
rect 482020 150452 482026 150454
rect 482645 150451 482711 150454
rect 483790 150452 483796 150516
rect 483860 150514 483866 150516
rect 484117 150514 484183 150517
rect 483860 150512 484183 150514
rect 483860 150456 484122 150512
rect 484178 150456 484183 150512
rect 483860 150454 484183 150456
rect 483860 150452 483866 150454
rect 484117 150451 484183 150454
rect 482502 150378 482508 150380
rect 477358 150352 482508 150378
rect 476940 150318 482508 150352
rect 476940 150292 477418 150318
rect 482502 150316 482508 150318
rect 482572 150316 482578 150380
rect 484710 150316 484716 150380
rect 484780 150378 484786 150380
rect 486200 150378 487000 150408
rect 484780 150318 487000 150378
rect 484780 150316 484786 150318
rect 486200 150288 487000 150318
rect 480662 150106 480668 150108
rect 477358 150080 480668 150106
rect 476940 150046 480668 150080
rect 476940 150020 477418 150046
rect 480662 150044 480668 150046
rect 480732 150044 480738 150108
rect 477166 149808 477172 149810
rect 476940 149748 477172 149808
rect 477166 149746 477172 149748
rect 477236 149746 477242 149810
rect 484342 149636 484348 149700
rect 484412 149698 484418 149700
rect 486200 149698 487000 149728
rect 484412 149638 487000 149698
rect 484412 149636 484418 149638
rect 486200 149608 487000 149638
rect 479926 149562 479932 149564
rect 477174 149536 479932 149562
rect 476940 149502 479932 149536
rect 476940 149476 477234 149502
rect 479926 149500 479932 149502
rect 479996 149500 480002 149564
rect 482318 149426 482324 149428
rect 477358 149366 482324 149426
rect 477358 149264 477418 149366
rect 482318 149364 482324 149366
rect 482388 149364 482394 149428
rect 476940 149204 477418 149264
rect 481766 149228 481772 149292
rect 481836 149290 481842 149292
rect 482829 149290 482895 149293
rect 481836 149288 482895 149290
rect 481836 149232 482834 149288
rect 482890 149232 482895 149288
rect 481836 149230 482895 149232
rect 481836 149228 481842 149230
rect 482829 149227 482895 149230
rect 482134 149092 482140 149156
rect 482204 149154 482210 149156
rect 482737 149154 482803 149157
rect 482204 149152 482803 149154
rect 482204 149096 482742 149152
rect 482798 149096 482803 149152
rect 482204 149094 482803 149096
rect 482204 149092 482210 149094
rect 482737 149091 482803 149094
rect 485446 149018 485452 149020
rect 477358 148992 485452 149018
rect 476940 148958 485452 148992
rect 476940 148932 477418 148958
rect 485446 148956 485452 148958
rect 485516 148956 485522 149020
rect 485630 148956 485636 149020
rect 485700 149018 485706 149020
rect 486200 149018 487000 149048
rect 485700 148958 487000 149018
rect 485700 148956 485706 148958
rect 486200 148928 487000 148958
rect 479190 148820 479196 148884
rect 479260 148882 479266 148884
rect 480069 148882 480135 148885
rect 479260 148880 480135 148882
rect 479260 148824 480074 148880
rect 480130 148824 480135 148880
rect 479260 148822 480135 148824
rect 479260 148820 479266 148822
rect 480069 148819 480135 148822
rect 479977 148748 480043 148749
rect 479558 148746 479564 148748
rect 477358 148720 479564 148746
rect 476940 148686 479564 148720
rect 476940 148660 477418 148686
rect 479558 148684 479564 148686
rect 479628 148684 479634 148748
rect 479926 148684 479932 148748
rect 479996 148746 480043 148748
rect 479996 148744 480088 148746
rect 480038 148688 480088 148744
rect 479996 148686 480088 148688
rect 479996 148684 480043 148686
rect 479977 148683 480043 148684
rect 483606 148474 483612 148476
rect 477358 148448 483612 148474
rect 476940 148414 483612 148448
rect 476940 148388 477418 148414
rect 483606 148412 483612 148414
rect 483676 148412 483682 148476
rect 0 148338 800 148368
rect 0 148278 9506 148338
rect 0 148248 800 148278
rect 9446 148176 9506 148278
rect 484526 148276 484532 148340
rect 484596 148338 484602 148340
rect 486200 148338 487000 148368
rect 484596 148278 487000 148338
rect 484596 148276 484602 148278
rect 486200 148248 487000 148278
rect 484342 148202 484348 148204
rect 477358 148176 484348 148202
rect 9446 148116 10060 148176
rect 476940 148142 484348 148176
rect 476940 148116 477418 148142
rect 484342 148140 484348 148142
rect 484412 148140 484418 148204
rect 478086 147930 478092 147932
rect 477358 147904 478092 147930
rect 476940 147870 478092 147904
rect 476940 147844 477418 147870
rect 478086 147868 478092 147870
rect 478156 147868 478162 147932
rect 477902 147732 477908 147796
rect 477972 147794 477978 147796
rect 478689 147794 478755 147797
rect 477972 147792 478755 147794
rect 477972 147736 478694 147792
rect 478750 147736 478755 147792
rect 477972 147734 478755 147736
rect 477972 147732 477978 147734
rect 478689 147731 478755 147734
rect 483422 147732 483428 147796
rect 483492 147794 483498 147796
rect 484209 147794 484275 147797
rect 483492 147792 484275 147794
rect 483492 147736 484214 147792
rect 484270 147736 484275 147792
rect 483492 147734 484275 147736
rect 483492 147732 483498 147734
rect 484209 147731 484275 147734
rect 0 147658 800 147688
rect 486200 147658 487000 147688
rect 0 147598 9506 147658
rect 477358 147632 487000 147658
rect 0 147568 800 147598
rect 9446 147360 9506 147598
rect 476940 147598 487000 147632
rect 476940 147572 477418 147598
rect 486200 147568 487000 147598
rect 479374 147386 479380 147388
rect 477358 147360 479380 147386
rect 9446 147300 10060 147360
rect 476940 147326 479380 147360
rect 476940 147300 477418 147326
rect 479374 147324 479380 147326
rect 479444 147324 479450 147388
rect 479517 147114 479583 147117
rect 477358 147112 479583 147114
rect 477358 147088 479522 147112
rect 476940 147056 479522 147088
rect 479578 147056 479583 147112
rect 476940 147054 479583 147056
rect 476940 147028 477418 147054
rect 479517 147051 479583 147054
rect 480662 147052 480668 147116
rect 480732 147114 480738 147116
rect 481449 147114 481515 147117
rect 480732 147112 481515 147114
rect 480732 147056 481454 147112
rect 481510 147056 481515 147112
rect 480732 147054 481515 147056
rect 480732 147052 480738 147054
rect 481449 147051 481515 147054
rect 479742 146916 479748 146980
rect 479812 146978 479818 146980
rect 486200 146978 487000 147008
rect 479812 146918 487000 146978
rect 479812 146916 479818 146918
rect 486200 146888 487000 146918
rect 476940 146706 477418 146760
rect 484526 146706 484532 146708
rect 476940 146700 484532 146706
rect 477358 146646 484532 146700
rect 484526 146644 484532 146646
rect 484596 146644 484602 146708
rect 480110 146570 480116 146572
rect 477358 146544 480116 146570
rect 476940 146510 480116 146544
rect 9446 146434 10060 146488
rect 476940 146484 477418 146510
rect 480110 146508 480116 146510
rect 480180 146508 480186 146572
rect 480161 146434 480227 146437
rect 6870 146428 10060 146434
rect 480118 146432 480227 146434
rect 6870 146374 9506 146428
rect 480118 146376 480166 146432
rect 480222 146376 480227 146432
rect 0 146298 800 146328
rect 6870 146298 6930 146374
rect 480118 146371 480227 146376
rect 480118 146298 480178 146371
rect 0 146238 6930 146298
rect 477358 146272 480178 146298
rect 476940 146238 480178 146272
rect 0 146208 800 146238
rect 476940 146212 477418 146238
rect 482318 146236 482324 146300
rect 482388 146298 482394 146300
rect 482921 146298 482987 146301
rect 482388 146296 482987 146298
rect 482388 146240 482926 146296
rect 482982 146240 482987 146296
rect 482388 146238 482987 146240
rect 482388 146236 482394 146238
rect 482921 146235 482987 146238
rect 483606 146236 483612 146300
rect 483676 146298 483682 146300
rect 484301 146298 484367 146301
rect 483676 146296 484367 146298
rect 483676 146240 484306 146296
rect 484362 146240 484367 146296
rect 483676 146238 484367 146240
rect 483676 146236 483682 146238
rect 484301 146235 484367 146238
rect 484526 146236 484532 146300
rect 484596 146298 484602 146300
rect 486200 146298 487000 146328
rect 484596 146238 487000 146298
rect 484596 146236 484602 146238
rect 486200 146208 487000 146238
rect 479190 146026 479196 146028
rect 477358 146000 479196 146026
rect 476940 145966 479196 146000
rect 476940 145940 477418 145966
rect 479190 145964 479196 145966
rect 479260 145964 479266 146028
rect 479926 145754 479932 145756
rect 477358 145728 479932 145754
rect 476940 145694 479932 145728
rect 0 145618 800 145648
rect 9446 145618 10060 145672
rect 476940 145668 477418 145694
rect 479926 145692 479932 145694
rect 479996 145692 480002 145756
rect 0 145612 10060 145618
rect 0 145558 9506 145612
rect 0 145528 800 145558
rect 484342 145556 484348 145620
rect 484412 145618 484418 145620
rect 486200 145618 487000 145648
rect 484412 145558 487000 145618
rect 484412 145556 484418 145558
rect 486200 145528 487000 145558
rect 483238 145482 483244 145484
rect 477358 145456 483244 145482
rect 476940 145422 483244 145456
rect 476940 145396 477418 145422
rect 483238 145420 483244 145422
rect 483308 145420 483314 145484
rect 481582 145210 481588 145212
rect 477358 145184 481588 145210
rect 476940 145150 481588 145184
rect 476940 145124 477418 145150
rect 481582 145148 481588 145150
rect 481652 145148 481658 145212
rect 0 144938 800 144968
rect 486200 144938 487000 144968
rect 0 144906 9874 144938
rect 477174 144912 487000 144938
rect 0 144878 10060 144906
rect 0 144848 800 144878
rect 9814 144846 10060 144878
rect 476940 144878 487000 144912
rect 476940 144852 477234 144878
rect 486200 144848 487000 144878
rect 478638 144740 478644 144804
rect 478708 144802 478714 144804
rect 478781 144802 478847 144805
rect 478708 144800 478847 144802
rect 478708 144744 478786 144800
rect 478842 144744 478847 144800
rect 478708 144742 478847 144744
rect 478708 144740 478714 144742
rect 478781 144739 478847 144742
rect 478137 144666 478203 144669
rect 477358 144664 478203 144666
rect 477358 144640 478142 144664
rect 476940 144608 478142 144640
rect 478198 144608 478203 144664
rect 476940 144606 478203 144608
rect 476940 144580 477418 144606
rect 478137 144603 478203 144606
rect 481950 144394 481956 144396
rect 477358 144368 481956 144394
rect 476940 144334 481956 144368
rect 476940 144308 477418 144334
rect 481950 144332 481956 144334
rect 482020 144332 482026 144396
rect 0 144258 800 144288
rect 0 144198 9506 144258
rect 0 144168 800 144198
rect 9446 144096 9506 144198
rect 478822 144196 478828 144260
rect 478892 144258 478898 144260
rect 486200 144258 487000 144288
rect 478892 144198 487000 144258
rect 478892 144196 478898 144198
rect 486200 144168 487000 144198
rect 484526 144122 484532 144124
rect 477358 144096 484532 144122
rect 9446 144036 10060 144096
rect 476940 144062 484532 144096
rect 476940 144036 477418 144062
rect 484526 144060 484532 144062
rect 484596 144060 484602 144124
rect 478270 143850 478276 143852
rect 477174 143824 478276 143850
rect 476940 143790 478276 143824
rect 476940 143764 477234 143790
rect 478270 143788 478276 143790
rect 478340 143788 478346 143852
rect 484342 143714 484348 143716
rect 477358 143654 484348 143714
rect 0 143578 800 143608
rect 0 143518 4170 143578
rect 477358 143552 477418 143654
rect 484342 143652 484348 143654
rect 484412 143652 484418 143716
rect 0 143488 800 143518
rect 4110 143442 4170 143518
rect 476940 143492 477418 143552
rect 480110 143516 480116 143580
rect 480180 143578 480186 143580
rect 486200 143578 487000 143608
rect 480180 143518 487000 143578
rect 480180 143516 480186 143518
rect 486200 143488 487000 143518
rect 4110 143382 9506 143442
rect 9446 143280 9506 143382
rect 477718 143306 477724 143308
rect 477358 143280 477724 143306
rect 9446 143220 10060 143280
rect 476940 143246 477724 143280
rect 476940 143220 477418 143246
rect 477718 143244 477724 143246
rect 477788 143244 477794 143308
rect 477534 143034 477540 143036
rect 477358 143008 477540 143034
rect 476940 142974 477540 143008
rect 476940 142948 477418 142974
rect 477534 142972 477540 142974
rect 477604 142972 477610 143036
rect 480478 142836 480484 142900
rect 480548 142898 480554 142900
rect 486200 142898 487000 142928
rect 480548 142838 487000 142898
rect 480548 142836 480554 142838
rect 486200 142808 487000 142838
rect 478822 142762 478828 142764
rect 477358 142736 478828 142762
rect 476940 142702 478828 142736
rect 476940 142676 477418 142702
rect 478822 142700 478828 142702
rect 478892 142700 478898 142764
rect 484710 142490 484716 142492
rect 477358 142464 484716 142490
rect 476940 142430 484716 142464
rect 9446 142348 10060 142408
rect 476940 142404 477418 142430
rect 484710 142428 484716 142430
rect 484780 142428 484786 142492
rect 485998 142354 486004 142356
rect 0 142218 800 142248
rect 9446 142218 9506 142348
rect 478830 142294 486004 142354
rect 478830 142218 478890 142294
rect 485998 142292 486004 142294
rect 486068 142292 486074 142356
rect 0 142158 9506 142218
rect 477358 142192 478890 142218
rect 476940 142158 478890 142192
rect 0 142128 800 142158
rect 476940 142132 477418 142158
rect 480294 142156 480300 142220
rect 480364 142218 480370 142220
rect 486200 142218 487000 142248
rect 480364 142158 487000 142218
rect 480364 142156 480370 142158
rect 486200 142128 487000 142158
rect 480478 141946 480484 141948
rect 477358 141920 480484 141946
rect 476940 141886 480484 141920
rect 476940 141860 477418 141886
rect 480478 141884 480484 141886
rect 480548 141884 480554 141948
rect 480110 141674 480116 141676
rect 477174 141648 480116 141674
rect 476940 141614 480116 141648
rect 0 141538 800 141568
rect 9446 141538 10060 141592
rect 476940 141588 477234 141614
rect 480110 141612 480116 141614
rect 480180 141612 480186 141676
rect 486200 141538 487000 141568
rect 0 141532 10060 141538
rect 0 141478 9506 141532
rect 477358 141478 487000 141538
rect 0 141448 800 141478
rect 477358 141376 477418 141478
rect 486200 141448 487000 141478
rect 476940 141316 477418 141376
rect 480294 141130 480300 141132
rect 477358 141104 480300 141130
rect 476940 141070 480300 141104
rect 476940 141044 477418 141070
rect 480294 141068 480300 141070
rect 480364 141068 480370 141132
rect 0 140858 800 140888
rect 486200 140858 487000 140888
rect 0 140832 9506 140858
rect 477358 140832 487000 140858
rect 0 140798 10060 140832
rect 0 140768 800 140798
rect 9446 140772 10060 140798
rect 476940 140798 487000 140832
rect 476940 140772 477418 140798
rect 486200 140768 487000 140798
rect 478638 140586 478644 140588
rect 477358 140560 478644 140586
rect 476940 140526 478644 140560
rect 476940 140500 477418 140526
rect 478638 140524 478644 140526
rect 478708 140524 478714 140588
rect 477902 140314 477908 140316
rect 477174 140288 477908 140314
rect 476940 140254 477908 140288
rect 476940 140228 477234 140254
rect 477902 140252 477908 140254
rect 477972 140252 477978 140316
rect 0 140178 800 140208
rect 486200 140178 487000 140208
rect 0 140118 9506 140178
rect 0 140088 800 140118
rect 9446 140016 9506 140118
rect 477358 140118 487000 140178
rect 477358 140016 477418 140118
rect 486200 140088 487000 140118
rect 9446 139956 10060 140016
rect 476940 139956 477418 140016
rect 483790 139770 483796 139772
rect 477358 139744 483796 139770
rect 476940 139710 483796 139744
rect 476940 139684 477418 139710
rect 483790 139708 483796 139710
rect 483860 139708 483866 139772
rect 0 139498 800 139528
rect 486200 139498 487000 139528
rect 0 139438 4170 139498
rect 477358 139472 487000 139498
rect 0 139408 800 139438
rect 4110 139362 4170 139438
rect 476940 139438 487000 139472
rect 476940 139412 477418 139438
rect 486200 139408 487000 139438
rect 4110 139302 9506 139362
rect 9446 139200 9506 139302
rect 482134 139226 482140 139228
rect 477358 139200 482140 139226
rect 9446 139140 10060 139200
rect 476940 139166 482140 139200
rect 476940 139140 477418 139166
rect 482134 139164 482140 139166
rect 482204 139164 482210 139228
rect 483422 138954 483428 138956
rect 477358 138928 483428 138954
rect 476940 138894 483428 138928
rect 476940 138868 477418 138894
rect 483422 138892 483428 138894
rect 483492 138892 483498 138956
rect 484526 138756 484532 138820
rect 484596 138818 484602 138820
rect 486200 138818 487000 138848
rect 484596 138758 487000 138818
rect 484596 138756 484602 138758
rect 486200 138728 487000 138758
rect 485630 138682 485636 138684
rect 477358 138656 485636 138682
rect 476940 138622 485636 138656
rect 476940 138596 477418 138622
rect 485630 138620 485636 138622
rect 485700 138620 485706 138684
rect 481766 138410 481772 138412
rect 477358 138384 481772 138410
rect 476940 138350 481772 138384
rect 9446 138268 10060 138328
rect 476940 138324 477418 138350
rect 481766 138348 481772 138350
rect 481836 138348 481842 138412
rect 0 138138 800 138168
rect 9446 138138 9506 138268
rect 486200 138138 487000 138168
rect 0 138078 9506 138138
rect 477358 138112 487000 138138
rect 476940 138078 487000 138112
rect 0 138048 800 138078
rect 476940 138052 477418 138078
rect 486200 138048 487000 138078
rect 483606 137866 483612 137868
rect 477358 137840 483612 137866
rect 476940 137806 483612 137840
rect 476940 137780 477418 137806
rect 483606 137804 483612 137806
rect 483676 137804 483682 137868
rect 482318 137594 482324 137596
rect 477358 137568 482324 137594
rect 476940 137534 482324 137568
rect 0 137458 800 137488
rect 9446 137458 10060 137512
rect 476940 137508 477418 137534
rect 482318 137532 482324 137534
rect 482388 137532 482394 137596
rect 0 137452 10060 137458
rect 0 137398 9506 137452
rect 0 137368 800 137398
rect 484342 137396 484348 137460
rect 484412 137458 484418 137460
rect 486200 137458 487000 137488
rect 484412 137398 487000 137458
rect 484412 137396 484418 137398
rect 486200 137368 487000 137398
rect 480662 137322 480668 137324
rect 477358 137296 480668 137322
rect 476940 137262 480668 137296
rect 476940 137236 477418 137262
rect 480662 137260 480668 137262
rect 480732 137260 480738 137324
rect 484526 137050 484532 137052
rect 477358 137024 484532 137050
rect 476940 136990 484532 137024
rect 476940 136964 477418 136990
rect 484526 136988 484532 136990
rect 484596 136988 484602 137052
rect 0 136778 800 136808
rect 486200 136778 487000 136808
rect 0 136752 9506 136778
rect 477358 136752 487000 136778
rect 0 136718 10060 136752
rect 0 136688 800 136718
rect 9446 136692 10060 136718
rect 476940 136718 487000 136752
rect 476940 136692 477418 136718
rect 486200 136688 487000 136718
rect 484342 136506 484348 136508
rect 477358 136480 484348 136506
rect 476940 136446 484348 136480
rect 476940 136420 477418 136446
rect 484342 136444 484348 136446
rect 484412 136444 484418 136508
rect 483054 136234 483060 136236
rect 477358 136208 483060 136234
rect 476940 136174 483060 136208
rect 476940 136148 477418 136174
rect 483054 136172 483060 136174
rect 483124 136172 483130 136236
rect 0 136098 800 136128
rect 486200 136098 487000 136128
rect 0 136038 9506 136098
rect 0 136008 800 136038
rect 9446 135936 9506 136038
rect 480210 136038 487000 136098
rect 479742 135962 479748 135964
rect 477174 135936 479748 135962
rect 9446 135876 10060 135936
rect 476940 135902 479748 135936
rect 476940 135876 477234 135902
rect 479742 135900 479748 135902
rect 479812 135900 479818 135964
rect 480210 135826 480270 136038
rect 486200 136008 487000 136038
rect 477358 135766 480270 135826
rect 477358 135664 477418 135766
rect 476940 135604 477418 135664
rect 0 135418 800 135448
rect 486200 135418 487000 135448
rect 0 135358 4170 135418
rect 477358 135392 487000 135418
rect 0 135328 800 135358
rect 4110 135146 4170 135358
rect 476940 135358 487000 135392
rect 476940 135332 477418 135358
rect 486200 135328 487000 135358
rect 483657 135146 483723 135149
rect 4110 135120 9506 135146
rect 477358 135144 483723 135146
rect 477358 135120 483662 135144
rect 4110 135086 10060 135120
rect 9446 135060 10060 135086
rect 476940 135088 483662 135120
rect 483718 135088 483723 135144
rect 476940 135086 483723 135088
rect 476940 135060 477418 135086
rect 483657 135083 483723 135086
rect 476940 134738 477418 134792
rect 486200 134738 487000 134768
rect 476940 134732 487000 134738
rect 477358 134678 487000 134732
rect 486200 134648 487000 134678
rect 476940 134466 477418 134520
rect 485814 134466 485820 134468
rect 476940 134460 485820 134466
rect 477358 134406 485820 134460
rect 485814 134404 485820 134406
rect 485884 134404 485890 134468
rect 477358 134304 483306 134330
rect 476940 134270 483306 134304
rect 9446 134188 10060 134248
rect 476940 134244 477418 134270
rect 0 134058 800 134088
rect 9446 134058 9506 134188
rect 0 133998 9506 134058
rect 483246 134058 483306 134270
rect 486200 134058 487000 134088
rect 483246 133998 487000 134058
rect 0 133968 800 133998
rect 476940 133922 477418 133976
rect 486200 133968 487000 133998
rect 485998 133922 486004 133924
rect 476940 133916 486004 133922
rect 477358 133862 486004 133916
rect 485998 133860 486004 133862
rect 486068 133860 486074 133924
rect 476940 133650 477418 133704
rect 478270 133650 478276 133652
rect 476940 133644 478276 133650
rect 477358 133590 478276 133644
rect 478270 133588 478276 133590
rect 478340 133588 478346 133652
rect 0 133378 800 133408
rect 9446 133378 10060 133432
rect 0 133372 10060 133378
rect 476940 133378 477418 133432
rect 486200 133378 487000 133408
rect 476940 133372 487000 133378
rect 0 133318 9506 133372
rect 477358 133318 487000 133372
rect 0 133288 800 133318
rect 486200 133288 487000 133318
rect 476940 133106 477418 133160
rect 478086 133106 478092 133108
rect 476940 133100 478092 133106
rect 477358 133046 478092 133100
rect 478086 133044 478092 133046
rect 478156 133044 478162 133108
rect 476940 132834 477418 132888
rect 476940 132828 480270 132834
rect 477358 132774 480270 132828
rect 0 132698 800 132728
rect 480210 132698 480270 132774
rect 486200 132698 487000 132728
rect 0 132672 9506 132698
rect 0 132638 10060 132672
rect 480210 132638 487000 132698
rect 0 132608 800 132638
rect 9446 132612 10060 132638
rect 476940 132562 477418 132616
rect 486200 132608 487000 132638
rect 485998 132562 486004 132564
rect 476940 132556 486004 132562
rect 477358 132502 486004 132556
rect 485998 132500 486004 132502
rect 486068 132500 486074 132564
rect 477350 132344 477356 132346
rect 476940 132284 477356 132344
rect 477350 132282 477356 132284
rect 477420 132282 477426 132346
rect 0 132018 800 132048
rect 476940 132018 477418 132072
rect 486200 132018 487000 132048
rect 0 131958 9506 132018
rect 476940 132012 487000 132018
rect 477358 131958 487000 132012
rect 0 131928 800 131958
rect 9446 131856 9506 131958
rect 486200 131928 487000 131958
rect 9446 131796 10060 131856
rect 476940 131746 477418 131800
rect 481398 131746 481404 131748
rect 476940 131740 481404 131746
rect 477358 131686 481404 131740
rect 481398 131684 481404 131686
rect 481468 131684 481474 131748
rect 476940 131474 477418 131528
rect 476940 131468 480270 131474
rect 477358 131414 480270 131468
rect 0 131338 800 131368
rect 480210 131338 480270 131414
rect 486200 131338 487000 131368
rect 0 131278 4170 131338
rect 480210 131278 487000 131338
rect 0 131248 800 131278
rect 4110 131066 4170 131278
rect 476940 131202 477418 131256
rect 486200 131248 487000 131278
rect 481582 131202 481588 131204
rect 476940 131196 481588 131202
rect 477358 131142 481588 131196
rect 481582 131140 481588 131142
rect 481652 131140 481658 131204
rect 484526 131066 484532 131068
rect 4110 131040 9506 131066
rect 477358 131040 484532 131066
rect 4110 131006 10060 131040
rect 9446 130980 10060 131006
rect 476940 131006 484532 131040
rect 476940 130980 477418 131006
rect 484526 131004 484532 131006
rect 484596 131004 484602 131068
rect 476940 130658 477418 130712
rect 486200 130658 487000 130688
rect 476940 130652 487000 130658
rect 477358 130598 487000 130652
rect 486200 130568 487000 130598
rect 476940 130386 477418 130440
rect 484342 130386 484348 130388
rect 476940 130380 484348 130386
rect 477358 130326 484348 130380
rect 484342 130324 484348 130326
rect 484412 130324 484418 130388
rect 477358 130224 483306 130250
rect 476940 130190 483306 130224
rect 9446 130108 10060 130168
rect 476940 130164 477418 130190
rect 0 129978 800 130008
rect 9446 129978 9506 130108
rect 483054 129978 483060 129980
rect 0 129918 9506 129978
rect 477358 129952 483060 129978
rect 476940 129918 483060 129952
rect 0 129888 800 129918
rect 476940 129892 477418 129918
rect 483054 129916 483060 129918
rect 483124 129916 483130 129980
rect 483246 129978 483306 130190
rect 486200 129978 487000 130008
rect 483246 129918 487000 129978
rect 486200 129888 487000 129918
rect 476940 129570 477418 129624
rect 478822 129570 478828 129572
rect 476940 129564 478828 129570
rect 477358 129510 478828 129564
rect 478822 129508 478828 129510
rect 478892 129508 478898 129572
rect 0 129298 800 129328
rect 9446 129298 10060 129352
rect 0 129292 10060 129298
rect 476940 129298 477418 129352
rect 486200 129298 487000 129328
rect 476940 129292 487000 129298
rect 0 129238 9506 129292
rect 477358 129238 487000 129292
rect 0 129208 800 129238
rect 486200 129208 487000 129238
rect 477358 129136 483306 129162
rect 476940 129102 483306 129136
rect 476940 129076 477418 129102
rect 476940 128748 477418 128808
rect 0 128618 800 128648
rect 0 128592 9506 128618
rect 0 128558 10060 128592
rect 0 128528 800 128558
rect 9446 128532 10060 128558
rect 477358 128482 477418 128748
rect 483246 128618 483306 129102
rect 486200 128618 487000 128648
rect 483246 128558 487000 128618
rect 486200 128528 487000 128558
rect 483790 128482 483796 128484
rect 477358 128422 483796 128482
rect 483790 128420 483796 128422
rect 483860 128420 483866 128484
rect 0 127938 800 127968
rect 0 127878 9506 127938
rect 0 127848 800 127878
rect 9446 127776 9506 127878
rect 478822 127876 478828 127940
rect 478892 127938 478898 127940
rect 486200 127938 487000 127968
rect 478892 127878 487000 127938
rect 478892 127876 478898 127878
rect 486200 127848 487000 127878
rect 9446 127716 10060 127776
rect 0 127258 800 127288
rect 0 127198 4170 127258
rect 0 127168 800 127198
rect 4110 126986 4170 127198
rect 483054 127196 483060 127260
rect 483124 127258 483130 127260
rect 486200 127258 487000 127288
rect 483124 127198 487000 127258
rect 483124 127196 483130 127198
rect 486200 127168 487000 127198
rect 4110 126960 9506 126986
rect 4110 126926 10060 126960
rect 9446 126900 10060 126926
rect 484342 126516 484348 126580
rect 484412 126578 484418 126580
rect 486200 126578 487000 126608
rect 484412 126518 487000 126578
rect 484412 126516 484418 126518
rect 486200 126488 487000 126518
rect 9446 126028 10060 126088
rect 0 125898 800 125928
rect 9446 125898 9506 126028
rect 0 125838 9506 125898
rect 0 125808 800 125838
rect 484526 125836 484532 125900
rect 484596 125898 484602 125900
rect 486200 125898 487000 125928
rect 484596 125838 487000 125898
rect 484596 125836 484602 125838
rect 486200 125808 487000 125838
rect 0 125218 800 125248
rect 9446 125218 10060 125272
rect 0 125212 10060 125218
rect 0 125158 9506 125212
rect 0 125128 800 125158
rect 481582 125156 481588 125220
rect 481652 125218 481658 125220
rect 486200 125218 487000 125248
rect 481652 125158 487000 125218
rect 481652 125156 481658 125158
rect 486200 125128 487000 125158
rect 0 124538 800 124568
rect 0 124512 9506 124538
rect 0 124478 10060 124512
rect 0 124448 800 124478
rect 9446 124452 10060 124478
rect 481398 124476 481404 124540
rect 481468 124538 481474 124540
rect 486200 124538 487000 124568
rect 481468 124478 487000 124538
rect 481468 124476 481474 124478
rect 486200 124448 487000 124478
rect 0 123858 800 123888
rect 0 123798 9506 123858
rect 0 123768 800 123798
rect 9446 123696 9506 123798
rect 477350 123796 477356 123860
rect 477420 123858 477426 123860
rect 486200 123858 487000 123888
rect 477420 123798 487000 123858
rect 477420 123796 477426 123798
rect 486200 123768 487000 123798
rect 9446 123636 10060 123696
rect 0 123178 800 123208
rect 0 123118 6930 123178
rect 0 123088 800 123118
rect 6870 122906 6930 123118
rect 485998 123116 486004 123180
rect 486068 123178 486074 123180
rect 486200 123178 487000 123208
rect 486068 123118 487000 123178
rect 486068 123116 486074 123118
rect 486200 123088 487000 123118
rect 6870 122880 9506 122906
rect 6870 122846 10060 122880
rect 9446 122820 10060 122846
rect 478086 122436 478092 122500
rect 478156 122498 478162 122500
rect 486200 122498 487000 122528
rect 478156 122438 487000 122498
rect 478156 122436 478162 122438
rect 486200 122408 487000 122438
rect 9446 121948 10060 122008
rect 0 121818 800 121848
rect 9446 121818 9506 121948
rect 0 121758 9506 121818
rect 0 121728 800 121758
rect 478270 121756 478276 121820
rect 478340 121818 478346 121820
rect 486200 121818 487000 121848
rect 478340 121758 487000 121818
rect 478340 121756 478346 121758
rect 486200 121728 487000 121758
rect 0 121138 800 121168
rect 9446 121138 10060 121192
rect 0 121132 10060 121138
rect 486200 121140 487000 121168
rect 0 121078 9506 121132
rect 0 121048 800 121078
rect 486200 121076 486372 121140
rect 486436 121076 487000 121140
rect 486200 121048 487000 121076
rect 0 120458 800 120488
rect 486200 120460 487000 120488
rect 0 120432 9506 120458
rect 0 120398 10060 120432
rect 0 120368 800 120398
rect 9446 120372 10060 120398
rect 486200 120396 486372 120460
rect 486436 120396 487000 120460
rect 486200 120368 487000 120396
rect 0 119778 800 119808
rect 483657 119778 483723 119781
rect 486200 119778 487000 119808
rect 0 119718 9506 119778
rect 0 119688 800 119718
rect 9446 119616 9506 119718
rect 483657 119776 487000 119778
rect 483657 119720 483662 119776
rect 483718 119720 487000 119776
rect 483657 119718 487000 119720
rect 483657 119715 483723 119718
rect 486200 119688 487000 119718
rect 9446 119556 10060 119616
rect 0 119098 800 119128
rect 0 119038 9506 119098
rect 0 119008 800 119038
rect 9446 118800 9506 119038
rect 483790 119036 483796 119100
rect 483860 119098 483866 119100
rect 486200 119098 487000 119128
rect 483860 119038 487000 119098
rect 483860 119036 483866 119038
rect 486200 119008 487000 119038
rect 9446 118740 10060 118800
rect 9446 117868 10060 117928
rect 0 117738 800 117768
rect 9446 117738 9506 117868
rect 0 117678 9506 117738
rect 0 117648 800 117678
rect 0 117058 800 117088
rect 9446 117058 10060 117112
rect 0 117052 10060 117058
rect 0 116998 9506 117052
rect 0 116968 800 116998
rect 0 116378 800 116408
rect 0 116352 9506 116378
rect 0 116318 10060 116352
rect 0 116288 800 116318
rect 9446 116292 10060 116318
rect 0 115698 800 115728
rect 0 115638 9506 115698
rect 0 115608 800 115638
rect 9446 115536 9506 115638
rect 9446 115476 10060 115536
rect 0 115018 800 115048
rect 0 114958 9506 115018
rect 0 114928 800 114958
rect 9446 114720 9506 114958
rect 9446 114660 10060 114720
rect 9446 113788 10060 113848
rect 0 113658 800 113688
rect 9446 113658 9506 113788
rect 0 113598 9506 113658
rect 0 113568 800 113598
rect 0 112978 800 113008
rect 9446 112978 10060 113032
rect 0 112972 10060 112978
rect 0 112918 9506 112972
rect 0 112888 800 112918
rect 0 112298 800 112328
rect 0 112272 9506 112298
rect 0 112238 10060 112272
rect 0 112208 800 112238
rect 9446 112212 10060 112238
rect 0 111618 800 111648
rect 0 111558 9506 111618
rect 0 111528 800 111558
rect 9446 111456 9506 111558
rect 9446 111396 10060 111456
rect 0 103458 800 103488
rect 0 103398 9506 103458
rect 0 103368 800 103398
rect 9446 103176 9506 103398
rect 9446 103116 10060 103176
rect 9446 102242 10060 102302
rect 9446 102234 9506 102242
rect 6870 102174 9506 102234
rect 0 102098 800 102128
rect 6870 102098 6930 102174
rect 0 102038 6930 102098
rect 0 102008 800 102038
rect 0 101418 800 101448
rect 9446 101426 10060 101486
rect 9446 101418 9506 101426
rect 0 101358 9506 101418
rect 0 101328 800 101358
rect 0 100738 800 100768
rect 0 100678 10032 100738
rect 0 100648 800 100678
rect 0 100058 800 100088
rect 0 99998 6930 100058
rect 0 99968 800 99998
rect 6870 99922 6930 99998
rect 6870 99862 10032 99922
rect 0 99378 800 99408
rect 0 99318 6930 99378
rect 0 99288 800 99318
rect 6870 99106 6930 99318
rect 6870 99046 10032 99106
rect 9446 98162 10060 98222
rect 0 98018 800 98048
rect 9446 98018 9506 98162
rect 0 97958 9506 98018
rect 0 97928 800 97958
rect 0 97338 800 97368
rect 9446 97346 10060 97406
rect 9446 97338 9506 97346
rect 0 97278 9506 97338
rect 0 97248 800 97278
rect 0 96658 800 96688
rect 0 96598 10032 96658
rect 0 96568 800 96598
rect 0 95978 800 96008
rect 0 95918 6930 95978
rect 0 95888 800 95918
rect 6870 95842 6930 95918
rect 6870 95782 10032 95842
rect 0 95298 800 95328
rect 0 95238 4170 95298
rect 0 95208 800 95238
rect 4110 95162 4170 95238
rect 4110 95102 6930 95162
rect 6870 95026 6930 95102
rect 6870 94966 10032 95026
rect 9446 94082 10060 94142
rect 0 93938 800 93968
rect 9446 93938 9506 94082
rect 0 93878 9506 93938
rect 0 93848 800 93878
rect 0 93258 800 93288
rect 9446 93266 10060 93326
rect 9446 93258 9506 93266
rect 0 93198 9506 93258
rect 0 93168 800 93198
rect 0 92578 800 92608
rect 0 92518 10032 92578
rect 0 92488 800 92518
rect 0 91898 800 91928
rect 0 91838 6930 91898
rect 0 91808 800 91838
rect 6870 91762 6930 91838
rect 6870 91702 10032 91762
rect 6310 90884 6316 90948
rect 6380 90946 6386 90948
rect 6380 90886 10032 90946
rect 6380 90884 6386 90886
rect 481541 90538 481607 90541
rect 486200 90538 487000 90568
rect 481541 90536 487000 90538
rect 481541 90480 481546 90536
rect 481602 90480 487000 90536
rect 481541 90478 487000 90480
rect 481541 90475 481607 90478
rect 486200 90448 487000 90478
rect 7598 90068 7604 90132
rect 7668 90130 7674 90132
rect 7668 90070 10032 90130
rect 7668 90068 7674 90070
rect 484301 89858 484367 89861
rect 486200 89858 487000 89888
rect 484301 89856 487000 89858
rect 484301 89800 484306 89856
rect 484362 89800 487000 89856
rect 484301 89798 487000 89800
rect 484301 89795 484367 89798
rect 486200 89768 487000 89798
rect 54 89252 60 89316
rect 124 89314 130 89316
rect 124 89254 10032 89314
rect 124 89252 130 89254
rect 482921 89178 482987 89181
rect 486200 89178 487000 89208
rect 482921 89176 487000 89178
rect 482921 89120 482926 89176
rect 482982 89120 487000 89176
rect 482921 89118 487000 89120
rect 482921 89115 482987 89118
rect 486200 89088 487000 89118
rect 8886 88436 8892 88500
rect 8956 88498 8962 88500
rect 481449 88498 481515 88501
rect 486200 88498 487000 88528
rect 8956 88438 10032 88498
rect 481449 88496 487000 88498
rect 481449 88440 481454 88496
rect 481510 88440 487000 88496
rect 481449 88438 487000 88440
rect 8956 88436 8962 88438
rect 481449 88435 481515 88438
rect 486200 88408 487000 88438
rect 484209 87818 484275 87821
rect 486200 87818 487000 87848
rect 484209 87816 487000 87818
rect 484209 87760 484214 87816
rect 484270 87760 487000 87816
rect 484209 87758 487000 87760
rect 484209 87755 484275 87758
rect 486200 87728 487000 87758
rect 3550 87620 3556 87684
rect 3620 87682 3626 87684
rect 3620 87622 10032 87682
rect 3620 87620 3626 87622
rect 482829 87138 482895 87141
rect 486200 87138 487000 87168
rect 482829 87136 487000 87138
rect 482829 87080 482834 87136
rect 482890 87080 487000 87136
rect 482829 87078 487000 87080
rect 482829 87075 482895 87078
rect 486200 87048 487000 87078
rect 6494 86804 6500 86868
rect 6564 86866 6570 86868
rect 6564 86806 10032 86866
rect 6564 86804 6570 86806
rect 480846 86396 480852 86460
rect 480916 86458 480922 86460
rect 486200 86458 487000 86488
rect 480916 86398 487000 86458
rect 480916 86396 480922 86398
rect 486200 86368 487000 86398
rect 4654 85988 4660 86052
rect 4724 86050 4730 86052
rect 4724 85990 10032 86050
rect 4724 85988 4730 85990
rect 483606 85716 483612 85780
rect 483676 85778 483682 85780
rect 486200 85778 487000 85808
rect 483676 85718 487000 85778
rect 483676 85716 483682 85718
rect 486200 85688 487000 85718
rect 7414 85172 7420 85236
rect 7484 85234 7490 85236
rect 7484 85174 10032 85234
rect 7484 85172 7490 85174
rect 478689 85098 478755 85101
rect 486200 85098 487000 85128
rect 478689 85096 487000 85098
rect 478689 85040 478694 85096
rect 478750 85040 487000 85096
rect 478689 85038 487000 85040
rect 478689 85035 478755 85038
rect 486200 85008 487000 85038
rect 7782 84356 7788 84420
rect 7852 84418 7858 84420
rect 478781 84418 478847 84421
rect 486200 84418 487000 84448
rect 7852 84358 10032 84418
rect 478781 84416 487000 84418
rect 478781 84360 478786 84416
rect 478842 84360 487000 84416
rect 478781 84358 487000 84360
rect 7852 84356 7858 84358
rect 478781 84355 478847 84358
rect 486200 84328 487000 84358
rect 478086 83676 478092 83740
rect 478156 83738 478162 83740
rect 486200 83738 487000 83768
rect 478156 83678 487000 83738
rect 478156 83676 478162 83678
rect 486200 83648 487000 83678
rect 6126 83540 6132 83604
rect 6196 83602 6202 83604
rect 6196 83542 10032 83602
rect 6196 83540 6202 83542
rect 478270 82996 478276 83060
rect 478340 83058 478346 83060
rect 486200 83058 487000 83088
rect 478340 82998 487000 83058
rect 478340 82996 478346 82998
rect 486200 82968 487000 82998
rect 5206 82724 5212 82788
rect 5276 82786 5282 82788
rect 5276 82726 10032 82786
rect 5276 82724 5282 82726
rect 482134 82316 482140 82380
rect 482204 82378 482210 82380
rect 486200 82378 487000 82408
rect 482204 82318 487000 82378
rect 482204 82316 482210 82318
rect 486200 82288 487000 82318
rect 1894 81908 1900 81972
rect 1964 81970 1970 81972
rect 1964 81910 10032 81970
rect 1964 81908 1970 81910
rect 478454 81636 478460 81700
rect 478524 81698 478530 81700
rect 486200 81698 487000 81728
rect 478524 81638 487000 81698
rect 478524 81636 478530 81638
rect 486200 81608 487000 81638
rect 7966 81092 7972 81156
rect 8036 81154 8042 81156
rect 8036 81094 10032 81154
rect 8036 81092 8042 81094
rect 480161 81018 480227 81021
rect 486200 81018 487000 81048
rect 480161 81016 487000 81018
rect 480161 80960 480166 81016
rect 480222 80960 487000 81016
rect 480161 80958 487000 80960
rect 480161 80955 480227 80958
rect 486200 80928 487000 80958
rect 238 80276 244 80340
rect 308 80338 314 80340
rect 308 80278 10032 80338
rect 308 80276 314 80278
rect 485814 80276 485820 80340
rect 485884 80338 485890 80340
rect 486200 80338 487000 80368
rect 485884 80278 487000 80338
rect 485884 80276 485890 80278
rect 486200 80248 487000 80278
rect 482277 79658 482343 79661
rect 486200 79658 487000 79688
rect 482277 79656 487000 79658
rect 482277 79600 482282 79656
rect 482338 79600 487000 79656
rect 482277 79598 487000 79600
rect 482277 79595 482343 79598
rect 486200 79568 487000 79598
rect 4838 79460 4844 79524
rect 4908 79522 4914 79524
rect 4908 79462 10032 79522
rect 4908 79460 4914 79462
rect 479558 78916 479564 78980
rect 479628 78978 479634 78980
rect 486200 78978 487000 79008
rect 479628 78918 487000 78978
rect 479628 78916 479634 78918
rect 486200 78888 487000 78918
rect 9070 78644 9076 78708
rect 9140 78706 9146 78708
rect 9140 78646 10032 78706
rect 9140 78644 9146 78646
rect 486200 78300 487000 78328
rect 486200 78236 486556 78300
rect 486620 78236 487000 78300
rect 486200 78208 487000 78236
rect 3366 77828 3372 77892
rect 3436 77890 3442 77892
rect 3436 77830 10032 77890
rect 3436 77828 3442 77830
rect 479374 77556 479380 77620
rect 479444 77618 479450 77620
rect 486200 77618 487000 77648
rect 479444 77558 487000 77618
rect 479444 77556 479450 77558
rect 486200 77528 487000 77558
rect 5022 77012 5028 77076
rect 5092 77074 5098 77076
rect 5092 77014 10032 77074
rect 5092 77012 5098 77014
rect 481030 76876 481036 76940
rect 481100 76938 481106 76940
rect 486200 76938 487000 76968
rect 481100 76878 487000 76938
rect 481100 76876 481106 76878
rect 486200 76848 487000 76878
rect 0 76258 800 76288
rect 6310 76258 6316 76260
rect 0 76198 6316 76258
rect 0 76168 800 76198
rect 6310 76196 6316 76198
rect 6380 76196 6386 76260
rect 482318 76196 482324 76260
rect 482388 76258 482394 76260
rect 486200 76258 487000 76288
rect 482388 76198 487000 76258
rect 482388 76196 482394 76198
rect 9446 76130 10060 76190
rect 486200 76168 487000 76198
rect 790 75924 796 75988
rect 860 75986 866 75988
rect 9446 75986 9506 76130
rect 860 75926 9506 75986
rect 860 75924 866 75926
rect 54 75788 60 75852
rect 124 75850 130 75852
rect 124 75790 1042 75850
rect 124 75788 130 75790
rect 0 75578 800 75608
rect 982 75578 1042 75790
rect 0 75518 1042 75578
rect 0 75488 800 75518
rect 479742 75516 479748 75580
rect 479812 75578 479818 75580
rect 486200 75578 487000 75608
rect 479812 75518 487000 75578
rect 479812 75516 479818 75518
rect 486200 75488 487000 75518
rect 8334 75380 8340 75444
rect 8404 75442 8410 75444
rect 8404 75382 10032 75442
rect 8404 75380 8410 75382
rect 0 74898 800 74928
rect 7782 74898 7788 74900
rect 0 74838 7788 74898
rect 0 74808 800 74838
rect 7782 74836 7788 74838
rect 7852 74836 7858 74900
rect 484342 74836 484348 74900
rect 484412 74898 484418 74900
rect 486200 74898 487000 74928
rect 484412 74838 487000 74898
rect 484412 74836 484418 74838
rect 486200 74808 487000 74838
rect 6310 74564 6316 74628
rect 6380 74626 6386 74628
rect 6380 74566 10032 74626
rect 6380 74564 6386 74566
rect 0 74218 800 74248
rect 7966 74218 7972 74220
rect 0 74158 7972 74218
rect 0 74128 800 74158
rect 7966 74156 7972 74158
rect 8036 74156 8042 74220
rect 479926 74156 479932 74220
rect 479996 74218 480002 74220
rect 486200 74218 487000 74248
rect 479996 74158 487000 74218
rect 479996 74156 480002 74158
rect 486200 74128 487000 74158
rect 7782 73748 7788 73812
rect 7852 73810 7858 73812
rect 7852 73750 10032 73810
rect 7852 73748 7858 73750
rect 0 73538 800 73568
rect 5206 73538 5212 73540
rect 0 73478 5212 73538
rect 0 73448 800 73478
rect 5206 73476 5212 73478
rect 5276 73476 5282 73540
rect 484894 73476 484900 73540
rect 484964 73538 484970 73540
rect 486200 73538 487000 73568
rect 484964 73478 487000 73538
rect 484964 73476 484970 73478
rect 486200 73448 487000 73478
rect 4102 72932 4108 72996
rect 4172 72994 4178 72996
rect 4172 72934 10032 72994
rect 4172 72932 4178 72934
rect 0 72858 800 72888
rect 6494 72858 6500 72860
rect 0 72798 6500 72858
rect 0 72768 800 72798
rect 6494 72796 6500 72798
rect 6564 72796 6570 72860
rect 481398 72796 481404 72860
rect 481468 72858 481474 72860
rect 486200 72858 487000 72888
rect 481468 72798 487000 72858
rect 481468 72796 481474 72798
rect 486200 72768 487000 72798
rect 0 72178 800 72208
rect 3550 72178 3556 72180
rect 0 72118 3556 72178
rect 0 72088 800 72118
rect 3550 72116 3556 72118
rect 3620 72116 3626 72180
rect 6678 72116 6684 72180
rect 6748 72178 6754 72180
rect 6748 72118 10032 72178
rect 6748 72116 6754 72118
rect 484710 72116 484716 72180
rect 484780 72178 484786 72180
rect 486200 72178 487000 72208
rect 484780 72118 487000 72178
rect 484780 72116 484786 72118
rect 486200 72088 487000 72118
rect 0 71498 800 71528
rect 8334 71498 8340 71500
rect 0 71438 8340 71498
rect 0 71408 800 71438
rect 8334 71436 8340 71438
rect 8404 71436 8410 71500
rect 484526 71436 484532 71500
rect 484596 71498 484602 71500
rect 486200 71498 487000 71528
rect 484596 71438 487000 71498
rect 484596 71436 484602 71438
rect 486200 71408 487000 71438
rect 9446 71234 10060 71294
rect 0 70818 800 70848
rect 9446 70818 9506 71234
rect 0 70758 9506 70818
rect 0 70728 800 70758
rect 484342 70756 484348 70820
rect 484412 70818 484418 70820
rect 486200 70818 487000 70848
rect 484412 70758 487000 70818
rect 484412 70756 484418 70758
rect 486200 70728 487000 70758
rect 9446 70418 10060 70478
rect 0 70138 800 70168
rect 9446 70138 9506 70418
rect 0 70078 9506 70138
rect 0 70048 800 70078
rect 483422 70076 483428 70140
rect 483492 70138 483498 70140
rect 486200 70138 487000 70168
rect 483492 70078 487000 70138
rect 483492 70076 483498 70078
rect 486200 70048 487000 70078
rect 9446 69602 10060 69662
rect 0 69458 800 69488
rect 9446 69458 9506 69602
rect 0 69398 9506 69458
rect 0 69368 800 69398
rect 481582 69396 481588 69460
rect 481652 69458 481658 69460
rect 486200 69458 487000 69488
rect 481652 69398 487000 69458
rect 481652 69396 481658 69398
rect 486200 69368 487000 69398
rect 2078 68852 2084 68916
rect 2148 68914 2154 68916
rect 2148 68854 10032 68914
rect 2148 68852 2154 68854
rect 0 68778 800 68808
rect 0 68718 1042 68778
rect 0 68688 800 68718
rect 238 68444 244 68508
rect 308 68506 314 68508
rect 982 68506 1042 68718
rect 483238 68716 483244 68780
rect 483308 68778 483314 68780
rect 486200 68778 487000 68808
rect 483308 68718 487000 68778
rect 483308 68716 483314 68718
rect 486200 68688 487000 68718
rect 308 68446 1042 68506
rect 308 68444 314 68446
rect 481398 68234 481404 68236
rect 476968 68174 481404 68234
rect 481398 68172 481404 68174
rect 481468 68172 481474 68236
rect 0 68098 800 68128
rect 5022 68098 5028 68100
rect 0 68038 5028 68098
rect 0 68008 800 68038
rect 5022 68036 5028 68038
rect 5092 68036 5098 68100
rect 9254 68036 9260 68100
rect 9324 68098 9330 68100
rect 9324 68038 10032 68098
rect 9324 68036 9330 68038
rect 478638 68036 478644 68100
rect 478708 68098 478714 68100
rect 486200 68098 487000 68128
rect 478708 68038 487000 68098
rect 478708 68036 478714 68038
rect 486200 68008 487000 68038
rect 484158 67962 484164 67964
rect 476968 67902 484164 67962
rect 484158 67900 484164 67902
rect 484228 67900 484234 67964
rect 481582 67690 481588 67692
rect 476968 67630 481588 67690
rect 481582 67628 481588 67630
rect 481652 67628 481658 67692
rect 480294 67492 480300 67556
rect 480364 67554 480370 67556
rect 481449 67554 481515 67557
rect 480364 67552 481515 67554
rect 480364 67496 481454 67552
rect 481510 67496 481515 67552
rect 480364 67494 481515 67496
rect 480364 67492 480370 67494
rect 481449 67491 481515 67494
rect 481582 67492 481588 67556
rect 481652 67554 481658 67556
rect 482829 67554 482895 67557
rect 481652 67552 482895 67554
rect 481652 67496 482834 67552
rect 482890 67496 482895 67552
rect 481652 67494 482895 67496
rect 481652 67492 481658 67494
rect 482829 67491 482895 67494
rect 483054 67492 483060 67556
rect 483124 67554 483130 67556
rect 484209 67554 484275 67557
rect 483124 67552 484275 67554
rect 483124 67496 484214 67552
rect 484270 67496 484275 67552
rect 483124 67494 484275 67496
rect 483124 67492 483130 67494
rect 484209 67491 484275 67494
rect 0 67418 800 67448
rect 7598 67418 7604 67420
rect 0 67358 7604 67418
rect 0 67328 800 67358
rect 7598 67356 7604 67358
rect 7668 67356 7674 67420
rect 481766 67356 481772 67420
rect 481836 67418 481842 67420
rect 486200 67418 487000 67448
rect 481836 67358 487000 67418
rect 481836 67356 481842 67358
rect 476940 67290 477418 67350
rect 486200 67328 487000 67358
rect 5574 67220 5580 67284
rect 5644 67282 5650 67284
rect 477358 67282 477418 67290
rect 483238 67282 483244 67284
rect 5644 67222 10032 67282
rect 477358 67222 483244 67282
rect 5644 67220 5650 67222
rect 483238 67220 483244 67222
rect 483308 67220 483314 67284
rect 483422 67146 483428 67148
rect 476968 67086 483428 67146
rect 483422 67084 483428 67086
rect 483492 67084 483498 67148
rect 484342 66874 484348 66876
rect 476968 66814 484348 66874
rect 484342 66812 484348 66814
rect 484412 66812 484418 66876
rect 0 66738 800 66768
rect 4654 66738 4660 66740
rect 0 66678 4660 66738
rect 0 66648 800 66678
rect 4654 66676 4660 66678
rect 4724 66676 4730 66740
rect 483238 66676 483244 66740
rect 483308 66738 483314 66740
rect 486200 66738 487000 66768
rect 483308 66678 487000 66738
rect 483308 66676 483314 66678
rect 486200 66648 487000 66678
rect 476940 66474 477418 66534
rect 3550 66404 3556 66468
rect 3620 66466 3626 66468
rect 477358 66466 477418 66474
rect 486182 66466 486188 66468
rect 3620 66406 10032 66466
rect 477358 66406 486188 66466
rect 3620 66404 3626 66406
rect 486182 66404 486188 66406
rect 486252 66404 486258 66468
rect 484526 66330 484532 66332
rect 476968 66270 484532 66330
rect 484526 66268 484532 66270
rect 484596 66268 484602 66332
rect 480161 66196 480227 66197
rect 480110 66194 480116 66196
rect 480070 66134 480116 66194
rect 480180 66192 480227 66196
rect 480222 66136 480227 66192
rect 480110 66132 480116 66134
rect 480180 66132 480227 66136
rect 480161 66131 480227 66132
rect 0 66058 800 66088
rect 5574 66058 5580 66060
rect 0 65998 5580 66058
rect 0 65968 800 65998
rect 5574 65996 5580 65998
rect 5644 65996 5650 66060
rect 483238 66058 483244 66060
rect 476968 65998 483244 66058
rect 483238 65996 483244 65998
rect 483308 65996 483314 66060
rect 484158 65996 484164 66060
rect 484228 66058 484234 66060
rect 486200 66058 487000 66088
rect 484228 65998 487000 66058
rect 484228 65996 484234 65998
rect 486200 65968 487000 65998
rect 483238 65860 483244 65924
rect 483308 65922 483314 65924
rect 484301 65922 484367 65925
rect 483308 65920 484367 65922
rect 483308 65864 484306 65920
rect 484362 65864 484367 65920
rect 483308 65862 484367 65864
rect 483308 65860 483314 65862
rect 484301 65859 484367 65862
rect 484710 65786 484716 65788
rect 476968 65726 484716 65786
rect 484710 65724 484716 65726
rect 484780 65724 484786 65788
rect 479558 65514 479564 65516
rect 476968 65454 479564 65514
rect 479558 65452 479564 65454
rect 479628 65452 479634 65516
rect 0 65378 800 65408
rect 4102 65378 4108 65380
rect 0 65318 4108 65378
rect 0 65288 800 65318
rect 4102 65316 4108 65318
rect 4172 65316 4178 65380
rect 477350 65316 477356 65380
rect 477420 65378 477426 65380
rect 486200 65378 487000 65408
rect 477420 65318 487000 65378
rect 477420 65316 477426 65318
rect 486200 65288 487000 65318
rect 478638 65242 478644 65244
rect 476968 65182 478644 65242
rect 478638 65180 478644 65182
rect 478708 65180 478714 65244
rect 484894 64970 484900 64972
rect 476968 64910 484900 64970
rect 484894 64908 484900 64910
rect 484964 64908 484970 64972
rect 0 64698 800 64728
rect 9254 64698 9260 64700
rect 0 64638 9260 64698
rect 0 64608 800 64638
rect 9254 64636 9260 64638
rect 9324 64636 9330 64700
rect 481766 64698 481772 64700
rect 476968 64638 481772 64698
rect 481766 64636 481772 64638
rect 481836 64636 481842 64700
rect 484342 64636 484348 64700
rect 484412 64698 484418 64700
rect 486200 64698 487000 64728
rect 484412 64638 487000 64698
rect 484412 64636 484418 64638
rect 486200 64608 487000 64638
rect 479926 64426 479932 64428
rect 476968 64366 479932 64426
rect 479926 64364 479932 64366
rect 479996 64364 480002 64428
rect 482277 64154 482343 64157
rect 484158 64154 484164 64156
rect 476968 64152 482343 64154
rect 476968 64096 482282 64152
rect 482338 64096 482343 64152
rect 476968 64094 482343 64096
rect 482277 64091 482343 64094
rect 482510 64094 484164 64154
rect 0 64018 800 64048
rect 6678 64018 6684 64020
rect 0 63958 6684 64018
rect 0 63928 800 63958
rect 6678 63956 6684 63958
rect 6748 63956 6754 64020
rect 482510 63882 482570 64094
rect 484158 64092 484164 64094
rect 484228 64092 484234 64156
rect 486200 64018 487000 64048
rect 476968 63822 482570 63882
rect 483062 63958 487000 64018
rect 478689 63748 478755 63749
rect 478638 63684 478644 63748
rect 478708 63746 478755 63748
rect 478708 63744 478800 63746
rect 478750 63688 478800 63744
rect 478708 63686 478800 63688
rect 478708 63684 478755 63686
rect 478689 63683 478755 63684
rect 479742 63610 479748 63612
rect 476968 63550 479748 63610
rect 479742 63548 479748 63550
rect 479812 63548 479818 63612
rect 0 63338 800 63368
rect 7782 63338 7788 63340
rect 0 63278 7788 63338
rect 0 63248 800 63278
rect 7782 63276 7788 63278
rect 7852 63276 7858 63340
rect 483062 63338 483122 63958
rect 486200 63928 487000 63958
rect 486200 63338 487000 63368
rect 476968 63278 483122 63338
rect 483246 63278 487000 63338
rect 477166 63140 477172 63204
rect 477236 63202 477242 63204
rect 483246 63202 483306 63278
rect 486200 63248 487000 63278
rect 477236 63142 483306 63202
rect 477236 63140 477242 63142
rect 482318 63066 482324 63068
rect 476968 63006 482324 63066
rect 482318 63004 482324 63006
rect 482388 63004 482394 63068
rect 481030 62794 481036 62796
rect 476968 62734 481036 62794
rect 481030 62732 481036 62734
rect 481100 62732 481106 62796
rect 0 62658 800 62688
rect 4838 62658 4844 62660
rect 0 62598 4844 62658
rect 0 62568 800 62598
rect 4838 62596 4844 62598
rect 4908 62596 4914 62660
rect 483422 62596 483428 62660
rect 483492 62658 483498 62660
rect 486200 62658 487000 62688
rect 483492 62598 487000 62658
rect 483492 62596 483498 62598
rect 486200 62568 487000 62598
rect 477350 62522 477356 62524
rect 476968 62462 477356 62522
rect 477350 62460 477356 62462
rect 477420 62460 477426 62524
rect 485262 62386 485268 62388
rect 480210 62326 485268 62386
rect 480210 62250 480270 62326
rect 485262 62324 485268 62326
rect 485332 62324 485338 62388
rect 476968 62190 480270 62250
rect 480478 62188 480484 62252
rect 480548 62250 480554 62252
rect 481541 62250 481607 62253
rect 480548 62248 481607 62250
rect 480548 62192 481546 62248
rect 481602 62192 481607 62248
rect 480548 62190 481607 62192
rect 480548 62188 480554 62190
rect 481541 62187 481607 62190
rect 481766 62188 481772 62252
rect 481836 62250 481842 62252
rect 482921 62250 482987 62253
rect 481836 62248 482987 62250
rect 481836 62192 482926 62248
rect 482982 62192 482987 62248
rect 481836 62190 482987 62192
rect 481836 62188 481842 62190
rect 482921 62187 482987 62190
rect 0 61978 800 62008
rect 6310 61978 6316 61980
rect 0 61918 6316 61978
rect 0 61888 800 61918
rect 6310 61916 6316 61918
rect 6380 61916 6386 61980
rect 480110 61978 480116 61980
rect 476968 61918 480116 61978
rect 480110 61916 480116 61918
rect 480180 61916 480186 61980
rect 481582 61916 481588 61980
rect 481652 61978 481658 61980
rect 486200 61978 487000 62008
rect 481652 61918 487000 61978
rect 481652 61916 481658 61918
rect 486200 61888 487000 61918
rect 484342 61706 484348 61708
rect 476968 61646 484348 61706
rect 484342 61644 484348 61646
rect 484412 61644 484418 61708
rect 479374 61434 479380 61436
rect 476968 61374 479380 61434
rect 479374 61372 479380 61374
rect 479444 61372 479450 61436
rect 0 61300 800 61328
rect 0 61236 796 61300
rect 860 61236 866 61300
rect 486200 61298 487000 61328
rect 480210 61238 487000 61298
rect 0 61208 800 61236
rect 480210 61162 480270 61238
rect 486200 61208 487000 61238
rect 476968 61102 480270 61162
rect 483422 60890 483428 60892
rect 476968 60830 483428 60890
rect 483422 60828 483428 60830
rect 483492 60828 483498 60892
rect 1342 60692 1348 60756
rect 1412 60754 1418 60756
rect 7414 60754 7420 60756
rect 1412 60694 7420 60754
rect 1412 60692 1418 60694
rect 7414 60692 7420 60694
rect 7484 60692 7490 60756
rect 0 60618 800 60648
rect 9070 60618 9076 60620
rect 0 60558 9076 60618
rect 0 60528 800 60558
rect 9070 60556 9076 60558
rect 9140 60556 9146 60620
rect 477902 60556 477908 60620
rect 477972 60618 477978 60620
rect 478781 60618 478847 60621
rect 486200 60618 487000 60648
rect 477972 60616 478847 60618
rect 477972 60560 478786 60616
rect 478842 60560 478847 60616
rect 477972 60558 478847 60560
rect 477972 60556 477978 60558
rect 478781 60555 478847 60558
rect 483246 60558 487000 60618
rect 476940 60490 477418 60550
rect 477358 60482 477418 60490
rect 481582 60482 481588 60484
rect 477358 60422 481588 60482
rect 481582 60420 481588 60422
rect 481652 60420 481658 60484
rect 477166 60346 477172 60348
rect 476968 60286 477172 60346
rect 477166 60284 477172 60286
rect 477236 60284 477242 60348
rect 483246 60074 483306 60558
rect 486200 60528 487000 60558
rect 476968 60014 483306 60074
rect 0 59938 800 59968
rect 1894 59938 1900 59940
rect 0 59878 1900 59938
rect 0 59848 800 59878
rect 1894 59876 1900 59878
rect 1964 59876 1970 59940
rect 486200 59938 487000 59968
rect 480210 59878 487000 59938
rect 480210 59802 480270 59878
rect 486200 59848 487000 59878
rect 476968 59742 480270 59802
rect 478454 59530 478460 59532
rect 476968 59470 478460 59530
rect 478454 59468 478460 59470
rect 478524 59468 478530 59532
rect 0 59258 800 59288
rect 6126 59258 6132 59260
rect 0 59198 6132 59258
rect 0 59168 800 59198
rect 6126 59196 6132 59198
rect 6196 59196 6202 59260
rect 486200 59258 487000 59288
rect 476968 59198 487000 59258
rect 486200 59168 487000 59198
rect 482134 58986 482140 58988
rect 476968 58926 482140 58986
rect 482134 58924 482140 58926
rect 482204 58924 482210 58988
rect 478270 58714 478276 58716
rect 476968 58654 478276 58714
rect 478270 58652 478276 58654
rect 478340 58652 478346 58716
rect 0 58578 800 58608
rect 1342 58578 1348 58580
rect 0 58518 1348 58578
rect 0 58488 800 58518
rect 1342 58516 1348 58518
rect 1412 58516 1418 58580
rect 486200 58578 487000 58608
rect 480210 58518 487000 58578
rect 480210 58442 480270 58518
rect 486200 58488 487000 58518
rect 476968 58382 480270 58442
rect 478086 58170 478092 58172
rect 476968 58110 478092 58170
rect 478086 58108 478092 58110
rect 478156 58108 478162 58172
rect 9446 58042 10060 58102
rect 9446 58034 9506 58042
rect 6870 57974 9506 58034
rect 0 57898 800 57928
rect 6870 57898 6930 57974
rect 486200 57898 487000 57928
rect 0 57838 6930 57898
rect 476968 57838 487000 57898
rect 0 57808 800 57838
rect 486200 57808 487000 57838
rect 477902 57626 477908 57628
rect 476968 57566 477908 57626
rect 477902 57564 477908 57566
rect 477972 57564 477978 57628
rect 478638 57354 478644 57356
rect 476968 57294 478644 57354
rect 478638 57292 478644 57294
rect 478708 57292 478714 57356
rect 0 57218 800 57248
rect 9446 57226 10060 57286
rect 9446 57218 9506 57226
rect 486200 57218 487000 57248
rect 0 57158 9506 57218
rect 480210 57158 487000 57218
rect 0 57128 800 57158
rect 480210 57082 480270 57158
rect 486200 57128 487000 57158
rect 476968 57022 480270 57082
rect 483606 56810 483612 56812
rect 476968 56750 483612 56810
rect 483606 56748 483612 56750
rect 483676 56748 483682 56812
rect 8886 56674 8892 56676
rect 1350 56614 8892 56674
rect 0 56538 800 56568
rect 1350 56538 1410 56614
rect 8886 56612 8892 56614
rect 8956 56612 8962 56676
rect 486200 56538 487000 56568
rect 0 56478 1410 56538
rect 476968 56478 487000 56538
rect 0 56448 800 56478
rect 9446 56410 10060 56470
rect 486200 56448 487000 56478
rect 0 55858 800 55888
rect 9446 55858 9506 56410
rect 480846 56266 480852 56268
rect 476968 56206 480852 56266
rect 480846 56204 480852 56206
rect 480916 56204 480922 56268
rect 481950 55994 481956 55996
rect 476968 55934 481956 55994
rect 481950 55932 481956 55934
rect 482020 55932 482026 55996
rect 486200 55858 487000 55888
rect 0 55798 9506 55858
rect 480210 55798 487000 55858
rect 0 55768 800 55798
rect 480210 55722 480270 55798
rect 486200 55768 487000 55798
rect 476968 55662 480270 55722
rect 9446 55594 10060 55654
rect 9446 55314 9506 55594
rect 483054 55450 483060 55452
rect 476968 55390 483060 55450
rect 483054 55388 483060 55390
rect 483124 55388 483130 55452
rect 5582 55254 9506 55314
rect 0 55178 800 55208
rect 5582 55178 5642 55254
rect 486200 55178 487000 55208
rect 0 55118 5642 55178
rect 476968 55118 487000 55178
rect 0 55088 800 55118
rect 486200 55088 487000 55118
rect 480294 54906 480300 54908
rect 476968 54846 480300 54906
rect 480294 54844 480300 54846
rect 480364 54844 480370 54908
rect 9446 54778 10060 54838
rect 0 54498 800 54528
rect 9446 54498 9506 54778
rect 481766 54634 481772 54636
rect 476968 54574 481772 54634
rect 481766 54572 481772 54574
rect 481836 54572 481842 54636
rect 486200 54498 487000 54528
rect 0 54438 9506 54498
rect 480210 54438 487000 54498
rect 0 54408 800 54438
rect 480210 54362 480270 54438
rect 486200 54408 487000 54438
rect 476968 54302 480270 54362
rect 483238 54090 483244 54092
rect 476968 54030 483244 54090
rect 483238 54028 483244 54030
rect 483308 54028 483314 54092
rect 9446 53962 10060 54022
rect 9446 53954 9506 53962
rect 6870 53894 9506 53954
rect 0 53818 800 53848
rect 6870 53818 6930 53894
rect 486200 53818 487000 53848
rect 0 53758 6930 53818
rect 476968 53758 487000 53818
rect 0 53728 800 53758
rect 486200 53728 487000 53758
rect 480478 53546 480484 53548
rect 476968 53486 480484 53546
rect 480478 53484 480484 53486
rect 480548 53484 480554 53548
rect 0 53138 800 53168
rect 9446 53146 10060 53206
rect 476940 53146 477418 53206
rect 9446 53138 9506 53146
rect 0 53078 9506 53138
rect 477358 53138 477418 53146
rect 486200 53138 487000 53168
rect 477358 53078 487000 53138
rect 0 53048 800 53078
rect 486200 53048 487000 53078
rect 483054 53002 483060 53004
rect 476968 52942 483060 53002
rect 483054 52940 483060 52942
rect 483124 52940 483130 53004
rect 476968 52670 483306 52730
rect 0 52458 800 52488
rect 3550 52458 3556 52460
rect 0 52398 3556 52458
rect 0 52368 800 52398
rect 3550 52396 3556 52398
rect 3620 52396 3626 52460
rect 480846 52458 480852 52460
rect 476968 52398 480852 52458
rect 480846 52396 480852 52398
rect 480916 52396 480922 52460
rect 483246 52458 483306 52670
rect 486200 52458 487000 52488
rect 483246 52398 487000 52458
rect 9446 52330 10060 52390
rect 486200 52368 487000 52398
rect 0 51778 800 51808
rect 9446 51778 9506 52330
rect 483238 52186 483244 52188
rect 476968 52126 483244 52186
rect 483238 52124 483244 52126
rect 483308 52124 483314 52188
rect 476940 51786 477418 51846
rect 0 51718 9506 51778
rect 477358 51778 477418 51786
rect 486200 51778 487000 51808
rect 477358 51718 487000 51778
rect 0 51688 800 51718
rect 486200 51688 487000 51718
rect 481766 51642 481772 51644
rect 476968 51582 481772 51642
rect 481766 51580 481772 51582
rect 481836 51580 481842 51644
rect 9446 51514 10060 51574
rect 0 51098 800 51128
rect 9446 51098 9506 51514
rect 476968 51310 483306 51370
rect 483246 51098 483306 51310
rect 486200 51098 487000 51128
rect 0 51038 9506 51098
rect 476968 51038 483122 51098
rect 483246 51038 487000 51098
rect 0 51008 800 51038
rect 483062 50962 483122 51038
rect 486200 51008 487000 51038
rect 483606 50962 483612 50964
rect 483062 50902 483612 50962
rect 483606 50900 483612 50902
rect 483676 50900 483682 50964
rect 481582 50826 481588 50828
rect 476968 50766 481588 50826
rect 481582 50764 481588 50766
rect 481652 50764 481658 50828
rect 9446 50698 10060 50758
rect 0 50418 800 50448
rect 9446 50418 9506 50698
rect 476940 50426 477418 50486
rect 0 50358 9506 50418
rect 477358 50418 477418 50426
rect 486200 50418 487000 50448
rect 477358 50358 487000 50418
rect 0 50328 800 50358
rect 486200 50328 487000 50358
rect 481030 50282 481036 50284
rect 476968 50222 481036 50282
rect 481030 50220 481036 50222
rect 481100 50220 481106 50284
rect 476968 49950 483306 50010
rect 9446 49882 10060 49942
rect 0 49738 800 49768
rect 9446 49738 9506 49882
rect 482134 49738 482140 49740
rect 0 49678 9506 49738
rect 476968 49678 482140 49738
rect 0 49648 800 49678
rect 482134 49676 482140 49678
rect 482204 49676 482210 49740
rect 483246 49738 483306 49950
rect 486200 49738 487000 49768
rect 483246 49678 487000 49738
rect 486200 49648 487000 49678
rect 483790 49466 483796 49468
rect 476968 49406 483796 49466
rect 483790 49404 483796 49406
rect 483860 49404 483866 49468
rect 0 49058 800 49088
rect 9446 49066 10060 49126
rect 476940 49066 477418 49126
rect 9446 49058 9506 49066
rect 0 48998 9506 49058
rect 477358 49058 477418 49066
rect 486200 49058 487000 49088
rect 477358 48998 487000 49058
rect 0 48968 800 48998
rect 486200 48968 487000 48998
rect 481214 48922 481220 48924
rect 476968 48862 481220 48922
rect 481214 48860 481220 48862
rect 481284 48860 481290 48924
rect 476968 48590 483306 48650
rect 0 48378 800 48408
rect 2078 48378 2084 48380
rect 0 48318 2084 48378
rect 0 48288 800 48318
rect 2078 48316 2084 48318
rect 2148 48316 2154 48380
rect 482318 48378 482324 48380
rect 6870 48318 10032 48378
rect 476968 48318 482324 48378
rect 1342 48180 1348 48244
rect 1412 48242 1418 48244
rect 3366 48242 3372 48244
rect 1412 48182 3372 48242
rect 1412 48180 1418 48182
rect 3366 48180 3372 48182
rect 3436 48180 3442 48244
rect 0 47698 800 47728
rect 6870 47698 6930 48318
rect 482318 48316 482324 48318
rect 482388 48316 482394 48380
rect 483246 48378 483306 48590
rect 486200 48378 487000 48408
rect 483246 48318 487000 48378
rect 486200 48288 487000 48318
rect 480846 48180 480852 48244
rect 480916 48242 480922 48244
rect 481541 48242 481607 48245
rect 480916 48240 481607 48242
rect 480916 48184 481546 48240
rect 481602 48184 481607 48240
rect 480916 48182 481607 48184
rect 480916 48180 480922 48182
rect 481541 48179 481607 48182
rect 481398 48106 481404 48108
rect 476968 48046 481404 48106
rect 481398 48044 481404 48046
rect 481468 48044 481474 48108
rect 476940 47706 477418 47766
rect 0 47638 6930 47698
rect 477358 47698 477418 47706
rect 486200 47698 487000 47728
rect 477358 47638 487000 47698
rect 0 47608 800 47638
rect 486200 47608 487000 47638
rect 480846 47562 480852 47564
rect 476968 47502 480852 47562
rect 480846 47500 480852 47502
rect 480916 47500 480922 47564
rect 9446 47434 10060 47494
rect 0 47018 800 47048
rect 9446 47018 9506 47434
rect 477217 47426 477283 47429
rect 479926 47426 479932 47428
rect 477217 47424 479932 47426
rect 477217 47368 477222 47424
rect 477278 47368 479932 47424
rect 477217 47366 479932 47368
rect 477217 47363 477283 47366
rect 479926 47364 479932 47366
rect 479996 47364 480002 47428
rect 476940 47162 477418 47222
rect 477217 47018 477283 47021
rect 0 46958 9506 47018
rect 476968 47016 477283 47018
rect 476968 46960 477222 47016
rect 477278 46960 477283 47016
rect 476968 46958 477283 46960
rect 477358 47018 477418 47162
rect 486200 47018 487000 47048
rect 477358 46958 487000 47018
rect 0 46928 800 46958
rect 477217 46955 477283 46958
rect 486200 46928 487000 46958
rect 479190 46746 479196 46748
rect 476968 46686 479196 46746
rect 479190 46684 479196 46686
rect 479260 46684 479266 46748
rect 9446 46618 10060 46678
rect 0 46338 800 46368
rect 9446 46338 9506 46618
rect 476940 46346 477418 46406
rect 0 46278 9506 46338
rect 477358 46338 477418 46346
rect 486200 46338 487000 46368
rect 477358 46278 487000 46338
rect 0 46248 800 46278
rect 486200 46248 487000 46278
rect 479558 46202 479564 46204
rect 476968 46142 479564 46202
rect 479558 46140 479564 46142
rect 479628 46140 479634 46204
rect 9446 45802 10060 45862
rect 476940 45802 477418 45862
rect 0 45658 800 45688
rect 9446 45658 9506 45802
rect 477358 45794 477418 45802
rect 477358 45734 480270 45794
rect 479374 45658 479380 45660
rect 0 45598 9506 45658
rect 476968 45598 479380 45658
rect 0 45568 800 45598
rect 479374 45596 479380 45598
rect 479444 45596 479450 45660
rect 480210 45658 480270 45734
rect 486200 45658 487000 45688
rect 480210 45598 487000 45658
rect 486200 45568 487000 45598
rect 479742 45386 479748 45388
rect 476968 45326 479748 45386
rect 479742 45324 479748 45326
rect 479812 45324 479818 45388
rect 0 44978 800 45008
rect 9446 44986 10060 45046
rect 476940 44986 477418 45046
rect 9446 44978 9506 44986
rect 0 44918 9506 44978
rect 477358 44978 477418 44986
rect 486200 44978 487000 45008
rect 477358 44918 487000 44978
rect 0 44888 800 44918
rect 486200 44888 487000 44918
rect 476940 44714 477418 44774
rect 477358 44706 477418 44714
rect 486417 44706 486483 44709
rect 477358 44704 486483 44706
rect 477358 44648 486422 44704
rect 486478 44648 486483 44704
rect 477358 44646 486483 44648
rect 486417 44643 486483 44646
rect 476968 44510 483306 44570
rect 479926 44372 479932 44436
rect 479996 44434 480002 44436
rect 480161 44434 480227 44437
rect 479996 44432 480227 44434
rect 479996 44376 480166 44432
rect 480222 44376 480227 44432
rect 479996 44374 480227 44376
rect 479996 44372 480002 44374
rect 480161 44371 480227 44374
rect 0 44298 800 44328
rect 1342 44298 1348 44300
rect 0 44238 1348 44298
rect 0 44208 800 44238
rect 1342 44236 1348 44238
rect 1412 44236 1418 44300
rect 483105 44298 483171 44301
rect 6870 44238 10032 44298
rect 476968 44296 483171 44298
rect 476968 44240 483110 44296
rect 483166 44240 483171 44296
rect 476968 44238 483171 44240
rect 483246 44298 483306 44510
rect 486200 44298 487000 44328
rect 483246 44238 487000 44298
rect 0 43618 800 43648
rect 6870 43618 6930 44238
rect 483105 44235 483171 44238
rect 486200 44208 487000 44238
rect 485630 44026 485636 44028
rect 476968 43966 485636 44026
rect 485630 43964 485636 43966
rect 485700 43964 485706 44028
rect 476940 43626 477418 43686
rect 0 43558 6930 43618
rect 477358 43618 477418 43626
rect 486200 43618 487000 43648
rect 477358 43558 487000 43618
rect 0 43528 800 43558
rect 486200 43528 487000 43558
rect 478086 43482 478092 43484
rect 476968 43422 478092 43482
rect 478086 43420 478092 43422
rect 478156 43420 478162 43484
rect 9446 43354 10060 43414
rect 0 42938 800 42968
rect 9446 42938 9506 43354
rect 483054 43284 483060 43348
rect 483124 43346 483130 43348
rect 484301 43346 484367 43349
rect 483124 43344 484367 43346
rect 483124 43288 484306 43344
rect 484362 43288 484367 43344
rect 483124 43286 484367 43288
rect 483124 43284 483130 43286
rect 484301 43283 484367 43286
rect 483289 43210 483355 43213
rect 476968 43208 483355 43210
rect 476968 43152 483294 43208
rect 483350 43152 483355 43208
rect 476968 43150 483355 43152
rect 483289 43147 483355 43150
rect 485998 43074 486004 43076
rect 480210 43014 486004 43074
rect 480210 42938 480270 43014
rect 485998 43012 486004 43014
rect 486068 43012 486074 43076
rect 0 42878 9506 42938
rect 476968 42878 480270 42938
rect 483289 42938 483355 42941
rect 486200 42938 487000 42968
rect 483289 42936 487000 42938
rect 483289 42880 483294 42936
rect 483350 42880 487000 42936
rect 483289 42878 487000 42880
rect 0 42848 800 42878
rect 483289 42875 483355 42878
rect 486200 42848 487000 42878
rect 478270 42666 478276 42668
rect 476968 42606 478276 42666
rect 478270 42604 478276 42606
rect 478340 42604 478346 42668
rect 9446 42538 10060 42598
rect 0 42258 800 42288
rect 9446 42258 9506 42538
rect 476940 42266 477418 42326
rect 0 42198 9506 42258
rect 477358 42258 477418 42266
rect 486200 42258 487000 42288
rect 477358 42198 487000 42258
rect 0 42168 800 42198
rect 486200 42168 487000 42198
rect 485998 42122 486004 42124
rect 476968 42062 486004 42122
rect 485998 42060 486004 42062
rect 486068 42060 486074 42124
rect 9446 41722 10060 41782
rect 476940 41722 477418 41782
rect 0 41578 800 41608
rect 9446 41578 9506 41722
rect 0 41518 9506 41578
rect 477358 41578 477418 41722
rect 486200 41578 487000 41608
rect 477358 41518 487000 41578
rect 0 41488 800 41518
rect 476902 41448 476908 41512
rect 476972 41448 476978 41512
rect 486200 41488 487000 41518
rect 481766 41380 481772 41444
rect 481836 41442 481842 41444
rect 482921 41442 482987 41445
rect 481836 41440 482987 41442
rect 481836 41384 482926 41440
rect 482982 41384 482987 41440
rect 481836 41382 482987 41384
rect 481836 41380 481842 41382
rect 482921 41379 482987 41382
rect 483238 41380 483244 41444
rect 483308 41442 483314 41444
rect 484209 41442 484275 41445
rect 483308 41440 484275 41442
rect 483308 41384 484214 41440
rect 484270 41384 484275 41440
rect 483308 41382 484275 41384
rect 483308 41380 483314 41382
rect 484209 41379 484275 41382
rect 485446 41306 485452 41308
rect 476968 41246 485452 41306
rect 485446 41244 485452 41246
rect 485516 41244 485522 41308
rect 0 40898 800 40928
rect 9446 40906 10060 40966
rect 476940 40906 477418 40966
rect 9446 40898 9506 40906
rect 0 40838 9506 40898
rect 477358 40898 477418 40906
rect 486200 40898 487000 40928
rect 477358 40838 487000 40898
rect 0 40808 800 40838
rect 486200 40808 487000 40838
rect 484894 40762 484900 40764
rect 476968 40702 484900 40762
rect 484894 40700 484900 40702
rect 484964 40700 484970 40764
rect 476940 40362 477418 40422
rect 477358 40354 477418 40362
rect 477358 40294 480270 40354
rect 0 40218 800 40248
rect 480210 40218 480270 40294
rect 486200 40218 487000 40248
rect 0 40158 10032 40218
rect 480210 40158 487000 40218
rect 0 40128 800 40158
rect 476940 40090 477418 40150
rect 486200 40128 487000 40158
rect 477358 40082 477418 40090
rect 484710 40082 484716 40084
rect 477358 40022 484716 40082
rect 484710 40020 484716 40022
rect 484780 40020 484786 40084
rect 479190 39884 479196 39948
rect 479260 39946 479266 39948
rect 480069 39946 480135 39949
rect 479260 39944 480135 39946
rect 479260 39888 480074 39944
rect 480130 39888 480135 39944
rect 479260 39886 480135 39888
rect 479260 39884 479266 39886
rect 480069 39883 480135 39886
rect 481582 39884 481588 39948
rect 481652 39946 481658 39948
rect 482829 39946 482895 39949
rect 481652 39944 482895 39946
rect 481652 39888 482834 39944
rect 482890 39888 482895 39944
rect 481652 39886 482895 39888
rect 481652 39884 481658 39886
rect 482829 39883 482895 39886
rect 476940 39818 477418 39878
rect 477358 39810 477418 39818
rect 484526 39810 484532 39812
rect 477358 39750 484532 39810
rect 484526 39748 484532 39750
rect 484596 39748 484602 39812
rect 0 39538 800 39568
rect 476940 39546 477418 39606
rect 477358 39538 477418 39546
rect 486200 39538 487000 39568
rect 0 39478 6930 39538
rect 477358 39478 487000 39538
rect 0 39448 800 39478
rect 6870 39402 6930 39478
rect 486200 39448 487000 39478
rect 6870 39342 10032 39402
rect 476940 39274 477418 39334
rect 477358 39266 477418 39274
rect 484342 39266 484348 39268
rect 477358 39206 484348 39266
rect 484342 39204 484348 39206
rect 484412 39204 484418 39268
rect 476940 39002 477418 39062
rect 477358 38994 477418 39002
rect 477358 38934 480270 38994
rect 0 38858 800 38888
rect 480210 38858 480270 38934
rect 486200 38858 487000 38888
rect 0 38798 4170 38858
rect 480210 38798 487000 38858
rect 0 38768 800 38798
rect 4110 38586 4170 38798
rect 476940 38730 477418 38790
rect 486200 38768 487000 38798
rect 477358 38722 477418 38730
rect 485078 38722 485084 38724
rect 477358 38662 485084 38722
rect 485078 38660 485084 38662
rect 485148 38660 485154 38724
rect 4110 38526 10032 38586
rect 0 38178 800 38208
rect 0 38118 6930 38178
rect 0 38088 800 38118
rect 6870 37770 6930 38118
rect 484342 38116 484348 38180
rect 484412 38178 484418 38180
rect 486200 38178 487000 38208
rect 484412 38118 487000 38178
rect 484412 38116 484418 38118
rect 486200 38088 487000 38118
rect 6870 37710 10032 37770
rect 0 37498 800 37528
rect 0 37438 4170 37498
rect 0 37408 800 37438
rect 4110 37226 4170 37438
rect 484526 37436 484532 37500
rect 484596 37498 484602 37500
rect 486200 37498 487000 37528
rect 484596 37438 487000 37498
rect 484596 37436 484602 37438
rect 486200 37408 487000 37438
rect 4110 37166 6930 37226
rect 6870 36954 6930 37166
rect 6870 36894 10032 36954
rect 0 36818 800 36848
rect 8334 36818 8340 36820
rect 0 36758 8340 36818
rect 0 36728 800 36758
rect 8334 36756 8340 36758
rect 8404 36756 8410 36820
rect 484710 36756 484716 36820
rect 484780 36818 484786 36820
rect 486200 36818 487000 36848
rect 484780 36758 487000 36818
rect 484780 36756 484786 36758
rect 486200 36728 487000 36758
rect 0 36138 800 36168
rect 0 36078 10032 36138
rect 0 36048 800 36078
rect 484894 36076 484900 36140
rect 484964 36138 484970 36140
rect 486200 36138 487000 36168
rect 484964 36078 487000 36138
rect 484964 36076 484970 36078
rect 486200 36048 487000 36078
rect 0 35458 800 35488
rect 0 35398 6930 35458
rect 0 35368 800 35398
rect 6870 35322 6930 35398
rect 485446 35396 485452 35460
rect 485516 35458 485522 35460
rect 486200 35458 487000 35488
rect 485516 35398 487000 35458
rect 485516 35396 485522 35398
rect 486200 35368 487000 35398
rect 6870 35262 10032 35322
rect 0 34778 800 34808
rect 0 34718 4170 34778
rect 0 34688 800 34718
rect 4110 34506 4170 34718
rect 476982 34716 476988 34780
rect 477052 34778 477058 34780
rect 486200 34778 487000 34808
rect 477052 34718 487000 34778
rect 477052 34716 477058 34718
rect 486200 34688 487000 34718
rect 4110 34446 10032 34506
rect 0 34098 800 34128
rect 0 34038 6930 34098
rect 0 34008 800 34038
rect 6870 33690 6930 34038
rect 485998 34036 486004 34100
rect 486068 34098 486074 34100
rect 486200 34098 487000 34128
rect 486068 34038 487000 34098
rect 486068 34036 486074 34038
rect 486200 34008 487000 34038
rect 6870 33630 10032 33690
rect 0 33418 800 33448
rect 1342 33418 1348 33420
rect 0 33358 1348 33418
rect 0 33328 800 33358
rect 1342 33356 1348 33358
rect 1412 33356 1418 33420
rect 478270 33356 478276 33420
rect 478340 33418 478346 33420
rect 486200 33418 487000 33448
rect 478340 33358 487000 33418
rect 478340 33356 478346 33358
rect 486200 33328 487000 33358
rect 8334 32812 8340 32876
rect 8404 32874 8410 32876
rect 8404 32814 10032 32874
rect 8404 32812 8410 32814
rect 0 32738 800 32768
rect 486200 32740 487000 32768
rect 1158 32738 1164 32740
rect 0 32678 1164 32738
rect 0 32648 800 32678
rect 1158 32676 1164 32678
rect 1228 32676 1234 32740
rect 486200 32676 486372 32740
rect 486436 32676 487000 32740
rect 486200 32648 487000 32676
rect 0 32058 800 32088
rect 6177 32058 6243 32061
rect 0 32056 6243 32058
rect 0 32000 6182 32056
rect 6238 32000 6243 32056
rect 0 31998 6243 32000
rect 0 31968 800 31998
rect 6177 31995 6243 31998
rect 8518 31996 8524 32060
rect 8588 32058 8594 32060
rect 8588 31998 10032 32058
rect 8588 31996 8594 31998
rect 478086 31996 478092 32060
rect 478156 32058 478162 32060
rect 486200 32058 487000 32088
rect 478156 31998 487000 32058
rect 478156 31996 478162 31998
rect 486200 31968 487000 31998
rect 1158 31588 1164 31652
rect 1228 31650 1234 31652
rect 6126 31650 6132 31652
rect 1228 31590 6132 31650
rect 1228 31588 1234 31590
rect 6126 31588 6132 31590
rect 6196 31588 6202 31652
rect 0 31378 800 31408
rect 4797 31378 4863 31381
rect 0 31376 4863 31378
rect 0 31320 4802 31376
rect 4858 31320 4863 31376
rect 0 31318 4863 31320
rect 0 31288 800 31318
rect 4797 31315 4863 31318
rect 485630 31316 485636 31380
rect 485700 31378 485706 31380
rect 486200 31378 487000 31408
rect 485700 31318 487000 31378
rect 485700 31316 485706 31318
rect 486200 31288 487000 31318
rect 7097 31242 7163 31245
rect 7097 31240 10032 31242
rect 7097 31184 7102 31240
rect 7158 31184 10032 31240
rect 7097 31182 10032 31184
rect 7097 31179 7163 31182
rect 0 30698 800 30728
rect 1117 30698 1183 30701
rect 0 30696 1183 30698
rect 0 30640 1122 30696
rect 1178 30640 1183 30696
rect 0 30638 1183 30640
rect 0 30608 800 30638
rect 1117 30635 1183 30638
rect 483105 30698 483171 30701
rect 486200 30698 487000 30728
rect 483105 30696 487000 30698
rect 483105 30640 483110 30696
rect 483166 30640 487000 30696
rect 483105 30638 487000 30640
rect 483105 30635 483171 30638
rect 486200 30608 487000 30638
rect 9305 30426 9371 30429
rect 9305 30424 10032 30426
rect 9305 30368 9310 30424
rect 9366 30368 10032 30424
rect 9305 30366 10032 30368
rect 9305 30363 9371 30366
rect 1342 30228 1348 30292
rect 1412 30290 1418 30292
rect 3366 30290 3372 30292
rect 1412 30230 3372 30290
rect 1412 30228 1418 30230
rect 3366 30228 3372 30230
rect 3436 30228 3442 30292
rect 0 30018 800 30048
rect 486200 30021 487000 30048
rect 7557 30018 7623 30021
rect 0 30016 7623 30018
rect 0 29960 7562 30016
rect 7618 29960 7623 30016
rect 0 29958 7623 29960
rect 0 29928 800 29958
rect 7557 29955 7623 29958
rect 486141 30016 487000 30021
rect 486141 29960 486146 30016
rect 486202 29960 487000 30016
rect 486141 29955 487000 29960
rect 486200 29928 487000 29955
rect 9581 29542 9647 29545
rect 9581 29540 10060 29542
rect 9581 29484 9586 29540
rect 9642 29484 10060 29540
rect 9581 29482 10060 29484
rect 9581 29479 9647 29482
rect 0 29338 800 29368
rect 4889 29338 4955 29341
rect 0 29336 4955 29338
rect 0 29280 4894 29336
rect 4950 29280 4955 29336
rect 0 29278 4955 29280
rect 0 29248 800 29278
rect 4889 29275 4955 29278
rect 479742 29276 479748 29340
rect 479812 29338 479818 29340
rect 486200 29338 487000 29368
rect 479812 29278 487000 29338
rect 479812 29276 479818 29278
rect 486200 29248 487000 29278
rect 1117 28930 1183 28933
rect 5073 28930 5139 28933
rect 1117 28928 5139 28930
rect 1117 28872 1122 28928
rect 1178 28872 5078 28928
rect 5134 28872 5139 28928
rect 1117 28870 5139 28872
rect 1117 28867 1183 28870
rect 5073 28867 5139 28870
rect 8661 28794 8727 28797
rect 8661 28792 10032 28794
rect 8661 28736 8666 28792
rect 8722 28736 10032 28792
rect 8661 28734 10032 28736
rect 8661 28731 8727 28734
rect 0 28658 800 28688
rect 0 28598 1042 28658
rect 0 28568 800 28598
rect 197 28386 263 28389
rect 982 28386 1042 28598
rect 479374 28596 479380 28660
rect 479444 28658 479450 28660
rect 486200 28658 487000 28688
rect 479444 28598 487000 28658
rect 479444 28596 479450 28598
rect 486200 28568 487000 28598
rect 197 28384 1042 28386
rect 197 28328 202 28384
rect 258 28328 1042 28384
rect 197 28326 1042 28328
rect 197 28323 263 28326
rect 0 27978 800 28008
rect 1301 27978 1367 27981
rect 0 27976 1367 27978
rect 0 27920 1306 27976
rect 1362 27920 1367 27976
rect 0 27918 1367 27920
rect 0 27888 800 27918
rect 1301 27915 1367 27918
rect 8201 27978 8267 27981
rect 8201 27976 10032 27978
rect 8201 27920 8206 27976
rect 8262 27920 10032 27976
rect 8201 27918 10032 27920
rect 8201 27915 8267 27918
rect 479558 27916 479564 27980
rect 479628 27978 479634 27980
rect 486200 27978 487000 28008
rect 479628 27918 487000 27978
rect 479628 27916 479634 27918
rect 486200 27888 487000 27918
rect 0 27298 800 27328
rect 7649 27298 7715 27301
rect 0 27296 7715 27298
rect 0 27240 7654 27296
rect 7710 27240 7715 27296
rect 0 27238 7715 27240
rect 0 27208 800 27238
rect 7649 27235 7715 27238
rect 480069 27298 480135 27301
rect 486200 27298 487000 27328
rect 480069 27296 487000 27298
rect 480069 27240 480074 27296
rect 480130 27240 487000 27296
rect 480069 27238 487000 27240
rect 480069 27235 480135 27238
rect 486200 27208 487000 27238
rect 8017 27162 8083 27165
rect 8017 27160 10032 27162
rect 8017 27104 8022 27160
rect 8078 27104 10032 27160
rect 8017 27102 10032 27104
rect 8017 27099 8083 27102
rect 0 26618 800 26648
rect 1209 26618 1275 26621
rect 0 26616 1275 26618
rect 0 26560 1214 26616
rect 1270 26560 1275 26616
rect 0 26558 1275 26560
rect 0 26528 800 26558
rect 1209 26555 1275 26558
rect 480161 26618 480227 26621
rect 486200 26618 487000 26648
rect 480161 26616 487000 26618
rect 480161 26560 480166 26616
rect 480222 26560 487000 26616
rect 480161 26558 487000 26560
rect 480161 26555 480227 26558
rect 486200 26528 487000 26558
rect 9397 26346 9463 26349
rect 9397 26344 10032 26346
rect 9397 26288 9402 26344
rect 9458 26288 10032 26344
rect 9397 26286 10032 26288
rect 9397 26283 9463 26286
rect 0 25938 800 25968
rect 1342 25938 1348 25940
rect 0 25878 1348 25938
rect 0 25848 800 25878
rect 1342 25876 1348 25878
rect 1412 25876 1418 25940
rect 484894 25876 484900 25940
rect 484964 25938 484970 25940
rect 486200 25938 487000 25968
rect 484964 25878 487000 25938
rect 484964 25876 484970 25878
rect 486200 25848 487000 25878
rect 9438 25468 9444 25532
rect 9508 25530 9514 25532
rect 9508 25470 10032 25530
rect 9508 25468 9514 25470
rect 0 25258 800 25288
rect 8937 25258 9003 25261
rect 0 25256 9003 25258
rect 0 25200 8942 25256
rect 8998 25200 9003 25256
rect 0 25198 9003 25200
rect 0 25168 800 25198
rect 8937 25195 9003 25198
rect 481398 25196 481404 25260
rect 481468 25258 481474 25260
rect 486200 25258 487000 25288
rect 481468 25198 487000 25258
rect 481468 25196 481474 25198
rect 486200 25168 487000 25198
rect 9029 24714 9095 24717
rect 9029 24712 10032 24714
rect 9029 24656 9034 24712
rect 9090 24656 10032 24712
rect 9029 24654 10032 24656
rect 9029 24651 9095 24654
rect 0 24578 800 24608
rect 4102 24578 4108 24580
rect 0 24518 4108 24578
rect 0 24488 800 24518
rect 4102 24516 4108 24518
rect 4172 24516 4178 24580
rect 482318 24516 482324 24580
rect 482388 24578 482394 24580
rect 486200 24578 487000 24608
rect 482388 24518 487000 24578
rect 482388 24516 482394 24518
rect 486200 24488 487000 24518
rect 0 23898 800 23928
rect 3417 23898 3483 23901
rect 0 23896 3483 23898
rect 0 23840 3422 23896
rect 3478 23840 3483 23896
rect 0 23838 3483 23840
rect 0 23808 800 23838
rect 3417 23835 3483 23838
rect 7741 23898 7807 23901
rect 7741 23896 10032 23898
rect 7741 23840 7746 23896
rect 7802 23840 10032 23896
rect 7741 23838 10032 23840
rect 7741 23835 7807 23838
rect 481214 23836 481220 23900
rect 481284 23898 481290 23900
rect 486200 23898 487000 23928
rect 481284 23838 487000 23898
rect 481284 23836 481290 23838
rect 486200 23808 487000 23838
rect 1301 23762 1367 23765
rect 7373 23762 7439 23765
rect 1301 23760 7439 23762
rect 1301 23704 1306 23760
rect 1362 23704 7378 23760
rect 7434 23704 7439 23760
rect 1301 23702 7439 23704
rect 1301 23699 1367 23702
rect 7373 23699 7439 23702
rect 0 23218 800 23248
rect 5533 23218 5599 23221
rect 0 23216 5599 23218
rect 0 23160 5538 23216
rect 5594 23160 5599 23216
rect 0 23158 5599 23160
rect 0 23128 800 23158
rect 5533 23155 5599 23158
rect 483790 23156 483796 23220
rect 483860 23218 483866 23220
rect 486200 23218 487000 23248
rect 483860 23158 487000 23218
rect 483860 23156 483866 23158
rect 486200 23128 487000 23158
rect 6453 23082 6519 23085
rect 6453 23080 10032 23082
rect 6453 23024 6458 23080
rect 6514 23024 10032 23080
rect 6453 23022 10032 23024
rect 6453 23019 6519 23022
rect 0 22538 800 22568
rect 9622 22538 9628 22540
rect 0 22478 9628 22538
rect 0 22448 800 22478
rect 9622 22476 9628 22478
rect 9692 22476 9698 22540
rect 482134 22476 482140 22540
rect 482204 22538 482210 22540
rect 486200 22538 487000 22568
rect 482204 22478 487000 22538
rect 482204 22476 482210 22478
rect 486200 22448 487000 22478
rect 4102 22204 4108 22268
rect 4172 22266 4178 22268
rect 4172 22206 10032 22266
rect 4172 22204 4178 22206
rect 1209 21994 1275 21997
rect 8845 21994 8911 21997
rect 1209 21992 8911 21994
rect 1209 21936 1214 21992
rect 1270 21936 8850 21992
rect 8906 21936 8911 21992
rect 1209 21934 8911 21936
rect 1209 21931 1275 21934
rect 8845 21931 8911 21934
rect 0 21858 800 21888
rect 0 21798 6930 21858
rect 0 21768 800 21798
rect 6870 21450 6930 21798
rect 481030 21796 481036 21860
rect 481100 21858 481106 21860
rect 486200 21858 487000 21888
rect 481100 21798 487000 21858
rect 481100 21796 481106 21798
rect 486200 21768 487000 21798
rect 6870 21390 10032 21450
rect 0 21178 800 21208
rect 8150 21178 8156 21180
rect 0 21118 8156 21178
rect 0 21088 800 21118
rect 8150 21116 8156 21118
rect 8220 21116 8226 21180
rect 482829 21178 482895 21181
rect 486200 21178 487000 21208
rect 482829 21176 487000 21178
rect 482829 21120 482834 21176
rect 482890 21120 487000 21176
rect 482829 21118 487000 21120
rect 482829 21115 482895 21118
rect 486200 21088 487000 21118
rect 0 20498 800 20528
rect 9121 20498 9187 20501
rect 0 20496 9187 20498
rect 0 20440 9126 20496
rect 9182 20440 9187 20496
rect 0 20438 9187 20440
rect 0 20408 800 20438
rect 9121 20435 9187 20438
rect 483606 20436 483612 20500
rect 483676 20498 483682 20500
rect 486200 20498 487000 20528
rect 483676 20438 487000 20498
rect 483676 20436 483682 20438
rect 486200 20408 487000 20438
rect 0 19818 800 19848
rect 9489 19818 9555 19821
rect 0 19816 9555 19818
rect 0 19760 9494 19816
rect 9550 19760 9555 19816
rect 0 19758 9555 19760
rect 0 19728 800 19758
rect 9489 19755 9555 19758
rect 482921 19818 482987 19821
rect 486200 19818 487000 19848
rect 482921 19816 487000 19818
rect 482921 19760 482926 19816
rect 482982 19760 487000 19816
rect 482921 19758 487000 19760
rect 482921 19755 482987 19758
rect 486200 19728 487000 19758
rect 0 19138 800 19168
rect 9806 19138 9812 19140
rect 0 19078 9812 19138
rect 0 19048 800 19078
rect 9806 19076 9812 19078
rect 9876 19076 9882 19140
rect 484209 19138 484275 19141
rect 486200 19138 487000 19168
rect 484209 19136 487000 19138
rect 484209 19080 484214 19136
rect 484270 19080 487000 19136
rect 484209 19078 487000 19080
rect 484209 19075 484275 19078
rect 486200 19048 487000 19078
rect 0 18458 800 18488
rect 6678 18458 6684 18460
rect 0 18398 6684 18458
rect 0 18368 800 18398
rect 6678 18396 6684 18398
rect 6748 18396 6754 18460
rect 481541 18458 481607 18461
rect 486200 18458 487000 18488
rect 481541 18456 487000 18458
rect 481541 18400 481546 18456
rect 481602 18400 487000 18456
rect 481541 18398 487000 18400
rect 481541 18395 481607 18398
rect 486200 18368 487000 18398
rect 1342 18124 1348 18188
rect 1412 18186 1418 18188
rect 11094 18186 11100 18188
rect 1412 18126 11100 18186
rect 1412 18124 1418 18126
rect 11094 18124 11100 18126
rect 11164 18124 11170 18188
rect 197 18050 263 18053
rect 8477 18050 8543 18053
rect 197 18048 8543 18050
rect 197 17992 202 18048
rect 258 17992 8482 18048
rect 8538 17992 8543 18048
rect 197 17990 8543 17992
rect 197 17987 263 17990
rect 8477 17987 8543 17990
rect 5073 17914 5139 17917
rect 9213 17914 9279 17917
rect 5073 17912 9279 17914
rect 5073 17856 5078 17912
rect 5134 17856 9218 17912
rect 9274 17856 9279 17912
rect 5073 17854 9279 17856
rect 5073 17851 5139 17854
rect 9213 17851 9279 17854
rect 0 17778 800 17808
rect 484301 17778 484367 17781
rect 486200 17778 487000 17808
rect 0 17718 6930 17778
rect 0 17688 800 17718
rect 0 17098 800 17128
rect 4838 17098 4844 17100
rect 0 17038 4844 17098
rect 0 17008 800 17038
rect 4838 17036 4844 17038
rect 4908 17036 4914 17100
rect 6870 17098 6930 17718
rect 484301 17776 487000 17778
rect 484301 17720 484306 17776
rect 484362 17720 487000 17776
rect 484301 17718 487000 17720
rect 484301 17715 484367 17718
rect 486200 17688 487000 17718
rect 9622 17580 9628 17644
rect 9692 17642 9698 17644
rect 9692 17582 18154 17642
rect 9692 17580 9698 17582
rect 9121 17506 9187 17509
rect 12566 17506 12572 17508
rect 9121 17504 12572 17506
rect 9121 17448 9126 17504
rect 9182 17448 12572 17504
rect 9121 17446 12572 17448
rect 9121 17443 9187 17446
rect 12566 17444 12572 17446
rect 12636 17444 12642 17508
rect 8150 17308 8156 17372
rect 8220 17370 8226 17372
rect 8220 17310 16590 17370
rect 8220 17308 8226 17310
rect 11094 17172 11100 17236
rect 11164 17234 11170 17236
rect 11164 17174 13738 17234
rect 11164 17172 11170 17174
rect 13678 17101 13738 17174
rect 13215 17098 13281 17101
rect 6870 17096 13281 17098
rect 6870 17040 13220 17096
rect 13276 17040 13281 17096
rect 6870 17038 13281 17040
rect 13215 17035 13281 17038
rect 13675 17096 13741 17101
rect 13675 17040 13680 17096
rect 13736 17040 13741 17096
rect 13675 17035 13741 17040
rect 16530 17098 16590 17310
rect 17815 17098 17881 17101
rect 16530 17096 17881 17098
rect 16530 17040 17820 17096
rect 17876 17040 17881 17096
rect 16530 17038 17881 17040
rect 18094 17098 18154 17582
rect 18735 17098 18801 17101
rect 18094 17096 18801 17098
rect 18094 17040 18740 17096
rect 18796 17040 18801 17096
rect 18094 17038 18801 17040
rect 17815 17035 17881 17038
rect 18735 17035 18801 17038
rect 480846 17036 480852 17100
rect 480916 17098 480922 17100
rect 486200 17098 487000 17128
rect 480916 17038 487000 17098
rect 480916 17036 480922 17038
rect 486200 17008 487000 17038
rect 9489 16962 9555 16965
rect 12341 16962 12407 16965
rect 9489 16960 12407 16962
rect 9489 16904 9494 16960
rect 9550 16904 12346 16960
rect 12402 16904 12407 16960
rect 9489 16902 12407 16904
rect 9489 16899 9555 16902
rect 12341 16899 12407 16902
rect 12566 16900 12572 16964
rect 12636 16962 12642 16964
rect 17401 16962 17467 16965
rect 12636 16960 17467 16962
rect 12636 16904 17406 16960
rect 17462 16904 17467 16960
rect 12636 16902 17467 16904
rect 12636 16900 12642 16902
rect 17401 16899 17467 16902
rect 4889 16826 4955 16829
rect 11881 16826 11947 16829
rect 4889 16824 11947 16826
rect 4889 16768 4894 16824
rect 4950 16768 11886 16824
rect 11942 16768 11947 16824
rect 4889 16766 11947 16768
rect 4889 16763 4955 16766
rect 11881 16763 11947 16766
rect 5533 16690 5599 16693
rect 14181 16690 14247 16693
rect 5533 16688 14247 16690
rect 5533 16632 5538 16688
rect 5594 16632 14186 16688
rect 14242 16632 14247 16688
rect 5533 16630 14247 16632
rect 5533 16627 5599 16630
rect 14181 16627 14247 16630
rect 4797 16554 4863 16557
rect 8109 16554 8175 16557
rect 4797 16552 8175 16554
rect 4797 16496 4802 16552
rect 4858 16496 8114 16552
rect 8170 16496 8175 16552
rect 4797 16494 8175 16496
rect 4797 16491 4863 16494
rect 8109 16491 8175 16494
rect 9806 16492 9812 16556
rect 9876 16554 9882 16556
rect 16941 16554 17007 16557
rect 9876 16552 17007 16554
rect 9876 16496 16946 16552
rect 17002 16496 17007 16552
rect 9876 16494 17007 16496
rect 9876 16492 9882 16494
rect 16941 16491 17007 16494
rect 0 16418 800 16448
rect 0 16358 20730 16418
rect 0 16328 800 16358
rect 8937 16282 9003 16285
rect 16021 16282 16087 16285
rect 8937 16280 16087 16282
rect 8937 16224 8942 16280
rect 8998 16224 16026 16280
rect 16082 16224 16087 16280
rect 8937 16222 16087 16224
rect 8937 16219 9003 16222
rect 16021 16219 16087 16222
rect 3417 16146 3483 16149
rect 15561 16146 15627 16149
rect 3417 16144 15627 16146
rect 3417 16088 3422 16144
rect 3478 16088 15566 16144
rect 15622 16088 15627 16144
rect 3417 16086 15627 16088
rect 3417 16083 3483 16086
rect 15561 16083 15627 16086
rect 6862 15948 6868 16012
rect 6932 16010 6938 16012
rect 12801 16010 12867 16013
rect 6932 16008 12867 16010
rect 6932 15952 12806 16008
rect 12862 15952 12867 16008
rect 6932 15950 12867 15952
rect 6932 15948 6938 15950
rect 12801 15947 12867 15950
rect 20670 15942 20730 16358
rect 20670 15882 21310 15942
rect 0 15738 800 15768
rect 0 15678 20730 15738
rect 0 15648 800 15678
rect 20670 15670 20730 15678
rect 20670 15610 21310 15670
rect 4838 15268 4844 15332
rect 4908 15330 4914 15332
rect 4908 15270 21282 15330
rect 4908 15268 4914 15270
rect 6126 15132 6132 15196
rect 6196 15194 6202 15196
rect 6196 15134 16590 15194
rect 6196 15132 6202 15134
rect 0 15058 800 15088
rect 16530 15058 16590 15134
rect 0 14998 6930 15058
rect 16530 14998 21282 15058
rect 0 14968 800 14998
rect 6870 14922 6930 14998
rect 6870 14862 20730 14922
rect 20670 14854 20730 14862
rect 20670 14794 21310 14854
rect 3366 14452 3372 14516
rect 3436 14514 3442 14516
rect 3436 14454 21282 14514
rect 3436 14452 3442 14454
rect 0 14378 800 14408
rect 0 14318 20730 14378
rect 0 14288 800 14318
rect 20670 14310 20730 14318
rect 20670 14250 21310 14310
rect 20670 13898 21310 13958
rect 20670 13834 20730 13898
rect 13862 13774 20730 13834
rect 0 13698 800 13728
rect 13862 13698 13922 13774
rect 0 13638 13922 13698
rect 18873 13698 18939 13701
rect 18873 13696 21282 13698
rect 18873 13640 18878 13696
rect 18934 13640 21282 13696
rect 18873 13638 21282 13640
rect 0 13608 800 13638
rect 18873 13635 18939 13638
rect 790 13364 796 13428
rect 860 13426 866 13428
rect 860 13366 21282 13426
rect 860 13364 866 13366
rect 54 13228 60 13292
rect 124 13290 130 13292
rect 124 13230 20730 13290
rect 124 13228 130 13230
rect 20670 13222 20730 13230
rect 20670 13162 21310 13222
rect 0 13018 800 13048
rect 18873 13018 18939 13021
rect 0 13016 18939 13018
rect 0 12960 18878 13016
rect 18934 12960 18939 13016
rect 0 12958 18939 12960
rect 0 12928 800 12958
rect 18873 12955 18939 12958
rect 18822 12820 18828 12884
rect 18892 12882 18898 12884
rect 18892 12822 21282 12882
rect 18892 12820 18898 12822
rect 19558 12548 19564 12612
rect 19628 12610 19634 12612
rect 19628 12550 21282 12610
rect 19628 12548 19634 12550
rect 0 12338 800 12368
rect 11513 12338 11579 12341
rect 0 12336 11579 12338
rect 0 12280 11518 12336
rect 11574 12280 11579 12336
rect 0 12278 11579 12280
rect 0 12248 800 12278
rect 11513 12275 11579 12278
rect 11654 12278 21282 12338
rect 3366 12140 3372 12204
rect 3436 12202 3442 12204
rect 11654 12202 11714 12278
rect 3436 12142 11714 12202
rect 11789 12202 11855 12205
rect 18822 12202 18828 12204
rect 11789 12200 18828 12202
rect 11789 12144 11794 12200
rect 11850 12144 18828 12200
rect 11789 12142 18828 12144
rect 3436 12140 3442 12142
rect 11789 12139 11855 12142
rect 18822 12140 18828 12142
rect 18892 12140 18898 12204
rect 6870 12006 21282 12066
rect 0 11658 800 11688
rect 6870 11658 6930 12006
rect 15326 11732 15332 11796
rect 15396 11794 15402 11796
rect 15396 11734 21282 11794
rect 15396 11732 15402 11734
rect 0 11598 6930 11658
rect 0 11568 800 11598
rect 18822 11460 18828 11524
rect 18892 11522 18898 11524
rect 18892 11462 21282 11522
rect 18892 11460 18898 11462
rect 18454 11188 18460 11252
rect 18524 11250 18530 11252
rect 18524 11190 21282 11250
rect 18524 11188 18530 11190
rect 0 10978 800 11008
rect 0 10918 6930 10978
rect 0 10888 800 10918
rect 6870 10842 6930 10918
rect 17166 10916 17172 10980
rect 17236 10978 17242 10980
rect 17236 10918 21282 10978
rect 17236 10916 17242 10918
rect 18822 10842 18828 10844
rect 6870 10782 18828 10842
rect 18822 10780 18828 10782
rect 18892 10780 18898 10844
rect 17350 10644 17356 10708
rect 17420 10706 17426 10708
rect 17420 10646 21282 10706
rect 17420 10644 17426 10646
rect 6870 10374 21282 10434
rect 0 10298 800 10328
rect 6870 10298 6930 10374
rect 0 10238 6930 10298
rect 0 10208 800 10238
rect 20110 10100 20116 10164
rect 20180 10162 20186 10164
rect 20180 10102 21282 10162
rect 20180 10100 20186 10102
rect 19926 9828 19932 9892
rect 19996 9890 20002 9892
rect 19996 9830 21282 9890
rect 19996 9828 20002 9830
rect 0 9618 800 9648
rect 0 9558 21282 9618
rect 0 9528 800 9558
rect 18638 9284 18644 9348
rect 18708 9346 18714 9348
rect 18708 9286 21282 9346
rect 18708 9284 18714 9286
rect 20345 9074 20411 9077
rect 20345 9072 21282 9074
rect 20345 9016 20350 9072
rect 20406 9016 21282 9072
rect 20345 9014 21282 9016
rect 20345 9011 20411 9014
rect 0 8938 800 8968
rect 19558 8938 19564 8940
rect 0 8878 19564 8938
rect 0 8848 800 8878
rect 19558 8876 19564 8878
rect 19628 8876 19634 8940
rect 15142 8740 15148 8804
rect 15212 8802 15218 8804
rect 15212 8742 21282 8802
rect 15212 8740 15218 8742
rect 14406 8468 14412 8532
rect 14476 8530 14482 8532
rect 14476 8470 21282 8530
rect 14476 8468 14482 8470
rect 0 8258 800 8288
rect 10961 8258 11027 8261
rect 14181 8258 14247 8261
rect 0 8198 6930 8258
rect 0 8168 800 8198
rect 6870 8122 6930 8198
rect 10961 8256 14247 8258
rect 10961 8200 10966 8256
rect 11022 8200 14186 8256
rect 14242 8200 14247 8256
rect 10961 8198 14247 8200
rect 10961 8195 11027 8198
rect 14181 8195 14247 8198
rect 21081 8258 21147 8261
rect 21081 8256 21282 8258
rect 21081 8200 21086 8256
rect 21142 8200 21282 8256
rect 21081 8198 21282 8200
rect 21081 8195 21147 8198
rect 15326 8122 15332 8124
rect 6870 8062 15332 8122
rect 15326 8060 15332 8062
rect 15396 8060 15402 8124
rect 20345 7988 20411 7989
rect 20294 7986 20300 7988
rect 20254 7926 20300 7986
rect 20364 7984 20411 7988
rect 20406 7928 20411 7984
rect 20294 7924 20300 7926
rect 20364 7924 20411 7928
rect 20345 7923 20411 7924
rect 20529 7986 20595 7989
rect 20529 7984 21282 7986
rect 20529 7928 20534 7984
rect 20590 7928 21282 7984
rect 20529 7926 21282 7928
rect 20529 7923 20595 7926
rect 21081 7714 21147 7717
rect 21081 7712 21282 7714
rect 21081 7656 21086 7712
rect 21142 7656 21282 7712
rect 21081 7654 21282 7656
rect 21081 7651 21147 7654
rect 0 7578 800 7608
rect 15142 7578 15148 7580
rect 0 7518 15148 7578
rect 0 7488 800 7518
rect 15142 7516 15148 7518
rect 15212 7516 15218 7580
rect 20621 7442 20687 7445
rect 20621 7440 21282 7442
rect 20621 7384 20626 7440
rect 20682 7384 21282 7440
rect 20621 7382 21282 7384
rect 20621 7379 20687 7382
rect 0 6898 800 6928
rect 17166 6898 17172 6900
rect 0 6838 17172 6898
rect 0 6808 800 6838
rect 17166 6836 17172 6838
rect 17236 6836 17242 6900
rect 0 6218 800 6248
rect 17350 6218 17356 6220
rect 0 6158 17356 6218
rect 0 6128 800 6158
rect 17350 6156 17356 6158
rect 17420 6156 17426 6220
rect 14181 5946 14247 5949
rect 29177 5946 29243 5949
rect 72371 5946 72437 5949
rect 104643 5946 104709 5949
rect 177103 5946 177169 5949
rect 218099 5946 218165 5949
rect 259131 5946 259197 5949
rect 276551 5946 276617 5949
rect 345105 5946 345171 5949
rect 378915 5946 378981 5949
rect 414407 5946 414473 5949
rect 444459 5946 444525 5949
rect 14181 5944 444525 5946
rect 14181 5888 14186 5944
rect 14242 5888 29182 5944
rect 29238 5888 72376 5944
rect 72432 5888 104648 5944
rect 104704 5888 177108 5944
rect 177164 5888 218104 5944
rect 218160 5888 259136 5944
rect 259192 5888 276556 5944
rect 276612 5888 345110 5944
rect 345166 5888 378920 5944
rect 378976 5888 414412 5944
rect 414468 5888 444464 5944
rect 444520 5888 444525 5944
rect 14181 5886 444525 5888
rect 14181 5883 14247 5886
rect 29177 5883 29243 5886
rect 72371 5883 72437 5886
rect 104643 5883 104709 5886
rect 177103 5883 177169 5886
rect 218099 5883 218165 5886
rect 259131 5883 259197 5886
rect 276551 5883 276617 5886
rect 345105 5883 345171 5886
rect 378915 5883 378981 5886
rect 414407 5883 414473 5886
rect 444459 5883 444525 5886
rect 383343 5810 383409 5813
rect 392853 5810 392919 5813
rect 383343 5808 392919 5810
rect 383343 5752 383348 5808
rect 383404 5752 392858 5808
rect 392914 5752 392919 5808
rect 383343 5750 392919 5752
rect 383343 5747 383409 5750
rect 392853 5747 392919 5750
rect 9438 5612 9444 5676
rect 9508 5674 9514 5676
rect 11605 5674 11671 5677
rect 9508 5672 11671 5674
rect 9508 5616 11610 5672
rect 11666 5616 11671 5672
rect 9508 5614 11671 5616
rect 9508 5612 9514 5614
rect 11605 5611 11671 5614
rect 0 5538 800 5568
rect 20110 5538 20116 5540
rect 0 5478 20116 5538
rect 0 5448 800 5478
rect 20110 5476 20116 5478
rect 20180 5476 20186 5540
rect 0 4858 800 4888
rect 14406 4858 14412 4860
rect 0 4798 14412 4858
rect 0 4768 800 4798
rect 14406 4796 14412 4798
rect 14476 4796 14482 4860
rect 54 4388 60 4452
rect 124 4450 130 4452
rect 124 4390 1042 4450
rect 124 4388 130 4390
rect 0 4178 800 4208
rect 982 4178 1042 4390
rect 0 4118 1042 4178
rect 9305 4178 9371 4181
rect 12893 4178 12959 4181
rect 9305 4176 12959 4178
rect 9305 4120 9310 4176
rect 9366 4120 12898 4176
rect 12954 4120 12959 4176
rect 9305 4118 12959 4120
rect 0 4088 800 4118
rect 9305 4115 9371 4118
rect 12893 4115 12959 4118
rect 20621 3634 20687 3637
rect 22553 3634 22619 3637
rect 20621 3632 22619 3634
rect 20621 3576 20626 3632
rect 20682 3576 22558 3632
rect 22614 3576 22619 3632
rect 20621 3574 22619 3576
rect 20621 3571 20687 3574
rect 22553 3571 22619 3574
rect 0 3498 800 3528
rect 19926 3498 19932 3500
rect 0 3438 19932 3498
rect 0 3408 800 3438
rect 19926 3436 19932 3438
rect 19996 3436 20002 3500
rect 238 3028 244 3092
rect 308 3090 314 3092
rect 308 3030 1042 3090
rect 308 3028 314 3030
rect 0 2818 800 2848
rect 982 2818 1042 3030
rect 1158 2892 1164 2956
rect 1228 2954 1234 2956
rect 3366 2954 3372 2956
rect 1228 2894 3372 2954
rect 1228 2892 1234 2894
rect 3366 2892 3372 2894
rect 3436 2892 3442 2956
rect 0 2758 1042 2818
rect 0 2728 800 2758
rect 1342 2348 1348 2412
rect 1412 2410 1418 2412
rect 18638 2410 18644 2412
rect 1412 2350 18644 2410
rect 1412 2348 1418 2350
rect 18638 2348 18644 2350
rect 18708 2348 18714 2412
rect 0 2138 800 2168
rect 18454 2138 18460 2140
rect 0 2078 18460 2138
rect 0 2048 800 2078
rect 18454 2076 18460 2078
rect 18524 2076 18530 2140
rect 0 1458 800 1488
rect 1158 1458 1164 1460
rect 0 1398 1164 1458
rect 0 1368 800 1398
rect 1158 1396 1164 1398
rect 1228 1396 1234 1460
rect 8385 1322 8451 1325
rect 8518 1322 8524 1324
rect 8385 1320 8524 1322
rect 8385 1264 8390 1320
rect 8446 1264 8524 1320
rect 8385 1262 8524 1264
rect 8385 1259 8451 1262
rect 8518 1260 8524 1262
rect 8588 1260 8594 1324
rect 9397 1322 9463 1325
rect 10317 1322 10383 1325
rect 9397 1320 10383 1322
rect 9397 1264 9402 1320
rect 9458 1264 10322 1320
rect 10378 1264 10383 1320
rect 9397 1262 10383 1264
rect 9397 1259 9463 1262
rect 10317 1259 10383 1262
rect 385585 1322 385651 1325
rect 386413 1322 386479 1325
rect 385585 1320 386479 1322
rect 385585 1264 385590 1320
rect 385646 1264 386418 1320
rect 386474 1264 386479 1320
rect 385585 1262 386479 1264
rect 385585 1259 385651 1262
rect 386413 1259 386479 1262
rect 388897 1322 388963 1325
rect 389633 1322 389699 1325
rect 388897 1320 389699 1322
rect 388897 1264 388902 1320
rect 388958 1264 389638 1320
rect 389694 1264 389699 1320
rect 388897 1262 389699 1264
rect 388897 1259 388963 1262
rect 389633 1259 389699 1262
rect 8661 1186 8727 1189
rect 10961 1186 11027 1189
rect 8661 1184 11027 1186
rect 8661 1128 8666 1184
rect 8722 1128 10966 1184
rect 11022 1128 11027 1184
rect 8661 1126 11027 1128
rect 8661 1123 8727 1126
rect 10961 1123 11027 1126
rect 384481 1186 384547 1189
rect 387701 1186 387767 1189
rect 384481 1184 387767 1186
rect 384481 1128 384486 1184
rect 384542 1128 387706 1184
rect 387762 1128 387767 1184
rect 384481 1126 387767 1128
rect 384481 1123 384547 1126
rect 387701 1123 387767 1126
rect 8017 1050 8083 1053
rect 12249 1050 12315 1053
rect 8017 1048 12315 1050
rect 8017 992 8022 1048
rect 8078 992 12254 1048
rect 12310 992 12315 1048
rect 8017 990 12315 992
rect 8017 987 8083 990
rect 12249 987 12315 990
rect 386689 1050 386755 1053
rect 390921 1050 390987 1053
rect 386689 1048 390987 1050
rect 386689 992 386694 1048
rect 386750 992 390926 1048
rect 390982 992 390987 1048
rect 386689 990 390987 992
rect 386689 987 386755 990
rect 390921 987 390987 990
rect 8109 914 8175 917
rect 13537 914 13603 917
rect 8109 912 13603 914
rect 8109 856 8114 912
rect 8170 856 13542 912
rect 13598 856 13603 912
rect 8109 854 13603 856
rect 8109 851 8175 854
rect 13537 851 13603 854
rect 0 778 800 808
rect 1342 778 1348 780
rect 0 718 1348 778
rect 0 688 800 718
rect 1342 716 1348 718
rect 1412 716 1418 780
rect 382273 506 382339 509
rect 388253 506 388319 509
rect 382273 504 388319 506
rect 382273 448 382278 504
rect 382334 448 388258 504
rect 388314 448 388319 504
rect 382273 446 388319 448
rect 382273 443 382339 446
rect 388253 443 388319 446
rect 380065 370 380131 373
rect 394049 370 394115 373
rect 380065 368 394115 370
rect 380065 312 380070 368
rect 380126 312 394054 368
rect 394110 312 394115 368
rect 380065 310 394115 312
rect 380065 307 380131 310
rect 394049 307 394115 310
rect 20294 234 20300 236
rect 6870 174 20300 234
rect 0 98 800 128
rect 6870 98 6930 174
rect 20294 172 20300 174
rect 20364 172 20370 236
rect 381169 234 381235 237
rect 386965 234 387031 237
rect 381169 232 387031 234
rect 381169 176 381174 232
rect 381230 176 386970 232
rect 387026 176 387031 232
rect 381169 174 387031 176
rect 381169 171 381235 174
rect 386965 171 387031 174
rect 0 38 6930 98
rect 0 8 800 38
<< via3 >>
rect 21220 755788 21284 755852
rect 19932 754972 19996 755036
rect 20668 749396 20732 749460
rect 20484 748580 20548 748644
rect 21278 746834 21342 746898
rect 19932 743276 19996 743340
rect 20668 741394 20732 741458
rect 20484 740012 20548 740076
rect 480116 737156 480180 737220
rect 482876 735116 482940 735180
rect 483612 725596 483676 725660
rect 483980 722876 484044 722940
rect 484900 720836 484964 720900
rect 483796 719476 483860 719540
rect 479380 716076 479444 716140
rect 480852 715396 480916 715460
rect 481036 714716 481100 714780
rect 486372 712676 486436 712740
rect 478092 711316 478156 711380
rect 484164 710636 484228 710700
rect 477172 709956 477236 710020
rect 478276 709276 478340 709340
rect 486004 708596 486068 708660
rect 485820 707916 485884 707980
rect 478460 707236 478524 707300
rect 485084 706556 485148 706620
rect 485268 705876 485332 705940
rect 481404 705196 481468 705260
rect 485636 704516 485700 704580
rect 482876 703700 482940 703764
rect 485452 703156 485516 703220
rect 479748 702476 479812 702540
rect 486372 701116 486436 701180
rect 479932 700436 479996 700500
rect 478644 699348 478708 699412
rect 484900 699348 484964 699412
rect 482876 699076 482940 699140
rect 482324 698396 482388 698460
rect 480116 698260 480180 698324
rect 478644 698124 478708 698188
rect 485268 697852 485332 697916
rect 483612 697308 483676 697372
rect 483980 697172 484044 697236
rect 483428 697036 483492 697100
rect 477540 696900 477604 696964
rect 483612 696900 483676 696964
rect 483796 696764 483860 696828
rect 485820 696492 485884 696556
rect 481588 696356 481652 696420
rect 482876 696220 482940 696284
rect 485268 695676 485332 695740
rect 478828 695540 478892 695604
rect 485452 695132 485516 695196
rect 478276 694860 478340 694924
rect 485636 694452 485700 694516
rect 477724 694180 477788 694244
rect 483980 694044 484044 694108
rect 486004 693772 486068 693836
rect 480484 693500 480548 693564
rect 481036 693500 481100 693564
rect 480852 693364 480916 693428
rect 476930 693228 476994 693292
rect 480852 693092 480916 693156
rect 482140 692956 482204 693020
rect 481220 692684 481284 692748
rect 477172 692276 477236 692340
rect 478644 692276 478708 692340
rect 486004 692140 486068 692204
rect 478092 691868 478156 691932
rect 481588 691596 481652 691660
rect 485820 691596 485884 691660
rect 477908 691324 477972 691388
rect 478644 691052 478708 691116
rect 484348 690916 484412 690980
rect 483980 690780 484044 690844
rect 483612 690508 483676 690572
rect 483612 690236 483676 690300
rect 480300 689964 480364 690028
rect 483060 689964 483124 690028
rect 484164 689692 484228 689756
rect 481220 689012 481284 689076
rect 481036 688196 481100 688260
rect 485268 688060 485332 688124
rect 480484 687516 480548 687580
rect 481220 687108 481284 687172
rect 485636 687108 485700 687172
rect 480852 686972 480916 687036
rect 485452 686836 485516 686900
rect 482324 686700 482388 686764
rect 479380 686428 479444 686492
rect 483244 686156 483308 686220
rect 479564 685748 479628 685812
rect 481588 685748 481652 685812
rect 478828 685612 478892 685676
rect 480116 685476 480180 685540
rect 479748 685340 479812 685404
rect 479380 684796 479444 684860
rect 483244 684660 483308 684724
rect 483244 684524 483308 684588
rect 483612 684524 483676 684588
rect 478276 684388 478340 684452
rect 483612 684388 483676 684452
rect 479748 684116 479812 684180
rect 479932 683980 479996 684044
rect 479564 683708 479628 683772
rect 477540 683436 477604 683500
rect 484716 683436 484780 683500
rect 484348 683164 484412 683228
rect 477724 682892 477788 682956
rect 484532 682756 484596 682820
rect 481404 682620 481468 682684
rect 484348 682076 484412 682140
rect 484716 681940 484780 682004
rect 478092 681804 478156 681868
rect 485636 681396 485700 681460
rect 484348 681260 484412 681324
rect 480300 681124 480364 681188
rect 482140 680852 482204 680916
rect 481404 680716 481468 680780
rect 480116 680444 480180 680508
rect 479196 680308 479260 680372
rect 482140 680308 482204 680372
rect 486372 680036 486436 680100
rect 478276 679900 478340 679964
rect 477724 679628 477788 679692
rect 485084 679628 485148 679692
rect 485820 679492 485884 679556
rect 478460 679084 478524 679148
rect 483060 679084 483124 679148
rect 483796 679084 483860 679148
rect 481956 678948 482020 679012
rect 477908 678812 477972 678876
rect 478460 678404 478524 678468
rect 483060 678404 483124 678468
rect 483428 678404 483492 678468
rect 481772 678132 481836 678196
rect 478092 677996 478156 678060
rect 481404 677724 481468 677788
rect 479012 677452 479076 677516
rect 481036 677180 481100 677244
rect 485452 676772 485516 676836
rect 483060 676500 483124 676564
rect 483060 676228 483124 676292
rect 480668 676092 480732 676156
rect 483612 676092 483676 676156
rect 479380 675820 479444 675884
rect 479564 675820 479628 675884
rect 482140 675548 482204 675612
rect 483796 675412 483860 675476
rect 479748 674732 479812 674796
rect 483796 674732 483860 674796
rect 484532 674596 484596 674660
rect 486372 674324 486436 674388
rect 483060 674052 483124 674116
rect 478460 673644 478524 673708
rect 479196 673372 479260 673436
rect 480668 673100 480732 673164
rect 481956 672828 482020 672892
rect 480852 672556 480916 672620
rect 485636 672420 485700 672484
rect 483612 672012 483676 672076
rect 483244 671604 483308 671668
rect 477724 670924 477788 670988
rect 476908 670448 476972 670512
rect 481588 670108 481652 670172
rect 479564 669836 479628 669900
rect 479012 669564 479076 669628
rect 481772 669292 481836 669356
rect 483796 669156 483860 669220
rect 483428 668884 483492 668948
rect 482140 626316 482204 626380
rect 480852 625636 480916 625700
rect 478092 623596 478156 623660
rect 478276 622916 478340 622980
rect 483612 622236 483676 622300
rect 478460 621556 478524 621620
rect 479380 620876 479444 620940
rect 485820 619516 485884 619580
rect 483796 618836 483860 618900
rect 479564 618156 479628 618220
rect 481036 617476 481100 617540
rect 479932 616116 479996 616180
rect 485268 615436 485332 615500
rect 486004 614756 486068 614820
rect 481220 614076 481284 614140
rect 478644 613396 478708 613460
rect 482876 612716 482940 612780
rect 479748 612036 479812 612100
rect 482692 611356 482756 611420
rect 483428 610676 483492 610740
rect 477356 609996 477420 610060
rect 486372 609316 486436 609380
rect 485636 608636 485700 608700
rect 482876 608092 482940 608156
rect 484716 607956 484780 608020
rect 479932 607820 479996 607884
rect 486372 607684 486436 607748
rect 477356 607362 477420 607426
rect 481772 607276 481836 607340
rect 481588 607140 481652 607204
rect 483244 607140 483308 607204
rect 483060 607004 483124 607068
rect 483428 606868 483492 606932
rect 482692 606188 482756 606252
rect 479564 605916 479628 605980
rect 484900 605916 484964 605980
rect 481772 605644 481836 605708
rect 483796 605508 483860 605572
rect 478644 604828 478708 604892
rect 481220 604556 481284 604620
rect 484532 604556 484596 604620
rect 480300 604420 480364 604484
rect 484716 604284 484780 604348
rect 486004 604148 486068 604212
rect 485268 603604 485332 603668
rect 485820 603332 485884 603396
rect 484348 603196 484412 603260
rect 480484 603060 480548 603124
rect 484532 602924 484596 602988
rect 481404 602516 481468 602580
rect 479748 602380 479812 602444
rect 481036 602108 481100 602172
rect 479380 601836 479444 601900
rect 483428 601836 483492 601900
rect 477724 601700 477788 601764
rect 481772 601700 481836 601764
rect 484900 601564 484964 601628
rect 484348 601428 484412 601492
rect 481404 601020 481468 601084
rect 483428 601292 483492 601356
rect 483428 600476 483492 600540
rect 485636 600204 485700 600268
rect 483428 600068 483492 600132
rect 478460 599388 478524 599452
rect 483612 599252 483676 599316
rect 477908 599116 477972 599180
rect 478276 598572 478340 598636
rect 478092 598028 478156 598092
rect 477724 597756 477788 597820
rect 477908 597212 477972 597276
rect 480852 596668 480916 596732
rect 482140 596396 482204 596460
rect 483244 595988 483308 596052
rect 481588 595308 481652 595372
rect 480300 595036 480364 595100
rect 483060 594628 483124 594692
rect 481772 593948 481836 594012
rect 480484 593676 480548 593740
rect 483060 592996 483124 593060
rect 480668 592588 480732 592652
rect 483612 592180 483676 592244
rect 481772 591500 481836 591564
rect 483796 591364 483860 591428
rect 481588 590684 481652 590748
rect 480300 590140 480364 590204
rect 482140 589868 482204 589932
rect 483980 589460 484044 589524
rect 480852 588780 480916 588844
rect 482324 588508 482388 588572
rect 481036 587964 481100 588028
rect 480668 587828 480732 587892
rect 481220 587420 481284 587484
rect 479748 586604 479812 586668
rect 486188 585924 486252 585988
rect 486372 585788 486436 585852
rect 478092 585244 478156 585308
rect 478276 583884 478340 583948
rect 478644 583340 478708 583404
rect 478460 583068 478524 583132
rect 485452 582524 485516 582588
rect 481772 582388 481836 582452
rect 486004 581980 486068 582044
rect 485268 581844 485332 581908
rect 479748 581572 479812 581636
rect 483060 581572 483124 581636
rect 485820 581300 485884 581364
rect 481220 580892 481284 580956
rect 485084 580620 485148 580684
rect 485636 580484 485700 580548
rect 477356 579804 477420 579868
rect 481588 579532 481652 579596
rect 482876 579260 482940 579324
rect 480300 578988 480364 579052
rect 482508 578716 482572 578780
rect 482876 578036 482940 578100
rect 477356 577356 477420 577420
rect 485636 576676 485700 576740
rect 485084 575996 485148 576060
rect 485820 575316 485884 575380
rect 485268 574636 485332 574700
rect 486004 573956 486068 574020
rect 485452 573276 485516 573340
rect 478460 572596 478524 572660
rect 478644 571916 478708 571980
rect 478276 571236 478340 571300
rect 478092 569196 478156 569260
rect 486372 568516 486436 568580
rect 486372 567836 486436 567900
rect 482508 565796 482572 565860
rect 481036 565116 481100 565180
rect 482324 564436 482388 564500
rect 480852 563756 480916 563820
rect 483980 563076 484044 563140
rect 482140 562396 482204 562460
rect 483796 560356 483860 560420
rect 483612 558996 483676 559060
rect 480852 536556 480916 536620
rect 482140 535196 482204 535260
rect 478092 533836 478156 533900
rect 478276 532476 478340 532540
rect 483612 531796 483676 531860
rect 481036 531116 481100 531180
rect 479564 529756 479628 529820
rect 485084 529076 485148 529140
rect 486372 528396 486436 528460
rect 485268 527716 485332 527780
rect 481220 527036 481284 527100
rect 479380 526356 479444 526420
rect 483980 525676 484044 525740
rect 486004 524996 486068 525060
rect 479748 524316 479812 524380
rect 483796 523636 483860 523700
rect 480668 522956 480732 523020
rect 486372 522276 486436 522340
rect 485820 521596 485884 521660
rect 484532 520916 484596 520980
rect 484716 520236 484780 520300
rect 484348 519556 484412 519620
rect 484900 518876 484964 518940
rect 479564 518196 479628 518260
rect 479932 518196 479996 518260
rect 483980 517924 484044 517988
rect 484348 517652 484412 517716
rect 486188 517244 486252 517308
rect 484716 517108 484780 517172
rect 478460 516700 478524 516764
rect 484532 516564 484596 516628
rect 483060 516292 483124 516356
rect 481588 516156 481652 516220
rect 486004 515748 486068 515812
rect 484900 515612 484964 515676
rect 483428 515476 483492 515540
rect 480668 515204 480732 515268
rect 483796 515068 483860 515132
rect 483244 514932 483308 514996
rect 480484 514796 480548 514860
rect 479748 514388 479812 514452
rect 483428 514116 483492 514180
rect 484348 514116 484412 514180
rect 485820 513844 485884 513908
rect 481772 513708 481836 513772
rect 485084 513572 485148 513636
rect 484532 513436 484596 513500
rect 477540 513300 477604 513364
rect 480668 513300 480732 513364
rect 479932 513164 479996 513228
rect 479380 513028 479444 513092
rect 484348 512892 484412 512956
rect 478828 512756 478892 512820
rect 481220 512484 481284 512548
rect 485268 512212 485332 512276
rect 484348 512076 484412 512140
rect 481036 511940 481100 512004
rect 478644 511804 478708 511868
rect 478460 511668 478524 511732
rect 485636 511532 485700 511596
rect 481404 511396 481468 511460
rect 484348 511124 484412 511188
rect 484532 510852 484596 510916
rect 478828 510580 478892 510644
rect 481404 510036 481468 510100
rect 483612 509492 483676 509556
rect 478276 508948 478340 509012
rect 477540 508404 477604 508468
rect 478092 508132 478156 508196
rect 478644 507588 478708 507652
rect 482140 507044 482204 507108
rect 483060 506772 483124 506836
rect 480852 506228 480916 506292
rect 481588 505684 481652 505748
rect 483244 505412 483308 505476
rect 480484 504868 480548 504932
rect 481772 504324 481836 504388
rect 480668 504052 480732 504116
rect 483060 503236 483124 503300
rect 481772 502828 481836 502892
rect 477540 502420 477604 502484
rect 480668 501740 480732 501804
rect 483428 501604 483492 501668
rect 481588 500924 481652 500988
rect 480852 500380 480916 500444
rect 483612 500244 483676 500308
rect 482140 499564 482204 499628
rect 481036 499020 481100 499084
rect 483796 498884 483860 498948
rect 482324 498204 482388 498268
rect 481220 497660 481284 497724
rect 480300 497388 480364 497452
rect 480116 496844 480180 496908
rect 480668 496844 480732 496908
rect 479564 496300 479628 496364
rect 478092 495484 478156 495548
rect 478276 494940 478340 495004
rect 486004 494804 486068 494868
rect 481772 494668 481836 494732
rect 483060 494668 483124 494732
rect 480116 494320 480180 494324
rect 480116 494264 480166 494320
rect 480166 494264 480180 494320
rect 480116 494260 480180 494264
rect 486188 494124 486252 494188
rect 483428 493988 483492 494052
rect 483980 493444 484044 493508
rect 478460 492764 478524 492828
rect 477540 492628 477604 492692
rect 481588 492628 481652 492692
rect 478828 492220 478892 492284
rect 481956 491948 482020 492012
rect 481772 491540 481836 491604
rect 479564 491132 479628 491196
rect 484900 490860 484964 490924
rect 484532 490724 484596 490788
rect 477356 490106 477420 490170
rect 484348 489500 484412 489564
rect 483244 489364 483308 489428
rect 485452 488684 485516 488748
rect 480300 488548 480364 488612
rect 483244 488276 483308 488340
rect 484348 487596 484412 487660
rect 477356 486916 477420 486980
rect 484532 486236 484596 486300
rect 484900 485556 484964 485620
rect 481772 484876 481836 484940
rect 481956 484196 482020 484260
rect 478828 483516 478892 483580
rect 478460 482836 478524 482900
rect 483980 482156 484044 482220
rect 486372 480796 486436 480860
rect 486004 480116 486068 480180
rect 478276 479436 478340 479500
rect 478092 478756 478156 478820
rect 485452 476036 485516 476100
rect 481220 475356 481284 475420
rect 482324 474676 482388 474740
rect 483796 473996 483860 474060
rect 481036 473316 481100 473380
rect 482140 472636 482204 472700
rect 483612 471956 483676 472020
rect 480852 471276 480916 471340
rect 483612 452916 483676 452980
rect 478092 447476 478156 447540
rect 479380 443396 479444 443460
rect 479564 442716 479628 442780
rect 478276 442036 478340 442100
rect 478644 441356 478708 441420
rect 482140 440676 482204 440740
rect 480852 439996 480916 440060
rect 485636 439316 485700 439380
rect 483796 438636 483860 438700
rect 485268 437276 485332 437340
rect 486372 436596 486436 436660
rect 485084 435916 485148 435980
rect 485820 435236 485884 435300
rect 484532 434556 484596 434620
rect 486004 433876 486068 433940
rect 480116 433196 480180 433260
rect 477356 432516 477420 432580
rect 484716 431836 484780 431900
rect 481588 431156 481652 431220
rect 483244 430476 483308 430540
rect 484348 429796 484412 429860
rect 483060 429116 483124 429180
rect 484900 428436 484964 428500
rect 484532 428164 484596 428228
rect 485636 427892 485700 427956
rect 484348 427348 484412 427412
rect 477540 427212 477604 427276
rect 479932 427272 479996 427276
rect 479932 427216 479946 427272
rect 479946 427216 479996 427272
rect 479932 427212 479996 427216
rect 483244 426804 483308 426868
rect 481588 426532 481652 426596
rect 481956 426184 482020 426188
rect 481956 426128 482006 426184
rect 482006 426128 482020 426184
rect 481956 426124 482020 426128
rect 482508 426124 482572 426188
rect 484716 425988 484780 426052
rect 480852 425716 480916 425780
rect 486372 425716 486436 425780
rect 477356 425458 477420 425522
rect 480116 425172 480180 425236
rect 482876 425036 482940 425100
rect 483244 424900 483308 424964
rect 486372 424764 486436 424828
rect 483612 424628 483676 424692
rect 479748 424492 479812 424556
rect 484348 424356 484412 424420
rect 485820 423812 485884 423876
rect 484532 423676 484596 423740
rect 481220 423540 481284 423604
rect 483428 423540 483492 423604
rect 482876 423404 482940 423468
rect 483060 423268 483124 423332
rect 485084 423132 485148 423196
rect 480852 422996 480916 423060
rect 486188 422724 486252 422788
rect 485268 422452 485332 422516
rect 484716 422316 484780 422380
rect 484348 422180 484412 422244
rect 478644 421908 478708 421972
rect 486004 421772 486068 421836
rect 484716 421228 484780 421292
rect 477908 420956 477972 421020
rect 482140 420412 482204 420476
rect 485820 420276 485884 420340
rect 481220 420004 481284 420068
rect 484900 420004 484964 420068
rect 481404 419868 481468 419932
rect 481588 419732 481652 419796
rect 481956 419596 482020 419660
rect 480116 419520 480180 419524
rect 480116 419464 480166 419520
rect 480166 419464 480180 419520
rect 480116 419460 480180 419464
rect 484532 419324 484596 419388
rect 478276 419188 478340 419252
rect 479564 418644 479628 418708
rect 479380 418372 479444 418436
rect 478276 418236 478340 418300
rect 483244 418236 483308 418300
rect 479932 417828 479996 417892
rect 479748 417012 479812 417076
rect 484348 416876 484412 416940
rect 483244 416740 483308 416804
rect 478644 416664 478708 416668
rect 478644 416608 478694 416664
rect 478694 416608 478708 416664
rect 478644 416604 478708 416608
rect 482324 416604 482388 416668
rect 483060 416604 483124 416668
rect 480116 416468 480180 416532
rect 483796 416196 483860 416260
rect 484532 416196 484596 416260
rect 481772 415924 481836 415988
rect 478092 415652 478156 415716
rect 484716 415516 484780 415580
rect 484348 415380 484412 415444
rect 478460 415244 478524 415308
rect 483612 415244 483676 415308
rect 482876 415108 482940 415172
rect 482508 414564 482572 414628
rect 477540 414292 477604 414356
rect 479932 414156 479996 414220
rect 484532 414020 484596 414084
rect 478276 413748 478340 413812
rect 481404 413476 481468 413540
rect 484164 413476 484228 413540
rect 477908 413204 477972 413268
rect 478644 412932 478708 412996
rect 480300 412796 480364 412860
rect 484716 412660 484780 412724
rect 485820 412388 485884 412452
rect 480852 412116 480916 412180
rect 484348 412116 484412 412180
rect 480300 411844 480364 411908
rect 479932 411572 479996 411636
rect 484532 411436 484596 411500
rect 484164 411300 484228 411364
rect 484348 411028 484412 411092
rect 478460 410484 478524 410548
rect 483428 410212 483492 410276
rect 482876 410076 482940 410140
rect 484532 409940 484596 410004
rect 481588 409668 481652 409732
rect 483060 409124 483124 409188
rect 481956 408852 482020 408916
rect 484348 408716 484412 408780
rect 482876 408580 482940 408644
rect 483612 408308 483676 408372
rect 484348 407764 484412 407828
rect 482324 407492 482388 407556
rect 477540 406540 477604 406604
rect 477724 406404 477788 406468
rect 486188 405724 486252 405788
rect 479380 405180 479444 405244
rect 486004 405044 486068 405108
rect 486188 404364 486252 404428
rect 479564 403820 479628 403884
rect 479748 403684 479812 403748
rect 480852 403140 480916 403204
rect 478092 402460 478156 402524
rect 483244 402324 483308 402388
rect 477356 401712 477420 401776
rect 484900 401100 484964 401164
rect 484716 400964 484780 401028
rect 484532 400284 484596 400348
rect 484348 399740 484412 399804
rect 478644 399604 478708 399668
rect 477540 399468 477604 399532
rect 477724 398788 477788 398852
rect 478644 397836 478708 397900
rect 484348 397156 484412 397220
rect 484532 396476 484596 396540
rect 484716 395796 484780 395860
rect 484900 395116 484964 395180
rect 477356 394436 477420 394500
rect 483244 393756 483308 393820
rect 478092 393076 478156 393140
rect 480852 392396 480916 392460
rect 479748 391716 479812 391780
rect 479564 391036 479628 391100
rect 486372 390356 486436 390420
rect 486004 389676 486068 389740
rect 479380 388996 479444 389060
rect 486556 388316 486620 388380
rect 482140 357036 482204 357100
rect 483612 356356 483676 356420
rect 480852 355676 480916 355740
rect 478092 354316 478156 354380
rect 478276 352956 478340 353020
rect 478460 352276 478524 352340
rect 481036 351596 481100 351660
rect 482324 350916 482388 350980
rect 477908 350236 477972 350300
rect 481220 348876 481284 348940
rect 482692 348196 482756 348260
rect 482508 347516 482572 347580
rect 483796 346156 483860 346220
rect 479380 345476 479444 345540
rect 486004 344796 486068 344860
rect 481404 344116 481468 344180
rect 479748 343436 479812 343500
rect 483980 342756 484044 342820
rect 483428 342076 483492 342140
rect 484348 341396 484412 341460
rect 477356 340716 477420 340780
rect 478828 340036 478892 340100
rect 483244 339356 483308 339420
rect 479564 338676 479628 338740
rect 483428 338132 483492 338196
rect 483244 337588 483308 337652
rect 478828 337452 478892 337516
rect 477356 336840 477420 336904
rect 480300 336636 480364 336700
rect 481772 336636 481836 336700
rect 483060 336636 483124 336700
rect 484716 336636 484780 336700
rect 482692 336500 482756 336564
rect 484348 336228 484412 336292
rect 481220 335956 481284 336020
rect 477356 335820 477420 335884
rect 483980 335412 484044 335476
rect 484348 335276 484412 335340
rect 477908 335140 477972 335204
rect 479748 334868 479812 334932
rect 481404 334732 481468 334796
rect 479012 334596 479076 334660
rect 484716 334324 484780 334388
rect 486004 334188 486068 334252
rect 478644 334112 478708 334116
rect 478644 334056 478694 334112
rect 478694 334056 478708 334112
rect 478644 334052 478708 334056
rect 480484 334052 480548 334116
rect 483244 334052 483308 334116
rect 478828 333916 478892 333980
rect 477356 333848 477420 333912
rect 479380 333508 479444 333572
rect 483796 333372 483860 333436
rect 483428 333236 483492 333300
rect 484348 332964 484412 333028
rect 477356 332556 477420 332620
rect 479012 332420 479076 332484
rect 482508 332148 482572 332212
rect 482324 332012 482388 332076
rect 482876 331876 482940 331940
rect 478828 331604 478892 331668
rect 483428 331332 483492 331396
rect 477356 331128 477420 331192
rect 479564 330788 479628 330852
rect 482876 330516 482940 330580
rect 477908 329564 477972 329628
rect 481036 329428 481100 329492
rect 478460 329292 478524 329356
rect 478276 328612 478340 328676
rect 478644 328068 478708 328132
rect 478092 327932 478156 327996
rect 477908 327252 477972 327316
rect 480852 326708 480916 326772
rect 483612 326572 483676 326636
rect 482140 325892 482204 325956
rect 483060 325348 483124 325412
rect 480300 325076 480364 325140
rect 481772 324532 481836 324596
rect 483244 323988 483308 324052
rect 480484 323716 480548 323780
rect 481772 322900 481836 322964
rect 480668 322628 480732 322692
rect 483060 322084 483124 322148
rect 481588 321540 481652 321604
rect 480852 321268 480916 321332
rect 483612 320724 483676 320788
rect 483796 320180 483860 320244
rect 483980 319908 484044 319972
rect 481036 319364 481100 319428
rect 482140 318820 482204 318884
rect 480668 318684 480732 318748
rect 482324 318548 482388 318612
rect 481220 318004 481284 318068
rect 481404 317596 481468 317660
rect 479380 317188 479444 317252
rect 479748 316644 479812 316708
rect 479932 316100 479996 316164
rect 478092 315828 478156 315892
rect 478276 315284 478340 315348
rect 479380 314876 479444 314940
rect 486188 313924 486252 313988
rect 485084 313380 485148 313444
rect 486004 313108 486068 313172
rect 485820 312564 485884 312628
rect 485636 312020 485700 312084
rect 481772 311884 481836 311948
rect 484900 311748 484964 311812
rect 479748 311204 479812 311268
rect 483060 311204 483124 311268
rect 485268 311068 485332 311132
rect 485452 310660 485516 310724
rect 478644 310388 478708 310452
rect 479932 310448 479996 310452
rect 479932 310392 479982 310448
rect 479982 310392 479996 310448
rect 479932 310388 479996 310392
rect 481404 310448 481468 310452
rect 481404 310392 481454 310448
rect 481454 310392 481468 310448
rect 481404 310388 481468 310392
rect 482876 309844 482940 309908
rect 484348 309300 484412 309364
rect 481588 308892 481652 308956
rect 486188 308484 486252 308548
rect 484348 308076 484412 308140
rect 482876 307396 482940 307460
rect 478644 306716 478708 306780
rect 485452 306036 485516 306100
rect 485268 305356 485332 305420
rect 484900 304676 484964 304740
rect 485636 303996 485700 304060
rect 485820 303316 485884 303380
rect 486004 302636 486068 302700
rect 485084 301956 485148 302020
rect 486372 301276 486436 301340
rect 478276 299236 478340 299300
rect 478092 298556 478156 298620
rect 486372 295836 486436 295900
rect 481220 295156 481284 295220
rect 482324 294476 482388 294540
rect 482140 293796 482204 293860
rect 481036 293116 481100 293180
rect 483980 292436 484044 292500
rect 483796 291756 483860 291820
rect 483612 291076 483676 291140
rect 480852 290396 480916 290460
rect 483612 267276 483676 267340
rect 483796 265916 483860 265980
rect 480852 265236 480916 265300
rect 478092 262516 478156 262580
rect 482140 261836 482204 261900
rect 478276 261156 478340 261220
rect 482324 260476 482388 260540
rect 485636 259796 485700 259860
rect 481036 259116 481100 259180
rect 479564 258436 479628 258500
rect 483980 257756 484044 257820
rect 485452 257076 485516 257140
rect 479380 256396 479444 256460
rect 479748 255036 479812 255100
rect 486372 254356 486436 254420
rect 485820 253676 485884 253740
rect 479932 252996 479996 253060
rect 481220 252316 481284 252380
rect 486004 251636 486068 251700
rect 484532 250956 484596 251020
rect 484716 250276 484780 250340
rect 481588 249596 481652 249660
rect 484348 248916 484412 248980
rect 486004 248100 486068 248164
rect 477540 247964 477604 248028
rect 481220 247828 481284 247892
rect 481588 247692 481652 247756
rect 482876 247556 482940 247620
rect 484348 247420 484412 247484
rect 484716 247148 484780 247212
rect 477540 247012 477604 247076
rect 480300 247012 480364 247076
rect 481772 247012 481836 247076
rect 477172 246818 477236 246882
rect 477356 246876 477420 246940
rect 484532 246604 484596 246668
rect 479564 246332 479628 246396
rect 483244 246196 483308 246260
rect 482876 246060 482940 246124
rect 481036 245788 481100 245852
rect 477724 245652 477788 245716
rect 481588 245652 481652 245716
rect 477356 245458 477420 245522
rect 484532 245516 484596 245580
rect 479932 245244 479996 245308
rect 485820 244972 485884 245036
rect 484348 244836 484412 244900
rect 483244 244700 483308 244764
rect 486188 244428 486252 244492
rect 480484 244292 480548 244356
rect 484900 244156 484964 244220
rect 485636 244020 485700 244084
rect 479748 243884 479812 243948
rect 482324 243612 482388 243676
rect 483060 243476 483124 243540
rect 484716 243476 484780 243540
rect 484532 243204 484596 243268
rect 479380 243068 479444 243132
rect 477908 242796 477972 242860
rect 483244 242796 483308 242860
rect 484348 242660 484412 242724
rect 485452 242524 485516 242588
rect 483980 242252 484044 242316
rect 484348 242116 484412 242180
rect 478276 241980 478340 242044
rect 484900 241300 484964 241364
rect 484716 241164 484780 241228
rect 483244 241028 483308 241092
rect 484348 240892 484412 240956
rect 482140 239532 482204 239596
rect 478092 238988 478156 239052
rect 477540 238444 477604 238508
rect 477908 238172 477972 238236
rect 477724 237628 477788 237692
rect 480852 237084 480916 237148
rect 483796 236812 483860 236876
rect 481772 236268 481836 236332
rect 483612 235724 483676 235788
rect 480300 235452 480364 235516
rect 483060 234908 483124 234972
rect 481588 234364 481652 234428
rect 480484 234092 480548 234156
rect 483060 233140 483124 233204
rect 477724 232732 477788 232796
rect 477540 232324 477604 232388
rect 480668 231780 480732 231844
rect 483428 231644 483492 231708
rect 482876 230964 482940 231028
rect 480852 230420 480916 230484
rect 481588 230148 481652 230212
rect 483612 229740 483676 229804
rect 483796 229060 483860 229124
rect 482140 228788 482204 228852
rect 480484 228244 480548 228308
rect 482324 227700 482388 227764
rect 481036 227428 481100 227492
rect 480116 226884 480180 226948
rect 480668 226340 480732 226404
rect 481220 226204 481284 226268
rect 479564 225524 479628 225588
rect 479380 224980 479444 225044
rect 486188 224708 486252 224772
rect 482508 224164 482572 224228
rect 485452 224028 485516 224092
rect 480116 223680 480180 223684
rect 480116 223624 480166 223680
rect 480166 223624 480180 223680
rect 480116 223620 480180 223624
rect 482876 223680 482940 223684
rect 482876 223624 482926 223680
rect 482926 223624 482940 223680
rect 482876 223620 482940 223624
rect 483060 223620 483124 223684
rect 486188 223348 486252 223412
rect 483980 222804 484044 222868
rect 483428 222260 483492 222324
rect 486004 222260 486068 222324
rect 485268 221988 485332 222052
rect 485084 221444 485148 221508
rect 484716 221308 484780 221372
rect 477724 220900 477788 220964
rect 481036 220900 481100 220964
rect 481588 220900 481652 220964
rect 484532 220628 484596 220692
rect 484348 220084 484412 220148
rect 480484 219948 480548 220012
rect 481036 219948 481100 220012
rect 483060 219540 483124 219604
rect 477540 219268 477604 219332
rect 481404 218724 481468 218788
rect 483060 217636 483124 217700
rect 484348 216956 484412 217020
rect 484532 216276 484596 216340
rect 484716 215596 484780 215660
rect 485084 214916 485148 214980
rect 485268 214236 485332 214300
rect 486004 213556 486068 213620
rect 483980 212876 484044 212940
rect 486372 212196 486436 212260
rect 485452 211516 485516 211580
rect 482508 210836 482572 210900
rect 486556 210156 486620 210220
rect 479380 209476 479444 209540
rect 479564 208796 479628 208860
rect 481220 207436 481284 207500
rect 481404 206076 481468 206140
rect 482324 205396 482388 205460
rect 481036 204716 481100 204780
rect 482140 204036 482204 204100
rect 483796 203356 483860 203420
rect 483612 202676 483676 202740
rect 480852 201316 480916 201380
rect 482140 181596 482204 181660
rect 478276 180236 478340 180300
rect 479380 174796 479444 174860
rect 478092 174116 478156 174180
rect 483612 173436 483676 173500
rect 479564 172756 479628 172820
rect 482324 172076 482388 172140
rect 477908 171396 477972 171460
rect 482508 170716 482572 170780
rect 485268 170036 485332 170100
rect 483796 169356 483860 169420
rect 486004 168676 486068 168740
rect 485452 167316 485516 167380
rect 479748 165956 479812 166020
rect 485820 165276 485884 165340
rect 486372 164596 486436 164660
rect 480852 163916 480916 163980
rect 480300 163236 480364 163300
rect 484164 162556 484228 162620
rect 484716 161876 484780 161940
rect 485636 161196 485700 161260
rect 482876 160516 482940 160580
rect 483244 159836 483308 159900
rect 480484 159156 480548 159220
rect 477172 158476 477236 158540
rect 486188 158204 486252 158268
rect 483796 157932 483860 157996
rect 483244 157524 483308 157588
rect 483060 157388 483124 157452
rect 482876 156844 482940 156908
rect 480116 156708 480180 156772
rect 486004 156572 486068 156636
rect 484716 156028 484780 156092
rect 481588 155952 481652 155956
rect 481588 155896 481638 155952
rect 481638 155896 481652 155952
rect 481588 155892 481652 155896
rect 483244 155892 483308 155956
rect 485268 155892 485332 155956
rect 484348 155756 484412 155820
rect 484164 155484 484228 155548
rect 480300 155212 480364 155276
rect 484532 155076 484596 155140
rect 478644 154396 478708 154460
rect 484348 154260 484412 154324
rect 485820 153852 485884 153916
rect 479932 153716 479996 153780
rect 484532 153444 484596 153508
rect 479748 153308 479812 153372
rect 480484 153036 480548 153100
rect 480668 153036 480732 153100
rect 486004 153036 486068 153100
rect 477724 152900 477788 152964
rect 477540 152628 477604 152692
rect 485452 152492 485516 152556
rect 484716 152356 484780 152420
rect 478644 152220 478708 152284
rect 477908 151948 477972 152012
rect 480852 151676 480916 151740
rect 482140 151404 482204 151468
rect 484716 151132 484780 151196
rect 481956 150452 482020 150516
rect 483796 150452 483860 150516
rect 482508 150316 482572 150380
rect 484716 150316 484780 150380
rect 480668 150044 480732 150108
rect 477172 149746 477236 149810
rect 484348 149636 484412 149700
rect 479932 149500 479996 149564
rect 482324 149364 482388 149428
rect 481772 149228 481836 149292
rect 482140 149092 482204 149156
rect 485452 148956 485516 149020
rect 485636 148956 485700 149020
rect 479196 148820 479260 148884
rect 479564 148684 479628 148748
rect 479932 148744 479996 148748
rect 479932 148688 479982 148744
rect 479982 148688 479996 148744
rect 479932 148684 479996 148688
rect 483612 148412 483676 148476
rect 484532 148276 484596 148340
rect 484348 148140 484412 148204
rect 478092 147868 478156 147932
rect 477908 147732 477972 147796
rect 483428 147732 483492 147796
rect 479380 147324 479444 147388
rect 480668 147052 480732 147116
rect 479748 146916 479812 146980
rect 484532 146644 484596 146708
rect 480116 146508 480180 146572
rect 482324 146236 482388 146300
rect 483612 146236 483676 146300
rect 484532 146236 484596 146300
rect 479196 145964 479260 146028
rect 479932 145692 479996 145756
rect 484348 145556 484412 145620
rect 483244 145420 483308 145484
rect 481588 145148 481652 145212
rect 478644 144740 478708 144804
rect 481956 144332 482020 144396
rect 478828 144196 478892 144260
rect 484532 144060 484596 144124
rect 478276 143788 478340 143852
rect 484348 143652 484412 143716
rect 480116 143516 480180 143580
rect 477724 143244 477788 143308
rect 477540 142972 477604 143036
rect 480484 142836 480548 142900
rect 478828 142700 478892 142764
rect 484716 142428 484780 142492
rect 486004 142292 486068 142356
rect 480300 142156 480364 142220
rect 480484 141884 480548 141948
rect 480116 141612 480180 141676
rect 480300 141068 480364 141132
rect 478644 140524 478708 140588
rect 477908 140252 477972 140316
rect 483796 139708 483860 139772
rect 482140 139164 482204 139228
rect 483428 138892 483492 138956
rect 484532 138756 484596 138820
rect 485636 138620 485700 138684
rect 481772 138348 481836 138412
rect 483612 137804 483676 137868
rect 482324 137532 482388 137596
rect 484348 137396 484412 137460
rect 480668 137260 480732 137324
rect 484532 136988 484596 137052
rect 484348 136444 484412 136508
rect 483060 136172 483124 136236
rect 479748 135900 479812 135964
rect 485820 134404 485884 134468
rect 486004 133860 486068 133924
rect 478276 133588 478340 133652
rect 478092 133044 478156 133108
rect 486004 132500 486068 132564
rect 477356 132282 477420 132346
rect 481404 131684 481468 131748
rect 481588 131140 481652 131204
rect 484532 131004 484596 131068
rect 484348 130324 484412 130388
rect 483060 129916 483124 129980
rect 478828 129508 478892 129572
rect 483796 128420 483860 128484
rect 478828 127876 478892 127940
rect 483060 127196 483124 127260
rect 484348 126516 484412 126580
rect 484532 125836 484596 125900
rect 481588 125156 481652 125220
rect 481404 124476 481468 124540
rect 477356 123796 477420 123860
rect 486004 123116 486068 123180
rect 478092 122436 478156 122500
rect 478276 121756 478340 121820
rect 486372 121076 486436 121140
rect 486372 120396 486436 120460
rect 483796 119036 483860 119100
rect 6316 90884 6380 90948
rect 7604 90068 7668 90132
rect 60 89252 124 89316
rect 8892 88436 8956 88500
rect 3556 87620 3620 87684
rect 6500 86804 6564 86868
rect 480852 86396 480916 86460
rect 4660 85988 4724 86052
rect 483612 85716 483676 85780
rect 7420 85172 7484 85236
rect 7788 84356 7852 84420
rect 478092 83676 478156 83740
rect 6132 83540 6196 83604
rect 478276 82996 478340 83060
rect 5212 82724 5276 82788
rect 482140 82316 482204 82380
rect 1900 81908 1964 81972
rect 478460 81636 478524 81700
rect 7972 81092 8036 81156
rect 244 80276 308 80340
rect 485820 80276 485884 80340
rect 4844 79460 4908 79524
rect 479564 78916 479628 78980
rect 9076 78644 9140 78708
rect 486556 78236 486620 78300
rect 3372 77828 3436 77892
rect 479380 77556 479444 77620
rect 5028 77012 5092 77076
rect 481036 76876 481100 76940
rect 6316 76196 6380 76260
rect 482324 76196 482388 76260
rect 796 75924 860 75988
rect 60 75788 124 75852
rect 479748 75516 479812 75580
rect 8340 75380 8404 75444
rect 7788 74836 7852 74900
rect 484348 74836 484412 74900
rect 6316 74564 6380 74628
rect 7972 74156 8036 74220
rect 479932 74156 479996 74220
rect 7788 73748 7852 73812
rect 5212 73476 5276 73540
rect 484900 73476 484964 73540
rect 4108 72932 4172 72996
rect 6500 72796 6564 72860
rect 481404 72796 481468 72860
rect 3556 72116 3620 72180
rect 6684 72116 6748 72180
rect 484716 72116 484780 72180
rect 8340 71436 8404 71500
rect 484532 71436 484596 71500
rect 484348 70756 484412 70820
rect 483428 70076 483492 70140
rect 481588 69396 481652 69460
rect 2084 68852 2148 68916
rect 244 68444 308 68508
rect 483244 68716 483308 68780
rect 481404 68172 481468 68236
rect 5028 68036 5092 68100
rect 9260 68036 9324 68100
rect 478644 68036 478708 68100
rect 484164 67900 484228 67964
rect 481588 67628 481652 67692
rect 480300 67492 480364 67556
rect 481588 67492 481652 67556
rect 483060 67492 483124 67556
rect 7604 67356 7668 67420
rect 481772 67356 481836 67420
rect 5580 67220 5644 67284
rect 483244 67220 483308 67284
rect 483428 67084 483492 67148
rect 484348 66812 484412 66876
rect 4660 66676 4724 66740
rect 483244 66676 483308 66740
rect 3556 66404 3620 66468
rect 486188 66404 486252 66468
rect 484532 66268 484596 66332
rect 480116 66192 480180 66196
rect 480116 66136 480166 66192
rect 480166 66136 480180 66192
rect 480116 66132 480180 66136
rect 5580 65996 5644 66060
rect 483244 65996 483308 66060
rect 484164 65996 484228 66060
rect 483244 65860 483308 65924
rect 484716 65724 484780 65788
rect 479564 65452 479628 65516
rect 4108 65316 4172 65380
rect 477356 65316 477420 65380
rect 478644 65180 478708 65244
rect 484900 64908 484964 64972
rect 9260 64636 9324 64700
rect 481772 64636 481836 64700
rect 484348 64636 484412 64700
rect 479932 64364 479996 64428
rect 6684 63956 6748 64020
rect 484164 64092 484228 64156
rect 478644 63744 478708 63748
rect 478644 63688 478694 63744
rect 478694 63688 478708 63744
rect 478644 63684 478708 63688
rect 479748 63548 479812 63612
rect 7788 63276 7852 63340
rect 477172 63140 477236 63204
rect 482324 63004 482388 63068
rect 481036 62732 481100 62796
rect 4844 62596 4908 62660
rect 483428 62596 483492 62660
rect 477356 62460 477420 62524
rect 485268 62324 485332 62388
rect 480484 62188 480548 62252
rect 481772 62188 481836 62252
rect 6316 61916 6380 61980
rect 480116 61916 480180 61980
rect 481588 61916 481652 61980
rect 484348 61644 484412 61708
rect 479380 61372 479444 61436
rect 796 61236 860 61300
rect 483428 60828 483492 60892
rect 1348 60692 1412 60756
rect 7420 60692 7484 60756
rect 9076 60556 9140 60620
rect 477908 60556 477972 60620
rect 481588 60420 481652 60484
rect 477172 60284 477236 60348
rect 1900 59876 1964 59940
rect 478460 59468 478524 59532
rect 6132 59196 6196 59260
rect 482140 58924 482204 58988
rect 478276 58652 478340 58716
rect 1348 58516 1412 58580
rect 478092 58108 478156 58172
rect 477908 57564 477972 57628
rect 478644 57292 478708 57356
rect 483612 56748 483676 56812
rect 8892 56612 8956 56676
rect 480852 56204 480916 56268
rect 481956 55932 482020 55996
rect 483060 55388 483124 55452
rect 480300 54844 480364 54908
rect 481772 54572 481836 54636
rect 483244 54028 483308 54092
rect 480484 53484 480548 53548
rect 483060 52940 483124 53004
rect 3556 52396 3620 52460
rect 480852 52396 480916 52460
rect 483244 52124 483308 52188
rect 481772 51580 481836 51644
rect 483612 50900 483676 50964
rect 481588 50764 481652 50828
rect 481036 50220 481100 50284
rect 482140 49676 482204 49740
rect 483796 49404 483860 49468
rect 481220 48860 481284 48924
rect 2084 48316 2148 48380
rect 1348 48180 1412 48244
rect 3372 48180 3436 48244
rect 482324 48316 482388 48380
rect 480852 48180 480916 48244
rect 481404 48044 481468 48108
rect 480852 47500 480916 47564
rect 479932 47364 479996 47428
rect 479196 46684 479260 46748
rect 479564 46140 479628 46204
rect 479380 45596 479444 45660
rect 479748 45324 479812 45388
rect 479932 44372 479996 44436
rect 1348 44236 1412 44300
rect 485636 43964 485700 44028
rect 478092 43420 478156 43484
rect 483060 43284 483124 43348
rect 486004 43012 486068 43076
rect 478276 42604 478340 42668
rect 486004 42060 486068 42124
rect 476908 41448 476972 41512
rect 481772 41380 481836 41444
rect 483244 41380 483308 41444
rect 485452 41244 485516 41308
rect 484900 40700 484964 40764
rect 484716 40020 484780 40084
rect 479196 39884 479260 39948
rect 481588 39884 481652 39948
rect 484532 39748 484596 39812
rect 484348 39204 484412 39268
rect 485084 38660 485148 38724
rect 484348 38116 484412 38180
rect 484532 37436 484596 37500
rect 8340 36756 8404 36820
rect 484716 36756 484780 36820
rect 484900 36076 484964 36140
rect 485452 35396 485516 35460
rect 476988 34716 477052 34780
rect 486004 34036 486068 34100
rect 1348 33356 1412 33420
rect 478276 33356 478340 33420
rect 8340 32812 8404 32876
rect 1164 32676 1228 32740
rect 486372 32676 486436 32740
rect 8524 31996 8588 32060
rect 478092 31996 478156 32060
rect 1164 31588 1228 31652
rect 6132 31588 6196 31652
rect 485636 31316 485700 31380
rect 1348 30228 1412 30292
rect 3372 30228 3436 30292
rect 479748 29276 479812 29340
rect 479380 28596 479444 28660
rect 479564 27916 479628 27980
rect 1348 25876 1412 25940
rect 484900 25876 484964 25940
rect 9444 25468 9508 25532
rect 481404 25196 481468 25260
rect 4108 24516 4172 24580
rect 482324 24516 482388 24580
rect 481220 23836 481284 23900
rect 483796 23156 483860 23220
rect 9628 22476 9692 22540
rect 482140 22476 482204 22540
rect 4108 22204 4172 22268
rect 481036 21796 481100 21860
rect 8156 21116 8220 21180
rect 483612 20436 483676 20500
rect 9812 19076 9876 19140
rect 6684 18396 6748 18460
rect 1348 18124 1412 18188
rect 11100 18124 11164 18188
rect 4844 17036 4908 17100
rect 9628 17580 9692 17644
rect 12572 17444 12636 17508
rect 8156 17308 8220 17372
rect 11100 17172 11164 17236
rect 480852 17036 480916 17100
rect 12572 16900 12636 16964
rect 9812 16492 9876 16556
rect 6868 15948 6932 16012
rect 4844 15268 4908 15332
rect 6132 15132 6196 15196
rect 3372 14452 3436 14516
rect 796 13364 860 13428
rect 60 13228 124 13292
rect 18828 12820 18892 12884
rect 19564 12548 19628 12612
rect 3372 12140 3436 12204
rect 18828 12140 18892 12204
rect 15332 11732 15396 11796
rect 18828 11460 18892 11524
rect 18460 11188 18524 11252
rect 17172 10916 17236 10980
rect 18828 10780 18892 10844
rect 17356 10644 17420 10708
rect 20116 10100 20180 10164
rect 19932 9828 19996 9892
rect 18644 9284 18708 9348
rect 19564 8876 19628 8940
rect 15148 8740 15212 8804
rect 14412 8468 14476 8532
rect 15332 8060 15396 8124
rect 20300 7984 20364 7988
rect 20300 7928 20350 7984
rect 20350 7928 20364 7984
rect 20300 7924 20364 7928
rect 15148 7516 15212 7580
rect 17172 6836 17236 6900
rect 17356 6156 17420 6220
rect 9444 5612 9508 5676
rect 20116 5476 20180 5540
rect 14412 4796 14476 4860
rect 60 4388 124 4452
rect 19932 3436 19996 3500
rect 244 3028 308 3092
rect 1164 2892 1228 2956
rect 3372 2892 3436 2956
rect 1348 2348 1412 2412
rect 18644 2348 18708 2412
rect 18460 2076 18524 2140
rect 1164 1396 1228 1460
rect 8524 1260 8588 1324
rect 1348 716 1412 780
rect 20300 172 20364 236
<< metal4 >>
rect 21219 755852 21285 755853
rect 21219 755788 21220 755852
rect 21284 755788 21285 755852
rect 21219 755787 21285 755788
rect 19931 755036 19997 755037
rect 19931 754972 19932 755036
rect 19996 754972 19997 755036
rect 19931 754971 19997 754972
rect 6315 90948 6381 90949
rect 6315 90884 6316 90948
rect 6380 90884 6381 90948
rect 6315 90883 6381 90884
rect 59 89316 125 89317
rect 59 89252 60 89316
rect 124 89252 125 89316
rect 59 89251 125 89252
rect 62 75853 122 89251
rect 3555 87684 3621 87685
rect 3555 87620 3556 87684
rect 3620 87620 3621 87684
rect 3555 87619 3621 87620
rect 1899 81972 1965 81973
rect 1899 81908 1900 81972
rect 1964 81908 1965 81972
rect 1899 81907 1965 81908
rect 243 80340 309 80341
rect 243 80276 244 80340
rect 308 80276 309 80340
rect 243 80275 309 80276
rect 59 75852 125 75853
rect 59 75788 60 75852
rect 124 75788 125 75852
rect 59 75787 125 75788
rect 246 68509 306 80275
rect 795 75988 861 75989
rect 795 75924 796 75988
rect 860 75924 861 75988
rect 795 75923 861 75924
rect 243 68508 309 68509
rect 243 68444 244 68508
rect 308 68444 309 68508
rect 243 68443 309 68444
rect 798 61301 858 75923
rect 795 61300 861 61301
rect 795 61236 796 61300
rect 860 61236 861 61300
rect 795 61235 861 61236
rect 1347 60756 1413 60757
rect 1347 60692 1348 60756
rect 1412 60692 1413 60756
rect 1347 60691 1413 60692
rect 1350 58581 1410 60691
rect 1902 59941 1962 81907
rect 3371 77892 3437 77893
rect 3371 77828 3372 77892
rect 3436 77828 3437 77892
rect 3371 77827 3437 77828
rect 2083 68916 2149 68917
rect 2083 68852 2084 68916
rect 2148 68852 2149 68916
rect 2083 68851 2149 68852
rect 1899 59940 1965 59941
rect 1899 59876 1900 59940
rect 1964 59876 1965 59940
rect 1899 59875 1965 59876
rect 1347 58580 1413 58581
rect 1347 58516 1348 58580
rect 1412 58516 1413 58580
rect 1347 58515 1413 58516
rect 2086 48381 2146 68851
rect 2083 48380 2149 48381
rect 2083 48316 2084 48380
rect 2148 48316 2149 48380
rect 2083 48315 2149 48316
rect 3374 48245 3434 77827
rect 3558 72181 3618 87619
rect 4659 86052 4725 86053
rect 4659 85988 4660 86052
rect 4724 85988 4725 86052
rect 4659 85987 4725 85988
rect 4107 72996 4173 72997
rect 4107 72932 4108 72996
rect 4172 72932 4173 72996
rect 4107 72931 4173 72932
rect 3555 72180 3621 72181
rect 3555 72116 3556 72180
rect 3620 72116 3621 72180
rect 3555 72115 3621 72116
rect 3555 66468 3621 66469
rect 3555 66404 3556 66468
rect 3620 66404 3621 66468
rect 3555 66403 3621 66404
rect 3558 52461 3618 66403
rect 4110 65381 4170 72931
rect 4662 66741 4722 85987
rect 6131 83604 6197 83605
rect 6131 83540 6132 83604
rect 6196 83540 6197 83604
rect 6131 83539 6197 83540
rect 5211 82788 5277 82789
rect 5211 82724 5212 82788
rect 5276 82724 5277 82788
rect 5211 82723 5277 82724
rect 4843 79524 4909 79525
rect 4843 79460 4844 79524
rect 4908 79460 4909 79524
rect 4843 79459 4909 79460
rect 4659 66740 4725 66741
rect 4659 66676 4660 66740
rect 4724 66676 4725 66740
rect 4659 66675 4725 66676
rect 4107 65380 4173 65381
rect 4107 65316 4108 65380
rect 4172 65316 4173 65380
rect 4107 65315 4173 65316
rect 4846 62661 4906 79459
rect 5027 77076 5093 77077
rect 5027 77012 5028 77076
rect 5092 77012 5093 77076
rect 5027 77011 5093 77012
rect 5030 68101 5090 77011
rect 5214 73541 5274 82723
rect 5211 73540 5277 73541
rect 5211 73476 5212 73540
rect 5276 73476 5277 73540
rect 5211 73475 5277 73476
rect 5027 68100 5093 68101
rect 5027 68036 5028 68100
rect 5092 68036 5093 68100
rect 5027 68035 5093 68036
rect 5579 67284 5645 67285
rect 5579 67220 5580 67284
rect 5644 67220 5645 67284
rect 5579 67219 5645 67220
rect 5582 66061 5642 67219
rect 5579 66060 5645 66061
rect 5579 65996 5580 66060
rect 5644 65996 5645 66060
rect 5579 65995 5645 65996
rect 4843 62660 4909 62661
rect 4843 62596 4844 62660
rect 4908 62596 4909 62660
rect 4843 62595 4909 62596
rect 6134 59261 6194 83539
rect 6318 76261 6378 90883
rect 7603 90132 7669 90133
rect 7603 90068 7604 90132
rect 7668 90068 7669 90132
rect 7603 90067 7669 90068
rect 6499 86868 6565 86869
rect 6499 86804 6500 86868
rect 6564 86804 6565 86868
rect 6499 86803 6565 86804
rect 6315 76260 6381 76261
rect 6315 76196 6316 76260
rect 6380 76196 6381 76260
rect 6315 76195 6381 76196
rect 6315 74628 6381 74629
rect 6315 74564 6316 74628
rect 6380 74564 6381 74628
rect 6315 74563 6381 74564
rect 6318 61981 6378 74563
rect 6502 72861 6562 86803
rect 7419 85236 7485 85237
rect 7419 85172 7420 85236
rect 7484 85172 7485 85236
rect 7419 85171 7485 85172
rect 6499 72860 6565 72861
rect 6499 72796 6500 72860
rect 6564 72796 6565 72860
rect 6499 72795 6565 72796
rect 6683 72180 6749 72181
rect 6683 72116 6684 72180
rect 6748 72116 6749 72180
rect 6683 72115 6749 72116
rect 6686 64021 6746 72115
rect 6683 64020 6749 64021
rect 6683 63956 6684 64020
rect 6748 63956 6749 64020
rect 6683 63955 6749 63956
rect 6315 61980 6381 61981
rect 6315 61916 6316 61980
rect 6380 61916 6381 61980
rect 6315 61915 6381 61916
rect 7422 60757 7482 85171
rect 7606 67421 7666 90067
rect 8891 88500 8957 88501
rect 8891 88436 8892 88500
rect 8956 88436 8957 88500
rect 8891 88435 8957 88436
rect 7787 84420 7853 84421
rect 7787 84356 7788 84420
rect 7852 84356 7853 84420
rect 7787 84355 7853 84356
rect 7790 74901 7850 84355
rect 7971 81156 8037 81157
rect 7971 81092 7972 81156
rect 8036 81092 8037 81156
rect 7971 81091 8037 81092
rect 7787 74900 7853 74901
rect 7787 74836 7788 74900
rect 7852 74836 7853 74900
rect 7787 74835 7853 74836
rect 7974 74221 8034 81091
rect 8339 75444 8405 75445
rect 8339 75380 8340 75444
rect 8404 75380 8405 75444
rect 8339 75379 8405 75380
rect 7971 74220 8037 74221
rect 7971 74156 7972 74220
rect 8036 74156 8037 74220
rect 7971 74155 8037 74156
rect 7787 73812 7853 73813
rect 7787 73748 7788 73812
rect 7852 73748 7853 73812
rect 7787 73747 7853 73748
rect 7603 67420 7669 67421
rect 7603 67356 7604 67420
rect 7668 67356 7669 67420
rect 7603 67355 7669 67356
rect 7790 63341 7850 73747
rect 8342 71501 8402 75379
rect 8339 71500 8405 71501
rect 8339 71436 8340 71500
rect 8404 71436 8405 71500
rect 8339 71435 8405 71436
rect 7787 63340 7853 63341
rect 7787 63276 7788 63340
rect 7852 63276 7853 63340
rect 7787 63275 7853 63276
rect 7419 60756 7485 60757
rect 7419 60692 7420 60756
rect 7484 60692 7485 60756
rect 7419 60691 7485 60692
rect 6131 59260 6197 59261
rect 6131 59196 6132 59260
rect 6196 59196 6197 59260
rect 6131 59195 6197 59196
rect 8894 56677 8954 88435
rect 9075 78708 9141 78709
rect 9075 78644 9076 78708
rect 9140 78644 9141 78708
rect 9075 78643 9141 78644
rect 9078 60621 9138 78643
rect 9259 68100 9325 68101
rect 9259 68036 9260 68100
rect 9324 68036 9325 68100
rect 9259 68035 9325 68036
rect 9262 64701 9322 68035
rect 9259 64700 9325 64701
rect 9259 64636 9260 64700
rect 9324 64636 9325 64700
rect 9259 64635 9325 64636
rect 9075 60620 9141 60621
rect 9075 60556 9076 60620
rect 9140 60556 9141 60620
rect 9075 60555 9141 60556
rect 8891 56676 8957 56677
rect 8891 56612 8892 56676
rect 8956 56612 8957 56676
rect 8891 56611 8957 56612
rect 3555 52460 3621 52461
rect 3555 52396 3556 52460
rect 3620 52396 3621 52460
rect 3555 52395 3621 52396
rect 1347 48244 1413 48245
rect 1347 48180 1348 48244
rect 1412 48180 1413 48244
rect 1347 48179 1413 48180
rect 3371 48244 3437 48245
rect 3371 48180 3372 48244
rect 3436 48180 3437 48244
rect 3371 48179 3437 48180
rect 1350 44301 1410 48179
rect 1347 44300 1413 44301
rect 1347 44236 1348 44300
rect 1412 44236 1413 44300
rect 1347 44235 1413 44236
rect 8339 36820 8405 36821
rect 8339 36756 8340 36820
rect 8404 36756 8405 36820
rect 8339 36755 8405 36756
rect 1347 33420 1413 33421
rect 1347 33356 1348 33420
rect 1412 33356 1413 33420
rect 1347 33355 1413 33356
rect 1163 32740 1229 32741
rect 1163 32676 1164 32740
rect 1228 32676 1229 32740
rect 1163 32675 1229 32676
rect 1166 31653 1226 32675
rect 1163 31652 1229 31653
rect 1163 31588 1164 31652
rect 1228 31588 1229 31652
rect 1163 31587 1229 31588
rect 1350 30293 1410 33355
rect 8342 32877 8402 36755
rect 8339 32876 8405 32877
rect 8339 32812 8340 32876
rect 8404 32812 8405 32876
rect 8339 32811 8405 32812
rect 8523 32060 8589 32061
rect 8523 31996 8524 32060
rect 8588 31996 8589 32060
rect 8523 31995 8589 31996
rect 6131 31652 6197 31653
rect 6131 31588 6132 31652
rect 6196 31588 6197 31652
rect 6131 31587 6197 31588
rect 1347 30292 1413 30293
rect 1347 30228 1348 30292
rect 1412 30228 1413 30292
rect 1347 30227 1413 30228
rect 3371 30292 3437 30293
rect 3371 30228 3372 30292
rect 3436 30228 3437 30292
rect 3371 30227 3437 30228
rect 1347 25940 1413 25941
rect 1347 25876 1348 25940
rect 1412 25876 1413 25940
rect 1347 25875 1413 25876
rect 1350 18189 1410 25875
rect 1347 18188 1413 18189
rect 1347 18124 1348 18188
rect 1412 18124 1413 18188
rect 1347 18123 1413 18124
rect 3374 14517 3434 30227
rect 4107 24580 4173 24581
rect 4107 24516 4108 24580
rect 4172 24516 4173 24580
rect 4107 24515 4173 24516
rect 4110 22269 4170 24515
rect 4107 22268 4173 22269
rect 4107 22204 4108 22268
rect 4172 22204 4173 22268
rect 4107 22203 4173 22204
rect 4843 17100 4909 17101
rect 4843 17036 4844 17100
rect 4908 17036 4909 17100
rect 4843 17035 4909 17036
rect 4846 15333 4906 17035
rect 4843 15332 4909 15333
rect 4843 15268 4844 15332
rect 4908 15268 4909 15332
rect 4843 15267 4909 15268
rect 6134 15197 6194 31587
rect 8155 21180 8221 21181
rect 8155 21116 8156 21180
rect 8220 21116 8221 21180
rect 8155 21115 8221 21116
rect 6683 18460 6749 18461
rect 6683 18396 6684 18460
rect 6748 18396 6749 18460
rect 6683 18395 6749 18396
rect 6686 16010 6746 18395
rect 8158 17373 8218 21115
rect 8155 17372 8221 17373
rect 8155 17308 8156 17372
rect 8220 17308 8221 17372
rect 8155 17307 8221 17308
rect 6867 16012 6933 16013
rect 6867 16010 6868 16012
rect 6686 15950 6868 16010
rect 6867 15948 6868 15950
rect 6932 15948 6933 16012
rect 6867 15947 6933 15948
rect 6131 15196 6197 15197
rect 6131 15132 6132 15196
rect 6196 15132 6197 15196
rect 6131 15131 6197 15132
rect 3371 14516 3437 14517
rect 3371 14452 3372 14516
rect 3436 14452 3437 14516
rect 3371 14451 3437 14452
rect 795 13428 861 13429
rect 795 13364 796 13428
rect 860 13364 861 13428
rect 795 13363 861 13364
rect 59 13292 125 13293
rect 59 13228 60 13292
rect 124 13228 125 13292
rect 59 13227 125 13228
rect 62 4453 122 13227
rect 798 6930 858 13363
rect 3371 12204 3437 12205
rect 3371 12140 3372 12204
rect 3436 12140 3437 12204
rect 3371 12139 3437 12140
rect 246 6870 858 6930
rect 59 4452 125 4453
rect 59 4388 60 4452
rect 124 4388 125 4452
rect 59 4387 125 4388
rect 246 3093 306 6870
rect 243 3092 309 3093
rect 243 3028 244 3092
rect 308 3028 309 3092
rect 243 3027 309 3028
rect 3374 2957 3434 12139
rect 1163 2956 1229 2957
rect 1163 2892 1164 2956
rect 1228 2892 1229 2956
rect 1163 2891 1229 2892
rect 3371 2956 3437 2957
rect 3371 2892 3372 2956
rect 3436 2892 3437 2956
rect 3371 2891 3437 2892
rect 1166 1461 1226 2891
rect 1347 2412 1413 2413
rect 1347 2348 1348 2412
rect 1412 2348 1413 2412
rect 1347 2347 1413 2348
rect 1163 1460 1229 1461
rect 1163 1396 1164 1460
rect 1228 1396 1229 1460
rect 1163 1395 1229 1396
rect 1350 781 1410 2347
rect 8526 1325 8586 31995
rect 9443 25532 9509 25533
rect 9443 25468 9444 25532
rect 9508 25468 9509 25532
rect 9443 25467 9509 25468
rect 9446 5677 9506 25467
rect 9627 22540 9693 22541
rect 9627 22476 9628 22540
rect 9692 22476 9693 22540
rect 9627 22475 9693 22476
rect 9630 17645 9690 22475
rect 9811 19140 9877 19141
rect 9811 19076 9812 19140
rect 9876 19076 9877 19140
rect 9811 19075 9877 19076
rect 9627 17644 9693 17645
rect 9627 17580 9628 17644
rect 9692 17580 9693 17644
rect 9627 17579 9693 17580
rect 9814 16557 9874 19075
rect 11099 18188 11165 18189
rect 11099 18124 11100 18188
rect 11164 18124 11165 18188
rect 11099 18123 11165 18124
rect 11102 17237 11162 18123
rect 11099 17236 11165 17237
rect 11099 17172 11100 17236
rect 11164 17172 11165 17236
rect 11099 17171 11165 17172
rect 9811 16556 9877 16557
rect 9811 16492 9812 16556
rect 9876 16492 9877 16556
rect 9811 16491 9877 16492
rect 11944 6000 12264 748500
rect 12571 17508 12637 17509
rect 12571 17444 12572 17508
rect 12636 17444 12637 17508
rect 12571 17443 12637 17444
rect 12574 16965 12634 17443
rect 12571 16964 12637 16965
rect 12571 16900 12572 16964
rect 12636 16900 12637 16964
rect 12571 16899 12637 16900
rect 13004 6000 13324 748500
rect 15331 11796 15397 11797
rect 15331 11732 15332 11796
rect 15396 11732 15397 11796
rect 15331 11731 15397 11732
rect 15147 8804 15213 8805
rect 15147 8740 15148 8804
rect 15212 8740 15213 8804
rect 15147 8739 15213 8740
rect 14411 8532 14477 8533
rect 14411 8468 14412 8532
rect 14476 8468 14477 8532
rect 14411 8467 14477 8468
rect 9443 5676 9509 5677
rect 9443 5612 9444 5676
rect 9508 5612 9509 5676
rect 9443 5611 9509 5612
rect 14414 4861 14474 8467
rect 15150 7581 15210 8739
rect 15334 8125 15394 11731
rect 17171 10980 17237 10981
rect 17171 10916 17172 10980
rect 17236 10916 17237 10980
rect 17171 10915 17237 10916
rect 15331 8124 15397 8125
rect 15331 8060 15332 8124
rect 15396 8060 15397 8124
rect 15331 8059 15397 8060
rect 15147 7580 15213 7581
rect 15147 7516 15148 7580
rect 15212 7516 15213 7580
rect 15147 7515 15213 7516
rect 17174 6901 17234 10915
rect 17355 10708 17421 10709
rect 17355 10644 17356 10708
rect 17420 10644 17421 10708
rect 17355 10643 17421 10644
rect 17171 6900 17237 6901
rect 17171 6836 17172 6900
rect 17236 6836 17237 6900
rect 17171 6835 17237 6836
rect 17358 6221 17418 10643
rect 17355 6220 17421 6221
rect 17355 6156 17356 6220
rect 17420 6156 17421 6220
rect 17355 6155 17421 6156
rect 17944 6000 18264 748500
rect 18827 12884 18893 12885
rect 18827 12820 18828 12884
rect 18892 12820 18893 12884
rect 18827 12819 18893 12820
rect 18830 12205 18890 12819
rect 18827 12204 18893 12205
rect 18827 12140 18828 12204
rect 18892 12140 18893 12204
rect 18827 12139 18893 12140
rect 18827 11524 18893 11525
rect 18827 11460 18828 11524
rect 18892 11460 18893 11524
rect 18827 11459 18893 11460
rect 18459 11252 18525 11253
rect 18459 11188 18460 11252
rect 18524 11188 18525 11252
rect 18459 11187 18525 11188
rect 14411 4860 14477 4861
rect 14411 4796 14412 4860
rect 14476 4796 14477 4860
rect 14411 4795 14477 4796
rect 18462 2141 18522 11187
rect 18830 10845 18890 11459
rect 18827 10844 18893 10845
rect 18827 10780 18828 10844
rect 18892 10780 18893 10844
rect 18827 10779 18893 10780
rect 18643 9348 18709 9349
rect 18643 9284 18644 9348
rect 18708 9284 18709 9348
rect 18643 9283 18709 9284
rect 18646 2413 18706 9283
rect 19004 6000 19324 748500
rect 19934 743341 19994 754971
rect 20667 749460 20733 749461
rect 20667 749396 20668 749460
rect 20732 749396 20733 749460
rect 20667 749395 20733 749396
rect 20483 748644 20549 748645
rect 20483 748580 20484 748644
rect 20548 748580 20549 748644
rect 20483 748579 20549 748580
rect 19931 743340 19997 743341
rect 19931 743276 19932 743340
rect 19996 743276 19997 743340
rect 19931 743275 19997 743276
rect 20486 740077 20546 748579
rect 20670 741459 20730 749395
rect 21222 747690 21282 755787
rect 21222 747630 21340 747690
rect 21280 746899 21340 747630
rect 21277 746898 21343 746899
rect 21277 746834 21278 746898
rect 21342 746834 21343 746898
rect 21277 746833 21343 746834
rect 20667 741458 20733 741459
rect 20667 741394 20668 741458
rect 20732 741394 20733 741458
rect 20667 741393 20733 741394
rect 20483 740076 20549 740077
rect 20483 740012 20484 740076
rect 20548 740012 20549 740076
rect 20483 740011 20549 740012
rect 19563 12612 19629 12613
rect 19563 12548 19564 12612
rect 19628 12548 19629 12612
rect 19563 12547 19629 12548
rect 19566 8941 19626 12547
rect 20115 10164 20181 10165
rect 20115 10100 20116 10164
rect 20180 10100 20181 10164
rect 20115 10099 20181 10100
rect 19931 9892 19997 9893
rect 19931 9828 19932 9892
rect 19996 9828 19997 9892
rect 19931 9827 19997 9828
rect 19563 8940 19629 8941
rect 19563 8876 19564 8940
rect 19628 8876 19629 8940
rect 19563 8875 19629 8876
rect 19934 3501 19994 9827
rect 20118 5541 20178 10099
rect 20299 7988 20365 7989
rect 20299 7924 20300 7988
rect 20364 7924 20365 7988
rect 20299 7923 20365 7924
rect 20115 5540 20181 5541
rect 20115 5476 20116 5540
rect 20180 5476 20181 5540
rect 20115 5475 20181 5476
rect 19931 3500 19997 3501
rect 19931 3436 19932 3500
rect 19996 3436 19997 3500
rect 19931 3435 19997 3436
rect 18643 2412 18709 2413
rect 18643 2348 18644 2412
rect 18708 2348 18709 2412
rect 18643 2347 18709 2348
rect 18459 2140 18525 2141
rect 18459 2076 18460 2140
rect 18524 2076 18525 2140
rect 18459 2075 18525 2076
rect 8523 1324 8589 1325
rect 8523 1260 8524 1324
rect 8588 1260 8589 1324
rect 8523 1259 8589 1260
rect 1347 780 1413 781
rect 1347 716 1348 780
rect 1412 716 1413 780
rect 1347 715 1413 716
rect 20302 237 20362 7923
rect 23194 6000 23514 748500
rect 24254 6000 24574 748500
rect 29194 6000 29514 748500
rect 30254 6000 30574 748500
rect 35194 6000 35514 748500
rect 36254 6000 36574 748500
rect 41194 6000 41514 748500
rect 42254 6000 42574 748500
rect 47194 6000 47514 748500
rect 48254 6000 48574 748500
rect 53194 6000 53514 748500
rect 54254 6000 54574 748500
rect 59194 6000 59514 748500
rect 60254 6000 60574 748500
rect 64194 6000 64514 748500
rect 65254 6000 65574 748500
rect 70194 6000 70514 748500
rect 71254 6000 71574 748500
rect 76194 6000 76514 748500
rect 77254 6000 77574 748500
rect 82194 6000 82514 748500
rect 83254 6000 83574 748500
rect 88194 6000 88514 748500
rect 89254 6000 89574 748500
rect 94194 6000 94514 748500
rect 95254 6000 95574 748500
rect 100194 6000 100514 748500
rect 101254 6000 101574 748500
rect 105194 6000 105514 748500
rect 106254 6000 106574 748500
rect 111194 6000 111514 748500
rect 112254 6000 112574 748500
rect 117194 6000 117514 748500
rect 118254 6000 118574 748500
rect 123194 6000 123514 748500
rect 124254 6000 124574 748500
rect 129194 6000 129514 748500
rect 130254 6000 130574 748500
rect 135194 6000 135514 748500
rect 136254 6000 136574 748500
rect 141194 6000 141514 748500
rect 142254 6000 142574 748500
rect 147194 6000 147514 748500
rect 148254 6000 148574 748500
rect 154194 6000 154514 748500
rect 155254 6000 155574 748500
rect 160194 6000 160514 748500
rect 161254 6000 161574 748500
rect 166194 6000 166514 748500
rect 167254 6000 167574 748500
rect 172194 6000 172514 748500
rect 173254 6000 173574 748500
rect 178194 6000 178514 748500
rect 179254 6000 179574 748500
rect 184194 6000 184514 748500
rect 185254 6000 185574 748500
rect 190194 6000 190514 748500
rect 191254 6000 191574 748500
rect 195194 6000 195514 748500
rect 196254 6000 196574 748500
rect 201194 6000 201514 748500
rect 202254 6000 202574 748500
rect 207194 6000 207514 748500
rect 208254 6000 208574 748500
rect 213194 6000 213514 748500
rect 214254 6000 214574 748500
rect 219194 6000 219514 748500
rect 220254 6000 220574 748500
rect 225194 6000 225514 748500
rect 226254 6000 226574 748500
rect 231194 6000 231514 748500
rect 232254 6000 232574 748500
rect 236194 6000 236514 748500
rect 237254 6000 237574 748500
rect 242194 6000 242514 748500
rect 243254 6000 243574 748500
rect 248194 6000 248514 748500
rect 249254 6000 249574 748500
rect 254194 6000 254514 748500
rect 255254 6000 255574 748500
rect 260194 6000 260514 748500
rect 261254 6000 261574 748500
rect 266194 6000 266514 748500
rect 267254 6000 267574 748500
rect 272194 6000 272514 748500
rect 273254 6000 273574 748500
rect 277194 6000 277514 748500
rect 278254 6000 278574 748500
rect 283194 6000 283514 748500
rect 284254 6000 284574 748500
rect 289194 6000 289514 748500
rect 290254 6000 290574 748500
rect 295194 6000 295514 748500
rect 296254 6000 296574 748500
rect 301194 6000 301514 748500
rect 302254 6000 302574 748500
rect 307194 6000 307514 748500
rect 308254 6000 308574 748500
rect 313194 6000 313514 748500
rect 314254 6000 314574 748500
rect 322194 6000 322514 748500
rect 323254 6000 323574 748500
rect 328194 6000 328514 748500
rect 329254 6000 329574 748500
rect 334194 6000 334514 748500
rect 335254 6000 335574 748500
rect 340194 6000 340514 748500
rect 341254 6000 341574 748500
rect 346194 6000 346514 748500
rect 347254 6000 347574 748500
rect 352194 6000 352514 748500
rect 353254 6000 353574 748500
rect 358194 6000 358514 748500
rect 359254 6000 359574 748500
rect 363194 6000 363514 748500
rect 364254 6000 364574 748500
rect 369194 6000 369514 748500
rect 370254 6000 370574 748500
rect 375194 6000 375514 748500
rect 376254 6000 376574 748500
rect 381194 6000 381514 748500
rect 382254 6000 382574 748500
rect 387194 6000 387514 748500
rect 388254 6000 388574 748500
rect 393194 6000 393514 748500
rect 394254 6000 394574 748500
rect 399194 6000 399514 748500
rect 400254 6000 400574 748500
rect 404194 6000 404514 748500
rect 405254 6000 405574 748500
rect 410194 6000 410514 748500
rect 411254 6000 411574 748500
rect 416194 6000 416514 748500
rect 417254 6000 417574 748500
rect 422194 6000 422514 748500
rect 423254 6000 423574 748500
rect 428194 6000 428514 748500
rect 429254 6000 429574 748500
rect 434194 6000 434514 748500
rect 435254 6000 435574 748500
rect 440194 6000 440514 748500
rect 441254 6000 441574 748500
rect 445194 6000 445514 748500
rect 446254 6000 446574 748500
rect 451194 6000 451514 748500
rect 452254 6000 452574 748500
rect 457194 6000 457514 748500
rect 458254 6000 458574 748500
rect 463194 6000 463514 748500
rect 464254 6000 464574 748500
rect 469194 6000 469514 748500
rect 470254 6000 470574 748500
rect 475194 6000 475514 748500
rect 480115 737220 480181 737221
rect 480115 737156 480116 737220
rect 480180 737156 480181 737220
rect 480115 737155 480181 737156
rect 479379 716140 479445 716141
rect 479379 716076 479380 716140
rect 479444 716076 479445 716140
rect 479379 716075 479445 716076
rect 478091 711380 478157 711381
rect 478091 711316 478092 711380
rect 478156 711316 478157 711380
rect 478091 711315 478157 711316
rect 477171 710020 477237 710021
rect 477171 709956 477172 710020
rect 477236 709956 477237 710020
rect 477171 709955 477237 709956
rect 477174 702450 477234 709955
rect 476990 702390 477234 702450
rect 476990 693293 477050 702390
rect 477539 696964 477605 696965
rect 477539 696900 477540 696964
rect 477604 696900 477605 696964
rect 477539 696899 477605 696900
rect 476929 693292 477050 693293
rect 476929 693228 476930 693292
rect 476994 693230 477050 693292
rect 476994 693228 476995 693230
rect 476929 693227 476995 693228
rect 477171 692340 477237 692341
rect 477171 692276 477172 692340
rect 477236 692276 477237 692340
rect 477171 692275 477237 692276
rect 477174 683130 477234 692275
rect 477542 683501 477602 696899
rect 477723 694244 477789 694245
rect 477723 694180 477724 694244
rect 477788 694180 477789 694244
rect 477723 694179 477789 694180
rect 477539 683500 477605 683501
rect 477539 683436 477540 683500
rect 477604 683436 477605 683500
rect 477539 683435 477605 683436
rect 476990 683070 477234 683130
rect 476990 670850 477050 683070
rect 477726 682957 477786 694179
rect 478094 691933 478154 711315
rect 478275 709340 478341 709341
rect 478275 709276 478276 709340
rect 478340 709276 478341 709340
rect 478275 709275 478341 709276
rect 478278 694925 478338 709275
rect 478459 707300 478525 707301
rect 478459 707236 478460 707300
rect 478524 707236 478525 707300
rect 478459 707235 478525 707236
rect 478275 694924 478341 694925
rect 478275 694860 478276 694924
rect 478340 694860 478341 694924
rect 478275 694859 478341 694860
rect 478091 691932 478157 691933
rect 478091 691868 478092 691932
rect 478156 691868 478157 691932
rect 478091 691867 478157 691868
rect 477907 691388 477973 691389
rect 477907 691324 477908 691388
rect 477972 691324 477973 691388
rect 477907 691323 477973 691324
rect 477723 682956 477789 682957
rect 477723 682892 477724 682956
rect 477788 682892 477789 682956
rect 477723 682891 477789 682892
rect 477723 679692 477789 679693
rect 477723 679628 477724 679692
rect 477788 679628 477789 679692
rect 477723 679627 477789 679628
rect 477726 670989 477786 679627
rect 477910 678877 477970 691323
rect 478275 684452 478341 684453
rect 478275 684388 478276 684452
rect 478340 684388 478341 684452
rect 478275 684387 478341 684388
rect 478091 681868 478157 681869
rect 478091 681804 478092 681868
rect 478156 681804 478157 681868
rect 478091 681803 478157 681804
rect 477907 678876 477973 678877
rect 477907 678812 477908 678876
rect 477972 678812 477973 678876
rect 477907 678811 477973 678812
rect 478094 678061 478154 681803
rect 478278 679965 478338 684387
rect 478275 679964 478341 679965
rect 478275 679900 478276 679964
rect 478340 679900 478341 679964
rect 478275 679899 478341 679900
rect 478462 679149 478522 707235
rect 478643 699412 478709 699413
rect 478643 699348 478644 699412
rect 478708 699348 478709 699412
rect 478643 699347 478709 699348
rect 478646 698189 478706 699347
rect 478643 698188 478709 698189
rect 478643 698124 478644 698188
rect 478708 698124 478709 698188
rect 478643 698123 478709 698124
rect 478827 695604 478893 695605
rect 478827 695540 478828 695604
rect 478892 695540 478893 695604
rect 478827 695539 478893 695540
rect 478643 692340 478709 692341
rect 478643 692276 478644 692340
rect 478708 692276 478709 692340
rect 478643 692275 478709 692276
rect 478646 691117 478706 692275
rect 478643 691116 478709 691117
rect 478643 691052 478644 691116
rect 478708 691052 478709 691116
rect 478643 691051 478709 691052
rect 478830 685677 478890 695539
rect 479382 686493 479442 716075
rect 479747 702540 479813 702541
rect 479747 702476 479748 702540
rect 479812 702476 479813 702540
rect 479747 702475 479813 702476
rect 479379 686492 479445 686493
rect 479379 686428 479380 686492
rect 479444 686428 479445 686492
rect 479379 686427 479445 686428
rect 479563 685812 479629 685813
rect 479563 685748 479564 685812
rect 479628 685748 479629 685812
rect 479563 685747 479629 685748
rect 478827 685676 478893 685677
rect 478827 685612 478828 685676
rect 478892 685612 478893 685676
rect 478827 685611 478893 685612
rect 479379 684860 479445 684861
rect 479379 684796 479380 684860
rect 479444 684796 479445 684860
rect 479379 684795 479445 684796
rect 479195 680372 479261 680373
rect 479195 680308 479196 680372
rect 479260 680308 479261 680372
rect 479195 680307 479261 680308
rect 478459 679148 478525 679149
rect 478459 679084 478460 679148
rect 478524 679084 478525 679148
rect 478459 679083 478525 679084
rect 478459 678468 478525 678469
rect 478459 678404 478460 678468
rect 478524 678404 478525 678468
rect 478459 678403 478525 678404
rect 478091 678060 478157 678061
rect 478091 677996 478092 678060
rect 478156 677996 478157 678060
rect 478091 677995 478157 677996
rect 478462 673709 478522 678403
rect 479011 677516 479077 677517
rect 479011 677452 479012 677516
rect 479076 677452 479077 677516
rect 479011 677451 479077 677452
rect 478459 673708 478525 673709
rect 478459 673644 478460 673708
rect 478524 673644 478525 673708
rect 478459 673643 478525 673644
rect 477723 670988 477789 670989
rect 477723 670924 477724 670988
rect 477788 670924 477789 670988
rect 477723 670923 477789 670924
rect 476910 670790 477050 670850
rect 476910 670513 476970 670790
rect 476907 670512 476973 670513
rect 476907 670448 476908 670512
rect 476972 670448 476973 670512
rect 476907 670447 476973 670448
rect 479014 669629 479074 677451
rect 479198 673437 479258 680307
rect 479382 675885 479442 684795
rect 479566 683773 479626 685747
rect 479750 685405 479810 702475
rect 479931 700500 479997 700501
rect 479931 700436 479932 700500
rect 479996 700436 479997 700500
rect 479931 700435 479997 700436
rect 479747 685404 479813 685405
rect 479747 685340 479748 685404
rect 479812 685340 479813 685404
rect 479747 685339 479813 685340
rect 479747 684180 479813 684181
rect 479747 684116 479748 684180
rect 479812 684116 479813 684180
rect 479747 684115 479813 684116
rect 479563 683772 479629 683773
rect 479563 683708 479564 683772
rect 479628 683708 479629 683772
rect 479563 683707 479629 683708
rect 479379 675884 479445 675885
rect 479379 675820 479380 675884
rect 479444 675820 479445 675884
rect 479379 675819 479445 675820
rect 479563 675884 479629 675885
rect 479563 675820 479564 675884
rect 479628 675820 479629 675884
rect 479563 675819 479629 675820
rect 479195 673436 479261 673437
rect 479195 673372 479196 673436
rect 479260 673372 479261 673436
rect 479195 673371 479261 673372
rect 479566 669901 479626 675819
rect 479750 674797 479810 684115
rect 479934 684045 479994 700435
rect 480118 698325 480178 737155
rect 482875 735180 482941 735181
rect 482875 735116 482876 735180
rect 482940 735116 482941 735180
rect 482875 735115 482941 735116
rect 480851 715460 480917 715461
rect 480851 715396 480852 715460
rect 480916 715396 480917 715460
rect 480851 715395 480917 715396
rect 480115 698324 480181 698325
rect 480115 698260 480116 698324
rect 480180 698260 480181 698324
rect 480115 698259 480181 698260
rect 480483 693564 480549 693565
rect 480483 693500 480484 693564
rect 480548 693500 480549 693564
rect 480483 693499 480549 693500
rect 480299 690028 480365 690029
rect 480299 689964 480300 690028
rect 480364 689964 480365 690028
rect 480299 689963 480365 689964
rect 480115 685540 480181 685541
rect 480115 685476 480116 685540
rect 480180 685476 480181 685540
rect 480115 685475 480181 685476
rect 479931 684044 479997 684045
rect 479931 683980 479932 684044
rect 479996 683980 479997 684044
rect 479931 683979 479997 683980
rect 480118 680509 480178 685475
rect 480302 681189 480362 689963
rect 480486 687581 480546 693499
rect 480854 693429 480914 715395
rect 481035 714780 481101 714781
rect 481035 714716 481036 714780
rect 481100 714716 481101 714780
rect 481035 714715 481101 714716
rect 481038 693565 481098 714715
rect 481403 705260 481469 705261
rect 481403 705196 481404 705260
rect 481468 705196 481469 705260
rect 481403 705195 481469 705196
rect 481035 693564 481101 693565
rect 481035 693500 481036 693564
rect 481100 693500 481101 693564
rect 481035 693499 481101 693500
rect 480851 693428 480917 693429
rect 480851 693364 480852 693428
rect 480916 693364 480917 693428
rect 480851 693363 480917 693364
rect 480851 693156 480917 693157
rect 480851 693092 480852 693156
rect 480916 693092 480917 693156
rect 480851 693091 480917 693092
rect 480483 687580 480549 687581
rect 480483 687516 480484 687580
rect 480548 687516 480549 687580
rect 480483 687515 480549 687516
rect 480854 687037 480914 693091
rect 481219 692748 481285 692749
rect 481219 692684 481220 692748
rect 481284 692684 481285 692748
rect 481219 692683 481285 692684
rect 481222 689077 481282 692683
rect 481219 689076 481285 689077
rect 481219 689012 481220 689076
rect 481284 689012 481285 689076
rect 481219 689011 481285 689012
rect 481035 688260 481101 688261
rect 481035 688196 481036 688260
rect 481100 688196 481101 688260
rect 481035 688195 481101 688196
rect 480851 687036 480917 687037
rect 480851 686972 480852 687036
rect 480916 686972 480917 687036
rect 480851 686971 480917 686972
rect 481038 685810 481098 688195
rect 481219 687172 481285 687173
rect 481219 687108 481220 687172
rect 481284 687108 481285 687172
rect 481219 687107 481285 687108
rect 480854 685750 481098 685810
rect 480299 681188 480365 681189
rect 480299 681124 480300 681188
rect 480364 681124 480365 681188
rect 480299 681123 480365 681124
rect 480115 680508 480181 680509
rect 480115 680444 480116 680508
rect 480180 680444 480181 680508
rect 480115 680443 480181 680444
rect 480667 676156 480733 676157
rect 480667 676092 480668 676156
rect 480732 676092 480733 676156
rect 480667 676091 480733 676092
rect 479747 674796 479813 674797
rect 479747 674732 479748 674796
rect 479812 674732 479813 674796
rect 479747 674731 479813 674732
rect 480670 673165 480730 676091
rect 480667 673164 480733 673165
rect 480667 673100 480668 673164
rect 480732 673100 480733 673164
rect 480667 673099 480733 673100
rect 480854 672621 480914 685750
rect 481222 683130 481282 687107
rect 481038 683070 481282 683130
rect 481038 677245 481098 683070
rect 481406 682685 481466 705195
rect 482878 703765 482938 735115
rect 483611 725660 483677 725661
rect 483611 725596 483612 725660
rect 483676 725596 483677 725660
rect 483611 725595 483677 725596
rect 482875 703764 482941 703765
rect 482875 703700 482876 703764
rect 482940 703700 482941 703764
rect 482875 703699 482941 703700
rect 482875 699140 482941 699141
rect 482875 699076 482876 699140
rect 482940 699076 482941 699140
rect 482875 699075 482941 699076
rect 482323 698460 482389 698461
rect 482323 698396 482324 698460
rect 482388 698396 482389 698460
rect 482323 698395 482389 698396
rect 481587 696420 481653 696421
rect 481587 696356 481588 696420
rect 481652 696356 481653 696420
rect 481587 696355 481653 696356
rect 481590 691661 481650 696355
rect 482139 693020 482205 693021
rect 482139 692956 482140 693020
rect 482204 692956 482205 693020
rect 482139 692955 482205 692956
rect 481587 691660 481653 691661
rect 481587 691596 481588 691660
rect 481652 691596 481653 691660
rect 481587 691595 481653 691596
rect 481587 685812 481653 685813
rect 481587 685748 481588 685812
rect 481652 685748 481653 685812
rect 481587 685747 481653 685748
rect 481403 682684 481469 682685
rect 481403 682620 481404 682684
rect 481468 682620 481469 682684
rect 481403 682619 481469 682620
rect 481403 680780 481469 680781
rect 481403 680716 481404 680780
rect 481468 680716 481469 680780
rect 481403 680715 481469 680716
rect 481406 677789 481466 680715
rect 481403 677788 481469 677789
rect 481403 677724 481404 677788
rect 481468 677724 481469 677788
rect 481403 677723 481469 677724
rect 481035 677244 481101 677245
rect 481035 677180 481036 677244
rect 481100 677180 481101 677244
rect 481035 677179 481101 677180
rect 480851 672620 480917 672621
rect 480851 672556 480852 672620
rect 480916 672556 480917 672620
rect 480851 672555 480917 672556
rect 481590 670173 481650 685747
rect 482142 680917 482202 692955
rect 482326 686765 482386 698395
rect 482878 696285 482938 699075
rect 483614 697373 483674 725595
rect 483979 722940 484045 722941
rect 483979 722876 483980 722940
rect 484044 722876 484045 722940
rect 483979 722875 484045 722876
rect 483795 719540 483861 719541
rect 483795 719476 483796 719540
rect 483860 719476 483861 719540
rect 483795 719475 483861 719476
rect 483611 697372 483677 697373
rect 483611 697308 483612 697372
rect 483676 697308 483677 697372
rect 483611 697307 483677 697308
rect 483427 697100 483493 697101
rect 483427 697036 483428 697100
rect 483492 697036 483493 697100
rect 483427 697035 483493 697036
rect 482875 696284 482941 696285
rect 482875 696220 482876 696284
rect 482940 696220 482941 696284
rect 482875 696219 482941 696220
rect 483059 690028 483125 690029
rect 483059 689964 483060 690028
rect 483124 689964 483125 690028
rect 483059 689963 483125 689964
rect 482323 686764 482389 686765
rect 482323 686700 482324 686764
rect 482388 686700 482389 686764
rect 482323 686699 482389 686700
rect 482139 680916 482205 680917
rect 482139 680852 482140 680916
rect 482204 680852 482205 680916
rect 482139 680851 482205 680852
rect 482139 680372 482205 680373
rect 482139 680308 482140 680372
rect 482204 680308 482205 680372
rect 482139 680307 482205 680308
rect 481955 679012 482021 679013
rect 481955 678948 481956 679012
rect 482020 678948 482021 679012
rect 481955 678947 482021 678948
rect 481771 678196 481837 678197
rect 481771 678132 481772 678196
rect 481836 678132 481837 678196
rect 481771 678131 481837 678132
rect 481587 670172 481653 670173
rect 481587 670108 481588 670172
rect 481652 670108 481653 670172
rect 481587 670107 481653 670108
rect 479563 669900 479629 669901
rect 479563 669836 479564 669900
rect 479628 669836 479629 669900
rect 479563 669835 479629 669836
rect 479011 669628 479077 669629
rect 479011 669564 479012 669628
rect 479076 669564 479077 669628
rect 479011 669563 479077 669564
rect 481774 669357 481834 678131
rect 481958 672893 482018 678947
rect 482142 675613 482202 680307
rect 483062 679149 483122 689963
rect 483243 686220 483309 686221
rect 483243 686156 483244 686220
rect 483308 686156 483309 686220
rect 483243 686155 483309 686156
rect 483246 684725 483306 686155
rect 483243 684724 483309 684725
rect 483243 684660 483244 684724
rect 483308 684660 483309 684724
rect 483243 684659 483309 684660
rect 483243 684588 483309 684589
rect 483243 684524 483244 684588
rect 483308 684524 483309 684588
rect 483243 684523 483309 684524
rect 483059 679148 483125 679149
rect 483059 679084 483060 679148
rect 483124 679084 483125 679148
rect 483059 679083 483125 679084
rect 483059 678468 483125 678469
rect 483059 678404 483060 678468
rect 483124 678404 483125 678468
rect 483059 678403 483125 678404
rect 483062 676565 483122 678403
rect 483059 676564 483125 676565
rect 483059 676500 483060 676564
rect 483124 676500 483125 676564
rect 483059 676499 483125 676500
rect 483059 676292 483125 676293
rect 483059 676228 483060 676292
rect 483124 676228 483125 676292
rect 483059 676227 483125 676228
rect 482139 675612 482205 675613
rect 482139 675548 482140 675612
rect 482204 675548 482205 675612
rect 482139 675547 482205 675548
rect 483062 674117 483122 676227
rect 483059 674116 483125 674117
rect 483059 674052 483060 674116
rect 483124 674052 483125 674116
rect 483059 674051 483125 674052
rect 481955 672892 482021 672893
rect 481955 672828 481956 672892
rect 482020 672828 482021 672892
rect 481955 672827 482021 672828
rect 483246 671669 483306 684523
rect 483430 678469 483490 697035
rect 483611 696964 483677 696965
rect 483611 696900 483612 696964
rect 483676 696900 483677 696964
rect 483611 696899 483677 696900
rect 483614 690573 483674 696899
rect 483798 696829 483858 719475
rect 483982 697237 484042 722875
rect 484899 720900 484965 720901
rect 484899 720836 484900 720900
rect 484964 720836 484965 720900
rect 484899 720835 484965 720836
rect 484163 710700 484229 710701
rect 484163 710636 484164 710700
rect 484228 710636 484229 710700
rect 484163 710635 484229 710636
rect 483979 697236 484045 697237
rect 483979 697172 483980 697236
rect 484044 697172 484045 697236
rect 483979 697171 484045 697172
rect 483795 696828 483861 696829
rect 483795 696764 483796 696828
rect 483860 696764 483861 696828
rect 483795 696763 483861 696764
rect 483979 694108 484045 694109
rect 483979 694044 483980 694108
rect 484044 694044 484045 694108
rect 483979 694043 484045 694044
rect 483982 690845 484042 694043
rect 483979 690844 484045 690845
rect 483979 690780 483980 690844
rect 484044 690780 484045 690844
rect 483979 690779 484045 690780
rect 483611 690572 483677 690573
rect 483611 690508 483612 690572
rect 483676 690508 483677 690572
rect 483611 690507 483677 690508
rect 483611 690300 483677 690301
rect 483611 690236 483612 690300
rect 483676 690236 483677 690300
rect 483611 690235 483677 690236
rect 483614 684589 483674 690235
rect 484166 689757 484226 710635
rect 484902 699413 484962 720835
rect 486371 712740 486437 712741
rect 486371 712676 486372 712740
rect 486436 712676 486437 712740
rect 486371 712675 486437 712676
rect 486003 708660 486069 708661
rect 486003 708596 486004 708660
rect 486068 708596 486069 708660
rect 486003 708595 486069 708596
rect 485819 707980 485885 707981
rect 485819 707916 485820 707980
rect 485884 707916 485885 707980
rect 485819 707915 485885 707916
rect 485083 706620 485149 706621
rect 485083 706556 485084 706620
rect 485148 706556 485149 706620
rect 485083 706555 485149 706556
rect 484899 699412 484965 699413
rect 484899 699348 484900 699412
rect 484964 699348 484965 699412
rect 484899 699347 484965 699348
rect 484347 690980 484413 690981
rect 484347 690916 484348 690980
rect 484412 690916 484413 690980
rect 484347 690915 484413 690916
rect 484163 689756 484229 689757
rect 484163 689692 484164 689756
rect 484228 689692 484229 689756
rect 484163 689691 484229 689692
rect 483611 684588 483677 684589
rect 483611 684524 483612 684588
rect 483676 684524 483677 684588
rect 483611 684523 483677 684524
rect 483611 684452 483677 684453
rect 483611 684388 483612 684452
rect 483676 684388 483677 684452
rect 483611 684387 483677 684388
rect 483427 678468 483493 678469
rect 483427 678404 483428 678468
rect 483492 678404 483493 678468
rect 483427 678403 483493 678404
rect 483614 678330 483674 684387
rect 484350 683229 484410 690915
rect 484715 683500 484781 683501
rect 484715 683436 484716 683500
rect 484780 683436 484781 683500
rect 484715 683435 484781 683436
rect 484347 683228 484413 683229
rect 484347 683164 484348 683228
rect 484412 683164 484413 683228
rect 484347 683163 484413 683164
rect 484531 682820 484597 682821
rect 484531 682756 484532 682820
rect 484596 682756 484597 682820
rect 484531 682755 484597 682756
rect 484347 682140 484413 682141
rect 484347 682076 484348 682140
rect 484412 682076 484413 682140
rect 484347 682075 484413 682076
rect 484350 681325 484410 682075
rect 484347 681324 484413 681325
rect 484347 681260 484348 681324
rect 484412 681260 484413 681324
rect 484347 681259 484413 681260
rect 483795 679148 483861 679149
rect 483795 679084 483796 679148
rect 483860 679084 483861 679148
rect 483795 679083 483861 679084
rect 483430 678270 483674 678330
rect 483243 671668 483309 671669
rect 483243 671604 483244 671668
rect 483308 671604 483309 671668
rect 483243 671603 483309 671604
rect 481771 669356 481837 669357
rect 481771 669292 481772 669356
rect 481836 669292 481837 669356
rect 481771 669291 481837 669292
rect 483430 668949 483490 678270
rect 483611 676156 483677 676157
rect 483611 676092 483612 676156
rect 483676 676092 483677 676156
rect 483611 676091 483677 676092
rect 483614 672077 483674 676091
rect 483798 675477 483858 679083
rect 483795 675476 483861 675477
rect 483795 675412 483796 675476
rect 483860 675412 483861 675476
rect 483795 675411 483861 675412
rect 483795 674796 483861 674797
rect 483795 674732 483796 674796
rect 483860 674732 483861 674796
rect 483795 674731 483861 674732
rect 483611 672076 483677 672077
rect 483611 672012 483612 672076
rect 483676 672012 483677 672076
rect 483611 672011 483677 672012
rect 483798 669221 483858 674731
rect 484534 674661 484594 682755
rect 484718 682005 484778 683435
rect 484715 682004 484781 682005
rect 484715 681940 484716 682004
rect 484780 681940 484781 682004
rect 484715 681939 484781 681940
rect 485086 679693 485146 706555
rect 485267 705940 485333 705941
rect 485267 705876 485268 705940
rect 485332 705876 485333 705940
rect 485267 705875 485333 705876
rect 485270 697917 485330 705875
rect 485635 704580 485701 704581
rect 485635 704516 485636 704580
rect 485700 704516 485701 704580
rect 485635 704515 485701 704516
rect 485451 703220 485517 703221
rect 485451 703156 485452 703220
rect 485516 703156 485517 703220
rect 485451 703155 485517 703156
rect 485267 697916 485333 697917
rect 485267 697852 485268 697916
rect 485332 697852 485333 697916
rect 485267 697851 485333 697852
rect 485267 695740 485333 695741
rect 485267 695676 485268 695740
rect 485332 695676 485333 695740
rect 485267 695675 485333 695676
rect 485270 688125 485330 695675
rect 485454 695197 485514 703155
rect 485451 695196 485517 695197
rect 485451 695132 485452 695196
rect 485516 695132 485517 695196
rect 485451 695131 485517 695132
rect 485638 694517 485698 704515
rect 485822 696557 485882 707915
rect 485819 696556 485885 696557
rect 485819 696492 485820 696556
rect 485884 696492 485885 696556
rect 485819 696491 485885 696492
rect 485635 694516 485701 694517
rect 485635 694452 485636 694516
rect 485700 694452 485701 694516
rect 485635 694451 485701 694452
rect 486006 693837 486066 708595
rect 486374 702450 486434 712675
rect 486190 702390 486434 702450
rect 486003 693836 486069 693837
rect 486003 693772 486004 693836
rect 486068 693772 486069 693836
rect 486003 693771 486069 693772
rect 486190 693290 486250 702390
rect 486371 701180 486437 701181
rect 486371 701116 486372 701180
rect 486436 701116 486437 701180
rect 486371 701115 486437 701116
rect 485638 693230 486250 693290
rect 485267 688124 485333 688125
rect 485267 688060 485268 688124
rect 485332 688060 485333 688124
rect 485267 688059 485333 688060
rect 485638 687173 485698 693230
rect 486374 692610 486434 701115
rect 486006 692550 486434 692610
rect 486006 692205 486066 692550
rect 486003 692204 486069 692205
rect 486003 692140 486004 692204
rect 486068 692140 486069 692204
rect 486003 692139 486069 692140
rect 485819 691660 485885 691661
rect 485819 691596 485820 691660
rect 485884 691596 485885 691660
rect 485819 691595 485885 691596
rect 485635 687172 485701 687173
rect 485635 687108 485636 687172
rect 485700 687108 485701 687172
rect 485635 687107 485701 687108
rect 485451 686900 485517 686901
rect 485451 686836 485452 686900
rect 485516 686836 485517 686900
rect 485451 686835 485517 686836
rect 485083 679692 485149 679693
rect 485083 679628 485084 679692
rect 485148 679628 485149 679692
rect 485083 679627 485149 679628
rect 485454 676837 485514 686835
rect 485635 681460 485701 681461
rect 485635 681396 485636 681460
rect 485700 681396 485701 681460
rect 485635 681395 485701 681396
rect 485451 676836 485517 676837
rect 485451 676772 485452 676836
rect 485516 676772 485517 676836
rect 485451 676771 485517 676772
rect 484531 674660 484597 674661
rect 484531 674596 484532 674660
rect 484596 674596 484597 674660
rect 484531 674595 484597 674596
rect 485638 672485 485698 681395
rect 485822 679557 485882 691595
rect 486371 680100 486437 680101
rect 486371 680036 486372 680100
rect 486436 680036 486437 680100
rect 486371 680035 486437 680036
rect 485819 679556 485885 679557
rect 485819 679492 485820 679556
rect 485884 679492 485885 679556
rect 485819 679491 485885 679492
rect 486374 674389 486434 680035
rect 486371 674388 486437 674389
rect 486371 674324 486372 674388
rect 486436 674324 486437 674388
rect 486371 674323 486437 674324
rect 485635 672484 485701 672485
rect 485635 672420 485636 672484
rect 485700 672420 485701 672484
rect 485635 672419 485701 672420
rect 483795 669220 483861 669221
rect 483795 669156 483796 669220
rect 483860 669156 483861 669220
rect 483795 669155 483861 669156
rect 483427 668948 483493 668949
rect 483427 668884 483428 668948
rect 483492 668884 483493 668948
rect 483427 668883 483493 668884
rect 482139 626380 482205 626381
rect 482139 626316 482140 626380
rect 482204 626316 482205 626380
rect 482139 626315 482205 626316
rect 480851 625700 480917 625701
rect 480851 625636 480852 625700
rect 480916 625636 480917 625700
rect 480851 625635 480917 625636
rect 478091 623660 478157 623661
rect 478091 623596 478092 623660
rect 478156 623596 478157 623660
rect 478091 623595 478157 623596
rect 477355 610060 477421 610061
rect 477355 609996 477356 610060
rect 477420 609996 477421 610060
rect 477355 609995 477421 609996
rect 477358 607427 477418 609995
rect 477355 607426 477421 607427
rect 477355 607362 477356 607426
rect 477420 607362 477421 607426
rect 477355 607361 477421 607362
rect 477723 601764 477789 601765
rect 477723 601700 477724 601764
rect 477788 601700 477789 601764
rect 477723 601699 477789 601700
rect 477726 597821 477786 601699
rect 477907 599180 477973 599181
rect 477907 599116 477908 599180
rect 477972 599116 477973 599180
rect 477907 599115 477973 599116
rect 477723 597820 477789 597821
rect 477723 597756 477724 597820
rect 477788 597756 477789 597820
rect 477723 597755 477789 597756
rect 477910 597277 477970 599115
rect 478094 598093 478154 623595
rect 478275 622980 478341 622981
rect 478275 622916 478276 622980
rect 478340 622916 478341 622980
rect 478275 622915 478341 622916
rect 478278 598637 478338 622915
rect 478459 621620 478525 621621
rect 478459 621556 478460 621620
rect 478524 621556 478525 621620
rect 478459 621555 478525 621556
rect 478462 599453 478522 621555
rect 479379 620940 479445 620941
rect 479379 620876 479380 620940
rect 479444 620876 479445 620940
rect 479379 620875 479445 620876
rect 478643 613460 478709 613461
rect 478643 613396 478644 613460
rect 478708 613396 478709 613460
rect 478643 613395 478709 613396
rect 478646 604893 478706 613395
rect 478643 604892 478709 604893
rect 478643 604828 478644 604892
rect 478708 604828 478709 604892
rect 478643 604827 478709 604828
rect 479382 601901 479442 620875
rect 479563 618220 479629 618221
rect 479563 618156 479564 618220
rect 479628 618156 479629 618220
rect 479563 618155 479629 618156
rect 479566 605981 479626 618155
rect 479931 616180 479997 616181
rect 479931 616116 479932 616180
rect 479996 616116 479997 616180
rect 479931 616115 479997 616116
rect 479747 612100 479813 612101
rect 479747 612036 479748 612100
rect 479812 612036 479813 612100
rect 479747 612035 479813 612036
rect 479563 605980 479629 605981
rect 479563 605916 479564 605980
rect 479628 605916 479629 605980
rect 479563 605915 479629 605916
rect 479750 602445 479810 612035
rect 479934 607885 479994 616115
rect 479931 607884 479997 607885
rect 479931 607820 479932 607884
rect 479996 607820 479997 607884
rect 479931 607819 479997 607820
rect 480299 604484 480365 604485
rect 480299 604420 480300 604484
rect 480364 604420 480365 604484
rect 480299 604419 480365 604420
rect 479747 602444 479813 602445
rect 479747 602380 479748 602444
rect 479812 602380 479813 602444
rect 479747 602379 479813 602380
rect 479379 601900 479445 601901
rect 479379 601836 479380 601900
rect 479444 601836 479445 601900
rect 479379 601835 479445 601836
rect 478459 599452 478525 599453
rect 478459 599388 478460 599452
rect 478524 599388 478525 599452
rect 478459 599387 478525 599388
rect 478275 598636 478341 598637
rect 478275 598572 478276 598636
rect 478340 598572 478341 598636
rect 478275 598571 478341 598572
rect 478091 598092 478157 598093
rect 478091 598028 478092 598092
rect 478156 598028 478157 598092
rect 478091 598027 478157 598028
rect 477907 597276 477973 597277
rect 477907 597212 477908 597276
rect 477972 597212 477973 597276
rect 477907 597211 477973 597212
rect 480302 595101 480362 604419
rect 480483 603124 480549 603125
rect 480483 603060 480484 603124
rect 480548 603060 480549 603124
rect 480483 603059 480549 603060
rect 480299 595100 480365 595101
rect 480299 595036 480300 595100
rect 480364 595036 480365 595100
rect 480299 595035 480365 595036
rect 480486 593741 480546 603059
rect 480854 596733 480914 625635
rect 481035 617540 481101 617541
rect 481035 617476 481036 617540
rect 481100 617476 481101 617540
rect 481035 617475 481101 617476
rect 481038 602173 481098 617475
rect 481219 614140 481285 614141
rect 481219 614076 481220 614140
rect 481284 614076 481285 614140
rect 481219 614075 481285 614076
rect 481222 604621 481282 614075
rect 481771 607340 481837 607341
rect 481771 607276 481772 607340
rect 481836 607276 481837 607340
rect 481771 607275 481837 607276
rect 481587 607204 481653 607205
rect 481587 607140 481588 607204
rect 481652 607140 481653 607204
rect 481587 607139 481653 607140
rect 481219 604620 481285 604621
rect 481219 604556 481220 604620
rect 481284 604556 481285 604620
rect 481219 604555 481285 604556
rect 481403 602580 481469 602581
rect 481403 602516 481404 602580
rect 481468 602516 481469 602580
rect 481403 602515 481469 602516
rect 481035 602172 481101 602173
rect 481035 602108 481036 602172
rect 481100 602108 481101 602172
rect 481035 602107 481101 602108
rect 481406 601085 481466 602515
rect 481403 601084 481469 601085
rect 481403 601020 481404 601084
rect 481468 601020 481469 601084
rect 481403 601019 481469 601020
rect 480851 596732 480917 596733
rect 480851 596668 480852 596732
rect 480916 596668 480917 596732
rect 480851 596667 480917 596668
rect 481590 595373 481650 607139
rect 481774 605709 481834 607275
rect 481771 605708 481837 605709
rect 481771 605644 481772 605708
rect 481836 605644 481837 605708
rect 481771 605643 481837 605644
rect 481771 601764 481837 601765
rect 481771 601700 481772 601764
rect 481836 601700 481837 601764
rect 481771 601699 481837 601700
rect 481587 595372 481653 595373
rect 481587 595308 481588 595372
rect 481652 595308 481653 595372
rect 481587 595307 481653 595308
rect 481774 594013 481834 601699
rect 482142 596461 482202 626315
rect 483611 622300 483677 622301
rect 483611 622236 483612 622300
rect 483676 622236 483677 622300
rect 483611 622235 483677 622236
rect 482875 612780 482941 612781
rect 482875 612716 482876 612780
rect 482940 612716 482941 612780
rect 482875 612715 482941 612716
rect 482691 611420 482757 611421
rect 482691 611356 482692 611420
rect 482756 611356 482757 611420
rect 482691 611355 482757 611356
rect 482694 606253 482754 611355
rect 482878 608157 482938 612715
rect 483427 610740 483493 610741
rect 483427 610676 483428 610740
rect 483492 610676 483493 610740
rect 483427 610675 483493 610676
rect 482875 608156 482941 608157
rect 482875 608092 482876 608156
rect 482940 608092 482941 608156
rect 482875 608091 482941 608092
rect 483243 607204 483309 607205
rect 483243 607140 483244 607204
rect 483308 607140 483309 607204
rect 483243 607139 483309 607140
rect 483059 607068 483125 607069
rect 483059 607004 483060 607068
rect 483124 607004 483125 607068
rect 483059 607003 483125 607004
rect 482691 606252 482757 606253
rect 482691 606188 482692 606252
rect 482756 606188 482757 606252
rect 482691 606187 482757 606188
rect 482139 596460 482205 596461
rect 482139 596396 482140 596460
rect 482204 596396 482205 596460
rect 482139 596395 482205 596396
rect 483062 594693 483122 607003
rect 483246 596053 483306 607139
rect 483430 606933 483490 610675
rect 483427 606932 483493 606933
rect 483427 606868 483428 606932
rect 483492 606868 483493 606932
rect 483427 606867 483493 606868
rect 483427 601900 483493 601901
rect 483427 601836 483428 601900
rect 483492 601836 483493 601900
rect 483427 601835 483493 601836
rect 483430 601357 483490 601835
rect 483427 601356 483493 601357
rect 483427 601292 483428 601356
rect 483492 601292 483493 601356
rect 483427 601291 483493 601292
rect 483427 600540 483493 600541
rect 483427 600476 483428 600540
rect 483492 600476 483493 600540
rect 483427 600475 483493 600476
rect 483430 600133 483490 600475
rect 483427 600132 483493 600133
rect 483427 600068 483428 600132
rect 483492 600068 483493 600132
rect 483427 600067 483493 600068
rect 483614 599317 483674 622235
rect 485819 619580 485885 619581
rect 485819 619516 485820 619580
rect 485884 619516 485885 619580
rect 485819 619515 485885 619516
rect 483795 618900 483861 618901
rect 483795 618836 483796 618900
rect 483860 618836 483861 618900
rect 483795 618835 483861 618836
rect 483798 605573 483858 618835
rect 485267 615500 485333 615501
rect 485267 615436 485268 615500
rect 485332 615436 485333 615500
rect 485267 615435 485333 615436
rect 484715 608020 484781 608021
rect 484715 607956 484716 608020
rect 484780 607956 484781 608020
rect 484715 607955 484781 607956
rect 483795 605572 483861 605573
rect 483795 605508 483796 605572
rect 483860 605508 483861 605572
rect 483795 605507 483861 605508
rect 484531 604620 484597 604621
rect 484531 604556 484532 604620
rect 484596 604556 484597 604620
rect 484531 604555 484597 604556
rect 484347 603260 484413 603261
rect 484347 603196 484348 603260
rect 484412 603196 484413 603260
rect 484347 603195 484413 603196
rect 484350 601493 484410 603195
rect 484534 602989 484594 604555
rect 484718 604349 484778 607955
rect 484899 605980 484965 605981
rect 484899 605916 484900 605980
rect 484964 605916 484965 605980
rect 484899 605915 484965 605916
rect 484715 604348 484781 604349
rect 484715 604284 484716 604348
rect 484780 604284 484781 604348
rect 484715 604283 484781 604284
rect 484531 602988 484597 602989
rect 484531 602924 484532 602988
rect 484596 602924 484597 602988
rect 484531 602923 484597 602924
rect 484902 601629 484962 605915
rect 485270 603669 485330 615435
rect 485635 608700 485701 608701
rect 485635 608636 485636 608700
rect 485700 608636 485701 608700
rect 485635 608635 485701 608636
rect 485267 603668 485333 603669
rect 485267 603604 485268 603668
rect 485332 603604 485333 603668
rect 485267 603603 485333 603604
rect 484899 601628 484965 601629
rect 484899 601564 484900 601628
rect 484964 601564 484965 601628
rect 484899 601563 484965 601564
rect 484347 601492 484413 601493
rect 484347 601428 484348 601492
rect 484412 601428 484413 601492
rect 484347 601427 484413 601428
rect 485638 600269 485698 608635
rect 485822 603397 485882 619515
rect 486003 614820 486069 614821
rect 486003 614756 486004 614820
rect 486068 614756 486069 614820
rect 486003 614755 486069 614756
rect 486006 604213 486066 614755
rect 486371 609380 486437 609381
rect 486371 609316 486372 609380
rect 486436 609316 486437 609380
rect 486371 609315 486437 609316
rect 486374 607749 486434 609315
rect 486371 607748 486437 607749
rect 486371 607684 486372 607748
rect 486436 607684 486437 607748
rect 486371 607683 486437 607684
rect 486003 604212 486069 604213
rect 486003 604148 486004 604212
rect 486068 604148 486069 604212
rect 486003 604147 486069 604148
rect 485819 603396 485885 603397
rect 485819 603332 485820 603396
rect 485884 603332 485885 603396
rect 485819 603331 485885 603332
rect 485635 600268 485701 600269
rect 485635 600204 485636 600268
rect 485700 600204 485701 600268
rect 485635 600203 485701 600204
rect 483611 599316 483677 599317
rect 483611 599252 483612 599316
rect 483676 599252 483677 599316
rect 483611 599251 483677 599252
rect 483243 596052 483309 596053
rect 483243 595988 483244 596052
rect 483308 595988 483309 596052
rect 483243 595987 483309 595988
rect 483059 594692 483125 594693
rect 483059 594628 483060 594692
rect 483124 594628 483125 594692
rect 483059 594627 483125 594628
rect 481771 594012 481837 594013
rect 481771 593948 481772 594012
rect 481836 593948 481837 594012
rect 481771 593947 481837 593948
rect 480483 593740 480549 593741
rect 480483 593676 480484 593740
rect 480548 593676 480549 593740
rect 480483 593675 480549 593676
rect 483059 593060 483125 593061
rect 483059 592996 483060 593060
rect 483124 592996 483125 593060
rect 483059 592995 483125 592996
rect 480667 592652 480733 592653
rect 480667 592588 480668 592652
rect 480732 592588 480733 592652
rect 480667 592587 480733 592588
rect 480299 590204 480365 590205
rect 480299 590140 480300 590204
rect 480364 590140 480365 590204
rect 480299 590139 480365 590140
rect 479747 586668 479813 586669
rect 479747 586604 479748 586668
rect 479812 586604 479813 586668
rect 479747 586603 479813 586604
rect 478091 585308 478157 585309
rect 478091 585244 478092 585308
rect 478156 585244 478157 585308
rect 478091 585243 478157 585244
rect 477355 579868 477421 579869
rect 477355 579804 477356 579868
rect 477420 579804 477421 579868
rect 477355 579803 477421 579804
rect 477358 577421 477418 579803
rect 477355 577420 477421 577421
rect 477355 577356 477356 577420
rect 477420 577356 477421 577420
rect 477355 577355 477421 577356
rect 478094 569261 478154 585243
rect 478275 583948 478341 583949
rect 478275 583884 478276 583948
rect 478340 583884 478341 583948
rect 478275 583883 478341 583884
rect 478278 571301 478338 583883
rect 478643 583404 478709 583405
rect 478643 583340 478644 583404
rect 478708 583340 478709 583404
rect 478643 583339 478709 583340
rect 478459 583132 478525 583133
rect 478459 583068 478460 583132
rect 478524 583068 478525 583132
rect 478459 583067 478525 583068
rect 478462 572661 478522 583067
rect 478459 572660 478525 572661
rect 478459 572596 478460 572660
rect 478524 572596 478525 572660
rect 478459 572595 478525 572596
rect 478646 571981 478706 583339
rect 479750 581637 479810 586603
rect 479747 581636 479813 581637
rect 479747 581572 479748 581636
rect 479812 581572 479813 581636
rect 479747 581571 479813 581572
rect 480302 579053 480362 590139
rect 480670 587893 480730 592587
rect 481771 591564 481837 591565
rect 481771 591500 481772 591564
rect 481836 591500 481837 591564
rect 481771 591499 481837 591500
rect 481587 590748 481653 590749
rect 481587 590684 481588 590748
rect 481652 590684 481653 590748
rect 481587 590683 481653 590684
rect 480851 588844 480917 588845
rect 480851 588780 480852 588844
rect 480916 588780 480917 588844
rect 480851 588779 480917 588780
rect 480667 587892 480733 587893
rect 480667 587828 480668 587892
rect 480732 587828 480733 587892
rect 480667 587827 480733 587828
rect 480299 579052 480365 579053
rect 480299 578988 480300 579052
rect 480364 578988 480365 579052
rect 480299 578987 480365 578988
rect 478643 571980 478709 571981
rect 478643 571916 478644 571980
rect 478708 571916 478709 571980
rect 478643 571915 478709 571916
rect 478275 571300 478341 571301
rect 478275 571236 478276 571300
rect 478340 571236 478341 571300
rect 478275 571235 478341 571236
rect 478091 569260 478157 569261
rect 478091 569196 478092 569260
rect 478156 569196 478157 569260
rect 478091 569195 478157 569196
rect 480854 563821 480914 588779
rect 481035 588028 481101 588029
rect 481035 587964 481036 588028
rect 481100 587964 481101 588028
rect 481035 587963 481101 587964
rect 481038 565181 481098 587963
rect 481219 587484 481285 587485
rect 481219 587420 481220 587484
rect 481284 587420 481285 587484
rect 481219 587419 481285 587420
rect 481222 580957 481282 587419
rect 481219 580956 481285 580957
rect 481219 580892 481220 580956
rect 481284 580892 481285 580956
rect 481219 580891 481285 580892
rect 481590 579597 481650 590683
rect 481774 582453 481834 591499
rect 482139 589932 482205 589933
rect 482139 589868 482140 589932
rect 482204 589868 482205 589932
rect 482139 589867 482205 589868
rect 481771 582452 481837 582453
rect 481771 582388 481772 582452
rect 481836 582388 481837 582452
rect 481771 582387 481837 582388
rect 481587 579596 481653 579597
rect 481587 579532 481588 579596
rect 481652 579532 481653 579596
rect 481587 579531 481653 579532
rect 481035 565180 481101 565181
rect 481035 565116 481036 565180
rect 481100 565116 481101 565180
rect 481035 565115 481101 565116
rect 480851 563820 480917 563821
rect 480851 563756 480852 563820
rect 480916 563756 480917 563820
rect 480851 563755 480917 563756
rect 482142 562461 482202 589867
rect 482323 588572 482389 588573
rect 482323 588508 482324 588572
rect 482388 588508 482389 588572
rect 482323 588507 482389 588508
rect 482326 564501 482386 588507
rect 483062 581637 483122 592995
rect 483611 592244 483677 592245
rect 483611 592180 483612 592244
rect 483676 592180 483677 592244
rect 483611 592179 483677 592180
rect 483059 581636 483125 581637
rect 483059 581572 483060 581636
rect 483124 581572 483125 581636
rect 483059 581571 483125 581572
rect 482875 579324 482941 579325
rect 482875 579260 482876 579324
rect 482940 579260 482941 579324
rect 482875 579259 482941 579260
rect 482507 578780 482573 578781
rect 482507 578716 482508 578780
rect 482572 578716 482573 578780
rect 482507 578715 482573 578716
rect 482510 565861 482570 578715
rect 482878 578101 482938 579259
rect 482875 578100 482941 578101
rect 482875 578036 482876 578100
rect 482940 578036 482941 578100
rect 482875 578035 482941 578036
rect 482507 565860 482573 565861
rect 482507 565796 482508 565860
rect 482572 565796 482573 565860
rect 482507 565795 482573 565796
rect 482323 564500 482389 564501
rect 482323 564436 482324 564500
rect 482388 564436 482389 564500
rect 482323 564435 482389 564436
rect 482139 562460 482205 562461
rect 482139 562396 482140 562460
rect 482204 562396 482205 562460
rect 482139 562395 482205 562396
rect 483614 559061 483674 592179
rect 483795 591428 483861 591429
rect 483795 591364 483796 591428
rect 483860 591364 483861 591428
rect 483795 591363 483861 591364
rect 483798 560421 483858 591363
rect 483979 589524 484045 589525
rect 483979 589460 483980 589524
rect 484044 589460 484045 589524
rect 483979 589459 484045 589460
rect 483982 563141 484042 589459
rect 486187 585988 486253 585989
rect 486187 585924 486188 585988
rect 486252 585924 486253 585988
rect 486187 585923 486253 585924
rect 485451 582588 485517 582589
rect 485451 582524 485452 582588
rect 485516 582524 485517 582588
rect 485451 582523 485517 582524
rect 485267 581908 485333 581909
rect 485267 581844 485268 581908
rect 485332 581844 485333 581908
rect 485267 581843 485333 581844
rect 485083 580684 485149 580685
rect 485083 580620 485084 580684
rect 485148 580620 485149 580684
rect 485083 580619 485149 580620
rect 485086 576061 485146 580619
rect 485083 576060 485149 576061
rect 485083 575996 485084 576060
rect 485148 575996 485149 576060
rect 485083 575995 485149 575996
rect 485270 574701 485330 581843
rect 485267 574700 485333 574701
rect 485267 574636 485268 574700
rect 485332 574636 485333 574700
rect 485267 574635 485333 574636
rect 485454 573341 485514 582523
rect 486003 582044 486069 582045
rect 486003 581980 486004 582044
rect 486068 581980 486069 582044
rect 486003 581979 486069 581980
rect 485819 581364 485885 581365
rect 485819 581300 485820 581364
rect 485884 581300 485885 581364
rect 485819 581299 485885 581300
rect 485635 580548 485701 580549
rect 485635 580484 485636 580548
rect 485700 580484 485701 580548
rect 485635 580483 485701 580484
rect 485638 576741 485698 580483
rect 485635 576740 485701 576741
rect 485635 576676 485636 576740
rect 485700 576676 485701 576740
rect 485635 576675 485701 576676
rect 485822 575381 485882 581299
rect 485819 575380 485885 575381
rect 485819 575316 485820 575380
rect 485884 575316 485885 575380
rect 485819 575315 485885 575316
rect 486006 574021 486066 581979
rect 486003 574020 486069 574021
rect 486003 573956 486004 574020
rect 486068 573956 486069 574020
rect 486003 573955 486069 573956
rect 485451 573340 485517 573341
rect 485451 573276 485452 573340
rect 485516 573276 485517 573340
rect 485451 573275 485517 573276
rect 486190 568170 486250 585923
rect 486371 585852 486437 585853
rect 486371 585788 486372 585852
rect 486436 585788 486437 585852
rect 486371 585787 486437 585788
rect 486374 568581 486434 585787
rect 486371 568580 486437 568581
rect 486371 568516 486372 568580
rect 486436 568516 486437 568580
rect 486371 568515 486437 568516
rect 486190 568110 486434 568170
rect 486374 567901 486434 568110
rect 486371 567900 486437 567901
rect 486371 567836 486372 567900
rect 486436 567836 486437 567900
rect 486371 567835 486437 567836
rect 483979 563140 484045 563141
rect 483979 563076 483980 563140
rect 484044 563076 484045 563140
rect 483979 563075 484045 563076
rect 483795 560420 483861 560421
rect 483795 560356 483796 560420
rect 483860 560356 483861 560420
rect 483795 560355 483861 560356
rect 483611 559060 483677 559061
rect 483611 558996 483612 559060
rect 483676 558996 483677 559060
rect 483611 558995 483677 558996
rect 480851 536620 480917 536621
rect 480851 536556 480852 536620
rect 480916 536556 480917 536620
rect 480851 536555 480917 536556
rect 478091 533900 478157 533901
rect 478091 533836 478092 533900
rect 478156 533836 478157 533900
rect 478091 533835 478157 533836
rect 477539 513364 477605 513365
rect 477539 513300 477540 513364
rect 477604 513300 477605 513364
rect 477539 513299 477605 513300
rect 477542 508469 477602 513299
rect 477539 508468 477605 508469
rect 477539 508404 477540 508468
rect 477604 508404 477605 508468
rect 477539 508403 477605 508404
rect 478094 508197 478154 533835
rect 478275 532540 478341 532541
rect 478275 532476 478276 532540
rect 478340 532476 478341 532540
rect 478275 532475 478341 532476
rect 478278 509013 478338 532475
rect 479563 529820 479629 529821
rect 479563 529756 479564 529820
rect 479628 529756 479629 529820
rect 479563 529755 479629 529756
rect 479379 526420 479445 526421
rect 479379 526356 479380 526420
rect 479444 526356 479445 526420
rect 479379 526355 479445 526356
rect 478459 516764 478525 516765
rect 478459 516700 478460 516764
rect 478524 516700 478525 516764
rect 478459 516699 478525 516700
rect 478462 511733 478522 516699
rect 479382 513093 479442 526355
rect 479566 518261 479626 529755
rect 479747 524380 479813 524381
rect 479747 524316 479748 524380
rect 479812 524316 479813 524380
rect 479747 524315 479813 524316
rect 479563 518260 479629 518261
rect 479563 518196 479564 518260
rect 479628 518196 479629 518260
rect 479563 518195 479629 518196
rect 479750 514453 479810 524315
rect 480667 523020 480733 523021
rect 480667 522956 480668 523020
rect 480732 522956 480733 523020
rect 480667 522955 480733 522956
rect 479931 518260 479997 518261
rect 479931 518196 479932 518260
rect 479996 518196 479997 518260
rect 479931 518195 479997 518196
rect 479747 514452 479813 514453
rect 479747 514388 479748 514452
rect 479812 514388 479813 514452
rect 479747 514387 479813 514388
rect 479934 513229 479994 518195
rect 480670 515269 480730 522955
rect 480667 515268 480733 515269
rect 480667 515204 480668 515268
rect 480732 515204 480733 515268
rect 480667 515203 480733 515204
rect 480483 514860 480549 514861
rect 480483 514796 480484 514860
rect 480548 514796 480549 514860
rect 480483 514795 480549 514796
rect 479931 513228 479997 513229
rect 479931 513164 479932 513228
rect 479996 513164 479997 513228
rect 479931 513163 479997 513164
rect 479379 513092 479445 513093
rect 479379 513028 479380 513092
rect 479444 513028 479445 513092
rect 479379 513027 479445 513028
rect 478827 512820 478893 512821
rect 478827 512756 478828 512820
rect 478892 512756 478893 512820
rect 478827 512755 478893 512756
rect 478643 511868 478709 511869
rect 478643 511804 478644 511868
rect 478708 511804 478709 511868
rect 478643 511803 478709 511804
rect 478459 511732 478525 511733
rect 478459 511668 478460 511732
rect 478524 511668 478525 511732
rect 478459 511667 478525 511668
rect 478275 509012 478341 509013
rect 478275 508948 478276 509012
rect 478340 508948 478341 509012
rect 478275 508947 478341 508948
rect 478091 508196 478157 508197
rect 478091 508132 478092 508196
rect 478156 508132 478157 508196
rect 478091 508131 478157 508132
rect 478646 507653 478706 511803
rect 478830 510645 478890 512755
rect 478827 510644 478893 510645
rect 478827 510580 478828 510644
rect 478892 510580 478893 510644
rect 478827 510579 478893 510580
rect 478643 507652 478709 507653
rect 478643 507588 478644 507652
rect 478708 507588 478709 507652
rect 478643 507587 478709 507588
rect 480486 504933 480546 514795
rect 480667 513364 480733 513365
rect 480667 513300 480668 513364
rect 480732 513300 480733 513364
rect 480667 513299 480733 513300
rect 480483 504932 480549 504933
rect 480483 504868 480484 504932
rect 480548 504868 480549 504932
rect 480483 504867 480549 504868
rect 480670 504117 480730 513299
rect 480854 506293 480914 536555
rect 482139 535260 482205 535261
rect 482139 535196 482140 535260
rect 482204 535196 482205 535260
rect 482139 535195 482205 535196
rect 481035 531180 481101 531181
rect 481035 531116 481036 531180
rect 481100 531116 481101 531180
rect 481035 531115 481101 531116
rect 481038 512005 481098 531115
rect 481219 527100 481285 527101
rect 481219 527036 481220 527100
rect 481284 527036 481285 527100
rect 481219 527035 481285 527036
rect 481222 512549 481282 527035
rect 481587 516220 481653 516221
rect 481587 516156 481588 516220
rect 481652 516156 481653 516220
rect 481587 516155 481653 516156
rect 481219 512548 481285 512549
rect 481219 512484 481220 512548
rect 481284 512484 481285 512548
rect 481219 512483 481285 512484
rect 481035 512004 481101 512005
rect 481035 511940 481036 512004
rect 481100 511940 481101 512004
rect 481035 511939 481101 511940
rect 481403 511460 481469 511461
rect 481403 511396 481404 511460
rect 481468 511396 481469 511460
rect 481403 511395 481469 511396
rect 481406 510101 481466 511395
rect 481403 510100 481469 510101
rect 481403 510036 481404 510100
rect 481468 510036 481469 510100
rect 481403 510035 481469 510036
rect 480851 506292 480917 506293
rect 480851 506228 480852 506292
rect 480916 506228 480917 506292
rect 480851 506227 480917 506228
rect 481590 505749 481650 516155
rect 481771 513772 481837 513773
rect 481771 513708 481772 513772
rect 481836 513708 481837 513772
rect 481771 513707 481837 513708
rect 481587 505748 481653 505749
rect 481587 505684 481588 505748
rect 481652 505684 481653 505748
rect 481587 505683 481653 505684
rect 481774 504389 481834 513707
rect 482142 507109 482202 535195
rect 483611 531860 483677 531861
rect 483611 531796 483612 531860
rect 483676 531796 483677 531860
rect 483611 531795 483677 531796
rect 483059 516356 483125 516357
rect 483059 516292 483060 516356
rect 483124 516292 483125 516356
rect 483059 516291 483125 516292
rect 482139 507108 482205 507109
rect 482139 507044 482140 507108
rect 482204 507044 482205 507108
rect 482139 507043 482205 507044
rect 483062 506837 483122 516291
rect 483427 515540 483493 515541
rect 483427 515476 483428 515540
rect 483492 515476 483493 515540
rect 483427 515475 483493 515476
rect 483243 514996 483309 514997
rect 483243 514932 483244 514996
rect 483308 514932 483309 514996
rect 483243 514931 483309 514932
rect 483059 506836 483125 506837
rect 483059 506772 483060 506836
rect 483124 506772 483125 506836
rect 483059 506771 483125 506772
rect 483246 505477 483306 514931
rect 483430 514181 483490 515475
rect 483427 514180 483493 514181
rect 483427 514116 483428 514180
rect 483492 514116 483493 514180
rect 483427 514115 483493 514116
rect 483614 509557 483674 531795
rect 485083 529140 485149 529141
rect 485083 529076 485084 529140
rect 485148 529076 485149 529140
rect 485083 529075 485149 529076
rect 483979 525740 484045 525741
rect 483979 525676 483980 525740
rect 484044 525676 484045 525740
rect 483979 525675 484045 525676
rect 483795 523700 483861 523701
rect 483795 523636 483796 523700
rect 483860 523636 483861 523700
rect 483795 523635 483861 523636
rect 483798 515133 483858 523635
rect 483982 517989 484042 525675
rect 484531 520980 484597 520981
rect 484531 520916 484532 520980
rect 484596 520916 484597 520980
rect 484531 520915 484597 520916
rect 484347 519620 484413 519621
rect 484347 519556 484348 519620
rect 484412 519556 484413 519620
rect 484347 519555 484413 519556
rect 483979 517988 484045 517989
rect 483979 517924 483980 517988
rect 484044 517924 484045 517988
rect 483979 517923 484045 517924
rect 484350 517717 484410 519555
rect 484347 517716 484413 517717
rect 484347 517652 484348 517716
rect 484412 517652 484413 517716
rect 484347 517651 484413 517652
rect 484534 516629 484594 520915
rect 484715 520300 484781 520301
rect 484715 520236 484716 520300
rect 484780 520236 484781 520300
rect 484715 520235 484781 520236
rect 484718 517173 484778 520235
rect 484899 518940 484965 518941
rect 484899 518876 484900 518940
rect 484964 518876 484965 518940
rect 484899 518875 484965 518876
rect 484715 517172 484781 517173
rect 484715 517108 484716 517172
rect 484780 517108 484781 517172
rect 484715 517107 484781 517108
rect 484531 516628 484597 516629
rect 484531 516564 484532 516628
rect 484596 516564 484597 516628
rect 484531 516563 484597 516564
rect 484902 515677 484962 518875
rect 484899 515676 484965 515677
rect 484899 515612 484900 515676
rect 484964 515612 484965 515676
rect 484899 515611 484965 515612
rect 483795 515132 483861 515133
rect 483795 515068 483796 515132
rect 483860 515068 483861 515132
rect 483795 515067 483861 515068
rect 484347 514180 484413 514181
rect 484347 514116 484348 514180
rect 484412 514116 484413 514180
rect 484347 514115 484413 514116
rect 484350 512957 484410 514115
rect 485086 513637 485146 529075
rect 486371 528460 486437 528461
rect 486371 528396 486372 528460
rect 486436 528396 486437 528460
rect 486371 528395 486437 528396
rect 485267 527780 485333 527781
rect 485267 527716 485268 527780
rect 485332 527716 485333 527780
rect 485267 527715 485333 527716
rect 485083 513636 485149 513637
rect 485083 513572 485084 513636
rect 485148 513572 485149 513636
rect 485083 513571 485149 513572
rect 484531 513500 484597 513501
rect 484531 513436 484532 513500
rect 484596 513436 484597 513500
rect 484531 513435 484597 513436
rect 484347 512956 484413 512957
rect 484347 512892 484348 512956
rect 484412 512892 484413 512956
rect 484347 512891 484413 512892
rect 484347 512140 484413 512141
rect 484347 512076 484348 512140
rect 484412 512076 484413 512140
rect 484347 512075 484413 512076
rect 484350 511189 484410 512075
rect 484347 511188 484413 511189
rect 484347 511124 484348 511188
rect 484412 511124 484413 511188
rect 484347 511123 484413 511124
rect 484534 510917 484594 513435
rect 485270 512277 485330 527715
rect 486003 525060 486069 525061
rect 486003 524996 486004 525060
rect 486068 524996 486069 525060
rect 486003 524995 486069 524996
rect 485819 521660 485885 521661
rect 485819 521596 485820 521660
rect 485884 521596 485885 521660
rect 485819 521595 485885 521596
rect 485822 518910 485882 521595
rect 485638 518850 485882 518910
rect 485267 512276 485333 512277
rect 485267 512212 485268 512276
rect 485332 512212 485333 512276
rect 485267 512211 485333 512212
rect 485638 511597 485698 518850
rect 486006 518530 486066 524995
rect 486374 523970 486434 528395
rect 485822 518470 486066 518530
rect 486190 523910 486434 523970
rect 485822 513909 485882 518470
rect 486190 517850 486250 523910
rect 486371 522340 486437 522341
rect 486371 522276 486372 522340
rect 486436 522276 486437 522340
rect 486371 522275 486437 522276
rect 486006 517790 486250 517850
rect 486006 515813 486066 517790
rect 486187 517308 486253 517309
rect 486187 517244 486188 517308
rect 486252 517244 486253 517308
rect 486187 517243 486253 517244
rect 486190 517170 486250 517243
rect 486374 517170 486434 522275
rect 486190 517110 486434 517170
rect 486003 515812 486069 515813
rect 486003 515748 486004 515812
rect 486068 515748 486069 515812
rect 486003 515747 486069 515748
rect 485819 513908 485885 513909
rect 485819 513844 485820 513908
rect 485884 513844 485885 513908
rect 485819 513843 485885 513844
rect 485635 511596 485701 511597
rect 485635 511532 485636 511596
rect 485700 511532 485701 511596
rect 485635 511531 485701 511532
rect 484531 510916 484597 510917
rect 484531 510852 484532 510916
rect 484596 510852 484597 510916
rect 484531 510851 484597 510852
rect 483611 509556 483677 509557
rect 483611 509492 483612 509556
rect 483676 509492 483677 509556
rect 483611 509491 483677 509492
rect 483243 505476 483309 505477
rect 483243 505412 483244 505476
rect 483308 505412 483309 505476
rect 483243 505411 483309 505412
rect 481771 504388 481837 504389
rect 481771 504324 481772 504388
rect 481836 504324 481837 504388
rect 481771 504323 481837 504324
rect 480667 504116 480733 504117
rect 480667 504052 480668 504116
rect 480732 504052 480733 504116
rect 480667 504051 480733 504052
rect 483059 503300 483125 503301
rect 483059 503236 483060 503300
rect 483124 503236 483125 503300
rect 483059 503235 483125 503236
rect 481771 502892 481837 502893
rect 481771 502828 481772 502892
rect 481836 502828 481837 502892
rect 481771 502827 481837 502828
rect 477539 502484 477605 502485
rect 477539 502420 477540 502484
rect 477604 502420 477605 502484
rect 477539 502419 477605 502420
rect 477542 492693 477602 502419
rect 480667 501804 480733 501805
rect 480667 501740 480668 501804
rect 480732 501740 480733 501804
rect 480667 501739 480733 501740
rect 480299 497452 480365 497453
rect 480299 497388 480300 497452
rect 480364 497388 480365 497452
rect 480299 497387 480365 497388
rect 480115 496908 480181 496909
rect 480115 496844 480116 496908
rect 480180 496844 480181 496908
rect 480115 496843 480181 496844
rect 479563 496364 479629 496365
rect 479563 496300 479564 496364
rect 479628 496300 479629 496364
rect 479563 496299 479629 496300
rect 478091 495548 478157 495549
rect 478091 495484 478092 495548
rect 478156 495484 478157 495548
rect 478091 495483 478157 495484
rect 477539 492692 477605 492693
rect 477539 492628 477540 492692
rect 477604 492628 477605 492692
rect 477539 492627 477605 492628
rect 477355 490170 477421 490171
rect 477355 490106 477356 490170
rect 477420 490106 477421 490170
rect 477355 490105 477421 490106
rect 477358 486981 477418 490105
rect 477355 486980 477421 486981
rect 477355 486916 477356 486980
rect 477420 486916 477421 486980
rect 477355 486915 477421 486916
rect 478094 478821 478154 495483
rect 478275 495004 478341 495005
rect 478275 494940 478276 495004
rect 478340 494940 478341 495004
rect 478275 494939 478341 494940
rect 478278 479501 478338 494939
rect 478459 492828 478525 492829
rect 478459 492764 478460 492828
rect 478524 492764 478525 492828
rect 478459 492763 478525 492764
rect 478462 482901 478522 492763
rect 478827 492284 478893 492285
rect 478827 492220 478828 492284
rect 478892 492220 478893 492284
rect 478827 492219 478893 492220
rect 478830 483581 478890 492219
rect 479566 491197 479626 496299
rect 480118 494325 480178 496843
rect 480115 494324 480181 494325
rect 480115 494260 480116 494324
rect 480180 494260 480181 494324
rect 480115 494259 480181 494260
rect 479563 491196 479629 491197
rect 479563 491132 479564 491196
rect 479628 491132 479629 491196
rect 479563 491131 479629 491132
rect 480302 488613 480362 497387
rect 480670 496909 480730 501739
rect 481587 500988 481653 500989
rect 481587 500924 481588 500988
rect 481652 500924 481653 500988
rect 481587 500923 481653 500924
rect 480851 500444 480917 500445
rect 480851 500380 480852 500444
rect 480916 500380 480917 500444
rect 480851 500379 480917 500380
rect 480667 496908 480733 496909
rect 480667 496844 480668 496908
rect 480732 496844 480733 496908
rect 480667 496843 480733 496844
rect 480299 488612 480365 488613
rect 480299 488548 480300 488612
rect 480364 488548 480365 488612
rect 480299 488547 480365 488548
rect 478827 483580 478893 483581
rect 478827 483516 478828 483580
rect 478892 483516 478893 483580
rect 478827 483515 478893 483516
rect 478459 482900 478525 482901
rect 478459 482836 478460 482900
rect 478524 482836 478525 482900
rect 478459 482835 478525 482836
rect 478275 479500 478341 479501
rect 478275 479436 478276 479500
rect 478340 479436 478341 479500
rect 478275 479435 478341 479436
rect 478091 478820 478157 478821
rect 478091 478756 478092 478820
rect 478156 478756 478157 478820
rect 478091 478755 478157 478756
rect 480854 471341 480914 500379
rect 481035 499084 481101 499085
rect 481035 499020 481036 499084
rect 481100 499020 481101 499084
rect 481035 499019 481101 499020
rect 481038 473381 481098 499019
rect 481219 497724 481285 497725
rect 481219 497660 481220 497724
rect 481284 497660 481285 497724
rect 481219 497659 481285 497660
rect 481222 475421 481282 497659
rect 481590 492693 481650 500923
rect 481774 494733 481834 502827
rect 482139 499628 482205 499629
rect 482139 499564 482140 499628
rect 482204 499564 482205 499628
rect 482139 499563 482205 499564
rect 481771 494732 481837 494733
rect 481771 494668 481772 494732
rect 481836 494668 481837 494732
rect 481771 494667 481837 494668
rect 481587 492692 481653 492693
rect 481587 492628 481588 492692
rect 481652 492628 481653 492692
rect 481587 492627 481653 492628
rect 481955 492012 482021 492013
rect 481955 491948 481956 492012
rect 482020 491948 482021 492012
rect 481955 491947 482021 491948
rect 481771 491604 481837 491605
rect 481771 491540 481772 491604
rect 481836 491540 481837 491604
rect 481771 491539 481837 491540
rect 481774 484941 481834 491539
rect 481771 484940 481837 484941
rect 481771 484876 481772 484940
rect 481836 484876 481837 484940
rect 481771 484875 481837 484876
rect 481958 484261 482018 491947
rect 481955 484260 482021 484261
rect 481955 484196 481956 484260
rect 482020 484196 482021 484260
rect 481955 484195 482021 484196
rect 481219 475420 481285 475421
rect 481219 475356 481220 475420
rect 481284 475356 481285 475420
rect 481219 475355 481285 475356
rect 481035 473380 481101 473381
rect 481035 473316 481036 473380
rect 481100 473316 481101 473380
rect 481035 473315 481101 473316
rect 482142 472701 482202 499563
rect 482323 498268 482389 498269
rect 482323 498204 482324 498268
rect 482388 498204 482389 498268
rect 482323 498203 482389 498204
rect 482326 474741 482386 498203
rect 483062 494733 483122 503235
rect 483427 501668 483493 501669
rect 483427 501604 483428 501668
rect 483492 501604 483493 501668
rect 483427 501603 483493 501604
rect 483059 494732 483125 494733
rect 483059 494668 483060 494732
rect 483124 494668 483125 494732
rect 483059 494667 483125 494668
rect 483430 494053 483490 501603
rect 483611 500308 483677 500309
rect 483611 500244 483612 500308
rect 483676 500244 483677 500308
rect 483611 500243 483677 500244
rect 483427 494052 483493 494053
rect 483427 493988 483428 494052
rect 483492 493988 483493 494052
rect 483427 493987 483493 493988
rect 483243 489428 483309 489429
rect 483243 489364 483244 489428
rect 483308 489364 483309 489428
rect 483243 489363 483309 489364
rect 483246 488341 483306 489363
rect 483243 488340 483309 488341
rect 483243 488276 483244 488340
rect 483308 488276 483309 488340
rect 483243 488275 483309 488276
rect 482323 474740 482389 474741
rect 482323 474676 482324 474740
rect 482388 474676 482389 474740
rect 482323 474675 482389 474676
rect 482139 472700 482205 472701
rect 482139 472636 482140 472700
rect 482204 472636 482205 472700
rect 482139 472635 482205 472636
rect 483614 472021 483674 500243
rect 483795 498948 483861 498949
rect 483795 498884 483796 498948
rect 483860 498884 483861 498948
rect 483795 498883 483861 498884
rect 483798 474061 483858 498883
rect 486003 494868 486069 494869
rect 486003 494804 486004 494868
rect 486068 494804 486069 494868
rect 486003 494803 486069 494804
rect 483979 493508 484045 493509
rect 483979 493444 483980 493508
rect 484044 493444 484045 493508
rect 483979 493443 484045 493444
rect 483982 482221 484042 493443
rect 484899 490924 484965 490925
rect 484899 490860 484900 490924
rect 484964 490860 484965 490924
rect 484899 490859 484965 490860
rect 484531 490788 484597 490789
rect 484531 490724 484532 490788
rect 484596 490724 484597 490788
rect 484531 490723 484597 490724
rect 484347 489564 484413 489565
rect 484347 489500 484348 489564
rect 484412 489500 484413 489564
rect 484347 489499 484413 489500
rect 484350 487661 484410 489499
rect 484347 487660 484413 487661
rect 484347 487596 484348 487660
rect 484412 487596 484413 487660
rect 484347 487595 484413 487596
rect 484534 486301 484594 490723
rect 484531 486300 484597 486301
rect 484531 486236 484532 486300
rect 484596 486236 484597 486300
rect 484531 486235 484597 486236
rect 484902 485621 484962 490859
rect 485451 488748 485517 488749
rect 485451 488684 485452 488748
rect 485516 488684 485517 488748
rect 485451 488683 485517 488684
rect 484899 485620 484965 485621
rect 484899 485556 484900 485620
rect 484964 485556 484965 485620
rect 484899 485555 484965 485556
rect 483979 482220 484045 482221
rect 483979 482156 483980 482220
rect 484044 482156 484045 482220
rect 483979 482155 484045 482156
rect 485454 476101 485514 488683
rect 486006 480181 486066 494803
rect 486187 494188 486253 494189
rect 486187 494124 486188 494188
rect 486252 494124 486253 494188
rect 486187 494123 486253 494124
rect 486190 489930 486250 494123
rect 486190 489870 486434 489930
rect 486374 480861 486434 489870
rect 486371 480860 486437 480861
rect 486371 480796 486372 480860
rect 486436 480796 486437 480860
rect 486371 480795 486437 480796
rect 486003 480180 486069 480181
rect 486003 480116 486004 480180
rect 486068 480116 486069 480180
rect 486003 480115 486069 480116
rect 485451 476100 485517 476101
rect 485451 476036 485452 476100
rect 485516 476036 485517 476100
rect 485451 476035 485517 476036
rect 483795 474060 483861 474061
rect 483795 473996 483796 474060
rect 483860 473996 483861 474060
rect 483795 473995 483861 473996
rect 483611 472020 483677 472021
rect 483611 471956 483612 472020
rect 483676 471956 483677 472020
rect 483611 471955 483677 471956
rect 480851 471340 480917 471341
rect 480851 471276 480852 471340
rect 480916 471276 480917 471340
rect 480851 471275 480917 471276
rect 483611 452980 483677 452981
rect 483611 452916 483612 452980
rect 483676 452916 483677 452980
rect 483611 452915 483677 452916
rect 478091 447540 478157 447541
rect 478091 447476 478092 447540
rect 478156 447476 478157 447540
rect 478091 447475 478157 447476
rect 477355 432580 477421 432581
rect 477355 432516 477356 432580
rect 477420 432516 477421 432580
rect 477355 432515 477421 432516
rect 477358 425523 477418 432515
rect 477539 427276 477605 427277
rect 477539 427212 477540 427276
rect 477604 427212 477605 427276
rect 477539 427211 477605 427212
rect 477355 425522 477421 425523
rect 477355 425458 477356 425522
rect 477420 425458 477421 425522
rect 477355 425457 477421 425458
rect 477542 414357 477602 427211
rect 477907 421020 477973 421021
rect 477907 420956 477908 421020
rect 477972 420956 477973 421020
rect 477907 420955 477973 420956
rect 477539 414356 477605 414357
rect 477539 414292 477540 414356
rect 477604 414292 477605 414356
rect 477539 414291 477605 414292
rect 477910 413269 477970 420955
rect 478094 415717 478154 447475
rect 479379 443460 479445 443461
rect 479379 443396 479380 443460
rect 479444 443396 479445 443460
rect 479379 443395 479445 443396
rect 478275 442100 478341 442101
rect 478275 442036 478276 442100
rect 478340 442036 478341 442100
rect 478275 442035 478341 442036
rect 478278 419253 478338 442035
rect 478643 441420 478709 441421
rect 478643 441356 478644 441420
rect 478708 441356 478709 441420
rect 478643 441355 478709 441356
rect 478646 421973 478706 441355
rect 478643 421972 478709 421973
rect 478643 421908 478644 421972
rect 478708 421908 478709 421972
rect 478643 421907 478709 421908
rect 478275 419252 478341 419253
rect 478275 419188 478276 419252
rect 478340 419188 478341 419252
rect 478275 419187 478341 419188
rect 479382 418437 479442 443395
rect 479563 442780 479629 442781
rect 479563 442716 479564 442780
rect 479628 442716 479629 442780
rect 479563 442715 479629 442716
rect 479566 418709 479626 442715
rect 482139 440740 482205 440741
rect 482139 440676 482140 440740
rect 482204 440676 482205 440740
rect 482139 440675 482205 440676
rect 480851 440060 480917 440061
rect 480851 439996 480852 440060
rect 480916 439996 480917 440060
rect 480851 439995 480917 439996
rect 480115 433260 480181 433261
rect 480115 433196 480116 433260
rect 480180 433196 480181 433260
rect 480115 433195 480181 433196
rect 479931 427276 479997 427277
rect 479931 427212 479932 427276
rect 479996 427212 479997 427276
rect 479931 427211 479997 427212
rect 479747 424556 479813 424557
rect 479747 424492 479748 424556
rect 479812 424492 479813 424556
rect 479747 424491 479813 424492
rect 479563 418708 479629 418709
rect 479563 418644 479564 418708
rect 479628 418644 479629 418708
rect 479563 418643 479629 418644
rect 479379 418436 479445 418437
rect 479379 418372 479380 418436
rect 479444 418372 479445 418436
rect 479379 418371 479445 418372
rect 478275 418300 478341 418301
rect 478275 418236 478276 418300
rect 478340 418236 478341 418300
rect 478275 418235 478341 418236
rect 478091 415716 478157 415717
rect 478091 415652 478092 415716
rect 478156 415652 478157 415716
rect 478091 415651 478157 415652
rect 478278 413813 478338 418235
rect 479750 417077 479810 424491
rect 479934 417893 479994 427211
rect 480118 425237 480178 433195
rect 480854 425781 480914 439995
rect 481587 431220 481653 431221
rect 481587 431156 481588 431220
rect 481652 431156 481653 431220
rect 481587 431155 481653 431156
rect 481590 426597 481650 431155
rect 481587 426596 481653 426597
rect 481587 426532 481588 426596
rect 481652 426532 481653 426596
rect 481587 426531 481653 426532
rect 481955 426188 482021 426189
rect 481955 426124 481956 426188
rect 482020 426124 482021 426188
rect 481955 426123 482021 426124
rect 480851 425780 480917 425781
rect 480851 425716 480852 425780
rect 480916 425716 480917 425780
rect 480851 425715 480917 425716
rect 480115 425236 480181 425237
rect 480115 425172 480116 425236
rect 480180 425172 480181 425236
rect 480115 425171 480181 425172
rect 481219 423604 481285 423605
rect 481219 423540 481220 423604
rect 481284 423540 481285 423604
rect 481219 423539 481285 423540
rect 480851 423060 480917 423061
rect 480851 422996 480852 423060
rect 480916 422996 480917 423060
rect 480851 422995 480917 422996
rect 480115 419524 480181 419525
rect 480115 419460 480116 419524
rect 480180 419460 480181 419524
rect 480115 419459 480181 419460
rect 479931 417892 479997 417893
rect 479931 417828 479932 417892
rect 479996 417828 479997 417892
rect 479931 417827 479997 417828
rect 479747 417076 479813 417077
rect 479747 417012 479748 417076
rect 479812 417012 479813 417076
rect 479747 417011 479813 417012
rect 478643 416668 478709 416669
rect 478643 416604 478644 416668
rect 478708 416604 478709 416668
rect 478643 416603 478709 416604
rect 478459 415308 478525 415309
rect 478459 415244 478460 415308
rect 478524 415244 478525 415308
rect 478459 415243 478525 415244
rect 478275 413812 478341 413813
rect 478275 413748 478276 413812
rect 478340 413748 478341 413812
rect 478275 413747 478341 413748
rect 477907 413268 477973 413269
rect 477907 413204 477908 413268
rect 477972 413204 477973 413268
rect 477907 413203 477973 413204
rect 478462 410549 478522 415243
rect 478646 412997 478706 416603
rect 480118 416533 480178 419459
rect 480115 416532 480181 416533
rect 480115 416468 480116 416532
rect 480180 416468 480181 416532
rect 480115 416467 480181 416468
rect 479931 414220 479997 414221
rect 479931 414156 479932 414220
rect 479996 414156 479997 414220
rect 479931 414155 479997 414156
rect 478643 412996 478709 412997
rect 478643 412932 478644 412996
rect 478708 412932 478709 412996
rect 478643 412931 478709 412932
rect 479934 411637 479994 414155
rect 480299 412860 480365 412861
rect 480299 412796 480300 412860
rect 480364 412796 480365 412860
rect 480299 412795 480365 412796
rect 480302 411909 480362 412795
rect 480854 412181 480914 422995
rect 481222 420069 481282 423539
rect 481958 422310 482018 426123
rect 481774 422250 482018 422310
rect 481219 420068 481285 420069
rect 481219 420004 481220 420068
rect 481284 420004 481285 420068
rect 481219 420003 481285 420004
rect 481403 419932 481469 419933
rect 481403 419868 481404 419932
rect 481468 419868 481469 419932
rect 481403 419867 481469 419868
rect 481406 413541 481466 419867
rect 481587 419796 481653 419797
rect 481587 419732 481588 419796
rect 481652 419732 481653 419796
rect 481587 419731 481653 419732
rect 481403 413540 481469 413541
rect 481403 413476 481404 413540
rect 481468 413476 481469 413540
rect 481403 413475 481469 413476
rect 480851 412180 480917 412181
rect 480851 412116 480852 412180
rect 480916 412116 480917 412180
rect 480851 412115 480917 412116
rect 480299 411908 480365 411909
rect 480299 411844 480300 411908
rect 480364 411844 480365 411908
rect 480299 411843 480365 411844
rect 479931 411636 479997 411637
rect 479931 411572 479932 411636
rect 479996 411572 479997 411636
rect 479931 411571 479997 411572
rect 478459 410548 478525 410549
rect 478459 410484 478460 410548
rect 478524 410484 478525 410548
rect 478459 410483 478525 410484
rect 481590 409733 481650 419731
rect 481774 415989 481834 422250
rect 482142 420477 482202 440675
rect 483243 430540 483309 430541
rect 483243 430476 483244 430540
rect 483308 430476 483309 430540
rect 483243 430475 483309 430476
rect 483059 429180 483125 429181
rect 483059 429116 483060 429180
rect 483124 429116 483125 429180
rect 483059 429115 483125 429116
rect 482507 426188 482573 426189
rect 482507 426124 482508 426188
rect 482572 426124 482573 426188
rect 482507 426123 482573 426124
rect 482139 420476 482205 420477
rect 482139 420412 482140 420476
rect 482204 420412 482205 420476
rect 482139 420411 482205 420412
rect 481955 419660 482021 419661
rect 481955 419596 481956 419660
rect 482020 419596 482021 419660
rect 481955 419595 482021 419596
rect 481771 415988 481837 415989
rect 481771 415924 481772 415988
rect 481836 415924 481837 415988
rect 481771 415923 481837 415924
rect 481587 409732 481653 409733
rect 481587 409668 481588 409732
rect 481652 409668 481653 409732
rect 481587 409667 481653 409668
rect 481958 408917 482018 419595
rect 482323 416668 482389 416669
rect 482323 416604 482324 416668
rect 482388 416604 482389 416668
rect 482323 416603 482389 416604
rect 481955 408916 482021 408917
rect 481955 408852 481956 408916
rect 482020 408852 482021 408916
rect 481955 408851 482021 408852
rect 482326 407557 482386 416603
rect 482510 414629 482570 426123
rect 482875 425100 482941 425101
rect 482875 425036 482876 425100
rect 482940 425036 482941 425100
rect 482875 425035 482941 425036
rect 482878 423469 482938 425035
rect 482875 423468 482941 423469
rect 482875 423404 482876 423468
rect 482940 423404 482941 423468
rect 482875 423403 482941 423404
rect 483062 423333 483122 429115
rect 483246 426869 483306 430475
rect 483243 426868 483309 426869
rect 483243 426804 483244 426868
rect 483308 426804 483309 426868
rect 483243 426803 483309 426804
rect 483243 424964 483309 424965
rect 483243 424900 483244 424964
rect 483308 424900 483309 424964
rect 483243 424899 483309 424900
rect 483059 423332 483125 423333
rect 483059 423268 483060 423332
rect 483124 423268 483125 423332
rect 483059 423267 483125 423268
rect 483246 422310 483306 424899
rect 483614 424693 483674 452915
rect 485635 439380 485701 439381
rect 485635 439316 485636 439380
rect 485700 439316 485701 439380
rect 485635 439315 485701 439316
rect 483795 438700 483861 438701
rect 483795 438636 483796 438700
rect 483860 438636 483861 438700
rect 483795 438635 483861 438636
rect 483611 424692 483677 424693
rect 483611 424628 483612 424692
rect 483676 424628 483677 424692
rect 483611 424627 483677 424628
rect 483427 423604 483493 423605
rect 483427 423540 483428 423604
rect 483492 423540 483493 423604
rect 483427 423539 483493 423540
rect 483062 422250 483306 422310
rect 483062 417210 483122 422250
rect 483243 418300 483309 418301
rect 483243 418236 483244 418300
rect 483308 418236 483309 418300
rect 483243 418235 483309 418236
rect 482878 417150 483122 417210
rect 482878 415173 482938 417150
rect 483246 416805 483306 418235
rect 483243 416804 483309 416805
rect 483243 416740 483244 416804
rect 483308 416740 483309 416804
rect 483243 416739 483309 416740
rect 483059 416668 483125 416669
rect 483059 416604 483060 416668
rect 483124 416604 483125 416668
rect 483059 416603 483125 416604
rect 482875 415172 482941 415173
rect 482875 415108 482876 415172
rect 482940 415108 482941 415172
rect 482875 415107 482941 415108
rect 482507 414628 482573 414629
rect 482507 414564 482508 414628
rect 482572 414564 482573 414628
rect 482507 414563 482573 414564
rect 482875 410140 482941 410141
rect 482875 410076 482876 410140
rect 482940 410076 482941 410140
rect 482875 410075 482941 410076
rect 482878 408645 482938 410075
rect 483062 409189 483122 416603
rect 483430 410277 483490 423539
rect 483798 416261 483858 438635
rect 485267 437340 485333 437341
rect 485267 437276 485268 437340
rect 485332 437276 485333 437340
rect 485267 437275 485333 437276
rect 485083 435980 485149 435981
rect 485083 435916 485084 435980
rect 485148 435916 485149 435980
rect 485083 435915 485149 435916
rect 484531 434620 484597 434621
rect 484531 434556 484532 434620
rect 484596 434556 484597 434620
rect 484531 434555 484597 434556
rect 484347 429860 484413 429861
rect 484347 429796 484348 429860
rect 484412 429796 484413 429860
rect 484347 429795 484413 429796
rect 484350 427413 484410 429795
rect 484534 428229 484594 434555
rect 484715 431900 484781 431901
rect 484715 431836 484716 431900
rect 484780 431836 484781 431900
rect 484715 431835 484781 431836
rect 484531 428228 484597 428229
rect 484531 428164 484532 428228
rect 484596 428164 484597 428228
rect 484531 428163 484597 428164
rect 484347 427412 484413 427413
rect 484347 427348 484348 427412
rect 484412 427348 484413 427412
rect 484347 427347 484413 427348
rect 484718 426053 484778 431835
rect 484899 428500 484965 428501
rect 484899 428436 484900 428500
rect 484964 428436 484965 428500
rect 484899 428435 484965 428436
rect 484715 426052 484781 426053
rect 484715 425988 484716 426052
rect 484780 425988 484781 426052
rect 484715 425987 484781 425988
rect 484347 424420 484413 424421
rect 484347 424356 484348 424420
rect 484412 424356 484413 424420
rect 484347 424355 484413 424356
rect 484350 422245 484410 424355
rect 484531 423740 484597 423741
rect 484531 423676 484532 423740
rect 484596 423676 484597 423740
rect 484531 423675 484597 423676
rect 484347 422244 484413 422245
rect 484347 422180 484348 422244
rect 484412 422180 484413 422244
rect 484347 422179 484413 422180
rect 484534 419389 484594 423675
rect 484715 422380 484781 422381
rect 484715 422316 484716 422380
rect 484780 422316 484781 422380
rect 484715 422315 484781 422316
rect 484718 421293 484778 422315
rect 484715 421292 484781 421293
rect 484715 421228 484716 421292
rect 484780 421228 484781 421292
rect 484715 421227 484781 421228
rect 484902 420069 484962 428435
rect 485086 423197 485146 435915
rect 485083 423196 485149 423197
rect 485083 423132 485084 423196
rect 485148 423132 485149 423196
rect 485083 423131 485149 423132
rect 485270 422517 485330 437275
rect 485638 427957 485698 439315
rect 486371 436660 486437 436661
rect 486371 436596 486372 436660
rect 486436 436596 486437 436660
rect 486371 436595 486437 436596
rect 485819 435300 485885 435301
rect 485819 435236 485820 435300
rect 485884 435236 485885 435300
rect 485819 435235 485885 435236
rect 485635 427956 485701 427957
rect 485635 427892 485636 427956
rect 485700 427892 485701 427956
rect 485635 427891 485701 427892
rect 485822 423877 485882 435235
rect 486003 433940 486069 433941
rect 486003 433876 486004 433940
rect 486068 433876 486069 433940
rect 486003 433875 486069 433876
rect 485819 423876 485885 423877
rect 485819 423812 485820 423876
rect 485884 423812 485885 423876
rect 485819 423811 485885 423812
rect 485267 422516 485333 422517
rect 485267 422452 485268 422516
rect 485332 422452 485333 422516
rect 485267 422451 485333 422452
rect 486006 421837 486066 433875
rect 486374 431970 486434 436595
rect 486190 431910 486434 431970
rect 486190 422789 486250 431910
rect 486371 425780 486437 425781
rect 486371 425716 486372 425780
rect 486436 425716 486437 425780
rect 486371 425715 486437 425716
rect 486374 424829 486434 425715
rect 486371 424828 486437 424829
rect 486371 424764 486372 424828
rect 486436 424764 486437 424828
rect 486371 424763 486437 424764
rect 486187 422788 486253 422789
rect 486187 422724 486188 422788
rect 486252 422724 486253 422788
rect 486187 422723 486253 422724
rect 486003 421836 486069 421837
rect 486003 421772 486004 421836
rect 486068 421772 486069 421836
rect 486003 421771 486069 421772
rect 485819 420340 485885 420341
rect 485819 420276 485820 420340
rect 485884 420276 485885 420340
rect 485819 420275 485885 420276
rect 484899 420068 484965 420069
rect 484899 420004 484900 420068
rect 484964 420004 484965 420068
rect 484899 420003 484965 420004
rect 484531 419388 484597 419389
rect 484531 419324 484532 419388
rect 484596 419324 484597 419388
rect 484531 419323 484597 419324
rect 484347 416940 484413 416941
rect 484347 416876 484348 416940
rect 484412 416876 484413 416940
rect 484347 416875 484413 416876
rect 483795 416260 483861 416261
rect 483795 416196 483796 416260
rect 483860 416196 483861 416260
rect 483795 416195 483861 416196
rect 484350 415445 484410 416875
rect 484531 416260 484597 416261
rect 484531 416196 484532 416260
rect 484596 416196 484597 416260
rect 484531 416195 484597 416196
rect 484347 415444 484413 415445
rect 484347 415380 484348 415444
rect 484412 415380 484413 415444
rect 484347 415379 484413 415380
rect 483611 415308 483677 415309
rect 483611 415244 483612 415308
rect 483676 415244 483677 415308
rect 483611 415243 483677 415244
rect 483427 410276 483493 410277
rect 483427 410212 483428 410276
rect 483492 410212 483493 410276
rect 483427 410211 483493 410212
rect 483059 409188 483125 409189
rect 483059 409124 483060 409188
rect 483124 409124 483125 409188
rect 483059 409123 483125 409124
rect 482875 408644 482941 408645
rect 482875 408580 482876 408644
rect 482940 408580 482941 408644
rect 482875 408579 482941 408580
rect 483614 408373 483674 415243
rect 484534 414085 484594 416195
rect 484715 415580 484781 415581
rect 484715 415516 484716 415580
rect 484780 415516 484781 415580
rect 484715 415515 484781 415516
rect 484531 414084 484597 414085
rect 484531 414020 484532 414084
rect 484596 414020 484597 414084
rect 484531 414019 484597 414020
rect 484163 413540 484229 413541
rect 484163 413476 484164 413540
rect 484228 413476 484229 413540
rect 484163 413475 484229 413476
rect 484166 411365 484226 413475
rect 484718 412725 484778 415515
rect 484715 412724 484781 412725
rect 484715 412660 484716 412724
rect 484780 412660 484781 412724
rect 484715 412659 484781 412660
rect 485822 412453 485882 420275
rect 485819 412452 485885 412453
rect 485819 412388 485820 412452
rect 485884 412388 485885 412452
rect 485819 412387 485885 412388
rect 484347 412180 484413 412181
rect 484347 412116 484348 412180
rect 484412 412116 484413 412180
rect 484347 412115 484413 412116
rect 484163 411364 484229 411365
rect 484163 411300 484164 411364
rect 484228 411300 484229 411364
rect 484163 411299 484229 411300
rect 484350 411093 484410 412115
rect 484531 411500 484597 411501
rect 484531 411436 484532 411500
rect 484596 411436 484597 411500
rect 484531 411435 484597 411436
rect 484347 411092 484413 411093
rect 484347 411028 484348 411092
rect 484412 411028 484413 411092
rect 484347 411027 484413 411028
rect 484534 410005 484594 411435
rect 484531 410004 484597 410005
rect 484531 409940 484532 410004
rect 484596 409940 484597 410004
rect 484531 409939 484597 409940
rect 484347 408780 484413 408781
rect 484347 408716 484348 408780
rect 484412 408716 484413 408780
rect 484347 408715 484413 408716
rect 483611 408372 483677 408373
rect 483611 408308 483612 408372
rect 483676 408308 483677 408372
rect 483611 408307 483677 408308
rect 484350 407829 484410 408715
rect 484347 407828 484413 407829
rect 484347 407764 484348 407828
rect 484412 407764 484413 407828
rect 484347 407763 484413 407764
rect 482323 407556 482389 407557
rect 482323 407492 482324 407556
rect 482388 407492 482389 407556
rect 482323 407491 482389 407492
rect 477539 406604 477605 406605
rect 477539 406540 477540 406604
rect 477604 406540 477605 406604
rect 477539 406539 477605 406540
rect 477355 401776 477421 401777
rect 477355 401712 477356 401776
rect 477420 401712 477421 401776
rect 477355 401711 477421 401712
rect 477358 394501 477418 401711
rect 477542 399533 477602 406539
rect 477723 406468 477789 406469
rect 477723 406404 477724 406468
rect 477788 406404 477789 406468
rect 477723 406403 477789 406404
rect 477539 399532 477605 399533
rect 477539 399468 477540 399532
rect 477604 399468 477605 399532
rect 477539 399467 477605 399468
rect 477726 398853 477786 406403
rect 486187 405788 486253 405789
rect 486187 405724 486188 405788
rect 486252 405724 486253 405788
rect 486187 405723 486253 405724
rect 486190 405650 486250 405723
rect 486190 405590 486434 405650
rect 479379 405244 479445 405245
rect 479379 405180 479380 405244
rect 479444 405180 479445 405244
rect 479379 405179 479445 405180
rect 478091 402524 478157 402525
rect 478091 402460 478092 402524
rect 478156 402460 478157 402524
rect 478091 402459 478157 402460
rect 477723 398852 477789 398853
rect 477723 398788 477724 398852
rect 477788 398788 477789 398852
rect 477723 398787 477789 398788
rect 477355 394500 477421 394501
rect 477355 394436 477356 394500
rect 477420 394436 477421 394500
rect 477355 394435 477421 394436
rect 478094 393141 478154 402459
rect 478643 399668 478709 399669
rect 478643 399604 478644 399668
rect 478708 399604 478709 399668
rect 478643 399603 478709 399604
rect 478646 397901 478706 399603
rect 478643 397900 478709 397901
rect 478643 397836 478644 397900
rect 478708 397836 478709 397900
rect 478643 397835 478709 397836
rect 478091 393140 478157 393141
rect 478091 393076 478092 393140
rect 478156 393076 478157 393140
rect 478091 393075 478157 393076
rect 479382 389061 479442 405179
rect 486003 405108 486069 405109
rect 486003 405044 486004 405108
rect 486068 405044 486069 405108
rect 486003 405043 486069 405044
rect 479563 403884 479629 403885
rect 479563 403820 479564 403884
rect 479628 403820 479629 403884
rect 479563 403819 479629 403820
rect 479566 391101 479626 403819
rect 479747 403748 479813 403749
rect 479747 403684 479748 403748
rect 479812 403684 479813 403748
rect 479747 403683 479813 403684
rect 479750 391781 479810 403683
rect 480851 403204 480917 403205
rect 480851 403140 480852 403204
rect 480916 403140 480917 403204
rect 480851 403139 480917 403140
rect 480854 392461 480914 403139
rect 483243 402388 483309 402389
rect 483243 402324 483244 402388
rect 483308 402324 483309 402388
rect 483243 402323 483309 402324
rect 483246 393821 483306 402323
rect 484899 401164 484965 401165
rect 484899 401100 484900 401164
rect 484964 401100 484965 401164
rect 484899 401099 484965 401100
rect 484715 401028 484781 401029
rect 484715 400964 484716 401028
rect 484780 400964 484781 401028
rect 484715 400963 484781 400964
rect 484531 400348 484597 400349
rect 484531 400284 484532 400348
rect 484596 400284 484597 400348
rect 484531 400283 484597 400284
rect 484347 399804 484413 399805
rect 484347 399740 484348 399804
rect 484412 399740 484413 399804
rect 484347 399739 484413 399740
rect 484350 397221 484410 399739
rect 484347 397220 484413 397221
rect 484347 397156 484348 397220
rect 484412 397156 484413 397220
rect 484347 397155 484413 397156
rect 484534 396541 484594 400283
rect 484531 396540 484597 396541
rect 484531 396476 484532 396540
rect 484596 396476 484597 396540
rect 484531 396475 484597 396476
rect 484718 395861 484778 400963
rect 484715 395860 484781 395861
rect 484715 395796 484716 395860
rect 484780 395796 484781 395860
rect 484715 395795 484781 395796
rect 484902 395181 484962 401099
rect 484899 395180 484965 395181
rect 484899 395116 484900 395180
rect 484964 395116 484965 395180
rect 484899 395115 484965 395116
rect 483243 393820 483309 393821
rect 483243 393756 483244 393820
rect 483308 393756 483309 393820
rect 483243 393755 483309 393756
rect 480851 392460 480917 392461
rect 480851 392396 480852 392460
rect 480916 392396 480917 392460
rect 480851 392395 480917 392396
rect 479747 391780 479813 391781
rect 479747 391716 479748 391780
rect 479812 391716 479813 391780
rect 479747 391715 479813 391716
rect 479563 391100 479629 391101
rect 479563 391036 479564 391100
rect 479628 391036 479629 391100
rect 479563 391035 479629 391036
rect 486006 389741 486066 405043
rect 486187 404428 486253 404429
rect 486187 404364 486188 404428
rect 486252 404364 486253 404428
rect 486187 404363 486253 404364
rect 486190 393330 486250 404363
rect 486374 402990 486434 405590
rect 486374 402930 486618 402990
rect 486190 393270 486434 393330
rect 486374 390421 486434 393270
rect 486371 390420 486437 390421
rect 486371 390356 486372 390420
rect 486436 390356 486437 390420
rect 486371 390355 486437 390356
rect 486003 389740 486069 389741
rect 486003 389676 486004 389740
rect 486068 389676 486069 389740
rect 486003 389675 486069 389676
rect 479379 389060 479445 389061
rect 479379 388996 479380 389060
rect 479444 388996 479445 389060
rect 479379 388995 479445 388996
rect 486558 388381 486618 402930
rect 486555 388380 486621 388381
rect 486555 388316 486556 388380
rect 486620 388316 486621 388380
rect 486555 388315 486621 388316
rect 482139 357100 482205 357101
rect 482139 357036 482140 357100
rect 482204 357036 482205 357100
rect 482139 357035 482205 357036
rect 480851 355740 480917 355741
rect 480851 355676 480852 355740
rect 480916 355676 480917 355740
rect 480851 355675 480917 355676
rect 478091 354380 478157 354381
rect 478091 354316 478092 354380
rect 478156 354316 478157 354380
rect 478091 354315 478157 354316
rect 477907 350300 477973 350301
rect 477907 350236 477908 350300
rect 477972 350236 477973 350300
rect 477907 350235 477973 350236
rect 477355 340780 477421 340781
rect 477355 340716 477356 340780
rect 477420 340716 477421 340780
rect 477355 340715 477421 340716
rect 477358 336905 477418 340715
rect 477355 336904 477421 336905
rect 477355 336840 477356 336904
rect 477420 336840 477421 336904
rect 477355 336839 477421 336840
rect 477355 335884 477421 335885
rect 477355 335820 477356 335884
rect 477420 335820 477421 335884
rect 477355 335819 477421 335820
rect 477358 333913 477418 335819
rect 477910 335205 477970 350235
rect 477907 335204 477973 335205
rect 477907 335140 477908 335204
rect 477972 335140 477973 335204
rect 477907 335139 477973 335140
rect 477355 333912 477421 333913
rect 477355 333848 477356 333912
rect 477420 333848 477421 333912
rect 477355 333847 477421 333848
rect 477355 332620 477421 332621
rect 477355 332556 477356 332620
rect 477420 332556 477421 332620
rect 477355 332555 477421 332556
rect 477358 331193 477418 332555
rect 477355 331192 477421 331193
rect 477355 331128 477356 331192
rect 477420 331128 477421 331192
rect 477355 331127 477421 331128
rect 477907 329628 477973 329629
rect 477907 329564 477908 329628
rect 477972 329564 477973 329628
rect 477907 329563 477973 329564
rect 477910 327317 477970 329563
rect 478094 327997 478154 354315
rect 478275 353020 478341 353021
rect 478275 352956 478276 353020
rect 478340 352956 478341 353020
rect 478275 352955 478341 352956
rect 478278 328677 478338 352955
rect 478459 352340 478525 352341
rect 478459 352276 478460 352340
rect 478524 352276 478525 352340
rect 478459 352275 478525 352276
rect 478462 329357 478522 352275
rect 479379 345540 479445 345541
rect 479379 345476 479380 345540
rect 479444 345476 479445 345540
rect 479379 345475 479445 345476
rect 478827 340100 478893 340101
rect 478827 340036 478828 340100
rect 478892 340036 478893 340100
rect 478827 340035 478893 340036
rect 478830 337517 478890 340035
rect 478827 337516 478893 337517
rect 478827 337452 478828 337516
rect 478892 337452 478893 337516
rect 478827 337451 478893 337452
rect 479011 334660 479077 334661
rect 479011 334596 479012 334660
rect 479076 334596 479077 334660
rect 479011 334595 479077 334596
rect 478643 334116 478709 334117
rect 478643 334052 478644 334116
rect 478708 334052 478709 334116
rect 478643 334051 478709 334052
rect 478459 329356 478525 329357
rect 478459 329292 478460 329356
rect 478524 329292 478525 329356
rect 478459 329291 478525 329292
rect 478275 328676 478341 328677
rect 478275 328612 478276 328676
rect 478340 328612 478341 328676
rect 478275 328611 478341 328612
rect 478646 328133 478706 334051
rect 478827 333980 478893 333981
rect 478827 333916 478828 333980
rect 478892 333916 478893 333980
rect 478827 333915 478893 333916
rect 478830 331669 478890 333915
rect 479014 332485 479074 334595
rect 479382 333573 479442 345475
rect 479747 343500 479813 343501
rect 479747 343436 479748 343500
rect 479812 343436 479813 343500
rect 479747 343435 479813 343436
rect 479563 338740 479629 338741
rect 479563 338676 479564 338740
rect 479628 338676 479629 338740
rect 479563 338675 479629 338676
rect 479379 333572 479445 333573
rect 479379 333508 479380 333572
rect 479444 333508 479445 333572
rect 479379 333507 479445 333508
rect 479011 332484 479077 332485
rect 479011 332420 479012 332484
rect 479076 332420 479077 332484
rect 479011 332419 479077 332420
rect 478827 331668 478893 331669
rect 478827 331604 478828 331668
rect 478892 331604 478893 331668
rect 478827 331603 478893 331604
rect 479566 330853 479626 338675
rect 479750 334933 479810 343435
rect 480299 336700 480365 336701
rect 480299 336636 480300 336700
rect 480364 336636 480365 336700
rect 480299 336635 480365 336636
rect 479747 334932 479813 334933
rect 479747 334868 479748 334932
rect 479812 334868 479813 334932
rect 479747 334867 479813 334868
rect 479563 330852 479629 330853
rect 479563 330788 479564 330852
rect 479628 330788 479629 330852
rect 479563 330787 479629 330788
rect 478643 328132 478709 328133
rect 478643 328068 478644 328132
rect 478708 328068 478709 328132
rect 478643 328067 478709 328068
rect 478091 327996 478157 327997
rect 478091 327932 478092 327996
rect 478156 327932 478157 327996
rect 478091 327931 478157 327932
rect 477907 327316 477973 327317
rect 477907 327252 477908 327316
rect 477972 327252 477973 327316
rect 477907 327251 477973 327252
rect 480302 325141 480362 336635
rect 480483 334116 480549 334117
rect 480483 334052 480484 334116
rect 480548 334052 480549 334116
rect 480483 334051 480549 334052
rect 480299 325140 480365 325141
rect 480299 325076 480300 325140
rect 480364 325076 480365 325140
rect 480299 325075 480365 325076
rect 480486 323781 480546 334051
rect 480854 326773 480914 355675
rect 481035 351660 481101 351661
rect 481035 351596 481036 351660
rect 481100 351596 481101 351660
rect 481035 351595 481101 351596
rect 481038 329493 481098 351595
rect 481219 348940 481285 348941
rect 481219 348876 481220 348940
rect 481284 348876 481285 348940
rect 481219 348875 481285 348876
rect 481222 336021 481282 348875
rect 481403 344180 481469 344181
rect 481403 344116 481404 344180
rect 481468 344116 481469 344180
rect 481403 344115 481469 344116
rect 481219 336020 481285 336021
rect 481219 335956 481220 336020
rect 481284 335956 481285 336020
rect 481219 335955 481285 335956
rect 481406 334797 481466 344115
rect 481771 336700 481837 336701
rect 481771 336636 481772 336700
rect 481836 336636 481837 336700
rect 481771 336635 481837 336636
rect 481403 334796 481469 334797
rect 481403 334732 481404 334796
rect 481468 334732 481469 334796
rect 481403 334731 481469 334732
rect 481035 329492 481101 329493
rect 481035 329428 481036 329492
rect 481100 329428 481101 329492
rect 481035 329427 481101 329428
rect 480851 326772 480917 326773
rect 480851 326708 480852 326772
rect 480916 326708 480917 326772
rect 480851 326707 480917 326708
rect 481774 324597 481834 336635
rect 482142 325957 482202 357035
rect 483611 356420 483677 356421
rect 483611 356356 483612 356420
rect 483676 356356 483677 356420
rect 483611 356355 483677 356356
rect 482323 350980 482389 350981
rect 482323 350916 482324 350980
rect 482388 350916 482389 350980
rect 482323 350915 482389 350916
rect 482326 332077 482386 350915
rect 482691 348260 482757 348261
rect 482691 348196 482692 348260
rect 482756 348196 482757 348260
rect 482691 348195 482757 348196
rect 482507 347580 482573 347581
rect 482507 347516 482508 347580
rect 482572 347516 482573 347580
rect 482507 347515 482573 347516
rect 482510 332213 482570 347515
rect 482694 336565 482754 348195
rect 483427 342140 483493 342141
rect 483427 342076 483428 342140
rect 483492 342076 483493 342140
rect 483427 342075 483493 342076
rect 483243 339420 483309 339421
rect 483243 339356 483244 339420
rect 483308 339356 483309 339420
rect 483243 339355 483309 339356
rect 483246 337653 483306 339355
rect 483430 338197 483490 342075
rect 483427 338196 483493 338197
rect 483427 338132 483428 338196
rect 483492 338132 483493 338196
rect 483427 338131 483493 338132
rect 483243 337652 483309 337653
rect 483243 337588 483244 337652
rect 483308 337588 483309 337652
rect 483243 337587 483309 337588
rect 483059 336700 483125 336701
rect 483059 336636 483060 336700
rect 483124 336636 483125 336700
rect 483059 336635 483125 336636
rect 482691 336564 482757 336565
rect 482691 336500 482692 336564
rect 482756 336500 482757 336564
rect 482691 336499 482757 336500
rect 482507 332212 482573 332213
rect 482507 332148 482508 332212
rect 482572 332148 482573 332212
rect 482507 332147 482573 332148
rect 482323 332076 482389 332077
rect 482323 332012 482324 332076
rect 482388 332012 482389 332076
rect 482323 332011 482389 332012
rect 482875 331940 482941 331941
rect 482875 331876 482876 331940
rect 482940 331876 482941 331940
rect 482875 331875 482941 331876
rect 482878 330581 482938 331875
rect 482875 330580 482941 330581
rect 482875 330516 482876 330580
rect 482940 330516 482941 330580
rect 482875 330515 482941 330516
rect 482139 325956 482205 325957
rect 482139 325892 482140 325956
rect 482204 325892 482205 325956
rect 482139 325891 482205 325892
rect 483062 325413 483122 336635
rect 483243 334116 483309 334117
rect 483243 334052 483244 334116
rect 483308 334052 483309 334116
rect 483243 334051 483309 334052
rect 483059 325412 483125 325413
rect 483059 325348 483060 325412
rect 483124 325348 483125 325412
rect 483059 325347 483125 325348
rect 481771 324596 481837 324597
rect 481771 324532 481772 324596
rect 481836 324532 481837 324596
rect 481771 324531 481837 324532
rect 483246 324053 483306 334051
rect 483427 333300 483493 333301
rect 483427 333236 483428 333300
rect 483492 333236 483493 333300
rect 483427 333235 483493 333236
rect 483430 331397 483490 333235
rect 483427 331396 483493 331397
rect 483427 331332 483428 331396
rect 483492 331332 483493 331396
rect 483427 331331 483493 331332
rect 483614 326637 483674 356355
rect 483795 346220 483861 346221
rect 483795 346156 483796 346220
rect 483860 346156 483861 346220
rect 483795 346155 483861 346156
rect 483798 333437 483858 346155
rect 486003 344860 486069 344861
rect 486003 344796 486004 344860
rect 486068 344796 486069 344860
rect 486003 344795 486069 344796
rect 483979 342820 484045 342821
rect 483979 342756 483980 342820
rect 484044 342756 484045 342820
rect 483979 342755 484045 342756
rect 483982 335477 484042 342755
rect 484347 341460 484413 341461
rect 484347 341396 484348 341460
rect 484412 341396 484413 341460
rect 484347 341395 484413 341396
rect 484350 336293 484410 341395
rect 484715 336700 484781 336701
rect 484715 336636 484716 336700
rect 484780 336636 484781 336700
rect 484715 336635 484781 336636
rect 484347 336292 484413 336293
rect 484347 336228 484348 336292
rect 484412 336228 484413 336292
rect 484347 336227 484413 336228
rect 483979 335476 484045 335477
rect 483979 335412 483980 335476
rect 484044 335412 484045 335476
rect 483979 335411 484045 335412
rect 484347 335340 484413 335341
rect 484347 335276 484348 335340
rect 484412 335276 484413 335340
rect 484347 335275 484413 335276
rect 483795 333436 483861 333437
rect 483795 333372 483796 333436
rect 483860 333372 483861 333436
rect 483795 333371 483861 333372
rect 484350 333029 484410 335275
rect 484718 334389 484778 336635
rect 484715 334388 484781 334389
rect 484715 334324 484716 334388
rect 484780 334324 484781 334388
rect 484715 334323 484781 334324
rect 486006 334253 486066 344795
rect 486003 334252 486069 334253
rect 486003 334188 486004 334252
rect 486068 334188 486069 334252
rect 486003 334187 486069 334188
rect 484347 333028 484413 333029
rect 484347 332964 484348 333028
rect 484412 332964 484413 333028
rect 484347 332963 484413 332964
rect 483611 326636 483677 326637
rect 483611 326572 483612 326636
rect 483676 326572 483677 326636
rect 483611 326571 483677 326572
rect 483243 324052 483309 324053
rect 483243 323988 483244 324052
rect 483308 323988 483309 324052
rect 483243 323987 483309 323988
rect 480483 323780 480549 323781
rect 480483 323716 480484 323780
rect 480548 323716 480549 323780
rect 480483 323715 480549 323716
rect 481771 322964 481837 322965
rect 481771 322900 481772 322964
rect 481836 322900 481837 322964
rect 481771 322899 481837 322900
rect 480667 322692 480733 322693
rect 480667 322628 480668 322692
rect 480732 322628 480733 322692
rect 480667 322627 480733 322628
rect 480670 318749 480730 322627
rect 481587 321604 481653 321605
rect 481587 321540 481588 321604
rect 481652 321540 481653 321604
rect 481587 321539 481653 321540
rect 480851 321332 480917 321333
rect 480851 321268 480852 321332
rect 480916 321268 480917 321332
rect 480851 321267 480917 321268
rect 480667 318748 480733 318749
rect 480667 318684 480668 318748
rect 480732 318684 480733 318748
rect 480667 318683 480733 318684
rect 479379 317252 479445 317253
rect 479379 317188 479380 317252
rect 479444 317188 479445 317252
rect 479379 317187 479445 317188
rect 478091 315892 478157 315893
rect 478091 315828 478092 315892
rect 478156 315828 478157 315892
rect 478091 315827 478157 315828
rect 478094 298621 478154 315827
rect 478275 315348 478341 315349
rect 478275 315284 478276 315348
rect 478340 315284 478341 315348
rect 478275 315283 478341 315284
rect 478278 299301 478338 315283
rect 479382 314941 479442 317187
rect 479747 316708 479813 316709
rect 479747 316644 479748 316708
rect 479812 316644 479813 316708
rect 479747 316643 479813 316644
rect 479379 314940 479445 314941
rect 479379 314876 479380 314940
rect 479444 314876 479445 314940
rect 479379 314875 479445 314876
rect 479750 311269 479810 316643
rect 479931 316164 479997 316165
rect 479931 316100 479932 316164
rect 479996 316100 479997 316164
rect 479931 316099 479997 316100
rect 479747 311268 479813 311269
rect 479747 311204 479748 311268
rect 479812 311204 479813 311268
rect 479747 311203 479813 311204
rect 479934 310453 479994 316099
rect 478643 310452 478709 310453
rect 478643 310388 478644 310452
rect 478708 310388 478709 310452
rect 478643 310387 478709 310388
rect 479931 310452 479997 310453
rect 479931 310388 479932 310452
rect 479996 310388 479997 310452
rect 479931 310387 479997 310388
rect 478646 306781 478706 310387
rect 478643 306780 478709 306781
rect 478643 306716 478644 306780
rect 478708 306716 478709 306780
rect 478643 306715 478709 306716
rect 478275 299300 478341 299301
rect 478275 299236 478276 299300
rect 478340 299236 478341 299300
rect 478275 299235 478341 299236
rect 478091 298620 478157 298621
rect 478091 298556 478092 298620
rect 478156 298556 478157 298620
rect 478091 298555 478157 298556
rect 480854 290461 480914 321267
rect 481035 319428 481101 319429
rect 481035 319364 481036 319428
rect 481100 319364 481101 319428
rect 481035 319363 481101 319364
rect 481038 293181 481098 319363
rect 481219 318068 481285 318069
rect 481219 318004 481220 318068
rect 481284 318004 481285 318068
rect 481219 318003 481285 318004
rect 481222 295221 481282 318003
rect 481403 317660 481469 317661
rect 481403 317596 481404 317660
rect 481468 317596 481469 317660
rect 481403 317595 481469 317596
rect 481406 310453 481466 317595
rect 481403 310452 481469 310453
rect 481403 310388 481404 310452
rect 481468 310388 481469 310452
rect 481403 310387 481469 310388
rect 481590 308957 481650 321539
rect 481774 311949 481834 322899
rect 483059 322148 483125 322149
rect 483059 322084 483060 322148
rect 483124 322084 483125 322148
rect 483059 322083 483125 322084
rect 482139 318884 482205 318885
rect 482139 318820 482140 318884
rect 482204 318820 482205 318884
rect 482139 318819 482205 318820
rect 481771 311948 481837 311949
rect 481771 311884 481772 311948
rect 481836 311884 481837 311948
rect 481771 311883 481837 311884
rect 481587 308956 481653 308957
rect 481587 308892 481588 308956
rect 481652 308892 481653 308956
rect 481587 308891 481653 308892
rect 481219 295220 481285 295221
rect 481219 295156 481220 295220
rect 481284 295156 481285 295220
rect 481219 295155 481285 295156
rect 482142 293861 482202 318819
rect 482323 318612 482389 318613
rect 482323 318548 482324 318612
rect 482388 318548 482389 318612
rect 482323 318547 482389 318548
rect 482326 294541 482386 318547
rect 483062 311269 483122 322083
rect 483611 320788 483677 320789
rect 483611 320724 483612 320788
rect 483676 320724 483677 320788
rect 483611 320723 483677 320724
rect 483059 311268 483125 311269
rect 483059 311204 483060 311268
rect 483124 311204 483125 311268
rect 483059 311203 483125 311204
rect 482875 309908 482941 309909
rect 482875 309844 482876 309908
rect 482940 309844 482941 309908
rect 482875 309843 482941 309844
rect 482878 307461 482938 309843
rect 482875 307460 482941 307461
rect 482875 307396 482876 307460
rect 482940 307396 482941 307460
rect 482875 307395 482941 307396
rect 482323 294540 482389 294541
rect 482323 294476 482324 294540
rect 482388 294476 482389 294540
rect 482323 294475 482389 294476
rect 482139 293860 482205 293861
rect 482139 293796 482140 293860
rect 482204 293796 482205 293860
rect 482139 293795 482205 293796
rect 481035 293180 481101 293181
rect 481035 293116 481036 293180
rect 481100 293116 481101 293180
rect 481035 293115 481101 293116
rect 483614 291141 483674 320723
rect 483795 320244 483861 320245
rect 483795 320180 483796 320244
rect 483860 320180 483861 320244
rect 483795 320179 483861 320180
rect 483798 291821 483858 320179
rect 483979 319972 484045 319973
rect 483979 319908 483980 319972
rect 484044 319908 484045 319972
rect 483979 319907 484045 319908
rect 483982 292501 484042 319907
rect 486187 313988 486253 313989
rect 486187 313924 486188 313988
rect 486252 313924 486253 313988
rect 486187 313923 486253 313924
rect 486190 313850 486250 313923
rect 486190 313790 486434 313850
rect 485083 313444 485149 313445
rect 485083 313380 485084 313444
rect 485148 313380 485149 313444
rect 485083 313379 485149 313380
rect 484899 311812 484965 311813
rect 484899 311748 484900 311812
rect 484964 311748 484965 311812
rect 484899 311747 484965 311748
rect 484347 309364 484413 309365
rect 484347 309300 484348 309364
rect 484412 309300 484413 309364
rect 484347 309299 484413 309300
rect 484350 308141 484410 309299
rect 484347 308140 484413 308141
rect 484347 308076 484348 308140
rect 484412 308076 484413 308140
rect 484347 308075 484413 308076
rect 484902 304741 484962 311747
rect 484899 304740 484965 304741
rect 484899 304676 484900 304740
rect 484964 304676 484965 304740
rect 484899 304675 484965 304676
rect 485086 302021 485146 313379
rect 486003 313172 486069 313173
rect 486003 313108 486004 313172
rect 486068 313108 486069 313172
rect 486003 313107 486069 313108
rect 485819 312628 485885 312629
rect 485819 312564 485820 312628
rect 485884 312564 485885 312628
rect 485819 312563 485885 312564
rect 485635 312084 485701 312085
rect 485635 312020 485636 312084
rect 485700 312020 485701 312084
rect 485635 312019 485701 312020
rect 485267 311132 485333 311133
rect 485267 311068 485268 311132
rect 485332 311068 485333 311132
rect 485267 311067 485333 311068
rect 485270 305421 485330 311067
rect 485451 310724 485517 310725
rect 485451 310660 485452 310724
rect 485516 310660 485517 310724
rect 485451 310659 485517 310660
rect 485454 306101 485514 310659
rect 485451 306100 485517 306101
rect 485451 306036 485452 306100
rect 485516 306036 485517 306100
rect 485451 306035 485517 306036
rect 485267 305420 485333 305421
rect 485267 305356 485268 305420
rect 485332 305356 485333 305420
rect 485267 305355 485333 305356
rect 485638 304061 485698 312019
rect 485635 304060 485701 304061
rect 485635 303996 485636 304060
rect 485700 303996 485701 304060
rect 485635 303995 485701 303996
rect 485822 303381 485882 312563
rect 485819 303380 485885 303381
rect 485819 303316 485820 303380
rect 485884 303316 485885 303380
rect 485819 303315 485885 303316
rect 486006 302701 486066 313107
rect 486187 308548 486253 308549
rect 486187 308484 486188 308548
rect 486252 308484 486253 308548
rect 486187 308483 486253 308484
rect 486003 302700 486069 302701
rect 486003 302636 486004 302700
rect 486068 302636 486069 302700
rect 486003 302635 486069 302636
rect 485083 302020 485149 302021
rect 485083 301956 485084 302020
rect 485148 301956 485149 302020
rect 485083 301955 485149 301956
rect 486190 296730 486250 308483
rect 486374 301341 486434 313790
rect 486371 301340 486437 301341
rect 486371 301276 486372 301340
rect 486436 301276 486437 301340
rect 486371 301275 486437 301276
rect 486190 296670 486434 296730
rect 486374 295901 486434 296670
rect 486371 295900 486437 295901
rect 486371 295836 486372 295900
rect 486436 295836 486437 295900
rect 486371 295835 486437 295836
rect 483979 292500 484045 292501
rect 483979 292436 483980 292500
rect 484044 292436 484045 292500
rect 483979 292435 484045 292436
rect 483795 291820 483861 291821
rect 483795 291756 483796 291820
rect 483860 291756 483861 291820
rect 483795 291755 483861 291756
rect 483611 291140 483677 291141
rect 483611 291076 483612 291140
rect 483676 291076 483677 291140
rect 483611 291075 483677 291076
rect 480851 290460 480917 290461
rect 480851 290396 480852 290460
rect 480916 290396 480917 290460
rect 480851 290395 480917 290396
rect 483611 267340 483677 267341
rect 483611 267276 483612 267340
rect 483676 267276 483677 267340
rect 483611 267275 483677 267276
rect 480851 265300 480917 265301
rect 480851 265236 480852 265300
rect 480916 265236 480917 265300
rect 480851 265235 480917 265236
rect 478091 262580 478157 262581
rect 478091 262516 478092 262580
rect 478156 262516 478157 262580
rect 478091 262515 478157 262516
rect 477539 248028 477605 248029
rect 477539 247964 477540 248028
rect 477604 247964 477605 248028
rect 477539 247963 477605 247964
rect 477542 247890 477602 247963
rect 477174 247830 477602 247890
rect 477174 246883 477234 247830
rect 477539 247076 477605 247077
rect 477539 247012 477540 247076
rect 477604 247012 477605 247076
rect 477539 247011 477605 247012
rect 477355 246940 477421 246941
rect 477171 246882 477237 246883
rect 477171 246818 477172 246882
rect 477236 246818 477237 246882
rect 477355 246876 477356 246940
rect 477420 246876 477421 246940
rect 477355 246875 477421 246876
rect 477171 246817 477237 246818
rect 477358 245523 477418 246875
rect 477355 245522 477421 245523
rect 477355 245458 477356 245522
rect 477420 245458 477421 245522
rect 477355 245457 477421 245458
rect 477542 238509 477602 247011
rect 477723 245716 477789 245717
rect 477723 245652 477724 245716
rect 477788 245652 477789 245716
rect 477723 245651 477789 245652
rect 477539 238508 477605 238509
rect 477539 238444 477540 238508
rect 477604 238444 477605 238508
rect 477539 238443 477605 238444
rect 477726 237693 477786 245651
rect 477907 242860 477973 242861
rect 477907 242796 477908 242860
rect 477972 242796 477973 242860
rect 477907 242795 477973 242796
rect 477910 238237 477970 242795
rect 478094 239053 478154 262515
rect 478275 261220 478341 261221
rect 478275 261156 478276 261220
rect 478340 261156 478341 261220
rect 478275 261155 478341 261156
rect 478278 242045 478338 261155
rect 479563 258500 479629 258501
rect 479563 258436 479564 258500
rect 479628 258436 479629 258500
rect 479563 258435 479629 258436
rect 479379 256460 479445 256461
rect 479379 256396 479380 256460
rect 479444 256396 479445 256460
rect 479379 256395 479445 256396
rect 479382 243133 479442 256395
rect 479566 246397 479626 258435
rect 479747 255100 479813 255101
rect 479747 255036 479748 255100
rect 479812 255036 479813 255100
rect 479747 255035 479813 255036
rect 479563 246396 479629 246397
rect 479563 246332 479564 246396
rect 479628 246332 479629 246396
rect 479563 246331 479629 246332
rect 479750 243949 479810 255035
rect 479931 253060 479997 253061
rect 479931 252996 479932 253060
rect 479996 252996 479997 253060
rect 479931 252995 479997 252996
rect 479934 245309 479994 252995
rect 480299 247076 480365 247077
rect 480299 247012 480300 247076
rect 480364 247012 480365 247076
rect 480299 247011 480365 247012
rect 479931 245308 479997 245309
rect 479931 245244 479932 245308
rect 479996 245244 479997 245308
rect 479931 245243 479997 245244
rect 479747 243948 479813 243949
rect 479747 243884 479748 243948
rect 479812 243884 479813 243948
rect 479747 243883 479813 243884
rect 479379 243132 479445 243133
rect 479379 243068 479380 243132
rect 479444 243068 479445 243132
rect 479379 243067 479445 243068
rect 478275 242044 478341 242045
rect 478275 241980 478276 242044
rect 478340 241980 478341 242044
rect 478275 241979 478341 241980
rect 478091 239052 478157 239053
rect 478091 238988 478092 239052
rect 478156 238988 478157 239052
rect 478091 238987 478157 238988
rect 477907 238236 477973 238237
rect 477907 238172 477908 238236
rect 477972 238172 477973 238236
rect 477907 238171 477973 238172
rect 477723 237692 477789 237693
rect 477723 237628 477724 237692
rect 477788 237628 477789 237692
rect 477723 237627 477789 237628
rect 480302 235517 480362 247011
rect 480483 244356 480549 244357
rect 480483 244292 480484 244356
rect 480548 244292 480549 244356
rect 480483 244291 480549 244292
rect 480299 235516 480365 235517
rect 480299 235452 480300 235516
rect 480364 235452 480365 235516
rect 480299 235451 480365 235452
rect 480486 234157 480546 244291
rect 480854 237149 480914 265235
rect 482139 261900 482205 261901
rect 482139 261836 482140 261900
rect 482204 261836 482205 261900
rect 482139 261835 482205 261836
rect 481035 259180 481101 259181
rect 481035 259116 481036 259180
rect 481100 259116 481101 259180
rect 481035 259115 481101 259116
rect 481038 245853 481098 259115
rect 481219 252380 481285 252381
rect 481219 252316 481220 252380
rect 481284 252316 481285 252380
rect 481219 252315 481285 252316
rect 481222 247893 481282 252315
rect 481587 249660 481653 249661
rect 481587 249596 481588 249660
rect 481652 249596 481653 249660
rect 481587 249595 481653 249596
rect 481219 247892 481285 247893
rect 481219 247828 481220 247892
rect 481284 247828 481285 247892
rect 481219 247827 481285 247828
rect 481590 247757 481650 249595
rect 481587 247756 481653 247757
rect 481587 247692 481588 247756
rect 481652 247692 481653 247756
rect 481587 247691 481653 247692
rect 481771 247076 481837 247077
rect 481771 247012 481772 247076
rect 481836 247012 481837 247076
rect 481771 247011 481837 247012
rect 481035 245852 481101 245853
rect 481035 245788 481036 245852
rect 481100 245788 481101 245852
rect 481035 245787 481101 245788
rect 481587 245716 481653 245717
rect 481587 245652 481588 245716
rect 481652 245652 481653 245716
rect 481587 245651 481653 245652
rect 480851 237148 480917 237149
rect 480851 237084 480852 237148
rect 480916 237084 480917 237148
rect 480851 237083 480917 237084
rect 481590 234429 481650 245651
rect 481774 236333 481834 247011
rect 482142 239597 482202 261835
rect 482323 260540 482389 260541
rect 482323 260476 482324 260540
rect 482388 260476 482389 260540
rect 482323 260475 482389 260476
rect 482326 243677 482386 260475
rect 482875 247620 482941 247621
rect 482875 247556 482876 247620
rect 482940 247556 482941 247620
rect 482875 247555 482941 247556
rect 482878 246125 482938 247555
rect 483243 246260 483309 246261
rect 483243 246196 483244 246260
rect 483308 246196 483309 246260
rect 483243 246195 483309 246196
rect 482875 246124 482941 246125
rect 482875 246060 482876 246124
rect 482940 246060 482941 246124
rect 482875 246059 482941 246060
rect 483246 244765 483306 246195
rect 483243 244764 483309 244765
rect 483243 244700 483244 244764
rect 483308 244700 483309 244764
rect 483243 244699 483309 244700
rect 482323 243676 482389 243677
rect 482323 243612 482324 243676
rect 482388 243612 482389 243676
rect 482323 243611 482389 243612
rect 483059 243540 483125 243541
rect 483059 243476 483060 243540
rect 483124 243476 483125 243540
rect 483059 243475 483125 243476
rect 482139 239596 482205 239597
rect 482139 239532 482140 239596
rect 482204 239532 482205 239596
rect 482139 239531 482205 239532
rect 481771 236332 481837 236333
rect 481771 236268 481772 236332
rect 481836 236268 481837 236332
rect 481771 236267 481837 236268
rect 483062 234973 483122 243475
rect 483243 242860 483309 242861
rect 483243 242796 483244 242860
rect 483308 242796 483309 242860
rect 483243 242795 483309 242796
rect 483246 241093 483306 242795
rect 483243 241092 483309 241093
rect 483243 241028 483244 241092
rect 483308 241028 483309 241092
rect 483243 241027 483309 241028
rect 483614 235789 483674 267275
rect 483795 265980 483861 265981
rect 483795 265916 483796 265980
rect 483860 265916 483861 265980
rect 483795 265915 483861 265916
rect 483798 236877 483858 265915
rect 485635 259860 485701 259861
rect 485635 259796 485636 259860
rect 485700 259796 485701 259860
rect 485635 259795 485701 259796
rect 483979 257820 484045 257821
rect 483979 257756 483980 257820
rect 484044 257756 484045 257820
rect 483979 257755 484045 257756
rect 483982 242317 484042 257755
rect 485451 257140 485517 257141
rect 485451 257076 485452 257140
rect 485516 257076 485517 257140
rect 485451 257075 485517 257076
rect 484531 251020 484597 251021
rect 484531 250956 484532 251020
rect 484596 250956 484597 251020
rect 484531 250955 484597 250956
rect 484347 248980 484413 248981
rect 484347 248916 484348 248980
rect 484412 248916 484413 248980
rect 484347 248915 484413 248916
rect 484350 247485 484410 248915
rect 484347 247484 484413 247485
rect 484347 247420 484348 247484
rect 484412 247420 484413 247484
rect 484347 247419 484413 247420
rect 484534 246669 484594 250955
rect 484715 250340 484781 250341
rect 484715 250276 484716 250340
rect 484780 250276 484781 250340
rect 484715 250275 484781 250276
rect 484718 247213 484778 250275
rect 484715 247212 484781 247213
rect 484715 247148 484716 247212
rect 484780 247148 484781 247212
rect 484715 247147 484781 247148
rect 484531 246668 484597 246669
rect 484531 246604 484532 246668
rect 484596 246604 484597 246668
rect 484531 246603 484597 246604
rect 484531 245580 484597 245581
rect 484531 245516 484532 245580
rect 484596 245516 484597 245580
rect 484531 245515 484597 245516
rect 484347 244900 484413 244901
rect 484347 244836 484348 244900
rect 484412 244836 484413 244900
rect 484347 244835 484413 244836
rect 484350 242725 484410 244835
rect 484534 243269 484594 245515
rect 484899 244220 484965 244221
rect 484899 244156 484900 244220
rect 484964 244156 484965 244220
rect 484899 244155 484965 244156
rect 484715 243540 484781 243541
rect 484715 243476 484716 243540
rect 484780 243476 484781 243540
rect 484715 243475 484781 243476
rect 484531 243268 484597 243269
rect 484531 243204 484532 243268
rect 484596 243204 484597 243268
rect 484531 243203 484597 243204
rect 484347 242724 484413 242725
rect 484347 242660 484348 242724
rect 484412 242660 484413 242724
rect 484347 242659 484413 242660
rect 483979 242316 484045 242317
rect 483979 242252 483980 242316
rect 484044 242252 484045 242316
rect 483979 242251 484045 242252
rect 484347 242180 484413 242181
rect 484347 242116 484348 242180
rect 484412 242116 484413 242180
rect 484347 242115 484413 242116
rect 484350 240957 484410 242115
rect 484718 241229 484778 243475
rect 484902 241365 484962 244155
rect 485454 242589 485514 257075
rect 485638 244085 485698 259795
rect 486371 254420 486437 254421
rect 486371 254356 486372 254420
rect 486436 254356 486437 254420
rect 486371 254355 486437 254356
rect 485819 253740 485885 253741
rect 485819 253676 485820 253740
rect 485884 253676 485885 253740
rect 485819 253675 485885 253676
rect 485822 245037 485882 253675
rect 486003 251700 486069 251701
rect 486003 251636 486004 251700
rect 486068 251636 486069 251700
rect 486003 251635 486069 251636
rect 486006 248165 486066 251635
rect 486003 248164 486069 248165
rect 486003 248100 486004 248164
rect 486068 248100 486069 248164
rect 486003 248099 486069 248100
rect 485819 245036 485885 245037
rect 485819 244972 485820 245036
rect 485884 244972 485885 245036
rect 485819 244971 485885 244972
rect 486187 244492 486253 244493
rect 486187 244428 486188 244492
rect 486252 244490 486253 244492
rect 486374 244490 486434 254355
rect 486252 244430 486434 244490
rect 486252 244428 486253 244430
rect 486187 244427 486253 244428
rect 485635 244084 485701 244085
rect 485635 244020 485636 244084
rect 485700 244020 485701 244084
rect 485635 244019 485701 244020
rect 485451 242588 485517 242589
rect 485451 242524 485452 242588
rect 485516 242524 485517 242588
rect 485451 242523 485517 242524
rect 484899 241364 484965 241365
rect 484899 241300 484900 241364
rect 484964 241300 484965 241364
rect 484899 241299 484965 241300
rect 484715 241228 484781 241229
rect 484715 241164 484716 241228
rect 484780 241164 484781 241228
rect 484715 241163 484781 241164
rect 484347 240956 484413 240957
rect 484347 240892 484348 240956
rect 484412 240892 484413 240956
rect 484347 240891 484413 240892
rect 483795 236876 483861 236877
rect 483795 236812 483796 236876
rect 483860 236812 483861 236876
rect 483795 236811 483861 236812
rect 483611 235788 483677 235789
rect 483611 235724 483612 235788
rect 483676 235724 483677 235788
rect 483611 235723 483677 235724
rect 483059 234972 483125 234973
rect 483059 234908 483060 234972
rect 483124 234908 483125 234972
rect 483059 234907 483125 234908
rect 481587 234428 481653 234429
rect 481587 234364 481588 234428
rect 481652 234364 481653 234428
rect 481587 234363 481653 234364
rect 480483 234156 480549 234157
rect 480483 234092 480484 234156
rect 480548 234092 480549 234156
rect 480483 234091 480549 234092
rect 483059 233204 483125 233205
rect 483059 233140 483060 233204
rect 483124 233140 483125 233204
rect 483059 233139 483125 233140
rect 477723 232796 477789 232797
rect 477723 232732 477724 232796
rect 477788 232732 477789 232796
rect 477723 232731 477789 232732
rect 477539 232388 477605 232389
rect 477539 232324 477540 232388
rect 477604 232324 477605 232388
rect 477539 232323 477605 232324
rect 477542 219333 477602 232323
rect 477726 220965 477786 232731
rect 480667 231844 480733 231845
rect 480667 231780 480668 231844
rect 480732 231780 480733 231844
rect 480667 231779 480733 231780
rect 480483 228308 480549 228309
rect 480483 228244 480484 228308
rect 480548 228244 480549 228308
rect 480483 228243 480549 228244
rect 480115 226948 480181 226949
rect 480115 226884 480116 226948
rect 480180 226884 480181 226948
rect 480115 226883 480181 226884
rect 479563 225588 479629 225589
rect 479563 225524 479564 225588
rect 479628 225524 479629 225588
rect 479563 225523 479629 225524
rect 479379 225044 479445 225045
rect 479379 224980 479380 225044
rect 479444 224980 479445 225044
rect 479379 224979 479445 224980
rect 477723 220964 477789 220965
rect 477723 220900 477724 220964
rect 477788 220900 477789 220964
rect 477723 220899 477789 220900
rect 477539 219332 477605 219333
rect 477539 219268 477540 219332
rect 477604 219268 477605 219332
rect 477539 219267 477605 219268
rect 479382 209541 479442 224979
rect 479379 209540 479445 209541
rect 479379 209476 479380 209540
rect 479444 209476 479445 209540
rect 479379 209475 479445 209476
rect 479566 208861 479626 225523
rect 480118 223685 480178 226883
rect 480115 223684 480181 223685
rect 480115 223620 480116 223684
rect 480180 223620 480181 223684
rect 480115 223619 480181 223620
rect 480486 220013 480546 228243
rect 480670 226405 480730 231779
rect 482875 231028 482941 231029
rect 482875 230964 482876 231028
rect 482940 230964 482941 231028
rect 482875 230963 482941 230964
rect 480851 230484 480917 230485
rect 480851 230420 480852 230484
rect 480916 230420 480917 230484
rect 480851 230419 480917 230420
rect 480667 226404 480733 226405
rect 480667 226340 480668 226404
rect 480732 226340 480733 226404
rect 480667 226339 480733 226340
rect 480483 220012 480549 220013
rect 480483 219948 480484 220012
rect 480548 219948 480549 220012
rect 480483 219947 480549 219948
rect 479563 208860 479629 208861
rect 479563 208796 479564 208860
rect 479628 208796 479629 208860
rect 479563 208795 479629 208796
rect 480854 201381 480914 230419
rect 481587 230212 481653 230213
rect 481587 230148 481588 230212
rect 481652 230148 481653 230212
rect 481587 230147 481653 230148
rect 481035 227492 481101 227493
rect 481035 227428 481036 227492
rect 481100 227428 481101 227492
rect 481035 227427 481101 227428
rect 481038 220965 481098 227427
rect 481219 226268 481285 226269
rect 481219 226204 481220 226268
rect 481284 226204 481285 226268
rect 481219 226203 481285 226204
rect 481035 220964 481101 220965
rect 481035 220900 481036 220964
rect 481100 220900 481101 220964
rect 481035 220899 481101 220900
rect 481035 220012 481101 220013
rect 481035 219948 481036 220012
rect 481100 219948 481101 220012
rect 481035 219947 481101 219948
rect 481038 204781 481098 219947
rect 481222 207501 481282 226203
rect 481590 220965 481650 230147
rect 482139 228852 482205 228853
rect 482139 228788 482140 228852
rect 482204 228788 482205 228852
rect 482139 228787 482205 228788
rect 481587 220964 481653 220965
rect 481587 220900 481588 220964
rect 481652 220900 481653 220964
rect 481587 220899 481653 220900
rect 481403 218788 481469 218789
rect 481403 218724 481404 218788
rect 481468 218724 481469 218788
rect 481403 218723 481469 218724
rect 481219 207500 481285 207501
rect 481219 207436 481220 207500
rect 481284 207436 481285 207500
rect 481219 207435 481285 207436
rect 481406 206141 481466 218723
rect 481403 206140 481469 206141
rect 481403 206076 481404 206140
rect 481468 206076 481469 206140
rect 481403 206075 481469 206076
rect 481035 204780 481101 204781
rect 481035 204716 481036 204780
rect 481100 204716 481101 204780
rect 481035 204715 481101 204716
rect 482142 204101 482202 228787
rect 482323 227764 482389 227765
rect 482323 227700 482324 227764
rect 482388 227700 482389 227764
rect 482323 227699 482389 227700
rect 482326 205461 482386 227699
rect 482507 224228 482573 224229
rect 482507 224164 482508 224228
rect 482572 224164 482573 224228
rect 482507 224163 482573 224164
rect 482510 210901 482570 224163
rect 482878 223685 482938 230963
rect 483062 223685 483122 233139
rect 483427 231708 483493 231709
rect 483427 231644 483428 231708
rect 483492 231644 483493 231708
rect 483427 231643 483493 231644
rect 482875 223684 482941 223685
rect 482875 223620 482876 223684
rect 482940 223620 482941 223684
rect 482875 223619 482941 223620
rect 483059 223684 483125 223685
rect 483059 223620 483060 223684
rect 483124 223620 483125 223684
rect 483059 223619 483125 223620
rect 483430 222325 483490 231643
rect 483611 229804 483677 229805
rect 483611 229740 483612 229804
rect 483676 229740 483677 229804
rect 483611 229739 483677 229740
rect 483427 222324 483493 222325
rect 483427 222260 483428 222324
rect 483492 222260 483493 222324
rect 483427 222259 483493 222260
rect 483059 219604 483125 219605
rect 483059 219540 483060 219604
rect 483124 219540 483125 219604
rect 483059 219539 483125 219540
rect 483062 217701 483122 219539
rect 483059 217700 483125 217701
rect 483059 217636 483060 217700
rect 483124 217636 483125 217700
rect 483059 217635 483125 217636
rect 482507 210900 482573 210901
rect 482507 210836 482508 210900
rect 482572 210836 482573 210900
rect 482507 210835 482573 210836
rect 482323 205460 482389 205461
rect 482323 205396 482324 205460
rect 482388 205396 482389 205460
rect 482323 205395 482389 205396
rect 482139 204100 482205 204101
rect 482139 204036 482140 204100
rect 482204 204036 482205 204100
rect 482139 204035 482205 204036
rect 483614 202741 483674 229739
rect 483795 229124 483861 229125
rect 483795 229060 483796 229124
rect 483860 229060 483861 229124
rect 483795 229059 483861 229060
rect 483798 203421 483858 229059
rect 486187 224772 486253 224773
rect 486187 224708 486188 224772
rect 486252 224770 486253 224772
rect 486252 224710 486618 224770
rect 486252 224708 486253 224710
rect 486187 224707 486253 224708
rect 485451 224092 485517 224093
rect 485451 224028 485452 224092
rect 485516 224028 485517 224092
rect 485451 224027 485517 224028
rect 483979 222868 484045 222869
rect 483979 222804 483980 222868
rect 484044 222804 484045 222868
rect 483979 222803 484045 222804
rect 483982 212941 484042 222803
rect 485267 222052 485333 222053
rect 485267 221988 485268 222052
rect 485332 221988 485333 222052
rect 485267 221987 485333 221988
rect 485083 221508 485149 221509
rect 485083 221444 485084 221508
rect 485148 221444 485149 221508
rect 485083 221443 485149 221444
rect 484715 221372 484781 221373
rect 484715 221308 484716 221372
rect 484780 221308 484781 221372
rect 484715 221307 484781 221308
rect 484531 220692 484597 220693
rect 484531 220628 484532 220692
rect 484596 220628 484597 220692
rect 484531 220627 484597 220628
rect 484347 220148 484413 220149
rect 484347 220084 484348 220148
rect 484412 220084 484413 220148
rect 484347 220083 484413 220084
rect 484350 217021 484410 220083
rect 484347 217020 484413 217021
rect 484347 216956 484348 217020
rect 484412 216956 484413 217020
rect 484347 216955 484413 216956
rect 484534 216341 484594 220627
rect 484531 216340 484597 216341
rect 484531 216276 484532 216340
rect 484596 216276 484597 216340
rect 484531 216275 484597 216276
rect 484718 215661 484778 221307
rect 484715 215660 484781 215661
rect 484715 215596 484716 215660
rect 484780 215596 484781 215660
rect 484715 215595 484781 215596
rect 485086 214981 485146 221443
rect 485083 214980 485149 214981
rect 485083 214916 485084 214980
rect 485148 214916 485149 214980
rect 485083 214915 485149 214916
rect 485270 214301 485330 221987
rect 485267 214300 485333 214301
rect 485267 214236 485268 214300
rect 485332 214236 485333 214300
rect 485267 214235 485333 214236
rect 483979 212940 484045 212941
rect 483979 212876 483980 212940
rect 484044 212876 484045 212940
rect 483979 212875 484045 212876
rect 485454 211581 485514 224027
rect 486187 223412 486253 223413
rect 486187 223348 486188 223412
rect 486252 223348 486253 223412
rect 486187 223347 486253 223348
rect 486003 222324 486069 222325
rect 486003 222260 486004 222324
rect 486068 222260 486069 222324
rect 486003 222259 486069 222260
rect 486006 213621 486066 222259
rect 486190 215310 486250 223347
rect 486190 215250 486434 215310
rect 486003 213620 486069 213621
rect 486003 213556 486004 213620
rect 486068 213556 486069 213620
rect 486003 213555 486069 213556
rect 486374 212261 486434 215250
rect 486371 212260 486437 212261
rect 486371 212196 486372 212260
rect 486436 212196 486437 212260
rect 486371 212195 486437 212196
rect 485451 211580 485517 211581
rect 485451 211516 485452 211580
rect 485516 211516 485517 211580
rect 485451 211515 485517 211516
rect 486558 210221 486618 224710
rect 486555 210220 486621 210221
rect 486555 210156 486556 210220
rect 486620 210156 486621 210220
rect 486555 210155 486621 210156
rect 483795 203420 483861 203421
rect 483795 203356 483796 203420
rect 483860 203356 483861 203420
rect 483795 203355 483861 203356
rect 483611 202740 483677 202741
rect 483611 202676 483612 202740
rect 483676 202676 483677 202740
rect 483611 202675 483677 202676
rect 480851 201380 480917 201381
rect 480851 201316 480852 201380
rect 480916 201316 480917 201380
rect 480851 201315 480917 201316
rect 482139 181660 482205 181661
rect 482139 181596 482140 181660
rect 482204 181596 482205 181660
rect 482139 181595 482205 181596
rect 478275 180300 478341 180301
rect 478275 180236 478276 180300
rect 478340 180236 478341 180300
rect 478275 180235 478341 180236
rect 478091 174180 478157 174181
rect 478091 174116 478092 174180
rect 478156 174116 478157 174180
rect 478091 174115 478157 174116
rect 477907 171460 477973 171461
rect 477907 171396 477908 171460
rect 477972 171396 477973 171460
rect 477907 171395 477973 171396
rect 477171 158540 477237 158541
rect 477171 158476 477172 158540
rect 477236 158476 477237 158540
rect 477171 158475 477237 158476
rect 477174 149811 477234 158475
rect 477723 152964 477789 152965
rect 477723 152900 477724 152964
rect 477788 152900 477789 152964
rect 477723 152899 477789 152900
rect 477539 152692 477605 152693
rect 477539 152628 477540 152692
rect 477604 152628 477605 152692
rect 477539 152627 477605 152628
rect 477171 149810 477237 149811
rect 477171 149746 477172 149810
rect 477236 149746 477237 149810
rect 477171 149745 477237 149746
rect 477542 143037 477602 152627
rect 477726 143309 477786 152899
rect 477910 152013 477970 171395
rect 477907 152012 477973 152013
rect 477907 151948 477908 152012
rect 477972 151948 477973 152012
rect 477907 151947 477973 151948
rect 478094 147933 478154 174115
rect 478091 147932 478157 147933
rect 478091 147868 478092 147932
rect 478156 147868 478157 147932
rect 478091 147867 478157 147868
rect 477907 147796 477973 147797
rect 477907 147732 477908 147796
rect 477972 147732 477973 147796
rect 477907 147731 477973 147732
rect 477723 143308 477789 143309
rect 477723 143244 477724 143308
rect 477788 143244 477789 143308
rect 477723 143243 477789 143244
rect 477539 143036 477605 143037
rect 477539 142972 477540 143036
rect 477604 142972 477605 143036
rect 477539 142971 477605 142972
rect 477910 140317 477970 147731
rect 478278 143853 478338 180235
rect 479379 174860 479445 174861
rect 479379 174796 479380 174860
rect 479444 174796 479445 174860
rect 479379 174795 479445 174796
rect 478643 154460 478709 154461
rect 478643 154396 478644 154460
rect 478708 154396 478709 154460
rect 478643 154395 478709 154396
rect 478646 152285 478706 154395
rect 478643 152284 478709 152285
rect 478643 152220 478644 152284
rect 478708 152220 478709 152284
rect 478643 152219 478709 152220
rect 479195 148884 479261 148885
rect 479195 148820 479196 148884
rect 479260 148820 479261 148884
rect 479195 148819 479261 148820
rect 479198 146029 479258 148819
rect 479382 147389 479442 174795
rect 479563 172820 479629 172821
rect 479563 172756 479564 172820
rect 479628 172756 479629 172820
rect 479563 172755 479629 172756
rect 479566 148749 479626 172755
rect 479747 166020 479813 166021
rect 479747 165956 479748 166020
rect 479812 165956 479813 166020
rect 479747 165955 479813 165956
rect 479750 153373 479810 165955
rect 480851 163980 480917 163981
rect 480851 163916 480852 163980
rect 480916 163916 480917 163980
rect 480851 163915 480917 163916
rect 480299 163300 480365 163301
rect 480299 163236 480300 163300
rect 480364 163236 480365 163300
rect 480299 163235 480365 163236
rect 480115 156772 480181 156773
rect 480115 156708 480116 156772
rect 480180 156708 480181 156772
rect 480115 156707 480181 156708
rect 479931 153780 479997 153781
rect 479931 153716 479932 153780
rect 479996 153716 479997 153780
rect 479931 153715 479997 153716
rect 479747 153372 479813 153373
rect 479747 153308 479748 153372
rect 479812 153308 479813 153372
rect 479747 153307 479813 153308
rect 479934 149565 479994 153715
rect 479931 149564 479997 149565
rect 479931 149500 479932 149564
rect 479996 149500 479997 149564
rect 479931 149499 479997 149500
rect 479563 148748 479629 148749
rect 479563 148684 479564 148748
rect 479628 148684 479629 148748
rect 479563 148683 479629 148684
rect 479931 148748 479997 148749
rect 479931 148684 479932 148748
rect 479996 148684 479997 148748
rect 479931 148683 479997 148684
rect 479379 147388 479445 147389
rect 479379 147324 479380 147388
rect 479444 147324 479445 147388
rect 479379 147323 479445 147324
rect 479747 146980 479813 146981
rect 479747 146916 479748 146980
rect 479812 146916 479813 146980
rect 479747 146915 479813 146916
rect 479195 146028 479261 146029
rect 479195 145964 479196 146028
rect 479260 145964 479261 146028
rect 479195 145963 479261 145964
rect 478643 144804 478709 144805
rect 478643 144740 478644 144804
rect 478708 144740 478709 144804
rect 478643 144739 478709 144740
rect 478275 143852 478341 143853
rect 478275 143788 478276 143852
rect 478340 143788 478341 143852
rect 478275 143787 478341 143788
rect 478646 140589 478706 144739
rect 478827 144260 478893 144261
rect 478827 144196 478828 144260
rect 478892 144196 478893 144260
rect 478827 144195 478893 144196
rect 478830 142765 478890 144195
rect 478827 142764 478893 142765
rect 478827 142700 478828 142764
rect 478892 142700 478893 142764
rect 478827 142699 478893 142700
rect 478643 140588 478709 140589
rect 478643 140524 478644 140588
rect 478708 140524 478709 140588
rect 478643 140523 478709 140524
rect 477907 140316 477973 140317
rect 477907 140252 477908 140316
rect 477972 140252 477973 140316
rect 477907 140251 477973 140252
rect 479750 135965 479810 146915
rect 479934 145757 479994 148683
rect 480118 146573 480178 156707
rect 480302 155277 480362 163235
rect 480483 159220 480549 159221
rect 480483 159156 480484 159220
rect 480548 159156 480549 159220
rect 480483 159155 480549 159156
rect 480299 155276 480365 155277
rect 480299 155212 480300 155276
rect 480364 155212 480365 155276
rect 480299 155211 480365 155212
rect 480486 153101 480546 159155
rect 480483 153100 480549 153101
rect 480483 153036 480484 153100
rect 480548 153036 480549 153100
rect 480483 153035 480549 153036
rect 480667 153100 480733 153101
rect 480667 153036 480668 153100
rect 480732 153036 480733 153100
rect 480667 153035 480733 153036
rect 480670 150109 480730 153035
rect 480854 151741 480914 163915
rect 481587 155956 481653 155957
rect 481587 155892 481588 155956
rect 481652 155892 481653 155956
rect 481587 155891 481653 155892
rect 480851 151740 480917 151741
rect 480851 151676 480852 151740
rect 480916 151676 480917 151740
rect 480851 151675 480917 151676
rect 480667 150108 480733 150109
rect 480667 150044 480668 150108
rect 480732 150044 480733 150108
rect 480667 150043 480733 150044
rect 480667 147116 480733 147117
rect 480667 147052 480668 147116
rect 480732 147052 480733 147116
rect 480667 147051 480733 147052
rect 480115 146572 480181 146573
rect 480115 146508 480116 146572
rect 480180 146508 480181 146572
rect 480115 146507 480181 146508
rect 479931 145756 479997 145757
rect 479931 145692 479932 145756
rect 479996 145692 479997 145756
rect 479931 145691 479997 145692
rect 480115 143580 480181 143581
rect 480115 143516 480116 143580
rect 480180 143516 480181 143580
rect 480115 143515 480181 143516
rect 480118 141677 480178 143515
rect 480483 142900 480549 142901
rect 480483 142836 480484 142900
rect 480548 142836 480549 142900
rect 480483 142835 480549 142836
rect 480299 142220 480365 142221
rect 480299 142156 480300 142220
rect 480364 142156 480365 142220
rect 480299 142155 480365 142156
rect 480115 141676 480181 141677
rect 480115 141612 480116 141676
rect 480180 141612 480181 141676
rect 480115 141611 480181 141612
rect 480302 141133 480362 142155
rect 480486 141949 480546 142835
rect 480483 141948 480549 141949
rect 480483 141884 480484 141948
rect 480548 141884 480549 141948
rect 480483 141883 480549 141884
rect 480299 141132 480365 141133
rect 480299 141068 480300 141132
rect 480364 141068 480365 141132
rect 480299 141067 480365 141068
rect 480670 137325 480730 147051
rect 481590 145213 481650 155891
rect 482142 151469 482202 181595
rect 483611 173500 483677 173501
rect 483611 173436 483612 173500
rect 483676 173436 483677 173500
rect 483611 173435 483677 173436
rect 482323 172140 482389 172141
rect 482323 172076 482324 172140
rect 482388 172076 482389 172140
rect 482323 172075 482389 172076
rect 482139 151468 482205 151469
rect 482139 151404 482140 151468
rect 482204 151404 482205 151468
rect 482139 151403 482205 151404
rect 481955 150516 482021 150517
rect 481955 150452 481956 150516
rect 482020 150452 482021 150516
rect 481955 150451 482021 150452
rect 481771 149292 481837 149293
rect 481771 149228 481772 149292
rect 481836 149228 481837 149292
rect 481771 149227 481837 149228
rect 481587 145212 481653 145213
rect 481587 145148 481588 145212
rect 481652 145148 481653 145212
rect 481587 145147 481653 145148
rect 481774 138413 481834 149227
rect 481958 144397 482018 150451
rect 482326 149429 482386 172075
rect 482507 170780 482573 170781
rect 482507 170716 482508 170780
rect 482572 170716 482573 170780
rect 482507 170715 482573 170716
rect 482510 150381 482570 170715
rect 482875 160580 482941 160581
rect 482875 160516 482876 160580
rect 482940 160516 482941 160580
rect 482875 160515 482941 160516
rect 482878 156909 482938 160515
rect 483243 159900 483309 159901
rect 483243 159836 483244 159900
rect 483308 159836 483309 159900
rect 483243 159835 483309 159836
rect 483246 157589 483306 159835
rect 483243 157588 483309 157589
rect 483243 157524 483244 157588
rect 483308 157524 483309 157588
rect 483243 157523 483309 157524
rect 483059 157452 483125 157453
rect 483059 157388 483060 157452
rect 483124 157388 483125 157452
rect 483059 157387 483125 157388
rect 482875 156908 482941 156909
rect 482875 156844 482876 156908
rect 482940 156844 482941 156908
rect 482875 156843 482941 156844
rect 482507 150380 482573 150381
rect 482507 150316 482508 150380
rect 482572 150316 482573 150380
rect 482507 150315 482573 150316
rect 482323 149428 482389 149429
rect 482323 149364 482324 149428
rect 482388 149364 482389 149428
rect 482323 149363 482389 149364
rect 482139 149156 482205 149157
rect 482139 149092 482140 149156
rect 482204 149092 482205 149156
rect 482139 149091 482205 149092
rect 481955 144396 482021 144397
rect 481955 144332 481956 144396
rect 482020 144332 482021 144396
rect 481955 144331 482021 144332
rect 482142 139229 482202 149091
rect 482323 146300 482389 146301
rect 482323 146236 482324 146300
rect 482388 146236 482389 146300
rect 482323 146235 482389 146236
rect 482139 139228 482205 139229
rect 482139 139164 482140 139228
rect 482204 139164 482205 139228
rect 482139 139163 482205 139164
rect 481771 138412 481837 138413
rect 481771 138348 481772 138412
rect 481836 138348 481837 138412
rect 481771 138347 481837 138348
rect 482326 137597 482386 146235
rect 482323 137596 482389 137597
rect 482323 137532 482324 137596
rect 482388 137532 482389 137596
rect 482323 137531 482389 137532
rect 480667 137324 480733 137325
rect 480667 137260 480668 137324
rect 480732 137260 480733 137324
rect 480667 137259 480733 137260
rect 483062 136237 483122 157387
rect 483243 155956 483309 155957
rect 483243 155892 483244 155956
rect 483308 155892 483309 155956
rect 483243 155891 483309 155892
rect 483246 145485 483306 155891
rect 483614 148477 483674 173435
rect 485267 170100 485333 170101
rect 485267 170036 485268 170100
rect 485332 170036 485333 170100
rect 485267 170035 485333 170036
rect 483795 169420 483861 169421
rect 483795 169356 483796 169420
rect 483860 169356 483861 169420
rect 483795 169355 483861 169356
rect 483798 157997 483858 169355
rect 484163 162620 484229 162621
rect 484163 162556 484164 162620
rect 484228 162556 484229 162620
rect 484163 162555 484229 162556
rect 483795 157996 483861 157997
rect 483795 157932 483796 157996
rect 483860 157932 483861 157996
rect 483795 157931 483861 157932
rect 484166 155549 484226 162555
rect 484715 161940 484781 161941
rect 484715 161876 484716 161940
rect 484780 161876 484781 161940
rect 484715 161875 484781 161876
rect 484718 156093 484778 161875
rect 484715 156092 484781 156093
rect 484715 156028 484716 156092
rect 484780 156028 484781 156092
rect 484715 156027 484781 156028
rect 485270 155957 485330 170035
rect 486003 168740 486069 168741
rect 486003 168676 486004 168740
rect 486068 168676 486069 168740
rect 486003 168675 486069 168676
rect 485451 167380 485517 167381
rect 485451 167316 485452 167380
rect 485516 167316 485517 167380
rect 485451 167315 485517 167316
rect 485267 155956 485333 155957
rect 485267 155892 485268 155956
rect 485332 155892 485333 155956
rect 485267 155891 485333 155892
rect 484347 155820 484413 155821
rect 484347 155756 484348 155820
rect 484412 155756 484413 155820
rect 484347 155755 484413 155756
rect 484163 155548 484229 155549
rect 484163 155484 484164 155548
rect 484228 155484 484229 155548
rect 484163 155483 484229 155484
rect 484350 154325 484410 155755
rect 484531 155140 484597 155141
rect 484531 155076 484532 155140
rect 484596 155076 484597 155140
rect 484531 155075 484597 155076
rect 484347 154324 484413 154325
rect 484347 154260 484348 154324
rect 484412 154260 484413 154324
rect 484347 154259 484413 154260
rect 484534 153509 484594 155075
rect 484531 153508 484597 153509
rect 484531 153444 484532 153508
rect 484596 153444 484597 153508
rect 484531 153443 484597 153444
rect 485454 152557 485514 167315
rect 485819 165340 485885 165341
rect 485819 165276 485820 165340
rect 485884 165276 485885 165340
rect 485819 165275 485885 165276
rect 485635 161260 485701 161261
rect 485635 161196 485636 161260
rect 485700 161196 485701 161260
rect 485635 161195 485701 161196
rect 485451 152556 485517 152557
rect 485451 152492 485452 152556
rect 485516 152492 485517 152556
rect 485451 152491 485517 152492
rect 484715 152420 484781 152421
rect 484715 152356 484716 152420
rect 484780 152356 484781 152420
rect 484715 152355 484781 152356
rect 484718 151197 484778 152355
rect 485638 151830 485698 161195
rect 485822 153917 485882 165275
rect 486006 156637 486066 168675
rect 486371 164660 486437 164661
rect 486371 164596 486372 164660
rect 486436 164596 486437 164660
rect 486371 164595 486437 164596
rect 486374 161490 486434 164595
rect 486190 161430 486434 161490
rect 486190 158269 486250 161430
rect 486187 158268 486253 158269
rect 486187 158204 486188 158268
rect 486252 158204 486253 158268
rect 486187 158203 486253 158204
rect 486003 156636 486069 156637
rect 486003 156572 486004 156636
rect 486068 156572 486069 156636
rect 486003 156571 486069 156572
rect 485819 153916 485885 153917
rect 485819 153852 485820 153916
rect 485884 153852 485885 153916
rect 485819 153851 485885 153852
rect 486003 153100 486069 153101
rect 486003 153036 486004 153100
rect 486068 153036 486069 153100
rect 486003 153035 486069 153036
rect 485454 151770 485698 151830
rect 484715 151196 484781 151197
rect 484715 151132 484716 151196
rect 484780 151132 484781 151196
rect 484715 151131 484781 151132
rect 483795 150516 483861 150517
rect 483795 150452 483796 150516
rect 483860 150452 483861 150516
rect 483795 150451 483861 150452
rect 483611 148476 483677 148477
rect 483611 148412 483612 148476
rect 483676 148412 483677 148476
rect 483611 148411 483677 148412
rect 483427 147796 483493 147797
rect 483427 147732 483428 147796
rect 483492 147732 483493 147796
rect 483427 147731 483493 147732
rect 483243 145484 483309 145485
rect 483243 145420 483244 145484
rect 483308 145420 483309 145484
rect 483243 145419 483309 145420
rect 483430 138957 483490 147731
rect 483611 146300 483677 146301
rect 483611 146236 483612 146300
rect 483676 146236 483677 146300
rect 483611 146235 483677 146236
rect 483427 138956 483493 138957
rect 483427 138892 483428 138956
rect 483492 138892 483493 138956
rect 483427 138891 483493 138892
rect 483614 137869 483674 146235
rect 483798 139773 483858 150451
rect 484715 150380 484781 150381
rect 484715 150316 484716 150380
rect 484780 150316 484781 150380
rect 484715 150315 484781 150316
rect 484347 149700 484413 149701
rect 484347 149636 484348 149700
rect 484412 149636 484413 149700
rect 484347 149635 484413 149636
rect 484350 148205 484410 149635
rect 484531 148340 484597 148341
rect 484531 148276 484532 148340
rect 484596 148276 484597 148340
rect 484531 148275 484597 148276
rect 484347 148204 484413 148205
rect 484347 148140 484348 148204
rect 484412 148140 484413 148204
rect 484347 148139 484413 148140
rect 484534 146709 484594 148275
rect 484531 146708 484597 146709
rect 484531 146644 484532 146708
rect 484596 146644 484597 146708
rect 484531 146643 484597 146644
rect 484531 146300 484597 146301
rect 484531 146236 484532 146300
rect 484596 146236 484597 146300
rect 484531 146235 484597 146236
rect 484347 145620 484413 145621
rect 484347 145556 484348 145620
rect 484412 145556 484413 145620
rect 484347 145555 484413 145556
rect 484350 143717 484410 145555
rect 484534 144125 484594 146235
rect 484531 144124 484597 144125
rect 484531 144060 484532 144124
rect 484596 144060 484597 144124
rect 484531 144059 484597 144060
rect 484347 143716 484413 143717
rect 484347 143652 484348 143716
rect 484412 143652 484413 143716
rect 484347 143651 484413 143652
rect 484718 142493 484778 150315
rect 485454 149021 485514 151770
rect 485451 149020 485517 149021
rect 485451 148956 485452 149020
rect 485516 148956 485517 149020
rect 485451 148955 485517 148956
rect 485635 149020 485701 149021
rect 485635 148956 485636 149020
rect 485700 148956 485701 149020
rect 485635 148955 485701 148956
rect 484715 142492 484781 142493
rect 484715 142428 484716 142492
rect 484780 142428 484781 142492
rect 484715 142427 484781 142428
rect 483795 139772 483861 139773
rect 483795 139708 483796 139772
rect 483860 139708 483861 139772
rect 483795 139707 483861 139708
rect 484531 138820 484597 138821
rect 484531 138756 484532 138820
rect 484596 138756 484597 138820
rect 484531 138755 484597 138756
rect 483611 137868 483677 137869
rect 483611 137804 483612 137868
rect 483676 137804 483677 137868
rect 483611 137803 483677 137804
rect 484347 137460 484413 137461
rect 484347 137396 484348 137460
rect 484412 137396 484413 137460
rect 484347 137395 484413 137396
rect 484350 136509 484410 137395
rect 484534 137053 484594 138755
rect 485638 138685 485698 148955
rect 486006 142357 486066 153035
rect 486003 142356 486069 142357
rect 486003 142292 486004 142356
rect 486068 142292 486069 142356
rect 486003 142291 486069 142292
rect 485635 138684 485701 138685
rect 485635 138620 485636 138684
rect 485700 138620 485701 138684
rect 485635 138619 485701 138620
rect 484531 137052 484597 137053
rect 484531 136988 484532 137052
rect 484596 136988 484597 137052
rect 484531 136987 484597 136988
rect 484347 136508 484413 136509
rect 484347 136444 484348 136508
rect 484412 136444 484413 136508
rect 484347 136443 484413 136444
rect 483059 136236 483125 136237
rect 483059 136172 483060 136236
rect 483124 136172 483125 136236
rect 483059 136171 483125 136172
rect 479747 135964 479813 135965
rect 479747 135900 479748 135964
rect 479812 135900 479813 135964
rect 479747 135899 479813 135900
rect 485819 134468 485885 134469
rect 485819 134404 485820 134468
rect 485884 134404 485885 134468
rect 485819 134403 485885 134404
rect 478275 133652 478341 133653
rect 478275 133588 478276 133652
rect 478340 133588 478341 133652
rect 478275 133587 478341 133588
rect 478091 133108 478157 133109
rect 478091 133044 478092 133108
rect 478156 133044 478157 133108
rect 478091 133043 478157 133044
rect 477355 132346 477421 132347
rect 477355 132282 477356 132346
rect 477420 132282 477421 132346
rect 477355 132281 477421 132282
rect 477358 123861 477418 132281
rect 477355 123860 477421 123861
rect 477355 123796 477356 123860
rect 477420 123796 477421 123860
rect 477355 123795 477421 123796
rect 478094 122501 478154 133043
rect 478091 122500 478157 122501
rect 478091 122436 478092 122500
rect 478156 122436 478157 122500
rect 478091 122435 478157 122436
rect 478278 121821 478338 133587
rect 485822 132970 485882 134403
rect 486003 133924 486069 133925
rect 486003 133860 486004 133924
rect 486068 133860 486069 133924
rect 486003 133859 486069 133860
rect 486006 133650 486066 133859
rect 486006 133590 486434 133650
rect 485822 132910 486250 132970
rect 486003 132564 486069 132565
rect 486003 132500 486004 132564
rect 486068 132500 486069 132564
rect 486003 132499 486069 132500
rect 481403 131748 481469 131749
rect 481403 131684 481404 131748
rect 481468 131684 481469 131748
rect 481403 131683 481469 131684
rect 478827 129572 478893 129573
rect 478827 129508 478828 129572
rect 478892 129508 478893 129572
rect 478827 129507 478893 129508
rect 478830 127941 478890 129507
rect 478827 127940 478893 127941
rect 478827 127876 478828 127940
rect 478892 127876 478893 127940
rect 478827 127875 478893 127876
rect 481406 124541 481466 131683
rect 481587 131204 481653 131205
rect 481587 131140 481588 131204
rect 481652 131140 481653 131204
rect 481587 131139 481653 131140
rect 481590 125221 481650 131139
rect 484531 131068 484597 131069
rect 484531 131004 484532 131068
rect 484596 131004 484597 131068
rect 484531 131003 484597 131004
rect 484347 130388 484413 130389
rect 484347 130324 484348 130388
rect 484412 130324 484413 130388
rect 484347 130323 484413 130324
rect 483059 129980 483125 129981
rect 483059 129916 483060 129980
rect 483124 129916 483125 129980
rect 483059 129915 483125 129916
rect 483062 127261 483122 129915
rect 483795 128484 483861 128485
rect 483795 128420 483796 128484
rect 483860 128420 483861 128484
rect 483795 128419 483861 128420
rect 483059 127260 483125 127261
rect 483059 127196 483060 127260
rect 483124 127196 483125 127260
rect 483059 127195 483125 127196
rect 481587 125220 481653 125221
rect 481587 125156 481588 125220
rect 481652 125156 481653 125220
rect 481587 125155 481653 125156
rect 481403 124540 481469 124541
rect 481403 124476 481404 124540
rect 481468 124476 481469 124540
rect 481403 124475 481469 124476
rect 478275 121820 478341 121821
rect 478275 121756 478276 121820
rect 478340 121756 478341 121820
rect 478275 121755 478341 121756
rect 483798 119101 483858 128419
rect 484350 126581 484410 130323
rect 484347 126580 484413 126581
rect 484347 126516 484348 126580
rect 484412 126516 484413 126580
rect 484347 126515 484413 126516
rect 484534 125901 484594 131003
rect 484531 125900 484597 125901
rect 484531 125836 484532 125900
rect 484596 125836 484597 125900
rect 484531 125835 484597 125836
rect 486006 123181 486066 132499
rect 486003 123180 486069 123181
rect 486003 123116 486004 123180
rect 486068 123116 486069 123180
rect 486003 123115 486069 123116
rect 486190 120730 486250 132910
rect 486374 121141 486434 133590
rect 486371 121140 486437 121141
rect 486371 121076 486372 121140
rect 486436 121076 486437 121140
rect 486371 121075 486437 121076
rect 486190 120670 486434 120730
rect 486374 120461 486434 120670
rect 486371 120460 486437 120461
rect 486371 120396 486372 120460
rect 486436 120396 486437 120460
rect 486371 120395 486437 120396
rect 483795 119100 483861 119101
rect 483795 119036 483796 119100
rect 483860 119036 483861 119100
rect 483795 119035 483861 119036
rect 480851 86460 480917 86461
rect 480851 86396 480852 86460
rect 480916 86396 480917 86460
rect 480851 86395 480917 86396
rect 478091 83740 478157 83741
rect 478091 83676 478092 83740
rect 478156 83676 478157 83740
rect 478091 83675 478157 83676
rect 477355 65380 477421 65381
rect 477355 65316 477356 65380
rect 477420 65316 477421 65380
rect 477355 65315 477421 65316
rect 477171 63204 477237 63205
rect 477171 63140 477172 63204
rect 477236 63140 477237 63204
rect 477171 63139 477237 63140
rect 477174 60349 477234 63139
rect 477358 62525 477418 65315
rect 477355 62524 477421 62525
rect 477355 62460 477356 62524
rect 477420 62460 477421 62524
rect 477355 62459 477421 62460
rect 477907 60620 477973 60621
rect 477907 60556 477908 60620
rect 477972 60556 477973 60620
rect 477907 60555 477973 60556
rect 477171 60348 477237 60349
rect 477171 60284 477172 60348
rect 477236 60284 477237 60348
rect 477171 60283 477237 60284
rect 477910 57629 477970 60555
rect 478094 58173 478154 83675
rect 478275 83060 478341 83061
rect 478275 82996 478276 83060
rect 478340 82996 478341 83060
rect 478275 82995 478341 82996
rect 478278 58717 478338 82995
rect 478459 81700 478525 81701
rect 478459 81636 478460 81700
rect 478524 81636 478525 81700
rect 478459 81635 478525 81636
rect 478462 59533 478522 81635
rect 479563 78980 479629 78981
rect 479563 78916 479564 78980
rect 479628 78916 479629 78980
rect 479563 78915 479629 78916
rect 479379 77620 479445 77621
rect 479379 77556 479380 77620
rect 479444 77556 479445 77620
rect 479379 77555 479445 77556
rect 478643 68100 478709 68101
rect 478643 68036 478644 68100
rect 478708 68036 478709 68100
rect 478643 68035 478709 68036
rect 478646 65245 478706 68035
rect 478643 65244 478709 65245
rect 478643 65180 478644 65244
rect 478708 65180 478709 65244
rect 478643 65179 478709 65180
rect 478643 63748 478709 63749
rect 478643 63684 478644 63748
rect 478708 63684 478709 63748
rect 478643 63683 478709 63684
rect 478459 59532 478525 59533
rect 478459 59468 478460 59532
rect 478524 59468 478525 59532
rect 478459 59467 478525 59468
rect 478275 58716 478341 58717
rect 478275 58652 478276 58716
rect 478340 58652 478341 58716
rect 478275 58651 478341 58652
rect 478091 58172 478157 58173
rect 478091 58108 478092 58172
rect 478156 58108 478157 58172
rect 478091 58107 478157 58108
rect 477907 57628 477973 57629
rect 477907 57564 477908 57628
rect 477972 57564 477973 57628
rect 477907 57563 477973 57564
rect 478646 57357 478706 63683
rect 479382 61437 479442 77555
rect 479566 65517 479626 78915
rect 479747 75580 479813 75581
rect 479747 75516 479748 75580
rect 479812 75516 479813 75580
rect 479747 75515 479813 75516
rect 479563 65516 479629 65517
rect 479563 65452 479564 65516
rect 479628 65452 479629 65516
rect 479563 65451 479629 65452
rect 479750 63613 479810 75515
rect 479931 74220 479997 74221
rect 479931 74156 479932 74220
rect 479996 74156 479997 74220
rect 479931 74155 479997 74156
rect 479934 64429 479994 74155
rect 480299 67556 480365 67557
rect 480299 67492 480300 67556
rect 480364 67492 480365 67556
rect 480299 67491 480365 67492
rect 480115 66196 480181 66197
rect 480115 66132 480116 66196
rect 480180 66132 480181 66196
rect 480115 66131 480181 66132
rect 479931 64428 479997 64429
rect 479931 64364 479932 64428
rect 479996 64364 479997 64428
rect 479931 64363 479997 64364
rect 479747 63612 479813 63613
rect 479747 63548 479748 63612
rect 479812 63548 479813 63612
rect 479747 63547 479813 63548
rect 480118 61981 480178 66131
rect 480115 61980 480181 61981
rect 480115 61916 480116 61980
rect 480180 61916 480181 61980
rect 480115 61915 480181 61916
rect 479379 61436 479445 61437
rect 479379 61372 479380 61436
rect 479444 61372 479445 61436
rect 479379 61371 479445 61372
rect 478643 57356 478709 57357
rect 478643 57292 478644 57356
rect 478708 57292 478709 57356
rect 478643 57291 478709 57292
rect 480302 54909 480362 67491
rect 480483 62252 480549 62253
rect 480483 62188 480484 62252
rect 480548 62188 480549 62252
rect 480483 62187 480549 62188
rect 480299 54908 480365 54909
rect 480299 54844 480300 54908
rect 480364 54844 480365 54908
rect 480299 54843 480365 54844
rect 480486 53549 480546 62187
rect 480854 56269 480914 86395
rect 483611 85780 483677 85781
rect 483611 85716 483612 85780
rect 483676 85716 483677 85780
rect 483611 85715 483677 85716
rect 482139 82380 482205 82381
rect 482139 82316 482140 82380
rect 482204 82316 482205 82380
rect 482139 82315 482205 82316
rect 481035 76940 481101 76941
rect 481035 76876 481036 76940
rect 481100 76876 481101 76940
rect 481035 76875 481101 76876
rect 481038 62797 481098 76875
rect 481403 72860 481469 72861
rect 481403 72796 481404 72860
rect 481468 72796 481469 72860
rect 481403 72795 481469 72796
rect 481406 68237 481466 72795
rect 481587 69460 481653 69461
rect 481587 69396 481588 69460
rect 481652 69396 481653 69460
rect 481587 69395 481653 69396
rect 481403 68236 481469 68237
rect 481403 68172 481404 68236
rect 481468 68172 481469 68236
rect 481403 68171 481469 68172
rect 481590 67693 481650 69395
rect 481587 67692 481653 67693
rect 481587 67628 481588 67692
rect 481652 67628 481653 67692
rect 481587 67627 481653 67628
rect 481587 67556 481653 67557
rect 481587 67492 481588 67556
rect 481652 67492 481653 67556
rect 481587 67491 481653 67492
rect 481590 62930 481650 67491
rect 481771 67420 481837 67421
rect 481771 67356 481772 67420
rect 481836 67356 481837 67420
rect 481771 67355 481837 67356
rect 481774 64701 481834 67355
rect 481771 64700 481837 64701
rect 481771 64636 481772 64700
rect 481836 64636 481837 64700
rect 481771 64635 481837 64636
rect 481590 62870 482018 62930
rect 481035 62796 481101 62797
rect 481035 62732 481036 62796
rect 481100 62732 481101 62796
rect 481035 62731 481101 62732
rect 481771 62252 481837 62253
rect 481771 62188 481772 62252
rect 481836 62188 481837 62252
rect 481771 62187 481837 62188
rect 481587 61980 481653 61981
rect 481587 61916 481588 61980
rect 481652 61916 481653 61980
rect 481587 61915 481653 61916
rect 481590 60485 481650 61915
rect 481587 60484 481653 60485
rect 481587 60420 481588 60484
rect 481652 60420 481653 60484
rect 481587 60419 481653 60420
rect 480851 56268 480917 56269
rect 480851 56204 480852 56268
rect 480916 56204 480917 56268
rect 480851 56203 480917 56204
rect 481774 54637 481834 62187
rect 481958 55997 482018 62870
rect 482142 58989 482202 82315
rect 482323 76260 482389 76261
rect 482323 76196 482324 76260
rect 482388 76196 482389 76260
rect 482323 76195 482389 76196
rect 482326 63069 482386 76195
rect 483427 70140 483493 70141
rect 483427 70076 483428 70140
rect 483492 70076 483493 70140
rect 483427 70075 483493 70076
rect 483243 68780 483309 68781
rect 483243 68716 483244 68780
rect 483308 68716 483309 68780
rect 483243 68715 483309 68716
rect 483059 67556 483125 67557
rect 483059 67492 483060 67556
rect 483124 67492 483125 67556
rect 483059 67491 483125 67492
rect 482323 63068 482389 63069
rect 482323 63004 482324 63068
rect 482388 63004 482389 63068
rect 482323 63003 482389 63004
rect 482139 58988 482205 58989
rect 482139 58924 482140 58988
rect 482204 58924 482205 58988
rect 482139 58923 482205 58924
rect 481955 55996 482021 55997
rect 481955 55932 481956 55996
rect 482020 55932 482021 55996
rect 481955 55931 482021 55932
rect 483062 55453 483122 67491
rect 483246 67285 483306 68715
rect 483243 67284 483309 67285
rect 483243 67220 483244 67284
rect 483308 67220 483309 67284
rect 483243 67219 483309 67220
rect 483430 67149 483490 70075
rect 483427 67148 483493 67149
rect 483427 67084 483428 67148
rect 483492 67084 483493 67148
rect 483427 67083 483493 67084
rect 483243 66740 483309 66741
rect 483243 66676 483244 66740
rect 483308 66676 483309 66740
rect 483243 66675 483309 66676
rect 483246 66061 483306 66675
rect 483243 66060 483309 66061
rect 483243 65996 483244 66060
rect 483308 65996 483309 66060
rect 483243 65995 483309 65996
rect 483243 65924 483309 65925
rect 483243 65860 483244 65924
rect 483308 65860 483309 65924
rect 483243 65859 483309 65860
rect 483059 55452 483125 55453
rect 483059 55388 483060 55452
rect 483124 55388 483125 55452
rect 483059 55387 483125 55388
rect 481771 54636 481837 54637
rect 481771 54572 481772 54636
rect 481836 54572 481837 54636
rect 481771 54571 481837 54572
rect 483246 54093 483306 65859
rect 483427 62660 483493 62661
rect 483427 62596 483428 62660
rect 483492 62596 483493 62660
rect 483427 62595 483493 62596
rect 483430 60893 483490 62595
rect 483427 60892 483493 60893
rect 483427 60828 483428 60892
rect 483492 60828 483493 60892
rect 483427 60827 483493 60828
rect 483614 56813 483674 85715
rect 485819 80340 485885 80341
rect 485819 80276 485820 80340
rect 485884 80276 485885 80340
rect 485819 80275 485885 80276
rect 484347 74900 484413 74901
rect 484347 74836 484348 74900
rect 484412 74836 484413 74900
rect 484347 74835 484413 74836
rect 484350 74550 484410 74835
rect 484166 74490 484410 74550
rect 484166 67965 484226 74490
rect 484899 73540 484965 73541
rect 484899 73476 484900 73540
rect 484964 73476 484965 73540
rect 484899 73475 484965 73476
rect 484715 72180 484781 72181
rect 484715 72116 484716 72180
rect 484780 72116 484781 72180
rect 484715 72115 484781 72116
rect 484531 71500 484597 71501
rect 484531 71436 484532 71500
rect 484596 71436 484597 71500
rect 484531 71435 484597 71436
rect 484347 70820 484413 70821
rect 484347 70756 484348 70820
rect 484412 70756 484413 70820
rect 484347 70755 484413 70756
rect 484163 67964 484229 67965
rect 484163 67900 484164 67964
rect 484228 67900 484229 67964
rect 484163 67899 484229 67900
rect 484350 66877 484410 70755
rect 484347 66876 484413 66877
rect 484347 66812 484348 66876
rect 484412 66812 484413 66876
rect 484347 66811 484413 66812
rect 484534 66333 484594 71435
rect 484531 66332 484597 66333
rect 484531 66268 484532 66332
rect 484596 66268 484597 66332
rect 484531 66267 484597 66268
rect 484163 66060 484229 66061
rect 484163 65996 484164 66060
rect 484228 65996 484229 66060
rect 484163 65995 484229 65996
rect 484166 64157 484226 65995
rect 484718 65789 484778 72115
rect 484715 65788 484781 65789
rect 484715 65724 484716 65788
rect 484780 65724 484781 65788
rect 484715 65723 484781 65724
rect 484902 64973 484962 73475
rect 484899 64972 484965 64973
rect 484899 64908 484900 64972
rect 484964 64908 484965 64972
rect 484899 64907 484965 64908
rect 485822 64890 485882 80275
rect 486555 78300 486621 78301
rect 486555 78236 486556 78300
rect 486620 78236 486621 78300
rect 486555 78235 486621 78236
rect 486558 74550 486618 78235
rect 486190 74490 486618 74550
rect 486190 66469 486250 74490
rect 486187 66468 486253 66469
rect 486187 66404 486188 66468
rect 486252 66404 486253 66468
rect 486187 66403 486253 66404
rect 485270 64830 485882 64890
rect 484347 64700 484413 64701
rect 484347 64636 484348 64700
rect 484412 64636 484413 64700
rect 484347 64635 484413 64636
rect 484163 64156 484229 64157
rect 484163 64092 484164 64156
rect 484228 64092 484229 64156
rect 484163 64091 484229 64092
rect 484350 61709 484410 64635
rect 485270 62389 485330 64830
rect 485267 62388 485333 62389
rect 485267 62324 485268 62388
rect 485332 62324 485333 62388
rect 485267 62323 485333 62324
rect 484347 61708 484413 61709
rect 484347 61644 484348 61708
rect 484412 61644 484413 61708
rect 484347 61643 484413 61644
rect 483611 56812 483677 56813
rect 483611 56748 483612 56812
rect 483676 56748 483677 56812
rect 483611 56747 483677 56748
rect 483243 54092 483309 54093
rect 483243 54028 483244 54092
rect 483308 54028 483309 54092
rect 483243 54027 483309 54028
rect 480483 53548 480549 53549
rect 480483 53484 480484 53548
rect 480548 53484 480549 53548
rect 480483 53483 480549 53484
rect 483059 53004 483125 53005
rect 483059 52940 483060 53004
rect 483124 52940 483125 53004
rect 483059 52939 483125 52940
rect 480851 52460 480917 52461
rect 480851 52396 480852 52460
rect 480916 52396 480917 52460
rect 480851 52395 480917 52396
rect 480854 48245 480914 52395
rect 481771 51644 481837 51645
rect 481771 51580 481772 51644
rect 481836 51580 481837 51644
rect 481771 51579 481837 51580
rect 481587 50828 481653 50829
rect 481587 50764 481588 50828
rect 481652 50764 481653 50828
rect 481587 50763 481653 50764
rect 481035 50284 481101 50285
rect 481035 50220 481036 50284
rect 481100 50220 481101 50284
rect 481035 50219 481101 50220
rect 480851 48244 480917 48245
rect 480851 48180 480852 48244
rect 480916 48180 480917 48244
rect 480851 48179 480917 48180
rect 480851 47564 480917 47565
rect 480851 47500 480852 47564
rect 480916 47500 480917 47564
rect 480851 47499 480917 47500
rect 479931 47428 479997 47429
rect 479931 47364 479932 47428
rect 479996 47364 479997 47428
rect 479931 47363 479997 47364
rect 479195 46748 479261 46749
rect 479195 46684 479196 46748
rect 479260 46684 479261 46748
rect 479195 46683 479261 46684
rect 478091 43484 478157 43485
rect 478091 43420 478092 43484
rect 478156 43420 478157 43484
rect 478091 43419 478157 43420
rect 476907 41512 476973 41513
rect 476907 41448 476908 41512
rect 476972 41448 476973 41512
rect 476907 41447 476973 41448
rect 476910 41170 476970 41447
rect 476910 41110 477050 41170
rect 476990 34781 477050 41110
rect 476987 34780 477053 34781
rect 476987 34716 476988 34780
rect 477052 34716 477053 34780
rect 476987 34715 477053 34716
rect 478094 32061 478154 43419
rect 478275 42668 478341 42669
rect 478275 42604 478276 42668
rect 478340 42604 478341 42668
rect 478275 42603 478341 42604
rect 478278 33421 478338 42603
rect 479198 39949 479258 46683
rect 479563 46204 479629 46205
rect 479563 46140 479564 46204
rect 479628 46140 479629 46204
rect 479563 46139 479629 46140
rect 479379 45660 479445 45661
rect 479379 45596 479380 45660
rect 479444 45596 479445 45660
rect 479379 45595 479445 45596
rect 479195 39948 479261 39949
rect 479195 39884 479196 39948
rect 479260 39884 479261 39948
rect 479195 39883 479261 39884
rect 478275 33420 478341 33421
rect 478275 33356 478276 33420
rect 478340 33356 478341 33420
rect 478275 33355 478341 33356
rect 478091 32060 478157 32061
rect 478091 31996 478092 32060
rect 478156 31996 478157 32060
rect 478091 31995 478157 31996
rect 479382 28661 479442 45595
rect 479379 28660 479445 28661
rect 479379 28596 479380 28660
rect 479444 28596 479445 28660
rect 479379 28595 479445 28596
rect 479566 27981 479626 46139
rect 479747 45388 479813 45389
rect 479747 45324 479748 45388
rect 479812 45324 479813 45388
rect 479747 45323 479813 45324
rect 479750 29341 479810 45323
rect 479934 44437 479994 47363
rect 479931 44436 479997 44437
rect 479931 44372 479932 44436
rect 479996 44372 479997 44436
rect 479931 44371 479997 44372
rect 479747 29340 479813 29341
rect 479747 29276 479748 29340
rect 479812 29276 479813 29340
rect 479747 29275 479813 29276
rect 479563 27980 479629 27981
rect 479563 27916 479564 27980
rect 479628 27916 479629 27980
rect 479563 27915 479629 27916
rect 480854 17101 480914 47499
rect 481038 21861 481098 50219
rect 481219 48924 481285 48925
rect 481219 48860 481220 48924
rect 481284 48860 481285 48924
rect 481219 48859 481285 48860
rect 481222 23901 481282 48859
rect 481403 48108 481469 48109
rect 481403 48044 481404 48108
rect 481468 48044 481469 48108
rect 481403 48043 481469 48044
rect 481406 25261 481466 48043
rect 481590 39949 481650 50763
rect 481774 41445 481834 51579
rect 483062 51370 483122 52939
rect 483243 52188 483309 52189
rect 483243 52124 483244 52188
rect 483308 52124 483309 52188
rect 483243 52123 483309 52124
rect 482878 51310 483122 51370
rect 482878 50010 482938 51310
rect 482878 49950 483122 50010
rect 482139 49740 482205 49741
rect 482139 49676 482140 49740
rect 482204 49676 482205 49740
rect 482139 49675 482205 49676
rect 481771 41444 481837 41445
rect 481771 41380 481772 41444
rect 481836 41380 481837 41444
rect 481771 41379 481837 41380
rect 481587 39948 481653 39949
rect 481587 39884 481588 39948
rect 481652 39884 481653 39948
rect 481587 39883 481653 39884
rect 481403 25260 481469 25261
rect 481403 25196 481404 25260
rect 481468 25196 481469 25260
rect 481403 25195 481469 25196
rect 481219 23900 481285 23901
rect 481219 23836 481220 23900
rect 481284 23836 481285 23900
rect 481219 23835 481285 23836
rect 482142 22541 482202 49675
rect 482323 48380 482389 48381
rect 482323 48316 482324 48380
rect 482388 48316 482389 48380
rect 482323 48315 482389 48316
rect 482326 24581 482386 48315
rect 483062 43349 483122 49950
rect 483059 43348 483125 43349
rect 483059 43284 483060 43348
rect 483124 43284 483125 43348
rect 483059 43283 483125 43284
rect 483246 41445 483306 52123
rect 483611 50964 483677 50965
rect 483611 50900 483612 50964
rect 483676 50900 483677 50964
rect 483611 50899 483677 50900
rect 483243 41444 483309 41445
rect 483243 41380 483244 41444
rect 483308 41380 483309 41444
rect 483243 41379 483309 41380
rect 482323 24580 482389 24581
rect 482323 24516 482324 24580
rect 482388 24516 482389 24580
rect 482323 24515 482389 24516
rect 482139 22540 482205 22541
rect 482139 22476 482140 22540
rect 482204 22476 482205 22540
rect 482139 22475 482205 22476
rect 481035 21860 481101 21861
rect 481035 21796 481036 21860
rect 481100 21796 481101 21860
rect 481035 21795 481101 21796
rect 483614 20501 483674 50899
rect 483795 49468 483861 49469
rect 483795 49404 483796 49468
rect 483860 49404 483861 49468
rect 483795 49403 483861 49404
rect 483798 23221 483858 49403
rect 485635 44028 485701 44029
rect 485635 43964 485636 44028
rect 485700 43964 485701 44028
rect 485635 43963 485701 43964
rect 485451 41308 485517 41309
rect 485451 41244 485452 41308
rect 485516 41244 485517 41308
rect 485451 41243 485517 41244
rect 484899 40764 484965 40765
rect 484899 40700 484900 40764
rect 484964 40700 484965 40764
rect 484899 40699 484965 40700
rect 484715 40084 484781 40085
rect 484715 40020 484716 40084
rect 484780 40020 484781 40084
rect 484715 40019 484781 40020
rect 484531 39812 484597 39813
rect 484531 39748 484532 39812
rect 484596 39748 484597 39812
rect 484531 39747 484597 39748
rect 484347 39268 484413 39269
rect 484347 39204 484348 39268
rect 484412 39204 484413 39268
rect 484347 39203 484413 39204
rect 484350 38181 484410 39203
rect 484347 38180 484413 38181
rect 484347 38116 484348 38180
rect 484412 38116 484413 38180
rect 484347 38115 484413 38116
rect 484534 37501 484594 39747
rect 484531 37500 484597 37501
rect 484531 37436 484532 37500
rect 484596 37436 484597 37500
rect 484531 37435 484597 37436
rect 484718 36821 484778 40019
rect 484715 36820 484781 36821
rect 484715 36756 484716 36820
rect 484780 36756 484781 36820
rect 484715 36755 484781 36756
rect 484902 36141 484962 40699
rect 485083 38724 485149 38725
rect 485083 38660 485084 38724
rect 485148 38660 485149 38724
rect 485083 38659 485149 38660
rect 484899 36140 484965 36141
rect 484899 36076 484900 36140
rect 484964 36076 484965 36140
rect 484899 36075 484965 36076
rect 485086 26250 485146 38659
rect 485454 35461 485514 41243
rect 485451 35460 485517 35461
rect 485451 35396 485452 35460
rect 485516 35396 485517 35460
rect 485451 35395 485517 35396
rect 485638 31381 485698 43963
rect 486003 43076 486069 43077
rect 486003 43012 486004 43076
rect 486068 43012 486069 43076
rect 486003 43011 486069 43012
rect 486006 42530 486066 43011
rect 486006 42470 486250 42530
rect 486003 42124 486069 42125
rect 486003 42060 486004 42124
rect 486068 42060 486069 42124
rect 486003 42059 486069 42060
rect 486006 34101 486066 42059
rect 486190 35910 486250 42470
rect 486190 35850 486434 35910
rect 486003 34100 486069 34101
rect 486003 34036 486004 34100
rect 486068 34036 486069 34100
rect 486003 34035 486069 34036
rect 486374 32741 486434 35850
rect 486371 32740 486437 32741
rect 486371 32676 486372 32740
rect 486436 32676 486437 32740
rect 486371 32675 486437 32676
rect 485635 31380 485701 31381
rect 485635 31316 485636 31380
rect 485700 31316 485701 31380
rect 485635 31315 485701 31316
rect 484902 26190 485146 26250
rect 484902 25941 484962 26190
rect 484899 25940 484965 25941
rect 484899 25876 484900 25940
rect 484964 25876 484965 25940
rect 484899 25875 484965 25876
rect 483795 23220 483861 23221
rect 483795 23156 483796 23220
rect 483860 23156 483861 23220
rect 483795 23155 483861 23156
rect 483611 20500 483677 20501
rect 483611 20436 483612 20500
rect 483676 20436 483677 20500
rect 483611 20435 483677 20436
rect 480851 17100 480917 17101
rect 480851 17036 480852 17100
rect 480916 17036 480917 17100
rect 480851 17035 480917 17036
rect 20299 236 20365 237
rect 20299 172 20300 236
rect 20364 172 20365 236
rect 20299 171 20365 172
use W_IO  Tile_X0Y1_W_IO
timestamp 0
transform 1 0 10000 0 1 692250
box 0 0 1 1
use W_IO  Tile_X0Y2_W_IO
timestamp 0
transform 1 0 10000 0 1 647250
box 0 0 1 1
use W_IO  Tile_X0Y3_W_IO
timestamp 0
transform 1 0 10000 0 1 602250
box 0 0 1 1
use W_IO  Tile_X0Y4_W_IO
timestamp 0
transform 1 0 10000 0 1 557250
box 0 0 1 1
use W_IO  Tile_X0Y5_W_IO
timestamp 0
transform 1 0 10000 0 1 512250
box 0 0 1 1
use W_IO  Tile_X0Y6_W_IO
timestamp 0
transform 1 0 10000 0 1 467250
box 0 0 1 1
use W_IO  Tile_X0Y7_W_IO
timestamp 0
transform 1 0 10000 0 1 422250
box 0 0 1 1
use W_IO  Tile_X0Y8_W_IO
timestamp 0
transform 1 0 10000 0 1 377250
box 0 0 1 1
use W_IO  Tile_X0Y9_W_IO
timestamp 0
transform 1 0 10000 0 1 332250
box 0 0 1 1
use W_IO  Tile_X0Y10_W_IO
timestamp 0
transform 1 0 10000 0 1 287250
box 0 0 1 1
use W_IO  Tile_X0Y11_W_IO
timestamp 0
transform 1 0 10000 0 1 242250
box 0 0 1 1
use W_IO  Tile_X0Y12_W_IO
timestamp 0
transform 1 0 10000 0 1 197250
box 0 0 1 1
use W_IO  Tile_X0Y13_W_IO
timestamp 0
transform 1 0 10000 0 1 152250
box 0 0 1 1
use W_IO  Tile_X0Y14_W_IO
timestamp 0
transform 1 0 10000 0 1 107250
box 0 0 1 1
use W_IO  Tile_X0Y15_W_IO
timestamp 0
transform 1 0 10000 0 1 62250
box 0 0 1 1
use W_IO  Tile_X0Y16_W_IO
timestamp 0
transform 1 0 10000 0 1 17250
box 0 0 1 1
use N_IO  Tile_X1Y0_N_IO
timestamp 0
transform 1 0 21250 0 1 737250
box 0 0 1 1
use LUT4AB  Tile_X1Y1_LUT4AB
timestamp 0
transform 1 0 21250 0 1 692250
box 0 0 1 1
use LUT4AB  Tile_X1Y2_LUT4AB
timestamp 0
transform 1 0 21250 0 1 647250
box 0 0 1 1
use LUT4AB  Tile_X1Y3_LUT4AB
timestamp 0
transform 1 0 21250 0 1 602250
box 0 0 1 1
use LUT4AB  Tile_X1Y4_LUT4AB
timestamp 0
transform 1 0 21250 0 1 557250
box 0 0 1 1
use LUT4AB  Tile_X1Y5_LUT4AB
timestamp 0
transform 1 0 21250 0 1 512250
box 0 0 1 1
use LUT4AB  Tile_X1Y6_LUT4AB
timestamp 0
transform 1 0 21250 0 1 467250
box 0 0 1 1
use LUT4AB  Tile_X1Y7_LUT4AB
timestamp 0
transform 1 0 21250 0 1 422250
box 0 0 1 1
use LUT4AB  Tile_X1Y8_LUT4AB
timestamp 0
transform 1 0 21250 0 1 377250
box 0 0 1 1
use LUT4AB  Tile_X1Y9_LUT4AB
timestamp 0
transform 1 0 21250 0 1 332250
box 0 0 1 1
use LUT4AB  Tile_X1Y10_LUT4AB
timestamp 0
transform 1 0 21250 0 1 287250
box 0 0 1 1
use LUT4AB  Tile_X1Y11_LUT4AB
timestamp 0
transform 1 0 21250 0 1 242250
box 0 0 1 1
use LUT4AB  Tile_X1Y12_LUT4AB
timestamp 0
transform 1 0 21250 0 1 197250
box 0 0 1 1
use LUT4AB  Tile_X1Y13_LUT4AB
timestamp 0
transform 1 0 21250 0 1 152250
box 0 0 1 1
use LUT4AB  Tile_X1Y14_LUT4AB
timestamp 0
transform 1 0 21250 0 1 107250
box 0 0 1 1
use LUT4AB  Tile_X1Y15_LUT4AB
timestamp 0
transform 1 0 21250 0 1 62250
box 0 0 1 1
use LUT4AB  Tile_X1Y16_LUT4AB
timestamp 0
transform 1 0 21250 0 1 17250
box 0 0 1 1
use S_CPU_IRQ  Tile_X1Y17_S_CPU_IRQ
timestamp 0
transform 1 0 21250 0 1 6000
box 0 0 1 1
use N_IO  Tile_X2Y0_N_IO
timestamp 0
transform 1 0 62250 0 1 737250
box 0 0 1 1
use LUT4AB  Tile_X2Y1_LUT4AB
timestamp 0
transform 1 0 62250 0 1 692250
box 0 0 1 1
use LUT4AB  Tile_X2Y2_LUT4AB
timestamp 0
transform 1 0 62250 0 1 647250
box 0 0 1 1
use LUT4AB  Tile_X2Y3_LUT4AB
timestamp 0
transform 1 0 62250 0 1 602250
box 0 0 1 1
use LUT4AB  Tile_X2Y4_LUT4AB
timestamp 0
transform 1 0 62250 0 1 557250
box 0 0 1 1
use LUT4AB  Tile_X2Y5_LUT4AB
timestamp 0
transform 1 0 62250 0 1 512250
box 0 0 1 1
use LUT4AB  Tile_X2Y6_LUT4AB
timestamp 0
transform 1 0 62250 0 1 467250
box 0 0 1 1
use LUT4AB  Tile_X2Y7_LUT4AB
timestamp 0
transform 1 0 62250 0 1 422250
box 0 0 1 1
use LUT4AB  Tile_X2Y8_LUT4AB
timestamp 0
transform 1 0 62250 0 1 377250
box 0 0 1 1
use LUT4AB  Tile_X2Y9_LUT4AB
timestamp 0
transform 1 0 62250 0 1 332250
box 0 0 1 1
use LUT4AB  Tile_X2Y10_LUT4AB
timestamp 0
transform 1 0 62250 0 1 287250
box 0 0 1 1
use LUT4AB  Tile_X2Y11_LUT4AB
timestamp 0
transform 1 0 62250 0 1 242250
box 0 0 1 1
use LUT4AB  Tile_X2Y12_LUT4AB
timestamp 0
transform 1 0 62250 0 1 197250
box 0 0 1 1
use LUT4AB  Tile_X2Y13_LUT4AB
timestamp 0
transform 1 0 62250 0 1 152250
box 0 0 1 1
use LUT4AB  Tile_X2Y14_LUT4AB
timestamp 0
transform 1 0 62250 0 1 107250
box 0 0 1 1
use LUT4AB  Tile_X2Y15_LUT4AB
timestamp 0
transform 1 0 62250 0 1 62250
box 0 0 1 1
use LUT4AB  Tile_X2Y16_LUT4AB
timestamp 0
transform 1 0 62250 0 1 17250
box 0 0 1 1
use S_WARMBOOT  Tile_X2Y17_S_WARMBOOT
timestamp 0
transform 1 0 62250 0 1 6000
box 0 0 1 1
use N_term_single2  Tile_X3Y0_N_term_single2
timestamp 0
transform 1 0 103250 0 1 737250
box 0 0 1 1
use RegFile  Tile_X3Y1_RegFile
timestamp 0
transform 1 0 103250 0 1 692250
box 0 0 1 1
use RegFile  Tile_X3Y2_RegFile
timestamp 0
transform 1 0 103250 0 1 647250
box 0 0 1 1
use RegFile  Tile_X3Y3_RegFile
timestamp 0
transform 1 0 103250 0 1 602250
box 0 0 1 1
use RegFile  Tile_X3Y4_RegFile
timestamp 0
transform 1 0 103250 0 1 557250
box 0 0 1 1
use RegFile  Tile_X3Y5_RegFile
timestamp 0
transform 1 0 103250 0 1 512250
box 0 0 1 1
use RegFile  Tile_X3Y6_RegFile
timestamp 0
transform 1 0 103250 0 1 467250
box 0 0 1 1
use RegFile  Tile_X3Y7_RegFile
timestamp 0
transform 1 0 103250 0 1 422250
box 0 0 1 1
use RegFile  Tile_X3Y8_RegFile
timestamp 0
transform 1 0 103250 0 1 377250
box 0 0 1 1
use RegFile  Tile_X3Y9_RegFile
timestamp 0
transform 1 0 103250 0 1 332250
box 0 0 1 1
use RegFile  Tile_X3Y10_RegFile
timestamp 0
transform 1 0 103250 0 1 287250
box 0 0 1 1
use RegFile  Tile_X3Y11_RegFile
timestamp 0
transform 1 0 103250 0 1 242250
box 0 0 1 1
use RegFile  Tile_X3Y12_RegFile
timestamp 0
transform 1 0 103250 0 1 197250
box 0 0 1 1
use RegFile  Tile_X3Y13_RegFile
timestamp 0
transform 1 0 103250 0 1 152250
box 0 0 1 1
use RegFile  Tile_X3Y14_RegFile
timestamp 0
transform 1 0 103250 0 1 107250
box 0 0 1 1
use RegFile  Tile_X3Y15_RegFile
timestamp 0
transform 1 0 103250 0 1 62250
box 0 0 1 1
use RegFile  Tile_X3Y16_RegFile
timestamp 0
transform 1 0 103250 0 1 17250
box 0 0 1 1
use S_term_single2  Tile_X3Y17_S_term_single2
timestamp 0
transform 1 0 103250 0 1 6000
box 0 0 1 1
use N_IO  Tile_X4Y0_N_IO
timestamp 0
transform 1 0 152250 0 1 737250
box 0 0 1 1
use LUT4AB  Tile_X4Y1_LUT4AB
timestamp 0
transform 1 0 152250 0 1 692250
box 0 0 1 1
use LUT4AB  Tile_X4Y2_LUT4AB
timestamp 0
transform 1 0 152250 0 1 647250
box 0 0 1 1
use LUT4AB  Tile_X4Y3_LUT4AB
timestamp 0
transform 1 0 152250 0 1 602250
box 0 0 1 1
use LUT4AB  Tile_X4Y4_LUT4AB
timestamp 0
transform 1 0 152250 0 1 557250
box 0 0 1 1
use LUT4AB  Tile_X4Y5_LUT4AB
timestamp 0
transform 1 0 152250 0 1 512250
box 0 0 1 1
use LUT4AB  Tile_X4Y6_LUT4AB
timestamp 0
transform 1 0 152250 0 1 467250
box 0 0 1 1
use LUT4AB  Tile_X4Y7_LUT4AB
timestamp 0
transform 1 0 152250 0 1 422250
box 0 0 1 1
use LUT4AB  Tile_X4Y8_LUT4AB
timestamp 0
transform 1 0 152250 0 1 377250
box 0 0 1 1
use LUT4AB  Tile_X4Y9_LUT4AB
timestamp 0
transform 1 0 152250 0 1 332250
box 0 0 1 1
use LUT4AB  Tile_X4Y10_LUT4AB
timestamp 0
transform 1 0 152250 0 1 287250
box 0 0 1 1
use LUT4AB  Tile_X4Y11_LUT4AB
timestamp 0
transform 1 0 152250 0 1 242250
box 0 0 1 1
use LUT4AB  Tile_X4Y12_LUT4AB
timestamp 0
transform 1 0 152250 0 1 197250
box 0 0 1 1
use LUT4AB  Tile_X4Y13_LUT4AB
timestamp 0
transform 1 0 152250 0 1 152250
box 0 0 1 1
use LUT4AB  Tile_X4Y14_LUT4AB
timestamp 0
transform 1 0 152250 0 1 107250
box 0 0 1 1
use LUT4AB  Tile_X4Y15_LUT4AB
timestamp 0
transform 1 0 152250 0 1 62250
box 0 0 1 1
use LUT4AB  Tile_X4Y16_LUT4AB
timestamp 0
transform 1 0 152250 0 1 17250
box 0 0 1 1
use S_CPU_IF  Tile_X4Y17_S_CPU_IF
timestamp 0
transform 1 0 152250 0 1 6000
box 0 0 1 1
use N_IO  Tile_X5Y0_N_IO
timestamp 0
transform 1 0 193250 0 1 737250
box 0 0 1 1
use LUT4AB  Tile_X5Y1_LUT4AB
timestamp 0
transform 1 0 193250 0 1 692250
box 0 0 1 1
use LUT4AB  Tile_X5Y2_LUT4AB
timestamp 0
transform 1 0 193250 0 1 647250
box 0 0 1 1
use LUT4AB  Tile_X5Y3_LUT4AB
timestamp 0
transform 1 0 193250 0 1 602250
box 0 0 1 1
use LUT4AB  Tile_X5Y4_LUT4AB
timestamp 0
transform 1 0 193250 0 1 557250
box 0 0 1 1
use LUT4AB  Tile_X5Y5_LUT4AB
timestamp 0
transform 1 0 193250 0 1 512250
box 0 0 1 1
use LUT4AB  Tile_X5Y6_LUT4AB
timestamp 0
transform 1 0 193250 0 1 467250
box 0 0 1 1
use LUT4AB  Tile_X5Y7_LUT4AB
timestamp 0
transform 1 0 193250 0 1 422250
box 0 0 1 1
use LUT4AB  Tile_X5Y8_LUT4AB
timestamp 0
transform 1 0 193250 0 1 377250
box 0 0 1 1
use LUT4AB  Tile_X5Y9_LUT4AB
timestamp 0
transform 1 0 193250 0 1 332250
box 0 0 1 1
use LUT4AB  Tile_X5Y10_LUT4AB
timestamp 0
transform 1 0 193250 0 1 287250
box 0 0 1 1
use LUT4AB  Tile_X5Y11_LUT4AB
timestamp 0
transform 1 0 193250 0 1 242250
box 0 0 1 1
use LUT4AB  Tile_X5Y12_LUT4AB
timestamp 0
transform 1 0 193250 0 1 197250
box 0 0 1 1
use LUT4AB  Tile_X5Y13_LUT4AB
timestamp 0
transform 1 0 193250 0 1 152250
box 0 0 1 1
use LUT4AB  Tile_X5Y14_LUT4AB
timestamp 0
transform 1 0 193250 0 1 107250
box 0 0 1 1
use LUT4AB  Tile_X5Y15_LUT4AB
timestamp 0
transform 1 0 193250 0 1 62250
box 0 0 1 1
use LUT4AB  Tile_X5Y16_LUT4AB
timestamp 0
transform 1 0 193250 0 1 17250
box 0 0 1 1
use S_CPU_IF  Tile_X5Y17_S_CPU_IF
timestamp 0
transform 1 0 193250 0 1 6000
box 0 0 1 1
use N_IO  Tile_X6Y0_N_IO
timestamp 0
transform 1 0 234250 0 1 737250
box 0 0 1 1
use LUT4AB  Tile_X6Y1_LUT4AB
timestamp 0
transform 1 0 234250 0 1 692250
box 0 0 1 1
use LUT4AB  Tile_X6Y2_LUT4AB
timestamp 0
transform 1 0 234250 0 1 647250
box 0 0 1 1
use LUT4AB  Tile_X6Y3_LUT4AB
timestamp 0
transform 1 0 234250 0 1 602250
box 0 0 1 1
use LUT4AB  Tile_X6Y4_LUT4AB
timestamp 0
transform 1 0 234250 0 1 557250
box 0 0 1 1
use LUT4AB  Tile_X6Y5_LUT4AB
timestamp 0
transform 1 0 234250 0 1 512250
box 0 0 1 1
use LUT4AB  Tile_X6Y6_LUT4AB
timestamp 0
transform 1 0 234250 0 1 467250
box 0 0 1 1
use LUT4AB  Tile_X6Y7_LUT4AB
timestamp 0
transform 1 0 234250 0 1 422250
box 0 0 1 1
use LUT4AB  Tile_X6Y8_LUT4AB
timestamp 0
transform 1 0 234250 0 1 377250
box 0 0 1 1
use LUT4AB  Tile_X6Y9_LUT4AB
timestamp 0
transform 1 0 234250 0 1 332250
box 0 0 1 1
use LUT4AB  Tile_X6Y10_LUT4AB
timestamp 0
transform 1 0 234250 0 1 287250
box 0 0 1 1
use LUT4AB  Tile_X6Y11_LUT4AB
timestamp 0
transform 1 0 234250 0 1 242250
box 0 0 1 1
use LUT4AB  Tile_X6Y12_LUT4AB
timestamp 0
transform 1 0 234250 0 1 197250
box 0 0 1 1
use LUT4AB  Tile_X6Y13_LUT4AB
timestamp 0
transform 1 0 234250 0 1 152250
box 0 0 1 1
use LUT4AB  Tile_X6Y14_LUT4AB
timestamp 0
transform 1 0 234250 0 1 107250
box 0 0 1 1
use LUT4AB  Tile_X6Y15_LUT4AB
timestamp 0
transform 1 0 234250 0 1 62250
box 0 0 1 1
use LUT4AB  Tile_X6Y16_LUT4AB
timestamp 0
transform 1 0 234250 0 1 17250
box 0 0 1 1
use S_CPU_IF  Tile_X6Y17_S_CPU_IF
timestamp 0
transform 1 0 234250 0 1 6000
box 0 0 1 1
use N_term_DSP  Tile_X7Y0_N_term_DSP
timestamp 0
transform 1 0 275250 0 1 737250
box 0 0 1 1
use DSP  Tile_X7Y1_DSP
timestamp 0
transform 1 0 275250 0 1 647250
box 0 0 1 1
use DSP  Tile_X7Y3_DSP
timestamp 0
transform 1 0 275250 0 1 557250
box 0 0 1 1
use DSP  Tile_X7Y5_DSP
timestamp 0
transform 1 0 275250 0 1 467250
box 0 0 1 1
use DSP  Tile_X7Y7_DSP
timestamp 0
transform 1 0 275250 0 1 377250
box 0 0 1 1
use DSP  Tile_X7Y9_DSP
timestamp 0
transform 1 0 275250 0 1 287250
box 0 0 1 1
use DSP  Tile_X7Y11_DSP
timestamp 0
transform 1 0 275250 0 1 197250
box 0 0 1 1
use DSP  Tile_X7Y13_DSP
timestamp 0
transform 1 0 275250 0 1 107250
box 0 0 1 1
use DSP  Tile_X7Y15_DSP
timestamp 0
transform 1 0 275250 0 1 17250
box 0 0 1 1
use S_term_DSP  Tile_X7Y17_S_term_DSP
timestamp 0
transform 1 0 275250 0 1 6000
box 0 0 1 1
use N_IO  Tile_X8Y0_N_IO
timestamp 0
transform 1 0 320250 0 1 737250
box 0 0 1 1
use LUT4AB  Tile_X8Y1_LUT4AB
timestamp 0
transform 1 0 320250 0 1 692250
box 0 0 1 1
use LUT4AB  Tile_X8Y2_LUT4AB
timestamp 0
transform 1 0 320250 0 1 647250
box 0 0 1 1
use LUT4AB  Tile_X8Y3_LUT4AB
timestamp 0
transform 1 0 320250 0 1 602250
box 0 0 1 1
use LUT4AB  Tile_X8Y4_LUT4AB
timestamp 0
transform 1 0 320250 0 1 557250
box 0 0 1 1
use LUT4AB  Tile_X8Y5_LUT4AB
timestamp 0
transform 1 0 320250 0 1 512250
box 0 0 1 1
use LUT4AB  Tile_X8Y6_LUT4AB
timestamp 0
transform 1 0 320250 0 1 467250
box 0 0 1 1
use LUT4AB  Tile_X8Y7_LUT4AB
timestamp 0
transform 1 0 320250 0 1 422250
box 0 0 1 1
use LUT4AB  Tile_X8Y8_LUT4AB
timestamp 0
transform 1 0 320250 0 1 377250
box 0 0 1 1
use LUT4AB  Tile_X8Y9_LUT4AB
timestamp 0
transform 1 0 320250 0 1 332250
box 0 0 1 1
use LUT4AB  Tile_X8Y10_LUT4AB
timestamp 0
transform 1 0 320250 0 1 287250
box 0 0 1 1
use LUT4AB  Tile_X8Y11_LUT4AB
timestamp 0
transform 1 0 320250 0 1 242250
box 0 0 1 1
use LUT4AB  Tile_X8Y12_LUT4AB
timestamp 0
transform 1 0 320250 0 1 197250
box 0 0 1 1
use LUT4AB  Tile_X8Y13_LUT4AB
timestamp 0
transform 1 0 320250 0 1 152250
box 0 0 1 1
use LUT4AB  Tile_X8Y14_LUT4AB
timestamp 0
transform 1 0 320250 0 1 107250
box 0 0 1 1
use LUT4AB  Tile_X8Y15_LUT4AB
timestamp 0
transform 1 0 320250 0 1 62250
box 0 0 1 1
use LUT4AB  Tile_X8Y16_LUT4AB
timestamp 0
transform 1 0 320250 0 1 17250
box 0 0 1 1
use S_CPU_IF  Tile_X8Y17_S_CPU_IF
timestamp 0
transform 1 0 320250 0 1 6000
box 0 0 1 1
use N_IO  Tile_X9Y0_N_IO
timestamp 0
transform 1 0 361250 0 1 737250
box 0 0 1 1
use LUT4AB  Tile_X9Y1_LUT4AB
timestamp 0
transform 1 0 361250 0 1 692250
box 0 0 1 1
use LUT4AB  Tile_X9Y2_LUT4AB
timestamp 0
transform 1 0 361250 0 1 647250
box 0 0 1 1
use LUT4AB  Tile_X9Y3_LUT4AB
timestamp 0
transform 1 0 361250 0 1 602250
box 0 0 1 1
use LUT4AB  Tile_X9Y4_LUT4AB
timestamp 0
transform 1 0 361250 0 1 557250
box 0 0 1 1
use LUT4AB  Tile_X9Y5_LUT4AB
timestamp 0
transform 1 0 361250 0 1 512250
box 0 0 1 1
use LUT4AB  Tile_X9Y6_LUT4AB
timestamp 0
transform 1 0 361250 0 1 467250
box 0 0 1 1
use LUT4AB  Tile_X9Y7_LUT4AB
timestamp 0
transform 1 0 361250 0 1 422250
box 0 0 1 1
use LUT4AB  Tile_X9Y8_LUT4AB
timestamp 0
transform 1 0 361250 0 1 377250
box 0 0 1 1
use LUT4AB  Tile_X9Y9_LUT4AB
timestamp 0
transform 1 0 361250 0 1 332250
box 0 0 1 1
use LUT4AB  Tile_X9Y10_LUT4AB
timestamp 0
transform 1 0 361250 0 1 287250
box 0 0 1 1
use LUT4AB  Tile_X9Y11_LUT4AB
timestamp 0
transform 1 0 361250 0 1 242250
box 0 0 1 1
use LUT4AB  Tile_X9Y12_LUT4AB
timestamp 0
transform 1 0 361250 0 1 197250
box 0 0 1 1
use LUT4AB  Tile_X9Y13_LUT4AB
timestamp 0
transform 1 0 361250 0 1 152250
box 0 0 1 1
use LUT4AB  Tile_X9Y14_LUT4AB
timestamp 0
transform 1 0 361250 0 1 107250
box 0 0 1 1
use LUT4AB  Tile_X9Y15_LUT4AB
timestamp 0
transform 1 0 361250 0 1 62250
box 0 0 1 1
use LUT4AB  Tile_X9Y16_LUT4AB
timestamp 0
transform 1 0 361250 0 1 17250
box 0 0 1 1
use S_EF_ADC12  Tile_X9Y17_S_EF_ADC12
timestamp 0
transform 1 0 361250 0 1 6000
box 0 0 1 1
use N_IO  Tile_X10Y0_N_IO
timestamp 0
transform 1 0 402250 0 1 737250
box 0 0 1 1
use LUT4AB  Tile_X10Y1_LUT4AB
timestamp 0
transform 1 0 402250 0 1 692250
box 0 0 1 1
use LUT4AB  Tile_X10Y2_LUT4AB
timestamp 0
transform 1 0 402250 0 1 647250
box 0 0 1 1
use LUT4AB  Tile_X10Y3_LUT4AB
timestamp 0
transform 1 0 402250 0 1 602250
box 0 0 1 1
use LUT4AB  Tile_X10Y4_LUT4AB
timestamp 0
transform 1 0 402250 0 1 557250
box 0 0 1 1
use LUT4AB  Tile_X10Y5_LUT4AB
timestamp 0
transform 1 0 402250 0 1 512250
box 0 0 1 1
use LUT4AB  Tile_X10Y6_LUT4AB
timestamp 0
transform 1 0 402250 0 1 467250
box 0 0 1 1
use LUT4AB  Tile_X10Y7_LUT4AB
timestamp 0
transform 1 0 402250 0 1 422250
box 0 0 1 1
use LUT4AB  Tile_X10Y8_LUT4AB
timestamp 0
transform 1 0 402250 0 1 377250
box 0 0 1 1
use LUT4AB  Tile_X10Y9_LUT4AB
timestamp 0
transform 1 0 402250 0 1 332250
box 0 0 1 1
use LUT4AB  Tile_X10Y10_LUT4AB
timestamp 0
transform 1 0 402250 0 1 287250
box 0 0 1 1
use LUT4AB  Tile_X10Y11_LUT4AB
timestamp 0
transform 1 0 402250 0 1 242250
box 0 0 1 1
use LUT4AB  Tile_X10Y12_LUT4AB
timestamp 0
transform 1 0 402250 0 1 197250
box 0 0 1 1
use LUT4AB  Tile_X10Y13_LUT4AB
timestamp 0
transform 1 0 402250 0 1 152250
box 0 0 1 1
use LUT4AB  Tile_X10Y14_LUT4AB
timestamp 0
transform 1 0 402250 0 1 107250
box 0 0 1 1
use LUT4AB  Tile_X10Y15_LUT4AB
timestamp 0
transform 1 0 402250 0 1 62250
box 0 0 1 1
use LUT4AB  Tile_X10Y16_LUT4AB
timestamp 0
transform 1 0 402250 0 1 17250
box 0 0 1 1
use S_EF_DAC8  Tile_X10Y17_S_EF_DAC8
timestamp 0
transform 1 0 402250 0 1 6000
box 0 0 1 1
use N_term_EF_SRAM  Tile_X11Y0_N_term_EF_SRAM
timestamp 0
transform 1 0 443250 0 1 737250
box 0 0 1 1
use EF_SRAM  Tile_X11Y1_EF_SRAM
timestamp 0
transform 1 0 443250 0 1 647250
box 0 0 1 1
use EF_SRAM  Tile_X11Y3_EF_SRAM
timestamp 0
transform 1 0 443250 0 1 557250
box 0 0 1 1
use EF_SRAM  Tile_X11Y5_EF_SRAM
timestamp 0
transform 1 0 443250 0 1 467250
box 0 0 1 1
use EF_SRAM  Tile_X11Y7_EF_SRAM
timestamp 0
transform 1 0 443250 0 1 377250
box 0 0 1 1
use EF_SRAM  Tile_X11Y9_EF_SRAM
timestamp 0
transform 1 0 443250 0 1 287250
box 0 0 1 1
use EF_SRAM  Tile_X11Y11_EF_SRAM
timestamp 0
transform 1 0 443250 0 1 197250
box 0 0 1 1
use EF_SRAM  Tile_X11Y13_EF_SRAM
timestamp 0
transform 1 0 443250 0 1 107250
box 0 0 1 1
use EF_SRAM  Tile_X11Y15_EF_SRAM
timestamp 0
transform 1 0 443250 0 1 17250
box 0 0 1 1
use S_term_EF_SRAM  Tile_X11Y17_S_term_EF_SRAM
timestamp 0
transform 1 0 443250 0 1 6000
box 0 0 1 1
<< labels >>
flabel metal2 s 7746 755700 7802 756500 0 FreeSans 224 90 0 0 FrameData[0]
port 0 nsew signal input
flabel metal3 s 0 620848 800 620968 0 FreeSans 480 0 0 0 FrameData[100]
port 1 nsew signal input
flabel metal3 s 0 621528 800 621648 0 FreeSans 480 0 0 0 FrameData[101]
port 2 nsew signal input
flabel metal3 s 0 622888 800 623008 0 FreeSans 480 0 0 0 FrameData[102]
port 3 nsew signal input
flabel metal3 s 0 623568 800 623688 0 FreeSans 480 0 0 0 FrameData[103]
port 4 nsew signal input
flabel metal3 s 0 624248 800 624368 0 FreeSans 480 0 0 0 FrameData[104]
port 5 nsew signal input
flabel metal3 s 0 624928 800 625048 0 FreeSans 480 0 0 0 FrameData[105]
port 6 nsew signal input
flabel metal3 s 0 625608 800 625728 0 FreeSans 480 0 0 0 FrameData[106]
port 7 nsew signal input
flabel metal3 s 0 626968 800 627088 0 FreeSans 480 0 0 0 FrameData[107]
port 8 nsew signal input
flabel metal3 s 0 627648 800 627768 0 FreeSans 480 0 0 0 FrameData[108]
port 9 nsew signal input
flabel metal3 s 0 628328 800 628448 0 FreeSans 480 0 0 0 FrameData[109]
port 10 nsew signal input
flabel metal2 s 21270 755700 21326 756500 0 FreeSans 224 90 0 0 FrameData[10]
port 11 nsew signal input
flabel metal3 s 0 629008 800 629128 0 FreeSans 480 0 0 0 FrameData[110]
port 12 nsew signal input
flabel metal3 s 0 629688 800 629808 0 FreeSans 480 0 0 0 FrameData[111]
port 13 nsew signal input
flabel metal3 s 0 631048 800 631168 0 FreeSans 480 0 0 0 FrameData[112]
port 14 nsew signal input
flabel metal3 s 0 631728 800 631848 0 FreeSans 480 0 0 0 FrameData[113]
port 15 nsew signal input
flabel metal3 s 0 632408 800 632528 0 FreeSans 480 0 0 0 FrameData[114]
port 16 nsew signal input
flabel metal3 s 0 633088 800 633208 0 FreeSans 480 0 0 0 FrameData[115]
port 17 nsew signal input
flabel metal3 s 0 633768 800 633888 0 FreeSans 480 0 0 0 FrameData[116]
port 18 nsew signal input
flabel metal3 s 0 635128 800 635248 0 FreeSans 480 0 0 0 FrameData[117]
port 19 nsew signal input
flabel metal3 s 0 635808 800 635928 0 FreeSans 480 0 0 0 FrameData[118]
port 20 nsew signal input
flabel metal3 s 0 636488 800 636608 0 FreeSans 480 0 0 0 FrameData[119]
port 21 nsew signal input
flabel metal2 s 15474 755700 15530 756500 0 FreeSans 224 90 0 0 FrameData[11]
port 22 nsew signal input
flabel metal3 s 0 637168 800 637288 0 FreeSans 480 0 0 0 FrameData[120]
port 23 nsew signal input
flabel metal3 s 0 637848 800 637968 0 FreeSans 480 0 0 0 FrameData[121]
port 24 nsew signal input
flabel metal3 s 0 639208 800 639328 0 FreeSans 480 0 0 0 FrameData[122]
port 25 nsew signal input
flabel metal3 s 0 639888 800 640008 0 FreeSans 480 0 0 0 FrameData[123]
port 26 nsew signal input
flabel metal3 s 0 640568 800 640688 0 FreeSans 480 0 0 0 FrameData[124]
port 27 nsew signal input
flabel metal3 s 0 641248 800 641368 0 FreeSans 480 0 0 0 FrameData[125]
port 28 nsew signal input
flabel metal3 s 0 641928 800 642048 0 FreeSans 480 0 0 0 FrameData[126]
port 29 nsew signal input
flabel metal3 s 0 643288 800 643408 0 FreeSans 480 0 0 0 FrameData[127]
port 30 nsew signal input
flabel metal3 s 0 572568 800 572688 0 FreeSans 480 0 0 0 FrameData[128]
port 31 nsew signal input
flabel metal3 s 0 573248 800 573368 0 FreeSans 480 0 0 0 FrameData[129]
port 32 nsew signal input
flabel metal2 s 12254 755700 12310 756500 0 FreeSans 224 90 0 0 FrameData[12]
port 33 nsew signal input
flabel metal3 s 0 574608 800 574728 0 FreeSans 480 0 0 0 FrameData[130]
port 34 nsew signal input
flabel metal3 s 0 575288 800 575408 0 FreeSans 480 0 0 0 FrameData[131]
port 35 nsew signal input
flabel metal3 s 0 575968 800 576088 0 FreeSans 480 0 0 0 FrameData[132]
port 36 nsew signal input
flabel metal3 s 0 576648 800 576768 0 FreeSans 480 0 0 0 FrameData[133]
port 37 nsew signal input
flabel metal3 s 0 577328 800 577448 0 FreeSans 480 0 0 0 FrameData[134]
port 38 nsew signal input
flabel metal3 s 0 578688 800 578808 0 FreeSans 480 0 0 0 FrameData[135]
port 39 nsew signal input
flabel metal3 s 0 579368 800 579488 0 FreeSans 480 0 0 0 FrameData[136]
port 40 nsew signal input
flabel metal3 s 0 580048 800 580168 0 FreeSans 480 0 0 0 FrameData[137]
port 41 nsew signal input
flabel metal3 s 0 580728 800 580848 0 FreeSans 480 0 0 0 FrameData[138]
port 42 nsew signal input
flabel metal3 s 0 581408 800 581528 0 FreeSans 480 0 0 0 FrameData[139]
port 43 nsew signal input
flabel metal2 s 19982 755700 20038 756500 0 FreeSans 224 90 0 0 FrameData[13]
port 44 nsew signal input
flabel metal3 s 0 582768 800 582888 0 FreeSans 480 0 0 0 FrameData[140]
port 45 nsew signal input
flabel metal3 s 0 583448 800 583568 0 FreeSans 480 0 0 0 FrameData[141]
port 46 nsew signal input
flabel metal3 s 0 584128 800 584248 0 FreeSans 480 0 0 0 FrameData[142]
port 47 nsew signal input
flabel metal3 s 0 584808 800 584928 0 FreeSans 480 0 0 0 FrameData[143]
port 48 nsew signal input
flabel metal3 s 0 585488 800 585608 0 FreeSans 480 0 0 0 FrameData[144]
port 49 nsew signal input
flabel metal3 s 0 586848 800 586968 0 FreeSans 480 0 0 0 FrameData[145]
port 50 nsew signal input
flabel metal3 s 0 587528 800 587648 0 FreeSans 480 0 0 0 FrameData[146]
port 51 nsew signal input
flabel metal3 s 0 588208 800 588328 0 FreeSans 480 0 0 0 FrameData[147]
port 52 nsew signal input
flabel metal3 s 0 588888 800 589008 0 FreeSans 480 0 0 0 FrameData[148]
port 53 nsew signal input
flabel metal3 s 0 589568 800 589688 0 FreeSans 480 0 0 0 FrameData[149]
port 54 nsew signal input
flabel metal2 s 20626 755700 20682 756500 0 FreeSans 224 90 0 0 FrameData[14]
port 55 nsew signal input
flabel metal3 s 0 590928 800 591048 0 FreeSans 480 0 0 0 FrameData[150]
port 56 nsew signal input
flabel metal3 s 0 591608 800 591728 0 FreeSans 480 0 0 0 FrameData[151]
port 57 nsew signal input
flabel metal3 s 0 592288 800 592408 0 FreeSans 480 0 0 0 FrameData[152]
port 58 nsew signal input
flabel metal3 s 0 592968 800 593088 0 FreeSans 480 0 0 0 FrameData[153]
port 59 nsew signal input
flabel metal3 s 0 593648 800 593768 0 FreeSans 480 0 0 0 FrameData[154]
port 60 nsew signal input
flabel metal3 s 0 595008 800 595128 0 FreeSans 480 0 0 0 FrameData[155]
port 61 nsew signal input
flabel metal3 s 0 595688 800 595808 0 FreeSans 480 0 0 0 FrameData[156]
port 62 nsew signal input
flabel metal3 s 0 596368 800 596488 0 FreeSans 480 0 0 0 FrameData[157]
port 63 nsew signal input
flabel metal3 s 0 597048 800 597168 0 FreeSans 480 0 0 0 FrameData[158]
port 64 nsew signal input
flabel metal3 s 0 597728 800 597848 0 FreeSans 480 0 0 0 FrameData[159]
port 65 nsew signal input
flabel metal2 s 14830 755700 14886 756500 0 FreeSans 224 90 0 0 FrameData[15]
port 66 nsew signal input
flabel metal3 s 0 527688 800 527808 0 FreeSans 480 0 0 0 FrameData[160]
port 67 nsew signal input
flabel metal3 s 0 528368 800 528488 0 FreeSans 480 0 0 0 FrameData[161]
port 68 nsew signal input
flabel metal3 s 0 529728 800 529848 0 FreeSans 480 0 0 0 FrameData[162]
port 69 nsew signal input
flabel metal3 s 0 530408 800 530528 0 FreeSans 480 0 0 0 FrameData[163]
port 70 nsew signal input
flabel metal3 s 0 531088 800 531208 0 FreeSans 480 0 0 0 FrameData[164]
port 71 nsew signal input
flabel metal3 s 0 531768 800 531888 0 FreeSans 480 0 0 0 FrameData[165]
port 72 nsew signal input
flabel metal3 s 0 532448 800 532568 0 FreeSans 480 0 0 0 FrameData[166]
port 73 nsew signal input
flabel metal3 s 0 533808 800 533928 0 FreeSans 480 0 0 0 FrameData[167]
port 74 nsew signal input
flabel metal3 s 0 534488 800 534608 0 FreeSans 480 0 0 0 FrameData[168]
port 75 nsew signal input
flabel metal3 s 0 535168 800 535288 0 FreeSans 480 0 0 0 FrameData[169]
port 76 nsew signal input
flabel metal2 s 10322 755700 10378 756500 0 FreeSans 224 90 0 0 FrameData[16]
port 77 nsew signal input
flabel metal3 s 0 535848 800 535968 0 FreeSans 480 0 0 0 FrameData[170]
port 78 nsew signal input
flabel metal3 s 0 536528 800 536648 0 FreeSans 480 0 0 0 FrameData[171]
port 79 nsew signal input
flabel metal3 s 0 537888 800 538008 0 FreeSans 480 0 0 0 FrameData[172]
port 80 nsew signal input
flabel metal3 s 0 538568 800 538688 0 FreeSans 480 0 0 0 FrameData[173]
port 81 nsew signal input
flabel metal3 s 0 539248 800 539368 0 FreeSans 480 0 0 0 FrameData[174]
port 82 nsew signal input
flabel metal3 s 0 539928 800 540048 0 FreeSans 480 0 0 0 FrameData[175]
port 83 nsew signal input
flabel metal3 s 0 540608 800 540728 0 FreeSans 480 0 0 0 FrameData[176]
port 84 nsew signal input
flabel metal3 s 0 541968 800 542088 0 FreeSans 480 0 0 0 FrameData[177]
port 85 nsew signal input
flabel metal3 s 0 542648 800 542768 0 FreeSans 480 0 0 0 FrameData[178]
port 86 nsew signal input
flabel metal3 s 0 543328 800 543448 0 FreeSans 480 0 0 0 FrameData[179]
port 87 nsew signal input
flabel metal2 s 28354 755700 28410 756500 0 FreeSans 224 90 0 0 FrameData[17]
port 88 nsew signal input
flabel metal3 s 0 544008 800 544128 0 FreeSans 480 0 0 0 FrameData[180]
port 89 nsew signal input
flabel metal3 s 0 544688 800 544808 0 FreeSans 480 0 0 0 FrameData[181]
port 90 nsew signal input
flabel metal3 s 0 546048 800 546168 0 FreeSans 480 0 0 0 FrameData[182]
port 91 nsew signal input
flabel metal3 s 0 546728 800 546848 0 FreeSans 480 0 0 0 FrameData[183]
port 92 nsew signal input
flabel metal3 s 0 547408 800 547528 0 FreeSans 480 0 0 0 FrameData[184]
port 93 nsew signal input
flabel metal3 s 0 548088 800 548208 0 FreeSans 480 0 0 0 FrameData[185]
port 94 nsew signal input
flabel metal3 s 0 548768 800 548888 0 FreeSans 480 0 0 0 FrameData[186]
port 95 nsew signal input
flabel metal3 s 0 550128 800 550248 0 FreeSans 480 0 0 0 FrameData[187]
port 96 nsew signal input
flabel metal3 s 0 550808 800 550928 0 FreeSans 480 0 0 0 FrameData[188]
port 97 nsew signal input
flabel metal3 s 0 551488 800 551608 0 FreeSans 480 0 0 0 FrameData[189]
port 98 nsew signal input
flabel metal2 s 17406 755700 17462 756500 0 FreeSans 224 90 0 0 FrameData[18]
port 99 nsew signal input
flabel metal3 s 0 552168 800 552288 0 FreeSans 480 0 0 0 FrameData[190]
port 100 nsew signal input
flabel metal3 s 0 552848 800 552968 0 FreeSans 480 0 0 0 FrameData[191]
port 101 nsew signal input
flabel metal3 s 0 482808 800 482928 0 FreeSans 480 0 0 0 FrameData[192]
port 102 nsew signal input
flabel metal3 s 0 483488 800 483608 0 FreeSans 480 0 0 0 FrameData[193]
port 103 nsew signal input
flabel metal3 s 0 484168 800 484288 0 FreeSans 480 0 0 0 FrameData[194]
port 104 nsew signal input
flabel metal3 s 0 485528 800 485648 0 FreeSans 480 0 0 0 FrameData[195]
port 105 nsew signal input
flabel metal3 s 0 486208 800 486328 0 FreeSans 480 0 0 0 FrameData[196]
port 106 nsew signal input
flabel metal3 s 0 486888 800 487008 0 FreeSans 480 0 0 0 FrameData[197]
port 107 nsew signal input
flabel metal3 s 0 487568 800 487688 0 FreeSans 480 0 0 0 FrameData[198]
port 108 nsew signal input
flabel metal3 s 0 488248 800 488368 0 FreeSans 480 0 0 0 FrameData[199]
port 109 nsew signal input
flabel metal2 s 11610 755700 11666 756500 0 FreeSans 224 90 0 0 FrameData[19]
port 110 nsew signal input
flabel metal2 s 14186 755700 14242 756500 0 FreeSans 224 90 0 0 FrameData[1]
port 111 nsew signal input
flabel metal3 s 0 489608 800 489728 0 FreeSans 480 0 0 0 FrameData[200]
port 112 nsew signal input
flabel metal3 s 0 490288 800 490408 0 FreeSans 480 0 0 0 FrameData[201]
port 113 nsew signal input
flabel metal3 s 0 490968 800 491088 0 FreeSans 480 0 0 0 FrameData[202]
port 114 nsew signal input
flabel metal3 s 0 491648 800 491768 0 FreeSans 480 0 0 0 FrameData[203]
port 115 nsew signal input
flabel metal3 s 0 492328 800 492448 0 FreeSans 480 0 0 0 FrameData[204]
port 116 nsew signal input
flabel metal3 s 0 493688 800 493808 0 FreeSans 480 0 0 0 FrameData[205]
port 117 nsew signal input
flabel metal3 s 0 494368 800 494488 0 FreeSans 480 0 0 0 FrameData[206]
port 118 nsew signal input
flabel metal3 s 0 495048 800 495168 0 FreeSans 480 0 0 0 FrameData[207]
port 119 nsew signal input
flabel metal3 s 0 495728 800 495848 0 FreeSans 480 0 0 0 FrameData[208]
port 120 nsew signal input
flabel metal3 s 0 496408 800 496528 0 FreeSans 480 0 0 0 FrameData[209]
port 121 nsew signal input
flabel metal2 s 19338 755700 19394 756500 0 FreeSans 224 90 0 0 FrameData[20]
port 122 nsew signal input
flabel metal3 s 0 497768 800 497888 0 FreeSans 480 0 0 0 FrameData[210]
port 123 nsew signal input
flabel metal3 s 0 498448 800 498568 0 FreeSans 480 0 0 0 FrameData[211]
port 124 nsew signal input
flabel metal3 s 0 499128 800 499248 0 FreeSans 480 0 0 0 FrameData[212]
port 125 nsew signal input
flabel metal3 s 0 499808 800 499928 0 FreeSans 480 0 0 0 FrameData[213]
port 126 nsew signal input
flabel metal3 s 0 500488 800 500608 0 FreeSans 480 0 0 0 FrameData[214]
port 127 nsew signal input
flabel metal3 s 0 501848 800 501968 0 FreeSans 480 0 0 0 FrameData[215]
port 128 nsew signal input
flabel metal3 s 0 502528 800 502648 0 FreeSans 480 0 0 0 FrameData[216]
port 129 nsew signal input
flabel metal3 s 0 503208 800 503328 0 FreeSans 480 0 0 0 FrameData[217]
port 130 nsew signal input
flabel metal3 s 0 503888 800 504008 0 FreeSans 480 0 0 0 FrameData[218]
port 131 nsew signal input
flabel metal3 s 0 504568 800 504688 0 FreeSans 480 0 0 0 FrameData[219]
port 132 nsew signal input
flabel metal2 s 22558 755700 22614 756500 0 FreeSans 224 90 0 0 FrameData[21]
port 133 nsew signal input
flabel metal3 s 0 505928 800 506048 0 FreeSans 480 0 0 0 FrameData[220]
port 134 nsew signal input
flabel metal3 s 0 506608 800 506728 0 FreeSans 480 0 0 0 FrameData[221]
port 135 nsew signal input
flabel metal3 s 0 507288 800 507408 0 FreeSans 480 0 0 0 FrameData[222]
port 136 nsew signal input
flabel metal3 s 0 507968 800 508088 0 FreeSans 480 0 0 0 FrameData[223]
port 137 nsew signal input
flabel metal3 s 0 437928 800 438048 0 FreeSans 480 0 0 0 FrameData[224]
port 138 nsew signal input
flabel metal3 s 0 438608 800 438728 0 FreeSans 480 0 0 0 FrameData[225]
port 139 nsew signal input
flabel metal3 s 0 439288 800 439408 0 FreeSans 480 0 0 0 FrameData[226]
port 140 nsew signal input
flabel metal3 s 0 439968 800 440088 0 FreeSans 480 0 0 0 FrameData[227]
port 141 nsew signal input
flabel metal3 s 0 441328 800 441448 0 FreeSans 480 0 0 0 FrameData[228]
port 142 nsew signal input
flabel metal3 s 0 442008 800 442128 0 FreeSans 480 0 0 0 FrameData[229]
port 143 nsew signal input
flabel metal2 s 23846 755700 23902 756500 0 FreeSans 224 90 0 0 FrameData[22]
port 144 nsew signal input
flabel metal3 s 0 442688 800 442808 0 FreeSans 480 0 0 0 FrameData[230]
port 145 nsew signal input
flabel metal3 s 0 443368 800 443488 0 FreeSans 480 0 0 0 FrameData[231]
port 146 nsew signal input
flabel metal3 s 0 444048 800 444168 0 FreeSans 480 0 0 0 FrameData[232]
port 147 nsew signal input
flabel metal3 s 0 445408 800 445528 0 FreeSans 480 0 0 0 FrameData[233]
port 148 nsew signal input
flabel metal3 s 0 446088 800 446208 0 FreeSans 480 0 0 0 FrameData[234]
port 149 nsew signal input
flabel metal3 s 0 446768 800 446888 0 FreeSans 480 0 0 0 FrameData[235]
port 150 nsew signal input
flabel metal3 s 0 447448 800 447568 0 FreeSans 480 0 0 0 FrameData[236]
port 151 nsew signal input
flabel metal3 s 0 448128 800 448248 0 FreeSans 480 0 0 0 FrameData[237]
port 152 nsew signal input
flabel metal3 s 0 449488 800 449608 0 FreeSans 480 0 0 0 FrameData[238]
port 153 nsew signal input
flabel metal3 s 0 450168 800 450288 0 FreeSans 480 0 0 0 FrameData[239]
port 154 nsew signal input
flabel metal2 s 13542 755700 13598 756500 0 FreeSans 224 90 0 0 FrameData[23]
port 155 nsew signal input
flabel metal3 s 0 450848 800 450968 0 FreeSans 480 0 0 0 FrameData[240]
port 156 nsew signal input
flabel metal3 s 0 451528 800 451648 0 FreeSans 480 0 0 0 FrameData[241]
port 157 nsew signal input
flabel metal3 s 0 452208 800 452328 0 FreeSans 480 0 0 0 FrameData[242]
port 158 nsew signal input
flabel metal3 s 0 453568 800 453688 0 FreeSans 480 0 0 0 FrameData[243]
port 159 nsew signal input
flabel metal3 s 0 454248 800 454368 0 FreeSans 480 0 0 0 FrameData[244]
port 160 nsew signal input
flabel metal3 s 0 454928 800 455048 0 FreeSans 480 0 0 0 FrameData[245]
port 161 nsew signal input
flabel metal3 s 0 455608 800 455728 0 FreeSans 480 0 0 0 FrameData[246]
port 162 nsew signal input
flabel metal3 s 0 456288 800 456408 0 FreeSans 480 0 0 0 FrameData[247]
port 163 nsew signal input
flabel metal3 s 0 457648 800 457768 0 FreeSans 480 0 0 0 FrameData[248]
port 164 nsew signal input
flabel metal3 s 0 458328 800 458448 0 FreeSans 480 0 0 0 FrameData[249]
port 165 nsew signal input
flabel metal2 s 18694 755700 18750 756500 0 FreeSans 224 90 0 0 FrameData[24]
port 166 nsew signal input
flabel metal3 s 0 459008 800 459128 0 FreeSans 480 0 0 0 FrameData[250]
port 167 nsew signal input
flabel metal3 s 0 459688 800 459808 0 FreeSans 480 0 0 0 FrameData[251]
port 168 nsew signal input
flabel metal3 s 0 460368 800 460488 0 FreeSans 480 0 0 0 FrameData[252]
port 169 nsew signal input
flabel metal3 s 0 461728 800 461848 0 FreeSans 480 0 0 0 FrameData[253]
port 170 nsew signal input
flabel metal3 s 0 462408 800 462528 0 FreeSans 480 0 0 0 FrameData[254]
port 171 nsew signal input
flabel metal3 s 0 463088 800 463208 0 FreeSans 480 0 0 0 FrameData[255]
port 172 nsew signal input
flabel metal3 s 0 393048 800 393168 0 FreeSans 480 0 0 0 FrameData[256]
port 173 nsew signal input
flabel metal3 s 0 393728 800 393848 0 FreeSans 480 0 0 0 FrameData[257]
port 174 nsew signal input
flabel metal3 s 0 394408 800 394528 0 FreeSans 480 0 0 0 FrameData[258]
port 175 nsew signal input
flabel metal3 s 0 395088 800 395208 0 FreeSans 480 0 0 0 FrameData[259]
port 176 nsew signal input
flabel metal2 s 8390 755700 8446 756500 0 FreeSans 224 90 0 0 FrameData[25]
port 177 nsew signal input
flabel metal3 s 0 395768 800 395888 0 FreeSans 480 0 0 0 FrameData[260]
port 178 nsew signal input
flabel metal3 s 0 397128 800 397248 0 FreeSans 480 0 0 0 FrameData[261]
port 179 nsew signal input
flabel metal3 s 0 397808 800 397928 0 FreeSans 480 0 0 0 FrameData[262]
port 180 nsew signal input
flabel metal3 s 0 398488 800 398608 0 FreeSans 480 0 0 0 FrameData[263]
port 181 nsew signal input
flabel metal3 s 0 399168 800 399288 0 FreeSans 480 0 0 0 FrameData[264]
port 182 nsew signal input
flabel metal3 s 0 399848 800 399968 0 FreeSans 480 0 0 0 FrameData[265]
port 183 nsew signal input
flabel metal3 s 0 401208 800 401328 0 FreeSans 480 0 0 0 FrameData[266]
port 184 nsew signal input
flabel metal3 s 0 401888 800 402008 0 FreeSans 480 0 0 0 FrameData[267]
port 185 nsew signal input
flabel metal3 s 0 402568 800 402688 0 FreeSans 480 0 0 0 FrameData[268]
port 186 nsew signal input
flabel metal3 s 0 403248 800 403368 0 FreeSans 480 0 0 0 FrameData[269]
port 187 nsew signal input
flabel metal2 s 31574 755700 31630 756500 0 FreeSans 224 90 0 0 FrameData[26]
port 188 nsew signal input
flabel metal3 s 0 403928 800 404048 0 FreeSans 480 0 0 0 FrameData[270]
port 189 nsew signal input
flabel metal3 s 0 405288 800 405408 0 FreeSans 480 0 0 0 FrameData[271]
port 190 nsew signal input
flabel metal3 s 0 405968 800 406088 0 FreeSans 480 0 0 0 FrameData[272]
port 191 nsew signal input
flabel metal3 s 0 406648 800 406768 0 FreeSans 480 0 0 0 FrameData[273]
port 192 nsew signal input
flabel metal3 s 0 407328 800 407448 0 FreeSans 480 0 0 0 FrameData[274]
port 193 nsew signal input
flabel metal3 s 0 408008 800 408128 0 FreeSans 480 0 0 0 FrameData[275]
port 194 nsew signal input
flabel metal3 s 0 409368 800 409488 0 FreeSans 480 0 0 0 FrameData[276]
port 195 nsew signal input
flabel metal3 s 0 410048 800 410168 0 FreeSans 480 0 0 0 FrameData[277]
port 196 nsew signal input
flabel metal3 s 0 410728 800 410848 0 FreeSans 480 0 0 0 FrameData[278]
port 197 nsew signal input
flabel metal3 s 0 411408 800 411528 0 FreeSans 480 0 0 0 FrameData[279]
port 198 nsew signal input
flabel metal2 s 18050 755700 18106 756500 0 FreeSans 224 90 0 0 FrameData[27]
port 199 nsew signal input
flabel metal3 s 0 412088 800 412208 0 FreeSans 480 0 0 0 FrameData[280]
port 200 nsew signal input
flabel metal3 s 0 413448 800 413568 0 FreeSans 480 0 0 0 FrameData[281]
port 201 nsew signal input
flabel metal3 s 0 414128 800 414248 0 FreeSans 480 0 0 0 FrameData[282]
port 202 nsew signal input
flabel metal3 s 0 414808 800 414928 0 FreeSans 480 0 0 0 FrameData[283]
port 203 nsew signal input
flabel metal3 s 0 415488 800 415608 0 FreeSans 480 0 0 0 FrameData[284]
port 204 nsew signal input
flabel metal3 s 0 416168 800 416288 0 FreeSans 480 0 0 0 FrameData[285]
port 205 nsew signal input
flabel metal3 s 0 417528 800 417648 0 FreeSans 480 0 0 0 FrameData[286]
port 206 nsew signal input
flabel metal3 s 0 418208 800 418328 0 FreeSans 480 0 0 0 FrameData[287]
port 207 nsew signal input
flabel metal3 s 0 347488 800 347608 0 FreeSans 480 0 0 0 FrameData[288]
port 208 nsew signal input
flabel metal3 s 0 348168 800 348288 0 FreeSans 480 0 0 0 FrameData[289]
port 209 nsew signal input
flabel metal2 s 9678 755700 9734 756500 0 FreeSans 224 90 0 0 FrameData[28]
port 210 nsew signal input
flabel metal3 s 0 349528 800 349648 0 FreeSans 480 0 0 0 FrameData[290]
port 211 nsew signal input
flabel metal3 s 0 350208 800 350328 0 FreeSans 480 0 0 0 FrameData[291]
port 212 nsew signal input
flabel metal3 s 0 350888 800 351008 0 FreeSans 480 0 0 0 FrameData[292]
port 213 nsew signal input
flabel metal3 s 0 351568 800 351688 0 FreeSans 480 0 0 0 FrameData[293]
port 214 nsew signal input
flabel metal3 s 0 352928 800 353048 0 FreeSans 480 0 0 0 FrameData[294]
port 215 nsew signal input
flabel metal3 s 0 353608 800 353728 0 FreeSans 480 0 0 0 FrameData[295]
port 216 nsew signal input
flabel metal3 s 0 354288 800 354408 0 FreeSans 480 0 0 0 FrameData[296]
port 217 nsew signal input
flabel metal3 s 0 354968 800 355088 0 FreeSans 480 0 0 0 FrameData[297]
port 218 nsew signal input
flabel metal3 s 0 355648 800 355768 0 FreeSans 480 0 0 0 FrameData[298]
port 219 nsew signal input
flabel metal3 s 0 357008 800 357128 0 FreeSans 480 0 0 0 FrameData[299]
port 220 nsew signal input
flabel metal2 s 12898 755700 12954 756500 0 FreeSans 224 90 0 0 FrameData[29]
port 221 nsew signal input
flabel metal2 s 10966 755700 11022 756500 0 FreeSans 224 90 0 0 FrameData[2]
port 222 nsew signal input
flabel metal3 s 0 357688 800 357808 0 FreeSans 480 0 0 0 FrameData[300]
port 223 nsew signal input
flabel metal3 s 0 358368 800 358488 0 FreeSans 480 0 0 0 FrameData[301]
port 224 nsew signal input
flabel metal3 s 0 359048 800 359168 0 FreeSans 480 0 0 0 FrameData[302]
port 225 nsew signal input
flabel metal3 s 0 359728 800 359848 0 FreeSans 480 0 0 0 FrameData[303]
port 226 nsew signal input
flabel metal3 s 0 361088 800 361208 0 FreeSans 480 0 0 0 FrameData[304]
port 227 nsew signal input
flabel metal3 s 0 361768 800 361888 0 FreeSans 480 0 0 0 FrameData[305]
port 228 nsew signal input
flabel metal3 s 0 362448 800 362568 0 FreeSans 480 0 0 0 FrameData[306]
port 229 nsew signal input
flabel metal3 s 0 363128 800 363248 0 FreeSans 480 0 0 0 FrameData[307]
port 230 nsew signal input
flabel metal3 s 0 363808 800 363928 0 FreeSans 480 0 0 0 FrameData[308]
port 231 nsew signal input
flabel metal3 s 0 365168 800 365288 0 FreeSans 480 0 0 0 FrameData[309]
port 232 nsew signal input
flabel metal2 s 27066 755700 27122 756500 0 FreeSans 224 90 0 0 FrameData[30]
port 233 nsew signal input
flabel metal3 s 0 365848 800 365968 0 FreeSans 480 0 0 0 FrameData[310]
port 234 nsew signal input
flabel metal3 s 0 366528 800 366648 0 FreeSans 480 0 0 0 FrameData[311]
port 235 nsew signal input
flabel metal3 s 0 367208 800 367328 0 FreeSans 480 0 0 0 FrameData[312]
port 236 nsew signal input
flabel metal3 s 0 367888 800 368008 0 FreeSans 480 0 0 0 FrameData[313]
port 237 nsew signal input
flabel metal3 s 0 369248 800 369368 0 FreeSans 480 0 0 0 FrameData[314]
port 238 nsew signal input
flabel metal3 s 0 369928 800 370048 0 FreeSans 480 0 0 0 FrameData[315]
port 239 nsew signal input
flabel metal3 s 0 370608 800 370728 0 FreeSans 480 0 0 0 FrameData[316]
port 240 nsew signal input
flabel metal3 s 0 371288 800 371408 0 FreeSans 480 0 0 0 FrameData[317]
port 241 nsew signal input
flabel metal3 s 0 371968 800 372088 0 FreeSans 480 0 0 0 FrameData[318]
port 242 nsew signal input
flabel metal3 s 0 373328 800 373448 0 FreeSans 480 0 0 0 FrameData[319]
port 243 nsew signal input
flabel metal2 s 9034 755700 9090 756500 0 FreeSans 224 90 0 0 FrameData[31]
port 244 nsew signal input
flabel metal3 s 0 302608 800 302728 0 FreeSans 480 0 0 0 FrameData[320]
port 245 nsew signal input
flabel metal3 s 0 303288 800 303408 0 FreeSans 480 0 0 0 FrameData[321]
port 246 nsew signal input
flabel metal3 s 0 304648 800 304768 0 FreeSans 480 0 0 0 FrameData[322]
port 247 nsew signal input
flabel metal3 s 0 305328 800 305448 0 FreeSans 480 0 0 0 FrameData[323]
port 248 nsew signal input
flabel metal3 s 0 306008 800 306128 0 FreeSans 480 0 0 0 FrameData[324]
port 249 nsew signal input
flabel metal3 s 0 306688 800 306808 0 FreeSans 480 0 0 0 FrameData[325]
port 250 nsew signal input
flabel metal3 s 0 307368 800 307488 0 FreeSans 480 0 0 0 FrameData[326]
port 251 nsew signal input
flabel metal3 s 0 308728 800 308848 0 FreeSans 480 0 0 0 FrameData[327]
port 252 nsew signal input
flabel metal3 s 0 309408 800 309528 0 FreeSans 480 0 0 0 FrameData[328]
port 253 nsew signal input
flabel metal3 s 0 310088 800 310208 0 FreeSans 480 0 0 0 FrameData[329]
port 254 nsew signal input
flabel metal3 s 0 707888 800 708008 0 FreeSans 480 0 0 0 FrameData[32]
port 255 nsew signal input
flabel metal3 s 0 310768 800 310888 0 FreeSans 480 0 0 0 FrameData[330]
port 256 nsew signal input
flabel metal3 s 0 311448 800 311568 0 FreeSans 480 0 0 0 FrameData[331]
port 257 nsew signal input
flabel metal3 s 0 312808 800 312928 0 FreeSans 480 0 0 0 FrameData[332]
port 258 nsew signal input
flabel metal3 s 0 313488 800 313608 0 FreeSans 480 0 0 0 FrameData[333]
port 259 nsew signal input
flabel metal3 s 0 314168 800 314288 0 FreeSans 480 0 0 0 FrameData[334]
port 260 nsew signal input
flabel metal3 s 0 314848 800 314968 0 FreeSans 480 0 0 0 FrameData[335]
port 261 nsew signal input
flabel metal3 s 0 315528 800 315648 0 FreeSans 480 0 0 0 FrameData[336]
port 262 nsew signal input
flabel metal3 s 0 316888 800 317008 0 FreeSans 480 0 0 0 FrameData[337]
port 263 nsew signal input
flabel metal3 s 0 317568 800 317688 0 FreeSans 480 0 0 0 FrameData[338]
port 264 nsew signal input
flabel metal3 s 0 318248 800 318368 0 FreeSans 480 0 0 0 FrameData[339]
port 265 nsew signal input
flabel metal3 s 0 708568 800 708688 0 FreeSans 480 0 0 0 FrameData[33]
port 266 nsew signal input
flabel metal3 s 0 318928 800 319048 0 FreeSans 480 0 0 0 FrameData[340]
port 267 nsew signal input
flabel metal3 s 0 319608 800 319728 0 FreeSans 480 0 0 0 FrameData[341]
port 268 nsew signal input
flabel metal3 s 0 320968 800 321088 0 FreeSans 480 0 0 0 FrameData[342]
port 269 nsew signal input
flabel metal3 s 0 321648 800 321768 0 FreeSans 480 0 0 0 FrameData[343]
port 270 nsew signal input
flabel metal3 s 0 322328 800 322448 0 FreeSans 480 0 0 0 FrameData[344]
port 271 nsew signal input
flabel metal3 s 0 323008 800 323128 0 FreeSans 480 0 0 0 FrameData[345]
port 272 nsew signal input
flabel metal3 s 0 323688 800 323808 0 FreeSans 480 0 0 0 FrameData[346]
port 273 nsew signal input
flabel metal3 s 0 325048 800 325168 0 FreeSans 480 0 0 0 FrameData[347]
port 274 nsew signal input
flabel metal3 s 0 325728 800 325848 0 FreeSans 480 0 0 0 FrameData[348]
port 275 nsew signal input
flabel metal3 s 0 326408 800 326528 0 FreeSans 480 0 0 0 FrameData[349]
port 276 nsew signal input
flabel metal3 s 0 709248 800 709368 0 FreeSans 480 0 0 0 FrameData[34]
port 277 nsew signal input
flabel metal3 s 0 327088 800 327208 0 FreeSans 480 0 0 0 FrameData[350]
port 278 nsew signal input
flabel metal3 s 0 327768 800 327888 0 FreeSans 480 0 0 0 FrameData[351]
port 279 nsew signal input
flabel metal3 s 0 257728 800 257848 0 FreeSans 480 0 0 0 FrameData[352]
port 280 nsew signal input
flabel metal3 s 0 258408 800 258528 0 FreeSans 480 0 0 0 FrameData[353]
port 281 nsew signal input
flabel metal3 s 0 259088 800 259208 0 FreeSans 480 0 0 0 FrameData[354]
port 282 nsew signal input
flabel metal3 s 0 260448 800 260568 0 FreeSans 480 0 0 0 FrameData[355]
port 283 nsew signal input
flabel metal3 s 0 261128 800 261248 0 FreeSans 480 0 0 0 FrameData[356]
port 284 nsew signal input
flabel metal3 s 0 261808 800 261928 0 FreeSans 480 0 0 0 FrameData[357]
port 285 nsew signal input
flabel metal3 s 0 262488 800 262608 0 FreeSans 480 0 0 0 FrameData[358]
port 286 nsew signal input
flabel metal3 s 0 263168 800 263288 0 FreeSans 480 0 0 0 FrameData[359]
port 287 nsew signal input
flabel metal3 s 0 709928 800 710048 0 FreeSans 480 0 0 0 FrameData[35]
port 288 nsew signal input
flabel metal3 s 0 264528 800 264648 0 FreeSans 480 0 0 0 FrameData[360]
port 289 nsew signal input
flabel metal3 s 0 265208 800 265328 0 FreeSans 480 0 0 0 FrameData[361]
port 290 nsew signal input
flabel metal3 s 0 265888 800 266008 0 FreeSans 480 0 0 0 FrameData[362]
port 291 nsew signal input
flabel metal3 s 0 266568 800 266688 0 FreeSans 480 0 0 0 FrameData[363]
port 292 nsew signal input
flabel metal3 s 0 267248 800 267368 0 FreeSans 480 0 0 0 FrameData[364]
port 293 nsew signal input
flabel metal3 s 0 268608 800 268728 0 FreeSans 480 0 0 0 FrameData[365]
port 294 nsew signal input
flabel metal3 s 0 269288 800 269408 0 FreeSans 480 0 0 0 FrameData[366]
port 295 nsew signal input
flabel metal3 s 0 269968 800 270088 0 FreeSans 480 0 0 0 FrameData[367]
port 296 nsew signal input
flabel metal3 s 0 270648 800 270768 0 FreeSans 480 0 0 0 FrameData[368]
port 297 nsew signal input
flabel metal3 s 0 271328 800 271448 0 FreeSans 480 0 0 0 FrameData[369]
port 298 nsew signal input
flabel metal3 s 0 711288 800 711408 0 FreeSans 480 0 0 0 FrameData[36]
port 299 nsew signal input
flabel metal3 s 0 272688 800 272808 0 FreeSans 480 0 0 0 FrameData[370]
port 300 nsew signal input
flabel metal3 s 0 273368 800 273488 0 FreeSans 480 0 0 0 FrameData[371]
port 301 nsew signal input
flabel metal3 s 0 274048 800 274168 0 FreeSans 480 0 0 0 FrameData[372]
port 302 nsew signal input
flabel metal3 s 0 274728 800 274848 0 FreeSans 480 0 0 0 FrameData[373]
port 303 nsew signal input
flabel metal3 s 0 275408 800 275528 0 FreeSans 480 0 0 0 FrameData[374]
port 304 nsew signal input
flabel metal3 s 0 276768 800 276888 0 FreeSans 480 0 0 0 FrameData[375]
port 305 nsew signal input
flabel metal3 s 0 277448 800 277568 0 FreeSans 480 0 0 0 FrameData[376]
port 306 nsew signal input
flabel metal3 s 0 278128 800 278248 0 FreeSans 480 0 0 0 FrameData[377]
port 307 nsew signal input
flabel metal3 s 0 278808 800 278928 0 FreeSans 480 0 0 0 FrameData[378]
port 308 nsew signal input
flabel metal3 s 0 279488 800 279608 0 FreeSans 480 0 0 0 FrameData[379]
port 309 nsew signal input
flabel metal3 s 0 711968 800 712088 0 FreeSans 480 0 0 0 FrameData[37]
port 310 nsew signal input
flabel metal3 s 0 280848 800 280968 0 FreeSans 480 0 0 0 FrameData[380]
port 311 nsew signal input
flabel metal3 s 0 281528 800 281648 0 FreeSans 480 0 0 0 FrameData[381]
port 312 nsew signal input
flabel metal3 s 0 282208 800 282328 0 FreeSans 480 0 0 0 FrameData[382]
port 313 nsew signal input
flabel metal3 s 0 282888 800 283008 0 FreeSans 480 0 0 0 FrameData[383]
port 314 nsew signal input
flabel metal3 s 0 212168 800 212288 0 FreeSans 480 0 0 0 FrameData[384]
port 315 nsew signal input
flabel metal3 s 0 213528 800 213648 0 FreeSans 480 0 0 0 FrameData[385]
port 316 nsew signal input
flabel metal3 s 0 214208 800 214328 0 FreeSans 480 0 0 0 FrameData[386]
port 317 nsew signal input
flabel metal3 s 0 214888 800 215008 0 FreeSans 480 0 0 0 FrameData[387]
port 318 nsew signal input
flabel metal3 s 0 216248 800 216368 0 FreeSans 480 0 0 0 FrameData[388]
port 319 nsew signal input
flabel metal3 s 0 216928 800 217048 0 FreeSans 480 0 0 0 FrameData[389]
port 320 nsew signal input
flabel metal3 s 0 712648 800 712768 0 FreeSans 480 0 0 0 FrameData[38]
port 321 nsew signal input
flabel metal3 s 0 217608 800 217728 0 FreeSans 480 0 0 0 FrameData[390]
port 322 nsew signal input
flabel metal3 s 0 218288 800 218408 0 FreeSans 480 0 0 0 FrameData[391]
port 323 nsew signal input
flabel metal3 s 0 218968 800 219088 0 FreeSans 480 0 0 0 FrameData[392]
port 324 nsew signal input
flabel metal3 s 0 220328 800 220448 0 FreeSans 480 0 0 0 FrameData[393]
port 325 nsew signal input
flabel metal3 s 0 221008 800 221128 0 FreeSans 480 0 0 0 FrameData[394]
port 326 nsew signal input
flabel metal3 s 0 221688 800 221808 0 FreeSans 480 0 0 0 FrameData[395]
port 327 nsew signal input
flabel metal3 s 0 222368 800 222488 0 FreeSans 480 0 0 0 FrameData[396]
port 328 nsew signal input
flabel metal3 s 0 223048 800 223168 0 FreeSans 480 0 0 0 FrameData[397]
port 329 nsew signal input
flabel metal3 s 0 224408 800 224528 0 FreeSans 480 0 0 0 FrameData[398]
port 330 nsew signal input
flabel metal3 s 0 225088 800 225208 0 FreeSans 480 0 0 0 FrameData[399]
port 331 nsew signal input
flabel metal3 s 0 713328 800 713448 0 FreeSans 480 0 0 0 FrameData[39]
port 332 nsew signal input
flabel metal2 s 21914 755700 21970 756500 0 FreeSans 224 90 0 0 FrameData[3]
port 333 nsew signal input
flabel metal3 s 0 225768 800 225888 0 FreeSans 480 0 0 0 FrameData[400]
port 334 nsew signal input
flabel metal3 s 0 226448 800 226568 0 FreeSans 480 0 0 0 FrameData[401]
port 335 nsew signal input
flabel metal3 s 0 227128 800 227248 0 FreeSans 480 0 0 0 FrameData[402]
port 336 nsew signal input
flabel metal3 s 0 228488 800 228608 0 FreeSans 480 0 0 0 FrameData[403]
port 337 nsew signal input
flabel metal3 s 0 229168 800 229288 0 FreeSans 480 0 0 0 FrameData[404]
port 338 nsew signal input
flabel metal3 s 0 229848 800 229968 0 FreeSans 480 0 0 0 FrameData[405]
port 339 nsew signal input
flabel metal3 s 0 230528 800 230648 0 FreeSans 480 0 0 0 FrameData[406]
port 340 nsew signal input
flabel metal3 s 0 231208 800 231328 0 FreeSans 480 0 0 0 FrameData[407]
port 341 nsew signal input
flabel metal3 s 0 232568 800 232688 0 FreeSans 480 0 0 0 FrameData[408]
port 342 nsew signal input
flabel metal3 s 0 233248 800 233368 0 FreeSans 480 0 0 0 FrameData[409]
port 343 nsew signal input
flabel metal3 s 0 714008 800 714128 0 FreeSans 480 0 0 0 FrameData[40]
port 344 nsew signal input
flabel metal3 s 0 233928 800 234048 0 FreeSans 480 0 0 0 FrameData[410]
port 345 nsew signal input
flabel metal3 s 0 234608 800 234728 0 FreeSans 480 0 0 0 FrameData[411]
port 346 nsew signal input
flabel metal3 s 0 235288 800 235408 0 FreeSans 480 0 0 0 FrameData[412]
port 347 nsew signal input
flabel metal3 s 0 236648 800 236768 0 FreeSans 480 0 0 0 FrameData[413]
port 348 nsew signal input
flabel metal3 s 0 237328 800 237448 0 FreeSans 480 0 0 0 FrameData[414]
port 349 nsew signal input
flabel metal3 s 0 238008 800 238128 0 FreeSans 480 0 0 0 FrameData[415]
port 350 nsew signal input
flabel metal3 s 0 167968 800 168088 0 FreeSans 480 0 0 0 FrameData[416]
port 351 nsew signal input
flabel metal3 s 0 168648 800 168768 0 FreeSans 480 0 0 0 FrameData[417]
port 352 nsew signal input
flabel metal3 s 0 169328 800 169448 0 FreeSans 480 0 0 0 FrameData[418]
port 353 nsew signal input
flabel metal3 s 0 170008 800 170128 0 FreeSans 480 0 0 0 FrameData[419]
port 354 nsew signal input
flabel metal3 s 0 715368 800 715488 0 FreeSans 480 0 0 0 FrameData[41]
port 355 nsew signal input
flabel metal3 s 0 170688 800 170808 0 FreeSans 480 0 0 0 FrameData[420]
port 356 nsew signal input
flabel metal3 s 0 172048 800 172168 0 FreeSans 480 0 0 0 FrameData[421]
port 357 nsew signal input
flabel metal3 s 0 172728 800 172848 0 FreeSans 480 0 0 0 FrameData[422]
port 358 nsew signal input
flabel metal3 s 0 173408 800 173528 0 FreeSans 480 0 0 0 FrameData[423]
port 359 nsew signal input
flabel metal3 s 0 174088 800 174208 0 FreeSans 480 0 0 0 FrameData[424]
port 360 nsew signal input
flabel metal3 s 0 174768 800 174888 0 FreeSans 480 0 0 0 FrameData[425]
port 361 nsew signal input
flabel metal3 s 0 176128 800 176248 0 FreeSans 480 0 0 0 FrameData[426]
port 362 nsew signal input
flabel metal3 s 0 176808 800 176928 0 FreeSans 480 0 0 0 FrameData[427]
port 363 nsew signal input
flabel metal3 s 0 177488 800 177608 0 FreeSans 480 0 0 0 FrameData[428]
port 364 nsew signal input
flabel metal3 s 0 178168 800 178288 0 FreeSans 480 0 0 0 FrameData[429]
port 365 nsew signal input
flabel metal3 s 0 716048 800 716168 0 FreeSans 480 0 0 0 FrameData[42]
port 366 nsew signal input
flabel metal3 s 0 178848 800 178968 0 FreeSans 480 0 0 0 FrameData[430]
port 367 nsew signal input
flabel metal3 s 0 180208 800 180328 0 FreeSans 480 0 0 0 FrameData[431]
port 368 nsew signal input
flabel metal3 s 0 180888 800 181008 0 FreeSans 480 0 0 0 FrameData[432]
port 369 nsew signal input
flabel metal3 s 0 181568 800 181688 0 FreeSans 480 0 0 0 FrameData[433]
port 370 nsew signal input
flabel metal3 s 0 182248 800 182368 0 FreeSans 480 0 0 0 FrameData[434]
port 371 nsew signal input
flabel metal3 s 0 182928 800 183048 0 FreeSans 480 0 0 0 FrameData[435]
port 372 nsew signal input
flabel metal3 s 0 184288 800 184408 0 FreeSans 480 0 0 0 FrameData[436]
port 373 nsew signal input
flabel metal3 s 0 184968 800 185088 0 FreeSans 480 0 0 0 FrameData[437]
port 374 nsew signal input
flabel metal3 s 0 185648 800 185768 0 FreeSans 480 0 0 0 FrameData[438]
port 375 nsew signal input
flabel metal3 s 0 186328 800 186448 0 FreeSans 480 0 0 0 FrameData[439]
port 376 nsew signal input
flabel metal3 s 0 716728 800 716848 0 FreeSans 480 0 0 0 FrameData[43]
port 377 nsew signal input
flabel metal3 s 0 187008 800 187128 0 FreeSans 480 0 0 0 FrameData[440]
port 378 nsew signal input
flabel metal3 s 0 188368 800 188488 0 FreeSans 480 0 0 0 FrameData[441]
port 379 nsew signal input
flabel metal3 s 0 189048 800 189168 0 FreeSans 480 0 0 0 FrameData[442]
port 380 nsew signal input
flabel metal3 s 0 189728 800 189848 0 FreeSans 480 0 0 0 FrameData[443]
port 381 nsew signal input
flabel metal3 s 0 190408 800 190528 0 FreeSans 480 0 0 0 FrameData[444]
port 382 nsew signal input
flabel metal3 s 0 191088 800 191208 0 FreeSans 480 0 0 0 FrameData[445]
port 383 nsew signal input
flabel metal3 s 0 192448 800 192568 0 FreeSans 480 0 0 0 FrameData[446]
port 384 nsew signal input
flabel metal3 s 0 193128 800 193248 0 FreeSans 480 0 0 0 FrameData[447]
port 385 nsew signal input
flabel metal3 s 0 123088 800 123208 0 FreeSans 480 0 0 0 FrameData[448]
port 386 nsew signal input
flabel metal3 s 0 123768 800 123888 0 FreeSans 480 0 0 0 FrameData[449]
port 387 nsew signal input
flabel metal3 s 0 717408 800 717528 0 FreeSans 480 0 0 0 FrameData[44]
port 388 nsew signal input
flabel metal3 s 0 124448 800 124568 0 FreeSans 480 0 0 0 FrameData[450]
port 389 nsew signal input
flabel metal3 s 0 125128 800 125248 0 FreeSans 480 0 0 0 FrameData[451]
port 390 nsew signal input
flabel metal3 s 0 125808 800 125928 0 FreeSans 480 0 0 0 FrameData[452]
port 391 nsew signal input
flabel metal3 s 0 127168 800 127288 0 FreeSans 480 0 0 0 FrameData[453]
port 392 nsew signal input
flabel metal3 s 0 127848 800 127968 0 FreeSans 480 0 0 0 FrameData[454]
port 393 nsew signal input
flabel metal3 s 0 128528 800 128648 0 FreeSans 480 0 0 0 FrameData[455]
port 394 nsew signal input
flabel metal3 s 0 129208 800 129328 0 FreeSans 480 0 0 0 FrameData[456]
port 395 nsew signal input
flabel metal3 s 0 129888 800 130008 0 FreeSans 480 0 0 0 FrameData[457]
port 396 nsew signal input
flabel metal3 s 0 131248 800 131368 0 FreeSans 480 0 0 0 FrameData[458]
port 397 nsew signal input
flabel metal3 s 0 131928 800 132048 0 FreeSans 480 0 0 0 FrameData[459]
port 398 nsew signal input
flabel metal3 s 0 718088 800 718208 0 FreeSans 480 0 0 0 FrameData[45]
port 399 nsew signal input
flabel metal3 s 0 132608 800 132728 0 FreeSans 480 0 0 0 FrameData[460]
port 400 nsew signal input
flabel metal3 s 0 133288 800 133408 0 FreeSans 480 0 0 0 FrameData[461]
port 401 nsew signal input
flabel metal3 s 0 133968 800 134088 0 FreeSans 480 0 0 0 FrameData[462]
port 402 nsew signal input
flabel metal3 s 0 135328 800 135448 0 FreeSans 480 0 0 0 FrameData[463]
port 403 nsew signal input
flabel metal3 s 0 136008 800 136128 0 FreeSans 480 0 0 0 FrameData[464]
port 404 nsew signal input
flabel metal3 s 0 136688 800 136808 0 FreeSans 480 0 0 0 FrameData[465]
port 405 nsew signal input
flabel metal3 s 0 137368 800 137488 0 FreeSans 480 0 0 0 FrameData[466]
port 406 nsew signal input
flabel metal3 s 0 138048 800 138168 0 FreeSans 480 0 0 0 FrameData[467]
port 407 nsew signal input
flabel metal3 s 0 139408 800 139528 0 FreeSans 480 0 0 0 FrameData[468]
port 408 nsew signal input
flabel metal3 s 0 140088 800 140208 0 FreeSans 480 0 0 0 FrameData[469]
port 409 nsew signal input
flabel metal3 s 0 719448 800 719568 0 FreeSans 480 0 0 0 FrameData[46]
port 410 nsew signal input
flabel metal3 s 0 140768 800 140888 0 FreeSans 480 0 0 0 FrameData[470]
port 411 nsew signal input
flabel metal3 s 0 141448 800 141568 0 FreeSans 480 0 0 0 FrameData[471]
port 412 nsew signal input
flabel metal3 s 0 142128 800 142248 0 FreeSans 480 0 0 0 FrameData[472]
port 413 nsew signal input
flabel metal3 s 0 143488 800 143608 0 FreeSans 480 0 0 0 FrameData[473]
port 414 nsew signal input
flabel metal3 s 0 144168 800 144288 0 FreeSans 480 0 0 0 FrameData[474]
port 415 nsew signal input
flabel metal3 s 0 144848 800 144968 0 FreeSans 480 0 0 0 FrameData[475]
port 416 nsew signal input
flabel metal3 s 0 145528 800 145648 0 FreeSans 480 0 0 0 FrameData[476]
port 417 nsew signal input
flabel metal3 s 0 146208 800 146328 0 FreeSans 480 0 0 0 FrameData[477]
port 418 nsew signal input
flabel metal3 s 0 147568 800 147688 0 FreeSans 480 0 0 0 FrameData[478]
port 419 nsew signal input
flabel metal3 s 0 148248 800 148368 0 FreeSans 480 0 0 0 FrameData[479]
port 420 nsew signal input
flabel metal3 s 0 720128 800 720248 0 FreeSans 480 0 0 0 FrameData[47]
port 421 nsew signal input
flabel metal3 s 0 44208 800 44328 0 FreeSans 480 0 0 0 FrameData[480]
port 422 nsew signal input
flabel metal3 s 0 60528 800 60648 0 FreeSans 480 0 0 0 FrameData[481]
port 423 nsew signal input
flabel metal3 s 0 62568 800 62688 0 FreeSans 480 0 0 0 FrameData[482]
port 424 nsew signal input
flabel metal3 s 0 68688 800 68808 0 FreeSans 480 0 0 0 FrameData[483]
port 425 nsew signal input
flabel metal3 s 0 74128 800 74248 0 FreeSans 480 0 0 0 FrameData[484]
port 426 nsew signal input
flabel metal3 s 0 59848 800 59968 0 FreeSans 480 0 0 0 FrameData[485]
port 427 nsew signal input
flabel metal3 s 0 73448 800 73568 0 FreeSans 480 0 0 0 FrameData[486]
port 428 nsew signal input
flabel metal3 s 0 59168 800 59288 0 FreeSans 480 0 0 0 FrameData[487]
port 429 nsew signal input
flabel metal3 s 0 74808 800 74928 0 FreeSans 480 0 0 0 FrameData[488]
port 430 nsew signal input
flabel metal3 s 0 58488 800 58608 0 FreeSans 480 0 0 0 FrameData[489]
port 431 nsew signal input
flabel metal3 s 0 720808 800 720928 0 FreeSans 480 0 0 0 FrameData[48]
port 432 nsew signal input
flabel metal3 s 0 66648 800 66768 0 FreeSans 480 0 0 0 FrameData[490]
port 433 nsew signal input
flabel metal3 s 0 72768 800 72888 0 FreeSans 480 0 0 0 FrameData[491]
port 434 nsew signal input
flabel metal3 s 0 72088 800 72208 0 FreeSans 480 0 0 0 FrameData[492]
port 435 nsew signal input
flabel metal3 s 0 56448 800 56568 0 FreeSans 480 0 0 0 FrameData[493]
port 436 nsew signal input
flabel metal3 s 0 75488 800 75608 0 FreeSans 480 0 0 0 FrameData[494]
port 437 nsew signal input
flabel metal3 s 0 67328 800 67448 0 FreeSans 480 0 0 0 FrameData[495]
port 438 nsew signal input
flabel metal3 s 0 76168 800 76288 0 FreeSans 480 0 0 0 FrameData[496]
port 439 nsew signal input
flabel metal3 s 0 91808 800 91928 0 FreeSans 480 0 0 0 FrameData[497]
port 440 nsew signal input
flabel metal3 s 0 92488 800 92608 0 FreeSans 480 0 0 0 FrameData[498]
port 441 nsew signal input
flabel metal3 s 0 93168 800 93288 0 FreeSans 480 0 0 0 FrameData[499]
port 442 nsew signal input
flabel metal3 s 0 721488 800 721608 0 FreeSans 480 0 0 0 FrameData[49]
port 443 nsew signal input
flabel metal2 s 16762 755700 16818 756500 0 FreeSans 224 90 0 0 FrameData[4]
port 444 nsew signal input
flabel metal3 s 0 93848 800 93968 0 FreeSans 480 0 0 0 FrameData[500]
port 445 nsew signal input
flabel metal3 s 0 95208 800 95328 0 FreeSans 480 0 0 0 FrameData[501]
port 446 nsew signal input
flabel metal3 s 0 95888 800 96008 0 FreeSans 480 0 0 0 FrameData[502]
port 447 nsew signal input
flabel metal3 s 0 96568 800 96688 0 FreeSans 480 0 0 0 FrameData[503]
port 448 nsew signal input
flabel metal3 s 0 97248 800 97368 0 FreeSans 480 0 0 0 FrameData[504]
port 449 nsew signal input
flabel metal3 s 0 97928 800 98048 0 FreeSans 480 0 0 0 FrameData[505]
port 450 nsew signal input
flabel metal3 s 0 99288 800 99408 0 FreeSans 480 0 0 0 FrameData[506]
port 451 nsew signal input
flabel metal3 s 0 99968 800 100088 0 FreeSans 480 0 0 0 FrameData[507]
port 452 nsew signal input
flabel metal3 s 0 100648 800 100768 0 FreeSans 480 0 0 0 FrameData[508]
port 453 nsew signal input
flabel metal3 s 0 101328 800 101448 0 FreeSans 480 0 0 0 FrameData[509]
port 454 nsew signal input
flabel metal3 s 0 722168 800 722288 0 FreeSans 480 0 0 0 FrameData[50]
port 455 nsew signal input
flabel metal3 s 0 102008 800 102128 0 FreeSans 480 0 0 0 FrameData[510]
port 456 nsew signal input
flabel metal3 s 0 103368 800 103488 0 FreeSans 480 0 0 0 FrameData[511]
port 457 nsew signal input
flabel metal3 s 0 36728 800 36848 0 FreeSans 480 0 0 0 FrameData[512]
port 458 nsew signal input
flabel metal3 s 0 34008 800 34128 0 FreeSans 480 0 0 0 FrameData[513]
port 459 nsew signal input
flabel metal3 s 0 34688 800 34808 0 FreeSans 480 0 0 0 FrameData[514]
port 460 nsew signal input
flabel metal3 s 0 35368 800 35488 0 FreeSans 480 0 0 0 FrameData[515]
port 461 nsew signal input
flabel metal3 s 0 36048 800 36168 0 FreeSans 480 0 0 0 FrameData[516]
port 462 nsew signal input
flabel metal3 s 0 37408 800 37528 0 FreeSans 480 0 0 0 FrameData[517]
port 463 nsew signal input
flabel metal3 s 0 38088 800 38208 0 FreeSans 480 0 0 0 FrameData[518]
port 464 nsew signal input
flabel metal3 s 0 38768 800 38888 0 FreeSans 480 0 0 0 FrameData[519]
port 465 nsew signal input
flabel metal3 s 0 723528 800 723648 0 FreeSans 480 0 0 0 FrameData[51]
port 466 nsew signal input
flabel metal3 s 0 39448 800 39568 0 FreeSans 480 0 0 0 FrameData[520]
port 467 nsew signal input
flabel metal3 s 0 40128 800 40248 0 FreeSans 480 0 0 0 FrameData[521]
port 468 nsew signal input
flabel metal3 s 0 40808 800 40928 0 FreeSans 480 0 0 0 FrameData[522]
port 469 nsew signal input
flabel metal3 s 0 41488 800 41608 0 FreeSans 480 0 0 0 FrameData[523]
port 470 nsew signal input
flabel metal3 s 0 42168 800 42288 0 FreeSans 480 0 0 0 FrameData[524]
port 471 nsew signal input
flabel metal3 s 0 42848 800 42968 0 FreeSans 480 0 0 0 FrameData[525]
port 472 nsew signal input
flabel metal3 s 0 43528 800 43648 0 FreeSans 480 0 0 0 FrameData[526]
port 473 nsew signal input
flabel metal3 s 0 44888 800 45008 0 FreeSans 480 0 0 0 FrameData[527]
port 474 nsew signal input
flabel metal3 s 0 45568 800 45688 0 FreeSans 480 0 0 0 FrameData[528]
port 475 nsew signal input
flabel metal3 s 0 46248 800 46368 0 FreeSans 480 0 0 0 FrameData[529]
port 476 nsew signal input
flabel metal3 s 0 724208 800 724328 0 FreeSans 480 0 0 0 FrameData[52]
port 477 nsew signal input
flabel metal3 s 0 46928 800 47048 0 FreeSans 480 0 0 0 FrameData[530]
port 478 nsew signal input
flabel metal3 s 0 47608 800 47728 0 FreeSans 480 0 0 0 FrameData[531]
port 479 nsew signal input
flabel metal3 s 0 48968 800 49088 0 FreeSans 480 0 0 0 FrameData[532]
port 480 nsew signal input
flabel metal3 s 0 49648 800 49768 0 FreeSans 480 0 0 0 FrameData[533]
port 481 nsew signal input
flabel metal3 s 0 50328 800 50448 0 FreeSans 480 0 0 0 FrameData[534]
port 482 nsew signal input
flabel metal3 s 0 51008 800 51128 0 FreeSans 480 0 0 0 FrameData[535]
port 483 nsew signal input
flabel metal3 s 0 51688 800 51808 0 FreeSans 480 0 0 0 FrameData[536]
port 484 nsew signal input
flabel metal3 s 0 53048 800 53168 0 FreeSans 480 0 0 0 FrameData[537]
port 485 nsew signal input
flabel metal3 s 0 53728 800 53848 0 FreeSans 480 0 0 0 FrameData[538]
port 486 nsew signal input
flabel metal3 s 0 54408 800 54528 0 FreeSans 480 0 0 0 FrameData[539]
port 487 nsew signal input
flabel metal3 s 0 724888 800 725008 0 FreeSans 480 0 0 0 FrameData[53]
port 488 nsew signal input
flabel metal3 s 0 55088 800 55208 0 FreeSans 480 0 0 0 FrameData[540]
port 489 nsew signal input
flabel metal3 s 0 55768 800 55888 0 FreeSans 480 0 0 0 FrameData[541]
port 490 nsew signal input
flabel metal3 s 0 57128 800 57248 0 FreeSans 480 0 0 0 FrameData[542]
port 491 nsew signal input
flabel metal3 s 0 57808 800 57928 0 FreeSans 480 0 0 0 FrameData[543]
port 492 nsew signal input
flabel metal2 s 22558 0 22614 800 0 FreeSans 224 90 0 0 FrameData[544]
port 493 nsew signal input
flabel metal2 s 21270 0 21326 800 0 FreeSans 224 90 0 0 FrameData[545]
port 494 nsew signal input
flabel metal2 s 20626 0 20682 800 0 FreeSans 224 90 0 0 FrameData[546]
port 495 nsew signal input
flabel metal2 s 21914 0 21970 800 0 FreeSans 224 90 0 0 FrameData[547]
port 496 nsew signal input
flabel metal3 s 0 4768 800 4888 0 FreeSans 480 0 0 0 FrameData[548]
port 497 nsew signal input
flabel metal3 s 0 7488 800 7608 0 FreeSans 480 0 0 0 FrameData[549]
port 498 nsew signal input
flabel metal3 s 0 725568 800 725688 0 FreeSans 480 0 0 0 FrameData[54]
port 499 nsew signal input
flabel metal3 s 0 8 800 128 0 FreeSans 480 0 0 0 FrameData[550]
port 500 nsew signal input
flabel metal3 s 0 688 800 808 0 FreeSans 480 0 0 0 FrameData[551]
port 501 nsew signal input
flabel metal3 s 0 9528 800 9648 0 FreeSans 480 0 0 0 FrameData[552]
port 502 nsew signal input
flabel metal3 s 0 3408 800 3528 0 FreeSans 480 0 0 0 FrameData[553]
port 503 nsew signal input
flabel metal3 s 0 5448 800 5568 0 FreeSans 480 0 0 0 FrameData[554]
port 504 nsew signal input
flabel metal3 s 0 10208 800 10328 0 FreeSans 480 0 0 0 FrameData[555]
port 505 nsew signal input
flabel metal3 s 0 6128 800 6248 0 FreeSans 480 0 0 0 FrameData[556]
port 506 nsew signal input
flabel metal3 s 0 6808 800 6928 0 FreeSans 480 0 0 0 FrameData[557]
port 507 nsew signal input
flabel metal3 s 0 2048 800 2168 0 FreeSans 480 0 0 0 FrameData[558]
port 508 nsew signal input
flabel metal3 s 0 10888 800 11008 0 FreeSans 480 0 0 0 FrameData[559]
port 509 nsew signal input
flabel metal3 s 0 726248 800 726368 0 FreeSans 480 0 0 0 FrameData[55]
port 510 nsew signal input
flabel metal3 s 0 8168 800 8288 0 FreeSans 480 0 0 0 FrameData[560]
port 511 nsew signal input
flabel metal3 s 0 11568 800 11688 0 FreeSans 480 0 0 0 FrameData[561]
port 512 nsew signal input
flabel metal3 s 0 1368 800 1488 0 FreeSans 480 0 0 0 FrameData[562]
port 513 nsew signal input
flabel metal3 s 0 8848 800 8968 0 FreeSans 480 0 0 0 FrameData[563]
port 514 nsew signal input
flabel metal3 s 0 12248 800 12368 0 FreeSans 480 0 0 0 FrameData[564]
port 515 nsew signal input
flabel metal3 s 0 4088 800 4208 0 FreeSans 480 0 0 0 FrameData[565]
port 516 nsew signal input
flabel metal3 s 0 2728 800 2848 0 FreeSans 480 0 0 0 FrameData[566]
port 517 nsew signal input
flabel metal3 s 0 12928 800 13048 0 FreeSans 480 0 0 0 FrameData[567]
port 518 nsew signal input
flabel metal3 s 0 13608 800 13728 0 FreeSans 480 0 0 0 FrameData[568]
port 519 nsew signal input
flabel metal3 s 0 14288 800 14408 0 FreeSans 480 0 0 0 FrameData[569]
port 520 nsew signal input
flabel metal3 s 0 727608 800 727728 0 FreeSans 480 0 0 0 FrameData[56]
port 521 nsew signal input
flabel metal3 s 0 33328 800 33448 0 FreeSans 480 0 0 0 FrameData[570]
port 522 nsew signal input
flabel metal3 s 0 14968 800 15088 0 FreeSans 480 0 0 0 FrameData[571]
port 523 nsew signal input
flabel metal3 s 0 32648 800 32768 0 FreeSans 480 0 0 0 FrameData[572]
port 524 nsew signal input
flabel metal3 s 0 17008 800 17128 0 FreeSans 480 0 0 0 FrameData[573]
port 525 nsew signal input
flabel metal3 s 0 15648 800 15768 0 FreeSans 480 0 0 0 FrameData[574]
port 526 nsew signal input
flabel metal3 s 0 16328 800 16448 0 FreeSans 480 0 0 0 FrameData[575]
port 527 nsew signal input
flabel metal3 s 0 728288 800 728408 0 FreeSans 480 0 0 0 FrameData[57]
port 528 nsew signal input
flabel metal3 s 0 728968 800 729088 0 FreeSans 480 0 0 0 FrameData[58]
port 529 nsew signal input
flabel metal3 s 0 729648 800 729768 0 FreeSans 480 0 0 0 FrameData[59]
port 530 nsew signal input
flabel metal2 s 25778 755700 25834 756500 0 FreeSans 224 90 0 0 FrameData[5]
port 531 nsew signal input
flabel metal3 s 0 730328 800 730448 0 FreeSans 480 0 0 0 FrameData[60]
port 532 nsew signal input
flabel metal3 s 0 731688 800 731808 0 FreeSans 480 0 0 0 FrameData[61]
port 533 nsew signal input
flabel metal3 s 0 732368 800 732488 0 FreeSans 480 0 0 0 FrameData[62]
port 534 nsew signal input
flabel metal3 s 0 733048 800 733168 0 FreeSans 480 0 0 0 FrameData[63]
port 535 nsew signal input
flabel metal3 s 0 663008 800 663128 0 FreeSans 480 0 0 0 FrameData[64]
port 536 nsew signal input
flabel metal3 s 0 663688 800 663808 0 FreeSans 480 0 0 0 FrameData[65]
port 537 nsew signal input
flabel metal3 s 0 664368 800 664488 0 FreeSans 480 0 0 0 FrameData[66]
port 538 nsew signal input
flabel metal3 s 0 665048 800 665168 0 FreeSans 480 0 0 0 FrameData[67]
port 539 nsew signal input
flabel metal3 s 0 665728 800 665848 0 FreeSans 480 0 0 0 FrameData[68]
port 540 nsew signal input
flabel metal3 s 0 667088 800 667208 0 FreeSans 480 0 0 0 FrameData[69]
port 541 nsew signal input
flabel metal2 s 34794 755700 34850 756500 0 FreeSans 224 90 0 0 FrameData[6]
port 542 nsew signal input
flabel metal3 s 0 667768 800 667888 0 FreeSans 480 0 0 0 FrameData[70]
port 543 nsew signal input
flabel metal3 s 0 668448 800 668568 0 FreeSans 480 0 0 0 FrameData[71]
port 544 nsew signal input
flabel metal3 s 0 669128 800 669248 0 FreeSans 480 0 0 0 FrameData[72]
port 545 nsew signal input
flabel metal3 s 0 669808 800 669928 0 FreeSans 480 0 0 0 FrameData[73]
port 546 nsew signal input
flabel metal3 s 0 671168 800 671288 0 FreeSans 480 0 0 0 FrameData[74]
port 547 nsew signal input
flabel metal3 s 0 671848 800 671968 0 FreeSans 480 0 0 0 FrameData[75]
port 548 nsew signal input
flabel metal3 s 0 672528 800 672648 0 FreeSans 480 0 0 0 FrameData[76]
port 549 nsew signal input
flabel metal3 s 0 673208 800 673328 0 FreeSans 480 0 0 0 FrameData[77]
port 550 nsew signal input
flabel metal3 s 0 673888 800 674008 0 FreeSans 480 0 0 0 FrameData[78]
port 551 nsew signal input
flabel metal3 s 0 675248 800 675368 0 FreeSans 480 0 0 0 FrameData[79]
port 552 nsew signal input
flabel metal2 s 16118 755700 16174 756500 0 FreeSans 224 90 0 0 FrameData[7]
port 553 nsew signal input
flabel metal3 s 0 675928 800 676048 0 FreeSans 480 0 0 0 FrameData[80]
port 554 nsew signal input
flabel metal3 s 0 676608 800 676728 0 FreeSans 480 0 0 0 FrameData[81]
port 555 nsew signal input
flabel metal3 s 0 677288 800 677408 0 FreeSans 480 0 0 0 FrameData[82]
port 556 nsew signal input
flabel metal3 s 0 677968 800 678088 0 FreeSans 480 0 0 0 FrameData[83]
port 557 nsew signal input
flabel metal3 s 0 679328 800 679448 0 FreeSans 480 0 0 0 FrameData[84]
port 558 nsew signal input
flabel metal3 s 0 680008 800 680128 0 FreeSans 480 0 0 0 FrameData[85]
port 559 nsew signal input
flabel metal3 s 0 680688 800 680808 0 FreeSans 480 0 0 0 FrameData[86]
port 560 nsew signal input
flabel metal3 s 0 681368 800 681488 0 FreeSans 480 0 0 0 FrameData[87]
port 561 nsew signal input
flabel metal3 s 0 682048 800 682168 0 FreeSans 480 0 0 0 FrameData[88]
port 562 nsew signal input
flabel metal3 s 0 683408 800 683528 0 FreeSans 480 0 0 0 FrameData[89]
port 563 nsew signal input
flabel metal2 s 30286 755700 30342 756500 0 FreeSans 224 90 0 0 FrameData[8]
port 564 nsew signal input
flabel metal3 s 0 684088 800 684208 0 FreeSans 480 0 0 0 FrameData[90]
port 565 nsew signal input
flabel metal3 s 0 684768 800 684888 0 FreeSans 480 0 0 0 FrameData[91]
port 566 nsew signal input
flabel metal3 s 0 685448 800 685568 0 FreeSans 480 0 0 0 FrameData[92]
port 567 nsew signal input
flabel metal3 s 0 686128 800 686248 0 FreeSans 480 0 0 0 FrameData[93]
port 568 nsew signal input
flabel metal3 s 0 687488 800 687608 0 FreeSans 480 0 0 0 FrameData[94]
port 569 nsew signal input
flabel metal3 s 0 688168 800 688288 0 FreeSans 480 0 0 0 FrameData[95]
port 570 nsew signal input
flabel metal3 s 0 617448 800 617568 0 FreeSans 480 0 0 0 FrameData[96]
port 571 nsew signal input
flabel metal3 s 0 618808 800 618928 0 FreeSans 480 0 0 0 FrameData[97]
port 572 nsew signal input
flabel metal3 s 0 619488 800 619608 0 FreeSans 480 0 0 0 FrameData[98]
port 573 nsew signal input
flabel metal3 s 0 620168 800 620288 0 FreeSans 480 0 0 0 FrameData[99]
port 574 nsew signal input
flabel metal2 s 33506 755700 33562 756500 0 FreeSans 224 90 0 0 FrameData[9]
port 575 nsew signal input
flabel metal3 s 0 31968 800 32088 0 FreeSans 480 0 0 0 FrameStrobe[0]
port 576 nsew signal input
flabel metal2 s 218978 0 219034 800 0 FreeSans 224 90 0 0 FrameStrobe[100]
port 577 nsew signal input
flabel metal2 s 219622 0 219678 800 0 FreeSans 224 90 0 0 FrameStrobe[101]
port 578 nsew signal input
flabel metal2 s 220266 0 220322 800 0 FreeSans 224 90 0 0 FrameStrobe[102]
port 579 nsew signal input
flabel metal2 s 220910 0 220966 800 0 FreeSans 224 90 0 0 FrameStrobe[103]
port 580 nsew signal input
flabel metal2 s 221554 0 221610 800 0 FreeSans 224 90 0 0 FrameStrobe[104]
port 581 nsew signal input
flabel metal2 s 222842 0 222898 800 0 FreeSans 224 90 0 0 FrameStrobe[105]
port 582 nsew signal input
flabel metal2 s 223486 0 223542 800 0 FreeSans 224 90 0 0 FrameStrobe[106]
port 583 nsew signal input
flabel metal2 s 224130 0 224186 800 0 FreeSans 224 90 0 0 FrameStrobe[107]
port 584 nsew signal input
flabel metal2 s 224774 0 224830 800 0 FreeSans 224 90 0 0 FrameStrobe[108]
port 585 nsew signal input
flabel metal2 s 225418 0 225474 800 0 FreeSans 224 90 0 0 FrameStrobe[109]
port 586 nsew signal input
flabel metal3 s 0 25168 800 25288 0 FreeSans 480 0 0 0 FrameStrobe[10]
port 587 nsew signal input
flabel metal2 s 226062 0 226118 800 0 FreeSans 224 90 0 0 FrameStrobe[110]
port 588 nsew signal input
flabel metal2 s 226706 0 226762 800 0 FreeSans 224 90 0 0 FrameStrobe[111]
port 589 nsew signal input
flabel metal2 s 227994 0 228050 800 0 FreeSans 224 90 0 0 FrameStrobe[112]
port 590 nsew signal input
flabel metal2 s 228638 0 228694 800 0 FreeSans 224 90 0 0 FrameStrobe[113]
port 591 nsew signal input
flabel metal2 s 229282 0 229338 800 0 FreeSans 224 90 0 0 FrameStrobe[114]
port 592 nsew signal input
flabel metal2 s 229926 0 229982 800 0 FreeSans 224 90 0 0 FrameStrobe[115]
port 593 nsew signal input
flabel metal2 s 230570 0 230626 800 0 FreeSans 224 90 0 0 FrameStrobe[116]
port 594 nsew signal input
flabel metal2 s 231214 0 231270 800 0 FreeSans 224 90 0 0 FrameStrobe[117]
port 595 nsew signal input
flabel metal2 s 231858 0 231914 800 0 FreeSans 224 90 0 0 FrameStrobe[118]
port 596 nsew signal input
flabel metal2 s 233146 0 233202 800 0 FreeSans 224 90 0 0 FrameStrobe[119]
port 597 nsew signal input
flabel metal3 s 0 31288 800 31408 0 FreeSans 480 0 0 0 FrameStrobe[11]
port 598 nsew signal input
flabel metal2 s 259550 0 259606 800 0 FreeSans 224 90 0 0 FrameStrobe[120]
port 599 nsew signal input
flabel metal2 s 260838 0 260894 800 0 FreeSans 224 90 0 0 FrameStrobe[121]
port 600 nsew signal input
flabel metal2 s 261482 0 261538 800 0 FreeSans 224 90 0 0 FrameStrobe[122]
port 601 nsew signal input
flabel metal2 s 262126 0 262182 800 0 FreeSans 224 90 0 0 FrameStrobe[123]
port 602 nsew signal input
flabel metal2 s 262770 0 262826 800 0 FreeSans 224 90 0 0 FrameStrobe[124]
port 603 nsew signal input
flabel metal2 s 263414 0 263470 800 0 FreeSans 224 90 0 0 FrameStrobe[125]
port 604 nsew signal input
flabel metal2 s 264058 0 264114 800 0 FreeSans 224 90 0 0 FrameStrobe[126]
port 605 nsew signal input
flabel metal2 s 264702 0 264758 800 0 FreeSans 224 90 0 0 FrameStrobe[127]
port 606 nsew signal input
flabel metal2 s 265990 0 266046 800 0 FreeSans 224 90 0 0 FrameStrobe[128]
port 607 nsew signal input
flabel metal2 s 266634 0 266690 800 0 FreeSans 224 90 0 0 FrameStrobe[129]
port 608 nsew signal input
flabel metal3 s 0 19048 800 19168 0 FreeSans 480 0 0 0 FrameStrobe[12]
port 609 nsew signal input
flabel metal2 s 267278 0 267334 800 0 FreeSans 224 90 0 0 FrameStrobe[130]
port 610 nsew signal input
flabel metal2 s 267922 0 267978 800 0 FreeSans 224 90 0 0 FrameStrobe[131]
port 611 nsew signal input
flabel metal2 s 268566 0 268622 800 0 FreeSans 224 90 0 0 FrameStrobe[132]
port 612 nsew signal input
flabel metal2 s 269210 0 269266 800 0 FreeSans 224 90 0 0 FrameStrobe[133]
port 613 nsew signal input
flabel metal2 s 269854 0 269910 800 0 FreeSans 224 90 0 0 FrameStrobe[134]
port 614 nsew signal input
flabel metal2 s 271142 0 271198 800 0 FreeSans 224 90 0 0 FrameStrobe[135]
port 615 nsew signal input
flabel metal2 s 271786 0 271842 800 0 FreeSans 224 90 0 0 FrameStrobe[136]
port 616 nsew signal input
flabel metal2 s 272430 0 272486 800 0 FreeSans 224 90 0 0 FrameStrobe[137]
port 617 nsew signal input
flabel metal2 s 273074 0 273130 800 0 FreeSans 224 90 0 0 FrameStrobe[138]
port 618 nsew signal input
flabel metal2 s 273718 0 273774 800 0 FreeSans 224 90 0 0 FrameStrobe[139]
port 619 nsew signal input
flabel metal3 s 0 20408 800 20528 0 FreeSans 480 0 0 0 FrameStrobe[13]
port 620 nsew signal input
flabel metal2 s 278870 0 278926 800 0 FreeSans 224 90 0 0 FrameStrobe[140]
port 621 nsew signal input
flabel metal2 s 280802 0 280858 800 0 FreeSans 224 90 0 0 FrameStrobe[141]
port 622 nsew signal input
flabel metal2 s 282734 0 282790 800 0 FreeSans 224 90 0 0 FrameStrobe[142]
port 623 nsew signal input
flabel metal2 s 285310 0 285366 800 0 FreeSans 224 90 0 0 FrameStrobe[143]
port 624 nsew signal input
flabel metal2 s 287242 0 287298 800 0 FreeSans 224 90 0 0 FrameStrobe[144]
port 625 nsew signal input
flabel metal2 s 289174 0 289230 800 0 FreeSans 224 90 0 0 FrameStrobe[145]
port 626 nsew signal input
flabel metal2 s 291106 0 291162 800 0 FreeSans 224 90 0 0 FrameStrobe[146]
port 627 nsew signal input
flabel metal2 s 293682 0 293738 800 0 FreeSans 224 90 0 0 FrameStrobe[147]
port 628 nsew signal input
flabel metal2 s 295614 0 295670 800 0 FreeSans 224 90 0 0 FrameStrobe[148]
port 629 nsew signal input
flabel metal2 s 297546 0 297602 800 0 FreeSans 224 90 0 0 FrameStrobe[149]
port 630 nsew signal input
flabel metal3 s 0 21088 800 21208 0 FreeSans 480 0 0 0 FrameStrobe[14]
port 631 nsew signal input
flabel metal2 s 300122 0 300178 800 0 FreeSans 224 90 0 0 FrameStrobe[150]
port 632 nsew signal input
flabel metal2 s 302054 0 302110 800 0 FreeSans 224 90 0 0 FrameStrobe[151]
port 633 nsew signal input
flabel metal2 s 303986 0 304042 800 0 FreeSans 224 90 0 0 FrameStrobe[152]
port 634 nsew signal input
flabel metal2 s 305918 0 305974 800 0 FreeSans 224 90 0 0 FrameStrobe[153]
port 635 nsew signal input
flabel metal2 s 308494 0 308550 800 0 FreeSans 224 90 0 0 FrameStrobe[154]
port 636 nsew signal input
flabel metal2 s 310426 0 310482 800 0 FreeSans 224 90 0 0 FrameStrobe[155]
port 637 nsew signal input
flabel metal2 s 312358 0 312414 800 0 FreeSans 224 90 0 0 FrameStrobe[156]
port 638 nsew signal input
flabel metal2 s 314934 0 314990 800 0 FreeSans 224 90 0 0 FrameStrobe[157]
port 639 nsew signal input
flabel metal2 s 316866 0 316922 800 0 FreeSans 224 90 0 0 FrameStrobe[158]
port 640 nsew signal input
flabel metal2 s 318798 0 318854 800 0 FreeSans 224 90 0 0 FrameStrobe[159]
port 641 nsew signal input
flabel metal3 s 0 26528 800 26648 0 FreeSans 480 0 0 0 FrameStrobe[15]
port 642 nsew signal input
flabel metal2 s 345846 0 345902 800 0 FreeSans 224 90 0 0 FrameStrobe[160]
port 643 nsew signal input
flabel metal2 s 346490 0 346546 800 0 FreeSans 224 90 0 0 FrameStrobe[161]
port 644 nsew signal input
flabel metal2 s 347134 0 347190 800 0 FreeSans 224 90 0 0 FrameStrobe[162]
port 645 nsew signal input
flabel metal2 s 347778 0 347834 800 0 FreeSans 224 90 0 0 FrameStrobe[163]
port 646 nsew signal input
flabel metal2 s 349066 0 349122 800 0 FreeSans 224 90 0 0 FrameStrobe[164]
port 647 nsew signal input
flabel metal2 s 349710 0 349766 800 0 FreeSans 224 90 0 0 FrameStrobe[165]
port 648 nsew signal input
flabel metal2 s 350354 0 350410 800 0 FreeSans 224 90 0 0 FrameStrobe[166]
port 649 nsew signal input
flabel metal2 s 350998 0 351054 800 0 FreeSans 224 90 0 0 FrameStrobe[167]
port 650 nsew signal input
flabel metal2 s 351642 0 351698 800 0 FreeSans 224 90 0 0 FrameStrobe[168]
port 651 nsew signal input
flabel metal2 s 352286 0 352342 800 0 FreeSans 224 90 0 0 FrameStrobe[169]
port 652 nsew signal input
flabel metal3 s 0 22448 800 22568 0 FreeSans 480 0 0 0 FrameStrobe[16]
port 653 nsew signal input
flabel metal2 s 352930 0 352986 800 0 FreeSans 224 90 0 0 FrameStrobe[170]
port 654 nsew signal input
flabel metal2 s 354218 0 354274 800 0 FreeSans 224 90 0 0 FrameStrobe[171]
port 655 nsew signal input
flabel metal2 s 354862 0 354918 800 0 FreeSans 224 90 0 0 FrameStrobe[172]
port 656 nsew signal input
flabel metal2 s 355506 0 355562 800 0 FreeSans 224 90 0 0 FrameStrobe[173]
port 657 nsew signal input
flabel metal2 s 356150 0 356206 800 0 FreeSans 224 90 0 0 FrameStrobe[174]
port 658 nsew signal input
flabel metal2 s 356794 0 356850 800 0 FreeSans 224 90 0 0 FrameStrobe[175]
port 659 nsew signal input
flabel metal2 s 357438 0 357494 800 0 FreeSans 224 90 0 0 FrameStrobe[176]
port 660 nsew signal input
flabel metal2 s 358082 0 358138 800 0 FreeSans 224 90 0 0 FrameStrobe[177]
port 661 nsew signal input
flabel metal2 s 359370 0 359426 800 0 FreeSans 224 90 0 0 FrameStrobe[178]
port 662 nsew signal input
flabel metal2 s 360014 0 360070 800 0 FreeSans 224 90 0 0 FrameStrobe[179]
port 663 nsew signal input
flabel metal3 s 0 27888 800 28008 0 FreeSans 480 0 0 0 FrameStrobe[17]
port 664 nsew signal input
flabel metal2 s 394146 0 394202 800 0 FreeSans 224 90 0 0 FrameStrobe[180]
port 665 nsew signal input
flabel metal2 s 387062 0 387118 800 0 FreeSans 224 90 0 0 FrameStrobe[181]
port 666 nsew signal input
flabel metal2 s 388350 0 388406 800 0 FreeSans 224 90 0 0 FrameStrobe[182]
port 667 nsew signal input
flabel metal2 s 392858 0 392914 800 0 FreeSans 224 90 0 0 FrameStrobe[183]
port 668 nsew signal input
flabel metal2 s 387706 0 387762 800 0 FreeSans 224 90 0 0 FrameStrobe[184]
port 669 nsew signal input
flabel metal2 s 386418 0 386474 800 0 FreeSans 224 90 0 0 FrameStrobe[185]
port 670 nsew signal input
flabel metal2 s 390926 0 390982 800 0 FreeSans 224 90 0 0 FrameStrobe[186]
port 671 nsew signal input
flabel metal2 s 388994 0 389050 800 0 FreeSans 224 90 0 0 FrameStrobe[187]
port 672 nsew signal input
flabel metal2 s 389638 0 389694 800 0 FreeSans 224 90 0 0 FrameStrobe[188]
port 673 nsew signal input
flabel metal2 s 390282 0 390338 800 0 FreeSans 224 90 0 0 FrameStrobe[189]
port 674 nsew signal input
flabel metal3 s 0 28568 800 28688 0 FreeSans 480 0 0 0 FrameStrobe[18]
port 675 nsew signal input
flabel metal2 s 391570 0 391626 800 0 FreeSans 224 90 0 0 FrameStrobe[190]
port 676 nsew signal input
flabel metal2 s 392214 0 392270 800 0 FreeSans 224 90 0 0 FrameStrobe[191]
port 677 nsew signal input
flabel metal2 s 393502 0 393558 800 0 FreeSans 224 90 0 0 FrameStrobe[192]
port 678 nsew signal input
flabel metal2 s 394790 0 394846 800 0 FreeSans 224 90 0 0 FrameStrobe[193]
port 679 nsew signal input
flabel metal2 s 395434 0 395490 800 0 FreeSans 224 90 0 0 FrameStrobe[194]
port 680 nsew signal input
flabel metal2 s 396722 0 396778 800 0 FreeSans 224 90 0 0 FrameStrobe[195]
port 681 nsew signal input
flabel metal2 s 398010 0 398066 800 0 FreeSans 224 90 0 0 FrameStrobe[196]
port 682 nsew signal input
flabel metal2 s 398654 0 398710 800 0 FreeSans 224 90 0 0 FrameStrobe[197]
port 683 nsew signal input
flabel metal2 s 399942 0 399998 800 0 FreeSans 224 90 0 0 FrameStrobe[198]
port 684 nsew signal input
flabel metal2 s 401230 0 401286 800 0 FreeSans 224 90 0 0 FrameStrobe[199]
port 685 nsew signal input
flabel metal3 s 0 29928 800 30048 0 FreeSans 480 0 0 0 FrameStrobe[19]
port 686 nsew signal input
flabel metal3 s 0 29248 800 29368 0 FreeSans 480 0 0 0 FrameStrobe[1]
port 687 nsew signal input
flabel metal2 s 416042 0 416098 800 0 FreeSans 224 90 0 0 FrameStrobe[200]
port 688 nsew signal input
flabel metal2 s 417330 0 417386 800 0 FreeSans 224 90 0 0 FrameStrobe[201]
port 689 nsew signal input
flabel metal2 s 418618 0 418674 800 0 FreeSans 224 90 0 0 FrameStrobe[202]
port 690 nsew signal input
flabel metal2 s 419906 0 419962 800 0 FreeSans 224 90 0 0 FrameStrobe[203]
port 691 nsew signal input
flabel metal2 s 421194 0 421250 800 0 FreeSans 224 90 0 0 FrameStrobe[204]
port 692 nsew signal input
flabel metal2 s 422482 0 422538 800 0 FreeSans 224 90 0 0 FrameStrobe[205]
port 693 nsew signal input
flabel metal2 s 423770 0 423826 800 0 FreeSans 224 90 0 0 FrameStrobe[206]
port 694 nsew signal input
flabel metal2 s 425702 0 425758 800 0 FreeSans 224 90 0 0 FrameStrobe[207]
port 695 nsew signal input
flabel metal2 s 426990 0 427046 800 0 FreeSans 224 90 0 0 FrameStrobe[208]
port 696 nsew signal input
flabel metal2 s 428278 0 428334 800 0 FreeSans 224 90 0 0 FrameStrobe[209]
port 697 nsew signal input
flabel metal2 s 30930 0 30986 800 0 FreeSans 224 90 0 0 FrameStrobe[20]
port 698 nsew signal input
flabel metal2 s 429566 0 429622 800 0 FreeSans 224 90 0 0 FrameStrobe[210]
port 699 nsew signal input
flabel metal2 s 430854 0 430910 800 0 FreeSans 224 90 0 0 FrameStrobe[211]
port 700 nsew signal input
flabel metal2 s 432142 0 432198 800 0 FreeSans 224 90 0 0 FrameStrobe[212]
port 701 nsew signal input
flabel metal2 s 433430 0 433486 800 0 FreeSans 224 90 0 0 FrameStrobe[213]
port 702 nsew signal input
flabel metal2 s 435362 0 435418 800 0 FreeSans 224 90 0 0 FrameStrobe[214]
port 703 nsew signal input
flabel metal2 s 436650 0 436706 800 0 FreeSans 224 90 0 0 FrameStrobe[215]
port 704 nsew signal input
flabel metal2 s 437938 0 437994 800 0 FreeSans 224 90 0 0 FrameStrobe[216]
port 705 nsew signal input
flabel metal2 s 439226 0 439282 800 0 FreeSans 224 90 0 0 FrameStrobe[217]
port 706 nsew signal input
flabel metal2 s 440514 0 440570 800 0 FreeSans 224 90 0 0 FrameStrobe[218]
port 707 nsew signal input
flabel metal2 s 441802 0 441858 800 0 FreeSans 224 90 0 0 FrameStrobe[219]
port 708 nsew signal input
flabel metal2 s 32218 0 32274 800 0 FreeSans 224 90 0 0 FrameStrobe[21]
port 709 nsew signal input
flabel metal2 s 446310 0 446366 800 0 FreeSans 224 90 0 0 FrameStrobe[220]
port 710 nsew signal input
flabel metal2 s 447598 0 447654 800 0 FreeSans 224 90 0 0 FrameStrobe[221]
port 711 nsew signal input
flabel metal2 s 448886 0 448942 800 0 FreeSans 224 90 0 0 FrameStrobe[222]
port 712 nsew signal input
flabel metal2 s 450818 0 450874 800 0 FreeSans 224 90 0 0 FrameStrobe[223]
port 713 nsew signal input
flabel metal2 s 452106 0 452162 800 0 FreeSans 224 90 0 0 FrameStrobe[224]
port 714 nsew signal input
flabel metal2 s 454038 0 454094 800 0 FreeSans 224 90 0 0 FrameStrobe[225]
port 715 nsew signal input
flabel metal2 s 455326 0 455382 800 0 FreeSans 224 90 0 0 FrameStrobe[226]
port 716 nsew signal input
flabel metal2 s 457258 0 457314 800 0 FreeSans 224 90 0 0 FrameStrobe[227]
port 717 nsew signal input
flabel metal2 s 458546 0 458602 800 0 FreeSans 224 90 0 0 FrameStrobe[228]
port 718 nsew signal input
flabel metal2 s 459834 0 459890 800 0 FreeSans 224 90 0 0 FrameStrobe[229]
port 719 nsew signal input
flabel metal2 s 34150 0 34206 800 0 FreeSans 224 90 0 0 FrameStrobe[22]
port 720 nsew signal input
flabel metal2 s 461766 0 461822 800 0 FreeSans 224 90 0 0 FrameStrobe[230]
port 721 nsew signal input
flabel metal2 s 463054 0 463110 800 0 FreeSans 224 90 0 0 FrameStrobe[231]
port 722 nsew signal input
flabel metal2 s 464986 0 465042 800 0 FreeSans 224 90 0 0 FrameStrobe[232]
port 723 nsew signal input
flabel metal2 s 466274 0 466330 800 0 FreeSans 224 90 0 0 FrameStrobe[233]
port 724 nsew signal input
flabel metal2 s 468206 0 468262 800 0 FreeSans 224 90 0 0 FrameStrobe[234]
port 725 nsew signal input
flabel metal2 s 469494 0 469550 800 0 FreeSans 224 90 0 0 FrameStrobe[235]
port 726 nsew signal input
flabel metal2 s 470782 0 470838 800 0 FreeSans 224 90 0 0 FrameStrobe[236]
port 727 nsew signal input
flabel metal2 s 472714 0 472770 800 0 FreeSans 224 90 0 0 FrameStrobe[237]
port 728 nsew signal input
flabel metal2 s 474002 0 474058 800 0 FreeSans 224 90 0 0 FrameStrobe[238]
port 729 nsew signal input
flabel metal2 s 475934 0 475990 800 0 FreeSans 224 90 0 0 FrameStrobe[239]
port 730 nsew signal input
flabel metal2 s 35438 0 35494 800 0 FreeSans 224 90 0 0 FrameStrobe[23]
port 731 nsew signal input
flabel metal2 s 36726 0 36782 800 0 FreeSans 224 90 0 0 FrameStrobe[24]
port 732 nsew signal input
flabel metal2 s 38658 0 38714 800 0 FreeSans 224 90 0 0 FrameStrobe[25]
port 733 nsew signal input
flabel metal2 s 39946 0 40002 800 0 FreeSans 224 90 0 0 FrameStrobe[26]
port 734 nsew signal input
flabel metal2 s 41878 0 41934 800 0 FreeSans 224 90 0 0 FrameStrobe[27]
port 735 nsew signal input
flabel metal2 s 43166 0 43222 800 0 FreeSans 224 90 0 0 FrameStrobe[28]
port 736 nsew signal input
flabel metal2 s 45098 0 45154 800 0 FreeSans 224 90 0 0 FrameStrobe[29]
port 737 nsew signal input
flabel metal3 s 0 19728 800 19848 0 FreeSans 480 0 0 0 FrameStrobe[2]
port 738 nsew signal input
flabel metal2 s 46386 0 46442 800 0 FreeSans 224 90 0 0 FrameStrobe[30]
port 739 nsew signal input
flabel metal2 s 47674 0 47730 800 0 FreeSans 224 90 0 0 FrameStrobe[31]
port 740 nsew signal input
flabel metal2 s 49606 0 49662 800 0 FreeSans 224 90 0 0 FrameStrobe[32]
port 741 nsew signal input
flabel metal2 s 50894 0 50950 800 0 FreeSans 224 90 0 0 FrameStrobe[33]
port 742 nsew signal input
flabel metal2 s 52826 0 52882 800 0 FreeSans 224 90 0 0 FrameStrobe[34]
port 743 nsew signal input
flabel metal2 s 54114 0 54170 800 0 FreeSans 224 90 0 0 FrameStrobe[35]
port 744 nsew signal input
flabel metal2 s 56046 0 56102 800 0 FreeSans 224 90 0 0 FrameStrobe[36]
port 745 nsew signal input
flabel metal2 s 57334 0 57390 800 0 FreeSans 224 90 0 0 FrameStrobe[37]
port 746 nsew signal input
flabel metal2 s 58622 0 58678 800 0 FreeSans 224 90 0 0 FrameStrobe[38]
port 747 nsew signal input
flabel metal2 s 60554 0 60610 800 0 FreeSans 224 90 0 0 FrameStrobe[39]
port 748 nsew signal input
flabel metal3 s 0 18368 800 18488 0 FreeSans 480 0 0 0 FrameStrobe[3]
port 749 nsew signal input
flabel metal2 s 74078 0 74134 800 0 FreeSans 224 90 0 0 FrameStrobe[40]
port 750 nsew signal input
flabel metal2 s 75366 0 75422 800 0 FreeSans 224 90 0 0 FrameStrobe[41]
port 751 nsew signal input
flabel metal2 s 76654 0 76710 800 0 FreeSans 224 90 0 0 FrameStrobe[42]
port 752 nsew signal input
flabel metal2 s 78586 0 78642 800 0 FreeSans 224 90 0 0 FrameStrobe[43]
port 753 nsew signal input
flabel metal2 s 79874 0 79930 800 0 FreeSans 224 90 0 0 FrameStrobe[44]
port 754 nsew signal input
flabel metal2 s 81162 0 81218 800 0 FreeSans 224 90 0 0 FrameStrobe[45]
port 755 nsew signal input
flabel metal2 s 82450 0 82506 800 0 FreeSans 224 90 0 0 FrameStrobe[46]
port 756 nsew signal input
flabel metal2 s 84382 0 84438 800 0 FreeSans 224 90 0 0 FrameStrobe[47]
port 757 nsew signal input
flabel metal2 s 85670 0 85726 800 0 FreeSans 224 90 0 0 FrameStrobe[48]
port 758 nsew signal input
flabel metal2 s 86958 0 87014 800 0 FreeSans 224 90 0 0 FrameStrobe[49]
port 759 nsew signal input
flabel metal3 s 0 17688 800 17808 0 FreeSans 480 0 0 0 FrameStrobe[4]
port 760 nsew signal input
flabel metal2 s 88890 0 88946 800 0 FreeSans 224 90 0 0 FrameStrobe[50]
port 761 nsew signal input
flabel metal2 s 90178 0 90234 800 0 FreeSans 224 90 0 0 FrameStrobe[51]
port 762 nsew signal input
flabel metal2 s 91466 0 91522 800 0 FreeSans 224 90 0 0 FrameStrobe[52]
port 763 nsew signal input
flabel metal2 s 92754 0 92810 800 0 FreeSans 224 90 0 0 FrameStrobe[53]
port 764 nsew signal input
flabel metal2 s 94686 0 94742 800 0 FreeSans 224 90 0 0 FrameStrobe[54]
port 765 nsew signal input
flabel metal2 s 95974 0 96030 800 0 FreeSans 224 90 0 0 FrameStrobe[55]
port 766 nsew signal input
flabel metal2 s 97262 0 97318 800 0 FreeSans 224 90 0 0 FrameStrobe[56]
port 767 nsew signal input
flabel metal2 s 99194 0 99250 800 0 FreeSans 224 90 0 0 FrameStrobe[57]
port 768 nsew signal input
flabel metal2 s 100482 0 100538 800 0 FreeSans 224 90 0 0 FrameStrobe[58]
port 769 nsew signal input
flabel metal2 s 101770 0 101826 800 0 FreeSans 224 90 0 0 FrameStrobe[59]
port 770 nsew signal input
flabel metal3 s 0 25848 800 25968 0 FreeSans 480 0 0 0 FrameStrobe[5]
port 771 nsew signal input
flabel metal2 s 106922 0 106978 800 0 FreeSans 224 90 0 0 FrameStrobe[60]
port 772 nsew signal input
flabel metal2 s 109498 0 109554 800 0 FreeSans 224 90 0 0 FrameStrobe[61]
port 773 nsew signal input
flabel metal2 s 111430 0 111486 800 0 FreeSans 224 90 0 0 FrameStrobe[62]
port 774 nsew signal input
flabel metal2 s 114006 0 114062 800 0 FreeSans 224 90 0 0 FrameStrobe[63]
port 775 nsew signal input
flabel metal2 s 115938 0 115994 800 0 FreeSans 224 90 0 0 FrameStrobe[64]
port 776 nsew signal input
flabel metal2 s 118514 0 118570 800 0 FreeSans 224 90 0 0 FrameStrobe[65]
port 777 nsew signal input
flabel metal2 s 120446 0 120502 800 0 FreeSans 224 90 0 0 FrameStrobe[66]
port 778 nsew signal input
flabel metal2 s 123022 0 123078 800 0 FreeSans 224 90 0 0 FrameStrobe[67]
port 779 nsew signal input
flabel metal2 s 125598 0 125654 800 0 FreeSans 224 90 0 0 FrameStrobe[68]
port 780 nsew signal input
flabel metal2 s 127530 0 127586 800 0 FreeSans 224 90 0 0 FrameStrobe[69]
port 781 nsew signal input
flabel metal3 s 0 23128 800 23248 0 FreeSans 480 0 0 0 FrameStrobe[6]
port 782 nsew signal input
flabel metal2 s 130106 0 130162 800 0 FreeSans 224 90 0 0 FrameStrobe[70]
port 783 nsew signal input
flabel metal2 s 132038 0 132094 800 0 FreeSans 224 90 0 0 FrameStrobe[71]
port 784 nsew signal input
flabel metal2 s 134614 0 134670 800 0 FreeSans 224 90 0 0 FrameStrobe[72]
port 785 nsew signal input
flabel metal2 s 136546 0 136602 800 0 FreeSans 224 90 0 0 FrameStrobe[73]
port 786 nsew signal input
flabel metal2 s 139122 0 139178 800 0 FreeSans 224 90 0 0 FrameStrobe[74]
port 787 nsew signal input
flabel metal2 s 141698 0 141754 800 0 FreeSans 224 90 0 0 FrameStrobe[75]
port 788 nsew signal input
flabel metal2 s 143630 0 143686 800 0 FreeSans 224 90 0 0 FrameStrobe[76]
port 789 nsew signal input
flabel metal2 s 146206 0 146262 800 0 FreeSans 224 90 0 0 FrameStrobe[77]
port 790 nsew signal input
flabel metal2 s 148138 0 148194 800 0 FreeSans 224 90 0 0 FrameStrobe[78]
port 791 nsew signal input
flabel metal2 s 150714 0 150770 800 0 FreeSans 224 90 0 0 FrameStrobe[79]
port 792 nsew signal input
flabel metal3 s 0 30608 800 30728 0 FreeSans 480 0 0 0 FrameStrobe[7]
port 793 nsew signal input
flabel metal2 s 177762 0 177818 800 0 FreeSans 224 90 0 0 FrameStrobe[80]
port 794 nsew signal input
flabel metal2 s 178406 0 178462 800 0 FreeSans 224 90 0 0 FrameStrobe[81]
port 795 nsew signal input
flabel metal2 s 179050 0 179106 800 0 FreeSans 224 90 0 0 FrameStrobe[82]
port 796 nsew signal input
flabel metal2 s 180338 0 180394 800 0 FreeSans 224 90 0 0 FrameStrobe[83]
port 797 nsew signal input
flabel metal2 s 180982 0 181038 800 0 FreeSans 224 90 0 0 FrameStrobe[84]
port 798 nsew signal input
flabel metal2 s 181626 0 181682 800 0 FreeSans 224 90 0 0 FrameStrobe[85]
port 799 nsew signal input
flabel metal2 s 182270 0 182326 800 0 FreeSans 224 90 0 0 FrameStrobe[86]
port 800 nsew signal input
flabel metal2 s 182914 0 182970 800 0 FreeSans 224 90 0 0 FrameStrobe[87]
port 801 nsew signal input
flabel metal2 s 183558 0 183614 800 0 FreeSans 224 90 0 0 FrameStrobe[88]
port 802 nsew signal input
flabel metal2 s 184202 0 184258 800 0 FreeSans 224 90 0 0 FrameStrobe[89]
port 803 nsew signal input
flabel metal3 s 0 27208 800 27328 0 FreeSans 480 0 0 0 FrameStrobe[8]
port 804 nsew signal input
flabel metal2 s 185490 0 185546 800 0 FreeSans 224 90 0 0 FrameStrobe[90]
port 805 nsew signal input
flabel metal2 s 186134 0 186190 800 0 FreeSans 224 90 0 0 FrameStrobe[91]
port 806 nsew signal input
flabel metal2 s 186778 0 186834 800 0 FreeSans 224 90 0 0 FrameStrobe[92]
port 807 nsew signal input
flabel metal2 s 187422 0 187478 800 0 FreeSans 224 90 0 0 FrameStrobe[93]
port 808 nsew signal input
flabel metal2 s 188066 0 188122 800 0 FreeSans 224 90 0 0 FrameStrobe[94]
port 809 nsew signal input
flabel metal2 s 188710 0 188766 800 0 FreeSans 224 90 0 0 FrameStrobe[95]
port 810 nsew signal input
flabel metal2 s 189354 0 189410 800 0 FreeSans 224 90 0 0 FrameStrobe[96]
port 811 nsew signal input
flabel metal2 s 190642 0 190698 800 0 FreeSans 224 90 0 0 FrameStrobe[97]
port 812 nsew signal input
flabel metal2 s 191286 0 191342 800 0 FreeSans 224 90 0 0 FrameStrobe[98]
port 813 nsew signal input
flabel metal2 s 191930 0 191986 800 0 FreeSans 224 90 0 0 FrameStrobe[99]
port 814 nsew signal input
flabel metal3 s 0 23808 800 23928 0 FreeSans 480 0 0 0 FrameStrobe[9]
port 815 nsew signal input
flabel metal3 s 0 292408 800 292528 0 FreeSans 480 0 0 0 Tile_X0Y10_A_I_top
port 816 nsew signal output
flabel metal3 s 0 291048 800 291168 0 FreeSans 480 0 0 0 Tile_X0Y10_A_O_top
port 817 nsew signal input
flabel metal3 s 0 293088 800 293208 0 FreeSans 480 0 0 0 Tile_X0Y10_A_T_top
port 818 nsew signal output
flabel metal3 s 0 296488 800 296608 0 FreeSans 480 0 0 0 Tile_X0Y10_A_config_C_bit0
port 819 nsew signal output
flabel metal3 s 0 297168 800 297288 0 FreeSans 480 0 0 0 Tile_X0Y10_A_config_C_bit1
port 820 nsew signal output
flabel metal3 s 0 297848 800 297968 0 FreeSans 480 0 0 0 Tile_X0Y10_A_config_C_bit2
port 821 nsew signal output
flabel metal3 s 0 298528 800 298648 0 FreeSans 480 0 0 0 Tile_X0Y10_A_config_C_bit3
port 822 nsew signal output
flabel metal3 s 0 294448 800 294568 0 FreeSans 480 0 0 0 Tile_X0Y10_B_I_top
port 823 nsew signal output
flabel metal3 s 0 293768 800 293888 0 FreeSans 480 0 0 0 Tile_X0Y10_B_O_top
port 824 nsew signal input
flabel metal3 s 0 295128 800 295248 0 FreeSans 480 0 0 0 Tile_X0Y10_B_T_top
port 825 nsew signal output
flabel metal3 s 0 299208 800 299328 0 FreeSans 480 0 0 0 Tile_X0Y10_B_config_C_bit0
port 826 nsew signal output
flabel metal3 s 0 300568 800 300688 0 FreeSans 480 0 0 0 Tile_X0Y10_B_config_C_bit1
port 827 nsew signal output
flabel metal3 s 0 301248 800 301368 0 FreeSans 480 0 0 0 Tile_X0Y10_B_config_C_bit2
port 828 nsew signal output
flabel metal3 s 0 301928 800 302048 0 FreeSans 480 0 0 0 Tile_X0Y10_B_config_C_bit3
port 829 nsew signal output
flabel metal3 s 0 246848 800 246968 0 FreeSans 480 0 0 0 Tile_X0Y11_A_I_top
port 830 nsew signal output
flabel metal3 s 0 246168 800 246288 0 FreeSans 480 0 0 0 Tile_X0Y11_A_O_top
port 831 nsew signal input
flabel metal3 s 0 248208 800 248328 0 FreeSans 480 0 0 0 Tile_X0Y11_A_T_top
port 832 nsew signal output
flabel metal3 s 0 250928 800 251048 0 FreeSans 480 0 0 0 Tile_X0Y11_A_config_C_bit0
port 833 nsew signal output
flabel metal3 s 0 252288 800 252408 0 FreeSans 480 0 0 0 Tile_X0Y11_A_config_C_bit1
port 834 nsew signal output
flabel metal3 s 0 252968 800 253088 0 FreeSans 480 0 0 0 Tile_X0Y11_A_config_C_bit2
port 835 nsew signal output
flabel metal3 s 0 253648 800 253768 0 FreeSans 480 0 0 0 Tile_X0Y11_A_config_C_bit3
port 836 nsew signal output
flabel metal3 s 0 249568 800 249688 0 FreeSans 480 0 0 0 Tile_X0Y11_B_I_top
port 837 nsew signal output
flabel metal3 s 0 248888 800 249008 0 FreeSans 480 0 0 0 Tile_X0Y11_B_O_top
port 838 nsew signal input
flabel metal3 s 0 250248 800 250368 0 FreeSans 480 0 0 0 Tile_X0Y11_B_T_top
port 839 nsew signal output
flabel metal3 s 0 254328 800 254448 0 FreeSans 480 0 0 0 Tile_X0Y11_B_config_C_bit0
port 840 nsew signal output
flabel metal3 s 0 255008 800 255128 0 FreeSans 480 0 0 0 Tile_X0Y11_B_config_C_bit1
port 841 nsew signal output
flabel metal3 s 0 256368 800 256488 0 FreeSans 480 0 0 0 Tile_X0Y11_B_config_C_bit2
port 842 nsew signal output
flabel metal3 s 0 257048 800 257168 0 FreeSans 480 0 0 0 Tile_X0Y11_B_config_C_bit3
port 843 nsew signal output
flabel metal3 s 0 201968 800 202088 0 FreeSans 480 0 0 0 Tile_X0Y12_A_I_top
port 844 nsew signal output
flabel metal3 s 0 201288 800 201408 0 FreeSans 480 0 0 0 Tile_X0Y12_A_O_top
port 845 nsew signal input
flabel metal3 s 0 202648 800 202768 0 FreeSans 480 0 0 0 Tile_X0Y12_A_T_top
port 846 nsew signal output
flabel metal3 s 0 206048 800 206168 0 FreeSans 480 0 0 0 Tile_X0Y12_A_config_C_bit0
port 847 nsew signal output
flabel metal3 s 0 206728 800 206848 0 FreeSans 480 0 0 0 Tile_X0Y12_A_config_C_bit1
port 848 nsew signal output
flabel metal3 s 0 208088 800 208208 0 FreeSans 480 0 0 0 Tile_X0Y12_A_config_C_bit2
port 849 nsew signal output
flabel metal3 s 0 208768 800 208888 0 FreeSans 480 0 0 0 Tile_X0Y12_A_config_C_bit3
port 850 nsew signal output
flabel metal3 s 0 204688 800 204808 0 FreeSans 480 0 0 0 Tile_X0Y12_B_I_top
port 851 nsew signal output
flabel metal3 s 0 204008 800 204128 0 FreeSans 480 0 0 0 Tile_X0Y12_B_O_top
port 852 nsew signal input
flabel metal3 s 0 205368 800 205488 0 FreeSans 480 0 0 0 Tile_X0Y12_B_T_top
port 853 nsew signal output
flabel metal3 s 0 209448 800 209568 0 FreeSans 480 0 0 0 Tile_X0Y12_B_config_C_bit0
port 854 nsew signal output
flabel metal3 s 0 210128 800 210248 0 FreeSans 480 0 0 0 Tile_X0Y12_B_config_C_bit1
port 855 nsew signal output
flabel metal3 s 0 210808 800 210928 0 FreeSans 480 0 0 0 Tile_X0Y12_B_config_C_bit2
port 856 nsew signal output
flabel metal3 s 0 211488 800 211608 0 FreeSans 480 0 0 0 Tile_X0Y12_B_config_C_bit3
port 857 nsew signal output
flabel metal3 s 0 157088 800 157208 0 FreeSans 480 0 0 0 Tile_X0Y13_A_I_top
port 858 nsew signal output
flabel metal3 s 0 156408 800 156528 0 FreeSans 480 0 0 0 Tile_X0Y13_A_O_top
port 859 nsew signal input
flabel metal3 s 0 157768 800 157888 0 FreeSans 480 0 0 0 Tile_X0Y13_A_T_top
port 860 nsew signal output
flabel metal3 s 0 161168 800 161288 0 FreeSans 480 0 0 0 Tile_X0Y13_A_config_C_bit0
port 861 nsew signal output
flabel metal3 s 0 161848 800 161968 0 FreeSans 480 0 0 0 Tile_X0Y13_A_config_C_bit1
port 862 nsew signal output
flabel metal3 s 0 162528 800 162648 0 FreeSans 480 0 0 0 Tile_X0Y13_A_config_C_bit2
port 863 nsew signal output
flabel metal3 s 0 163888 800 164008 0 FreeSans 480 0 0 0 Tile_X0Y13_A_config_C_bit3
port 864 nsew signal output
flabel metal3 s 0 159808 800 159928 0 FreeSans 480 0 0 0 Tile_X0Y13_B_I_top
port 865 nsew signal output
flabel metal3 s 0 158448 800 158568 0 FreeSans 480 0 0 0 Tile_X0Y13_B_O_top
port 866 nsew signal input
flabel metal3 s 0 160488 800 160608 0 FreeSans 480 0 0 0 Tile_X0Y13_B_T_top
port 867 nsew signal output
flabel metal3 s 0 164568 800 164688 0 FreeSans 480 0 0 0 Tile_X0Y13_B_config_C_bit0
port 868 nsew signal output
flabel metal3 s 0 165248 800 165368 0 FreeSans 480 0 0 0 Tile_X0Y13_B_config_C_bit1
port 869 nsew signal output
flabel metal3 s 0 165928 800 166048 0 FreeSans 480 0 0 0 Tile_X0Y13_B_config_C_bit2
port 870 nsew signal output
flabel metal3 s 0 166608 800 166728 0 FreeSans 480 0 0 0 Tile_X0Y13_B_config_C_bit3
port 871 nsew signal output
flabel metal3 s 0 112208 800 112328 0 FreeSans 480 0 0 0 Tile_X0Y14_A_I_top
port 872 nsew signal output
flabel metal3 s 0 111528 800 111648 0 FreeSans 480 0 0 0 Tile_X0Y14_A_O_top
port 873 nsew signal input
flabel metal3 s 0 112888 800 113008 0 FreeSans 480 0 0 0 Tile_X0Y14_A_T_top
port 874 nsew signal output
flabel metal3 s 0 116288 800 116408 0 FreeSans 480 0 0 0 Tile_X0Y14_A_config_C_bit0
port 875 nsew signal output
flabel metal3 s 0 116968 800 117088 0 FreeSans 480 0 0 0 Tile_X0Y14_A_config_C_bit1
port 876 nsew signal output
flabel metal3 s 0 117648 800 117768 0 FreeSans 480 0 0 0 Tile_X0Y14_A_config_C_bit2
port 877 nsew signal output
flabel metal3 s 0 119008 800 119128 0 FreeSans 480 0 0 0 Tile_X0Y14_A_config_C_bit3
port 878 nsew signal output
flabel metal3 s 0 114928 800 115048 0 FreeSans 480 0 0 0 Tile_X0Y14_B_I_top
port 879 nsew signal output
flabel metal3 s 0 113568 800 113688 0 FreeSans 480 0 0 0 Tile_X0Y14_B_O_top
port 880 nsew signal input
flabel metal3 s 0 115608 800 115728 0 FreeSans 480 0 0 0 Tile_X0Y14_B_T_top
port 881 nsew signal output
flabel metal3 s 0 119688 800 119808 0 FreeSans 480 0 0 0 Tile_X0Y14_B_config_C_bit0
port 882 nsew signal output
flabel metal3 s 0 120368 800 120488 0 FreeSans 480 0 0 0 Tile_X0Y14_B_config_C_bit1
port 883 nsew signal output
flabel metal3 s 0 121048 800 121168 0 FreeSans 480 0 0 0 Tile_X0Y14_B_config_C_bit2
port 884 nsew signal output
flabel metal3 s 0 121728 800 121848 0 FreeSans 480 0 0 0 Tile_X0Y14_B_config_C_bit3
port 885 nsew signal output
flabel metal3 s 0 65968 800 66088 0 FreeSans 480 0 0 0 Tile_X0Y15_A_I_top
port 886 nsew signal output
flabel metal3 s 0 52368 800 52488 0 FreeSans 480 0 0 0 Tile_X0Y15_A_O_top
port 887 nsew signal input
flabel metal3 s 0 64608 800 64728 0 FreeSans 480 0 0 0 Tile_X0Y15_A_T_top
port 888 nsew signal output
flabel metal3 s 0 70728 800 70848 0 FreeSans 480 0 0 0 Tile_X0Y15_A_config_C_bit0
port 889 nsew signal output
flabel metal3 s 0 63928 800 64048 0 FreeSans 480 0 0 0 Tile_X0Y15_A_config_C_bit1
port 890 nsew signal output
flabel metal3 s 0 65288 800 65408 0 FreeSans 480 0 0 0 Tile_X0Y15_A_config_C_bit2
port 891 nsew signal output
flabel metal3 s 0 63248 800 63368 0 FreeSans 480 0 0 0 Tile_X0Y15_A_config_C_bit3
port 892 nsew signal output
flabel metal3 s 0 69368 800 69488 0 FreeSans 480 0 0 0 Tile_X0Y15_B_I_top
port 893 nsew signal output
flabel metal3 s 0 48288 800 48408 0 FreeSans 480 0 0 0 Tile_X0Y15_B_O_top
port 894 nsew signal input
flabel metal3 s 0 70048 800 70168 0 FreeSans 480 0 0 0 Tile_X0Y15_B_T_top
port 895 nsew signal output
flabel metal3 s 0 61888 800 62008 0 FreeSans 480 0 0 0 Tile_X0Y15_B_config_C_bit0
port 896 nsew signal output
flabel metal3 s 0 71408 800 71528 0 FreeSans 480 0 0 0 Tile_X0Y15_B_config_C_bit1
port 897 nsew signal output
flabel metal3 s 0 61208 800 61328 0 FreeSans 480 0 0 0 Tile_X0Y15_B_config_C_bit2
port 898 nsew signal output
flabel metal3 s 0 68008 800 68128 0 FreeSans 480 0 0 0 Tile_X0Y15_B_config_C_bit3
port 899 nsew signal output
flabel metal3 s 0 24488 800 24608 0 FreeSans 480 0 0 0 Tile_X0Y16_A_I_top
port 900 nsew signal output
flabel metal3 s 0 21768 800 21888 0 FreeSans 480 0 0 0 Tile_X0Y16_A_O_top
port 901 nsew signal input
flabel metal2 s 6458 0 6514 800 0 FreeSans 224 90 0 0 Tile_X0Y16_A_T_top
port 902 nsew signal output
flabel metal2 s 10322 0 10378 800 0 FreeSans 224 90 0 0 Tile_X0Y16_A_config_C_bit0
port 903 nsew signal output
flabel metal2 s 12254 0 12310 800 0 FreeSans 224 90 0 0 Tile_X0Y16_A_config_C_bit1
port 904 nsew signal output
flabel metal2 s 13542 0 13598 800 0 FreeSans 224 90 0 0 Tile_X0Y16_A_config_C_bit2
port 905 nsew signal output
flabel metal2 s 10966 0 11022 800 0 FreeSans 224 90 0 0 Tile_X0Y16_A_config_C_bit3
port 906 nsew signal output
flabel metal2 s 9034 0 9090 800 0 FreeSans 224 90 0 0 Tile_X0Y16_B_I_top
port 907 nsew signal output
flabel metal2 s 7746 0 7802 800 0 FreeSans 224 90 0 0 Tile_X0Y16_B_O_top
port 908 nsew signal input
flabel metal2 s 11610 0 11666 800 0 FreeSans 224 90 0 0 Tile_X0Y16_B_T_top
port 909 nsew signal output
flabel metal2 s 9678 0 9734 800 0 FreeSans 224 90 0 0 Tile_X0Y16_B_config_C_bit0
port 910 nsew signal output
flabel metal2 s 12898 0 12954 800 0 FreeSans 224 90 0 0 Tile_X0Y16_B_config_C_bit1
port 911 nsew signal output
flabel metal2 s 7102 0 7158 800 0 FreeSans 224 90 0 0 Tile_X0Y16_B_config_C_bit2
port 912 nsew signal output
flabel metal2 s 8390 0 8446 800 0 FreeSans 224 90 0 0 Tile_X0Y16_B_config_C_bit3
port 913 nsew signal output
flabel metal3 s 0 697008 800 697128 0 FreeSans 480 0 0 0 Tile_X0Y1_A_I_top
port 914 nsew signal output
flabel metal3 s 0 696328 800 696448 0 FreeSans 480 0 0 0 Tile_X0Y1_A_O_top
port 915 nsew signal input
flabel metal3 s 0 697688 800 697808 0 FreeSans 480 0 0 0 Tile_X0Y1_A_T_top
port 916 nsew signal output
flabel metal3 s 0 701088 800 701208 0 FreeSans 480 0 0 0 Tile_X0Y1_A_config_C_bit0
port 917 nsew signal output
flabel metal3 s 0 701768 800 701888 0 FreeSans 480 0 0 0 Tile_X0Y1_A_config_C_bit1
port 918 nsew signal output
flabel metal3 s 0 703128 800 703248 0 FreeSans 480 0 0 0 Tile_X0Y1_A_config_C_bit2
port 919 nsew signal output
flabel metal3 s 0 703808 800 703928 0 FreeSans 480 0 0 0 Tile_X0Y1_A_config_C_bit3
port 920 nsew signal output
flabel metal3 s 0 699728 800 699848 0 FreeSans 480 0 0 0 Tile_X0Y1_B_I_top
port 921 nsew signal output
flabel metal3 s 0 699048 800 699168 0 FreeSans 480 0 0 0 Tile_X0Y1_B_O_top
port 922 nsew signal input
flabel metal3 s 0 700408 800 700528 0 FreeSans 480 0 0 0 Tile_X0Y1_B_T_top
port 923 nsew signal output
flabel metal3 s 0 704488 800 704608 0 FreeSans 480 0 0 0 Tile_X0Y1_B_config_C_bit0
port 924 nsew signal output
flabel metal3 s 0 705168 800 705288 0 FreeSans 480 0 0 0 Tile_X0Y1_B_config_C_bit1
port 925 nsew signal output
flabel metal3 s 0 705848 800 705968 0 FreeSans 480 0 0 0 Tile_X0Y1_B_config_C_bit2
port 926 nsew signal output
flabel metal3 s 0 707208 800 707328 0 FreeSans 480 0 0 0 Tile_X0Y1_B_config_C_bit3
port 927 nsew signal output
flabel metal3 s 0 652128 800 652248 0 FreeSans 480 0 0 0 Tile_X0Y2_A_I_top
port 928 nsew signal output
flabel metal3 s 0 651448 800 651568 0 FreeSans 480 0 0 0 Tile_X0Y2_A_O_top
port 929 nsew signal input
flabel metal3 s 0 652808 800 652928 0 FreeSans 480 0 0 0 Tile_X0Y2_A_T_top
port 930 nsew signal output
flabel metal3 s 0 656208 800 656328 0 FreeSans 480 0 0 0 Tile_X0Y2_A_config_C_bit0
port 931 nsew signal output
flabel metal3 s 0 656888 800 657008 0 FreeSans 480 0 0 0 Tile_X0Y2_A_config_C_bit1
port 932 nsew signal output
flabel metal3 s 0 657568 800 657688 0 FreeSans 480 0 0 0 Tile_X0Y2_A_config_C_bit2
port 933 nsew signal output
flabel metal3 s 0 658928 800 659048 0 FreeSans 480 0 0 0 Tile_X0Y2_A_config_C_bit3
port 934 nsew signal output
flabel metal3 s 0 654848 800 654968 0 FreeSans 480 0 0 0 Tile_X0Y2_B_I_top
port 935 nsew signal output
flabel metal3 s 0 653488 800 653608 0 FreeSans 480 0 0 0 Tile_X0Y2_B_O_top
port 936 nsew signal input
flabel metal3 s 0 655528 800 655648 0 FreeSans 480 0 0 0 Tile_X0Y2_B_T_top
port 937 nsew signal output
flabel metal3 s 0 659608 800 659728 0 FreeSans 480 0 0 0 Tile_X0Y2_B_config_C_bit0
port 938 nsew signal output
flabel metal3 s 0 660288 800 660408 0 FreeSans 480 0 0 0 Tile_X0Y2_B_config_C_bit1
port 939 nsew signal output
flabel metal3 s 0 660968 800 661088 0 FreeSans 480 0 0 0 Tile_X0Y2_B_config_C_bit2
port 940 nsew signal output
flabel metal3 s 0 661648 800 661768 0 FreeSans 480 0 0 0 Tile_X0Y2_B_config_C_bit3
port 941 nsew signal output
flabel metal3 s 0 607248 800 607368 0 FreeSans 480 0 0 0 Tile_X0Y3_A_I_top
port 942 nsew signal output
flabel metal3 s 0 606568 800 606688 0 FreeSans 480 0 0 0 Tile_X0Y3_A_O_top
port 943 nsew signal input
flabel metal3 s 0 607928 800 608048 0 FreeSans 480 0 0 0 Tile_X0Y3_A_T_top
port 944 nsew signal output
flabel metal3 s 0 611328 800 611448 0 FreeSans 480 0 0 0 Tile_X0Y3_A_config_C_bit0
port 945 nsew signal output
flabel metal3 s 0 612008 800 612128 0 FreeSans 480 0 0 0 Tile_X0Y3_A_config_C_bit1
port 946 nsew signal output
flabel metal3 s 0 612688 800 612808 0 FreeSans 480 0 0 0 Tile_X0Y3_A_config_C_bit2
port 947 nsew signal output
flabel metal3 s 0 613368 800 613488 0 FreeSans 480 0 0 0 Tile_X0Y3_A_config_C_bit3
port 948 nsew signal output
flabel metal3 s 0 609288 800 609408 0 FreeSans 480 0 0 0 Tile_X0Y3_B_I_top
port 949 nsew signal output
flabel metal3 s 0 608608 800 608728 0 FreeSans 480 0 0 0 Tile_X0Y3_B_O_top
port 950 nsew signal input
flabel metal3 s 0 610648 800 610768 0 FreeSans 480 0 0 0 Tile_X0Y3_B_T_top
port 951 nsew signal output
flabel metal3 s 0 614728 800 614848 0 FreeSans 480 0 0 0 Tile_X0Y3_B_config_C_bit0
port 952 nsew signal output
flabel metal3 s 0 615408 800 615528 0 FreeSans 480 0 0 0 Tile_X0Y3_B_config_C_bit1
port 953 nsew signal output
flabel metal3 s 0 616088 800 616208 0 FreeSans 480 0 0 0 Tile_X0Y3_B_config_C_bit2
port 954 nsew signal output
flabel metal3 s 0 616768 800 616888 0 FreeSans 480 0 0 0 Tile_X0Y3_B_config_C_bit3
port 955 nsew signal output
flabel metal3 s 0 562368 800 562488 0 FreeSans 480 0 0 0 Tile_X0Y4_A_I_top
port 956 nsew signal output
flabel metal3 s 0 561008 800 561128 0 FreeSans 480 0 0 0 Tile_X0Y4_A_O_top
port 957 nsew signal input
flabel metal3 s 0 563048 800 563168 0 FreeSans 480 0 0 0 Tile_X0Y4_A_T_top
port 958 nsew signal output
flabel metal3 s 0 566448 800 566568 0 FreeSans 480 0 0 0 Tile_X0Y4_A_config_C_bit0
port 959 nsew signal output
flabel metal3 s 0 567128 800 567248 0 FreeSans 480 0 0 0 Tile_X0Y4_A_config_C_bit1
port 960 nsew signal output
flabel metal3 s 0 567808 800 567928 0 FreeSans 480 0 0 0 Tile_X0Y4_A_config_C_bit2
port 961 nsew signal output
flabel metal3 s 0 568488 800 568608 0 FreeSans 480 0 0 0 Tile_X0Y4_A_config_C_bit3
port 962 nsew signal output
flabel metal3 s 0 564408 800 564528 0 FreeSans 480 0 0 0 Tile_X0Y4_B_I_top
port 963 nsew signal output
flabel metal3 s 0 563728 800 563848 0 FreeSans 480 0 0 0 Tile_X0Y4_B_O_top
port 964 nsew signal input
flabel metal3 s 0 565088 800 565208 0 FreeSans 480 0 0 0 Tile_X0Y4_B_T_top
port 965 nsew signal output
flabel metal3 s 0 569168 800 569288 0 FreeSans 480 0 0 0 Tile_X0Y4_B_config_C_bit0
port 966 nsew signal output
flabel metal3 s 0 570528 800 570648 0 FreeSans 480 0 0 0 Tile_X0Y4_B_config_C_bit1
port 967 nsew signal output
flabel metal3 s 0 571208 800 571328 0 FreeSans 480 0 0 0 Tile_X0Y4_B_config_C_bit2
port 968 nsew signal output
flabel metal3 s 0 571888 800 572008 0 FreeSans 480 0 0 0 Tile_X0Y4_B_config_C_bit3
port 969 nsew signal output
flabel metal3 s 0 517488 800 517608 0 FreeSans 480 0 0 0 Tile_X0Y5_A_I_top
port 970 nsew signal output
flabel metal3 s 0 516128 800 516248 0 FreeSans 480 0 0 0 Tile_X0Y5_A_O_top
port 971 nsew signal input
flabel metal3 s 0 518168 800 518288 0 FreeSans 480 0 0 0 Tile_X0Y5_A_T_top
port 972 nsew signal output
flabel metal3 s 0 521568 800 521688 0 FreeSans 480 0 0 0 Tile_X0Y5_A_config_C_bit0
port 973 nsew signal output
flabel metal3 s 0 522248 800 522368 0 FreeSans 480 0 0 0 Tile_X0Y5_A_config_C_bit1
port 974 nsew signal output
flabel metal3 s 0 522928 800 523048 0 FreeSans 480 0 0 0 Tile_X0Y5_A_config_C_bit2
port 975 nsew signal output
flabel metal3 s 0 523608 800 523728 0 FreeSans 480 0 0 0 Tile_X0Y5_A_config_C_bit3
port 976 nsew signal output
flabel metal3 s 0 519528 800 519648 0 FreeSans 480 0 0 0 Tile_X0Y5_B_I_top
port 977 nsew signal output
flabel metal3 s 0 518848 800 518968 0 FreeSans 480 0 0 0 Tile_X0Y5_B_O_top
port 978 nsew signal input
flabel metal3 s 0 520208 800 520328 0 FreeSans 480 0 0 0 Tile_X0Y5_B_T_top
port 979 nsew signal output
flabel metal3 s 0 524288 800 524408 0 FreeSans 480 0 0 0 Tile_X0Y5_B_config_C_bit0
port 980 nsew signal output
flabel metal3 s 0 525648 800 525768 0 FreeSans 480 0 0 0 Tile_X0Y5_B_config_C_bit1
port 981 nsew signal output
flabel metal3 s 0 526328 800 526448 0 FreeSans 480 0 0 0 Tile_X0Y5_B_config_C_bit2
port 982 nsew signal output
flabel metal3 s 0 527008 800 527128 0 FreeSans 480 0 0 0 Tile_X0Y5_B_config_C_bit3
port 983 nsew signal output
flabel metal3 s 0 471928 800 472048 0 FreeSans 480 0 0 0 Tile_X0Y6_A_I_top
port 984 nsew signal output
flabel metal3 s 0 471248 800 471368 0 FreeSans 480 0 0 0 Tile_X0Y6_A_O_top
port 985 nsew signal input
flabel metal3 s 0 473288 800 473408 0 FreeSans 480 0 0 0 Tile_X0Y6_A_T_top
port 986 nsew signal output
flabel metal3 s 0 476008 800 476128 0 FreeSans 480 0 0 0 Tile_X0Y6_A_config_C_bit0
port 987 nsew signal output
flabel metal3 s 0 477368 800 477488 0 FreeSans 480 0 0 0 Tile_X0Y6_A_config_C_bit1
port 988 nsew signal output
flabel metal3 s 0 478048 800 478168 0 FreeSans 480 0 0 0 Tile_X0Y6_A_config_C_bit2
port 989 nsew signal output
flabel metal3 s 0 478728 800 478848 0 FreeSans 480 0 0 0 Tile_X0Y6_A_config_C_bit3
port 990 nsew signal output
flabel metal3 s 0 474648 800 474768 0 FreeSans 480 0 0 0 Tile_X0Y6_B_I_top
port 991 nsew signal output
flabel metal3 s 0 473968 800 474088 0 FreeSans 480 0 0 0 Tile_X0Y6_B_O_top
port 992 nsew signal input
flabel metal3 s 0 475328 800 475448 0 FreeSans 480 0 0 0 Tile_X0Y6_B_T_top
port 993 nsew signal output
flabel metal3 s 0 479408 800 479528 0 FreeSans 480 0 0 0 Tile_X0Y6_B_config_C_bit0
port 994 nsew signal output
flabel metal3 s 0 480088 800 480208 0 FreeSans 480 0 0 0 Tile_X0Y6_B_config_C_bit1
port 995 nsew signal output
flabel metal3 s 0 481448 800 481568 0 FreeSans 480 0 0 0 Tile_X0Y6_B_config_C_bit2
port 996 nsew signal output
flabel metal3 s 0 482128 800 482248 0 FreeSans 480 0 0 0 Tile_X0Y6_B_config_C_bit3
port 997 nsew signal output
flabel metal3 s 0 427048 800 427168 0 FreeSans 480 0 0 0 Tile_X0Y7_A_I_top
port 998 nsew signal output
flabel metal3 s 0 426368 800 426488 0 FreeSans 480 0 0 0 Tile_X0Y7_A_O_top
port 999 nsew signal input
flabel metal3 s 0 427728 800 427848 0 FreeSans 480 0 0 0 Tile_X0Y7_A_T_top
port 1000 nsew signal output
flabel metal3 s 0 431128 800 431248 0 FreeSans 480 0 0 0 Tile_X0Y7_A_config_C_bit0
port 1001 nsew signal output
flabel metal3 s 0 431808 800 431928 0 FreeSans 480 0 0 0 Tile_X0Y7_A_config_C_bit1
port 1002 nsew signal output
flabel metal3 s 0 433168 800 433288 0 FreeSans 480 0 0 0 Tile_X0Y7_A_config_C_bit2
port 1003 nsew signal output
flabel metal3 s 0 433848 800 433968 0 FreeSans 480 0 0 0 Tile_X0Y7_A_config_C_bit3
port 1004 nsew signal output
flabel metal3 s 0 429768 800 429888 0 FreeSans 480 0 0 0 Tile_X0Y7_B_I_top
port 1005 nsew signal output
flabel metal3 s 0 429088 800 429208 0 FreeSans 480 0 0 0 Tile_X0Y7_B_O_top
port 1006 nsew signal input
flabel metal3 s 0 430448 800 430568 0 FreeSans 480 0 0 0 Tile_X0Y7_B_T_top
port 1007 nsew signal output
flabel metal3 s 0 434528 800 434648 0 FreeSans 480 0 0 0 Tile_X0Y7_B_config_C_bit0
port 1008 nsew signal output
flabel metal3 s 0 435208 800 435328 0 FreeSans 480 0 0 0 Tile_X0Y7_B_config_C_bit1
port 1009 nsew signal output
flabel metal3 s 0 435888 800 436008 0 FreeSans 480 0 0 0 Tile_X0Y7_B_config_C_bit2
port 1010 nsew signal output
flabel metal3 s 0 437248 800 437368 0 FreeSans 480 0 0 0 Tile_X0Y7_B_config_C_bit3
port 1011 nsew signal output
flabel metal3 s 0 382168 800 382288 0 FreeSans 480 0 0 0 Tile_X0Y8_A_I_top
port 1012 nsew signal output
flabel metal3 s 0 381488 800 381608 0 FreeSans 480 0 0 0 Tile_X0Y8_A_O_top
port 1013 nsew signal input
flabel metal3 s 0 382848 800 382968 0 FreeSans 480 0 0 0 Tile_X0Y8_A_T_top
port 1014 nsew signal output
flabel metal3 s 0 386248 800 386368 0 FreeSans 480 0 0 0 Tile_X0Y8_A_config_C_bit0
port 1015 nsew signal output
flabel metal3 s 0 386928 800 387048 0 FreeSans 480 0 0 0 Tile_X0Y8_A_config_C_bit1
port 1016 nsew signal output
flabel metal3 s 0 387608 800 387728 0 FreeSans 480 0 0 0 Tile_X0Y8_A_config_C_bit2
port 1017 nsew signal output
flabel metal3 s 0 388968 800 389088 0 FreeSans 480 0 0 0 Tile_X0Y8_A_config_C_bit3
port 1018 nsew signal output
flabel metal3 s 0 384888 800 385008 0 FreeSans 480 0 0 0 Tile_X0Y8_B_I_top
port 1019 nsew signal output
flabel metal3 s 0 383528 800 383648 0 FreeSans 480 0 0 0 Tile_X0Y8_B_O_top
port 1020 nsew signal input
flabel metal3 s 0 385568 800 385688 0 FreeSans 480 0 0 0 Tile_X0Y8_B_T_top
port 1021 nsew signal output
flabel metal3 s 0 389648 800 389768 0 FreeSans 480 0 0 0 Tile_X0Y8_B_config_C_bit0
port 1022 nsew signal output
flabel metal3 s 0 390328 800 390448 0 FreeSans 480 0 0 0 Tile_X0Y8_B_config_C_bit1
port 1023 nsew signal output
flabel metal3 s 0 391008 800 391128 0 FreeSans 480 0 0 0 Tile_X0Y8_B_config_C_bit2
port 1024 nsew signal output
flabel metal3 s 0 391688 800 391808 0 FreeSans 480 0 0 0 Tile_X0Y8_B_config_C_bit3
port 1025 nsew signal output
flabel metal3 s 0 337288 800 337408 0 FreeSans 480 0 0 0 Tile_X0Y9_A_I_top
port 1026 nsew signal output
flabel metal3 s 0 336608 800 336728 0 FreeSans 480 0 0 0 Tile_X0Y9_A_O_top
port 1027 nsew signal input
flabel metal3 s 0 337968 800 338088 0 FreeSans 480 0 0 0 Tile_X0Y9_A_T_top
port 1028 nsew signal output
flabel metal3 s 0 341368 800 341488 0 FreeSans 480 0 0 0 Tile_X0Y9_A_config_C_bit0
port 1029 nsew signal output
flabel metal3 s 0 342048 800 342168 0 FreeSans 480 0 0 0 Tile_X0Y9_A_config_C_bit1
port 1030 nsew signal output
flabel metal3 s 0 342728 800 342848 0 FreeSans 480 0 0 0 Tile_X0Y9_A_config_C_bit2
port 1031 nsew signal output
flabel metal3 s 0 343408 800 343528 0 FreeSans 480 0 0 0 Tile_X0Y9_A_config_C_bit3
port 1032 nsew signal output
flabel metal3 s 0 339328 800 339448 0 FreeSans 480 0 0 0 Tile_X0Y9_B_I_top
port 1033 nsew signal output
flabel metal3 s 0 338648 800 338768 0 FreeSans 480 0 0 0 Tile_X0Y9_B_O_top
port 1034 nsew signal input
flabel metal3 s 0 340688 800 340808 0 FreeSans 480 0 0 0 Tile_X0Y9_B_T_top
port 1035 nsew signal output
flabel metal3 s 0 344768 800 344888 0 FreeSans 480 0 0 0 Tile_X0Y9_B_config_C_bit0
port 1036 nsew signal output
flabel metal3 s 0 345448 800 345568 0 FreeSans 480 0 0 0 Tile_X0Y9_B_config_C_bit1
port 1037 nsew signal output
flabel metal3 s 0 346128 800 346248 0 FreeSans 480 0 0 0 Tile_X0Y9_B_config_C_bit2
port 1038 nsew signal output
flabel metal3 s 0 346808 800 346928 0 FreeSans 480 0 0 0 Tile_X0Y9_B_config_C_bit3
port 1039 nsew signal output
flabel metal2 s 405094 755700 405150 756500 0 FreeSans 224 90 0 0 Tile_X10Y0_A_I_top
port 1040 nsew signal output
flabel metal2 s 403806 755700 403862 756500 0 FreeSans 224 90 0 0 Tile_X10Y0_A_O_top
port 1041 nsew signal input
flabel metal2 s 406382 755700 406438 756500 0 FreeSans 224 90 0 0 Tile_X10Y0_A_T_top
port 1042 nsew signal output
flabel metal2 s 410246 755700 410302 756500 0 FreeSans 224 90 0 0 Tile_X10Y0_A_config_C_bit0
port 1043 nsew signal output
flabel metal2 s 411534 755700 411590 756500 0 FreeSans 224 90 0 0 Tile_X10Y0_A_config_C_bit1
port 1044 nsew signal output
flabel metal2 s 412822 755700 412878 756500 0 FreeSans 224 90 0 0 Tile_X10Y0_A_config_C_bit2
port 1045 nsew signal output
flabel metal2 s 414110 755700 414166 756500 0 FreeSans 224 90 0 0 Tile_X10Y0_A_config_C_bit3
port 1046 nsew signal output
flabel metal2 s 408314 755700 408370 756500 0 FreeSans 224 90 0 0 Tile_X10Y0_B_I_top
port 1047 nsew signal output
flabel metal2 s 407026 755700 407082 756500 0 FreeSans 224 90 0 0 Tile_X10Y0_B_O_top
port 1048 nsew signal input
flabel metal2 s 409602 755700 409658 756500 0 FreeSans 224 90 0 0 Tile_X10Y0_B_T_top
port 1049 nsew signal output
flabel metal2 s 414754 755700 414810 756500 0 FreeSans 224 90 0 0 Tile_X10Y0_B_config_C_bit0
port 1050 nsew signal output
flabel metal2 s 416042 755700 416098 756500 0 FreeSans 224 90 0 0 Tile_X10Y0_B_config_C_bit1
port 1051 nsew signal output
flabel metal2 s 417330 755700 417386 756500 0 FreeSans 224 90 0 0 Tile_X10Y0_B_config_C_bit2
port 1052 nsew signal output
flabel metal2 s 417974 755700 418030 756500 0 FreeSans 224 90 0 0 Tile_X10Y0_B_config_C_bit3
port 1053 nsew signal output
flabel metal2 s 403162 0 403218 800 0 FreeSans 224 90 0 0 Tile_X10Y17_VALUE_top0
port 1054 nsew signal output
flabel metal2 s 404450 0 404506 800 0 FreeSans 224 90 0 0 Tile_X10Y17_VALUE_top1
port 1055 nsew signal output
flabel metal2 s 406382 0 406438 800 0 FreeSans 224 90 0 0 Tile_X10Y17_VALUE_top2
port 1056 nsew signal output
flabel metal2 s 407670 0 407726 800 0 FreeSans 224 90 0 0 Tile_X10Y17_VALUE_top3
port 1057 nsew signal output
flabel metal2 s 408958 0 409014 800 0 FreeSans 224 90 0 0 Tile_X10Y17_VALUE_top4
port 1058 nsew signal output
flabel metal2 s 410246 0 410302 800 0 FreeSans 224 90 0 0 Tile_X10Y17_VALUE_top5
port 1059 nsew signal output
flabel metal2 s 411534 0 411590 800 0 FreeSans 224 90 0 0 Tile_X10Y17_VALUE_top6
port 1060 nsew signal output
flabel metal2 s 412822 0 412878 800 0 FreeSans 224 90 0 0 Tile_X10Y17_VALUE_top7
port 1061 nsew signal output
flabel metal3 s 486200 286968 487000 287088 0 FreeSans 480 0 0 0 Tile_X11Y10_AD_SRAM0
port 1062 nsew signal output
flabel metal3 s 486200 317568 487000 317688 0 FreeSans 480 0 0 0 Tile_X11Y10_AD_SRAM1
port 1063 nsew signal output
flabel metal3 s 486200 295128 487000 295248 0 FreeSans 480 0 0 0 Tile_X11Y10_AD_SRAM2
port 1064 nsew signal output
flabel metal3 s 486200 318248 487000 318368 0 FreeSans 480 0 0 0 Tile_X11Y10_AD_SRAM3
port 1065 nsew signal output
flabel metal3 s 486200 294448 487000 294568 0 FreeSans 480 0 0 0 Tile_X11Y10_AD_SRAM4
port 1066 nsew signal output
flabel metal3 s 486200 293768 487000 293888 0 FreeSans 480 0 0 0 Tile_X11Y10_AD_SRAM5
port 1067 nsew signal output
flabel metal3 s 486200 318928 487000 319048 0 FreeSans 480 0 0 0 Tile_X11Y10_AD_SRAM6
port 1068 nsew signal output
flabel metal3 s 486200 293088 487000 293208 0 FreeSans 480 0 0 0 Tile_X11Y10_AD_SRAM7
port 1069 nsew signal output
flabel metal3 s 486200 319608 487000 319728 0 FreeSans 480 0 0 0 Tile_X11Y10_AD_SRAM8
port 1070 nsew signal output
flabel metal3 s 486200 292408 487000 292528 0 FreeSans 480 0 0 0 Tile_X11Y10_AD_SRAM9
port 1071 nsew signal output
flabel metal3 s 486200 291728 487000 291848 0 FreeSans 480 0 0 0 Tile_X11Y10_BEN_SRAM0
port 1072 nsew signal output
flabel metal3 s 486200 320288 487000 320408 0 FreeSans 480 0 0 0 Tile_X11Y10_BEN_SRAM1
port 1073 nsew signal output
flabel metal3 s 486200 287648 487000 287768 0 FreeSans 480 0 0 0 Tile_X11Y10_BEN_SRAM10
port 1074 nsew signal output
flabel metal3 s 486200 323008 487000 323128 0 FreeSans 480 0 0 0 Tile_X11Y10_BEN_SRAM11
port 1075 nsew signal output
flabel metal3 s 486200 323688 487000 323808 0 FreeSans 480 0 0 0 Tile_X11Y10_BEN_SRAM12
port 1076 nsew signal output
flabel metal3 s 486200 360408 487000 360528 0 FreeSans 480 0 0 0 Tile_X11Y10_BEN_SRAM13
port 1077 nsew signal output
flabel metal3 s 486200 359728 487000 359848 0 FreeSans 480 0 0 0 Tile_X11Y10_BEN_SRAM14
port 1078 nsew signal output
flabel metal3 s 486200 324368 487000 324488 0 FreeSans 480 0 0 0 Tile_X11Y10_BEN_SRAM15
port 1079 nsew signal output
flabel metal3 s 486200 359048 487000 359168 0 FreeSans 480 0 0 0 Tile_X11Y10_BEN_SRAM16
port 1080 nsew signal output
flabel metal3 s 486200 325048 487000 325168 0 FreeSans 480 0 0 0 Tile_X11Y10_BEN_SRAM17
port 1081 nsew signal output
flabel metal3 s 486200 358368 487000 358488 0 FreeSans 480 0 0 0 Tile_X11Y10_BEN_SRAM18
port 1082 nsew signal output
flabel metal3 s 486200 357688 487000 357808 0 FreeSans 480 0 0 0 Tile_X11Y10_BEN_SRAM19
port 1083 nsew signal output
flabel metal3 s 486200 291048 487000 291168 0 FreeSans 480 0 0 0 Tile_X11Y10_BEN_SRAM2
port 1084 nsew signal output
flabel metal3 s 486200 325728 487000 325848 0 FreeSans 480 0 0 0 Tile_X11Y10_BEN_SRAM20
port 1085 nsew signal output
flabel metal3 s 486200 357008 487000 357128 0 FreeSans 480 0 0 0 Tile_X11Y10_BEN_SRAM21
port 1086 nsew signal output
flabel metal3 s 486200 326408 487000 326528 0 FreeSans 480 0 0 0 Tile_X11Y10_BEN_SRAM22
port 1087 nsew signal output
flabel metal3 s 486200 356328 487000 356448 0 FreeSans 480 0 0 0 Tile_X11Y10_BEN_SRAM23
port 1088 nsew signal output
flabel metal3 s 486200 355648 487000 355768 0 FreeSans 480 0 0 0 Tile_X11Y10_BEN_SRAM24
port 1089 nsew signal output
flabel metal3 s 486200 327088 487000 327208 0 FreeSans 480 0 0 0 Tile_X11Y10_BEN_SRAM25
port 1090 nsew signal output
flabel metal3 s 486200 354968 487000 355088 0 FreeSans 480 0 0 0 Tile_X11Y10_BEN_SRAM26
port 1091 nsew signal output
flabel metal3 s 486200 327768 487000 327888 0 FreeSans 480 0 0 0 Tile_X11Y10_BEN_SRAM27
port 1092 nsew signal output
flabel metal3 s 486200 354288 487000 354408 0 FreeSans 480 0 0 0 Tile_X11Y10_BEN_SRAM28
port 1093 nsew signal output
flabel metal3 s 486200 353608 487000 353728 0 FreeSans 480 0 0 0 Tile_X11Y10_BEN_SRAM29
port 1094 nsew signal output
flabel metal3 s 486200 320968 487000 321088 0 FreeSans 480 0 0 0 Tile_X11Y10_BEN_SRAM3
port 1095 nsew signal output
flabel metal3 s 486200 328448 487000 328568 0 FreeSans 480 0 0 0 Tile_X11Y10_BEN_SRAM30
port 1096 nsew signal output
flabel metal3 s 486200 352928 487000 353048 0 FreeSans 480 0 0 0 Tile_X11Y10_BEN_SRAM31
port 1097 nsew signal output
flabel metal3 s 486200 290368 487000 290488 0 FreeSans 480 0 0 0 Tile_X11Y10_BEN_SRAM4
port 1098 nsew signal output
flabel metal3 s 486200 289688 487000 289808 0 FreeSans 480 0 0 0 Tile_X11Y10_BEN_SRAM5
port 1099 nsew signal output
flabel metal3 s 486200 321648 487000 321768 0 FreeSans 480 0 0 0 Tile_X11Y10_BEN_SRAM6
port 1100 nsew signal output
flabel metal3 s 486200 289008 487000 289128 0 FreeSans 480 0 0 0 Tile_X11Y10_BEN_SRAM7
port 1101 nsew signal output
flabel metal3 s 486200 322328 487000 322448 0 FreeSans 480 0 0 0 Tile_X11Y10_BEN_SRAM8
port 1102 nsew signal output
flabel metal3 s 486200 288328 487000 288448 0 FreeSans 480 0 0 0 Tile_X11Y10_BEN_SRAM9
port 1103 nsew signal output
flabel metal3 s 486200 329128 487000 329248 0 FreeSans 480 0 0 0 Tile_X11Y10_CLOCK_SRAM
port 1104 nsew signal output
flabel metal3 s 486200 352248 487000 352368 0 FreeSans 480 0 0 0 Tile_X11Y10_DI_SRAM0
port 1105 nsew signal output
flabel metal3 s 486200 351568 487000 351688 0 FreeSans 480 0 0 0 Tile_X11Y10_DI_SRAM1
port 1106 nsew signal output
flabel metal3 s 486200 350888 487000 351008 0 FreeSans 480 0 0 0 Tile_X11Y10_DI_SRAM10
port 1107 nsew signal output
flabel metal3 s 486200 347488 487000 347608 0 FreeSans 480 0 0 0 Tile_X11Y10_DI_SRAM11
port 1108 nsew signal output
flabel metal3 s 486200 334568 487000 334688 0 FreeSans 480 0 0 0 Tile_X11Y10_DI_SRAM12
port 1109 nsew signal output
flabel metal3 s 486200 346808 487000 346928 0 FreeSans 480 0 0 0 Tile_X11Y10_DI_SRAM13
port 1110 nsew signal output
flabel metal3 s 486200 335248 487000 335368 0 FreeSans 480 0 0 0 Tile_X11Y10_DI_SRAM14
port 1111 nsew signal output
flabel metal3 s 486200 346128 487000 346248 0 FreeSans 480 0 0 0 Tile_X11Y10_DI_SRAM15
port 1112 nsew signal output
flabel metal3 s 486200 345448 487000 345568 0 FreeSans 480 0 0 0 Tile_X11Y10_DI_SRAM16
port 1113 nsew signal output
flabel metal3 s 486200 335928 487000 336048 0 FreeSans 480 0 0 0 Tile_X11Y10_DI_SRAM17
port 1114 nsew signal output
flabel metal3 s 486200 344768 487000 344888 0 FreeSans 480 0 0 0 Tile_X11Y10_DI_SRAM18
port 1115 nsew signal output
flabel metal3 s 486200 336608 487000 336728 0 FreeSans 480 0 0 0 Tile_X11Y10_DI_SRAM19
port 1116 nsew signal output
flabel metal3 s 486200 329808 487000 329928 0 FreeSans 480 0 0 0 Tile_X11Y10_DI_SRAM2
port 1117 nsew signal output
flabel metal3 s 486200 344088 487000 344208 0 FreeSans 480 0 0 0 Tile_X11Y10_DI_SRAM20
port 1118 nsew signal output
flabel metal3 s 486200 343408 487000 343528 0 FreeSans 480 0 0 0 Tile_X11Y10_DI_SRAM21
port 1119 nsew signal output
flabel metal3 s 486200 350208 487000 350328 0 FreeSans 480 0 0 0 Tile_X11Y10_DI_SRAM22
port 1120 nsew signal output
flabel metal3 s 486200 342728 487000 342848 0 FreeSans 480 0 0 0 Tile_X11Y10_DI_SRAM23
port 1121 nsew signal output
flabel metal3 s 486200 349528 487000 349648 0 FreeSans 480 0 0 0 Tile_X11Y10_DI_SRAM24
port 1122 nsew signal output
flabel metal3 s 486200 348848 487000 348968 0 FreeSans 480 0 0 0 Tile_X11Y10_DI_SRAM25
port 1123 nsew signal output
flabel metal3 s 486200 341368 487000 341488 0 FreeSans 480 0 0 0 Tile_X11Y10_DI_SRAM26
port 1124 nsew signal output
flabel metal3 s 486200 348168 487000 348288 0 FreeSans 480 0 0 0 Tile_X11Y10_DI_SRAM27
port 1125 nsew signal output
flabel metal3 s 486200 340688 487000 340808 0 FreeSans 480 0 0 0 Tile_X11Y10_DI_SRAM28
port 1126 nsew signal output
flabel metal3 s 486200 337288 487000 337408 0 FreeSans 480 0 0 0 Tile_X11Y10_DI_SRAM29
port 1127 nsew signal output
flabel metal3 s 486200 330488 487000 330608 0 FreeSans 480 0 0 0 Tile_X11Y10_DI_SRAM3
port 1128 nsew signal output
flabel metal3 s 486200 340008 487000 340128 0 FreeSans 480 0 0 0 Tile_X11Y10_DI_SRAM30
port 1129 nsew signal output
flabel metal3 s 486200 339328 487000 339448 0 FreeSans 480 0 0 0 Tile_X11Y10_DI_SRAM31
port 1130 nsew signal output
flabel metal3 s 486200 331168 487000 331288 0 FreeSans 480 0 0 0 Tile_X11Y10_DI_SRAM4
port 1131 nsew signal output
flabel metal3 s 486200 331848 487000 331968 0 FreeSans 480 0 0 0 Tile_X11Y10_DI_SRAM5
port 1132 nsew signal output
flabel metal3 s 486200 338648 487000 338768 0 FreeSans 480 0 0 0 Tile_X11Y10_DI_SRAM6
port 1133 nsew signal output
flabel metal3 s 486200 332528 487000 332648 0 FreeSans 480 0 0 0 Tile_X11Y10_DI_SRAM7
port 1134 nsew signal output
flabel metal3 s 486200 333208 487000 333328 0 FreeSans 480 0 0 0 Tile_X11Y10_DI_SRAM8
port 1135 nsew signal output
flabel metal3 s 486200 333888 487000 334008 0 FreeSans 480 0 0 0 Tile_X11Y10_DI_SRAM9
port 1136 nsew signal output
flabel metal3 s 486200 295808 487000 295928 0 FreeSans 480 0 0 0 Tile_X11Y10_DO_SRAM0
port 1137 nsew signal input
flabel metal3 s 486200 308728 487000 308848 0 FreeSans 480 0 0 0 Tile_X11Y10_DO_SRAM1
port 1138 nsew signal input
flabel metal3 s 486200 311448 487000 311568 0 FreeSans 480 0 0 0 Tile_X11Y10_DO_SRAM10
port 1139 nsew signal input
flabel metal3 s 486200 304648 487000 304768 0 FreeSans 480 0 0 0 Tile_X11Y10_DO_SRAM11
port 1140 nsew signal input
flabel metal3 s 486200 303968 487000 304088 0 FreeSans 480 0 0 0 Tile_X11Y10_DO_SRAM12
port 1141 nsew signal input
flabel metal3 s 486200 312128 487000 312248 0 FreeSans 480 0 0 0 Tile_X11Y10_DO_SRAM13
port 1142 nsew signal input
flabel metal3 s 486200 303288 487000 303408 0 FreeSans 480 0 0 0 Tile_X11Y10_DO_SRAM14
port 1143 nsew signal input
flabel metal3 s 486200 312808 487000 312928 0 FreeSans 480 0 0 0 Tile_X11Y10_DO_SRAM15
port 1144 nsew signal input
flabel metal3 s 486200 302608 487000 302728 0 FreeSans 480 0 0 0 Tile_X11Y10_DO_SRAM16
port 1145 nsew signal input
flabel metal3 s 486200 301928 487000 302048 0 FreeSans 480 0 0 0 Tile_X11Y10_DO_SRAM17
port 1146 nsew signal input
flabel metal3 s 486200 313488 487000 313608 0 FreeSans 480 0 0 0 Tile_X11Y10_DO_SRAM18
port 1147 nsew signal input
flabel metal3 s 486200 301248 487000 301368 0 FreeSans 480 0 0 0 Tile_X11Y10_DO_SRAM19
port 1148 nsew signal input
flabel metal3 s 486200 308048 487000 308168 0 FreeSans 480 0 0 0 Tile_X11Y10_DO_SRAM2
port 1149 nsew signal input
flabel metal3 s 486200 314168 487000 314288 0 FreeSans 480 0 0 0 Tile_X11Y10_DO_SRAM20
port 1150 nsew signal input
flabel metal3 s 486200 300568 487000 300688 0 FreeSans 480 0 0 0 Tile_X11Y10_DO_SRAM21
port 1151 nsew signal input
flabel metal3 s 486200 299888 487000 300008 0 FreeSans 480 0 0 0 Tile_X11Y10_DO_SRAM22
port 1152 nsew signal input
flabel metal3 s 486200 314848 487000 314968 0 FreeSans 480 0 0 0 Tile_X11Y10_DO_SRAM23
port 1153 nsew signal input
flabel metal3 s 486200 299208 487000 299328 0 FreeSans 480 0 0 0 Tile_X11Y10_DO_SRAM24
port 1154 nsew signal input
flabel metal3 s 486200 315528 487000 315648 0 FreeSans 480 0 0 0 Tile_X11Y10_DO_SRAM25
port 1155 nsew signal input
flabel metal3 s 486200 298528 487000 298648 0 FreeSans 480 0 0 0 Tile_X11Y10_DO_SRAM26
port 1156 nsew signal input
flabel metal3 s 486200 297848 487000 297968 0 FreeSans 480 0 0 0 Tile_X11Y10_DO_SRAM27
port 1157 nsew signal input
flabel metal3 s 486200 316208 487000 316328 0 FreeSans 480 0 0 0 Tile_X11Y10_DO_SRAM28
port 1158 nsew signal input
flabel metal3 s 486200 297168 487000 297288 0 FreeSans 480 0 0 0 Tile_X11Y10_DO_SRAM29
port 1159 nsew signal input
flabel metal3 s 486200 309408 487000 309528 0 FreeSans 480 0 0 0 Tile_X11Y10_DO_SRAM3
port 1160 nsew signal input
flabel metal3 s 486200 316888 487000 317008 0 FreeSans 480 0 0 0 Tile_X11Y10_DO_SRAM30
port 1161 nsew signal input
flabel metal3 s 486200 296488 487000 296608 0 FreeSans 480 0 0 0 Tile_X11Y10_DO_SRAM31
port 1162 nsew signal input
flabel metal3 s 486200 307368 487000 307488 0 FreeSans 480 0 0 0 Tile_X11Y10_DO_SRAM4
port 1163 nsew signal input
flabel metal3 s 486200 310088 487000 310208 0 FreeSans 480 0 0 0 Tile_X11Y10_DO_SRAM5
port 1164 nsew signal input
flabel metal3 s 486200 306688 487000 306808 0 FreeSans 480 0 0 0 Tile_X11Y10_DO_SRAM6
port 1165 nsew signal input
flabel metal3 s 486200 306008 487000 306128 0 FreeSans 480 0 0 0 Tile_X11Y10_DO_SRAM7
port 1166 nsew signal input
flabel metal3 s 486200 310768 487000 310888 0 FreeSans 480 0 0 0 Tile_X11Y10_DO_SRAM8
port 1167 nsew signal input
flabel metal3 s 486200 305328 487000 305448 0 FreeSans 480 0 0 0 Tile_X11Y10_DO_SRAM9
port 1168 nsew signal input
flabel metal3 s 486200 337968 487000 338088 0 FreeSans 480 0 0 0 Tile_X11Y10_EN_SRAM
port 1169 nsew signal output
flabel metal3 s 486200 342048 487000 342168 0 FreeSans 480 0 0 0 Tile_X11Y10_R_WB_SRAM
port 1170 nsew signal output
flabel metal3 s 486200 196528 487000 196648 0 FreeSans 480 0 0 0 Tile_X11Y12_AD_SRAM0
port 1171 nsew signal output
flabel metal3 s 486200 205368 487000 205488 0 FreeSans 480 0 0 0 Tile_X11Y12_AD_SRAM1
port 1172 nsew signal output
flabel metal3 s 486200 227808 487000 227928 0 FreeSans 480 0 0 0 Tile_X11Y12_AD_SRAM2
port 1173 nsew signal output
flabel metal3 s 486200 204688 487000 204808 0 FreeSans 480 0 0 0 Tile_X11Y12_AD_SRAM3
port 1174 nsew signal output
flabel metal3 s 486200 228488 487000 228608 0 FreeSans 480 0 0 0 Tile_X11Y12_AD_SRAM4
port 1175 nsew signal output
flabel metal3 s 486200 204008 487000 204128 0 FreeSans 480 0 0 0 Tile_X11Y12_AD_SRAM5
port 1176 nsew signal output
flabel metal3 s 486200 203328 487000 203448 0 FreeSans 480 0 0 0 Tile_X11Y12_AD_SRAM6
port 1177 nsew signal output
flabel metal3 s 486200 229168 487000 229288 0 FreeSans 480 0 0 0 Tile_X11Y12_AD_SRAM7
port 1178 nsew signal output
flabel metal3 s 486200 202648 487000 202768 0 FreeSans 480 0 0 0 Tile_X11Y12_AD_SRAM8
port 1179 nsew signal output
flabel metal3 s 486200 229848 487000 229968 0 FreeSans 480 0 0 0 Tile_X11Y12_AD_SRAM9
port 1180 nsew signal output
flabel metal3 s 486200 201968 487000 202088 0 FreeSans 480 0 0 0 Tile_X11Y12_BEN_SRAM0
port 1181 nsew signal output
flabel metal3 s 486200 201288 487000 201408 0 FreeSans 480 0 0 0 Tile_X11Y12_BEN_SRAM1
port 1182 nsew signal output
flabel metal3 s 486200 232568 487000 232688 0 FreeSans 480 0 0 0 Tile_X11Y12_BEN_SRAM10
port 1183 nsew signal output
flabel metal3 s 486200 197208 487000 197328 0 FreeSans 480 0 0 0 Tile_X11Y12_BEN_SRAM11
port 1184 nsew signal output
flabel metal3 s 486200 233248 487000 233368 0 FreeSans 480 0 0 0 Tile_X11Y12_BEN_SRAM12
port 1185 nsew signal output
flabel metal3 s 486200 233928 487000 234048 0 FreeSans 480 0 0 0 Tile_X11Y12_BEN_SRAM13
port 1186 nsew signal output
flabel metal3 s 486200 269968 487000 270088 0 FreeSans 480 0 0 0 Tile_X11Y12_BEN_SRAM14
port 1187 nsew signal output
flabel metal3 s 486200 269288 487000 269408 0 FreeSans 480 0 0 0 Tile_X11Y12_BEN_SRAM15
port 1188 nsew signal output
flabel metal3 s 486200 234608 487000 234728 0 FreeSans 480 0 0 0 Tile_X11Y12_BEN_SRAM16
port 1189 nsew signal output
flabel metal3 s 486200 268608 487000 268728 0 FreeSans 480 0 0 0 Tile_X11Y12_BEN_SRAM17
port 1190 nsew signal output
flabel metal3 s 486200 235288 487000 235408 0 FreeSans 480 0 0 0 Tile_X11Y12_BEN_SRAM18
port 1191 nsew signal output
flabel metal3 s 486200 267928 487000 268048 0 FreeSans 480 0 0 0 Tile_X11Y12_BEN_SRAM19
port 1192 nsew signal output
flabel metal3 s 486200 230528 487000 230648 0 FreeSans 480 0 0 0 Tile_X11Y12_BEN_SRAM2
port 1193 nsew signal output
flabel metal3 s 486200 267248 487000 267368 0 FreeSans 480 0 0 0 Tile_X11Y12_BEN_SRAM20
port 1194 nsew signal output
flabel metal3 s 486200 235968 487000 236088 0 FreeSans 480 0 0 0 Tile_X11Y12_BEN_SRAM21
port 1195 nsew signal output
flabel metal3 s 486200 266568 487000 266688 0 FreeSans 480 0 0 0 Tile_X11Y12_BEN_SRAM22
port 1196 nsew signal output
flabel metal3 s 486200 236648 487000 236768 0 FreeSans 480 0 0 0 Tile_X11Y12_BEN_SRAM23
port 1197 nsew signal output
flabel metal3 s 486200 265888 487000 266008 0 FreeSans 480 0 0 0 Tile_X11Y12_BEN_SRAM24
port 1198 nsew signal output
flabel metal3 s 486200 265208 487000 265328 0 FreeSans 480 0 0 0 Tile_X11Y12_BEN_SRAM25
port 1199 nsew signal output
flabel metal3 s 486200 237328 487000 237448 0 FreeSans 480 0 0 0 Tile_X11Y12_BEN_SRAM26
port 1200 nsew signal output
flabel metal3 s 486200 264528 487000 264648 0 FreeSans 480 0 0 0 Tile_X11Y12_BEN_SRAM27
port 1201 nsew signal output
flabel metal3 s 486200 238008 487000 238128 0 FreeSans 480 0 0 0 Tile_X11Y12_BEN_SRAM28
port 1202 nsew signal output
flabel metal3 s 486200 263848 487000 263968 0 FreeSans 480 0 0 0 Tile_X11Y12_BEN_SRAM29
port 1203 nsew signal output
flabel metal3 s 486200 200608 487000 200728 0 FreeSans 480 0 0 0 Tile_X11Y12_BEN_SRAM3
port 1204 nsew signal output
flabel metal3 s 486200 263168 487000 263288 0 FreeSans 480 0 0 0 Tile_X11Y12_BEN_SRAM30
port 1205 nsew signal output
flabel metal3 s 486200 238688 487000 238808 0 FreeSans 480 0 0 0 Tile_X11Y12_BEN_SRAM31
port 1206 nsew signal output
flabel metal3 s 486200 231208 487000 231328 0 FreeSans 480 0 0 0 Tile_X11Y12_BEN_SRAM4
port 1207 nsew signal output
flabel metal3 s 486200 199928 487000 200048 0 FreeSans 480 0 0 0 Tile_X11Y12_BEN_SRAM5
port 1208 nsew signal output
flabel metal3 s 486200 199248 487000 199368 0 FreeSans 480 0 0 0 Tile_X11Y12_BEN_SRAM6
port 1209 nsew signal output
flabel metal3 s 486200 231888 487000 232008 0 FreeSans 480 0 0 0 Tile_X11Y12_BEN_SRAM7
port 1210 nsew signal output
flabel metal3 s 486200 198568 487000 198688 0 FreeSans 480 0 0 0 Tile_X11Y12_BEN_SRAM8
port 1211 nsew signal output
flabel metal3 s 486200 197888 487000 198008 0 FreeSans 480 0 0 0 Tile_X11Y12_BEN_SRAM9
port 1212 nsew signal output
flabel metal3 s 486200 262488 487000 262608 0 FreeSans 480 0 0 0 Tile_X11Y12_CLOCK_SRAM
port 1213 nsew signal output
flabel metal3 s 486200 239368 487000 239488 0 FreeSans 480 0 0 0 Tile_X11Y12_DI_SRAM0
port 1214 nsew signal output
flabel metal3 s 486200 261808 487000 261928 0 FreeSans 480 0 0 0 Tile_X11Y12_DI_SRAM1
port 1215 nsew signal output
flabel metal3 s 486200 261128 487000 261248 0 FreeSans 480 0 0 0 Tile_X11Y12_DI_SRAM10
port 1216 nsew signal output
flabel metal3 s 486200 257728 487000 257848 0 FreeSans 480 0 0 0 Tile_X11Y12_DI_SRAM11
port 1217 nsew signal output
flabel metal3 s 486200 257048 487000 257168 0 FreeSans 480 0 0 0 Tile_X11Y12_DI_SRAM12
port 1218 nsew signal output
flabel metal3 s 486200 244808 487000 244928 0 FreeSans 480 0 0 0 Tile_X11Y12_DI_SRAM13
port 1219 nsew signal output
flabel metal3 s 486200 256368 487000 256488 0 FreeSans 480 0 0 0 Tile_X11Y12_DI_SRAM14
port 1220 nsew signal output
flabel metal3 s 486200 245488 487000 245608 0 FreeSans 480 0 0 0 Tile_X11Y12_DI_SRAM15
port 1221 nsew signal output
flabel metal3 s 486200 260448 487000 260568 0 FreeSans 480 0 0 0 Tile_X11Y12_DI_SRAM16
port 1222 nsew signal output
flabel metal3 s 486200 255008 487000 255128 0 FreeSans 480 0 0 0 Tile_X11Y12_DI_SRAM17
port 1223 nsew signal output
flabel metal3 s 486200 259768 487000 259888 0 FreeSans 480 0 0 0 Tile_X11Y12_DI_SRAM18
port 1224 nsew signal output
flabel metal3 s 486200 254328 487000 254448 0 FreeSans 480 0 0 0 Tile_X11Y12_DI_SRAM19
port 1225 nsew signal output
flabel metal3 s 486200 240048 487000 240168 0 FreeSans 480 0 0 0 Tile_X11Y12_DI_SRAM2
port 1226 nsew signal output
flabel metal3 s 486200 246168 487000 246288 0 FreeSans 480 0 0 0 Tile_X11Y12_DI_SRAM20
port 1227 nsew signal output
flabel metal3 s 486200 253648 487000 253768 0 FreeSans 480 0 0 0 Tile_X11Y12_DI_SRAM21
port 1228 nsew signal output
flabel metal3 s 486200 252968 487000 253088 0 FreeSans 480 0 0 0 Tile_X11Y12_DI_SRAM22
port 1229 nsew signal output
flabel metal3 s 486200 246848 487000 246968 0 FreeSans 480 0 0 0 Tile_X11Y12_DI_SRAM23
port 1230 nsew signal output
flabel metal3 s 486200 259088 487000 259208 0 FreeSans 480 0 0 0 Tile_X11Y12_DI_SRAM24
port 1231 nsew signal output
flabel metal3 s 486200 247528 487000 247648 0 FreeSans 480 0 0 0 Tile_X11Y12_DI_SRAM25
port 1232 nsew signal output
flabel metal3 s 486200 258408 487000 258528 0 FreeSans 480 0 0 0 Tile_X11Y12_DI_SRAM26
port 1233 nsew signal output
flabel metal3 s 486200 250928 487000 251048 0 FreeSans 480 0 0 0 Tile_X11Y12_DI_SRAM27
port 1234 nsew signal output
flabel metal3 s 486200 248208 487000 248328 0 FreeSans 480 0 0 0 Tile_X11Y12_DI_SRAM28
port 1235 nsew signal output
flabel metal3 s 486200 250248 487000 250368 0 FreeSans 480 0 0 0 Tile_X11Y12_DI_SRAM29
port 1236 nsew signal output
flabel metal3 s 486200 240728 487000 240848 0 FreeSans 480 0 0 0 Tile_X11Y12_DI_SRAM3
port 1237 nsew signal output
flabel metal3 s 486200 248888 487000 249008 0 FreeSans 480 0 0 0 Tile_X11Y12_DI_SRAM30
port 1238 nsew signal output
flabel metal3 s 486200 249568 487000 249688 0 FreeSans 480 0 0 0 Tile_X11Y12_DI_SRAM31
port 1239 nsew signal output
flabel metal3 s 486200 241408 487000 241528 0 FreeSans 480 0 0 0 Tile_X11Y12_DI_SRAM4
port 1240 nsew signal output
flabel metal3 s 486200 242088 487000 242208 0 FreeSans 480 0 0 0 Tile_X11Y12_DI_SRAM5
port 1241 nsew signal output
flabel metal3 s 486200 242768 487000 242888 0 FreeSans 480 0 0 0 Tile_X11Y12_DI_SRAM6
port 1242 nsew signal output
flabel metal3 s 486200 243448 487000 243568 0 FreeSans 480 0 0 0 Tile_X11Y12_DI_SRAM7
port 1243 nsew signal output
flabel metal3 s 486200 244128 487000 244248 0 FreeSans 480 0 0 0 Tile_X11Y12_DI_SRAM8
port 1244 nsew signal output
flabel metal3 s 486200 255688 487000 255808 0 FreeSans 480 0 0 0 Tile_X11Y12_DI_SRAM9
port 1245 nsew signal output
flabel metal3 s 486200 206048 487000 206168 0 FreeSans 480 0 0 0 Tile_X11Y12_DO_SRAM0
port 1246 nsew signal input
flabel metal3 s 486200 218968 487000 219088 0 FreeSans 480 0 0 0 Tile_X11Y12_DO_SRAM1
port 1247 nsew signal input
flabel metal3 s 486200 214888 487000 215008 0 FreeSans 480 0 0 0 Tile_X11Y12_DO_SRAM10
port 1248 nsew signal input
flabel metal3 s 486200 221688 487000 221808 0 FreeSans 480 0 0 0 Tile_X11Y12_DO_SRAM11
port 1249 nsew signal input
flabel metal3 s 486200 214208 487000 214328 0 FreeSans 480 0 0 0 Tile_X11Y12_DO_SRAM12
port 1250 nsew signal input
flabel metal3 s 486200 213528 487000 213648 0 FreeSans 480 0 0 0 Tile_X11Y12_DO_SRAM13
port 1251 nsew signal input
flabel metal3 s 486200 222368 487000 222488 0 FreeSans 480 0 0 0 Tile_X11Y12_DO_SRAM14
port 1252 nsew signal input
flabel metal3 s 486200 212848 487000 212968 0 FreeSans 480 0 0 0 Tile_X11Y12_DO_SRAM15
port 1253 nsew signal input
flabel metal3 s 486200 223048 487000 223168 0 FreeSans 480 0 0 0 Tile_X11Y12_DO_SRAM16
port 1254 nsew signal input
flabel metal3 s 486200 212168 487000 212288 0 FreeSans 480 0 0 0 Tile_X11Y12_DO_SRAM17
port 1255 nsew signal input
flabel metal3 s 486200 211488 487000 211608 0 FreeSans 480 0 0 0 Tile_X11Y12_DO_SRAM18
port 1256 nsew signal input
flabel metal3 s 486200 223728 487000 223848 0 FreeSans 480 0 0 0 Tile_X11Y12_DO_SRAM19
port 1257 nsew signal input
flabel metal3 s 486200 218288 487000 218408 0 FreeSans 480 0 0 0 Tile_X11Y12_DO_SRAM2
port 1258 nsew signal input
flabel metal3 s 486200 210808 487000 210928 0 FreeSans 480 0 0 0 Tile_X11Y12_DO_SRAM20
port 1259 nsew signal input
flabel metal3 s 486200 224408 487000 224528 0 FreeSans 480 0 0 0 Tile_X11Y12_DO_SRAM21
port 1260 nsew signal input
flabel metal3 s 486200 210128 487000 210248 0 FreeSans 480 0 0 0 Tile_X11Y12_DO_SRAM22
port 1261 nsew signal input
flabel metal3 s 486200 209448 487000 209568 0 FreeSans 480 0 0 0 Tile_X11Y12_DO_SRAM23
port 1262 nsew signal input
flabel metal3 s 486200 225088 487000 225208 0 FreeSans 480 0 0 0 Tile_X11Y12_DO_SRAM24
port 1263 nsew signal input
flabel metal3 s 486200 208768 487000 208888 0 FreeSans 480 0 0 0 Tile_X11Y12_DO_SRAM25
port 1264 nsew signal input
flabel metal3 s 486200 225768 487000 225888 0 FreeSans 480 0 0 0 Tile_X11Y12_DO_SRAM26
port 1265 nsew signal input
flabel metal3 s 486200 208088 487000 208208 0 FreeSans 480 0 0 0 Tile_X11Y12_DO_SRAM27
port 1266 nsew signal input
flabel metal3 s 486200 207408 487000 207528 0 FreeSans 480 0 0 0 Tile_X11Y12_DO_SRAM28
port 1267 nsew signal input
flabel metal3 s 486200 226448 487000 226568 0 FreeSans 480 0 0 0 Tile_X11Y12_DO_SRAM29
port 1268 nsew signal input
flabel metal3 s 486200 217608 487000 217728 0 FreeSans 480 0 0 0 Tile_X11Y12_DO_SRAM3
port 1269 nsew signal input
flabel metal3 s 486200 206728 487000 206848 0 FreeSans 480 0 0 0 Tile_X11Y12_DO_SRAM30
port 1270 nsew signal input
flabel metal3 s 486200 227128 487000 227248 0 FreeSans 480 0 0 0 Tile_X11Y12_DO_SRAM31
port 1271 nsew signal input
flabel metal3 s 486200 219648 487000 219768 0 FreeSans 480 0 0 0 Tile_X11Y12_DO_SRAM4
port 1272 nsew signal input
flabel metal3 s 486200 216928 487000 217048 0 FreeSans 480 0 0 0 Tile_X11Y12_DO_SRAM5
port 1273 nsew signal input
flabel metal3 s 486200 220328 487000 220448 0 FreeSans 480 0 0 0 Tile_X11Y12_DO_SRAM6
port 1274 nsew signal input
flabel metal3 s 486200 216248 487000 216368 0 FreeSans 480 0 0 0 Tile_X11Y12_DO_SRAM7
port 1275 nsew signal input
flabel metal3 s 486200 215568 487000 215688 0 FreeSans 480 0 0 0 Tile_X11Y12_DO_SRAM8
port 1276 nsew signal input
flabel metal3 s 486200 221008 487000 221128 0 FreeSans 480 0 0 0 Tile_X11Y12_DO_SRAM9
port 1277 nsew signal input
flabel metal3 s 486200 252288 487000 252408 0 FreeSans 480 0 0 0 Tile_X11Y12_EN_SRAM
port 1278 nsew signal output
flabel metal3 s 486200 251608 487000 251728 0 FreeSans 480 0 0 0 Tile_X11Y12_R_WB_SRAM
port 1279 nsew signal output
flabel metal3 s 486200 192448 487000 192568 0 FreeSans 480 0 0 0 Tile_X11Y14_AD_SRAM0
port 1280 nsew signal output
flabel metal3 s 486200 189048 487000 189168 0 FreeSans 480 0 0 0 Tile_X11Y14_AD_SRAM1
port 1281 nsew signal output
flabel metal3 s 486200 138048 487000 138168 0 FreeSans 480 0 0 0 Tile_X11Y14_AD_SRAM2
port 1282 nsew signal output
flabel metal3 s 486200 188368 487000 188488 0 FreeSans 480 0 0 0 Tile_X11Y14_AD_SRAM3
port 1283 nsew signal output
flabel metal3 s 486200 148928 487000 149048 0 FreeSans 480 0 0 0 Tile_X11Y14_AD_SRAM4
port 1284 nsew signal output
flabel metal3 s 486200 187688 487000 187808 0 FreeSans 480 0 0 0 Tile_X11Y14_AD_SRAM5
port 1285 nsew signal output
flabel metal3 s 486200 187008 487000 187128 0 FreeSans 480 0 0 0 Tile_X11Y14_AD_SRAM6
port 1286 nsew signal output
flabel metal3 s 486200 139408 487000 139528 0 FreeSans 480 0 0 0 Tile_X11Y14_AD_SRAM7
port 1287 nsew signal output
flabel metal3 s 486200 186328 487000 186448 0 FreeSans 480 0 0 0 Tile_X11Y14_AD_SRAM8
port 1288 nsew signal output
flabel metal3 s 486200 140088 487000 140208 0 FreeSans 480 0 0 0 Tile_X11Y14_AD_SRAM9
port 1289 nsew signal output
flabel metal3 s 486200 185648 487000 185768 0 FreeSans 480 0 0 0 Tile_X11Y14_BEN_SRAM0
port 1290 nsew signal output
flabel metal3 s 486200 184968 487000 185088 0 FreeSans 480 0 0 0 Tile_X11Y14_BEN_SRAM1
port 1291 nsew signal output
flabel metal3 s 486200 184288 487000 184408 0 FreeSans 480 0 0 0 Tile_X11Y14_BEN_SRAM10
port 1292 nsew signal output
flabel metal3 s 486200 180888 487000 181008 0 FreeSans 480 0 0 0 Tile_X11Y14_BEN_SRAM11
port 1293 nsew signal output
flabel metal3 s 486200 145528 487000 145648 0 FreeSans 480 0 0 0 Tile_X11Y14_BEN_SRAM12
port 1294 nsew signal output
flabel metal3 s 486200 180208 487000 180328 0 FreeSans 480 0 0 0 Tile_X11Y14_BEN_SRAM13
port 1295 nsew signal output
flabel metal3 s 486200 146208 487000 146328 0 FreeSans 480 0 0 0 Tile_X11Y14_BEN_SRAM14
port 1296 nsew signal output
flabel metal3 s 486200 179528 487000 179648 0 FreeSans 480 0 0 0 Tile_X11Y14_BEN_SRAM15
port 1297 nsew signal output
flabel metal3 s 486200 191768 487000 191888 0 FreeSans 480 0 0 0 Tile_X11Y14_BEN_SRAM16
port 1298 nsew signal output
flabel metal3 s 486200 144848 487000 144968 0 FreeSans 480 0 0 0 Tile_X11Y14_BEN_SRAM17
port 1299 nsew signal output
flabel metal3 s 486200 178168 487000 178288 0 FreeSans 480 0 0 0 Tile_X11Y14_BEN_SRAM18
port 1300 nsew signal output
flabel metal3 s 486200 191088 487000 191208 0 FreeSans 480 0 0 0 Tile_X11Y14_BEN_SRAM19
port 1301 nsew signal output
flabel metal3 s 486200 140768 487000 140888 0 FreeSans 480 0 0 0 Tile_X11Y14_BEN_SRAM2
port 1302 nsew signal output
flabel metal3 s 486200 177488 487000 177608 0 FreeSans 480 0 0 0 Tile_X11Y14_BEN_SRAM20
port 1303 nsew signal output
flabel metal3 s 486200 176808 487000 176928 0 FreeSans 480 0 0 0 Tile_X11Y14_BEN_SRAM21
port 1304 nsew signal output
flabel metal3 s 486200 190408 487000 190528 0 FreeSans 480 0 0 0 Tile_X11Y14_BEN_SRAM22
port 1305 nsew signal output
flabel metal3 s 486200 176128 487000 176248 0 FreeSans 480 0 0 0 Tile_X11Y14_BEN_SRAM23
port 1306 nsew signal output
flabel metal3 s 486200 148248 487000 148368 0 FreeSans 480 0 0 0 Tile_X11Y14_BEN_SRAM24
port 1307 nsew signal output
flabel metal3 s 486200 189728 487000 189848 0 FreeSans 480 0 0 0 Tile_X11Y14_BEN_SRAM25
port 1308 nsew signal output
flabel metal3 s 486200 174768 487000 174888 0 FreeSans 480 0 0 0 Tile_X11Y14_BEN_SRAM26
port 1309 nsew signal output
flabel metal3 s 486200 147568 487000 147688 0 FreeSans 480 0 0 0 Tile_X11Y14_BEN_SRAM27
port 1310 nsew signal output
flabel metal3 s 486200 174088 487000 174208 0 FreeSans 480 0 0 0 Tile_X11Y14_BEN_SRAM28
port 1311 nsew signal output
flabel metal3 s 486200 149608 487000 149728 0 FreeSans 480 0 0 0 Tile_X11Y14_BEN_SRAM29
port 1312 nsew signal output
flabel metal3 s 486200 142128 487000 142248 0 FreeSans 480 0 0 0 Tile_X11Y14_BEN_SRAM3
port 1313 nsew signal output
flabel metal3 s 486200 173408 487000 173528 0 FreeSans 480 0 0 0 Tile_X11Y14_BEN_SRAM30
port 1314 nsew signal output
flabel metal3 s 486200 172728 487000 172848 0 FreeSans 480 0 0 0 Tile_X11Y14_BEN_SRAM31
port 1315 nsew signal output
flabel metal3 s 486200 141448 487000 141568 0 FreeSans 480 0 0 0 Tile_X11Y14_BEN_SRAM4
port 1316 nsew signal output
flabel metal3 s 486200 143488 487000 143608 0 FreeSans 480 0 0 0 Tile_X11Y14_BEN_SRAM5
port 1317 nsew signal output
flabel metal3 s 486200 142808 487000 142928 0 FreeSans 480 0 0 0 Tile_X11Y14_BEN_SRAM6
port 1318 nsew signal output
flabel metal3 s 486200 153008 487000 153128 0 FreeSans 480 0 0 0 Tile_X11Y14_BEN_SRAM7
port 1319 nsew signal output
flabel metal3 s 486200 150288 487000 150408 0 FreeSans 480 0 0 0 Tile_X11Y14_BEN_SRAM8
port 1320 nsew signal output
flabel metal3 s 486200 144168 487000 144288 0 FreeSans 480 0 0 0 Tile_X11Y14_BEN_SRAM9
port 1321 nsew signal output
flabel metal3 s 486200 161168 487000 161288 0 FreeSans 480 0 0 0 Tile_X11Y14_CLOCK_SRAM
port 1322 nsew signal output
flabel metal3 s 486200 172048 487000 172168 0 FreeSans 480 0 0 0 Tile_X11Y14_DI_SRAM0
port 1323 nsew signal output
flabel metal3 s 486200 153688 487000 153808 0 FreeSans 480 0 0 0 Tile_X11Y14_DI_SRAM1
port 1324 nsew signal output
flabel metal3 s 486200 171368 487000 171488 0 FreeSans 480 0 0 0 Tile_X11Y14_DI_SRAM10
port 1325 nsew signal output
flabel metal3 s 486200 154368 487000 154488 0 FreeSans 480 0 0 0 Tile_X11Y14_DI_SRAM11
port 1326 nsew signal output
flabel metal3 s 486200 167288 487000 167408 0 FreeSans 480 0 0 0 Tile_X11Y14_DI_SRAM12
port 1327 nsew signal output
flabel metal3 s 486200 166608 487000 166728 0 FreeSans 480 0 0 0 Tile_X11Y14_DI_SRAM13
port 1328 nsew signal output
flabel metal3 s 486200 159128 487000 159248 0 FreeSans 480 0 0 0 Tile_X11Y14_DI_SRAM14
port 1329 nsew signal output
flabel metal3 s 486200 165928 487000 166048 0 FreeSans 480 0 0 0 Tile_X11Y14_DI_SRAM15
port 1330 nsew signal output
flabel metal3 s 486200 155048 487000 155168 0 FreeSans 480 0 0 0 Tile_X11Y14_DI_SRAM16
port 1331 nsew signal output
flabel metal3 s 486200 165248 487000 165368 0 FreeSans 480 0 0 0 Tile_X11Y14_DI_SRAM17
port 1332 nsew signal output
flabel metal3 s 486200 183608 487000 183728 0 FreeSans 480 0 0 0 Tile_X11Y14_DI_SRAM18
port 1333 nsew signal output
flabel metal3 s 486200 155728 487000 155848 0 FreeSans 480 0 0 0 Tile_X11Y14_DI_SRAM19
port 1334 nsew signal output
flabel metal3 s 486200 158448 487000 158568 0 FreeSans 480 0 0 0 Tile_X11Y14_DI_SRAM2
port 1335 nsew signal output
flabel metal3 s 486200 182928 487000 183048 0 FreeSans 480 0 0 0 Tile_X11Y14_DI_SRAM20
port 1336 nsew signal output
flabel metal3 s 486200 167968 487000 168088 0 FreeSans 480 0 0 0 Tile_X11Y14_DI_SRAM21
port 1337 nsew signal output
flabel metal3 s 486200 163208 487000 163328 0 FreeSans 480 0 0 0 Tile_X11Y14_DI_SRAM22
port 1338 nsew signal output
flabel metal3 s 486200 162528 487000 162648 0 FreeSans 480 0 0 0 Tile_X11Y14_DI_SRAM23
port 1339 nsew signal output
flabel metal3 s 486200 170008 487000 170128 0 FreeSans 480 0 0 0 Tile_X11Y14_DI_SRAM24
port 1340 nsew signal output
flabel metal3 s 486200 161848 487000 161968 0 FreeSans 480 0 0 0 Tile_X11Y14_DI_SRAM25
port 1341 nsew signal output
flabel metal3 s 486200 156408 487000 156528 0 FreeSans 480 0 0 0 Tile_X11Y14_DI_SRAM26
port 1342 nsew signal output
flabel metal3 s 486200 168648 487000 168768 0 FreeSans 480 0 0 0 Tile_X11Y14_DI_SRAM27
port 1343 nsew signal output
flabel metal3 s 486200 160488 487000 160608 0 FreeSans 480 0 0 0 Tile_X11Y14_DI_SRAM28
port 1344 nsew signal output
flabel metal3 s 486200 157088 487000 157208 0 FreeSans 480 0 0 0 Tile_X11Y14_DI_SRAM29
port 1345 nsew signal output
flabel metal3 s 486200 182248 487000 182368 0 FreeSans 480 0 0 0 Tile_X11Y14_DI_SRAM3
port 1346 nsew signal output
flabel metal3 s 486200 159808 487000 159928 0 FreeSans 480 0 0 0 Tile_X11Y14_DI_SRAM30
port 1347 nsew signal output
flabel metal3 s 486200 157768 487000 157888 0 FreeSans 480 0 0 0 Tile_X11Y14_DI_SRAM31
port 1348 nsew signal output
flabel metal3 s 486200 170688 487000 170808 0 FreeSans 480 0 0 0 Tile_X11Y14_DI_SRAM4
port 1349 nsew signal output
flabel metal3 s 486200 150968 487000 151088 0 FreeSans 480 0 0 0 Tile_X11Y14_DI_SRAM5
port 1350 nsew signal output
flabel metal3 s 486200 151648 487000 151768 0 FreeSans 480 0 0 0 Tile_X11Y14_DI_SRAM6
port 1351 nsew signal output
flabel metal3 s 486200 152328 487000 152448 0 FreeSans 480 0 0 0 Tile_X11Y14_DI_SRAM7
port 1352 nsew signal output
flabel metal3 s 486200 181568 487000 181688 0 FreeSans 480 0 0 0 Tile_X11Y14_DI_SRAM8
port 1353 nsew signal output
flabel metal3 s 486200 163888 487000 164008 0 FreeSans 480 0 0 0 Tile_X11Y14_DI_SRAM9
port 1354 nsew signal output
flabel metal3 s 486200 119008 487000 119128 0 FreeSans 480 0 0 0 Tile_X11Y14_DO_SRAM0
port 1355 nsew signal input
flabel metal3 s 486200 128528 487000 128648 0 FreeSans 480 0 0 0 Tile_X11Y14_DO_SRAM1
port 1356 nsew signal input
flabel metal3 s 486200 131248 487000 131368 0 FreeSans 480 0 0 0 Tile_X11Y14_DO_SRAM10
port 1357 nsew signal input
flabel metal3 s 486200 124448 487000 124568 0 FreeSans 480 0 0 0 Tile_X11Y14_DO_SRAM11
port 1358 nsew signal input
flabel metal3 s 486200 131928 487000 132048 0 FreeSans 480 0 0 0 Tile_X11Y14_DO_SRAM12
port 1359 nsew signal input
flabel metal3 s 486200 123768 487000 123888 0 FreeSans 480 0 0 0 Tile_X11Y14_DO_SRAM13
port 1360 nsew signal input
flabel metal3 s 486200 123088 487000 123208 0 FreeSans 480 0 0 0 Tile_X11Y14_DO_SRAM14
port 1361 nsew signal input
flabel metal3 s 486200 132608 487000 132728 0 FreeSans 480 0 0 0 Tile_X11Y14_DO_SRAM15
port 1362 nsew signal input
flabel metal3 s 486200 122408 487000 122528 0 FreeSans 480 0 0 0 Tile_X11Y14_DO_SRAM16
port 1363 nsew signal input
flabel metal3 s 486200 133288 487000 133408 0 FreeSans 480 0 0 0 Tile_X11Y14_DO_SRAM17
port 1364 nsew signal input
flabel metal3 s 486200 121728 487000 121848 0 FreeSans 480 0 0 0 Tile_X11Y14_DO_SRAM18
port 1365 nsew signal input
flabel metal3 s 486200 121048 487000 121168 0 FreeSans 480 0 0 0 Tile_X11Y14_DO_SRAM19
port 1366 nsew signal input
flabel metal3 s 486200 129208 487000 129328 0 FreeSans 480 0 0 0 Tile_X11Y14_DO_SRAM2
port 1367 nsew signal input
flabel metal3 s 486200 133968 487000 134088 0 FreeSans 480 0 0 0 Tile_X11Y14_DO_SRAM20
port 1368 nsew signal input
flabel metal3 s 486200 120368 487000 120488 0 FreeSans 480 0 0 0 Tile_X11Y14_DO_SRAM21
port 1369 nsew signal input
flabel metal3 s 486200 134648 487000 134768 0 FreeSans 480 0 0 0 Tile_X11Y14_DO_SRAM22
port 1370 nsew signal input
flabel metal3 s 486200 119688 487000 119808 0 FreeSans 480 0 0 0 Tile_X11Y14_DO_SRAM23
port 1371 nsew signal input
flabel metal3 s 486200 135328 487000 135448 0 FreeSans 480 0 0 0 Tile_X11Y14_DO_SRAM24
port 1372 nsew signal input
flabel metal3 s 486200 136008 487000 136128 0 FreeSans 480 0 0 0 Tile_X11Y14_DO_SRAM25
port 1373 nsew signal input
flabel metal3 s 486200 146888 487000 147008 0 FreeSans 480 0 0 0 Tile_X11Y14_DO_SRAM26
port 1374 nsew signal input
flabel metal3 s 486200 178848 487000 178968 0 FreeSans 480 0 0 0 Tile_X11Y14_DO_SRAM27
port 1375 nsew signal input
flabel metal3 s 486200 137368 487000 137488 0 FreeSans 480 0 0 0 Tile_X11Y14_DO_SRAM28
port 1376 nsew signal input
flabel metal3 s 486200 136688 487000 136808 0 FreeSans 480 0 0 0 Tile_X11Y14_DO_SRAM29
port 1377 nsew signal input
flabel metal3 s 486200 127848 487000 127968 0 FreeSans 480 0 0 0 Tile_X11Y14_DO_SRAM3
port 1378 nsew signal input
flabel metal3 s 486200 138728 487000 138848 0 FreeSans 480 0 0 0 Tile_X11Y14_DO_SRAM30
port 1379 nsew signal input
flabel metal3 s 486200 175448 487000 175568 0 FreeSans 480 0 0 0 Tile_X11Y14_DO_SRAM31
port 1380 nsew signal input
flabel metal3 s 486200 127168 487000 127288 0 FreeSans 480 0 0 0 Tile_X11Y14_DO_SRAM4
port 1381 nsew signal input
flabel metal3 s 486200 129888 487000 130008 0 FreeSans 480 0 0 0 Tile_X11Y14_DO_SRAM5
port 1382 nsew signal input
flabel metal3 s 486200 126488 487000 126608 0 FreeSans 480 0 0 0 Tile_X11Y14_DO_SRAM6
port 1383 nsew signal input
flabel metal3 s 486200 130568 487000 130688 0 FreeSans 480 0 0 0 Tile_X11Y14_DO_SRAM7
port 1384 nsew signal input
flabel metal3 s 486200 125808 487000 125928 0 FreeSans 480 0 0 0 Tile_X11Y14_DO_SRAM8
port 1385 nsew signal input
flabel metal3 s 486200 125128 487000 125248 0 FreeSans 480 0 0 0 Tile_X11Y14_DO_SRAM9
port 1386 nsew signal input
flabel metal3 s 486200 169328 487000 169448 0 FreeSans 480 0 0 0 Tile_X11Y14_EN_SRAM
port 1387 nsew signal output
flabel metal3 s 486200 164568 487000 164688 0 FreeSans 480 0 0 0 Tile_X11Y14_R_WB_SRAM
port 1388 nsew signal output
flabel metal3 s 486200 17008 487000 17128 0 FreeSans 480 0 0 0 Tile_X11Y16_AD_SRAM0
port 1389 nsew signal output
flabel metal3 s 486200 47608 487000 47728 0 FreeSans 480 0 0 0 Tile_X11Y16_AD_SRAM1
port 1390 nsew signal output
flabel metal3 s 486200 25168 487000 25288 0 FreeSans 480 0 0 0 Tile_X11Y16_AD_SRAM2
port 1391 nsew signal output
flabel metal3 s 486200 24488 487000 24608 0 FreeSans 480 0 0 0 Tile_X11Y16_AD_SRAM3
port 1392 nsew signal output
flabel metal3 s 486200 48288 487000 48408 0 FreeSans 480 0 0 0 Tile_X11Y16_AD_SRAM4
port 1393 nsew signal output
flabel metal3 s 486200 23808 487000 23928 0 FreeSans 480 0 0 0 Tile_X11Y16_AD_SRAM5
port 1394 nsew signal output
flabel metal3 s 486200 48968 487000 49088 0 FreeSans 480 0 0 0 Tile_X11Y16_AD_SRAM6
port 1395 nsew signal output
flabel metal3 s 486200 23128 487000 23248 0 FreeSans 480 0 0 0 Tile_X11Y16_AD_SRAM7
port 1396 nsew signal output
flabel metal3 s 486200 22448 487000 22568 0 FreeSans 480 0 0 0 Tile_X11Y16_AD_SRAM8
port 1397 nsew signal output
flabel metal3 s 486200 49648 487000 49768 0 FreeSans 480 0 0 0 Tile_X11Y16_AD_SRAM9
port 1398 nsew signal output
flabel metal3 s 486200 21768 487000 21888 0 FreeSans 480 0 0 0 Tile_X11Y16_BEN_SRAM0
port 1399 nsew signal output
flabel metal3 s 486200 50328 487000 50448 0 FreeSans 480 0 0 0 Tile_X11Y16_BEN_SRAM1
port 1400 nsew signal output
flabel metal3 s 486200 17688 487000 17808 0 FreeSans 480 0 0 0 Tile_X11Y16_BEN_SRAM10
port 1401 nsew signal output
flabel metal3 s 486200 53048 487000 53168 0 FreeSans 480 0 0 0 Tile_X11Y16_BEN_SRAM11
port 1402 nsew signal output
flabel metal3 s 486200 90448 487000 90568 0 FreeSans 480 0 0 0 Tile_X11Y16_BEN_SRAM12
port 1403 nsew signal output
flabel metal3 s 486200 53728 487000 53848 0 FreeSans 480 0 0 0 Tile_X11Y16_BEN_SRAM13
port 1404 nsew signal output
flabel metal3 s 486200 89768 487000 89888 0 FreeSans 480 0 0 0 Tile_X11Y16_BEN_SRAM14
port 1405 nsew signal output
flabel metal3 s 486200 54408 487000 54528 0 FreeSans 480 0 0 0 Tile_X11Y16_BEN_SRAM15
port 1406 nsew signal output
flabel metal3 s 486200 89088 487000 89208 0 FreeSans 480 0 0 0 Tile_X11Y16_BEN_SRAM16
port 1407 nsew signal output
flabel metal3 s 486200 88408 487000 88528 0 FreeSans 480 0 0 0 Tile_X11Y16_BEN_SRAM17
port 1408 nsew signal output
flabel metal3 s 486200 55088 487000 55208 0 FreeSans 480 0 0 0 Tile_X11Y16_BEN_SRAM18
port 1409 nsew signal output
flabel metal3 s 486200 87728 487000 87848 0 FreeSans 480 0 0 0 Tile_X11Y16_BEN_SRAM19
port 1410 nsew signal output
flabel metal3 s 486200 21088 487000 21208 0 FreeSans 480 0 0 0 Tile_X11Y16_BEN_SRAM2
port 1411 nsew signal output
flabel metal3 s 486200 55768 487000 55888 0 FreeSans 480 0 0 0 Tile_X11Y16_BEN_SRAM20
port 1412 nsew signal output
flabel metal3 s 486200 87048 487000 87168 0 FreeSans 480 0 0 0 Tile_X11Y16_BEN_SRAM21
port 1413 nsew signal output
flabel metal3 s 486200 86368 487000 86488 0 FreeSans 480 0 0 0 Tile_X11Y16_BEN_SRAM22
port 1414 nsew signal output
flabel metal3 s 486200 56448 487000 56568 0 FreeSans 480 0 0 0 Tile_X11Y16_BEN_SRAM23
port 1415 nsew signal output
flabel metal3 s 486200 85688 487000 85808 0 FreeSans 480 0 0 0 Tile_X11Y16_BEN_SRAM24
port 1416 nsew signal output
flabel metal3 s 486200 57128 487000 57248 0 FreeSans 480 0 0 0 Tile_X11Y16_BEN_SRAM25
port 1417 nsew signal output
flabel metal3 s 486200 85008 487000 85128 0 FreeSans 480 0 0 0 Tile_X11Y16_BEN_SRAM26
port 1418 nsew signal output
flabel metal3 s 486200 84328 487000 84448 0 FreeSans 480 0 0 0 Tile_X11Y16_BEN_SRAM27
port 1419 nsew signal output
flabel metal3 s 486200 57808 487000 57928 0 FreeSans 480 0 0 0 Tile_X11Y16_BEN_SRAM28
port 1420 nsew signal output
flabel metal3 s 486200 83648 487000 83768 0 FreeSans 480 0 0 0 Tile_X11Y16_BEN_SRAM29
port 1421 nsew signal output
flabel metal3 s 486200 20408 487000 20528 0 FreeSans 480 0 0 0 Tile_X11Y16_BEN_SRAM3
port 1422 nsew signal output
flabel metal3 s 486200 58488 487000 58608 0 FreeSans 480 0 0 0 Tile_X11Y16_BEN_SRAM30
port 1423 nsew signal output
flabel metal3 s 486200 82968 487000 83088 0 FreeSans 480 0 0 0 Tile_X11Y16_BEN_SRAM31
port 1424 nsew signal output
flabel metal3 s 486200 51008 487000 51128 0 FreeSans 480 0 0 0 Tile_X11Y16_BEN_SRAM4
port 1425 nsew signal output
flabel metal3 s 486200 19728 487000 19848 0 FreeSans 480 0 0 0 Tile_X11Y16_BEN_SRAM5
port 1426 nsew signal output
flabel metal3 s 486200 51688 487000 51808 0 FreeSans 480 0 0 0 Tile_X11Y16_BEN_SRAM6
port 1427 nsew signal output
flabel metal3 s 486200 19048 487000 19168 0 FreeSans 480 0 0 0 Tile_X11Y16_BEN_SRAM7
port 1428 nsew signal output
flabel metal3 s 486200 18368 487000 18488 0 FreeSans 480 0 0 0 Tile_X11Y16_BEN_SRAM8
port 1429 nsew signal output
flabel metal3 s 486200 52368 487000 52488 0 FreeSans 480 0 0 0 Tile_X11Y16_BEN_SRAM9
port 1430 nsew signal output
flabel metal3 s 486200 82288 487000 82408 0 FreeSans 480 0 0 0 Tile_X11Y16_CLOCK_SRAM
port 1431 nsew signal output
flabel metal3 s 486200 59168 487000 59288 0 FreeSans 480 0 0 0 Tile_X11Y16_DI_SRAM0
port 1432 nsew signal output
flabel metal3 s 486200 81608 487000 81728 0 FreeSans 480 0 0 0 Tile_X11Y16_DI_SRAM1
port 1433 nsew signal output
flabel metal3 s 486200 80928 487000 81048 0 FreeSans 480 0 0 0 Tile_X11Y16_DI_SRAM10
port 1434 nsew signal output
flabel metal3 s 486200 80248 487000 80368 0 FreeSans 480 0 0 0 Tile_X11Y16_DI_SRAM11
port 1435 nsew signal output
flabel metal3 s 486200 65288 487000 65408 0 FreeSans 480 0 0 0 Tile_X11Y16_DI_SRAM12
port 1436 nsew signal output
flabel metal3 s 486200 76848 487000 76968 0 FreeSans 480 0 0 0 Tile_X11Y16_DI_SRAM13
port 1437 nsew signal output
flabel metal3 s 486200 76168 487000 76288 0 FreeSans 480 0 0 0 Tile_X11Y16_DI_SRAM14
port 1438 nsew signal output
flabel metal3 s 486200 63928 487000 64048 0 FreeSans 480 0 0 0 Tile_X11Y16_DI_SRAM15
port 1439 nsew signal output
flabel metal3 s 486200 75488 487000 75608 0 FreeSans 480 0 0 0 Tile_X11Y16_DI_SRAM16
port 1440 nsew signal output
flabel metal3 s 486200 65968 487000 66088 0 FreeSans 480 0 0 0 Tile_X11Y16_DI_SRAM17
port 1441 nsew signal output
flabel metal3 s 486200 79568 487000 79688 0 FreeSans 480 0 0 0 Tile_X11Y16_DI_SRAM18
port 1442 nsew signal output
flabel metal3 s 486200 74128 487000 74248 0 FreeSans 480 0 0 0 Tile_X11Y16_DI_SRAM19
port 1443 nsew signal output
flabel metal3 s 486200 59848 487000 59968 0 FreeSans 480 0 0 0 Tile_X11Y16_DI_SRAM2
port 1444 nsew signal output
flabel metal3 s 486200 67328 487000 67448 0 FreeSans 480 0 0 0 Tile_X11Y16_DI_SRAM20
port 1445 nsew signal output
flabel metal3 s 486200 73448 487000 73568 0 FreeSans 480 0 0 0 Tile_X11Y16_DI_SRAM21
port 1446 nsew signal output
flabel metal3 s 486200 68008 487000 68128 0 FreeSans 480 0 0 0 Tile_X11Y16_DI_SRAM22
port 1447 nsew signal output
flabel metal3 s 486200 78888 487000 79008 0 FreeSans 480 0 0 0 Tile_X11Y16_DI_SRAM23
port 1448 nsew signal output
flabel metal3 s 486200 72088 487000 72208 0 FreeSans 480 0 0 0 Tile_X11Y16_DI_SRAM24
port 1449 nsew signal output
flabel metal3 s 486200 66648 487000 66768 0 FreeSans 480 0 0 0 Tile_X11Y16_DI_SRAM25
port 1450 nsew signal output
flabel metal3 s 486200 71408 487000 71528 0 FreeSans 480 0 0 0 Tile_X11Y16_DI_SRAM26
port 1451 nsew signal output
flabel metal3 s 486200 78208 487000 78328 0 FreeSans 480 0 0 0 Tile_X11Y16_DI_SRAM27
port 1452 nsew signal output
flabel metal3 s 486200 70728 487000 70848 0 FreeSans 480 0 0 0 Tile_X11Y16_DI_SRAM28
port 1453 nsew signal output
flabel metal3 s 486200 70048 487000 70168 0 FreeSans 480 0 0 0 Tile_X11Y16_DI_SRAM29
port 1454 nsew signal output
flabel metal3 s 486200 60528 487000 60648 0 FreeSans 480 0 0 0 Tile_X11Y16_DI_SRAM3
port 1455 nsew signal output
flabel metal3 s 486200 68688 487000 68808 0 FreeSans 480 0 0 0 Tile_X11Y16_DI_SRAM30
port 1456 nsew signal output
flabel metal3 s 486200 69368 487000 69488 0 FreeSans 480 0 0 0 Tile_X11Y16_DI_SRAM31
port 1457 nsew signal output
flabel metal3 s 486200 63248 487000 63368 0 FreeSans 480 0 0 0 Tile_X11Y16_DI_SRAM4
port 1458 nsew signal output
flabel metal3 s 486200 61888 487000 62008 0 FreeSans 480 0 0 0 Tile_X11Y16_DI_SRAM5
port 1459 nsew signal output
flabel metal3 s 486200 62568 487000 62688 0 FreeSans 480 0 0 0 Tile_X11Y16_DI_SRAM6
port 1460 nsew signal output
flabel metal3 s 486200 61208 487000 61328 0 FreeSans 480 0 0 0 Tile_X11Y16_DI_SRAM7
port 1461 nsew signal output
flabel metal3 s 486200 77528 487000 77648 0 FreeSans 480 0 0 0 Tile_X11Y16_DI_SRAM8
port 1462 nsew signal output
flabel metal3 s 486200 64608 487000 64728 0 FreeSans 480 0 0 0 Tile_X11Y16_DI_SRAM9
port 1463 nsew signal output
flabel metal3 s 486200 25848 487000 25968 0 FreeSans 480 0 0 0 Tile_X11Y16_DO_SRAM0
port 1464 nsew signal input
flabel metal3 s 486200 38768 487000 38888 0 FreeSans 480 0 0 0 Tile_X11Y16_DO_SRAM1
port 1465 nsew signal input
flabel metal3 s 486200 34688 487000 34808 0 FreeSans 480 0 0 0 Tile_X11Y16_DO_SRAM10
port 1466 nsew signal input
flabel metal3 s 486200 41488 487000 41608 0 FreeSans 480 0 0 0 Tile_X11Y16_DO_SRAM11
port 1467 nsew signal input
flabel metal3 s 486200 34008 487000 34128 0 FreeSans 480 0 0 0 Tile_X11Y16_DO_SRAM12
port 1468 nsew signal input
flabel metal3 s 486200 42168 487000 42288 0 FreeSans 480 0 0 0 Tile_X11Y16_DO_SRAM13
port 1469 nsew signal input
flabel metal3 s 486200 33328 487000 33448 0 FreeSans 480 0 0 0 Tile_X11Y16_DO_SRAM14
port 1470 nsew signal input
flabel metal3 s 486200 32648 487000 32768 0 FreeSans 480 0 0 0 Tile_X11Y16_DO_SRAM15
port 1471 nsew signal input
flabel metal3 s 486200 42848 487000 42968 0 FreeSans 480 0 0 0 Tile_X11Y16_DO_SRAM16
port 1472 nsew signal input
flabel metal3 s 486200 31968 487000 32088 0 FreeSans 480 0 0 0 Tile_X11Y16_DO_SRAM17
port 1473 nsew signal input
flabel metal3 s 486200 43528 487000 43648 0 FreeSans 480 0 0 0 Tile_X11Y16_DO_SRAM18
port 1474 nsew signal input
flabel metal3 s 486200 31288 487000 31408 0 FreeSans 480 0 0 0 Tile_X11Y16_DO_SRAM19
port 1475 nsew signal input
flabel metal3 s 486200 38088 487000 38208 0 FreeSans 480 0 0 0 Tile_X11Y16_DO_SRAM2
port 1476 nsew signal input
flabel metal3 s 486200 30608 487000 30728 0 FreeSans 480 0 0 0 Tile_X11Y16_DO_SRAM20
port 1477 nsew signal input
flabel metal3 s 486200 44208 487000 44328 0 FreeSans 480 0 0 0 Tile_X11Y16_DO_SRAM21
port 1478 nsew signal input
flabel metal3 s 486200 29928 487000 30048 0 FreeSans 480 0 0 0 Tile_X11Y16_DO_SRAM22
port 1479 nsew signal input
flabel metal3 s 486200 44888 487000 45008 0 FreeSans 480 0 0 0 Tile_X11Y16_DO_SRAM23
port 1480 nsew signal input
flabel metal3 s 486200 29248 487000 29368 0 FreeSans 480 0 0 0 Tile_X11Y16_DO_SRAM24
port 1481 nsew signal input
flabel metal3 s 486200 28568 487000 28688 0 FreeSans 480 0 0 0 Tile_X11Y16_DO_SRAM25
port 1482 nsew signal input
flabel metal3 s 486200 45568 487000 45688 0 FreeSans 480 0 0 0 Tile_X11Y16_DO_SRAM26
port 1483 nsew signal input
flabel metal3 s 486200 27888 487000 28008 0 FreeSans 480 0 0 0 Tile_X11Y16_DO_SRAM27
port 1484 nsew signal input
flabel metal3 s 486200 46248 487000 46368 0 FreeSans 480 0 0 0 Tile_X11Y16_DO_SRAM28
port 1485 nsew signal input
flabel metal3 s 486200 27208 487000 27328 0 FreeSans 480 0 0 0 Tile_X11Y16_DO_SRAM29
port 1486 nsew signal input
flabel metal3 s 486200 39448 487000 39568 0 FreeSans 480 0 0 0 Tile_X11Y16_DO_SRAM3
port 1487 nsew signal input
flabel metal3 s 486200 26528 487000 26648 0 FreeSans 480 0 0 0 Tile_X11Y16_DO_SRAM30
port 1488 nsew signal input
flabel metal3 s 486200 46928 487000 47048 0 FreeSans 480 0 0 0 Tile_X11Y16_DO_SRAM31
port 1489 nsew signal input
flabel metal3 s 486200 37408 487000 37528 0 FreeSans 480 0 0 0 Tile_X11Y16_DO_SRAM4
port 1490 nsew signal input
flabel metal3 s 486200 36728 487000 36848 0 FreeSans 480 0 0 0 Tile_X11Y16_DO_SRAM5
port 1491 nsew signal input
flabel metal3 s 486200 40128 487000 40248 0 FreeSans 480 0 0 0 Tile_X11Y16_DO_SRAM6
port 1492 nsew signal input
flabel metal3 s 486200 36048 487000 36168 0 FreeSans 480 0 0 0 Tile_X11Y16_DO_SRAM7
port 1493 nsew signal input
flabel metal3 s 486200 40808 487000 40928 0 FreeSans 480 0 0 0 Tile_X11Y16_DO_SRAM8
port 1494 nsew signal input
flabel metal3 s 486200 35368 487000 35488 0 FreeSans 480 0 0 0 Tile_X11Y16_DO_SRAM9
port 1495 nsew signal input
flabel metal3 s 486200 74808 487000 74928 0 FreeSans 480 0 0 0 Tile_X11Y16_EN_SRAM
port 1496 nsew signal output
flabel metal3 s 486200 72768 487000 72888 0 FreeSans 480 0 0 0 Tile_X11Y16_R_WB_SRAM
port 1497 nsew signal output
flabel metal3 s 486200 753448 487000 753568 0 FreeSans 480 0 0 0 Tile_X11Y2_AD_SRAM0
port 1498 nsew signal output
flabel metal3 s 486200 680688 487000 680808 0 FreeSans 480 0 0 0 Tile_X11Y2_AD_SRAM1
port 1499 nsew signal output
flabel metal3 s 486200 739168 487000 739288 0 FreeSans 480 0 0 0 Tile_X11Y2_AD_SRAM2
port 1500 nsew signal output
flabel metal3 s 486200 694968 487000 695088 0 FreeSans 480 0 0 0 Tile_X11Y2_AD_SRAM3
port 1501 nsew signal output
flabel metal3 s 486200 748688 487000 748808 0 FreeSans 480 0 0 0 Tile_X11Y2_AD_SRAM4
port 1502 nsew signal output
flabel metal3 s 486200 724208 487000 724328 0 FreeSans 480 0 0 0 Tile_X11Y2_AD_SRAM5
port 1503 nsew signal output
flabel metal3 s 486200 707208 487000 707328 0 FreeSans 480 0 0 0 Tile_X11Y2_AD_SRAM6
port 1504 nsew signal output
flabel metal3 s 486200 691568 487000 691688 0 FreeSans 480 0 0 0 Tile_X11Y2_AD_SRAM7
port 1505 nsew signal output
flabel metal3 s 486200 739848 487000 739968 0 FreeSans 480 0 0 0 Tile_X11Y2_AD_SRAM8
port 1506 nsew signal output
flabel metal3 s 486200 726928 487000 727048 0 FreeSans 480 0 0 0 Tile_X11Y2_AD_SRAM9
port 1507 nsew signal output
flabel metal3 s 486200 751408 487000 751528 0 FreeSans 480 0 0 0 Tile_X11Y2_BEN_SRAM0
port 1508 nsew signal output
flabel metal3 s 486200 685448 487000 685568 0 FreeSans 480 0 0 0 Tile_X11Y2_BEN_SRAM1
port 1509 nsew signal output
flabel metal3 s 486200 724888 487000 725008 0 FreeSans 480 0 0 0 Tile_X11Y2_BEN_SRAM10
port 1510 nsew signal output
flabel metal3 s 486200 690888 487000 691008 0 FreeSans 480 0 0 0 Tile_X11Y2_BEN_SRAM11
port 1511 nsew signal output
flabel metal3 s 486200 722168 487000 722288 0 FreeSans 480 0 0 0 Tile_X11Y2_BEN_SRAM12
port 1512 nsew signal output
flabel metal3 s 486200 740528 487000 740648 0 FreeSans 480 0 0 0 Tile_X11Y2_BEN_SRAM13
port 1513 nsew signal output
flabel metal3 s 486200 700408 487000 700528 0 FreeSans 480 0 0 0 Tile_X11Y2_BEN_SRAM14
port 1514 nsew signal output
flabel metal3 s 486200 749368 487000 749488 0 FreeSans 480 0 0 0 Tile_X11Y2_BEN_SRAM15
port 1515 nsew signal output
flabel metal3 s 486200 686128 487000 686248 0 FreeSans 480 0 0 0 Tile_X11Y2_BEN_SRAM16
port 1516 nsew signal output
flabel metal3 s 486200 741208 487000 741328 0 FreeSans 480 0 0 0 Tile_X11Y2_BEN_SRAM17
port 1517 nsew signal output
flabel metal3 s 486200 718088 487000 718208 0 FreeSans 480 0 0 0 Tile_X11Y2_BEN_SRAM18
port 1518 nsew signal output
flabel metal3 s 486200 702448 487000 702568 0 FreeSans 480 0 0 0 Tile_X11Y2_BEN_SRAM19
port 1519 nsew signal output
flabel metal3 s 486200 692928 487000 693048 0 FreeSans 480 0 0 0 Tile_X11Y2_BEN_SRAM2
port 1520 nsew signal output
flabel metal3 s 486200 717408 487000 717528 0 FreeSans 480 0 0 0 Tile_X11Y2_BEN_SRAM20
port 1521 nsew signal output
flabel metal3 s 486200 741888 487000 742008 0 FreeSans 480 0 0 0 Tile_X11Y2_BEN_SRAM21
port 1522 nsew signal output
flabel metal3 s 486200 729648 487000 729768 0 FreeSans 480 0 0 0 Tile_X11Y2_BEN_SRAM22
port 1523 nsew signal output
flabel metal3 s 486200 716048 487000 716168 0 FreeSans 480 0 0 0 Tile_X11Y2_BEN_SRAM23
port 1524 nsew signal output
flabel metal3 s 486200 698368 487000 698488 0 FreeSans 480 0 0 0 Tile_X11Y2_BEN_SRAM24
port 1525 nsew signal output
flabel metal3 s 486200 715368 487000 715488 0 FreeSans 480 0 0 0 Tile_X11Y2_BEN_SRAM25
port 1526 nsew signal output
flabel metal3 s 486200 687488 487000 687608 0 FreeSans 480 0 0 0 Tile_X11Y2_BEN_SRAM26
port 1527 nsew signal output
flabel metal3 s 486200 714688 487000 714808 0 FreeSans 480 0 0 0 Tile_X11Y2_BEN_SRAM27
port 1528 nsew signal output
flabel metal3 s 486200 742568 487000 742688 0 FreeSans 480 0 0 0 Tile_X11Y2_BEN_SRAM28
port 1529 nsew signal output
flabel metal3 s 486200 695648 487000 695768 0 FreeSans 480 0 0 0 Tile_X11Y2_BEN_SRAM29
port 1530 nsew signal output
flabel metal3 s 486200 727608 487000 727728 0 FreeSans 480 0 0 0 Tile_X11Y2_BEN_SRAM3
port 1531 nsew signal output
flabel metal3 s 486200 752088 487000 752208 0 FreeSans 480 0 0 0 Tile_X11Y2_BEN_SRAM30
port 1532 nsew signal output
flabel metal3 s 486200 688848 487000 688968 0 FreeSans 480 0 0 0 Tile_X11Y2_BEN_SRAM31
port 1533 nsew signal output
flabel metal3 s 486200 682048 487000 682168 0 FreeSans 480 0 0 0 Tile_X11Y2_BEN_SRAM4
port 1534 nsew signal output
flabel metal3 s 486200 728288 487000 728408 0 FreeSans 480 0 0 0 Tile_X11Y2_BEN_SRAM5
port 1535 nsew signal output
flabel metal3 s 486200 683408 487000 683528 0 FreeSans 480 0 0 0 Tile_X11Y2_BEN_SRAM6
port 1536 nsew signal output
flabel metal3 s 486200 743248 487000 743368 0 FreeSans 480 0 0 0 Tile_X11Y2_BEN_SRAM7
port 1537 nsew signal output
flabel metal3 s 486200 728968 487000 729088 0 FreeSans 480 0 0 0 Tile_X11Y2_BEN_SRAM8
port 1538 nsew signal output
flabel metal3 s 486200 705168 487000 705288 0 FreeSans 480 0 0 0 Tile_X11Y2_BEN_SRAM9
port 1539 nsew signal output
flabel metal3 s 486200 732368 487000 732488 0 FreeSans 480 0 0 0 Tile_X11Y2_CLOCK_SRAM
port 1540 nsew signal output
flabel metal3 s 486200 711968 487000 712088 0 FreeSans 480 0 0 0 Tile_X11Y2_DI_SRAM0
port 1541 nsew signal output
flabel metal3 s 486200 689528 487000 689648 0 FreeSans 480 0 0 0 Tile_X11Y2_DI_SRAM1
port 1542 nsew signal output
flabel metal3 s 486200 711288 487000 711408 0 FreeSans 480 0 0 0 Tile_X11Y2_DI_SRAM10
port 1543 nsew signal output
flabel metal3 s 486200 701088 487000 701208 0 FreeSans 480 0 0 0 Tile_X11Y2_DI_SRAM11
port 1544 nsew signal output
flabel metal3 s 486200 750048 487000 750168 0 FreeSans 480 0 0 0 Tile_X11Y2_DI_SRAM12
port 1545 nsew signal output
flabel metal3 s 486200 743928 487000 744048 0 FreeSans 480 0 0 0 Tile_X11Y2_DI_SRAM13
port 1546 nsew signal output
flabel metal3 s 486200 726248 487000 726368 0 FreeSans 480 0 0 0 Tile_X11Y2_DI_SRAM14
port 1547 nsew signal output
flabel metal3 s 486200 709928 487000 710048 0 FreeSans 480 0 0 0 Tile_X11Y2_DI_SRAM15
port 1548 nsew signal output
flabel metal3 s 486200 693608 487000 693728 0 FreeSans 480 0 0 0 Tile_X11Y2_DI_SRAM16
port 1549 nsew signal output
flabel metal3 s 486200 708568 487000 708688 0 FreeSans 480 0 0 0 Tile_X11Y2_DI_SRAM17
port 1550 nsew signal output
flabel metal3 s 486200 744608 487000 744728 0 FreeSans 480 0 0 0 Tile_X11Y2_DI_SRAM18
port 1551 nsew signal output
flabel metal3 s 486200 704488 487000 704608 0 FreeSans 480 0 0 0 Tile_X11Y2_DI_SRAM19
port 1552 nsew signal output
flabel metal3 s 486200 723528 487000 723648 0 FreeSans 480 0 0 0 Tile_X11Y2_DI_SRAM2
port 1553 nsew signal output
flabel metal3 s 486200 730328 487000 730448 0 FreeSans 480 0 0 0 Tile_X11Y2_DI_SRAM20
port 1554 nsew signal output
flabel metal3 s 486200 709248 487000 709368 0 FreeSans 480 0 0 0 Tile_X11Y2_DI_SRAM21
port 1555 nsew signal output
flabel metal3 s 486200 703128 487000 703248 0 FreeSans 480 0 0 0 Tile_X11Y2_DI_SRAM22
port 1556 nsew signal output
flabel metal3 s 486200 731008 487000 731128 0 FreeSans 480 0 0 0 Tile_X11Y2_DI_SRAM23
port 1557 nsew signal output
flabel metal3 s 486200 713328 487000 713448 0 FreeSans 480 0 0 0 Tile_X11Y2_DI_SRAM24
port 1558 nsew signal output
flabel metal3 s 486200 745288 487000 745408 0 FreeSans 480 0 0 0 Tile_X11Y2_DI_SRAM25
port 1559 nsew signal output
flabel metal3 s 486200 699048 487000 699168 0 FreeSans 480 0 0 0 Tile_X11Y2_DI_SRAM26
port 1560 nsew signal output
flabel metal3 s 486200 707888 487000 708008 0 FreeSans 480 0 0 0 Tile_X11Y2_DI_SRAM27
port 1561 nsew signal output
flabel metal3 s 486200 719448 487000 719568 0 FreeSans 480 0 0 0 Tile_X11Y2_DI_SRAM28
port 1562 nsew signal output
flabel metal3 s 486200 722848 487000 722968 0 FreeSans 480 0 0 0 Tile_X11Y2_DI_SRAM29
port 1563 nsew signal output
flabel metal3 s 486200 710608 487000 710728 0 FreeSans 480 0 0 0 Tile_X11Y2_DI_SRAM3
port 1564 nsew signal output
flabel metal3 s 486200 725568 487000 725688 0 FreeSans 480 0 0 0 Tile_X11Y2_DI_SRAM30
port 1565 nsew signal output
flabel metal3 s 486200 697688 487000 697808 0 FreeSans 480 0 0 0 Tile_X11Y2_DI_SRAM31
port 1566 nsew signal output
flabel metal3 s 486200 745968 487000 746088 0 FreeSans 480 0 0 0 Tile_X11Y2_DI_SRAM4
port 1567 nsew signal output
flabel metal3 s 486200 731688 487000 731808 0 FreeSans 480 0 0 0 Tile_X11Y2_DI_SRAM5
port 1568 nsew signal output
flabel metal3 s 486200 733048 487000 733168 0 FreeSans 480 0 0 0 Tile_X11Y2_DI_SRAM6
port 1569 nsew signal output
flabel metal3 s 486200 692248 487000 692368 0 FreeSans 480 0 0 0 Tile_X11Y2_DI_SRAM7
port 1570 nsew signal output
flabel metal3 s 486200 750728 487000 750848 0 FreeSans 480 0 0 0 Tile_X11Y2_DI_SRAM8
port 1571 nsew signal output
flabel metal3 s 486200 696328 487000 696448 0 FreeSans 480 0 0 0 Tile_X11Y2_DI_SRAM9
port 1572 nsew signal output
flabel metal3 s 486200 701768 487000 701888 0 FreeSans 480 0 0 0 Tile_X11Y2_DO_SRAM0
port 1573 nsew signal input
flabel metal3 s 486200 736448 487000 736568 0 FreeSans 480 0 0 0 Tile_X11Y2_DO_SRAM1
port 1574 nsew signal input
flabel metal3 s 486200 690208 487000 690328 0 FreeSans 480 0 0 0 Tile_X11Y2_DO_SRAM10
port 1575 nsew signal input
flabel metal3 s 486200 746648 487000 746768 0 FreeSans 480 0 0 0 Tile_X11Y2_DO_SRAM11
port 1576 nsew signal input
flabel metal3 s 486200 733728 487000 733848 0 FreeSans 480 0 0 0 Tile_X11Y2_DO_SRAM12
port 1577 nsew signal input
flabel metal3 s 486200 681368 487000 681488 0 FreeSans 480 0 0 0 Tile_X11Y2_DO_SRAM13
port 1578 nsew signal input
flabel metal3 s 486200 688168 487000 688288 0 FreeSans 480 0 0 0 Tile_X11Y2_DO_SRAM14
port 1579 nsew signal input
flabel metal3 s 486200 718768 487000 718888 0 FreeSans 480 0 0 0 Tile_X11Y2_DO_SRAM15
port 1580 nsew signal input
flabel metal3 s 486200 734408 487000 734528 0 FreeSans 480 0 0 0 Tile_X11Y2_DO_SRAM16
port 1581 nsew signal input
flabel metal3 s 486200 720128 487000 720248 0 FreeSans 480 0 0 0 Tile_X11Y2_DO_SRAM17
port 1582 nsew signal input
flabel metal3 s 486200 747328 487000 747448 0 FreeSans 480 0 0 0 Tile_X11Y2_DO_SRAM18
port 1583 nsew signal input
flabel metal3 s 486200 714008 487000 714128 0 FreeSans 480 0 0 0 Tile_X11Y2_DO_SRAM19
port 1584 nsew signal input
flabel metal3 s 486200 735088 487000 735208 0 FreeSans 480 0 0 0 Tile_X11Y2_DO_SRAM2
port 1585 nsew signal input
flabel metal3 s 486200 680008 487000 680128 0 FreeSans 480 0 0 0 Tile_X11Y2_DO_SRAM20
port 1586 nsew signal input
flabel metal3 s 486200 682728 487000 682848 0 FreeSans 480 0 0 0 Tile_X11Y2_DO_SRAM21
port 1587 nsew signal input
flabel metal3 s 486200 684088 487000 684208 0 FreeSans 480 0 0 0 Tile_X11Y2_DO_SRAM22
port 1588 nsew signal input
flabel metal3 s 486200 735768 487000 735888 0 FreeSans 480 0 0 0 Tile_X11Y2_DO_SRAM23
port 1589 nsew signal input
flabel metal3 s 486200 699728 487000 699848 0 FreeSans 480 0 0 0 Tile_X11Y2_DO_SRAM24
port 1590 nsew signal input
flabel metal3 s 486200 703808 487000 703928 0 FreeSans 480 0 0 0 Tile_X11Y2_DO_SRAM25
port 1591 nsew signal input
flabel metal3 s 486200 684768 487000 684888 0 FreeSans 480 0 0 0 Tile_X11Y2_DO_SRAM26
port 1592 nsew signal input
flabel metal3 s 486200 748008 487000 748128 0 FreeSans 480 0 0 0 Tile_X11Y2_DO_SRAM27
port 1593 nsew signal input
flabel metal3 s 486200 697008 487000 697128 0 FreeSans 480 0 0 0 Tile_X11Y2_DO_SRAM28
port 1594 nsew signal input
flabel metal3 s 486200 686808 487000 686928 0 FreeSans 480 0 0 0 Tile_X11Y2_DO_SRAM29
port 1595 nsew signal input
flabel metal3 s 486200 737128 487000 737248 0 FreeSans 480 0 0 0 Tile_X11Y2_DO_SRAM3
port 1596 nsew signal input
flabel metal3 s 486200 752768 487000 752888 0 FreeSans 480 0 0 0 Tile_X11Y2_DO_SRAM30
port 1597 nsew signal input
flabel metal3 s 486200 712648 487000 712768 0 FreeSans 480 0 0 0 Tile_X11Y2_DO_SRAM31
port 1598 nsew signal input
flabel metal3 s 486200 737808 487000 737928 0 FreeSans 480 0 0 0 Tile_X11Y2_DO_SRAM4
port 1599 nsew signal input
flabel metal3 s 486200 694288 487000 694408 0 FreeSans 480 0 0 0 Tile_X11Y2_DO_SRAM5
port 1600 nsew signal input
flabel metal3 s 486200 716728 487000 716848 0 FreeSans 480 0 0 0 Tile_X11Y2_DO_SRAM6
port 1601 nsew signal input
flabel metal3 s 486200 721488 487000 721608 0 FreeSans 480 0 0 0 Tile_X11Y2_DO_SRAM7
port 1602 nsew signal input
flabel metal3 s 486200 706528 487000 706648 0 FreeSans 480 0 0 0 Tile_X11Y2_DO_SRAM8
port 1603 nsew signal input
flabel metal3 s 486200 738488 487000 738608 0 FreeSans 480 0 0 0 Tile_X11Y2_DO_SRAM9
port 1604 nsew signal input
flabel metal3 s 486200 705848 487000 705968 0 FreeSans 480 0 0 0 Tile_X11Y2_EN_SRAM
port 1605 nsew signal output
flabel metal3 s 486200 720808 487000 720928 0 FreeSans 480 0 0 0 Tile_X11Y2_R_WB_SRAM
port 1606 nsew signal output
flabel metal3 s 486200 556928 487000 557048 0 FreeSans 480 0 0 0 Tile_X11Y4_AD_SRAM0
port 1607 nsew signal output
flabel metal3 s 486200 587528 487000 587648 0 FreeSans 480 0 0 0 Tile_X11Y4_AD_SRAM1
port 1608 nsew signal output
flabel metal3 s 486200 565088 487000 565208 0 FreeSans 480 0 0 0 Tile_X11Y4_AD_SRAM2
port 1609 nsew signal output
flabel metal3 s 486200 588208 487000 588328 0 FreeSans 480 0 0 0 Tile_X11Y4_AD_SRAM3
port 1610 nsew signal output
flabel metal3 s 486200 564408 487000 564528 0 FreeSans 480 0 0 0 Tile_X11Y4_AD_SRAM4
port 1611 nsew signal output
flabel metal3 s 486200 563728 487000 563848 0 FreeSans 480 0 0 0 Tile_X11Y4_AD_SRAM5
port 1612 nsew signal output
flabel metal3 s 486200 588888 487000 589008 0 FreeSans 480 0 0 0 Tile_X11Y4_AD_SRAM6
port 1613 nsew signal output
flabel metal3 s 486200 563048 487000 563168 0 FreeSans 480 0 0 0 Tile_X11Y4_AD_SRAM7
port 1614 nsew signal output
flabel metal3 s 486200 589568 487000 589688 0 FreeSans 480 0 0 0 Tile_X11Y4_AD_SRAM8
port 1615 nsew signal output
flabel metal3 s 486200 562368 487000 562488 0 FreeSans 480 0 0 0 Tile_X11Y4_AD_SRAM9
port 1616 nsew signal output
flabel metal3 s 486200 561688 487000 561808 0 FreeSans 480 0 0 0 Tile_X11Y4_BEN_SRAM0
port 1617 nsew signal output
flabel metal3 s 486200 590248 487000 590368 0 FreeSans 480 0 0 0 Tile_X11Y4_BEN_SRAM1
port 1618 nsew signal output
flabel metal3 s 486200 557608 487000 557728 0 FreeSans 480 0 0 0 Tile_X11Y4_BEN_SRAM10
port 1619 nsew signal output
flabel metal3 s 486200 592968 487000 593088 0 FreeSans 480 0 0 0 Tile_X11Y4_BEN_SRAM11
port 1620 nsew signal output
flabel metal3 s 486200 593648 487000 593768 0 FreeSans 480 0 0 0 Tile_X11Y4_BEN_SRAM12
port 1621 nsew signal output
flabel metal3 s 486200 630368 487000 630488 0 FreeSans 480 0 0 0 Tile_X11Y4_BEN_SRAM13
port 1622 nsew signal output
flabel metal3 s 486200 629688 487000 629808 0 FreeSans 480 0 0 0 Tile_X11Y4_BEN_SRAM14
port 1623 nsew signal output
flabel metal3 s 486200 594328 487000 594448 0 FreeSans 480 0 0 0 Tile_X11Y4_BEN_SRAM15
port 1624 nsew signal output
flabel metal3 s 486200 629008 487000 629128 0 FreeSans 480 0 0 0 Tile_X11Y4_BEN_SRAM16
port 1625 nsew signal output
flabel metal3 s 486200 595008 487000 595128 0 FreeSans 480 0 0 0 Tile_X11Y4_BEN_SRAM17
port 1626 nsew signal output
flabel metal3 s 486200 628328 487000 628448 0 FreeSans 480 0 0 0 Tile_X11Y4_BEN_SRAM18
port 1627 nsew signal output
flabel metal3 s 486200 627648 487000 627768 0 FreeSans 480 0 0 0 Tile_X11Y4_BEN_SRAM19
port 1628 nsew signal output
flabel metal3 s 486200 561008 487000 561128 0 FreeSans 480 0 0 0 Tile_X11Y4_BEN_SRAM2
port 1629 nsew signal output
flabel metal3 s 486200 595688 487000 595808 0 FreeSans 480 0 0 0 Tile_X11Y4_BEN_SRAM20
port 1630 nsew signal output
flabel metal3 s 486200 626968 487000 627088 0 FreeSans 480 0 0 0 Tile_X11Y4_BEN_SRAM21
port 1631 nsew signal output
flabel metal3 s 486200 596368 487000 596488 0 FreeSans 480 0 0 0 Tile_X11Y4_BEN_SRAM22
port 1632 nsew signal output
flabel metal3 s 486200 626288 487000 626408 0 FreeSans 480 0 0 0 Tile_X11Y4_BEN_SRAM23
port 1633 nsew signal output
flabel metal3 s 486200 625608 487000 625728 0 FreeSans 480 0 0 0 Tile_X11Y4_BEN_SRAM24
port 1634 nsew signal output
flabel metal3 s 486200 597048 487000 597168 0 FreeSans 480 0 0 0 Tile_X11Y4_BEN_SRAM25
port 1635 nsew signal output
flabel metal3 s 486200 624928 487000 625048 0 FreeSans 480 0 0 0 Tile_X11Y4_BEN_SRAM26
port 1636 nsew signal output
flabel metal3 s 486200 597728 487000 597848 0 FreeSans 480 0 0 0 Tile_X11Y4_BEN_SRAM27
port 1637 nsew signal output
flabel metal3 s 486200 624248 487000 624368 0 FreeSans 480 0 0 0 Tile_X11Y4_BEN_SRAM28
port 1638 nsew signal output
flabel metal3 s 486200 623568 487000 623688 0 FreeSans 480 0 0 0 Tile_X11Y4_BEN_SRAM29
port 1639 nsew signal output
flabel metal3 s 486200 590928 487000 591048 0 FreeSans 480 0 0 0 Tile_X11Y4_BEN_SRAM3
port 1640 nsew signal output
flabel metal3 s 486200 598408 487000 598528 0 FreeSans 480 0 0 0 Tile_X11Y4_BEN_SRAM30
port 1641 nsew signal output
flabel metal3 s 486200 622888 487000 623008 0 FreeSans 480 0 0 0 Tile_X11Y4_BEN_SRAM31
port 1642 nsew signal output
flabel metal3 s 486200 560328 487000 560448 0 FreeSans 480 0 0 0 Tile_X11Y4_BEN_SRAM4
port 1643 nsew signal output
flabel metal3 s 486200 559648 487000 559768 0 FreeSans 480 0 0 0 Tile_X11Y4_BEN_SRAM5
port 1644 nsew signal output
flabel metal3 s 486200 591608 487000 591728 0 FreeSans 480 0 0 0 Tile_X11Y4_BEN_SRAM6
port 1645 nsew signal output
flabel metal3 s 486200 558968 487000 559088 0 FreeSans 480 0 0 0 Tile_X11Y4_BEN_SRAM7
port 1646 nsew signal output
flabel metal3 s 486200 592288 487000 592408 0 FreeSans 480 0 0 0 Tile_X11Y4_BEN_SRAM8
port 1647 nsew signal output
flabel metal3 s 486200 558288 487000 558408 0 FreeSans 480 0 0 0 Tile_X11Y4_BEN_SRAM9
port 1648 nsew signal output
flabel metal3 s 486200 599088 487000 599208 0 FreeSans 480 0 0 0 Tile_X11Y4_CLOCK_SRAM
port 1649 nsew signal output
flabel metal3 s 486200 622208 487000 622328 0 FreeSans 480 0 0 0 Tile_X11Y4_DI_SRAM0
port 1650 nsew signal output
flabel metal3 s 486200 621528 487000 621648 0 FreeSans 480 0 0 0 Tile_X11Y4_DI_SRAM1
port 1651 nsew signal output
flabel metal3 s 486200 620848 487000 620968 0 FreeSans 480 0 0 0 Tile_X11Y4_DI_SRAM10
port 1652 nsew signal output
flabel metal3 s 486200 617448 487000 617568 0 FreeSans 480 0 0 0 Tile_X11Y4_DI_SRAM11
port 1653 nsew signal output
flabel metal3 s 486200 612008 487000 612128 0 FreeSans 480 0 0 0 Tile_X11Y4_DI_SRAM12
port 1654 nsew signal output
flabel metal3 s 486200 616768 487000 616888 0 FreeSans 480 0 0 0 Tile_X11Y4_DI_SRAM13
port 1655 nsew signal output
flabel metal3 s 486200 604528 487000 604648 0 FreeSans 480 0 0 0 Tile_X11Y4_DI_SRAM14
port 1656 nsew signal output
flabel metal3 s 486200 619488 487000 619608 0 FreeSans 480 0 0 0 Tile_X11Y4_DI_SRAM15
port 1657 nsew signal output
flabel metal3 s 486200 615408 487000 615528 0 FreeSans 480 0 0 0 Tile_X11Y4_DI_SRAM16
port 1658 nsew signal output
flabel metal3 s 486200 603848 487000 603968 0 FreeSans 480 0 0 0 Tile_X11Y4_DI_SRAM17
port 1659 nsew signal output
flabel metal3 s 486200 614728 487000 614848 0 FreeSans 480 0 0 0 Tile_X11Y4_DI_SRAM18
port 1660 nsew signal output
flabel metal3 s 486200 607928 487000 608048 0 FreeSans 480 0 0 0 Tile_X11Y4_DI_SRAM19
port 1661 nsew signal output
flabel metal3 s 486200 599768 487000 599888 0 FreeSans 480 0 0 0 Tile_X11Y4_DI_SRAM2
port 1662 nsew signal output
flabel metal3 s 486200 614048 487000 614168 0 FreeSans 480 0 0 0 Tile_X11Y4_DI_SRAM20
port 1663 nsew signal output
flabel metal3 s 486200 613368 487000 613488 0 FreeSans 480 0 0 0 Tile_X11Y4_DI_SRAM21
port 1664 nsew signal output
flabel metal3 s 486200 605208 487000 605328 0 FreeSans 480 0 0 0 Tile_X11Y4_DI_SRAM22
port 1665 nsew signal output
flabel metal3 s 486200 618808 487000 618928 0 FreeSans 480 0 0 0 Tile_X11Y4_DI_SRAM23
port 1666 nsew signal output
flabel metal3 s 486200 607248 487000 607368 0 FreeSans 480 0 0 0 Tile_X11Y4_DI_SRAM24
port 1667 nsew signal output
flabel metal3 s 486200 618128 487000 618248 0 FreeSans 480 0 0 0 Tile_X11Y4_DI_SRAM25
port 1668 nsew signal output
flabel metal3 s 486200 611328 487000 611448 0 FreeSans 480 0 0 0 Tile_X11Y4_DI_SRAM26
port 1669 nsew signal output
flabel metal3 s 486200 606568 487000 606688 0 FreeSans 480 0 0 0 Tile_X11Y4_DI_SRAM27
port 1670 nsew signal output
flabel metal3 s 486200 610648 487000 610768 0 FreeSans 480 0 0 0 Tile_X11Y4_DI_SRAM28
port 1671 nsew signal output
flabel metal3 s 486200 620168 487000 620288 0 FreeSans 480 0 0 0 Tile_X11Y4_DI_SRAM29
port 1672 nsew signal output
flabel metal3 s 486200 600448 487000 600568 0 FreeSans 480 0 0 0 Tile_X11Y4_DI_SRAM3
port 1673 nsew signal output
flabel metal3 s 486200 609968 487000 610088 0 FreeSans 480 0 0 0 Tile_X11Y4_DI_SRAM30
port 1674 nsew signal output
flabel metal3 s 486200 609288 487000 609408 0 FreeSans 480 0 0 0 Tile_X11Y4_DI_SRAM31
port 1675 nsew signal output
flabel metal3 s 486200 608608 487000 608728 0 FreeSans 480 0 0 0 Tile_X11Y4_DI_SRAM4
port 1676 nsew signal output
flabel metal3 s 486200 601128 487000 601248 0 FreeSans 480 0 0 0 Tile_X11Y4_DI_SRAM5
port 1677 nsew signal output
flabel metal3 s 486200 601808 487000 601928 0 FreeSans 480 0 0 0 Tile_X11Y4_DI_SRAM6
port 1678 nsew signal output
flabel metal3 s 486200 602488 487000 602608 0 FreeSans 480 0 0 0 Tile_X11Y4_DI_SRAM7
port 1679 nsew signal output
flabel metal3 s 486200 603168 487000 603288 0 FreeSans 480 0 0 0 Tile_X11Y4_DI_SRAM8
port 1680 nsew signal output
flabel metal3 s 486200 605888 487000 606008 0 FreeSans 480 0 0 0 Tile_X11Y4_DI_SRAM9
port 1681 nsew signal output
flabel metal3 s 486200 565768 487000 565888 0 FreeSans 480 0 0 0 Tile_X11Y4_DO_SRAM0
port 1682 nsew signal input
flabel metal3 s 486200 578688 487000 578808 0 FreeSans 480 0 0 0 Tile_X11Y4_DO_SRAM1
port 1683 nsew signal input
flabel metal3 s 486200 581408 487000 581528 0 FreeSans 480 0 0 0 Tile_X11Y4_DO_SRAM10
port 1684 nsew signal input
flabel metal3 s 486200 574608 487000 574728 0 FreeSans 480 0 0 0 Tile_X11Y4_DO_SRAM11
port 1685 nsew signal input
flabel metal3 s 486200 573928 487000 574048 0 FreeSans 480 0 0 0 Tile_X11Y4_DO_SRAM12
port 1686 nsew signal input
flabel metal3 s 486200 582088 487000 582208 0 FreeSans 480 0 0 0 Tile_X11Y4_DO_SRAM13
port 1687 nsew signal input
flabel metal3 s 486200 573248 487000 573368 0 FreeSans 480 0 0 0 Tile_X11Y4_DO_SRAM14
port 1688 nsew signal input
flabel metal3 s 486200 582768 487000 582888 0 FreeSans 480 0 0 0 Tile_X11Y4_DO_SRAM15
port 1689 nsew signal input
flabel metal3 s 486200 572568 487000 572688 0 FreeSans 480 0 0 0 Tile_X11Y4_DO_SRAM16
port 1690 nsew signal input
flabel metal3 s 486200 571888 487000 572008 0 FreeSans 480 0 0 0 Tile_X11Y4_DO_SRAM17
port 1691 nsew signal input
flabel metal3 s 486200 583448 487000 583568 0 FreeSans 480 0 0 0 Tile_X11Y4_DO_SRAM18
port 1692 nsew signal input
flabel metal3 s 486200 571208 487000 571328 0 FreeSans 480 0 0 0 Tile_X11Y4_DO_SRAM19
port 1693 nsew signal input
flabel metal3 s 486200 578008 487000 578128 0 FreeSans 480 0 0 0 Tile_X11Y4_DO_SRAM2
port 1694 nsew signal input
flabel metal3 s 486200 584128 487000 584248 0 FreeSans 480 0 0 0 Tile_X11Y4_DO_SRAM20
port 1695 nsew signal input
flabel metal3 s 486200 570528 487000 570648 0 FreeSans 480 0 0 0 Tile_X11Y4_DO_SRAM21
port 1696 nsew signal input
flabel metal3 s 486200 569848 487000 569968 0 FreeSans 480 0 0 0 Tile_X11Y4_DO_SRAM22
port 1697 nsew signal input
flabel metal3 s 486200 584808 487000 584928 0 FreeSans 480 0 0 0 Tile_X11Y4_DO_SRAM23
port 1698 nsew signal input
flabel metal3 s 486200 569168 487000 569288 0 FreeSans 480 0 0 0 Tile_X11Y4_DO_SRAM24
port 1699 nsew signal input
flabel metal3 s 486200 585488 487000 585608 0 FreeSans 480 0 0 0 Tile_X11Y4_DO_SRAM25
port 1700 nsew signal input
flabel metal3 s 486200 568488 487000 568608 0 FreeSans 480 0 0 0 Tile_X11Y4_DO_SRAM26
port 1701 nsew signal input
flabel metal3 s 486200 567808 487000 567928 0 FreeSans 480 0 0 0 Tile_X11Y4_DO_SRAM27
port 1702 nsew signal input
flabel metal3 s 486200 586168 487000 586288 0 FreeSans 480 0 0 0 Tile_X11Y4_DO_SRAM28
port 1703 nsew signal input
flabel metal3 s 486200 567128 487000 567248 0 FreeSans 480 0 0 0 Tile_X11Y4_DO_SRAM29
port 1704 nsew signal input
flabel metal3 s 486200 579368 487000 579488 0 FreeSans 480 0 0 0 Tile_X11Y4_DO_SRAM3
port 1705 nsew signal input
flabel metal3 s 486200 586848 487000 586968 0 FreeSans 480 0 0 0 Tile_X11Y4_DO_SRAM30
port 1706 nsew signal input
flabel metal3 s 486200 566448 487000 566568 0 FreeSans 480 0 0 0 Tile_X11Y4_DO_SRAM31
port 1707 nsew signal input
flabel metal3 s 486200 577328 487000 577448 0 FreeSans 480 0 0 0 Tile_X11Y4_DO_SRAM4
port 1708 nsew signal input
flabel metal3 s 486200 580048 487000 580168 0 FreeSans 480 0 0 0 Tile_X11Y4_DO_SRAM5
port 1709 nsew signal input
flabel metal3 s 486200 576648 487000 576768 0 FreeSans 480 0 0 0 Tile_X11Y4_DO_SRAM6
port 1710 nsew signal input
flabel metal3 s 486200 575968 487000 576088 0 FreeSans 480 0 0 0 Tile_X11Y4_DO_SRAM7
port 1711 nsew signal input
flabel metal3 s 486200 580728 487000 580848 0 FreeSans 480 0 0 0 Tile_X11Y4_DO_SRAM8
port 1712 nsew signal input
flabel metal3 s 486200 575288 487000 575408 0 FreeSans 480 0 0 0 Tile_X11Y4_DO_SRAM9
port 1713 nsew signal input
flabel metal3 s 486200 616088 487000 616208 0 FreeSans 480 0 0 0 Tile_X11Y4_EN_SRAM
port 1714 nsew signal output
flabel metal3 s 486200 612688 487000 612808 0 FreeSans 480 0 0 0 Tile_X11Y4_R_WB_SRAM
port 1715 nsew signal output
flabel metal3 s 486200 466488 487000 466608 0 FreeSans 480 0 0 0 Tile_X11Y6_AD_SRAM0
port 1716 nsew signal output
flabel metal3 s 486200 475328 487000 475448 0 FreeSans 480 0 0 0 Tile_X11Y6_AD_SRAM1
port 1717 nsew signal output
flabel metal3 s 486200 497768 487000 497888 0 FreeSans 480 0 0 0 Tile_X11Y6_AD_SRAM2
port 1718 nsew signal output
flabel metal3 s 486200 474648 487000 474768 0 FreeSans 480 0 0 0 Tile_X11Y6_AD_SRAM3
port 1719 nsew signal output
flabel metal3 s 486200 498448 487000 498568 0 FreeSans 480 0 0 0 Tile_X11Y6_AD_SRAM4
port 1720 nsew signal output
flabel metal3 s 486200 473968 487000 474088 0 FreeSans 480 0 0 0 Tile_X11Y6_AD_SRAM5
port 1721 nsew signal output
flabel metal3 s 486200 473288 487000 473408 0 FreeSans 480 0 0 0 Tile_X11Y6_AD_SRAM6
port 1722 nsew signal output
flabel metal3 s 486200 499128 487000 499248 0 FreeSans 480 0 0 0 Tile_X11Y6_AD_SRAM7
port 1723 nsew signal output
flabel metal3 s 486200 472608 487000 472728 0 FreeSans 480 0 0 0 Tile_X11Y6_AD_SRAM8
port 1724 nsew signal output
flabel metal3 s 486200 499808 487000 499928 0 FreeSans 480 0 0 0 Tile_X11Y6_AD_SRAM9
port 1725 nsew signal output
flabel metal3 s 486200 471928 487000 472048 0 FreeSans 480 0 0 0 Tile_X11Y6_BEN_SRAM0
port 1726 nsew signal output
flabel metal3 s 486200 471248 487000 471368 0 FreeSans 480 0 0 0 Tile_X11Y6_BEN_SRAM1
port 1727 nsew signal output
flabel metal3 s 486200 467848 487000 467968 0 FreeSans 480 0 0 0 Tile_X11Y6_BEN_SRAM10
port 1728 nsew signal output
flabel metal3 s 486200 467168 487000 467288 0 FreeSans 480 0 0 0 Tile_X11Y6_BEN_SRAM11
port 1729 nsew signal output
flabel metal3 s 486200 503208 487000 503328 0 FreeSans 480 0 0 0 Tile_X11Y6_BEN_SRAM12
port 1730 nsew signal output
flabel metal3 s 486200 503888 487000 504008 0 FreeSans 480 0 0 0 Tile_X11Y6_BEN_SRAM13
port 1731 nsew signal output
flabel metal3 s 486200 539928 487000 540048 0 FreeSans 480 0 0 0 Tile_X11Y6_BEN_SRAM14
port 1732 nsew signal output
flabel metal3 s 486200 539248 487000 539368 0 FreeSans 480 0 0 0 Tile_X11Y6_BEN_SRAM15
port 1733 nsew signal output
flabel metal3 s 486200 504568 487000 504688 0 FreeSans 480 0 0 0 Tile_X11Y6_BEN_SRAM16
port 1734 nsew signal output
flabel metal3 s 486200 538568 487000 538688 0 FreeSans 480 0 0 0 Tile_X11Y6_BEN_SRAM17
port 1735 nsew signal output
flabel metal3 s 486200 505248 487000 505368 0 FreeSans 480 0 0 0 Tile_X11Y6_BEN_SRAM18
port 1736 nsew signal output
flabel metal3 s 486200 537888 487000 538008 0 FreeSans 480 0 0 0 Tile_X11Y6_BEN_SRAM19
port 1737 nsew signal output
flabel metal3 s 486200 500488 487000 500608 0 FreeSans 480 0 0 0 Tile_X11Y6_BEN_SRAM2
port 1738 nsew signal output
flabel metal3 s 486200 537208 487000 537328 0 FreeSans 480 0 0 0 Tile_X11Y6_BEN_SRAM20
port 1739 nsew signal output
flabel metal3 s 486200 505928 487000 506048 0 FreeSans 480 0 0 0 Tile_X11Y6_BEN_SRAM21
port 1740 nsew signal output
flabel metal3 s 486200 536528 487000 536648 0 FreeSans 480 0 0 0 Tile_X11Y6_BEN_SRAM22
port 1741 nsew signal output
flabel metal3 s 486200 506608 487000 506728 0 FreeSans 480 0 0 0 Tile_X11Y6_BEN_SRAM23
port 1742 nsew signal output
flabel metal3 s 486200 535848 487000 535968 0 FreeSans 480 0 0 0 Tile_X11Y6_BEN_SRAM24
port 1743 nsew signal output
flabel metal3 s 486200 535168 487000 535288 0 FreeSans 480 0 0 0 Tile_X11Y6_BEN_SRAM25
port 1744 nsew signal output
flabel metal3 s 486200 507288 487000 507408 0 FreeSans 480 0 0 0 Tile_X11Y6_BEN_SRAM26
port 1745 nsew signal output
flabel metal3 s 486200 534488 487000 534608 0 FreeSans 480 0 0 0 Tile_X11Y6_BEN_SRAM27
port 1746 nsew signal output
flabel metal3 s 486200 507968 487000 508088 0 FreeSans 480 0 0 0 Tile_X11Y6_BEN_SRAM28
port 1747 nsew signal output
flabel metal3 s 486200 533808 487000 533928 0 FreeSans 480 0 0 0 Tile_X11Y6_BEN_SRAM29
port 1748 nsew signal output
flabel metal3 s 486200 470568 487000 470688 0 FreeSans 480 0 0 0 Tile_X11Y6_BEN_SRAM3
port 1749 nsew signal output
flabel metal3 s 486200 533128 487000 533248 0 FreeSans 480 0 0 0 Tile_X11Y6_BEN_SRAM30
port 1750 nsew signal output
flabel metal3 s 486200 508648 487000 508768 0 FreeSans 480 0 0 0 Tile_X11Y6_BEN_SRAM31
port 1751 nsew signal output
flabel metal3 s 486200 501168 487000 501288 0 FreeSans 480 0 0 0 Tile_X11Y6_BEN_SRAM4
port 1752 nsew signal output
flabel metal3 s 486200 469888 487000 470008 0 FreeSans 480 0 0 0 Tile_X11Y6_BEN_SRAM5
port 1753 nsew signal output
flabel metal3 s 486200 469208 487000 469328 0 FreeSans 480 0 0 0 Tile_X11Y6_BEN_SRAM6
port 1754 nsew signal output
flabel metal3 s 486200 501848 487000 501968 0 FreeSans 480 0 0 0 Tile_X11Y6_BEN_SRAM7
port 1755 nsew signal output
flabel metal3 s 486200 468528 487000 468648 0 FreeSans 480 0 0 0 Tile_X11Y6_BEN_SRAM8
port 1756 nsew signal output
flabel metal3 s 486200 502528 487000 502648 0 FreeSans 480 0 0 0 Tile_X11Y6_BEN_SRAM9
port 1757 nsew signal output
flabel metal3 s 486200 532448 487000 532568 0 FreeSans 480 0 0 0 Tile_X11Y6_CLOCK_SRAM
port 1758 nsew signal output
flabel metal3 s 486200 509328 487000 509448 0 FreeSans 480 0 0 0 Tile_X11Y6_DI_SRAM0
port 1759 nsew signal output
flabel metal3 s 486200 531768 487000 531888 0 FreeSans 480 0 0 0 Tile_X11Y6_DI_SRAM1
port 1760 nsew signal output
flabel metal3 s 486200 531088 487000 531208 0 FreeSans 480 0 0 0 Tile_X11Y6_DI_SRAM10
port 1761 nsew signal output
flabel metal3 s 486200 527688 487000 527808 0 FreeSans 480 0 0 0 Tile_X11Y6_DI_SRAM11
port 1762 nsew signal output
flabel metal3 s 486200 527008 487000 527128 0 FreeSans 480 0 0 0 Tile_X11Y6_DI_SRAM12
port 1763 nsew signal output
flabel metal3 s 486200 514088 487000 514208 0 FreeSans 480 0 0 0 Tile_X11Y6_DI_SRAM13
port 1764 nsew signal output
flabel metal3 s 486200 526328 487000 526448 0 FreeSans 480 0 0 0 Tile_X11Y6_DI_SRAM14
port 1765 nsew signal output
flabel metal3 s 486200 518168 487000 518288 0 FreeSans 480 0 0 0 Tile_X11Y6_DI_SRAM15
port 1766 nsew signal output
flabel metal3 s 486200 529048 487000 529168 0 FreeSans 480 0 0 0 Tile_X11Y6_DI_SRAM16
port 1767 nsew signal output
flabel metal3 s 486200 524968 487000 525088 0 FreeSans 480 0 0 0 Tile_X11Y6_DI_SRAM17
port 1768 nsew signal output
flabel metal3 s 486200 515448 487000 515568 0 FreeSans 480 0 0 0 Tile_X11Y6_DI_SRAM18
port 1769 nsew signal output
flabel metal3 s 486200 524288 487000 524408 0 FreeSans 480 0 0 0 Tile_X11Y6_DI_SRAM19
port 1770 nsew signal output
flabel metal3 s 486200 510008 487000 510128 0 FreeSans 480 0 0 0 Tile_X11Y6_DI_SRAM2
port 1771 nsew signal output
flabel metal3 s 486200 514768 487000 514888 0 FreeSans 480 0 0 0 Tile_X11Y6_DI_SRAM20
port 1772 nsew signal output
flabel metal3 s 486200 523608 487000 523728 0 FreeSans 480 0 0 0 Tile_X11Y6_DI_SRAM21
port 1773 nsew signal output
flabel metal3 s 486200 522928 487000 523048 0 FreeSans 480 0 0 0 Tile_X11Y6_DI_SRAM22
port 1774 nsew signal output
flabel metal3 s 486200 518848 487000 518968 0 FreeSans 480 0 0 0 Tile_X11Y6_DI_SRAM23
port 1775 nsew signal output
flabel metal3 s 486200 528368 487000 528488 0 FreeSans 480 0 0 0 Tile_X11Y6_DI_SRAM24
port 1776 nsew signal output
flabel metal3 s 486200 516128 487000 516248 0 FreeSans 480 0 0 0 Tile_X11Y6_DI_SRAM25
port 1777 nsew signal output
flabel metal3 s 486200 530408 487000 530528 0 FreeSans 480 0 0 0 Tile_X11Y6_DI_SRAM26
port 1778 nsew signal output
flabel metal3 s 486200 520888 487000 521008 0 FreeSans 480 0 0 0 Tile_X11Y6_DI_SRAM27
port 1779 nsew signal output
flabel metal3 s 486200 522248 487000 522368 0 FreeSans 480 0 0 0 Tile_X11Y6_DI_SRAM28
port 1780 nsew signal output
flabel metal3 s 486200 520208 487000 520328 0 FreeSans 480 0 0 0 Tile_X11Y6_DI_SRAM29
port 1781 nsew signal output
flabel metal3 s 486200 511368 487000 511488 0 FreeSans 480 0 0 0 Tile_X11Y6_DI_SRAM3
port 1782 nsew signal output
flabel metal3 s 486200 517488 487000 517608 0 FreeSans 480 0 0 0 Tile_X11Y6_DI_SRAM30
port 1783 nsew signal output
flabel metal3 s 486200 519528 487000 519648 0 FreeSans 480 0 0 0 Tile_X11Y6_DI_SRAM31
port 1784 nsew signal output
flabel metal3 s 486200 510688 487000 510808 0 FreeSans 480 0 0 0 Tile_X11Y6_DI_SRAM4
port 1785 nsew signal output
flabel metal3 s 486200 512728 487000 512848 0 FreeSans 480 0 0 0 Tile_X11Y6_DI_SRAM5
port 1786 nsew signal output
flabel metal3 s 486200 513408 487000 513528 0 FreeSans 480 0 0 0 Tile_X11Y6_DI_SRAM6
port 1787 nsew signal output
flabel metal3 s 486200 512048 487000 512168 0 FreeSans 480 0 0 0 Tile_X11Y6_DI_SRAM7
port 1788 nsew signal output
flabel metal3 s 486200 521568 487000 521688 0 FreeSans 480 0 0 0 Tile_X11Y6_DI_SRAM8
port 1789 nsew signal output
flabel metal3 s 486200 516808 487000 516928 0 FreeSans 480 0 0 0 Tile_X11Y6_DI_SRAM9
port 1790 nsew signal output
flabel metal3 s 486200 476008 487000 476128 0 FreeSans 480 0 0 0 Tile_X11Y6_DO_SRAM0
port 1791 nsew signal input
flabel metal3 s 486200 488928 487000 489048 0 FreeSans 480 0 0 0 Tile_X11Y6_DO_SRAM1
port 1792 nsew signal input
flabel metal3 s 486200 484848 487000 484968 0 FreeSans 480 0 0 0 Tile_X11Y6_DO_SRAM10
port 1793 nsew signal input
flabel metal3 s 486200 491648 487000 491768 0 FreeSans 480 0 0 0 Tile_X11Y6_DO_SRAM11
port 1794 nsew signal input
flabel metal3 s 486200 484168 487000 484288 0 FreeSans 480 0 0 0 Tile_X11Y6_DO_SRAM12
port 1795 nsew signal input
flabel metal3 s 486200 483488 487000 483608 0 FreeSans 480 0 0 0 Tile_X11Y6_DO_SRAM13
port 1796 nsew signal input
flabel metal3 s 486200 492328 487000 492448 0 FreeSans 480 0 0 0 Tile_X11Y6_DO_SRAM14
port 1797 nsew signal input
flabel metal3 s 486200 482808 487000 482928 0 FreeSans 480 0 0 0 Tile_X11Y6_DO_SRAM15
port 1798 nsew signal input
flabel metal3 s 486200 493008 487000 493128 0 FreeSans 480 0 0 0 Tile_X11Y6_DO_SRAM16
port 1799 nsew signal input
flabel metal3 s 486200 482128 487000 482248 0 FreeSans 480 0 0 0 Tile_X11Y6_DO_SRAM17
port 1800 nsew signal input
flabel metal3 s 486200 481448 487000 481568 0 FreeSans 480 0 0 0 Tile_X11Y6_DO_SRAM18
port 1801 nsew signal input
flabel metal3 s 486200 493688 487000 493808 0 FreeSans 480 0 0 0 Tile_X11Y6_DO_SRAM19
port 1802 nsew signal input
flabel metal3 s 486200 488248 487000 488368 0 FreeSans 480 0 0 0 Tile_X11Y6_DO_SRAM2
port 1803 nsew signal input
flabel metal3 s 486200 480768 487000 480888 0 FreeSans 480 0 0 0 Tile_X11Y6_DO_SRAM20
port 1804 nsew signal input
flabel metal3 s 486200 494368 487000 494488 0 FreeSans 480 0 0 0 Tile_X11Y6_DO_SRAM21
port 1805 nsew signal input
flabel metal3 s 486200 480088 487000 480208 0 FreeSans 480 0 0 0 Tile_X11Y6_DO_SRAM22
port 1806 nsew signal input
flabel metal3 s 486200 479408 487000 479528 0 FreeSans 480 0 0 0 Tile_X11Y6_DO_SRAM23
port 1807 nsew signal input
flabel metal3 s 486200 495048 487000 495168 0 FreeSans 480 0 0 0 Tile_X11Y6_DO_SRAM24
port 1808 nsew signal input
flabel metal3 s 486200 478728 487000 478848 0 FreeSans 480 0 0 0 Tile_X11Y6_DO_SRAM25
port 1809 nsew signal input
flabel metal3 s 486200 495728 487000 495848 0 FreeSans 480 0 0 0 Tile_X11Y6_DO_SRAM26
port 1810 nsew signal input
flabel metal3 s 486200 478048 487000 478168 0 FreeSans 480 0 0 0 Tile_X11Y6_DO_SRAM27
port 1811 nsew signal input
flabel metal3 s 486200 477368 487000 477488 0 FreeSans 480 0 0 0 Tile_X11Y6_DO_SRAM28
port 1812 nsew signal input
flabel metal3 s 486200 496408 487000 496528 0 FreeSans 480 0 0 0 Tile_X11Y6_DO_SRAM29
port 1813 nsew signal input
flabel metal3 s 486200 487568 487000 487688 0 FreeSans 480 0 0 0 Tile_X11Y6_DO_SRAM3
port 1814 nsew signal input
flabel metal3 s 486200 476688 487000 476808 0 FreeSans 480 0 0 0 Tile_X11Y6_DO_SRAM30
port 1815 nsew signal input
flabel metal3 s 486200 497088 487000 497208 0 FreeSans 480 0 0 0 Tile_X11Y6_DO_SRAM31
port 1816 nsew signal input
flabel metal3 s 486200 489608 487000 489728 0 FreeSans 480 0 0 0 Tile_X11Y6_DO_SRAM4
port 1817 nsew signal input
flabel metal3 s 486200 486888 487000 487008 0 FreeSans 480 0 0 0 Tile_X11Y6_DO_SRAM5
port 1818 nsew signal input
flabel metal3 s 486200 490288 487000 490408 0 FreeSans 480 0 0 0 Tile_X11Y6_DO_SRAM6
port 1819 nsew signal input
flabel metal3 s 486200 486208 487000 486328 0 FreeSans 480 0 0 0 Tile_X11Y6_DO_SRAM7
port 1820 nsew signal input
flabel metal3 s 486200 485528 487000 485648 0 FreeSans 480 0 0 0 Tile_X11Y6_DO_SRAM8
port 1821 nsew signal input
flabel metal3 s 486200 490968 487000 491088 0 FreeSans 480 0 0 0 Tile_X11Y6_DO_SRAM9
port 1822 nsew signal input
flabel metal3 s 486200 525648 487000 525768 0 FreeSans 480 0 0 0 Tile_X11Y6_EN_SRAM
port 1823 nsew signal output
flabel metal3 s 486200 529728 487000 529848 0 FreeSans 480 0 0 0 Tile_X11Y6_R_WB_SRAM
port 1824 nsew signal output
flabel metal3 s 486200 459688 487000 459808 0 FreeSans 480 0 0 0 Tile_X11Y8_AD_SRAM0
port 1825 nsew signal output
flabel metal3 s 486200 408688 487000 408808 0 FreeSans 480 0 0 0 Tile_X11Y8_AD_SRAM1
port 1826 nsew signal output
flabel metal3 s 486200 408008 487000 408128 0 FreeSans 480 0 0 0 Tile_X11Y8_AD_SRAM2
port 1827 nsew signal output
flabel metal3 s 486200 458328 487000 458448 0 FreeSans 480 0 0 0 Tile_X11Y8_AD_SRAM3
port 1828 nsew signal output
flabel metal3 s 486200 410048 487000 410168 0 FreeSans 480 0 0 0 Tile_X11Y8_AD_SRAM4
port 1829 nsew signal output
flabel metal3 s 486200 457648 487000 457768 0 FreeSans 480 0 0 0 Tile_X11Y8_AD_SRAM5
port 1830 nsew signal output
flabel metal3 s 486200 456968 487000 457088 0 FreeSans 480 0 0 0 Tile_X11Y8_AD_SRAM6
port 1831 nsew signal output
flabel metal3 s 486200 409368 487000 409488 0 FreeSans 480 0 0 0 Tile_X11Y8_AD_SRAM7
port 1832 nsew signal output
flabel metal3 s 486200 456288 487000 456408 0 FreeSans 480 0 0 0 Tile_X11Y8_AD_SRAM8
port 1833 nsew signal output
flabel metal3 s 486200 411408 487000 411528 0 FreeSans 480 0 0 0 Tile_X11Y8_AD_SRAM9
port 1834 nsew signal output
flabel metal3 s 486200 455608 487000 455728 0 FreeSans 480 0 0 0 Tile_X11Y8_BEN_SRAM0
port 1835 nsew signal output
flabel metal3 s 486200 454928 487000 455048 0 FreeSans 480 0 0 0 Tile_X11Y8_BEN_SRAM1
port 1836 nsew signal output
flabel metal3 s 486200 454248 487000 454368 0 FreeSans 480 0 0 0 Tile_X11Y8_BEN_SRAM10
port 1837 nsew signal output
flabel metal3 s 486200 450848 487000 450968 0 FreeSans 480 0 0 0 Tile_X11Y8_BEN_SRAM11
port 1838 nsew signal output
flabel metal3 s 486200 419568 487000 419688 0 FreeSans 480 0 0 0 Tile_X11Y8_BEN_SRAM12
port 1839 nsew signal output
flabel metal3 s 486200 450168 487000 450288 0 FreeSans 480 0 0 0 Tile_X11Y8_BEN_SRAM13
port 1840 nsew signal output
flabel metal3 s 486200 416168 487000 416288 0 FreeSans 480 0 0 0 Tile_X11Y8_BEN_SRAM14
port 1841 nsew signal output
flabel metal3 s 486200 449488 487000 449608 0 FreeSans 480 0 0 0 Tile_X11Y8_BEN_SRAM15
port 1842 nsew signal output
flabel metal3 s 486200 448808 487000 448928 0 FreeSans 480 0 0 0 Tile_X11Y8_BEN_SRAM16
port 1843 nsew signal output
flabel metal3 s 486200 414808 487000 414928 0 FreeSans 480 0 0 0 Tile_X11Y8_BEN_SRAM17
port 1844 nsew signal output
flabel metal3 s 486200 448128 487000 448248 0 FreeSans 480 0 0 0 Tile_X11Y8_BEN_SRAM18
port 1845 nsew signal output
flabel metal3 s 486200 416848 487000 416968 0 FreeSans 480 0 0 0 Tile_X11Y8_BEN_SRAM19
port 1846 nsew signal output
flabel metal3 s 486200 410728 487000 410848 0 FreeSans 480 0 0 0 Tile_X11Y8_BEN_SRAM2
port 1847 nsew signal output
flabel metal3 s 486200 447448 487000 447568 0 FreeSans 480 0 0 0 Tile_X11Y8_BEN_SRAM20
port 1848 nsew signal output
flabel metal3 s 486200 446768 487000 446888 0 FreeSans 480 0 0 0 Tile_X11Y8_BEN_SRAM21
port 1849 nsew signal output
flabel metal3 s 486200 438608 487000 438728 0 FreeSans 480 0 0 0 Tile_X11Y8_BEN_SRAM22
port 1850 nsew signal output
flabel metal3 s 486200 446088 487000 446208 0 FreeSans 480 0 0 0 Tile_X11Y8_BEN_SRAM23
port 1851 nsew signal output
flabel metal3 s 486200 418208 487000 418328 0 FreeSans 480 0 0 0 Tile_X11Y8_BEN_SRAM24
port 1852 nsew signal output
flabel metal3 s 486200 445408 487000 445528 0 FreeSans 480 0 0 0 Tile_X11Y8_BEN_SRAM25
port 1853 nsew signal output
flabel metal3 s 486200 444728 487000 444848 0 FreeSans 480 0 0 0 Tile_X11Y8_BEN_SRAM26
port 1854 nsew signal output
flabel metal3 s 486200 417528 487000 417648 0 FreeSans 480 0 0 0 Tile_X11Y8_BEN_SRAM27
port 1855 nsew signal output
flabel metal3 s 486200 444048 487000 444168 0 FreeSans 480 0 0 0 Tile_X11Y8_BEN_SRAM28
port 1856 nsew signal output
flabel metal3 s 486200 459008 487000 459128 0 FreeSans 480 0 0 0 Tile_X11Y8_BEN_SRAM29
port 1857 nsew signal output
flabel metal3 s 486200 412088 487000 412208 0 FreeSans 480 0 0 0 Tile_X11Y8_BEN_SRAM3
port 1858 nsew signal output
flabel metal3 s 486200 443368 487000 443488 0 FreeSans 480 0 0 0 Tile_X11Y8_BEN_SRAM30
port 1859 nsew signal output
flabel metal3 s 486200 442688 487000 442808 0 FreeSans 480 0 0 0 Tile_X11Y8_BEN_SRAM31
port 1860 nsew signal output
flabel metal3 s 486200 413448 487000 413568 0 FreeSans 480 0 0 0 Tile_X11Y8_BEN_SRAM4
port 1861 nsew signal output
flabel metal3 s 486200 414128 487000 414248 0 FreeSans 480 0 0 0 Tile_X11Y8_BEN_SRAM5
port 1862 nsew signal output
flabel metal3 s 486200 412768 487000 412888 0 FreeSans 480 0 0 0 Tile_X11Y8_BEN_SRAM6
port 1863 nsew signal output
flabel metal3 s 486200 422968 487000 423088 0 FreeSans 480 0 0 0 Tile_X11Y8_BEN_SRAM7
port 1864 nsew signal output
flabel metal3 s 486200 420248 487000 420368 0 FreeSans 480 0 0 0 Tile_X11Y8_BEN_SRAM8
port 1865 nsew signal output
flabel metal3 s 486200 415488 487000 415608 0 FreeSans 480 0 0 0 Tile_X11Y8_BEN_SRAM9
port 1866 nsew signal output
flabel metal3 s 486200 418888 487000 419008 0 FreeSans 480 0 0 0 Tile_X11Y8_CLOCK_SRAM
port 1867 nsew signal output
flabel metal3 s 486200 442008 487000 442128 0 FreeSans 480 0 0 0 Tile_X11Y8_DI_SRAM0
port 1868 nsew signal output
flabel metal3 s 486200 423648 487000 423768 0 FreeSans 480 0 0 0 Tile_X11Y8_DI_SRAM1
port 1869 nsew signal output
flabel metal3 s 486200 441328 487000 441448 0 FreeSans 480 0 0 0 Tile_X11Y8_DI_SRAM10
port 1870 nsew signal output
flabel metal3 s 486200 424328 487000 424448 0 FreeSans 480 0 0 0 Tile_X11Y8_DI_SRAM11
port 1871 nsew signal output
flabel metal3 s 486200 437248 487000 437368 0 FreeSans 480 0 0 0 Tile_X11Y8_DI_SRAM12
port 1872 nsew signal output
flabel metal3 s 486200 436568 487000 436688 0 FreeSans 480 0 0 0 Tile_X11Y8_DI_SRAM13
port 1873 nsew signal output
flabel metal3 s 486200 429088 487000 429208 0 FreeSans 480 0 0 0 Tile_X11Y8_DI_SRAM14
port 1874 nsew signal output
flabel metal3 s 486200 435888 487000 436008 0 FreeSans 480 0 0 0 Tile_X11Y8_DI_SRAM15
port 1875 nsew signal output
flabel metal3 s 486200 425008 487000 425128 0 FreeSans 480 0 0 0 Tile_X11Y8_DI_SRAM16
port 1876 nsew signal output
flabel metal3 s 486200 435208 487000 435328 0 FreeSans 480 0 0 0 Tile_X11Y8_DI_SRAM17
port 1877 nsew signal output
flabel metal3 s 486200 453568 487000 453688 0 FreeSans 480 0 0 0 Tile_X11Y8_DI_SRAM18
port 1878 nsew signal output
flabel metal3 s 486200 425688 487000 425808 0 FreeSans 480 0 0 0 Tile_X11Y8_DI_SRAM19
port 1879 nsew signal output
flabel metal3 s 486200 428408 487000 428528 0 FreeSans 480 0 0 0 Tile_X11Y8_DI_SRAM2
port 1880 nsew signal output
flabel metal3 s 486200 452888 487000 453008 0 FreeSans 480 0 0 0 Tile_X11Y8_DI_SRAM20
port 1881 nsew signal output
flabel metal3 s 486200 437928 487000 438048 0 FreeSans 480 0 0 0 Tile_X11Y8_DI_SRAM21
port 1882 nsew signal output
flabel metal3 s 486200 433168 487000 433288 0 FreeSans 480 0 0 0 Tile_X11Y8_DI_SRAM22
port 1883 nsew signal output
flabel metal3 s 486200 432488 487000 432608 0 FreeSans 480 0 0 0 Tile_X11Y8_DI_SRAM23
port 1884 nsew signal output
flabel metal3 s 486200 439968 487000 440088 0 FreeSans 480 0 0 0 Tile_X11Y8_DI_SRAM24
port 1885 nsew signal output
flabel metal3 s 486200 431808 487000 431928 0 FreeSans 480 0 0 0 Tile_X11Y8_DI_SRAM25
port 1886 nsew signal output
flabel metal3 s 486200 426368 487000 426488 0 FreeSans 480 0 0 0 Tile_X11Y8_DI_SRAM26
port 1887 nsew signal output
flabel metal3 s 486200 431128 487000 431248 0 FreeSans 480 0 0 0 Tile_X11Y8_DI_SRAM27
port 1888 nsew signal output
flabel metal3 s 486200 430448 487000 430568 0 FreeSans 480 0 0 0 Tile_X11Y8_DI_SRAM28
port 1889 nsew signal output
flabel metal3 s 486200 427048 487000 427168 0 FreeSans 480 0 0 0 Tile_X11Y8_DI_SRAM29
port 1890 nsew signal output
flabel metal3 s 486200 452208 487000 452328 0 FreeSans 480 0 0 0 Tile_X11Y8_DI_SRAM3
port 1891 nsew signal output
flabel metal3 s 486200 429768 487000 429888 0 FreeSans 480 0 0 0 Tile_X11Y8_DI_SRAM30
port 1892 nsew signal output
flabel metal3 s 486200 427728 487000 427848 0 FreeSans 480 0 0 0 Tile_X11Y8_DI_SRAM31
port 1893 nsew signal output
flabel metal3 s 486200 440648 487000 440768 0 FreeSans 480 0 0 0 Tile_X11Y8_DI_SRAM4
port 1894 nsew signal output
flabel metal3 s 486200 420928 487000 421048 0 FreeSans 480 0 0 0 Tile_X11Y8_DI_SRAM5
port 1895 nsew signal output
flabel metal3 s 486200 421608 487000 421728 0 FreeSans 480 0 0 0 Tile_X11Y8_DI_SRAM6
port 1896 nsew signal output
flabel metal3 s 486200 422288 487000 422408 0 FreeSans 480 0 0 0 Tile_X11Y8_DI_SRAM7
port 1897 nsew signal output
flabel metal3 s 486200 451528 487000 451648 0 FreeSans 480 0 0 0 Tile_X11Y8_DI_SRAM8
port 1898 nsew signal output
flabel metal3 s 486200 433848 487000 433968 0 FreeSans 480 0 0 0 Tile_X11Y8_DI_SRAM9
port 1899 nsew signal output
flabel metal3 s 486200 386248 487000 386368 0 FreeSans 480 0 0 0 Tile_X11Y8_DO_SRAM0
port 1900 nsew signal input
flabel metal3 s 486200 398488 487000 398608 0 FreeSans 480 0 0 0 Tile_X11Y8_DO_SRAM1
port 1901 nsew signal input
flabel metal3 s 486200 401208 487000 401328 0 FreeSans 480 0 0 0 Tile_X11Y8_DO_SRAM10
port 1902 nsew signal input
flabel metal3 s 486200 394408 487000 394528 0 FreeSans 480 0 0 0 Tile_X11Y8_DO_SRAM11
port 1903 nsew signal input
flabel metal3 s 486200 401888 487000 402008 0 FreeSans 480 0 0 0 Tile_X11Y8_DO_SRAM12
port 1904 nsew signal input
flabel metal3 s 486200 393728 487000 393848 0 FreeSans 480 0 0 0 Tile_X11Y8_DO_SRAM13
port 1905 nsew signal input
flabel metal3 s 486200 393048 487000 393168 0 FreeSans 480 0 0 0 Tile_X11Y8_DO_SRAM14
port 1906 nsew signal input
flabel metal3 s 486200 402568 487000 402688 0 FreeSans 480 0 0 0 Tile_X11Y8_DO_SRAM15
port 1907 nsew signal input
flabel metal3 s 486200 392368 487000 392488 0 FreeSans 480 0 0 0 Tile_X11Y8_DO_SRAM16
port 1908 nsew signal input
flabel metal3 s 486200 403248 487000 403368 0 FreeSans 480 0 0 0 Tile_X11Y8_DO_SRAM17
port 1909 nsew signal input
flabel metal3 s 486200 391688 487000 391808 0 FreeSans 480 0 0 0 Tile_X11Y8_DO_SRAM18
port 1910 nsew signal input
flabel metal3 s 486200 391008 487000 391128 0 FreeSans 480 0 0 0 Tile_X11Y8_DO_SRAM19
port 1911 nsew signal input
flabel metal3 s 486200 399168 487000 399288 0 FreeSans 480 0 0 0 Tile_X11Y8_DO_SRAM2
port 1912 nsew signal input
flabel metal3 s 486200 403928 487000 404048 0 FreeSans 480 0 0 0 Tile_X11Y8_DO_SRAM20
port 1913 nsew signal input
flabel metal3 s 486200 390328 487000 390448 0 FreeSans 480 0 0 0 Tile_X11Y8_DO_SRAM21
port 1914 nsew signal input
flabel metal3 s 486200 404608 487000 404728 0 FreeSans 480 0 0 0 Tile_X11Y8_DO_SRAM22
port 1915 nsew signal input
flabel metal3 s 486200 389648 487000 389768 0 FreeSans 480 0 0 0 Tile_X11Y8_DO_SRAM23
port 1916 nsew signal input
flabel metal3 s 486200 388968 487000 389088 0 FreeSans 480 0 0 0 Tile_X11Y8_DO_SRAM24
port 1917 nsew signal input
flabel metal3 s 486200 405288 487000 405408 0 FreeSans 480 0 0 0 Tile_X11Y8_DO_SRAM25
port 1918 nsew signal input
flabel metal3 s 486200 388288 487000 388408 0 FreeSans 480 0 0 0 Tile_X11Y8_DO_SRAM26
port 1919 nsew signal input
flabel metal3 s 486200 405968 487000 406088 0 FreeSans 480 0 0 0 Tile_X11Y8_DO_SRAM27
port 1920 nsew signal input
flabel metal3 s 486200 387608 487000 387728 0 FreeSans 480 0 0 0 Tile_X11Y8_DO_SRAM28
port 1921 nsew signal input
flabel metal3 s 486200 386928 487000 387048 0 FreeSans 480 0 0 0 Tile_X11Y8_DO_SRAM29
port 1922 nsew signal input
flabel metal3 s 486200 397808 487000 397928 0 FreeSans 480 0 0 0 Tile_X11Y8_DO_SRAM3
port 1923 nsew signal input
flabel metal3 s 486200 406648 487000 406768 0 FreeSans 480 0 0 0 Tile_X11Y8_DO_SRAM30
port 1924 nsew signal input
flabel metal3 s 486200 407328 487000 407448 0 FreeSans 480 0 0 0 Tile_X11Y8_DO_SRAM31
port 1925 nsew signal input
flabel metal3 s 486200 397128 487000 397248 0 FreeSans 480 0 0 0 Tile_X11Y8_DO_SRAM4
port 1926 nsew signal input
flabel metal3 s 486200 399848 487000 399968 0 FreeSans 480 0 0 0 Tile_X11Y8_DO_SRAM5
port 1927 nsew signal input
flabel metal3 s 486200 396448 487000 396568 0 FreeSans 480 0 0 0 Tile_X11Y8_DO_SRAM6
port 1928 nsew signal input
flabel metal3 s 486200 400528 487000 400648 0 FreeSans 480 0 0 0 Tile_X11Y8_DO_SRAM7
port 1929 nsew signal input
flabel metal3 s 486200 395768 487000 395888 0 FreeSans 480 0 0 0 Tile_X11Y8_DO_SRAM8
port 1930 nsew signal input
flabel metal3 s 486200 395088 487000 395208 0 FreeSans 480 0 0 0 Tile_X11Y8_DO_SRAM9
port 1931 nsew signal input
flabel metal3 s 486200 439288 487000 439408 0 FreeSans 480 0 0 0 Tile_X11Y8_EN_SRAM
port 1932 nsew signal output
flabel metal3 s 486200 434528 487000 434648 0 FreeSans 480 0 0 0 Tile_X11Y8_R_WB_SRAM
port 1933 nsew signal output
flabel metal2 s 24490 755700 24546 756500 0 FreeSans 224 90 0 0 Tile_X1Y0_A_I_top
port 1934 nsew signal output
flabel metal2 s 23202 755700 23258 756500 0 FreeSans 224 90 0 0 Tile_X1Y0_A_O_top
port 1935 nsew signal input
flabel metal2 s 25134 755700 25190 756500 0 FreeSans 224 90 0 0 Tile_X1Y0_A_T_top
port 1936 nsew signal output
flabel metal2 s 29642 755700 29698 756500 0 FreeSans 224 90 0 0 Tile_X1Y0_A_config_C_bit0
port 1937 nsew signal output
flabel metal2 s 30930 755700 30986 756500 0 FreeSans 224 90 0 0 Tile_X1Y0_A_config_C_bit1
port 1938 nsew signal output
flabel metal2 s 32218 755700 32274 756500 0 FreeSans 224 90 0 0 Tile_X1Y0_A_config_C_bit2
port 1939 nsew signal output
flabel metal2 s 32862 755700 32918 756500 0 FreeSans 224 90 0 0 Tile_X1Y0_A_config_C_bit3
port 1940 nsew signal output
flabel metal2 s 27710 755700 27766 756500 0 FreeSans 224 90 0 0 Tile_X1Y0_B_I_top
port 1941 nsew signal output
flabel metal2 s 26422 755700 26478 756500 0 FreeSans 224 90 0 0 Tile_X1Y0_B_O_top
port 1942 nsew signal input
flabel metal2 s 28998 755700 29054 756500 0 FreeSans 224 90 0 0 Tile_X1Y0_B_T_top
port 1943 nsew signal output
flabel metal2 s 34150 755700 34206 756500 0 FreeSans 224 90 0 0 Tile_X1Y0_B_config_C_bit0
port 1944 nsew signal output
flabel metal2 s 35438 755700 35494 756500 0 FreeSans 224 90 0 0 Tile_X1Y0_B_config_C_bit1
port 1945 nsew signal output
flabel metal2 s 36082 755700 36138 756500 0 FreeSans 224 90 0 0 Tile_X1Y0_B_config_C_bit2
port 1946 nsew signal output
flabel metal2 s 37370 755700 37426 756500 0 FreeSans 224 90 0 0 Tile_X1Y0_B_config_C_bit3
port 1947 nsew signal output
flabel metal2 s 23202 0 23258 800 0 FreeSans 224 90 0 0 Tile_X1Y17_IRQ_top0
port 1948 nsew signal output
flabel metal2 s 24490 0 24546 800 0 FreeSans 224 90 0 0 Tile_X1Y17_IRQ_top1
port 1949 nsew signal output
flabel metal2 s 25778 0 25834 800 0 FreeSans 224 90 0 0 Tile_X1Y17_IRQ_top2
port 1950 nsew signal output
flabel metal2 s 27710 0 27766 800 0 FreeSans 224 90 0 0 Tile_X1Y17_IRQ_top3
port 1951 nsew signal output
flabel metal2 s 65062 755700 65118 756500 0 FreeSans 224 90 0 0 Tile_X2Y0_A_I_top
port 1952 nsew signal output
flabel metal2 s 63774 755700 63830 756500 0 FreeSans 224 90 0 0 Tile_X2Y0_A_O_top
port 1953 nsew signal input
flabel metal2 s 66350 755700 66406 756500 0 FreeSans 224 90 0 0 Tile_X2Y0_A_T_top
port 1954 nsew signal output
flabel metal2 s 70858 755700 70914 756500 0 FreeSans 224 90 0 0 Tile_X2Y0_A_config_C_bit0
port 1955 nsew signal output
flabel metal2 s 71502 755700 71558 756500 0 FreeSans 224 90 0 0 Tile_X2Y0_A_config_C_bit1
port 1956 nsew signal output
flabel metal2 s 72790 755700 72846 756500 0 FreeSans 224 90 0 0 Tile_X2Y0_A_config_C_bit2
port 1957 nsew signal output
flabel metal2 s 74078 755700 74134 756500 0 FreeSans 224 90 0 0 Tile_X2Y0_A_config_C_bit3
port 1958 nsew signal output
flabel metal2 s 68282 755700 68338 756500 0 FreeSans 224 90 0 0 Tile_X2Y0_B_I_top
port 1959 nsew signal output
flabel metal2 s 66994 755700 67050 756500 0 FreeSans 224 90 0 0 Tile_X2Y0_B_O_top
port 1960 nsew signal input
flabel metal2 s 69570 755700 69626 756500 0 FreeSans 224 90 0 0 Tile_X2Y0_B_T_top
port 1961 nsew signal output
flabel metal2 s 74722 755700 74778 756500 0 FreeSans 224 90 0 0 Tile_X2Y0_B_config_C_bit0
port 1962 nsew signal output
flabel metal2 s 76010 755700 76066 756500 0 FreeSans 224 90 0 0 Tile_X2Y0_B_config_C_bit1
port 1963 nsew signal output
flabel metal2 s 77298 755700 77354 756500 0 FreeSans 224 90 0 0 Tile_X2Y0_B_config_C_bit2
port 1964 nsew signal output
flabel metal2 s 78586 755700 78642 756500 0 FreeSans 224 90 0 0 Tile_X2Y0_B_config_C_bit3
port 1965 nsew signal output
flabel metal2 s 65062 0 65118 800 0 FreeSans 224 90 0 0 Tile_X2Y17_BOOT_top
port 1966 nsew signal output
flabel metal2 s 63774 0 63830 800 0 FreeSans 224 90 0 0 Tile_X2Y17_RESET_top
port 1967 nsew signal input
flabel metal2 s 66350 0 66406 800 0 FreeSans 224 90 0 0 Tile_X2Y17_SLOT_top0
port 1968 nsew signal output
flabel metal2 s 68282 0 68338 800 0 FreeSans 224 90 0 0 Tile_X2Y17_SLOT_top1
port 1969 nsew signal output
flabel metal2 s 69570 0 69626 800 0 FreeSans 224 90 0 0 Tile_X2Y17_SLOT_top2
port 1970 nsew signal output
flabel metal2 s 70858 0 70914 800 0 FreeSans 224 90 0 0 Tile_X2Y17_SLOT_top3
port 1971 nsew signal output
flabel metal2 s 155222 755700 155278 756500 0 FreeSans 224 90 0 0 Tile_X4Y0_A_I_top
port 1972 nsew signal output
flabel metal2 s 153934 755700 153990 756500 0 FreeSans 224 90 0 0 Tile_X4Y0_A_O_top
port 1973 nsew signal input
flabel metal2 s 155866 755700 155922 756500 0 FreeSans 224 90 0 0 Tile_X4Y0_A_T_top
port 1974 nsew signal output
flabel metal2 s 160374 755700 160430 756500 0 FreeSans 224 90 0 0 Tile_X4Y0_A_config_C_bit0
port 1975 nsew signal output
flabel metal2 s 161662 755700 161718 756500 0 FreeSans 224 90 0 0 Tile_X4Y0_A_config_C_bit1
port 1976 nsew signal output
flabel metal2 s 162950 755700 163006 756500 0 FreeSans 224 90 0 0 Tile_X4Y0_A_config_C_bit2
port 1977 nsew signal output
flabel metal2 s 163594 755700 163650 756500 0 FreeSans 224 90 0 0 Tile_X4Y0_A_config_C_bit3
port 1978 nsew signal output
flabel metal2 s 158442 755700 158498 756500 0 FreeSans 224 90 0 0 Tile_X4Y0_B_I_top
port 1979 nsew signal output
flabel metal2 s 157154 755700 157210 756500 0 FreeSans 224 90 0 0 Tile_X4Y0_B_O_top
port 1980 nsew signal input
flabel metal2 s 159730 755700 159786 756500 0 FreeSans 224 90 0 0 Tile_X4Y0_B_T_top
port 1981 nsew signal output
flabel metal2 s 164882 755700 164938 756500 0 FreeSans 224 90 0 0 Tile_X4Y0_B_config_C_bit0
port 1982 nsew signal output
flabel metal2 s 166170 755700 166226 756500 0 FreeSans 224 90 0 0 Tile_X4Y0_B_config_C_bit1
port 1983 nsew signal output
flabel metal2 s 167458 755700 167514 756500 0 FreeSans 224 90 0 0 Tile_X4Y0_B_config_C_bit2
port 1984 nsew signal output
flabel metal2 s 168102 755700 168158 756500 0 FreeSans 224 90 0 0 Tile_X4Y0_B_config_C_bit3
port 1985 nsew signal output
flabel metal2 s 165526 0 165582 800 0 FreeSans 224 90 0 0 Tile_X4Y17_I_top0
port 1986 nsew signal output
flabel metal2 s 166170 0 166226 800 0 FreeSans 224 90 0 0 Tile_X4Y17_I_top1
port 1987 nsew signal output
flabel metal2 s 172610 0 172666 800 0 FreeSans 224 90 0 0 Tile_X4Y17_I_top10
port 1988 nsew signal output
flabel metal2 s 173254 0 173310 800 0 FreeSans 224 90 0 0 Tile_X4Y17_I_top11
port 1989 nsew signal output
flabel metal2 s 173898 0 173954 800 0 FreeSans 224 90 0 0 Tile_X4Y17_I_top12
port 1990 nsew signal output
flabel metal2 s 175186 0 175242 800 0 FreeSans 224 90 0 0 Tile_X4Y17_I_top13
port 1991 nsew signal output
flabel metal2 s 175830 0 175886 800 0 FreeSans 224 90 0 0 Tile_X4Y17_I_top14
port 1992 nsew signal output
flabel metal2 s 176474 0 176530 800 0 FreeSans 224 90 0 0 Tile_X4Y17_I_top15
port 1993 nsew signal output
flabel metal2 s 166814 0 166870 800 0 FreeSans 224 90 0 0 Tile_X4Y17_I_top2
port 1994 nsew signal output
flabel metal2 s 167458 0 167514 800 0 FreeSans 224 90 0 0 Tile_X4Y17_I_top3
port 1995 nsew signal output
flabel metal2 s 168102 0 168158 800 0 FreeSans 224 90 0 0 Tile_X4Y17_I_top4
port 1996 nsew signal output
flabel metal2 s 168746 0 168802 800 0 FreeSans 224 90 0 0 Tile_X4Y17_I_top5
port 1997 nsew signal output
flabel metal2 s 170034 0 170090 800 0 FreeSans 224 90 0 0 Tile_X4Y17_I_top6
port 1998 nsew signal output
flabel metal2 s 170678 0 170734 800 0 FreeSans 224 90 0 0 Tile_X4Y17_I_top7
port 1999 nsew signal output
flabel metal2 s 171322 0 171378 800 0 FreeSans 224 90 0 0 Tile_X4Y17_I_top8
port 2000 nsew signal output
flabel metal2 s 171966 0 172022 800 0 FreeSans 224 90 0 0 Tile_X4Y17_I_top9
port 2001 nsew signal output
flabel metal2 s 153290 0 153346 800 0 FreeSans 224 90 0 0 Tile_X4Y17_O_top0
port 2002 nsew signal input
flabel metal2 s 154578 0 154634 800 0 FreeSans 224 90 0 0 Tile_X4Y17_O_top1
port 2003 nsew signal input
flabel metal2 s 161018 0 161074 800 0 FreeSans 224 90 0 0 Tile_X4Y17_O_top10
port 2004 nsew signal input
flabel metal2 s 161662 0 161718 800 0 FreeSans 224 90 0 0 Tile_X4Y17_O_top11
port 2005 nsew signal input
flabel metal2 s 162306 0 162362 800 0 FreeSans 224 90 0 0 Tile_X4Y17_O_top12
port 2006 nsew signal input
flabel metal2 s 162950 0 163006 800 0 FreeSans 224 90 0 0 Tile_X4Y17_O_top13
port 2007 nsew signal input
flabel metal2 s 163594 0 163650 800 0 FreeSans 224 90 0 0 Tile_X4Y17_O_top14
port 2008 nsew signal input
flabel metal2 s 164882 0 164938 800 0 FreeSans 224 90 0 0 Tile_X4Y17_O_top15
port 2009 nsew signal input
flabel metal2 s 155222 0 155278 800 0 FreeSans 224 90 0 0 Tile_X4Y17_O_top2
port 2010 nsew signal input
flabel metal2 s 155866 0 155922 800 0 FreeSans 224 90 0 0 Tile_X4Y17_O_top3
port 2011 nsew signal input
flabel metal2 s 156510 0 156566 800 0 FreeSans 224 90 0 0 Tile_X4Y17_O_top4
port 2012 nsew signal input
flabel metal2 s 157154 0 157210 800 0 FreeSans 224 90 0 0 Tile_X4Y17_O_top5
port 2013 nsew signal input
flabel metal2 s 157798 0 157854 800 0 FreeSans 224 90 0 0 Tile_X4Y17_O_top6
port 2014 nsew signal input
flabel metal2 s 158442 0 158498 800 0 FreeSans 224 90 0 0 Tile_X4Y17_O_top7
port 2015 nsew signal input
flabel metal2 s 159730 0 159786 800 0 FreeSans 224 90 0 0 Tile_X4Y17_O_top8
port 2016 nsew signal input
flabel metal2 s 160374 0 160430 800 0 FreeSans 224 90 0 0 Tile_X4Y17_O_top9
port 2017 nsew signal input
flabel metal2 s 195794 755700 195850 756500 0 FreeSans 224 90 0 0 Tile_X5Y0_A_I_top
port 2018 nsew signal output
flabel metal2 s 195150 755700 195206 756500 0 FreeSans 224 90 0 0 Tile_X5Y0_A_O_top
port 2019 nsew signal input
flabel metal2 s 197082 755700 197138 756500 0 FreeSans 224 90 0 0 Tile_X5Y0_A_T_top
port 2020 nsew signal output
flabel metal2 s 201590 755700 201646 756500 0 FreeSans 224 90 0 0 Tile_X5Y0_A_config_C_bit0
port 2021 nsew signal output
flabel metal2 s 202878 755700 202934 756500 0 FreeSans 224 90 0 0 Tile_X5Y0_A_config_C_bit1
port 2022 nsew signal output
flabel metal2 s 203522 755700 203578 756500 0 FreeSans 224 90 0 0 Tile_X5Y0_A_config_C_bit2
port 2023 nsew signal output
flabel metal2 s 204810 755700 204866 756500 0 FreeSans 224 90 0 0 Tile_X5Y0_A_config_C_bit3
port 2024 nsew signal output
flabel metal2 s 199658 755700 199714 756500 0 FreeSans 224 90 0 0 Tile_X5Y0_B_I_top
port 2025 nsew signal output
flabel metal2 s 198370 755700 198426 756500 0 FreeSans 224 90 0 0 Tile_X5Y0_B_O_top
port 2026 nsew signal input
flabel metal2 s 200302 755700 200358 756500 0 FreeSans 224 90 0 0 Tile_X5Y0_B_T_top
port 2027 nsew signal output
flabel metal2 s 206098 755700 206154 756500 0 FreeSans 224 90 0 0 Tile_X5Y0_B_config_C_bit0
port 2028 nsew signal output
flabel metal2 s 207386 755700 207442 756500 0 FreeSans 224 90 0 0 Tile_X5Y0_B_config_C_bit1
port 2029 nsew signal output
flabel metal2 s 208030 755700 208086 756500 0 FreeSans 224 90 0 0 Tile_X5Y0_B_config_C_bit2
port 2030 nsew signal output
flabel metal2 s 209318 755700 209374 756500 0 FreeSans 224 90 0 0 Tile_X5Y0_B_config_C_bit3
port 2031 nsew signal output
flabel metal2 s 206098 0 206154 800 0 FreeSans 224 90 0 0 Tile_X5Y17_I_top0
port 2032 nsew signal output
flabel metal2 s 207386 0 207442 800 0 FreeSans 224 90 0 0 Tile_X5Y17_I_top1
port 2033 nsew signal output
flabel metal2 s 213826 0 213882 800 0 FreeSans 224 90 0 0 Tile_X5Y17_I_top10
port 2034 nsew signal output
flabel metal2 s 214470 0 214526 800 0 FreeSans 224 90 0 0 Tile_X5Y17_I_top11
port 2035 nsew signal output
flabel metal2 s 215114 0 215170 800 0 FreeSans 224 90 0 0 Tile_X5Y17_I_top12
port 2036 nsew signal output
flabel metal2 s 215758 0 215814 800 0 FreeSans 224 90 0 0 Tile_X5Y17_I_top13
port 2037 nsew signal output
flabel metal2 s 216402 0 216458 800 0 FreeSans 224 90 0 0 Tile_X5Y17_I_top14
port 2038 nsew signal output
flabel metal2 s 217690 0 217746 800 0 FreeSans 224 90 0 0 Tile_X5Y17_I_top15
port 2039 nsew signal output
flabel metal2 s 208030 0 208086 800 0 FreeSans 224 90 0 0 Tile_X5Y17_I_top2
port 2040 nsew signal output
flabel metal2 s 208674 0 208730 800 0 FreeSans 224 90 0 0 Tile_X5Y17_I_top3
port 2041 nsew signal output
flabel metal2 s 209318 0 209374 800 0 FreeSans 224 90 0 0 Tile_X5Y17_I_top4
port 2042 nsew signal output
flabel metal2 s 209962 0 210018 800 0 FreeSans 224 90 0 0 Tile_X5Y17_I_top5
port 2043 nsew signal output
flabel metal2 s 210606 0 210662 800 0 FreeSans 224 90 0 0 Tile_X5Y17_I_top6
port 2044 nsew signal output
flabel metal2 s 211250 0 211306 800 0 FreeSans 224 90 0 0 Tile_X5Y17_I_top7
port 2045 nsew signal output
flabel metal2 s 212538 0 212594 800 0 FreeSans 224 90 0 0 Tile_X5Y17_I_top8
port 2046 nsew signal output
flabel metal2 s 213182 0 213238 800 0 FreeSans 224 90 0 0 Tile_X5Y17_I_top9
port 2047 nsew signal output
flabel metal2 s 194506 0 194562 800 0 FreeSans 224 90 0 0 Tile_X5Y17_O_top0
port 2048 nsew signal input
flabel metal2 s 195150 0 195206 800 0 FreeSans 224 90 0 0 Tile_X5Y17_O_top1
port 2049 nsew signal input
flabel metal2 s 202234 0 202290 800 0 FreeSans 224 90 0 0 Tile_X5Y17_O_top10
port 2050 nsew signal input
flabel metal2 s 202878 0 202934 800 0 FreeSans 224 90 0 0 Tile_X5Y17_O_top11
port 2051 nsew signal input
flabel metal2 s 203522 0 203578 800 0 FreeSans 224 90 0 0 Tile_X5Y17_O_top12
port 2052 nsew signal input
flabel metal2 s 204166 0 204222 800 0 FreeSans 224 90 0 0 Tile_X5Y17_O_top13
port 2053 nsew signal input
flabel metal2 s 204810 0 204866 800 0 FreeSans 224 90 0 0 Tile_X5Y17_O_top14
port 2054 nsew signal input
flabel metal2 s 205454 0 205510 800 0 FreeSans 224 90 0 0 Tile_X5Y17_O_top15
port 2055 nsew signal input
flabel metal2 s 195794 0 195850 800 0 FreeSans 224 90 0 0 Tile_X5Y17_O_top2
port 2056 nsew signal input
flabel metal2 s 197082 0 197138 800 0 FreeSans 224 90 0 0 Tile_X5Y17_O_top3
port 2057 nsew signal input
flabel metal2 s 197726 0 197782 800 0 FreeSans 224 90 0 0 Tile_X5Y17_O_top4
port 2058 nsew signal input
flabel metal2 s 198370 0 198426 800 0 FreeSans 224 90 0 0 Tile_X5Y17_O_top5
port 2059 nsew signal input
flabel metal2 s 199014 0 199070 800 0 FreeSans 224 90 0 0 Tile_X5Y17_O_top6
port 2060 nsew signal input
flabel metal2 s 199658 0 199714 800 0 FreeSans 224 90 0 0 Tile_X5Y17_O_top7
port 2061 nsew signal input
flabel metal2 s 200302 0 200358 800 0 FreeSans 224 90 0 0 Tile_X5Y17_O_top8
port 2062 nsew signal input
flabel metal2 s 200946 0 201002 800 0 FreeSans 224 90 0 0 Tile_X5Y17_O_top9
port 2063 nsew signal input
flabel metal2 s 237010 755700 237066 756500 0 FreeSans 224 90 0 0 Tile_X6Y0_A_I_top
port 2064 nsew signal output
flabel metal2 s 235722 755700 235778 756500 0 FreeSans 224 90 0 0 Tile_X6Y0_A_O_top
port 2065 nsew signal input
flabel metal2 s 238298 755700 238354 756500 0 FreeSans 224 90 0 0 Tile_X6Y0_A_T_top
port 2066 nsew signal output
flabel metal2 s 242806 755700 242862 756500 0 FreeSans 224 90 0 0 Tile_X6Y0_A_config_C_bit0
port 2067 nsew signal output
flabel metal2 s 243450 755700 243506 756500 0 FreeSans 224 90 0 0 Tile_X6Y0_A_config_C_bit1
port 2068 nsew signal output
flabel metal2 s 244738 755700 244794 756500 0 FreeSans 224 90 0 0 Tile_X6Y0_A_config_C_bit2
port 2069 nsew signal output
flabel metal2 s 246026 755700 246082 756500 0 FreeSans 224 90 0 0 Tile_X6Y0_A_config_C_bit3
port 2070 nsew signal output
flabel metal2 s 240230 755700 240286 756500 0 FreeSans 224 90 0 0 Tile_X6Y0_B_I_top
port 2071 nsew signal output
flabel metal2 s 238942 755700 238998 756500 0 FreeSans 224 90 0 0 Tile_X6Y0_B_O_top
port 2072 nsew signal input
flabel metal2 s 241518 755700 241574 756500 0 FreeSans 224 90 0 0 Tile_X6Y0_B_T_top
port 2073 nsew signal output
flabel metal2 s 246670 755700 246726 756500 0 FreeSans 224 90 0 0 Tile_X6Y0_B_config_C_bit0
port 2074 nsew signal output
flabel metal2 s 247958 755700 248014 756500 0 FreeSans 224 90 0 0 Tile_X6Y0_B_config_C_bit1
port 2075 nsew signal output
flabel metal2 s 249246 755700 249302 756500 0 FreeSans 224 90 0 0 Tile_X6Y0_B_config_C_bit2
port 2076 nsew signal output
flabel metal2 s 250534 755700 250590 756500 0 FreeSans 224 90 0 0 Tile_X6Y0_B_config_C_bit3
port 2077 nsew signal output
flabel metal2 s 247314 0 247370 800 0 FreeSans 224 90 0 0 Tile_X6Y17_I_top0
port 2078 nsew signal output
flabel metal2 s 247958 0 248014 800 0 FreeSans 224 90 0 0 Tile_X6Y17_I_top1
port 2079 nsew signal output
flabel metal2 s 254398 0 254454 800 0 FreeSans 224 90 0 0 Tile_X6Y17_I_top10
port 2080 nsew signal output
flabel metal2 s 255686 0 255742 800 0 FreeSans 224 90 0 0 Tile_X6Y17_I_top11
port 2081 nsew signal output
flabel metal2 s 256330 0 256386 800 0 FreeSans 224 90 0 0 Tile_X6Y17_I_top12
port 2082 nsew signal output
flabel metal2 s 256974 0 257030 800 0 FreeSans 224 90 0 0 Tile_X6Y17_I_top13
port 2083 nsew signal output
flabel metal2 s 257618 0 257674 800 0 FreeSans 224 90 0 0 Tile_X6Y17_I_top14
port 2084 nsew signal output
flabel metal2 s 258262 0 258318 800 0 FreeSans 224 90 0 0 Tile_X6Y17_I_top15
port 2085 nsew signal output
flabel metal2 s 248602 0 248658 800 0 FreeSans 224 90 0 0 Tile_X6Y17_I_top2
port 2086 nsew signal output
flabel metal2 s 249246 0 249302 800 0 FreeSans 224 90 0 0 Tile_X6Y17_I_top3
port 2087 nsew signal output
flabel metal2 s 250534 0 250590 800 0 FreeSans 224 90 0 0 Tile_X6Y17_I_top4
port 2088 nsew signal output
flabel metal2 s 251178 0 251234 800 0 FreeSans 224 90 0 0 Tile_X6Y17_I_top5
port 2089 nsew signal output
flabel metal2 s 251822 0 251878 800 0 FreeSans 224 90 0 0 Tile_X6Y17_I_top6
port 2090 nsew signal output
flabel metal2 s 252466 0 252522 800 0 FreeSans 224 90 0 0 Tile_X6Y17_I_top7
port 2091 nsew signal output
flabel metal2 s 253110 0 253166 800 0 FreeSans 224 90 0 0 Tile_X6Y17_I_top8
port 2092 nsew signal output
flabel metal2 s 253754 0 253810 800 0 FreeSans 224 90 0 0 Tile_X6Y17_I_top9
port 2093 nsew signal output
flabel metal2 s 235722 0 235778 800 0 FreeSans 224 90 0 0 Tile_X6Y17_O_top0
port 2094 nsew signal input
flabel metal2 s 236366 0 236422 800 0 FreeSans 224 90 0 0 Tile_X6Y17_O_top1
port 2095 nsew signal input
flabel metal2 s 242806 0 242862 800 0 FreeSans 224 90 0 0 Tile_X6Y17_O_top10
port 2096 nsew signal input
flabel metal2 s 243450 0 243506 800 0 FreeSans 224 90 0 0 Tile_X6Y17_O_top11
port 2097 nsew signal input
flabel metal2 s 244094 0 244150 800 0 FreeSans 224 90 0 0 Tile_X6Y17_O_top12
port 2098 nsew signal input
flabel metal2 s 245382 0 245438 800 0 FreeSans 224 90 0 0 Tile_X6Y17_O_top13
port 2099 nsew signal input
flabel metal2 s 246026 0 246082 800 0 FreeSans 224 90 0 0 Tile_X6Y17_O_top14
port 2100 nsew signal input
flabel metal2 s 246670 0 246726 800 0 FreeSans 224 90 0 0 Tile_X6Y17_O_top15
port 2101 nsew signal input
flabel metal2 s 237010 0 237066 800 0 FreeSans 224 90 0 0 Tile_X6Y17_O_top2
port 2102 nsew signal input
flabel metal2 s 237654 0 237710 800 0 FreeSans 224 90 0 0 Tile_X6Y17_O_top3
port 2103 nsew signal input
flabel metal2 s 238298 0 238354 800 0 FreeSans 224 90 0 0 Tile_X6Y17_O_top4
port 2104 nsew signal input
flabel metal2 s 238942 0 238998 800 0 FreeSans 224 90 0 0 Tile_X6Y17_O_top5
port 2105 nsew signal input
flabel metal2 s 240230 0 240286 800 0 FreeSans 224 90 0 0 Tile_X6Y17_O_top6
port 2106 nsew signal input
flabel metal2 s 240874 0 240930 800 0 FreeSans 224 90 0 0 Tile_X6Y17_O_top7
port 2107 nsew signal input
flabel metal2 s 241518 0 241574 800 0 FreeSans 224 90 0 0 Tile_X6Y17_O_top8
port 2108 nsew signal input
flabel metal2 s 242162 0 242218 800 0 FreeSans 224 90 0 0 Tile_X6Y17_O_top9
port 2109 nsew signal input
flabel metal2 s 323306 755700 323362 756500 0 FreeSans 224 90 0 0 Tile_X8Y0_A_I_top
port 2110 nsew signal output
flabel metal2 s 322018 755700 322074 756500 0 FreeSans 224 90 0 0 Tile_X8Y0_A_O_top
port 2111 nsew signal input
flabel metal2 s 323950 755700 324006 756500 0 FreeSans 224 90 0 0 Tile_X8Y0_A_T_top
port 2112 nsew signal output
flabel metal2 s 328458 755700 328514 756500 0 FreeSans 224 90 0 0 Tile_X8Y0_A_config_C_bit0
port 2113 nsew signal output
flabel metal2 s 329746 755700 329802 756500 0 FreeSans 224 90 0 0 Tile_X8Y0_A_config_C_bit1
port 2114 nsew signal output
flabel metal2 s 331034 755700 331090 756500 0 FreeSans 224 90 0 0 Tile_X8Y0_A_config_C_bit2
port 2115 nsew signal output
flabel metal2 s 331678 755700 331734 756500 0 FreeSans 224 90 0 0 Tile_X8Y0_A_config_C_bit3
port 2116 nsew signal output
flabel metal2 s 326526 755700 326582 756500 0 FreeSans 224 90 0 0 Tile_X8Y0_B_I_top
port 2117 nsew signal output
flabel metal2 s 325238 755700 325294 756500 0 FreeSans 224 90 0 0 Tile_X8Y0_B_O_top
port 2118 nsew signal input
flabel metal2 s 327170 755700 327226 756500 0 FreeSans 224 90 0 0 Tile_X8Y0_B_T_top
port 2119 nsew signal output
flabel metal2 s 332966 755700 333022 756500 0 FreeSans 224 90 0 0 Tile_X8Y0_B_config_C_bit0
port 2120 nsew signal output
flabel metal2 s 334254 755700 334310 756500 0 FreeSans 224 90 0 0 Tile_X8Y0_B_config_C_bit1
port 2121 nsew signal output
flabel metal2 s 334898 755700 334954 756500 0 FreeSans 224 90 0 0 Tile_X8Y0_B_config_C_bit2
port 2122 nsew signal output
flabel metal2 s 336186 755700 336242 756500 0 FreeSans 224 90 0 0 Tile_X8Y0_B_config_C_bit3
port 2123 nsew signal output
flabel metal2 s 333610 0 333666 800 0 FreeSans 224 90 0 0 Tile_X8Y17_I_top0
port 2124 nsew signal output
flabel metal2 s 334254 0 334310 800 0 FreeSans 224 90 0 0 Tile_X8Y17_I_top1
port 2125 nsew signal output
flabel metal2 s 340694 0 340750 800 0 FreeSans 224 90 0 0 Tile_X8Y17_I_top10
port 2126 nsew signal output
flabel metal2 s 341338 0 341394 800 0 FreeSans 224 90 0 0 Tile_X8Y17_I_top11
port 2127 nsew signal output
flabel metal2 s 341982 0 342038 800 0 FreeSans 224 90 0 0 Tile_X8Y17_I_top12
port 2128 nsew signal output
flabel metal2 s 342626 0 342682 800 0 FreeSans 224 90 0 0 Tile_X8Y17_I_top13
port 2129 nsew signal output
flabel metal2 s 343914 0 343970 800 0 FreeSans 224 90 0 0 Tile_X8Y17_I_top14
port 2130 nsew signal output
flabel metal2 s 344558 0 344614 800 0 FreeSans 224 90 0 0 Tile_X8Y17_I_top15
port 2131 nsew signal output
flabel metal2 s 334898 0 334954 800 0 FreeSans 224 90 0 0 Tile_X8Y17_I_top2
port 2132 nsew signal output
flabel metal2 s 335542 0 335598 800 0 FreeSans 224 90 0 0 Tile_X8Y17_I_top3
port 2133 nsew signal output
flabel metal2 s 336186 0 336242 800 0 FreeSans 224 90 0 0 Tile_X8Y17_I_top4
port 2134 nsew signal output
flabel metal2 s 336830 0 336886 800 0 FreeSans 224 90 0 0 Tile_X8Y17_I_top5
port 2135 nsew signal output
flabel metal2 s 337474 0 337530 800 0 FreeSans 224 90 0 0 Tile_X8Y17_I_top6
port 2136 nsew signal output
flabel metal2 s 338762 0 338818 800 0 FreeSans 224 90 0 0 Tile_X8Y17_I_top7
port 2137 nsew signal output
flabel metal2 s 339406 0 339462 800 0 FreeSans 224 90 0 0 Tile_X8Y17_I_top8
port 2138 nsew signal output
flabel metal2 s 340050 0 340106 800 0 FreeSans 224 90 0 0 Tile_X8Y17_I_top9
port 2139 nsew signal output
flabel metal2 s 321374 0 321430 800 0 FreeSans 224 90 0 0 Tile_X8Y17_O_top0
port 2140 nsew signal input
flabel metal2 s 322018 0 322074 800 0 FreeSans 224 90 0 0 Tile_X8Y17_O_top1
port 2141 nsew signal input
flabel metal2 s 329102 0 329158 800 0 FreeSans 224 90 0 0 Tile_X8Y17_O_top10
port 2142 nsew signal input
flabel metal2 s 329746 0 329802 800 0 FreeSans 224 90 0 0 Tile_X8Y17_O_top11
port 2143 nsew signal input
flabel metal2 s 330390 0 330446 800 0 FreeSans 224 90 0 0 Tile_X8Y17_O_top12
port 2144 nsew signal input
flabel metal2 s 331034 0 331090 800 0 FreeSans 224 90 0 0 Tile_X8Y17_O_top13
port 2145 nsew signal input
flabel metal2 s 331678 0 331734 800 0 FreeSans 224 90 0 0 Tile_X8Y17_O_top14
port 2146 nsew signal input
flabel metal2 s 332322 0 332378 800 0 FreeSans 224 90 0 0 Tile_X8Y17_O_top15
port 2147 nsew signal input
flabel metal2 s 323306 0 323362 800 0 FreeSans 224 90 0 0 Tile_X8Y17_O_top2
port 2148 nsew signal input
flabel metal2 s 323950 0 324006 800 0 FreeSans 224 90 0 0 Tile_X8Y17_O_top3
port 2149 nsew signal input
flabel metal2 s 324594 0 324650 800 0 FreeSans 224 90 0 0 Tile_X8Y17_O_top4
port 2150 nsew signal input
flabel metal2 s 325238 0 325294 800 0 FreeSans 224 90 0 0 Tile_X8Y17_O_top5
port 2151 nsew signal input
flabel metal2 s 325882 0 325938 800 0 FreeSans 224 90 0 0 Tile_X8Y17_O_top6
port 2152 nsew signal input
flabel metal2 s 326526 0 326582 800 0 FreeSans 224 90 0 0 Tile_X8Y17_O_top7
port 2153 nsew signal input
flabel metal2 s 327170 0 327226 800 0 FreeSans 224 90 0 0 Tile_X8Y17_O_top8
port 2154 nsew signal input
flabel metal2 s 328458 0 328514 800 0 FreeSans 224 90 0 0 Tile_X8Y17_O_top9
port 2155 nsew signal input
flabel metal2 s 363878 755700 363934 756500 0 FreeSans 224 90 0 0 Tile_X9Y0_A_I_top
port 2156 nsew signal output
flabel metal2 s 363234 755700 363290 756500 0 FreeSans 224 90 0 0 Tile_X9Y0_A_O_top
port 2157 nsew signal input
flabel metal2 s 365166 755700 365222 756500 0 FreeSans 224 90 0 0 Tile_X9Y0_A_T_top
port 2158 nsew signal output
flabel metal2 s 369674 755700 369730 756500 0 FreeSans 224 90 0 0 Tile_X9Y0_A_config_C_bit0
port 2159 nsew signal output
flabel metal2 s 370962 755700 371018 756500 0 FreeSans 224 90 0 0 Tile_X9Y0_A_config_C_bit1
port 2160 nsew signal output
flabel metal2 s 371606 755700 371662 756500 0 FreeSans 224 90 0 0 Tile_X9Y0_A_config_C_bit2
port 2161 nsew signal output
flabel metal2 s 372894 755700 372950 756500 0 FreeSans 224 90 0 0 Tile_X9Y0_A_config_C_bit3
port 2162 nsew signal output
flabel metal2 s 367098 755700 367154 756500 0 FreeSans 224 90 0 0 Tile_X9Y0_B_I_top
port 2163 nsew signal output
flabel metal2 s 366454 755700 366510 756500 0 FreeSans 224 90 0 0 Tile_X9Y0_B_O_top
port 2164 nsew signal input
flabel metal2 s 368386 755700 368442 756500 0 FreeSans 224 90 0 0 Tile_X9Y0_B_T_top
port 2165 nsew signal output
flabel metal2 s 374182 755700 374238 756500 0 FreeSans 224 90 0 0 Tile_X9Y0_B_config_C_bit0
port 2166 nsew signal output
flabel metal2 s 374826 755700 374882 756500 0 FreeSans 224 90 0 0 Tile_X9Y0_B_config_C_bit1
port 2167 nsew signal output
flabel metal2 s 376114 755700 376170 756500 0 FreeSans 224 90 0 0 Tile_X9Y0_B_config_C_bit2
port 2168 nsew signal output
flabel metal2 s 377402 755700 377458 756500 0 FreeSans 224 90 0 0 Tile_X9Y0_B_config_C_bit3
port 2169 nsew signal output
flabel metal2 s 362590 0 362646 800 0 FreeSans 224 90 0 0 Tile_X9Y17_CMP_top
port 2170 nsew signal input
flabel metal2 s 363234 0 363290 800 0 FreeSans 224 90 0 0 Tile_X9Y17_HOLD_top
port 2171 nsew signal output
flabel metal2 s 364522 0 364578 800 0 FreeSans 224 90 0 0 Tile_X9Y17_RESET_top
port 2172 nsew signal output
flabel metal2 s 365810 0 365866 800 0 FreeSans 224 90 0 0 Tile_X9Y17_VALUE_top0
port 2173 nsew signal output
flabel metal2 s 367098 0 367154 800 0 FreeSans 224 90 0 0 Tile_X9Y17_VALUE_top1
port 2174 nsew signal output
flabel metal2 s 376758 0 376814 800 0 FreeSans 224 90 0 0 Tile_X9Y17_VALUE_top10
port 2175 nsew signal output
flabel metal2 s 378046 0 378102 800 0 FreeSans 224 90 0 0 Tile_X9Y17_VALUE_top11
port 2176 nsew signal output
flabel metal2 s 367742 0 367798 800 0 FreeSans 224 90 0 0 Tile_X9Y17_VALUE_top2
port 2177 nsew signal output
flabel metal2 s 369030 0 369086 800 0 FreeSans 224 90 0 0 Tile_X9Y17_VALUE_top3
port 2178 nsew signal output
flabel metal2 s 370318 0 370374 800 0 FreeSans 224 90 0 0 Tile_X9Y17_VALUE_top4
port 2179 nsew signal output
flabel metal2 s 370962 0 371018 800 0 FreeSans 224 90 0 0 Tile_X9Y17_VALUE_top5
port 2180 nsew signal output
flabel metal2 s 372250 0 372306 800 0 FreeSans 224 90 0 0 Tile_X9Y17_VALUE_top6
port 2181 nsew signal output
flabel metal2 s 373538 0 373594 800 0 FreeSans 224 90 0 0 Tile_X9Y17_VALUE_top7
port 2182 nsew signal output
flabel metal2 s 374826 0 374882 800 0 FreeSans 224 90 0 0 Tile_X9Y17_VALUE_top8
port 2183 nsew signal output
flabel metal2 s 375470 0 375526 800 0 FreeSans 224 90 0 0 Tile_X9Y17_VALUE_top9
port 2184 nsew signal output
flabel metal2 s 14186 0 14242 800 0 FreeSans 224 90 0 0 UserCLK
port 2185 nsew signal input
flabel metal4 s 13004 6000 13324 748500 0 FreeSans 1920 90 0 0 VGND
port 2186 nsew ground bidirectional
flabel metal4 s 19004 6000 19324 748500 0 FreeSans 1920 90 0 0 VGND
port 2186 nsew ground bidirectional
flabel metal4 s 24254 6000 24574 748500 0 FreeSans 1920 90 0 0 VGND
port 2186 nsew ground bidirectional
flabel metal4 s 30254 6000 30574 748500 0 FreeSans 1920 90 0 0 VGND
port 2186 nsew ground bidirectional
flabel metal4 s 36254 6000 36574 748500 0 FreeSans 1920 90 0 0 VGND
port 2186 nsew ground bidirectional
flabel metal4 s 42254 6000 42574 748500 0 FreeSans 1920 90 0 0 VGND
port 2186 nsew ground bidirectional
flabel metal4 s 48254 6000 48574 748500 0 FreeSans 1920 90 0 0 VGND
port 2186 nsew ground bidirectional
flabel metal4 s 54254 6000 54574 748500 0 FreeSans 1920 90 0 0 VGND
port 2186 nsew ground bidirectional
flabel metal4 s 60254 6000 60574 748500 0 FreeSans 1920 90 0 0 VGND
port 2186 nsew ground bidirectional
flabel metal4 s 65254 6000 65574 748500 0 FreeSans 1920 90 0 0 VGND
port 2186 nsew ground bidirectional
flabel metal4 s 71254 6000 71574 748500 0 FreeSans 1920 90 0 0 VGND
port 2186 nsew ground bidirectional
flabel metal4 s 77254 6000 77574 748500 0 FreeSans 1920 90 0 0 VGND
port 2186 nsew ground bidirectional
flabel metal4 s 83254 6000 83574 748500 0 FreeSans 1920 90 0 0 VGND
port 2186 nsew ground bidirectional
flabel metal4 s 89254 6000 89574 748500 0 FreeSans 1920 90 0 0 VGND
port 2186 nsew ground bidirectional
flabel metal4 s 95254 6000 95574 748500 0 FreeSans 1920 90 0 0 VGND
port 2186 nsew ground bidirectional
flabel metal4 s 101254 6000 101574 748500 0 FreeSans 1920 90 0 0 VGND
port 2186 nsew ground bidirectional
flabel metal4 s 106254 6000 106574 748500 0 FreeSans 1920 90 0 0 VGND
port 2186 nsew ground bidirectional
flabel metal4 s 112254 6000 112574 748500 0 FreeSans 1920 90 0 0 VGND
port 2186 nsew ground bidirectional
flabel metal4 s 118254 6000 118574 748500 0 FreeSans 1920 90 0 0 VGND
port 2186 nsew ground bidirectional
flabel metal4 s 124254 6000 124574 748500 0 FreeSans 1920 90 0 0 VGND
port 2186 nsew ground bidirectional
flabel metal4 s 130254 6000 130574 748500 0 FreeSans 1920 90 0 0 VGND
port 2186 nsew ground bidirectional
flabel metal4 s 136254 6000 136574 748500 0 FreeSans 1920 90 0 0 VGND
port 2186 nsew ground bidirectional
flabel metal4 s 142254 6000 142574 748500 0 FreeSans 1920 90 0 0 VGND
port 2186 nsew ground bidirectional
flabel metal4 s 148254 6000 148574 748500 0 FreeSans 1920 90 0 0 VGND
port 2186 nsew ground bidirectional
flabel metal4 s 155254 6000 155574 748500 0 FreeSans 1920 90 0 0 VGND
port 2186 nsew ground bidirectional
flabel metal4 s 161254 6000 161574 748500 0 FreeSans 1920 90 0 0 VGND
port 2186 nsew ground bidirectional
flabel metal4 s 167254 6000 167574 748500 0 FreeSans 1920 90 0 0 VGND
port 2186 nsew ground bidirectional
flabel metal4 s 173254 6000 173574 748500 0 FreeSans 1920 90 0 0 VGND
port 2186 nsew ground bidirectional
flabel metal4 s 179254 6000 179574 748500 0 FreeSans 1920 90 0 0 VGND
port 2186 nsew ground bidirectional
flabel metal4 s 185254 6000 185574 748500 0 FreeSans 1920 90 0 0 VGND
port 2186 nsew ground bidirectional
flabel metal4 s 191254 6000 191574 748500 0 FreeSans 1920 90 0 0 VGND
port 2186 nsew ground bidirectional
flabel metal4 s 196254 6000 196574 748500 0 FreeSans 1920 90 0 0 VGND
port 2186 nsew ground bidirectional
flabel metal4 s 202254 6000 202574 748500 0 FreeSans 1920 90 0 0 VGND
port 2186 nsew ground bidirectional
flabel metal4 s 208254 6000 208574 748500 0 FreeSans 1920 90 0 0 VGND
port 2186 nsew ground bidirectional
flabel metal4 s 214254 6000 214574 748500 0 FreeSans 1920 90 0 0 VGND
port 2186 nsew ground bidirectional
flabel metal4 s 220254 6000 220574 748500 0 FreeSans 1920 90 0 0 VGND
port 2186 nsew ground bidirectional
flabel metal4 s 226254 6000 226574 748500 0 FreeSans 1920 90 0 0 VGND
port 2186 nsew ground bidirectional
flabel metal4 s 232254 6000 232574 748500 0 FreeSans 1920 90 0 0 VGND
port 2186 nsew ground bidirectional
flabel metal4 s 237254 6000 237574 748500 0 FreeSans 1920 90 0 0 VGND
port 2186 nsew ground bidirectional
flabel metal4 s 243254 6000 243574 748500 0 FreeSans 1920 90 0 0 VGND
port 2186 nsew ground bidirectional
flabel metal4 s 249254 6000 249574 748500 0 FreeSans 1920 90 0 0 VGND
port 2186 nsew ground bidirectional
flabel metal4 s 255254 6000 255574 748500 0 FreeSans 1920 90 0 0 VGND
port 2186 nsew ground bidirectional
flabel metal4 s 261254 6000 261574 748500 0 FreeSans 1920 90 0 0 VGND
port 2186 nsew ground bidirectional
flabel metal4 s 267254 6000 267574 748500 0 FreeSans 1920 90 0 0 VGND
port 2186 nsew ground bidirectional
flabel metal4 s 273254 6000 273574 748500 0 FreeSans 1920 90 0 0 VGND
port 2186 nsew ground bidirectional
flabel metal4 s 278254 6000 278574 748500 0 FreeSans 1920 90 0 0 VGND
port 2186 nsew ground bidirectional
flabel metal4 s 284254 6000 284574 748500 0 FreeSans 1920 90 0 0 VGND
port 2186 nsew ground bidirectional
flabel metal4 s 290254 6000 290574 748500 0 FreeSans 1920 90 0 0 VGND
port 2186 nsew ground bidirectional
flabel metal4 s 296254 6000 296574 748500 0 FreeSans 1920 90 0 0 VGND
port 2186 nsew ground bidirectional
flabel metal4 s 302254 6000 302574 748500 0 FreeSans 1920 90 0 0 VGND
port 2186 nsew ground bidirectional
flabel metal4 s 308254 6000 308574 748500 0 FreeSans 1920 90 0 0 VGND
port 2186 nsew ground bidirectional
flabel metal4 s 314254 6000 314574 748500 0 FreeSans 1920 90 0 0 VGND
port 2186 nsew ground bidirectional
flabel metal4 s 323254 6000 323574 748500 0 FreeSans 1920 90 0 0 VGND
port 2186 nsew ground bidirectional
flabel metal4 s 329254 6000 329574 748500 0 FreeSans 1920 90 0 0 VGND
port 2186 nsew ground bidirectional
flabel metal4 s 335254 6000 335574 748500 0 FreeSans 1920 90 0 0 VGND
port 2186 nsew ground bidirectional
flabel metal4 s 341254 6000 341574 748500 0 FreeSans 1920 90 0 0 VGND
port 2186 nsew ground bidirectional
flabel metal4 s 347254 6000 347574 748500 0 FreeSans 1920 90 0 0 VGND
port 2186 nsew ground bidirectional
flabel metal4 s 353254 6000 353574 748500 0 FreeSans 1920 90 0 0 VGND
port 2186 nsew ground bidirectional
flabel metal4 s 359254 6000 359574 748500 0 FreeSans 1920 90 0 0 VGND
port 2186 nsew ground bidirectional
flabel metal4 s 364254 6000 364574 748500 0 FreeSans 1920 90 0 0 VGND
port 2186 nsew ground bidirectional
flabel metal4 s 370254 6000 370574 748500 0 FreeSans 1920 90 0 0 VGND
port 2186 nsew ground bidirectional
flabel metal4 s 376254 6000 376574 748500 0 FreeSans 1920 90 0 0 VGND
port 2186 nsew ground bidirectional
flabel metal4 s 382254 6000 382574 748500 0 FreeSans 1920 90 0 0 VGND
port 2186 nsew ground bidirectional
flabel metal4 s 388254 6000 388574 748500 0 FreeSans 1920 90 0 0 VGND
port 2186 nsew ground bidirectional
flabel metal4 s 394254 6000 394574 748500 0 FreeSans 1920 90 0 0 VGND
port 2186 nsew ground bidirectional
flabel metal4 s 400254 6000 400574 748500 0 FreeSans 1920 90 0 0 VGND
port 2186 nsew ground bidirectional
flabel metal4 s 405254 6000 405574 748500 0 FreeSans 1920 90 0 0 VGND
port 2186 nsew ground bidirectional
flabel metal4 s 411254 6000 411574 748500 0 FreeSans 1920 90 0 0 VGND
port 2186 nsew ground bidirectional
flabel metal4 s 417254 6000 417574 748500 0 FreeSans 1920 90 0 0 VGND
port 2186 nsew ground bidirectional
flabel metal4 s 423254 6000 423574 748500 0 FreeSans 1920 90 0 0 VGND
port 2186 nsew ground bidirectional
flabel metal4 s 429254 6000 429574 748500 0 FreeSans 1920 90 0 0 VGND
port 2186 nsew ground bidirectional
flabel metal4 s 435254 6000 435574 748500 0 FreeSans 1920 90 0 0 VGND
port 2186 nsew ground bidirectional
flabel metal4 s 441254 6000 441574 748500 0 FreeSans 1920 90 0 0 VGND
port 2186 nsew ground bidirectional
flabel metal4 s 446254 6000 446574 748500 0 FreeSans 1920 90 0 0 VGND
port 2186 nsew ground bidirectional
flabel metal4 s 452254 6000 452574 748500 0 FreeSans 1920 90 0 0 VGND
port 2186 nsew ground bidirectional
flabel metal4 s 458254 6000 458574 748500 0 FreeSans 1920 90 0 0 VGND
port 2186 nsew ground bidirectional
flabel metal4 s 464254 6000 464574 748500 0 FreeSans 1920 90 0 0 VGND
port 2186 nsew ground bidirectional
flabel metal4 s 470254 6000 470574 748500 0 FreeSans 1920 90 0 0 VGND
port 2186 nsew ground bidirectional
flabel metal4 s 11944 6000 12264 748500 0 FreeSans 1920 90 0 0 VPWR
port 2187 nsew power bidirectional
flabel metal4 s 17944 6000 18264 748500 0 FreeSans 1920 90 0 0 VPWR
port 2187 nsew power bidirectional
flabel metal4 s 23194 6000 23514 748500 0 FreeSans 1920 90 0 0 VPWR
port 2187 nsew power bidirectional
flabel metal4 s 29194 6000 29514 748500 0 FreeSans 1920 90 0 0 VPWR
port 2187 nsew power bidirectional
flabel metal4 s 35194 6000 35514 748500 0 FreeSans 1920 90 0 0 VPWR
port 2187 nsew power bidirectional
flabel metal4 s 41194 6000 41514 748500 0 FreeSans 1920 90 0 0 VPWR
port 2187 nsew power bidirectional
flabel metal4 s 47194 6000 47514 748500 0 FreeSans 1920 90 0 0 VPWR
port 2187 nsew power bidirectional
flabel metal4 s 53194 6000 53514 748500 0 FreeSans 1920 90 0 0 VPWR
port 2187 nsew power bidirectional
flabel metal4 s 59194 6000 59514 748500 0 FreeSans 1920 90 0 0 VPWR
port 2187 nsew power bidirectional
flabel metal4 s 64194 6000 64514 748500 0 FreeSans 1920 90 0 0 VPWR
port 2187 nsew power bidirectional
flabel metal4 s 70194 6000 70514 748500 0 FreeSans 1920 90 0 0 VPWR
port 2187 nsew power bidirectional
flabel metal4 s 76194 6000 76514 748500 0 FreeSans 1920 90 0 0 VPWR
port 2187 nsew power bidirectional
flabel metal4 s 82194 6000 82514 748500 0 FreeSans 1920 90 0 0 VPWR
port 2187 nsew power bidirectional
flabel metal4 s 88194 6000 88514 748500 0 FreeSans 1920 90 0 0 VPWR
port 2187 nsew power bidirectional
flabel metal4 s 94194 6000 94514 748500 0 FreeSans 1920 90 0 0 VPWR
port 2187 nsew power bidirectional
flabel metal4 s 100194 6000 100514 748500 0 FreeSans 1920 90 0 0 VPWR
port 2187 nsew power bidirectional
flabel metal4 s 105194 6000 105514 748500 0 FreeSans 1920 90 0 0 VPWR
port 2187 nsew power bidirectional
flabel metal4 s 111194 6000 111514 748500 0 FreeSans 1920 90 0 0 VPWR
port 2187 nsew power bidirectional
flabel metal4 s 117194 6000 117514 748500 0 FreeSans 1920 90 0 0 VPWR
port 2187 nsew power bidirectional
flabel metal4 s 123194 6000 123514 748500 0 FreeSans 1920 90 0 0 VPWR
port 2187 nsew power bidirectional
flabel metal4 s 129194 6000 129514 748500 0 FreeSans 1920 90 0 0 VPWR
port 2187 nsew power bidirectional
flabel metal4 s 135194 6000 135514 748500 0 FreeSans 1920 90 0 0 VPWR
port 2187 nsew power bidirectional
flabel metal4 s 141194 6000 141514 748500 0 FreeSans 1920 90 0 0 VPWR
port 2187 nsew power bidirectional
flabel metal4 s 147194 6000 147514 748500 0 FreeSans 1920 90 0 0 VPWR
port 2187 nsew power bidirectional
flabel metal4 s 154194 6000 154514 748500 0 FreeSans 1920 90 0 0 VPWR
port 2187 nsew power bidirectional
flabel metal4 s 160194 6000 160514 748500 0 FreeSans 1920 90 0 0 VPWR
port 2187 nsew power bidirectional
flabel metal4 s 166194 6000 166514 748500 0 FreeSans 1920 90 0 0 VPWR
port 2187 nsew power bidirectional
flabel metal4 s 172194 6000 172514 748500 0 FreeSans 1920 90 0 0 VPWR
port 2187 nsew power bidirectional
flabel metal4 s 178194 6000 178514 748500 0 FreeSans 1920 90 0 0 VPWR
port 2187 nsew power bidirectional
flabel metal4 s 184194 6000 184514 748500 0 FreeSans 1920 90 0 0 VPWR
port 2187 nsew power bidirectional
flabel metal4 s 190194 6000 190514 748500 0 FreeSans 1920 90 0 0 VPWR
port 2187 nsew power bidirectional
flabel metal4 s 195194 6000 195514 748500 0 FreeSans 1920 90 0 0 VPWR
port 2187 nsew power bidirectional
flabel metal4 s 201194 6000 201514 748500 0 FreeSans 1920 90 0 0 VPWR
port 2187 nsew power bidirectional
flabel metal4 s 207194 6000 207514 748500 0 FreeSans 1920 90 0 0 VPWR
port 2187 nsew power bidirectional
flabel metal4 s 213194 6000 213514 748500 0 FreeSans 1920 90 0 0 VPWR
port 2187 nsew power bidirectional
flabel metal4 s 219194 6000 219514 748500 0 FreeSans 1920 90 0 0 VPWR
port 2187 nsew power bidirectional
flabel metal4 s 225194 6000 225514 748500 0 FreeSans 1920 90 0 0 VPWR
port 2187 nsew power bidirectional
flabel metal4 s 231194 6000 231514 748500 0 FreeSans 1920 90 0 0 VPWR
port 2187 nsew power bidirectional
flabel metal4 s 236194 6000 236514 748500 0 FreeSans 1920 90 0 0 VPWR
port 2187 nsew power bidirectional
flabel metal4 s 242194 6000 242514 748500 0 FreeSans 1920 90 0 0 VPWR
port 2187 nsew power bidirectional
flabel metal4 s 248194 6000 248514 748500 0 FreeSans 1920 90 0 0 VPWR
port 2187 nsew power bidirectional
flabel metal4 s 254194 6000 254514 748500 0 FreeSans 1920 90 0 0 VPWR
port 2187 nsew power bidirectional
flabel metal4 s 260194 6000 260514 748500 0 FreeSans 1920 90 0 0 VPWR
port 2187 nsew power bidirectional
flabel metal4 s 266194 6000 266514 748500 0 FreeSans 1920 90 0 0 VPWR
port 2187 nsew power bidirectional
flabel metal4 s 272194 6000 272514 748500 0 FreeSans 1920 90 0 0 VPWR
port 2187 nsew power bidirectional
flabel metal4 s 277194 6000 277514 748500 0 FreeSans 1920 90 0 0 VPWR
port 2187 nsew power bidirectional
flabel metal4 s 283194 6000 283514 748500 0 FreeSans 1920 90 0 0 VPWR
port 2187 nsew power bidirectional
flabel metal4 s 289194 6000 289514 748500 0 FreeSans 1920 90 0 0 VPWR
port 2187 nsew power bidirectional
flabel metal4 s 295194 6000 295514 748500 0 FreeSans 1920 90 0 0 VPWR
port 2187 nsew power bidirectional
flabel metal4 s 301194 6000 301514 748500 0 FreeSans 1920 90 0 0 VPWR
port 2187 nsew power bidirectional
flabel metal4 s 307194 6000 307514 748500 0 FreeSans 1920 90 0 0 VPWR
port 2187 nsew power bidirectional
flabel metal4 s 313194 6000 313514 748500 0 FreeSans 1920 90 0 0 VPWR
port 2187 nsew power bidirectional
flabel metal4 s 322194 6000 322514 748500 0 FreeSans 1920 90 0 0 VPWR
port 2187 nsew power bidirectional
flabel metal4 s 328194 6000 328514 748500 0 FreeSans 1920 90 0 0 VPWR
port 2187 nsew power bidirectional
flabel metal4 s 334194 6000 334514 748500 0 FreeSans 1920 90 0 0 VPWR
port 2187 nsew power bidirectional
flabel metal4 s 340194 6000 340514 748500 0 FreeSans 1920 90 0 0 VPWR
port 2187 nsew power bidirectional
flabel metal4 s 346194 6000 346514 748500 0 FreeSans 1920 90 0 0 VPWR
port 2187 nsew power bidirectional
flabel metal4 s 352194 6000 352514 748500 0 FreeSans 1920 90 0 0 VPWR
port 2187 nsew power bidirectional
flabel metal4 s 358194 6000 358514 748500 0 FreeSans 1920 90 0 0 VPWR
port 2187 nsew power bidirectional
flabel metal4 s 363194 6000 363514 748500 0 FreeSans 1920 90 0 0 VPWR
port 2187 nsew power bidirectional
flabel metal4 s 369194 6000 369514 748500 0 FreeSans 1920 90 0 0 VPWR
port 2187 nsew power bidirectional
flabel metal4 s 375194 6000 375514 748500 0 FreeSans 1920 90 0 0 VPWR
port 2187 nsew power bidirectional
flabel metal4 s 381194 6000 381514 748500 0 FreeSans 1920 90 0 0 VPWR
port 2187 nsew power bidirectional
flabel metal4 s 387194 6000 387514 748500 0 FreeSans 1920 90 0 0 VPWR
port 2187 nsew power bidirectional
flabel metal4 s 393194 6000 393514 748500 0 FreeSans 1920 90 0 0 VPWR
port 2187 nsew power bidirectional
flabel metal4 s 399194 6000 399514 748500 0 FreeSans 1920 90 0 0 VPWR
port 2187 nsew power bidirectional
flabel metal4 s 404194 6000 404514 748500 0 FreeSans 1920 90 0 0 VPWR
port 2187 nsew power bidirectional
flabel metal4 s 410194 6000 410514 748500 0 FreeSans 1920 90 0 0 VPWR
port 2187 nsew power bidirectional
flabel metal4 s 416194 6000 416514 748500 0 FreeSans 1920 90 0 0 VPWR
port 2187 nsew power bidirectional
flabel metal4 s 422194 6000 422514 748500 0 FreeSans 1920 90 0 0 VPWR
port 2187 nsew power bidirectional
flabel metal4 s 428194 6000 428514 748500 0 FreeSans 1920 90 0 0 VPWR
port 2187 nsew power bidirectional
flabel metal4 s 434194 6000 434514 748500 0 FreeSans 1920 90 0 0 VPWR
port 2187 nsew power bidirectional
flabel metal4 s 440194 6000 440514 748500 0 FreeSans 1920 90 0 0 VPWR
port 2187 nsew power bidirectional
flabel metal4 s 445194 6000 445514 748500 0 FreeSans 1920 90 0 0 VPWR
port 2187 nsew power bidirectional
flabel metal4 s 451194 6000 451514 748500 0 FreeSans 1920 90 0 0 VPWR
port 2187 nsew power bidirectional
flabel metal4 s 457194 6000 457514 748500 0 FreeSans 1920 90 0 0 VPWR
port 2187 nsew power bidirectional
flabel metal4 s 463194 6000 463514 748500 0 FreeSans 1920 90 0 0 VPWR
port 2187 nsew power bidirectional
flabel metal4 s 469194 6000 469514 748500 0 FreeSans 1920 90 0 0 VPWR
port 2187 nsew power bidirectional
flabel metal4 s 475194 6000 475514 748500 0 FreeSans 1920 90 0 0 VPWR
port 2187 nsew power bidirectional
rlabel metal4 470414 377250 470414 377250 0 VGND
rlabel metal4 475354 377250 475354 377250 0 VPWR
rlabel metal3 14513 738684 14513 738684 0 FrameData[0]
rlabel metal3 3787 620908 3787 620908 0 FrameData[100]
rlabel metal3 3787 621588 3787 621588 0 FrameData[101]
rlabel metal3 9476 622847 9476 622847 0 FrameData[102]
rlabel metal3 9476 623595 9476 623595 0 FrameData[103]
rlabel metal3 5341 624308 5341 624308 0 FrameData[104]
rlabel metal3 3787 624988 3787 624988 0 FrameData[105]
rlabel metal3 3787 625668 3787 625668 0 FrameData[106]
rlabel metal3 9476 626927 9476 626927 0 FrameData[107]
rlabel metal3 9476 627675 9476 627675 0 FrameData[108]
rlabel metal3 5341 628388 5341 628388 0 FrameData[109]
rlabel metal2 21245 755820 21245 755820 0 FrameData[10]
rlabel metal3 3787 629068 3787 629068 0 FrameData[110]
rlabel metal3 3787 629748 3787 629748 0 FrameData[111]
rlabel metal3 9476 631007 9476 631007 0 FrameData[112]
rlabel metal3 9476 631755 9476 631755 0 FrameData[113]
rlabel metal3 5341 632468 5341 632468 0 FrameData[114]
rlabel metal3 3787 633148 3787 633148 0 FrameData[115]
rlabel metal3 3787 633828 3787 633828 0 FrameData[116]
rlabel metal3 9476 635087 9476 635087 0 FrameData[117]
rlabel metal3 9476 635835 9476 635835 0 FrameData[118]
rlabel metal3 5341 636548 5341 636548 0 FrameData[119]
rlabel metal2 15555 755820 15555 755820 0 FrameData[11]
rlabel metal3 3787 637228 3787 637228 0 FrameData[120]
rlabel metal3 3787 637908 3787 637908 0 FrameData[121]
rlabel metal3 9476 639167 9476 639167 0 FrameData[122]
rlabel metal3 9476 639915 9476 639915 0 FrameData[123]
rlabel metal3 5341 640628 5341 640628 0 FrameData[124]
rlabel metal3 3787 641308 3787 641308 0 FrameData[125]
rlabel metal3 3787 641988 3787 641988 0 FrameData[126]
rlabel metal3 2407 643348 2407 643348 0 FrameData[127]
rlabel metal3 3787 572628 3787 572628 0 FrameData[128]
rlabel metal3 9476 573459 9476 573459 0 FrameData[129]
rlabel metal2 12229 755820 12229 755820 0 FrameData[12]
rlabel metal3 9476 574575 9476 574575 0 FrameData[130]
rlabel metal3 9476 575323 9476 575323 0 FrameData[131]
rlabel metal3 9476 576043 9476 576043 0 FrameData[132]
rlabel metal3 3143 576708 3143 576708 0 FrameData[133]
rlabel metal3 9476 577539 9476 577539 0 FrameData[134]
rlabel metal3 9476 578655 9476 578655 0 FrameData[135]
rlabel metal3 9476 579403 9476 579403 0 FrameData[136]
rlabel metal3 9476 580123 9476 580123 0 FrameData[137]
rlabel metal3 9476 580871 9476 580871 0 FrameData[138]
rlabel metal3 9476 581619 9476 581619 0 FrameData[139]
rlabel metal2 19957 755820 19957 755820 0 FrameData[13]
rlabel metal3 9476 582735 9476 582735 0 FrameData[140]
rlabel metal3 9476 583483 9476 583483 0 FrameData[141]
rlabel metal3 9476 584203 9476 584203 0 FrameData[142]
rlabel metal3 9476 584951 9476 584951 0 FrameData[143]
rlabel metal3 9476 585699 9476 585699 0 FrameData[144]
rlabel metal3 9476 586815 9476 586815 0 FrameData[145]
rlabel metal3 9476 587563 9476 587563 0 FrameData[146]
rlabel metal3 9476 588283 9476 588283 0 FrameData[147]
rlabel metal3 9476 589031 9476 589031 0 FrameData[148]
rlabel metal3 9476 589779 9476 589779 0 FrameData[149]
rlabel metal2 20608 753236 20608 753236 0 FrameData[14]
rlabel metal3 9476 590895 9476 590895 0 FrameData[150]
rlabel metal3 9476 591643 9476 591643 0 FrameData[151]
rlabel metal3 9476 592363 9476 592363 0 FrameData[152]
rlabel metal3 9476 593111 9476 593111 0 FrameData[153]
rlabel metal3 9476 593859 9476 593859 0 FrameData[154]
rlabel metal3 9476 594975 9476 594975 0 FrameData[155]
rlabel metal3 9476 595723 9476 595723 0 FrameData[156]
rlabel metal3 9476 596443 9476 596443 0 FrameData[157]
rlabel metal3 9476 597191 9476 597191 0 FrameData[158]
rlabel metal3 9476 597939 9476 597939 0 FrameData[159]
rlabel metal2 14805 755820 14805 755820 0 FrameData[15]
rlabel metal3 9476 527771 9476 527771 0 FrameData[160]
rlabel metal3 3143 528428 3143 528428 0 FrameData[161]
rlabel metal3 9476 529635 9476 529635 0 FrameData[162]
rlabel metal3 9476 530383 9476 530383 0 FrameData[163]
rlabel metal3 9476 531131 9476 531131 0 FrameData[164]
rlabel metal3 9476 531851 9476 531851 0 FrameData[165]
rlabel metal3 3787 532508 3787 532508 0 FrameData[166]
rlabel metal3 9476 533715 9476 533715 0 FrameData[167]
rlabel metal3 9476 534463 9476 534463 0 FrameData[168]
rlabel metal3 9476 535211 9476 535211 0 FrameData[169]
rlabel metal2 10403 755820 10403 755820 0 FrameData[16]
rlabel metal3 9476 535931 9476 535931 0 FrameData[170]
rlabel metal3 9476 536679 9476 536679 0 FrameData[171]
rlabel metal3 9476 537795 9476 537795 0 FrameData[172]
rlabel metal3 9476 538543 9476 538543 0 FrameData[173]
rlabel metal3 9476 539291 9476 539291 0 FrameData[174]
rlabel metal3 9476 540011 9476 540011 0 FrameData[175]
rlabel metal3 9476 540759 9476 540759 0 FrameData[176]
rlabel metal3 9476 541875 9476 541875 0 FrameData[177]
rlabel metal3 9476 542623 9476 542623 0 FrameData[178]
rlabel metal3 9476 543371 9476 543371 0 FrameData[179]
rlabel metal3 20608 743308 20608 743308 0 FrameData[17]
rlabel metal3 9476 544091 9476 544091 0 FrameData[180]
rlabel metal3 9476 544839 9476 544839 0 FrameData[181]
rlabel metal3 9476 545955 9476 545955 0 FrameData[182]
rlabel metal3 9476 546703 9476 546703 0 FrameData[183]
rlabel metal3 9476 547451 9476 547451 0 FrameData[184]
rlabel metal3 9476 548171 9476 548171 0 FrameData[185]
rlabel metal3 9476 548919 9476 548919 0 FrameData[186]
rlabel metal3 9476 550035 9476 550035 0 FrameData[187]
rlabel metal3 9476 550783 9476 550783 0 FrameData[188]
rlabel metal3 9476 551531 9476 551531 0 FrameData[189]
rlabel metal2 17381 755820 17381 755820 0 FrameData[18]
rlabel metal3 9476 552251 9476 552251 0 FrameData[190]
rlabel metal3 9476 552999 9476 552999 0 FrameData[191]
rlabel metal3 9476 482859 9476 482859 0 FrameData[192]
rlabel metal3 9476 483579 9476 483579 0 FrameData[193]
rlabel metal3 3787 484228 3787 484228 0 FrameData[194]
rlabel metal3 9476 485443 9476 485443 0 FrameData[195]
rlabel metal3 9476 486191 9476 486191 0 FrameData[196]
rlabel metal3 9476 486939 9476 486939 0 FrameData[197]
rlabel metal3 9476 487659 9476 487659 0 FrameData[198]
rlabel metal3 3787 488308 3787 488308 0 FrameData[199]
rlabel metal2 11691 755820 11691 755820 0 FrameData[19]
rlabel metal3 17733 738956 17733 738956 0 FrameData[1]
rlabel metal3 9476 489523 9476 489523 0 FrameData[200]
rlabel metal3 9476 490271 9476 490271 0 FrameData[201]
rlabel metal3 9476 491019 9476 491019 0 FrameData[202]
rlabel metal3 9476 491739 9476 491739 0 FrameData[203]
rlabel metal3 3787 492388 3787 492388 0 FrameData[204]
rlabel metal3 9476 493603 9476 493603 0 FrameData[205]
rlabel metal3 9476 494351 9476 494351 0 FrameData[206]
rlabel metal3 9476 495099 9476 495099 0 FrameData[207]
rlabel metal3 9476 495819 9476 495819 0 FrameData[208]
rlabel metal3 9476 496567 9476 496567 0 FrameData[209]
rlabel metal2 19419 755820 19419 755820 0 FrameData[20]
rlabel metal3 9476 497683 9476 497683 0 FrameData[210]
rlabel metal3 9476 498431 9476 498431 0 FrameData[211]
rlabel metal3 9476 499179 9476 499179 0 FrameData[212]
rlabel metal3 9476 499899 9476 499899 0 FrameData[213]
rlabel metal3 9476 500647 9476 500647 0 FrameData[214]
rlabel metal3 9476 501763 9476 501763 0 FrameData[215]
rlabel metal3 9476 502511 9476 502511 0 FrameData[216]
rlabel metal3 9476 503259 9476 503259 0 FrameData[217]
rlabel metal3 9476 503979 9476 503979 0 FrameData[218]
rlabel metal3 9476 504727 9476 504727 0 FrameData[219]
rlabel metal3 21896 753508 21896 753508 0 FrameData[21]
rlabel metal3 9476 505843 9476 505843 0 FrameData[220]
rlabel metal3 9476 506591 9476 506591 0 FrameData[221]
rlabel metal3 9476 507339 9476 507339 0 FrameData[222]
rlabel metal3 9476 508062 9476 508062 0 FrameData[223]
rlabel metal3 3787 437988 3787 437988 0 FrameData[224]
rlabel metal3 5338 438668 5338 438668 0 FrameData[225]
rlabel metal3 9476 439382 9476 439382 0 FrameData[226]
rlabel metal3 3787 440028 3787 440028 0 FrameData[227]
rlabel metal3 3787 441388 3787 441388 0 FrameData[228]
rlabel metal3 3787 442068 3787 442068 0 FrameData[229]
rlabel metal3 21942 754868 21942 754868 0 FrameData[22]
rlabel metal3 5338 442748 5338 442748 0 FrameData[230]
rlabel metal3 9476 443462 9476 443462 0 FrameData[231]
rlabel metal3 3787 444108 3787 444108 0 FrameData[232]
rlabel metal3 3787 445468 3787 445468 0 FrameData[233]
rlabel metal3 3787 446148 3787 446148 0 FrameData[234]
rlabel metal3 5338 446828 5338 446828 0 FrameData[235]
rlabel metal3 9476 447542 9476 447542 0 FrameData[236]
rlabel metal3 9476 448290 9476 448290 0 FrameData[237]
rlabel metal3 3787 449548 3787 449548 0 FrameData[238]
rlabel metal3 3787 450228 3787 450228 0 FrameData[239]
rlabel metal2 13517 755820 13517 755820 0 FrameData[23]
rlabel metal3 5338 450908 5338 450908 0 FrameData[240]
rlabel metal3 9476 451622 9476 451622 0 FrameData[241]
rlabel metal3 9476 452370 9476 452370 0 FrameData[242]
rlabel metal3 3787 453628 3787 453628 0 FrameData[243]
rlabel metal3 3787 454308 3787 454308 0 FrameData[244]
rlabel metal3 5338 454988 5338 454988 0 FrameData[245]
rlabel metal3 9476 455702 9476 455702 0 FrameData[246]
rlabel metal3 9476 456450 9476 456450 0 FrameData[247]
rlabel metal3 3787 457708 3787 457708 0 FrameData[248]
rlabel metal3 3787 458388 3787 458388 0 FrameData[249]
rlabel metal2 18669 755820 18669 755820 0 FrameData[24]
rlabel metal3 5338 459068 5338 459068 0 FrameData[250]
rlabel metal3 9476 459782 9476 459782 0 FrameData[251]
rlabel metal3 9476 460530 9476 460530 0 FrameData[252]
rlabel metal3 3787 461788 3787 461788 0 FrameData[253]
rlabel metal3 3787 462468 3787 462468 0 FrameData[254]
rlabel metal3 5338 463148 5338 463148 0 FrameData[255]
rlabel metal3 9476 392979 9476 392979 0 FrameData[256]
rlabel metal3 9476 393727 9476 393727 0 FrameData[257]
rlabel metal3 5338 394468 5338 394468 0 FrameData[258]
rlabel metal3 9476 395195 9476 395195 0 FrameData[259]
rlabel metal2 8365 755820 8365 755820 0 FrameData[25]
rlabel metal3 3787 395828 3787 395828 0 FrameData[260]
rlabel metal3 9476 397059 9476 397059 0 FrameData[261]
rlabel metal3 9476 397807 9476 397807 0 FrameData[262]
rlabel metal3 5338 398548 5338 398548 0 FrameData[263]
rlabel metal3 9476 399275 9476 399275 0 FrameData[264]
rlabel metal3 9476 400023 9476 400023 0 FrameData[265]
rlabel metal3 9476 401139 9476 401139 0 FrameData[266]
rlabel metal3 9476 401887 9476 401887 0 FrameData[267]
rlabel metal3 5338 402628 5338 402628 0 FrameData[268]
rlabel metal3 9476 403355 9476 403355 0 FrameData[269]
rlabel metal2 20516 753100 20516 753100 0 FrameData[26]
rlabel metal3 9476 404103 9476 404103 0 FrameData[270]
rlabel metal3 9476 405219 9476 405219 0 FrameData[271]
rlabel metal3 9476 405967 9476 405967 0 FrameData[272]
rlabel metal3 5338 406708 5338 406708 0 FrameData[273]
rlabel metal3 9476 407435 9476 407435 0 FrameData[274]
rlabel metal3 9476 408183 9476 408183 0 FrameData[275]
rlabel metal3 9476 409299 9476 409299 0 FrameData[276]
rlabel metal3 9476 410047 9476 410047 0 FrameData[277]
rlabel metal3 5338 410788 5338 410788 0 FrameData[278]
rlabel metal3 9476 411515 9476 411515 0 FrameData[279]
rlabel metal2 18131 755820 18131 755820 0 FrameData[27]
rlabel metal3 9476 412263 9476 412263 0 FrameData[280]
rlabel metal3 9476 413379 9476 413379 0 FrameData[281]
rlabel metal3 9476 414127 9476 414127 0 FrameData[282]
rlabel metal3 5338 414868 5338 414868 0 FrameData[283]
rlabel metal3 9476 415595 9476 415595 0 FrameData[284]
rlabel metal3 9476 416343 9476 416343 0 FrameData[285]
rlabel metal3 9476 417459 9476 417459 0 FrameData[286]
rlabel metal3 2407 418268 2407 418268 0 FrameData[287]
rlabel metal3 3787 347548 3787 347548 0 FrameData[288]
rlabel metal3 9476 348419 9476 348419 0 FrameData[289]
rlabel metal2 9759 755820 9759 755820 0 FrameData[28]
rlabel metal3 9476 349535 9476 349535 0 FrameData[290]
rlabel metal3 5338 350268 5338 350268 0 FrameData[291]
rlabel metal3 9476 351003 9476 351003 0 FrameData[292]
rlabel metal3 3787 351628 3787 351628 0 FrameData[293]
rlabel metal3 9476 352867 9476 352867 0 FrameData[294]
rlabel metal3 9476 353615 9476 353615 0 FrameData[295]
rlabel metal3 5338 354348 5338 354348 0 FrameData[296]
rlabel metal3 9476 355083 9476 355083 0 FrameData[297]
rlabel metal3 9476 355831 9476 355831 0 FrameData[298]
rlabel metal3 9476 356947 9476 356947 0 FrameData[299]
rlabel metal2 12979 755820 12979 755820 0 FrameData[29]
rlabel metal3 16123 739228 16123 739228 0 FrameData[2]
rlabel metal3 9476 357695 9476 357695 0 FrameData[300]
rlabel metal3 5338 358428 5338 358428 0 FrameData[301]
rlabel metal3 9476 359163 9476 359163 0 FrameData[302]
rlabel metal3 9476 359911 9476 359911 0 FrameData[303]
rlabel metal3 9476 361027 9476 361027 0 FrameData[304]
rlabel metal3 9476 361775 9476 361775 0 FrameData[305]
rlabel metal3 5338 362508 5338 362508 0 FrameData[306]
rlabel metal3 9476 363243 9476 363243 0 FrameData[307]
rlabel metal3 9476 363991 9476 363991 0 FrameData[308]
rlabel metal3 9476 365107 9476 365107 0 FrameData[309]
rlabel metal4 21281 747660 21281 747660 0 FrameData[30]
rlabel metal3 9476 365855 9476 365855 0 FrameData[310]
rlabel metal3 5338 366588 5338 366588 0 FrameData[311]
rlabel metal3 9476 367323 9476 367323 0 FrameData[312]
rlabel metal3 9476 368071 9476 368071 0 FrameData[313]
rlabel metal3 9476 369187 9476 369187 0 FrameData[314]
rlabel metal3 9476 369935 9476 369935 0 FrameData[315]
rlabel metal3 5338 370668 5338 370668 0 FrameData[316]
rlabel metal3 9476 371403 9476 371403 0 FrameData[317]
rlabel metal3 9476 372151 9476 372151 0 FrameData[318]
rlabel metal3 9476 373267 9476 373267 0 FrameData[319]
rlabel metal2 9115 755820 9115 755820 0 FrameData[31]
rlabel metal3 9476 302731 9476 302731 0 FrameData[320]
rlabel metal3 3787 303348 3787 303348 0 FrameData[321]
rlabel metal3 9476 304606 9476 304606 0 FrameData[322]
rlabel metal3 9476 305354 9476 305354 0 FrameData[323]
rlabel metal3 5338 306068 5338 306068 0 FrameData[324]
rlabel metal3 9476 306811 9476 306811 0 FrameData[325]
rlabel metal3 9476 307559 9476 307559 0 FrameData[326]
rlabel metal3 9476 308686 9476 308686 0 FrameData[327]
rlabel metal3 9476 309434 9476 309434 0 FrameData[328]
rlabel metal3 5338 310148 5338 310148 0 FrameData[329]
rlabel metal3 2407 707948 2407 707948 0 FrameData[32]
rlabel metal3 9476 310891 9476 310891 0 FrameData[330]
rlabel metal3 9476 311639 9476 311639 0 FrameData[331]
rlabel metal3 9476 312766 9476 312766 0 FrameData[332]
rlabel metal3 9476 313514 9476 313514 0 FrameData[333]
rlabel metal3 5338 314228 5338 314228 0 FrameData[334]
rlabel metal3 9476 314971 9476 314971 0 FrameData[335]
rlabel metal3 9476 315719 9476 315719 0 FrameData[336]
rlabel metal3 9476 316846 9476 316846 0 FrameData[337]
rlabel metal3 9476 317594 9476 317594 0 FrameData[338]
rlabel metal3 5338 318308 5338 318308 0 FrameData[339]
rlabel metal3 5338 708628 5338 708628 0 FrameData[33]
rlabel metal3 9476 319051 9476 319051 0 FrameData[340]
rlabel metal3 9476 319799 9476 319799 0 FrameData[341]
rlabel metal3 9476 320926 9476 320926 0 FrameData[342]
rlabel metal3 9476 321674 9476 321674 0 FrameData[343]
rlabel metal3 5338 322388 5338 322388 0 FrameData[344]
rlabel metal3 9476 323131 9476 323131 0 FrameData[345]
rlabel metal3 9476 323879 9476 323879 0 FrameData[346]
rlabel metal3 9476 325006 9476 325006 0 FrameData[347]
rlabel metal3 2775 325788 2775 325788 0 FrameData[348]
rlabel metal3 5338 326468 5338 326468 0 FrameData[349]
rlabel metal3 3787 709308 3787 709308 0 FrameData[34]
rlabel metal3 9476 327211 9476 327211 0 FrameData[350]
rlabel metal3 9476 327959 9476 327959 0 FrameData[351]
rlabel metal3 5352 257788 5352 257788 0 FrameData[352]
rlabel metal3 3787 258468 3787 258468 0 FrameData[353]
rlabel metal3 3787 259148 3787 259148 0 FrameData[354]
rlabel metal3 3787 260508 3787 260508 0 FrameData[355]
rlabel metal3 9753 261120 9753 261120 0 FrameData[356]
rlabel metal3 5352 261868 5352 261868 0 FrameData[357]
rlabel metal3 3787 262548 3787 262548 0 FrameData[358]
rlabel metal3 3787 263228 3787 263228 0 FrameData[359]
rlabel metal3 9476 710115 9476 710115 0 FrameData[35]
rlabel metal3 3787 264588 3787 264588 0 FrameData[360]
rlabel metal3 9753 265200 9753 265200 0 FrameData[361]
rlabel metal3 5352 265948 5352 265948 0 FrameData[362]
rlabel metal3 3787 266628 3787 266628 0 FrameData[363]
rlabel metal3 3787 267308 3787 267308 0 FrameData[364]
rlabel metal3 3787 268668 3787 268668 0 FrameData[365]
rlabel metal3 9753 269280 9753 269280 0 FrameData[366]
rlabel metal3 5352 270028 5352 270028 0 FrameData[367]
rlabel metal3 3787 270708 3787 270708 0 FrameData[368]
rlabel metal3 3787 271388 3787 271388 0 FrameData[369]
rlabel metal3 9476 711231 9476 711231 0 FrameData[36]
rlabel metal3 3787 272748 3787 272748 0 FrameData[370]
rlabel metal3 9753 273360 9753 273360 0 FrameData[371]
rlabel metal3 5352 274108 5352 274108 0 FrameData[372]
rlabel metal3 3787 274788 3787 274788 0 FrameData[373]
rlabel metal3 3787 275468 3787 275468 0 FrameData[374]
rlabel metal3 3787 276828 3787 276828 0 FrameData[375]
rlabel metal3 2775 277508 2775 277508 0 FrameData[376]
rlabel metal3 5352 278188 5352 278188 0 FrameData[377]
rlabel metal3 3787 278868 3787 278868 0 FrameData[378]
rlabel metal3 3787 279548 3787 279548 0 FrameData[379]
rlabel metal3 9476 711979 9476 711979 0 FrameData[37]
rlabel metal3 3787 280908 3787 280908 0 FrameData[380]
rlabel metal3 2407 281588 2407 281588 0 FrameData[381]
rlabel metal3 5352 282268 5352 282268 0 FrameData[382]
rlabel metal3 3787 282948 3787 282948 0 FrameData[383]
rlabel metal3 3787 212228 3787 212228 0 FrameData[384]
rlabel metal3 5352 213588 5352 213588 0 FrameData[385]
rlabel metal3 3787 214268 3787 214268 0 FrameData[386]
rlabel metal3 3787 214948 3787 214948 0 FrameData[387]
rlabel metal3 9476 216211 9476 216211 0 FrameData[388]
rlabel metal3 9476 216959 9476 216959 0 FrameData[389]
rlabel metal3 5338 712708 5338 712708 0 FrameData[38]
rlabel metal3 5352 217668 5352 217668 0 FrameData[390]
rlabel metal3 3787 218348 3787 218348 0 FrameData[391]
rlabel metal3 3787 219028 3787 219028 0 FrameData[392]
rlabel metal3 9476 220291 9476 220291 0 FrameData[393]
rlabel metal3 9476 221039 9476 221039 0 FrameData[394]
rlabel metal3 5352 221748 5352 221748 0 FrameData[395]
rlabel metal3 3787 222428 3787 222428 0 FrameData[396]
rlabel metal3 3787 223108 3787 223108 0 FrameData[397]
rlabel metal3 9476 224371 9476 224371 0 FrameData[398]
rlabel metal3 9476 225119 9476 225119 0 FrameData[399]
rlabel metal3 3787 713388 3787 713388 0 FrameData[39]
rlabel metal3 20723 739500 20723 739500 0 FrameData[3]
rlabel metal3 5352 225828 5352 225828 0 FrameData[400]
rlabel metal3 3787 226508 3787 226508 0 FrameData[401]
rlabel metal3 3787 227188 3787 227188 0 FrameData[402]
rlabel metal3 9476 228451 9476 228451 0 FrameData[403]
rlabel metal3 9476 229199 9476 229199 0 FrameData[404]
rlabel metal3 5352 229908 5352 229908 0 FrameData[405]
rlabel metal3 3787 230588 3787 230588 0 FrameData[406]
rlabel metal3 3787 231268 3787 231268 0 FrameData[407]
rlabel metal3 9476 232531 9476 232531 0 FrameData[408]
rlabel metal3 2407 233308 2407 233308 0 FrameData[409]
rlabel metal3 9476 714195 9476 714195 0 FrameData[40]
rlabel metal3 5352 233988 5352 233988 0 FrameData[410]
rlabel metal3 3787 234668 3787 234668 0 FrameData[411]
rlabel metal3 3787 235348 3787 235348 0 FrameData[412]
rlabel metal3 9476 236611 9476 236611 0 FrameData[413]
rlabel metal3 2407 237388 2407 237388 0 FrameData[414]
rlabel metal3 5352 238068 5352 238068 0 FrameData[415]
rlabel metal3 9476 167939 9476 167939 0 FrameData[416]
rlabel metal3 9476 168687 9476 168687 0 FrameData[417]
rlabel metal3 9476 169407 9476 169407 0 FrameData[418]
rlabel metal3 9476 170155 9476 170155 0 FrameData[419]
rlabel metal3 9476 715311 9476 715311 0 FrameData[41]
rlabel metal3 9476 170903 9476 170903 0 FrameData[420]
rlabel metal3 9476 172019 9476 172019 0 FrameData[421]
rlabel metal3 9476 172767 9476 172767 0 FrameData[422]
rlabel metal3 9476 173487 9476 173487 0 FrameData[423]
rlabel metal3 9476 174235 9476 174235 0 FrameData[424]
rlabel metal3 9476 174983 9476 174983 0 FrameData[425]
rlabel metal3 9476 176099 9476 176099 0 FrameData[426]
rlabel metal3 9476 176847 9476 176847 0 FrameData[427]
rlabel metal3 9476 177567 9476 177567 0 FrameData[428]
rlabel metal3 9476 178315 9476 178315 0 FrameData[429]
rlabel metal3 9476 716059 9476 716059 0 FrameData[42]
rlabel metal3 9476 179063 9476 179063 0 FrameData[430]
rlabel metal3 9476 180179 9476 180179 0 FrameData[431]
rlabel metal3 9476 180927 9476 180927 0 FrameData[432]
rlabel metal3 9476 181647 9476 181647 0 FrameData[433]
rlabel metal3 9476 182395 9476 182395 0 FrameData[434]
rlabel metal3 9476 183143 9476 183143 0 FrameData[435]
rlabel metal3 9476 184259 9476 184259 0 FrameData[436]
rlabel metal3 9476 185007 9476 185007 0 FrameData[437]
rlabel metal3 9476 185727 9476 185727 0 FrameData[438]
rlabel metal3 9476 186475 9476 186475 0 FrameData[439]
rlabel metal3 5338 716788 5338 716788 0 FrameData[43]
rlabel metal3 9476 187223 9476 187223 0 FrameData[440]
rlabel metal3 9476 188339 9476 188339 0 FrameData[441]
rlabel metal3 2407 189108 2407 189108 0 FrameData[442]
rlabel metal3 9476 189807 9476 189807 0 FrameData[443]
rlabel metal3 9476 190555 9476 190555 0 FrameData[444]
rlabel metal3 9476 191303 9476 191303 0 FrameData[445]
rlabel metal3 9476 192419 9476 192419 0 FrameData[446]
rlabel metal3 9476 193167 9476 193167 0 FrameData[447]
rlabel metal3 3787 123148 3787 123148 0 FrameData[448]
rlabel metal3 9476 123747 9476 123747 0 FrameData[449]
rlabel metal3 3787 717468 3787 717468 0 FrameData[44]
rlabel metal3 9476 124495 9476 124495 0 FrameData[450]
rlabel metal3 9476 125215 9476 125215 0 FrameData[451]
rlabel metal3 9476 125963 9476 125963 0 FrameData[452]
rlabel metal3 2407 127228 2407 127228 0 FrameData[453]
rlabel metal3 9476 127827 9476 127827 0 FrameData[454]
rlabel metal3 9476 128575 9476 128575 0 FrameData[455]
rlabel metal3 9476 129295 9476 129295 0 FrameData[456]
rlabel metal3 9476 130043 9476 130043 0 FrameData[457]
rlabel metal3 2407 131308 2407 131308 0 FrameData[458]
rlabel metal3 9476 131907 9476 131907 0 FrameData[459]
rlabel metal3 9476 718275 9476 718275 0 FrameData[45]
rlabel metal3 9476 132655 9476 132655 0 FrameData[460]
rlabel metal3 9476 133375 9476 133375 0 FrameData[461]
rlabel metal3 9476 134123 9476 134123 0 FrameData[462]
rlabel metal3 2407 135388 2407 135388 0 FrameData[463]
rlabel metal3 9476 135987 9476 135987 0 FrameData[464]
rlabel metal3 9476 136735 9476 136735 0 FrameData[465]
rlabel metal3 9476 137455 9476 137455 0 FrameData[466]
rlabel metal3 9476 138203 9476 138203 0 FrameData[467]
rlabel metal3 2407 139468 2407 139468 0 FrameData[468]
rlabel metal3 9476 140067 9476 140067 0 FrameData[469]
rlabel metal3 9476 719391 9476 719391 0 FrameData[46]
rlabel metal3 9476 140815 9476 140815 0 FrameData[470]
rlabel metal3 9476 141535 9476 141535 0 FrameData[471]
rlabel metal3 9476 142283 9476 142283 0 FrameData[472]
rlabel metal3 2407 143548 2407 143548 0 FrameData[473]
rlabel metal3 9476 144147 9476 144147 0 FrameData[474]
rlabel metal3 9844 144892 9844 144892 0 FrameData[475]
rlabel metal3 9476 145615 9476 145615 0 FrameData[476]
rlabel metal3 3787 146268 3787 146268 0 FrameData[477]
rlabel metal3 9476 147479 9476 147479 0 FrameData[478]
rlabel metal3 9476 148227 9476 148227 0 FrameData[479]
rlabel metal3 9476 720139 9476 720139 0 FrameData[47]
rlabel metal3 1027 44268 1027 44268 0 FrameData[480]
rlabel metal3 4891 60588 4891 60588 0 FrameData[481]
rlabel metal3 2775 62628 2775 62628 0 FrameData[482]
rlabel metal3 644 68476 644 68476 0 FrameData[483]
rlabel metal3 9003 81124 9003 81124 0 FrameData[484]
rlabel metal3 1303 59908 1303 59908 0 FrameData[485]
rlabel metal3 2959 73508 2959 73508 0 FrameData[486]
rlabel metal3 3419 59228 3419 59228 0 FrameData[487]
rlabel metal3 4247 74868 4247 74868 0 FrameData[488]
rlabel metal3 1027 58548 1027 58548 0 FrameData[489]
rlabel metal3 5338 720868 5338 720868 0 FrameData[48]
rlabel metal3 2683 66708 2683 66708 0 FrameData[490]
rlabel metal3 3603 72828 3603 72828 0 FrameData[491]
rlabel metal3 2131 72148 2131 72148 0 FrameData[492]
rlabel metal3 1027 56508 1027 56508 0 FrameData[493]
rlabel metal3 552 75820 552 75820 0 FrameData[494]
rlabel metal3 4155 67388 4155 67388 0 FrameData[495]
rlabel metal3 3511 76228 3511 76228 0 FrameData[496]
rlabel metal3 3787 91868 3787 91868 0 FrameData[497]
rlabel metal3 5338 92548 5338 92548 0 FrameData[498]
rlabel metal3 9476 93262 9476 93262 0 FrameData[499]
rlabel metal3 9476 721607 9476 721607 0 FrameData[49]
rlabel metal3 19021 739772 19021 739772 0 FrameData[4]
rlabel metal3 9476 94010 9476 94010 0 FrameData[500]
rlabel metal3 2407 95268 2407 95268 0 FrameData[501]
rlabel metal3 3787 95948 3787 95948 0 FrameData[502]
rlabel metal3 5338 96628 5338 96628 0 FrameData[503]
rlabel metal3 9476 97342 9476 97342 0 FrameData[504]
rlabel metal3 9476 98090 9476 98090 0 FrameData[505]
rlabel metal3 3787 99348 3787 99348 0 FrameData[506]
rlabel metal3 3787 100028 3787 100028 0 FrameData[507]
rlabel metal3 5338 100708 5338 100708 0 FrameData[508]
rlabel metal3 9476 101422 9476 101422 0 FrameData[509]
rlabel metal3 9476 722355 9476 722355 0 FrameData[50]
rlabel metal3 3787 102068 3787 102068 0 FrameData[510]
rlabel metal3 9476 103287 9476 103287 0 FrameData[511]
rlabel metal3 4523 36788 4523 36788 0 FrameData[512]
rlabel metal3 3787 34068 3787 34068 0 FrameData[513]
rlabel metal3 2407 34748 2407 34748 0 FrameData[514]
rlabel metal3 3787 35428 3787 35428 0 FrameData[515]
rlabel metal3 5338 36108 5338 36108 0 FrameData[516]
rlabel metal3 2407 37468 2407 37468 0 FrameData[517]
rlabel metal3 3787 38148 3787 38148 0 FrameData[518]
rlabel metal3 2407 38828 2407 38828 0 FrameData[519]
rlabel metal3 9476 723471 9476 723471 0 FrameData[51]
rlabel metal3 3787 39508 3787 39508 0 FrameData[520]
rlabel metal3 5338 40188 5338 40188 0 FrameData[521]
rlabel metal3 9476 40902 9476 40902 0 FrameData[522]
rlabel metal3 9476 41650 9476 41650 0 FrameData[523]
rlabel metal3 9476 42398 9476 42398 0 FrameData[524]
rlabel metal3 9476 43146 9476 43146 0 FrameData[525]
rlabel metal3 3787 43588 3787 43588 0 FrameData[526]
rlabel metal3 9476 44982 9476 44982 0 FrameData[527]
rlabel metal3 9476 45730 9476 45730 0 FrameData[528]
rlabel metal3 9476 46478 9476 46478 0 FrameData[529]
rlabel metal3 9476 724219 9476 724219 0 FrameData[52]
rlabel metal3 9476 47226 9476 47226 0 FrameData[530]
rlabel metal3 3787 47668 3787 47668 0 FrameData[531]
rlabel metal3 9476 49062 9476 49062 0 FrameData[532]
rlabel metal3 9476 49810 9476 49810 0 FrameData[533]
rlabel metal3 9476 50558 9476 50558 0 FrameData[534]
rlabel metal3 9476 51306 9476 51306 0 FrameData[535]
rlabel metal3 9476 52054 9476 52054 0 FrameData[536]
rlabel metal3 9476 53142 9476 53142 0 FrameData[537]
rlabel metal3 3787 53788 3787 53788 0 FrameData[538]
rlabel metal3 9476 54638 9476 54638 0 FrameData[539]
rlabel metal3 5338 724948 5338 724948 0 FrameData[53]
rlabel metal3 3143 55148 3143 55148 0 FrameData[540]
rlabel metal3 9476 56134 9476 56134 0 FrameData[541]
rlabel metal3 9476 57222 9476 57222 0 FrameData[542]
rlabel metal3 3787 57868 3787 57868 0 FrameData[543]
rlabel metal2 22586 2183 22586 2183 0 FrameData[544]
rlabel metal2 21298 3831 21298 3831 0 FrameData[545]
rlabel metal2 20654 2115 20654 2115 0 FrameData[546]
rlabel metal2 21942 823 21942 823 0 FrameData[547]
rlabel metal3 7559 4828 7559 4828 0 FrameData[548]
rlabel metal4 15180 8160 15180 8160 0 FrameData[549]
rlabel metal3 9476 725687 9476 725687 0 FrameData[54]
rlabel via3 20355 7956 20355 7956 0 FrameData[550]
rlabel metal3 1027 748 1027 748 0 FrameData[551]
rlabel metal3 10963 9588 10963 9588 0 FrameData[552]
rlabel metal3 20608 9860 20608 9860 0 FrameData[553]
rlabel metal3 20700 10132 20700 10132 0 FrameData[554]
rlabel metal3 3787 10268 3787 10268 0 FrameData[555]
rlabel metal3 19320 10676 19320 10676 0 FrameData[556]
rlabel metal3 19228 10948 19228 10948 0 FrameData[557]
rlabel metal3 19872 11220 19872 11220 0 FrameData[558]
rlabel metal4 18860 11152 18860 11152 0 FrameData[559]
rlabel metal3 9476 726435 9476 726435 0 FrameData[55]
rlabel metal3 3787 8228 3787 8228 0 FrameData[560]
rlabel metal3 3787 11628 3787 11628 0 FrameData[561]
rlabel metal3 935 1428 935 1428 0 FrameData[562]
rlabel metal4 19596 10744 19596 10744 0 FrameData[563]
rlabel metal4 18860 12512 18860 12512 0 FrameData[564]
rlabel metal3 552 4420 552 4420 0 FrameData[565]
rlabel metal3 644 3060 644 3060 0 FrameData[566]
rlabel metal2 18906 13328 18906 13328 0 FrameData[567]
rlabel metal3 20700 13866 20700 13866 0 FrameData[568]
rlabel metal3 20700 14314 20700 14314 0 FrameData[569]
rlabel metal3 9476 727551 9476 727551 0 FrameData[56]
rlabel metal3 1027 33388 1027 33388 0 FrameData[570]
rlabel metal3 20700 14858 20700 14858 0 FrameData[571]
rlabel metal3 935 32708 935 32708 0 FrameData[572]
rlabel metal3 2775 17068 2775 17068 0 FrameData[573]
rlabel metal3 20700 15674 20700 15674 0 FrameData[574]
rlabel metal3 20700 16150 20700 16150 0 FrameData[575]
rlabel metal3 9476 728299 9476 728299 0 FrameData[57]
rlabel metal3 5338 729028 5338 729028 0 FrameData[58]
rlabel metal3 9476 729767 9476 729767 0 FrameData[59]
rlabel metal3 20884 740044 20884 740044 0 FrameData[5]
rlabel metal3 9476 730515 9476 730515 0 FrameData[60]
rlabel metal3 9476 731631 9476 731631 0 FrameData[61]
rlabel metal3 9476 732379 9476 732379 0 FrameData[62]
rlabel metal3 5338 733108 5338 733108 0 FrameData[63]
rlabel metal3 9476 662966 9476 662966 0 FrameData[64]
rlabel metal3 9476 663714 9476 663714 0 FrameData[65]
rlabel metal3 5338 664428 5338 664428 0 FrameData[66]
rlabel metal3 3787 665108 3787 665108 0 FrameData[67]
rlabel metal3 3787 665788 3787 665788 0 FrameData[68]
rlabel metal3 9476 667046 9476 667046 0 FrameData[69]
rlabel metal3 20677 740316 20677 740316 0 FrameData[6]
rlabel metal3 9476 667794 9476 667794 0 FrameData[70]
rlabel metal3 5338 668508 5338 668508 0 FrameData[71]
rlabel metal3 3787 669188 3787 669188 0 FrameData[72]
rlabel metal3 3787 669868 3787 669868 0 FrameData[73]
rlabel metal3 9476 671126 9476 671126 0 FrameData[74]
rlabel metal3 9476 671874 9476 671874 0 FrameData[75]
rlabel metal3 5338 672588 5338 672588 0 FrameData[76]
rlabel metal3 3787 673268 3787 673268 0 FrameData[77]
rlabel metal3 3787 673948 3787 673948 0 FrameData[78]
rlabel metal3 9476 675206 9476 675206 0 FrameData[79]
rlabel metal3 18699 740588 18699 740588 0 FrameData[7]
rlabel metal3 9476 675954 9476 675954 0 FrameData[80]
rlabel metal3 5338 676668 5338 676668 0 FrameData[81]
rlabel metal3 3787 677348 3787 677348 0 FrameData[82]
rlabel metal3 3787 678028 3787 678028 0 FrameData[83]
rlabel metal3 9476 679286 9476 679286 0 FrameData[84]
rlabel metal3 9476 680034 9476 680034 0 FrameData[85]
rlabel metal3 5338 680748 5338 680748 0 FrameData[86]
rlabel metal3 3787 681428 3787 681428 0 FrameData[87]
rlabel metal3 3787 682108 3787 682108 0 FrameData[88]
rlabel metal3 9476 683366 9476 683366 0 FrameData[89]
rlabel metal3 20861 740860 20861 740860 0 FrameData[8]
rlabel metal3 9476 684114 9476 684114 0 FrameData[90]
rlabel metal3 5338 684828 5338 684828 0 FrameData[91]
rlabel metal3 3787 685508 3787 685508 0 FrameData[92]
rlabel metal3 3787 686188 3787 686188 0 FrameData[93]
rlabel metal3 9476 687446 9476 687446 0 FrameData[94]
rlabel metal3 9476 688187 9476 688187 0 FrameData[95]
rlabel metal3 3787 617508 3787 617508 0 FrameData[96]
rlabel metal3 9476 618767 9476 618767 0 FrameData[97]
rlabel metal3 9476 619515 9476 619515 0 FrameData[98]
rlabel metal3 5341 620228 5341 620228 0 FrameData[99]
rlabel metal3 20815 741132 20815 741132 0 FrameData[9]
rlabel metal3 3442 32028 3442 32028 0 FrameStrobe[0]
rlabel metal2 218872 5897 218872 5897 0 FrameStrobe[100]
rlabel metal2 219608 5897 219608 5897 0 FrameStrobe[101]
rlabel metal2 220294 3271 220294 3271 0 FrameStrobe[102]
rlabel metal2 220938 3271 220938 3271 0 FrameStrobe[103]
rlabel metal2 221582 3271 221582 3271 0 FrameStrobe[104]
rlabel metal2 222552 5897 222552 5897 0 FrameStrobe[105]
rlabel metal2 223288 5897 223288 5897 0 FrameStrobe[106]
rlabel metal2 224024 5897 224024 5897 0 FrameStrobe[107]
rlabel metal2 224760 5897 224760 5897 0 FrameStrobe[108]
rlabel metal2 225446 3271 225446 3271 0 FrameStrobe[109]
rlabel metal3 4822 25228 4822 25228 0 FrameStrobe[10]
rlabel metal2 226090 3271 226090 3271 0 FrameStrobe[110]
rlabel metal2 226734 3271 226734 3271 0 FrameStrobe[111]
rlabel metal2 227704 5897 227704 5897 0 FrameStrobe[112]
rlabel metal2 228440 5897 228440 5897 0 FrameStrobe[113]
rlabel metal2 229176 5897 229176 5897 0 FrameStrobe[114]
rlabel metal2 229912 5897 229912 5897 0 FrameStrobe[115]
rlabel metal2 230598 3271 230598 3271 0 FrameStrobe[116]
rlabel metal2 231242 3271 231242 3271 0 FrameStrobe[117]
rlabel metal2 231886 3271 231886 3271 0 FrameStrobe[118]
rlabel metal2 232856 5897 232856 5897 0 FrameStrobe[119]
rlabel metal3 2752 31348 2752 31348 0 FrameStrobe[11]
rlabel metal2 259578 823 259578 823 0 FrameStrobe[120]
rlabel metal2 260636 5897 260636 5897 0 FrameStrobe[121]
rlabel metal2 261372 5897 261372 5897 0 FrameStrobe[122]
rlabel metal2 262108 5897 262108 5897 0 FrameStrobe[123]
rlabel metal2 262798 3388 262798 3388 0 FrameStrobe[124]
rlabel metal2 263442 1911 263442 1911 0 FrameStrobe[125]
rlabel metal2 264086 1231 264086 1231 0 FrameStrobe[126]
rlabel metal2 264730 3203 264730 3203 0 FrameStrobe[127]
rlabel metal2 265788 5897 265788 5897 0 FrameStrobe[128]
rlabel metal2 266524 5897 266524 5897 0 FrameStrobe[129]
rlabel metal2 16974 16894 16974 16894 0 FrameStrobe[12]
rlabel metal2 267260 5897 267260 5897 0 FrameStrobe[130]
rlabel metal2 267950 3388 267950 3388 0 FrameStrobe[131]
rlabel metal2 268594 1911 268594 1911 0 FrameStrobe[132]
rlabel metal2 269238 1231 269238 1231 0 FrameStrobe[133]
rlabel metal2 269882 823 269882 823 0 FrameStrobe[134]
rlabel metal2 270940 5897 270940 5897 0 FrameStrobe[135]
rlabel metal2 271676 5897 271676 5897 0 FrameStrobe[136]
rlabel metal2 272412 5897 272412 5897 0 FrameStrobe[137]
rlabel metal2 273102 3388 273102 3388 0 FrameStrobe[138]
rlabel metal2 273746 1911 273746 1911 0 FrameStrobe[139]
rlabel metal2 17434 17098 17434 17098 0 FrameStrobe[13]
rlabel metal2 278898 1027 278898 1027 0 FrameStrobe[140]
rlabel metal2 280830 3388 280830 3388 0 FrameStrobe[141]
rlabel metal2 282932 5897 282932 5897 0 FrameStrobe[142]
rlabel metal2 285338 823 285338 823 0 FrameStrobe[143]
rlabel metal2 287270 1911 287270 1911 0 FrameStrobe[144]
rlabel metal2 289280 5897 289280 5897 0 FrameStrobe[145]
rlabel metal2 291396 5897 291396 5897 0 FrameStrobe[146]
rlabel metal2 293710 1911 293710 1911 0 FrameStrobe[147]
rlabel metal2 295642 3388 295642 3388 0 FrameStrobe[148]
rlabel metal2 297744 5897 297744 5897 0 FrameStrobe[149]
rlabel metal2 17848 17163 17848 17163 0 FrameStrobe[14]
rlabel metal2 300150 823 300150 823 0 FrameStrobe[150]
rlabel metal2 302082 959 302082 959 0 FrameStrobe[151]
rlabel metal2 304092 5897 304092 5897 0 FrameStrobe[152]
rlabel metal2 306222 3381 306222 3381 0 FrameStrobe[153]
rlabel metal2 308522 1911 308522 1911 0 FrameStrobe[154]
rlabel metal2 310454 3388 310454 3388 0 FrameStrobe[155]
rlabel metal2 312556 5897 312556 5897 0 FrameStrobe[156]
rlabel metal2 314962 823 314962 823 0 FrameStrobe[157]
rlabel metal2 316894 1911 316894 1911 0 FrameStrobe[158]
rlabel metal2 318904 5897 318904 5897 0 FrameStrobe[159]
rlabel metal2 18354 17115 18354 17115 0 FrameStrobe[15]
rlabel metal2 345874 3388 345874 3388 0 FrameStrobe[160]
rlabel metal2 346608 5897 346608 5897 0 FrameStrobe[161]
rlabel metal2 347344 5897 347344 5897 0 FrameStrobe[162]
rlabel metal2 348082 3381 348082 3381 0 FrameStrobe[163]
rlabel metal2 349094 823 349094 823 0 FrameStrobe[164]
rlabel metal2 349738 1911 349738 1911 0 FrameStrobe[165]
rlabel metal2 350382 1911 350382 1911 0 FrameStrobe[166]
rlabel metal2 351026 3388 351026 3388 0 FrameStrobe[167]
rlabel metal2 351760 5897 351760 5897 0 FrameStrobe[168]
rlabel metal2 352496 5897 352496 5897 0 FrameStrobe[169]
rlabel metal3 18124 17340 18124 17340 0 FrameStrobe[16]
rlabel metal2 353234 3381 353234 3381 0 FrameStrobe[170]
rlabel metal2 354246 823 354246 823 0 FrameStrobe[171]
rlabel metal2 354890 1911 354890 1911 0 FrameStrobe[172]
rlabel metal2 355534 1911 355534 1911 0 FrameStrobe[173]
rlabel metal2 356178 3388 356178 3388 0 FrameStrobe[174]
rlabel metal2 356912 5897 356912 5897 0 FrameStrobe[175]
rlabel metal2 357648 5897 357648 5897 0 FrameStrobe[176]
rlabel metal2 358386 3381 358386 3381 0 FrameStrobe[177]
rlabel metal2 359398 823 359398 823 0 FrameStrobe[178]
rlabel metal2 360042 1911 360042 1911 0 FrameStrobe[179]
rlabel metal2 19274 17081 19274 17081 0 FrameStrobe[17]
rlabel metal2 380064 5897 380064 5897 0 FrameStrobe[180]
rlabel metal2 386998 544 386998 544 0 FrameStrobe[181]
rlabel metal2 388286 680 388286 680 0 FrameStrobe[182]
rlabel metal2 392886 3271 392886 3271 0 FrameStrobe[183]
rlabel metal2 384480 5897 384480 5897 0 FrameStrobe[184]
rlabel metal2 385584 5897 385584 5897 0 FrameStrobe[185]
rlabel metal2 386688 5897 386688 5897 0 FrameStrobe[186]
rlabel metal2 387792 5897 387792 5897 0 FrameStrobe[187]
rlabel metal2 388896 5897 388896 5897 0 FrameStrobe[188]
rlabel metal2 390000 5897 390000 5897 0 FrameStrobe[189]
rlabel metal2 19734 17047 19734 17047 0 FrameStrobe[18]
rlabel metal2 391104 5897 391104 5897 0 FrameStrobe[190]
rlabel metal2 392208 5897 392208 5897 0 FrameStrobe[191]
rlabel metal2 393312 5897 393312 5897 0 FrameStrobe[192]
rlabel metal2 394416 5897 394416 5897 0 FrameStrobe[193]
rlabel metal2 395462 3271 395462 3271 0 FrameStrobe[194]
rlabel metal2 396624 5897 396624 5897 0 FrameStrobe[195]
rlabel metal2 397728 5897 397728 5897 0 FrameStrobe[196]
rlabel metal2 398682 3271 398682 3271 0 FrameStrobe[197]
rlabel metal2 399936 5897 399936 5897 0 FrameStrobe[198]
rlabel metal2 401040 5897 401040 5897 0 FrameStrobe[199]
rlabel metal2 20148 17146 20148 17146 0 FrameStrobe[19]
rlabel metal3 2798 29308 2798 29308 0 FrameStrobe[1]
rlabel metal2 415820 5897 415820 5897 0 FrameStrobe[200]
rlabel metal2 417200 5897 417200 5897 0 FrameStrobe[201]
rlabel metal2 418580 5897 418580 5897 0 FrameStrobe[202]
rlabel metal2 419960 5897 419960 5897 0 FrameStrobe[203]
rlabel metal2 421340 5897 421340 5897 0 FrameStrobe[204]
rlabel metal2 422720 5897 422720 5897 0 FrameStrobe[205]
rlabel metal2 424100 5897 424100 5897 0 FrameStrobe[206]
rlabel metal2 425480 5897 425480 5897 0 FrameStrobe[207]
rlabel metal2 426860 5897 426860 5897 0 FrameStrobe[208]
rlabel metal2 428240 5897 428240 5897 0 FrameStrobe[209]
rlabel metal2 30958 1911 30958 1911 0 FrameStrobe[20]
rlabel metal2 429620 5897 429620 5897 0 FrameStrobe[210]
rlabel metal2 431000 5897 431000 5897 0 FrameStrobe[211]
rlabel metal2 432380 5897 432380 5897 0 FrameStrobe[212]
rlabel metal2 433760 5897 433760 5897 0 FrameStrobe[213]
rlabel metal2 435140 5897 435140 5897 0 FrameStrobe[214]
rlabel metal2 436520 5897 436520 5897 0 FrameStrobe[215]
rlabel metal2 437900 5897 437900 5897 0 FrameStrobe[216]
rlabel metal2 439280 5897 439280 5897 0 FrameStrobe[217]
rlabel metal2 440660 5897 440660 5897 0 FrameStrobe[218]
rlabel metal2 442040 5897 442040 5897 0 FrameStrobe[219]
rlabel metal2 32336 5897 32336 5897 0 FrameStrobe[21]
rlabel metal2 446338 823 446338 823 0 FrameStrobe[220]
rlabel metal2 447626 3388 447626 3388 0 FrameStrobe[221]
rlabel metal2 449190 3381 449190 3381 0 FrameStrobe[222]
rlabel metal2 450846 1911 450846 1911 0 FrameStrobe[223]
rlabel metal2 452312 5897 452312 5897 0 FrameStrobe[224]
rlabel metal2 454066 1027 454066 1027 0 FrameStrobe[225]
rlabel metal2 455440 5897 455440 5897 0 FrameStrobe[226]
rlabel metal2 457286 823 457286 823 0 FrameStrobe[227]
rlabel metal2 458574 3388 458574 3388 0 FrameStrobe[228]
rlabel metal2 460138 3381 460138 3381 0 FrameStrobe[229]
rlabel metal2 34178 823 34178 823 0 FrameStrobe[22]
rlabel metal2 461794 1911 461794 1911 0 FrameStrobe[230]
rlabel metal2 463260 5897 463260 5897 0 FrameStrobe[231]
rlabel metal2 465014 1911 465014 1911 0 FrameStrobe[232]
rlabel metal2 466388 5897 466388 5897 0 FrameStrobe[233]
rlabel metal2 468234 823 468234 823 0 FrameStrobe[234]
rlabel metal2 469522 3388 469522 3388 0 FrameStrobe[235]
rlabel metal2 471086 3381 471086 3381 0 FrameStrobe[236]
rlabel metal2 472742 1911 472742 1911 0 FrameStrobe[237]
rlabel metal2 474208 5897 474208 5897 0 FrameStrobe[238]
rlabel metal2 475962 1911 475962 1911 0 FrameStrobe[239]
rlabel metal2 35466 3388 35466 3388 0 FrameStrobe[23]
rlabel metal2 37030 3381 37030 3381 0 FrameStrobe[24]
rlabel metal2 38686 1027 38686 1027 0 FrameStrobe[25]
rlabel metal2 40156 5897 40156 5897 0 FrameStrobe[26]
rlabel metal2 41906 1911 41906 1911 0 FrameStrobe[27]
rlabel metal2 43284 5897 43284 5897 0 FrameStrobe[28]
rlabel metal2 45126 823 45126 823 0 FrameStrobe[29]
rlabel metal2 9522 18360 9522 18360 0 FrameStrobe[2]
rlabel metal2 46414 3388 46414 3388 0 FrameStrobe[30]
rlabel metal2 47978 3381 47978 3381 0 FrameStrobe[31]
rlabel metal2 49634 1911 49634 1911 0 FrameStrobe[32]
rlabel metal2 51104 5897 51104 5897 0 FrameStrobe[33]
rlabel metal2 52854 1911 52854 1911 0 FrameStrobe[34]
rlabel metal2 54232 5897 54232 5897 0 FrameStrobe[35]
rlabel metal2 56074 823 56074 823 0 FrameStrobe[36]
rlabel metal2 57362 3388 57362 3388 0 FrameStrobe[37]
rlabel metal2 58926 3381 58926 3381 0 FrameStrobe[38]
rlabel metal2 60582 1911 60582 1911 0 FrameStrobe[39]
rlabel metal3 3695 18428 3695 18428 0 FrameStrobe[3]
rlabel metal2 73888 5897 73888 5897 0 FrameStrobe[40]
rlabel metal2 75360 5897 75360 5897 0 FrameStrobe[41]
rlabel metal2 76682 3271 76682 3271 0 FrameStrobe[42]
rlabel metal2 78304 5897 78304 5897 0 FrameStrobe[43]
rlabel metal2 79776 5897 79776 5897 0 FrameStrobe[44]
rlabel metal2 81190 3271 81190 3271 0 FrameStrobe[45]
rlabel metal2 82478 3271 82478 3271 0 FrameStrobe[46]
rlabel metal2 84192 5897 84192 5897 0 FrameStrobe[47]
rlabel metal2 85664 5897 85664 5897 0 FrameStrobe[48]
rlabel metal2 86986 3271 86986 3271 0 FrameStrobe[49]
rlabel metal3 3787 17748 3787 17748 0 FrameStrobe[4]
rlabel metal2 88608 5897 88608 5897 0 FrameStrobe[50]
rlabel metal2 90080 5897 90080 5897 0 FrameStrobe[51]
rlabel metal2 91494 3271 91494 3271 0 FrameStrobe[52]
rlabel metal2 92782 3271 92782 3271 0 FrameStrobe[53]
rlabel metal2 94496 5897 94496 5897 0 FrameStrobe[54]
rlabel metal2 95968 5897 95968 5897 0 FrameStrobe[55]
rlabel metal2 97290 3271 97290 3271 0 FrameStrobe[56]
rlabel metal2 98912 5897 98912 5897 0 FrameStrobe[57]
rlabel metal2 100384 5897 100384 5897 0 FrameStrobe[58]
rlabel metal2 101798 3271 101798 3271 0 FrameStrobe[59]
rlabel metal3 1027 25908 1027 25908 0 FrameStrobe[5]
rlabel metal2 106976 5897 106976 5897 0 FrameStrobe[60]
rlabel metal2 109276 5897 109276 5897 0 FrameStrobe[61]
rlabel metal2 111576 5897 111576 5897 0 FrameStrobe[62]
rlabel metal2 113876 5897 113876 5897 0 FrameStrobe[63]
rlabel metal2 116176 5897 116176 5897 0 FrameStrobe[64]
rlabel metal2 118476 5897 118476 5897 0 FrameStrobe[65]
rlabel metal2 120776 5897 120776 5897 0 FrameStrobe[66]
rlabel metal2 123076 5897 123076 5897 0 FrameStrobe[67]
rlabel metal2 125376 5897 125376 5897 0 FrameStrobe[68]
rlabel metal2 127676 5897 127676 5897 0 FrameStrobe[69]
rlabel metal3 3120 23188 3120 23188 0 FrameStrobe[6]
rlabel metal2 129976 5897 129976 5897 0 FrameStrobe[70]
rlabel metal2 132276 5897 132276 5897 0 FrameStrobe[71]
rlabel metal2 134576 5897 134576 5897 0 FrameStrobe[72]
rlabel metal2 136876 5897 136876 5897 0 FrameStrobe[73]
rlabel metal2 139176 5897 139176 5897 0 FrameStrobe[74]
rlabel metal2 141476 5897 141476 5897 0 FrameStrobe[75]
rlabel metal2 143776 5897 143776 5897 0 FrameStrobe[76]
rlabel metal2 146076 5897 146076 5897 0 FrameStrobe[77]
rlabel metal2 148376 5897 148376 5897 0 FrameStrobe[78]
rlabel metal2 150742 3271 150742 3271 0 FrameStrobe[79]
rlabel metal3 912 30668 912 30668 0 FrameStrobe[7]
rlabel metal2 177872 5897 177872 5897 0 FrameStrobe[80]
rlabel metal2 178608 5897 178608 5897 0 FrameStrobe[81]
rlabel metal2 179354 3381 179354 3381 0 FrameStrobe[82]
rlabel metal2 180366 823 180366 823 0 FrameStrobe[83]
rlabel metal2 181010 1911 181010 1911 0 FrameStrobe[84]
rlabel metal2 181654 1911 181654 1911 0 FrameStrobe[85]
rlabel metal2 182298 3388 182298 3388 0 FrameStrobe[86]
rlabel metal2 183024 5897 183024 5897 0 FrameStrobe[87]
rlabel metal2 183760 5897 183760 5897 0 FrameStrobe[88]
rlabel metal2 184506 3381 184506 3381 0 FrameStrobe[89]
rlabel metal1 11385 17238 11385 17238 0 FrameStrobe[8]
rlabel metal2 185518 823 185518 823 0 FrameStrobe[90]
rlabel metal2 186162 1911 186162 1911 0 FrameStrobe[91]
rlabel metal2 186806 1911 186806 1911 0 FrameStrobe[92]
rlabel metal2 187450 3388 187450 3388 0 FrameStrobe[93]
rlabel metal2 188176 5897 188176 5897 0 FrameStrobe[94]
rlabel metal2 188912 5897 188912 5897 0 FrameStrobe[95]
rlabel metal2 189658 3381 189658 3381 0 FrameStrobe[96]
rlabel metal2 190670 823 190670 823 0 FrameStrobe[97]
rlabel metal2 191314 1911 191314 1911 0 FrameStrobe[98]
rlabel metal2 191958 1095 191958 1095 0 FrameStrobe[99]
rlabel metal3 2062 23868 2062 23868 0 FrameStrobe[9]
rlabel metal3 9476 292366 9476 292366 0 Tile_X0Y10_A_I_top
rlabel metal3 3787 291108 3787 291108 0 Tile_X0Y10_A_O_top
rlabel metal3 9476 293114 9476 293114 0 Tile_X0Y10_A_T_top
rlabel metal3 9476 296446 9476 296446 0 Tile_X0Y10_A_config_C_bit0
rlabel metal3 9476 297194 9476 297194 0 Tile_X0Y10_A_config_C_bit1
rlabel metal3 5338 297908 5338 297908 0 Tile_X0Y10_A_config_C_bit2
rlabel metal3 9476 298651 9476 298651 0 Tile_X0Y10_A_config_C_bit3
rlabel metal3 9476 294571 9476 294571 0 Tile_X0Y10_B_I_top
rlabel metal3 5338 293828 5338 293828 0 Tile_X0Y10_B_O_top
rlabel metal3 3787 295188 3787 295188 0 Tile_X0Y10_B_T_top
rlabel metal3 3787 299268 3787 299268 0 Tile_X0Y10_B_config_C_bit0
rlabel metal3 9476 300526 9476 300526 0 Tile_X0Y10_B_config_C_bit1
rlabel metal3 9476 301274 9476 301274 0 Tile_X0Y10_B_config_C_bit2
rlabel metal3 5338 301988 5338 301988 0 Tile_X0Y10_B_config_C_bit3
rlabel metal3 3787 246908 3787 246908 0 Tile_X0Y11_A_I_top
rlabel metal3 9476 246299 9476 246299 0 Tile_X0Y11_A_O_top
rlabel metal3 3787 248268 3787 248268 0 Tile_X0Y11_A_T_top
rlabel metal3 3787 250988 3787 250988 0 Tile_X0Y11_A_config_C_bit0
rlabel metal3 3787 252348 3787 252348 0 Tile_X0Y11_A_config_C_bit1
rlabel metal3 9753 252960 9753 252960 0 Tile_X0Y11_A_config_C_bit2
rlabel metal3 5352 253708 5352 253708 0 Tile_X0Y11_A_config_C_bit3
rlabel metal3 5352 249628 5352 249628 0 Tile_X0Y11_B_I_top
rlabel metal3 9753 248880 9753 248880 0 Tile_X0Y11_B_O_top
rlabel metal3 3787 250308 3787 250308 0 Tile_X0Y11_B_T_top
rlabel metal3 3787 254388 3787 254388 0 Tile_X0Y11_B_config_C_bit0
rlabel metal3 3787 255068 3787 255068 0 Tile_X0Y11_B_config_C_bit1
rlabel metal3 3787 256428 3787 256428 0 Tile_X0Y11_B_config_C_bit2
rlabel metal3 9753 257040 9753 257040 0 Tile_X0Y11_B_config_C_bit3
rlabel metal3 3787 202028 3787 202028 0 Tile_X0Y12_A_I_top
rlabel metal3 9476 201359 9476 201359 0 Tile_X0Y12_A_O_top
rlabel metal3 3787 202708 3787 202708 0 Tile_X0Y12_A_T_top
rlabel metal3 3787 206108 3787 206108 0 Tile_X0Y12_A_config_C_bit0
rlabel metal3 3787 206788 3787 206788 0 Tile_X0Y12_A_config_C_bit1
rlabel metal3 9476 208051 9476 208051 0 Tile_X0Y12_A_config_C_bit2
rlabel metal3 9476 208799 9476 208799 0 Tile_X0Y12_A_config_C_bit3
rlabel metal3 9476 204719 9476 204719 0 Tile_X0Y12_B_I_top
rlabel metal3 9476 203971 9476 203971 0 Tile_X0Y12_B_O_top
rlabel metal3 5352 205428 5352 205428 0 Tile_X0Y12_B_T_top
rlabel metal3 5352 209508 5352 209508 0 Tile_X0Y12_B_config_C_bit0
rlabel metal3 3787 210188 3787 210188 0 Tile_X0Y12_B_config_C_bit1
rlabel metal3 3787 210868 3787 210868 0 Tile_X0Y12_B_config_C_bit2
rlabel metal3 3787 211548 3787 211548 0 Tile_X0Y12_B_config_C_bit3
rlabel metal3 9476 157167 9476 157167 0 Tile_X0Y13_A_I_top
rlabel metal3 9476 156447 9476 156447 0 Tile_X0Y13_A_O_top
rlabel metal3 9476 157915 9476 157915 0 Tile_X0Y13_A_T_top
rlabel metal3 9476 161247 9476 161247 0 Tile_X0Y13_A_config_C_bit0
rlabel metal3 9476 161995 9476 161995 0 Tile_X0Y13_A_config_C_bit1
rlabel metal3 3787 162588 3787 162588 0 Tile_X0Y13_A_config_C_bit2
rlabel metal3 9476 163859 9476 163859 0 Tile_X0Y13_A_config_C_bit3
rlabel metal3 9476 159779 9476 159779 0 Tile_X0Y13_B_I_top
rlabel metal3 3787 158508 3787 158508 0 Tile_X0Y13_B_O_top
rlabel metal3 9476 160527 9476 160527 0 Tile_X0Y13_B_T_top
rlabel metal3 9476 164607 9476 164607 0 Tile_X0Y13_B_config_C_bit0
rlabel metal3 9476 165327 9476 165327 0 Tile_X0Y13_B_config_C_bit1
rlabel metal3 9476 166075 9476 166075 0 Tile_X0Y13_B_config_C_bit2
rlabel metal3 3787 166668 3787 166668 0 Tile_X0Y13_B_config_C_bit3
rlabel metal3 9476 112255 9476 112255 0 Tile_X0Y14_A_I_top
rlabel metal3 9476 111507 9476 111507 0 Tile_X0Y14_A_O_top
rlabel metal3 9476 112975 9476 112975 0 Tile_X0Y14_A_T_top
rlabel metal3 9476 116335 9476 116335 0 Tile_X0Y14_A_config_C_bit0
rlabel metal3 9476 117055 9476 117055 0 Tile_X0Y14_A_config_C_bit1
rlabel metal3 9476 117803 9476 117803 0 Tile_X0Y14_A_config_C_bit2
rlabel metal3 9476 118919 9476 118919 0 Tile_X0Y14_A_config_C_bit3
rlabel metal3 9476 114839 9476 114839 0 Tile_X0Y14_B_I_top
rlabel metal3 9476 113723 9476 113723 0 Tile_X0Y14_B_O_top
rlabel metal3 9476 115587 9476 115587 0 Tile_X0Y14_B_T_top
rlabel metal3 9476 119667 9476 119667 0 Tile_X0Y14_B_config_C_bit0
rlabel metal3 9476 120415 9476 120415 0 Tile_X0Y14_B_config_C_bit1
rlabel metal3 9476 121135 9476 121135 0 Tile_X0Y14_B_config_C_bit2
rlabel metal3 9476 121883 9476 121883 0 Tile_X0Y14_B_config_C_bit3
rlabel metal3 3143 66028 3143 66028 0 Tile_X0Y15_A_I_top
rlabel metal3 2131 52428 2131 52428 0 Tile_X0Y15_A_O_top
rlabel metal3 4983 64668 4983 64668 0 Tile_X0Y15_A_T_top
rlabel metal3 9476 71026 9476 71026 0 Tile_X0Y15_A_config_C_bit0
rlabel metal3 3695 63988 3695 63988 0 Tile_X0Y15_A_config_C_bit1
rlabel metal3 2407 65348 2407 65348 0 Tile_X0Y15_A_config_C_bit2
rlabel metal3 4247 63308 4247 63308 0 Tile_X0Y15_A_config_C_bit3
rlabel metal3 9476 69530 9476 69530 0 Tile_X0Y15_B_I_top
rlabel metal3 1395 48348 1395 48348 0 Tile_X0Y15_B_O_top
rlabel metal3 9476 70278 9476 70278 0 Tile_X0Y15_B_T_top
rlabel metal3 3511 61948 3511 61948 0 Tile_X0Y15_B_config_C_bit0
rlabel metal3 9187 75412 9187 75412 0 Tile_X0Y15_B_config_C_bit1
rlabel metal3 751 61268 751 61268 0 Tile_X0Y15_B_config_C_bit2
rlabel metal3 2867 68068 2867 68068 0 Tile_X0Y15_B_config_C_bit3
rlabel metal3 2407 24548 2407 24548 0 Tile_X0Y16_A_I_top
rlabel metal3 3787 21828 3787 21828 0 Tile_X0Y16_A_O_top
rlabel metal2 6486 11907 6486 11907 0 Tile_X0Y16_A_T_top
rlabel metal2 10350 1027 10350 1027 0 Tile_X0Y16_A_config_C_bit0
rlabel metal2 12282 891 12282 891 0 Tile_X0Y16_A_config_C_bit1
rlabel metal2 13570 823 13570 823 0 Tile_X0Y16_A_config_C_bit2
rlabel metal2 10994 959 10994 959 0 Tile_X0Y16_A_config_C_bit3
rlabel metal3 9532 24684 9532 24684 0 Tile_X0Y16_B_I_top
rlabel metal3 8888 23868 8888 23868 0 Tile_X0Y16_B_O_top
rlabel metal2 11638 3203 11638 3203 0 Tile_X0Y16_B_T_top
rlabel metal2 9706 1027 9706 1027 0 Tile_X0Y16_B_config_C_bit0
rlabel metal2 12926 2455 12926 2455 0 Tile_X0Y16_B_config_C_bit1
rlabel metal3 8566 31212 8566 31212 0 Tile_X0Y16_B_config_C_bit2
rlabel metal2 8418 1027 8418 1027 0 Tile_X0Y16_B_config_C_bit3
rlabel metal3 9476 697127 9476 697127 0 Tile_X0Y1_A_I_top
rlabel metal3 5338 696388 5338 696388 0 Tile_X0Y1_A_O_top
rlabel metal3 9476 697875 9476 697875 0 Tile_X0Y1_A_T_top
rlabel metal3 9476 701207 9476 701207 0 Tile_X0Y1_A_config_C_bit0
rlabel metal3 9476 701955 9476 701955 0 Tile_X0Y1_A_config_C_bit1
rlabel metal3 9476 703071 9476 703071 0 Tile_X0Y1_A_config_C_bit2
rlabel metal3 2407 703868 2407 703868 0 Tile_X0Y1_A_config_C_bit3
rlabel metal3 2407 699788 2407 699788 0 Tile_X0Y1_B_I_top
rlabel metal3 9476 698991 9476 698991 0 Tile_X0Y1_B_O_top
rlabel metal3 5338 700468 5338 700468 0 Tile_X0Y1_B_T_top
rlabel metal3 5338 704548 5338 704548 0 Tile_X0Y1_B_config_C_bit0
rlabel metal3 9476 705287 9476 705287 0 Tile_X0Y1_B_config_C_bit1
rlabel metal3 9476 706035 9476 706035 0 Tile_X0Y1_B_config_C_bit2
rlabel metal3 9476 707151 9476 707151 0 Tile_X0Y1_B_config_C_bit3
rlabel metal3 5338 652188 5338 652188 0 Tile_X0Y2_A_I_top
rlabel metal3 9476 651474 9476 651474 0 Tile_X0Y2_A_O_top
rlabel metal3 3787 652868 3787 652868 0 Tile_X0Y2_A_T_top
rlabel metal3 5338 656268 5338 656268 0 Tile_X0Y2_A_config_C_bit0
rlabel metal3 3787 656948 3787 656948 0 Tile_X0Y2_A_config_C_bit1
rlabel metal3 3787 657628 3787 657628 0 Tile_X0Y2_A_config_C_bit2
rlabel metal3 9476 658886 9476 658886 0 Tile_X0Y2_A_config_C_bit3
rlabel metal3 9476 654806 9476 654806 0 Tile_X0Y2_B_I_top
rlabel metal3 3787 653548 3787 653548 0 Tile_X0Y2_B_O_top
rlabel metal3 2407 655588 2407 655588 0 Tile_X0Y2_B_T_top
rlabel metal3 2407 659668 2407 659668 0 Tile_X0Y2_B_config_C_bit0
rlabel metal3 5338 660348 5338 660348 0 Tile_X0Y2_B_config_C_bit1
rlabel metal3 3787 661028 3787 661028 0 Tile_X0Y2_B_config_C_bit2
rlabel metal3 3787 661708 3787 661708 0 Tile_X0Y2_B_config_C_bit3
rlabel metal3 2407 607308 2407 607308 0 Tile_X0Y3_A_I_top
rlabel metal3 9476 606526 9476 606526 0 Tile_X0Y3_A_O_top
rlabel metal3 5341 607988 5341 607988 0 Tile_X0Y3_A_T_top
rlabel metal3 2407 611388 2407 611388 0 Tile_X0Y3_A_config_C_bit0
rlabel metal3 5341 612068 5341 612068 0 Tile_X0Y3_A_config_C_bit1
rlabel metal3 3787 612748 3787 612748 0 Tile_X0Y3_A_config_C_bit2
rlabel metal3 3787 613428 3787 613428 0 Tile_X0Y3_A_config_C_bit3
rlabel metal3 3787 609348 3787 609348 0 Tile_X0Y3_B_I_top
rlabel metal3 3787 608668 3787 608668 0 Tile_X0Y3_B_O_top
rlabel metal3 9476 610607 9476 610607 0 Tile_X0Y3_B_T_top
rlabel metal3 9476 614687 9476 614687 0 Tile_X0Y3_B_config_C_bit0
rlabel metal3 9476 615435 9476 615435 0 Tile_X0Y3_B_config_C_bit1
rlabel metal3 5341 616148 5341 616148 0 Tile_X0Y3_B_config_C_bit2
rlabel metal3 3787 616828 3787 616828 0 Tile_X0Y3_B_config_C_bit3
rlabel metal3 9476 562335 9476 562335 0 Tile_X0Y4_A_I_top
rlabel metal3 9476 561219 9476 561219 0 Tile_X0Y4_A_O_top
rlabel metal3 2407 563108 2407 563108 0 Tile_X0Y4_A_T_top
rlabel metal3 9476 566415 9476 566415 0 Tile_X0Y4_A_config_C_bit0
rlabel metal3 2775 567188 2775 567188 0 Tile_X0Y4_A_config_C_bit1
rlabel metal3 9476 567883 9476 567883 0 Tile_X0Y4_A_config_C_bit2
rlabel metal3 3787 568548 3787 568548 0 Tile_X0Y4_A_config_C_bit3
rlabel metal3 9476 564551 9476 564551 0 Tile_X0Y4_B_I_top
rlabel metal3 9476 563803 9476 563803 0 Tile_X0Y4_B_O_top
rlabel metal3 9476 565299 9476 565299 0 Tile_X0Y4_B_T_top
rlabel metal3 9476 569379 9476 569379 0 Tile_X0Y4_B_config_C_bit0
rlabel metal3 9476 570495 9476 570495 0 Tile_X0Y4_B_config_C_bit1
rlabel metal3 9476 571243 9476 571243 0 Tile_X0Y4_B_config_C_bit2
rlabel metal3 9476 571963 9476 571963 0 Tile_X0Y4_B_config_C_bit3
rlabel metal3 2407 517548 2407 517548 0 Tile_X0Y5_A_I_top
rlabel metal3 9476 516279 9476 516279 0 Tile_X0Y5_A_O_top
rlabel metal3 9476 518143 9476 518143 0 Tile_X0Y5_A_T_top
rlabel metal3 9476 521475 9476 521475 0 Tile_X0Y5_A_config_C_bit0
rlabel metal3 9476 522223 9476 522223 0 Tile_X0Y5_A_config_C_bit1
rlabel metal3 9476 522971 9476 522971 0 Tile_X0Y5_A_config_C_bit2
rlabel metal3 9476 523691 9476 523691 0 Tile_X0Y5_A_config_C_bit3
rlabel metal3 9476 519611 9476 519611 0 Tile_X0Y5_B_I_top
rlabel metal3 2775 518908 2775 518908 0 Tile_X0Y5_B_O_top
rlabel metal3 9476 520359 9476 520359 0 Tile_X0Y5_B_T_top
rlabel metal3 3787 524348 3787 524348 0 Tile_X0Y5_B_config_C_bit0
rlabel metal3 9476 525555 9476 525555 0 Tile_X0Y5_B_config_C_bit1
rlabel metal3 9476 526303 9476 526303 0 Tile_X0Y5_B_config_C_bit2
rlabel metal3 9476 527051 9476 527051 0 Tile_X0Y5_B_config_C_bit3
rlabel metal3 9476 472087 9476 472087 0 Tile_X0Y6_A_I_top
rlabel metal3 9476 471339 9476 471339 0 Tile_X0Y6_A_O_top
rlabel metal3 2407 473348 2407 473348 0 Tile_X0Y6_A_T_top
rlabel metal3 3787 476068 3787 476068 0 Tile_X0Y6_A_config_C_bit0
rlabel metal3 9476 477283 9476 477283 0 Tile_X0Y6_A_config_C_bit1
rlabel metal3 9476 478031 9476 478031 0 Tile_X0Y6_A_config_C_bit2
rlabel metal3 9476 478779 9476 478779 0 Tile_X0Y6_A_config_C_bit3
rlabel metal3 9476 474699 9476 474699 0 Tile_X0Y6_B_I_top
rlabel metal3 9476 473951 9476 473951 0 Tile_X0Y6_B_O_top
rlabel metal3 9476 475419 9476 475419 0 Tile_X0Y6_B_T_top
rlabel metal3 9476 479499 9476 479499 0 Tile_X0Y6_B_config_C_bit0
rlabel metal3 3143 480148 3143 480148 0 Tile_X0Y6_B_config_C_bit1
rlabel metal3 9476 481363 9476 481363 0 Tile_X0Y6_B_config_C_bit2
rlabel metal3 9476 482111 9476 482111 0 Tile_X0Y6_B_config_C_bit3
rlabel metal3 9476 427142 9476 427142 0 Tile_X0Y7_A_I_top
rlabel metal3 5338 426428 5338 426428 0 Tile_X0Y7_A_O_top
rlabel metal3 3787 427788 3787 427788 0 Tile_X0Y7_A_T_top
rlabel metal3 9476 431222 9476 431222 0 Tile_X0Y7_A_config_C_bit0
rlabel metal3 3143 431868 3143 431868 0 Tile_X0Y7_A_config_C_bit1
rlabel metal3 3787 433228 3787 433228 0 Tile_X0Y7_A_config_C_bit2
rlabel metal3 3787 433908 3787 433908 0 Tile_X0Y7_A_config_C_bit3
rlabel metal3 3787 429828 3787 429828 0 Tile_X0Y7_B_I_top
rlabel metal3 3787 429148 3787 429148 0 Tile_X0Y7_B_O_top
rlabel metal3 5338 430508 5338 430508 0 Tile_X0Y7_B_T_top
rlabel metal3 5338 434588 5338 434588 0 Tile_X0Y7_B_config_C_bit0
rlabel metal3 9476 435302 9476 435302 0 Tile_X0Y7_B_config_C_bit1
rlabel metal3 3787 435948 3787 435948 0 Tile_X0Y7_B_config_C_bit2
rlabel metal3 3787 437308 3787 437308 0 Tile_X0Y7_B_config_C_bit3
rlabel metal3 5338 382228 5338 382228 0 Tile_X0Y8_A_I_top
rlabel metal3 9476 381487 9476 381487 0 Tile_X0Y8_A_O_top
rlabel metal3 9476 382955 9476 382955 0 Tile_X0Y8_A_T_top
rlabel metal3 5338 386308 5338 386308 0 Tile_X0Y8_A_config_C_bit0
rlabel metal3 9476 387035 9476 387035 0 Tile_X0Y8_A_config_C_bit1
rlabel metal3 3787 387668 3787 387668 0 Tile_X0Y8_A_config_C_bit2
rlabel metal3 9476 388899 9476 388899 0 Tile_X0Y8_A_config_C_bit3
rlabel metal3 9476 384819 9476 384819 0 Tile_X0Y8_B_I_top
rlabel metal3 3143 383588 3143 383588 0 Tile_X0Y8_B_O_top
rlabel metal3 9476 385567 9476 385567 0 Tile_X0Y8_B_T_top
rlabel metal3 9476 389647 9476 389647 0 Tile_X0Y8_B_config_C_bit0
rlabel metal3 5338 390388 5338 390388 0 Tile_X0Y8_B_config_C_bit1
rlabel metal3 9476 391115 9476 391115 0 Tile_X0Y8_B_config_C_bit2
rlabel metal3 3787 391748 3787 391748 0 Tile_X0Y8_B_config_C_bit3
rlabel metal3 9476 337295 9476 337295 0 Tile_X0Y9_A_I_top
rlabel metal3 9476 336547 9476 336547 0 Tile_X0Y9_A_O_top
rlabel metal3 5338 338028 5338 338028 0 Tile_X0Y9_A_T_top
rlabel metal3 9476 341375 9476 341375 0 Tile_X0Y9_A_config_C_bit0
rlabel metal3 5338 342108 5338 342108 0 Tile_X0Y9_A_config_C_bit1
rlabel metal3 9476 342843 9476 342843 0 Tile_X0Y9_A_config_C_bit2
rlabel metal3 3787 343468 3787 343468 0 Tile_X0Y9_A_config_C_bit3
rlabel metal3 3787 339388 3787 339388 0 Tile_X0Y9_B_I_top
rlabel metal3 9476 338763 9476 338763 0 Tile_X0Y9_B_O_top
rlabel metal3 9476 340627 9476 340627 0 Tile_X0Y9_B_T_top
rlabel metal3 9476 344707 9476 344707 0 Tile_X0Y9_B_config_C_bit0
rlabel metal3 9476 345455 9476 345455 0 Tile_X0Y9_B_config_C_bit1
rlabel metal3 5338 346188 5338 346188 0 Tile_X0Y9_B_config_C_bit2
rlabel metal3 9476 346923 9476 346923 0 Tile_X0Y9_B_config_C_bit3
rlabel metal2 405069 755820 405069 755820 0 Tile_X10Y0_A_I_top
rlabel metal2 403933 755820 403933 755820 0 Tile_X10Y0_A_O_top
rlabel metal2 406311 755820 406311 755820 0 Tile_X10Y0_A_T_top
rlabel metal2 410465 755820 410465 755820 0 Tile_X10Y0_A_config_C_bit0
rlabel metal2 411661 755820 411661 755820 0 Tile_X10Y0_A_config_C_bit1
rlabel metal2 412797 755820 412797 755820 0 Tile_X10Y0_A_config_C_bit2
rlabel metal2 414039 755820 414039 755820 0 Tile_X10Y0_A_config_C_bit3
rlabel metal2 408395 755820 408395 755820 0 Tile_X10Y0_B_I_top
rlabel metal2 407001 755820 407001 755820 0 Tile_X10Y0_B_O_top
rlabel metal2 409577 755820 409577 755820 0 Tile_X10Y0_B_T_top
rlabel metal2 414927 755820 414927 755820 0 Tile_X10Y0_B_config_C_bit0
rlabel metal2 416123 755820 416123 755820 0 Tile_X10Y0_B_config_C_bit1
rlabel metal2 417305 755820 417305 755820 0 Tile_X10Y0_B_config_C_bit2
rlabel metal2 417949 755820 417949 755820 0 Tile_X10Y0_B_config_C_bit3
rlabel metal2 403400 5897 403400 5897 0 Tile_X10Y17_VALUE_top0
rlabel metal2 404780 5897 404780 5897 0 Tile_X10Y17_VALUE_top1
rlabel metal2 406160 5897 406160 5897 0 Tile_X10Y17_VALUE_top2
rlabel metal2 407540 5897 407540 5897 0 Tile_X10Y17_VALUE_top3
rlabel metal2 408920 5897 408920 5897 0 Tile_X10Y17_VALUE_top4
rlabel metal2 410300 5897 410300 5897 0 Tile_X10Y17_VALUE_top5
rlabel metal2 411680 5897 411680 5897 0 Tile_X10Y17_VALUE_top6
rlabel metal2 413060 5897 413060 5897 0 Tile_X10Y17_VALUE_top7
rlabel via3 481459 310420 481459 310420 0 Tile_X11Y10_AD_SRAM0
rlabel metal3 483276 317696 483276 317696 0 Tile_X11Y10_AD_SRAM1
rlabel metal3 483813 295188 483813 295188 0 Tile_X11Y10_AD_SRAM2
rlabel metal3 481686 318308 481686 318308 0 Tile_X11Y10_AD_SRAM3
rlabel metal3 484365 294508 484365 294508 0 Tile_X11Y10_AD_SRAM4
rlabel metal3 484273 293828 484273 293828 0 Tile_X11Y10_AD_SRAM5
rlabel metal3 477388 319051 477388 319051 0 Tile_X11Y10_AD_SRAM6
rlabel metal3 483721 293148 483721 293148 0 Tile_X11Y10_AD_SRAM7
rlabel metal3 481686 319668 481686 319668 0 Tile_X11Y10_AD_SRAM8
rlabel metal3 485193 292468 485193 292468 0 Tile_X11Y10_AD_SRAM9
rlabel metal3 485101 291788 485101 291788 0 Tile_X11Y10_BEN_SRAM0
rlabel metal3 477388 320411 477388 320411 0 Tile_X11Y10_BEN_SRAM1
rlabel metal3 484664 287708 484664 287708 0 Tile_X11Y10_BEN_SRAM10
rlabel metal3 477388 323131 477388 323131 0 Tile_X11Y10_BEN_SRAM11
rlabel metal3 483276 323612 483276 323612 0 Tile_X11Y10_BEN_SRAM12
rlabel metal3 481045 334084 481045 334084 0 Tile_X11Y10_BEN_SRAM13
rlabel metal3 483805 334084 483805 334084 0 Tile_X11Y10_BEN_SRAM14
rlabel metal3 483000 324360 483000 324360 0 Tile_X11Y10_BEN_SRAM15
rlabel metal3 482379 336668 482379 336668 0 Tile_X11Y10_BEN_SRAM16
rlabel metal3 483276 324972 483276 324972 0 Tile_X11Y10_BEN_SRAM17
rlabel metal3 480907 336668 480907 336668 0 Tile_X11Y10_BEN_SRAM18
rlabel metal3 483667 336668 483667 336668 0 Tile_X11Y10_BEN_SRAM19
rlabel metal3 485009 291108 485009 291108 0 Tile_X11Y10_BEN_SRAM2
rlabel metal3 484687 325788 484687 325788 0 Tile_X11Y10_BEN_SRAM20
rlabel metal3 484273 357068 484273 357068 0 Tile_X11Y10_BEN_SRAM21
rlabel metal3 483276 326332 483276 326332 0 Tile_X11Y10_BEN_SRAM22
rlabel metal3 485009 356388 485009 356388 0 Tile_X11Y10_BEN_SRAM23
rlabel metal3 483629 355708 483629 355708 0 Tile_X11Y10_BEN_SRAM24
rlabel metal3 484380 327080 484380 327080 0 Tile_X11Y10_BEN_SRAM25
rlabel metal3 478377 329596 478377 329596 0 Tile_X11Y10_BEN_SRAM26
rlabel metal3 477388 327726 477388 327726 0 Tile_X11Y10_BEN_SRAM27
rlabel metal3 477664 327964 477664 327964 0 Tile_X11Y10_BEN_SRAM28
rlabel via3 478699 334084 478699 334084 0 Tile_X11Y10_BEN_SRAM29
rlabel metal3 481686 321028 481686 321028 0 Tile_X11Y10_BEN_SRAM3
rlabel metal3 483000 328440 483000 328440 0 Tile_X11Y10_BEN_SRAM30
rlabel metal3 477653 328644 477653 328644 0 Tile_X11Y10_BEN_SRAM31
rlabel metal3 483629 290428 483629 290428 0 Tile_X11Y10_BEN_SRAM4
rlabel metal3 484618 289748 484618 289748 0 Tile_X11Y10_BEN_SRAM5
rlabel metal3 477388 321771 477388 321771 0 Tile_X11Y10_BEN_SRAM6
rlabel metal3 485354 289068 485354 289068 0 Tile_X11Y10_BEN_SRAM7
rlabel metal3 481686 322388 481686 322388 0 Tile_X11Y10_BEN_SRAM8
rlabel metal3 483974 288388 483974 288388 0 Tile_X11Y10_BEN_SRAM9
rlabel metal3 477388 329086 477388 329086 0 Tile_X11Y10_CLOCK_SRAM
rlabel metal3 477848 329324 477848 329324 0 Tile_X11Y10_DI_SRAM0
rlabel metal3 483721 351628 483721 351628 0 Tile_X11Y10_DI_SRAM1
rlabel metal3 484365 350948 484365 350948 0 Tile_X11Y10_DI_SRAM10
rlabel metal3 484457 347548 484457 347548 0 Tile_X11Y10_DI_SRAM11
rlabel metal4 479044 333540 479044 333540 0 Tile_X11Y10_DI_SRAM12
rlabel metal3 484342 346868 484342 346868 0 Tile_X11Y10_DI_SRAM13
rlabel metal4 484380 334152 484380 334152 0 Tile_X11Y10_DI_SRAM14
rlabel metal3 485101 346188 485101 346188 0 Tile_X11Y10_DI_SRAM15
rlabel metal3 478205 333540 478205 333540 0 Tile_X11Y10_DI_SRAM16
rlabel metal3 483276 335920 483276 335920 0 Tile_X11Y10_DI_SRAM17
rlabel metal3 486205 344828 486205 344828 0 Tile_X11Y10_DI_SRAM18
rlabel metal3 485561 336668 485561 336668 0 Tile_X11Y10_DI_SRAM19
rlabel metal3 484380 329800 484380 329800 0 Tile_X11Y10_DI_SRAM2
rlabel metal3 483905 344148 483905 344148 0 Tile_X11Y10_DI_SRAM20
rlabel metal3 478389 334900 478389 334900 0 Tile_X11Y10_DI_SRAM21
rlabel metal3 477469 335172 477469 335172 0 Tile_X11Y10_DI_SRAM22
rlabel metal4 484012 339116 484012 339116 0 Tile_X11Y10_DI_SRAM23
rlabel metal3 481766 349588 481766 349588 0 Tile_X11Y10_DI_SRAM24
rlabel metal3 483813 348908 483813 348908 0 Tile_X11Y10_DI_SRAM25
rlabel metal4 484380 338844 484380 338844 0 Tile_X11Y10_DI_SRAM26
rlabel metal3 484549 348228 484549 348228 0 Tile_X11Y10_DI_SRAM27
rlabel metal4 477388 338810 477388 338810 0 Tile_X11Y10_DI_SRAM28
rlabel metal3 477388 337246 477388 337246 0 Tile_X11Y10_DI_SRAM29
rlabel metal3 483276 330276 483276 330276 0 Tile_X11Y10_DI_SRAM3
rlabel metal4 478860 338776 478860 338776 0 Tile_X11Y10_DI_SRAM30
rlabel metal4 483276 338504 483276 338504 0 Tile_X11Y10_DI_SRAM31
rlabel metal3 483092 330752 483092 330752 0 Tile_X11Y10_DI_SRAM4
rlabel metal4 482908 331228 482908 331228 0 Tile_X11Y10_DI_SRAM5
rlabel metal3 478297 330820 478297 330820 0 Tile_X11Y10_DI_SRAM6
rlabel metal4 477388 331874 477388 331874 0 Tile_X11Y10_DI_SRAM7
rlabel metal4 483460 332316 483460 332316 0 Tile_X11Y10_DI_SRAM8
rlabel metal4 478860 332792 478860 332792 0 Tile_X11Y10_DI_SRAM9
rlabel metal4 486404 296284 486404 296284 0 Tile_X11Y10_DO_SRAM0
rlabel metal3 483276 308924 483276 308924 0 Tile_X11Y10_DO_SRAM1
rlabel metal3 481686 311508 481686 311508 0 Tile_X11Y10_DO_SRAM10
rlabel metal3 485653 304708 485653 304708 0 Tile_X11Y10_DO_SRAM11
rlabel metal3 486021 304028 486021 304028 0 Tile_X11Y10_DO_SRAM12
rlabel metal3 477388 312251 477388 312251 0 Tile_X11Y10_DO_SRAM13
rlabel metal3 486113 303348 486113 303348 0 Tile_X11Y10_DO_SRAM14
rlabel metal3 481686 312868 481686 312868 0 Tile_X11Y10_DO_SRAM15
rlabel metal3 486205 302668 486205 302668 0 Tile_X11Y10_DO_SRAM16
rlabel metal3 485745 301988 485745 301988 0 Tile_X11Y10_DO_SRAM17
rlabel metal3 477388 313611 477388 313611 0 Tile_X11Y10_DO_SRAM18
rlabel metal4 486220 313888 486220 313888 0 Tile_X11Y10_DO_SRAM19
rlabel metal4 484380 308720 484380 308720 0 Tile_X11Y10_DO_SRAM2
rlabel metal3 481686 314228 481686 314228 0 Tile_X11Y10_DO_SRAM20
rlabel metal3 484342 300628 484342 300628 0 Tile_X11Y10_DO_SRAM21
rlabel metal3 486228 299948 486228 299948 0 Tile_X11Y10_DO_SRAM22
rlabel metal3 483276 314976 483276 314976 0 Tile_X11Y10_DO_SRAM23
rlabel metal3 477653 315316 477653 315316 0 Tile_X11Y10_DO_SRAM24
rlabel metal3 481686 315588 481686 315588 0 Tile_X11Y10_DO_SRAM25
rlabel metal3 477561 315860 477561 315860 0 Tile_X11Y10_DO_SRAM26
rlabel via3 479987 310420 479987 310420 0 Tile_X11Y10_DO_SRAM27
rlabel metal3 477388 316331 477388 316331 0 Tile_X11Y10_DO_SRAM28
rlabel metal3 479941 311236 479941 311236 0 Tile_X11Y10_DO_SRAM29
rlabel metal3 477388 309531 477388 309531 0 Tile_X11Y10_DO_SRAM3
rlabel metal3 481686 316948 481686 316948 0 Tile_X11Y10_DO_SRAM30
rlabel metal3 483284 296548 483284 296548 0 Tile_X11Y10_DO_SRAM31
rlabel metal4 482908 308652 482908 308652 0 Tile_X11Y10_DO_SRAM4
rlabel metal3 481686 310148 481686 310148 0 Tile_X11Y10_DO_SRAM5
rlabel metal4 478676 308584 478676 308584 0 Tile_X11Y10_DO_SRAM6
rlabel metal3 485929 306068 485929 306068 0 Tile_X11Y10_DO_SRAM7
rlabel metal3 477388 310891 477388 310891 0 Tile_X11Y10_DO_SRAM8
rlabel metal3 485837 305388 485837 305388 0 Tile_X11Y10_DO_SRAM9
rlabel metal3 477388 337994 477388 337994 0 Tile_X11Y10_EN_SRAM
rlabel metal4 483460 340136 483460 340136 0 Tile_X11Y10_R_WB_SRAM
rlabel metal3 483928 196588 483928 196588 0 Tile_X11Y12_AD_SRAM0
rlabel metal3 484365 205428 484365 205428 0 Tile_X11Y12_AD_SRAM1
rlabel metal3 483307 227868 483307 227868 0 Tile_X11Y12_AD_SRAM2
rlabel metal3 483721 204748 483721 204748 0 Tile_X11Y12_AD_SRAM3
rlabel metal3 477388 228559 477388 228559 0 Tile_X11Y12_AD_SRAM4
rlabel metal3 484273 204068 484273 204068 0 Tile_X11Y12_AD_SRAM5
rlabel metal3 485101 203388 485101 203388 0 Tile_X11Y12_AD_SRAM6
rlabel metal3 483276 229364 483276 229364 0 Tile_X11Y12_AD_SRAM7
rlabel metal3 485009 202708 485009 202708 0 Tile_X11Y12_AD_SRAM8
rlabel metal3 477388 229919 477388 229919 0 Tile_X11Y12_AD_SRAM9
rlabel metal3 484618 202028 484618 202028 0 Tile_X11Y12_BEN_SRAM0
rlabel metal3 483629 201348 483629 201348 0 Tile_X11Y12_BEN_SRAM1
rlabel metal3 483307 232628 483307 232628 0 Tile_X11Y12_BEN_SRAM10
rlabel metal3 485354 197268 485354 197268 0 Tile_X11Y12_BEN_SRAM11
rlabel metal3 483307 233308 483307 233308 0 Tile_X11Y12_BEN_SRAM12
rlabel metal3 483307 233988 483307 233988 0 Tile_X11Y12_BEN_SRAM13
rlabel metal3 483974 270028 483974 270028 0 Tile_X11Y12_BEN_SRAM14
rlabel metal3 484664 269348 484664 269348 0 Tile_X11Y12_BEN_SRAM15
rlabel metal3 483000 234600 483000 234600 0 Tile_X11Y12_BEN_SRAM16
rlabel metal3 485354 268668 485354 268668 0 Tile_X11Y12_BEN_SRAM17
rlabel metal3 483307 235348 483307 235348 0 Tile_X11Y12_BEN_SRAM18
rlabel metal3 483928 267988 483928 267988 0 Tile_X11Y12_BEN_SRAM19
rlabel metal3 477388 230667 477388 230667 0 Tile_X11Y12_BEN_SRAM2
rlabel metal3 485009 267308 485009 267308 0 Tile_X11Y12_BEN_SRAM20
rlabel metal3 483000 235960 483000 235960 0 Tile_X11Y12_BEN_SRAM21
rlabel metal3 482333 247044 482333 247044 0 Tile_X11Y12_BEN_SRAM22
rlabel metal3 483307 236708 483307 236708 0 Tile_X11Y12_BEN_SRAM23
rlabel metal3 485101 265948 485101 265948 0 Tile_X11Y12_BEN_SRAM24
rlabel metal3 483629 265268 483629 265268 0 Tile_X11Y12_BEN_SRAM25
rlabel metal3 484380 237320 484380 237320 0 Tile_X11Y12_BEN_SRAM26
rlabel metal3 477572 237660 477572 237660 0 Tile_X11Y12_BEN_SRAM27
rlabel metal3 477388 237971 477388 237971 0 Tile_X11Y12_BEN_SRAM28
rlabel metal3 477572 238204 477572 238204 0 Tile_X11Y12_BEN_SRAM29
rlabel metal3 484664 200668 484664 200668 0 Tile_X11Y12_BEN_SRAM3
rlabel metal3 477480 238476 477480 238476 0 Tile_X11Y12_BEN_SRAM30
rlabel metal3 485561 238748 485561 238748 0 Tile_X11Y12_BEN_SRAM31
rlabel metal3 477388 231279 477388 231279 0 Tile_X11Y12_BEN_SRAM4
rlabel metal3 485308 199988 485308 199988 0 Tile_X11Y12_BEN_SRAM5
rlabel metal3 483974 199308 483974 199308 0 Tile_X11Y12_BEN_SRAM6
rlabel metal3 483307 231948 483307 231948 0 Tile_X11Y12_BEN_SRAM7
rlabel metal3 482548 198628 482548 198628 0 Tile_X11Y12_BEN_SRAM8
rlabel metal3 482594 197948 482594 197948 0 Tile_X11Y12_BEN_SRAM9
rlabel metal3 477756 239020 477756 239020 0 Tile_X11Y12_CLOCK_SRAM
rlabel metal3 483307 239428 483307 239428 0 Tile_X11Y12_DI_SRAM0
rlabel metal3 484273 261868 484273 261868 0 Tile_X11Y12_DI_SRAM1
rlabel metal3 477848 242012 477848 242012 0 Tile_X11Y12_DI_SRAM10
rlabel metal3 485193 257788 485193 257788 0 Tile_X11Y12_DI_SRAM11
rlabel metal3 485929 257108 485929 257108 0 Tile_X11Y12_DI_SRAM12
rlabel metal4 484380 243780 484380 243780 0 Tile_X11Y12_DI_SRAM13
rlabel metal3 482893 256428 482893 256428 0 Tile_X11Y12_DI_SRAM14
rlabel metal4 484564 244392 484564 244392 0 Tile_X11Y12_DI_SRAM15
rlabel metal3 484365 260508 484365 260508 0 Tile_X11Y12_DI_SRAM16
rlabel metal3 483077 255068 483077 255068 0 Tile_X11Y12_DI_SRAM17
rlabel metal3 486021 259828 486021 259828 0 Tile_X11Y12_DI_SRAM18
rlabel metal4 486312 244460 486312 244460 0 Tile_X11Y12_DI_SRAM19
rlabel metal3 483276 239972 483276 239972 0 Tile_X11Y12_DI_SRAM2
rlabel metal4 483276 245480 483276 245480 0 Tile_X11Y12_DI_SRAM20
rlabel metal3 486113 253708 486113 253708 0 Tile_X11Y12_DI_SRAM21
rlabel metal3 483169 253028 483169 253028 0 Tile_X11Y12_DI_SRAM22
rlabel metal4 477388 246199 477388 246199 0 Tile_X11Y12_DI_SRAM23
rlabel metal3 483721 259148 483721 259148 0 Tile_X11Y12_DI_SRAM24
rlabel metal4 482908 246840 482908 246840 0 Tile_X11Y12_DI_SRAM25
rlabel metal3 478492 246364 478492 246364 0 Tile_X11Y12_DI_SRAM26
rlabel metal3 485469 250988 485469 250988 0 Tile_X11Y12_DI_SRAM27
rlabel metal2 483230 248132 483230 248132 0 Tile_X11Y12_DI_SRAM28
rlabel metal3 485561 250308 485561 250308 0 Tile_X11Y12_DI_SRAM29
rlabel metal3 483092 240448 483092 240448 0 Tile_X11Y12_DI_SRAM3
rlabel metal3 485377 248948 485377 248948 0 Tile_X11Y12_DI_SRAM30
rlabel metal3 483997 249628 483997 249628 0 Tile_X11Y12_DI_SRAM31
rlabel metal2 482954 240924 482954 240924 0 Tile_X11Y12_DI_SRAM4
rlabel metal3 482724 240720 482724 240720 0 Tile_X11Y12_DI_SRAM5
rlabel metal4 483276 241944 483276 241944 0 Tile_X11Y12_DI_SRAM6
rlabel metal4 484748 242352 484748 242352 0 Tile_X11Y12_DI_SRAM7
rlabel metal4 484932 242760 484932 242760 0 Tile_X11Y12_DI_SRAM8
rlabel metal3 485032 255748 485032 255748 0 Tile_X11Y12_DI_SRAM9
rlabel metal3 483905 206108 483905 206108 0 Tile_X11Y12_DO_SRAM0
rlabel metal3 477179 219050 477179 219050 0 Tile_X11Y12_DO_SRAM1
rlabel metal3 485745 214948 485745 214948 0 Tile_X11Y12_DO_SRAM10
rlabel metal3 477179 221770 477179 221770 0 Tile_X11Y12_DO_SRAM11
rlabel metal3 485837 214268 485837 214268 0 Tile_X11Y12_DO_SRAM12
rlabel metal3 486205 213588 486205 213588 0 Tile_X11Y12_DO_SRAM13
rlabel metal3 477179 222586 477179 222586 0 Tile_X11Y12_DO_SRAM14
rlabel metal3 485193 212908 485193 212908 0 Tile_X11Y12_DO_SRAM15
rlabel metal3 477179 223130 477179 223130 0 Tile_X11Y12_DO_SRAM16
rlabel metal4 486404 213754 486404 213754 0 Tile_X11Y12_DO_SRAM17
rlabel metal3 485929 211548 485929 211548 0 Tile_X11Y12_DO_SRAM18
rlabel metal3 477179 223946 477179 223946 0 Tile_X11Y12_DO_SRAM19
rlabel metal3 477202 219322 477202 219322 0 Tile_X11Y12_DO_SRAM2
rlabel metal3 484457 210868 484457 210868 0 Tile_X11Y12_DO_SRAM20
rlabel metal3 477179 224490 477179 224490 0 Tile_X11Y12_DO_SRAM21
rlabel metal4 486404 224740 486404 224740 0 Tile_X11Y12_DO_SRAM22
rlabel metal3 482893 209508 482893 209508 0 Tile_X11Y12_DO_SRAM23
rlabel metal3 477388 225227 477388 225227 0 Tile_X11Y12_DO_SRAM24
rlabel metal3 482985 208828 482985 208828 0 Tile_X11Y12_DO_SRAM25
rlabel metal3 477388 225839 477388 225839 0 Tile_X11Y12_DO_SRAM26
rlabel metal2 486312 209760 486312 209760 0 Tile_X11Y12_DO_SRAM27
rlabel metal3 483813 207468 483813 207468 0 Tile_X11Y12_DO_SRAM28
rlabel metal3 483307 226508 483307 226508 0 Tile_X11Y12_DO_SRAM29
rlabel metal3 477179 219594 477179 219594 0 Tile_X11Y12_DO_SRAM3
rlabel metal3 483284 206788 483284 206788 0 Tile_X11Y12_DO_SRAM30
rlabel metal3 477388 227199 477388 227199 0 Tile_X11Y12_DO_SRAM31
rlabel metal3 477179 219866 477179 219866 0 Tile_X11Y12_DO_SRAM4
rlabel metal3 477179 220138 477179 220138 0 Tile_X11Y12_DO_SRAM5
rlabel metal3 477179 220410 477179 220410 0 Tile_X11Y12_DO_SRAM6
rlabel metal3 477179 220682 477179 220682 0 Tile_X11Y12_DO_SRAM7
rlabel metal3 477179 221010 477179 221010 0 Tile_X11Y12_DO_SRAM8
rlabel metal3 477179 221226 477179 221226 0 Tile_X11Y12_DO_SRAM9
rlabel metal3 483813 252348 483813 252348 0 Tile_X11Y12_EN_SRAM
rlabel metal3 486205 251668 486205 251668 0 Tile_X11Y12_R_WB_SRAM
rlabel metal3 484664 192508 484664 192508 0 Tile_X11Y14_AD_SRAM0
rlabel metal3 483989 146268 483989 146268 0 Tile_X11Y14_AD_SRAM1
rlabel metal3 477388 138095 477388 138095 0 Tile_X11Y14_AD_SRAM2
rlabel metal3 482333 149260 482333 149260 0 Tile_X11Y14_AD_SRAM3
rlabel metal3 486021 148988 486021 148988 0 Tile_X11Y14_AD_SRAM4
rlabel metal3 483851 147764 483851 147764 0 Tile_X11Y14_AD_SRAM5
rlabel metal3 482471 149124 482471 149124 0 Tile_X11Y14_AD_SRAM6
rlabel metal3 477388 139455 477388 139455 0 Tile_X11Y14_AD_SRAM7
rlabel metal3 483989 150484 483989 150484 0 Tile_X11Y14_AD_SRAM8
rlabel metal3 477388 140067 477388 140067 0 Tile_X11Y14_AD_SRAM9
rlabel metal3 477572 140284 477572 140284 0 Tile_X11Y14_BEN_SRAM0
rlabel metal3 478032 140556 478032 140556 0 Tile_X11Y14_BEN_SRAM1
rlabel metal3 478101 152660 478101 152660 0 Tile_X11Y14_BEN_SRAM10
rlabel metal3 478147 152932 478147 152932 0 Tile_X11Y14_BEN_SRAM11
rlabel metal4 484380 144636 484380 144636 0 Tile_X11Y14_BEN_SRAM12
rlabel metal3 482341 180268 482341 180268 0 Tile_X11Y14_BEN_SRAM13
rlabel metal4 484564 145180 484564 145180 0 Tile_X11Y14_BEN_SRAM14
rlabel metal3 484526 179588 484526 179588 0 Tile_X11Y14_BEN_SRAM15
rlabel metal3 482272 191828 482272 191828 0 Tile_X11Y14_BEN_SRAM16
rlabel metal3 477204 144895 477204 144895 0 Tile_X11Y14_BEN_SRAM17
rlabel via3 481643 155924 481643 155924 0 Tile_X11Y14_BEN_SRAM18
rlabel metal3 483667 155924 483667 155924 0 Tile_X11Y14_BEN_SRAM19
rlabel metal3 477388 140815 477388 140815 0 Tile_X11Y14_BEN_SRAM2
rlabel metal3 483192 177548 483192 177548 0 Tile_X11Y14_BEN_SRAM20
rlabel metal3 483238 176868 483238 176868 0 Tile_X11Y14_BEN_SRAM21
rlabel metal3 483284 190468 483284 190468 0 Tile_X11Y14_BEN_SRAM22
rlabel metal3 480033 156740 480033 156740 0 Tile_X11Y14_BEN_SRAM23
rlabel metal4 484564 147492 484564 147492 0 Tile_X11Y14_BEN_SRAM24
rlabel metal3 478469 147084 478469 147084 0 Tile_X11Y14_BEN_SRAM25
rlabel metal3 482893 174828 482893 174828 0 Tile_X11Y14_BEN_SRAM26
rlabel metal3 477388 147615 477388 147615 0 Tile_X11Y14_BEN_SRAM27
rlabel metal3 482249 174148 482249 174148 0 Tile_X11Y14_BEN_SRAM28
rlabel metal4 484380 148920 484380 148920 0 Tile_X11Y14_BEN_SRAM29
rlabel metal3 483353 142188 483353 142188 0 Tile_X11Y14_BEN_SRAM3
rlabel metal3 485009 173468 485009 173468 0 Tile_X11Y14_BEN_SRAM30
rlabel metal3 482985 172788 482985 172788 0 Tile_X11Y14_BEN_SRAM31
rlabel metal3 477388 141427 477388 141427 0 Tile_X11Y14_BEN_SRAM4
rlabel metal3 478676 141644 478676 141644 0 Tile_X11Y14_BEN_SRAM5
rlabel metal3 483445 142868 483445 142868 0 Tile_X11Y14_BEN_SRAM6
rlabel metal3 486205 153068 486205 153068 0 Tile_X11Y14_BEN_SRAM7
rlabel metal4 484748 146404 484748 146404 0 Tile_X11Y14_BEN_SRAM8
rlabel metal4 478860 143480 478860 143480 0 Tile_X11Y14_BEN_SRAM9
rlabel metal3 486021 161228 486021 161228 0 Tile_X11Y14_CLOCK_SRAM
rlabel metal3 484365 172108 484365 172108 0 Tile_X11Y14_DI_SRAM0
rlabel metal3 483169 153748 483169 153748 0 Tile_X11Y14_DI_SRAM1
rlabel metal3 477664 151980 477664 151980 0 Tile_X11Y14_DI_SRAM10
rlabel metal4 478676 153340 478676 153340 0 Tile_X11Y14_DI_SRAM11
rlabel metal3 485929 167348 485929 167348 0 Tile_X11Y14_DI_SRAM12
rlabel metal3 485032 166668 485032 166668 0 Tile_X11Y14_DI_SRAM13
rlabel metal4 480516 156128 480516 156128 0 Tile_X11Y14_DI_SRAM14
rlabel metal3 478584 153340 478584 153340 0 Tile_X11Y14_DI_SRAM15
rlabel metal4 484564 154292 484564 154292 0 Tile_X11Y14_DI_SRAM16
rlabel metal3 486113 165308 486113 165308 0 Tile_X11Y14_DI_SRAM17
rlabel metal3 483652 183668 483652 183668 0 Tile_X11Y14_DI_SRAM18
rlabel metal4 484380 155040 484380 155040 0 Tile_X11Y14_DI_SRAM19
rlabel metal3 481789 158508 481789 158508 0 Tile_X11Y14_DI_SRAM2
rlabel metal3 483698 182988 483698 182988 0 Tile_X11Y14_DI_SRAM20
rlabel metal2 486266 158148 486266 158148 0 Tile_X11Y14_DI_SRAM21
rlabel metal3 483353 163268 483353 163268 0 Tile_X11Y14_DI_SRAM22
rlabel metal3 485285 162588 485285 162588 0 Tile_X11Y14_DI_SRAM23
rlabel metal3 484196 155856 484196 155856 0 Tile_X11Y14_DI_SRAM24
rlabel metal3 485561 161908 485561 161908 0 Tile_X11Y14_DI_SRAM25
rlabel metal3 483307 156468 483307 156468 0 Tile_X11Y14_DI_SRAM26
rlabel metal3 486205 168708 486205 168708 0 Tile_X11Y14_DI_SRAM27
rlabel metal4 482908 158712 482908 158712 0 Tile_X11Y14_DI_SRAM28
rlabel metal3 477388 157135 477388 157135 0 Tile_X11Y14_DI_SRAM29
rlabel metal3 481137 153068 481137 153068 0 Tile_X11Y14_DI_SRAM3
rlabel metal4 483276 158712 483276 158712 0 Tile_X11Y14_DI_SRAM30
rlabel metal3 483307 157828 483307 157828 0 Tile_X11Y14_DI_SRAM31
rlabel metal3 484457 170748 484457 170748 0 Tile_X11Y14_DI_SRAM4
rlabel metal3 483276 150824 483276 150824 0 Tile_X11Y14_DI_SRAM5
rlabel metal2 483138 151300 483138 151300 0 Tile_X11Y14_DI_SRAM6
rlabel metal3 485561 152388 485561 152388 0 Tile_X11Y14_DI_SRAM7
rlabel metal3 484273 181628 484273 181628 0 Tile_X11Y14_DI_SRAM8
rlabel metal3 483629 163948 483629 163948 0 Tile_X11Y14_DI_SRAM9
rlabel metal3 485101 119068 485101 119068 0 Tile_X11Y14_DO_SRAM0
rlabel metal3 483276 128860 483276 128860 0 Tile_X11Y14_DO_SRAM1
rlabel metal3 483307 131308 483307 131308 0 Tile_X11Y14_DO_SRAM10
rlabel metal4 481436 128112 481436 128112 0 Tile_X11Y14_DO_SRAM11
rlabel metal3 477388 132015 477388 132015 0 Tile_X11Y14_DO_SRAM12
rlabel metal4 477388 128071 477388 128071 0 Tile_X11Y14_DO_SRAM13
rlabel metal3 486205 123148 486205 123148 0 Tile_X11Y14_DO_SRAM14
rlabel metal3 483307 132668 483307 132668 0 Tile_X11Y14_DO_SRAM15
rlabel metal3 482249 122468 482249 122468 0 Tile_X11Y14_DO_SRAM16
rlabel metal3 477388 133375 477388 133375 0 Tile_X11Y14_DO_SRAM17
rlabel metal3 482341 121788 482341 121788 0 Tile_X11Y14_DO_SRAM18
rlabel metal4 486036 133756 486036 133756 0 Tile_X11Y14_DO_SRAM19
rlabel metal3 477388 129295 477388 129295 0 Tile_X11Y14_DO_SRAM2
rlabel metal3 483276 134164 483276 134164 0 Tile_X11Y14_DO_SRAM20
rlabel metal4 486312 120700 486312 120700 0 Tile_X11Y14_DO_SRAM21
rlabel metal3 477388 134735 477388 134735 0 Tile_X11Y14_DO_SRAM22
rlabel metal3 485032 119748 485032 119748 0 Tile_X11Y14_DO_SRAM23
rlabel metal3 477388 135375 477388 135375 0 Tile_X11Y14_DO_SRAM24
rlabel metal3 483307 136068 483307 136068 0 Tile_X11Y14_DO_SRAM25
rlabel metal3 478492 135932 478492 135932 0 Tile_X11Y14_DO_SRAM26
rlabel metal3 483529 157420 483529 157420 0 Tile_X11Y14_DO_SRAM27
rlabel metal4 484380 136952 484380 136952 0 Tile_X11Y14_DO_SRAM28
rlabel metal3 477388 136735 477388 136735 0 Tile_X11Y14_DO_SRAM29
rlabel metal4 478860 128724 478860 128724 0 Tile_X11Y14_DO_SRAM3
rlabel metal4 484564 137904 484564 137904 0 Tile_X11Y14_DO_SRAM30
rlabel metal3 483928 175508 483928 175508 0 Tile_X11Y14_DO_SRAM31
rlabel metal4 483092 128588 483092 128588 0 Tile_X11Y14_DO_SRAM4
rlabel metal3 483276 130084 483276 130084 0 Tile_X11Y14_DO_SRAM5
rlabel metal4 484380 128452 484380 128452 0 Tile_X11Y14_DO_SRAM6
rlabel metal3 477388 130655 477388 130655 0 Tile_X11Y14_DO_SRAM7
rlabel metal4 484564 128452 484564 128452 0 Tile_X11Y14_DO_SRAM8
rlabel metal4 481620 128180 481620 128180 0 Tile_X11Y14_DO_SRAM9
rlabel metal3 485101 169388 485101 169388 0 Tile_X11Y14_EN_SRAM
rlabel metal4 486220 159848 486220 159848 0 Tile_X11Y14_R_WB_SRAM
rlabel metal3 483629 17068 483629 17068 0 Tile_X11Y16_AD_SRAM0
rlabel metal3 477388 47702 477388 47702 0 Tile_X11Y16_AD_SRAM1
rlabel metal3 483905 25228 483905 25228 0 Tile_X11Y16_AD_SRAM2
rlabel metal3 484365 24548 484365 24548 0 Tile_X11Y16_AD_SRAM3
rlabel metal3 483276 48484 483276 48484 0 Tile_X11Y16_AD_SRAM4
rlabel metal3 483813 23868 483813 23868 0 Tile_X11Y16_AD_SRAM5
rlabel metal3 477388 49062 477388 49062 0 Tile_X11Y16_AD_SRAM6
rlabel metal3 485101 23188 485101 23188 0 Tile_X11Y16_AD_SRAM7
rlabel metal3 484273 22508 484273 22508 0 Tile_X11Y16_AD_SRAM8
rlabel metal3 483276 49844 483276 49844 0 Tile_X11Y16_AD_SRAM9
rlabel metal3 483721 21828 483721 21828 0 Tile_X11Y16_BEN_SRAM0
rlabel metal3 477388 50422 477388 50422 0 Tile_X11Y16_BEN_SRAM1
rlabel metal3 485354 17748 485354 17748 0 Tile_X11Y16_BEN_SRAM10
rlabel metal3 477388 53142 477388 53142 0 Tile_X11Y16_BEN_SRAM11
rlabel metal3 481045 62220 481045 62220 0 Tile_X11Y16_BEN_SRAM12
rlabel metal3 481686 53788 481686 53788 0 Tile_X11Y16_BEN_SRAM13
rlabel metal3 483805 65892 483805 65892 0 Tile_X11Y16_BEN_SRAM14
rlabel metal3 483307 54468 483307 54468 0 Tile_X11Y16_BEN_SRAM15
rlabel metal3 482379 62220 482379 62220 0 Tile_X11Y16_BEN_SRAM16
rlabel metal3 480907 67524 480907 67524 0 Tile_X11Y16_BEN_SRAM17
rlabel metal3 481686 55148 481686 55148 0 Tile_X11Y16_BEN_SRAM18
rlabel metal3 483667 67524 483667 67524 0 Tile_X11Y16_BEN_SRAM19
rlabel metal3 484618 21148 484618 21148 0 Tile_X11Y16_BEN_SRAM2
rlabel metal3 483307 55828 483307 55828 0 Tile_X11Y16_BEN_SRAM20
rlabel metal4 481988 59432 481988 59432 0 Tile_X11Y16_BEN_SRAM21
rlabel metal3 483629 86428 483629 86428 0 Tile_X11Y16_BEN_SRAM22
rlabel metal3 481686 56508 481686 56508 0 Tile_X11Y16_BEN_SRAM23
rlabel metal3 485009 85748 485009 85748 0 Tile_X11Y16_BEN_SRAM24
rlabel metal3 483307 57188 483307 57188 0 Tile_X11Y16_BEN_SRAM25
rlabel via3 478699 63716 478699 63716 0 Tile_X11Y16_BEN_SRAM26
rlabel metal3 478377 60588 478377 60588 0 Tile_X11Y16_BEN_SRAM27
rlabel metal3 481686 57868 481686 57868 0 Tile_X11Y16_BEN_SRAM28
rlabel metal3 477561 58140 477561 58140 0 Tile_X11Y16_BEN_SRAM29
rlabel metal3 485009 20468 485009 20468 0 Tile_X11Y16_BEN_SRAM3
rlabel metal3 483307 58548 483307 58548 0 Tile_X11Y16_BEN_SRAM30
rlabel metal3 477653 58684 477653 58684 0 Tile_X11Y16_BEN_SRAM31
rlabel metal3 483276 51204 483276 51204 0 Tile_X11Y16_BEN_SRAM4
rlabel metal3 484664 19788 484664 19788 0 Tile_X11Y16_BEN_SRAM5
rlabel metal3 477388 51782 477388 51782 0 Tile_X11Y16_BEN_SRAM6
rlabel metal3 485308 19108 485308 19108 0 Tile_X11Y16_BEN_SRAM7
rlabel metal3 483974 18428 483974 18428 0 Tile_X11Y16_BEN_SRAM8
rlabel metal3 483276 52564 483276 52564 0 Tile_X11Y16_BEN_SRAM9
rlabel metal3 484273 82348 484273 82348 0 Tile_X11Y16_CLOCK_SRAM
rlabel metal3 481686 59228 481686 59228 0 Tile_X11Y16_DI_SRAM0
rlabel metal3 477745 59500 477745 59500 0 Tile_X11Y16_DI_SRAM1
rlabel metal3 478573 61948 478573 61948 0 Tile_X11Y16_DI_SRAM10
rlabel metal3 486113 80308 486113 80308 0 Tile_X11Y16_DI_SRAM11
rlabel metal3 477193 62492 477193 62492 0 Tile_X11Y16_DI_SRAM12
rlabel metal3 483721 76908 483721 76908 0 Tile_X11Y16_DI_SRAM13
rlabel metal3 484365 76228 484365 76228 0 Tile_X11Y16_DI_SRAM14
rlabel metal3 483092 63648 483092 63648 0 Tile_X11Y16_DI_SRAM15
rlabel metal3 478389 63580 478389 63580 0 Tile_X11Y16_DI_SRAM16
rlabel metal3 482540 63988 482540 63988 0 Tile_X11Y16_DI_SRAM17
rlabel metal3 484342 79628 484342 79628 0 Tile_X11Y16_DI_SRAM18
rlabel metal3 478481 64396 478481 64396 0 Tile_X11Y16_DI_SRAM19
rlabel metal3 483307 59908 483307 59908 0 Tile_X11Y16_DI_SRAM2
rlabel metal3 484089 67388 484089 67388 0 Tile_X11Y16_DI_SRAM20
rlabel metal4 484932 69224 484932 69224 0 Tile_X11Y16_DI_SRAM21
rlabel metal4 478676 66640 478676 66640 0 Tile_X11Y16_DI_SRAM22
rlabel metal3 482985 78948 482985 78948 0 Tile_X11Y16_DI_SRAM23
rlabel metal4 484748 68952 484748 68952 0 Tile_X11Y16_DI_SRAM24
rlabel metal4 483276 66368 483276 66368 0 Tile_X11Y16_DI_SRAM25
rlabel metal4 484564 68884 484564 68884 0 Tile_X11Y16_DI_SRAM26
rlabel metal4 486588 76394 486588 76394 0 Tile_X11Y16_DI_SRAM27
rlabel metal4 484380 68816 484380 68816 0 Tile_X11Y16_DI_SRAM28
rlabel metal4 483460 68612 483460 68612 0 Tile_X11Y16_DI_SRAM29
rlabel metal3 483276 60316 483276 60316 0 Tile_X11Y16_DI_SRAM3
rlabel metal4 483276 68000 483276 68000 0 Tile_X11Y16_DI_SRAM30
rlabel metal4 481620 68544 481620 68544 0 Tile_X11Y16_DI_SRAM31
rlabel metal3 483276 63240 483276 63240 0 Tile_X11Y16_DI_SRAM4
rlabel metal4 481620 61200 481620 61200 0 Tile_X11Y16_DI_SRAM5
rlabel metal4 483460 61744 483460 61744 0 Tile_X11Y16_DI_SRAM6
rlabel metal3 483307 61268 483307 61268 0 Tile_X11Y16_DI_SRAM7
rlabel metal3 478205 61404 478205 61404 0 Tile_X11Y16_DI_SRAM8
rlabel metal4 484380 63172 484380 63172 0 Tile_X11Y16_DI_SRAM9
rlabel metal3 485653 25908 485653 25908 0 Tile_X11Y16_DO_SRAM0
rlabel metal3 483307 38828 483307 38828 0 Tile_X11Y16_DO_SRAM1
rlabel metal4 476980 41140 476980 41140 0 Tile_X11Y16_DO_SRAM10
rlabel metal3 477388 41650 477388 41650 0 Tile_X11Y16_DO_SRAM11
rlabel metal3 486205 34068 486205 34068 0 Tile_X11Y16_DO_SRAM12
rlabel metal3 477388 42262 477388 42262 0 Tile_X11Y16_DO_SRAM13
rlabel metal3 477653 42636 477653 42636 0 Tile_X11Y16_DO_SRAM14
rlabel metal4 486036 42772 486036 42772 0 Tile_X11Y16_DO_SRAM15
rlabel metal2 483322 43044 483322 43044 0 Tile_X11Y16_DO_SRAM16
rlabel metal3 477561 43452 477561 43452 0 Tile_X11Y16_DO_SRAM17
rlabel metal3 477388 43622 477388 43622 0 Tile_X11Y16_DO_SRAM18
rlabel metal3 486021 31348 486021 31348 0 Tile_X11Y16_DO_SRAM19
rlabel metal4 484380 38692 484380 38692 0 Tile_X11Y16_DO_SRAM2
rlabel metal3 484756 30668 484756 30668 0 Tile_X11Y16_DO_SRAM20
rlabel metal3 483276 44404 483276 44404 0 Tile_X11Y16_DO_SRAM21
rlabel metal2 486450 40278 486450 40278 0 Tile_X11Y16_DO_SRAM22
rlabel metal3 477388 44982 477388 44982 0 Tile_X11Y16_DO_SRAM23
rlabel metal3 478389 45356 478389 45356 0 Tile_X11Y16_DO_SRAM24
rlabel metal3 482893 28628 482893 28628 0 Tile_X11Y16_DO_SRAM25
rlabel metal3 483307 45628 483307 45628 0 Tile_X11Y16_DO_SRAM26
rlabel metal3 482985 27948 482985 27948 0 Tile_X11Y16_DO_SRAM27
rlabel metal3 477388 46342 477388 46342 0 Tile_X11Y16_DO_SRAM28
rlabel metal3 479665 39916 479665 39916 0 Tile_X11Y16_DO_SRAM29
rlabel metal3 477388 39542 477388 39542 0 Tile_X11Y16_DO_SRAM3
rlabel metal3 480079 44404 480079 44404 0 Tile_X11Y16_DO_SRAM30
rlabel metal3 477388 47090 477388 47090 0 Tile_X11Y16_DO_SRAM31
rlabel metal4 484564 38624 484564 38624 0 Tile_X11Y16_DO_SRAM4
rlabel metal4 484748 38420 484748 38420 0 Tile_X11Y16_DO_SRAM5
rlabel metal3 483307 40188 483307 40188 0 Tile_X11Y16_DO_SRAM6
rlabel metal4 484932 38420 484932 38420 0 Tile_X11Y16_DO_SRAM7
rlabel metal3 477388 40902 477388 40902 0 Tile_X11Y16_DO_SRAM8
rlabel metal3 485929 35428 485929 35428 0 Tile_X11Y16_DO_SRAM9
rlabel metal3 485377 74868 485377 74868 0 Tile_X11Y16_EN_SRAM
rlabel metal4 481436 70516 481436 70516 0 Tile_X11Y16_R_WB_SRAM
rlabel metal3 478193 677620 478193 677620 0 Tile_X11Y2_AD_SRAM0
rlabel metal4 481436 679252 481436 679252 0 Tile_X11Y2_AD_SRAM1
rlabel metal3 478331 681836 478331 681836 0 Tile_X11Y2_AD_SRAM2
rlabel metal3 479516 678300 479516 678300 0 Tile_X11Y2_AD_SRAM3
rlabel via2 478699 678980 478699 678980 0 Tile_X11Y2_AD_SRAM4
rlabel metal3 477469 678844 477469 678844 0 Tile_X11Y2_AD_SRAM5
rlabel metal3 477745 679116 477745 679116 0 Tile_X11Y2_AD_SRAM6
rlabel metal3 477388 679490 477388 679490 0 Tile_X11Y2_AD_SRAM7
rlabel metal3 477871 679796 477871 679796 0 Tile_X11Y2_AD_SRAM8
rlabel metal3 477653 679932 477653 679932 0 Tile_X11Y2_AD_SRAM9
rlabel metal3 477584 680204 477584 680204 0 Tile_X11Y2_BEN_SRAM0
rlabel metal3 478573 680476 478573 680476 0 Tile_X11Y2_BEN_SRAM1
rlabel metal3 477377 682924 477377 682924 0 Tile_X11Y2_BEN_SRAM10
rlabel metal3 480689 683196 480689 683196 0 Tile_X11Y2_BEN_SRAM11
rlabel metal3 477285 683468 477285 683468 0 Tile_X11Y2_BEN_SRAM12
rlabel metal3 483284 740588 483284 740588 0 Tile_X11Y2_BEN_SRAM13
rlabel metal3 483169 700468 483169 700468 0 Tile_X11Y2_BEN_SRAM14
rlabel metal3 478274 684284 478274 684284 0 Tile_X11Y2_BEN_SRAM15
rlabel metal4 483276 685440 483276 685440 0 Tile_X11Y2_BEN_SRAM16
rlabel metal3 478515 684964 478515 684964 0 Tile_X11Y2_BEN_SRAM17
rlabel metal3 483146 718148 483146 718148 0 Tile_X11Y2_BEN_SRAM18
rlabel metal3 478389 685372 478389 685372 0 Tile_X11Y2_BEN_SRAM19
rlabel metal3 477388 680850 477388 680850 0 Tile_X11Y2_BEN_SRAM2
rlabel metal3 482870 717468 482870 717468 0 Tile_X11Y2_BEN_SRAM20
rlabel metal3 478412 685916 478412 685916 0 Tile_X11Y2_BEN_SRAM21
rlabel metal3 478504 686188 478504 686188 0 Tile_X11Y2_BEN_SRAM22
rlabel metal3 482893 716108 482893 716108 0 Tile_X11Y2_BEN_SRAM23
rlabel metal3 484365 698428 484365 698428 0 Tile_X11Y2_BEN_SRAM24
rlabel metal3 483629 715428 483629 715428 0 Tile_X11Y2_BEN_SRAM25
rlabel metal3 483276 687480 483276 687480 0 Tile_X11Y2_BEN_SRAM26
rlabel metal3 483721 714748 483721 714748 0 Tile_X11Y2_BEN_SRAM27
rlabel metal3 483790 742628 483790 742628 0 Tile_X11Y2_BEN_SRAM28
rlabel metal3 481149 688092 481149 688092 0 Tile_X11Y2_BEN_SRAM29
rlabel metal3 483606 727668 483606 727668 0 Tile_X11Y2_BEN_SRAM3
rlabel metal3 483652 752148 483652 752148 0 Tile_X11Y2_BEN_SRAM30
rlabel metal3 477179 688704 477179 688704 0 Tile_X11Y2_BEN_SRAM31
rlabel metal4 484380 681700 484380 681700 0 Tile_X11Y2_BEN_SRAM4
rlabel metal3 483744 728348 483744 728348 0 Tile_X11Y2_BEN_SRAM5
rlabel metal3 485561 683468 485561 683468 0 Tile_X11Y2_BEN_SRAM6
rlabel metal3 483698 743308 483698 743308 0 Tile_X11Y2_BEN_SRAM7
rlabel metal3 483836 729028 483836 729028 0 Tile_X11Y2_BEN_SRAM8
rlabel metal3 483905 705228 483905 705228 0 Tile_X11Y2_BEN_SRAM9
rlabel metal3 483882 732428 483882 732428 0 Tile_X11Y2_CLOCK_SRAM
rlabel metal3 484250 712028 484250 712028 0 Tile_X11Y2_DI_SRAM0
rlabel metal3 477179 689520 477179 689520 0 Tile_X11Y2_DI_SRAM1
rlabel metal3 482249 711348 482249 711348 0 Tile_X11Y2_DI_SRAM10
rlabel metal4 486220 692580 486220 692580 0 Tile_X11Y2_DI_SRAM11
rlabel metal3 484342 750108 484342 750108 0 Tile_X11Y2_DI_SRAM12
rlabel metal3 484664 743988 484664 743988 0 Tile_X11Y2_DI_SRAM13
rlabel metal3 483054 726308 483054 726308 0 Tile_X11Y2_DI_SRAM14
rlabel metal4 477112 702420 477112 702420 0 Tile_X11Y2_DI_SRAM15
rlabel metal3 477179 693600 477179 693600 0 Tile_X11Y2_DI_SRAM16
rlabel metal3 486205 708628 486205 708628 0 Tile_X11Y2_DI_SRAM17
rlabel metal3 484618 744668 484618 744668 0 Tile_X11Y2_DI_SRAM18
rlabel metal3 486021 704548 486021 704548 0 Tile_X11Y2_DI_SRAM19
rlabel metal3 484480 723588 484480 723588 0 Tile_X11Y2_DI_SRAM2
rlabel metal3 484434 730388 484434 730388 0 Tile_X11Y2_DI_SRAM20
rlabel metal3 482341 709308 482341 709308 0 Tile_X11Y2_DI_SRAM21
rlabel metal3 485929 703188 485929 703188 0 Tile_X11Y2_DI_SRAM22
rlabel metal3 484526 731068 484526 731068 0 Tile_X11Y2_DI_SRAM23
rlabel metal3 481858 713388 481858 713388 0 Tile_X11Y2_DI_SRAM24
rlabel metal3 484388 745348 484388 745348 0 Tile_X11Y2_DI_SRAM25
rlabel metal3 484641 699108 484641 699108 0 Tile_X11Y2_DI_SRAM26
rlabel metal3 486113 707948 486113 707948 0 Tile_X11Y2_DI_SRAM27
rlabel metal3 485101 719508 485101 719508 0 Tile_X11Y2_DI_SRAM28
rlabel metal3 485193 722908 485193 722908 0 Tile_X11Y2_DI_SRAM29
rlabel metal3 485285 710668 485285 710668 0 Tile_X11Y2_DI_SRAM3
rlabel metal3 485009 725628 485009 725628 0 Tile_X11Y2_DI_SRAM30
rlabel metal3 477179 697680 477179 697680 0 Tile_X11Y2_DI_SRAM31
rlabel metal3 485170 746028 485170 746028 0 Tile_X11Y2_DI_SRAM4
rlabel metal3 485124 731748 485124 731748 0 Tile_X11Y2_DI_SRAM5
rlabel metal3 485262 733108 485262 733108 0 Tile_X11Y2_DI_SRAM6
rlabel metal3 477837 691084 477837 691084 0 Tile_X11Y2_DI_SRAM7
rlabel metal3 485078 750788 485078 750788 0 Tile_X11Y2_DI_SRAM8
rlabel metal3 479309 691628 479309 691628 0 Tile_X11Y2_DI_SRAM9
rlabel metal4 483552 678300 483552 678300 0 Tile_X11Y2_DO_SRAM0
rlabel metal3 484081 674764 484081 674764 0 Tile_X11Y2_DO_SRAM1
rlabel metal3 483460 684556 483460 684556 0 Tile_X11Y2_DO_SRAM10
rlabel metal3 485032 746708 485032 746708 0 Tile_X11Y2_DO_SRAM11
rlabel metal3 483943 676124 483943 676124 0 Tile_X11Y2_DO_SRAM12
rlabel metal3 486021 681428 486021 681428 0 Tile_X11Y2_DO_SRAM13
rlabel metal4 480976 685780 480976 685780 0 Tile_X11Y2_DO_SRAM14
rlabel metal3 482379 678980 482379 678980 0 Tile_X11Y2_DO_SRAM15
rlabel metal3 481137 676124 481137 676124 0 Tile_X11Y2_DO_SRAM16
rlabel metal3 479665 680340 479665 680340 0 Tile_X11Y2_DO_SRAM17
rlabel metal3 478561 678436 478561 678436 0 Tile_X11Y2_DO_SRAM18
rlabel metal4 483092 675172 483092 675172 0 Tile_X11Y2_DO_SRAM19
rlabel metal3 482011 678164 482011 678164 0 Tile_X11Y2_DO_SRAM2
rlabel metal4 486404 677212 486404 677212 0 Tile_X11Y2_DO_SRAM20
rlabel metal4 484564 678708 484564 678708 0 Tile_X11Y2_DO_SRAM21
rlabel metal3 478389 674764 478389 674764 0 Tile_X11Y2_DO_SRAM22
rlabel metal3 483928 735828 483928 735828 0 Tile_X11Y2_DO_SRAM23
rlabel metal4 483828 677280 483828 677280 0 Tile_X11Y2_DO_SRAM24
rlabel metal4 482172 677960 482172 677960 0 Tile_X11Y2_DO_SRAM25
rlabel metal3 478205 675852 478205 675852 0 Tile_X11Y2_DO_SRAM26
rlabel metal2 486266 741060 486266 741060 0 Tile_X11Y2_DO_SRAM27
rlabel metal4 483092 677484 483092 677484 0 Tile_X11Y2_DO_SRAM28
rlabel metal3 485929 686868 485929 686868 0 Tile_X11Y2_DO_SRAM29
rlabel metal3 479251 677484 479251 677484 0 Tile_X11Y2_DO_SRAM3
rlabel metal3 486274 752828 486274 752828 0 Tile_X11Y2_DO_SRAM30
rlabel metal4 481068 680156 481068 680156 0 Tile_X11Y2_DO_SRAM31
rlabel metal3 486274 737868 486274 737868 0 Tile_X11Y2_DO_SRAM4
rlabel metal3 482241 685780 482241 685780 0 Tile_X11Y2_DO_SRAM5
rlabel metal3 484296 716788 484296 716788 0 Tile_X11Y2_DO_SRAM6
rlabel metal2 482126 716856 482126 716856 0 Tile_X11Y2_DO_SRAM7
rlabel metal3 485745 706588 485745 706588 0 Tile_X11Y2_DO_SRAM8
rlabel metal3 478262 716924 478262 716924 0 Tile_X11Y2_DO_SRAM9
rlabel metal3 485837 705908 485837 705908 0 Tile_X11Y2_EN_SRAM
rlabel metal3 485653 720868 485653 720868 0 Tile_X11Y2_R_WB_SRAM
rlabel metal3 481367 580924 481367 580924 0 Tile_X11Y4_AD_SRAM0
rlabel metal3 483307 587588 483307 587588 0 Tile_X11Y4_AD_SRAM1
rlabel metal3 483721 565148 483721 565148 0 Tile_X11Y4_AD_SRAM2
rlabel metal3 481672 588268 481672 588268 0 Tile_X11Y4_AD_SRAM3
rlabel metal3 484365 564468 484365 564468 0 Tile_X11Y4_AD_SRAM4
rlabel metal3 483629 563788 483629 563788 0 Tile_X11Y4_AD_SRAM5
rlabel metal3 483307 588948 483307 588948 0 Tile_X11Y4_AD_SRAM6
rlabel metal3 485193 563108 485193 563108 0 Tile_X11Y4_AD_SRAM7
rlabel metal3 481672 589628 481672 589628 0 Tile_X11Y4_AD_SRAM8
rlabel metal3 484273 562428 484273 562428 0 Tile_X11Y4_AD_SRAM9
rlabel metal3 483882 561748 483882 561748 0 Tile_X11Y4_BEN_SRAM0
rlabel metal3 483307 590308 483307 590308 0 Tile_X11Y4_BEN_SRAM1
rlabel metal3 485354 557668 485354 557668 0 Tile_X11Y4_BEN_SRAM10
rlabel metal3 483276 593164 483276 593164 0 Tile_X11Y4_BEN_SRAM11
rlabel metal3 483276 593640 483276 593640 0 Tile_X11Y4_BEN_SRAM12
rlabel metal3 481045 603092 481045 603092 0 Tile_X11Y4_BEN_SRAM13
rlabel metal3 482379 601732 482379 601732 0 Tile_X11Y4_BEN_SRAM14
rlabel metal3 477173 594338 477173 594338 0 Tile_X11Y4_BEN_SRAM15
rlabel metal3 483713 607036 483713 607036 0 Tile_X11Y4_BEN_SRAM16
rlabel metal3 483276 595000 483276 595000 0 Tile_X11Y4_BEN_SRAM17
rlabel metal3 480907 604452 480907 604452 0 Tile_X11Y4_BEN_SRAM18
rlabel metal3 482241 607172 482241 607172 0 Tile_X11Y4_BEN_SRAM19
rlabel metal3 484618 561068 484618 561068 0 Tile_X11Y4_BEN_SRAM2
rlabel metal3 477173 595698 477173 595698 0 Tile_X11Y4_BEN_SRAM20
rlabel metal3 483759 607172 483759 607172 0 Tile_X11Y4_BEN_SRAM21
rlabel metal3 485561 596428 485561 596428 0 Tile_X11Y4_BEN_SRAM22
rlabel metal3 484273 626348 484273 626348 0 Tile_X11Y4_BEN_SRAM23
rlabel metal3 483629 625668 483629 625668 0 Tile_X11Y4_BEN_SRAM24
rlabel metal3 477173 597058 477173 597058 0 Tile_X11Y4_BEN_SRAM25
rlabel metal3 477455 597244 477455 597244 0 Tile_X11Y4_BEN_SRAM26
rlabel metal3 481804 597652 481804 597652 0 Tile_X11Y4_BEN_SRAM27
rlabel metal3 477363 597788 477363 597788 0 Tile_X11Y4_BEN_SRAM28
rlabel metal3 477547 598060 477547 598060 0 Tile_X11Y4_BEN_SRAM29
rlabel metal3 481672 590988 481672 590988 0 Tile_X11Y4_BEN_SRAM3
rlabel metal3 477173 598418 477173 598418 0 Tile_X11Y4_BEN_SRAM30
rlabel metal3 477639 598604 477639 598604 0 Tile_X11Y4_BEN_SRAM31
rlabel metal3 485101 560388 485101 560388 0 Tile_X11Y4_BEN_SRAM4
rlabel metal3 484664 559708 484664 559708 0 Tile_X11Y4_BEN_SRAM5
rlabel metal3 483307 591668 483307 591668 0 Tile_X11Y4_BEN_SRAM6
rlabel metal3 485009 559028 485009 559028 0 Tile_X11Y4_BEN_SRAM7
rlabel metal3 481672 592348 481672 592348 0 Tile_X11Y4_BEN_SRAM8
rlabel metal3 483974 558348 483974 558348 0 Tile_X11Y4_BEN_SRAM9
rlabel metal3 484564 599012 484564 599012 0 Tile_X11Y4_CLOCK_SRAM
rlabel metal3 485009 622268 485009 622268 0 Tile_X11Y4_DI_SRAM0
rlabel metal3 477731 599420 477731 599420 0 Tile_X11Y4_DI_SRAM1
rlabel metal3 478191 601868 478191 601868 0 Tile_X11Y4_DI_SRAM10
rlabel metal3 483721 617508 483721 617508 0 Tile_X11Y4_DI_SRAM11
rlabel metal3 478375 602412 478375 602412 0 Tile_X11Y4_DI_SRAM12
rlabel metal3 485032 616828 485032 616828 0 Tile_X11Y4_DI_SRAM13
rlabel metal4 484564 603772 484564 603772 0 Tile_X11Y4_DI_SRAM14
rlabel metal3 486113 619548 486113 619548 0 Tile_X11Y4_DI_SRAM15
rlabel metal3 485837 615468 485837 615468 0 Tile_X11Y4_DI_SRAM16
rlabel metal3 477173 603858 477173 603858 0 Tile_X11Y4_DI_SRAM17
rlabel metal3 486205 614788 486205 614788 0 Tile_X11Y4_DI_SRAM18
rlabel metal3 485561 607988 485561 607988 0 Tile_X11Y4_DI_SRAM19
rlabel metal3 477173 599778 477173 599778 0 Tile_X11Y4_DI_SRAM2
rlabel metal3 483813 614108 483813 614108 0 Tile_X11Y4_DI_SRAM20
rlabel metal3 477823 604860 477823 604860 0 Tile_X11Y4_DI_SRAM21
rlabel metal3 477173 605218 477173 605218 0 Tile_X11Y4_DI_SRAM22
rlabel metal3 485101 618868 485101 618868 0 Tile_X11Y4_DI_SRAM23
rlabel metal3 484089 607308 484089 607308 0 Tile_X11Y4_DI_SRAM24
rlabel metal3 482985 618188 482985 618188 0 Tile_X11Y4_DI_SRAM25
rlabel metal4 482724 608804 482724 608804 0 Tile_X11Y4_DI_SRAM26
rlabel metal3 477173 606578 477173 606578 0 Tile_X11Y4_DI_SRAM27
rlabel metal4 483460 608804 483460 608804 0 Tile_X11Y4_DI_SRAM28
rlabel metal3 484342 620228 484342 620228 0 Tile_X11Y4_DI_SRAM29
rlabel metal4 483460 600304 483460 600304 0 Tile_X11Y4_DI_SRAM3
rlabel metal3 477173 607394 477173 607394 0 Tile_X11Y4_DI_SRAM30
rlabel metal4 486404 608532 486404 608532 0 Tile_X11Y4_DI_SRAM31
rlabel metal3 486021 608668 486021 608668 0 Tile_X11Y4_DI_SRAM4
rlabel metal3 483276 600916 483276 600916 0 Tile_X11Y4_DI_SRAM5
rlabel metal3 483092 601120 483092 601120 0 Tile_X11Y4_DI_SRAM6
rlabel metal4 481436 601800 481436 601800 0 Tile_X11Y4_DI_SRAM7
rlabel metal4 484380 602344 484380 602344 0 Tile_X11Y4_DI_SRAM8
rlabel metal3 485653 605948 485653 605948 0 Tile_X11Y4_DI_SRAM9
rlabel metal3 484457 565828 484457 565828 0 Tile_X11Y4_DO_SRAM0
rlabel metal3 483276 578952 483276 578952 0 Tile_X11Y4_DO_SRAM1
rlabel metal3 481672 581468 481672 581468 0 Tile_X11Y4_DO_SRAM10
rlabel metal3 485837 574668 485837 574668 0 Tile_X11Y4_DO_SRAM11
rlabel metal3 486205 573988 486205 573988 0 Tile_X11Y4_DO_SRAM12
rlabel metal3 483276 582216 483276 582216 0 Tile_X11Y4_DO_SRAM13
rlabel metal3 485929 573308 485929 573308 0 Tile_X11Y4_DO_SRAM14
rlabel metal3 481672 582828 481672 582828 0 Tile_X11Y4_DO_SRAM15
rlabel metal3 477731 583100 477731 583100 0 Tile_X11Y4_DO_SRAM16
rlabel metal3 477823 583372 477823 583372 0 Tile_X11Y4_DO_SRAM17
rlabel metal3 483307 583508 483307 583508 0 Tile_X11Y4_DO_SRAM18
rlabel metal3 477639 583916 477639 583916 0 Tile_X11Y4_DO_SRAM19
rlabel metal4 482908 578680 482908 578680 0 Tile_X11Y4_DO_SRAM2
rlabel metal3 481672 584188 481672 584188 0 Tile_X11Y4_DO_SRAM20
rlabel metal3 485032 570588 485032 570588 0 Tile_X11Y4_DO_SRAM21
rlabel metal3 477064 584732 477064 584732 0 Tile_X11Y4_DO_SRAM22
rlabel metal3 483307 584868 483307 584868 0 Tile_X11Y4_DO_SRAM23
rlabel metal3 477547 585276 477547 585276 0 Tile_X11Y4_DO_SRAM24
rlabel metal3 481672 585548 481672 585548 0 Tile_X11Y4_DO_SRAM25
rlabel metal4 486404 577184 486404 577184 0 Tile_X11Y4_DO_SRAM26
rlabel metal3 482908 586092 482908 586092 0 Tile_X11Y4_DO_SRAM27
rlabel metal3 483276 586296 483276 586296 0 Tile_X11Y4_DO_SRAM28
rlabel metal3 479941 581604 479941 581604 0 Tile_X11Y4_DO_SRAM29
rlabel metal3 483307 579428 483307 579428 0 Tile_X11Y4_DO_SRAM3
rlabel metal3 481672 586908 481672 586908 0 Tile_X11Y4_DO_SRAM30
rlabel metal3 483284 566508 483284 566508 0 Tile_X11Y4_DO_SRAM31
rlabel metal4 477388 578612 477388 578612 0 Tile_X11Y4_DO_SRAM4
rlabel metal3 481672 580108 481672 580108 0 Tile_X11Y4_DO_SRAM5
rlabel metal3 486021 576708 486021 576708 0 Tile_X11Y4_DO_SRAM6
rlabel metal3 485745 576028 485745 576028 0 Tile_X11Y4_DO_SRAM7
rlabel metal3 483307 580788 483307 580788 0 Tile_X11Y4_DO_SRAM8
rlabel metal3 486113 575348 486113 575348 0 Tile_X11Y4_DO_SRAM9
rlabel metal3 483169 616148 483169 616148 0 Tile_X11Y4_EN_SRAM
rlabel metal4 482908 610436 482908 610436 0 Tile_X11Y4_R_WB_SRAM
rlabel metal3 483928 466548 483928 466548 0 Tile_X11Y6_AD_SRAM0
rlabel metal3 483813 475388 483813 475388 0 Tile_X11Y6_AD_SRAM1
rlabel metal3 483307 497828 483307 497828 0 Tile_X11Y6_AD_SRAM2
rlabel metal3 484365 474708 484365 474708 0 Tile_X11Y6_AD_SRAM3
rlabel metal3 477388 498539 477388 498539 0 Tile_X11Y6_AD_SRAM4
rlabel metal3 485101 474028 485101 474028 0 Tile_X11Y6_AD_SRAM5
rlabel metal3 483721 473348 483721 473348 0 Tile_X11Y6_AD_SRAM6
rlabel metal3 483307 499188 483307 499188 0 Tile_X11Y6_AD_SRAM7
rlabel metal3 484273 472668 484273 472668 0 Tile_X11Y6_AD_SRAM8
rlabel metal3 477388 499899 477388 499899 0 Tile_X11Y6_AD_SRAM9
rlabel metal3 485009 471988 485009 471988 0 Tile_X11Y6_BEN_SRAM0
rlabel metal3 483629 471308 483629 471308 0 Tile_X11Y6_BEN_SRAM1
rlabel metal3 484664 467908 484664 467908 0 Tile_X11Y6_BEN_SRAM10
rlabel metal3 485354 467228 485354 467228 0 Tile_X11Y6_BEN_SRAM11
rlabel metal3 483276 503404 483276 503404 0 Tile_X11Y6_BEN_SRAM12
rlabel metal3 483307 503948 483307 503948 0 Tile_X11Y6_BEN_SRAM13
rlabel metal3 483974 539988 483974 539988 0 Tile_X11Y6_BEN_SRAM14
rlabel metal3 484664 539308 484664 539308 0 Tile_X11Y6_BEN_SRAM15
rlabel metal3 477388 504619 477388 504619 0 Tile_X11Y6_BEN_SRAM16
rlabel metal3 483928 538628 483928 538628 0 Tile_X11Y6_BEN_SRAM17
rlabel metal3 483307 505308 483307 505308 0 Tile_X11Y6_BEN_SRAM18
rlabel metal3 483805 514964 483805 514964 0 Tile_X11Y6_BEN_SRAM19
rlabel metal3 483307 500548 483307 500548 0 Tile_X11Y6_BEN_SRAM2
rlabel metal3 482241 516188 482241 516188 0 Tile_X11Y6_BEN_SRAM20
rlabel metal3 477388 505979 477388 505979 0 Tile_X11Y6_BEN_SRAM21
rlabel metal3 483629 536588 483629 536588 0 Tile_X11Y6_BEN_SRAM22
rlabel metal3 483307 506668 483307 506668 0 Tile_X11Y6_BEN_SRAM23
rlabel metal3 483667 516324 483667 516324 0 Tile_X11Y6_BEN_SRAM24
rlabel metal3 484273 535228 484273 535228 0 Tile_X11Y6_BEN_SRAM25
rlabel metal3 477388 507339 477388 507339 0 Tile_X11Y6_BEN_SRAM26
rlabel metal3 478032 507620 478032 507620 0 Tile_X11Y6_BEN_SRAM27
rlabel metal3 477388 507951 477388 507951 0 Tile_X11Y6_BEN_SRAM28
rlabel metal3 477664 508164 477664 508164 0 Tile_X11Y6_BEN_SRAM29
rlabel metal3 484618 470628 484618 470628 0 Tile_X11Y6_BEN_SRAM3
rlabel metal3 477480 508436 477480 508436 0 Tile_X11Y6_BEN_SRAM30
rlabel metal3 477388 508699 477388 508699 0 Tile_X11Y6_BEN_SRAM31
rlabel metal3 477388 501259 477388 501259 0 Tile_X11Y6_BEN_SRAM4
rlabel metal3 485308 469948 485308 469948 0 Tile_X11Y6_BEN_SRAM5
rlabel metal3 483974 469268 483974 469268 0 Tile_X11Y6_BEN_SRAM6
rlabel metal3 483307 501908 483307 501908 0 Tile_X11Y6_BEN_SRAM7
rlabel metal3 482594 468588 482594 468588 0 Tile_X11Y6_BEN_SRAM8
rlabel metal3 477388 502619 477388 502619 0 Tile_X11Y6_BEN_SRAM9
rlabel metal3 477848 508980 477848 508980 0 Tile_X11Y6_CLOCK_SRAM
rlabel metal3 483307 509388 483307 509388 0 Tile_X11Y6_DI_SRAM0
rlabel metal3 485009 531828 485009 531828 0 Tile_X11Y6_DI_SRAM1
rlabel metal3 483721 531148 483721 531148 0 Tile_X11Y6_DI_SRAM10
rlabel metal3 485837 527748 485837 527748 0 Tile_X11Y6_DI_SRAM11
rlabel metal3 483813 527068 483813 527068 0 Tile_X11Y6_DI_SRAM12
rlabel metal4 484380 513536 484380 513536 0 Tile_X11Y6_DI_SRAM13
rlabel metal3 482893 526388 482893 526388 0 Tile_X11Y6_DI_SRAM14
rlabel metal4 479964 515712 479964 515712 0 Tile_X11Y6_DI_SRAM15
rlabel metal3 485745 529108 485745 529108 0 Tile_X11Y6_DI_SRAM16
rlabel metal3 486205 525028 486205 525028 0 Tile_X11Y6_DI_SRAM17
rlabel metal4 483460 514828 483460 514828 0 Tile_X11Y6_DI_SRAM18
rlabel metal3 483077 524348 483077 524348 0 Tile_X11Y6_DI_SRAM19
rlabel metal3 483276 509932 483276 509932 0 Tile_X11Y6_DI_SRAM2
rlabel metal3 482908 514760 482908 514760 0 Tile_X11Y6_DI_SRAM20
rlabel metal3 485101 523668 485101 523668 0 Tile_X11Y6_DI_SRAM21
rlabel metal3 483537 522988 483537 522988 0 Tile_X11Y6_DI_SRAM22
rlabel metal3 485653 518908 485653 518908 0 Tile_X11Y6_DI_SRAM23
rlabel metal4 486312 523940 486312 523940 0 Tile_X11Y6_DI_SRAM24
rlabel metal3 483276 516120 483276 516120 0 Tile_X11Y6_DI_SRAM25
rlabel metal3 485032 530468 485032 530468 0 Tile_X11Y6_DI_SRAM26
rlabel metal3 485469 520948 485469 520948 0 Tile_X11Y6_DI_SRAM27
rlabel metal4 486220 517208 486220 517208 0 Tile_X11Y6_DI_SRAM28
rlabel metal3 485561 520268 485561 520268 0 Tile_X11Y6_DI_SRAM29
rlabel metal4 481436 510748 481436 510748 0 Tile_X11Y6_DI_SRAM3
rlabel metal3 483276 517480 483276 517480 0 Tile_X11Y6_DI_SRAM30
rlabel metal3 485377 519588 485377 519588 0 Tile_X11Y6_DI_SRAM31
rlabel metal3 483276 510544 483276 510544 0 Tile_X11Y6_DI_SRAM4
rlabel metal4 478860 511700 478860 511700 0 Tile_X11Y6_DI_SRAM5
rlabel metal4 484564 512176 484564 512176 0 Tile_X11Y6_DI_SRAM6
rlabel metal4 484380 511632 484380 511632 0 Tile_X11Y6_DI_SRAM7
rlabel metal3 486113 521628 486113 521628 0 Tile_X11Y6_DI_SRAM8
rlabel metal3 483307 516868 483307 516868 0 Tile_X11Y6_DI_SRAM9
rlabel metal3 485929 476068 485929 476068 0 Tile_X11Y6_DO_SRAM0
rlabel metal3 477388 489019 477388 489019 0 Tile_X11Y6_DO_SRAM1
rlabel metal3 484089 484908 484089 484908 0 Tile_X11Y6_DO_SRAM10
rlabel metal3 477388 491739 477388 491739 0 Tile_X11Y6_DO_SRAM11
rlabel metal3 484181 484228 484181 484228 0 Tile_X11Y6_DO_SRAM12
rlabel metal3 482617 483548 482617 483548 0 Tile_X11Y6_DO_SRAM13
rlabel metal3 477388 492487 477388 492487 0 Tile_X11Y6_DO_SRAM14
rlabel metal3 482433 482868 482433 482868 0 Tile_X11Y6_DO_SRAM15
rlabel metal3 477388 493099 477388 493099 0 Tile_X11Y6_DO_SRAM16
rlabel metal3 485193 482188 485193 482188 0 Tile_X11Y6_DO_SRAM17
rlabel metal3 484342 481508 484342 481508 0 Tile_X11Y6_DO_SRAM18
rlabel metal3 483307 493748 483307 493748 0 Tile_X11Y6_DO_SRAM19
rlabel metal4 483276 488852 483276 488852 0 Tile_X11Y6_DO_SRAM2
rlabel metal4 486404 485364 486404 485364 0 Tile_X11Y6_DO_SRAM20
rlabel metal3 477388 494459 477388 494459 0 Tile_X11Y6_DO_SRAM21
rlabel metal3 486205 480148 486205 480148 0 Tile_X11Y6_DO_SRAM22
rlabel metal3 482341 479468 482341 479468 0 Tile_X11Y6_DO_SRAM23
rlabel metal3 477388 495207 477388 495207 0 Tile_X11Y6_DO_SRAM24
rlabel metal3 482249 478788 482249 478788 0 Tile_X11Y6_DO_SRAM25
rlabel metal3 477388 495819 477388 495819 0 Tile_X11Y6_DO_SRAM26
rlabel metal2 486312 480240 486312 480240 0 Tile_X11Y6_DO_SRAM27
rlabel metal3 483238 477428 483238 477428 0 Tile_X11Y6_DO_SRAM28
rlabel metal3 477388 496567 477388 496567 0 Tile_X11Y6_DO_SRAM29
rlabel metal4 484380 488580 484380 488580 0 Tile_X11Y6_DO_SRAM3
rlabel metal3 483284 476748 483284 476748 0 Tile_X11Y6_DO_SRAM30
rlabel metal3 477388 497179 477388 497179 0 Tile_X11Y6_DO_SRAM31
rlabel metal3 485561 489668 485561 489668 0 Tile_X11Y6_DO_SRAM4
rlabel metal3 481881 486948 481881 486948 0 Tile_X11Y6_DO_SRAM5
rlabel metal3 477388 490379 477388 490379 0 Tile_X11Y6_DO_SRAM6
rlabel metal3 485469 486268 485469 486268 0 Tile_X11Y6_DO_SRAM7
rlabel metal3 485653 485588 485653 485588 0 Tile_X11Y6_DO_SRAM8
rlabel metal3 483276 491164 483276 491164 0 Tile_X11Y6_DO_SRAM9
rlabel metal3 485193 525708 485193 525708 0 Tile_X11Y6_EN_SRAM
rlabel metal3 478492 518228 478492 518228 0 Tile_X11Y6_R_WB_SRAM
rlabel metal3 482655 416636 482655 416636 0 Tile_X11Y8_AD_SRAM0
rlabel metal4 484380 408272 484380 408272 0 Tile_X11Y8_AD_SRAM1
rlabel metal3 481672 408068 481672 408068 0 Tile_X11Y8_AD_SRAM2
rlabel metal3 483989 415276 483989 415276 0 Tile_X11Y8_AD_SRAM3
rlabel metal4 482908 409360 482908 409360 0 Tile_X11Y8_AD_SRAM4
rlabel metal3 482425 419628 482425 419628 0 Tile_X11Y8_AD_SRAM5
rlabel metal3 483667 416636 483667 416636 0 Tile_X11Y8_AD_SRAM6
rlabel metal3 481672 409428 481672 409428 0 Tile_X11Y8_AD_SRAM7
rlabel metal3 482195 419764 482195 419764 0 Tile_X11Y8_AD_SRAM8
rlabel metal4 484564 410720 484564 410720 0 Tile_X11Y8_AD_SRAM9
rlabel metal3 483805 423572 483805 423572 0 Tile_X11Y8_BEN_SRAM0
rlabel metal3 477731 410516 477731 410516 0 Tile_X11Y8_BEN_SRAM1
rlabel via3 478699 416636 478699 416636 0 Tile_X11Y8_BEN_SRAM10
rlabel metal3 482456 450908 482456 450908 0 Tile_X11Y8_BEN_SRAM11
rlabel metal4 481436 416704 481436 416704 0 Tile_X11Y8_BEN_SRAM12
rlabel metal3 482502 450228 482502 450228 0 Tile_X11Y8_BEN_SRAM13
rlabel metal4 484564 415140 484564 415140 0 Tile_X11Y8_BEN_SRAM14
rlabel metal3 478009 427244 478009 427244 0 Tile_X11Y8_BEN_SRAM15
rlabel metal3 482609 426156 482609 426156 0 Tile_X11Y8_BEN_SRAM16
rlabel metal3 481672 414868 481672 414868 0 Tile_X11Y8_BEN_SRAM17
rlabel metal3 483667 424932 483667 424932 0 Tile_X11Y8_BEN_SRAM18
rlabel metal4 484380 416160 484380 416160 0 Tile_X11Y8_BEN_SRAM19
rlabel metal3 481672 410788 481672 410788 0 Tile_X11Y8_BEN_SRAM2
rlabel metal3 482249 447508 482249 447508 0 Tile_X11Y8_BEN_SRAM20
rlabel via3 482011 426156 482011 426156 0 Tile_X11Y8_BEN_SRAM21
rlabel metal3 485101 438668 485101 438668 0 Tile_X11Y8_BEN_SRAM22
rlabel metal3 483284 446148 483284 446148 0 Tile_X11Y8_BEN_SRAM23
rlabel metal4 483276 417520 483276 417520 0 Tile_X11Y8_BEN_SRAM24
rlabel metal3 479895 424524 479895 424524 0 Tile_X11Y8_BEN_SRAM25
rlabel metal3 483238 444788 483238 444788 0 Tile_X11Y8_BEN_SRAM26
rlabel metal3 481672 417588 481672 417588 0 Tile_X11Y8_BEN_SRAM27
rlabel via3 479941 427244 479941 427244 0 Tile_X11Y8_BEN_SRAM28
rlabel metal3 478260 418132 478260 418132 0 Tile_X11Y8_BEN_SRAM29
rlabel metal4 484380 411604 484380 411604 0 Tile_X11Y8_BEN_SRAM3
rlabel metal3 482893 443428 482893 443428 0 Tile_X11Y8_BEN_SRAM30
rlabel metal3 482985 442748 482985 442748 0 Tile_X11Y8_BEN_SRAM31
rlabel metal3 485285 413508 485285 413508 0 Tile_X11Y8_BEN_SRAM4
rlabel metal3 478467 411604 478467 411604 0 Tile_X11Y8_BEN_SRAM5
rlabel metal3 483353 412828 483353 412828 0 Tile_X11Y8_BEN_SRAM6
rlabel metal3 483629 423028 483629 423028 0 Tile_X11Y8_BEN_SRAM7
rlabel metal3 486113 420308 486113 420308 0 Tile_X11Y8_BEN_SRAM8
rlabel metal4 484748 414120 484748 414120 0 Tile_X11Y8_BEN_SRAM9
rlabel metal3 481672 418948 481672 418948 0 Tile_X11Y8_CLOCK_SRAM
rlabel metal3 482341 442068 482341 442068 0 Tile_X11Y8_DI_SRAM0
rlabel metal3 485469 423708 485469 423708 0 Tile_X11Y8_DI_SRAM1
rlabel metal3 477823 421940 477823 421940 0 Tile_X11Y8_DI_SRAM10
rlabel metal3 485377 424388 485377 424388 0 Tile_X11Y8_DI_SRAM11
rlabel metal3 485837 437308 485837 437308 0 Tile_X11Y8_DI_SRAM12
rlabel metal4 486220 427348 486220 427348 0 Tile_X11Y8_DI_SRAM13
rlabel metal3 480884 423368 480884 423368 0 Tile_X11Y8_DI_SRAM14
rlabel metal3 485745 435948 485745 435948 0 Tile_X11Y8_DI_SRAM15
rlabel metal3 481068 423504 481068 423504 0 Tile_X11Y8_DI_SRAM16
rlabel metal3 486113 435268 486113 435268 0 Tile_X11Y8_DI_SRAM17
rlabel metal3 483652 453628 483652 453628 0 Tile_X11Y8_DI_SRAM18
rlabel metal4 486404 425272 486404 425272 0 Tile_X11Y8_DI_SRAM19
rlabel metal3 485653 428468 485653 428468 0 Tile_X11Y8_DI_SRAM2
rlabel metal3 485009 452948 485009 452948 0 Tile_X11Y8_DI_SRAM20
rlabel metal2 483138 424728 483138 424728 0 Tile_X11Y8_DI_SRAM21
rlabel metal3 478559 425204 478559 425204 0 Tile_X11Y8_DI_SRAM22
rlabel metal3 477173 425490 477173 425490 0 Tile_X11Y8_DI_SRAM23
rlabel metal3 483629 440028 483629 440028 0 Tile_X11Y8_DI_SRAM24
rlabel metal4 484748 428944 484748 428944 0 Tile_X11Y8_DI_SRAM25
rlabel metal3 484380 426360 484380 426360 0 Tile_X11Y8_DI_SRAM26
rlabel metal4 481620 428876 481620 428876 0 Tile_X11Y8_DI_SRAM27
rlabel metal4 483276 428672 483276 428672 0 Tile_X11Y8_DI_SRAM28
rlabel metal3 481672 427108 481672 427108 0 Tile_X11Y8_DI_SRAM29
rlabel metal3 481413 423572 481413 423572 0 Tile_X11Y8_DI_SRAM3
rlabel metal4 484380 428604 484380 428604 0 Tile_X11Y8_DI_SRAM30
rlabel metal3 477388 427727 477388 427727 0 Tile_X11Y8_DI_SRAM31
rlabel metal3 484273 440708 484273 440708 0 Tile_X11Y8_DI_SRAM4
rlabel metal3 482908 420784 482908 420784 0 Tile_X11Y8_DI_SRAM5
rlabel metal3 482724 420988 482724 420988 0 Tile_X11Y8_DI_SRAM6
rlabel metal3 485561 422348 485561 422348 0 Tile_X11Y8_DI_SRAM7
rlabel metal3 483928 451588 483928 451588 0 Tile_X11Y8_DI_SRAM8
rlabel metal3 486205 433908 486205 433908 0 Tile_X11Y8_DI_SRAM9
rlabel metal3 482962 386308 482962 386308 0 Tile_X11Y8_DO_SRAM0
rlabel metal3 483307 398548 483307 398548 0 Tile_X11Y8_DO_SRAM1
rlabel metal3 483307 401268 483307 401268 0 Tile_X11Y8_DO_SRAM10
rlabel metal4 477388 398106 477388 398106 0 Tile_X11Y8_DO_SRAM11
rlabel metal3 477572 401982 477572 401982 0 Tile_X11Y8_DO_SRAM12
rlabel metal4 483276 398072 483276 398072 0 Tile_X11Y8_DO_SRAM13
rlabel metal3 482249 393108 482249 393108 0 Tile_X11Y8_DO_SRAM14
rlabel metal3 477572 402730 477572 402730 0 Tile_X11Y8_DO_SRAM15
rlabel metal3 483629 392428 483629 392428 0 Tile_X11Y8_DO_SRAM16
rlabel metal3 477572 403342 477572 403342 0 Tile_X11Y8_DO_SRAM17
rlabel metal3 483077 391748 483077 391748 0 Tile_X11Y8_DO_SRAM18
rlabel metal3 482985 391068 482985 391068 0 Tile_X11Y8_DO_SRAM19
rlabel metal3 477572 399262 477572 399262 0 Tile_X11Y8_DO_SRAM2
rlabel metal3 477572 404090 477572 404090 0 Tile_X11Y8_DO_SRAM20
rlabel metal4 486404 391844 486404 391844 0 Tile_X11Y8_DO_SRAM21
rlabel metal3 477572 404702 477572 404702 0 Tile_X11Y8_DO_SRAM22
rlabel metal3 486205 389708 486205 389708 0 Tile_X11Y8_DO_SRAM23
rlabel metal3 482893 389028 482893 389028 0 Tile_X11Y8_DO_SRAM24
rlabel metal3 477572 405450 477572 405450 0 Tile_X11Y8_DO_SRAM25
rlabel metal4 486220 405688 486220 405688 0 Tile_X11Y8_DO_SRAM26
rlabel metal3 477572 406062 477572 406062 0 Tile_X11Y8_DO_SRAM27
rlabel metal3 482548 387668 482548 387668 0 Tile_X11Y8_DO_SRAM28
rlabel metal3 482594 386988 482594 386988 0 Tile_X11Y8_DO_SRAM29
rlabel metal4 478676 398752 478676 398752 0 Tile_X11Y8_DO_SRAM3
rlabel metal3 477572 406810 477572 406810 0 Tile_X11Y8_DO_SRAM30
rlabel metal3 477388 407327 477388 407327 0 Tile_X11Y8_DO_SRAM31
rlabel metal4 484380 398480 484380 398480 0 Tile_X11Y8_DO_SRAM4
rlabel metal3 483307 399908 483307 399908 0 Tile_X11Y8_DO_SRAM5
rlabel metal4 484564 398412 484564 398412 0 Tile_X11Y8_DO_SRAM6
rlabel metal3 477572 400622 477572 400622 0 Tile_X11Y8_DO_SRAM7
rlabel metal4 484748 398412 484748 398412 0 Tile_X11Y8_DO_SRAM8
rlabel metal4 484932 398140 484932 398140 0 Tile_X11Y8_DO_SRAM9
rlabel metal3 486021 439348 486021 439348 0 Tile_X11Y8_EN_SRAM
rlabel metal3 485469 434588 485469 434588 0 Tile_X11Y8_R_WB_SRAM
rlabel metal2 24281 755820 24281 755820 0 Tile_X1Y0_A_I_top
rlabel metal2 23085 755820 23085 755820 0 Tile_X1Y0_A_O_top
rlabel metal2 25109 755820 25109 755820 0 Tile_X1Y0_A_T_top
rlabel metal2 29617 755820 29617 755820 0 Tile_X1Y0_A_config_C_bit0
rlabel metal2 30813 755820 30813 755820 0 Tile_X1Y0_A_config_C_bit1
rlabel metal2 32009 755820 32009 755820 0 Tile_X1Y0_A_config_C_bit2
rlabel metal2 32837 755820 32837 755820 0 Tile_X1Y0_A_config_C_bit3
rlabel metal2 27547 755820 27547 755820 0 Tile_X1Y0_B_I_top
rlabel metal2 26351 755820 26351 755820 0 Tile_X1Y0_B_O_top
rlabel metal2 28743 755820 28743 755820 0 Tile_X1Y0_B_T_top
rlabel metal2 34079 755820 34079 755820 0 Tile_X1Y0_B_config_C_bit0
rlabel metal2 35275 755820 35275 755820 0 Tile_X1Y0_B_config_C_bit1
rlabel metal2 36163 755820 36163 755820 0 Tile_X1Y0_B_config_C_bit2
rlabel metal2 37345 755820 37345 755820 0 Tile_X1Y0_B_config_C_bit3
rlabel metal2 23230 823 23230 823 0 Tile_X1Y17_IRQ_top0
rlabel metal2 24518 3388 24518 3388 0 Tile_X1Y17_IRQ_top1
rlabel metal2 26082 3381 26082 3381 0 Tile_X1Y17_IRQ_top2
rlabel metal2 27738 1163 27738 1163 0 Tile_X1Y17_IRQ_top3
rlabel metal2 65037 755820 65037 755820 0 Tile_X2Y0_A_I_top
rlabel metal2 63901 755820 63901 755820 0 Tile_X2Y0_A_O_top
rlabel metal2 66279 755820 66279 755820 0 Tile_X2Y0_A_T_top
rlabel metal2 70741 755820 70741 755820 0 Tile_X2Y0_A_config_C_bit0
rlabel metal2 71629 755820 71629 755820 0 Tile_X2Y0_A_config_C_bit1
rlabel metal2 72765 755820 72765 755820 0 Tile_X2Y0_A_config_C_bit2
rlabel metal2 74007 755820 74007 755820 0 Tile_X2Y0_A_config_C_bit3
rlabel metal2 68363 755820 68363 755820 0 Tile_X2Y0_B_I_top
rlabel metal2 67167 755820 67167 755820 0 Tile_X2Y0_B_O_top
rlabel metal2 69545 755820 69545 755820 0 Tile_X2Y0_B_T_top
rlabel metal2 74895 755820 74895 755820 0 Tile_X2Y0_B_config_C_bit0
rlabel metal2 76091 755820 76091 755820 0 Tile_X2Y0_B_config_C_bit1
rlabel metal2 77273 755820 77273 755820 0 Tile_X2Y0_B_config_C_bit2
rlabel metal2 78469 755820 78469 755820 0 Tile_X2Y0_B_config_C_bit3
rlabel metal2 65056 5897 65056 5897 0 Tile_X2Y17_BOOT_top
rlabel metal2 63584 5897 63584 5897 0 Tile_X2Y17_RESET_top
rlabel metal2 66378 3271 66378 3271 0 Tile_X2Y17_SLOT_top0
rlabel metal2 68000 5897 68000 5897 0 Tile_X2Y17_SLOT_top1
rlabel metal2 69472 5897 69472 5897 0 Tile_X2Y17_SLOT_top2
rlabel metal2 70886 3271 70886 3271 0 Tile_X2Y17_SLOT_top3
rlabel metal2 155151 755820 155151 755820 0 Tile_X4Y0_A_I_top
rlabel metal2 153909 755820 153909 755820 0 Tile_X4Y0_A_O_top
rlabel metal2 155841 755820 155841 755820 0 Tile_X4Y0_A_T_top
rlabel metal2 160501 755820 160501 755820 0 Tile_X4Y0_A_config_C_bit0
rlabel metal2 161637 755820 161637 755820 0 Tile_X4Y0_A_config_C_bit1
rlabel metal2 162879 755820 162879 755820 0 Tile_X4Y0_A_config_C_bit2
rlabel metal2 163767 755820 163767 755820 0 Tile_X4Y0_A_config_C_bit3
rlabel metal2 158417 755820 158417 755820 0 Tile_X4Y0_B_I_top
rlabel metal2 157235 755820 157235 755820 0 Tile_X4Y0_B_O_top
rlabel metal2 159613 755820 159613 755820 0 Tile_X4Y0_B_T_top
rlabel metal2 164963 755820 164963 755820 0 Tile_X4Y0_B_config_C_bit0
rlabel metal2 166145 755820 166145 755820 0 Tile_X4Y0_B_config_C_bit1
rlabel metal2 167341 755820 167341 755820 0 Tile_X4Y0_B_config_C_bit2
rlabel metal2 168229 755820 168229 755820 0 Tile_X4Y0_B_config_C_bit3
rlabel metal2 165554 1911 165554 1911 0 Tile_X4Y17_I_top0
rlabel metal2 166198 1911 166198 1911 0 Tile_X4Y17_I_top1
rlabel metal2 172720 5897 172720 5897 0 Tile_X4Y17_I_top10
rlabel metal2 173456 5897 173456 5897 0 Tile_X4Y17_I_top11
rlabel metal2 174202 3381 174202 3381 0 Tile_X4Y17_I_top12
rlabel metal2 175214 823 175214 823 0 Tile_X4Y17_I_top13
rlabel metal2 175858 1911 175858 1911 0 Tile_X4Y17_I_top14
rlabel metal2 176502 1911 176502 1911 0 Tile_X4Y17_I_top15
rlabel metal2 166842 3388 166842 3388 0 Tile_X4Y17_I_top2
rlabel metal2 167568 5897 167568 5897 0 Tile_X4Y17_I_top3
rlabel metal2 168304 5897 168304 5897 0 Tile_X4Y17_I_top4
rlabel metal2 169050 3381 169050 3381 0 Tile_X4Y17_I_top5
rlabel metal2 170062 823 170062 823 0 Tile_X4Y17_I_top6
rlabel metal2 170706 1911 170706 1911 0 Tile_X4Y17_I_top7
rlabel metal2 171350 1911 171350 1911 0 Tile_X4Y17_I_top8
rlabel metal2 171994 3388 171994 3388 0 Tile_X4Y17_I_top9
rlabel metal2 153594 3381 153594 3381 0 Tile_X4Y17_O_top0
rlabel metal2 154606 823 154606 823 0 Tile_X4Y17_O_top1
rlabel metal2 161046 1911 161046 1911 0 Tile_X4Y17_O_top10
rlabel metal2 161690 3388 161690 3388 0 Tile_X4Y17_O_top11
rlabel metal2 162416 5897 162416 5897 0 Tile_X4Y17_O_top12
rlabel metal2 163152 5897 163152 5897 0 Tile_X4Y17_O_top13
rlabel metal2 163898 3381 163898 3381 0 Tile_X4Y17_O_top14
rlabel metal2 164910 823 164910 823 0 Tile_X4Y17_O_top15
rlabel metal2 155250 1911 155250 1911 0 Tile_X4Y17_O_top2
rlabel metal2 155894 1911 155894 1911 0 Tile_X4Y17_O_top3
rlabel metal2 156538 3388 156538 3388 0 Tile_X4Y17_O_top4
rlabel metal2 157264 5897 157264 5897 0 Tile_X4Y17_O_top5
rlabel metal2 158000 5897 158000 5897 0 Tile_X4Y17_O_top6
rlabel metal2 158736 5897 158736 5897 0 Tile_X4Y17_O_top7
rlabel metal2 159758 823 159758 823 0 Tile_X4Y17_O_top8
rlabel metal2 160402 1911 160402 1911 0 Tile_X4Y17_O_top9
rlabel metal2 195875 755820 195875 755820 0 Tile_X5Y0_A_I_top
rlabel metal2 195079 755820 195079 755820 0 Tile_X5Y0_A_O_top
rlabel metal2 197163 755820 197163 755820 0 Tile_X5Y0_A_T_top
rlabel metal2 201565 755820 201565 755820 0 Tile_X5Y0_A_config_C_bit0
rlabel metal2 202807 755820 202807 755820 0 Tile_X5Y0_A_config_C_bit1
rlabel metal2 203695 755820 203695 755820 0 Tile_X5Y0_A_config_C_bit2
rlabel metal2 204891 755820 204891 755820 0 Tile_X5Y0_A_config_C_bit3
rlabel metal2 199541 755820 199541 755820 0 Tile_X5Y0_B_I_top
rlabel metal2 198345 755820 198345 755820 0 Tile_X5Y0_B_O_top
rlabel metal2 200429 755820 200429 755820 0 Tile_X5Y0_B_T_top
rlabel metal2 206073 755820 206073 755820 0 Tile_X5Y0_B_config_C_bit0
rlabel metal2 207269 755820 207269 755820 0 Tile_X5Y0_B_config_C_bit1
rlabel metal2 208157 755820 208157 755820 0 Tile_X5Y0_B_config_C_bit2
rlabel metal2 209293 755820 209293 755820 0 Tile_X5Y0_B_config_C_bit3
rlabel metal2 206126 3271 206126 3271 0 Tile_X5Y17_I_top0
rlabel metal2 207096 5897 207096 5897 0 Tile_X5Y17_I_top1
rlabel metal2 213720 5897 213720 5897 0 Tile_X5Y17_I_top10
rlabel metal2 214456 5897 214456 5897 0 Tile_X5Y17_I_top11
rlabel metal2 215142 3271 215142 3271 0 Tile_X5Y17_I_top12
rlabel metal2 215786 3271 215786 3271 0 Tile_X5Y17_I_top13
rlabel metal2 216430 3271 216430 3271 0 Tile_X5Y17_I_top14
rlabel metal2 217400 5897 217400 5897 0 Tile_X5Y17_I_top15
rlabel metal2 207832 5897 207832 5897 0 Tile_X5Y17_I_top2
rlabel metal2 208568 5897 208568 5897 0 Tile_X5Y17_I_top3
rlabel metal2 209304 5897 209304 5897 0 Tile_X5Y17_I_top4
rlabel metal2 209990 3271 209990 3271 0 Tile_X5Y17_I_top5
rlabel metal2 210634 3271 210634 3271 0 Tile_X5Y17_I_top6
rlabel metal2 211278 3271 211278 3271 0 Tile_X5Y17_I_top7
rlabel metal2 212248 5897 212248 5897 0 Tile_X5Y17_I_top8
rlabel metal2 212984 5897 212984 5897 0 Tile_X5Y17_I_top9
rlabel metal2 194534 3271 194534 3271 0 Tile_X5Y17_O_top0
rlabel metal2 195178 3271 195178 3271 0 Tile_X5Y17_O_top1
rlabel metal2 201944 5897 201944 5897 0 Tile_X5Y17_O_top10
rlabel metal2 202680 5897 202680 5897 0 Tile_X5Y17_O_top11
rlabel metal2 203416 5897 203416 5897 0 Tile_X5Y17_O_top12
rlabel metal2 204152 5897 204152 5897 0 Tile_X5Y17_O_top13
rlabel metal2 204838 3271 204838 3271 0 Tile_X5Y17_O_top14
rlabel metal2 205482 3271 205482 3271 0 Tile_X5Y17_O_top15
rlabel metal2 195822 3271 195822 3271 0 Tile_X5Y17_O_top2
rlabel metal2 196792 5897 196792 5897 0 Tile_X5Y17_O_top3
rlabel metal2 197528 5897 197528 5897 0 Tile_X5Y17_O_top4
rlabel metal2 198264 5897 198264 5897 0 Tile_X5Y17_O_top5
rlabel metal2 199000 5897 199000 5897 0 Tile_X5Y17_O_top6
rlabel metal2 199686 3271 199686 3271 0 Tile_X5Y17_O_top7
rlabel metal2 200330 3271 200330 3271 0 Tile_X5Y17_O_top8
rlabel metal2 200974 3271 200974 3271 0 Tile_X5Y17_O_top9
rlabel metal2 237091 755820 237091 755820 0 Tile_X6Y0_A_I_top
rlabel metal2 235849 755820 235849 755820 0 Tile_X6Y0_A_O_top
rlabel metal2 238273 755820 238273 755820 0 Tile_X6Y0_A_T_top
rlabel metal2 242735 755820 242735 755820 0 Tile_X6Y0_A_config_C_bit0
rlabel metal2 243623 755820 243623 755820 0 Tile_X6Y0_A_config_C_bit1
rlabel metal2 244819 755820 244819 755820 0 Tile_X6Y0_A_config_C_bit2
rlabel metal2 246001 755820 246001 755820 0 Tile_X6Y0_A_config_C_bit3
rlabel metal2 240357 755820 240357 755820 0 Tile_X6Y0_B_I_top
rlabel metal2 239161 755820 239161 755820 0 Tile_X6Y0_B_O_top
rlabel metal2 241493 755820 241493 755820 0 Tile_X6Y0_B_T_top
rlabel metal2 246843 755820 246843 755820 0 Tile_X6Y0_B_config_C_bit0
rlabel metal2 248085 755820 248085 755820 0 Tile_X6Y0_B_config_C_bit1
rlabel metal2 249221 755820 249221 755820 0 Tile_X6Y0_B_config_C_bit2
rlabel metal2 250463 755820 250463 755820 0 Tile_X6Y0_B_config_C_bit3
rlabel metal2 247342 3388 247342 3388 0 Tile_X6Y17_I_top0
rlabel metal2 247986 1911 247986 1911 0 Tile_X6Y17_I_top1
rlabel metal2 254426 823 254426 823 0 Tile_X6Y17_I_top10
rlabel metal2 255484 5897 255484 5897 0 Tile_X6Y17_I_top11
rlabel metal2 256220 5897 256220 5897 0 Tile_X6Y17_I_top12
rlabel metal2 256956 5897 256956 5897 0 Tile_X6Y17_I_top13
rlabel metal2 257646 3388 257646 3388 0 Tile_X6Y17_I_top14
rlabel metal2 258290 1911 258290 1911 0 Tile_X6Y17_I_top15
rlabel metal2 248630 1231 248630 1231 0 Tile_X6Y17_I_top2
rlabel metal2 249274 823 249274 823 0 Tile_X6Y17_I_top3
rlabel metal2 250332 5897 250332 5897 0 Tile_X6Y17_I_top4
rlabel metal2 251068 5897 251068 5897 0 Tile_X6Y17_I_top5
rlabel metal2 251804 5897 251804 5897 0 Tile_X6Y17_I_top6
rlabel metal2 252494 3388 252494 3388 0 Tile_X6Y17_I_top7
rlabel metal2 253138 1911 253138 1911 0 Tile_X6Y17_I_top8
rlabel metal2 253782 3203 253782 3203 0 Tile_X6Y17_I_top9
rlabel metal2 235750 3271 235750 3271 0 Tile_X6Y17_O_top0
rlabel metal2 236348 5897 236348 5897 0 Tile_X6Y17_O_top1
rlabel metal2 242834 3203 242834 3203 0 Tile_X6Y17_O_top10
rlabel metal2 243478 1231 243478 1231 0 Tile_X6Y17_O_top11
rlabel metal2 244122 3203 244122 3203 0 Tile_X6Y17_O_top12
rlabel metal2 245180 5897 245180 5897 0 Tile_X6Y17_O_top13
rlabel metal2 245916 5897 245916 5897 0 Tile_X6Y17_O_top14
rlabel metal2 246652 5897 246652 5897 0 Tile_X6Y17_O_top15
rlabel metal2 237038 3388 237038 3388 0 Tile_X6Y17_O_top2
rlabel metal2 237682 1911 237682 1911 0 Tile_X6Y17_O_top3
rlabel metal2 238326 1231 238326 1231 0 Tile_X6Y17_O_top4
rlabel metal2 238970 823 238970 823 0 Tile_X6Y17_O_top5
rlabel metal2 240028 5897 240028 5897 0 Tile_X6Y17_O_top6
rlabel metal2 240764 5897 240764 5897 0 Tile_X6Y17_O_top7
rlabel metal2 241454 3653 241454 3653 0 Tile_X6Y17_O_top8
rlabel metal2 242190 3388 242190 3388 0 Tile_X6Y17_O_top9
rlabel metal2 323189 755820 323189 755820 0 Tile_X8Y0_A_I_top
rlabel metal2 321993 755820 321993 755820 0 Tile_X8Y0_A_O_top
rlabel metal2 324077 755820 324077 755820 0 Tile_X8Y0_A_T_top
rlabel metal2 328539 755820 328539 755820 0 Tile_X8Y0_A_config_C_bit0
rlabel metal2 329721 755820 329721 755820 0 Tile_X8Y0_A_config_C_bit1
rlabel metal2 330917 755820 330917 755820 0 Tile_X8Y0_A_config_C_bit2
rlabel metal2 331805 755820 331805 755820 0 Tile_X8Y0_A_config_C_bit3
rlabel metal2 326455 755820 326455 755820 0 Tile_X8Y0_B_I_top
rlabel metal2 325213 755820 325213 755820 0 Tile_X8Y0_B_O_top
rlabel metal2 327343 755820 327343 755820 0 Tile_X8Y0_B_T_top
rlabel metal2 332941 755820 332941 755820 0 Tile_X8Y0_B_config_C_bit0
rlabel metal2 334183 755820 334183 755820 0 Tile_X8Y0_B_config_C_bit1
rlabel metal2 335071 755820 335071 755820 0 Tile_X8Y0_B_config_C_bit2
rlabel metal2 336267 755820 336267 755820 0 Tile_X8Y0_B_config_C_bit3
rlabel metal2 333638 823 333638 823 0 Tile_X8Y17_I_top0
rlabel metal2 334282 1911 334282 1911 0 Tile_X8Y17_I_top1
rlabel metal2 340722 3388 340722 3388 0 Tile_X8Y17_I_top10
rlabel metal2 341456 5897 341456 5897 0 Tile_X8Y17_I_top11
rlabel metal2 342192 5897 342192 5897 0 Tile_X8Y17_I_top12
rlabel metal2 342930 3381 342930 3381 0 Tile_X8Y17_I_top13
rlabel metal2 343942 823 343942 823 0 Tile_X8Y17_I_top14
rlabel metal2 344586 1911 344586 1911 0 Tile_X8Y17_I_top15
rlabel metal2 334926 1911 334926 1911 0 Tile_X8Y17_I_top2
rlabel metal2 335570 3388 335570 3388 0 Tile_X8Y17_I_top3
rlabel metal2 336304 5897 336304 5897 0 Tile_X8Y17_I_top4
rlabel metal2 337040 5897 337040 5897 0 Tile_X8Y17_I_top5
rlabel metal2 337778 3381 337778 3381 0 Tile_X8Y17_I_top6
rlabel metal2 338790 823 338790 823 0 Tile_X8Y17_I_top7
rlabel metal2 339434 1911 339434 1911 0 Tile_X8Y17_I_top8
rlabel metal2 340078 1911 340078 1911 0 Tile_X8Y17_I_top9
rlabel metal2 321584 5897 321584 5897 0 Tile_X8Y17_O_top0
rlabel metal2 322322 3381 322322 3381 0 Tile_X8Y17_O_top1
rlabel metal2 329130 1911 329130 1911 0 Tile_X8Y17_O_top10
rlabel metal2 329774 1911 329774 1911 0 Tile_X8Y17_O_top11
rlabel metal2 330418 3388 330418 3388 0 Tile_X8Y17_O_top12
rlabel metal2 331152 5897 331152 5897 0 Tile_X8Y17_O_top13
rlabel metal2 331888 5897 331888 5897 0 Tile_X8Y17_O_top14
rlabel metal2 332624 5897 332624 5897 0 Tile_X8Y17_O_top15
rlabel metal2 323334 823 323334 823 0 Tile_X8Y17_O_top2
rlabel metal2 323978 1911 323978 1911 0 Tile_X8Y17_O_top3
rlabel metal2 324622 1911 324622 1911 0 Tile_X8Y17_O_top4
rlabel metal2 325266 3388 325266 3388 0 Tile_X8Y17_O_top5
rlabel metal2 326000 5897 326000 5897 0 Tile_X8Y17_O_top6
rlabel metal2 326736 5897 326736 5897 0 Tile_X8Y17_O_top7
rlabel metal2 327474 3381 327474 3381 0 Tile_X8Y17_O_top8
rlabel metal2 328486 823 328486 823 0 Tile_X8Y17_O_top9
rlabel metal2 364005 755820 364005 755820 0 Tile_X9Y0_A_I_top
rlabel metal2 363117 755820 363117 755820 0 Tile_X9Y0_A_O_top
rlabel metal2 365141 755820 365141 755820 0 Tile_X9Y0_A_T_top
rlabel metal2 369649 755820 369649 755820 0 Tile_X9Y0_A_config_C_bit0
rlabel metal2 370845 755820 370845 755820 0 Tile_X9Y0_A_config_C_bit1
rlabel metal2 371733 755820 371733 755820 0 Tile_X9Y0_A_config_C_bit2
rlabel metal2 372869 755820 372869 755820 0 Tile_X9Y0_A_config_C_bit3
rlabel metal2 367271 755820 367271 755820 0 Tile_X9Y0_B_I_top
rlabel metal2 366383 755820 366383 755820 0 Tile_X9Y0_B_O_top
rlabel metal2 368361 755820 368361 755820 0 Tile_X9Y0_B_T_top
rlabel metal2 374111 755820 374111 755820 0 Tile_X9Y0_B_config_C_bit0
rlabel metal2 374999 755820 374999 755820 0 Tile_X9Y0_B_config_C_bit1
rlabel metal2 376195 755820 376195 755820 0 Tile_X9Y0_B_config_C_bit2
rlabel metal2 377377 755820 377377 755820 0 Tile_X9Y0_B_config_C_bit3
rlabel metal2 362400 5897 362400 5897 0 Tile_X9Y17_CMP_top
rlabel metal2 363262 3271 363262 3271 0 Tile_X9Y17_HOLD_top
rlabel metal2 364550 3271 364550 3271 0 Tile_X9Y17_RESET_top
rlabel metal2 365712 5897 365712 5897 0 Tile_X9Y17_VALUE_top0
rlabel metal2 366816 5897 366816 5897 0 Tile_X9Y17_VALUE_top1
rlabel metal2 376752 5897 376752 5897 0 Tile_X9Y17_VALUE_top10
rlabel metal2 377856 5897 377856 5897 0 Tile_X9Y17_VALUE_top11
rlabel metal2 367770 3271 367770 3271 0 Tile_X9Y17_VALUE_top2
rlabel metal2 369024 5897 369024 5897 0 Tile_X9Y17_VALUE_top3
rlabel metal2 370128 5897 370128 5897 0 Tile_X9Y17_VALUE_top4
rlabel metal2 370990 3271 370990 3271 0 Tile_X9Y17_VALUE_top5
rlabel metal2 372278 3271 372278 3271 0 Tile_X9Y17_VALUE_top6
rlabel metal2 373440 5897 373440 5897 0 Tile_X9Y17_VALUE_top7
rlabel metal2 374544 5897 374544 5897 0 Tile_X9Y17_VALUE_top8
rlabel metal2 375498 3271 375498 3271 0 Tile_X9Y17_VALUE_top9
rlabel metal2 177136 5965 177136 5965 0 UserCLK
<< properties >>
string FIXED_BBOX 0 0 487000 756500
<< end >>
