`default_nettype none

module fabric_wrapper #(
    	parameter FrameBitsPerRow = 32,
	parameter MaxFramesPerCol = 20,
	
	parameter NumColumns = 12,
	parameter NumRows = 18,
	
    parameter FABRIC_NUM_IO_WEST = 32,
    parameter FABRIC_NUM_IO_NORTH = 16
)(
    input clk_i,
    
    // Configuration
    input  logic [(FrameBitsPerRow*NumRows)-1:0]    FrameData_i,
    input  logic [(MaxFramesPerCol*NumColumns)-1:0] FrameStrobe_i,
    
    // I/Os West
    input  [FABRIC_NUM_IO_WEST-1:0]      fabric_io_west_in_i,
    output [FABRIC_NUM_IO_WEST-1:0]      fabric_io_west_out_o,
    output [FABRIC_NUM_IO_WEST-1:0]      fabric_io_west_oeb_o,

    // I/O West config
    output [FABRIC_NUM_IO_WEST-1:0]      fabric_io_west_config_bit0_o,
    output [FABRIC_NUM_IO_WEST-1:0]      fabric_io_west_config_bit1_o,
    output [FABRIC_NUM_IO_WEST-1:0]      fabric_io_west_config_bit2_o,
    output [FABRIC_NUM_IO_WEST-1:0]      fabric_io_west_config_bit3_o,

    // I/Os North
    input  [FABRIC_NUM_IO_NORTH-1:0]      fabric_io_north_in_i,
    output [FABRIC_NUM_IO_NORTH-1:0]      fabric_io_north_out_o,
    output [FABRIC_NUM_IO_NORTH-1:0]      fabric_io_north_oeb_o,

    // I/O North config
    output [FABRIC_NUM_IO_NORTH-1:0]      fabric_io_north_config_bit0_o,
    output [FABRIC_NUM_IO_NORTH-1:0]      fabric_io_north_config_bit1_o,
    output [FABRIC_NUM_IO_NORTH-1:0]      fabric_io_north_config_bit2_o,
    output [FABRIC_NUM_IO_NORTH-1:0]      fabric_io_north_config_bit3_o,

    // ADC
    input         fabric_adc0_cmp_i,
    output        fabric_adc0_hold_o,
    output        fabric_adc0_reset_o,
    output [11:0] fabric_adc0_value_o,

    // DAC
    output [7:0] fabric_dac0_value_o,

    // SRAM 0
    input  [31:0] fabric_sram0_do_i,
    output [9 :0] fabric_sram0_ad_o,
    output [31:0] fabric_sram0_ben_o,
    output [31:0] fabric_sram0_di_o,
    output        fabric_sram0_en_o,
    output        fabric_sram0_rw_no,
    output        fabric_sram0_clk_o,

    // SRAM 1
    input  [31:0] fabric_sram1_do_i,
    output [9 :0] fabric_sram1_ad_o,
    output [31:0] fabric_sram1_ben_o,
    output [31:0] fabric_sram1_di_o,
    output        fabric_sram1_en_o,
    output        fabric_sram1_rw_no,
    output        fabric_sram1_clk_o,

    // SRAM 2
    input  [31:0] fabric_sram2_do_i,
    output [9 :0] fabric_sram2_ad_o,
    output [31:0] fabric_sram2_ben_o,
    output [31:0] fabric_sram2_di_o,
    output        fabric_sram2_en_o,
    output        fabric_sram2_rw_no,
    output        fabric_sram2_clk_o,

    // SRAM 3
    input  [31:0] fabric_sram3_do_i,
    output [9 :0] fabric_sram3_ad_o,
    output [31:0] fabric_sram3_ben_o,
    output [31:0] fabric_sram3_di_o,
    output        fabric_sram3_en_o,
    output        fabric_sram3_rw_no,
    output        fabric_sram3_clk_o,

    // SRAM 4
    input  [31:0] fabric_sram4_do_i,
    output [9 :0] fabric_sram4_ad_o,
    output [31:0] fabric_sram4_ben_o,
    output [31:0] fabric_sram4_di_o,
    output        fabric_sram4_en_o,
    output        fabric_sram4_rw_no,
    output        fabric_sram4_clk_o,

    // SRAM 5
    input  [31:0] fabric_sram5_do_i,
    output [9 :0] fabric_sram5_ad_o,
    output [31:0] fabric_sram5_ben_o,
    output [31:0] fabric_sram5_di_o,
    output        fabric_sram5_en_o,
    output        fabric_sram5_rw_no,
    output        fabric_sram5_clk_o,

    // SRAM 6
    input  [31:0] fabric_sram6_do_i,
    output [9 :0] fabric_sram6_ad_o,
    output [31:0] fabric_sram6_ben_o,
    output [31:0] fabric_sram6_di_o,
    output        fabric_sram6_en_o,
    output        fabric_sram6_rw_no,
    output        fabric_sram6_clk_o,

    // SRAM 7
    input  [31:0] fabric_sram7_do_i,
    output [9 :0] fabric_sram7_ad_o,
    output [31:0] fabric_sram7_ben_o,
    output [31:0] fabric_sram7_di_o,
    output        fabric_sram7_en_o,
    output        fabric_sram7_rw_no,
    output        fabric_sram7_clk_o,

    // WARMBOOT
    output        fabric_warmboot_boot_o,
    output  [3:0] fabric_warmboot_slot_o,
    input         fabric_warmboot_reset_i,

    // CPU_IRQ
    output  [3:0] fabric_irq_o,
    
    // CPU_IF - Selector
    input  logic            fabric_xif_or_periph_i,
    
    // Custom instruction interface
    input  logic [31:0]     fabric_rs1_i,
    input  logic [31:0]     fabric_rs2_i,
    output logic [31:0]     fabric_result_o,
    
    // Bus interface
    output logic            fabric_gnt_o,
    input  logic            fabric_req_i,
    output logic            fabric_rvalid_o,
    input  logic            fabric_we_i,
    input  logic [ 3:0]     fabric_be_i,
    input  logic [23:0]     fabric_addr_i,
    input  logic [31:0]     fabric_wdata_i,
    output logic [31:0]     fabric_rdata_o
);
    
    logic [63:0] fabric_cpu_i;
    logic [63:0] fabric_cpu_o;
    
    // CPU_IF muxing
    always_comb begin
        // Custom instruction interface selected
        if (fabric_xif_or_periph_i == 1'b0) begin
            // XIF connected to CPU_IF
            fabric_cpu_i    = {fabric_rs2_i, fabric_rs1_i};
            fabric_result_o = fabric_cpu_o[31:0];

            // Default values for peripheral
            fabric_gnt_o    = fabric_req_i;
            fabric_rvalid_o = fabric_req_i;
            fabric_rdata_o  = 32'hDEADBEEF;

        // Bus interface selected
        end else begin
            // Periperhal connected to CPU_IF
            fabric_cpu_i = {2'b0, fabric_req_i, fabric_we_i, fabric_be_i, fabric_addr_i, fabric_wdata_i};

            fabric_gnt_o    = fabric_cpu_o[33];
            fabric_rvalid_o = fabric_cpu_o[32];
            fabric_rdata_o  = fabric_cpu_o[31:0];

            // Default value for XIF
            fabric_result_o = 32'hDEADBEEF;
        end
    end
    
    // Gated signals:
    // Make sure those signals can not trigger
    // while the fabric is configured
    
    logic fabric_sram0_en;
    logic fabric_sram1_en;
    logic fabric_sram2_en;
    logic fabric_sram3_en;
    logic fabric_sram4_en;
    logic fabric_sram5_en;
    logic fabric_sram6_en;
    logic fabric_sram7_en;
    
    assign fabric_sram0_en_o = fabric_sram0_en && !fabric_warmboot_reset_i;
    assign fabric_sram1_en_o = fabric_sram1_en && !fabric_warmboot_reset_i;
    assign fabric_sram2_en_o = fabric_sram2_en && !fabric_warmboot_reset_i;
    assign fabric_sram3_en_o = fabric_sram3_en && !fabric_warmboot_reset_i;
    assign fabric_sram4_en_o = fabric_sram4_en && !fabric_warmboot_reset_i;
    assign fabric_sram5_en_o = fabric_sram5_en && !fabric_warmboot_reset_i;
    assign fabric_sram6_en_o = fabric_sram6_en && !fabric_warmboot_reset_i;
    assign fabric_sram7_en_o = fabric_sram7_en && !fabric_warmboot_reset_i;
    
    logic [3:0] fabric_irq;
    
    assign fabric_irq_o[0] = fabric_irq[0] && !fabric_warmboot_reset_i;
    assign fabric_irq_o[1] = fabric_irq[1] && !fabric_warmboot_reset_i;
    assign fabric_irq_o[2] = fabric_irq[2] && !fabric_warmboot_reset_i;
    assign fabric_irq_o[3] = fabric_irq[3] && !fabric_warmboot_reset_i;
    
    logic fabric_warmboot_boot;
    
    assign fabric_warmboot_boot_o = fabric_warmboot_boot && !fabric_warmboot_reset_i;
    
    eFPGA
    //#(
    //    .MaxFramesPerCol(MaxFramesPerCol),
    //    .FrameBitsPerRow(FrameBitsPerRow)
    //)
    eFPGA
    (
        .FrameData      (FrameData_i),
        .FrameStrobe    (FrameStrobe_i),
        .UserCLK        (clk_i),
        
        // West I/Os
        .Tile_X0Y1_A_O_top(fabric_io_west_in_i[31]),
        .Tile_X0Y1_A_I_top(fabric_io_west_out_o[31]),
        .Tile_X0Y1_A_T_top(fabric_io_west_oeb_o[31]),

        .Tile_X0Y1_B_O_top(fabric_io_west_in_i[30]),
        .Tile_X0Y1_B_I_top(fabric_io_west_out_o[30]),
        .Tile_X0Y1_B_T_top(fabric_io_west_oeb_o[30]),

        .Tile_X0Y1_A_config_C_bit0(fabric_io_west_config_bit0_o[31]),
        .Tile_X0Y1_A_config_C_bit1(fabric_io_west_config_bit1_o[31]),
        .Tile_X0Y1_A_config_C_bit2(fabric_io_west_config_bit2_o[31]),
        .Tile_X0Y1_A_config_C_bit3(fabric_io_west_config_bit3_o[31]),

        .Tile_X0Y1_B_config_C_bit0(fabric_io_west_config_bit0_o[30]),
        .Tile_X0Y1_B_config_C_bit1(fabric_io_west_config_bit1_o[30]),
        .Tile_X0Y1_B_config_C_bit2(fabric_io_west_config_bit2_o[30]),
        .Tile_X0Y1_B_config_C_bit3(fabric_io_west_config_bit3_o[30]),

        .Tile_X0Y2_A_O_top(fabric_io_west_in_i[29]),
        .Tile_X0Y2_A_I_top(fabric_io_west_out_o[29]),
        .Tile_X0Y2_A_T_top(fabric_io_west_oeb_o[29]),

        .Tile_X0Y2_B_O_top(fabric_io_west_in_i[28]),
        .Tile_X0Y2_B_I_top(fabric_io_west_out_o[28]),
        .Tile_X0Y2_B_T_top(fabric_io_west_oeb_o[28]),

        .Tile_X0Y2_A_config_C_bit0(fabric_io_west_config_bit0_o[29]),
        .Tile_X0Y2_A_config_C_bit1(fabric_io_west_config_bit1_o[29]),
        .Tile_X0Y2_A_config_C_bit2(fabric_io_west_config_bit2_o[29]),
        .Tile_X0Y2_A_config_C_bit3(fabric_io_west_config_bit3_o[29]),

        .Tile_X0Y2_B_config_C_bit0(fabric_io_west_config_bit0_o[28]),
        .Tile_X0Y2_B_config_C_bit1(fabric_io_west_config_bit1_o[28]),
        .Tile_X0Y2_B_config_C_bit2(fabric_io_west_config_bit2_o[28]),
        .Tile_X0Y2_B_config_C_bit3(fabric_io_west_config_bit3_o[28]),

        .Tile_X0Y3_A_O_top(fabric_io_west_in_i[27]),
        .Tile_X0Y3_A_I_top(fabric_io_west_out_o[27]),
        .Tile_X0Y3_A_T_top(fabric_io_west_oeb_o[27]),

        .Tile_X0Y3_B_O_top(fabric_io_west_in_i[26]),
        .Tile_X0Y3_B_I_top(fabric_io_west_out_o[26]),
        .Tile_X0Y3_B_T_top(fabric_io_west_oeb_o[26]),

        .Tile_X0Y3_A_config_C_bit0(fabric_io_west_config_bit0_o[27]),
        .Tile_X0Y3_A_config_C_bit1(fabric_io_west_config_bit1_o[27]),
        .Tile_X0Y3_A_config_C_bit2(fabric_io_west_config_bit2_o[27]),
        .Tile_X0Y3_A_config_C_bit3(fabric_io_west_config_bit3_o[27]),

        .Tile_X0Y3_B_config_C_bit0(fabric_io_west_config_bit0_o[26]),
        .Tile_X0Y3_B_config_C_bit1(fabric_io_west_config_bit1_o[26]),
        .Tile_X0Y3_B_config_C_bit2(fabric_io_west_config_bit2_o[26]),
        .Tile_X0Y3_B_config_C_bit3(fabric_io_west_config_bit3_o[26]),

        .Tile_X0Y4_A_O_top(fabric_io_west_in_i[25]),
        .Tile_X0Y4_A_I_top(fabric_io_west_out_o[25]),
        .Tile_X0Y4_A_T_top(fabric_io_west_oeb_o[25]),

        .Tile_X0Y4_B_O_top(fabric_io_west_in_i[24]),
        .Tile_X0Y4_B_I_top(fabric_io_west_out_o[24]),
        .Tile_X0Y4_B_T_top(fabric_io_west_oeb_o[24]),

        .Tile_X0Y4_A_config_C_bit0(fabric_io_west_config_bit0_o[25]),
        .Tile_X0Y4_A_config_C_bit1(fabric_io_west_config_bit1_o[25]),
        .Tile_X0Y4_A_config_C_bit2(fabric_io_west_config_bit2_o[25]),
        .Tile_X0Y4_A_config_C_bit3(fabric_io_west_config_bit3_o[25]),

        .Tile_X0Y4_B_config_C_bit0(fabric_io_west_config_bit0_o[24]),
        .Tile_X0Y4_B_config_C_bit1(fabric_io_west_config_bit1_o[24]),
        .Tile_X0Y4_B_config_C_bit2(fabric_io_west_config_bit2_o[24]),
        .Tile_X0Y4_B_config_C_bit3(fabric_io_west_config_bit3_o[24]),

        .Tile_X0Y5_A_O_top(fabric_io_west_in_i[23]),
        .Tile_X0Y5_A_I_top(fabric_io_west_out_o[23]),
        .Tile_X0Y5_A_T_top(fabric_io_west_oeb_o[23]),

        .Tile_X0Y5_B_O_top(fabric_io_west_in_i[22]),
        .Tile_X0Y5_B_I_top(fabric_io_west_out_o[22]),
        .Tile_X0Y5_B_T_top(fabric_io_west_oeb_o[22]),

        .Tile_X0Y5_A_config_C_bit0(fabric_io_west_config_bit0_o[23]),
        .Tile_X0Y5_A_config_C_bit1(fabric_io_west_config_bit1_o[23]),
        .Tile_X0Y5_A_config_C_bit2(fabric_io_west_config_bit2_o[23]),
        .Tile_X0Y5_A_config_C_bit3(fabric_io_west_config_bit3_o[23]),

        .Tile_X0Y5_B_config_C_bit0(fabric_io_west_config_bit0_o[22]),
        .Tile_X0Y5_B_config_C_bit1(fabric_io_west_config_bit1_o[22]),
        .Tile_X0Y5_B_config_C_bit2(fabric_io_west_config_bit2_o[22]),
        .Tile_X0Y5_B_config_C_bit3(fabric_io_west_config_bit3_o[22]),

        .Tile_X0Y6_A_O_top(fabric_io_west_in_i[21]),
        .Tile_X0Y6_A_I_top(fabric_io_west_out_o[21]),
        .Tile_X0Y6_A_T_top(fabric_io_west_oeb_o[21]),

        .Tile_X0Y6_B_O_top(fabric_io_west_in_i[20]),
        .Tile_X0Y6_B_I_top(fabric_io_west_out_o[20]),
        .Tile_X0Y6_B_T_top(fabric_io_west_oeb_o[20]),

        .Tile_X0Y6_A_config_C_bit0(fabric_io_west_config_bit0_o[21]),
        .Tile_X0Y6_A_config_C_bit1(fabric_io_west_config_bit1_o[21]),
        .Tile_X0Y6_A_config_C_bit2(fabric_io_west_config_bit2_o[21]),
        .Tile_X0Y6_A_config_C_bit3(fabric_io_west_config_bit3_o[21]),

        .Tile_X0Y6_B_config_C_bit0(fabric_io_west_config_bit0_o[20]),
        .Tile_X0Y6_B_config_C_bit1(fabric_io_west_config_bit1_o[20]),
        .Tile_X0Y6_B_config_C_bit2(fabric_io_west_config_bit2_o[20]),
        .Tile_X0Y6_B_config_C_bit3(fabric_io_west_config_bit3_o[20]),

        .Tile_X0Y7_A_O_top(fabric_io_west_in_i[19]),
        .Tile_X0Y7_A_I_top(fabric_io_west_out_o[19]),
        .Tile_X0Y7_A_T_top(fabric_io_west_oeb_o[19]),

        .Tile_X0Y7_B_O_top(fabric_io_west_in_i[18]),
        .Tile_X0Y7_B_I_top(fabric_io_west_out_o[18]),
        .Tile_X0Y7_B_T_top(fabric_io_west_oeb_o[18]),

        .Tile_X0Y7_A_config_C_bit0(fabric_io_west_config_bit0_o[19]),
        .Tile_X0Y7_A_config_C_bit1(fabric_io_west_config_bit1_o[19]),
        .Tile_X0Y7_A_config_C_bit2(fabric_io_west_config_bit2_o[19]),
        .Tile_X0Y7_A_config_C_bit3(fabric_io_west_config_bit3_o[19]),

        .Tile_X0Y7_B_config_C_bit0(fabric_io_west_config_bit0_o[18]),
        .Tile_X0Y7_B_config_C_bit1(fabric_io_west_config_bit1_o[18]),
        .Tile_X0Y7_B_config_C_bit2(fabric_io_west_config_bit2_o[18]),
        .Tile_X0Y7_B_config_C_bit3(fabric_io_west_config_bit3_o[18]),

        .Tile_X0Y8_A_O_top(fabric_io_west_in_i[17]),
        .Tile_X0Y8_A_I_top(fabric_io_west_out_o[17]),
        .Tile_X0Y8_A_T_top(fabric_io_west_oeb_o[17]),

        .Tile_X0Y8_B_O_top(fabric_io_west_in_i[16]),
        .Tile_X0Y8_B_I_top(fabric_io_west_out_o[16]),
        .Tile_X0Y8_B_T_top(fabric_io_west_oeb_o[16]),

        .Tile_X0Y8_A_config_C_bit0(fabric_io_west_config_bit0_o[17]),
        .Tile_X0Y8_A_config_C_bit1(fabric_io_west_config_bit1_o[17]),
        .Tile_X0Y8_A_config_C_bit2(fabric_io_west_config_bit2_o[17]),
        .Tile_X0Y8_A_config_C_bit3(fabric_io_west_config_bit3_o[17]),

        .Tile_X0Y8_B_config_C_bit0(fabric_io_west_config_bit0_o[16]),
        .Tile_X0Y8_B_config_C_bit1(fabric_io_west_config_bit1_o[16]),
        .Tile_X0Y8_B_config_C_bit2(fabric_io_west_config_bit2_o[16]),
        .Tile_X0Y8_B_config_C_bit3(fabric_io_west_config_bit3_o[16]),

        .Tile_X0Y9_A_O_top(fabric_io_west_in_i[15]),
        .Tile_X0Y9_A_I_top(fabric_io_west_out_o[15]),
        .Tile_X0Y9_A_T_top(fabric_io_west_oeb_o[15]),

        .Tile_X0Y9_B_O_top(fabric_io_west_in_i[14]),
        .Tile_X0Y9_B_I_top(fabric_io_west_out_o[14]),
        .Tile_X0Y9_B_T_top(fabric_io_west_oeb_o[14]),

        .Tile_X0Y9_A_config_C_bit0(fabric_io_west_config_bit0_o[15]),
        .Tile_X0Y9_A_config_C_bit1(fabric_io_west_config_bit1_o[15]),
        .Tile_X0Y9_A_config_C_bit2(fabric_io_west_config_bit2_o[15]),
        .Tile_X0Y9_A_config_C_bit3(fabric_io_west_config_bit3_o[15]),

        .Tile_X0Y9_B_config_C_bit0(fabric_io_west_config_bit0_o[14]),
        .Tile_X0Y9_B_config_C_bit1(fabric_io_west_config_bit1_o[14]),
        .Tile_X0Y9_B_config_C_bit2(fabric_io_west_config_bit2_o[14]),
        .Tile_X0Y9_B_config_C_bit3(fabric_io_west_config_bit3_o[14]),

        .Tile_X0Y10_A_O_top(fabric_io_west_in_i[13]),
        .Tile_X0Y10_A_I_top(fabric_io_west_out_o[13]),
        .Tile_X0Y10_A_T_top(fabric_io_west_oeb_o[13]),

        .Tile_X0Y10_B_O_top(fabric_io_west_in_i[12]),
        .Tile_X0Y10_B_I_top(fabric_io_west_out_o[12]),
        .Tile_X0Y10_B_T_top(fabric_io_west_oeb_o[12]),

        .Tile_X0Y10_A_config_C_bit0(fabric_io_west_config_bit0_o[13]),
        .Tile_X0Y10_A_config_C_bit1(fabric_io_west_config_bit1_o[13]),
        .Tile_X0Y10_A_config_C_bit2(fabric_io_west_config_bit2_o[13]),
        .Tile_X0Y10_A_config_C_bit3(fabric_io_west_config_bit3_o[13]),

        .Tile_X0Y10_B_config_C_bit0(fabric_io_west_config_bit0_o[12]),
        .Tile_X0Y10_B_config_C_bit1(fabric_io_west_config_bit1_o[12]),
        .Tile_X0Y10_B_config_C_bit2(fabric_io_west_config_bit2_o[12]),
        .Tile_X0Y10_B_config_C_bit3(fabric_io_west_config_bit3_o[12]),

        .Tile_X0Y11_A_O_top(fabric_io_west_in_i[11]),
        .Tile_X0Y11_A_I_top(fabric_io_west_out_o[11]),
        .Tile_X0Y11_A_T_top(fabric_io_west_oeb_o[11]),

        .Tile_X0Y11_B_O_top(fabric_io_west_in_i[10]),
        .Tile_X0Y11_B_I_top(fabric_io_west_out_o[10]),
        .Tile_X0Y11_B_T_top(fabric_io_west_oeb_o[10]),

        .Tile_X0Y11_A_config_C_bit0(fabric_io_west_config_bit0_o[11]),
        .Tile_X0Y11_A_config_C_bit1(fabric_io_west_config_bit1_o[11]),
        .Tile_X0Y11_A_config_C_bit2(fabric_io_west_config_bit2_o[11]),
        .Tile_X0Y11_A_config_C_bit3(fabric_io_west_config_bit3_o[11]),

        .Tile_X0Y11_B_config_C_bit0(fabric_io_west_config_bit0_o[10]),
        .Tile_X0Y11_B_config_C_bit1(fabric_io_west_config_bit1_o[10]),
        .Tile_X0Y11_B_config_C_bit2(fabric_io_west_config_bit2_o[10]),
        .Tile_X0Y11_B_config_C_bit3(fabric_io_west_config_bit3_o[10]),

        .Tile_X0Y12_A_O_top(fabric_io_west_in_i[9]),
        .Tile_X0Y12_A_I_top(fabric_io_west_out_o[9]),
        .Tile_X0Y12_A_T_top(fabric_io_west_oeb_o[9]),

        .Tile_X0Y12_B_O_top(fabric_io_west_in_i[8]),
        .Tile_X0Y12_B_I_top(fabric_io_west_out_o[8]),
        .Tile_X0Y12_B_T_top(fabric_io_west_oeb_o[8]),

        .Tile_X0Y12_A_config_C_bit0(fabric_io_west_config_bit0_o[9]),
        .Tile_X0Y12_A_config_C_bit1(fabric_io_west_config_bit1_o[9]),
        .Tile_X0Y12_A_config_C_bit2(fabric_io_west_config_bit2_o[9]),
        .Tile_X0Y12_A_config_C_bit3(fabric_io_west_config_bit3_o[9]),

        .Tile_X0Y12_B_config_C_bit0(fabric_io_west_config_bit0_o[8]),
        .Tile_X0Y12_B_config_C_bit1(fabric_io_west_config_bit1_o[8]),
        .Tile_X0Y12_B_config_C_bit2(fabric_io_west_config_bit2_o[8]),
        .Tile_X0Y12_B_config_C_bit3(fabric_io_west_config_bit3_o[8]),

        .Tile_X0Y13_A_O_top(fabric_io_west_in_i[7]),
        .Tile_X0Y13_A_I_top(fabric_io_west_out_o[7]),
        .Tile_X0Y13_A_T_top(fabric_io_west_oeb_o[7]),

        .Tile_X0Y13_B_O_top(fabric_io_west_in_i[6]),
        .Tile_X0Y13_B_I_top(fabric_io_west_out_o[6]),
        .Tile_X0Y13_B_T_top(fabric_io_west_oeb_o[6]),

        .Tile_X0Y13_A_config_C_bit0(fabric_io_west_config_bit0_o[7]),
        .Tile_X0Y13_A_config_C_bit1(fabric_io_west_config_bit1_o[7]),
        .Tile_X0Y13_A_config_C_bit2(fabric_io_west_config_bit2_o[7]),
        .Tile_X0Y13_A_config_C_bit3(fabric_io_west_config_bit3_o[7]),

        .Tile_X0Y13_B_config_C_bit0(fabric_io_west_config_bit0_o[6]),
        .Tile_X0Y13_B_config_C_bit1(fabric_io_west_config_bit1_o[6]),
        .Tile_X0Y13_B_config_C_bit2(fabric_io_west_config_bit2_o[6]),
        .Tile_X0Y13_B_config_C_bit3(fabric_io_west_config_bit3_o[6]),

        .Tile_X0Y14_A_O_top(fabric_io_west_in_i[5]),
        .Tile_X0Y14_A_I_top(fabric_io_west_out_o[5]),
        .Tile_X0Y14_A_T_top(fabric_io_west_oeb_o[5]),

        .Tile_X0Y14_B_O_top(fabric_io_west_in_i[4]),
        .Tile_X0Y14_B_I_top(fabric_io_west_out_o[4]),
        .Tile_X0Y14_B_T_top(fabric_io_west_oeb_o[4]),

        .Tile_X0Y14_A_config_C_bit0(fabric_io_west_config_bit0_o[5]),
        .Tile_X0Y14_A_config_C_bit1(fabric_io_west_config_bit1_o[5]),
        .Tile_X0Y14_A_config_C_bit2(fabric_io_west_config_bit2_o[5]),
        .Tile_X0Y14_A_config_C_bit3(fabric_io_west_config_bit3_o[5]),

        .Tile_X0Y14_B_config_C_bit0(fabric_io_west_config_bit0_o[4]),
        .Tile_X0Y14_B_config_C_bit1(fabric_io_west_config_bit1_o[4]),
        .Tile_X0Y14_B_config_C_bit2(fabric_io_west_config_bit2_o[4]),
        .Tile_X0Y14_B_config_C_bit3(fabric_io_west_config_bit3_o[4]),

        .Tile_X0Y15_A_O_top(fabric_io_west_in_i[3]),
        .Tile_X0Y15_A_I_top(fabric_io_west_out_o[3]),
        .Tile_X0Y15_A_T_top(fabric_io_west_oeb_o[3]),

        .Tile_X0Y15_B_O_top(fabric_io_west_in_i[2]),
        .Tile_X0Y15_B_I_top(fabric_io_west_out_o[2]),
        .Tile_X0Y15_B_T_top(fabric_io_west_oeb_o[2]),

        .Tile_X0Y15_A_config_C_bit0(fabric_io_west_config_bit0_o[3]),
        .Tile_X0Y15_A_config_C_bit1(fabric_io_west_config_bit1_o[3]),
        .Tile_X0Y15_A_config_C_bit2(fabric_io_west_config_bit2_o[3]),
        .Tile_X0Y15_A_config_C_bit3(fabric_io_west_config_bit3_o[3]),

        .Tile_X0Y15_B_config_C_bit0(fabric_io_west_config_bit0_o[2]),
        .Tile_X0Y15_B_config_C_bit1(fabric_io_west_config_bit1_o[2]),
        .Tile_X0Y15_B_config_C_bit2(fabric_io_west_config_bit2_o[2]),
        .Tile_X0Y15_B_config_C_bit3(fabric_io_west_config_bit3_o[2]),

        .Tile_X0Y16_A_O_top(fabric_io_west_in_i[1]),
        .Tile_X0Y16_A_I_top(fabric_io_west_out_o[1]),
        .Tile_X0Y16_A_T_top(fabric_io_west_oeb_o[1]),

        .Tile_X0Y16_B_O_top(fabric_io_west_in_i[0]),
        .Tile_X0Y16_B_I_top(fabric_io_west_out_o[0]),
        .Tile_X0Y16_B_T_top(fabric_io_west_oeb_o[0]),

        .Tile_X0Y16_A_config_C_bit0(fabric_io_west_config_bit0_o[1]),
        .Tile_X0Y16_A_config_C_bit1(fabric_io_west_config_bit1_o[1]),
        .Tile_X0Y16_A_config_C_bit2(fabric_io_west_config_bit2_o[1]),
        .Tile_X0Y16_A_config_C_bit3(fabric_io_west_config_bit3_o[1]),

        .Tile_X0Y16_B_config_C_bit0(fabric_io_west_config_bit0_o[0]),
        .Tile_X0Y16_B_config_C_bit1(fabric_io_west_config_bit1_o[0]),
        .Tile_X0Y16_B_config_C_bit2(fabric_io_west_config_bit2_o[0]),
        .Tile_X0Y16_B_config_C_bit3(fabric_io_west_config_bit3_o[0]),

        // North I/Os
        .Tile_X1Y0_A_O_top(fabric_io_north_in_i[1]),
        .Tile_X1Y0_A_I_top(fabric_io_north_out_o[1]),
        .Tile_X1Y0_A_T_top(fabric_io_north_oeb_o[1]),

        .Tile_X1Y0_B_O_top(fabric_io_north_in_i[0]),
        .Tile_X1Y0_B_I_top(fabric_io_north_out_o[0]),
        .Tile_X1Y0_B_T_top(fabric_io_north_oeb_o[0]),

        .Tile_X1Y0_A_config_C_bit0(fabric_io_north_config_bit0_o[1]),
        .Tile_X1Y0_A_config_C_bit1(fabric_io_north_config_bit1_o[1]),
        .Tile_X1Y0_A_config_C_bit2(fabric_io_north_config_bit2_o[1]),
        .Tile_X1Y0_A_config_C_bit3(fabric_io_north_config_bit3_o[1]),

        .Tile_X1Y0_B_config_C_bit0(fabric_io_north_config_bit0_o[0]),
        .Tile_X1Y0_B_config_C_bit1(fabric_io_north_config_bit1_o[0]),
        .Tile_X1Y0_B_config_C_bit2(fabric_io_north_config_bit2_o[0]),
        .Tile_X1Y0_B_config_C_bit3(fabric_io_north_config_bit3_o[0]),

        .Tile_X2Y0_A_O_top(fabric_io_north_in_i[3]),
        .Tile_X2Y0_A_I_top(fabric_io_north_out_o[3]),
        .Tile_X2Y0_A_T_top(fabric_io_north_oeb_o[3]),

        .Tile_X2Y0_B_O_top(fabric_io_north_in_i[2]),
        .Tile_X2Y0_B_I_top(fabric_io_north_out_o[2]),
        .Tile_X2Y0_B_T_top(fabric_io_north_oeb_o[2]),

        .Tile_X2Y0_A_config_C_bit0(fabric_io_north_config_bit0_o[3]),
        .Tile_X2Y0_A_config_C_bit1(fabric_io_north_config_bit1_o[3]),
        .Tile_X2Y0_A_config_C_bit2(fabric_io_north_config_bit2_o[3]),
        .Tile_X2Y0_A_config_C_bit3(fabric_io_north_config_bit3_o[3]),

        .Tile_X2Y0_B_config_C_bit0(fabric_io_north_config_bit0_o[2]),
        .Tile_X2Y0_B_config_C_bit1(fabric_io_north_config_bit1_o[2]),
        .Tile_X2Y0_B_config_C_bit2(fabric_io_north_config_bit2_o[2]),
        .Tile_X2Y0_B_config_C_bit3(fabric_io_north_config_bit3_o[2]),

        .Tile_X4Y0_A_O_top(fabric_io_north_in_i[5]),
        .Tile_X4Y0_A_I_top(fabric_io_north_out_o[5]),
        .Tile_X4Y0_A_T_top(fabric_io_north_oeb_o[5]),

        .Tile_X4Y0_B_O_top(fabric_io_north_in_i[4]),
        .Tile_X4Y0_B_I_top(fabric_io_north_out_o[4]),
        .Tile_X4Y0_B_T_top(fabric_io_north_oeb_o[4]),

        .Tile_X4Y0_A_config_C_bit0(fabric_io_north_config_bit0_o[5]),
        .Tile_X4Y0_A_config_C_bit1(fabric_io_north_config_bit1_o[5]),
        .Tile_X4Y0_A_config_C_bit2(fabric_io_north_config_bit2_o[5]),
        .Tile_X4Y0_A_config_C_bit3(fabric_io_north_config_bit3_o[5]),

        .Tile_X4Y0_B_config_C_bit0(fabric_io_north_config_bit0_o[4]),
        .Tile_X4Y0_B_config_C_bit1(fabric_io_north_config_bit1_o[4]),
        .Tile_X4Y0_B_config_C_bit2(fabric_io_north_config_bit2_o[4]),
        .Tile_X4Y0_B_config_C_bit3(fabric_io_north_config_bit3_o[4]),

        .Tile_X5Y0_A_O_top(fabric_io_north_in_i[7]),
        .Tile_X5Y0_A_I_top(fabric_io_north_out_o[7]),
        .Tile_X5Y0_A_T_top(fabric_io_north_oeb_o[7]),

        .Tile_X5Y0_B_O_top(fabric_io_north_in_i[6]),
        .Tile_X5Y0_B_I_top(fabric_io_north_out_o[6]),
        .Tile_X5Y0_B_T_top(fabric_io_north_oeb_o[6]),

        .Tile_X5Y0_A_config_C_bit0(fabric_io_north_config_bit0_o[7]),
        .Tile_X5Y0_A_config_C_bit1(fabric_io_north_config_bit1_o[7]),
        .Tile_X5Y0_A_config_C_bit2(fabric_io_north_config_bit2_o[7]),
        .Tile_X5Y0_A_config_C_bit3(fabric_io_north_config_bit3_o[7]),

        .Tile_X5Y0_B_config_C_bit0(fabric_io_north_config_bit0_o[6]),
        .Tile_X5Y0_B_config_C_bit1(fabric_io_north_config_bit1_o[6]),
        .Tile_X5Y0_B_config_C_bit2(fabric_io_north_config_bit2_o[6]),
        .Tile_X5Y0_B_config_C_bit3(fabric_io_north_config_bit3_o[6]),

        .Tile_X6Y0_A_O_top(fabric_io_north_in_i[9]),
        .Tile_X6Y0_A_I_top(fabric_io_north_out_o[9]),
        .Tile_X6Y0_A_T_top(fabric_io_north_oeb_o[9]),

        .Tile_X6Y0_B_O_top(fabric_io_north_in_i[8]),
        .Tile_X6Y0_B_I_top(fabric_io_north_out_o[8]),
        .Tile_X6Y0_B_T_top(fabric_io_north_oeb_o[8]),

        .Tile_X6Y0_A_config_C_bit0(fabric_io_north_config_bit0_o[9]),
        .Tile_X6Y0_A_config_C_bit1(fabric_io_north_config_bit1_o[9]),
        .Tile_X6Y0_A_config_C_bit2(fabric_io_north_config_bit2_o[9]),
        .Tile_X6Y0_A_config_C_bit3(fabric_io_north_config_bit3_o[9]),

        .Tile_X6Y0_B_config_C_bit0(fabric_io_north_config_bit0_o[8]),
        .Tile_X6Y0_B_config_C_bit1(fabric_io_north_config_bit1_o[8]),
        .Tile_X6Y0_B_config_C_bit2(fabric_io_north_config_bit2_o[8]),
        .Tile_X6Y0_B_config_C_bit3(fabric_io_north_config_bit3_o[8]),

        .Tile_X8Y0_A_O_top(fabric_io_north_in_i[11]),
        .Tile_X8Y0_A_I_top(fabric_io_north_out_o[11]),
        .Tile_X8Y0_A_T_top(fabric_io_north_oeb_o[11]),

        .Tile_X8Y0_B_O_top(fabric_io_north_in_i[10]),
        .Tile_X8Y0_B_I_top(fabric_io_north_out_o[10]),
        .Tile_X8Y0_B_T_top(fabric_io_north_oeb_o[10]),

        .Tile_X8Y0_A_config_C_bit0(fabric_io_north_config_bit0_o[11]),
        .Tile_X8Y0_A_config_C_bit1(fabric_io_north_config_bit1_o[11]),
        .Tile_X8Y0_A_config_C_bit2(fabric_io_north_config_bit2_o[11]),
        .Tile_X8Y0_A_config_C_bit3(fabric_io_north_config_bit3_o[11]),

        .Tile_X8Y0_B_config_C_bit0(fabric_io_north_config_bit0_o[10]),
        .Tile_X8Y0_B_config_C_bit1(fabric_io_north_config_bit1_o[10]),
        .Tile_X8Y0_B_config_C_bit2(fabric_io_north_config_bit2_o[10]),
        .Tile_X8Y0_B_config_C_bit3(fabric_io_north_config_bit3_o[10]),

        .Tile_X9Y0_A_O_top(fabric_io_north_in_i[13]),
        .Tile_X9Y0_A_I_top(fabric_io_north_out_o[13]),
        .Tile_X9Y0_A_T_top(fabric_io_north_oeb_o[13]),

        .Tile_X9Y0_B_O_top(fabric_io_north_in_i[12]),
        .Tile_X9Y0_B_I_top(fabric_io_north_out_o[12]),
        .Tile_X9Y0_B_T_top(fabric_io_north_oeb_o[12]),

        .Tile_X9Y0_A_config_C_bit0(fabric_io_north_config_bit0_o[13]),
        .Tile_X9Y0_A_config_C_bit1(fabric_io_north_config_bit1_o[13]),
        .Tile_X9Y0_A_config_C_bit2(fabric_io_north_config_bit2_o[13]),
        .Tile_X9Y0_A_config_C_bit3(fabric_io_north_config_bit3_o[13]),

        .Tile_X9Y0_B_config_C_bit0(fabric_io_north_config_bit0_o[12]),
        .Tile_X9Y0_B_config_C_bit1(fabric_io_north_config_bit1_o[12]),
        .Tile_X9Y0_B_config_C_bit2(fabric_io_north_config_bit2_o[12]),
        .Tile_X9Y0_B_config_C_bit3(fabric_io_north_config_bit3_o[12]),

        .Tile_X10Y0_A_O_top(fabric_io_north_in_i[15]),
        .Tile_X10Y0_A_I_top(fabric_io_north_out_o[15]),
        .Tile_X10Y0_A_T_top(fabric_io_north_oeb_o[15]),

        .Tile_X10Y0_B_O_top(fabric_io_north_in_i[14]),
        .Tile_X10Y0_B_I_top(fabric_io_north_out_o[14]),
        .Tile_X10Y0_B_T_top(fabric_io_north_oeb_o[14]),

        .Tile_X10Y0_A_config_C_bit0(fabric_io_north_config_bit0_o[15]),
        .Tile_X10Y0_A_config_C_bit1(fabric_io_north_config_bit1_o[15]),
        .Tile_X10Y0_A_config_C_bit2(fabric_io_north_config_bit2_o[15]),
        .Tile_X10Y0_A_config_C_bit3(fabric_io_north_config_bit3_o[15]),

        .Tile_X10Y0_B_config_C_bit0(fabric_io_north_config_bit0_o[14]),
        .Tile_X10Y0_B_config_C_bit1(fabric_io_north_config_bit1_o[14]),
        .Tile_X10Y0_B_config_C_bit2(fabric_io_north_config_bit2_o[14]),
        .Tile_X10Y0_B_config_C_bit3(fabric_io_north_config_bit3_o[14]),

        // ADC
        .Tile_X9Y17_CMP_top(fabric_adc0_cmp_i),
        .Tile_X9Y17_HOLD_top(fabric_adc0_hold_o),
        .Tile_X9Y17_RESET_top(fabric_adc0_reset_o),
        .Tile_X9Y17_VALUE_top0(fabric_adc0_value_o[0]),
        .Tile_X9Y17_VALUE_top1(fabric_adc0_value_o[1]),
        .Tile_X9Y17_VALUE_top2(fabric_adc0_value_o[2]),
        .Tile_X9Y17_VALUE_top3(fabric_adc0_value_o[3]),
        .Tile_X9Y17_VALUE_top4(fabric_adc0_value_o[4]),
        .Tile_X9Y17_VALUE_top5(fabric_adc0_value_o[5]),
        .Tile_X9Y17_VALUE_top6(fabric_adc0_value_o[6]),
        .Tile_X9Y17_VALUE_top7(fabric_adc0_value_o[7]),
        .Tile_X9Y17_VALUE_top8(fabric_adc0_value_o[8]),
        .Tile_X9Y17_VALUE_top9(fabric_adc0_value_o[9]),
        .Tile_X9Y17_VALUE_top10(fabric_adc0_value_o[10]),
        .Tile_X9Y17_VALUE_top11(fabric_adc0_value_o[11]),

        // DAC
        .Tile_X10Y17_VALUE_top0(fabric_dac0_value_o[0]),
        .Tile_X10Y17_VALUE_top1(fabric_dac0_value_o[1]),
        .Tile_X10Y17_VALUE_top2(fabric_dac0_value_o[2]),
        .Tile_X10Y17_VALUE_top3(fabric_dac0_value_o[3]),
        .Tile_X10Y17_VALUE_top4(fabric_dac0_value_o[4]),
        .Tile_X10Y17_VALUE_top5(fabric_dac0_value_o[5]),
        .Tile_X10Y17_VALUE_top6(fabric_dac0_value_o[6]),
        .Tile_X10Y17_VALUE_top7(fabric_dac0_value_o[7]),

        // SRAM 0
        .Tile_X11Y2_DO_SRAM0(fabric_sram0_do_i[0]),
        .Tile_X11Y2_DO_SRAM1(fabric_sram0_do_i[1]),
        .Tile_X11Y2_DO_SRAM2(fabric_sram0_do_i[2]),
        .Tile_X11Y2_DO_SRAM3(fabric_sram0_do_i[3]),
        .Tile_X11Y2_DO_SRAM4(fabric_sram0_do_i[4]),
        .Tile_X11Y2_DO_SRAM5(fabric_sram0_do_i[5]),
        .Tile_X11Y2_DO_SRAM6(fabric_sram0_do_i[6]),
        .Tile_X11Y2_DO_SRAM7(fabric_sram0_do_i[7]),
        .Tile_X11Y2_DO_SRAM8(fabric_sram0_do_i[8]),
        .Tile_X11Y2_DO_SRAM9(fabric_sram0_do_i[9]),
        .Tile_X11Y2_DO_SRAM10(fabric_sram0_do_i[10]),
        .Tile_X11Y2_DO_SRAM11(fabric_sram0_do_i[11]),
        .Tile_X11Y2_DO_SRAM12(fabric_sram0_do_i[12]),
        .Tile_X11Y2_DO_SRAM13(fabric_sram0_do_i[13]),
        .Tile_X11Y2_DO_SRAM14(fabric_sram0_do_i[14]),
        .Tile_X11Y2_DO_SRAM15(fabric_sram0_do_i[15]),
        .Tile_X11Y2_DO_SRAM16(fabric_sram0_do_i[16]),
        .Tile_X11Y2_DO_SRAM17(fabric_sram0_do_i[17]),
        .Tile_X11Y2_DO_SRAM18(fabric_sram0_do_i[18]),
        .Tile_X11Y2_DO_SRAM19(fabric_sram0_do_i[19]),
        .Tile_X11Y2_DO_SRAM20(fabric_sram0_do_i[20]),
        .Tile_X11Y2_DO_SRAM21(fabric_sram0_do_i[21]),
        .Tile_X11Y2_DO_SRAM22(fabric_sram0_do_i[22]),
        .Tile_X11Y2_DO_SRAM23(fabric_sram0_do_i[23]),
        .Tile_X11Y2_DO_SRAM24(fabric_sram0_do_i[24]),
        .Tile_X11Y2_DO_SRAM25(fabric_sram0_do_i[25]),
        .Tile_X11Y2_DO_SRAM26(fabric_sram0_do_i[26]),
        .Tile_X11Y2_DO_SRAM27(fabric_sram0_do_i[27]),
        .Tile_X11Y2_DO_SRAM28(fabric_sram0_do_i[28]),
        .Tile_X11Y2_DO_SRAM29(fabric_sram0_do_i[29]),
        .Tile_X11Y2_DO_SRAM30(fabric_sram0_do_i[30]),
        .Tile_X11Y2_DO_SRAM31(fabric_sram0_do_i[31]),
        .Tile_X11Y2_AD_SRAM0(fabric_sram0_ad_o[0]),
        .Tile_X11Y2_AD_SRAM1(fabric_sram0_ad_o[1]),
        .Tile_X11Y2_AD_SRAM2(fabric_sram0_ad_o[2]),
        .Tile_X11Y2_AD_SRAM3(fabric_sram0_ad_o[3]),
        .Tile_X11Y2_AD_SRAM4(fabric_sram0_ad_o[4]),
        .Tile_X11Y2_AD_SRAM5(fabric_sram0_ad_o[5]),
        .Tile_X11Y2_AD_SRAM6(fabric_sram0_ad_o[6]),
        .Tile_X11Y2_AD_SRAM7(fabric_sram0_ad_o[7]),
        .Tile_X11Y2_AD_SRAM8(fabric_sram0_ad_o[8]),
        .Tile_X11Y2_AD_SRAM9(fabric_sram0_ad_o[9]),
        .Tile_X11Y2_BEN_SRAM0(fabric_sram0_ben_o[0]),
        .Tile_X11Y2_BEN_SRAM1(fabric_sram0_ben_o[1]),
        .Tile_X11Y2_BEN_SRAM2(fabric_sram0_ben_o[2]),
        .Tile_X11Y2_BEN_SRAM3(fabric_sram0_ben_o[3]),
        .Tile_X11Y2_BEN_SRAM4(fabric_sram0_ben_o[4]),
        .Tile_X11Y2_BEN_SRAM5(fabric_sram0_ben_o[5]),
        .Tile_X11Y2_BEN_SRAM6(fabric_sram0_ben_o[6]),
        .Tile_X11Y2_BEN_SRAM7(fabric_sram0_ben_o[7]),
        .Tile_X11Y2_BEN_SRAM8(fabric_sram0_ben_o[8]),
        .Tile_X11Y2_BEN_SRAM9(fabric_sram0_ben_o[9]),
        .Tile_X11Y2_BEN_SRAM10(fabric_sram0_ben_o[10]),
        .Tile_X11Y2_BEN_SRAM11(fabric_sram0_ben_o[11]),
        .Tile_X11Y2_BEN_SRAM12(fabric_sram0_ben_o[12]),
        .Tile_X11Y2_BEN_SRAM13(fabric_sram0_ben_o[13]),
        .Tile_X11Y2_BEN_SRAM14(fabric_sram0_ben_o[14]),
        .Tile_X11Y2_BEN_SRAM15(fabric_sram0_ben_o[15]),
        .Tile_X11Y2_BEN_SRAM16(fabric_sram0_ben_o[16]),
        .Tile_X11Y2_BEN_SRAM17(fabric_sram0_ben_o[17]),
        .Tile_X11Y2_BEN_SRAM18(fabric_sram0_ben_o[18]),
        .Tile_X11Y2_BEN_SRAM19(fabric_sram0_ben_o[19]),
        .Tile_X11Y2_BEN_SRAM20(fabric_sram0_ben_o[20]),
        .Tile_X11Y2_BEN_SRAM21(fabric_sram0_ben_o[21]),
        .Tile_X11Y2_BEN_SRAM22(fabric_sram0_ben_o[22]),
        .Tile_X11Y2_BEN_SRAM23(fabric_sram0_ben_o[23]),
        .Tile_X11Y2_BEN_SRAM24(fabric_sram0_ben_o[24]),
        .Tile_X11Y2_BEN_SRAM25(fabric_sram0_ben_o[25]),
        .Tile_X11Y2_BEN_SRAM26(fabric_sram0_ben_o[26]),
        .Tile_X11Y2_BEN_SRAM27(fabric_sram0_ben_o[27]),
        .Tile_X11Y2_BEN_SRAM28(fabric_sram0_ben_o[28]),
        .Tile_X11Y2_BEN_SRAM29(fabric_sram0_ben_o[29]),
        .Tile_X11Y2_BEN_SRAM30(fabric_sram0_ben_o[30]),
        .Tile_X11Y2_BEN_SRAM31(fabric_sram0_ben_o[31]),
        .Tile_X11Y2_DI_SRAM0(fabric_sram0_di_o[0]),
        .Tile_X11Y2_DI_SRAM1(fabric_sram0_di_o[1]),
        .Tile_X11Y2_DI_SRAM2(fabric_sram0_di_o[2]),
        .Tile_X11Y2_DI_SRAM3(fabric_sram0_di_o[3]),
        .Tile_X11Y2_DI_SRAM4(fabric_sram0_di_o[4]),
        .Tile_X11Y2_DI_SRAM5(fabric_sram0_di_o[5]),
        .Tile_X11Y2_DI_SRAM6(fabric_sram0_di_o[6]),
        .Tile_X11Y2_DI_SRAM7(fabric_sram0_di_o[7]),
        .Tile_X11Y2_DI_SRAM8(fabric_sram0_di_o[8]),
        .Tile_X11Y2_DI_SRAM9(fabric_sram0_di_o[9]),
        .Tile_X11Y2_DI_SRAM10(fabric_sram0_di_o[10]),
        .Tile_X11Y2_DI_SRAM11(fabric_sram0_di_o[11]),
        .Tile_X11Y2_DI_SRAM12(fabric_sram0_di_o[12]),
        .Tile_X11Y2_DI_SRAM13(fabric_sram0_di_o[13]),
        .Tile_X11Y2_DI_SRAM14(fabric_sram0_di_o[14]),
        .Tile_X11Y2_DI_SRAM15(fabric_sram0_di_o[15]),
        .Tile_X11Y2_DI_SRAM16(fabric_sram0_di_o[16]),
        .Tile_X11Y2_DI_SRAM17(fabric_sram0_di_o[17]),
        .Tile_X11Y2_DI_SRAM18(fabric_sram0_di_o[18]),
        .Tile_X11Y2_DI_SRAM19(fabric_sram0_di_o[19]),
        .Tile_X11Y2_DI_SRAM20(fabric_sram0_di_o[20]),
        .Tile_X11Y2_DI_SRAM21(fabric_sram0_di_o[21]),
        .Tile_X11Y2_DI_SRAM22(fabric_sram0_di_o[22]),
        .Tile_X11Y2_DI_SRAM23(fabric_sram0_di_o[23]),
        .Tile_X11Y2_DI_SRAM24(fabric_sram0_di_o[24]),
        .Tile_X11Y2_DI_SRAM25(fabric_sram0_di_o[25]),
        .Tile_X11Y2_DI_SRAM26(fabric_sram0_di_o[26]),
        .Tile_X11Y2_DI_SRAM27(fabric_sram0_di_o[27]),
        .Tile_X11Y2_DI_SRAM28(fabric_sram0_di_o[28]),
        .Tile_X11Y2_DI_SRAM29(fabric_sram0_di_o[29]),
        .Tile_X11Y2_DI_SRAM30(fabric_sram0_di_o[30]),
        .Tile_X11Y2_DI_SRAM31(fabric_sram0_di_o[31]),
        .Tile_X11Y2_EN_SRAM(fabric_sram0_en),
        .Tile_X11Y2_R_WB_SRAM(fabric_sram0_rw_no),
        .Tile_X11Y2_CLOCK_SRAM(fabric_sram0_clk_o),

        // SRAM 1
        .Tile_X11Y4_DO_SRAM0(fabric_sram1_do_i[0]),
        .Tile_X11Y4_DO_SRAM1(fabric_sram1_do_i[1]),
        .Tile_X11Y4_DO_SRAM2(fabric_sram1_do_i[2]),
        .Tile_X11Y4_DO_SRAM3(fabric_sram1_do_i[3]),
        .Tile_X11Y4_DO_SRAM4(fabric_sram1_do_i[4]),
        .Tile_X11Y4_DO_SRAM5(fabric_sram1_do_i[5]),
        .Tile_X11Y4_DO_SRAM6(fabric_sram1_do_i[6]),
        .Tile_X11Y4_DO_SRAM7(fabric_sram1_do_i[7]),
        .Tile_X11Y4_DO_SRAM8(fabric_sram1_do_i[8]),
        .Tile_X11Y4_DO_SRAM9(fabric_sram1_do_i[9]),
        .Tile_X11Y4_DO_SRAM10(fabric_sram1_do_i[10]),
        .Tile_X11Y4_DO_SRAM11(fabric_sram1_do_i[11]),
        .Tile_X11Y4_DO_SRAM12(fabric_sram1_do_i[12]),
        .Tile_X11Y4_DO_SRAM13(fabric_sram1_do_i[13]),
        .Tile_X11Y4_DO_SRAM14(fabric_sram1_do_i[14]),
        .Tile_X11Y4_DO_SRAM15(fabric_sram1_do_i[15]),
        .Tile_X11Y4_DO_SRAM16(fabric_sram1_do_i[16]),
        .Tile_X11Y4_DO_SRAM17(fabric_sram1_do_i[17]),
        .Tile_X11Y4_DO_SRAM18(fabric_sram1_do_i[18]),
        .Tile_X11Y4_DO_SRAM19(fabric_sram1_do_i[19]),
        .Tile_X11Y4_DO_SRAM20(fabric_sram1_do_i[20]),
        .Tile_X11Y4_DO_SRAM21(fabric_sram1_do_i[21]),
        .Tile_X11Y4_DO_SRAM22(fabric_sram1_do_i[22]),
        .Tile_X11Y4_DO_SRAM23(fabric_sram1_do_i[23]),
        .Tile_X11Y4_DO_SRAM24(fabric_sram1_do_i[24]),
        .Tile_X11Y4_DO_SRAM25(fabric_sram1_do_i[25]),
        .Tile_X11Y4_DO_SRAM26(fabric_sram1_do_i[26]),
        .Tile_X11Y4_DO_SRAM27(fabric_sram1_do_i[27]),
        .Tile_X11Y4_DO_SRAM28(fabric_sram1_do_i[28]),
        .Tile_X11Y4_DO_SRAM29(fabric_sram1_do_i[29]),
        .Tile_X11Y4_DO_SRAM30(fabric_sram1_do_i[30]),
        .Tile_X11Y4_DO_SRAM31(fabric_sram1_do_i[31]),
        .Tile_X11Y4_AD_SRAM0(fabric_sram1_ad_o[0]),
        .Tile_X11Y4_AD_SRAM1(fabric_sram1_ad_o[1]),
        .Tile_X11Y4_AD_SRAM2(fabric_sram1_ad_o[2]),
        .Tile_X11Y4_AD_SRAM3(fabric_sram1_ad_o[3]),
        .Tile_X11Y4_AD_SRAM4(fabric_sram1_ad_o[4]),
        .Tile_X11Y4_AD_SRAM5(fabric_sram1_ad_o[5]),
        .Tile_X11Y4_AD_SRAM6(fabric_sram1_ad_o[6]),
        .Tile_X11Y4_AD_SRAM7(fabric_sram1_ad_o[7]),
        .Tile_X11Y4_AD_SRAM8(fabric_sram1_ad_o[8]),
        .Tile_X11Y4_AD_SRAM9(fabric_sram1_ad_o[9]),
        .Tile_X11Y4_BEN_SRAM0(fabric_sram1_ben_o[0]),
        .Tile_X11Y4_BEN_SRAM1(fabric_sram1_ben_o[1]),
        .Tile_X11Y4_BEN_SRAM2(fabric_sram1_ben_o[2]),
        .Tile_X11Y4_BEN_SRAM3(fabric_sram1_ben_o[3]),
        .Tile_X11Y4_BEN_SRAM4(fabric_sram1_ben_o[4]),
        .Tile_X11Y4_BEN_SRAM5(fabric_sram1_ben_o[5]),
        .Tile_X11Y4_BEN_SRAM6(fabric_sram1_ben_o[6]),
        .Tile_X11Y4_BEN_SRAM7(fabric_sram1_ben_o[7]),
        .Tile_X11Y4_BEN_SRAM8(fabric_sram1_ben_o[8]),
        .Tile_X11Y4_BEN_SRAM9(fabric_sram1_ben_o[9]),
        .Tile_X11Y4_BEN_SRAM10(fabric_sram1_ben_o[10]),
        .Tile_X11Y4_BEN_SRAM11(fabric_sram1_ben_o[11]),
        .Tile_X11Y4_BEN_SRAM12(fabric_sram1_ben_o[12]),
        .Tile_X11Y4_BEN_SRAM13(fabric_sram1_ben_o[13]),
        .Tile_X11Y4_BEN_SRAM14(fabric_sram1_ben_o[14]),
        .Tile_X11Y4_BEN_SRAM15(fabric_sram1_ben_o[15]),
        .Tile_X11Y4_BEN_SRAM16(fabric_sram1_ben_o[16]),
        .Tile_X11Y4_BEN_SRAM17(fabric_sram1_ben_o[17]),
        .Tile_X11Y4_BEN_SRAM18(fabric_sram1_ben_o[18]),
        .Tile_X11Y4_BEN_SRAM19(fabric_sram1_ben_o[19]),
        .Tile_X11Y4_BEN_SRAM20(fabric_sram1_ben_o[20]),
        .Tile_X11Y4_BEN_SRAM21(fabric_sram1_ben_o[21]),
        .Tile_X11Y4_BEN_SRAM22(fabric_sram1_ben_o[22]),
        .Tile_X11Y4_BEN_SRAM23(fabric_sram1_ben_o[23]),
        .Tile_X11Y4_BEN_SRAM24(fabric_sram1_ben_o[24]),
        .Tile_X11Y4_BEN_SRAM25(fabric_sram1_ben_o[25]),
        .Tile_X11Y4_BEN_SRAM26(fabric_sram1_ben_o[26]),
        .Tile_X11Y4_BEN_SRAM27(fabric_sram1_ben_o[27]),
        .Tile_X11Y4_BEN_SRAM28(fabric_sram1_ben_o[28]),
        .Tile_X11Y4_BEN_SRAM29(fabric_sram1_ben_o[29]),
        .Tile_X11Y4_BEN_SRAM30(fabric_sram1_ben_o[30]),
        .Tile_X11Y4_BEN_SRAM31(fabric_sram1_ben_o[31]),
        .Tile_X11Y4_DI_SRAM0(fabric_sram1_di_o[0]),
        .Tile_X11Y4_DI_SRAM1(fabric_sram1_di_o[1]),
        .Tile_X11Y4_DI_SRAM2(fabric_sram1_di_o[2]),
        .Tile_X11Y4_DI_SRAM3(fabric_sram1_di_o[3]),
        .Tile_X11Y4_DI_SRAM4(fabric_sram1_di_o[4]),
        .Tile_X11Y4_DI_SRAM5(fabric_sram1_di_o[5]),
        .Tile_X11Y4_DI_SRAM6(fabric_sram1_di_o[6]),
        .Tile_X11Y4_DI_SRAM7(fabric_sram1_di_o[7]),
        .Tile_X11Y4_DI_SRAM8(fabric_sram1_di_o[8]),
        .Tile_X11Y4_DI_SRAM9(fabric_sram1_di_o[9]),
        .Tile_X11Y4_DI_SRAM10(fabric_sram1_di_o[10]),
        .Tile_X11Y4_DI_SRAM11(fabric_sram1_di_o[11]),
        .Tile_X11Y4_DI_SRAM12(fabric_sram1_di_o[12]),
        .Tile_X11Y4_DI_SRAM13(fabric_sram1_di_o[13]),
        .Tile_X11Y4_DI_SRAM14(fabric_sram1_di_o[14]),
        .Tile_X11Y4_DI_SRAM15(fabric_sram1_di_o[15]),
        .Tile_X11Y4_DI_SRAM16(fabric_sram1_di_o[16]),
        .Tile_X11Y4_DI_SRAM17(fabric_sram1_di_o[17]),
        .Tile_X11Y4_DI_SRAM18(fabric_sram1_di_o[18]),
        .Tile_X11Y4_DI_SRAM19(fabric_sram1_di_o[19]),
        .Tile_X11Y4_DI_SRAM20(fabric_sram1_di_o[20]),
        .Tile_X11Y4_DI_SRAM21(fabric_sram1_di_o[21]),
        .Tile_X11Y4_DI_SRAM22(fabric_sram1_di_o[22]),
        .Tile_X11Y4_DI_SRAM23(fabric_sram1_di_o[23]),
        .Tile_X11Y4_DI_SRAM24(fabric_sram1_di_o[24]),
        .Tile_X11Y4_DI_SRAM25(fabric_sram1_di_o[25]),
        .Tile_X11Y4_DI_SRAM26(fabric_sram1_di_o[26]),
        .Tile_X11Y4_DI_SRAM27(fabric_sram1_di_o[27]),
        .Tile_X11Y4_DI_SRAM28(fabric_sram1_di_o[28]),
        .Tile_X11Y4_DI_SRAM29(fabric_sram1_di_o[29]),
        .Tile_X11Y4_DI_SRAM30(fabric_sram1_di_o[30]),
        .Tile_X11Y4_DI_SRAM31(fabric_sram1_di_o[31]),
        .Tile_X11Y4_EN_SRAM(fabric_sram1_en),
        .Tile_X11Y4_R_WB_SRAM(fabric_sram1_rw_no),
        .Tile_X11Y4_CLOCK_SRAM(fabric_sram1_clk_o),

        // SRAM 2
        .Tile_X11Y6_DO_SRAM0(fabric_sram2_do_i[0]),
        .Tile_X11Y6_DO_SRAM1(fabric_sram2_do_i[1]),
        .Tile_X11Y6_DO_SRAM2(fabric_sram2_do_i[2]),
        .Tile_X11Y6_DO_SRAM3(fabric_sram2_do_i[3]),
        .Tile_X11Y6_DO_SRAM4(fabric_sram2_do_i[4]),
        .Tile_X11Y6_DO_SRAM5(fabric_sram2_do_i[5]),
        .Tile_X11Y6_DO_SRAM6(fabric_sram2_do_i[6]),
        .Tile_X11Y6_DO_SRAM7(fabric_sram2_do_i[7]),
        .Tile_X11Y6_DO_SRAM8(fabric_sram2_do_i[8]),
        .Tile_X11Y6_DO_SRAM9(fabric_sram2_do_i[9]),
        .Tile_X11Y6_DO_SRAM10(fabric_sram2_do_i[10]),
        .Tile_X11Y6_DO_SRAM11(fabric_sram2_do_i[11]),
        .Tile_X11Y6_DO_SRAM12(fabric_sram2_do_i[12]),
        .Tile_X11Y6_DO_SRAM13(fabric_sram2_do_i[13]),
        .Tile_X11Y6_DO_SRAM14(fabric_sram2_do_i[14]),
        .Tile_X11Y6_DO_SRAM15(fabric_sram2_do_i[15]),
        .Tile_X11Y6_DO_SRAM16(fabric_sram2_do_i[16]),
        .Tile_X11Y6_DO_SRAM17(fabric_sram2_do_i[17]),
        .Tile_X11Y6_DO_SRAM18(fabric_sram2_do_i[18]),
        .Tile_X11Y6_DO_SRAM19(fabric_sram2_do_i[19]),
        .Tile_X11Y6_DO_SRAM20(fabric_sram2_do_i[20]),
        .Tile_X11Y6_DO_SRAM21(fabric_sram2_do_i[21]),
        .Tile_X11Y6_DO_SRAM22(fabric_sram2_do_i[22]),
        .Tile_X11Y6_DO_SRAM23(fabric_sram2_do_i[23]),
        .Tile_X11Y6_DO_SRAM24(fabric_sram2_do_i[24]),
        .Tile_X11Y6_DO_SRAM25(fabric_sram2_do_i[25]),
        .Tile_X11Y6_DO_SRAM26(fabric_sram2_do_i[26]),
        .Tile_X11Y6_DO_SRAM27(fabric_sram2_do_i[27]),
        .Tile_X11Y6_DO_SRAM28(fabric_sram2_do_i[28]),
        .Tile_X11Y6_DO_SRAM29(fabric_sram2_do_i[29]),
        .Tile_X11Y6_DO_SRAM30(fabric_sram2_do_i[30]),
        .Tile_X11Y6_DO_SRAM31(fabric_sram2_do_i[31]),
        .Tile_X11Y6_AD_SRAM0(fabric_sram2_ad_o[0]),
        .Tile_X11Y6_AD_SRAM1(fabric_sram2_ad_o[1]),
        .Tile_X11Y6_AD_SRAM2(fabric_sram2_ad_o[2]),
        .Tile_X11Y6_AD_SRAM3(fabric_sram2_ad_o[3]),
        .Tile_X11Y6_AD_SRAM4(fabric_sram2_ad_o[4]),
        .Tile_X11Y6_AD_SRAM5(fabric_sram2_ad_o[5]),
        .Tile_X11Y6_AD_SRAM6(fabric_sram2_ad_o[6]),
        .Tile_X11Y6_AD_SRAM7(fabric_sram2_ad_o[7]),
        .Tile_X11Y6_AD_SRAM8(fabric_sram2_ad_o[8]),
        .Tile_X11Y6_AD_SRAM9(fabric_sram2_ad_o[9]),
        .Tile_X11Y6_BEN_SRAM0(fabric_sram2_ben_o[0]),
        .Tile_X11Y6_BEN_SRAM1(fabric_sram2_ben_o[1]),
        .Tile_X11Y6_BEN_SRAM2(fabric_sram2_ben_o[2]),
        .Tile_X11Y6_BEN_SRAM3(fabric_sram2_ben_o[3]),
        .Tile_X11Y6_BEN_SRAM4(fabric_sram2_ben_o[4]),
        .Tile_X11Y6_BEN_SRAM5(fabric_sram2_ben_o[5]),
        .Tile_X11Y6_BEN_SRAM6(fabric_sram2_ben_o[6]),
        .Tile_X11Y6_BEN_SRAM7(fabric_sram2_ben_o[7]),
        .Tile_X11Y6_BEN_SRAM8(fabric_sram2_ben_o[8]),
        .Tile_X11Y6_BEN_SRAM9(fabric_sram2_ben_o[9]),
        .Tile_X11Y6_BEN_SRAM10(fabric_sram2_ben_o[10]),
        .Tile_X11Y6_BEN_SRAM11(fabric_sram2_ben_o[11]),
        .Tile_X11Y6_BEN_SRAM12(fabric_sram2_ben_o[12]),
        .Tile_X11Y6_BEN_SRAM13(fabric_sram2_ben_o[13]),
        .Tile_X11Y6_BEN_SRAM14(fabric_sram2_ben_o[14]),
        .Tile_X11Y6_BEN_SRAM15(fabric_sram2_ben_o[15]),
        .Tile_X11Y6_BEN_SRAM16(fabric_sram2_ben_o[16]),
        .Tile_X11Y6_BEN_SRAM17(fabric_sram2_ben_o[17]),
        .Tile_X11Y6_BEN_SRAM18(fabric_sram2_ben_o[18]),
        .Tile_X11Y6_BEN_SRAM19(fabric_sram2_ben_o[19]),
        .Tile_X11Y6_BEN_SRAM20(fabric_sram2_ben_o[20]),
        .Tile_X11Y6_BEN_SRAM21(fabric_sram2_ben_o[21]),
        .Tile_X11Y6_BEN_SRAM22(fabric_sram2_ben_o[22]),
        .Tile_X11Y6_BEN_SRAM23(fabric_sram2_ben_o[23]),
        .Tile_X11Y6_BEN_SRAM24(fabric_sram2_ben_o[24]),
        .Tile_X11Y6_BEN_SRAM25(fabric_sram2_ben_o[25]),
        .Tile_X11Y6_BEN_SRAM26(fabric_sram2_ben_o[26]),
        .Tile_X11Y6_BEN_SRAM27(fabric_sram2_ben_o[27]),
        .Tile_X11Y6_BEN_SRAM28(fabric_sram2_ben_o[28]),
        .Tile_X11Y6_BEN_SRAM29(fabric_sram2_ben_o[29]),
        .Tile_X11Y6_BEN_SRAM30(fabric_sram2_ben_o[30]),
        .Tile_X11Y6_BEN_SRAM31(fabric_sram2_ben_o[31]),
        .Tile_X11Y6_DI_SRAM0(fabric_sram2_di_o[0]),
        .Tile_X11Y6_DI_SRAM1(fabric_sram2_di_o[1]),
        .Tile_X11Y6_DI_SRAM2(fabric_sram2_di_o[2]),
        .Tile_X11Y6_DI_SRAM3(fabric_sram2_di_o[3]),
        .Tile_X11Y6_DI_SRAM4(fabric_sram2_di_o[4]),
        .Tile_X11Y6_DI_SRAM5(fabric_sram2_di_o[5]),
        .Tile_X11Y6_DI_SRAM6(fabric_sram2_di_o[6]),
        .Tile_X11Y6_DI_SRAM7(fabric_sram2_di_o[7]),
        .Tile_X11Y6_DI_SRAM8(fabric_sram2_di_o[8]),
        .Tile_X11Y6_DI_SRAM9(fabric_sram2_di_o[9]),
        .Tile_X11Y6_DI_SRAM10(fabric_sram2_di_o[10]),
        .Tile_X11Y6_DI_SRAM11(fabric_sram2_di_o[11]),
        .Tile_X11Y6_DI_SRAM12(fabric_sram2_di_o[12]),
        .Tile_X11Y6_DI_SRAM13(fabric_sram2_di_o[13]),
        .Tile_X11Y6_DI_SRAM14(fabric_sram2_di_o[14]),
        .Tile_X11Y6_DI_SRAM15(fabric_sram2_di_o[15]),
        .Tile_X11Y6_DI_SRAM16(fabric_sram2_di_o[16]),
        .Tile_X11Y6_DI_SRAM17(fabric_sram2_di_o[17]),
        .Tile_X11Y6_DI_SRAM18(fabric_sram2_di_o[18]),
        .Tile_X11Y6_DI_SRAM19(fabric_sram2_di_o[19]),
        .Tile_X11Y6_DI_SRAM20(fabric_sram2_di_o[20]),
        .Tile_X11Y6_DI_SRAM21(fabric_sram2_di_o[21]),
        .Tile_X11Y6_DI_SRAM22(fabric_sram2_di_o[22]),
        .Tile_X11Y6_DI_SRAM23(fabric_sram2_di_o[23]),
        .Tile_X11Y6_DI_SRAM24(fabric_sram2_di_o[24]),
        .Tile_X11Y6_DI_SRAM25(fabric_sram2_di_o[25]),
        .Tile_X11Y6_DI_SRAM26(fabric_sram2_di_o[26]),
        .Tile_X11Y6_DI_SRAM27(fabric_sram2_di_o[27]),
        .Tile_X11Y6_DI_SRAM28(fabric_sram2_di_o[28]),
        .Tile_X11Y6_DI_SRAM29(fabric_sram2_di_o[29]),
        .Tile_X11Y6_DI_SRAM30(fabric_sram2_di_o[30]),
        .Tile_X11Y6_DI_SRAM31(fabric_sram2_di_o[31]),
        .Tile_X11Y6_EN_SRAM(fabric_sram2_en),
        .Tile_X11Y6_R_WB_SRAM(fabric_sram2_rw_no),
        .Tile_X11Y6_CLOCK_SRAM(fabric_sram2_clk_o),

        // SRAM 3
        .Tile_X11Y8_DO_SRAM0(fabric_sram3_do_i[0]),
        .Tile_X11Y8_DO_SRAM1(fabric_sram3_do_i[1]),
        .Tile_X11Y8_DO_SRAM2(fabric_sram3_do_i[2]),
        .Tile_X11Y8_DO_SRAM3(fabric_sram3_do_i[3]),
        .Tile_X11Y8_DO_SRAM4(fabric_sram3_do_i[4]),
        .Tile_X11Y8_DO_SRAM5(fabric_sram3_do_i[5]),
        .Tile_X11Y8_DO_SRAM6(fabric_sram3_do_i[6]),
        .Tile_X11Y8_DO_SRAM7(fabric_sram3_do_i[7]),
        .Tile_X11Y8_DO_SRAM8(fabric_sram3_do_i[8]),
        .Tile_X11Y8_DO_SRAM9(fabric_sram3_do_i[9]),
        .Tile_X11Y8_DO_SRAM10(fabric_sram3_do_i[10]),
        .Tile_X11Y8_DO_SRAM11(fabric_sram3_do_i[11]),
        .Tile_X11Y8_DO_SRAM12(fabric_sram3_do_i[12]),
        .Tile_X11Y8_DO_SRAM13(fabric_sram3_do_i[13]),
        .Tile_X11Y8_DO_SRAM14(fabric_sram3_do_i[14]),
        .Tile_X11Y8_DO_SRAM15(fabric_sram3_do_i[15]),
        .Tile_X11Y8_DO_SRAM16(fabric_sram3_do_i[16]),
        .Tile_X11Y8_DO_SRAM17(fabric_sram3_do_i[17]),
        .Tile_X11Y8_DO_SRAM18(fabric_sram3_do_i[18]),
        .Tile_X11Y8_DO_SRAM19(fabric_sram3_do_i[19]),
        .Tile_X11Y8_DO_SRAM20(fabric_sram3_do_i[20]),
        .Tile_X11Y8_DO_SRAM21(fabric_sram3_do_i[21]),
        .Tile_X11Y8_DO_SRAM22(fabric_sram3_do_i[22]),
        .Tile_X11Y8_DO_SRAM23(fabric_sram3_do_i[23]),
        .Tile_X11Y8_DO_SRAM24(fabric_sram3_do_i[24]),
        .Tile_X11Y8_DO_SRAM25(fabric_sram3_do_i[25]),
        .Tile_X11Y8_DO_SRAM26(fabric_sram3_do_i[26]),
        .Tile_X11Y8_DO_SRAM27(fabric_sram3_do_i[27]),
        .Tile_X11Y8_DO_SRAM28(fabric_sram3_do_i[28]),
        .Tile_X11Y8_DO_SRAM29(fabric_sram3_do_i[29]),
        .Tile_X11Y8_DO_SRAM30(fabric_sram3_do_i[30]),
        .Tile_X11Y8_DO_SRAM31(fabric_sram3_do_i[31]),
        .Tile_X11Y8_AD_SRAM0(fabric_sram3_ad_o[0]),
        .Tile_X11Y8_AD_SRAM1(fabric_sram3_ad_o[1]),
        .Tile_X11Y8_AD_SRAM2(fabric_sram3_ad_o[2]),
        .Tile_X11Y8_AD_SRAM3(fabric_sram3_ad_o[3]),
        .Tile_X11Y8_AD_SRAM4(fabric_sram3_ad_o[4]),
        .Tile_X11Y8_AD_SRAM5(fabric_sram3_ad_o[5]),
        .Tile_X11Y8_AD_SRAM6(fabric_sram3_ad_o[6]),
        .Tile_X11Y8_AD_SRAM7(fabric_sram3_ad_o[7]),
        .Tile_X11Y8_AD_SRAM8(fabric_sram3_ad_o[8]),
        .Tile_X11Y8_AD_SRAM9(fabric_sram3_ad_o[9]),
        .Tile_X11Y8_BEN_SRAM0(fabric_sram3_ben_o[0]),
        .Tile_X11Y8_BEN_SRAM1(fabric_sram3_ben_o[1]),
        .Tile_X11Y8_BEN_SRAM2(fabric_sram3_ben_o[2]),
        .Tile_X11Y8_BEN_SRAM3(fabric_sram3_ben_o[3]),
        .Tile_X11Y8_BEN_SRAM4(fabric_sram3_ben_o[4]),
        .Tile_X11Y8_BEN_SRAM5(fabric_sram3_ben_o[5]),
        .Tile_X11Y8_BEN_SRAM6(fabric_sram3_ben_o[6]),
        .Tile_X11Y8_BEN_SRAM7(fabric_sram3_ben_o[7]),
        .Tile_X11Y8_BEN_SRAM8(fabric_sram3_ben_o[8]),
        .Tile_X11Y8_BEN_SRAM9(fabric_sram3_ben_o[9]),
        .Tile_X11Y8_BEN_SRAM10(fabric_sram3_ben_o[10]),
        .Tile_X11Y8_BEN_SRAM11(fabric_sram3_ben_o[11]),
        .Tile_X11Y8_BEN_SRAM12(fabric_sram3_ben_o[12]),
        .Tile_X11Y8_BEN_SRAM13(fabric_sram3_ben_o[13]),
        .Tile_X11Y8_BEN_SRAM14(fabric_sram3_ben_o[14]),
        .Tile_X11Y8_BEN_SRAM15(fabric_sram3_ben_o[15]),
        .Tile_X11Y8_BEN_SRAM16(fabric_sram3_ben_o[16]),
        .Tile_X11Y8_BEN_SRAM17(fabric_sram3_ben_o[17]),
        .Tile_X11Y8_BEN_SRAM18(fabric_sram3_ben_o[18]),
        .Tile_X11Y8_BEN_SRAM19(fabric_sram3_ben_o[19]),
        .Tile_X11Y8_BEN_SRAM20(fabric_sram3_ben_o[20]),
        .Tile_X11Y8_BEN_SRAM21(fabric_sram3_ben_o[21]),
        .Tile_X11Y8_BEN_SRAM22(fabric_sram3_ben_o[22]),
        .Tile_X11Y8_BEN_SRAM23(fabric_sram3_ben_o[23]),
        .Tile_X11Y8_BEN_SRAM24(fabric_sram3_ben_o[24]),
        .Tile_X11Y8_BEN_SRAM25(fabric_sram3_ben_o[25]),
        .Tile_X11Y8_BEN_SRAM26(fabric_sram3_ben_o[26]),
        .Tile_X11Y8_BEN_SRAM27(fabric_sram3_ben_o[27]),
        .Tile_X11Y8_BEN_SRAM28(fabric_sram3_ben_o[28]),
        .Tile_X11Y8_BEN_SRAM29(fabric_sram3_ben_o[29]),
        .Tile_X11Y8_BEN_SRAM30(fabric_sram3_ben_o[30]),
        .Tile_X11Y8_BEN_SRAM31(fabric_sram3_ben_o[31]),
        .Tile_X11Y8_DI_SRAM0(fabric_sram3_di_o[0]),
        .Tile_X11Y8_DI_SRAM1(fabric_sram3_di_o[1]),
        .Tile_X11Y8_DI_SRAM2(fabric_sram3_di_o[2]),
        .Tile_X11Y8_DI_SRAM3(fabric_sram3_di_o[3]),
        .Tile_X11Y8_DI_SRAM4(fabric_sram3_di_o[4]),
        .Tile_X11Y8_DI_SRAM5(fabric_sram3_di_o[5]),
        .Tile_X11Y8_DI_SRAM6(fabric_sram3_di_o[6]),
        .Tile_X11Y8_DI_SRAM7(fabric_sram3_di_o[7]),
        .Tile_X11Y8_DI_SRAM8(fabric_sram3_di_o[8]),
        .Tile_X11Y8_DI_SRAM9(fabric_sram3_di_o[9]),
        .Tile_X11Y8_DI_SRAM10(fabric_sram3_di_o[10]),
        .Tile_X11Y8_DI_SRAM11(fabric_sram3_di_o[11]),
        .Tile_X11Y8_DI_SRAM12(fabric_sram3_di_o[12]),
        .Tile_X11Y8_DI_SRAM13(fabric_sram3_di_o[13]),
        .Tile_X11Y8_DI_SRAM14(fabric_sram3_di_o[14]),
        .Tile_X11Y8_DI_SRAM15(fabric_sram3_di_o[15]),
        .Tile_X11Y8_DI_SRAM16(fabric_sram3_di_o[16]),
        .Tile_X11Y8_DI_SRAM17(fabric_sram3_di_o[17]),
        .Tile_X11Y8_DI_SRAM18(fabric_sram3_di_o[18]),
        .Tile_X11Y8_DI_SRAM19(fabric_sram3_di_o[19]),
        .Tile_X11Y8_DI_SRAM20(fabric_sram3_di_o[20]),
        .Tile_X11Y8_DI_SRAM21(fabric_sram3_di_o[21]),
        .Tile_X11Y8_DI_SRAM22(fabric_sram3_di_o[22]),
        .Tile_X11Y8_DI_SRAM23(fabric_sram3_di_o[23]),
        .Tile_X11Y8_DI_SRAM24(fabric_sram3_di_o[24]),
        .Tile_X11Y8_DI_SRAM25(fabric_sram3_di_o[25]),
        .Tile_X11Y8_DI_SRAM26(fabric_sram3_di_o[26]),
        .Tile_X11Y8_DI_SRAM27(fabric_sram3_di_o[27]),
        .Tile_X11Y8_DI_SRAM28(fabric_sram3_di_o[28]),
        .Tile_X11Y8_DI_SRAM29(fabric_sram3_di_o[29]),
        .Tile_X11Y8_DI_SRAM30(fabric_sram3_di_o[30]),
        .Tile_X11Y8_DI_SRAM31(fabric_sram3_di_o[31]),
        .Tile_X11Y8_EN_SRAM(fabric_sram3_en),
        .Tile_X11Y8_R_WB_SRAM(fabric_sram3_rw_no),
        .Tile_X11Y8_CLOCK_SRAM(fabric_sram3_clk_o),

        // SRAM 4
        .Tile_X11Y10_DO_SRAM0(fabric_sram4_do_i[0]),
        .Tile_X11Y10_DO_SRAM1(fabric_sram4_do_i[1]),
        .Tile_X11Y10_DO_SRAM2(fabric_sram4_do_i[2]),
        .Tile_X11Y10_DO_SRAM3(fabric_sram4_do_i[3]),
        .Tile_X11Y10_DO_SRAM4(fabric_sram4_do_i[4]),
        .Tile_X11Y10_DO_SRAM5(fabric_sram4_do_i[5]),
        .Tile_X11Y10_DO_SRAM6(fabric_sram4_do_i[6]),
        .Tile_X11Y10_DO_SRAM7(fabric_sram4_do_i[7]),
        .Tile_X11Y10_DO_SRAM8(fabric_sram4_do_i[8]),
        .Tile_X11Y10_DO_SRAM9(fabric_sram4_do_i[9]),
        .Tile_X11Y10_DO_SRAM10(fabric_sram4_do_i[10]),
        .Tile_X11Y10_DO_SRAM11(fabric_sram4_do_i[11]),
        .Tile_X11Y10_DO_SRAM12(fabric_sram4_do_i[12]),
        .Tile_X11Y10_DO_SRAM13(fabric_sram4_do_i[13]),
        .Tile_X11Y10_DO_SRAM14(fabric_sram4_do_i[14]),
        .Tile_X11Y10_DO_SRAM15(fabric_sram4_do_i[15]),
        .Tile_X11Y10_DO_SRAM16(fabric_sram4_do_i[16]),
        .Tile_X11Y10_DO_SRAM17(fabric_sram4_do_i[17]),
        .Tile_X11Y10_DO_SRAM18(fabric_sram4_do_i[18]),
        .Tile_X11Y10_DO_SRAM19(fabric_sram4_do_i[19]),
        .Tile_X11Y10_DO_SRAM20(fabric_sram4_do_i[20]),
        .Tile_X11Y10_DO_SRAM21(fabric_sram4_do_i[21]),
        .Tile_X11Y10_DO_SRAM22(fabric_sram4_do_i[22]),
        .Tile_X11Y10_DO_SRAM23(fabric_sram4_do_i[23]),
        .Tile_X11Y10_DO_SRAM24(fabric_sram4_do_i[24]),
        .Tile_X11Y10_DO_SRAM25(fabric_sram4_do_i[25]),
        .Tile_X11Y10_DO_SRAM26(fabric_sram4_do_i[26]),
        .Tile_X11Y10_DO_SRAM27(fabric_sram4_do_i[27]),
        .Tile_X11Y10_DO_SRAM28(fabric_sram4_do_i[28]),
        .Tile_X11Y10_DO_SRAM29(fabric_sram4_do_i[29]),
        .Tile_X11Y10_DO_SRAM30(fabric_sram4_do_i[30]),
        .Tile_X11Y10_DO_SRAM31(fabric_sram4_do_i[31]),
        .Tile_X11Y10_AD_SRAM0(fabric_sram4_ad_o[0]),
        .Tile_X11Y10_AD_SRAM1(fabric_sram4_ad_o[1]),
        .Tile_X11Y10_AD_SRAM2(fabric_sram4_ad_o[2]),
        .Tile_X11Y10_AD_SRAM3(fabric_sram4_ad_o[3]),
        .Tile_X11Y10_AD_SRAM4(fabric_sram4_ad_o[4]),
        .Tile_X11Y10_AD_SRAM5(fabric_sram4_ad_o[5]),
        .Tile_X11Y10_AD_SRAM6(fabric_sram4_ad_o[6]),
        .Tile_X11Y10_AD_SRAM7(fabric_sram4_ad_o[7]),
        .Tile_X11Y10_AD_SRAM8(fabric_sram4_ad_o[8]),
        .Tile_X11Y10_AD_SRAM9(fabric_sram4_ad_o[9]),
        .Tile_X11Y10_BEN_SRAM0(fabric_sram4_ben_o[0]),
        .Tile_X11Y10_BEN_SRAM1(fabric_sram4_ben_o[1]),
        .Tile_X11Y10_BEN_SRAM2(fabric_sram4_ben_o[2]),
        .Tile_X11Y10_BEN_SRAM3(fabric_sram4_ben_o[3]),
        .Tile_X11Y10_BEN_SRAM4(fabric_sram4_ben_o[4]),
        .Tile_X11Y10_BEN_SRAM5(fabric_sram4_ben_o[5]),
        .Tile_X11Y10_BEN_SRAM6(fabric_sram4_ben_o[6]),
        .Tile_X11Y10_BEN_SRAM7(fabric_sram4_ben_o[7]),
        .Tile_X11Y10_BEN_SRAM8(fabric_sram4_ben_o[8]),
        .Tile_X11Y10_BEN_SRAM9(fabric_sram4_ben_o[9]),
        .Tile_X11Y10_BEN_SRAM10(fabric_sram4_ben_o[10]),
        .Tile_X11Y10_BEN_SRAM11(fabric_sram4_ben_o[11]),
        .Tile_X11Y10_BEN_SRAM12(fabric_sram4_ben_o[12]),
        .Tile_X11Y10_BEN_SRAM13(fabric_sram4_ben_o[13]),
        .Tile_X11Y10_BEN_SRAM14(fabric_sram4_ben_o[14]),
        .Tile_X11Y10_BEN_SRAM15(fabric_sram4_ben_o[15]),
        .Tile_X11Y10_BEN_SRAM16(fabric_sram4_ben_o[16]),
        .Tile_X11Y10_BEN_SRAM17(fabric_sram4_ben_o[17]),
        .Tile_X11Y10_BEN_SRAM18(fabric_sram4_ben_o[18]),
        .Tile_X11Y10_BEN_SRAM19(fabric_sram4_ben_o[19]),
        .Tile_X11Y10_BEN_SRAM20(fabric_sram4_ben_o[20]),
        .Tile_X11Y10_BEN_SRAM21(fabric_sram4_ben_o[21]),
        .Tile_X11Y10_BEN_SRAM22(fabric_sram4_ben_o[22]),
        .Tile_X11Y10_BEN_SRAM23(fabric_sram4_ben_o[23]),
        .Tile_X11Y10_BEN_SRAM24(fabric_sram4_ben_o[24]),
        .Tile_X11Y10_BEN_SRAM25(fabric_sram4_ben_o[25]),
        .Tile_X11Y10_BEN_SRAM26(fabric_sram4_ben_o[26]),
        .Tile_X11Y10_BEN_SRAM27(fabric_sram4_ben_o[27]),
        .Tile_X11Y10_BEN_SRAM28(fabric_sram4_ben_o[28]),
        .Tile_X11Y10_BEN_SRAM29(fabric_sram4_ben_o[29]),
        .Tile_X11Y10_BEN_SRAM30(fabric_sram4_ben_o[30]),
        .Tile_X11Y10_BEN_SRAM31(fabric_sram4_ben_o[31]),
        .Tile_X11Y10_DI_SRAM0(fabric_sram4_di_o[0]),
        .Tile_X11Y10_DI_SRAM1(fabric_sram4_di_o[1]),
        .Tile_X11Y10_DI_SRAM2(fabric_sram4_di_o[2]),
        .Tile_X11Y10_DI_SRAM3(fabric_sram4_di_o[3]),
        .Tile_X11Y10_DI_SRAM4(fabric_sram4_di_o[4]),
        .Tile_X11Y10_DI_SRAM5(fabric_sram4_di_o[5]),
        .Tile_X11Y10_DI_SRAM6(fabric_sram4_di_o[6]),
        .Tile_X11Y10_DI_SRAM7(fabric_sram4_di_o[7]),
        .Tile_X11Y10_DI_SRAM8(fabric_sram4_di_o[8]),
        .Tile_X11Y10_DI_SRAM9(fabric_sram4_di_o[9]),
        .Tile_X11Y10_DI_SRAM10(fabric_sram4_di_o[10]),
        .Tile_X11Y10_DI_SRAM11(fabric_sram4_di_o[11]),
        .Tile_X11Y10_DI_SRAM12(fabric_sram4_di_o[12]),
        .Tile_X11Y10_DI_SRAM13(fabric_sram4_di_o[13]),
        .Tile_X11Y10_DI_SRAM14(fabric_sram4_di_o[14]),
        .Tile_X11Y10_DI_SRAM15(fabric_sram4_di_o[15]),
        .Tile_X11Y10_DI_SRAM16(fabric_sram4_di_o[16]),
        .Tile_X11Y10_DI_SRAM17(fabric_sram4_di_o[17]),
        .Tile_X11Y10_DI_SRAM18(fabric_sram4_di_o[18]),
        .Tile_X11Y10_DI_SRAM19(fabric_sram4_di_o[19]),
        .Tile_X11Y10_DI_SRAM20(fabric_sram4_di_o[20]),
        .Tile_X11Y10_DI_SRAM21(fabric_sram4_di_o[21]),
        .Tile_X11Y10_DI_SRAM22(fabric_sram4_di_o[22]),
        .Tile_X11Y10_DI_SRAM23(fabric_sram4_di_o[23]),
        .Tile_X11Y10_DI_SRAM24(fabric_sram4_di_o[24]),
        .Tile_X11Y10_DI_SRAM25(fabric_sram4_di_o[25]),
        .Tile_X11Y10_DI_SRAM26(fabric_sram4_di_o[26]),
        .Tile_X11Y10_DI_SRAM27(fabric_sram4_di_o[27]),
        .Tile_X11Y10_DI_SRAM28(fabric_sram4_di_o[28]),
        .Tile_X11Y10_DI_SRAM29(fabric_sram4_di_o[29]),
        .Tile_X11Y10_DI_SRAM30(fabric_sram4_di_o[30]),
        .Tile_X11Y10_DI_SRAM31(fabric_sram4_di_o[31]),
        .Tile_X11Y10_EN_SRAM(fabric_sram4_en),
        .Tile_X11Y10_R_WB_SRAM(fabric_sram4_rw_no),
        .Tile_X11Y10_CLOCK_SRAM(fabric_sram4_clk_o),

        // SRAM 5
        .Tile_X11Y12_DO_SRAM0(fabric_sram5_do_i[0]),
        .Tile_X11Y12_DO_SRAM1(fabric_sram5_do_i[1]),
        .Tile_X11Y12_DO_SRAM2(fabric_sram5_do_i[2]),
        .Tile_X11Y12_DO_SRAM3(fabric_sram5_do_i[3]),
        .Tile_X11Y12_DO_SRAM4(fabric_sram5_do_i[4]),
        .Tile_X11Y12_DO_SRAM5(fabric_sram5_do_i[5]),
        .Tile_X11Y12_DO_SRAM6(fabric_sram5_do_i[6]),
        .Tile_X11Y12_DO_SRAM7(fabric_sram5_do_i[7]),
        .Tile_X11Y12_DO_SRAM8(fabric_sram5_do_i[8]),
        .Tile_X11Y12_DO_SRAM9(fabric_sram5_do_i[9]),
        .Tile_X11Y12_DO_SRAM10(fabric_sram5_do_i[10]),
        .Tile_X11Y12_DO_SRAM11(fabric_sram5_do_i[11]),
        .Tile_X11Y12_DO_SRAM12(fabric_sram5_do_i[12]),
        .Tile_X11Y12_DO_SRAM13(fabric_sram5_do_i[13]),
        .Tile_X11Y12_DO_SRAM14(fabric_sram5_do_i[14]),
        .Tile_X11Y12_DO_SRAM15(fabric_sram5_do_i[15]),
        .Tile_X11Y12_DO_SRAM16(fabric_sram5_do_i[16]),
        .Tile_X11Y12_DO_SRAM17(fabric_sram5_do_i[17]),
        .Tile_X11Y12_DO_SRAM18(fabric_sram5_do_i[18]),
        .Tile_X11Y12_DO_SRAM19(fabric_sram5_do_i[19]),
        .Tile_X11Y12_DO_SRAM20(fabric_sram5_do_i[20]),
        .Tile_X11Y12_DO_SRAM21(fabric_sram5_do_i[21]),
        .Tile_X11Y12_DO_SRAM22(fabric_sram5_do_i[22]),
        .Tile_X11Y12_DO_SRAM23(fabric_sram5_do_i[23]),
        .Tile_X11Y12_DO_SRAM24(fabric_sram5_do_i[24]),
        .Tile_X11Y12_DO_SRAM25(fabric_sram5_do_i[25]),
        .Tile_X11Y12_DO_SRAM26(fabric_sram5_do_i[26]),
        .Tile_X11Y12_DO_SRAM27(fabric_sram5_do_i[27]),
        .Tile_X11Y12_DO_SRAM28(fabric_sram5_do_i[28]),
        .Tile_X11Y12_DO_SRAM29(fabric_sram5_do_i[29]),
        .Tile_X11Y12_DO_SRAM30(fabric_sram5_do_i[30]),
        .Tile_X11Y12_DO_SRAM31(fabric_sram5_do_i[31]),
        .Tile_X11Y12_AD_SRAM0(fabric_sram5_ad_o[0]),
        .Tile_X11Y12_AD_SRAM1(fabric_sram5_ad_o[1]),
        .Tile_X11Y12_AD_SRAM2(fabric_sram5_ad_o[2]),
        .Tile_X11Y12_AD_SRAM3(fabric_sram5_ad_o[3]),
        .Tile_X11Y12_AD_SRAM4(fabric_sram5_ad_o[4]),
        .Tile_X11Y12_AD_SRAM5(fabric_sram5_ad_o[5]),
        .Tile_X11Y12_AD_SRAM6(fabric_sram5_ad_o[6]),
        .Tile_X11Y12_AD_SRAM7(fabric_sram5_ad_o[7]),
        .Tile_X11Y12_AD_SRAM8(fabric_sram5_ad_o[8]),
        .Tile_X11Y12_AD_SRAM9(fabric_sram5_ad_o[9]),
        .Tile_X11Y12_BEN_SRAM0(fabric_sram5_ben_o[0]),
        .Tile_X11Y12_BEN_SRAM1(fabric_sram5_ben_o[1]),
        .Tile_X11Y12_BEN_SRAM2(fabric_sram5_ben_o[2]),
        .Tile_X11Y12_BEN_SRAM3(fabric_sram5_ben_o[3]),
        .Tile_X11Y12_BEN_SRAM4(fabric_sram5_ben_o[4]),
        .Tile_X11Y12_BEN_SRAM5(fabric_sram5_ben_o[5]),
        .Tile_X11Y12_BEN_SRAM6(fabric_sram5_ben_o[6]),
        .Tile_X11Y12_BEN_SRAM7(fabric_sram5_ben_o[7]),
        .Tile_X11Y12_BEN_SRAM8(fabric_sram5_ben_o[8]),
        .Tile_X11Y12_BEN_SRAM9(fabric_sram5_ben_o[9]),
        .Tile_X11Y12_BEN_SRAM10(fabric_sram5_ben_o[10]),
        .Tile_X11Y12_BEN_SRAM11(fabric_sram5_ben_o[11]),
        .Tile_X11Y12_BEN_SRAM12(fabric_sram5_ben_o[12]),
        .Tile_X11Y12_BEN_SRAM13(fabric_sram5_ben_o[13]),
        .Tile_X11Y12_BEN_SRAM14(fabric_sram5_ben_o[14]),
        .Tile_X11Y12_BEN_SRAM15(fabric_sram5_ben_o[15]),
        .Tile_X11Y12_BEN_SRAM16(fabric_sram5_ben_o[16]),
        .Tile_X11Y12_BEN_SRAM17(fabric_sram5_ben_o[17]),
        .Tile_X11Y12_BEN_SRAM18(fabric_sram5_ben_o[18]),
        .Tile_X11Y12_BEN_SRAM19(fabric_sram5_ben_o[19]),
        .Tile_X11Y12_BEN_SRAM20(fabric_sram5_ben_o[20]),
        .Tile_X11Y12_BEN_SRAM21(fabric_sram5_ben_o[21]),
        .Tile_X11Y12_BEN_SRAM22(fabric_sram5_ben_o[22]),
        .Tile_X11Y12_BEN_SRAM23(fabric_sram5_ben_o[23]),
        .Tile_X11Y12_BEN_SRAM24(fabric_sram5_ben_o[24]),
        .Tile_X11Y12_BEN_SRAM25(fabric_sram5_ben_o[25]),
        .Tile_X11Y12_BEN_SRAM26(fabric_sram5_ben_o[26]),
        .Tile_X11Y12_BEN_SRAM27(fabric_sram5_ben_o[27]),
        .Tile_X11Y12_BEN_SRAM28(fabric_sram5_ben_o[28]),
        .Tile_X11Y12_BEN_SRAM29(fabric_sram5_ben_o[29]),
        .Tile_X11Y12_BEN_SRAM30(fabric_sram5_ben_o[30]),
        .Tile_X11Y12_BEN_SRAM31(fabric_sram5_ben_o[31]),
        .Tile_X11Y12_DI_SRAM0(fabric_sram5_di_o[0]),
        .Tile_X11Y12_DI_SRAM1(fabric_sram5_di_o[1]),
        .Tile_X11Y12_DI_SRAM2(fabric_sram5_di_o[2]),
        .Tile_X11Y12_DI_SRAM3(fabric_sram5_di_o[3]),
        .Tile_X11Y12_DI_SRAM4(fabric_sram5_di_o[4]),
        .Tile_X11Y12_DI_SRAM5(fabric_sram5_di_o[5]),
        .Tile_X11Y12_DI_SRAM6(fabric_sram5_di_o[6]),
        .Tile_X11Y12_DI_SRAM7(fabric_sram5_di_o[7]),
        .Tile_X11Y12_DI_SRAM8(fabric_sram5_di_o[8]),
        .Tile_X11Y12_DI_SRAM9(fabric_sram5_di_o[9]),
        .Tile_X11Y12_DI_SRAM10(fabric_sram5_di_o[10]),
        .Tile_X11Y12_DI_SRAM11(fabric_sram5_di_o[11]),
        .Tile_X11Y12_DI_SRAM12(fabric_sram5_di_o[12]),
        .Tile_X11Y12_DI_SRAM13(fabric_sram5_di_o[13]),
        .Tile_X11Y12_DI_SRAM14(fabric_sram5_di_o[14]),
        .Tile_X11Y12_DI_SRAM15(fabric_sram5_di_o[15]),
        .Tile_X11Y12_DI_SRAM16(fabric_sram5_di_o[16]),
        .Tile_X11Y12_DI_SRAM17(fabric_sram5_di_o[17]),
        .Tile_X11Y12_DI_SRAM18(fabric_sram5_di_o[18]),
        .Tile_X11Y12_DI_SRAM19(fabric_sram5_di_o[19]),
        .Tile_X11Y12_DI_SRAM20(fabric_sram5_di_o[20]),
        .Tile_X11Y12_DI_SRAM21(fabric_sram5_di_o[21]),
        .Tile_X11Y12_DI_SRAM22(fabric_sram5_di_o[22]),
        .Tile_X11Y12_DI_SRAM23(fabric_sram5_di_o[23]),
        .Tile_X11Y12_DI_SRAM24(fabric_sram5_di_o[24]),
        .Tile_X11Y12_DI_SRAM25(fabric_sram5_di_o[25]),
        .Tile_X11Y12_DI_SRAM26(fabric_sram5_di_o[26]),
        .Tile_X11Y12_DI_SRAM27(fabric_sram5_di_o[27]),
        .Tile_X11Y12_DI_SRAM28(fabric_sram5_di_o[28]),
        .Tile_X11Y12_DI_SRAM29(fabric_sram5_di_o[29]),
        .Tile_X11Y12_DI_SRAM30(fabric_sram5_di_o[30]),
        .Tile_X11Y12_DI_SRAM31(fabric_sram5_di_o[31]),
        .Tile_X11Y12_EN_SRAM(fabric_sram5_en),
        .Tile_X11Y12_R_WB_SRAM(fabric_sram5_rw_no),
        .Tile_X11Y12_CLOCK_SRAM(fabric_sram5_clk_o),

        // SRAM 6
        .Tile_X11Y14_DO_SRAM0(fabric_sram6_do_i[0]),
        .Tile_X11Y14_DO_SRAM1(fabric_sram6_do_i[1]),
        .Tile_X11Y14_DO_SRAM2(fabric_sram6_do_i[2]),
        .Tile_X11Y14_DO_SRAM3(fabric_sram6_do_i[3]),
        .Tile_X11Y14_DO_SRAM4(fabric_sram6_do_i[4]),
        .Tile_X11Y14_DO_SRAM5(fabric_sram6_do_i[5]),
        .Tile_X11Y14_DO_SRAM6(fabric_sram6_do_i[6]),
        .Tile_X11Y14_DO_SRAM7(fabric_sram6_do_i[7]),
        .Tile_X11Y14_DO_SRAM8(fabric_sram6_do_i[8]),
        .Tile_X11Y14_DO_SRAM9(fabric_sram6_do_i[9]),
        .Tile_X11Y14_DO_SRAM10(fabric_sram6_do_i[10]),
        .Tile_X11Y14_DO_SRAM11(fabric_sram6_do_i[11]),
        .Tile_X11Y14_DO_SRAM12(fabric_sram6_do_i[12]),
        .Tile_X11Y14_DO_SRAM13(fabric_sram6_do_i[13]),
        .Tile_X11Y14_DO_SRAM14(fabric_sram6_do_i[14]),
        .Tile_X11Y14_DO_SRAM15(fabric_sram6_do_i[15]),
        .Tile_X11Y14_DO_SRAM16(fabric_sram6_do_i[16]),
        .Tile_X11Y14_DO_SRAM17(fabric_sram6_do_i[17]),
        .Tile_X11Y14_DO_SRAM18(fabric_sram6_do_i[18]),
        .Tile_X11Y14_DO_SRAM19(fabric_sram6_do_i[19]),
        .Tile_X11Y14_DO_SRAM20(fabric_sram6_do_i[20]),
        .Tile_X11Y14_DO_SRAM21(fabric_sram6_do_i[21]),
        .Tile_X11Y14_DO_SRAM22(fabric_sram6_do_i[22]),
        .Tile_X11Y14_DO_SRAM23(fabric_sram6_do_i[23]),
        .Tile_X11Y14_DO_SRAM24(fabric_sram6_do_i[24]),
        .Tile_X11Y14_DO_SRAM25(fabric_sram6_do_i[25]),
        .Tile_X11Y14_DO_SRAM26(fabric_sram6_do_i[26]),
        .Tile_X11Y14_DO_SRAM27(fabric_sram6_do_i[27]),
        .Tile_X11Y14_DO_SRAM28(fabric_sram6_do_i[28]),
        .Tile_X11Y14_DO_SRAM29(fabric_sram6_do_i[29]),
        .Tile_X11Y14_DO_SRAM30(fabric_sram6_do_i[30]),
        .Tile_X11Y14_DO_SRAM31(fabric_sram6_do_i[31]),
        .Tile_X11Y14_AD_SRAM0(fabric_sram6_ad_o[0]),
        .Tile_X11Y14_AD_SRAM1(fabric_sram6_ad_o[1]),
        .Tile_X11Y14_AD_SRAM2(fabric_sram6_ad_o[2]),
        .Tile_X11Y14_AD_SRAM3(fabric_sram6_ad_o[3]),
        .Tile_X11Y14_AD_SRAM4(fabric_sram6_ad_o[4]),
        .Tile_X11Y14_AD_SRAM5(fabric_sram6_ad_o[5]),
        .Tile_X11Y14_AD_SRAM6(fabric_sram6_ad_o[6]),
        .Tile_X11Y14_AD_SRAM7(fabric_sram6_ad_o[7]),
        .Tile_X11Y14_AD_SRAM8(fabric_sram6_ad_o[8]),
        .Tile_X11Y14_AD_SRAM9(fabric_sram6_ad_o[9]),
        .Tile_X11Y14_BEN_SRAM0(fabric_sram6_ben_o[0]),
        .Tile_X11Y14_BEN_SRAM1(fabric_sram6_ben_o[1]),
        .Tile_X11Y14_BEN_SRAM2(fabric_sram6_ben_o[2]),
        .Tile_X11Y14_BEN_SRAM3(fabric_sram6_ben_o[3]),
        .Tile_X11Y14_BEN_SRAM4(fabric_sram6_ben_o[4]),
        .Tile_X11Y14_BEN_SRAM5(fabric_sram6_ben_o[5]),
        .Tile_X11Y14_BEN_SRAM6(fabric_sram6_ben_o[6]),
        .Tile_X11Y14_BEN_SRAM7(fabric_sram6_ben_o[7]),
        .Tile_X11Y14_BEN_SRAM8(fabric_sram6_ben_o[8]),
        .Tile_X11Y14_BEN_SRAM9(fabric_sram6_ben_o[9]),
        .Tile_X11Y14_BEN_SRAM10(fabric_sram6_ben_o[10]),
        .Tile_X11Y14_BEN_SRAM11(fabric_sram6_ben_o[11]),
        .Tile_X11Y14_BEN_SRAM12(fabric_sram6_ben_o[12]),
        .Tile_X11Y14_BEN_SRAM13(fabric_sram6_ben_o[13]),
        .Tile_X11Y14_BEN_SRAM14(fabric_sram6_ben_o[14]),
        .Tile_X11Y14_BEN_SRAM15(fabric_sram6_ben_o[15]),
        .Tile_X11Y14_BEN_SRAM16(fabric_sram6_ben_o[16]),
        .Tile_X11Y14_BEN_SRAM17(fabric_sram6_ben_o[17]),
        .Tile_X11Y14_BEN_SRAM18(fabric_sram6_ben_o[18]),
        .Tile_X11Y14_BEN_SRAM19(fabric_sram6_ben_o[19]),
        .Tile_X11Y14_BEN_SRAM20(fabric_sram6_ben_o[20]),
        .Tile_X11Y14_BEN_SRAM21(fabric_sram6_ben_o[21]),
        .Tile_X11Y14_BEN_SRAM22(fabric_sram6_ben_o[22]),
        .Tile_X11Y14_BEN_SRAM23(fabric_sram6_ben_o[23]),
        .Tile_X11Y14_BEN_SRAM24(fabric_sram6_ben_o[24]),
        .Tile_X11Y14_BEN_SRAM25(fabric_sram6_ben_o[25]),
        .Tile_X11Y14_BEN_SRAM26(fabric_sram6_ben_o[26]),
        .Tile_X11Y14_BEN_SRAM27(fabric_sram6_ben_o[27]),
        .Tile_X11Y14_BEN_SRAM28(fabric_sram6_ben_o[28]),
        .Tile_X11Y14_BEN_SRAM29(fabric_sram6_ben_o[29]),
        .Tile_X11Y14_BEN_SRAM30(fabric_sram6_ben_o[30]),
        .Tile_X11Y14_BEN_SRAM31(fabric_sram6_ben_o[31]),
        .Tile_X11Y14_DI_SRAM0(fabric_sram6_di_o[0]),
        .Tile_X11Y14_DI_SRAM1(fabric_sram6_di_o[1]),
        .Tile_X11Y14_DI_SRAM2(fabric_sram6_di_o[2]),
        .Tile_X11Y14_DI_SRAM3(fabric_sram6_di_o[3]),
        .Tile_X11Y14_DI_SRAM4(fabric_sram6_di_o[4]),
        .Tile_X11Y14_DI_SRAM5(fabric_sram6_di_o[5]),
        .Tile_X11Y14_DI_SRAM6(fabric_sram6_di_o[6]),
        .Tile_X11Y14_DI_SRAM7(fabric_sram6_di_o[7]),
        .Tile_X11Y14_DI_SRAM8(fabric_sram6_di_o[8]),
        .Tile_X11Y14_DI_SRAM9(fabric_sram6_di_o[9]),
        .Tile_X11Y14_DI_SRAM10(fabric_sram6_di_o[10]),
        .Tile_X11Y14_DI_SRAM11(fabric_sram6_di_o[11]),
        .Tile_X11Y14_DI_SRAM12(fabric_sram6_di_o[12]),
        .Tile_X11Y14_DI_SRAM13(fabric_sram6_di_o[13]),
        .Tile_X11Y14_DI_SRAM14(fabric_sram6_di_o[14]),
        .Tile_X11Y14_DI_SRAM15(fabric_sram6_di_o[15]),
        .Tile_X11Y14_DI_SRAM16(fabric_sram6_di_o[16]),
        .Tile_X11Y14_DI_SRAM17(fabric_sram6_di_o[17]),
        .Tile_X11Y14_DI_SRAM18(fabric_sram6_di_o[18]),
        .Tile_X11Y14_DI_SRAM19(fabric_sram6_di_o[19]),
        .Tile_X11Y14_DI_SRAM20(fabric_sram6_di_o[20]),
        .Tile_X11Y14_DI_SRAM21(fabric_sram6_di_o[21]),
        .Tile_X11Y14_DI_SRAM22(fabric_sram6_di_o[22]),
        .Tile_X11Y14_DI_SRAM23(fabric_sram6_di_o[23]),
        .Tile_X11Y14_DI_SRAM24(fabric_sram6_di_o[24]),
        .Tile_X11Y14_DI_SRAM25(fabric_sram6_di_o[25]),
        .Tile_X11Y14_DI_SRAM26(fabric_sram6_di_o[26]),
        .Tile_X11Y14_DI_SRAM27(fabric_sram6_di_o[27]),
        .Tile_X11Y14_DI_SRAM28(fabric_sram6_di_o[28]),
        .Tile_X11Y14_DI_SRAM29(fabric_sram6_di_o[29]),
        .Tile_X11Y14_DI_SRAM30(fabric_sram6_di_o[30]),
        .Tile_X11Y14_DI_SRAM31(fabric_sram6_di_o[31]),
        .Tile_X11Y14_EN_SRAM(fabric_sram6_en),
        .Tile_X11Y14_R_WB_SRAM(fabric_sram6_rw_no),
        .Tile_X11Y14_CLOCK_SRAM(fabric_sram6_clk_o),

        // SRAM 7
        .Tile_X11Y16_DO_SRAM0(fabric_sram7_do_i[0]),
        .Tile_X11Y16_DO_SRAM1(fabric_sram7_do_i[1]),
        .Tile_X11Y16_DO_SRAM2(fabric_sram7_do_i[2]),
        .Tile_X11Y16_DO_SRAM3(fabric_sram7_do_i[3]),
        .Tile_X11Y16_DO_SRAM4(fabric_sram7_do_i[4]),
        .Tile_X11Y16_DO_SRAM5(fabric_sram7_do_i[5]),
        .Tile_X11Y16_DO_SRAM6(fabric_sram7_do_i[6]),
        .Tile_X11Y16_DO_SRAM7(fabric_sram7_do_i[7]),
        .Tile_X11Y16_DO_SRAM8(fabric_sram7_do_i[8]),
        .Tile_X11Y16_DO_SRAM9(fabric_sram7_do_i[9]),
        .Tile_X11Y16_DO_SRAM10(fabric_sram7_do_i[10]),
        .Tile_X11Y16_DO_SRAM11(fabric_sram7_do_i[11]),
        .Tile_X11Y16_DO_SRAM12(fabric_sram7_do_i[12]),
        .Tile_X11Y16_DO_SRAM13(fabric_sram7_do_i[13]),
        .Tile_X11Y16_DO_SRAM14(fabric_sram7_do_i[14]),
        .Tile_X11Y16_DO_SRAM15(fabric_sram7_do_i[15]),
        .Tile_X11Y16_DO_SRAM16(fabric_sram7_do_i[16]),
        .Tile_X11Y16_DO_SRAM17(fabric_sram7_do_i[17]),
        .Tile_X11Y16_DO_SRAM18(fabric_sram7_do_i[18]),
        .Tile_X11Y16_DO_SRAM19(fabric_sram7_do_i[19]),
        .Tile_X11Y16_DO_SRAM20(fabric_sram7_do_i[20]),
        .Tile_X11Y16_DO_SRAM21(fabric_sram7_do_i[21]),
        .Tile_X11Y16_DO_SRAM22(fabric_sram7_do_i[22]),
        .Tile_X11Y16_DO_SRAM23(fabric_sram7_do_i[23]),
        .Tile_X11Y16_DO_SRAM24(fabric_sram7_do_i[24]),
        .Tile_X11Y16_DO_SRAM25(fabric_sram7_do_i[25]),
        .Tile_X11Y16_DO_SRAM26(fabric_sram7_do_i[26]),
        .Tile_X11Y16_DO_SRAM27(fabric_sram7_do_i[27]),
        .Tile_X11Y16_DO_SRAM28(fabric_sram7_do_i[28]),
        .Tile_X11Y16_DO_SRAM29(fabric_sram7_do_i[29]),
        .Tile_X11Y16_DO_SRAM30(fabric_sram7_do_i[30]),
        .Tile_X11Y16_DO_SRAM31(fabric_sram7_do_i[31]),
        .Tile_X11Y16_AD_SRAM0(fabric_sram7_ad_o[0]),
        .Tile_X11Y16_AD_SRAM1(fabric_sram7_ad_o[1]),
        .Tile_X11Y16_AD_SRAM2(fabric_sram7_ad_o[2]),
        .Tile_X11Y16_AD_SRAM3(fabric_sram7_ad_o[3]),
        .Tile_X11Y16_AD_SRAM4(fabric_sram7_ad_o[4]),
        .Tile_X11Y16_AD_SRAM5(fabric_sram7_ad_o[5]),
        .Tile_X11Y16_AD_SRAM6(fabric_sram7_ad_o[6]),
        .Tile_X11Y16_AD_SRAM7(fabric_sram7_ad_o[7]),
        .Tile_X11Y16_AD_SRAM8(fabric_sram7_ad_o[8]),
        .Tile_X11Y16_AD_SRAM9(fabric_sram7_ad_o[9]),
        .Tile_X11Y16_BEN_SRAM0(fabric_sram7_ben_o[0]),
        .Tile_X11Y16_BEN_SRAM1(fabric_sram7_ben_o[1]),
        .Tile_X11Y16_BEN_SRAM2(fabric_sram7_ben_o[2]),
        .Tile_X11Y16_BEN_SRAM3(fabric_sram7_ben_o[3]),
        .Tile_X11Y16_BEN_SRAM4(fabric_sram7_ben_o[4]),
        .Tile_X11Y16_BEN_SRAM5(fabric_sram7_ben_o[5]),
        .Tile_X11Y16_BEN_SRAM6(fabric_sram7_ben_o[6]),
        .Tile_X11Y16_BEN_SRAM7(fabric_sram7_ben_o[7]),
        .Tile_X11Y16_BEN_SRAM8(fabric_sram7_ben_o[8]),
        .Tile_X11Y16_BEN_SRAM9(fabric_sram7_ben_o[9]),
        .Tile_X11Y16_BEN_SRAM10(fabric_sram7_ben_o[10]),
        .Tile_X11Y16_BEN_SRAM11(fabric_sram7_ben_o[11]),
        .Tile_X11Y16_BEN_SRAM12(fabric_sram7_ben_o[12]),
        .Tile_X11Y16_BEN_SRAM13(fabric_sram7_ben_o[13]),
        .Tile_X11Y16_BEN_SRAM14(fabric_sram7_ben_o[14]),
        .Tile_X11Y16_BEN_SRAM15(fabric_sram7_ben_o[15]),
        .Tile_X11Y16_BEN_SRAM16(fabric_sram7_ben_o[16]),
        .Tile_X11Y16_BEN_SRAM17(fabric_sram7_ben_o[17]),
        .Tile_X11Y16_BEN_SRAM18(fabric_sram7_ben_o[18]),
        .Tile_X11Y16_BEN_SRAM19(fabric_sram7_ben_o[19]),
        .Tile_X11Y16_BEN_SRAM20(fabric_sram7_ben_o[20]),
        .Tile_X11Y16_BEN_SRAM21(fabric_sram7_ben_o[21]),
        .Tile_X11Y16_BEN_SRAM22(fabric_sram7_ben_o[22]),
        .Tile_X11Y16_BEN_SRAM23(fabric_sram7_ben_o[23]),
        .Tile_X11Y16_BEN_SRAM24(fabric_sram7_ben_o[24]),
        .Tile_X11Y16_BEN_SRAM25(fabric_sram7_ben_o[25]),
        .Tile_X11Y16_BEN_SRAM26(fabric_sram7_ben_o[26]),
        .Tile_X11Y16_BEN_SRAM27(fabric_sram7_ben_o[27]),
        .Tile_X11Y16_BEN_SRAM28(fabric_sram7_ben_o[28]),
        .Tile_X11Y16_BEN_SRAM29(fabric_sram7_ben_o[29]),
        .Tile_X11Y16_BEN_SRAM30(fabric_sram7_ben_o[30]),
        .Tile_X11Y16_BEN_SRAM31(fabric_sram7_ben_o[31]),
        .Tile_X11Y16_DI_SRAM0(fabric_sram7_di_o[0]),
        .Tile_X11Y16_DI_SRAM1(fabric_sram7_di_o[1]),
        .Tile_X11Y16_DI_SRAM2(fabric_sram7_di_o[2]),
        .Tile_X11Y16_DI_SRAM3(fabric_sram7_di_o[3]),
        .Tile_X11Y16_DI_SRAM4(fabric_sram7_di_o[4]),
        .Tile_X11Y16_DI_SRAM5(fabric_sram7_di_o[5]),
        .Tile_X11Y16_DI_SRAM6(fabric_sram7_di_o[6]),
        .Tile_X11Y16_DI_SRAM7(fabric_sram7_di_o[7]),
        .Tile_X11Y16_DI_SRAM8(fabric_sram7_di_o[8]),
        .Tile_X11Y16_DI_SRAM9(fabric_sram7_di_o[9]),
        .Tile_X11Y16_DI_SRAM10(fabric_sram7_di_o[10]),
        .Tile_X11Y16_DI_SRAM11(fabric_sram7_di_o[11]),
        .Tile_X11Y16_DI_SRAM12(fabric_sram7_di_o[12]),
        .Tile_X11Y16_DI_SRAM13(fabric_sram7_di_o[13]),
        .Tile_X11Y16_DI_SRAM14(fabric_sram7_di_o[14]),
        .Tile_X11Y16_DI_SRAM15(fabric_sram7_di_o[15]),
        .Tile_X11Y16_DI_SRAM16(fabric_sram7_di_o[16]),
        .Tile_X11Y16_DI_SRAM17(fabric_sram7_di_o[17]),
        .Tile_X11Y16_DI_SRAM18(fabric_sram7_di_o[18]),
        .Tile_X11Y16_DI_SRAM19(fabric_sram7_di_o[19]),
        .Tile_X11Y16_DI_SRAM20(fabric_sram7_di_o[20]),
        .Tile_X11Y16_DI_SRAM21(fabric_sram7_di_o[21]),
        .Tile_X11Y16_DI_SRAM22(fabric_sram7_di_o[22]),
        .Tile_X11Y16_DI_SRAM23(fabric_sram7_di_o[23]),
        .Tile_X11Y16_DI_SRAM24(fabric_sram7_di_o[24]),
        .Tile_X11Y16_DI_SRAM25(fabric_sram7_di_o[25]),
        .Tile_X11Y16_DI_SRAM26(fabric_sram7_di_o[26]),
        .Tile_X11Y16_DI_SRAM27(fabric_sram7_di_o[27]),
        .Tile_X11Y16_DI_SRAM28(fabric_sram7_di_o[28]),
        .Tile_X11Y16_DI_SRAM29(fabric_sram7_di_o[29]),
        .Tile_X11Y16_DI_SRAM30(fabric_sram7_di_o[30]),
        .Tile_X11Y16_DI_SRAM31(fabric_sram7_di_o[31]),
        .Tile_X11Y16_EN_SRAM(fabric_sram7_en),
        .Tile_X11Y16_R_WB_SRAM(fabric_sram7_rw_no),
        .Tile_X11Y16_CLOCK_SRAM(fabric_sram7_clk_o),

        // WARMBOOT
        .Tile_X2Y17_RESET_top(fabric_warmboot_reset_i),
        .Tile_X2Y17_BOOT_top(fabric_warmboot_boot),
        .Tile_X2Y17_SLOT_top0(fabric_warmboot_slot_o[0]),
        .Tile_X2Y17_SLOT_top1(fabric_warmboot_slot_o[1]),
        .Tile_X2Y17_SLOT_top2(fabric_warmboot_slot_o[2]),
        .Tile_X2Y17_SLOT_top3(fabric_warmboot_slot_o[3]),

        // IRQ
        .Tile_X1Y17_IRQ_top0(fabric_irq[0]),
        .Tile_X1Y17_IRQ_top1(fabric_irq[1]),
        .Tile_X1Y17_IRQ_top2(fabric_irq[2]),
        .Tile_X1Y17_IRQ_top3(fabric_irq[3]),

        // CPU_IF 0
        .Tile_X4Y17_I_top0(fabric_cpu_o[0]),
        .Tile_X4Y17_I_top1(fabric_cpu_o[1]),
        .Tile_X4Y17_I_top2(fabric_cpu_o[2]),
        .Tile_X4Y17_I_top3(fabric_cpu_o[3]),
        .Tile_X4Y17_I_top4(fabric_cpu_o[4]),
        .Tile_X4Y17_I_top5(fabric_cpu_o[5]),
        .Tile_X4Y17_I_top6(fabric_cpu_o[6]),
        .Tile_X4Y17_I_top7(fabric_cpu_o[7]),
        .Tile_X4Y17_I_top8(fabric_cpu_o[8]),
        .Tile_X4Y17_I_top9(fabric_cpu_o[9]),
        .Tile_X4Y17_I_top10(fabric_cpu_o[10]),
        .Tile_X4Y17_I_top11(fabric_cpu_o[11]),
        .Tile_X4Y17_I_top12(fabric_cpu_o[12]),
        .Tile_X4Y17_I_top13(fabric_cpu_o[13]),
        .Tile_X4Y17_I_top14(fabric_cpu_o[14]),
        .Tile_X4Y17_I_top15(fabric_cpu_o[15]),
        .Tile_X4Y17_O_top0(fabric_cpu_i[0]),
        .Tile_X4Y17_O_top1(fabric_cpu_i[1]),
        .Tile_X4Y17_O_top2(fabric_cpu_i[2]),
        .Tile_X4Y17_O_top3(fabric_cpu_i[3]),
        .Tile_X4Y17_O_top4(fabric_cpu_i[4]),
        .Tile_X4Y17_O_top5(fabric_cpu_i[5]),
        .Tile_X4Y17_O_top6(fabric_cpu_i[6]),
        .Tile_X4Y17_O_top7(fabric_cpu_i[7]),
        .Tile_X4Y17_O_top8(fabric_cpu_i[8]),
        .Tile_X4Y17_O_top9(fabric_cpu_i[9]),
        .Tile_X4Y17_O_top10(fabric_cpu_i[10]),
        .Tile_X4Y17_O_top11(fabric_cpu_i[11]),
        .Tile_X4Y17_O_top12(fabric_cpu_i[12]),
        .Tile_X4Y17_O_top13(fabric_cpu_i[13]),
        .Tile_X4Y17_O_top14(fabric_cpu_i[14]),
        .Tile_X4Y17_O_top15(fabric_cpu_i[15]),

        // CPU_IF 1
        .Tile_X5Y17_I_top0(fabric_cpu_o[16]),
        .Tile_X5Y17_I_top1(fabric_cpu_o[17]),
        .Tile_X5Y17_I_top2(fabric_cpu_o[18]),
        .Tile_X5Y17_I_top3(fabric_cpu_o[19]),
        .Tile_X5Y17_I_top4(fabric_cpu_o[20]),
        .Tile_X5Y17_I_top5(fabric_cpu_o[21]),
        .Tile_X5Y17_I_top6(fabric_cpu_o[22]),
        .Tile_X5Y17_I_top7(fabric_cpu_o[23]),
        .Tile_X5Y17_I_top8(fabric_cpu_o[24]),
        .Tile_X5Y17_I_top9(fabric_cpu_o[25]),
        .Tile_X5Y17_I_top10(fabric_cpu_o[26]),
        .Tile_X5Y17_I_top11(fabric_cpu_o[27]),
        .Tile_X5Y17_I_top12(fabric_cpu_o[28]),
        .Tile_X5Y17_I_top13(fabric_cpu_o[29]),
        .Tile_X5Y17_I_top14(fabric_cpu_o[30]),
        .Tile_X5Y17_I_top15(fabric_cpu_o[31]),
        .Tile_X5Y17_O_top0(fabric_cpu_i[16]),
        .Tile_X5Y17_O_top1(fabric_cpu_i[17]),
        .Tile_X5Y17_O_top2(fabric_cpu_i[18]),
        .Tile_X5Y17_O_top3(fabric_cpu_i[19]),
        .Tile_X5Y17_O_top4(fabric_cpu_i[20]),
        .Tile_X5Y17_O_top5(fabric_cpu_i[21]),
        .Tile_X5Y17_O_top6(fabric_cpu_i[22]),
        .Tile_X5Y17_O_top7(fabric_cpu_i[23]),
        .Tile_X5Y17_O_top8(fabric_cpu_i[24]),
        .Tile_X5Y17_O_top9(fabric_cpu_i[25]),
        .Tile_X5Y17_O_top10(fabric_cpu_i[26]),
        .Tile_X5Y17_O_top11(fabric_cpu_i[27]),
        .Tile_X5Y17_O_top12(fabric_cpu_i[28]),
        .Tile_X5Y17_O_top13(fabric_cpu_i[29]),
        .Tile_X5Y17_O_top14(fabric_cpu_i[30]),
        .Tile_X5Y17_O_top15(fabric_cpu_i[31]),

        // CPU_IF 2
        .Tile_X6Y17_I_top0(fabric_cpu_o[32]),
        .Tile_X6Y17_I_top1(fabric_cpu_o[33]),
        .Tile_X6Y17_I_top2(fabric_cpu_o[34]),
        .Tile_X6Y17_I_top3(fabric_cpu_o[35]),
        .Tile_X6Y17_I_top4(fabric_cpu_o[36]),
        .Tile_X6Y17_I_top5(fabric_cpu_o[37]),
        .Tile_X6Y17_I_top6(fabric_cpu_o[38]),
        .Tile_X6Y17_I_top7(fabric_cpu_o[39]),
        .Tile_X6Y17_I_top8(fabric_cpu_o[40]),
        .Tile_X6Y17_I_top9(fabric_cpu_o[41]),
        .Tile_X6Y17_I_top10(fabric_cpu_o[42]),
        .Tile_X6Y17_I_top11(fabric_cpu_o[43]),
        .Tile_X6Y17_I_top12(fabric_cpu_o[44]),
        .Tile_X6Y17_I_top13(fabric_cpu_o[45]),
        .Tile_X6Y17_I_top14(fabric_cpu_o[46]),
        .Tile_X6Y17_I_top15(fabric_cpu_o[47]),
        .Tile_X6Y17_O_top0(fabric_cpu_i[32]),
        .Tile_X6Y17_O_top1(fabric_cpu_i[33]),
        .Tile_X6Y17_O_top2(fabric_cpu_i[34]),
        .Tile_X6Y17_O_top3(fabric_cpu_i[35]),
        .Tile_X6Y17_O_top4(fabric_cpu_i[36]),
        .Tile_X6Y17_O_top5(fabric_cpu_i[37]),
        .Tile_X6Y17_O_top6(fabric_cpu_i[38]),
        .Tile_X6Y17_O_top7(fabric_cpu_i[39]),
        .Tile_X6Y17_O_top8(fabric_cpu_i[40]),
        .Tile_X6Y17_O_top9(fabric_cpu_i[41]),
        .Tile_X6Y17_O_top10(fabric_cpu_i[42]),
        .Tile_X6Y17_O_top11(fabric_cpu_i[43]),
        .Tile_X6Y17_O_top12(fabric_cpu_i[44]),
        .Tile_X6Y17_O_top13(fabric_cpu_i[45]),
        .Tile_X6Y17_O_top14(fabric_cpu_i[46]),
        .Tile_X6Y17_O_top15(fabric_cpu_i[47]),

        // CPU_IF 3
        .Tile_X8Y17_I_top0(fabric_cpu_o[48]),
        .Tile_X8Y17_I_top1(fabric_cpu_o[49]),
        .Tile_X8Y17_I_top2(fabric_cpu_o[50]),
        .Tile_X8Y17_I_top3(fabric_cpu_o[51]),
        .Tile_X8Y17_I_top4(fabric_cpu_o[52]),
        .Tile_X8Y17_I_top5(fabric_cpu_o[53]),
        .Tile_X8Y17_I_top6(fabric_cpu_o[54]),
        .Tile_X8Y17_I_top7(fabric_cpu_o[55]),
        .Tile_X8Y17_I_top8(fabric_cpu_o[56]),
        .Tile_X8Y17_I_top9(fabric_cpu_o[57]),
        .Tile_X8Y17_I_top10(fabric_cpu_o[58]),
        .Tile_X8Y17_I_top11(fabric_cpu_o[59]),
        .Tile_X8Y17_I_top12(fabric_cpu_o[60]),
        .Tile_X8Y17_I_top13(fabric_cpu_o[61]),
        .Tile_X8Y17_I_top14(fabric_cpu_o[62]),
        .Tile_X8Y17_I_top15(fabric_cpu_o[63]),
        .Tile_X8Y17_O_top0(fabric_cpu_i[48]),
        .Tile_X8Y17_O_top1(fabric_cpu_i[49]),
        .Tile_X8Y17_O_top2(fabric_cpu_i[50]),
        .Tile_X8Y17_O_top3(fabric_cpu_i[51]),
        .Tile_X8Y17_O_top4(fabric_cpu_i[52]),
        .Tile_X8Y17_O_top5(fabric_cpu_i[53]),
        .Tile_X8Y17_O_top6(fabric_cpu_i[54]),
        .Tile_X8Y17_O_top7(fabric_cpu_i[55]),
        .Tile_X8Y17_O_top8(fabric_cpu_i[56]),
        .Tile_X8Y17_O_top9(fabric_cpu_i[57]),
        .Tile_X8Y17_O_top10(fabric_cpu_i[58]),
        .Tile_X8Y17_O_top11(fabric_cpu_i[59]),
        .Tile_X8Y17_O_top12(fabric_cpu_i[60]),
        .Tile_X8Y17_O_top13(fabric_cpu_i[61]),
        .Tile_X8Y17_O_top14(fabric_cpu_i[62]),
        .Tile_X8Y17_O_top15(fabric_cpu_i[63])
    );

endmodule

`default_nettype wire
