module eFPGA (Tile_X0Y10_A_I_top,
    Tile_X0Y10_A_O_top,
    Tile_X0Y10_A_T_top,
    Tile_X0Y10_A_config_C_bit0,
    Tile_X0Y10_A_config_C_bit1,
    Tile_X0Y10_A_config_C_bit2,
    Tile_X0Y10_A_config_C_bit3,
    Tile_X0Y10_B_I_top,
    Tile_X0Y10_B_O_top,
    Tile_X0Y10_B_T_top,
    Tile_X0Y10_B_config_C_bit0,
    Tile_X0Y10_B_config_C_bit1,
    Tile_X0Y10_B_config_C_bit2,
    Tile_X0Y10_B_config_C_bit3,
    Tile_X0Y11_A_I_top,
    Tile_X0Y11_A_O_top,
    Tile_X0Y11_A_T_top,
    Tile_X0Y11_A_config_C_bit0,
    Tile_X0Y11_A_config_C_bit1,
    Tile_X0Y11_A_config_C_bit2,
    Tile_X0Y11_A_config_C_bit3,
    Tile_X0Y11_B_I_top,
    Tile_X0Y11_B_O_top,
    Tile_X0Y11_B_T_top,
    Tile_X0Y11_B_config_C_bit0,
    Tile_X0Y11_B_config_C_bit1,
    Tile_X0Y11_B_config_C_bit2,
    Tile_X0Y11_B_config_C_bit3,
    Tile_X0Y12_A_I_top,
    Tile_X0Y12_A_O_top,
    Tile_X0Y12_A_T_top,
    Tile_X0Y12_A_config_C_bit0,
    Tile_X0Y12_A_config_C_bit1,
    Tile_X0Y12_A_config_C_bit2,
    Tile_X0Y12_A_config_C_bit3,
    Tile_X0Y12_B_I_top,
    Tile_X0Y12_B_O_top,
    Tile_X0Y12_B_T_top,
    Tile_X0Y12_B_config_C_bit0,
    Tile_X0Y12_B_config_C_bit1,
    Tile_X0Y12_B_config_C_bit2,
    Tile_X0Y12_B_config_C_bit3,
    Tile_X0Y13_A_I_top,
    Tile_X0Y13_A_O_top,
    Tile_X0Y13_A_T_top,
    Tile_X0Y13_A_config_C_bit0,
    Tile_X0Y13_A_config_C_bit1,
    Tile_X0Y13_A_config_C_bit2,
    Tile_X0Y13_A_config_C_bit3,
    Tile_X0Y13_B_I_top,
    Tile_X0Y13_B_O_top,
    Tile_X0Y13_B_T_top,
    Tile_X0Y13_B_config_C_bit0,
    Tile_X0Y13_B_config_C_bit1,
    Tile_X0Y13_B_config_C_bit2,
    Tile_X0Y13_B_config_C_bit3,
    Tile_X0Y14_A_I_top,
    Tile_X0Y14_A_O_top,
    Tile_X0Y14_A_T_top,
    Tile_X0Y14_A_config_C_bit0,
    Tile_X0Y14_A_config_C_bit1,
    Tile_X0Y14_A_config_C_bit2,
    Tile_X0Y14_A_config_C_bit3,
    Tile_X0Y14_B_I_top,
    Tile_X0Y14_B_O_top,
    Tile_X0Y14_B_T_top,
    Tile_X0Y14_B_config_C_bit0,
    Tile_X0Y14_B_config_C_bit1,
    Tile_X0Y14_B_config_C_bit2,
    Tile_X0Y14_B_config_C_bit3,
    Tile_X0Y1_A_I_top,
    Tile_X0Y1_A_O_top,
    Tile_X0Y1_A_T_top,
    Tile_X0Y1_A_config_C_bit0,
    Tile_X0Y1_A_config_C_bit1,
    Tile_X0Y1_A_config_C_bit2,
    Tile_X0Y1_A_config_C_bit3,
    Tile_X0Y1_B_I_top,
    Tile_X0Y1_B_O_top,
    Tile_X0Y1_B_T_top,
    Tile_X0Y1_B_config_C_bit0,
    Tile_X0Y1_B_config_C_bit1,
    Tile_X0Y1_B_config_C_bit2,
    Tile_X0Y1_B_config_C_bit3,
    Tile_X0Y2_A_I_top,
    Tile_X0Y2_A_O_top,
    Tile_X0Y2_A_T_top,
    Tile_X0Y2_A_config_C_bit0,
    Tile_X0Y2_A_config_C_bit1,
    Tile_X0Y2_A_config_C_bit2,
    Tile_X0Y2_A_config_C_bit3,
    Tile_X0Y2_B_I_top,
    Tile_X0Y2_B_O_top,
    Tile_X0Y2_B_T_top,
    Tile_X0Y2_B_config_C_bit0,
    Tile_X0Y2_B_config_C_bit1,
    Tile_X0Y2_B_config_C_bit2,
    Tile_X0Y2_B_config_C_bit3,
    Tile_X0Y3_A_I_top,
    Tile_X0Y3_A_O_top,
    Tile_X0Y3_A_T_top,
    Tile_X0Y3_A_config_C_bit0,
    Tile_X0Y3_A_config_C_bit1,
    Tile_X0Y3_A_config_C_bit2,
    Tile_X0Y3_A_config_C_bit3,
    Tile_X0Y3_B_I_top,
    Tile_X0Y3_B_O_top,
    Tile_X0Y3_B_T_top,
    Tile_X0Y3_B_config_C_bit0,
    Tile_X0Y3_B_config_C_bit1,
    Tile_X0Y3_B_config_C_bit2,
    Tile_X0Y3_B_config_C_bit3,
    Tile_X0Y4_A_I_top,
    Tile_X0Y4_A_O_top,
    Tile_X0Y4_A_T_top,
    Tile_X0Y4_A_config_C_bit0,
    Tile_X0Y4_A_config_C_bit1,
    Tile_X0Y4_A_config_C_bit2,
    Tile_X0Y4_A_config_C_bit3,
    Tile_X0Y4_B_I_top,
    Tile_X0Y4_B_O_top,
    Tile_X0Y4_B_T_top,
    Tile_X0Y4_B_config_C_bit0,
    Tile_X0Y4_B_config_C_bit1,
    Tile_X0Y4_B_config_C_bit2,
    Tile_X0Y4_B_config_C_bit3,
    Tile_X0Y5_A_I_top,
    Tile_X0Y5_A_O_top,
    Tile_X0Y5_A_T_top,
    Tile_X0Y5_A_config_C_bit0,
    Tile_X0Y5_A_config_C_bit1,
    Tile_X0Y5_A_config_C_bit2,
    Tile_X0Y5_A_config_C_bit3,
    Tile_X0Y5_B_I_top,
    Tile_X0Y5_B_O_top,
    Tile_X0Y5_B_T_top,
    Tile_X0Y5_B_config_C_bit0,
    Tile_X0Y5_B_config_C_bit1,
    Tile_X0Y5_B_config_C_bit2,
    Tile_X0Y5_B_config_C_bit3,
    Tile_X0Y6_A_I_top,
    Tile_X0Y6_A_O_top,
    Tile_X0Y6_A_T_top,
    Tile_X0Y6_A_config_C_bit0,
    Tile_X0Y6_A_config_C_bit1,
    Tile_X0Y6_A_config_C_bit2,
    Tile_X0Y6_A_config_C_bit3,
    Tile_X0Y6_B_I_top,
    Tile_X0Y6_B_O_top,
    Tile_X0Y6_B_T_top,
    Tile_X0Y6_B_config_C_bit0,
    Tile_X0Y6_B_config_C_bit1,
    Tile_X0Y6_B_config_C_bit2,
    Tile_X0Y6_B_config_C_bit3,
    Tile_X0Y7_A_I_top,
    Tile_X0Y7_A_O_top,
    Tile_X0Y7_A_T_top,
    Tile_X0Y7_A_config_C_bit0,
    Tile_X0Y7_A_config_C_bit1,
    Tile_X0Y7_A_config_C_bit2,
    Tile_X0Y7_A_config_C_bit3,
    Tile_X0Y7_B_I_top,
    Tile_X0Y7_B_O_top,
    Tile_X0Y7_B_T_top,
    Tile_X0Y7_B_config_C_bit0,
    Tile_X0Y7_B_config_C_bit1,
    Tile_X0Y7_B_config_C_bit2,
    Tile_X0Y7_B_config_C_bit3,
    Tile_X0Y8_A_I_top,
    Tile_X0Y8_A_O_top,
    Tile_X0Y8_A_T_top,
    Tile_X0Y8_A_config_C_bit0,
    Tile_X0Y8_A_config_C_bit1,
    Tile_X0Y8_A_config_C_bit2,
    Tile_X0Y8_A_config_C_bit3,
    Tile_X0Y8_B_I_top,
    Tile_X0Y8_B_O_top,
    Tile_X0Y8_B_T_top,
    Tile_X0Y8_B_config_C_bit0,
    Tile_X0Y8_B_config_C_bit1,
    Tile_X0Y8_B_config_C_bit2,
    Tile_X0Y8_B_config_C_bit3,
    Tile_X0Y9_A_I_top,
    Tile_X0Y9_A_O_top,
    Tile_X0Y9_A_T_top,
    Tile_X0Y9_A_config_C_bit0,
    Tile_X0Y9_A_config_C_bit1,
    Tile_X0Y9_A_config_C_bit2,
    Tile_X0Y9_A_config_C_bit3,
    Tile_X0Y9_B_I_top,
    Tile_X0Y9_B_O_top,
    Tile_X0Y9_B_T_top,
    Tile_X0Y9_B_config_C_bit0,
    Tile_X0Y9_B_config_C_bit1,
    Tile_X0Y9_B_config_C_bit2,
    Tile_X0Y9_B_config_C_bit3,
    Tile_X10Y10_ADDR_SRAM0,
    Tile_X10Y10_ADDR_SRAM1,
    Tile_X10Y10_ADDR_SRAM2,
    Tile_X10Y10_ADDR_SRAM3,
    Tile_X10Y10_ADDR_SRAM4,
    Tile_X10Y10_ADDR_SRAM5,
    Tile_X10Y10_ADDR_SRAM6,
    Tile_X10Y10_ADDR_SRAM7,
    Tile_X10Y10_ADDR_SRAM8,
    Tile_X10Y10_ADDR_SRAM9,
    Tile_X10Y10_BM_SRAM0,
    Tile_X10Y10_BM_SRAM1,
    Tile_X10Y10_BM_SRAM10,
    Tile_X10Y10_BM_SRAM11,
    Tile_X10Y10_BM_SRAM12,
    Tile_X10Y10_BM_SRAM13,
    Tile_X10Y10_BM_SRAM14,
    Tile_X10Y10_BM_SRAM15,
    Tile_X10Y10_BM_SRAM16,
    Tile_X10Y10_BM_SRAM17,
    Tile_X10Y10_BM_SRAM18,
    Tile_X10Y10_BM_SRAM19,
    Tile_X10Y10_BM_SRAM2,
    Tile_X10Y10_BM_SRAM20,
    Tile_X10Y10_BM_SRAM21,
    Tile_X10Y10_BM_SRAM22,
    Tile_X10Y10_BM_SRAM23,
    Tile_X10Y10_BM_SRAM24,
    Tile_X10Y10_BM_SRAM25,
    Tile_X10Y10_BM_SRAM26,
    Tile_X10Y10_BM_SRAM27,
    Tile_X10Y10_BM_SRAM28,
    Tile_X10Y10_BM_SRAM29,
    Tile_X10Y10_BM_SRAM3,
    Tile_X10Y10_BM_SRAM30,
    Tile_X10Y10_BM_SRAM31,
    Tile_X10Y10_BM_SRAM4,
    Tile_X10Y10_BM_SRAM5,
    Tile_X10Y10_BM_SRAM6,
    Tile_X10Y10_BM_SRAM7,
    Tile_X10Y10_BM_SRAM8,
    Tile_X10Y10_BM_SRAM9,
    Tile_X10Y10_CLK_SRAM,
    Tile_X10Y10_CONFIGURED_top,
    Tile_X10Y10_DIN_SRAM0,
    Tile_X10Y10_DIN_SRAM1,
    Tile_X10Y10_DIN_SRAM10,
    Tile_X10Y10_DIN_SRAM11,
    Tile_X10Y10_DIN_SRAM12,
    Tile_X10Y10_DIN_SRAM13,
    Tile_X10Y10_DIN_SRAM14,
    Tile_X10Y10_DIN_SRAM15,
    Tile_X10Y10_DIN_SRAM16,
    Tile_X10Y10_DIN_SRAM17,
    Tile_X10Y10_DIN_SRAM18,
    Tile_X10Y10_DIN_SRAM19,
    Tile_X10Y10_DIN_SRAM2,
    Tile_X10Y10_DIN_SRAM20,
    Tile_X10Y10_DIN_SRAM21,
    Tile_X10Y10_DIN_SRAM22,
    Tile_X10Y10_DIN_SRAM23,
    Tile_X10Y10_DIN_SRAM24,
    Tile_X10Y10_DIN_SRAM25,
    Tile_X10Y10_DIN_SRAM26,
    Tile_X10Y10_DIN_SRAM27,
    Tile_X10Y10_DIN_SRAM28,
    Tile_X10Y10_DIN_SRAM29,
    Tile_X10Y10_DIN_SRAM3,
    Tile_X10Y10_DIN_SRAM30,
    Tile_X10Y10_DIN_SRAM31,
    Tile_X10Y10_DIN_SRAM4,
    Tile_X10Y10_DIN_SRAM5,
    Tile_X10Y10_DIN_SRAM6,
    Tile_X10Y10_DIN_SRAM7,
    Tile_X10Y10_DIN_SRAM8,
    Tile_X10Y10_DIN_SRAM9,
    Tile_X10Y10_DOUT_SRAM0,
    Tile_X10Y10_DOUT_SRAM1,
    Tile_X10Y10_DOUT_SRAM10,
    Tile_X10Y10_DOUT_SRAM11,
    Tile_X10Y10_DOUT_SRAM12,
    Tile_X10Y10_DOUT_SRAM13,
    Tile_X10Y10_DOUT_SRAM14,
    Tile_X10Y10_DOUT_SRAM15,
    Tile_X10Y10_DOUT_SRAM16,
    Tile_X10Y10_DOUT_SRAM17,
    Tile_X10Y10_DOUT_SRAM18,
    Tile_X10Y10_DOUT_SRAM19,
    Tile_X10Y10_DOUT_SRAM2,
    Tile_X10Y10_DOUT_SRAM20,
    Tile_X10Y10_DOUT_SRAM21,
    Tile_X10Y10_DOUT_SRAM22,
    Tile_X10Y10_DOUT_SRAM23,
    Tile_X10Y10_DOUT_SRAM24,
    Tile_X10Y10_DOUT_SRAM25,
    Tile_X10Y10_DOUT_SRAM26,
    Tile_X10Y10_DOUT_SRAM27,
    Tile_X10Y10_DOUT_SRAM28,
    Tile_X10Y10_DOUT_SRAM29,
    Tile_X10Y10_DOUT_SRAM3,
    Tile_X10Y10_DOUT_SRAM30,
    Tile_X10Y10_DOUT_SRAM31,
    Tile_X10Y10_DOUT_SRAM4,
    Tile_X10Y10_DOUT_SRAM5,
    Tile_X10Y10_DOUT_SRAM6,
    Tile_X10Y10_DOUT_SRAM7,
    Tile_X10Y10_DOUT_SRAM8,
    Tile_X10Y10_DOUT_SRAM9,
    Tile_X10Y10_MEN_SRAM,
    Tile_X10Y10_REN_SRAM,
    Tile_X10Y10_TIE_HIGH_SRAM,
    Tile_X10Y10_TIE_LOW_SRAM,
    Tile_X10Y10_WEN_SRAM,
    Tile_X10Y12_ADDR_SRAM0,
    Tile_X10Y12_ADDR_SRAM1,
    Tile_X10Y12_ADDR_SRAM2,
    Tile_X10Y12_ADDR_SRAM3,
    Tile_X10Y12_ADDR_SRAM4,
    Tile_X10Y12_ADDR_SRAM5,
    Tile_X10Y12_ADDR_SRAM6,
    Tile_X10Y12_ADDR_SRAM7,
    Tile_X10Y12_ADDR_SRAM8,
    Tile_X10Y12_ADDR_SRAM9,
    Tile_X10Y12_BM_SRAM0,
    Tile_X10Y12_BM_SRAM1,
    Tile_X10Y12_BM_SRAM10,
    Tile_X10Y12_BM_SRAM11,
    Tile_X10Y12_BM_SRAM12,
    Tile_X10Y12_BM_SRAM13,
    Tile_X10Y12_BM_SRAM14,
    Tile_X10Y12_BM_SRAM15,
    Tile_X10Y12_BM_SRAM16,
    Tile_X10Y12_BM_SRAM17,
    Tile_X10Y12_BM_SRAM18,
    Tile_X10Y12_BM_SRAM19,
    Tile_X10Y12_BM_SRAM2,
    Tile_X10Y12_BM_SRAM20,
    Tile_X10Y12_BM_SRAM21,
    Tile_X10Y12_BM_SRAM22,
    Tile_X10Y12_BM_SRAM23,
    Tile_X10Y12_BM_SRAM24,
    Tile_X10Y12_BM_SRAM25,
    Tile_X10Y12_BM_SRAM26,
    Tile_X10Y12_BM_SRAM27,
    Tile_X10Y12_BM_SRAM28,
    Tile_X10Y12_BM_SRAM29,
    Tile_X10Y12_BM_SRAM3,
    Tile_X10Y12_BM_SRAM30,
    Tile_X10Y12_BM_SRAM31,
    Tile_X10Y12_BM_SRAM4,
    Tile_X10Y12_BM_SRAM5,
    Tile_X10Y12_BM_SRAM6,
    Tile_X10Y12_BM_SRAM7,
    Tile_X10Y12_BM_SRAM8,
    Tile_X10Y12_BM_SRAM9,
    Tile_X10Y12_CLK_SRAM,
    Tile_X10Y12_CONFIGURED_top,
    Tile_X10Y12_DIN_SRAM0,
    Tile_X10Y12_DIN_SRAM1,
    Tile_X10Y12_DIN_SRAM10,
    Tile_X10Y12_DIN_SRAM11,
    Tile_X10Y12_DIN_SRAM12,
    Tile_X10Y12_DIN_SRAM13,
    Tile_X10Y12_DIN_SRAM14,
    Tile_X10Y12_DIN_SRAM15,
    Tile_X10Y12_DIN_SRAM16,
    Tile_X10Y12_DIN_SRAM17,
    Tile_X10Y12_DIN_SRAM18,
    Tile_X10Y12_DIN_SRAM19,
    Tile_X10Y12_DIN_SRAM2,
    Tile_X10Y12_DIN_SRAM20,
    Tile_X10Y12_DIN_SRAM21,
    Tile_X10Y12_DIN_SRAM22,
    Tile_X10Y12_DIN_SRAM23,
    Tile_X10Y12_DIN_SRAM24,
    Tile_X10Y12_DIN_SRAM25,
    Tile_X10Y12_DIN_SRAM26,
    Tile_X10Y12_DIN_SRAM27,
    Tile_X10Y12_DIN_SRAM28,
    Tile_X10Y12_DIN_SRAM29,
    Tile_X10Y12_DIN_SRAM3,
    Tile_X10Y12_DIN_SRAM30,
    Tile_X10Y12_DIN_SRAM31,
    Tile_X10Y12_DIN_SRAM4,
    Tile_X10Y12_DIN_SRAM5,
    Tile_X10Y12_DIN_SRAM6,
    Tile_X10Y12_DIN_SRAM7,
    Tile_X10Y12_DIN_SRAM8,
    Tile_X10Y12_DIN_SRAM9,
    Tile_X10Y12_DOUT_SRAM0,
    Tile_X10Y12_DOUT_SRAM1,
    Tile_X10Y12_DOUT_SRAM10,
    Tile_X10Y12_DOUT_SRAM11,
    Tile_X10Y12_DOUT_SRAM12,
    Tile_X10Y12_DOUT_SRAM13,
    Tile_X10Y12_DOUT_SRAM14,
    Tile_X10Y12_DOUT_SRAM15,
    Tile_X10Y12_DOUT_SRAM16,
    Tile_X10Y12_DOUT_SRAM17,
    Tile_X10Y12_DOUT_SRAM18,
    Tile_X10Y12_DOUT_SRAM19,
    Tile_X10Y12_DOUT_SRAM2,
    Tile_X10Y12_DOUT_SRAM20,
    Tile_X10Y12_DOUT_SRAM21,
    Tile_X10Y12_DOUT_SRAM22,
    Tile_X10Y12_DOUT_SRAM23,
    Tile_X10Y12_DOUT_SRAM24,
    Tile_X10Y12_DOUT_SRAM25,
    Tile_X10Y12_DOUT_SRAM26,
    Tile_X10Y12_DOUT_SRAM27,
    Tile_X10Y12_DOUT_SRAM28,
    Tile_X10Y12_DOUT_SRAM29,
    Tile_X10Y12_DOUT_SRAM3,
    Tile_X10Y12_DOUT_SRAM30,
    Tile_X10Y12_DOUT_SRAM31,
    Tile_X10Y12_DOUT_SRAM4,
    Tile_X10Y12_DOUT_SRAM5,
    Tile_X10Y12_DOUT_SRAM6,
    Tile_X10Y12_DOUT_SRAM7,
    Tile_X10Y12_DOUT_SRAM8,
    Tile_X10Y12_DOUT_SRAM9,
    Tile_X10Y12_MEN_SRAM,
    Tile_X10Y12_REN_SRAM,
    Tile_X10Y12_TIE_HIGH_SRAM,
    Tile_X10Y12_TIE_LOW_SRAM,
    Tile_X10Y12_WEN_SRAM,
    Tile_X10Y14_ADDR_SRAM0,
    Tile_X10Y14_ADDR_SRAM1,
    Tile_X10Y14_ADDR_SRAM2,
    Tile_X10Y14_ADDR_SRAM3,
    Tile_X10Y14_ADDR_SRAM4,
    Tile_X10Y14_ADDR_SRAM5,
    Tile_X10Y14_ADDR_SRAM6,
    Tile_X10Y14_ADDR_SRAM7,
    Tile_X10Y14_ADDR_SRAM8,
    Tile_X10Y14_ADDR_SRAM9,
    Tile_X10Y14_BM_SRAM0,
    Tile_X10Y14_BM_SRAM1,
    Tile_X10Y14_BM_SRAM10,
    Tile_X10Y14_BM_SRAM11,
    Tile_X10Y14_BM_SRAM12,
    Tile_X10Y14_BM_SRAM13,
    Tile_X10Y14_BM_SRAM14,
    Tile_X10Y14_BM_SRAM15,
    Tile_X10Y14_BM_SRAM16,
    Tile_X10Y14_BM_SRAM17,
    Tile_X10Y14_BM_SRAM18,
    Tile_X10Y14_BM_SRAM19,
    Tile_X10Y14_BM_SRAM2,
    Tile_X10Y14_BM_SRAM20,
    Tile_X10Y14_BM_SRAM21,
    Tile_X10Y14_BM_SRAM22,
    Tile_X10Y14_BM_SRAM23,
    Tile_X10Y14_BM_SRAM24,
    Tile_X10Y14_BM_SRAM25,
    Tile_X10Y14_BM_SRAM26,
    Tile_X10Y14_BM_SRAM27,
    Tile_X10Y14_BM_SRAM28,
    Tile_X10Y14_BM_SRAM29,
    Tile_X10Y14_BM_SRAM3,
    Tile_X10Y14_BM_SRAM30,
    Tile_X10Y14_BM_SRAM31,
    Tile_X10Y14_BM_SRAM4,
    Tile_X10Y14_BM_SRAM5,
    Tile_X10Y14_BM_SRAM6,
    Tile_X10Y14_BM_SRAM7,
    Tile_X10Y14_BM_SRAM8,
    Tile_X10Y14_BM_SRAM9,
    Tile_X10Y14_CLK_SRAM,
    Tile_X10Y14_CONFIGURED_top,
    Tile_X10Y14_DIN_SRAM0,
    Tile_X10Y14_DIN_SRAM1,
    Tile_X10Y14_DIN_SRAM10,
    Tile_X10Y14_DIN_SRAM11,
    Tile_X10Y14_DIN_SRAM12,
    Tile_X10Y14_DIN_SRAM13,
    Tile_X10Y14_DIN_SRAM14,
    Tile_X10Y14_DIN_SRAM15,
    Tile_X10Y14_DIN_SRAM16,
    Tile_X10Y14_DIN_SRAM17,
    Tile_X10Y14_DIN_SRAM18,
    Tile_X10Y14_DIN_SRAM19,
    Tile_X10Y14_DIN_SRAM2,
    Tile_X10Y14_DIN_SRAM20,
    Tile_X10Y14_DIN_SRAM21,
    Tile_X10Y14_DIN_SRAM22,
    Tile_X10Y14_DIN_SRAM23,
    Tile_X10Y14_DIN_SRAM24,
    Tile_X10Y14_DIN_SRAM25,
    Tile_X10Y14_DIN_SRAM26,
    Tile_X10Y14_DIN_SRAM27,
    Tile_X10Y14_DIN_SRAM28,
    Tile_X10Y14_DIN_SRAM29,
    Tile_X10Y14_DIN_SRAM3,
    Tile_X10Y14_DIN_SRAM30,
    Tile_X10Y14_DIN_SRAM31,
    Tile_X10Y14_DIN_SRAM4,
    Tile_X10Y14_DIN_SRAM5,
    Tile_X10Y14_DIN_SRAM6,
    Tile_X10Y14_DIN_SRAM7,
    Tile_X10Y14_DIN_SRAM8,
    Tile_X10Y14_DIN_SRAM9,
    Tile_X10Y14_DOUT_SRAM0,
    Tile_X10Y14_DOUT_SRAM1,
    Tile_X10Y14_DOUT_SRAM10,
    Tile_X10Y14_DOUT_SRAM11,
    Tile_X10Y14_DOUT_SRAM12,
    Tile_X10Y14_DOUT_SRAM13,
    Tile_X10Y14_DOUT_SRAM14,
    Tile_X10Y14_DOUT_SRAM15,
    Tile_X10Y14_DOUT_SRAM16,
    Tile_X10Y14_DOUT_SRAM17,
    Tile_X10Y14_DOUT_SRAM18,
    Tile_X10Y14_DOUT_SRAM19,
    Tile_X10Y14_DOUT_SRAM2,
    Tile_X10Y14_DOUT_SRAM20,
    Tile_X10Y14_DOUT_SRAM21,
    Tile_X10Y14_DOUT_SRAM22,
    Tile_X10Y14_DOUT_SRAM23,
    Tile_X10Y14_DOUT_SRAM24,
    Tile_X10Y14_DOUT_SRAM25,
    Tile_X10Y14_DOUT_SRAM26,
    Tile_X10Y14_DOUT_SRAM27,
    Tile_X10Y14_DOUT_SRAM28,
    Tile_X10Y14_DOUT_SRAM29,
    Tile_X10Y14_DOUT_SRAM3,
    Tile_X10Y14_DOUT_SRAM30,
    Tile_X10Y14_DOUT_SRAM31,
    Tile_X10Y14_DOUT_SRAM4,
    Tile_X10Y14_DOUT_SRAM5,
    Tile_X10Y14_DOUT_SRAM6,
    Tile_X10Y14_DOUT_SRAM7,
    Tile_X10Y14_DOUT_SRAM8,
    Tile_X10Y14_DOUT_SRAM9,
    Tile_X10Y14_MEN_SRAM,
    Tile_X10Y14_REN_SRAM,
    Tile_X10Y14_TIE_HIGH_SRAM,
    Tile_X10Y14_TIE_LOW_SRAM,
    Tile_X10Y14_WEN_SRAM,
    Tile_X10Y2_ADDR_SRAM0,
    Tile_X10Y2_ADDR_SRAM1,
    Tile_X10Y2_ADDR_SRAM2,
    Tile_X10Y2_ADDR_SRAM3,
    Tile_X10Y2_ADDR_SRAM4,
    Tile_X10Y2_ADDR_SRAM5,
    Tile_X10Y2_ADDR_SRAM6,
    Tile_X10Y2_ADDR_SRAM7,
    Tile_X10Y2_ADDR_SRAM8,
    Tile_X10Y2_ADDR_SRAM9,
    Tile_X10Y2_BM_SRAM0,
    Tile_X10Y2_BM_SRAM1,
    Tile_X10Y2_BM_SRAM10,
    Tile_X10Y2_BM_SRAM11,
    Tile_X10Y2_BM_SRAM12,
    Tile_X10Y2_BM_SRAM13,
    Tile_X10Y2_BM_SRAM14,
    Tile_X10Y2_BM_SRAM15,
    Tile_X10Y2_BM_SRAM16,
    Tile_X10Y2_BM_SRAM17,
    Tile_X10Y2_BM_SRAM18,
    Tile_X10Y2_BM_SRAM19,
    Tile_X10Y2_BM_SRAM2,
    Tile_X10Y2_BM_SRAM20,
    Tile_X10Y2_BM_SRAM21,
    Tile_X10Y2_BM_SRAM22,
    Tile_X10Y2_BM_SRAM23,
    Tile_X10Y2_BM_SRAM24,
    Tile_X10Y2_BM_SRAM25,
    Tile_X10Y2_BM_SRAM26,
    Tile_X10Y2_BM_SRAM27,
    Tile_X10Y2_BM_SRAM28,
    Tile_X10Y2_BM_SRAM29,
    Tile_X10Y2_BM_SRAM3,
    Tile_X10Y2_BM_SRAM30,
    Tile_X10Y2_BM_SRAM31,
    Tile_X10Y2_BM_SRAM4,
    Tile_X10Y2_BM_SRAM5,
    Tile_X10Y2_BM_SRAM6,
    Tile_X10Y2_BM_SRAM7,
    Tile_X10Y2_BM_SRAM8,
    Tile_X10Y2_BM_SRAM9,
    Tile_X10Y2_CLK_SRAM,
    Tile_X10Y2_CONFIGURED_top,
    Tile_X10Y2_DIN_SRAM0,
    Tile_X10Y2_DIN_SRAM1,
    Tile_X10Y2_DIN_SRAM10,
    Tile_X10Y2_DIN_SRAM11,
    Tile_X10Y2_DIN_SRAM12,
    Tile_X10Y2_DIN_SRAM13,
    Tile_X10Y2_DIN_SRAM14,
    Tile_X10Y2_DIN_SRAM15,
    Tile_X10Y2_DIN_SRAM16,
    Tile_X10Y2_DIN_SRAM17,
    Tile_X10Y2_DIN_SRAM18,
    Tile_X10Y2_DIN_SRAM19,
    Tile_X10Y2_DIN_SRAM2,
    Tile_X10Y2_DIN_SRAM20,
    Tile_X10Y2_DIN_SRAM21,
    Tile_X10Y2_DIN_SRAM22,
    Tile_X10Y2_DIN_SRAM23,
    Tile_X10Y2_DIN_SRAM24,
    Tile_X10Y2_DIN_SRAM25,
    Tile_X10Y2_DIN_SRAM26,
    Tile_X10Y2_DIN_SRAM27,
    Tile_X10Y2_DIN_SRAM28,
    Tile_X10Y2_DIN_SRAM29,
    Tile_X10Y2_DIN_SRAM3,
    Tile_X10Y2_DIN_SRAM30,
    Tile_X10Y2_DIN_SRAM31,
    Tile_X10Y2_DIN_SRAM4,
    Tile_X10Y2_DIN_SRAM5,
    Tile_X10Y2_DIN_SRAM6,
    Tile_X10Y2_DIN_SRAM7,
    Tile_X10Y2_DIN_SRAM8,
    Tile_X10Y2_DIN_SRAM9,
    Tile_X10Y2_DOUT_SRAM0,
    Tile_X10Y2_DOUT_SRAM1,
    Tile_X10Y2_DOUT_SRAM10,
    Tile_X10Y2_DOUT_SRAM11,
    Tile_X10Y2_DOUT_SRAM12,
    Tile_X10Y2_DOUT_SRAM13,
    Tile_X10Y2_DOUT_SRAM14,
    Tile_X10Y2_DOUT_SRAM15,
    Tile_X10Y2_DOUT_SRAM16,
    Tile_X10Y2_DOUT_SRAM17,
    Tile_X10Y2_DOUT_SRAM18,
    Tile_X10Y2_DOUT_SRAM19,
    Tile_X10Y2_DOUT_SRAM2,
    Tile_X10Y2_DOUT_SRAM20,
    Tile_X10Y2_DOUT_SRAM21,
    Tile_X10Y2_DOUT_SRAM22,
    Tile_X10Y2_DOUT_SRAM23,
    Tile_X10Y2_DOUT_SRAM24,
    Tile_X10Y2_DOUT_SRAM25,
    Tile_X10Y2_DOUT_SRAM26,
    Tile_X10Y2_DOUT_SRAM27,
    Tile_X10Y2_DOUT_SRAM28,
    Tile_X10Y2_DOUT_SRAM29,
    Tile_X10Y2_DOUT_SRAM3,
    Tile_X10Y2_DOUT_SRAM30,
    Tile_X10Y2_DOUT_SRAM31,
    Tile_X10Y2_DOUT_SRAM4,
    Tile_X10Y2_DOUT_SRAM5,
    Tile_X10Y2_DOUT_SRAM6,
    Tile_X10Y2_DOUT_SRAM7,
    Tile_X10Y2_DOUT_SRAM8,
    Tile_X10Y2_DOUT_SRAM9,
    Tile_X10Y2_MEN_SRAM,
    Tile_X10Y2_REN_SRAM,
    Tile_X10Y2_TIE_HIGH_SRAM,
    Tile_X10Y2_TIE_LOW_SRAM,
    Tile_X10Y2_WEN_SRAM,
    Tile_X10Y4_ADDR_SRAM0,
    Tile_X10Y4_ADDR_SRAM1,
    Tile_X10Y4_ADDR_SRAM2,
    Tile_X10Y4_ADDR_SRAM3,
    Tile_X10Y4_ADDR_SRAM4,
    Tile_X10Y4_ADDR_SRAM5,
    Tile_X10Y4_ADDR_SRAM6,
    Tile_X10Y4_ADDR_SRAM7,
    Tile_X10Y4_ADDR_SRAM8,
    Tile_X10Y4_ADDR_SRAM9,
    Tile_X10Y4_BM_SRAM0,
    Tile_X10Y4_BM_SRAM1,
    Tile_X10Y4_BM_SRAM10,
    Tile_X10Y4_BM_SRAM11,
    Tile_X10Y4_BM_SRAM12,
    Tile_X10Y4_BM_SRAM13,
    Tile_X10Y4_BM_SRAM14,
    Tile_X10Y4_BM_SRAM15,
    Tile_X10Y4_BM_SRAM16,
    Tile_X10Y4_BM_SRAM17,
    Tile_X10Y4_BM_SRAM18,
    Tile_X10Y4_BM_SRAM19,
    Tile_X10Y4_BM_SRAM2,
    Tile_X10Y4_BM_SRAM20,
    Tile_X10Y4_BM_SRAM21,
    Tile_X10Y4_BM_SRAM22,
    Tile_X10Y4_BM_SRAM23,
    Tile_X10Y4_BM_SRAM24,
    Tile_X10Y4_BM_SRAM25,
    Tile_X10Y4_BM_SRAM26,
    Tile_X10Y4_BM_SRAM27,
    Tile_X10Y4_BM_SRAM28,
    Tile_X10Y4_BM_SRAM29,
    Tile_X10Y4_BM_SRAM3,
    Tile_X10Y4_BM_SRAM30,
    Tile_X10Y4_BM_SRAM31,
    Tile_X10Y4_BM_SRAM4,
    Tile_X10Y4_BM_SRAM5,
    Tile_X10Y4_BM_SRAM6,
    Tile_X10Y4_BM_SRAM7,
    Tile_X10Y4_BM_SRAM8,
    Tile_X10Y4_BM_SRAM9,
    Tile_X10Y4_CLK_SRAM,
    Tile_X10Y4_CONFIGURED_top,
    Tile_X10Y4_DIN_SRAM0,
    Tile_X10Y4_DIN_SRAM1,
    Tile_X10Y4_DIN_SRAM10,
    Tile_X10Y4_DIN_SRAM11,
    Tile_X10Y4_DIN_SRAM12,
    Tile_X10Y4_DIN_SRAM13,
    Tile_X10Y4_DIN_SRAM14,
    Tile_X10Y4_DIN_SRAM15,
    Tile_X10Y4_DIN_SRAM16,
    Tile_X10Y4_DIN_SRAM17,
    Tile_X10Y4_DIN_SRAM18,
    Tile_X10Y4_DIN_SRAM19,
    Tile_X10Y4_DIN_SRAM2,
    Tile_X10Y4_DIN_SRAM20,
    Tile_X10Y4_DIN_SRAM21,
    Tile_X10Y4_DIN_SRAM22,
    Tile_X10Y4_DIN_SRAM23,
    Tile_X10Y4_DIN_SRAM24,
    Tile_X10Y4_DIN_SRAM25,
    Tile_X10Y4_DIN_SRAM26,
    Tile_X10Y4_DIN_SRAM27,
    Tile_X10Y4_DIN_SRAM28,
    Tile_X10Y4_DIN_SRAM29,
    Tile_X10Y4_DIN_SRAM3,
    Tile_X10Y4_DIN_SRAM30,
    Tile_X10Y4_DIN_SRAM31,
    Tile_X10Y4_DIN_SRAM4,
    Tile_X10Y4_DIN_SRAM5,
    Tile_X10Y4_DIN_SRAM6,
    Tile_X10Y4_DIN_SRAM7,
    Tile_X10Y4_DIN_SRAM8,
    Tile_X10Y4_DIN_SRAM9,
    Tile_X10Y4_DOUT_SRAM0,
    Tile_X10Y4_DOUT_SRAM1,
    Tile_X10Y4_DOUT_SRAM10,
    Tile_X10Y4_DOUT_SRAM11,
    Tile_X10Y4_DOUT_SRAM12,
    Tile_X10Y4_DOUT_SRAM13,
    Tile_X10Y4_DOUT_SRAM14,
    Tile_X10Y4_DOUT_SRAM15,
    Tile_X10Y4_DOUT_SRAM16,
    Tile_X10Y4_DOUT_SRAM17,
    Tile_X10Y4_DOUT_SRAM18,
    Tile_X10Y4_DOUT_SRAM19,
    Tile_X10Y4_DOUT_SRAM2,
    Tile_X10Y4_DOUT_SRAM20,
    Tile_X10Y4_DOUT_SRAM21,
    Tile_X10Y4_DOUT_SRAM22,
    Tile_X10Y4_DOUT_SRAM23,
    Tile_X10Y4_DOUT_SRAM24,
    Tile_X10Y4_DOUT_SRAM25,
    Tile_X10Y4_DOUT_SRAM26,
    Tile_X10Y4_DOUT_SRAM27,
    Tile_X10Y4_DOUT_SRAM28,
    Tile_X10Y4_DOUT_SRAM29,
    Tile_X10Y4_DOUT_SRAM3,
    Tile_X10Y4_DOUT_SRAM30,
    Tile_X10Y4_DOUT_SRAM31,
    Tile_X10Y4_DOUT_SRAM4,
    Tile_X10Y4_DOUT_SRAM5,
    Tile_X10Y4_DOUT_SRAM6,
    Tile_X10Y4_DOUT_SRAM7,
    Tile_X10Y4_DOUT_SRAM8,
    Tile_X10Y4_DOUT_SRAM9,
    Tile_X10Y4_MEN_SRAM,
    Tile_X10Y4_REN_SRAM,
    Tile_X10Y4_TIE_HIGH_SRAM,
    Tile_X10Y4_TIE_LOW_SRAM,
    Tile_X10Y4_WEN_SRAM,
    Tile_X10Y6_ADDR_SRAM0,
    Tile_X10Y6_ADDR_SRAM1,
    Tile_X10Y6_ADDR_SRAM2,
    Tile_X10Y6_ADDR_SRAM3,
    Tile_X10Y6_ADDR_SRAM4,
    Tile_X10Y6_ADDR_SRAM5,
    Tile_X10Y6_ADDR_SRAM6,
    Tile_X10Y6_ADDR_SRAM7,
    Tile_X10Y6_ADDR_SRAM8,
    Tile_X10Y6_ADDR_SRAM9,
    Tile_X10Y6_BM_SRAM0,
    Tile_X10Y6_BM_SRAM1,
    Tile_X10Y6_BM_SRAM10,
    Tile_X10Y6_BM_SRAM11,
    Tile_X10Y6_BM_SRAM12,
    Tile_X10Y6_BM_SRAM13,
    Tile_X10Y6_BM_SRAM14,
    Tile_X10Y6_BM_SRAM15,
    Tile_X10Y6_BM_SRAM16,
    Tile_X10Y6_BM_SRAM17,
    Tile_X10Y6_BM_SRAM18,
    Tile_X10Y6_BM_SRAM19,
    Tile_X10Y6_BM_SRAM2,
    Tile_X10Y6_BM_SRAM20,
    Tile_X10Y6_BM_SRAM21,
    Tile_X10Y6_BM_SRAM22,
    Tile_X10Y6_BM_SRAM23,
    Tile_X10Y6_BM_SRAM24,
    Tile_X10Y6_BM_SRAM25,
    Tile_X10Y6_BM_SRAM26,
    Tile_X10Y6_BM_SRAM27,
    Tile_X10Y6_BM_SRAM28,
    Tile_X10Y6_BM_SRAM29,
    Tile_X10Y6_BM_SRAM3,
    Tile_X10Y6_BM_SRAM30,
    Tile_X10Y6_BM_SRAM31,
    Tile_X10Y6_BM_SRAM4,
    Tile_X10Y6_BM_SRAM5,
    Tile_X10Y6_BM_SRAM6,
    Tile_X10Y6_BM_SRAM7,
    Tile_X10Y6_BM_SRAM8,
    Tile_X10Y6_BM_SRAM9,
    Tile_X10Y6_CLK_SRAM,
    Tile_X10Y6_CONFIGURED_top,
    Tile_X10Y6_DIN_SRAM0,
    Tile_X10Y6_DIN_SRAM1,
    Tile_X10Y6_DIN_SRAM10,
    Tile_X10Y6_DIN_SRAM11,
    Tile_X10Y6_DIN_SRAM12,
    Tile_X10Y6_DIN_SRAM13,
    Tile_X10Y6_DIN_SRAM14,
    Tile_X10Y6_DIN_SRAM15,
    Tile_X10Y6_DIN_SRAM16,
    Tile_X10Y6_DIN_SRAM17,
    Tile_X10Y6_DIN_SRAM18,
    Tile_X10Y6_DIN_SRAM19,
    Tile_X10Y6_DIN_SRAM2,
    Tile_X10Y6_DIN_SRAM20,
    Tile_X10Y6_DIN_SRAM21,
    Tile_X10Y6_DIN_SRAM22,
    Tile_X10Y6_DIN_SRAM23,
    Tile_X10Y6_DIN_SRAM24,
    Tile_X10Y6_DIN_SRAM25,
    Tile_X10Y6_DIN_SRAM26,
    Tile_X10Y6_DIN_SRAM27,
    Tile_X10Y6_DIN_SRAM28,
    Tile_X10Y6_DIN_SRAM29,
    Tile_X10Y6_DIN_SRAM3,
    Tile_X10Y6_DIN_SRAM30,
    Tile_X10Y6_DIN_SRAM31,
    Tile_X10Y6_DIN_SRAM4,
    Tile_X10Y6_DIN_SRAM5,
    Tile_X10Y6_DIN_SRAM6,
    Tile_X10Y6_DIN_SRAM7,
    Tile_X10Y6_DIN_SRAM8,
    Tile_X10Y6_DIN_SRAM9,
    Tile_X10Y6_DOUT_SRAM0,
    Tile_X10Y6_DOUT_SRAM1,
    Tile_X10Y6_DOUT_SRAM10,
    Tile_X10Y6_DOUT_SRAM11,
    Tile_X10Y6_DOUT_SRAM12,
    Tile_X10Y6_DOUT_SRAM13,
    Tile_X10Y6_DOUT_SRAM14,
    Tile_X10Y6_DOUT_SRAM15,
    Tile_X10Y6_DOUT_SRAM16,
    Tile_X10Y6_DOUT_SRAM17,
    Tile_X10Y6_DOUT_SRAM18,
    Tile_X10Y6_DOUT_SRAM19,
    Tile_X10Y6_DOUT_SRAM2,
    Tile_X10Y6_DOUT_SRAM20,
    Tile_X10Y6_DOUT_SRAM21,
    Tile_X10Y6_DOUT_SRAM22,
    Tile_X10Y6_DOUT_SRAM23,
    Tile_X10Y6_DOUT_SRAM24,
    Tile_X10Y6_DOUT_SRAM25,
    Tile_X10Y6_DOUT_SRAM26,
    Tile_X10Y6_DOUT_SRAM27,
    Tile_X10Y6_DOUT_SRAM28,
    Tile_X10Y6_DOUT_SRAM29,
    Tile_X10Y6_DOUT_SRAM3,
    Tile_X10Y6_DOUT_SRAM30,
    Tile_X10Y6_DOUT_SRAM31,
    Tile_X10Y6_DOUT_SRAM4,
    Tile_X10Y6_DOUT_SRAM5,
    Tile_X10Y6_DOUT_SRAM6,
    Tile_X10Y6_DOUT_SRAM7,
    Tile_X10Y6_DOUT_SRAM8,
    Tile_X10Y6_DOUT_SRAM9,
    Tile_X10Y6_MEN_SRAM,
    Tile_X10Y6_REN_SRAM,
    Tile_X10Y6_TIE_HIGH_SRAM,
    Tile_X10Y6_TIE_LOW_SRAM,
    Tile_X10Y6_WEN_SRAM,
    Tile_X10Y8_ADDR_SRAM0,
    Tile_X10Y8_ADDR_SRAM1,
    Tile_X10Y8_ADDR_SRAM2,
    Tile_X10Y8_ADDR_SRAM3,
    Tile_X10Y8_ADDR_SRAM4,
    Tile_X10Y8_ADDR_SRAM5,
    Tile_X10Y8_ADDR_SRAM6,
    Tile_X10Y8_ADDR_SRAM7,
    Tile_X10Y8_ADDR_SRAM8,
    Tile_X10Y8_ADDR_SRAM9,
    Tile_X10Y8_BM_SRAM0,
    Tile_X10Y8_BM_SRAM1,
    Tile_X10Y8_BM_SRAM10,
    Tile_X10Y8_BM_SRAM11,
    Tile_X10Y8_BM_SRAM12,
    Tile_X10Y8_BM_SRAM13,
    Tile_X10Y8_BM_SRAM14,
    Tile_X10Y8_BM_SRAM15,
    Tile_X10Y8_BM_SRAM16,
    Tile_X10Y8_BM_SRAM17,
    Tile_X10Y8_BM_SRAM18,
    Tile_X10Y8_BM_SRAM19,
    Tile_X10Y8_BM_SRAM2,
    Tile_X10Y8_BM_SRAM20,
    Tile_X10Y8_BM_SRAM21,
    Tile_X10Y8_BM_SRAM22,
    Tile_X10Y8_BM_SRAM23,
    Tile_X10Y8_BM_SRAM24,
    Tile_X10Y8_BM_SRAM25,
    Tile_X10Y8_BM_SRAM26,
    Tile_X10Y8_BM_SRAM27,
    Tile_X10Y8_BM_SRAM28,
    Tile_X10Y8_BM_SRAM29,
    Tile_X10Y8_BM_SRAM3,
    Tile_X10Y8_BM_SRAM30,
    Tile_X10Y8_BM_SRAM31,
    Tile_X10Y8_BM_SRAM4,
    Tile_X10Y8_BM_SRAM5,
    Tile_X10Y8_BM_SRAM6,
    Tile_X10Y8_BM_SRAM7,
    Tile_X10Y8_BM_SRAM8,
    Tile_X10Y8_BM_SRAM9,
    Tile_X10Y8_CLK_SRAM,
    Tile_X10Y8_CONFIGURED_top,
    Tile_X10Y8_DIN_SRAM0,
    Tile_X10Y8_DIN_SRAM1,
    Tile_X10Y8_DIN_SRAM10,
    Tile_X10Y8_DIN_SRAM11,
    Tile_X10Y8_DIN_SRAM12,
    Tile_X10Y8_DIN_SRAM13,
    Tile_X10Y8_DIN_SRAM14,
    Tile_X10Y8_DIN_SRAM15,
    Tile_X10Y8_DIN_SRAM16,
    Tile_X10Y8_DIN_SRAM17,
    Tile_X10Y8_DIN_SRAM18,
    Tile_X10Y8_DIN_SRAM19,
    Tile_X10Y8_DIN_SRAM2,
    Tile_X10Y8_DIN_SRAM20,
    Tile_X10Y8_DIN_SRAM21,
    Tile_X10Y8_DIN_SRAM22,
    Tile_X10Y8_DIN_SRAM23,
    Tile_X10Y8_DIN_SRAM24,
    Tile_X10Y8_DIN_SRAM25,
    Tile_X10Y8_DIN_SRAM26,
    Tile_X10Y8_DIN_SRAM27,
    Tile_X10Y8_DIN_SRAM28,
    Tile_X10Y8_DIN_SRAM29,
    Tile_X10Y8_DIN_SRAM3,
    Tile_X10Y8_DIN_SRAM30,
    Tile_X10Y8_DIN_SRAM31,
    Tile_X10Y8_DIN_SRAM4,
    Tile_X10Y8_DIN_SRAM5,
    Tile_X10Y8_DIN_SRAM6,
    Tile_X10Y8_DIN_SRAM7,
    Tile_X10Y8_DIN_SRAM8,
    Tile_X10Y8_DIN_SRAM9,
    Tile_X10Y8_DOUT_SRAM0,
    Tile_X10Y8_DOUT_SRAM1,
    Tile_X10Y8_DOUT_SRAM10,
    Tile_X10Y8_DOUT_SRAM11,
    Tile_X10Y8_DOUT_SRAM12,
    Tile_X10Y8_DOUT_SRAM13,
    Tile_X10Y8_DOUT_SRAM14,
    Tile_X10Y8_DOUT_SRAM15,
    Tile_X10Y8_DOUT_SRAM16,
    Tile_X10Y8_DOUT_SRAM17,
    Tile_X10Y8_DOUT_SRAM18,
    Tile_X10Y8_DOUT_SRAM19,
    Tile_X10Y8_DOUT_SRAM2,
    Tile_X10Y8_DOUT_SRAM20,
    Tile_X10Y8_DOUT_SRAM21,
    Tile_X10Y8_DOUT_SRAM22,
    Tile_X10Y8_DOUT_SRAM23,
    Tile_X10Y8_DOUT_SRAM24,
    Tile_X10Y8_DOUT_SRAM25,
    Tile_X10Y8_DOUT_SRAM26,
    Tile_X10Y8_DOUT_SRAM27,
    Tile_X10Y8_DOUT_SRAM28,
    Tile_X10Y8_DOUT_SRAM29,
    Tile_X10Y8_DOUT_SRAM3,
    Tile_X10Y8_DOUT_SRAM30,
    Tile_X10Y8_DOUT_SRAM31,
    Tile_X10Y8_DOUT_SRAM4,
    Tile_X10Y8_DOUT_SRAM5,
    Tile_X10Y8_DOUT_SRAM6,
    Tile_X10Y8_DOUT_SRAM7,
    Tile_X10Y8_DOUT_SRAM8,
    Tile_X10Y8_DOUT_SRAM9,
    Tile_X10Y8_MEN_SRAM,
    Tile_X10Y8_REN_SRAM,
    Tile_X10Y8_TIE_HIGH_SRAM,
    Tile_X10Y8_TIE_LOW_SRAM,
    Tile_X10Y8_WEN_SRAM,
    Tile_X1Y0_A_I_top,
    Tile_X1Y0_A_O_top,
    Tile_X1Y0_A_T_top,
    Tile_X1Y0_A_config_C_bit0,
    Tile_X1Y0_A_config_C_bit1,
    Tile_X1Y0_A_config_C_bit2,
    Tile_X1Y0_A_config_C_bit3,
    Tile_X1Y0_B_I_top,
    Tile_X1Y0_B_O_top,
    Tile_X1Y0_B_T_top,
    Tile_X1Y0_B_config_C_bit0,
    Tile_X1Y0_B_config_C_bit1,
    Tile_X1Y0_B_config_C_bit2,
    Tile_X1Y0_B_config_C_bit3,
    Tile_X2Y0_A_I_top,
    Tile_X2Y0_A_O_top,
    Tile_X2Y0_A_T_top,
    Tile_X2Y0_A_config_C_bit0,
    Tile_X2Y0_A_config_C_bit1,
    Tile_X2Y0_A_config_C_bit2,
    Tile_X2Y0_A_config_C_bit3,
    Tile_X2Y0_B_I_top,
    Tile_X2Y0_B_O_top,
    Tile_X2Y0_B_T_top,
    Tile_X2Y0_B_config_C_bit0,
    Tile_X2Y0_B_config_C_bit1,
    Tile_X2Y0_B_config_C_bit2,
    Tile_X2Y0_B_config_C_bit3,
    Tile_X2Y15_BOOT_top,
    Tile_X2Y15_CONFIGURED_top,
    Tile_X2Y15_RESET_top,
    Tile_X2Y15_SLOT_top0,
    Tile_X2Y15_SLOT_top1,
    Tile_X2Y15_SLOT_top2,
    Tile_X2Y15_SLOT_top3,
    Tile_X3Y15_CONFIGURED_top,
    Tile_X3Y15_IRQ_top0,
    Tile_X3Y15_IRQ_top1,
    Tile_X3Y15_IRQ_top2,
    Tile_X3Y15_IRQ_top3,
    Tile_X5Y15_I_top0,
    Tile_X5Y15_I_top1,
    Tile_X5Y15_I_top10,
    Tile_X5Y15_I_top11,
    Tile_X5Y15_I_top12,
    Tile_X5Y15_I_top13,
    Tile_X5Y15_I_top14,
    Tile_X5Y15_I_top15,
    Tile_X5Y15_I_top2,
    Tile_X5Y15_I_top3,
    Tile_X5Y15_I_top4,
    Tile_X5Y15_I_top5,
    Tile_X5Y15_I_top6,
    Tile_X5Y15_I_top7,
    Tile_X5Y15_I_top8,
    Tile_X5Y15_I_top9,
    Tile_X5Y15_O_top0,
    Tile_X5Y15_O_top1,
    Tile_X5Y15_O_top10,
    Tile_X5Y15_O_top11,
    Tile_X5Y15_O_top12,
    Tile_X5Y15_O_top13,
    Tile_X5Y15_O_top14,
    Tile_X5Y15_O_top15,
    Tile_X5Y15_O_top2,
    Tile_X5Y15_O_top3,
    Tile_X5Y15_O_top4,
    Tile_X5Y15_O_top5,
    Tile_X5Y15_O_top6,
    Tile_X5Y15_O_top7,
    Tile_X5Y15_O_top8,
    Tile_X5Y15_O_top9,
    Tile_X6Y15_I_top0,
    Tile_X6Y15_I_top1,
    Tile_X6Y15_I_top10,
    Tile_X6Y15_I_top11,
    Tile_X6Y15_I_top12,
    Tile_X6Y15_I_top13,
    Tile_X6Y15_I_top14,
    Tile_X6Y15_I_top15,
    Tile_X6Y15_I_top2,
    Tile_X6Y15_I_top3,
    Tile_X6Y15_I_top4,
    Tile_X6Y15_I_top5,
    Tile_X6Y15_I_top6,
    Tile_X6Y15_I_top7,
    Tile_X6Y15_I_top8,
    Tile_X6Y15_I_top9,
    Tile_X6Y15_O_top0,
    Tile_X6Y15_O_top1,
    Tile_X6Y15_O_top10,
    Tile_X6Y15_O_top11,
    Tile_X6Y15_O_top12,
    Tile_X6Y15_O_top13,
    Tile_X6Y15_O_top14,
    Tile_X6Y15_O_top15,
    Tile_X6Y15_O_top2,
    Tile_X6Y15_O_top3,
    Tile_X6Y15_O_top4,
    Tile_X6Y15_O_top5,
    Tile_X6Y15_O_top6,
    Tile_X6Y15_O_top7,
    Tile_X6Y15_O_top8,
    Tile_X6Y15_O_top9,
    Tile_X8Y15_I_top0,
    Tile_X8Y15_I_top1,
    Tile_X8Y15_I_top10,
    Tile_X8Y15_I_top11,
    Tile_X8Y15_I_top12,
    Tile_X8Y15_I_top13,
    Tile_X8Y15_I_top14,
    Tile_X8Y15_I_top15,
    Tile_X8Y15_I_top2,
    Tile_X8Y15_I_top3,
    Tile_X8Y15_I_top4,
    Tile_X8Y15_I_top5,
    Tile_X8Y15_I_top6,
    Tile_X8Y15_I_top7,
    Tile_X8Y15_I_top8,
    Tile_X8Y15_I_top9,
    Tile_X8Y15_O_top0,
    Tile_X8Y15_O_top1,
    Tile_X8Y15_O_top10,
    Tile_X8Y15_O_top11,
    Tile_X8Y15_O_top12,
    Tile_X8Y15_O_top13,
    Tile_X8Y15_O_top14,
    Tile_X8Y15_O_top15,
    Tile_X8Y15_O_top2,
    Tile_X8Y15_O_top3,
    Tile_X8Y15_O_top4,
    Tile_X8Y15_O_top5,
    Tile_X8Y15_O_top6,
    Tile_X8Y15_O_top7,
    Tile_X8Y15_O_top8,
    Tile_X8Y15_O_top9,
    Tile_X9Y15_I_top0,
    Tile_X9Y15_I_top1,
    Tile_X9Y15_I_top10,
    Tile_X9Y15_I_top11,
    Tile_X9Y15_I_top12,
    Tile_X9Y15_I_top13,
    Tile_X9Y15_I_top14,
    Tile_X9Y15_I_top15,
    Tile_X9Y15_I_top2,
    Tile_X9Y15_I_top3,
    Tile_X9Y15_I_top4,
    Tile_X9Y15_I_top5,
    Tile_X9Y15_I_top6,
    Tile_X9Y15_I_top7,
    Tile_X9Y15_I_top8,
    Tile_X9Y15_I_top9,
    Tile_X9Y15_O_top0,
    Tile_X9Y15_O_top1,
    Tile_X9Y15_O_top10,
    Tile_X9Y15_O_top11,
    Tile_X9Y15_O_top12,
    Tile_X9Y15_O_top13,
    Tile_X9Y15_O_top14,
    Tile_X9Y15_O_top15,
    Tile_X9Y15_O_top2,
    Tile_X9Y15_O_top3,
    Tile_X9Y15_O_top4,
    Tile_X9Y15_O_top5,
    Tile_X9Y15_O_top6,
    Tile_X9Y15_O_top7,
    Tile_X9Y15_O_top8,
    Tile_X9Y15_O_top9,
    UserCLK,
    VPWR,
    VGND,
    FrameData,
    FrameStrobe);
 output Tile_X0Y10_A_I_top;
 input Tile_X0Y10_A_O_top;
 output Tile_X0Y10_A_T_top;
 output Tile_X0Y10_A_config_C_bit0;
 output Tile_X0Y10_A_config_C_bit1;
 output Tile_X0Y10_A_config_C_bit2;
 output Tile_X0Y10_A_config_C_bit3;
 output Tile_X0Y10_B_I_top;
 input Tile_X0Y10_B_O_top;
 output Tile_X0Y10_B_T_top;
 output Tile_X0Y10_B_config_C_bit0;
 output Tile_X0Y10_B_config_C_bit1;
 output Tile_X0Y10_B_config_C_bit2;
 output Tile_X0Y10_B_config_C_bit3;
 output Tile_X0Y11_A_I_top;
 input Tile_X0Y11_A_O_top;
 output Tile_X0Y11_A_T_top;
 output Tile_X0Y11_A_config_C_bit0;
 output Tile_X0Y11_A_config_C_bit1;
 output Tile_X0Y11_A_config_C_bit2;
 output Tile_X0Y11_A_config_C_bit3;
 output Tile_X0Y11_B_I_top;
 input Tile_X0Y11_B_O_top;
 output Tile_X0Y11_B_T_top;
 output Tile_X0Y11_B_config_C_bit0;
 output Tile_X0Y11_B_config_C_bit1;
 output Tile_X0Y11_B_config_C_bit2;
 output Tile_X0Y11_B_config_C_bit3;
 output Tile_X0Y12_A_I_top;
 input Tile_X0Y12_A_O_top;
 output Tile_X0Y12_A_T_top;
 output Tile_X0Y12_A_config_C_bit0;
 output Tile_X0Y12_A_config_C_bit1;
 output Tile_X0Y12_A_config_C_bit2;
 output Tile_X0Y12_A_config_C_bit3;
 output Tile_X0Y12_B_I_top;
 input Tile_X0Y12_B_O_top;
 output Tile_X0Y12_B_T_top;
 output Tile_X0Y12_B_config_C_bit0;
 output Tile_X0Y12_B_config_C_bit1;
 output Tile_X0Y12_B_config_C_bit2;
 output Tile_X0Y12_B_config_C_bit3;
 output Tile_X0Y13_A_I_top;
 input Tile_X0Y13_A_O_top;
 output Tile_X0Y13_A_T_top;
 output Tile_X0Y13_A_config_C_bit0;
 output Tile_X0Y13_A_config_C_bit1;
 output Tile_X0Y13_A_config_C_bit2;
 output Tile_X0Y13_A_config_C_bit3;
 output Tile_X0Y13_B_I_top;
 input Tile_X0Y13_B_O_top;
 output Tile_X0Y13_B_T_top;
 output Tile_X0Y13_B_config_C_bit0;
 output Tile_X0Y13_B_config_C_bit1;
 output Tile_X0Y13_B_config_C_bit2;
 output Tile_X0Y13_B_config_C_bit3;
 output Tile_X0Y14_A_I_top;
 input Tile_X0Y14_A_O_top;
 output Tile_X0Y14_A_T_top;
 output Tile_X0Y14_A_config_C_bit0;
 output Tile_X0Y14_A_config_C_bit1;
 output Tile_X0Y14_A_config_C_bit2;
 output Tile_X0Y14_A_config_C_bit3;
 output Tile_X0Y14_B_I_top;
 input Tile_X0Y14_B_O_top;
 output Tile_X0Y14_B_T_top;
 output Tile_X0Y14_B_config_C_bit0;
 output Tile_X0Y14_B_config_C_bit1;
 output Tile_X0Y14_B_config_C_bit2;
 output Tile_X0Y14_B_config_C_bit3;
 output Tile_X0Y1_A_I_top;
 input Tile_X0Y1_A_O_top;
 output Tile_X0Y1_A_T_top;
 output Tile_X0Y1_A_config_C_bit0;
 output Tile_X0Y1_A_config_C_bit1;
 output Tile_X0Y1_A_config_C_bit2;
 output Tile_X0Y1_A_config_C_bit3;
 output Tile_X0Y1_B_I_top;
 input Tile_X0Y1_B_O_top;
 output Tile_X0Y1_B_T_top;
 output Tile_X0Y1_B_config_C_bit0;
 output Tile_X0Y1_B_config_C_bit1;
 output Tile_X0Y1_B_config_C_bit2;
 output Tile_X0Y1_B_config_C_bit3;
 output Tile_X0Y2_A_I_top;
 input Tile_X0Y2_A_O_top;
 output Tile_X0Y2_A_T_top;
 output Tile_X0Y2_A_config_C_bit0;
 output Tile_X0Y2_A_config_C_bit1;
 output Tile_X0Y2_A_config_C_bit2;
 output Tile_X0Y2_A_config_C_bit3;
 output Tile_X0Y2_B_I_top;
 input Tile_X0Y2_B_O_top;
 output Tile_X0Y2_B_T_top;
 output Tile_X0Y2_B_config_C_bit0;
 output Tile_X0Y2_B_config_C_bit1;
 output Tile_X0Y2_B_config_C_bit2;
 output Tile_X0Y2_B_config_C_bit3;
 output Tile_X0Y3_A_I_top;
 input Tile_X0Y3_A_O_top;
 output Tile_X0Y3_A_T_top;
 output Tile_X0Y3_A_config_C_bit0;
 output Tile_X0Y3_A_config_C_bit1;
 output Tile_X0Y3_A_config_C_bit2;
 output Tile_X0Y3_A_config_C_bit3;
 output Tile_X0Y3_B_I_top;
 input Tile_X0Y3_B_O_top;
 output Tile_X0Y3_B_T_top;
 output Tile_X0Y3_B_config_C_bit0;
 output Tile_X0Y3_B_config_C_bit1;
 output Tile_X0Y3_B_config_C_bit2;
 output Tile_X0Y3_B_config_C_bit3;
 output Tile_X0Y4_A_I_top;
 input Tile_X0Y4_A_O_top;
 output Tile_X0Y4_A_T_top;
 output Tile_X0Y4_A_config_C_bit0;
 output Tile_X0Y4_A_config_C_bit1;
 output Tile_X0Y4_A_config_C_bit2;
 output Tile_X0Y4_A_config_C_bit3;
 output Tile_X0Y4_B_I_top;
 input Tile_X0Y4_B_O_top;
 output Tile_X0Y4_B_T_top;
 output Tile_X0Y4_B_config_C_bit0;
 output Tile_X0Y4_B_config_C_bit1;
 output Tile_X0Y4_B_config_C_bit2;
 output Tile_X0Y4_B_config_C_bit3;
 output Tile_X0Y5_A_I_top;
 input Tile_X0Y5_A_O_top;
 output Tile_X0Y5_A_T_top;
 output Tile_X0Y5_A_config_C_bit0;
 output Tile_X0Y5_A_config_C_bit1;
 output Tile_X0Y5_A_config_C_bit2;
 output Tile_X0Y5_A_config_C_bit3;
 output Tile_X0Y5_B_I_top;
 input Tile_X0Y5_B_O_top;
 output Tile_X0Y5_B_T_top;
 output Tile_X0Y5_B_config_C_bit0;
 output Tile_X0Y5_B_config_C_bit1;
 output Tile_X0Y5_B_config_C_bit2;
 output Tile_X0Y5_B_config_C_bit3;
 output Tile_X0Y6_A_I_top;
 input Tile_X0Y6_A_O_top;
 output Tile_X0Y6_A_T_top;
 output Tile_X0Y6_A_config_C_bit0;
 output Tile_X0Y6_A_config_C_bit1;
 output Tile_X0Y6_A_config_C_bit2;
 output Tile_X0Y6_A_config_C_bit3;
 output Tile_X0Y6_B_I_top;
 input Tile_X0Y6_B_O_top;
 output Tile_X0Y6_B_T_top;
 output Tile_X0Y6_B_config_C_bit0;
 output Tile_X0Y6_B_config_C_bit1;
 output Tile_X0Y6_B_config_C_bit2;
 output Tile_X0Y6_B_config_C_bit3;
 output Tile_X0Y7_A_I_top;
 input Tile_X0Y7_A_O_top;
 output Tile_X0Y7_A_T_top;
 output Tile_X0Y7_A_config_C_bit0;
 output Tile_X0Y7_A_config_C_bit1;
 output Tile_X0Y7_A_config_C_bit2;
 output Tile_X0Y7_A_config_C_bit3;
 output Tile_X0Y7_B_I_top;
 input Tile_X0Y7_B_O_top;
 output Tile_X0Y7_B_T_top;
 output Tile_X0Y7_B_config_C_bit0;
 output Tile_X0Y7_B_config_C_bit1;
 output Tile_X0Y7_B_config_C_bit2;
 output Tile_X0Y7_B_config_C_bit3;
 output Tile_X0Y8_A_I_top;
 input Tile_X0Y8_A_O_top;
 output Tile_X0Y8_A_T_top;
 output Tile_X0Y8_A_config_C_bit0;
 output Tile_X0Y8_A_config_C_bit1;
 output Tile_X0Y8_A_config_C_bit2;
 output Tile_X0Y8_A_config_C_bit3;
 output Tile_X0Y8_B_I_top;
 input Tile_X0Y8_B_O_top;
 output Tile_X0Y8_B_T_top;
 output Tile_X0Y8_B_config_C_bit0;
 output Tile_X0Y8_B_config_C_bit1;
 output Tile_X0Y8_B_config_C_bit2;
 output Tile_X0Y8_B_config_C_bit3;
 output Tile_X0Y9_A_I_top;
 input Tile_X0Y9_A_O_top;
 output Tile_X0Y9_A_T_top;
 output Tile_X0Y9_A_config_C_bit0;
 output Tile_X0Y9_A_config_C_bit1;
 output Tile_X0Y9_A_config_C_bit2;
 output Tile_X0Y9_A_config_C_bit3;
 output Tile_X0Y9_B_I_top;
 input Tile_X0Y9_B_O_top;
 output Tile_X0Y9_B_T_top;
 output Tile_X0Y9_B_config_C_bit0;
 output Tile_X0Y9_B_config_C_bit1;
 output Tile_X0Y9_B_config_C_bit2;
 output Tile_X0Y9_B_config_C_bit3;
 output Tile_X10Y10_ADDR_SRAM0;
 output Tile_X10Y10_ADDR_SRAM1;
 output Tile_X10Y10_ADDR_SRAM2;
 output Tile_X10Y10_ADDR_SRAM3;
 output Tile_X10Y10_ADDR_SRAM4;
 output Tile_X10Y10_ADDR_SRAM5;
 output Tile_X10Y10_ADDR_SRAM6;
 output Tile_X10Y10_ADDR_SRAM7;
 output Tile_X10Y10_ADDR_SRAM8;
 output Tile_X10Y10_ADDR_SRAM9;
 output Tile_X10Y10_BM_SRAM0;
 output Tile_X10Y10_BM_SRAM1;
 output Tile_X10Y10_BM_SRAM10;
 output Tile_X10Y10_BM_SRAM11;
 output Tile_X10Y10_BM_SRAM12;
 output Tile_X10Y10_BM_SRAM13;
 output Tile_X10Y10_BM_SRAM14;
 output Tile_X10Y10_BM_SRAM15;
 output Tile_X10Y10_BM_SRAM16;
 output Tile_X10Y10_BM_SRAM17;
 output Tile_X10Y10_BM_SRAM18;
 output Tile_X10Y10_BM_SRAM19;
 output Tile_X10Y10_BM_SRAM2;
 output Tile_X10Y10_BM_SRAM20;
 output Tile_X10Y10_BM_SRAM21;
 output Tile_X10Y10_BM_SRAM22;
 output Tile_X10Y10_BM_SRAM23;
 output Tile_X10Y10_BM_SRAM24;
 output Tile_X10Y10_BM_SRAM25;
 output Tile_X10Y10_BM_SRAM26;
 output Tile_X10Y10_BM_SRAM27;
 output Tile_X10Y10_BM_SRAM28;
 output Tile_X10Y10_BM_SRAM29;
 output Tile_X10Y10_BM_SRAM3;
 output Tile_X10Y10_BM_SRAM30;
 output Tile_X10Y10_BM_SRAM31;
 output Tile_X10Y10_BM_SRAM4;
 output Tile_X10Y10_BM_SRAM5;
 output Tile_X10Y10_BM_SRAM6;
 output Tile_X10Y10_BM_SRAM7;
 output Tile_X10Y10_BM_SRAM8;
 output Tile_X10Y10_BM_SRAM9;
 output Tile_X10Y10_CLK_SRAM;
 input Tile_X10Y10_CONFIGURED_top;
 output Tile_X10Y10_DIN_SRAM0;
 output Tile_X10Y10_DIN_SRAM1;
 output Tile_X10Y10_DIN_SRAM10;
 output Tile_X10Y10_DIN_SRAM11;
 output Tile_X10Y10_DIN_SRAM12;
 output Tile_X10Y10_DIN_SRAM13;
 output Tile_X10Y10_DIN_SRAM14;
 output Tile_X10Y10_DIN_SRAM15;
 output Tile_X10Y10_DIN_SRAM16;
 output Tile_X10Y10_DIN_SRAM17;
 output Tile_X10Y10_DIN_SRAM18;
 output Tile_X10Y10_DIN_SRAM19;
 output Tile_X10Y10_DIN_SRAM2;
 output Tile_X10Y10_DIN_SRAM20;
 output Tile_X10Y10_DIN_SRAM21;
 output Tile_X10Y10_DIN_SRAM22;
 output Tile_X10Y10_DIN_SRAM23;
 output Tile_X10Y10_DIN_SRAM24;
 output Tile_X10Y10_DIN_SRAM25;
 output Tile_X10Y10_DIN_SRAM26;
 output Tile_X10Y10_DIN_SRAM27;
 output Tile_X10Y10_DIN_SRAM28;
 output Tile_X10Y10_DIN_SRAM29;
 output Tile_X10Y10_DIN_SRAM3;
 output Tile_X10Y10_DIN_SRAM30;
 output Tile_X10Y10_DIN_SRAM31;
 output Tile_X10Y10_DIN_SRAM4;
 output Tile_X10Y10_DIN_SRAM5;
 output Tile_X10Y10_DIN_SRAM6;
 output Tile_X10Y10_DIN_SRAM7;
 output Tile_X10Y10_DIN_SRAM8;
 output Tile_X10Y10_DIN_SRAM9;
 input Tile_X10Y10_DOUT_SRAM0;
 input Tile_X10Y10_DOUT_SRAM1;
 input Tile_X10Y10_DOUT_SRAM10;
 input Tile_X10Y10_DOUT_SRAM11;
 input Tile_X10Y10_DOUT_SRAM12;
 input Tile_X10Y10_DOUT_SRAM13;
 input Tile_X10Y10_DOUT_SRAM14;
 input Tile_X10Y10_DOUT_SRAM15;
 input Tile_X10Y10_DOUT_SRAM16;
 input Tile_X10Y10_DOUT_SRAM17;
 input Tile_X10Y10_DOUT_SRAM18;
 input Tile_X10Y10_DOUT_SRAM19;
 input Tile_X10Y10_DOUT_SRAM2;
 input Tile_X10Y10_DOUT_SRAM20;
 input Tile_X10Y10_DOUT_SRAM21;
 input Tile_X10Y10_DOUT_SRAM22;
 input Tile_X10Y10_DOUT_SRAM23;
 input Tile_X10Y10_DOUT_SRAM24;
 input Tile_X10Y10_DOUT_SRAM25;
 input Tile_X10Y10_DOUT_SRAM26;
 input Tile_X10Y10_DOUT_SRAM27;
 input Tile_X10Y10_DOUT_SRAM28;
 input Tile_X10Y10_DOUT_SRAM29;
 input Tile_X10Y10_DOUT_SRAM3;
 input Tile_X10Y10_DOUT_SRAM30;
 input Tile_X10Y10_DOUT_SRAM31;
 input Tile_X10Y10_DOUT_SRAM4;
 input Tile_X10Y10_DOUT_SRAM5;
 input Tile_X10Y10_DOUT_SRAM6;
 input Tile_X10Y10_DOUT_SRAM7;
 input Tile_X10Y10_DOUT_SRAM8;
 input Tile_X10Y10_DOUT_SRAM9;
 output Tile_X10Y10_MEN_SRAM;
 output Tile_X10Y10_REN_SRAM;
 output Tile_X10Y10_TIE_HIGH_SRAM;
 output Tile_X10Y10_TIE_LOW_SRAM;
 output Tile_X10Y10_WEN_SRAM;
 output Tile_X10Y12_ADDR_SRAM0;
 output Tile_X10Y12_ADDR_SRAM1;
 output Tile_X10Y12_ADDR_SRAM2;
 output Tile_X10Y12_ADDR_SRAM3;
 output Tile_X10Y12_ADDR_SRAM4;
 output Tile_X10Y12_ADDR_SRAM5;
 output Tile_X10Y12_ADDR_SRAM6;
 output Tile_X10Y12_ADDR_SRAM7;
 output Tile_X10Y12_ADDR_SRAM8;
 output Tile_X10Y12_ADDR_SRAM9;
 output Tile_X10Y12_BM_SRAM0;
 output Tile_X10Y12_BM_SRAM1;
 output Tile_X10Y12_BM_SRAM10;
 output Tile_X10Y12_BM_SRAM11;
 output Tile_X10Y12_BM_SRAM12;
 output Tile_X10Y12_BM_SRAM13;
 output Tile_X10Y12_BM_SRAM14;
 output Tile_X10Y12_BM_SRAM15;
 output Tile_X10Y12_BM_SRAM16;
 output Tile_X10Y12_BM_SRAM17;
 output Tile_X10Y12_BM_SRAM18;
 output Tile_X10Y12_BM_SRAM19;
 output Tile_X10Y12_BM_SRAM2;
 output Tile_X10Y12_BM_SRAM20;
 output Tile_X10Y12_BM_SRAM21;
 output Tile_X10Y12_BM_SRAM22;
 output Tile_X10Y12_BM_SRAM23;
 output Tile_X10Y12_BM_SRAM24;
 output Tile_X10Y12_BM_SRAM25;
 output Tile_X10Y12_BM_SRAM26;
 output Tile_X10Y12_BM_SRAM27;
 output Tile_X10Y12_BM_SRAM28;
 output Tile_X10Y12_BM_SRAM29;
 output Tile_X10Y12_BM_SRAM3;
 output Tile_X10Y12_BM_SRAM30;
 output Tile_X10Y12_BM_SRAM31;
 output Tile_X10Y12_BM_SRAM4;
 output Tile_X10Y12_BM_SRAM5;
 output Tile_X10Y12_BM_SRAM6;
 output Tile_X10Y12_BM_SRAM7;
 output Tile_X10Y12_BM_SRAM8;
 output Tile_X10Y12_BM_SRAM9;
 output Tile_X10Y12_CLK_SRAM;
 input Tile_X10Y12_CONFIGURED_top;
 output Tile_X10Y12_DIN_SRAM0;
 output Tile_X10Y12_DIN_SRAM1;
 output Tile_X10Y12_DIN_SRAM10;
 output Tile_X10Y12_DIN_SRAM11;
 output Tile_X10Y12_DIN_SRAM12;
 output Tile_X10Y12_DIN_SRAM13;
 output Tile_X10Y12_DIN_SRAM14;
 output Tile_X10Y12_DIN_SRAM15;
 output Tile_X10Y12_DIN_SRAM16;
 output Tile_X10Y12_DIN_SRAM17;
 output Tile_X10Y12_DIN_SRAM18;
 output Tile_X10Y12_DIN_SRAM19;
 output Tile_X10Y12_DIN_SRAM2;
 output Tile_X10Y12_DIN_SRAM20;
 output Tile_X10Y12_DIN_SRAM21;
 output Tile_X10Y12_DIN_SRAM22;
 output Tile_X10Y12_DIN_SRAM23;
 output Tile_X10Y12_DIN_SRAM24;
 output Tile_X10Y12_DIN_SRAM25;
 output Tile_X10Y12_DIN_SRAM26;
 output Tile_X10Y12_DIN_SRAM27;
 output Tile_X10Y12_DIN_SRAM28;
 output Tile_X10Y12_DIN_SRAM29;
 output Tile_X10Y12_DIN_SRAM3;
 output Tile_X10Y12_DIN_SRAM30;
 output Tile_X10Y12_DIN_SRAM31;
 output Tile_X10Y12_DIN_SRAM4;
 output Tile_X10Y12_DIN_SRAM5;
 output Tile_X10Y12_DIN_SRAM6;
 output Tile_X10Y12_DIN_SRAM7;
 output Tile_X10Y12_DIN_SRAM8;
 output Tile_X10Y12_DIN_SRAM9;
 input Tile_X10Y12_DOUT_SRAM0;
 input Tile_X10Y12_DOUT_SRAM1;
 input Tile_X10Y12_DOUT_SRAM10;
 input Tile_X10Y12_DOUT_SRAM11;
 input Tile_X10Y12_DOUT_SRAM12;
 input Tile_X10Y12_DOUT_SRAM13;
 input Tile_X10Y12_DOUT_SRAM14;
 input Tile_X10Y12_DOUT_SRAM15;
 input Tile_X10Y12_DOUT_SRAM16;
 input Tile_X10Y12_DOUT_SRAM17;
 input Tile_X10Y12_DOUT_SRAM18;
 input Tile_X10Y12_DOUT_SRAM19;
 input Tile_X10Y12_DOUT_SRAM2;
 input Tile_X10Y12_DOUT_SRAM20;
 input Tile_X10Y12_DOUT_SRAM21;
 input Tile_X10Y12_DOUT_SRAM22;
 input Tile_X10Y12_DOUT_SRAM23;
 input Tile_X10Y12_DOUT_SRAM24;
 input Tile_X10Y12_DOUT_SRAM25;
 input Tile_X10Y12_DOUT_SRAM26;
 input Tile_X10Y12_DOUT_SRAM27;
 input Tile_X10Y12_DOUT_SRAM28;
 input Tile_X10Y12_DOUT_SRAM29;
 input Tile_X10Y12_DOUT_SRAM3;
 input Tile_X10Y12_DOUT_SRAM30;
 input Tile_X10Y12_DOUT_SRAM31;
 input Tile_X10Y12_DOUT_SRAM4;
 input Tile_X10Y12_DOUT_SRAM5;
 input Tile_X10Y12_DOUT_SRAM6;
 input Tile_X10Y12_DOUT_SRAM7;
 input Tile_X10Y12_DOUT_SRAM8;
 input Tile_X10Y12_DOUT_SRAM9;
 output Tile_X10Y12_MEN_SRAM;
 output Tile_X10Y12_REN_SRAM;
 output Tile_X10Y12_TIE_HIGH_SRAM;
 output Tile_X10Y12_TIE_LOW_SRAM;
 output Tile_X10Y12_WEN_SRAM;
 output Tile_X10Y14_ADDR_SRAM0;
 output Tile_X10Y14_ADDR_SRAM1;
 output Tile_X10Y14_ADDR_SRAM2;
 output Tile_X10Y14_ADDR_SRAM3;
 output Tile_X10Y14_ADDR_SRAM4;
 output Tile_X10Y14_ADDR_SRAM5;
 output Tile_X10Y14_ADDR_SRAM6;
 output Tile_X10Y14_ADDR_SRAM7;
 output Tile_X10Y14_ADDR_SRAM8;
 output Tile_X10Y14_ADDR_SRAM9;
 output Tile_X10Y14_BM_SRAM0;
 output Tile_X10Y14_BM_SRAM1;
 output Tile_X10Y14_BM_SRAM10;
 output Tile_X10Y14_BM_SRAM11;
 output Tile_X10Y14_BM_SRAM12;
 output Tile_X10Y14_BM_SRAM13;
 output Tile_X10Y14_BM_SRAM14;
 output Tile_X10Y14_BM_SRAM15;
 output Tile_X10Y14_BM_SRAM16;
 output Tile_X10Y14_BM_SRAM17;
 output Tile_X10Y14_BM_SRAM18;
 output Tile_X10Y14_BM_SRAM19;
 output Tile_X10Y14_BM_SRAM2;
 output Tile_X10Y14_BM_SRAM20;
 output Tile_X10Y14_BM_SRAM21;
 output Tile_X10Y14_BM_SRAM22;
 output Tile_X10Y14_BM_SRAM23;
 output Tile_X10Y14_BM_SRAM24;
 output Tile_X10Y14_BM_SRAM25;
 output Tile_X10Y14_BM_SRAM26;
 output Tile_X10Y14_BM_SRAM27;
 output Tile_X10Y14_BM_SRAM28;
 output Tile_X10Y14_BM_SRAM29;
 output Tile_X10Y14_BM_SRAM3;
 output Tile_X10Y14_BM_SRAM30;
 output Tile_X10Y14_BM_SRAM31;
 output Tile_X10Y14_BM_SRAM4;
 output Tile_X10Y14_BM_SRAM5;
 output Tile_X10Y14_BM_SRAM6;
 output Tile_X10Y14_BM_SRAM7;
 output Tile_X10Y14_BM_SRAM8;
 output Tile_X10Y14_BM_SRAM9;
 output Tile_X10Y14_CLK_SRAM;
 input Tile_X10Y14_CONFIGURED_top;
 output Tile_X10Y14_DIN_SRAM0;
 output Tile_X10Y14_DIN_SRAM1;
 output Tile_X10Y14_DIN_SRAM10;
 output Tile_X10Y14_DIN_SRAM11;
 output Tile_X10Y14_DIN_SRAM12;
 output Tile_X10Y14_DIN_SRAM13;
 output Tile_X10Y14_DIN_SRAM14;
 output Tile_X10Y14_DIN_SRAM15;
 output Tile_X10Y14_DIN_SRAM16;
 output Tile_X10Y14_DIN_SRAM17;
 output Tile_X10Y14_DIN_SRAM18;
 output Tile_X10Y14_DIN_SRAM19;
 output Tile_X10Y14_DIN_SRAM2;
 output Tile_X10Y14_DIN_SRAM20;
 output Tile_X10Y14_DIN_SRAM21;
 output Tile_X10Y14_DIN_SRAM22;
 output Tile_X10Y14_DIN_SRAM23;
 output Tile_X10Y14_DIN_SRAM24;
 output Tile_X10Y14_DIN_SRAM25;
 output Tile_X10Y14_DIN_SRAM26;
 output Tile_X10Y14_DIN_SRAM27;
 output Tile_X10Y14_DIN_SRAM28;
 output Tile_X10Y14_DIN_SRAM29;
 output Tile_X10Y14_DIN_SRAM3;
 output Tile_X10Y14_DIN_SRAM30;
 output Tile_X10Y14_DIN_SRAM31;
 output Tile_X10Y14_DIN_SRAM4;
 output Tile_X10Y14_DIN_SRAM5;
 output Tile_X10Y14_DIN_SRAM6;
 output Tile_X10Y14_DIN_SRAM7;
 output Tile_X10Y14_DIN_SRAM8;
 output Tile_X10Y14_DIN_SRAM9;
 input Tile_X10Y14_DOUT_SRAM0;
 input Tile_X10Y14_DOUT_SRAM1;
 input Tile_X10Y14_DOUT_SRAM10;
 input Tile_X10Y14_DOUT_SRAM11;
 input Tile_X10Y14_DOUT_SRAM12;
 input Tile_X10Y14_DOUT_SRAM13;
 input Tile_X10Y14_DOUT_SRAM14;
 input Tile_X10Y14_DOUT_SRAM15;
 input Tile_X10Y14_DOUT_SRAM16;
 input Tile_X10Y14_DOUT_SRAM17;
 input Tile_X10Y14_DOUT_SRAM18;
 input Tile_X10Y14_DOUT_SRAM19;
 input Tile_X10Y14_DOUT_SRAM2;
 input Tile_X10Y14_DOUT_SRAM20;
 input Tile_X10Y14_DOUT_SRAM21;
 input Tile_X10Y14_DOUT_SRAM22;
 input Tile_X10Y14_DOUT_SRAM23;
 input Tile_X10Y14_DOUT_SRAM24;
 input Tile_X10Y14_DOUT_SRAM25;
 input Tile_X10Y14_DOUT_SRAM26;
 input Tile_X10Y14_DOUT_SRAM27;
 input Tile_X10Y14_DOUT_SRAM28;
 input Tile_X10Y14_DOUT_SRAM29;
 input Tile_X10Y14_DOUT_SRAM3;
 input Tile_X10Y14_DOUT_SRAM30;
 input Tile_X10Y14_DOUT_SRAM31;
 input Tile_X10Y14_DOUT_SRAM4;
 input Tile_X10Y14_DOUT_SRAM5;
 input Tile_X10Y14_DOUT_SRAM6;
 input Tile_X10Y14_DOUT_SRAM7;
 input Tile_X10Y14_DOUT_SRAM8;
 input Tile_X10Y14_DOUT_SRAM9;
 output Tile_X10Y14_MEN_SRAM;
 output Tile_X10Y14_REN_SRAM;
 output Tile_X10Y14_TIE_HIGH_SRAM;
 output Tile_X10Y14_TIE_LOW_SRAM;
 output Tile_X10Y14_WEN_SRAM;
 output Tile_X10Y2_ADDR_SRAM0;
 output Tile_X10Y2_ADDR_SRAM1;
 output Tile_X10Y2_ADDR_SRAM2;
 output Tile_X10Y2_ADDR_SRAM3;
 output Tile_X10Y2_ADDR_SRAM4;
 output Tile_X10Y2_ADDR_SRAM5;
 output Tile_X10Y2_ADDR_SRAM6;
 output Tile_X10Y2_ADDR_SRAM7;
 output Tile_X10Y2_ADDR_SRAM8;
 output Tile_X10Y2_ADDR_SRAM9;
 output Tile_X10Y2_BM_SRAM0;
 output Tile_X10Y2_BM_SRAM1;
 output Tile_X10Y2_BM_SRAM10;
 output Tile_X10Y2_BM_SRAM11;
 output Tile_X10Y2_BM_SRAM12;
 output Tile_X10Y2_BM_SRAM13;
 output Tile_X10Y2_BM_SRAM14;
 output Tile_X10Y2_BM_SRAM15;
 output Tile_X10Y2_BM_SRAM16;
 output Tile_X10Y2_BM_SRAM17;
 output Tile_X10Y2_BM_SRAM18;
 output Tile_X10Y2_BM_SRAM19;
 output Tile_X10Y2_BM_SRAM2;
 output Tile_X10Y2_BM_SRAM20;
 output Tile_X10Y2_BM_SRAM21;
 output Tile_X10Y2_BM_SRAM22;
 output Tile_X10Y2_BM_SRAM23;
 output Tile_X10Y2_BM_SRAM24;
 output Tile_X10Y2_BM_SRAM25;
 output Tile_X10Y2_BM_SRAM26;
 output Tile_X10Y2_BM_SRAM27;
 output Tile_X10Y2_BM_SRAM28;
 output Tile_X10Y2_BM_SRAM29;
 output Tile_X10Y2_BM_SRAM3;
 output Tile_X10Y2_BM_SRAM30;
 output Tile_X10Y2_BM_SRAM31;
 output Tile_X10Y2_BM_SRAM4;
 output Tile_X10Y2_BM_SRAM5;
 output Tile_X10Y2_BM_SRAM6;
 output Tile_X10Y2_BM_SRAM7;
 output Tile_X10Y2_BM_SRAM8;
 output Tile_X10Y2_BM_SRAM9;
 output Tile_X10Y2_CLK_SRAM;
 input Tile_X10Y2_CONFIGURED_top;
 output Tile_X10Y2_DIN_SRAM0;
 output Tile_X10Y2_DIN_SRAM1;
 output Tile_X10Y2_DIN_SRAM10;
 output Tile_X10Y2_DIN_SRAM11;
 output Tile_X10Y2_DIN_SRAM12;
 output Tile_X10Y2_DIN_SRAM13;
 output Tile_X10Y2_DIN_SRAM14;
 output Tile_X10Y2_DIN_SRAM15;
 output Tile_X10Y2_DIN_SRAM16;
 output Tile_X10Y2_DIN_SRAM17;
 output Tile_X10Y2_DIN_SRAM18;
 output Tile_X10Y2_DIN_SRAM19;
 output Tile_X10Y2_DIN_SRAM2;
 output Tile_X10Y2_DIN_SRAM20;
 output Tile_X10Y2_DIN_SRAM21;
 output Tile_X10Y2_DIN_SRAM22;
 output Tile_X10Y2_DIN_SRAM23;
 output Tile_X10Y2_DIN_SRAM24;
 output Tile_X10Y2_DIN_SRAM25;
 output Tile_X10Y2_DIN_SRAM26;
 output Tile_X10Y2_DIN_SRAM27;
 output Tile_X10Y2_DIN_SRAM28;
 output Tile_X10Y2_DIN_SRAM29;
 output Tile_X10Y2_DIN_SRAM3;
 output Tile_X10Y2_DIN_SRAM30;
 output Tile_X10Y2_DIN_SRAM31;
 output Tile_X10Y2_DIN_SRAM4;
 output Tile_X10Y2_DIN_SRAM5;
 output Tile_X10Y2_DIN_SRAM6;
 output Tile_X10Y2_DIN_SRAM7;
 output Tile_X10Y2_DIN_SRAM8;
 output Tile_X10Y2_DIN_SRAM9;
 input Tile_X10Y2_DOUT_SRAM0;
 input Tile_X10Y2_DOUT_SRAM1;
 input Tile_X10Y2_DOUT_SRAM10;
 input Tile_X10Y2_DOUT_SRAM11;
 input Tile_X10Y2_DOUT_SRAM12;
 input Tile_X10Y2_DOUT_SRAM13;
 input Tile_X10Y2_DOUT_SRAM14;
 input Tile_X10Y2_DOUT_SRAM15;
 input Tile_X10Y2_DOUT_SRAM16;
 input Tile_X10Y2_DOUT_SRAM17;
 input Tile_X10Y2_DOUT_SRAM18;
 input Tile_X10Y2_DOUT_SRAM19;
 input Tile_X10Y2_DOUT_SRAM2;
 input Tile_X10Y2_DOUT_SRAM20;
 input Tile_X10Y2_DOUT_SRAM21;
 input Tile_X10Y2_DOUT_SRAM22;
 input Tile_X10Y2_DOUT_SRAM23;
 input Tile_X10Y2_DOUT_SRAM24;
 input Tile_X10Y2_DOUT_SRAM25;
 input Tile_X10Y2_DOUT_SRAM26;
 input Tile_X10Y2_DOUT_SRAM27;
 input Tile_X10Y2_DOUT_SRAM28;
 input Tile_X10Y2_DOUT_SRAM29;
 input Tile_X10Y2_DOUT_SRAM3;
 input Tile_X10Y2_DOUT_SRAM30;
 input Tile_X10Y2_DOUT_SRAM31;
 input Tile_X10Y2_DOUT_SRAM4;
 input Tile_X10Y2_DOUT_SRAM5;
 input Tile_X10Y2_DOUT_SRAM6;
 input Tile_X10Y2_DOUT_SRAM7;
 input Tile_X10Y2_DOUT_SRAM8;
 input Tile_X10Y2_DOUT_SRAM9;
 output Tile_X10Y2_MEN_SRAM;
 output Tile_X10Y2_REN_SRAM;
 output Tile_X10Y2_TIE_HIGH_SRAM;
 output Tile_X10Y2_TIE_LOW_SRAM;
 output Tile_X10Y2_WEN_SRAM;
 output Tile_X10Y4_ADDR_SRAM0;
 output Tile_X10Y4_ADDR_SRAM1;
 output Tile_X10Y4_ADDR_SRAM2;
 output Tile_X10Y4_ADDR_SRAM3;
 output Tile_X10Y4_ADDR_SRAM4;
 output Tile_X10Y4_ADDR_SRAM5;
 output Tile_X10Y4_ADDR_SRAM6;
 output Tile_X10Y4_ADDR_SRAM7;
 output Tile_X10Y4_ADDR_SRAM8;
 output Tile_X10Y4_ADDR_SRAM9;
 output Tile_X10Y4_BM_SRAM0;
 output Tile_X10Y4_BM_SRAM1;
 output Tile_X10Y4_BM_SRAM10;
 output Tile_X10Y4_BM_SRAM11;
 output Tile_X10Y4_BM_SRAM12;
 output Tile_X10Y4_BM_SRAM13;
 output Tile_X10Y4_BM_SRAM14;
 output Tile_X10Y4_BM_SRAM15;
 output Tile_X10Y4_BM_SRAM16;
 output Tile_X10Y4_BM_SRAM17;
 output Tile_X10Y4_BM_SRAM18;
 output Tile_X10Y4_BM_SRAM19;
 output Tile_X10Y4_BM_SRAM2;
 output Tile_X10Y4_BM_SRAM20;
 output Tile_X10Y4_BM_SRAM21;
 output Tile_X10Y4_BM_SRAM22;
 output Tile_X10Y4_BM_SRAM23;
 output Tile_X10Y4_BM_SRAM24;
 output Tile_X10Y4_BM_SRAM25;
 output Tile_X10Y4_BM_SRAM26;
 output Tile_X10Y4_BM_SRAM27;
 output Tile_X10Y4_BM_SRAM28;
 output Tile_X10Y4_BM_SRAM29;
 output Tile_X10Y4_BM_SRAM3;
 output Tile_X10Y4_BM_SRAM30;
 output Tile_X10Y4_BM_SRAM31;
 output Tile_X10Y4_BM_SRAM4;
 output Tile_X10Y4_BM_SRAM5;
 output Tile_X10Y4_BM_SRAM6;
 output Tile_X10Y4_BM_SRAM7;
 output Tile_X10Y4_BM_SRAM8;
 output Tile_X10Y4_BM_SRAM9;
 output Tile_X10Y4_CLK_SRAM;
 input Tile_X10Y4_CONFIGURED_top;
 output Tile_X10Y4_DIN_SRAM0;
 output Tile_X10Y4_DIN_SRAM1;
 output Tile_X10Y4_DIN_SRAM10;
 output Tile_X10Y4_DIN_SRAM11;
 output Tile_X10Y4_DIN_SRAM12;
 output Tile_X10Y4_DIN_SRAM13;
 output Tile_X10Y4_DIN_SRAM14;
 output Tile_X10Y4_DIN_SRAM15;
 output Tile_X10Y4_DIN_SRAM16;
 output Tile_X10Y4_DIN_SRAM17;
 output Tile_X10Y4_DIN_SRAM18;
 output Tile_X10Y4_DIN_SRAM19;
 output Tile_X10Y4_DIN_SRAM2;
 output Tile_X10Y4_DIN_SRAM20;
 output Tile_X10Y4_DIN_SRAM21;
 output Tile_X10Y4_DIN_SRAM22;
 output Tile_X10Y4_DIN_SRAM23;
 output Tile_X10Y4_DIN_SRAM24;
 output Tile_X10Y4_DIN_SRAM25;
 output Tile_X10Y4_DIN_SRAM26;
 output Tile_X10Y4_DIN_SRAM27;
 output Tile_X10Y4_DIN_SRAM28;
 output Tile_X10Y4_DIN_SRAM29;
 output Tile_X10Y4_DIN_SRAM3;
 output Tile_X10Y4_DIN_SRAM30;
 output Tile_X10Y4_DIN_SRAM31;
 output Tile_X10Y4_DIN_SRAM4;
 output Tile_X10Y4_DIN_SRAM5;
 output Tile_X10Y4_DIN_SRAM6;
 output Tile_X10Y4_DIN_SRAM7;
 output Tile_X10Y4_DIN_SRAM8;
 output Tile_X10Y4_DIN_SRAM9;
 input Tile_X10Y4_DOUT_SRAM0;
 input Tile_X10Y4_DOUT_SRAM1;
 input Tile_X10Y4_DOUT_SRAM10;
 input Tile_X10Y4_DOUT_SRAM11;
 input Tile_X10Y4_DOUT_SRAM12;
 input Tile_X10Y4_DOUT_SRAM13;
 input Tile_X10Y4_DOUT_SRAM14;
 input Tile_X10Y4_DOUT_SRAM15;
 input Tile_X10Y4_DOUT_SRAM16;
 input Tile_X10Y4_DOUT_SRAM17;
 input Tile_X10Y4_DOUT_SRAM18;
 input Tile_X10Y4_DOUT_SRAM19;
 input Tile_X10Y4_DOUT_SRAM2;
 input Tile_X10Y4_DOUT_SRAM20;
 input Tile_X10Y4_DOUT_SRAM21;
 input Tile_X10Y4_DOUT_SRAM22;
 input Tile_X10Y4_DOUT_SRAM23;
 input Tile_X10Y4_DOUT_SRAM24;
 input Tile_X10Y4_DOUT_SRAM25;
 input Tile_X10Y4_DOUT_SRAM26;
 input Tile_X10Y4_DOUT_SRAM27;
 input Tile_X10Y4_DOUT_SRAM28;
 input Tile_X10Y4_DOUT_SRAM29;
 input Tile_X10Y4_DOUT_SRAM3;
 input Tile_X10Y4_DOUT_SRAM30;
 input Tile_X10Y4_DOUT_SRAM31;
 input Tile_X10Y4_DOUT_SRAM4;
 input Tile_X10Y4_DOUT_SRAM5;
 input Tile_X10Y4_DOUT_SRAM6;
 input Tile_X10Y4_DOUT_SRAM7;
 input Tile_X10Y4_DOUT_SRAM8;
 input Tile_X10Y4_DOUT_SRAM9;
 output Tile_X10Y4_MEN_SRAM;
 output Tile_X10Y4_REN_SRAM;
 output Tile_X10Y4_TIE_HIGH_SRAM;
 output Tile_X10Y4_TIE_LOW_SRAM;
 output Tile_X10Y4_WEN_SRAM;
 output Tile_X10Y6_ADDR_SRAM0;
 output Tile_X10Y6_ADDR_SRAM1;
 output Tile_X10Y6_ADDR_SRAM2;
 output Tile_X10Y6_ADDR_SRAM3;
 output Tile_X10Y6_ADDR_SRAM4;
 output Tile_X10Y6_ADDR_SRAM5;
 output Tile_X10Y6_ADDR_SRAM6;
 output Tile_X10Y6_ADDR_SRAM7;
 output Tile_X10Y6_ADDR_SRAM8;
 output Tile_X10Y6_ADDR_SRAM9;
 output Tile_X10Y6_BM_SRAM0;
 output Tile_X10Y6_BM_SRAM1;
 output Tile_X10Y6_BM_SRAM10;
 output Tile_X10Y6_BM_SRAM11;
 output Tile_X10Y6_BM_SRAM12;
 output Tile_X10Y6_BM_SRAM13;
 output Tile_X10Y6_BM_SRAM14;
 output Tile_X10Y6_BM_SRAM15;
 output Tile_X10Y6_BM_SRAM16;
 output Tile_X10Y6_BM_SRAM17;
 output Tile_X10Y6_BM_SRAM18;
 output Tile_X10Y6_BM_SRAM19;
 output Tile_X10Y6_BM_SRAM2;
 output Tile_X10Y6_BM_SRAM20;
 output Tile_X10Y6_BM_SRAM21;
 output Tile_X10Y6_BM_SRAM22;
 output Tile_X10Y6_BM_SRAM23;
 output Tile_X10Y6_BM_SRAM24;
 output Tile_X10Y6_BM_SRAM25;
 output Tile_X10Y6_BM_SRAM26;
 output Tile_X10Y6_BM_SRAM27;
 output Tile_X10Y6_BM_SRAM28;
 output Tile_X10Y6_BM_SRAM29;
 output Tile_X10Y6_BM_SRAM3;
 output Tile_X10Y6_BM_SRAM30;
 output Tile_X10Y6_BM_SRAM31;
 output Tile_X10Y6_BM_SRAM4;
 output Tile_X10Y6_BM_SRAM5;
 output Tile_X10Y6_BM_SRAM6;
 output Tile_X10Y6_BM_SRAM7;
 output Tile_X10Y6_BM_SRAM8;
 output Tile_X10Y6_BM_SRAM9;
 output Tile_X10Y6_CLK_SRAM;
 input Tile_X10Y6_CONFIGURED_top;
 output Tile_X10Y6_DIN_SRAM0;
 output Tile_X10Y6_DIN_SRAM1;
 output Tile_X10Y6_DIN_SRAM10;
 output Tile_X10Y6_DIN_SRAM11;
 output Tile_X10Y6_DIN_SRAM12;
 output Tile_X10Y6_DIN_SRAM13;
 output Tile_X10Y6_DIN_SRAM14;
 output Tile_X10Y6_DIN_SRAM15;
 output Tile_X10Y6_DIN_SRAM16;
 output Tile_X10Y6_DIN_SRAM17;
 output Tile_X10Y6_DIN_SRAM18;
 output Tile_X10Y6_DIN_SRAM19;
 output Tile_X10Y6_DIN_SRAM2;
 output Tile_X10Y6_DIN_SRAM20;
 output Tile_X10Y6_DIN_SRAM21;
 output Tile_X10Y6_DIN_SRAM22;
 output Tile_X10Y6_DIN_SRAM23;
 output Tile_X10Y6_DIN_SRAM24;
 output Tile_X10Y6_DIN_SRAM25;
 output Tile_X10Y6_DIN_SRAM26;
 output Tile_X10Y6_DIN_SRAM27;
 output Tile_X10Y6_DIN_SRAM28;
 output Tile_X10Y6_DIN_SRAM29;
 output Tile_X10Y6_DIN_SRAM3;
 output Tile_X10Y6_DIN_SRAM30;
 output Tile_X10Y6_DIN_SRAM31;
 output Tile_X10Y6_DIN_SRAM4;
 output Tile_X10Y6_DIN_SRAM5;
 output Tile_X10Y6_DIN_SRAM6;
 output Tile_X10Y6_DIN_SRAM7;
 output Tile_X10Y6_DIN_SRAM8;
 output Tile_X10Y6_DIN_SRAM9;
 input Tile_X10Y6_DOUT_SRAM0;
 input Tile_X10Y6_DOUT_SRAM1;
 input Tile_X10Y6_DOUT_SRAM10;
 input Tile_X10Y6_DOUT_SRAM11;
 input Tile_X10Y6_DOUT_SRAM12;
 input Tile_X10Y6_DOUT_SRAM13;
 input Tile_X10Y6_DOUT_SRAM14;
 input Tile_X10Y6_DOUT_SRAM15;
 input Tile_X10Y6_DOUT_SRAM16;
 input Tile_X10Y6_DOUT_SRAM17;
 input Tile_X10Y6_DOUT_SRAM18;
 input Tile_X10Y6_DOUT_SRAM19;
 input Tile_X10Y6_DOUT_SRAM2;
 input Tile_X10Y6_DOUT_SRAM20;
 input Tile_X10Y6_DOUT_SRAM21;
 input Tile_X10Y6_DOUT_SRAM22;
 input Tile_X10Y6_DOUT_SRAM23;
 input Tile_X10Y6_DOUT_SRAM24;
 input Tile_X10Y6_DOUT_SRAM25;
 input Tile_X10Y6_DOUT_SRAM26;
 input Tile_X10Y6_DOUT_SRAM27;
 input Tile_X10Y6_DOUT_SRAM28;
 input Tile_X10Y6_DOUT_SRAM29;
 input Tile_X10Y6_DOUT_SRAM3;
 input Tile_X10Y6_DOUT_SRAM30;
 input Tile_X10Y6_DOUT_SRAM31;
 input Tile_X10Y6_DOUT_SRAM4;
 input Tile_X10Y6_DOUT_SRAM5;
 input Tile_X10Y6_DOUT_SRAM6;
 input Tile_X10Y6_DOUT_SRAM7;
 input Tile_X10Y6_DOUT_SRAM8;
 input Tile_X10Y6_DOUT_SRAM9;
 output Tile_X10Y6_MEN_SRAM;
 output Tile_X10Y6_REN_SRAM;
 output Tile_X10Y6_TIE_HIGH_SRAM;
 output Tile_X10Y6_TIE_LOW_SRAM;
 output Tile_X10Y6_WEN_SRAM;
 output Tile_X10Y8_ADDR_SRAM0;
 output Tile_X10Y8_ADDR_SRAM1;
 output Tile_X10Y8_ADDR_SRAM2;
 output Tile_X10Y8_ADDR_SRAM3;
 output Tile_X10Y8_ADDR_SRAM4;
 output Tile_X10Y8_ADDR_SRAM5;
 output Tile_X10Y8_ADDR_SRAM6;
 output Tile_X10Y8_ADDR_SRAM7;
 output Tile_X10Y8_ADDR_SRAM8;
 output Tile_X10Y8_ADDR_SRAM9;
 output Tile_X10Y8_BM_SRAM0;
 output Tile_X10Y8_BM_SRAM1;
 output Tile_X10Y8_BM_SRAM10;
 output Tile_X10Y8_BM_SRAM11;
 output Tile_X10Y8_BM_SRAM12;
 output Tile_X10Y8_BM_SRAM13;
 output Tile_X10Y8_BM_SRAM14;
 output Tile_X10Y8_BM_SRAM15;
 output Tile_X10Y8_BM_SRAM16;
 output Tile_X10Y8_BM_SRAM17;
 output Tile_X10Y8_BM_SRAM18;
 output Tile_X10Y8_BM_SRAM19;
 output Tile_X10Y8_BM_SRAM2;
 output Tile_X10Y8_BM_SRAM20;
 output Tile_X10Y8_BM_SRAM21;
 output Tile_X10Y8_BM_SRAM22;
 output Tile_X10Y8_BM_SRAM23;
 output Tile_X10Y8_BM_SRAM24;
 output Tile_X10Y8_BM_SRAM25;
 output Tile_X10Y8_BM_SRAM26;
 output Tile_X10Y8_BM_SRAM27;
 output Tile_X10Y8_BM_SRAM28;
 output Tile_X10Y8_BM_SRAM29;
 output Tile_X10Y8_BM_SRAM3;
 output Tile_X10Y8_BM_SRAM30;
 output Tile_X10Y8_BM_SRAM31;
 output Tile_X10Y8_BM_SRAM4;
 output Tile_X10Y8_BM_SRAM5;
 output Tile_X10Y8_BM_SRAM6;
 output Tile_X10Y8_BM_SRAM7;
 output Tile_X10Y8_BM_SRAM8;
 output Tile_X10Y8_BM_SRAM9;
 output Tile_X10Y8_CLK_SRAM;
 input Tile_X10Y8_CONFIGURED_top;
 output Tile_X10Y8_DIN_SRAM0;
 output Tile_X10Y8_DIN_SRAM1;
 output Tile_X10Y8_DIN_SRAM10;
 output Tile_X10Y8_DIN_SRAM11;
 output Tile_X10Y8_DIN_SRAM12;
 output Tile_X10Y8_DIN_SRAM13;
 output Tile_X10Y8_DIN_SRAM14;
 output Tile_X10Y8_DIN_SRAM15;
 output Tile_X10Y8_DIN_SRAM16;
 output Tile_X10Y8_DIN_SRAM17;
 output Tile_X10Y8_DIN_SRAM18;
 output Tile_X10Y8_DIN_SRAM19;
 output Tile_X10Y8_DIN_SRAM2;
 output Tile_X10Y8_DIN_SRAM20;
 output Tile_X10Y8_DIN_SRAM21;
 output Tile_X10Y8_DIN_SRAM22;
 output Tile_X10Y8_DIN_SRAM23;
 output Tile_X10Y8_DIN_SRAM24;
 output Tile_X10Y8_DIN_SRAM25;
 output Tile_X10Y8_DIN_SRAM26;
 output Tile_X10Y8_DIN_SRAM27;
 output Tile_X10Y8_DIN_SRAM28;
 output Tile_X10Y8_DIN_SRAM29;
 output Tile_X10Y8_DIN_SRAM3;
 output Tile_X10Y8_DIN_SRAM30;
 output Tile_X10Y8_DIN_SRAM31;
 output Tile_X10Y8_DIN_SRAM4;
 output Tile_X10Y8_DIN_SRAM5;
 output Tile_X10Y8_DIN_SRAM6;
 output Tile_X10Y8_DIN_SRAM7;
 output Tile_X10Y8_DIN_SRAM8;
 output Tile_X10Y8_DIN_SRAM9;
 input Tile_X10Y8_DOUT_SRAM0;
 input Tile_X10Y8_DOUT_SRAM1;
 input Tile_X10Y8_DOUT_SRAM10;
 input Tile_X10Y8_DOUT_SRAM11;
 input Tile_X10Y8_DOUT_SRAM12;
 input Tile_X10Y8_DOUT_SRAM13;
 input Tile_X10Y8_DOUT_SRAM14;
 input Tile_X10Y8_DOUT_SRAM15;
 input Tile_X10Y8_DOUT_SRAM16;
 input Tile_X10Y8_DOUT_SRAM17;
 input Tile_X10Y8_DOUT_SRAM18;
 input Tile_X10Y8_DOUT_SRAM19;
 input Tile_X10Y8_DOUT_SRAM2;
 input Tile_X10Y8_DOUT_SRAM20;
 input Tile_X10Y8_DOUT_SRAM21;
 input Tile_X10Y8_DOUT_SRAM22;
 input Tile_X10Y8_DOUT_SRAM23;
 input Tile_X10Y8_DOUT_SRAM24;
 input Tile_X10Y8_DOUT_SRAM25;
 input Tile_X10Y8_DOUT_SRAM26;
 input Tile_X10Y8_DOUT_SRAM27;
 input Tile_X10Y8_DOUT_SRAM28;
 input Tile_X10Y8_DOUT_SRAM29;
 input Tile_X10Y8_DOUT_SRAM3;
 input Tile_X10Y8_DOUT_SRAM30;
 input Tile_X10Y8_DOUT_SRAM31;
 input Tile_X10Y8_DOUT_SRAM4;
 input Tile_X10Y8_DOUT_SRAM5;
 input Tile_X10Y8_DOUT_SRAM6;
 input Tile_X10Y8_DOUT_SRAM7;
 input Tile_X10Y8_DOUT_SRAM8;
 input Tile_X10Y8_DOUT_SRAM9;
 output Tile_X10Y8_MEN_SRAM;
 output Tile_X10Y8_REN_SRAM;
 output Tile_X10Y8_TIE_HIGH_SRAM;
 output Tile_X10Y8_TIE_LOW_SRAM;
 output Tile_X10Y8_WEN_SRAM;
 output Tile_X1Y0_A_I_top;
 input Tile_X1Y0_A_O_top;
 output Tile_X1Y0_A_T_top;
 output Tile_X1Y0_A_config_C_bit0;
 output Tile_X1Y0_A_config_C_bit1;
 output Tile_X1Y0_A_config_C_bit2;
 output Tile_X1Y0_A_config_C_bit3;
 output Tile_X1Y0_B_I_top;
 input Tile_X1Y0_B_O_top;
 output Tile_X1Y0_B_T_top;
 output Tile_X1Y0_B_config_C_bit0;
 output Tile_X1Y0_B_config_C_bit1;
 output Tile_X1Y0_B_config_C_bit2;
 output Tile_X1Y0_B_config_C_bit3;
 output Tile_X2Y0_A_I_top;
 input Tile_X2Y0_A_O_top;
 output Tile_X2Y0_A_T_top;
 output Tile_X2Y0_A_config_C_bit0;
 output Tile_X2Y0_A_config_C_bit1;
 output Tile_X2Y0_A_config_C_bit2;
 output Tile_X2Y0_A_config_C_bit3;
 output Tile_X2Y0_B_I_top;
 input Tile_X2Y0_B_O_top;
 output Tile_X2Y0_B_T_top;
 output Tile_X2Y0_B_config_C_bit0;
 output Tile_X2Y0_B_config_C_bit1;
 output Tile_X2Y0_B_config_C_bit2;
 output Tile_X2Y0_B_config_C_bit3;
 output Tile_X2Y15_BOOT_top;
 input Tile_X2Y15_CONFIGURED_top;
 input Tile_X2Y15_RESET_top;
 output Tile_X2Y15_SLOT_top0;
 output Tile_X2Y15_SLOT_top1;
 output Tile_X2Y15_SLOT_top2;
 output Tile_X2Y15_SLOT_top3;
 input Tile_X3Y15_CONFIGURED_top;
 output Tile_X3Y15_IRQ_top0;
 output Tile_X3Y15_IRQ_top1;
 output Tile_X3Y15_IRQ_top2;
 output Tile_X3Y15_IRQ_top3;
 output Tile_X5Y15_I_top0;
 output Tile_X5Y15_I_top1;
 output Tile_X5Y15_I_top10;
 output Tile_X5Y15_I_top11;
 output Tile_X5Y15_I_top12;
 output Tile_X5Y15_I_top13;
 output Tile_X5Y15_I_top14;
 output Tile_X5Y15_I_top15;
 output Tile_X5Y15_I_top2;
 output Tile_X5Y15_I_top3;
 output Tile_X5Y15_I_top4;
 output Tile_X5Y15_I_top5;
 output Tile_X5Y15_I_top6;
 output Tile_X5Y15_I_top7;
 output Tile_X5Y15_I_top8;
 output Tile_X5Y15_I_top9;
 input Tile_X5Y15_O_top0;
 input Tile_X5Y15_O_top1;
 input Tile_X5Y15_O_top10;
 input Tile_X5Y15_O_top11;
 input Tile_X5Y15_O_top12;
 input Tile_X5Y15_O_top13;
 input Tile_X5Y15_O_top14;
 input Tile_X5Y15_O_top15;
 input Tile_X5Y15_O_top2;
 input Tile_X5Y15_O_top3;
 input Tile_X5Y15_O_top4;
 input Tile_X5Y15_O_top5;
 input Tile_X5Y15_O_top6;
 input Tile_X5Y15_O_top7;
 input Tile_X5Y15_O_top8;
 input Tile_X5Y15_O_top9;
 output Tile_X6Y15_I_top0;
 output Tile_X6Y15_I_top1;
 output Tile_X6Y15_I_top10;
 output Tile_X6Y15_I_top11;
 output Tile_X6Y15_I_top12;
 output Tile_X6Y15_I_top13;
 output Tile_X6Y15_I_top14;
 output Tile_X6Y15_I_top15;
 output Tile_X6Y15_I_top2;
 output Tile_X6Y15_I_top3;
 output Tile_X6Y15_I_top4;
 output Tile_X6Y15_I_top5;
 output Tile_X6Y15_I_top6;
 output Tile_X6Y15_I_top7;
 output Tile_X6Y15_I_top8;
 output Tile_X6Y15_I_top9;
 input Tile_X6Y15_O_top0;
 input Tile_X6Y15_O_top1;
 input Tile_X6Y15_O_top10;
 input Tile_X6Y15_O_top11;
 input Tile_X6Y15_O_top12;
 input Tile_X6Y15_O_top13;
 input Tile_X6Y15_O_top14;
 input Tile_X6Y15_O_top15;
 input Tile_X6Y15_O_top2;
 input Tile_X6Y15_O_top3;
 input Tile_X6Y15_O_top4;
 input Tile_X6Y15_O_top5;
 input Tile_X6Y15_O_top6;
 input Tile_X6Y15_O_top7;
 input Tile_X6Y15_O_top8;
 input Tile_X6Y15_O_top9;
 output Tile_X8Y15_I_top0;
 output Tile_X8Y15_I_top1;
 output Tile_X8Y15_I_top10;
 output Tile_X8Y15_I_top11;
 output Tile_X8Y15_I_top12;
 output Tile_X8Y15_I_top13;
 output Tile_X8Y15_I_top14;
 output Tile_X8Y15_I_top15;
 output Tile_X8Y15_I_top2;
 output Tile_X8Y15_I_top3;
 output Tile_X8Y15_I_top4;
 output Tile_X8Y15_I_top5;
 output Tile_X8Y15_I_top6;
 output Tile_X8Y15_I_top7;
 output Tile_X8Y15_I_top8;
 output Tile_X8Y15_I_top9;
 input Tile_X8Y15_O_top0;
 input Tile_X8Y15_O_top1;
 input Tile_X8Y15_O_top10;
 input Tile_X8Y15_O_top11;
 input Tile_X8Y15_O_top12;
 input Tile_X8Y15_O_top13;
 input Tile_X8Y15_O_top14;
 input Tile_X8Y15_O_top15;
 input Tile_X8Y15_O_top2;
 input Tile_X8Y15_O_top3;
 input Tile_X8Y15_O_top4;
 input Tile_X8Y15_O_top5;
 input Tile_X8Y15_O_top6;
 input Tile_X8Y15_O_top7;
 input Tile_X8Y15_O_top8;
 input Tile_X8Y15_O_top9;
 output Tile_X9Y15_I_top0;
 output Tile_X9Y15_I_top1;
 output Tile_X9Y15_I_top10;
 output Tile_X9Y15_I_top11;
 output Tile_X9Y15_I_top12;
 output Tile_X9Y15_I_top13;
 output Tile_X9Y15_I_top14;
 output Tile_X9Y15_I_top15;
 output Tile_X9Y15_I_top2;
 output Tile_X9Y15_I_top3;
 output Tile_X9Y15_I_top4;
 output Tile_X9Y15_I_top5;
 output Tile_X9Y15_I_top6;
 output Tile_X9Y15_I_top7;
 output Tile_X9Y15_I_top8;
 output Tile_X9Y15_I_top9;
 input Tile_X9Y15_O_top0;
 input Tile_X9Y15_O_top1;
 input Tile_X9Y15_O_top10;
 input Tile_X9Y15_O_top11;
 input Tile_X9Y15_O_top12;
 input Tile_X9Y15_O_top13;
 input Tile_X9Y15_O_top14;
 input Tile_X9Y15_O_top15;
 input Tile_X9Y15_O_top2;
 input Tile_X9Y15_O_top3;
 input Tile_X9Y15_O_top4;
 input Tile_X9Y15_O_top5;
 input Tile_X9Y15_O_top6;
 input Tile_X9Y15_O_top7;
 input Tile_X9Y15_O_top8;
 input Tile_X9Y15_O_top9;
 input UserCLK;
 inout VPWR;
 inout VGND;
 input [511:0] FrameData;
 input [219:0] FrameStrobe;

 wire \Tile_X0Y10_E1BEG[0] ;
 wire \Tile_X0Y10_E1BEG[1] ;
 wire \Tile_X0Y10_E1BEG[2] ;
 wire \Tile_X0Y10_E1BEG[3] ;
 wire \Tile_X0Y10_E2BEG[0] ;
 wire \Tile_X0Y10_E2BEG[1] ;
 wire \Tile_X0Y10_E2BEG[2] ;
 wire \Tile_X0Y10_E2BEG[3] ;
 wire \Tile_X0Y10_E2BEG[4] ;
 wire \Tile_X0Y10_E2BEG[5] ;
 wire \Tile_X0Y10_E2BEG[6] ;
 wire \Tile_X0Y10_E2BEG[7] ;
 wire \Tile_X0Y10_E2BEGb[0] ;
 wire \Tile_X0Y10_E2BEGb[1] ;
 wire \Tile_X0Y10_E2BEGb[2] ;
 wire \Tile_X0Y10_E2BEGb[3] ;
 wire \Tile_X0Y10_E2BEGb[4] ;
 wire \Tile_X0Y10_E2BEGb[5] ;
 wire \Tile_X0Y10_E2BEGb[6] ;
 wire \Tile_X0Y10_E2BEGb[7] ;
 wire \Tile_X0Y10_E6BEG[0] ;
 wire \Tile_X0Y10_E6BEG[10] ;
 wire \Tile_X0Y10_E6BEG[11] ;
 wire \Tile_X0Y10_E6BEG[1] ;
 wire \Tile_X0Y10_E6BEG[2] ;
 wire \Tile_X0Y10_E6BEG[3] ;
 wire \Tile_X0Y10_E6BEG[4] ;
 wire \Tile_X0Y10_E6BEG[5] ;
 wire \Tile_X0Y10_E6BEG[6] ;
 wire \Tile_X0Y10_E6BEG[7] ;
 wire \Tile_X0Y10_E6BEG[8] ;
 wire \Tile_X0Y10_E6BEG[9] ;
 wire \Tile_X0Y10_EE4BEG[0] ;
 wire \Tile_X0Y10_EE4BEG[10] ;
 wire \Tile_X0Y10_EE4BEG[11] ;
 wire \Tile_X0Y10_EE4BEG[12] ;
 wire \Tile_X0Y10_EE4BEG[13] ;
 wire \Tile_X0Y10_EE4BEG[14] ;
 wire \Tile_X0Y10_EE4BEG[15] ;
 wire \Tile_X0Y10_EE4BEG[1] ;
 wire \Tile_X0Y10_EE4BEG[2] ;
 wire \Tile_X0Y10_EE4BEG[3] ;
 wire \Tile_X0Y10_EE4BEG[4] ;
 wire \Tile_X0Y10_EE4BEG[5] ;
 wire \Tile_X0Y10_EE4BEG[6] ;
 wire \Tile_X0Y10_EE4BEG[7] ;
 wire \Tile_X0Y10_EE4BEG[8] ;
 wire \Tile_X0Y10_EE4BEG[9] ;
 wire \Tile_X0Y10_FrameData_O[0] ;
 wire \Tile_X0Y10_FrameData_O[10] ;
 wire \Tile_X0Y10_FrameData_O[11] ;
 wire \Tile_X0Y10_FrameData_O[12] ;
 wire \Tile_X0Y10_FrameData_O[13] ;
 wire \Tile_X0Y10_FrameData_O[14] ;
 wire \Tile_X0Y10_FrameData_O[15] ;
 wire \Tile_X0Y10_FrameData_O[16] ;
 wire \Tile_X0Y10_FrameData_O[17] ;
 wire \Tile_X0Y10_FrameData_O[18] ;
 wire \Tile_X0Y10_FrameData_O[19] ;
 wire \Tile_X0Y10_FrameData_O[1] ;
 wire \Tile_X0Y10_FrameData_O[20] ;
 wire \Tile_X0Y10_FrameData_O[21] ;
 wire \Tile_X0Y10_FrameData_O[22] ;
 wire \Tile_X0Y10_FrameData_O[23] ;
 wire \Tile_X0Y10_FrameData_O[24] ;
 wire \Tile_X0Y10_FrameData_O[25] ;
 wire \Tile_X0Y10_FrameData_O[26] ;
 wire \Tile_X0Y10_FrameData_O[27] ;
 wire \Tile_X0Y10_FrameData_O[28] ;
 wire \Tile_X0Y10_FrameData_O[29] ;
 wire \Tile_X0Y10_FrameData_O[2] ;
 wire \Tile_X0Y10_FrameData_O[30] ;
 wire \Tile_X0Y10_FrameData_O[31] ;
 wire \Tile_X0Y10_FrameData_O[3] ;
 wire \Tile_X0Y10_FrameData_O[4] ;
 wire \Tile_X0Y10_FrameData_O[5] ;
 wire \Tile_X0Y10_FrameData_O[6] ;
 wire \Tile_X0Y10_FrameData_O[7] ;
 wire \Tile_X0Y10_FrameData_O[8] ;
 wire \Tile_X0Y10_FrameData_O[9] ;
 wire \Tile_X0Y10_FrameStrobe_O[0] ;
 wire \Tile_X0Y10_FrameStrobe_O[10] ;
 wire \Tile_X0Y10_FrameStrobe_O[11] ;
 wire \Tile_X0Y10_FrameStrobe_O[12] ;
 wire \Tile_X0Y10_FrameStrobe_O[13] ;
 wire \Tile_X0Y10_FrameStrobe_O[14] ;
 wire \Tile_X0Y10_FrameStrobe_O[15] ;
 wire \Tile_X0Y10_FrameStrobe_O[16] ;
 wire \Tile_X0Y10_FrameStrobe_O[17] ;
 wire \Tile_X0Y10_FrameStrobe_O[18] ;
 wire \Tile_X0Y10_FrameStrobe_O[19] ;
 wire \Tile_X0Y10_FrameStrobe_O[1] ;
 wire \Tile_X0Y10_FrameStrobe_O[2] ;
 wire \Tile_X0Y10_FrameStrobe_O[3] ;
 wire \Tile_X0Y10_FrameStrobe_O[4] ;
 wire \Tile_X0Y10_FrameStrobe_O[5] ;
 wire \Tile_X0Y10_FrameStrobe_O[6] ;
 wire \Tile_X0Y10_FrameStrobe_O[7] ;
 wire \Tile_X0Y10_FrameStrobe_O[8] ;
 wire \Tile_X0Y10_FrameStrobe_O[9] ;
 wire Tile_X0Y10_UserCLKo;
 wire \Tile_X0Y11_E1BEG[0] ;
 wire \Tile_X0Y11_E1BEG[1] ;
 wire \Tile_X0Y11_E1BEG[2] ;
 wire \Tile_X0Y11_E1BEG[3] ;
 wire \Tile_X0Y11_E2BEG[0] ;
 wire \Tile_X0Y11_E2BEG[1] ;
 wire \Tile_X0Y11_E2BEG[2] ;
 wire \Tile_X0Y11_E2BEG[3] ;
 wire \Tile_X0Y11_E2BEG[4] ;
 wire \Tile_X0Y11_E2BEG[5] ;
 wire \Tile_X0Y11_E2BEG[6] ;
 wire \Tile_X0Y11_E2BEG[7] ;
 wire \Tile_X0Y11_E2BEGb[0] ;
 wire \Tile_X0Y11_E2BEGb[1] ;
 wire \Tile_X0Y11_E2BEGb[2] ;
 wire \Tile_X0Y11_E2BEGb[3] ;
 wire \Tile_X0Y11_E2BEGb[4] ;
 wire \Tile_X0Y11_E2BEGb[5] ;
 wire \Tile_X0Y11_E2BEGb[6] ;
 wire \Tile_X0Y11_E2BEGb[7] ;
 wire \Tile_X0Y11_E6BEG[0] ;
 wire \Tile_X0Y11_E6BEG[10] ;
 wire \Tile_X0Y11_E6BEG[11] ;
 wire \Tile_X0Y11_E6BEG[1] ;
 wire \Tile_X0Y11_E6BEG[2] ;
 wire \Tile_X0Y11_E6BEG[3] ;
 wire \Tile_X0Y11_E6BEG[4] ;
 wire \Tile_X0Y11_E6BEG[5] ;
 wire \Tile_X0Y11_E6BEG[6] ;
 wire \Tile_X0Y11_E6BEG[7] ;
 wire \Tile_X0Y11_E6BEG[8] ;
 wire \Tile_X0Y11_E6BEG[9] ;
 wire \Tile_X0Y11_EE4BEG[0] ;
 wire \Tile_X0Y11_EE4BEG[10] ;
 wire \Tile_X0Y11_EE4BEG[11] ;
 wire \Tile_X0Y11_EE4BEG[12] ;
 wire \Tile_X0Y11_EE4BEG[13] ;
 wire \Tile_X0Y11_EE4BEG[14] ;
 wire \Tile_X0Y11_EE4BEG[15] ;
 wire \Tile_X0Y11_EE4BEG[1] ;
 wire \Tile_X0Y11_EE4BEG[2] ;
 wire \Tile_X0Y11_EE4BEG[3] ;
 wire \Tile_X0Y11_EE4BEG[4] ;
 wire \Tile_X0Y11_EE4BEG[5] ;
 wire \Tile_X0Y11_EE4BEG[6] ;
 wire \Tile_X0Y11_EE4BEG[7] ;
 wire \Tile_X0Y11_EE4BEG[8] ;
 wire \Tile_X0Y11_EE4BEG[9] ;
 wire \Tile_X0Y11_FrameData_O[0] ;
 wire \Tile_X0Y11_FrameData_O[10] ;
 wire \Tile_X0Y11_FrameData_O[11] ;
 wire \Tile_X0Y11_FrameData_O[12] ;
 wire \Tile_X0Y11_FrameData_O[13] ;
 wire \Tile_X0Y11_FrameData_O[14] ;
 wire \Tile_X0Y11_FrameData_O[15] ;
 wire \Tile_X0Y11_FrameData_O[16] ;
 wire \Tile_X0Y11_FrameData_O[17] ;
 wire \Tile_X0Y11_FrameData_O[18] ;
 wire \Tile_X0Y11_FrameData_O[19] ;
 wire \Tile_X0Y11_FrameData_O[1] ;
 wire \Tile_X0Y11_FrameData_O[20] ;
 wire \Tile_X0Y11_FrameData_O[21] ;
 wire \Tile_X0Y11_FrameData_O[22] ;
 wire \Tile_X0Y11_FrameData_O[23] ;
 wire \Tile_X0Y11_FrameData_O[24] ;
 wire \Tile_X0Y11_FrameData_O[25] ;
 wire \Tile_X0Y11_FrameData_O[26] ;
 wire \Tile_X0Y11_FrameData_O[27] ;
 wire \Tile_X0Y11_FrameData_O[28] ;
 wire \Tile_X0Y11_FrameData_O[29] ;
 wire \Tile_X0Y11_FrameData_O[2] ;
 wire \Tile_X0Y11_FrameData_O[30] ;
 wire \Tile_X0Y11_FrameData_O[31] ;
 wire \Tile_X0Y11_FrameData_O[3] ;
 wire \Tile_X0Y11_FrameData_O[4] ;
 wire \Tile_X0Y11_FrameData_O[5] ;
 wire \Tile_X0Y11_FrameData_O[6] ;
 wire \Tile_X0Y11_FrameData_O[7] ;
 wire \Tile_X0Y11_FrameData_O[8] ;
 wire \Tile_X0Y11_FrameData_O[9] ;
 wire \Tile_X0Y11_FrameStrobe_O[0] ;
 wire \Tile_X0Y11_FrameStrobe_O[10] ;
 wire \Tile_X0Y11_FrameStrobe_O[11] ;
 wire \Tile_X0Y11_FrameStrobe_O[12] ;
 wire \Tile_X0Y11_FrameStrobe_O[13] ;
 wire \Tile_X0Y11_FrameStrobe_O[14] ;
 wire \Tile_X0Y11_FrameStrobe_O[15] ;
 wire \Tile_X0Y11_FrameStrobe_O[16] ;
 wire \Tile_X0Y11_FrameStrobe_O[17] ;
 wire \Tile_X0Y11_FrameStrobe_O[18] ;
 wire \Tile_X0Y11_FrameStrobe_O[19] ;
 wire \Tile_X0Y11_FrameStrobe_O[1] ;
 wire \Tile_X0Y11_FrameStrobe_O[2] ;
 wire \Tile_X0Y11_FrameStrobe_O[3] ;
 wire \Tile_X0Y11_FrameStrobe_O[4] ;
 wire \Tile_X0Y11_FrameStrobe_O[5] ;
 wire \Tile_X0Y11_FrameStrobe_O[6] ;
 wire \Tile_X0Y11_FrameStrobe_O[7] ;
 wire \Tile_X0Y11_FrameStrobe_O[8] ;
 wire \Tile_X0Y11_FrameStrobe_O[9] ;
 wire Tile_X0Y11_UserCLKo;
 wire \Tile_X0Y12_E1BEG[0] ;
 wire \Tile_X0Y12_E1BEG[1] ;
 wire \Tile_X0Y12_E1BEG[2] ;
 wire \Tile_X0Y12_E1BEG[3] ;
 wire \Tile_X0Y12_E2BEG[0] ;
 wire \Tile_X0Y12_E2BEG[1] ;
 wire \Tile_X0Y12_E2BEG[2] ;
 wire \Tile_X0Y12_E2BEG[3] ;
 wire \Tile_X0Y12_E2BEG[4] ;
 wire \Tile_X0Y12_E2BEG[5] ;
 wire \Tile_X0Y12_E2BEG[6] ;
 wire \Tile_X0Y12_E2BEG[7] ;
 wire \Tile_X0Y12_E2BEGb[0] ;
 wire \Tile_X0Y12_E2BEGb[1] ;
 wire \Tile_X0Y12_E2BEGb[2] ;
 wire \Tile_X0Y12_E2BEGb[3] ;
 wire \Tile_X0Y12_E2BEGb[4] ;
 wire \Tile_X0Y12_E2BEGb[5] ;
 wire \Tile_X0Y12_E2BEGb[6] ;
 wire \Tile_X0Y12_E2BEGb[7] ;
 wire \Tile_X0Y12_E6BEG[0] ;
 wire \Tile_X0Y12_E6BEG[10] ;
 wire \Tile_X0Y12_E6BEG[11] ;
 wire \Tile_X0Y12_E6BEG[1] ;
 wire \Tile_X0Y12_E6BEG[2] ;
 wire \Tile_X0Y12_E6BEG[3] ;
 wire \Tile_X0Y12_E6BEG[4] ;
 wire \Tile_X0Y12_E6BEG[5] ;
 wire \Tile_X0Y12_E6BEG[6] ;
 wire \Tile_X0Y12_E6BEG[7] ;
 wire \Tile_X0Y12_E6BEG[8] ;
 wire \Tile_X0Y12_E6BEG[9] ;
 wire \Tile_X0Y12_EE4BEG[0] ;
 wire \Tile_X0Y12_EE4BEG[10] ;
 wire \Tile_X0Y12_EE4BEG[11] ;
 wire \Tile_X0Y12_EE4BEG[12] ;
 wire \Tile_X0Y12_EE4BEG[13] ;
 wire \Tile_X0Y12_EE4BEG[14] ;
 wire \Tile_X0Y12_EE4BEG[15] ;
 wire \Tile_X0Y12_EE4BEG[1] ;
 wire \Tile_X0Y12_EE4BEG[2] ;
 wire \Tile_X0Y12_EE4BEG[3] ;
 wire \Tile_X0Y12_EE4BEG[4] ;
 wire \Tile_X0Y12_EE4BEG[5] ;
 wire \Tile_X0Y12_EE4BEG[6] ;
 wire \Tile_X0Y12_EE4BEG[7] ;
 wire \Tile_X0Y12_EE4BEG[8] ;
 wire \Tile_X0Y12_EE4BEG[9] ;
 wire \Tile_X0Y12_FrameData_O[0] ;
 wire \Tile_X0Y12_FrameData_O[10] ;
 wire \Tile_X0Y12_FrameData_O[11] ;
 wire \Tile_X0Y12_FrameData_O[12] ;
 wire \Tile_X0Y12_FrameData_O[13] ;
 wire \Tile_X0Y12_FrameData_O[14] ;
 wire \Tile_X0Y12_FrameData_O[15] ;
 wire \Tile_X0Y12_FrameData_O[16] ;
 wire \Tile_X0Y12_FrameData_O[17] ;
 wire \Tile_X0Y12_FrameData_O[18] ;
 wire \Tile_X0Y12_FrameData_O[19] ;
 wire \Tile_X0Y12_FrameData_O[1] ;
 wire \Tile_X0Y12_FrameData_O[20] ;
 wire \Tile_X0Y12_FrameData_O[21] ;
 wire \Tile_X0Y12_FrameData_O[22] ;
 wire \Tile_X0Y12_FrameData_O[23] ;
 wire \Tile_X0Y12_FrameData_O[24] ;
 wire \Tile_X0Y12_FrameData_O[25] ;
 wire \Tile_X0Y12_FrameData_O[26] ;
 wire \Tile_X0Y12_FrameData_O[27] ;
 wire \Tile_X0Y12_FrameData_O[28] ;
 wire \Tile_X0Y12_FrameData_O[29] ;
 wire \Tile_X0Y12_FrameData_O[2] ;
 wire \Tile_X0Y12_FrameData_O[30] ;
 wire \Tile_X0Y12_FrameData_O[31] ;
 wire \Tile_X0Y12_FrameData_O[3] ;
 wire \Tile_X0Y12_FrameData_O[4] ;
 wire \Tile_X0Y12_FrameData_O[5] ;
 wire \Tile_X0Y12_FrameData_O[6] ;
 wire \Tile_X0Y12_FrameData_O[7] ;
 wire \Tile_X0Y12_FrameData_O[8] ;
 wire \Tile_X0Y12_FrameData_O[9] ;
 wire \Tile_X0Y12_FrameStrobe_O[0] ;
 wire \Tile_X0Y12_FrameStrobe_O[10] ;
 wire \Tile_X0Y12_FrameStrobe_O[11] ;
 wire \Tile_X0Y12_FrameStrobe_O[12] ;
 wire \Tile_X0Y12_FrameStrobe_O[13] ;
 wire \Tile_X0Y12_FrameStrobe_O[14] ;
 wire \Tile_X0Y12_FrameStrobe_O[15] ;
 wire \Tile_X0Y12_FrameStrobe_O[16] ;
 wire \Tile_X0Y12_FrameStrobe_O[17] ;
 wire \Tile_X0Y12_FrameStrobe_O[18] ;
 wire \Tile_X0Y12_FrameStrobe_O[19] ;
 wire \Tile_X0Y12_FrameStrobe_O[1] ;
 wire \Tile_X0Y12_FrameStrobe_O[2] ;
 wire \Tile_X0Y12_FrameStrobe_O[3] ;
 wire \Tile_X0Y12_FrameStrobe_O[4] ;
 wire \Tile_X0Y12_FrameStrobe_O[5] ;
 wire \Tile_X0Y12_FrameStrobe_O[6] ;
 wire \Tile_X0Y12_FrameStrobe_O[7] ;
 wire \Tile_X0Y12_FrameStrobe_O[8] ;
 wire \Tile_X0Y12_FrameStrobe_O[9] ;
 wire Tile_X0Y12_UserCLKo;
 wire \Tile_X0Y13_E1BEG[0] ;
 wire \Tile_X0Y13_E1BEG[1] ;
 wire \Tile_X0Y13_E1BEG[2] ;
 wire \Tile_X0Y13_E1BEG[3] ;
 wire \Tile_X0Y13_E2BEG[0] ;
 wire \Tile_X0Y13_E2BEG[1] ;
 wire \Tile_X0Y13_E2BEG[2] ;
 wire \Tile_X0Y13_E2BEG[3] ;
 wire \Tile_X0Y13_E2BEG[4] ;
 wire \Tile_X0Y13_E2BEG[5] ;
 wire \Tile_X0Y13_E2BEG[6] ;
 wire \Tile_X0Y13_E2BEG[7] ;
 wire \Tile_X0Y13_E2BEGb[0] ;
 wire \Tile_X0Y13_E2BEGb[1] ;
 wire \Tile_X0Y13_E2BEGb[2] ;
 wire \Tile_X0Y13_E2BEGb[3] ;
 wire \Tile_X0Y13_E2BEGb[4] ;
 wire \Tile_X0Y13_E2BEGb[5] ;
 wire \Tile_X0Y13_E2BEGb[6] ;
 wire \Tile_X0Y13_E2BEGb[7] ;
 wire \Tile_X0Y13_E6BEG[0] ;
 wire \Tile_X0Y13_E6BEG[10] ;
 wire \Tile_X0Y13_E6BEG[11] ;
 wire \Tile_X0Y13_E6BEG[1] ;
 wire \Tile_X0Y13_E6BEG[2] ;
 wire \Tile_X0Y13_E6BEG[3] ;
 wire \Tile_X0Y13_E6BEG[4] ;
 wire \Tile_X0Y13_E6BEG[5] ;
 wire \Tile_X0Y13_E6BEG[6] ;
 wire \Tile_X0Y13_E6BEG[7] ;
 wire \Tile_X0Y13_E6BEG[8] ;
 wire \Tile_X0Y13_E6BEG[9] ;
 wire \Tile_X0Y13_EE4BEG[0] ;
 wire \Tile_X0Y13_EE4BEG[10] ;
 wire \Tile_X0Y13_EE4BEG[11] ;
 wire \Tile_X0Y13_EE4BEG[12] ;
 wire \Tile_X0Y13_EE4BEG[13] ;
 wire \Tile_X0Y13_EE4BEG[14] ;
 wire \Tile_X0Y13_EE4BEG[15] ;
 wire \Tile_X0Y13_EE4BEG[1] ;
 wire \Tile_X0Y13_EE4BEG[2] ;
 wire \Tile_X0Y13_EE4BEG[3] ;
 wire \Tile_X0Y13_EE4BEG[4] ;
 wire \Tile_X0Y13_EE4BEG[5] ;
 wire \Tile_X0Y13_EE4BEG[6] ;
 wire \Tile_X0Y13_EE4BEG[7] ;
 wire \Tile_X0Y13_EE4BEG[8] ;
 wire \Tile_X0Y13_EE4BEG[9] ;
 wire \Tile_X0Y13_FrameData_O[0] ;
 wire \Tile_X0Y13_FrameData_O[10] ;
 wire \Tile_X0Y13_FrameData_O[11] ;
 wire \Tile_X0Y13_FrameData_O[12] ;
 wire \Tile_X0Y13_FrameData_O[13] ;
 wire \Tile_X0Y13_FrameData_O[14] ;
 wire \Tile_X0Y13_FrameData_O[15] ;
 wire \Tile_X0Y13_FrameData_O[16] ;
 wire \Tile_X0Y13_FrameData_O[17] ;
 wire \Tile_X0Y13_FrameData_O[18] ;
 wire \Tile_X0Y13_FrameData_O[19] ;
 wire \Tile_X0Y13_FrameData_O[1] ;
 wire \Tile_X0Y13_FrameData_O[20] ;
 wire \Tile_X0Y13_FrameData_O[21] ;
 wire \Tile_X0Y13_FrameData_O[22] ;
 wire \Tile_X0Y13_FrameData_O[23] ;
 wire \Tile_X0Y13_FrameData_O[24] ;
 wire \Tile_X0Y13_FrameData_O[25] ;
 wire \Tile_X0Y13_FrameData_O[26] ;
 wire \Tile_X0Y13_FrameData_O[27] ;
 wire \Tile_X0Y13_FrameData_O[28] ;
 wire \Tile_X0Y13_FrameData_O[29] ;
 wire \Tile_X0Y13_FrameData_O[2] ;
 wire \Tile_X0Y13_FrameData_O[30] ;
 wire \Tile_X0Y13_FrameData_O[31] ;
 wire \Tile_X0Y13_FrameData_O[3] ;
 wire \Tile_X0Y13_FrameData_O[4] ;
 wire \Tile_X0Y13_FrameData_O[5] ;
 wire \Tile_X0Y13_FrameData_O[6] ;
 wire \Tile_X0Y13_FrameData_O[7] ;
 wire \Tile_X0Y13_FrameData_O[8] ;
 wire \Tile_X0Y13_FrameData_O[9] ;
 wire \Tile_X0Y13_FrameStrobe_O[0] ;
 wire \Tile_X0Y13_FrameStrobe_O[10] ;
 wire \Tile_X0Y13_FrameStrobe_O[11] ;
 wire \Tile_X0Y13_FrameStrobe_O[12] ;
 wire \Tile_X0Y13_FrameStrobe_O[13] ;
 wire \Tile_X0Y13_FrameStrobe_O[14] ;
 wire \Tile_X0Y13_FrameStrobe_O[15] ;
 wire \Tile_X0Y13_FrameStrobe_O[16] ;
 wire \Tile_X0Y13_FrameStrobe_O[17] ;
 wire \Tile_X0Y13_FrameStrobe_O[18] ;
 wire \Tile_X0Y13_FrameStrobe_O[19] ;
 wire \Tile_X0Y13_FrameStrobe_O[1] ;
 wire \Tile_X0Y13_FrameStrobe_O[2] ;
 wire \Tile_X0Y13_FrameStrobe_O[3] ;
 wire \Tile_X0Y13_FrameStrobe_O[4] ;
 wire \Tile_X0Y13_FrameStrobe_O[5] ;
 wire \Tile_X0Y13_FrameStrobe_O[6] ;
 wire \Tile_X0Y13_FrameStrobe_O[7] ;
 wire \Tile_X0Y13_FrameStrobe_O[8] ;
 wire \Tile_X0Y13_FrameStrobe_O[9] ;
 wire Tile_X0Y13_UserCLKo;
 wire \Tile_X0Y14_E1BEG[0] ;
 wire \Tile_X0Y14_E1BEG[1] ;
 wire \Tile_X0Y14_E1BEG[2] ;
 wire \Tile_X0Y14_E1BEG[3] ;
 wire \Tile_X0Y14_E2BEG[0] ;
 wire \Tile_X0Y14_E2BEG[1] ;
 wire \Tile_X0Y14_E2BEG[2] ;
 wire \Tile_X0Y14_E2BEG[3] ;
 wire \Tile_X0Y14_E2BEG[4] ;
 wire \Tile_X0Y14_E2BEG[5] ;
 wire \Tile_X0Y14_E2BEG[6] ;
 wire \Tile_X0Y14_E2BEG[7] ;
 wire \Tile_X0Y14_E2BEGb[0] ;
 wire \Tile_X0Y14_E2BEGb[1] ;
 wire \Tile_X0Y14_E2BEGb[2] ;
 wire \Tile_X0Y14_E2BEGb[3] ;
 wire \Tile_X0Y14_E2BEGb[4] ;
 wire \Tile_X0Y14_E2BEGb[5] ;
 wire \Tile_X0Y14_E2BEGb[6] ;
 wire \Tile_X0Y14_E2BEGb[7] ;
 wire \Tile_X0Y14_E6BEG[0] ;
 wire \Tile_X0Y14_E6BEG[10] ;
 wire \Tile_X0Y14_E6BEG[11] ;
 wire \Tile_X0Y14_E6BEG[1] ;
 wire \Tile_X0Y14_E6BEG[2] ;
 wire \Tile_X0Y14_E6BEG[3] ;
 wire \Tile_X0Y14_E6BEG[4] ;
 wire \Tile_X0Y14_E6BEG[5] ;
 wire \Tile_X0Y14_E6BEG[6] ;
 wire \Tile_X0Y14_E6BEG[7] ;
 wire \Tile_X0Y14_E6BEG[8] ;
 wire \Tile_X0Y14_E6BEG[9] ;
 wire \Tile_X0Y14_EE4BEG[0] ;
 wire \Tile_X0Y14_EE4BEG[10] ;
 wire \Tile_X0Y14_EE4BEG[11] ;
 wire \Tile_X0Y14_EE4BEG[12] ;
 wire \Tile_X0Y14_EE4BEG[13] ;
 wire \Tile_X0Y14_EE4BEG[14] ;
 wire \Tile_X0Y14_EE4BEG[15] ;
 wire \Tile_X0Y14_EE4BEG[1] ;
 wire \Tile_X0Y14_EE4BEG[2] ;
 wire \Tile_X0Y14_EE4BEG[3] ;
 wire \Tile_X0Y14_EE4BEG[4] ;
 wire \Tile_X0Y14_EE4BEG[5] ;
 wire \Tile_X0Y14_EE4BEG[6] ;
 wire \Tile_X0Y14_EE4BEG[7] ;
 wire \Tile_X0Y14_EE4BEG[8] ;
 wire \Tile_X0Y14_EE4BEG[9] ;
 wire \Tile_X0Y14_FrameData_O[0] ;
 wire \Tile_X0Y14_FrameData_O[10] ;
 wire \Tile_X0Y14_FrameData_O[11] ;
 wire \Tile_X0Y14_FrameData_O[12] ;
 wire \Tile_X0Y14_FrameData_O[13] ;
 wire \Tile_X0Y14_FrameData_O[14] ;
 wire \Tile_X0Y14_FrameData_O[15] ;
 wire \Tile_X0Y14_FrameData_O[16] ;
 wire \Tile_X0Y14_FrameData_O[17] ;
 wire \Tile_X0Y14_FrameData_O[18] ;
 wire \Tile_X0Y14_FrameData_O[19] ;
 wire \Tile_X0Y14_FrameData_O[1] ;
 wire \Tile_X0Y14_FrameData_O[20] ;
 wire \Tile_X0Y14_FrameData_O[21] ;
 wire \Tile_X0Y14_FrameData_O[22] ;
 wire \Tile_X0Y14_FrameData_O[23] ;
 wire \Tile_X0Y14_FrameData_O[24] ;
 wire \Tile_X0Y14_FrameData_O[25] ;
 wire \Tile_X0Y14_FrameData_O[26] ;
 wire \Tile_X0Y14_FrameData_O[27] ;
 wire \Tile_X0Y14_FrameData_O[28] ;
 wire \Tile_X0Y14_FrameData_O[29] ;
 wire \Tile_X0Y14_FrameData_O[2] ;
 wire \Tile_X0Y14_FrameData_O[30] ;
 wire \Tile_X0Y14_FrameData_O[31] ;
 wire \Tile_X0Y14_FrameData_O[3] ;
 wire \Tile_X0Y14_FrameData_O[4] ;
 wire \Tile_X0Y14_FrameData_O[5] ;
 wire \Tile_X0Y14_FrameData_O[6] ;
 wire \Tile_X0Y14_FrameData_O[7] ;
 wire \Tile_X0Y14_FrameData_O[8] ;
 wire \Tile_X0Y14_FrameData_O[9] ;
 wire \Tile_X0Y14_FrameStrobe_O[0] ;
 wire \Tile_X0Y14_FrameStrobe_O[10] ;
 wire \Tile_X0Y14_FrameStrobe_O[11] ;
 wire \Tile_X0Y14_FrameStrobe_O[12] ;
 wire \Tile_X0Y14_FrameStrobe_O[13] ;
 wire \Tile_X0Y14_FrameStrobe_O[14] ;
 wire \Tile_X0Y14_FrameStrobe_O[15] ;
 wire \Tile_X0Y14_FrameStrobe_O[16] ;
 wire \Tile_X0Y14_FrameStrobe_O[17] ;
 wire \Tile_X0Y14_FrameStrobe_O[18] ;
 wire \Tile_X0Y14_FrameStrobe_O[19] ;
 wire \Tile_X0Y14_FrameStrobe_O[1] ;
 wire \Tile_X0Y14_FrameStrobe_O[2] ;
 wire \Tile_X0Y14_FrameStrobe_O[3] ;
 wire \Tile_X0Y14_FrameStrobe_O[4] ;
 wire \Tile_X0Y14_FrameStrobe_O[5] ;
 wire \Tile_X0Y14_FrameStrobe_O[6] ;
 wire \Tile_X0Y14_FrameStrobe_O[7] ;
 wire \Tile_X0Y14_FrameStrobe_O[8] ;
 wire \Tile_X0Y14_FrameStrobe_O[9] ;
 wire Tile_X0Y14_UserCLKo;
 wire \Tile_X0Y1_E1BEG[0] ;
 wire \Tile_X0Y1_E1BEG[1] ;
 wire \Tile_X0Y1_E1BEG[2] ;
 wire \Tile_X0Y1_E1BEG[3] ;
 wire \Tile_X0Y1_E2BEG[0] ;
 wire \Tile_X0Y1_E2BEG[1] ;
 wire \Tile_X0Y1_E2BEG[2] ;
 wire \Tile_X0Y1_E2BEG[3] ;
 wire \Tile_X0Y1_E2BEG[4] ;
 wire \Tile_X0Y1_E2BEG[5] ;
 wire \Tile_X0Y1_E2BEG[6] ;
 wire \Tile_X0Y1_E2BEG[7] ;
 wire \Tile_X0Y1_E2BEGb[0] ;
 wire \Tile_X0Y1_E2BEGb[1] ;
 wire \Tile_X0Y1_E2BEGb[2] ;
 wire \Tile_X0Y1_E2BEGb[3] ;
 wire \Tile_X0Y1_E2BEGb[4] ;
 wire \Tile_X0Y1_E2BEGb[5] ;
 wire \Tile_X0Y1_E2BEGb[6] ;
 wire \Tile_X0Y1_E2BEGb[7] ;
 wire \Tile_X0Y1_E6BEG[0] ;
 wire \Tile_X0Y1_E6BEG[10] ;
 wire \Tile_X0Y1_E6BEG[11] ;
 wire \Tile_X0Y1_E6BEG[1] ;
 wire \Tile_X0Y1_E6BEG[2] ;
 wire \Tile_X0Y1_E6BEG[3] ;
 wire \Tile_X0Y1_E6BEG[4] ;
 wire \Tile_X0Y1_E6BEG[5] ;
 wire \Tile_X0Y1_E6BEG[6] ;
 wire \Tile_X0Y1_E6BEG[7] ;
 wire \Tile_X0Y1_E6BEG[8] ;
 wire \Tile_X0Y1_E6BEG[9] ;
 wire \Tile_X0Y1_EE4BEG[0] ;
 wire \Tile_X0Y1_EE4BEG[10] ;
 wire \Tile_X0Y1_EE4BEG[11] ;
 wire \Tile_X0Y1_EE4BEG[12] ;
 wire \Tile_X0Y1_EE4BEG[13] ;
 wire \Tile_X0Y1_EE4BEG[14] ;
 wire \Tile_X0Y1_EE4BEG[15] ;
 wire \Tile_X0Y1_EE4BEG[1] ;
 wire \Tile_X0Y1_EE4BEG[2] ;
 wire \Tile_X0Y1_EE4BEG[3] ;
 wire \Tile_X0Y1_EE4BEG[4] ;
 wire \Tile_X0Y1_EE4BEG[5] ;
 wire \Tile_X0Y1_EE4BEG[6] ;
 wire \Tile_X0Y1_EE4BEG[7] ;
 wire \Tile_X0Y1_EE4BEG[8] ;
 wire \Tile_X0Y1_EE4BEG[9] ;
 wire \Tile_X0Y1_FrameData_O[0] ;
 wire \Tile_X0Y1_FrameData_O[10] ;
 wire \Tile_X0Y1_FrameData_O[11] ;
 wire \Tile_X0Y1_FrameData_O[12] ;
 wire \Tile_X0Y1_FrameData_O[13] ;
 wire \Tile_X0Y1_FrameData_O[14] ;
 wire \Tile_X0Y1_FrameData_O[15] ;
 wire \Tile_X0Y1_FrameData_O[16] ;
 wire \Tile_X0Y1_FrameData_O[17] ;
 wire \Tile_X0Y1_FrameData_O[18] ;
 wire \Tile_X0Y1_FrameData_O[19] ;
 wire \Tile_X0Y1_FrameData_O[1] ;
 wire \Tile_X0Y1_FrameData_O[20] ;
 wire \Tile_X0Y1_FrameData_O[21] ;
 wire \Tile_X0Y1_FrameData_O[22] ;
 wire \Tile_X0Y1_FrameData_O[23] ;
 wire \Tile_X0Y1_FrameData_O[24] ;
 wire \Tile_X0Y1_FrameData_O[25] ;
 wire \Tile_X0Y1_FrameData_O[26] ;
 wire \Tile_X0Y1_FrameData_O[27] ;
 wire \Tile_X0Y1_FrameData_O[28] ;
 wire \Tile_X0Y1_FrameData_O[29] ;
 wire \Tile_X0Y1_FrameData_O[2] ;
 wire \Tile_X0Y1_FrameData_O[30] ;
 wire \Tile_X0Y1_FrameData_O[31] ;
 wire \Tile_X0Y1_FrameData_O[3] ;
 wire \Tile_X0Y1_FrameData_O[4] ;
 wire \Tile_X0Y1_FrameData_O[5] ;
 wire \Tile_X0Y1_FrameData_O[6] ;
 wire \Tile_X0Y1_FrameData_O[7] ;
 wire \Tile_X0Y1_FrameData_O[8] ;
 wire \Tile_X0Y1_FrameData_O[9] ;
 wire \Tile_X0Y1_FrameStrobe_O[0] ;
 wire \Tile_X0Y1_FrameStrobe_O[10] ;
 wire \Tile_X0Y1_FrameStrobe_O[11] ;
 wire \Tile_X0Y1_FrameStrobe_O[12] ;
 wire \Tile_X0Y1_FrameStrobe_O[13] ;
 wire \Tile_X0Y1_FrameStrobe_O[14] ;
 wire \Tile_X0Y1_FrameStrobe_O[15] ;
 wire \Tile_X0Y1_FrameStrobe_O[16] ;
 wire \Tile_X0Y1_FrameStrobe_O[17] ;
 wire \Tile_X0Y1_FrameStrobe_O[18] ;
 wire \Tile_X0Y1_FrameStrobe_O[19] ;
 wire \Tile_X0Y1_FrameStrobe_O[1] ;
 wire \Tile_X0Y1_FrameStrobe_O[2] ;
 wire \Tile_X0Y1_FrameStrobe_O[3] ;
 wire \Tile_X0Y1_FrameStrobe_O[4] ;
 wire \Tile_X0Y1_FrameStrobe_O[5] ;
 wire \Tile_X0Y1_FrameStrobe_O[6] ;
 wire \Tile_X0Y1_FrameStrobe_O[7] ;
 wire \Tile_X0Y1_FrameStrobe_O[8] ;
 wire \Tile_X0Y1_FrameStrobe_O[9] ;
 wire Tile_X0Y1_UserCLKo;
 wire \Tile_X0Y2_E1BEG[0] ;
 wire \Tile_X0Y2_E1BEG[1] ;
 wire \Tile_X0Y2_E1BEG[2] ;
 wire \Tile_X0Y2_E1BEG[3] ;
 wire \Tile_X0Y2_E2BEG[0] ;
 wire \Tile_X0Y2_E2BEG[1] ;
 wire \Tile_X0Y2_E2BEG[2] ;
 wire \Tile_X0Y2_E2BEG[3] ;
 wire \Tile_X0Y2_E2BEG[4] ;
 wire \Tile_X0Y2_E2BEG[5] ;
 wire \Tile_X0Y2_E2BEG[6] ;
 wire \Tile_X0Y2_E2BEG[7] ;
 wire \Tile_X0Y2_E2BEGb[0] ;
 wire \Tile_X0Y2_E2BEGb[1] ;
 wire \Tile_X0Y2_E2BEGb[2] ;
 wire \Tile_X0Y2_E2BEGb[3] ;
 wire \Tile_X0Y2_E2BEGb[4] ;
 wire \Tile_X0Y2_E2BEGb[5] ;
 wire \Tile_X0Y2_E2BEGb[6] ;
 wire \Tile_X0Y2_E2BEGb[7] ;
 wire \Tile_X0Y2_E6BEG[0] ;
 wire \Tile_X0Y2_E6BEG[10] ;
 wire \Tile_X0Y2_E6BEG[11] ;
 wire \Tile_X0Y2_E6BEG[1] ;
 wire \Tile_X0Y2_E6BEG[2] ;
 wire \Tile_X0Y2_E6BEG[3] ;
 wire \Tile_X0Y2_E6BEG[4] ;
 wire \Tile_X0Y2_E6BEG[5] ;
 wire \Tile_X0Y2_E6BEG[6] ;
 wire \Tile_X0Y2_E6BEG[7] ;
 wire \Tile_X0Y2_E6BEG[8] ;
 wire \Tile_X0Y2_E6BEG[9] ;
 wire \Tile_X0Y2_EE4BEG[0] ;
 wire \Tile_X0Y2_EE4BEG[10] ;
 wire \Tile_X0Y2_EE4BEG[11] ;
 wire \Tile_X0Y2_EE4BEG[12] ;
 wire \Tile_X0Y2_EE4BEG[13] ;
 wire \Tile_X0Y2_EE4BEG[14] ;
 wire \Tile_X0Y2_EE4BEG[15] ;
 wire \Tile_X0Y2_EE4BEG[1] ;
 wire \Tile_X0Y2_EE4BEG[2] ;
 wire \Tile_X0Y2_EE4BEG[3] ;
 wire \Tile_X0Y2_EE4BEG[4] ;
 wire \Tile_X0Y2_EE4BEG[5] ;
 wire \Tile_X0Y2_EE4BEG[6] ;
 wire \Tile_X0Y2_EE4BEG[7] ;
 wire \Tile_X0Y2_EE4BEG[8] ;
 wire \Tile_X0Y2_EE4BEG[9] ;
 wire \Tile_X0Y2_FrameData_O[0] ;
 wire \Tile_X0Y2_FrameData_O[10] ;
 wire \Tile_X0Y2_FrameData_O[11] ;
 wire \Tile_X0Y2_FrameData_O[12] ;
 wire \Tile_X0Y2_FrameData_O[13] ;
 wire \Tile_X0Y2_FrameData_O[14] ;
 wire \Tile_X0Y2_FrameData_O[15] ;
 wire \Tile_X0Y2_FrameData_O[16] ;
 wire \Tile_X0Y2_FrameData_O[17] ;
 wire \Tile_X0Y2_FrameData_O[18] ;
 wire \Tile_X0Y2_FrameData_O[19] ;
 wire \Tile_X0Y2_FrameData_O[1] ;
 wire \Tile_X0Y2_FrameData_O[20] ;
 wire \Tile_X0Y2_FrameData_O[21] ;
 wire \Tile_X0Y2_FrameData_O[22] ;
 wire \Tile_X0Y2_FrameData_O[23] ;
 wire \Tile_X0Y2_FrameData_O[24] ;
 wire \Tile_X0Y2_FrameData_O[25] ;
 wire \Tile_X0Y2_FrameData_O[26] ;
 wire \Tile_X0Y2_FrameData_O[27] ;
 wire \Tile_X0Y2_FrameData_O[28] ;
 wire \Tile_X0Y2_FrameData_O[29] ;
 wire \Tile_X0Y2_FrameData_O[2] ;
 wire \Tile_X0Y2_FrameData_O[30] ;
 wire \Tile_X0Y2_FrameData_O[31] ;
 wire \Tile_X0Y2_FrameData_O[3] ;
 wire \Tile_X0Y2_FrameData_O[4] ;
 wire \Tile_X0Y2_FrameData_O[5] ;
 wire \Tile_X0Y2_FrameData_O[6] ;
 wire \Tile_X0Y2_FrameData_O[7] ;
 wire \Tile_X0Y2_FrameData_O[8] ;
 wire \Tile_X0Y2_FrameData_O[9] ;
 wire \Tile_X0Y2_FrameStrobe_O[0] ;
 wire \Tile_X0Y2_FrameStrobe_O[10] ;
 wire \Tile_X0Y2_FrameStrobe_O[11] ;
 wire \Tile_X0Y2_FrameStrobe_O[12] ;
 wire \Tile_X0Y2_FrameStrobe_O[13] ;
 wire \Tile_X0Y2_FrameStrobe_O[14] ;
 wire \Tile_X0Y2_FrameStrobe_O[15] ;
 wire \Tile_X0Y2_FrameStrobe_O[16] ;
 wire \Tile_X0Y2_FrameStrobe_O[17] ;
 wire \Tile_X0Y2_FrameStrobe_O[18] ;
 wire \Tile_X0Y2_FrameStrobe_O[19] ;
 wire \Tile_X0Y2_FrameStrobe_O[1] ;
 wire \Tile_X0Y2_FrameStrobe_O[2] ;
 wire \Tile_X0Y2_FrameStrobe_O[3] ;
 wire \Tile_X0Y2_FrameStrobe_O[4] ;
 wire \Tile_X0Y2_FrameStrobe_O[5] ;
 wire \Tile_X0Y2_FrameStrobe_O[6] ;
 wire \Tile_X0Y2_FrameStrobe_O[7] ;
 wire \Tile_X0Y2_FrameStrobe_O[8] ;
 wire \Tile_X0Y2_FrameStrobe_O[9] ;
 wire Tile_X0Y2_UserCLKo;
 wire \Tile_X0Y3_E1BEG[0] ;
 wire \Tile_X0Y3_E1BEG[1] ;
 wire \Tile_X0Y3_E1BEG[2] ;
 wire \Tile_X0Y3_E1BEG[3] ;
 wire \Tile_X0Y3_E2BEG[0] ;
 wire \Tile_X0Y3_E2BEG[1] ;
 wire \Tile_X0Y3_E2BEG[2] ;
 wire \Tile_X0Y3_E2BEG[3] ;
 wire \Tile_X0Y3_E2BEG[4] ;
 wire \Tile_X0Y3_E2BEG[5] ;
 wire \Tile_X0Y3_E2BEG[6] ;
 wire \Tile_X0Y3_E2BEG[7] ;
 wire \Tile_X0Y3_E2BEGb[0] ;
 wire \Tile_X0Y3_E2BEGb[1] ;
 wire \Tile_X0Y3_E2BEGb[2] ;
 wire \Tile_X0Y3_E2BEGb[3] ;
 wire \Tile_X0Y3_E2BEGb[4] ;
 wire \Tile_X0Y3_E2BEGb[5] ;
 wire \Tile_X0Y3_E2BEGb[6] ;
 wire \Tile_X0Y3_E2BEGb[7] ;
 wire \Tile_X0Y3_E6BEG[0] ;
 wire \Tile_X0Y3_E6BEG[10] ;
 wire \Tile_X0Y3_E6BEG[11] ;
 wire \Tile_X0Y3_E6BEG[1] ;
 wire \Tile_X0Y3_E6BEG[2] ;
 wire \Tile_X0Y3_E6BEG[3] ;
 wire \Tile_X0Y3_E6BEG[4] ;
 wire \Tile_X0Y3_E6BEG[5] ;
 wire \Tile_X0Y3_E6BEG[6] ;
 wire \Tile_X0Y3_E6BEG[7] ;
 wire \Tile_X0Y3_E6BEG[8] ;
 wire \Tile_X0Y3_E6BEG[9] ;
 wire \Tile_X0Y3_EE4BEG[0] ;
 wire \Tile_X0Y3_EE4BEG[10] ;
 wire \Tile_X0Y3_EE4BEG[11] ;
 wire \Tile_X0Y3_EE4BEG[12] ;
 wire \Tile_X0Y3_EE4BEG[13] ;
 wire \Tile_X0Y3_EE4BEG[14] ;
 wire \Tile_X0Y3_EE4BEG[15] ;
 wire \Tile_X0Y3_EE4BEG[1] ;
 wire \Tile_X0Y3_EE4BEG[2] ;
 wire \Tile_X0Y3_EE4BEG[3] ;
 wire \Tile_X0Y3_EE4BEG[4] ;
 wire \Tile_X0Y3_EE4BEG[5] ;
 wire \Tile_X0Y3_EE4BEG[6] ;
 wire \Tile_X0Y3_EE4BEG[7] ;
 wire \Tile_X0Y3_EE4BEG[8] ;
 wire \Tile_X0Y3_EE4BEG[9] ;
 wire \Tile_X0Y3_FrameData_O[0] ;
 wire \Tile_X0Y3_FrameData_O[10] ;
 wire \Tile_X0Y3_FrameData_O[11] ;
 wire \Tile_X0Y3_FrameData_O[12] ;
 wire \Tile_X0Y3_FrameData_O[13] ;
 wire \Tile_X0Y3_FrameData_O[14] ;
 wire \Tile_X0Y3_FrameData_O[15] ;
 wire \Tile_X0Y3_FrameData_O[16] ;
 wire \Tile_X0Y3_FrameData_O[17] ;
 wire \Tile_X0Y3_FrameData_O[18] ;
 wire \Tile_X0Y3_FrameData_O[19] ;
 wire \Tile_X0Y3_FrameData_O[1] ;
 wire \Tile_X0Y3_FrameData_O[20] ;
 wire \Tile_X0Y3_FrameData_O[21] ;
 wire \Tile_X0Y3_FrameData_O[22] ;
 wire \Tile_X0Y3_FrameData_O[23] ;
 wire \Tile_X0Y3_FrameData_O[24] ;
 wire \Tile_X0Y3_FrameData_O[25] ;
 wire \Tile_X0Y3_FrameData_O[26] ;
 wire \Tile_X0Y3_FrameData_O[27] ;
 wire \Tile_X0Y3_FrameData_O[28] ;
 wire \Tile_X0Y3_FrameData_O[29] ;
 wire \Tile_X0Y3_FrameData_O[2] ;
 wire \Tile_X0Y3_FrameData_O[30] ;
 wire \Tile_X0Y3_FrameData_O[31] ;
 wire \Tile_X0Y3_FrameData_O[3] ;
 wire \Tile_X0Y3_FrameData_O[4] ;
 wire \Tile_X0Y3_FrameData_O[5] ;
 wire \Tile_X0Y3_FrameData_O[6] ;
 wire \Tile_X0Y3_FrameData_O[7] ;
 wire \Tile_X0Y3_FrameData_O[8] ;
 wire \Tile_X0Y3_FrameData_O[9] ;
 wire \Tile_X0Y3_FrameStrobe_O[0] ;
 wire \Tile_X0Y3_FrameStrobe_O[10] ;
 wire \Tile_X0Y3_FrameStrobe_O[11] ;
 wire \Tile_X0Y3_FrameStrobe_O[12] ;
 wire \Tile_X0Y3_FrameStrobe_O[13] ;
 wire \Tile_X0Y3_FrameStrobe_O[14] ;
 wire \Tile_X0Y3_FrameStrobe_O[15] ;
 wire \Tile_X0Y3_FrameStrobe_O[16] ;
 wire \Tile_X0Y3_FrameStrobe_O[17] ;
 wire \Tile_X0Y3_FrameStrobe_O[18] ;
 wire \Tile_X0Y3_FrameStrobe_O[19] ;
 wire \Tile_X0Y3_FrameStrobe_O[1] ;
 wire \Tile_X0Y3_FrameStrobe_O[2] ;
 wire \Tile_X0Y3_FrameStrobe_O[3] ;
 wire \Tile_X0Y3_FrameStrobe_O[4] ;
 wire \Tile_X0Y3_FrameStrobe_O[5] ;
 wire \Tile_X0Y3_FrameStrobe_O[6] ;
 wire \Tile_X0Y3_FrameStrobe_O[7] ;
 wire \Tile_X0Y3_FrameStrobe_O[8] ;
 wire \Tile_X0Y3_FrameStrobe_O[9] ;
 wire Tile_X0Y3_UserCLKo;
 wire \Tile_X0Y4_E1BEG[0] ;
 wire \Tile_X0Y4_E1BEG[1] ;
 wire \Tile_X0Y4_E1BEG[2] ;
 wire \Tile_X0Y4_E1BEG[3] ;
 wire \Tile_X0Y4_E2BEG[0] ;
 wire \Tile_X0Y4_E2BEG[1] ;
 wire \Tile_X0Y4_E2BEG[2] ;
 wire \Tile_X0Y4_E2BEG[3] ;
 wire \Tile_X0Y4_E2BEG[4] ;
 wire \Tile_X0Y4_E2BEG[5] ;
 wire \Tile_X0Y4_E2BEG[6] ;
 wire \Tile_X0Y4_E2BEG[7] ;
 wire \Tile_X0Y4_E2BEGb[0] ;
 wire \Tile_X0Y4_E2BEGb[1] ;
 wire \Tile_X0Y4_E2BEGb[2] ;
 wire \Tile_X0Y4_E2BEGb[3] ;
 wire \Tile_X0Y4_E2BEGb[4] ;
 wire \Tile_X0Y4_E2BEGb[5] ;
 wire \Tile_X0Y4_E2BEGb[6] ;
 wire \Tile_X0Y4_E2BEGb[7] ;
 wire \Tile_X0Y4_E6BEG[0] ;
 wire \Tile_X0Y4_E6BEG[10] ;
 wire \Tile_X0Y4_E6BEG[11] ;
 wire \Tile_X0Y4_E6BEG[1] ;
 wire \Tile_X0Y4_E6BEG[2] ;
 wire \Tile_X0Y4_E6BEG[3] ;
 wire \Tile_X0Y4_E6BEG[4] ;
 wire \Tile_X0Y4_E6BEG[5] ;
 wire \Tile_X0Y4_E6BEG[6] ;
 wire \Tile_X0Y4_E6BEG[7] ;
 wire \Tile_X0Y4_E6BEG[8] ;
 wire \Tile_X0Y4_E6BEG[9] ;
 wire \Tile_X0Y4_EE4BEG[0] ;
 wire \Tile_X0Y4_EE4BEG[10] ;
 wire \Tile_X0Y4_EE4BEG[11] ;
 wire \Tile_X0Y4_EE4BEG[12] ;
 wire \Tile_X0Y4_EE4BEG[13] ;
 wire \Tile_X0Y4_EE4BEG[14] ;
 wire \Tile_X0Y4_EE4BEG[15] ;
 wire \Tile_X0Y4_EE4BEG[1] ;
 wire \Tile_X0Y4_EE4BEG[2] ;
 wire \Tile_X0Y4_EE4BEG[3] ;
 wire \Tile_X0Y4_EE4BEG[4] ;
 wire \Tile_X0Y4_EE4BEG[5] ;
 wire \Tile_X0Y4_EE4BEG[6] ;
 wire \Tile_X0Y4_EE4BEG[7] ;
 wire \Tile_X0Y4_EE4BEG[8] ;
 wire \Tile_X0Y4_EE4BEG[9] ;
 wire \Tile_X0Y4_FrameData_O[0] ;
 wire \Tile_X0Y4_FrameData_O[10] ;
 wire \Tile_X0Y4_FrameData_O[11] ;
 wire \Tile_X0Y4_FrameData_O[12] ;
 wire \Tile_X0Y4_FrameData_O[13] ;
 wire \Tile_X0Y4_FrameData_O[14] ;
 wire \Tile_X0Y4_FrameData_O[15] ;
 wire \Tile_X0Y4_FrameData_O[16] ;
 wire \Tile_X0Y4_FrameData_O[17] ;
 wire \Tile_X0Y4_FrameData_O[18] ;
 wire \Tile_X0Y4_FrameData_O[19] ;
 wire \Tile_X0Y4_FrameData_O[1] ;
 wire \Tile_X0Y4_FrameData_O[20] ;
 wire \Tile_X0Y4_FrameData_O[21] ;
 wire \Tile_X0Y4_FrameData_O[22] ;
 wire \Tile_X0Y4_FrameData_O[23] ;
 wire \Tile_X0Y4_FrameData_O[24] ;
 wire \Tile_X0Y4_FrameData_O[25] ;
 wire \Tile_X0Y4_FrameData_O[26] ;
 wire \Tile_X0Y4_FrameData_O[27] ;
 wire \Tile_X0Y4_FrameData_O[28] ;
 wire \Tile_X0Y4_FrameData_O[29] ;
 wire \Tile_X0Y4_FrameData_O[2] ;
 wire \Tile_X0Y4_FrameData_O[30] ;
 wire \Tile_X0Y4_FrameData_O[31] ;
 wire \Tile_X0Y4_FrameData_O[3] ;
 wire \Tile_X0Y4_FrameData_O[4] ;
 wire \Tile_X0Y4_FrameData_O[5] ;
 wire \Tile_X0Y4_FrameData_O[6] ;
 wire \Tile_X0Y4_FrameData_O[7] ;
 wire \Tile_X0Y4_FrameData_O[8] ;
 wire \Tile_X0Y4_FrameData_O[9] ;
 wire \Tile_X0Y4_FrameStrobe_O[0] ;
 wire \Tile_X0Y4_FrameStrobe_O[10] ;
 wire \Tile_X0Y4_FrameStrobe_O[11] ;
 wire \Tile_X0Y4_FrameStrobe_O[12] ;
 wire \Tile_X0Y4_FrameStrobe_O[13] ;
 wire \Tile_X0Y4_FrameStrobe_O[14] ;
 wire \Tile_X0Y4_FrameStrobe_O[15] ;
 wire \Tile_X0Y4_FrameStrobe_O[16] ;
 wire \Tile_X0Y4_FrameStrobe_O[17] ;
 wire \Tile_X0Y4_FrameStrobe_O[18] ;
 wire \Tile_X0Y4_FrameStrobe_O[19] ;
 wire \Tile_X0Y4_FrameStrobe_O[1] ;
 wire \Tile_X0Y4_FrameStrobe_O[2] ;
 wire \Tile_X0Y4_FrameStrobe_O[3] ;
 wire \Tile_X0Y4_FrameStrobe_O[4] ;
 wire \Tile_X0Y4_FrameStrobe_O[5] ;
 wire \Tile_X0Y4_FrameStrobe_O[6] ;
 wire \Tile_X0Y4_FrameStrobe_O[7] ;
 wire \Tile_X0Y4_FrameStrobe_O[8] ;
 wire \Tile_X0Y4_FrameStrobe_O[9] ;
 wire Tile_X0Y4_UserCLKo;
 wire \Tile_X0Y5_E1BEG[0] ;
 wire \Tile_X0Y5_E1BEG[1] ;
 wire \Tile_X0Y5_E1BEG[2] ;
 wire \Tile_X0Y5_E1BEG[3] ;
 wire \Tile_X0Y5_E2BEG[0] ;
 wire \Tile_X0Y5_E2BEG[1] ;
 wire \Tile_X0Y5_E2BEG[2] ;
 wire \Tile_X0Y5_E2BEG[3] ;
 wire \Tile_X0Y5_E2BEG[4] ;
 wire \Tile_X0Y5_E2BEG[5] ;
 wire \Tile_X0Y5_E2BEG[6] ;
 wire \Tile_X0Y5_E2BEG[7] ;
 wire \Tile_X0Y5_E2BEGb[0] ;
 wire \Tile_X0Y5_E2BEGb[1] ;
 wire \Tile_X0Y5_E2BEGb[2] ;
 wire \Tile_X0Y5_E2BEGb[3] ;
 wire \Tile_X0Y5_E2BEGb[4] ;
 wire \Tile_X0Y5_E2BEGb[5] ;
 wire \Tile_X0Y5_E2BEGb[6] ;
 wire \Tile_X0Y5_E2BEGb[7] ;
 wire \Tile_X0Y5_E6BEG[0] ;
 wire \Tile_X0Y5_E6BEG[10] ;
 wire \Tile_X0Y5_E6BEG[11] ;
 wire \Tile_X0Y5_E6BEG[1] ;
 wire \Tile_X0Y5_E6BEG[2] ;
 wire \Tile_X0Y5_E6BEG[3] ;
 wire \Tile_X0Y5_E6BEG[4] ;
 wire \Tile_X0Y5_E6BEG[5] ;
 wire \Tile_X0Y5_E6BEG[6] ;
 wire \Tile_X0Y5_E6BEG[7] ;
 wire \Tile_X0Y5_E6BEG[8] ;
 wire \Tile_X0Y5_E6BEG[9] ;
 wire \Tile_X0Y5_EE4BEG[0] ;
 wire \Tile_X0Y5_EE4BEG[10] ;
 wire \Tile_X0Y5_EE4BEG[11] ;
 wire \Tile_X0Y5_EE4BEG[12] ;
 wire \Tile_X0Y5_EE4BEG[13] ;
 wire \Tile_X0Y5_EE4BEG[14] ;
 wire \Tile_X0Y5_EE4BEG[15] ;
 wire \Tile_X0Y5_EE4BEG[1] ;
 wire \Tile_X0Y5_EE4BEG[2] ;
 wire \Tile_X0Y5_EE4BEG[3] ;
 wire \Tile_X0Y5_EE4BEG[4] ;
 wire \Tile_X0Y5_EE4BEG[5] ;
 wire \Tile_X0Y5_EE4BEG[6] ;
 wire \Tile_X0Y5_EE4BEG[7] ;
 wire \Tile_X0Y5_EE4BEG[8] ;
 wire \Tile_X0Y5_EE4BEG[9] ;
 wire \Tile_X0Y5_FrameData_O[0] ;
 wire \Tile_X0Y5_FrameData_O[10] ;
 wire \Tile_X0Y5_FrameData_O[11] ;
 wire \Tile_X0Y5_FrameData_O[12] ;
 wire \Tile_X0Y5_FrameData_O[13] ;
 wire \Tile_X0Y5_FrameData_O[14] ;
 wire \Tile_X0Y5_FrameData_O[15] ;
 wire \Tile_X0Y5_FrameData_O[16] ;
 wire \Tile_X0Y5_FrameData_O[17] ;
 wire \Tile_X0Y5_FrameData_O[18] ;
 wire \Tile_X0Y5_FrameData_O[19] ;
 wire \Tile_X0Y5_FrameData_O[1] ;
 wire \Tile_X0Y5_FrameData_O[20] ;
 wire \Tile_X0Y5_FrameData_O[21] ;
 wire \Tile_X0Y5_FrameData_O[22] ;
 wire \Tile_X0Y5_FrameData_O[23] ;
 wire \Tile_X0Y5_FrameData_O[24] ;
 wire \Tile_X0Y5_FrameData_O[25] ;
 wire \Tile_X0Y5_FrameData_O[26] ;
 wire \Tile_X0Y5_FrameData_O[27] ;
 wire \Tile_X0Y5_FrameData_O[28] ;
 wire \Tile_X0Y5_FrameData_O[29] ;
 wire \Tile_X0Y5_FrameData_O[2] ;
 wire \Tile_X0Y5_FrameData_O[30] ;
 wire \Tile_X0Y5_FrameData_O[31] ;
 wire \Tile_X0Y5_FrameData_O[3] ;
 wire \Tile_X0Y5_FrameData_O[4] ;
 wire \Tile_X0Y5_FrameData_O[5] ;
 wire \Tile_X0Y5_FrameData_O[6] ;
 wire \Tile_X0Y5_FrameData_O[7] ;
 wire \Tile_X0Y5_FrameData_O[8] ;
 wire \Tile_X0Y5_FrameData_O[9] ;
 wire \Tile_X0Y5_FrameStrobe_O[0] ;
 wire \Tile_X0Y5_FrameStrobe_O[10] ;
 wire \Tile_X0Y5_FrameStrobe_O[11] ;
 wire \Tile_X0Y5_FrameStrobe_O[12] ;
 wire \Tile_X0Y5_FrameStrobe_O[13] ;
 wire \Tile_X0Y5_FrameStrobe_O[14] ;
 wire \Tile_X0Y5_FrameStrobe_O[15] ;
 wire \Tile_X0Y5_FrameStrobe_O[16] ;
 wire \Tile_X0Y5_FrameStrobe_O[17] ;
 wire \Tile_X0Y5_FrameStrobe_O[18] ;
 wire \Tile_X0Y5_FrameStrobe_O[19] ;
 wire \Tile_X0Y5_FrameStrobe_O[1] ;
 wire \Tile_X0Y5_FrameStrobe_O[2] ;
 wire \Tile_X0Y5_FrameStrobe_O[3] ;
 wire \Tile_X0Y5_FrameStrobe_O[4] ;
 wire \Tile_X0Y5_FrameStrobe_O[5] ;
 wire \Tile_X0Y5_FrameStrobe_O[6] ;
 wire \Tile_X0Y5_FrameStrobe_O[7] ;
 wire \Tile_X0Y5_FrameStrobe_O[8] ;
 wire \Tile_X0Y5_FrameStrobe_O[9] ;
 wire Tile_X0Y5_UserCLKo;
 wire \Tile_X0Y6_E1BEG[0] ;
 wire \Tile_X0Y6_E1BEG[1] ;
 wire \Tile_X0Y6_E1BEG[2] ;
 wire \Tile_X0Y6_E1BEG[3] ;
 wire \Tile_X0Y6_E2BEG[0] ;
 wire \Tile_X0Y6_E2BEG[1] ;
 wire \Tile_X0Y6_E2BEG[2] ;
 wire \Tile_X0Y6_E2BEG[3] ;
 wire \Tile_X0Y6_E2BEG[4] ;
 wire \Tile_X0Y6_E2BEG[5] ;
 wire \Tile_X0Y6_E2BEG[6] ;
 wire \Tile_X0Y6_E2BEG[7] ;
 wire \Tile_X0Y6_E2BEGb[0] ;
 wire \Tile_X0Y6_E2BEGb[1] ;
 wire \Tile_X0Y6_E2BEGb[2] ;
 wire \Tile_X0Y6_E2BEGb[3] ;
 wire \Tile_X0Y6_E2BEGb[4] ;
 wire \Tile_X0Y6_E2BEGb[5] ;
 wire \Tile_X0Y6_E2BEGb[6] ;
 wire \Tile_X0Y6_E2BEGb[7] ;
 wire \Tile_X0Y6_E6BEG[0] ;
 wire \Tile_X0Y6_E6BEG[10] ;
 wire \Tile_X0Y6_E6BEG[11] ;
 wire \Tile_X0Y6_E6BEG[1] ;
 wire \Tile_X0Y6_E6BEG[2] ;
 wire \Tile_X0Y6_E6BEG[3] ;
 wire \Tile_X0Y6_E6BEG[4] ;
 wire \Tile_X0Y6_E6BEG[5] ;
 wire \Tile_X0Y6_E6BEG[6] ;
 wire \Tile_X0Y6_E6BEG[7] ;
 wire \Tile_X0Y6_E6BEG[8] ;
 wire \Tile_X0Y6_E6BEG[9] ;
 wire \Tile_X0Y6_EE4BEG[0] ;
 wire \Tile_X0Y6_EE4BEG[10] ;
 wire \Tile_X0Y6_EE4BEG[11] ;
 wire \Tile_X0Y6_EE4BEG[12] ;
 wire \Tile_X0Y6_EE4BEG[13] ;
 wire \Tile_X0Y6_EE4BEG[14] ;
 wire \Tile_X0Y6_EE4BEG[15] ;
 wire \Tile_X0Y6_EE4BEG[1] ;
 wire \Tile_X0Y6_EE4BEG[2] ;
 wire \Tile_X0Y6_EE4BEG[3] ;
 wire \Tile_X0Y6_EE4BEG[4] ;
 wire \Tile_X0Y6_EE4BEG[5] ;
 wire \Tile_X0Y6_EE4BEG[6] ;
 wire \Tile_X0Y6_EE4BEG[7] ;
 wire \Tile_X0Y6_EE4BEG[8] ;
 wire \Tile_X0Y6_EE4BEG[9] ;
 wire \Tile_X0Y6_FrameData_O[0] ;
 wire \Tile_X0Y6_FrameData_O[10] ;
 wire \Tile_X0Y6_FrameData_O[11] ;
 wire \Tile_X0Y6_FrameData_O[12] ;
 wire \Tile_X0Y6_FrameData_O[13] ;
 wire \Tile_X0Y6_FrameData_O[14] ;
 wire \Tile_X0Y6_FrameData_O[15] ;
 wire \Tile_X0Y6_FrameData_O[16] ;
 wire \Tile_X0Y6_FrameData_O[17] ;
 wire \Tile_X0Y6_FrameData_O[18] ;
 wire \Tile_X0Y6_FrameData_O[19] ;
 wire \Tile_X0Y6_FrameData_O[1] ;
 wire \Tile_X0Y6_FrameData_O[20] ;
 wire \Tile_X0Y6_FrameData_O[21] ;
 wire \Tile_X0Y6_FrameData_O[22] ;
 wire \Tile_X0Y6_FrameData_O[23] ;
 wire \Tile_X0Y6_FrameData_O[24] ;
 wire \Tile_X0Y6_FrameData_O[25] ;
 wire \Tile_X0Y6_FrameData_O[26] ;
 wire \Tile_X0Y6_FrameData_O[27] ;
 wire \Tile_X0Y6_FrameData_O[28] ;
 wire \Tile_X0Y6_FrameData_O[29] ;
 wire \Tile_X0Y6_FrameData_O[2] ;
 wire \Tile_X0Y6_FrameData_O[30] ;
 wire \Tile_X0Y6_FrameData_O[31] ;
 wire \Tile_X0Y6_FrameData_O[3] ;
 wire \Tile_X0Y6_FrameData_O[4] ;
 wire \Tile_X0Y6_FrameData_O[5] ;
 wire \Tile_X0Y6_FrameData_O[6] ;
 wire \Tile_X0Y6_FrameData_O[7] ;
 wire \Tile_X0Y6_FrameData_O[8] ;
 wire \Tile_X0Y6_FrameData_O[9] ;
 wire \Tile_X0Y6_FrameStrobe_O[0] ;
 wire \Tile_X0Y6_FrameStrobe_O[10] ;
 wire \Tile_X0Y6_FrameStrobe_O[11] ;
 wire \Tile_X0Y6_FrameStrobe_O[12] ;
 wire \Tile_X0Y6_FrameStrobe_O[13] ;
 wire \Tile_X0Y6_FrameStrobe_O[14] ;
 wire \Tile_X0Y6_FrameStrobe_O[15] ;
 wire \Tile_X0Y6_FrameStrobe_O[16] ;
 wire \Tile_X0Y6_FrameStrobe_O[17] ;
 wire \Tile_X0Y6_FrameStrobe_O[18] ;
 wire \Tile_X0Y6_FrameStrobe_O[19] ;
 wire \Tile_X0Y6_FrameStrobe_O[1] ;
 wire \Tile_X0Y6_FrameStrobe_O[2] ;
 wire \Tile_X0Y6_FrameStrobe_O[3] ;
 wire \Tile_X0Y6_FrameStrobe_O[4] ;
 wire \Tile_X0Y6_FrameStrobe_O[5] ;
 wire \Tile_X0Y6_FrameStrobe_O[6] ;
 wire \Tile_X0Y6_FrameStrobe_O[7] ;
 wire \Tile_X0Y6_FrameStrobe_O[8] ;
 wire \Tile_X0Y6_FrameStrobe_O[9] ;
 wire Tile_X0Y6_UserCLKo;
 wire \Tile_X0Y7_E1BEG[0] ;
 wire \Tile_X0Y7_E1BEG[1] ;
 wire \Tile_X0Y7_E1BEG[2] ;
 wire \Tile_X0Y7_E1BEG[3] ;
 wire \Tile_X0Y7_E2BEG[0] ;
 wire \Tile_X0Y7_E2BEG[1] ;
 wire \Tile_X0Y7_E2BEG[2] ;
 wire \Tile_X0Y7_E2BEG[3] ;
 wire \Tile_X0Y7_E2BEG[4] ;
 wire \Tile_X0Y7_E2BEG[5] ;
 wire \Tile_X0Y7_E2BEG[6] ;
 wire \Tile_X0Y7_E2BEG[7] ;
 wire \Tile_X0Y7_E2BEGb[0] ;
 wire \Tile_X0Y7_E2BEGb[1] ;
 wire \Tile_X0Y7_E2BEGb[2] ;
 wire \Tile_X0Y7_E2BEGb[3] ;
 wire \Tile_X0Y7_E2BEGb[4] ;
 wire \Tile_X0Y7_E2BEGb[5] ;
 wire \Tile_X0Y7_E2BEGb[6] ;
 wire \Tile_X0Y7_E2BEGb[7] ;
 wire \Tile_X0Y7_E6BEG[0] ;
 wire \Tile_X0Y7_E6BEG[10] ;
 wire \Tile_X0Y7_E6BEG[11] ;
 wire \Tile_X0Y7_E6BEG[1] ;
 wire \Tile_X0Y7_E6BEG[2] ;
 wire \Tile_X0Y7_E6BEG[3] ;
 wire \Tile_X0Y7_E6BEG[4] ;
 wire \Tile_X0Y7_E6BEG[5] ;
 wire \Tile_X0Y7_E6BEG[6] ;
 wire \Tile_X0Y7_E6BEG[7] ;
 wire \Tile_X0Y7_E6BEG[8] ;
 wire \Tile_X0Y7_E6BEG[9] ;
 wire \Tile_X0Y7_EE4BEG[0] ;
 wire \Tile_X0Y7_EE4BEG[10] ;
 wire \Tile_X0Y7_EE4BEG[11] ;
 wire \Tile_X0Y7_EE4BEG[12] ;
 wire \Tile_X0Y7_EE4BEG[13] ;
 wire \Tile_X0Y7_EE4BEG[14] ;
 wire \Tile_X0Y7_EE4BEG[15] ;
 wire \Tile_X0Y7_EE4BEG[1] ;
 wire \Tile_X0Y7_EE4BEG[2] ;
 wire \Tile_X0Y7_EE4BEG[3] ;
 wire \Tile_X0Y7_EE4BEG[4] ;
 wire \Tile_X0Y7_EE4BEG[5] ;
 wire \Tile_X0Y7_EE4BEG[6] ;
 wire \Tile_X0Y7_EE4BEG[7] ;
 wire \Tile_X0Y7_EE4BEG[8] ;
 wire \Tile_X0Y7_EE4BEG[9] ;
 wire \Tile_X0Y7_FrameData_O[0] ;
 wire \Tile_X0Y7_FrameData_O[10] ;
 wire \Tile_X0Y7_FrameData_O[11] ;
 wire \Tile_X0Y7_FrameData_O[12] ;
 wire \Tile_X0Y7_FrameData_O[13] ;
 wire \Tile_X0Y7_FrameData_O[14] ;
 wire \Tile_X0Y7_FrameData_O[15] ;
 wire \Tile_X0Y7_FrameData_O[16] ;
 wire \Tile_X0Y7_FrameData_O[17] ;
 wire \Tile_X0Y7_FrameData_O[18] ;
 wire \Tile_X0Y7_FrameData_O[19] ;
 wire \Tile_X0Y7_FrameData_O[1] ;
 wire \Tile_X0Y7_FrameData_O[20] ;
 wire \Tile_X0Y7_FrameData_O[21] ;
 wire \Tile_X0Y7_FrameData_O[22] ;
 wire \Tile_X0Y7_FrameData_O[23] ;
 wire \Tile_X0Y7_FrameData_O[24] ;
 wire \Tile_X0Y7_FrameData_O[25] ;
 wire \Tile_X0Y7_FrameData_O[26] ;
 wire \Tile_X0Y7_FrameData_O[27] ;
 wire \Tile_X0Y7_FrameData_O[28] ;
 wire \Tile_X0Y7_FrameData_O[29] ;
 wire \Tile_X0Y7_FrameData_O[2] ;
 wire \Tile_X0Y7_FrameData_O[30] ;
 wire \Tile_X0Y7_FrameData_O[31] ;
 wire \Tile_X0Y7_FrameData_O[3] ;
 wire \Tile_X0Y7_FrameData_O[4] ;
 wire \Tile_X0Y7_FrameData_O[5] ;
 wire \Tile_X0Y7_FrameData_O[6] ;
 wire \Tile_X0Y7_FrameData_O[7] ;
 wire \Tile_X0Y7_FrameData_O[8] ;
 wire \Tile_X0Y7_FrameData_O[9] ;
 wire \Tile_X0Y7_FrameStrobe_O[0] ;
 wire \Tile_X0Y7_FrameStrobe_O[10] ;
 wire \Tile_X0Y7_FrameStrobe_O[11] ;
 wire \Tile_X0Y7_FrameStrobe_O[12] ;
 wire \Tile_X0Y7_FrameStrobe_O[13] ;
 wire \Tile_X0Y7_FrameStrobe_O[14] ;
 wire \Tile_X0Y7_FrameStrobe_O[15] ;
 wire \Tile_X0Y7_FrameStrobe_O[16] ;
 wire \Tile_X0Y7_FrameStrobe_O[17] ;
 wire \Tile_X0Y7_FrameStrobe_O[18] ;
 wire \Tile_X0Y7_FrameStrobe_O[19] ;
 wire \Tile_X0Y7_FrameStrobe_O[1] ;
 wire \Tile_X0Y7_FrameStrobe_O[2] ;
 wire \Tile_X0Y7_FrameStrobe_O[3] ;
 wire \Tile_X0Y7_FrameStrobe_O[4] ;
 wire \Tile_X0Y7_FrameStrobe_O[5] ;
 wire \Tile_X0Y7_FrameStrobe_O[6] ;
 wire \Tile_X0Y7_FrameStrobe_O[7] ;
 wire \Tile_X0Y7_FrameStrobe_O[8] ;
 wire \Tile_X0Y7_FrameStrobe_O[9] ;
 wire Tile_X0Y7_UserCLKo;
 wire \Tile_X0Y8_E1BEG[0] ;
 wire \Tile_X0Y8_E1BEG[1] ;
 wire \Tile_X0Y8_E1BEG[2] ;
 wire \Tile_X0Y8_E1BEG[3] ;
 wire \Tile_X0Y8_E2BEG[0] ;
 wire \Tile_X0Y8_E2BEG[1] ;
 wire \Tile_X0Y8_E2BEG[2] ;
 wire \Tile_X0Y8_E2BEG[3] ;
 wire \Tile_X0Y8_E2BEG[4] ;
 wire \Tile_X0Y8_E2BEG[5] ;
 wire \Tile_X0Y8_E2BEG[6] ;
 wire \Tile_X0Y8_E2BEG[7] ;
 wire \Tile_X0Y8_E2BEGb[0] ;
 wire \Tile_X0Y8_E2BEGb[1] ;
 wire \Tile_X0Y8_E2BEGb[2] ;
 wire \Tile_X0Y8_E2BEGb[3] ;
 wire \Tile_X0Y8_E2BEGb[4] ;
 wire \Tile_X0Y8_E2BEGb[5] ;
 wire \Tile_X0Y8_E2BEGb[6] ;
 wire \Tile_X0Y8_E2BEGb[7] ;
 wire \Tile_X0Y8_E6BEG[0] ;
 wire \Tile_X0Y8_E6BEG[10] ;
 wire \Tile_X0Y8_E6BEG[11] ;
 wire \Tile_X0Y8_E6BEG[1] ;
 wire \Tile_X0Y8_E6BEG[2] ;
 wire \Tile_X0Y8_E6BEG[3] ;
 wire \Tile_X0Y8_E6BEG[4] ;
 wire \Tile_X0Y8_E6BEG[5] ;
 wire \Tile_X0Y8_E6BEG[6] ;
 wire \Tile_X0Y8_E6BEG[7] ;
 wire \Tile_X0Y8_E6BEG[8] ;
 wire \Tile_X0Y8_E6BEG[9] ;
 wire \Tile_X0Y8_EE4BEG[0] ;
 wire \Tile_X0Y8_EE4BEG[10] ;
 wire \Tile_X0Y8_EE4BEG[11] ;
 wire \Tile_X0Y8_EE4BEG[12] ;
 wire \Tile_X0Y8_EE4BEG[13] ;
 wire \Tile_X0Y8_EE4BEG[14] ;
 wire \Tile_X0Y8_EE4BEG[15] ;
 wire \Tile_X0Y8_EE4BEG[1] ;
 wire \Tile_X0Y8_EE4BEG[2] ;
 wire \Tile_X0Y8_EE4BEG[3] ;
 wire \Tile_X0Y8_EE4BEG[4] ;
 wire \Tile_X0Y8_EE4BEG[5] ;
 wire \Tile_X0Y8_EE4BEG[6] ;
 wire \Tile_X0Y8_EE4BEG[7] ;
 wire \Tile_X0Y8_EE4BEG[8] ;
 wire \Tile_X0Y8_EE4BEG[9] ;
 wire \Tile_X0Y8_FrameData_O[0] ;
 wire \Tile_X0Y8_FrameData_O[10] ;
 wire \Tile_X0Y8_FrameData_O[11] ;
 wire \Tile_X0Y8_FrameData_O[12] ;
 wire \Tile_X0Y8_FrameData_O[13] ;
 wire \Tile_X0Y8_FrameData_O[14] ;
 wire \Tile_X0Y8_FrameData_O[15] ;
 wire \Tile_X0Y8_FrameData_O[16] ;
 wire \Tile_X0Y8_FrameData_O[17] ;
 wire \Tile_X0Y8_FrameData_O[18] ;
 wire \Tile_X0Y8_FrameData_O[19] ;
 wire \Tile_X0Y8_FrameData_O[1] ;
 wire \Tile_X0Y8_FrameData_O[20] ;
 wire \Tile_X0Y8_FrameData_O[21] ;
 wire \Tile_X0Y8_FrameData_O[22] ;
 wire \Tile_X0Y8_FrameData_O[23] ;
 wire \Tile_X0Y8_FrameData_O[24] ;
 wire \Tile_X0Y8_FrameData_O[25] ;
 wire \Tile_X0Y8_FrameData_O[26] ;
 wire \Tile_X0Y8_FrameData_O[27] ;
 wire \Tile_X0Y8_FrameData_O[28] ;
 wire \Tile_X0Y8_FrameData_O[29] ;
 wire \Tile_X0Y8_FrameData_O[2] ;
 wire \Tile_X0Y8_FrameData_O[30] ;
 wire \Tile_X0Y8_FrameData_O[31] ;
 wire \Tile_X0Y8_FrameData_O[3] ;
 wire \Tile_X0Y8_FrameData_O[4] ;
 wire \Tile_X0Y8_FrameData_O[5] ;
 wire \Tile_X0Y8_FrameData_O[6] ;
 wire \Tile_X0Y8_FrameData_O[7] ;
 wire \Tile_X0Y8_FrameData_O[8] ;
 wire \Tile_X0Y8_FrameData_O[9] ;
 wire \Tile_X0Y8_FrameStrobe_O[0] ;
 wire \Tile_X0Y8_FrameStrobe_O[10] ;
 wire \Tile_X0Y8_FrameStrobe_O[11] ;
 wire \Tile_X0Y8_FrameStrobe_O[12] ;
 wire \Tile_X0Y8_FrameStrobe_O[13] ;
 wire \Tile_X0Y8_FrameStrobe_O[14] ;
 wire \Tile_X0Y8_FrameStrobe_O[15] ;
 wire \Tile_X0Y8_FrameStrobe_O[16] ;
 wire \Tile_X0Y8_FrameStrobe_O[17] ;
 wire \Tile_X0Y8_FrameStrobe_O[18] ;
 wire \Tile_X0Y8_FrameStrobe_O[19] ;
 wire \Tile_X0Y8_FrameStrobe_O[1] ;
 wire \Tile_X0Y8_FrameStrobe_O[2] ;
 wire \Tile_X0Y8_FrameStrobe_O[3] ;
 wire \Tile_X0Y8_FrameStrobe_O[4] ;
 wire \Tile_X0Y8_FrameStrobe_O[5] ;
 wire \Tile_X0Y8_FrameStrobe_O[6] ;
 wire \Tile_X0Y8_FrameStrobe_O[7] ;
 wire \Tile_X0Y8_FrameStrobe_O[8] ;
 wire \Tile_X0Y8_FrameStrobe_O[9] ;
 wire Tile_X0Y8_UserCLKo;
 wire \Tile_X0Y9_E1BEG[0] ;
 wire \Tile_X0Y9_E1BEG[1] ;
 wire \Tile_X0Y9_E1BEG[2] ;
 wire \Tile_X0Y9_E1BEG[3] ;
 wire \Tile_X0Y9_E2BEG[0] ;
 wire \Tile_X0Y9_E2BEG[1] ;
 wire \Tile_X0Y9_E2BEG[2] ;
 wire \Tile_X0Y9_E2BEG[3] ;
 wire \Tile_X0Y9_E2BEG[4] ;
 wire \Tile_X0Y9_E2BEG[5] ;
 wire \Tile_X0Y9_E2BEG[6] ;
 wire \Tile_X0Y9_E2BEG[7] ;
 wire \Tile_X0Y9_E2BEGb[0] ;
 wire \Tile_X0Y9_E2BEGb[1] ;
 wire \Tile_X0Y9_E2BEGb[2] ;
 wire \Tile_X0Y9_E2BEGb[3] ;
 wire \Tile_X0Y9_E2BEGb[4] ;
 wire \Tile_X0Y9_E2BEGb[5] ;
 wire \Tile_X0Y9_E2BEGb[6] ;
 wire \Tile_X0Y9_E2BEGb[7] ;
 wire \Tile_X0Y9_E6BEG[0] ;
 wire \Tile_X0Y9_E6BEG[10] ;
 wire \Tile_X0Y9_E6BEG[11] ;
 wire \Tile_X0Y9_E6BEG[1] ;
 wire \Tile_X0Y9_E6BEG[2] ;
 wire \Tile_X0Y9_E6BEG[3] ;
 wire \Tile_X0Y9_E6BEG[4] ;
 wire \Tile_X0Y9_E6BEG[5] ;
 wire \Tile_X0Y9_E6BEG[6] ;
 wire \Tile_X0Y9_E6BEG[7] ;
 wire \Tile_X0Y9_E6BEG[8] ;
 wire \Tile_X0Y9_E6BEG[9] ;
 wire \Tile_X0Y9_EE4BEG[0] ;
 wire \Tile_X0Y9_EE4BEG[10] ;
 wire \Tile_X0Y9_EE4BEG[11] ;
 wire \Tile_X0Y9_EE4BEG[12] ;
 wire \Tile_X0Y9_EE4BEG[13] ;
 wire \Tile_X0Y9_EE4BEG[14] ;
 wire \Tile_X0Y9_EE4BEG[15] ;
 wire \Tile_X0Y9_EE4BEG[1] ;
 wire \Tile_X0Y9_EE4BEG[2] ;
 wire \Tile_X0Y9_EE4BEG[3] ;
 wire \Tile_X0Y9_EE4BEG[4] ;
 wire \Tile_X0Y9_EE4BEG[5] ;
 wire \Tile_X0Y9_EE4BEG[6] ;
 wire \Tile_X0Y9_EE4BEG[7] ;
 wire \Tile_X0Y9_EE4BEG[8] ;
 wire \Tile_X0Y9_EE4BEG[9] ;
 wire \Tile_X0Y9_FrameData_O[0] ;
 wire \Tile_X0Y9_FrameData_O[10] ;
 wire \Tile_X0Y9_FrameData_O[11] ;
 wire \Tile_X0Y9_FrameData_O[12] ;
 wire \Tile_X0Y9_FrameData_O[13] ;
 wire \Tile_X0Y9_FrameData_O[14] ;
 wire \Tile_X0Y9_FrameData_O[15] ;
 wire \Tile_X0Y9_FrameData_O[16] ;
 wire \Tile_X0Y9_FrameData_O[17] ;
 wire \Tile_X0Y9_FrameData_O[18] ;
 wire \Tile_X0Y9_FrameData_O[19] ;
 wire \Tile_X0Y9_FrameData_O[1] ;
 wire \Tile_X0Y9_FrameData_O[20] ;
 wire \Tile_X0Y9_FrameData_O[21] ;
 wire \Tile_X0Y9_FrameData_O[22] ;
 wire \Tile_X0Y9_FrameData_O[23] ;
 wire \Tile_X0Y9_FrameData_O[24] ;
 wire \Tile_X0Y9_FrameData_O[25] ;
 wire \Tile_X0Y9_FrameData_O[26] ;
 wire \Tile_X0Y9_FrameData_O[27] ;
 wire \Tile_X0Y9_FrameData_O[28] ;
 wire \Tile_X0Y9_FrameData_O[29] ;
 wire \Tile_X0Y9_FrameData_O[2] ;
 wire \Tile_X0Y9_FrameData_O[30] ;
 wire \Tile_X0Y9_FrameData_O[31] ;
 wire \Tile_X0Y9_FrameData_O[3] ;
 wire \Tile_X0Y9_FrameData_O[4] ;
 wire \Tile_X0Y9_FrameData_O[5] ;
 wire \Tile_X0Y9_FrameData_O[6] ;
 wire \Tile_X0Y9_FrameData_O[7] ;
 wire \Tile_X0Y9_FrameData_O[8] ;
 wire \Tile_X0Y9_FrameData_O[9] ;
 wire \Tile_X0Y9_FrameStrobe_O[0] ;
 wire \Tile_X0Y9_FrameStrobe_O[10] ;
 wire \Tile_X0Y9_FrameStrobe_O[11] ;
 wire \Tile_X0Y9_FrameStrobe_O[12] ;
 wire \Tile_X0Y9_FrameStrobe_O[13] ;
 wire \Tile_X0Y9_FrameStrobe_O[14] ;
 wire \Tile_X0Y9_FrameStrobe_O[15] ;
 wire \Tile_X0Y9_FrameStrobe_O[16] ;
 wire \Tile_X0Y9_FrameStrobe_O[17] ;
 wire \Tile_X0Y9_FrameStrobe_O[18] ;
 wire \Tile_X0Y9_FrameStrobe_O[19] ;
 wire \Tile_X0Y9_FrameStrobe_O[1] ;
 wire \Tile_X0Y9_FrameStrobe_O[2] ;
 wire \Tile_X0Y9_FrameStrobe_O[3] ;
 wire \Tile_X0Y9_FrameStrobe_O[4] ;
 wire \Tile_X0Y9_FrameStrobe_O[5] ;
 wire \Tile_X0Y9_FrameStrobe_O[6] ;
 wire \Tile_X0Y9_FrameStrobe_O[7] ;
 wire \Tile_X0Y9_FrameStrobe_O[8] ;
 wire \Tile_X0Y9_FrameStrobe_O[9] ;
 wire Tile_X0Y9_UserCLKo;
 wire \Tile_X10Y0_FrameData_O[0] ;
 wire \Tile_X10Y0_FrameData_O[10] ;
 wire \Tile_X10Y0_FrameData_O[11] ;
 wire \Tile_X10Y0_FrameData_O[12] ;
 wire \Tile_X10Y0_FrameData_O[13] ;
 wire \Tile_X10Y0_FrameData_O[14] ;
 wire \Tile_X10Y0_FrameData_O[15] ;
 wire \Tile_X10Y0_FrameData_O[16] ;
 wire \Tile_X10Y0_FrameData_O[17] ;
 wire \Tile_X10Y0_FrameData_O[18] ;
 wire \Tile_X10Y0_FrameData_O[19] ;
 wire \Tile_X10Y0_FrameData_O[1] ;
 wire \Tile_X10Y0_FrameData_O[20] ;
 wire \Tile_X10Y0_FrameData_O[21] ;
 wire \Tile_X10Y0_FrameData_O[22] ;
 wire \Tile_X10Y0_FrameData_O[23] ;
 wire \Tile_X10Y0_FrameData_O[24] ;
 wire \Tile_X10Y0_FrameData_O[25] ;
 wire \Tile_X10Y0_FrameData_O[26] ;
 wire \Tile_X10Y0_FrameData_O[27] ;
 wire \Tile_X10Y0_FrameData_O[28] ;
 wire \Tile_X10Y0_FrameData_O[29] ;
 wire \Tile_X10Y0_FrameData_O[2] ;
 wire \Tile_X10Y0_FrameData_O[30] ;
 wire \Tile_X10Y0_FrameData_O[31] ;
 wire \Tile_X10Y0_FrameData_O[3] ;
 wire \Tile_X10Y0_FrameData_O[4] ;
 wire \Tile_X10Y0_FrameData_O[5] ;
 wire \Tile_X10Y0_FrameData_O[6] ;
 wire \Tile_X10Y0_FrameData_O[7] ;
 wire \Tile_X10Y0_FrameData_O[8] ;
 wire \Tile_X10Y0_FrameData_O[9] ;
 wire \Tile_X10Y0_FrameStrobe_O[0] ;
 wire \Tile_X10Y0_FrameStrobe_O[10] ;
 wire \Tile_X10Y0_FrameStrobe_O[11] ;
 wire \Tile_X10Y0_FrameStrobe_O[12] ;
 wire \Tile_X10Y0_FrameStrobe_O[13] ;
 wire \Tile_X10Y0_FrameStrobe_O[14] ;
 wire \Tile_X10Y0_FrameStrobe_O[15] ;
 wire \Tile_X10Y0_FrameStrobe_O[16] ;
 wire \Tile_X10Y0_FrameStrobe_O[17] ;
 wire \Tile_X10Y0_FrameStrobe_O[18] ;
 wire \Tile_X10Y0_FrameStrobe_O[19] ;
 wire \Tile_X10Y0_FrameStrobe_O[1] ;
 wire \Tile_X10Y0_FrameStrobe_O[2] ;
 wire \Tile_X10Y0_FrameStrobe_O[3] ;
 wire \Tile_X10Y0_FrameStrobe_O[4] ;
 wire \Tile_X10Y0_FrameStrobe_O[5] ;
 wire \Tile_X10Y0_FrameStrobe_O[6] ;
 wire \Tile_X10Y0_FrameStrobe_O[7] ;
 wire \Tile_X10Y0_FrameStrobe_O[8] ;
 wire \Tile_X10Y0_FrameStrobe_O[9] ;
 wire \Tile_X10Y0_S1BEG[0] ;
 wire \Tile_X10Y0_S1BEG[1] ;
 wire \Tile_X10Y0_S1BEG[2] ;
 wire \Tile_X10Y0_S1BEG[3] ;
 wire \Tile_X10Y0_S2BEG[0] ;
 wire \Tile_X10Y0_S2BEG[1] ;
 wire \Tile_X10Y0_S2BEG[2] ;
 wire \Tile_X10Y0_S2BEG[3] ;
 wire \Tile_X10Y0_S2BEG[4] ;
 wire \Tile_X10Y0_S2BEG[5] ;
 wire \Tile_X10Y0_S2BEG[6] ;
 wire \Tile_X10Y0_S2BEG[7] ;
 wire \Tile_X10Y0_S2BEGb[0] ;
 wire \Tile_X10Y0_S2BEGb[1] ;
 wire \Tile_X10Y0_S2BEGb[2] ;
 wire \Tile_X10Y0_S2BEGb[3] ;
 wire \Tile_X10Y0_S2BEGb[4] ;
 wire \Tile_X10Y0_S2BEGb[5] ;
 wire \Tile_X10Y0_S2BEGb[6] ;
 wire \Tile_X10Y0_S2BEGb[7] ;
 wire \Tile_X10Y0_S4BEG[0] ;
 wire \Tile_X10Y0_S4BEG[10] ;
 wire \Tile_X10Y0_S4BEG[11] ;
 wire \Tile_X10Y0_S4BEG[12] ;
 wire \Tile_X10Y0_S4BEG[13] ;
 wire \Tile_X10Y0_S4BEG[14] ;
 wire \Tile_X10Y0_S4BEG[15] ;
 wire \Tile_X10Y0_S4BEG[1] ;
 wire \Tile_X10Y0_S4BEG[2] ;
 wire \Tile_X10Y0_S4BEG[3] ;
 wire \Tile_X10Y0_S4BEG[4] ;
 wire \Tile_X10Y0_S4BEG[5] ;
 wire \Tile_X10Y0_S4BEG[6] ;
 wire \Tile_X10Y0_S4BEG[7] ;
 wire \Tile_X10Y0_S4BEG[8] ;
 wire \Tile_X10Y0_S4BEG[9] ;
 wire Tile_X10Y0_UserCLKo;
 wire \Tile_X10Y10_FrameData_O[0] ;
 wire \Tile_X10Y10_FrameData_O[10] ;
 wire \Tile_X10Y10_FrameData_O[11] ;
 wire \Tile_X10Y10_FrameData_O[12] ;
 wire \Tile_X10Y10_FrameData_O[13] ;
 wire \Tile_X10Y10_FrameData_O[14] ;
 wire \Tile_X10Y10_FrameData_O[15] ;
 wire \Tile_X10Y10_FrameData_O[16] ;
 wire \Tile_X10Y10_FrameData_O[17] ;
 wire \Tile_X10Y10_FrameData_O[18] ;
 wire \Tile_X10Y10_FrameData_O[19] ;
 wire \Tile_X10Y10_FrameData_O[1] ;
 wire \Tile_X10Y10_FrameData_O[20] ;
 wire \Tile_X10Y10_FrameData_O[21] ;
 wire \Tile_X10Y10_FrameData_O[22] ;
 wire \Tile_X10Y10_FrameData_O[23] ;
 wire \Tile_X10Y10_FrameData_O[24] ;
 wire \Tile_X10Y10_FrameData_O[25] ;
 wire \Tile_X10Y10_FrameData_O[26] ;
 wire \Tile_X10Y10_FrameData_O[27] ;
 wire \Tile_X10Y10_FrameData_O[28] ;
 wire \Tile_X10Y10_FrameData_O[29] ;
 wire \Tile_X10Y10_FrameData_O[2] ;
 wire \Tile_X10Y10_FrameData_O[30] ;
 wire \Tile_X10Y10_FrameData_O[31] ;
 wire \Tile_X10Y10_FrameData_O[3] ;
 wire \Tile_X10Y10_FrameData_O[4] ;
 wire \Tile_X10Y10_FrameData_O[5] ;
 wire \Tile_X10Y10_FrameData_O[6] ;
 wire \Tile_X10Y10_FrameData_O[7] ;
 wire \Tile_X10Y10_FrameData_O[8] ;
 wire \Tile_X10Y10_FrameData_O[9] ;
 wire \Tile_X10Y10_S1BEG[0] ;
 wire \Tile_X10Y10_S1BEG[1] ;
 wire \Tile_X10Y10_S1BEG[2] ;
 wire \Tile_X10Y10_S1BEG[3] ;
 wire \Tile_X10Y10_S2BEG[0] ;
 wire \Tile_X10Y10_S2BEG[1] ;
 wire \Tile_X10Y10_S2BEG[2] ;
 wire \Tile_X10Y10_S2BEG[3] ;
 wire \Tile_X10Y10_S2BEG[4] ;
 wire \Tile_X10Y10_S2BEG[5] ;
 wire \Tile_X10Y10_S2BEG[6] ;
 wire \Tile_X10Y10_S2BEG[7] ;
 wire \Tile_X10Y10_S2BEGb[0] ;
 wire \Tile_X10Y10_S2BEGb[1] ;
 wire \Tile_X10Y10_S2BEGb[2] ;
 wire \Tile_X10Y10_S2BEGb[3] ;
 wire \Tile_X10Y10_S2BEGb[4] ;
 wire \Tile_X10Y10_S2BEGb[5] ;
 wire \Tile_X10Y10_S2BEGb[6] ;
 wire \Tile_X10Y10_S2BEGb[7] ;
 wire \Tile_X10Y10_S4BEG[0] ;
 wire \Tile_X10Y10_S4BEG[10] ;
 wire \Tile_X10Y10_S4BEG[11] ;
 wire \Tile_X10Y10_S4BEG[12] ;
 wire \Tile_X10Y10_S4BEG[13] ;
 wire \Tile_X10Y10_S4BEG[14] ;
 wire \Tile_X10Y10_S4BEG[15] ;
 wire \Tile_X10Y10_S4BEG[1] ;
 wire \Tile_X10Y10_S4BEG[2] ;
 wire \Tile_X10Y10_S4BEG[3] ;
 wire \Tile_X10Y10_S4BEG[4] ;
 wire \Tile_X10Y10_S4BEG[5] ;
 wire \Tile_X10Y10_S4BEG[6] ;
 wire \Tile_X10Y10_S4BEG[7] ;
 wire \Tile_X10Y10_S4BEG[8] ;
 wire \Tile_X10Y10_S4BEG[9] ;
 wire \Tile_X10Y10_W1BEG[0] ;
 wire \Tile_X10Y10_W1BEG[1] ;
 wire \Tile_X10Y10_W1BEG[2] ;
 wire \Tile_X10Y10_W1BEG[3] ;
 wire \Tile_X10Y10_W2BEG[0] ;
 wire \Tile_X10Y10_W2BEG[1] ;
 wire \Tile_X10Y10_W2BEG[2] ;
 wire \Tile_X10Y10_W2BEG[3] ;
 wire \Tile_X10Y10_W2BEG[4] ;
 wire \Tile_X10Y10_W2BEG[5] ;
 wire \Tile_X10Y10_W2BEG[6] ;
 wire \Tile_X10Y10_W2BEG[7] ;
 wire \Tile_X10Y10_W2BEGb[0] ;
 wire \Tile_X10Y10_W2BEGb[1] ;
 wire \Tile_X10Y10_W2BEGb[2] ;
 wire \Tile_X10Y10_W2BEGb[3] ;
 wire \Tile_X10Y10_W2BEGb[4] ;
 wire \Tile_X10Y10_W2BEGb[5] ;
 wire \Tile_X10Y10_W2BEGb[6] ;
 wire \Tile_X10Y10_W2BEGb[7] ;
 wire \Tile_X10Y10_W6BEG[0] ;
 wire \Tile_X10Y10_W6BEG[10] ;
 wire \Tile_X10Y10_W6BEG[11] ;
 wire \Tile_X10Y10_W6BEG[1] ;
 wire \Tile_X10Y10_W6BEG[2] ;
 wire \Tile_X10Y10_W6BEG[3] ;
 wire \Tile_X10Y10_W6BEG[4] ;
 wire \Tile_X10Y10_W6BEG[5] ;
 wire \Tile_X10Y10_W6BEG[6] ;
 wire \Tile_X10Y10_W6BEG[7] ;
 wire \Tile_X10Y10_W6BEG[8] ;
 wire \Tile_X10Y10_W6BEG[9] ;
 wire \Tile_X10Y10_WW4BEG[0] ;
 wire \Tile_X10Y10_WW4BEG[10] ;
 wire \Tile_X10Y10_WW4BEG[11] ;
 wire \Tile_X10Y10_WW4BEG[12] ;
 wire \Tile_X10Y10_WW4BEG[13] ;
 wire \Tile_X10Y10_WW4BEG[14] ;
 wire \Tile_X10Y10_WW4BEG[15] ;
 wire \Tile_X10Y10_WW4BEG[1] ;
 wire \Tile_X10Y10_WW4BEG[2] ;
 wire \Tile_X10Y10_WW4BEG[3] ;
 wire \Tile_X10Y10_WW4BEG[4] ;
 wire \Tile_X10Y10_WW4BEG[5] ;
 wire \Tile_X10Y10_WW4BEG[6] ;
 wire \Tile_X10Y10_WW4BEG[7] ;
 wire \Tile_X10Y10_WW4BEG[8] ;
 wire \Tile_X10Y10_WW4BEG[9] ;
 wire \Tile_X10Y11_FrameData_O[0] ;
 wire \Tile_X10Y11_FrameData_O[10] ;
 wire \Tile_X10Y11_FrameData_O[11] ;
 wire \Tile_X10Y11_FrameData_O[12] ;
 wire \Tile_X10Y11_FrameData_O[13] ;
 wire \Tile_X10Y11_FrameData_O[14] ;
 wire \Tile_X10Y11_FrameData_O[15] ;
 wire \Tile_X10Y11_FrameData_O[16] ;
 wire \Tile_X10Y11_FrameData_O[17] ;
 wire \Tile_X10Y11_FrameData_O[18] ;
 wire \Tile_X10Y11_FrameData_O[19] ;
 wire \Tile_X10Y11_FrameData_O[1] ;
 wire \Tile_X10Y11_FrameData_O[20] ;
 wire \Tile_X10Y11_FrameData_O[21] ;
 wire \Tile_X10Y11_FrameData_O[22] ;
 wire \Tile_X10Y11_FrameData_O[23] ;
 wire \Tile_X10Y11_FrameData_O[24] ;
 wire \Tile_X10Y11_FrameData_O[25] ;
 wire \Tile_X10Y11_FrameData_O[26] ;
 wire \Tile_X10Y11_FrameData_O[27] ;
 wire \Tile_X10Y11_FrameData_O[28] ;
 wire \Tile_X10Y11_FrameData_O[29] ;
 wire \Tile_X10Y11_FrameData_O[2] ;
 wire \Tile_X10Y11_FrameData_O[30] ;
 wire \Tile_X10Y11_FrameData_O[31] ;
 wire \Tile_X10Y11_FrameData_O[3] ;
 wire \Tile_X10Y11_FrameData_O[4] ;
 wire \Tile_X10Y11_FrameData_O[5] ;
 wire \Tile_X10Y11_FrameData_O[6] ;
 wire \Tile_X10Y11_FrameData_O[7] ;
 wire \Tile_X10Y11_FrameData_O[8] ;
 wire \Tile_X10Y11_FrameData_O[9] ;
 wire \Tile_X10Y11_FrameStrobe_O[0] ;
 wire \Tile_X10Y11_FrameStrobe_O[10] ;
 wire \Tile_X10Y11_FrameStrobe_O[11] ;
 wire \Tile_X10Y11_FrameStrobe_O[12] ;
 wire \Tile_X10Y11_FrameStrobe_O[13] ;
 wire \Tile_X10Y11_FrameStrobe_O[14] ;
 wire \Tile_X10Y11_FrameStrobe_O[15] ;
 wire \Tile_X10Y11_FrameStrobe_O[16] ;
 wire \Tile_X10Y11_FrameStrobe_O[17] ;
 wire \Tile_X10Y11_FrameStrobe_O[18] ;
 wire \Tile_X10Y11_FrameStrobe_O[19] ;
 wire \Tile_X10Y11_FrameStrobe_O[1] ;
 wire \Tile_X10Y11_FrameStrobe_O[2] ;
 wire \Tile_X10Y11_FrameStrobe_O[3] ;
 wire \Tile_X10Y11_FrameStrobe_O[4] ;
 wire \Tile_X10Y11_FrameStrobe_O[5] ;
 wire \Tile_X10Y11_FrameStrobe_O[6] ;
 wire \Tile_X10Y11_FrameStrobe_O[7] ;
 wire \Tile_X10Y11_FrameStrobe_O[8] ;
 wire \Tile_X10Y11_FrameStrobe_O[9] ;
 wire \Tile_X10Y11_N1BEG[0] ;
 wire \Tile_X10Y11_N1BEG[1] ;
 wire \Tile_X10Y11_N1BEG[2] ;
 wire \Tile_X10Y11_N1BEG[3] ;
 wire \Tile_X10Y11_N2BEG[0] ;
 wire \Tile_X10Y11_N2BEG[1] ;
 wire \Tile_X10Y11_N2BEG[2] ;
 wire \Tile_X10Y11_N2BEG[3] ;
 wire \Tile_X10Y11_N2BEG[4] ;
 wire \Tile_X10Y11_N2BEG[5] ;
 wire \Tile_X10Y11_N2BEG[6] ;
 wire \Tile_X10Y11_N2BEG[7] ;
 wire \Tile_X10Y11_N2BEGb[0] ;
 wire \Tile_X10Y11_N2BEGb[1] ;
 wire \Tile_X10Y11_N2BEGb[2] ;
 wire \Tile_X10Y11_N2BEGb[3] ;
 wire \Tile_X10Y11_N2BEGb[4] ;
 wire \Tile_X10Y11_N2BEGb[5] ;
 wire \Tile_X10Y11_N2BEGb[6] ;
 wire \Tile_X10Y11_N2BEGb[7] ;
 wire \Tile_X10Y11_N4BEG[0] ;
 wire \Tile_X10Y11_N4BEG[10] ;
 wire \Tile_X10Y11_N4BEG[11] ;
 wire \Tile_X10Y11_N4BEG[12] ;
 wire \Tile_X10Y11_N4BEG[13] ;
 wire \Tile_X10Y11_N4BEG[14] ;
 wire \Tile_X10Y11_N4BEG[15] ;
 wire \Tile_X10Y11_N4BEG[1] ;
 wire \Tile_X10Y11_N4BEG[2] ;
 wire \Tile_X10Y11_N4BEG[3] ;
 wire \Tile_X10Y11_N4BEG[4] ;
 wire \Tile_X10Y11_N4BEG[5] ;
 wire \Tile_X10Y11_N4BEG[6] ;
 wire \Tile_X10Y11_N4BEG[7] ;
 wire \Tile_X10Y11_N4BEG[8] ;
 wire \Tile_X10Y11_N4BEG[9] ;
 wire Tile_X10Y11_UserCLKo;
 wire \Tile_X10Y11_W1BEG[0] ;
 wire \Tile_X10Y11_W1BEG[1] ;
 wire \Tile_X10Y11_W1BEG[2] ;
 wire \Tile_X10Y11_W1BEG[3] ;
 wire \Tile_X10Y11_W2BEG[0] ;
 wire \Tile_X10Y11_W2BEG[1] ;
 wire \Tile_X10Y11_W2BEG[2] ;
 wire \Tile_X10Y11_W2BEG[3] ;
 wire \Tile_X10Y11_W2BEG[4] ;
 wire \Tile_X10Y11_W2BEG[5] ;
 wire \Tile_X10Y11_W2BEG[6] ;
 wire \Tile_X10Y11_W2BEG[7] ;
 wire \Tile_X10Y11_W2BEGb[0] ;
 wire \Tile_X10Y11_W2BEGb[1] ;
 wire \Tile_X10Y11_W2BEGb[2] ;
 wire \Tile_X10Y11_W2BEGb[3] ;
 wire \Tile_X10Y11_W2BEGb[4] ;
 wire \Tile_X10Y11_W2BEGb[5] ;
 wire \Tile_X10Y11_W2BEGb[6] ;
 wire \Tile_X10Y11_W2BEGb[7] ;
 wire \Tile_X10Y11_W6BEG[0] ;
 wire \Tile_X10Y11_W6BEG[10] ;
 wire \Tile_X10Y11_W6BEG[11] ;
 wire \Tile_X10Y11_W6BEG[1] ;
 wire \Tile_X10Y11_W6BEG[2] ;
 wire \Tile_X10Y11_W6BEG[3] ;
 wire \Tile_X10Y11_W6BEG[4] ;
 wire \Tile_X10Y11_W6BEG[5] ;
 wire \Tile_X10Y11_W6BEG[6] ;
 wire \Tile_X10Y11_W6BEG[7] ;
 wire \Tile_X10Y11_W6BEG[8] ;
 wire \Tile_X10Y11_W6BEG[9] ;
 wire \Tile_X10Y11_WW4BEG[0] ;
 wire \Tile_X10Y11_WW4BEG[10] ;
 wire \Tile_X10Y11_WW4BEG[11] ;
 wire \Tile_X10Y11_WW4BEG[12] ;
 wire \Tile_X10Y11_WW4BEG[13] ;
 wire \Tile_X10Y11_WW4BEG[14] ;
 wire \Tile_X10Y11_WW4BEG[15] ;
 wire \Tile_X10Y11_WW4BEG[1] ;
 wire \Tile_X10Y11_WW4BEG[2] ;
 wire \Tile_X10Y11_WW4BEG[3] ;
 wire \Tile_X10Y11_WW4BEG[4] ;
 wire \Tile_X10Y11_WW4BEG[5] ;
 wire \Tile_X10Y11_WW4BEG[6] ;
 wire \Tile_X10Y11_WW4BEG[7] ;
 wire \Tile_X10Y11_WW4BEG[8] ;
 wire \Tile_X10Y11_WW4BEG[9] ;
 wire \Tile_X10Y12_FrameData_O[0] ;
 wire \Tile_X10Y12_FrameData_O[10] ;
 wire \Tile_X10Y12_FrameData_O[11] ;
 wire \Tile_X10Y12_FrameData_O[12] ;
 wire \Tile_X10Y12_FrameData_O[13] ;
 wire \Tile_X10Y12_FrameData_O[14] ;
 wire \Tile_X10Y12_FrameData_O[15] ;
 wire \Tile_X10Y12_FrameData_O[16] ;
 wire \Tile_X10Y12_FrameData_O[17] ;
 wire \Tile_X10Y12_FrameData_O[18] ;
 wire \Tile_X10Y12_FrameData_O[19] ;
 wire \Tile_X10Y12_FrameData_O[1] ;
 wire \Tile_X10Y12_FrameData_O[20] ;
 wire \Tile_X10Y12_FrameData_O[21] ;
 wire \Tile_X10Y12_FrameData_O[22] ;
 wire \Tile_X10Y12_FrameData_O[23] ;
 wire \Tile_X10Y12_FrameData_O[24] ;
 wire \Tile_X10Y12_FrameData_O[25] ;
 wire \Tile_X10Y12_FrameData_O[26] ;
 wire \Tile_X10Y12_FrameData_O[27] ;
 wire \Tile_X10Y12_FrameData_O[28] ;
 wire \Tile_X10Y12_FrameData_O[29] ;
 wire \Tile_X10Y12_FrameData_O[2] ;
 wire \Tile_X10Y12_FrameData_O[30] ;
 wire \Tile_X10Y12_FrameData_O[31] ;
 wire \Tile_X10Y12_FrameData_O[3] ;
 wire \Tile_X10Y12_FrameData_O[4] ;
 wire \Tile_X10Y12_FrameData_O[5] ;
 wire \Tile_X10Y12_FrameData_O[6] ;
 wire \Tile_X10Y12_FrameData_O[7] ;
 wire \Tile_X10Y12_FrameData_O[8] ;
 wire \Tile_X10Y12_FrameData_O[9] ;
 wire \Tile_X10Y12_S1BEG[0] ;
 wire \Tile_X10Y12_S1BEG[1] ;
 wire \Tile_X10Y12_S1BEG[2] ;
 wire \Tile_X10Y12_S1BEG[3] ;
 wire \Tile_X10Y12_S2BEG[0] ;
 wire \Tile_X10Y12_S2BEG[1] ;
 wire \Tile_X10Y12_S2BEG[2] ;
 wire \Tile_X10Y12_S2BEG[3] ;
 wire \Tile_X10Y12_S2BEG[4] ;
 wire \Tile_X10Y12_S2BEG[5] ;
 wire \Tile_X10Y12_S2BEG[6] ;
 wire \Tile_X10Y12_S2BEG[7] ;
 wire \Tile_X10Y12_S2BEGb[0] ;
 wire \Tile_X10Y12_S2BEGb[1] ;
 wire \Tile_X10Y12_S2BEGb[2] ;
 wire \Tile_X10Y12_S2BEGb[3] ;
 wire \Tile_X10Y12_S2BEGb[4] ;
 wire \Tile_X10Y12_S2BEGb[5] ;
 wire \Tile_X10Y12_S2BEGb[6] ;
 wire \Tile_X10Y12_S2BEGb[7] ;
 wire \Tile_X10Y12_S4BEG[0] ;
 wire \Tile_X10Y12_S4BEG[10] ;
 wire \Tile_X10Y12_S4BEG[11] ;
 wire \Tile_X10Y12_S4BEG[12] ;
 wire \Tile_X10Y12_S4BEG[13] ;
 wire \Tile_X10Y12_S4BEG[14] ;
 wire \Tile_X10Y12_S4BEG[15] ;
 wire \Tile_X10Y12_S4BEG[1] ;
 wire \Tile_X10Y12_S4BEG[2] ;
 wire \Tile_X10Y12_S4BEG[3] ;
 wire \Tile_X10Y12_S4BEG[4] ;
 wire \Tile_X10Y12_S4BEG[5] ;
 wire \Tile_X10Y12_S4BEG[6] ;
 wire \Tile_X10Y12_S4BEG[7] ;
 wire \Tile_X10Y12_S4BEG[8] ;
 wire \Tile_X10Y12_S4BEG[9] ;
 wire \Tile_X10Y12_W1BEG[0] ;
 wire \Tile_X10Y12_W1BEG[1] ;
 wire \Tile_X10Y12_W1BEG[2] ;
 wire \Tile_X10Y12_W1BEG[3] ;
 wire \Tile_X10Y12_W2BEG[0] ;
 wire \Tile_X10Y12_W2BEG[1] ;
 wire \Tile_X10Y12_W2BEG[2] ;
 wire \Tile_X10Y12_W2BEG[3] ;
 wire \Tile_X10Y12_W2BEG[4] ;
 wire \Tile_X10Y12_W2BEG[5] ;
 wire \Tile_X10Y12_W2BEG[6] ;
 wire \Tile_X10Y12_W2BEG[7] ;
 wire \Tile_X10Y12_W2BEGb[0] ;
 wire \Tile_X10Y12_W2BEGb[1] ;
 wire \Tile_X10Y12_W2BEGb[2] ;
 wire \Tile_X10Y12_W2BEGb[3] ;
 wire \Tile_X10Y12_W2BEGb[4] ;
 wire \Tile_X10Y12_W2BEGb[5] ;
 wire \Tile_X10Y12_W2BEGb[6] ;
 wire \Tile_X10Y12_W2BEGb[7] ;
 wire \Tile_X10Y12_W6BEG[0] ;
 wire \Tile_X10Y12_W6BEG[10] ;
 wire \Tile_X10Y12_W6BEG[11] ;
 wire \Tile_X10Y12_W6BEG[1] ;
 wire \Tile_X10Y12_W6BEG[2] ;
 wire \Tile_X10Y12_W6BEG[3] ;
 wire \Tile_X10Y12_W6BEG[4] ;
 wire \Tile_X10Y12_W6BEG[5] ;
 wire \Tile_X10Y12_W6BEG[6] ;
 wire \Tile_X10Y12_W6BEG[7] ;
 wire \Tile_X10Y12_W6BEG[8] ;
 wire \Tile_X10Y12_W6BEG[9] ;
 wire \Tile_X10Y12_WW4BEG[0] ;
 wire \Tile_X10Y12_WW4BEG[10] ;
 wire \Tile_X10Y12_WW4BEG[11] ;
 wire \Tile_X10Y12_WW4BEG[12] ;
 wire \Tile_X10Y12_WW4BEG[13] ;
 wire \Tile_X10Y12_WW4BEG[14] ;
 wire \Tile_X10Y12_WW4BEG[15] ;
 wire \Tile_X10Y12_WW4BEG[1] ;
 wire \Tile_X10Y12_WW4BEG[2] ;
 wire \Tile_X10Y12_WW4BEG[3] ;
 wire \Tile_X10Y12_WW4BEG[4] ;
 wire \Tile_X10Y12_WW4BEG[5] ;
 wire \Tile_X10Y12_WW4BEG[6] ;
 wire \Tile_X10Y12_WW4BEG[7] ;
 wire \Tile_X10Y12_WW4BEG[8] ;
 wire \Tile_X10Y12_WW4BEG[9] ;
 wire \Tile_X10Y13_FrameData_O[0] ;
 wire \Tile_X10Y13_FrameData_O[10] ;
 wire \Tile_X10Y13_FrameData_O[11] ;
 wire \Tile_X10Y13_FrameData_O[12] ;
 wire \Tile_X10Y13_FrameData_O[13] ;
 wire \Tile_X10Y13_FrameData_O[14] ;
 wire \Tile_X10Y13_FrameData_O[15] ;
 wire \Tile_X10Y13_FrameData_O[16] ;
 wire \Tile_X10Y13_FrameData_O[17] ;
 wire \Tile_X10Y13_FrameData_O[18] ;
 wire \Tile_X10Y13_FrameData_O[19] ;
 wire \Tile_X10Y13_FrameData_O[1] ;
 wire \Tile_X10Y13_FrameData_O[20] ;
 wire \Tile_X10Y13_FrameData_O[21] ;
 wire \Tile_X10Y13_FrameData_O[22] ;
 wire \Tile_X10Y13_FrameData_O[23] ;
 wire \Tile_X10Y13_FrameData_O[24] ;
 wire \Tile_X10Y13_FrameData_O[25] ;
 wire \Tile_X10Y13_FrameData_O[26] ;
 wire \Tile_X10Y13_FrameData_O[27] ;
 wire \Tile_X10Y13_FrameData_O[28] ;
 wire \Tile_X10Y13_FrameData_O[29] ;
 wire \Tile_X10Y13_FrameData_O[2] ;
 wire \Tile_X10Y13_FrameData_O[30] ;
 wire \Tile_X10Y13_FrameData_O[31] ;
 wire \Tile_X10Y13_FrameData_O[3] ;
 wire \Tile_X10Y13_FrameData_O[4] ;
 wire \Tile_X10Y13_FrameData_O[5] ;
 wire \Tile_X10Y13_FrameData_O[6] ;
 wire \Tile_X10Y13_FrameData_O[7] ;
 wire \Tile_X10Y13_FrameData_O[8] ;
 wire \Tile_X10Y13_FrameData_O[9] ;
 wire \Tile_X10Y13_FrameStrobe_O[0] ;
 wire \Tile_X10Y13_FrameStrobe_O[10] ;
 wire \Tile_X10Y13_FrameStrobe_O[11] ;
 wire \Tile_X10Y13_FrameStrobe_O[12] ;
 wire \Tile_X10Y13_FrameStrobe_O[13] ;
 wire \Tile_X10Y13_FrameStrobe_O[14] ;
 wire \Tile_X10Y13_FrameStrobe_O[15] ;
 wire \Tile_X10Y13_FrameStrobe_O[16] ;
 wire \Tile_X10Y13_FrameStrobe_O[17] ;
 wire \Tile_X10Y13_FrameStrobe_O[18] ;
 wire \Tile_X10Y13_FrameStrobe_O[19] ;
 wire \Tile_X10Y13_FrameStrobe_O[1] ;
 wire \Tile_X10Y13_FrameStrobe_O[2] ;
 wire \Tile_X10Y13_FrameStrobe_O[3] ;
 wire \Tile_X10Y13_FrameStrobe_O[4] ;
 wire \Tile_X10Y13_FrameStrobe_O[5] ;
 wire \Tile_X10Y13_FrameStrobe_O[6] ;
 wire \Tile_X10Y13_FrameStrobe_O[7] ;
 wire \Tile_X10Y13_FrameStrobe_O[8] ;
 wire \Tile_X10Y13_FrameStrobe_O[9] ;
 wire \Tile_X10Y13_N1BEG[0] ;
 wire \Tile_X10Y13_N1BEG[1] ;
 wire \Tile_X10Y13_N1BEG[2] ;
 wire \Tile_X10Y13_N1BEG[3] ;
 wire \Tile_X10Y13_N2BEG[0] ;
 wire \Tile_X10Y13_N2BEG[1] ;
 wire \Tile_X10Y13_N2BEG[2] ;
 wire \Tile_X10Y13_N2BEG[3] ;
 wire \Tile_X10Y13_N2BEG[4] ;
 wire \Tile_X10Y13_N2BEG[5] ;
 wire \Tile_X10Y13_N2BEG[6] ;
 wire \Tile_X10Y13_N2BEG[7] ;
 wire \Tile_X10Y13_N2BEGb[0] ;
 wire \Tile_X10Y13_N2BEGb[1] ;
 wire \Tile_X10Y13_N2BEGb[2] ;
 wire \Tile_X10Y13_N2BEGb[3] ;
 wire \Tile_X10Y13_N2BEGb[4] ;
 wire \Tile_X10Y13_N2BEGb[5] ;
 wire \Tile_X10Y13_N2BEGb[6] ;
 wire \Tile_X10Y13_N2BEGb[7] ;
 wire \Tile_X10Y13_N4BEG[0] ;
 wire \Tile_X10Y13_N4BEG[10] ;
 wire \Tile_X10Y13_N4BEG[11] ;
 wire \Tile_X10Y13_N4BEG[12] ;
 wire \Tile_X10Y13_N4BEG[13] ;
 wire \Tile_X10Y13_N4BEG[14] ;
 wire \Tile_X10Y13_N4BEG[15] ;
 wire \Tile_X10Y13_N4BEG[1] ;
 wire \Tile_X10Y13_N4BEG[2] ;
 wire \Tile_X10Y13_N4BEG[3] ;
 wire \Tile_X10Y13_N4BEG[4] ;
 wire \Tile_X10Y13_N4BEG[5] ;
 wire \Tile_X10Y13_N4BEG[6] ;
 wire \Tile_X10Y13_N4BEG[7] ;
 wire \Tile_X10Y13_N4BEG[8] ;
 wire \Tile_X10Y13_N4BEG[9] ;
 wire Tile_X10Y13_UserCLKo;
 wire \Tile_X10Y13_W1BEG[0] ;
 wire \Tile_X10Y13_W1BEG[1] ;
 wire \Tile_X10Y13_W1BEG[2] ;
 wire \Tile_X10Y13_W1BEG[3] ;
 wire \Tile_X10Y13_W2BEG[0] ;
 wire \Tile_X10Y13_W2BEG[1] ;
 wire \Tile_X10Y13_W2BEG[2] ;
 wire \Tile_X10Y13_W2BEG[3] ;
 wire \Tile_X10Y13_W2BEG[4] ;
 wire \Tile_X10Y13_W2BEG[5] ;
 wire \Tile_X10Y13_W2BEG[6] ;
 wire \Tile_X10Y13_W2BEG[7] ;
 wire \Tile_X10Y13_W2BEGb[0] ;
 wire \Tile_X10Y13_W2BEGb[1] ;
 wire \Tile_X10Y13_W2BEGb[2] ;
 wire \Tile_X10Y13_W2BEGb[3] ;
 wire \Tile_X10Y13_W2BEGb[4] ;
 wire \Tile_X10Y13_W2BEGb[5] ;
 wire \Tile_X10Y13_W2BEGb[6] ;
 wire \Tile_X10Y13_W2BEGb[7] ;
 wire \Tile_X10Y13_W6BEG[0] ;
 wire \Tile_X10Y13_W6BEG[10] ;
 wire \Tile_X10Y13_W6BEG[11] ;
 wire \Tile_X10Y13_W6BEG[1] ;
 wire \Tile_X10Y13_W6BEG[2] ;
 wire \Tile_X10Y13_W6BEG[3] ;
 wire \Tile_X10Y13_W6BEG[4] ;
 wire \Tile_X10Y13_W6BEG[5] ;
 wire \Tile_X10Y13_W6BEG[6] ;
 wire \Tile_X10Y13_W6BEG[7] ;
 wire \Tile_X10Y13_W6BEG[8] ;
 wire \Tile_X10Y13_W6BEG[9] ;
 wire \Tile_X10Y13_WW4BEG[0] ;
 wire \Tile_X10Y13_WW4BEG[10] ;
 wire \Tile_X10Y13_WW4BEG[11] ;
 wire \Tile_X10Y13_WW4BEG[12] ;
 wire \Tile_X10Y13_WW4BEG[13] ;
 wire \Tile_X10Y13_WW4BEG[14] ;
 wire \Tile_X10Y13_WW4BEG[15] ;
 wire \Tile_X10Y13_WW4BEG[1] ;
 wire \Tile_X10Y13_WW4BEG[2] ;
 wire \Tile_X10Y13_WW4BEG[3] ;
 wire \Tile_X10Y13_WW4BEG[4] ;
 wire \Tile_X10Y13_WW4BEG[5] ;
 wire \Tile_X10Y13_WW4BEG[6] ;
 wire \Tile_X10Y13_WW4BEG[7] ;
 wire \Tile_X10Y13_WW4BEG[8] ;
 wire \Tile_X10Y13_WW4BEG[9] ;
 wire \Tile_X10Y14_FrameData_O[0] ;
 wire \Tile_X10Y14_FrameData_O[10] ;
 wire \Tile_X10Y14_FrameData_O[11] ;
 wire \Tile_X10Y14_FrameData_O[12] ;
 wire \Tile_X10Y14_FrameData_O[13] ;
 wire \Tile_X10Y14_FrameData_O[14] ;
 wire \Tile_X10Y14_FrameData_O[15] ;
 wire \Tile_X10Y14_FrameData_O[16] ;
 wire \Tile_X10Y14_FrameData_O[17] ;
 wire \Tile_X10Y14_FrameData_O[18] ;
 wire \Tile_X10Y14_FrameData_O[19] ;
 wire \Tile_X10Y14_FrameData_O[1] ;
 wire \Tile_X10Y14_FrameData_O[20] ;
 wire \Tile_X10Y14_FrameData_O[21] ;
 wire \Tile_X10Y14_FrameData_O[22] ;
 wire \Tile_X10Y14_FrameData_O[23] ;
 wire \Tile_X10Y14_FrameData_O[24] ;
 wire \Tile_X10Y14_FrameData_O[25] ;
 wire \Tile_X10Y14_FrameData_O[26] ;
 wire \Tile_X10Y14_FrameData_O[27] ;
 wire \Tile_X10Y14_FrameData_O[28] ;
 wire \Tile_X10Y14_FrameData_O[29] ;
 wire \Tile_X10Y14_FrameData_O[2] ;
 wire \Tile_X10Y14_FrameData_O[30] ;
 wire \Tile_X10Y14_FrameData_O[31] ;
 wire \Tile_X10Y14_FrameData_O[3] ;
 wire \Tile_X10Y14_FrameData_O[4] ;
 wire \Tile_X10Y14_FrameData_O[5] ;
 wire \Tile_X10Y14_FrameData_O[6] ;
 wire \Tile_X10Y14_FrameData_O[7] ;
 wire \Tile_X10Y14_FrameData_O[8] ;
 wire \Tile_X10Y14_FrameData_O[9] ;
 wire \Tile_X10Y14_S1BEG[0] ;
 wire \Tile_X10Y14_S1BEG[1] ;
 wire \Tile_X10Y14_S1BEG[2] ;
 wire \Tile_X10Y14_S1BEG[3] ;
 wire \Tile_X10Y14_S2BEG[0] ;
 wire \Tile_X10Y14_S2BEG[1] ;
 wire \Tile_X10Y14_S2BEG[2] ;
 wire \Tile_X10Y14_S2BEG[3] ;
 wire \Tile_X10Y14_S2BEG[4] ;
 wire \Tile_X10Y14_S2BEG[5] ;
 wire \Tile_X10Y14_S2BEG[6] ;
 wire \Tile_X10Y14_S2BEG[7] ;
 wire \Tile_X10Y14_S2BEGb[0] ;
 wire \Tile_X10Y14_S2BEGb[1] ;
 wire \Tile_X10Y14_S2BEGb[2] ;
 wire \Tile_X10Y14_S2BEGb[3] ;
 wire \Tile_X10Y14_S2BEGb[4] ;
 wire \Tile_X10Y14_S2BEGb[5] ;
 wire \Tile_X10Y14_S2BEGb[6] ;
 wire \Tile_X10Y14_S2BEGb[7] ;
 wire \Tile_X10Y14_S4BEG[0] ;
 wire \Tile_X10Y14_S4BEG[10] ;
 wire \Tile_X10Y14_S4BEG[11] ;
 wire \Tile_X10Y14_S4BEG[12] ;
 wire \Tile_X10Y14_S4BEG[13] ;
 wire \Tile_X10Y14_S4BEG[14] ;
 wire \Tile_X10Y14_S4BEG[15] ;
 wire \Tile_X10Y14_S4BEG[1] ;
 wire \Tile_X10Y14_S4BEG[2] ;
 wire \Tile_X10Y14_S4BEG[3] ;
 wire \Tile_X10Y14_S4BEG[4] ;
 wire \Tile_X10Y14_S4BEG[5] ;
 wire \Tile_X10Y14_S4BEG[6] ;
 wire \Tile_X10Y14_S4BEG[7] ;
 wire \Tile_X10Y14_S4BEG[8] ;
 wire \Tile_X10Y14_S4BEG[9] ;
 wire \Tile_X10Y14_W1BEG[0] ;
 wire \Tile_X10Y14_W1BEG[1] ;
 wire \Tile_X10Y14_W1BEG[2] ;
 wire \Tile_X10Y14_W1BEG[3] ;
 wire \Tile_X10Y14_W2BEG[0] ;
 wire \Tile_X10Y14_W2BEG[1] ;
 wire \Tile_X10Y14_W2BEG[2] ;
 wire \Tile_X10Y14_W2BEG[3] ;
 wire \Tile_X10Y14_W2BEG[4] ;
 wire \Tile_X10Y14_W2BEG[5] ;
 wire \Tile_X10Y14_W2BEG[6] ;
 wire \Tile_X10Y14_W2BEG[7] ;
 wire \Tile_X10Y14_W2BEGb[0] ;
 wire \Tile_X10Y14_W2BEGb[1] ;
 wire \Tile_X10Y14_W2BEGb[2] ;
 wire \Tile_X10Y14_W2BEGb[3] ;
 wire \Tile_X10Y14_W2BEGb[4] ;
 wire \Tile_X10Y14_W2BEGb[5] ;
 wire \Tile_X10Y14_W2BEGb[6] ;
 wire \Tile_X10Y14_W2BEGb[7] ;
 wire \Tile_X10Y14_W6BEG[0] ;
 wire \Tile_X10Y14_W6BEG[10] ;
 wire \Tile_X10Y14_W6BEG[11] ;
 wire \Tile_X10Y14_W6BEG[1] ;
 wire \Tile_X10Y14_W6BEG[2] ;
 wire \Tile_X10Y14_W6BEG[3] ;
 wire \Tile_X10Y14_W6BEG[4] ;
 wire \Tile_X10Y14_W6BEG[5] ;
 wire \Tile_X10Y14_W6BEG[6] ;
 wire \Tile_X10Y14_W6BEG[7] ;
 wire \Tile_X10Y14_W6BEG[8] ;
 wire \Tile_X10Y14_W6BEG[9] ;
 wire \Tile_X10Y14_WW4BEG[0] ;
 wire \Tile_X10Y14_WW4BEG[10] ;
 wire \Tile_X10Y14_WW4BEG[11] ;
 wire \Tile_X10Y14_WW4BEG[12] ;
 wire \Tile_X10Y14_WW4BEG[13] ;
 wire \Tile_X10Y14_WW4BEG[14] ;
 wire \Tile_X10Y14_WW4BEG[15] ;
 wire \Tile_X10Y14_WW4BEG[1] ;
 wire \Tile_X10Y14_WW4BEG[2] ;
 wire \Tile_X10Y14_WW4BEG[3] ;
 wire \Tile_X10Y14_WW4BEG[4] ;
 wire \Tile_X10Y14_WW4BEG[5] ;
 wire \Tile_X10Y14_WW4BEG[6] ;
 wire \Tile_X10Y14_WW4BEG[7] ;
 wire \Tile_X10Y14_WW4BEG[8] ;
 wire \Tile_X10Y14_WW4BEG[9] ;
 wire \Tile_X10Y15_FrameData_O[0] ;
 wire \Tile_X10Y15_FrameData_O[10] ;
 wire \Tile_X10Y15_FrameData_O[11] ;
 wire \Tile_X10Y15_FrameData_O[12] ;
 wire \Tile_X10Y15_FrameData_O[13] ;
 wire \Tile_X10Y15_FrameData_O[14] ;
 wire \Tile_X10Y15_FrameData_O[15] ;
 wire \Tile_X10Y15_FrameData_O[16] ;
 wire \Tile_X10Y15_FrameData_O[17] ;
 wire \Tile_X10Y15_FrameData_O[18] ;
 wire \Tile_X10Y15_FrameData_O[19] ;
 wire \Tile_X10Y15_FrameData_O[1] ;
 wire \Tile_X10Y15_FrameData_O[20] ;
 wire \Tile_X10Y15_FrameData_O[21] ;
 wire \Tile_X10Y15_FrameData_O[22] ;
 wire \Tile_X10Y15_FrameData_O[23] ;
 wire \Tile_X10Y15_FrameData_O[24] ;
 wire \Tile_X10Y15_FrameData_O[25] ;
 wire \Tile_X10Y15_FrameData_O[26] ;
 wire \Tile_X10Y15_FrameData_O[27] ;
 wire \Tile_X10Y15_FrameData_O[28] ;
 wire \Tile_X10Y15_FrameData_O[29] ;
 wire \Tile_X10Y15_FrameData_O[2] ;
 wire \Tile_X10Y15_FrameData_O[30] ;
 wire \Tile_X10Y15_FrameData_O[31] ;
 wire \Tile_X10Y15_FrameData_O[3] ;
 wire \Tile_X10Y15_FrameData_O[4] ;
 wire \Tile_X10Y15_FrameData_O[5] ;
 wire \Tile_X10Y15_FrameData_O[6] ;
 wire \Tile_X10Y15_FrameData_O[7] ;
 wire \Tile_X10Y15_FrameData_O[8] ;
 wire \Tile_X10Y15_FrameData_O[9] ;
 wire \Tile_X10Y15_FrameStrobe_O[0] ;
 wire \Tile_X10Y15_FrameStrobe_O[10] ;
 wire \Tile_X10Y15_FrameStrobe_O[11] ;
 wire \Tile_X10Y15_FrameStrobe_O[12] ;
 wire \Tile_X10Y15_FrameStrobe_O[13] ;
 wire \Tile_X10Y15_FrameStrobe_O[14] ;
 wire \Tile_X10Y15_FrameStrobe_O[15] ;
 wire \Tile_X10Y15_FrameStrobe_O[16] ;
 wire \Tile_X10Y15_FrameStrobe_O[17] ;
 wire \Tile_X10Y15_FrameStrobe_O[18] ;
 wire \Tile_X10Y15_FrameStrobe_O[19] ;
 wire \Tile_X10Y15_FrameStrobe_O[1] ;
 wire \Tile_X10Y15_FrameStrobe_O[2] ;
 wire \Tile_X10Y15_FrameStrobe_O[3] ;
 wire \Tile_X10Y15_FrameStrobe_O[4] ;
 wire \Tile_X10Y15_FrameStrobe_O[5] ;
 wire \Tile_X10Y15_FrameStrobe_O[6] ;
 wire \Tile_X10Y15_FrameStrobe_O[7] ;
 wire \Tile_X10Y15_FrameStrobe_O[8] ;
 wire \Tile_X10Y15_FrameStrobe_O[9] ;
 wire \Tile_X10Y15_N1BEG[0] ;
 wire \Tile_X10Y15_N1BEG[1] ;
 wire \Tile_X10Y15_N1BEG[2] ;
 wire \Tile_X10Y15_N1BEG[3] ;
 wire \Tile_X10Y15_N2BEG[0] ;
 wire \Tile_X10Y15_N2BEG[1] ;
 wire \Tile_X10Y15_N2BEG[2] ;
 wire \Tile_X10Y15_N2BEG[3] ;
 wire \Tile_X10Y15_N2BEG[4] ;
 wire \Tile_X10Y15_N2BEG[5] ;
 wire \Tile_X10Y15_N2BEG[6] ;
 wire \Tile_X10Y15_N2BEG[7] ;
 wire \Tile_X10Y15_N2BEGb[0] ;
 wire \Tile_X10Y15_N2BEGb[1] ;
 wire \Tile_X10Y15_N2BEGb[2] ;
 wire \Tile_X10Y15_N2BEGb[3] ;
 wire \Tile_X10Y15_N2BEGb[4] ;
 wire \Tile_X10Y15_N2BEGb[5] ;
 wire \Tile_X10Y15_N2BEGb[6] ;
 wire \Tile_X10Y15_N2BEGb[7] ;
 wire \Tile_X10Y15_N4BEG[0] ;
 wire \Tile_X10Y15_N4BEG[10] ;
 wire \Tile_X10Y15_N4BEG[11] ;
 wire \Tile_X10Y15_N4BEG[12] ;
 wire \Tile_X10Y15_N4BEG[13] ;
 wire \Tile_X10Y15_N4BEG[14] ;
 wire \Tile_X10Y15_N4BEG[15] ;
 wire \Tile_X10Y15_N4BEG[1] ;
 wire \Tile_X10Y15_N4BEG[2] ;
 wire \Tile_X10Y15_N4BEG[3] ;
 wire \Tile_X10Y15_N4BEG[4] ;
 wire \Tile_X10Y15_N4BEG[5] ;
 wire \Tile_X10Y15_N4BEG[6] ;
 wire \Tile_X10Y15_N4BEG[7] ;
 wire \Tile_X10Y15_N4BEG[8] ;
 wire \Tile_X10Y15_N4BEG[9] ;
 wire Tile_X10Y15_UserCLKo;
 wire \Tile_X10Y1_FrameData_O[0] ;
 wire \Tile_X10Y1_FrameData_O[10] ;
 wire \Tile_X10Y1_FrameData_O[11] ;
 wire \Tile_X10Y1_FrameData_O[12] ;
 wire \Tile_X10Y1_FrameData_O[13] ;
 wire \Tile_X10Y1_FrameData_O[14] ;
 wire \Tile_X10Y1_FrameData_O[15] ;
 wire \Tile_X10Y1_FrameData_O[16] ;
 wire \Tile_X10Y1_FrameData_O[17] ;
 wire \Tile_X10Y1_FrameData_O[18] ;
 wire \Tile_X10Y1_FrameData_O[19] ;
 wire \Tile_X10Y1_FrameData_O[1] ;
 wire \Tile_X10Y1_FrameData_O[20] ;
 wire \Tile_X10Y1_FrameData_O[21] ;
 wire \Tile_X10Y1_FrameData_O[22] ;
 wire \Tile_X10Y1_FrameData_O[23] ;
 wire \Tile_X10Y1_FrameData_O[24] ;
 wire \Tile_X10Y1_FrameData_O[25] ;
 wire \Tile_X10Y1_FrameData_O[26] ;
 wire \Tile_X10Y1_FrameData_O[27] ;
 wire \Tile_X10Y1_FrameData_O[28] ;
 wire \Tile_X10Y1_FrameData_O[29] ;
 wire \Tile_X10Y1_FrameData_O[2] ;
 wire \Tile_X10Y1_FrameData_O[30] ;
 wire \Tile_X10Y1_FrameData_O[31] ;
 wire \Tile_X10Y1_FrameData_O[3] ;
 wire \Tile_X10Y1_FrameData_O[4] ;
 wire \Tile_X10Y1_FrameData_O[5] ;
 wire \Tile_X10Y1_FrameData_O[6] ;
 wire \Tile_X10Y1_FrameData_O[7] ;
 wire \Tile_X10Y1_FrameData_O[8] ;
 wire \Tile_X10Y1_FrameData_O[9] ;
 wire \Tile_X10Y1_FrameStrobe_O[0] ;
 wire \Tile_X10Y1_FrameStrobe_O[10] ;
 wire \Tile_X10Y1_FrameStrobe_O[11] ;
 wire \Tile_X10Y1_FrameStrobe_O[12] ;
 wire \Tile_X10Y1_FrameStrobe_O[13] ;
 wire \Tile_X10Y1_FrameStrobe_O[14] ;
 wire \Tile_X10Y1_FrameStrobe_O[15] ;
 wire \Tile_X10Y1_FrameStrobe_O[16] ;
 wire \Tile_X10Y1_FrameStrobe_O[17] ;
 wire \Tile_X10Y1_FrameStrobe_O[18] ;
 wire \Tile_X10Y1_FrameStrobe_O[19] ;
 wire \Tile_X10Y1_FrameStrobe_O[1] ;
 wire \Tile_X10Y1_FrameStrobe_O[2] ;
 wire \Tile_X10Y1_FrameStrobe_O[3] ;
 wire \Tile_X10Y1_FrameStrobe_O[4] ;
 wire \Tile_X10Y1_FrameStrobe_O[5] ;
 wire \Tile_X10Y1_FrameStrobe_O[6] ;
 wire \Tile_X10Y1_FrameStrobe_O[7] ;
 wire \Tile_X10Y1_FrameStrobe_O[8] ;
 wire \Tile_X10Y1_FrameStrobe_O[9] ;
 wire \Tile_X10Y1_N1BEG[0] ;
 wire \Tile_X10Y1_N1BEG[1] ;
 wire \Tile_X10Y1_N1BEG[2] ;
 wire \Tile_X10Y1_N1BEG[3] ;
 wire \Tile_X10Y1_N2BEG[0] ;
 wire \Tile_X10Y1_N2BEG[1] ;
 wire \Tile_X10Y1_N2BEG[2] ;
 wire \Tile_X10Y1_N2BEG[3] ;
 wire \Tile_X10Y1_N2BEG[4] ;
 wire \Tile_X10Y1_N2BEG[5] ;
 wire \Tile_X10Y1_N2BEG[6] ;
 wire \Tile_X10Y1_N2BEG[7] ;
 wire \Tile_X10Y1_N2BEGb[0] ;
 wire \Tile_X10Y1_N2BEGb[1] ;
 wire \Tile_X10Y1_N2BEGb[2] ;
 wire \Tile_X10Y1_N2BEGb[3] ;
 wire \Tile_X10Y1_N2BEGb[4] ;
 wire \Tile_X10Y1_N2BEGb[5] ;
 wire \Tile_X10Y1_N2BEGb[6] ;
 wire \Tile_X10Y1_N2BEGb[7] ;
 wire \Tile_X10Y1_N4BEG[0] ;
 wire \Tile_X10Y1_N4BEG[10] ;
 wire \Tile_X10Y1_N4BEG[11] ;
 wire \Tile_X10Y1_N4BEG[12] ;
 wire \Tile_X10Y1_N4BEG[13] ;
 wire \Tile_X10Y1_N4BEG[14] ;
 wire \Tile_X10Y1_N4BEG[15] ;
 wire \Tile_X10Y1_N4BEG[1] ;
 wire \Tile_X10Y1_N4BEG[2] ;
 wire \Tile_X10Y1_N4BEG[3] ;
 wire \Tile_X10Y1_N4BEG[4] ;
 wire \Tile_X10Y1_N4BEG[5] ;
 wire \Tile_X10Y1_N4BEG[6] ;
 wire \Tile_X10Y1_N4BEG[7] ;
 wire \Tile_X10Y1_N4BEG[8] ;
 wire \Tile_X10Y1_N4BEG[9] ;
 wire Tile_X10Y1_UserCLKo;
 wire \Tile_X10Y1_W1BEG[0] ;
 wire \Tile_X10Y1_W1BEG[1] ;
 wire \Tile_X10Y1_W1BEG[2] ;
 wire \Tile_X10Y1_W1BEG[3] ;
 wire \Tile_X10Y1_W2BEG[0] ;
 wire \Tile_X10Y1_W2BEG[1] ;
 wire \Tile_X10Y1_W2BEG[2] ;
 wire \Tile_X10Y1_W2BEG[3] ;
 wire \Tile_X10Y1_W2BEG[4] ;
 wire \Tile_X10Y1_W2BEG[5] ;
 wire \Tile_X10Y1_W2BEG[6] ;
 wire \Tile_X10Y1_W2BEG[7] ;
 wire \Tile_X10Y1_W2BEGb[0] ;
 wire \Tile_X10Y1_W2BEGb[1] ;
 wire \Tile_X10Y1_W2BEGb[2] ;
 wire \Tile_X10Y1_W2BEGb[3] ;
 wire \Tile_X10Y1_W2BEGb[4] ;
 wire \Tile_X10Y1_W2BEGb[5] ;
 wire \Tile_X10Y1_W2BEGb[6] ;
 wire \Tile_X10Y1_W2BEGb[7] ;
 wire \Tile_X10Y1_W6BEG[0] ;
 wire \Tile_X10Y1_W6BEG[10] ;
 wire \Tile_X10Y1_W6BEG[11] ;
 wire \Tile_X10Y1_W6BEG[1] ;
 wire \Tile_X10Y1_W6BEG[2] ;
 wire \Tile_X10Y1_W6BEG[3] ;
 wire \Tile_X10Y1_W6BEG[4] ;
 wire \Tile_X10Y1_W6BEG[5] ;
 wire \Tile_X10Y1_W6BEG[6] ;
 wire \Tile_X10Y1_W6BEG[7] ;
 wire \Tile_X10Y1_W6BEG[8] ;
 wire \Tile_X10Y1_W6BEG[9] ;
 wire \Tile_X10Y1_WW4BEG[0] ;
 wire \Tile_X10Y1_WW4BEG[10] ;
 wire \Tile_X10Y1_WW4BEG[11] ;
 wire \Tile_X10Y1_WW4BEG[12] ;
 wire \Tile_X10Y1_WW4BEG[13] ;
 wire \Tile_X10Y1_WW4BEG[14] ;
 wire \Tile_X10Y1_WW4BEG[15] ;
 wire \Tile_X10Y1_WW4BEG[1] ;
 wire \Tile_X10Y1_WW4BEG[2] ;
 wire \Tile_X10Y1_WW4BEG[3] ;
 wire \Tile_X10Y1_WW4BEG[4] ;
 wire \Tile_X10Y1_WW4BEG[5] ;
 wire \Tile_X10Y1_WW4BEG[6] ;
 wire \Tile_X10Y1_WW4BEG[7] ;
 wire \Tile_X10Y1_WW4BEG[8] ;
 wire \Tile_X10Y1_WW4BEG[9] ;
 wire \Tile_X10Y2_FrameData_O[0] ;
 wire \Tile_X10Y2_FrameData_O[10] ;
 wire \Tile_X10Y2_FrameData_O[11] ;
 wire \Tile_X10Y2_FrameData_O[12] ;
 wire \Tile_X10Y2_FrameData_O[13] ;
 wire \Tile_X10Y2_FrameData_O[14] ;
 wire \Tile_X10Y2_FrameData_O[15] ;
 wire \Tile_X10Y2_FrameData_O[16] ;
 wire \Tile_X10Y2_FrameData_O[17] ;
 wire \Tile_X10Y2_FrameData_O[18] ;
 wire \Tile_X10Y2_FrameData_O[19] ;
 wire \Tile_X10Y2_FrameData_O[1] ;
 wire \Tile_X10Y2_FrameData_O[20] ;
 wire \Tile_X10Y2_FrameData_O[21] ;
 wire \Tile_X10Y2_FrameData_O[22] ;
 wire \Tile_X10Y2_FrameData_O[23] ;
 wire \Tile_X10Y2_FrameData_O[24] ;
 wire \Tile_X10Y2_FrameData_O[25] ;
 wire \Tile_X10Y2_FrameData_O[26] ;
 wire \Tile_X10Y2_FrameData_O[27] ;
 wire \Tile_X10Y2_FrameData_O[28] ;
 wire \Tile_X10Y2_FrameData_O[29] ;
 wire \Tile_X10Y2_FrameData_O[2] ;
 wire \Tile_X10Y2_FrameData_O[30] ;
 wire \Tile_X10Y2_FrameData_O[31] ;
 wire \Tile_X10Y2_FrameData_O[3] ;
 wire \Tile_X10Y2_FrameData_O[4] ;
 wire \Tile_X10Y2_FrameData_O[5] ;
 wire \Tile_X10Y2_FrameData_O[6] ;
 wire \Tile_X10Y2_FrameData_O[7] ;
 wire \Tile_X10Y2_FrameData_O[8] ;
 wire \Tile_X10Y2_FrameData_O[9] ;
 wire \Tile_X10Y2_S1BEG[0] ;
 wire \Tile_X10Y2_S1BEG[1] ;
 wire \Tile_X10Y2_S1BEG[2] ;
 wire \Tile_X10Y2_S1BEG[3] ;
 wire \Tile_X10Y2_S2BEG[0] ;
 wire \Tile_X10Y2_S2BEG[1] ;
 wire \Tile_X10Y2_S2BEG[2] ;
 wire \Tile_X10Y2_S2BEG[3] ;
 wire \Tile_X10Y2_S2BEG[4] ;
 wire \Tile_X10Y2_S2BEG[5] ;
 wire \Tile_X10Y2_S2BEG[6] ;
 wire \Tile_X10Y2_S2BEG[7] ;
 wire \Tile_X10Y2_S2BEGb[0] ;
 wire \Tile_X10Y2_S2BEGb[1] ;
 wire \Tile_X10Y2_S2BEGb[2] ;
 wire \Tile_X10Y2_S2BEGb[3] ;
 wire \Tile_X10Y2_S2BEGb[4] ;
 wire \Tile_X10Y2_S2BEGb[5] ;
 wire \Tile_X10Y2_S2BEGb[6] ;
 wire \Tile_X10Y2_S2BEGb[7] ;
 wire \Tile_X10Y2_S4BEG[0] ;
 wire \Tile_X10Y2_S4BEG[10] ;
 wire \Tile_X10Y2_S4BEG[11] ;
 wire \Tile_X10Y2_S4BEG[12] ;
 wire \Tile_X10Y2_S4BEG[13] ;
 wire \Tile_X10Y2_S4BEG[14] ;
 wire \Tile_X10Y2_S4BEG[15] ;
 wire \Tile_X10Y2_S4BEG[1] ;
 wire \Tile_X10Y2_S4BEG[2] ;
 wire \Tile_X10Y2_S4BEG[3] ;
 wire \Tile_X10Y2_S4BEG[4] ;
 wire \Tile_X10Y2_S4BEG[5] ;
 wire \Tile_X10Y2_S4BEG[6] ;
 wire \Tile_X10Y2_S4BEG[7] ;
 wire \Tile_X10Y2_S4BEG[8] ;
 wire \Tile_X10Y2_S4BEG[9] ;
 wire \Tile_X10Y2_W1BEG[0] ;
 wire \Tile_X10Y2_W1BEG[1] ;
 wire \Tile_X10Y2_W1BEG[2] ;
 wire \Tile_X10Y2_W1BEG[3] ;
 wire \Tile_X10Y2_W2BEG[0] ;
 wire \Tile_X10Y2_W2BEG[1] ;
 wire \Tile_X10Y2_W2BEG[2] ;
 wire \Tile_X10Y2_W2BEG[3] ;
 wire \Tile_X10Y2_W2BEG[4] ;
 wire \Tile_X10Y2_W2BEG[5] ;
 wire \Tile_X10Y2_W2BEG[6] ;
 wire \Tile_X10Y2_W2BEG[7] ;
 wire \Tile_X10Y2_W2BEGb[0] ;
 wire \Tile_X10Y2_W2BEGb[1] ;
 wire \Tile_X10Y2_W2BEGb[2] ;
 wire \Tile_X10Y2_W2BEGb[3] ;
 wire \Tile_X10Y2_W2BEGb[4] ;
 wire \Tile_X10Y2_W2BEGb[5] ;
 wire \Tile_X10Y2_W2BEGb[6] ;
 wire \Tile_X10Y2_W2BEGb[7] ;
 wire \Tile_X10Y2_W6BEG[0] ;
 wire \Tile_X10Y2_W6BEG[10] ;
 wire \Tile_X10Y2_W6BEG[11] ;
 wire \Tile_X10Y2_W6BEG[1] ;
 wire \Tile_X10Y2_W6BEG[2] ;
 wire \Tile_X10Y2_W6BEG[3] ;
 wire \Tile_X10Y2_W6BEG[4] ;
 wire \Tile_X10Y2_W6BEG[5] ;
 wire \Tile_X10Y2_W6BEG[6] ;
 wire \Tile_X10Y2_W6BEG[7] ;
 wire \Tile_X10Y2_W6BEG[8] ;
 wire \Tile_X10Y2_W6BEG[9] ;
 wire \Tile_X10Y2_WW4BEG[0] ;
 wire \Tile_X10Y2_WW4BEG[10] ;
 wire \Tile_X10Y2_WW4BEG[11] ;
 wire \Tile_X10Y2_WW4BEG[12] ;
 wire \Tile_X10Y2_WW4BEG[13] ;
 wire \Tile_X10Y2_WW4BEG[14] ;
 wire \Tile_X10Y2_WW4BEG[15] ;
 wire \Tile_X10Y2_WW4BEG[1] ;
 wire \Tile_X10Y2_WW4BEG[2] ;
 wire \Tile_X10Y2_WW4BEG[3] ;
 wire \Tile_X10Y2_WW4BEG[4] ;
 wire \Tile_X10Y2_WW4BEG[5] ;
 wire \Tile_X10Y2_WW4BEG[6] ;
 wire \Tile_X10Y2_WW4BEG[7] ;
 wire \Tile_X10Y2_WW4BEG[8] ;
 wire \Tile_X10Y2_WW4BEG[9] ;
 wire \Tile_X10Y3_FrameData_O[0] ;
 wire \Tile_X10Y3_FrameData_O[10] ;
 wire \Tile_X10Y3_FrameData_O[11] ;
 wire \Tile_X10Y3_FrameData_O[12] ;
 wire \Tile_X10Y3_FrameData_O[13] ;
 wire \Tile_X10Y3_FrameData_O[14] ;
 wire \Tile_X10Y3_FrameData_O[15] ;
 wire \Tile_X10Y3_FrameData_O[16] ;
 wire \Tile_X10Y3_FrameData_O[17] ;
 wire \Tile_X10Y3_FrameData_O[18] ;
 wire \Tile_X10Y3_FrameData_O[19] ;
 wire \Tile_X10Y3_FrameData_O[1] ;
 wire \Tile_X10Y3_FrameData_O[20] ;
 wire \Tile_X10Y3_FrameData_O[21] ;
 wire \Tile_X10Y3_FrameData_O[22] ;
 wire \Tile_X10Y3_FrameData_O[23] ;
 wire \Tile_X10Y3_FrameData_O[24] ;
 wire \Tile_X10Y3_FrameData_O[25] ;
 wire \Tile_X10Y3_FrameData_O[26] ;
 wire \Tile_X10Y3_FrameData_O[27] ;
 wire \Tile_X10Y3_FrameData_O[28] ;
 wire \Tile_X10Y3_FrameData_O[29] ;
 wire \Tile_X10Y3_FrameData_O[2] ;
 wire \Tile_X10Y3_FrameData_O[30] ;
 wire \Tile_X10Y3_FrameData_O[31] ;
 wire \Tile_X10Y3_FrameData_O[3] ;
 wire \Tile_X10Y3_FrameData_O[4] ;
 wire \Tile_X10Y3_FrameData_O[5] ;
 wire \Tile_X10Y3_FrameData_O[6] ;
 wire \Tile_X10Y3_FrameData_O[7] ;
 wire \Tile_X10Y3_FrameData_O[8] ;
 wire \Tile_X10Y3_FrameData_O[9] ;
 wire \Tile_X10Y3_FrameStrobe_O[0] ;
 wire \Tile_X10Y3_FrameStrobe_O[10] ;
 wire \Tile_X10Y3_FrameStrobe_O[11] ;
 wire \Tile_X10Y3_FrameStrobe_O[12] ;
 wire \Tile_X10Y3_FrameStrobe_O[13] ;
 wire \Tile_X10Y3_FrameStrobe_O[14] ;
 wire \Tile_X10Y3_FrameStrobe_O[15] ;
 wire \Tile_X10Y3_FrameStrobe_O[16] ;
 wire \Tile_X10Y3_FrameStrobe_O[17] ;
 wire \Tile_X10Y3_FrameStrobe_O[18] ;
 wire \Tile_X10Y3_FrameStrobe_O[19] ;
 wire \Tile_X10Y3_FrameStrobe_O[1] ;
 wire \Tile_X10Y3_FrameStrobe_O[2] ;
 wire \Tile_X10Y3_FrameStrobe_O[3] ;
 wire \Tile_X10Y3_FrameStrobe_O[4] ;
 wire \Tile_X10Y3_FrameStrobe_O[5] ;
 wire \Tile_X10Y3_FrameStrobe_O[6] ;
 wire \Tile_X10Y3_FrameStrobe_O[7] ;
 wire \Tile_X10Y3_FrameStrobe_O[8] ;
 wire \Tile_X10Y3_FrameStrobe_O[9] ;
 wire \Tile_X10Y3_N1BEG[0] ;
 wire \Tile_X10Y3_N1BEG[1] ;
 wire \Tile_X10Y3_N1BEG[2] ;
 wire \Tile_X10Y3_N1BEG[3] ;
 wire \Tile_X10Y3_N2BEG[0] ;
 wire \Tile_X10Y3_N2BEG[1] ;
 wire \Tile_X10Y3_N2BEG[2] ;
 wire \Tile_X10Y3_N2BEG[3] ;
 wire \Tile_X10Y3_N2BEG[4] ;
 wire \Tile_X10Y3_N2BEG[5] ;
 wire \Tile_X10Y3_N2BEG[6] ;
 wire \Tile_X10Y3_N2BEG[7] ;
 wire \Tile_X10Y3_N2BEGb[0] ;
 wire \Tile_X10Y3_N2BEGb[1] ;
 wire \Tile_X10Y3_N2BEGb[2] ;
 wire \Tile_X10Y3_N2BEGb[3] ;
 wire \Tile_X10Y3_N2BEGb[4] ;
 wire \Tile_X10Y3_N2BEGb[5] ;
 wire \Tile_X10Y3_N2BEGb[6] ;
 wire \Tile_X10Y3_N2BEGb[7] ;
 wire \Tile_X10Y3_N4BEG[0] ;
 wire \Tile_X10Y3_N4BEG[10] ;
 wire \Tile_X10Y3_N4BEG[11] ;
 wire \Tile_X10Y3_N4BEG[12] ;
 wire \Tile_X10Y3_N4BEG[13] ;
 wire \Tile_X10Y3_N4BEG[14] ;
 wire \Tile_X10Y3_N4BEG[15] ;
 wire \Tile_X10Y3_N4BEG[1] ;
 wire \Tile_X10Y3_N4BEG[2] ;
 wire \Tile_X10Y3_N4BEG[3] ;
 wire \Tile_X10Y3_N4BEG[4] ;
 wire \Tile_X10Y3_N4BEG[5] ;
 wire \Tile_X10Y3_N4BEG[6] ;
 wire \Tile_X10Y3_N4BEG[7] ;
 wire \Tile_X10Y3_N4BEG[8] ;
 wire \Tile_X10Y3_N4BEG[9] ;
 wire Tile_X10Y3_UserCLKo;
 wire \Tile_X10Y3_W1BEG[0] ;
 wire \Tile_X10Y3_W1BEG[1] ;
 wire \Tile_X10Y3_W1BEG[2] ;
 wire \Tile_X10Y3_W1BEG[3] ;
 wire \Tile_X10Y3_W2BEG[0] ;
 wire \Tile_X10Y3_W2BEG[1] ;
 wire \Tile_X10Y3_W2BEG[2] ;
 wire \Tile_X10Y3_W2BEG[3] ;
 wire \Tile_X10Y3_W2BEG[4] ;
 wire \Tile_X10Y3_W2BEG[5] ;
 wire \Tile_X10Y3_W2BEG[6] ;
 wire \Tile_X10Y3_W2BEG[7] ;
 wire \Tile_X10Y3_W2BEGb[0] ;
 wire \Tile_X10Y3_W2BEGb[1] ;
 wire \Tile_X10Y3_W2BEGb[2] ;
 wire \Tile_X10Y3_W2BEGb[3] ;
 wire \Tile_X10Y3_W2BEGb[4] ;
 wire \Tile_X10Y3_W2BEGb[5] ;
 wire \Tile_X10Y3_W2BEGb[6] ;
 wire \Tile_X10Y3_W2BEGb[7] ;
 wire \Tile_X10Y3_W6BEG[0] ;
 wire \Tile_X10Y3_W6BEG[10] ;
 wire \Tile_X10Y3_W6BEG[11] ;
 wire \Tile_X10Y3_W6BEG[1] ;
 wire \Tile_X10Y3_W6BEG[2] ;
 wire \Tile_X10Y3_W6BEG[3] ;
 wire \Tile_X10Y3_W6BEG[4] ;
 wire \Tile_X10Y3_W6BEG[5] ;
 wire \Tile_X10Y3_W6BEG[6] ;
 wire \Tile_X10Y3_W6BEG[7] ;
 wire \Tile_X10Y3_W6BEG[8] ;
 wire \Tile_X10Y3_W6BEG[9] ;
 wire \Tile_X10Y3_WW4BEG[0] ;
 wire \Tile_X10Y3_WW4BEG[10] ;
 wire \Tile_X10Y3_WW4BEG[11] ;
 wire \Tile_X10Y3_WW4BEG[12] ;
 wire \Tile_X10Y3_WW4BEG[13] ;
 wire \Tile_X10Y3_WW4BEG[14] ;
 wire \Tile_X10Y3_WW4BEG[15] ;
 wire \Tile_X10Y3_WW4BEG[1] ;
 wire \Tile_X10Y3_WW4BEG[2] ;
 wire \Tile_X10Y3_WW4BEG[3] ;
 wire \Tile_X10Y3_WW4BEG[4] ;
 wire \Tile_X10Y3_WW4BEG[5] ;
 wire \Tile_X10Y3_WW4BEG[6] ;
 wire \Tile_X10Y3_WW4BEG[7] ;
 wire \Tile_X10Y3_WW4BEG[8] ;
 wire \Tile_X10Y3_WW4BEG[9] ;
 wire \Tile_X10Y4_FrameData_O[0] ;
 wire \Tile_X10Y4_FrameData_O[10] ;
 wire \Tile_X10Y4_FrameData_O[11] ;
 wire \Tile_X10Y4_FrameData_O[12] ;
 wire \Tile_X10Y4_FrameData_O[13] ;
 wire \Tile_X10Y4_FrameData_O[14] ;
 wire \Tile_X10Y4_FrameData_O[15] ;
 wire \Tile_X10Y4_FrameData_O[16] ;
 wire \Tile_X10Y4_FrameData_O[17] ;
 wire \Tile_X10Y4_FrameData_O[18] ;
 wire \Tile_X10Y4_FrameData_O[19] ;
 wire \Tile_X10Y4_FrameData_O[1] ;
 wire \Tile_X10Y4_FrameData_O[20] ;
 wire \Tile_X10Y4_FrameData_O[21] ;
 wire \Tile_X10Y4_FrameData_O[22] ;
 wire \Tile_X10Y4_FrameData_O[23] ;
 wire \Tile_X10Y4_FrameData_O[24] ;
 wire \Tile_X10Y4_FrameData_O[25] ;
 wire \Tile_X10Y4_FrameData_O[26] ;
 wire \Tile_X10Y4_FrameData_O[27] ;
 wire \Tile_X10Y4_FrameData_O[28] ;
 wire \Tile_X10Y4_FrameData_O[29] ;
 wire \Tile_X10Y4_FrameData_O[2] ;
 wire \Tile_X10Y4_FrameData_O[30] ;
 wire \Tile_X10Y4_FrameData_O[31] ;
 wire \Tile_X10Y4_FrameData_O[3] ;
 wire \Tile_X10Y4_FrameData_O[4] ;
 wire \Tile_X10Y4_FrameData_O[5] ;
 wire \Tile_X10Y4_FrameData_O[6] ;
 wire \Tile_X10Y4_FrameData_O[7] ;
 wire \Tile_X10Y4_FrameData_O[8] ;
 wire \Tile_X10Y4_FrameData_O[9] ;
 wire \Tile_X10Y4_S1BEG[0] ;
 wire \Tile_X10Y4_S1BEG[1] ;
 wire \Tile_X10Y4_S1BEG[2] ;
 wire \Tile_X10Y4_S1BEG[3] ;
 wire \Tile_X10Y4_S2BEG[0] ;
 wire \Tile_X10Y4_S2BEG[1] ;
 wire \Tile_X10Y4_S2BEG[2] ;
 wire \Tile_X10Y4_S2BEG[3] ;
 wire \Tile_X10Y4_S2BEG[4] ;
 wire \Tile_X10Y4_S2BEG[5] ;
 wire \Tile_X10Y4_S2BEG[6] ;
 wire \Tile_X10Y4_S2BEG[7] ;
 wire \Tile_X10Y4_S2BEGb[0] ;
 wire \Tile_X10Y4_S2BEGb[1] ;
 wire \Tile_X10Y4_S2BEGb[2] ;
 wire \Tile_X10Y4_S2BEGb[3] ;
 wire \Tile_X10Y4_S2BEGb[4] ;
 wire \Tile_X10Y4_S2BEGb[5] ;
 wire \Tile_X10Y4_S2BEGb[6] ;
 wire \Tile_X10Y4_S2BEGb[7] ;
 wire \Tile_X10Y4_S4BEG[0] ;
 wire \Tile_X10Y4_S4BEG[10] ;
 wire \Tile_X10Y4_S4BEG[11] ;
 wire \Tile_X10Y4_S4BEG[12] ;
 wire \Tile_X10Y4_S4BEG[13] ;
 wire \Tile_X10Y4_S4BEG[14] ;
 wire \Tile_X10Y4_S4BEG[15] ;
 wire \Tile_X10Y4_S4BEG[1] ;
 wire \Tile_X10Y4_S4BEG[2] ;
 wire \Tile_X10Y4_S4BEG[3] ;
 wire \Tile_X10Y4_S4BEG[4] ;
 wire \Tile_X10Y4_S4BEG[5] ;
 wire \Tile_X10Y4_S4BEG[6] ;
 wire \Tile_X10Y4_S4BEG[7] ;
 wire \Tile_X10Y4_S4BEG[8] ;
 wire \Tile_X10Y4_S4BEG[9] ;
 wire \Tile_X10Y4_W1BEG[0] ;
 wire \Tile_X10Y4_W1BEG[1] ;
 wire \Tile_X10Y4_W1BEG[2] ;
 wire \Tile_X10Y4_W1BEG[3] ;
 wire \Tile_X10Y4_W2BEG[0] ;
 wire \Tile_X10Y4_W2BEG[1] ;
 wire \Tile_X10Y4_W2BEG[2] ;
 wire \Tile_X10Y4_W2BEG[3] ;
 wire \Tile_X10Y4_W2BEG[4] ;
 wire \Tile_X10Y4_W2BEG[5] ;
 wire \Tile_X10Y4_W2BEG[6] ;
 wire \Tile_X10Y4_W2BEG[7] ;
 wire \Tile_X10Y4_W2BEGb[0] ;
 wire \Tile_X10Y4_W2BEGb[1] ;
 wire \Tile_X10Y4_W2BEGb[2] ;
 wire \Tile_X10Y4_W2BEGb[3] ;
 wire \Tile_X10Y4_W2BEGb[4] ;
 wire \Tile_X10Y4_W2BEGb[5] ;
 wire \Tile_X10Y4_W2BEGb[6] ;
 wire \Tile_X10Y4_W2BEGb[7] ;
 wire \Tile_X10Y4_W6BEG[0] ;
 wire \Tile_X10Y4_W6BEG[10] ;
 wire \Tile_X10Y4_W6BEG[11] ;
 wire \Tile_X10Y4_W6BEG[1] ;
 wire \Tile_X10Y4_W6BEG[2] ;
 wire \Tile_X10Y4_W6BEG[3] ;
 wire \Tile_X10Y4_W6BEG[4] ;
 wire \Tile_X10Y4_W6BEG[5] ;
 wire \Tile_X10Y4_W6BEG[6] ;
 wire \Tile_X10Y4_W6BEG[7] ;
 wire \Tile_X10Y4_W6BEG[8] ;
 wire \Tile_X10Y4_W6BEG[9] ;
 wire \Tile_X10Y4_WW4BEG[0] ;
 wire \Tile_X10Y4_WW4BEG[10] ;
 wire \Tile_X10Y4_WW4BEG[11] ;
 wire \Tile_X10Y4_WW4BEG[12] ;
 wire \Tile_X10Y4_WW4BEG[13] ;
 wire \Tile_X10Y4_WW4BEG[14] ;
 wire \Tile_X10Y4_WW4BEG[15] ;
 wire \Tile_X10Y4_WW4BEG[1] ;
 wire \Tile_X10Y4_WW4BEG[2] ;
 wire \Tile_X10Y4_WW4BEG[3] ;
 wire \Tile_X10Y4_WW4BEG[4] ;
 wire \Tile_X10Y4_WW4BEG[5] ;
 wire \Tile_X10Y4_WW4BEG[6] ;
 wire \Tile_X10Y4_WW4BEG[7] ;
 wire \Tile_X10Y4_WW4BEG[8] ;
 wire \Tile_X10Y4_WW4BEG[9] ;
 wire \Tile_X10Y5_FrameData_O[0] ;
 wire \Tile_X10Y5_FrameData_O[10] ;
 wire \Tile_X10Y5_FrameData_O[11] ;
 wire \Tile_X10Y5_FrameData_O[12] ;
 wire \Tile_X10Y5_FrameData_O[13] ;
 wire \Tile_X10Y5_FrameData_O[14] ;
 wire \Tile_X10Y5_FrameData_O[15] ;
 wire \Tile_X10Y5_FrameData_O[16] ;
 wire \Tile_X10Y5_FrameData_O[17] ;
 wire \Tile_X10Y5_FrameData_O[18] ;
 wire \Tile_X10Y5_FrameData_O[19] ;
 wire \Tile_X10Y5_FrameData_O[1] ;
 wire \Tile_X10Y5_FrameData_O[20] ;
 wire \Tile_X10Y5_FrameData_O[21] ;
 wire \Tile_X10Y5_FrameData_O[22] ;
 wire \Tile_X10Y5_FrameData_O[23] ;
 wire \Tile_X10Y5_FrameData_O[24] ;
 wire \Tile_X10Y5_FrameData_O[25] ;
 wire \Tile_X10Y5_FrameData_O[26] ;
 wire \Tile_X10Y5_FrameData_O[27] ;
 wire \Tile_X10Y5_FrameData_O[28] ;
 wire \Tile_X10Y5_FrameData_O[29] ;
 wire \Tile_X10Y5_FrameData_O[2] ;
 wire \Tile_X10Y5_FrameData_O[30] ;
 wire \Tile_X10Y5_FrameData_O[31] ;
 wire \Tile_X10Y5_FrameData_O[3] ;
 wire \Tile_X10Y5_FrameData_O[4] ;
 wire \Tile_X10Y5_FrameData_O[5] ;
 wire \Tile_X10Y5_FrameData_O[6] ;
 wire \Tile_X10Y5_FrameData_O[7] ;
 wire \Tile_X10Y5_FrameData_O[8] ;
 wire \Tile_X10Y5_FrameData_O[9] ;
 wire \Tile_X10Y5_FrameStrobe_O[0] ;
 wire \Tile_X10Y5_FrameStrobe_O[10] ;
 wire \Tile_X10Y5_FrameStrobe_O[11] ;
 wire \Tile_X10Y5_FrameStrobe_O[12] ;
 wire \Tile_X10Y5_FrameStrobe_O[13] ;
 wire \Tile_X10Y5_FrameStrobe_O[14] ;
 wire \Tile_X10Y5_FrameStrobe_O[15] ;
 wire \Tile_X10Y5_FrameStrobe_O[16] ;
 wire \Tile_X10Y5_FrameStrobe_O[17] ;
 wire \Tile_X10Y5_FrameStrobe_O[18] ;
 wire \Tile_X10Y5_FrameStrobe_O[19] ;
 wire \Tile_X10Y5_FrameStrobe_O[1] ;
 wire \Tile_X10Y5_FrameStrobe_O[2] ;
 wire \Tile_X10Y5_FrameStrobe_O[3] ;
 wire \Tile_X10Y5_FrameStrobe_O[4] ;
 wire \Tile_X10Y5_FrameStrobe_O[5] ;
 wire \Tile_X10Y5_FrameStrobe_O[6] ;
 wire \Tile_X10Y5_FrameStrobe_O[7] ;
 wire \Tile_X10Y5_FrameStrobe_O[8] ;
 wire \Tile_X10Y5_FrameStrobe_O[9] ;
 wire \Tile_X10Y5_N1BEG[0] ;
 wire \Tile_X10Y5_N1BEG[1] ;
 wire \Tile_X10Y5_N1BEG[2] ;
 wire \Tile_X10Y5_N1BEG[3] ;
 wire \Tile_X10Y5_N2BEG[0] ;
 wire \Tile_X10Y5_N2BEG[1] ;
 wire \Tile_X10Y5_N2BEG[2] ;
 wire \Tile_X10Y5_N2BEG[3] ;
 wire \Tile_X10Y5_N2BEG[4] ;
 wire \Tile_X10Y5_N2BEG[5] ;
 wire \Tile_X10Y5_N2BEG[6] ;
 wire \Tile_X10Y5_N2BEG[7] ;
 wire \Tile_X10Y5_N2BEGb[0] ;
 wire \Tile_X10Y5_N2BEGb[1] ;
 wire \Tile_X10Y5_N2BEGb[2] ;
 wire \Tile_X10Y5_N2BEGb[3] ;
 wire \Tile_X10Y5_N2BEGb[4] ;
 wire \Tile_X10Y5_N2BEGb[5] ;
 wire \Tile_X10Y5_N2BEGb[6] ;
 wire \Tile_X10Y5_N2BEGb[7] ;
 wire \Tile_X10Y5_N4BEG[0] ;
 wire \Tile_X10Y5_N4BEG[10] ;
 wire \Tile_X10Y5_N4BEG[11] ;
 wire \Tile_X10Y5_N4BEG[12] ;
 wire \Tile_X10Y5_N4BEG[13] ;
 wire \Tile_X10Y5_N4BEG[14] ;
 wire \Tile_X10Y5_N4BEG[15] ;
 wire \Tile_X10Y5_N4BEG[1] ;
 wire \Tile_X10Y5_N4BEG[2] ;
 wire \Tile_X10Y5_N4BEG[3] ;
 wire \Tile_X10Y5_N4BEG[4] ;
 wire \Tile_X10Y5_N4BEG[5] ;
 wire \Tile_X10Y5_N4BEG[6] ;
 wire \Tile_X10Y5_N4BEG[7] ;
 wire \Tile_X10Y5_N4BEG[8] ;
 wire \Tile_X10Y5_N4BEG[9] ;
 wire Tile_X10Y5_UserCLKo;
 wire \Tile_X10Y5_W1BEG[0] ;
 wire \Tile_X10Y5_W1BEG[1] ;
 wire \Tile_X10Y5_W1BEG[2] ;
 wire \Tile_X10Y5_W1BEG[3] ;
 wire \Tile_X10Y5_W2BEG[0] ;
 wire \Tile_X10Y5_W2BEG[1] ;
 wire \Tile_X10Y5_W2BEG[2] ;
 wire \Tile_X10Y5_W2BEG[3] ;
 wire \Tile_X10Y5_W2BEG[4] ;
 wire \Tile_X10Y5_W2BEG[5] ;
 wire \Tile_X10Y5_W2BEG[6] ;
 wire \Tile_X10Y5_W2BEG[7] ;
 wire \Tile_X10Y5_W2BEGb[0] ;
 wire \Tile_X10Y5_W2BEGb[1] ;
 wire \Tile_X10Y5_W2BEGb[2] ;
 wire \Tile_X10Y5_W2BEGb[3] ;
 wire \Tile_X10Y5_W2BEGb[4] ;
 wire \Tile_X10Y5_W2BEGb[5] ;
 wire \Tile_X10Y5_W2BEGb[6] ;
 wire \Tile_X10Y5_W2BEGb[7] ;
 wire \Tile_X10Y5_W6BEG[0] ;
 wire \Tile_X10Y5_W6BEG[10] ;
 wire \Tile_X10Y5_W6BEG[11] ;
 wire \Tile_X10Y5_W6BEG[1] ;
 wire \Tile_X10Y5_W6BEG[2] ;
 wire \Tile_X10Y5_W6BEG[3] ;
 wire \Tile_X10Y5_W6BEG[4] ;
 wire \Tile_X10Y5_W6BEG[5] ;
 wire \Tile_X10Y5_W6BEG[6] ;
 wire \Tile_X10Y5_W6BEG[7] ;
 wire \Tile_X10Y5_W6BEG[8] ;
 wire \Tile_X10Y5_W6BEG[9] ;
 wire \Tile_X10Y5_WW4BEG[0] ;
 wire \Tile_X10Y5_WW4BEG[10] ;
 wire \Tile_X10Y5_WW4BEG[11] ;
 wire \Tile_X10Y5_WW4BEG[12] ;
 wire \Tile_X10Y5_WW4BEG[13] ;
 wire \Tile_X10Y5_WW4BEG[14] ;
 wire \Tile_X10Y5_WW4BEG[15] ;
 wire \Tile_X10Y5_WW4BEG[1] ;
 wire \Tile_X10Y5_WW4BEG[2] ;
 wire \Tile_X10Y5_WW4BEG[3] ;
 wire \Tile_X10Y5_WW4BEG[4] ;
 wire \Tile_X10Y5_WW4BEG[5] ;
 wire \Tile_X10Y5_WW4BEG[6] ;
 wire \Tile_X10Y5_WW4BEG[7] ;
 wire \Tile_X10Y5_WW4BEG[8] ;
 wire \Tile_X10Y5_WW4BEG[9] ;
 wire \Tile_X10Y6_FrameData_O[0] ;
 wire \Tile_X10Y6_FrameData_O[10] ;
 wire \Tile_X10Y6_FrameData_O[11] ;
 wire \Tile_X10Y6_FrameData_O[12] ;
 wire \Tile_X10Y6_FrameData_O[13] ;
 wire \Tile_X10Y6_FrameData_O[14] ;
 wire \Tile_X10Y6_FrameData_O[15] ;
 wire \Tile_X10Y6_FrameData_O[16] ;
 wire \Tile_X10Y6_FrameData_O[17] ;
 wire \Tile_X10Y6_FrameData_O[18] ;
 wire \Tile_X10Y6_FrameData_O[19] ;
 wire \Tile_X10Y6_FrameData_O[1] ;
 wire \Tile_X10Y6_FrameData_O[20] ;
 wire \Tile_X10Y6_FrameData_O[21] ;
 wire \Tile_X10Y6_FrameData_O[22] ;
 wire \Tile_X10Y6_FrameData_O[23] ;
 wire \Tile_X10Y6_FrameData_O[24] ;
 wire \Tile_X10Y6_FrameData_O[25] ;
 wire \Tile_X10Y6_FrameData_O[26] ;
 wire \Tile_X10Y6_FrameData_O[27] ;
 wire \Tile_X10Y6_FrameData_O[28] ;
 wire \Tile_X10Y6_FrameData_O[29] ;
 wire \Tile_X10Y6_FrameData_O[2] ;
 wire \Tile_X10Y6_FrameData_O[30] ;
 wire \Tile_X10Y6_FrameData_O[31] ;
 wire \Tile_X10Y6_FrameData_O[3] ;
 wire \Tile_X10Y6_FrameData_O[4] ;
 wire \Tile_X10Y6_FrameData_O[5] ;
 wire \Tile_X10Y6_FrameData_O[6] ;
 wire \Tile_X10Y6_FrameData_O[7] ;
 wire \Tile_X10Y6_FrameData_O[8] ;
 wire \Tile_X10Y6_FrameData_O[9] ;
 wire \Tile_X10Y6_S1BEG[0] ;
 wire \Tile_X10Y6_S1BEG[1] ;
 wire \Tile_X10Y6_S1BEG[2] ;
 wire \Tile_X10Y6_S1BEG[3] ;
 wire \Tile_X10Y6_S2BEG[0] ;
 wire \Tile_X10Y6_S2BEG[1] ;
 wire \Tile_X10Y6_S2BEG[2] ;
 wire \Tile_X10Y6_S2BEG[3] ;
 wire \Tile_X10Y6_S2BEG[4] ;
 wire \Tile_X10Y6_S2BEG[5] ;
 wire \Tile_X10Y6_S2BEG[6] ;
 wire \Tile_X10Y6_S2BEG[7] ;
 wire \Tile_X10Y6_S2BEGb[0] ;
 wire \Tile_X10Y6_S2BEGb[1] ;
 wire \Tile_X10Y6_S2BEGb[2] ;
 wire \Tile_X10Y6_S2BEGb[3] ;
 wire \Tile_X10Y6_S2BEGb[4] ;
 wire \Tile_X10Y6_S2BEGb[5] ;
 wire \Tile_X10Y6_S2BEGb[6] ;
 wire \Tile_X10Y6_S2BEGb[7] ;
 wire \Tile_X10Y6_S4BEG[0] ;
 wire \Tile_X10Y6_S4BEG[10] ;
 wire \Tile_X10Y6_S4BEG[11] ;
 wire \Tile_X10Y6_S4BEG[12] ;
 wire \Tile_X10Y6_S4BEG[13] ;
 wire \Tile_X10Y6_S4BEG[14] ;
 wire \Tile_X10Y6_S4BEG[15] ;
 wire \Tile_X10Y6_S4BEG[1] ;
 wire \Tile_X10Y6_S4BEG[2] ;
 wire \Tile_X10Y6_S4BEG[3] ;
 wire \Tile_X10Y6_S4BEG[4] ;
 wire \Tile_X10Y6_S4BEG[5] ;
 wire \Tile_X10Y6_S4BEG[6] ;
 wire \Tile_X10Y6_S4BEG[7] ;
 wire \Tile_X10Y6_S4BEG[8] ;
 wire \Tile_X10Y6_S4BEG[9] ;
 wire \Tile_X10Y6_W1BEG[0] ;
 wire \Tile_X10Y6_W1BEG[1] ;
 wire \Tile_X10Y6_W1BEG[2] ;
 wire \Tile_X10Y6_W1BEG[3] ;
 wire \Tile_X10Y6_W2BEG[0] ;
 wire \Tile_X10Y6_W2BEG[1] ;
 wire \Tile_X10Y6_W2BEG[2] ;
 wire \Tile_X10Y6_W2BEG[3] ;
 wire \Tile_X10Y6_W2BEG[4] ;
 wire \Tile_X10Y6_W2BEG[5] ;
 wire \Tile_X10Y6_W2BEG[6] ;
 wire \Tile_X10Y6_W2BEG[7] ;
 wire \Tile_X10Y6_W2BEGb[0] ;
 wire \Tile_X10Y6_W2BEGb[1] ;
 wire \Tile_X10Y6_W2BEGb[2] ;
 wire \Tile_X10Y6_W2BEGb[3] ;
 wire \Tile_X10Y6_W2BEGb[4] ;
 wire \Tile_X10Y6_W2BEGb[5] ;
 wire \Tile_X10Y6_W2BEGb[6] ;
 wire \Tile_X10Y6_W2BEGb[7] ;
 wire \Tile_X10Y6_W6BEG[0] ;
 wire \Tile_X10Y6_W6BEG[10] ;
 wire \Tile_X10Y6_W6BEG[11] ;
 wire \Tile_X10Y6_W6BEG[1] ;
 wire \Tile_X10Y6_W6BEG[2] ;
 wire \Tile_X10Y6_W6BEG[3] ;
 wire \Tile_X10Y6_W6BEG[4] ;
 wire \Tile_X10Y6_W6BEG[5] ;
 wire \Tile_X10Y6_W6BEG[6] ;
 wire \Tile_X10Y6_W6BEG[7] ;
 wire \Tile_X10Y6_W6BEG[8] ;
 wire \Tile_X10Y6_W6BEG[9] ;
 wire \Tile_X10Y6_WW4BEG[0] ;
 wire \Tile_X10Y6_WW4BEG[10] ;
 wire \Tile_X10Y6_WW4BEG[11] ;
 wire \Tile_X10Y6_WW4BEG[12] ;
 wire \Tile_X10Y6_WW4BEG[13] ;
 wire \Tile_X10Y6_WW4BEG[14] ;
 wire \Tile_X10Y6_WW4BEG[15] ;
 wire \Tile_X10Y6_WW4BEG[1] ;
 wire \Tile_X10Y6_WW4BEG[2] ;
 wire \Tile_X10Y6_WW4BEG[3] ;
 wire \Tile_X10Y6_WW4BEG[4] ;
 wire \Tile_X10Y6_WW4BEG[5] ;
 wire \Tile_X10Y6_WW4BEG[6] ;
 wire \Tile_X10Y6_WW4BEG[7] ;
 wire \Tile_X10Y6_WW4BEG[8] ;
 wire \Tile_X10Y6_WW4BEG[9] ;
 wire \Tile_X10Y7_FrameData_O[0] ;
 wire \Tile_X10Y7_FrameData_O[10] ;
 wire \Tile_X10Y7_FrameData_O[11] ;
 wire \Tile_X10Y7_FrameData_O[12] ;
 wire \Tile_X10Y7_FrameData_O[13] ;
 wire \Tile_X10Y7_FrameData_O[14] ;
 wire \Tile_X10Y7_FrameData_O[15] ;
 wire \Tile_X10Y7_FrameData_O[16] ;
 wire \Tile_X10Y7_FrameData_O[17] ;
 wire \Tile_X10Y7_FrameData_O[18] ;
 wire \Tile_X10Y7_FrameData_O[19] ;
 wire \Tile_X10Y7_FrameData_O[1] ;
 wire \Tile_X10Y7_FrameData_O[20] ;
 wire \Tile_X10Y7_FrameData_O[21] ;
 wire \Tile_X10Y7_FrameData_O[22] ;
 wire \Tile_X10Y7_FrameData_O[23] ;
 wire \Tile_X10Y7_FrameData_O[24] ;
 wire \Tile_X10Y7_FrameData_O[25] ;
 wire \Tile_X10Y7_FrameData_O[26] ;
 wire \Tile_X10Y7_FrameData_O[27] ;
 wire \Tile_X10Y7_FrameData_O[28] ;
 wire \Tile_X10Y7_FrameData_O[29] ;
 wire \Tile_X10Y7_FrameData_O[2] ;
 wire \Tile_X10Y7_FrameData_O[30] ;
 wire \Tile_X10Y7_FrameData_O[31] ;
 wire \Tile_X10Y7_FrameData_O[3] ;
 wire \Tile_X10Y7_FrameData_O[4] ;
 wire \Tile_X10Y7_FrameData_O[5] ;
 wire \Tile_X10Y7_FrameData_O[6] ;
 wire \Tile_X10Y7_FrameData_O[7] ;
 wire \Tile_X10Y7_FrameData_O[8] ;
 wire \Tile_X10Y7_FrameData_O[9] ;
 wire \Tile_X10Y7_FrameStrobe_O[0] ;
 wire \Tile_X10Y7_FrameStrobe_O[10] ;
 wire \Tile_X10Y7_FrameStrobe_O[11] ;
 wire \Tile_X10Y7_FrameStrobe_O[12] ;
 wire \Tile_X10Y7_FrameStrobe_O[13] ;
 wire \Tile_X10Y7_FrameStrobe_O[14] ;
 wire \Tile_X10Y7_FrameStrobe_O[15] ;
 wire \Tile_X10Y7_FrameStrobe_O[16] ;
 wire \Tile_X10Y7_FrameStrobe_O[17] ;
 wire \Tile_X10Y7_FrameStrobe_O[18] ;
 wire \Tile_X10Y7_FrameStrobe_O[19] ;
 wire \Tile_X10Y7_FrameStrobe_O[1] ;
 wire \Tile_X10Y7_FrameStrobe_O[2] ;
 wire \Tile_X10Y7_FrameStrobe_O[3] ;
 wire \Tile_X10Y7_FrameStrobe_O[4] ;
 wire \Tile_X10Y7_FrameStrobe_O[5] ;
 wire \Tile_X10Y7_FrameStrobe_O[6] ;
 wire \Tile_X10Y7_FrameStrobe_O[7] ;
 wire \Tile_X10Y7_FrameStrobe_O[8] ;
 wire \Tile_X10Y7_FrameStrobe_O[9] ;
 wire \Tile_X10Y7_N1BEG[0] ;
 wire \Tile_X10Y7_N1BEG[1] ;
 wire \Tile_X10Y7_N1BEG[2] ;
 wire \Tile_X10Y7_N1BEG[3] ;
 wire \Tile_X10Y7_N2BEG[0] ;
 wire \Tile_X10Y7_N2BEG[1] ;
 wire \Tile_X10Y7_N2BEG[2] ;
 wire \Tile_X10Y7_N2BEG[3] ;
 wire \Tile_X10Y7_N2BEG[4] ;
 wire \Tile_X10Y7_N2BEG[5] ;
 wire \Tile_X10Y7_N2BEG[6] ;
 wire \Tile_X10Y7_N2BEG[7] ;
 wire \Tile_X10Y7_N2BEGb[0] ;
 wire \Tile_X10Y7_N2BEGb[1] ;
 wire \Tile_X10Y7_N2BEGb[2] ;
 wire \Tile_X10Y7_N2BEGb[3] ;
 wire \Tile_X10Y7_N2BEGb[4] ;
 wire \Tile_X10Y7_N2BEGb[5] ;
 wire \Tile_X10Y7_N2BEGb[6] ;
 wire \Tile_X10Y7_N2BEGb[7] ;
 wire \Tile_X10Y7_N4BEG[0] ;
 wire \Tile_X10Y7_N4BEG[10] ;
 wire \Tile_X10Y7_N4BEG[11] ;
 wire \Tile_X10Y7_N4BEG[12] ;
 wire \Tile_X10Y7_N4BEG[13] ;
 wire \Tile_X10Y7_N4BEG[14] ;
 wire \Tile_X10Y7_N4BEG[15] ;
 wire \Tile_X10Y7_N4BEG[1] ;
 wire \Tile_X10Y7_N4BEG[2] ;
 wire \Tile_X10Y7_N4BEG[3] ;
 wire \Tile_X10Y7_N4BEG[4] ;
 wire \Tile_X10Y7_N4BEG[5] ;
 wire \Tile_X10Y7_N4BEG[6] ;
 wire \Tile_X10Y7_N4BEG[7] ;
 wire \Tile_X10Y7_N4BEG[8] ;
 wire \Tile_X10Y7_N4BEG[9] ;
 wire Tile_X10Y7_UserCLKo;
 wire \Tile_X10Y7_W1BEG[0] ;
 wire \Tile_X10Y7_W1BEG[1] ;
 wire \Tile_X10Y7_W1BEG[2] ;
 wire \Tile_X10Y7_W1BEG[3] ;
 wire \Tile_X10Y7_W2BEG[0] ;
 wire \Tile_X10Y7_W2BEG[1] ;
 wire \Tile_X10Y7_W2BEG[2] ;
 wire \Tile_X10Y7_W2BEG[3] ;
 wire \Tile_X10Y7_W2BEG[4] ;
 wire \Tile_X10Y7_W2BEG[5] ;
 wire \Tile_X10Y7_W2BEG[6] ;
 wire \Tile_X10Y7_W2BEG[7] ;
 wire \Tile_X10Y7_W2BEGb[0] ;
 wire \Tile_X10Y7_W2BEGb[1] ;
 wire \Tile_X10Y7_W2BEGb[2] ;
 wire \Tile_X10Y7_W2BEGb[3] ;
 wire \Tile_X10Y7_W2BEGb[4] ;
 wire \Tile_X10Y7_W2BEGb[5] ;
 wire \Tile_X10Y7_W2BEGb[6] ;
 wire \Tile_X10Y7_W2BEGb[7] ;
 wire \Tile_X10Y7_W6BEG[0] ;
 wire \Tile_X10Y7_W6BEG[10] ;
 wire \Tile_X10Y7_W6BEG[11] ;
 wire \Tile_X10Y7_W6BEG[1] ;
 wire \Tile_X10Y7_W6BEG[2] ;
 wire \Tile_X10Y7_W6BEG[3] ;
 wire \Tile_X10Y7_W6BEG[4] ;
 wire \Tile_X10Y7_W6BEG[5] ;
 wire \Tile_X10Y7_W6BEG[6] ;
 wire \Tile_X10Y7_W6BEG[7] ;
 wire \Tile_X10Y7_W6BEG[8] ;
 wire \Tile_X10Y7_W6BEG[9] ;
 wire \Tile_X10Y7_WW4BEG[0] ;
 wire \Tile_X10Y7_WW4BEG[10] ;
 wire \Tile_X10Y7_WW4BEG[11] ;
 wire \Tile_X10Y7_WW4BEG[12] ;
 wire \Tile_X10Y7_WW4BEG[13] ;
 wire \Tile_X10Y7_WW4BEG[14] ;
 wire \Tile_X10Y7_WW4BEG[15] ;
 wire \Tile_X10Y7_WW4BEG[1] ;
 wire \Tile_X10Y7_WW4BEG[2] ;
 wire \Tile_X10Y7_WW4BEG[3] ;
 wire \Tile_X10Y7_WW4BEG[4] ;
 wire \Tile_X10Y7_WW4BEG[5] ;
 wire \Tile_X10Y7_WW4BEG[6] ;
 wire \Tile_X10Y7_WW4BEG[7] ;
 wire \Tile_X10Y7_WW4BEG[8] ;
 wire \Tile_X10Y7_WW4BEG[9] ;
 wire \Tile_X10Y8_FrameData_O[0] ;
 wire \Tile_X10Y8_FrameData_O[10] ;
 wire \Tile_X10Y8_FrameData_O[11] ;
 wire \Tile_X10Y8_FrameData_O[12] ;
 wire \Tile_X10Y8_FrameData_O[13] ;
 wire \Tile_X10Y8_FrameData_O[14] ;
 wire \Tile_X10Y8_FrameData_O[15] ;
 wire \Tile_X10Y8_FrameData_O[16] ;
 wire \Tile_X10Y8_FrameData_O[17] ;
 wire \Tile_X10Y8_FrameData_O[18] ;
 wire \Tile_X10Y8_FrameData_O[19] ;
 wire \Tile_X10Y8_FrameData_O[1] ;
 wire \Tile_X10Y8_FrameData_O[20] ;
 wire \Tile_X10Y8_FrameData_O[21] ;
 wire \Tile_X10Y8_FrameData_O[22] ;
 wire \Tile_X10Y8_FrameData_O[23] ;
 wire \Tile_X10Y8_FrameData_O[24] ;
 wire \Tile_X10Y8_FrameData_O[25] ;
 wire \Tile_X10Y8_FrameData_O[26] ;
 wire \Tile_X10Y8_FrameData_O[27] ;
 wire \Tile_X10Y8_FrameData_O[28] ;
 wire \Tile_X10Y8_FrameData_O[29] ;
 wire \Tile_X10Y8_FrameData_O[2] ;
 wire \Tile_X10Y8_FrameData_O[30] ;
 wire \Tile_X10Y8_FrameData_O[31] ;
 wire \Tile_X10Y8_FrameData_O[3] ;
 wire \Tile_X10Y8_FrameData_O[4] ;
 wire \Tile_X10Y8_FrameData_O[5] ;
 wire \Tile_X10Y8_FrameData_O[6] ;
 wire \Tile_X10Y8_FrameData_O[7] ;
 wire \Tile_X10Y8_FrameData_O[8] ;
 wire \Tile_X10Y8_FrameData_O[9] ;
 wire \Tile_X10Y8_S1BEG[0] ;
 wire \Tile_X10Y8_S1BEG[1] ;
 wire \Tile_X10Y8_S1BEG[2] ;
 wire \Tile_X10Y8_S1BEG[3] ;
 wire \Tile_X10Y8_S2BEG[0] ;
 wire \Tile_X10Y8_S2BEG[1] ;
 wire \Tile_X10Y8_S2BEG[2] ;
 wire \Tile_X10Y8_S2BEG[3] ;
 wire \Tile_X10Y8_S2BEG[4] ;
 wire \Tile_X10Y8_S2BEG[5] ;
 wire \Tile_X10Y8_S2BEG[6] ;
 wire \Tile_X10Y8_S2BEG[7] ;
 wire \Tile_X10Y8_S2BEGb[0] ;
 wire \Tile_X10Y8_S2BEGb[1] ;
 wire \Tile_X10Y8_S2BEGb[2] ;
 wire \Tile_X10Y8_S2BEGb[3] ;
 wire \Tile_X10Y8_S2BEGb[4] ;
 wire \Tile_X10Y8_S2BEGb[5] ;
 wire \Tile_X10Y8_S2BEGb[6] ;
 wire \Tile_X10Y8_S2BEGb[7] ;
 wire \Tile_X10Y8_S4BEG[0] ;
 wire \Tile_X10Y8_S4BEG[10] ;
 wire \Tile_X10Y8_S4BEG[11] ;
 wire \Tile_X10Y8_S4BEG[12] ;
 wire \Tile_X10Y8_S4BEG[13] ;
 wire \Tile_X10Y8_S4BEG[14] ;
 wire \Tile_X10Y8_S4BEG[15] ;
 wire \Tile_X10Y8_S4BEG[1] ;
 wire \Tile_X10Y8_S4BEG[2] ;
 wire \Tile_X10Y8_S4BEG[3] ;
 wire \Tile_X10Y8_S4BEG[4] ;
 wire \Tile_X10Y8_S4BEG[5] ;
 wire \Tile_X10Y8_S4BEG[6] ;
 wire \Tile_X10Y8_S4BEG[7] ;
 wire \Tile_X10Y8_S4BEG[8] ;
 wire \Tile_X10Y8_S4BEG[9] ;
 wire \Tile_X10Y8_W1BEG[0] ;
 wire \Tile_X10Y8_W1BEG[1] ;
 wire \Tile_X10Y8_W1BEG[2] ;
 wire \Tile_X10Y8_W1BEG[3] ;
 wire \Tile_X10Y8_W2BEG[0] ;
 wire \Tile_X10Y8_W2BEG[1] ;
 wire \Tile_X10Y8_W2BEG[2] ;
 wire \Tile_X10Y8_W2BEG[3] ;
 wire \Tile_X10Y8_W2BEG[4] ;
 wire \Tile_X10Y8_W2BEG[5] ;
 wire \Tile_X10Y8_W2BEG[6] ;
 wire \Tile_X10Y8_W2BEG[7] ;
 wire \Tile_X10Y8_W2BEGb[0] ;
 wire \Tile_X10Y8_W2BEGb[1] ;
 wire \Tile_X10Y8_W2BEGb[2] ;
 wire \Tile_X10Y8_W2BEGb[3] ;
 wire \Tile_X10Y8_W2BEGb[4] ;
 wire \Tile_X10Y8_W2BEGb[5] ;
 wire \Tile_X10Y8_W2BEGb[6] ;
 wire \Tile_X10Y8_W2BEGb[7] ;
 wire \Tile_X10Y8_W6BEG[0] ;
 wire \Tile_X10Y8_W6BEG[10] ;
 wire \Tile_X10Y8_W6BEG[11] ;
 wire \Tile_X10Y8_W6BEG[1] ;
 wire \Tile_X10Y8_W6BEG[2] ;
 wire \Tile_X10Y8_W6BEG[3] ;
 wire \Tile_X10Y8_W6BEG[4] ;
 wire \Tile_X10Y8_W6BEG[5] ;
 wire \Tile_X10Y8_W6BEG[6] ;
 wire \Tile_X10Y8_W6BEG[7] ;
 wire \Tile_X10Y8_W6BEG[8] ;
 wire \Tile_X10Y8_W6BEG[9] ;
 wire \Tile_X10Y8_WW4BEG[0] ;
 wire \Tile_X10Y8_WW4BEG[10] ;
 wire \Tile_X10Y8_WW4BEG[11] ;
 wire \Tile_X10Y8_WW4BEG[12] ;
 wire \Tile_X10Y8_WW4BEG[13] ;
 wire \Tile_X10Y8_WW4BEG[14] ;
 wire \Tile_X10Y8_WW4BEG[15] ;
 wire \Tile_X10Y8_WW4BEG[1] ;
 wire \Tile_X10Y8_WW4BEG[2] ;
 wire \Tile_X10Y8_WW4BEG[3] ;
 wire \Tile_X10Y8_WW4BEG[4] ;
 wire \Tile_X10Y8_WW4BEG[5] ;
 wire \Tile_X10Y8_WW4BEG[6] ;
 wire \Tile_X10Y8_WW4BEG[7] ;
 wire \Tile_X10Y8_WW4BEG[8] ;
 wire \Tile_X10Y8_WW4BEG[9] ;
 wire \Tile_X10Y9_FrameData_O[0] ;
 wire \Tile_X10Y9_FrameData_O[10] ;
 wire \Tile_X10Y9_FrameData_O[11] ;
 wire \Tile_X10Y9_FrameData_O[12] ;
 wire \Tile_X10Y9_FrameData_O[13] ;
 wire \Tile_X10Y9_FrameData_O[14] ;
 wire \Tile_X10Y9_FrameData_O[15] ;
 wire \Tile_X10Y9_FrameData_O[16] ;
 wire \Tile_X10Y9_FrameData_O[17] ;
 wire \Tile_X10Y9_FrameData_O[18] ;
 wire \Tile_X10Y9_FrameData_O[19] ;
 wire \Tile_X10Y9_FrameData_O[1] ;
 wire \Tile_X10Y9_FrameData_O[20] ;
 wire \Tile_X10Y9_FrameData_O[21] ;
 wire \Tile_X10Y9_FrameData_O[22] ;
 wire \Tile_X10Y9_FrameData_O[23] ;
 wire \Tile_X10Y9_FrameData_O[24] ;
 wire \Tile_X10Y9_FrameData_O[25] ;
 wire \Tile_X10Y9_FrameData_O[26] ;
 wire \Tile_X10Y9_FrameData_O[27] ;
 wire \Tile_X10Y9_FrameData_O[28] ;
 wire \Tile_X10Y9_FrameData_O[29] ;
 wire \Tile_X10Y9_FrameData_O[2] ;
 wire \Tile_X10Y9_FrameData_O[30] ;
 wire \Tile_X10Y9_FrameData_O[31] ;
 wire \Tile_X10Y9_FrameData_O[3] ;
 wire \Tile_X10Y9_FrameData_O[4] ;
 wire \Tile_X10Y9_FrameData_O[5] ;
 wire \Tile_X10Y9_FrameData_O[6] ;
 wire \Tile_X10Y9_FrameData_O[7] ;
 wire \Tile_X10Y9_FrameData_O[8] ;
 wire \Tile_X10Y9_FrameData_O[9] ;
 wire \Tile_X10Y9_FrameStrobe_O[0] ;
 wire \Tile_X10Y9_FrameStrobe_O[10] ;
 wire \Tile_X10Y9_FrameStrobe_O[11] ;
 wire \Tile_X10Y9_FrameStrobe_O[12] ;
 wire \Tile_X10Y9_FrameStrobe_O[13] ;
 wire \Tile_X10Y9_FrameStrobe_O[14] ;
 wire \Tile_X10Y9_FrameStrobe_O[15] ;
 wire \Tile_X10Y9_FrameStrobe_O[16] ;
 wire \Tile_X10Y9_FrameStrobe_O[17] ;
 wire \Tile_X10Y9_FrameStrobe_O[18] ;
 wire \Tile_X10Y9_FrameStrobe_O[19] ;
 wire \Tile_X10Y9_FrameStrobe_O[1] ;
 wire \Tile_X10Y9_FrameStrobe_O[2] ;
 wire \Tile_X10Y9_FrameStrobe_O[3] ;
 wire \Tile_X10Y9_FrameStrobe_O[4] ;
 wire \Tile_X10Y9_FrameStrobe_O[5] ;
 wire \Tile_X10Y9_FrameStrobe_O[6] ;
 wire \Tile_X10Y9_FrameStrobe_O[7] ;
 wire \Tile_X10Y9_FrameStrobe_O[8] ;
 wire \Tile_X10Y9_FrameStrobe_O[9] ;
 wire \Tile_X10Y9_N1BEG[0] ;
 wire \Tile_X10Y9_N1BEG[1] ;
 wire \Tile_X10Y9_N1BEG[2] ;
 wire \Tile_X10Y9_N1BEG[3] ;
 wire \Tile_X10Y9_N2BEG[0] ;
 wire \Tile_X10Y9_N2BEG[1] ;
 wire \Tile_X10Y9_N2BEG[2] ;
 wire \Tile_X10Y9_N2BEG[3] ;
 wire \Tile_X10Y9_N2BEG[4] ;
 wire \Tile_X10Y9_N2BEG[5] ;
 wire \Tile_X10Y9_N2BEG[6] ;
 wire \Tile_X10Y9_N2BEG[7] ;
 wire \Tile_X10Y9_N2BEGb[0] ;
 wire \Tile_X10Y9_N2BEGb[1] ;
 wire \Tile_X10Y9_N2BEGb[2] ;
 wire \Tile_X10Y9_N2BEGb[3] ;
 wire \Tile_X10Y9_N2BEGb[4] ;
 wire \Tile_X10Y9_N2BEGb[5] ;
 wire \Tile_X10Y9_N2BEGb[6] ;
 wire \Tile_X10Y9_N2BEGb[7] ;
 wire \Tile_X10Y9_N4BEG[0] ;
 wire \Tile_X10Y9_N4BEG[10] ;
 wire \Tile_X10Y9_N4BEG[11] ;
 wire \Tile_X10Y9_N4BEG[12] ;
 wire \Tile_X10Y9_N4BEG[13] ;
 wire \Tile_X10Y9_N4BEG[14] ;
 wire \Tile_X10Y9_N4BEG[15] ;
 wire \Tile_X10Y9_N4BEG[1] ;
 wire \Tile_X10Y9_N4BEG[2] ;
 wire \Tile_X10Y9_N4BEG[3] ;
 wire \Tile_X10Y9_N4BEG[4] ;
 wire \Tile_X10Y9_N4BEG[5] ;
 wire \Tile_X10Y9_N4BEG[6] ;
 wire \Tile_X10Y9_N4BEG[7] ;
 wire \Tile_X10Y9_N4BEG[8] ;
 wire \Tile_X10Y9_N4BEG[9] ;
 wire Tile_X10Y9_UserCLKo;
 wire \Tile_X10Y9_W1BEG[0] ;
 wire \Tile_X10Y9_W1BEG[1] ;
 wire \Tile_X10Y9_W1BEG[2] ;
 wire \Tile_X10Y9_W1BEG[3] ;
 wire \Tile_X10Y9_W2BEG[0] ;
 wire \Tile_X10Y9_W2BEG[1] ;
 wire \Tile_X10Y9_W2BEG[2] ;
 wire \Tile_X10Y9_W2BEG[3] ;
 wire \Tile_X10Y9_W2BEG[4] ;
 wire \Tile_X10Y9_W2BEG[5] ;
 wire \Tile_X10Y9_W2BEG[6] ;
 wire \Tile_X10Y9_W2BEG[7] ;
 wire \Tile_X10Y9_W2BEGb[0] ;
 wire \Tile_X10Y9_W2BEGb[1] ;
 wire \Tile_X10Y9_W2BEGb[2] ;
 wire \Tile_X10Y9_W2BEGb[3] ;
 wire \Tile_X10Y9_W2BEGb[4] ;
 wire \Tile_X10Y9_W2BEGb[5] ;
 wire \Tile_X10Y9_W2BEGb[6] ;
 wire \Tile_X10Y9_W2BEGb[7] ;
 wire \Tile_X10Y9_W6BEG[0] ;
 wire \Tile_X10Y9_W6BEG[10] ;
 wire \Tile_X10Y9_W6BEG[11] ;
 wire \Tile_X10Y9_W6BEG[1] ;
 wire \Tile_X10Y9_W6BEG[2] ;
 wire \Tile_X10Y9_W6BEG[3] ;
 wire \Tile_X10Y9_W6BEG[4] ;
 wire \Tile_X10Y9_W6BEG[5] ;
 wire \Tile_X10Y9_W6BEG[6] ;
 wire \Tile_X10Y9_W6BEG[7] ;
 wire \Tile_X10Y9_W6BEG[8] ;
 wire \Tile_X10Y9_W6BEG[9] ;
 wire \Tile_X10Y9_WW4BEG[0] ;
 wire \Tile_X10Y9_WW4BEG[10] ;
 wire \Tile_X10Y9_WW4BEG[11] ;
 wire \Tile_X10Y9_WW4BEG[12] ;
 wire \Tile_X10Y9_WW4BEG[13] ;
 wire \Tile_X10Y9_WW4BEG[14] ;
 wire \Tile_X10Y9_WW4BEG[15] ;
 wire \Tile_X10Y9_WW4BEG[1] ;
 wire \Tile_X10Y9_WW4BEG[2] ;
 wire \Tile_X10Y9_WW4BEG[3] ;
 wire \Tile_X10Y9_WW4BEG[4] ;
 wire \Tile_X10Y9_WW4BEG[5] ;
 wire \Tile_X10Y9_WW4BEG[6] ;
 wire \Tile_X10Y9_WW4BEG[7] ;
 wire \Tile_X10Y9_WW4BEG[8] ;
 wire \Tile_X10Y9_WW4BEG[9] ;
 wire \Tile_X1Y0_FrameData_O[0] ;
 wire \Tile_X1Y0_FrameData_O[10] ;
 wire \Tile_X1Y0_FrameData_O[11] ;
 wire \Tile_X1Y0_FrameData_O[12] ;
 wire \Tile_X1Y0_FrameData_O[13] ;
 wire \Tile_X1Y0_FrameData_O[14] ;
 wire \Tile_X1Y0_FrameData_O[15] ;
 wire \Tile_X1Y0_FrameData_O[16] ;
 wire \Tile_X1Y0_FrameData_O[17] ;
 wire \Tile_X1Y0_FrameData_O[18] ;
 wire \Tile_X1Y0_FrameData_O[19] ;
 wire \Tile_X1Y0_FrameData_O[1] ;
 wire \Tile_X1Y0_FrameData_O[20] ;
 wire \Tile_X1Y0_FrameData_O[21] ;
 wire \Tile_X1Y0_FrameData_O[22] ;
 wire \Tile_X1Y0_FrameData_O[23] ;
 wire \Tile_X1Y0_FrameData_O[24] ;
 wire \Tile_X1Y0_FrameData_O[25] ;
 wire \Tile_X1Y0_FrameData_O[26] ;
 wire \Tile_X1Y0_FrameData_O[27] ;
 wire \Tile_X1Y0_FrameData_O[28] ;
 wire \Tile_X1Y0_FrameData_O[29] ;
 wire \Tile_X1Y0_FrameData_O[2] ;
 wire \Tile_X1Y0_FrameData_O[30] ;
 wire \Tile_X1Y0_FrameData_O[31] ;
 wire \Tile_X1Y0_FrameData_O[3] ;
 wire \Tile_X1Y0_FrameData_O[4] ;
 wire \Tile_X1Y0_FrameData_O[5] ;
 wire \Tile_X1Y0_FrameData_O[6] ;
 wire \Tile_X1Y0_FrameData_O[7] ;
 wire \Tile_X1Y0_FrameData_O[8] ;
 wire \Tile_X1Y0_FrameData_O[9] ;
 wire \Tile_X1Y0_FrameStrobe_O[0] ;
 wire \Tile_X1Y0_FrameStrobe_O[10] ;
 wire \Tile_X1Y0_FrameStrobe_O[11] ;
 wire \Tile_X1Y0_FrameStrobe_O[12] ;
 wire \Tile_X1Y0_FrameStrobe_O[13] ;
 wire \Tile_X1Y0_FrameStrobe_O[14] ;
 wire \Tile_X1Y0_FrameStrobe_O[15] ;
 wire \Tile_X1Y0_FrameStrobe_O[16] ;
 wire \Tile_X1Y0_FrameStrobe_O[17] ;
 wire \Tile_X1Y0_FrameStrobe_O[18] ;
 wire \Tile_X1Y0_FrameStrobe_O[19] ;
 wire \Tile_X1Y0_FrameStrobe_O[1] ;
 wire \Tile_X1Y0_FrameStrobe_O[2] ;
 wire \Tile_X1Y0_FrameStrobe_O[3] ;
 wire \Tile_X1Y0_FrameStrobe_O[4] ;
 wire \Tile_X1Y0_FrameStrobe_O[5] ;
 wire \Tile_X1Y0_FrameStrobe_O[6] ;
 wire \Tile_X1Y0_FrameStrobe_O[7] ;
 wire \Tile_X1Y0_FrameStrobe_O[8] ;
 wire \Tile_X1Y0_FrameStrobe_O[9] ;
 wire \Tile_X1Y0_S1BEG[0] ;
 wire \Tile_X1Y0_S1BEG[1] ;
 wire \Tile_X1Y0_S1BEG[2] ;
 wire \Tile_X1Y0_S1BEG[3] ;
 wire \Tile_X1Y0_S2BEG[0] ;
 wire \Tile_X1Y0_S2BEG[1] ;
 wire \Tile_X1Y0_S2BEG[2] ;
 wire \Tile_X1Y0_S2BEG[3] ;
 wire \Tile_X1Y0_S2BEG[4] ;
 wire \Tile_X1Y0_S2BEG[5] ;
 wire \Tile_X1Y0_S2BEG[6] ;
 wire \Tile_X1Y0_S2BEG[7] ;
 wire \Tile_X1Y0_S2BEGb[0] ;
 wire \Tile_X1Y0_S2BEGb[1] ;
 wire \Tile_X1Y0_S2BEGb[2] ;
 wire \Tile_X1Y0_S2BEGb[3] ;
 wire \Tile_X1Y0_S2BEGb[4] ;
 wire \Tile_X1Y0_S2BEGb[5] ;
 wire \Tile_X1Y0_S2BEGb[6] ;
 wire \Tile_X1Y0_S2BEGb[7] ;
 wire \Tile_X1Y0_S4BEG[0] ;
 wire \Tile_X1Y0_S4BEG[10] ;
 wire \Tile_X1Y0_S4BEG[11] ;
 wire \Tile_X1Y0_S4BEG[12] ;
 wire \Tile_X1Y0_S4BEG[13] ;
 wire \Tile_X1Y0_S4BEG[14] ;
 wire \Tile_X1Y0_S4BEG[15] ;
 wire \Tile_X1Y0_S4BEG[1] ;
 wire \Tile_X1Y0_S4BEG[2] ;
 wire \Tile_X1Y0_S4BEG[3] ;
 wire \Tile_X1Y0_S4BEG[4] ;
 wire \Tile_X1Y0_S4BEG[5] ;
 wire \Tile_X1Y0_S4BEG[6] ;
 wire \Tile_X1Y0_S4BEG[7] ;
 wire \Tile_X1Y0_S4BEG[8] ;
 wire \Tile_X1Y0_S4BEG[9] ;
 wire \Tile_X1Y0_SS4BEG[0] ;
 wire \Tile_X1Y0_SS4BEG[10] ;
 wire \Tile_X1Y0_SS4BEG[11] ;
 wire \Tile_X1Y0_SS4BEG[12] ;
 wire \Tile_X1Y0_SS4BEG[13] ;
 wire \Tile_X1Y0_SS4BEG[14] ;
 wire \Tile_X1Y0_SS4BEG[15] ;
 wire \Tile_X1Y0_SS4BEG[1] ;
 wire \Tile_X1Y0_SS4BEG[2] ;
 wire \Tile_X1Y0_SS4BEG[3] ;
 wire \Tile_X1Y0_SS4BEG[4] ;
 wire \Tile_X1Y0_SS4BEG[5] ;
 wire \Tile_X1Y0_SS4BEG[6] ;
 wire \Tile_X1Y0_SS4BEG[7] ;
 wire \Tile_X1Y0_SS4BEG[8] ;
 wire \Tile_X1Y0_SS4BEG[9] ;
 wire Tile_X1Y0_UserCLKo;
 wire Tile_X1Y10_Co;
 wire \Tile_X1Y10_E1BEG[0] ;
 wire \Tile_X1Y10_E1BEG[1] ;
 wire \Tile_X1Y10_E1BEG[2] ;
 wire \Tile_X1Y10_E1BEG[3] ;
 wire \Tile_X1Y10_E2BEG[0] ;
 wire \Tile_X1Y10_E2BEG[1] ;
 wire \Tile_X1Y10_E2BEG[2] ;
 wire \Tile_X1Y10_E2BEG[3] ;
 wire \Tile_X1Y10_E2BEG[4] ;
 wire \Tile_X1Y10_E2BEG[5] ;
 wire \Tile_X1Y10_E2BEG[6] ;
 wire \Tile_X1Y10_E2BEG[7] ;
 wire \Tile_X1Y10_E2BEGb[0] ;
 wire \Tile_X1Y10_E2BEGb[1] ;
 wire \Tile_X1Y10_E2BEGb[2] ;
 wire \Tile_X1Y10_E2BEGb[3] ;
 wire \Tile_X1Y10_E2BEGb[4] ;
 wire \Tile_X1Y10_E2BEGb[5] ;
 wire \Tile_X1Y10_E2BEGb[6] ;
 wire \Tile_X1Y10_E2BEGb[7] ;
 wire \Tile_X1Y10_E6BEG[0] ;
 wire \Tile_X1Y10_E6BEG[10] ;
 wire \Tile_X1Y10_E6BEG[11] ;
 wire \Tile_X1Y10_E6BEG[1] ;
 wire \Tile_X1Y10_E6BEG[2] ;
 wire \Tile_X1Y10_E6BEG[3] ;
 wire \Tile_X1Y10_E6BEG[4] ;
 wire \Tile_X1Y10_E6BEG[5] ;
 wire \Tile_X1Y10_E6BEG[6] ;
 wire \Tile_X1Y10_E6BEG[7] ;
 wire \Tile_X1Y10_E6BEG[8] ;
 wire \Tile_X1Y10_E6BEG[9] ;
 wire \Tile_X1Y10_EE4BEG[0] ;
 wire \Tile_X1Y10_EE4BEG[10] ;
 wire \Tile_X1Y10_EE4BEG[11] ;
 wire \Tile_X1Y10_EE4BEG[12] ;
 wire \Tile_X1Y10_EE4BEG[13] ;
 wire \Tile_X1Y10_EE4BEG[14] ;
 wire \Tile_X1Y10_EE4BEG[15] ;
 wire \Tile_X1Y10_EE4BEG[1] ;
 wire \Tile_X1Y10_EE4BEG[2] ;
 wire \Tile_X1Y10_EE4BEG[3] ;
 wire \Tile_X1Y10_EE4BEG[4] ;
 wire \Tile_X1Y10_EE4BEG[5] ;
 wire \Tile_X1Y10_EE4BEG[6] ;
 wire \Tile_X1Y10_EE4BEG[7] ;
 wire \Tile_X1Y10_EE4BEG[8] ;
 wire \Tile_X1Y10_EE4BEG[9] ;
 wire \Tile_X1Y10_FrameData_O[0] ;
 wire \Tile_X1Y10_FrameData_O[10] ;
 wire \Tile_X1Y10_FrameData_O[11] ;
 wire \Tile_X1Y10_FrameData_O[12] ;
 wire \Tile_X1Y10_FrameData_O[13] ;
 wire \Tile_X1Y10_FrameData_O[14] ;
 wire \Tile_X1Y10_FrameData_O[15] ;
 wire \Tile_X1Y10_FrameData_O[16] ;
 wire \Tile_X1Y10_FrameData_O[17] ;
 wire \Tile_X1Y10_FrameData_O[18] ;
 wire \Tile_X1Y10_FrameData_O[19] ;
 wire \Tile_X1Y10_FrameData_O[1] ;
 wire \Tile_X1Y10_FrameData_O[20] ;
 wire \Tile_X1Y10_FrameData_O[21] ;
 wire \Tile_X1Y10_FrameData_O[22] ;
 wire \Tile_X1Y10_FrameData_O[23] ;
 wire \Tile_X1Y10_FrameData_O[24] ;
 wire \Tile_X1Y10_FrameData_O[25] ;
 wire \Tile_X1Y10_FrameData_O[26] ;
 wire \Tile_X1Y10_FrameData_O[27] ;
 wire \Tile_X1Y10_FrameData_O[28] ;
 wire \Tile_X1Y10_FrameData_O[29] ;
 wire \Tile_X1Y10_FrameData_O[2] ;
 wire \Tile_X1Y10_FrameData_O[30] ;
 wire \Tile_X1Y10_FrameData_O[31] ;
 wire \Tile_X1Y10_FrameData_O[3] ;
 wire \Tile_X1Y10_FrameData_O[4] ;
 wire \Tile_X1Y10_FrameData_O[5] ;
 wire \Tile_X1Y10_FrameData_O[6] ;
 wire \Tile_X1Y10_FrameData_O[7] ;
 wire \Tile_X1Y10_FrameData_O[8] ;
 wire \Tile_X1Y10_FrameData_O[9] ;
 wire \Tile_X1Y10_FrameStrobe_O[0] ;
 wire \Tile_X1Y10_FrameStrobe_O[10] ;
 wire \Tile_X1Y10_FrameStrobe_O[11] ;
 wire \Tile_X1Y10_FrameStrobe_O[12] ;
 wire \Tile_X1Y10_FrameStrobe_O[13] ;
 wire \Tile_X1Y10_FrameStrobe_O[14] ;
 wire \Tile_X1Y10_FrameStrobe_O[15] ;
 wire \Tile_X1Y10_FrameStrobe_O[16] ;
 wire \Tile_X1Y10_FrameStrobe_O[17] ;
 wire \Tile_X1Y10_FrameStrobe_O[18] ;
 wire \Tile_X1Y10_FrameStrobe_O[19] ;
 wire \Tile_X1Y10_FrameStrobe_O[1] ;
 wire \Tile_X1Y10_FrameStrobe_O[2] ;
 wire \Tile_X1Y10_FrameStrobe_O[3] ;
 wire \Tile_X1Y10_FrameStrobe_O[4] ;
 wire \Tile_X1Y10_FrameStrobe_O[5] ;
 wire \Tile_X1Y10_FrameStrobe_O[6] ;
 wire \Tile_X1Y10_FrameStrobe_O[7] ;
 wire \Tile_X1Y10_FrameStrobe_O[8] ;
 wire \Tile_X1Y10_FrameStrobe_O[9] ;
 wire \Tile_X1Y10_N1BEG[0] ;
 wire \Tile_X1Y10_N1BEG[1] ;
 wire \Tile_X1Y10_N1BEG[2] ;
 wire \Tile_X1Y10_N1BEG[3] ;
 wire \Tile_X1Y10_N2BEG[0] ;
 wire \Tile_X1Y10_N2BEG[1] ;
 wire \Tile_X1Y10_N2BEG[2] ;
 wire \Tile_X1Y10_N2BEG[3] ;
 wire \Tile_X1Y10_N2BEG[4] ;
 wire \Tile_X1Y10_N2BEG[5] ;
 wire \Tile_X1Y10_N2BEG[6] ;
 wire \Tile_X1Y10_N2BEG[7] ;
 wire \Tile_X1Y10_N2BEGb[0] ;
 wire \Tile_X1Y10_N2BEGb[1] ;
 wire \Tile_X1Y10_N2BEGb[2] ;
 wire \Tile_X1Y10_N2BEGb[3] ;
 wire \Tile_X1Y10_N2BEGb[4] ;
 wire \Tile_X1Y10_N2BEGb[5] ;
 wire \Tile_X1Y10_N2BEGb[6] ;
 wire \Tile_X1Y10_N2BEGb[7] ;
 wire \Tile_X1Y10_N4BEG[0] ;
 wire \Tile_X1Y10_N4BEG[10] ;
 wire \Tile_X1Y10_N4BEG[11] ;
 wire \Tile_X1Y10_N4BEG[12] ;
 wire \Tile_X1Y10_N4BEG[13] ;
 wire \Tile_X1Y10_N4BEG[14] ;
 wire \Tile_X1Y10_N4BEG[15] ;
 wire \Tile_X1Y10_N4BEG[1] ;
 wire \Tile_X1Y10_N4BEG[2] ;
 wire \Tile_X1Y10_N4BEG[3] ;
 wire \Tile_X1Y10_N4BEG[4] ;
 wire \Tile_X1Y10_N4BEG[5] ;
 wire \Tile_X1Y10_N4BEG[6] ;
 wire \Tile_X1Y10_N4BEG[7] ;
 wire \Tile_X1Y10_N4BEG[8] ;
 wire \Tile_X1Y10_N4BEG[9] ;
 wire \Tile_X1Y10_NN4BEG[0] ;
 wire \Tile_X1Y10_NN4BEG[10] ;
 wire \Tile_X1Y10_NN4BEG[11] ;
 wire \Tile_X1Y10_NN4BEG[12] ;
 wire \Tile_X1Y10_NN4BEG[13] ;
 wire \Tile_X1Y10_NN4BEG[14] ;
 wire \Tile_X1Y10_NN4BEG[15] ;
 wire \Tile_X1Y10_NN4BEG[1] ;
 wire \Tile_X1Y10_NN4BEG[2] ;
 wire \Tile_X1Y10_NN4BEG[3] ;
 wire \Tile_X1Y10_NN4BEG[4] ;
 wire \Tile_X1Y10_NN4BEG[5] ;
 wire \Tile_X1Y10_NN4BEG[6] ;
 wire \Tile_X1Y10_NN4BEG[7] ;
 wire \Tile_X1Y10_NN4BEG[8] ;
 wire \Tile_X1Y10_NN4BEG[9] ;
 wire \Tile_X1Y10_S1BEG[0] ;
 wire \Tile_X1Y10_S1BEG[1] ;
 wire \Tile_X1Y10_S1BEG[2] ;
 wire \Tile_X1Y10_S1BEG[3] ;
 wire \Tile_X1Y10_S2BEG[0] ;
 wire \Tile_X1Y10_S2BEG[1] ;
 wire \Tile_X1Y10_S2BEG[2] ;
 wire \Tile_X1Y10_S2BEG[3] ;
 wire \Tile_X1Y10_S2BEG[4] ;
 wire \Tile_X1Y10_S2BEG[5] ;
 wire \Tile_X1Y10_S2BEG[6] ;
 wire \Tile_X1Y10_S2BEG[7] ;
 wire \Tile_X1Y10_S2BEGb[0] ;
 wire \Tile_X1Y10_S2BEGb[1] ;
 wire \Tile_X1Y10_S2BEGb[2] ;
 wire \Tile_X1Y10_S2BEGb[3] ;
 wire \Tile_X1Y10_S2BEGb[4] ;
 wire \Tile_X1Y10_S2BEGb[5] ;
 wire \Tile_X1Y10_S2BEGb[6] ;
 wire \Tile_X1Y10_S2BEGb[7] ;
 wire \Tile_X1Y10_S4BEG[0] ;
 wire \Tile_X1Y10_S4BEG[10] ;
 wire \Tile_X1Y10_S4BEG[11] ;
 wire \Tile_X1Y10_S4BEG[12] ;
 wire \Tile_X1Y10_S4BEG[13] ;
 wire \Tile_X1Y10_S4BEG[14] ;
 wire \Tile_X1Y10_S4BEG[15] ;
 wire \Tile_X1Y10_S4BEG[1] ;
 wire \Tile_X1Y10_S4BEG[2] ;
 wire \Tile_X1Y10_S4BEG[3] ;
 wire \Tile_X1Y10_S4BEG[4] ;
 wire \Tile_X1Y10_S4BEG[5] ;
 wire \Tile_X1Y10_S4BEG[6] ;
 wire \Tile_X1Y10_S4BEG[7] ;
 wire \Tile_X1Y10_S4BEG[8] ;
 wire \Tile_X1Y10_S4BEG[9] ;
 wire \Tile_X1Y10_SS4BEG[0] ;
 wire \Tile_X1Y10_SS4BEG[10] ;
 wire \Tile_X1Y10_SS4BEG[11] ;
 wire \Tile_X1Y10_SS4BEG[12] ;
 wire \Tile_X1Y10_SS4BEG[13] ;
 wire \Tile_X1Y10_SS4BEG[14] ;
 wire \Tile_X1Y10_SS4BEG[15] ;
 wire \Tile_X1Y10_SS4BEG[1] ;
 wire \Tile_X1Y10_SS4BEG[2] ;
 wire \Tile_X1Y10_SS4BEG[3] ;
 wire \Tile_X1Y10_SS4BEG[4] ;
 wire \Tile_X1Y10_SS4BEG[5] ;
 wire \Tile_X1Y10_SS4BEG[6] ;
 wire \Tile_X1Y10_SS4BEG[7] ;
 wire \Tile_X1Y10_SS4BEG[8] ;
 wire \Tile_X1Y10_SS4BEG[9] ;
 wire Tile_X1Y10_UserCLKo;
 wire \Tile_X1Y10_W1BEG[0] ;
 wire \Tile_X1Y10_W1BEG[1] ;
 wire \Tile_X1Y10_W1BEG[2] ;
 wire \Tile_X1Y10_W1BEG[3] ;
 wire \Tile_X1Y10_W2BEG[0] ;
 wire \Tile_X1Y10_W2BEG[1] ;
 wire \Tile_X1Y10_W2BEG[2] ;
 wire \Tile_X1Y10_W2BEG[3] ;
 wire \Tile_X1Y10_W2BEG[4] ;
 wire \Tile_X1Y10_W2BEG[5] ;
 wire \Tile_X1Y10_W2BEG[6] ;
 wire \Tile_X1Y10_W2BEG[7] ;
 wire \Tile_X1Y10_W2BEGb[0] ;
 wire \Tile_X1Y10_W2BEGb[1] ;
 wire \Tile_X1Y10_W2BEGb[2] ;
 wire \Tile_X1Y10_W2BEGb[3] ;
 wire \Tile_X1Y10_W2BEGb[4] ;
 wire \Tile_X1Y10_W2BEGb[5] ;
 wire \Tile_X1Y10_W2BEGb[6] ;
 wire \Tile_X1Y10_W2BEGb[7] ;
 wire \Tile_X1Y10_W6BEG[0] ;
 wire \Tile_X1Y10_W6BEG[10] ;
 wire \Tile_X1Y10_W6BEG[11] ;
 wire \Tile_X1Y10_W6BEG[1] ;
 wire \Tile_X1Y10_W6BEG[2] ;
 wire \Tile_X1Y10_W6BEG[3] ;
 wire \Tile_X1Y10_W6BEG[4] ;
 wire \Tile_X1Y10_W6BEG[5] ;
 wire \Tile_X1Y10_W6BEG[6] ;
 wire \Tile_X1Y10_W6BEG[7] ;
 wire \Tile_X1Y10_W6BEG[8] ;
 wire \Tile_X1Y10_W6BEG[9] ;
 wire \Tile_X1Y10_WW4BEG[0] ;
 wire \Tile_X1Y10_WW4BEG[10] ;
 wire \Tile_X1Y10_WW4BEG[11] ;
 wire \Tile_X1Y10_WW4BEG[12] ;
 wire \Tile_X1Y10_WW4BEG[13] ;
 wire \Tile_X1Y10_WW4BEG[14] ;
 wire \Tile_X1Y10_WW4BEG[15] ;
 wire \Tile_X1Y10_WW4BEG[1] ;
 wire \Tile_X1Y10_WW4BEG[2] ;
 wire \Tile_X1Y10_WW4BEG[3] ;
 wire \Tile_X1Y10_WW4BEG[4] ;
 wire \Tile_X1Y10_WW4BEG[5] ;
 wire \Tile_X1Y10_WW4BEG[6] ;
 wire \Tile_X1Y10_WW4BEG[7] ;
 wire \Tile_X1Y10_WW4BEG[8] ;
 wire \Tile_X1Y10_WW4BEG[9] ;
 wire Tile_X1Y11_Co;
 wire \Tile_X1Y11_E1BEG[0] ;
 wire \Tile_X1Y11_E1BEG[1] ;
 wire \Tile_X1Y11_E1BEG[2] ;
 wire \Tile_X1Y11_E1BEG[3] ;
 wire \Tile_X1Y11_E2BEG[0] ;
 wire \Tile_X1Y11_E2BEG[1] ;
 wire \Tile_X1Y11_E2BEG[2] ;
 wire \Tile_X1Y11_E2BEG[3] ;
 wire \Tile_X1Y11_E2BEG[4] ;
 wire \Tile_X1Y11_E2BEG[5] ;
 wire \Tile_X1Y11_E2BEG[6] ;
 wire \Tile_X1Y11_E2BEG[7] ;
 wire \Tile_X1Y11_E2BEGb[0] ;
 wire \Tile_X1Y11_E2BEGb[1] ;
 wire \Tile_X1Y11_E2BEGb[2] ;
 wire \Tile_X1Y11_E2BEGb[3] ;
 wire \Tile_X1Y11_E2BEGb[4] ;
 wire \Tile_X1Y11_E2BEGb[5] ;
 wire \Tile_X1Y11_E2BEGb[6] ;
 wire \Tile_X1Y11_E2BEGb[7] ;
 wire \Tile_X1Y11_E6BEG[0] ;
 wire \Tile_X1Y11_E6BEG[10] ;
 wire \Tile_X1Y11_E6BEG[11] ;
 wire \Tile_X1Y11_E6BEG[1] ;
 wire \Tile_X1Y11_E6BEG[2] ;
 wire \Tile_X1Y11_E6BEG[3] ;
 wire \Tile_X1Y11_E6BEG[4] ;
 wire \Tile_X1Y11_E6BEG[5] ;
 wire \Tile_X1Y11_E6BEG[6] ;
 wire \Tile_X1Y11_E6BEG[7] ;
 wire \Tile_X1Y11_E6BEG[8] ;
 wire \Tile_X1Y11_E6BEG[9] ;
 wire \Tile_X1Y11_EE4BEG[0] ;
 wire \Tile_X1Y11_EE4BEG[10] ;
 wire \Tile_X1Y11_EE4BEG[11] ;
 wire \Tile_X1Y11_EE4BEG[12] ;
 wire \Tile_X1Y11_EE4BEG[13] ;
 wire \Tile_X1Y11_EE4BEG[14] ;
 wire \Tile_X1Y11_EE4BEG[15] ;
 wire \Tile_X1Y11_EE4BEG[1] ;
 wire \Tile_X1Y11_EE4BEG[2] ;
 wire \Tile_X1Y11_EE4BEG[3] ;
 wire \Tile_X1Y11_EE4BEG[4] ;
 wire \Tile_X1Y11_EE4BEG[5] ;
 wire \Tile_X1Y11_EE4BEG[6] ;
 wire \Tile_X1Y11_EE4BEG[7] ;
 wire \Tile_X1Y11_EE4BEG[8] ;
 wire \Tile_X1Y11_EE4BEG[9] ;
 wire \Tile_X1Y11_FrameData_O[0] ;
 wire \Tile_X1Y11_FrameData_O[10] ;
 wire \Tile_X1Y11_FrameData_O[11] ;
 wire \Tile_X1Y11_FrameData_O[12] ;
 wire \Tile_X1Y11_FrameData_O[13] ;
 wire \Tile_X1Y11_FrameData_O[14] ;
 wire \Tile_X1Y11_FrameData_O[15] ;
 wire \Tile_X1Y11_FrameData_O[16] ;
 wire \Tile_X1Y11_FrameData_O[17] ;
 wire \Tile_X1Y11_FrameData_O[18] ;
 wire \Tile_X1Y11_FrameData_O[19] ;
 wire \Tile_X1Y11_FrameData_O[1] ;
 wire \Tile_X1Y11_FrameData_O[20] ;
 wire \Tile_X1Y11_FrameData_O[21] ;
 wire \Tile_X1Y11_FrameData_O[22] ;
 wire \Tile_X1Y11_FrameData_O[23] ;
 wire \Tile_X1Y11_FrameData_O[24] ;
 wire \Tile_X1Y11_FrameData_O[25] ;
 wire \Tile_X1Y11_FrameData_O[26] ;
 wire \Tile_X1Y11_FrameData_O[27] ;
 wire \Tile_X1Y11_FrameData_O[28] ;
 wire \Tile_X1Y11_FrameData_O[29] ;
 wire \Tile_X1Y11_FrameData_O[2] ;
 wire \Tile_X1Y11_FrameData_O[30] ;
 wire \Tile_X1Y11_FrameData_O[31] ;
 wire \Tile_X1Y11_FrameData_O[3] ;
 wire \Tile_X1Y11_FrameData_O[4] ;
 wire \Tile_X1Y11_FrameData_O[5] ;
 wire \Tile_X1Y11_FrameData_O[6] ;
 wire \Tile_X1Y11_FrameData_O[7] ;
 wire \Tile_X1Y11_FrameData_O[8] ;
 wire \Tile_X1Y11_FrameData_O[9] ;
 wire \Tile_X1Y11_FrameStrobe_O[0] ;
 wire \Tile_X1Y11_FrameStrobe_O[10] ;
 wire \Tile_X1Y11_FrameStrobe_O[11] ;
 wire \Tile_X1Y11_FrameStrobe_O[12] ;
 wire \Tile_X1Y11_FrameStrobe_O[13] ;
 wire \Tile_X1Y11_FrameStrobe_O[14] ;
 wire \Tile_X1Y11_FrameStrobe_O[15] ;
 wire \Tile_X1Y11_FrameStrobe_O[16] ;
 wire \Tile_X1Y11_FrameStrobe_O[17] ;
 wire \Tile_X1Y11_FrameStrobe_O[18] ;
 wire \Tile_X1Y11_FrameStrobe_O[19] ;
 wire \Tile_X1Y11_FrameStrobe_O[1] ;
 wire \Tile_X1Y11_FrameStrobe_O[2] ;
 wire \Tile_X1Y11_FrameStrobe_O[3] ;
 wire \Tile_X1Y11_FrameStrobe_O[4] ;
 wire \Tile_X1Y11_FrameStrobe_O[5] ;
 wire \Tile_X1Y11_FrameStrobe_O[6] ;
 wire \Tile_X1Y11_FrameStrobe_O[7] ;
 wire \Tile_X1Y11_FrameStrobe_O[8] ;
 wire \Tile_X1Y11_FrameStrobe_O[9] ;
 wire \Tile_X1Y11_N1BEG[0] ;
 wire \Tile_X1Y11_N1BEG[1] ;
 wire \Tile_X1Y11_N1BEG[2] ;
 wire \Tile_X1Y11_N1BEG[3] ;
 wire \Tile_X1Y11_N2BEG[0] ;
 wire \Tile_X1Y11_N2BEG[1] ;
 wire \Tile_X1Y11_N2BEG[2] ;
 wire \Tile_X1Y11_N2BEG[3] ;
 wire \Tile_X1Y11_N2BEG[4] ;
 wire \Tile_X1Y11_N2BEG[5] ;
 wire \Tile_X1Y11_N2BEG[6] ;
 wire \Tile_X1Y11_N2BEG[7] ;
 wire \Tile_X1Y11_N2BEGb[0] ;
 wire \Tile_X1Y11_N2BEGb[1] ;
 wire \Tile_X1Y11_N2BEGb[2] ;
 wire \Tile_X1Y11_N2BEGb[3] ;
 wire \Tile_X1Y11_N2BEGb[4] ;
 wire \Tile_X1Y11_N2BEGb[5] ;
 wire \Tile_X1Y11_N2BEGb[6] ;
 wire \Tile_X1Y11_N2BEGb[7] ;
 wire \Tile_X1Y11_N4BEG[0] ;
 wire \Tile_X1Y11_N4BEG[10] ;
 wire \Tile_X1Y11_N4BEG[11] ;
 wire \Tile_X1Y11_N4BEG[12] ;
 wire \Tile_X1Y11_N4BEG[13] ;
 wire \Tile_X1Y11_N4BEG[14] ;
 wire \Tile_X1Y11_N4BEG[15] ;
 wire \Tile_X1Y11_N4BEG[1] ;
 wire \Tile_X1Y11_N4BEG[2] ;
 wire \Tile_X1Y11_N4BEG[3] ;
 wire \Tile_X1Y11_N4BEG[4] ;
 wire \Tile_X1Y11_N4BEG[5] ;
 wire \Tile_X1Y11_N4BEG[6] ;
 wire \Tile_X1Y11_N4BEG[7] ;
 wire \Tile_X1Y11_N4BEG[8] ;
 wire \Tile_X1Y11_N4BEG[9] ;
 wire \Tile_X1Y11_NN4BEG[0] ;
 wire \Tile_X1Y11_NN4BEG[10] ;
 wire \Tile_X1Y11_NN4BEG[11] ;
 wire \Tile_X1Y11_NN4BEG[12] ;
 wire \Tile_X1Y11_NN4BEG[13] ;
 wire \Tile_X1Y11_NN4BEG[14] ;
 wire \Tile_X1Y11_NN4BEG[15] ;
 wire \Tile_X1Y11_NN4BEG[1] ;
 wire \Tile_X1Y11_NN4BEG[2] ;
 wire \Tile_X1Y11_NN4BEG[3] ;
 wire \Tile_X1Y11_NN4BEG[4] ;
 wire \Tile_X1Y11_NN4BEG[5] ;
 wire \Tile_X1Y11_NN4BEG[6] ;
 wire \Tile_X1Y11_NN4BEG[7] ;
 wire \Tile_X1Y11_NN4BEG[8] ;
 wire \Tile_X1Y11_NN4BEG[9] ;
 wire \Tile_X1Y11_S1BEG[0] ;
 wire \Tile_X1Y11_S1BEG[1] ;
 wire \Tile_X1Y11_S1BEG[2] ;
 wire \Tile_X1Y11_S1BEG[3] ;
 wire \Tile_X1Y11_S2BEG[0] ;
 wire \Tile_X1Y11_S2BEG[1] ;
 wire \Tile_X1Y11_S2BEG[2] ;
 wire \Tile_X1Y11_S2BEG[3] ;
 wire \Tile_X1Y11_S2BEG[4] ;
 wire \Tile_X1Y11_S2BEG[5] ;
 wire \Tile_X1Y11_S2BEG[6] ;
 wire \Tile_X1Y11_S2BEG[7] ;
 wire \Tile_X1Y11_S2BEGb[0] ;
 wire \Tile_X1Y11_S2BEGb[1] ;
 wire \Tile_X1Y11_S2BEGb[2] ;
 wire \Tile_X1Y11_S2BEGb[3] ;
 wire \Tile_X1Y11_S2BEGb[4] ;
 wire \Tile_X1Y11_S2BEGb[5] ;
 wire \Tile_X1Y11_S2BEGb[6] ;
 wire \Tile_X1Y11_S2BEGb[7] ;
 wire \Tile_X1Y11_S4BEG[0] ;
 wire \Tile_X1Y11_S4BEG[10] ;
 wire \Tile_X1Y11_S4BEG[11] ;
 wire \Tile_X1Y11_S4BEG[12] ;
 wire \Tile_X1Y11_S4BEG[13] ;
 wire \Tile_X1Y11_S4BEG[14] ;
 wire \Tile_X1Y11_S4BEG[15] ;
 wire \Tile_X1Y11_S4BEG[1] ;
 wire \Tile_X1Y11_S4BEG[2] ;
 wire \Tile_X1Y11_S4BEG[3] ;
 wire \Tile_X1Y11_S4BEG[4] ;
 wire \Tile_X1Y11_S4BEG[5] ;
 wire \Tile_X1Y11_S4BEG[6] ;
 wire \Tile_X1Y11_S4BEG[7] ;
 wire \Tile_X1Y11_S4BEG[8] ;
 wire \Tile_X1Y11_S4BEG[9] ;
 wire \Tile_X1Y11_SS4BEG[0] ;
 wire \Tile_X1Y11_SS4BEG[10] ;
 wire \Tile_X1Y11_SS4BEG[11] ;
 wire \Tile_X1Y11_SS4BEG[12] ;
 wire \Tile_X1Y11_SS4BEG[13] ;
 wire \Tile_X1Y11_SS4BEG[14] ;
 wire \Tile_X1Y11_SS4BEG[15] ;
 wire \Tile_X1Y11_SS4BEG[1] ;
 wire \Tile_X1Y11_SS4BEG[2] ;
 wire \Tile_X1Y11_SS4BEG[3] ;
 wire \Tile_X1Y11_SS4BEG[4] ;
 wire \Tile_X1Y11_SS4BEG[5] ;
 wire \Tile_X1Y11_SS4BEG[6] ;
 wire \Tile_X1Y11_SS4BEG[7] ;
 wire \Tile_X1Y11_SS4BEG[8] ;
 wire \Tile_X1Y11_SS4BEG[9] ;
 wire Tile_X1Y11_UserCLKo;
 wire \Tile_X1Y11_W1BEG[0] ;
 wire \Tile_X1Y11_W1BEG[1] ;
 wire \Tile_X1Y11_W1BEG[2] ;
 wire \Tile_X1Y11_W1BEG[3] ;
 wire \Tile_X1Y11_W2BEG[0] ;
 wire \Tile_X1Y11_W2BEG[1] ;
 wire \Tile_X1Y11_W2BEG[2] ;
 wire \Tile_X1Y11_W2BEG[3] ;
 wire \Tile_X1Y11_W2BEG[4] ;
 wire \Tile_X1Y11_W2BEG[5] ;
 wire \Tile_X1Y11_W2BEG[6] ;
 wire \Tile_X1Y11_W2BEG[7] ;
 wire \Tile_X1Y11_W2BEGb[0] ;
 wire \Tile_X1Y11_W2BEGb[1] ;
 wire \Tile_X1Y11_W2BEGb[2] ;
 wire \Tile_X1Y11_W2BEGb[3] ;
 wire \Tile_X1Y11_W2BEGb[4] ;
 wire \Tile_X1Y11_W2BEGb[5] ;
 wire \Tile_X1Y11_W2BEGb[6] ;
 wire \Tile_X1Y11_W2BEGb[7] ;
 wire \Tile_X1Y11_W6BEG[0] ;
 wire \Tile_X1Y11_W6BEG[10] ;
 wire \Tile_X1Y11_W6BEG[11] ;
 wire \Tile_X1Y11_W6BEG[1] ;
 wire \Tile_X1Y11_W6BEG[2] ;
 wire \Tile_X1Y11_W6BEG[3] ;
 wire \Tile_X1Y11_W6BEG[4] ;
 wire \Tile_X1Y11_W6BEG[5] ;
 wire \Tile_X1Y11_W6BEG[6] ;
 wire \Tile_X1Y11_W6BEG[7] ;
 wire \Tile_X1Y11_W6BEG[8] ;
 wire \Tile_X1Y11_W6BEG[9] ;
 wire \Tile_X1Y11_WW4BEG[0] ;
 wire \Tile_X1Y11_WW4BEG[10] ;
 wire \Tile_X1Y11_WW4BEG[11] ;
 wire \Tile_X1Y11_WW4BEG[12] ;
 wire \Tile_X1Y11_WW4BEG[13] ;
 wire \Tile_X1Y11_WW4BEG[14] ;
 wire \Tile_X1Y11_WW4BEG[15] ;
 wire \Tile_X1Y11_WW4BEG[1] ;
 wire \Tile_X1Y11_WW4BEG[2] ;
 wire \Tile_X1Y11_WW4BEG[3] ;
 wire \Tile_X1Y11_WW4BEG[4] ;
 wire \Tile_X1Y11_WW4BEG[5] ;
 wire \Tile_X1Y11_WW4BEG[6] ;
 wire \Tile_X1Y11_WW4BEG[7] ;
 wire \Tile_X1Y11_WW4BEG[8] ;
 wire \Tile_X1Y11_WW4BEG[9] ;
 wire Tile_X1Y12_Co;
 wire \Tile_X1Y12_E1BEG[0] ;
 wire \Tile_X1Y12_E1BEG[1] ;
 wire \Tile_X1Y12_E1BEG[2] ;
 wire \Tile_X1Y12_E1BEG[3] ;
 wire \Tile_X1Y12_E2BEG[0] ;
 wire \Tile_X1Y12_E2BEG[1] ;
 wire \Tile_X1Y12_E2BEG[2] ;
 wire \Tile_X1Y12_E2BEG[3] ;
 wire \Tile_X1Y12_E2BEG[4] ;
 wire \Tile_X1Y12_E2BEG[5] ;
 wire \Tile_X1Y12_E2BEG[6] ;
 wire \Tile_X1Y12_E2BEG[7] ;
 wire \Tile_X1Y12_E2BEGb[0] ;
 wire \Tile_X1Y12_E2BEGb[1] ;
 wire \Tile_X1Y12_E2BEGb[2] ;
 wire \Tile_X1Y12_E2BEGb[3] ;
 wire \Tile_X1Y12_E2BEGb[4] ;
 wire \Tile_X1Y12_E2BEGb[5] ;
 wire \Tile_X1Y12_E2BEGb[6] ;
 wire \Tile_X1Y12_E2BEGb[7] ;
 wire \Tile_X1Y12_E6BEG[0] ;
 wire \Tile_X1Y12_E6BEG[10] ;
 wire \Tile_X1Y12_E6BEG[11] ;
 wire \Tile_X1Y12_E6BEG[1] ;
 wire \Tile_X1Y12_E6BEG[2] ;
 wire \Tile_X1Y12_E6BEG[3] ;
 wire \Tile_X1Y12_E6BEG[4] ;
 wire \Tile_X1Y12_E6BEG[5] ;
 wire \Tile_X1Y12_E6BEG[6] ;
 wire \Tile_X1Y12_E6BEG[7] ;
 wire \Tile_X1Y12_E6BEG[8] ;
 wire \Tile_X1Y12_E6BEG[9] ;
 wire \Tile_X1Y12_EE4BEG[0] ;
 wire \Tile_X1Y12_EE4BEG[10] ;
 wire \Tile_X1Y12_EE4BEG[11] ;
 wire \Tile_X1Y12_EE4BEG[12] ;
 wire \Tile_X1Y12_EE4BEG[13] ;
 wire \Tile_X1Y12_EE4BEG[14] ;
 wire \Tile_X1Y12_EE4BEG[15] ;
 wire \Tile_X1Y12_EE4BEG[1] ;
 wire \Tile_X1Y12_EE4BEG[2] ;
 wire \Tile_X1Y12_EE4BEG[3] ;
 wire \Tile_X1Y12_EE4BEG[4] ;
 wire \Tile_X1Y12_EE4BEG[5] ;
 wire \Tile_X1Y12_EE4BEG[6] ;
 wire \Tile_X1Y12_EE4BEG[7] ;
 wire \Tile_X1Y12_EE4BEG[8] ;
 wire \Tile_X1Y12_EE4BEG[9] ;
 wire \Tile_X1Y12_FrameData_O[0] ;
 wire \Tile_X1Y12_FrameData_O[10] ;
 wire \Tile_X1Y12_FrameData_O[11] ;
 wire \Tile_X1Y12_FrameData_O[12] ;
 wire \Tile_X1Y12_FrameData_O[13] ;
 wire \Tile_X1Y12_FrameData_O[14] ;
 wire \Tile_X1Y12_FrameData_O[15] ;
 wire \Tile_X1Y12_FrameData_O[16] ;
 wire \Tile_X1Y12_FrameData_O[17] ;
 wire \Tile_X1Y12_FrameData_O[18] ;
 wire \Tile_X1Y12_FrameData_O[19] ;
 wire \Tile_X1Y12_FrameData_O[1] ;
 wire \Tile_X1Y12_FrameData_O[20] ;
 wire \Tile_X1Y12_FrameData_O[21] ;
 wire \Tile_X1Y12_FrameData_O[22] ;
 wire \Tile_X1Y12_FrameData_O[23] ;
 wire \Tile_X1Y12_FrameData_O[24] ;
 wire \Tile_X1Y12_FrameData_O[25] ;
 wire \Tile_X1Y12_FrameData_O[26] ;
 wire \Tile_X1Y12_FrameData_O[27] ;
 wire \Tile_X1Y12_FrameData_O[28] ;
 wire \Tile_X1Y12_FrameData_O[29] ;
 wire \Tile_X1Y12_FrameData_O[2] ;
 wire \Tile_X1Y12_FrameData_O[30] ;
 wire \Tile_X1Y12_FrameData_O[31] ;
 wire \Tile_X1Y12_FrameData_O[3] ;
 wire \Tile_X1Y12_FrameData_O[4] ;
 wire \Tile_X1Y12_FrameData_O[5] ;
 wire \Tile_X1Y12_FrameData_O[6] ;
 wire \Tile_X1Y12_FrameData_O[7] ;
 wire \Tile_X1Y12_FrameData_O[8] ;
 wire \Tile_X1Y12_FrameData_O[9] ;
 wire \Tile_X1Y12_FrameStrobe_O[0] ;
 wire \Tile_X1Y12_FrameStrobe_O[10] ;
 wire \Tile_X1Y12_FrameStrobe_O[11] ;
 wire \Tile_X1Y12_FrameStrobe_O[12] ;
 wire \Tile_X1Y12_FrameStrobe_O[13] ;
 wire \Tile_X1Y12_FrameStrobe_O[14] ;
 wire \Tile_X1Y12_FrameStrobe_O[15] ;
 wire \Tile_X1Y12_FrameStrobe_O[16] ;
 wire \Tile_X1Y12_FrameStrobe_O[17] ;
 wire \Tile_X1Y12_FrameStrobe_O[18] ;
 wire \Tile_X1Y12_FrameStrobe_O[19] ;
 wire \Tile_X1Y12_FrameStrobe_O[1] ;
 wire \Tile_X1Y12_FrameStrobe_O[2] ;
 wire \Tile_X1Y12_FrameStrobe_O[3] ;
 wire \Tile_X1Y12_FrameStrobe_O[4] ;
 wire \Tile_X1Y12_FrameStrobe_O[5] ;
 wire \Tile_X1Y12_FrameStrobe_O[6] ;
 wire \Tile_X1Y12_FrameStrobe_O[7] ;
 wire \Tile_X1Y12_FrameStrobe_O[8] ;
 wire \Tile_X1Y12_FrameStrobe_O[9] ;
 wire \Tile_X1Y12_N1BEG[0] ;
 wire \Tile_X1Y12_N1BEG[1] ;
 wire \Tile_X1Y12_N1BEG[2] ;
 wire \Tile_X1Y12_N1BEG[3] ;
 wire \Tile_X1Y12_N2BEG[0] ;
 wire \Tile_X1Y12_N2BEG[1] ;
 wire \Tile_X1Y12_N2BEG[2] ;
 wire \Tile_X1Y12_N2BEG[3] ;
 wire \Tile_X1Y12_N2BEG[4] ;
 wire \Tile_X1Y12_N2BEG[5] ;
 wire \Tile_X1Y12_N2BEG[6] ;
 wire \Tile_X1Y12_N2BEG[7] ;
 wire \Tile_X1Y12_N2BEGb[0] ;
 wire \Tile_X1Y12_N2BEGb[1] ;
 wire \Tile_X1Y12_N2BEGb[2] ;
 wire \Tile_X1Y12_N2BEGb[3] ;
 wire \Tile_X1Y12_N2BEGb[4] ;
 wire \Tile_X1Y12_N2BEGb[5] ;
 wire \Tile_X1Y12_N2BEGb[6] ;
 wire \Tile_X1Y12_N2BEGb[7] ;
 wire \Tile_X1Y12_N4BEG[0] ;
 wire \Tile_X1Y12_N4BEG[10] ;
 wire \Tile_X1Y12_N4BEG[11] ;
 wire \Tile_X1Y12_N4BEG[12] ;
 wire \Tile_X1Y12_N4BEG[13] ;
 wire \Tile_X1Y12_N4BEG[14] ;
 wire \Tile_X1Y12_N4BEG[15] ;
 wire \Tile_X1Y12_N4BEG[1] ;
 wire \Tile_X1Y12_N4BEG[2] ;
 wire \Tile_X1Y12_N4BEG[3] ;
 wire \Tile_X1Y12_N4BEG[4] ;
 wire \Tile_X1Y12_N4BEG[5] ;
 wire \Tile_X1Y12_N4BEG[6] ;
 wire \Tile_X1Y12_N4BEG[7] ;
 wire \Tile_X1Y12_N4BEG[8] ;
 wire \Tile_X1Y12_N4BEG[9] ;
 wire \Tile_X1Y12_NN4BEG[0] ;
 wire \Tile_X1Y12_NN4BEG[10] ;
 wire \Tile_X1Y12_NN4BEG[11] ;
 wire \Tile_X1Y12_NN4BEG[12] ;
 wire \Tile_X1Y12_NN4BEG[13] ;
 wire \Tile_X1Y12_NN4BEG[14] ;
 wire \Tile_X1Y12_NN4BEG[15] ;
 wire \Tile_X1Y12_NN4BEG[1] ;
 wire \Tile_X1Y12_NN4BEG[2] ;
 wire \Tile_X1Y12_NN4BEG[3] ;
 wire \Tile_X1Y12_NN4BEG[4] ;
 wire \Tile_X1Y12_NN4BEG[5] ;
 wire \Tile_X1Y12_NN4BEG[6] ;
 wire \Tile_X1Y12_NN4BEG[7] ;
 wire \Tile_X1Y12_NN4BEG[8] ;
 wire \Tile_X1Y12_NN4BEG[9] ;
 wire \Tile_X1Y12_S1BEG[0] ;
 wire \Tile_X1Y12_S1BEG[1] ;
 wire \Tile_X1Y12_S1BEG[2] ;
 wire \Tile_X1Y12_S1BEG[3] ;
 wire \Tile_X1Y12_S2BEG[0] ;
 wire \Tile_X1Y12_S2BEG[1] ;
 wire \Tile_X1Y12_S2BEG[2] ;
 wire \Tile_X1Y12_S2BEG[3] ;
 wire \Tile_X1Y12_S2BEG[4] ;
 wire \Tile_X1Y12_S2BEG[5] ;
 wire \Tile_X1Y12_S2BEG[6] ;
 wire \Tile_X1Y12_S2BEG[7] ;
 wire \Tile_X1Y12_S2BEGb[0] ;
 wire \Tile_X1Y12_S2BEGb[1] ;
 wire \Tile_X1Y12_S2BEGb[2] ;
 wire \Tile_X1Y12_S2BEGb[3] ;
 wire \Tile_X1Y12_S2BEGb[4] ;
 wire \Tile_X1Y12_S2BEGb[5] ;
 wire \Tile_X1Y12_S2BEGb[6] ;
 wire \Tile_X1Y12_S2BEGb[7] ;
 wire \Tile_X1Y12_S4BEG[0] ;
 wire \Tile_X1Y12_S4BEG[10] ;
 wire \Tile_X1Y12_S4BEG[11] ;
 wire \Tile_X1Y12_S4BEG[12] ;
 wire \Tile_X1Y12_S4BEG[13] ;
 wire \Tile_X1Y12_S4BEG[14] ;
 wire \Tile_X1Y12_S4BEG[15] ;
 wire \Tile_X1Y12_S4BEG[1] ;
 wire \Tile_X1Y12_S4BEG[2] ;
 wire \Tile_X1Y12_S4BEG[3] ;
 wire \Tile_X1Y12_S4BEG[4] ;
 wire \Tile_X1Y12_S4BEG[5] ;
 wire \Tile_X1Y12_S4BEG[6] ;
 wire \Tile_X1Y12_S4BEG[7] ;
 wire \Tile_X1Y12_S4BEG[8] ;
 wire \Tile_X1Y12_S4BEG[9] ;
 wire \Tile_X1Y12_SS4BEG[0] ;
 wire \Tile_X1Y12_SS4BEG[10] ;
 wire \Tile_X1Y12_SS4BEG[11] ;
 wire \Tile_X1Y12_SS4BEG[12] ;
 wire \Tile_X1Y12_SS4BEG[13] ;
 wire \Tile_X1Y12_SS4BEG[14] ;
 wire \Tile_X1Y12_SS4BEG[15] ;
 wire \Tile_X1Y12_SS4BEG[1] ;
 wire \Tile_X1Y12_SS4BEG[2] ;
 wire \Tile_X1Y12_SS4BEG[3] ;
 wire \Tile_X1Y12_SS4BEG[4] ;
 wire \Tile_X1Y12_SS4BEG[5] ;
 wire \Tile_X1Y12_SS4BEG[6] ;
 wire \Tile_X1Y12_SS4BEG[7] ;
 wire \Tile_X1Y12_SS4BEG[8] ;
 wire \Tile_X1Y12_SS4BEG[9] ;
 wire Tile_X1Y12_UserCLKo;
 wire \Tile_X1Y12_W1BEG[0] ;
 wire \Tile_X1Y12_W1BEG[1] ;
 wire \Tile_X1Y12_W1BEG[2] ;
 wire \Tile_X1Y12_W1BEG[3] ;
 wire \Tile_X1Y12_W2BEG[0] ;
 wire \Tile_X1Y12_W2BEG[1] ;
 wire \Tile_X1Y12_W2BEG[2] ;
 wire \Tile_X1Y12_W2BEG[3] ;
 wire \Tile_X1Y12_W2BEG[4] ;
 wire \Tile_X1Y12_W2BEG[5] ;
 wire \Tile_X1Y12_W2BEG[6] ;
 wire \Tile_X1Y12_W2BEG[7] ;
 wire \Tile_X1Y12_W2BEGb[0] ;
 wire \Tile_X1Y12_W2BEGb[1] ;
 wire \Tile_X1Y12_W2BEGb[2] ;
 wire \Tile_X1Y12_W2BEGb[3] ;
 wire \Tile_X1Y12_W2BEGb[4] ;
 wire \Tile_X1Y12_W2BEGb[5] ;
 wire \Tile_X1Y12_W2BEGb[6] ;
 wire \Tile_X1Y12_W2BEGb[7] ;
 wire \Tile_X1Y12_W6BEG[0] ;
 wire \Tile_X1Y12_W6BEG[10] ;
 wire \Tile_X1Y12_W6BEG[11] ;
 wire \Tile_X1Y12_W6BEG[1] ;
 wire \Tile_X1Y12_W6BEG[2] ;
 wire \Tile_X1Y12_W6BEG[3] ;
 wire \Tile_X1Y12_W6BEG[4] ;
 wire \Tile_X1Y12_W6BEG[5] ;
 wire \Tile_X1Y12_W6BEG[6] ;
 wire \Tile_X1Y12_W6BEG[7] ;
 wire \Tile_X1Y12_W6BEG[8] ;
 wire \Tile_X1Y12_W6BEG[9] ;
 wire \Tile_X1Y12_WW4BEG[0] ;
 wire \Tile_X1Y12_WW4BEG[10] ;
 wire \Tile_X1Y12_WW4BEG[11] ;
 wire \Tile_X1Y12_WW4BEG[12] ;
 wire \Tile_X1Y12_WW4BEG[13] ;
 wire \Tile_X1Y12_WW4BEG[14] ;
 wire \Tile_X1Y12_WW4BEG[15] ;
 wire \Tile_X1Y12_WW4BEG[1] ;
 wire \Tile_X1Y12_WW4BEG[2] ;
 wire \Tile_X1Y12_WW4BEG[3] ;
 wire \Tile_X1Y12_WW4BEG[4] ;
 wire \Tile_X1Y12_WW4BEG[5] ;
 wire \Tile_X1Y12_WW4BEG[6] ;
 wire \Tile_X1Y12_WW4BEG[7] ;
 wire \Tile_X1Y12_WW4BEG[8] ;
 wire \Tile_X1Y12_WW4BEG[9] ;
 wire Tile_X1Y13_Co;
 wire \Tile_X1Y13_E1BEG[0] ;
 wire \Tile_X1Y13_E1BEG[1] ;
 wire \Tile_X1Y13_E1BEG[2] ;
 wire \Tile_X1Y13_E1BEG[3] ;
 wire \Tile_X1Y13_E2BEG[0] ;
 wire \Tile_X1Y13_E2BEG[1] ;
 wire \Tile_X1Y13_E2BEG[2] ;
 wire \Tile_X1Y13_E2BEG[3] ;
 wire \Tile_X1Y13_E2BEG[4] ;
 wire \Tile_X1Y13_E2BEG[5] ;
 wire \Tile_X1Y13_E2BEG[6] ;
 wire \Tile_X1Y13_E2BEG[7] ;
 wire \Tile_X1Y13_E2BEGb[0] ;
 wire \Tile_X1Y13_E2BEGb[1] ;
 wire \Tile_X1Y13_E2BEGb[2] ;
 wire \Tile_X1Y13_E2BEGb[3] ;
 wire \Tile_X1Y13_E2BEGb[4] ;
 wire \Tile_X1Y13_E2BEGb[5] ;
 wire \Tile_X1Y13_E2BEGb[6] ;
 wire \Tile_X1Y13_E2BEGb[7] ;
 wire \Tile_X1Y13_E6BEG[0] ;
 wire \Tile_X1Y13_E6BEG[10] ;
 wire \Tile_X1Y13_E6BEG[11] ;
 wire \Tile_X1Y13_E6BEG[1] ;
 wire \Tile_X1Y13_E6BEG[2] ;
 wire \Tile_X1Y13_E6BEG[3] ;
 wire \Tile_X1Y13_E6BEG[4] ;
 wire \Tile_X1Y13_E6BEG[5] ;
 wire \Tile_X1Y13_E6BEG[6] ;
 wire \Tile_X1Y13_E6BEG[7] ;
 wire \Tile_X1Y13_E6BEG[8] ;
 wire \Tile_X1Y13_E6BEG[9] ;
 wire \Tile_X1Y13_EE4BEG[0] ;
 wire \Tile_X1Y13_EE4BEG[10] ;
 wire \Tile_X1Y13_EE4BEG[11] ;
 wire \Tile_X1Y13_EE4BEG[12] ;
 wire \Tile_X1Y13_EE4BEG[13] ;
 wire \Tile_X1Y13_EE4BEG[14] ;
 wire \Tile_X1Y13_EE4BEG[15] ;
 wire \Tile_X1Y13_EE4BEG[1] ;
 wire \Tile_X1Y13_EE4BEG[2] ;
 wire \Tile_X1Y13_EE4BEG[3] ;
 wire \Tile_X1Y13_EE4BEG[4] ;
 wire \Tile_X1Y13_EE4BEG[5] ;
 wire \Tile_X1Y13_EE4BEG[6] ;
 wire \Tile_X1Y13_EE4BEG[7] ;
 wire \Tile_X1Y13_EE4BEG[8] ;
 wire \Tile_X1Y13_EE4BEG[9] ;
 wire \Tile_X1Y13_FrameData_O[0] ;
 wire \Tile_X1Y13_FrameData_O[10] ;
 wire \Tile_X1Y13_FrameData_O[11] ;
 wire \Tile_X1Y13_FrameData_O[12] ;
 wire \Tile_X1Y13_FrameData_O[13] ;
 wire \Tile_X1Y13_FrameData_O[14] ;
 wire \Tile_X1Y13_FrameData_O[15] ;
 wire \Tile_X1Y13_FrameData_O[16] ;
 wire \Tile_X1Y13_FrameData_O[17] ;
 wire \Tile_X1Y13_FrameData_O[18] ;
 wire \Tile_X1Y13_FrameData_O[19] ;
 wire \Tile_X1Y13_FrameData_O[1] ;
 wire \Tile_X1Y13_FrameData_O[20] ;
 wire \Tile_X1Y13_FrameData_O[21] ;
 wire \Tile_X1Y13_FrameData_O[22] ;
 wire \Tile_X1Y13_FrameData_O[23] ;
 wire \Tile_X1Y13_FrameData_O[24] ;
 wire \Tile_X1Y13_FrameData_O[25] ;
 wire \Tile_X1Y13_FrameData_O[26] ;
 wire \Tile_X1Y13_FrameData_O[27] ;
 wire \Tile_X1Y13_FrameData_O[28] ;
 wire \Tile_X1Y13_FrameData_O[29] ;
 wire \Tile_X1Y13_FrameData_O[2] ;
 wire \Tile_X1Y13_FrameData_O[30] ;
 wire \Tile_X1Y13_FrameData_O[31] ;
 wire \Tile_X1Y13_FrameData_O[3] ;
 wire \Tile_X1Y13_FrameData_O[4] ;
 wire \Tile_X1Y13_FrameData_O[5] ;
 wire \Tile_X1Y13_FrameData_O[6] ;
 wire \Tile_X1Y13_FrameData_O[7] ;
 wire \Tile_X1Y13_FrameData_O[8] ;
 wire \Tile_X1Y13_FrameData_O[9] ;
 wire \Tile_X1Y13_FrameStrobe_O[0] ;
 wire \Tile_X1Y13_FrameStrobe_O[10] ;
 wire \Tile_X1Y13_FrameStrobe_O[11] ;
 wire \Tile_X1Y13_FrameStrobe_O[12] ;
 wire \Tile_X1Y13_FrameStrobe_O[13] ;
 wire \Tile_X1Y13_FrameStrobe_O[14] ;
 wire \Tile_X1Y13_FrameStrobe_O[15] ;
 wire \Tile_X1Y13_FrameStrobe_O[16] ;
 wire \Tile_X1Y13_FrameStrobe_O[17] ;
 wire \Tile_X1Y13_FrameStrobe_O[18] ;
 wire \Tile_X1Y13_FrameStrobe_O[19] ;
 wire \Tile_X1Y13_FrameStrobe_O[1] ;
 wire \Tile_X1Y13_FrameStrobe_O[2] ;
 wire \Tile_X1Y13_FrameStrobe_O[3] ;
 wire \Tile_X1Y13_FrameStrobe_O[4] ;
 wire \Tile_X1Y13_FrameStrobe_O[5] ;
 wire \Tile_X1Y13_FrameStrobe_O[6] ;
 wire \Tile_X1Y13_FrameStrobe_O[7] ;
 wire \Tile_X1Y13_FrameStrobe_O[8] ;
 wire \Tile_X1Y13_FrameStrobe_O[9] ;
 wire \Tile_X1Y13_N1BEG[0] ;
 wire \Tile_X1Y13_N1BEG[1] ;
 wire \Tile_X1Y13_N1BEG[2] ;
 wire \Tile_X1Y13_N1BEG[3] ;
 wire \Tile_X1Y13_N2BEG[0] ;
 wire \Tile_X1Y13_N2BEG[1] ;
 wire \Tile_X1Y13_N2BEG[2] ;
 wire \Tile_X1Y13_N2BEG[3] ;
 wire \Tile_X1Y13_N2BEG[4] ;
 wire \Tile_X1Y13_N2BEG[5] ;
 wire \Tile_X1Y13_N2BEG[6] ;
 wire \Tile_X1Y13_N2BEG[7] ;
 wire \Tile_X1Y13_N2BEGb[0] ;
 wire \Tile_X1Y13_N2BEGb[1] ;
 wire \Tile_X1Y13_N2BEGb[2] ;
 wire \Tile_X1Y13_N2BEGb[3] ;
 wire \Tile_X1Y13_N2BEGb[4] ;
 wire \Tile_X1Y13_N2BEGb[5] ;
 wire \Tile_X1Y13_N2BEGb[6] ;
 wire \Tile_X1Y13_N2BEGb[7] ;
 wire \Tile_X1Y13_N4BEG[0] ;
 wire \Tile_X1Y13_N4BEG[10] ;
 wire \Tile_X1Y13_N4BEG[11] ;
 wire \Tile_X1Y13_N4BEG[12] ;
 wire \Tile_X1Y13_N4BEG[13] ;
 wire \Tile_X1Y13_N4BEG[14] ;
 wire \Tile_X1Y13_N4BEG[15] ;
 wire \Tile_X1Y13_N4BEG[1] ;
 wire \Tile_X1Y13_N4BEG[2] ;
 wire \Tile_X1Y13_N4BEG[3] ;
 wire \Tile_X1Y13_N4BEG[4] ;
 wire \Tile_X1Y13_N4BEG[5] ;
 wire \Tile_X1Y13_N4BEG[6] ;
 wire \Tile_X1Y13_N4BEG[7] ;
 wire \Tile_X1Y13_N4BEG[8] ;
 wire \Tile_X1Y13_N4BEG[9] ;
 wire \Tile_X1Y13_NN4BEG[0] ;
 wire \Tile_X1Y13_NN4BEG[10] ;
 wire \Tile_X1Y13_NN4BEG[11] ;
 wire \Tile_X1Y13_NN4BEG[12] ;
 wire \Tile_X1Y13_NN4BEG[13] ;
 wire \Tile_X1Y13_NN4BEG[14] ;
 wire \Tile_X1Y13_NN4BEG[15] ;
 wire \Tile_X1Y13_NN4BEG[1] ;
 wire \Tile_X1Y13_NN4BEG[2] ;
 wire \Tile_X1Y13_NN4BEG[3] ;
 wire \Tile_X1Y13_NN4BEG[4] ;
 wire \Tile_X1Y13_NN4BEG[5] ;
 wire \Tile_X1Y13_NN4BEG[6] ;
 wire \Tile_X1Y13_NN4BEG[7] ;
 wire \Tile_X1Y13_NN4BEG[8] ;
 wire \Tile_X1Y13_NN4BEG[9] ;
 wire \Tile_X1Y13_S1BEG[0] ;
 wire \Tile_X1Y13_S1BEG[1] ;
 wire \Tile_X1Y13_S1BEG[2] ;
 wire \Tile_X1Y13_S1BEG[3] ;
 wire \Tile_X1Y13_S2BEG[0] ;
 wire \Tile_X1Y13_S2BEG[1] ;
 wire \Tile_X1Y13_S2BEG[2] ;
 wire \Tile_X1Y13_S2BEG[3] ;
 wire \Tile_X1Y13_S2BEG[4] ;
 wire \Tile_X1Y13_S2BEG[5] ;
 wire \Tile_X1Y13_S2BEG[6] ;
 wire \Tile_X1Y13_S2BEG[7] ;
 wire \Tile_X1Y13_S2BEGb[0] ;
 wire \Tile_X1Y13_S2BEGb[1] ;
 wire \Tile_X1Y13_S2BEGb[2] ;
 wire \Tile_X1Y13_S2BEGb[3] ;
 wire \Tile_X1Y13_S2BEGb[4] ;
 wire \Tile_X1Y13_S2BEGb[5] ;
 wire \Tile_X1Y13_S2BEGb[6] ;
 wire \Tile_X1Y13_S2BEGb[7] ;
 wire \Tile_X1Y13_S4BEG[0] ;
 wire \Tile_X1Y13_S4BEG[10] ;
 wire \Tile_X1Y13_S4BEG[11] ;
 wire \Tile_X1Y13_S4BEG[12] ;
 wire \Tile_X1Y13_S4BEG[13] ;
 wire \Tile_X1Y13_S4BEG[14] ;
 wire \Tile_X1Y13_S4BEG[15] ;
 wire \Tile_X1Y13_S4BEG[1] ;
 wire \Tile_X1Y13_S4BEG[2] ;
 wire \Tile_X1Y13_S4BEG[3] ;
 wire \Tile_X1Y13_S4BEG[4] ;
 wire \Tile_X1Y13_S4BEG[5] ;
 wire \Tile_X1Y13_S4BEG[6] ;
 wire \Tile_X1Y13_S4BEG[7] ;
 wire \Tile_X1Y13_S4BEG[8] ;
 wire \Tile_X1Y13_S4BEG[9] ;
 wire \Tile_X1Y13_SS4BEG[0] ;
 wire \Tile_X1Y13_SS4BEG[10] ;
 wire \Tile_X1Y13_SS4BEG[11] ;
 wire \Tile_X1Y13_SS4BEG[12] ;
 wire \Tile_X1Y13_SS4BEG[13] ;
 wire \Tile_X1Y13_SS4BEG[14] ;
 wire \Tile_X1Y13_SS4BEG[15] ;
 wire \Tile_X1Y13_SS4BEG[1] ;
 wire \Tile_X1Y13_SS4BEG[2] ;
 wire \Tile_X1Y13_SS4BEG[3] ;
 wire \Tile_X1Y13_SS4BEG[4] ;
 wire \Tile_X1Y13_SS4BEG[5] ;
 wire \Tile_X1Y13_SS4BEG[6] ;
 wire \Tile_X1Y13_SS4BEG[7] ;
 wire \Tile_X1Y13_SS4BEG[8] ;
 wire \Tile_X1Y13_SS4BEG[9] ;
 wire Tile_X1Y13_UserCLKo;
 wire \Tile_X1Y13_W1BEG[0] ;
 wire \Tile_X1Y13_W1BEG[1] ;
 wire \Tile_X1Y13_W1BEG[2] ;
 wire \Tile_X1Y13_W1BEG[3] ;
 wire \Tile_X1Y13_W2BEG[0] ;
 wire \Tile_X1Y13_W2BEG[1] ;
 wire \Tile_X1Y13_W2BEG[2] ;
 wire \Tile_X1Y13_W2BEG[3] ;
 wire \Tile_X1Y13_W2BEG[4] ;
 wire \Tile_X1Y13_W2BEG[5] ;
 wire \Tile_X1Y13_W2BEG[6] ;
 wire \Tile_X1Y13_W2BEG[7] ;
 wire \Tile_X1Y13_W2BEGb[0] ;
 wire \Tile_X1Y13_W2BEGb[1] ;
 wire \Tile_X1Y13_W2BEGb[2] ;
 wire \Tile_X1Y13_W2BEGb[3] ;
 wire \Tile_X1Y13_W2BEGb[4] ;
 wire \Tile_X1Y13_W2BEGb[5] ;
 wire \Tile_X1Y13_W2BEGb[6] ;
 wire \Tile_X1Y13_W2BEGb[7] ;
 wire \Tile_X1Y13_W6BEG[0] ;
 wire \Tile_X1Y13_W6BEG[10] ;
 wire \Tile_X1Y13_W6BEG[11] ;
 wire \Tile_X1Y13_W6BEG[1] ;
 wire \Tile_X1Y13_W6BEG[2] ;
 wire \Tile_X1Y13_W6BEG[3] ;
 wire \Tile_X1Y13_W6BEG[4] ;
 wire \Tile_X1Y13_W6BEG[5] ;
 wire \Tile_X1Y13_W6BEG[6] ;
 wire \Tile_X1Y13_W6BEG[7] ;
 wire \Tile_X1Y13_W6BEG[8] ;
 wire \Tile_X1Y13_W6BEG[9] ;
 wire \Tile_X1Y13_WW4BEG[0] ;
 wire \Tile_X1Y13_WW4BEG[10] ;
 wire \Tile_X1Y13_WW4BEG[11] ;
 wire \Tile_X1Y13_WW4BEG[12] ;
 wire \Tile_X1Y13_WW4BEG[13] ;
 wire \Tile_X1Y13_WW4BEG[14] ;
 wire \Tile_X1Y13_WW4BEG[15] ;
 wire \Tile_X1Y13_WW4BEG[1] ;
 wire \Tile_X1Y13_WW4BEG[2] ;
 wire \Tile_X1Y13_WW4BEG[3] ;
 wire \Tile_X1Y13_WW4BEG[4] ;
 wire \Tile_X1Y13_WW4BEG[5] ;
 wire \Tile_X1Y13_WW4BEG[6] ;
 wire \Tile_X1Y13_WW4BEG[7] ;
 wire \Tile_X1Y13_WW4BEG[8] ;
 wire \Tile_X1Y13_WW4BEG[9] ;
 wire Tile_X1Y14_Co;
 wire \Tile_X1Y14_E1BEG[0] ;
 wire \Tile_X1Y14_E1BEG[1] ;
 wire \Tile_X1Y14_E1BEG[2] ;
 wire \Tile_X1Y14_E1BEG[3] ;
 wire \Tile_X1Y14_E2BEG[0] ;
 wire \Tile_X1Y14_E2BEG[1] ;
 wire \Tile_X1Y14_E2BEG[2] ;
 wire \Tile_X1Y14_E2BEG[3] ;
 wire \Tile_X1Y14_E2BEG[4] ;
 wire \Tile_X1Y14_E2BEG[5] ;
 wire \Tile_X1Y14_E2BEG[6] ;
 wire \Tile_X1Y14_E2BEG[7] ;
 wire \Tile_X1Y14_E2BEGb[0] ;
 wire \Tile_X1Y14_E2BEGb[1] ;
 wire \Tile_X1Y14_E2BEGb[2] ;
 wire \Tile_X1Y14_E2BEGb[3] ;
 wire \Tile_X1Y14_E2BEGb[4] ;
 wire \Tile_X1Y14_E2BEGb[5] ;
 wire \Tile_X1Y14_E2BEGb[6] ;
 wire \Tile_X1Y14_E2BEGb[7] ;
 wire \Tile_X1Y14_E6BEG[0] ;
 wire \Tile_X1Y14_E6BEG[10] ;
 wire \Tile_X1Y14_E6BEG[11] ;
 wire \Tile_X1Y14_E6BEG[1] ;
 wire \Tile_X1Y14_E6BEG[2] ;
 wire \Tile_X1Y14_E6BEG[3] ;
 wire \Tile_X1Y14_E6BEG[4] ;
 wire \Tile_X1Y14_E6BEG[5] ;
 wire \Tile_X1Y14_E6BEG[6] ;
 wire \Tile_X1Y14_E6BEG[7] ;
 wire \Tile_X1Y14_E6BEG[8] ;
 wire \Tile_X1Y14_E6BEG[9] ;
 wire \Tile_X1Y14_EE4BEG[0] ;
 wire \Tile_X1Y14_EE4BEG[10] ;
 wire \Tile_X1Y14_EE4BEG[11] ;
 wire \Tile_X1Y14_EE4BEG[12] ;
 wire \Tile_X1Y14_EE4BEG[13] ;
 wire \Tile_X1Y14_EE4BEG[14] ;
 wire \Tile_X1Y14_EE4BEG[15] ;
 wire \Tile_X1Y14_EE4BEG[1] ;
 wire \Tile_X1Y14_EE4BEG[2] ;
 wire \Tile_X1Y14_EE4BEG[3] ;
 wire \Tile_X1Y14_EE4BEG[4] ;
 wire \Tile_X1Y14_EE4BEG[5] ;
 wire \Tile_X1Y14_EE4BEG[6] ;
 wire \Tile_X1Y14_EE4BEG[7] ;
 wire \Tile_X1Y14_EE4BEG[8] ;
 wire \Tile_X1Y14_EE4BEG[9] ;
 wire \Tile_X1Y14_FrameData_O[0] ;
 wire \Tile_X1Y14_FrameData_O[10] ;
 wire \Tile_X1Y14_FrameData_O[11] ;
 wire \Tile_X1Y14_FrameData_O[12] ;
 wire \Tile_X1Y14_FrameData_O[13] ;
 wire \Tile_X1Y14_FrameData_O[14] ;
 wire \Tile_X1Y14_FrameData_O[15] ;
 wire \Tile_X1Y14_FrameData_O[16] ;
 wire \Tile_X1Y14_FrameData_O[17] ;
 wire \Tile_X1Y14_FrameData_O[18] ;
 wire \Tile_X1Y14_FrameData_O[19] ;
 wire \Tile_X1Y14_FrameData_O[1] ;
 wire \Tile_X1Y14_FrameData_O[20] ;
 wire \Tile_X1Y14_FrameData_O[21] ;
 wire \Tile_X1Y14_FrameData_O[22] ;
 wire \Tile_X1Y14_FrameData_O[23] ;
 wire \Tile_X1Y14_FrameData_O[24] ;
 wire \Tile_X1Y14_FrameData_O[25] ;
 wire \Tile_X1Y14_FrameData_O[26] ;
 wire \Tile_X1Y14_FrameData_O[27] ;
 wire \Tile_X1Y14_FrameData_O[28] ;
 wire \Tile_X1Y14_FrameData_O[29] ;
 wire \Tile_X1Y14_FrameData_O[2] ;
 wire \Tile_X1Y14_FrameData_O[30] ;
 wire \Tile_X1Y14_FrameData_O[31] ;
 wire \Tile_X1Y14_FrameData_O[3] ;
 wire \Tile_X1Y14_FrameData_O[4] ;
 wire \Tile_X1Y14_FrameData_O[5] ;
 wire \Tile_X1Y14_FrameData_O[6] ;
 wire \Tile_X1Y14_FrameData_O[7] ;
 wire \Tile_X1Y14_FrameData_O[8] ;
 wire \Tile_X1Y14_FrameData_O[9] ;
 wire \Tile_X1Y14_FrameStrobe_O[0] ;
 wire \Tile_X1Y14_FrameStrobe_O[10] ;
 wire \Tile_X1Y14_FrameStrobe_O[11] ;
 wire \Tile_X1Y14_FrameStrobe_O[12] ;
 wire \Tile_X1Y14_FrameStrobe_O[13] ;
 wire \Tile_X1Y14_FrameStrobe_O[14] ;
 wire \Tile_X1Y14_FrameStrobe_O[15] ;
 wire \Tile_X1Y14_FrameStrobe_O[16] ;
 wire \Tile_X1Y14_FrameStrobe_O[17] ;
 wire \Tile_X1Y14_FrameStrobe_O[18] ;
 wire \Tile_X1Y14_FrameStrobe_O[19] ;
 wire \Tile_X1Y14_FrameStrobe_O[1] ;
 wire \Tile_X1Y14_FrameStrobe_O[2] ;
 wire \Tile_X1Y14_FrameStrobe_O[3] ;
 wire \Tile_X1Y14_FrameStrobe_O[4] ;
 wire \Tile_X1Y14_FrameStrobe_O[5] ;
 wire \Tile_X1Y14_FrameStrobe_O[6] ;
 wire \Tile_X1Y14_FrameStrobe_O[7] ;
 wire \Tile_X1Y14_FrameStrobe_O[8] ;
 wire \Tile_X1Y14_FrameStrobe_O[9] ;
 wire \Tile_X1Y14_N1BEG[0] ;
 wire \Tile_X1Y14_N1BEG[1] ;
 wire \Tile_X1Y14_N1BEG[2] ;
 wire \Tile_X1Y14_N1BEG[3] ;
 wire \Tile_X1Y14_N2BEG[0] ;
 wire \Tile_X1Y14_N2BEG[1] ;
 wire \Tile_X1Y14_N2BEG[2] ;
 wire \Tile_X1Y14_N2BEG[3] ;
 wire \Tile_X1Y14_N2BEG[4] ;
 wire \Tile_X1Y14_N2BEG[5] ;
 wire \Tile_X1Y14_N2BEG[6] ;
 wire \Tile_X1Y14_N2BEG[7] ;
 wire \Tile_X1Y14_N2BEGb[0] ;
 wire \Tile_X1Y14_N2BEGb[1] ;
 wire \Tile_X1Y14_N2BEGb[2] ;
 wire \Tile_X1Y14_N2BEGb[3] ;
 wire \Tile_X1Y14_N2BEGb[4] ;
 wire \Tile_X1Y14_N2BEGb[5] ;
 wire \Tile_X1Y14_N2BEGb[6] ;
 wire \Tile_X1Y14_N2BEGb[7] ;
 wire \Tile_X1Y14_N4BEG[0] ;
 wire \Tile_X1Y14_N4BEG[10] ;
 wire \Tile_X1Y14_N4BEG[11] ;
 wire \Tile_X1Y14_N4BEG[12] ;
 wire \Tile_X1Y14_N4BEG[13] ;
 wire \Tile_X1Y14_N4BEG[14] ;
 wire \Tile_X1Y14_N4BEG[15] ;
 wire \Tile_X1Y14_N4BEG[1] ;
 wire \Tile_X1Y14_N4BEG[2] ;
 wire \Tile_X1Y14_N4BEG[3] ;
 wire \Tile_X1Y14_N4BEG[4] ;
 wire \Tile_X1Y14_N4BEG[5] ;
 wire \Tile_X1Y14_N4BEG[6] ;
 wire \Tile_X1Y14_N4BEG[7] ;
 wire \Tile_X1Y14_N4BEG[8] ;
 wire \Tile_X1Y14_N4BEG[9] ;
 wire \Tile_X1Y14_NN4BEG[0] ;
 wire \Tile_X1Y14_NN4BEG[10] ;
 wire \Tile_X1Y14_NN4BEG[11] ;
 wire \Tile_X1Y14_NN4BEG[12] ;
 wire \Tile_X1Y14_NN4BEG[13] ;
 wire \Tile_X1Y14_NN4BEG[14] ;
 wire \Tile_X1Y14_NN4BEG[15] ;
 wire \Tile_X1Y14_NN4BEG[1] ;
 wire \Tile_X1Y14_NN4BEG[2] ;
 wire \Tile_X1Y14_NN4BEG[3] ;
 wire \Tile_X1Y14_NN4BEG[4] ;
 wire \Tile_X1Y14_NN4BEG[5] ;
 wire \Tile_X1Y14_NN4BEG[6] ;
 wire \Tile_X1Y14_NN4BEG[7] ;
 wire \Tile_X1Y14_NN4BEG[8] ;
 wire \Tile_X1Y14_NN4BEG[9] ;
 wire \Tile_X1Y14_S1BEG[0] ;
 wire \Tile_X1Y14_S1BEG[1] ;
 wire \Tile_X1Y14_S1BEG[2] ;
 wire \Tile_X1Y14_S1BEG[3] ;
 wire \Tile_X1Y14_S2BEG[0] ;
 wire \Tile_X1Y14_S2BEG[1] ;
 wire \Tile_X1Y14_S2BEG[2] ;
 wire \Tile_X1Y14_S2BEG[3] ;
 wire \Tile_X1Y14_S2BEG[4] ;
 wire \Tile_X1Y14_S2BEG[5] ;
 wire \Tile_X1Y14_S2BEG[6] ;
 wire \Tile_X1Y14_S2BEG[7] ;
 wire \Tile_X1Y14_S2BEGb[0] ;
 wire \Tile_X1Y14_S2BEGb[1] ;
 wire \Tile_X1Y14_S2BEGb[2] ;
 wire \Tile_X1Y14_S2BEGb[3] ;
 wire \Tile_X1Y14_S2BEGb[4] ;
 wire \Tile_X1Y14_S2BEGb[5] ;
 wire \Tile_X1Y14_S2BEGb[6] ;
 wire \Tile_X1Y14_S2BEGb[7] ;
 wire \Tile_X1Y14_S4BEG[0] ;
 wire \Tile_X1Y14_S4BEG[10] ;
 wire \Tile_X1Y14_S4BEG[11] ;
 wire \Tile_X1Y14_S4BEG[12] ;
 wire \Tile_X1Y14_S4BEG[13] ;
 wire \Tile_X1Y14_S4BEG[14] ;
 wire \Tile_X1Y14_S4BEG[15] ;
 wire \Tile_X1Y14_S4BEG[1] ;
 wire \Tile_X1Y14_S4BEG[2] ;
 wire \Tile_X1Y14_S4BEG[3] ;
 wire \Tile_X1Y14_S4BEG[4] ;
 wire \Tile_X1Y14_S4BEG[5] ;
 wire \Tile_X1Y14_S4BEG[6] ;
 wire \Tile_X1Y14_S4BEG[7] ;
 wire \Tile_X1Y14_S4BEG[8] ;
 wire \Tile_X1Y14_S4BEG[9] ;
 wire \Tile_X1Y14_SS4BEG[0] ;
 wire \Tile_X1Y14_SS4BEG[10] ;
 wire \Tile_X1Y14_SS4BEG[11] ;
 wire \Tile_X1Y14_SS4BEG[12] ;
 wire \Tile_X1Y14_SS4BEG[13] ;
 wire \Tile_X1Y14_SS4BEG[14] ;
 wire \Tile_X1Y14_SS4BEG[15] ;
 wire \Tile_X1Y14_SS4BEG[1] ;
 wire \Tile_X1Y14_SS4BEG[2] ;
 wire \Tile_X1Y14_SS4BEG[3] ;
 wire \Tile_X1Y14_SS4BEG[4] ;
 wire \Tile_X1Y14_SS4BEG[5] ;
 wire \Tile_X1Y14_SS4BEG[6] ;
 wire \Tile_X1Y14_SS4BEG[7] ;
 wire \Tile_X1Y14_SS4BEG[8] ;
 wire \Tile_X1Y14_SS4BEG[9] ;
 wire Tile_X1Y14_UserCLKo;
 wire \Tile_X1Y14_W1BEG[0] ;
 wire \Tile_X1Y14_W1BEG[1] ;
 wire \Tile_X1Y14_W1BEG[2] ;
 wire \Tile_X1Y14_W1BEG[3] ;
 wire \Tile_X1Y14_W2BEG[0] ;
 wire \Tile_X1Y14_W2BEG[1] ;
 wire \Tile_X1Y14_W2BEG[2] ;
 wire \Tile_X1Y14_W2BEG[3] ;
 wire \Tile_X1Y14_W2BEG[4] ;
 wire \Tile_X1Y14_W2BEG[5] ;
 wire \Tile_X1Y14_W2BEG[6] ;
 wire \Tile_X1Y14_W2BEG[7] ;
 wire \Tile_X1Y14_W2BEGb[0] ;
 wire \Tile_X1Y14_W2BEGb[1] ;
 wire \Tile_X1Y14_W2BEGb[2] ;
 wire \Tile_X1Y14_W2BEGb[3] ;
 wire \Tile_X1Y14_W2BEGb[4] ;
 wire \Tile_X1Y14_W2BEGb[5] ;
 wire \Tile_X1Y14_W2BEGb[6] ;
 wire \Tile_X1Y14_W2BEGb[7] ;
 wire \Tile_X1Y14_W6BEG[0] ;
 wire \Tile_X1Y14_W6BEG[10] ;
 wire \Tile_X1Y14_W6BEG[11] ;
 wire \Tile_X1Y14_W6BEG[1] ;
 wire \Tile_X1Y14_W6BEG[2] ;
 wire \Tile_X1Y14_W6BEG[3] ;
 wire \Tile_X1Y14_W6BEG[4] ;
 wire \Tile_X1Y14_W6BEG[5] ;
 wire \Tile_X1Y14_W6BEG[6] ;
 wire \Tile_X1Y14_W6BEG[7] ;
 wire \Tile_X1Y14_W6BEG[8] ;
 wire \Tile_X1Y14_W6BEG[9] ;
 wire \Tile_X1Y14_WW4BEG[0] ;
 wire \Tile_X1Y14_WW4BEG[10] ;
 wire \Tile_X1Y14_WW4BEG[11] ;
 wire \Tile_X1Y14_WW4BEG[12] ;
 wire \Tile_X1Y14_WW4BEG[13] ;
 wire \Tile_X1Y14_WW4BEG[14] ;
 wire \Tile_X1Y14_WW4BEG[15] ;
 wire \Tile_X1Y14_WW4BEG[1] ;
 wire \Tile_X1Y14_WW4BEG[2] ;
 wire \Tile_X1Y14_WW4BEG[3] ;
 wire \Tile_X1Y14_WW4BEG[4] ;
 wire \Tile_X1Y14_WW4BEG[5] ;
 wire \Tile_X1Y14_WW4BEG[6] ;
 wire \Tile_X1Y14_WW4BEG[7] ;
 wire \Tile_X1Y14_WW4BEG[8] ;
 wire \Tile_X1Y14_WW4BEG[9] ;
 wire Tile_X1Y15_Co;
 wire \Tile_X1Y15_FrameData_O[0] ;
 wire \Tile_X1Y15_FrameData_O[10] ;
 wire \Tile_X1Y15_FrameData_O[11] ;
 wire \Tile_X1Y15_FrameData_O[12] ;
 wire \Tile_X1Y15_FrameData_O[13] ;
 wire \Tile_X1Y15_FrameData_O[14] ;
 wire \Tile_X1Y15_FrameData_O[15] ;
 wire \Tile_X1Y15_FrameData_O[16] ;
 wire \Tile_X1Y15_FrameData_O[17] ;
 wire \Tile_X1Y15_FrameData_O[18] ;
 wire \Tile_X1Y15_FrameData_O[19] ;
 wire \Tile_X1Y15_FrameData_O[1] ;
 wire \Tile_X1Y15_FrameData_O[20] ;
 wire \Tile_X1Y15_FrameData_O[21] ;
 wire \Tile_X1Y15_FrameData_O[22] ;
 wire \Tile_X1Y15_FrameData_O[23] ;
 wire \Tile_X1Y15_FrameData_O[24] ;
 wire \Tile_X1Y15_FrameData_O[25] ;
 wire \Tile_X1Y15_FrameData_O[26] ;
 wire \Tile_X1Y15_FrameData_O[27] ;
 wire \Tile_X1Y15_FrameData_O[28] ;
 wire \Tile_X1Y15_FrameData_O[29] ;
 wire \Tile_X1Y15_FrameData_O[2] ;
 wire \Tile_X1Y15_FrameData_O[30] ;
 wire \Tile_X1Y15_FrameData_O[31] ;
 wire \Tile_X1Y15_FrameData_O[3] ;
 wire \Tile_X1Y15_FrameData_O[4] ;
 wire \Tile_X1Y15_FrameData_O[5] ;
 wire \Tile_X1Y15_FrameData_O[6] ;
 wire \Tile_X1Y15_FrameData_O[7] ;
 wire \Tile_X1Y15_FrameData_O[8] ;
 wire \Tile_X1Y15_FrameData_O[9] ;
 wire \Tile_X1Y15_FrameStrobe_O[0] ;
 wire \Tile_X1Y15_FrameStrobe_O[10] ;
 wire \Tile_X1Y15_FrameStrobe_O[11] ;
 wire \Tile_X1Y15_FrameStrobe_O[12] ;
 wire \Tile_X1Y15_FrameStrobe_O[13] ;
 wire \Tile_X1Y15_FrameStrobe_O[14] ;
 wire \Tile_X1Y15_FrameStrobe_O[15] ;
 wire \Tile_X1Y15_FrameStrobe_O[16] ;
 wire \Tile_X1Y15_FrameStrobe_O[17] ;
 wire \Tile_X1Y15_FrameStrobe_O[18] ;
 wire \Tile_X1Y15_FrameStrobe_O[19] ;
 wire \Tile_X1Y15_FrameStrobe_O[1] ;
 wire \Tile_X1Y15_FrameStrobe_O[2] ;
 wire \Tile_X1Y15_FrameStrobe_O[3] ;
 wire \Tile_X1Y15_FrameStrobe_O[4] ;
 wire \Tile_X1Y15_FrameStrobe_O[5] ;
 wire \Tile_X1Y15_FrameStrobe_O[6] ;
 wire \Tile_X1Y15_FrameStrobe_O[7] ;
 wire \Tile_X1Y15_FrameStrobe_O[8] ;
 wire \Tile_X1Y15_FrameStrobe_O[9] ;
 wire \Tile_X1Y15_N1BEG[0] ;
 wire \Tile_X1Y15_N1BEG[1] ;
 wire \Tile_X1Y15_N1BEG[2] ;
 wire \Tile_X1Y15_N1BEG[3] ;
 wire \Tile_X1Y15_N2BEG[0] ;
 wire \Tile_X1Y15_N2BEG[1] ;
 wire \Tile_X1Y15_N2BEG[2] ;
 wire \Tile_X1Y15_N2BEG[3] ;
 wire \Tile_X1Y15_N2BEG[4] ;
 wire \Tile_X1Y15_N2BEG[5] ;
 wire \Tile_X1Y15_N2BEG[6] ;
 wire \Tile_X1Y15_N2BEG[7] ;
 wire \Tile_X1Y15_N2BEGb[0] ;
 wire \Tile_X1Y15_N2BEGb[1] ;
 wire \Tile_X1Y15_N2BEGb[2] ;
 wire \Tile_X1Y15_N2BEGb[3] ;
 wire \Tile_X1Y15_N2BEGb[4] ;
 wire \Tile_X1Y15_N2BEGb[5] ;
 wire \Tile_X1Y15_N2BEGb[6] ;
 wire \Tile_X1Y15_N2BEGb[7] ;
 wire \Tile_X1Y15_N4BEG[0] ;
 wire \Tile_X1Y15_N4BEG[10] ;
 wire \Tile_X1Y15_N4BEG[11] ;
 wire \Tile_X1Y15_N4BEG[12] ;
 wire \Tile_X1Y15_N4BEG[13] ;
 wire \Tile_X1Y15_N4BEG[14] ;
 wire \Tile_X1Y15_N4BEG[15] ;
 wire \Tile_X1Y15_N4BEG[1] ;
 wire \Tile_X1Y15_N4BEG[2] ;
 wire \Tile_X1Y15_N4BEG[3] ;
 wire \Tile_X1Y15_N4BEG[4] ;
 wire \Tile_X1Y15_N4BEG[5] ;
 wire \Tile_X1Y15_N4BEG[6] ;
 wire \Tile_X1Y15_N4BEG[7] ;
 wire \Tile_X1Y15_N4BEG[8] ;
 wire \Tile_X1Y15_N4BEG[9] ;
 wire \Tile_X1Y15_NN4BEG[0] ;
 wire \Tile_X1Y15_NN4BEG[10] ;
 wire \Tile_X1Y15_NN4BEG[11] ;
 wire \Tile_X1Y15_NN4BEG[12] ;
 wire \Tile_X1Y15_NN4BEG[13] ;
 wire \Tile_X1Y15_NN4BEG[14] ;
 wire \Tile_X1Y15_NN4BEG[15] ;
 wire \Tile_X1Y15_NN4BEG[1] ;
 wire \Tile_X1Y15_NN4BEG[2] ;
 wire \Tile_X1Y15_NN4BEG[3] ;
 wire \Tile_X1Y15_NN4BEG[4] ;
 wire \Tile_X1Y15_NN4BEG[5] ;
 wire \Tile_X1Y15_NN4BEG[6] ;
 wire \Tile_X1Y15_NN4BEG[7] ;
 wire \Tile_X1Y15_NN4BEG[8] ;
 wire \Tile_X1Y15_NN4BEG[9] ;
 wire Tile_X1Y15_UserCLKo;
 wire Tile_X1Y1_Co;
 wire \Tile_X1Y1_E1BEG[0] ;
 wire \Tile_X1Y1_E1BEG[1] ;
 wire \Tile_X1Y1_E1BEG[2] ;
 wire \Tile_X1Y1_E1BEG[3] ;
 wire \Tile_X1Y1_E2BEG[0] ;
 wire \Tile_X1Y1_E2BEG[1] ;
 wire \Tile_X1Y1_E2BEG[2] ;
 wire \Tile_X1Y1_E2BEG[3] ;
 wire \Tile_X1Y1_E2BEG[4] ;
 wire \Tile_X1Y1_E2BEG[5] ;
 wire \Tile_X1Y1_E2BEG[6] ;
 wire \Tile_X1Y1_E2BEG[7] ;
 wire \Tile_X1Y1_E2BEGb[0] ;
 wire \Tile_X1Y1_E2BEGb[1] ;
 wire \Tile_X1Y1_E2BEGb[2] ;
 wire \Tile_X1Y1_E2BEGb[3] ;
 wire \Tile_X1Y1_E2BEGb[4] ;
 wire \Tile_X1Y1_E2BEGb[5] ;
 wire \Tile_X1Y1_E2BEGb[6] ;
 wire \Tile_X1Y1_E2BEGb[7] ;
 wire \Tile_X1Y1_E6BEG[0] ;
 wire \Tile_X1Y1_E6BEG[10] ;
 wire \Tile_X1Y1_E6BEG[11] ;
 wire \Tile_X1Y1_E6BEG[1] ;
 wire \Tile_X1Y1_E6BEG[2] ;
 wire \Tile_X1Y1_E6BEG[3] ;
 wire \Tile_X1Y1_E6BEG[4] ;
 wire \Tile_X1Y1_E6BEG[5] ;
 wire \Tile_X1Y1_E6BEG[6] ;
 wire \Tile_X1Y1_E6BEG[7] ;
 wire \Tile_X1Y1_E6BEG[8] ;
 wire \Tile_X1Y1_E6BEG[9] ;
 wire \Tile_X1Y1_EE4BEG[0] ;
 wire \Tile_X1Y1_EE4BEG[10] ;
 wire \Tile_X1Y1_EE4BEG[11] ;
 wire \Tile_X1Y1_EE4BEG[12] ;
 wire \Tile_X1Y1_EE4BEG[13] ;
 wire \Tile_X1Y1_EE4BEG[14] ;
 wire \Tile_X1Y1_EE4BEG[15] ;
 wire \Tile_X1Y1_EE4BEG[1] ;
 wire \Tile_X1Y1_EE4BEG[2] ;
 wire \Tile_X1Y1_EE4BEG[3] ;
 wire \Tile_X1Y1_EE4BEG[4] ;
 wire \Tile_X1Y1_EE4BEG[5] ;
 wire \Tile_X1Y1_EE4BEG[6] ;
 wire \Tile_X1Y1_EE4BEG[7] ;
 wire \Tile_X1Y1_EE4BEG[8] ;
 wire \Tile_X1Y1_EE4BEG[9] ;
 wire \Tile_X1Y1_FrameData_O[0] ;
 wire \Tile_X1Y1_FrameData_O[10] ;
 wire \Tile_X1Y1_FrameData_O[11] ;
 wire \Tile_X1Y1_FrameData_O[12] ;
 wire \Tile_X1Y1_FrameData_O[13] ;
 wire \Tile_X1Y1_FrameData_O[14] ;
 wire \Tile_X1Y1_FrameData_O[15] ;
 wire \Tile_X1Y1_FrameData_O[16] ;
 wire \Tile_X1Y1_FrameData_O[17] ;
 wire \Tile_X1Y1_FrameData_O[18] ;
 wire \Tile_X1Y1_FrameData_O[19] ;
 wire \Tile_X1Y1_FrameData_O[1] ;
 wire \Tile_X1Y1_FrameData_O[20] ;
 wire \Tile_X1Y1_FrameData_O[21] ;
 wire \Tile_X1Y1_FrameData_O[22] ;
 wire \Tile_X1Y1_FrameData_O[23] ;
 wire \Tile_X1Y1_FrameData_O[24] ;
 wire \Tile_X1Y1_FrameData_O[25] ;
 wire \Tile_X1Y1_FrameData_O[26] ;
 wire \Tile_X1Y1_FrameData_O[27] ;
 wire \Tile_X1Y1_FrameData_O[28] ;
 wire \Tile_X1Y1_FrameData_O[29] ;
 wire \Tile_X1Y1_FrameData_O[2] ;
 wire \Tile_X1Y1_FrameData_O[30] ;
 wire \Tile_X1Y1_FrameData_O[31] ;
 wire \Tile_X1Y1_FrameData_O[3] ;
 wire \Tile_X1Y1_FrameData_O[4] ;
 wire \Tile_X1Y1_FrameData_O[5] ;
 wire \Tile_X1Y1_FrameData_O[6] ;
 wire \Tile_X1Y1_FrameData_O[7] ;
 wire \Tile_X1Y1_FrameData_O[8] ;
 wire \Tile_X1Y1_FrameData_O[9] ;
 wire \Tile_X1Y1_FrameStrobe_O[0] ;
 wire \Tile_X1Y1_FrameStrobe_O[10] ;
 wire \Tile_X1Y1_FrameStrobe_O[11] ;
 wire \Tile_X1Y1_FrameStrobe_O[12] ;
 wire \Tile_X1Y1_FrameStrobe_O[13] ;
 wire \Tile_X1Y1_FrameStrobe_O[14] ;
 wire \Tile_X1Y1_FrameStrobe_O[15] ;
 wire \Tile_X1Y1_FrameStrobe_O[16] ;
 wire \Tile_X1Y1_FrameStrobe_O[17] ;
 wire \Tile_X1Y1_FrameStrobe_O[18] ;
 wire \Tile_X1Y1_FrameStrobe_O[19] ;
 wire \Tile_X1Y1_FrameStrobe_O[1] ;
 wire \Tile_X1Y1_FrameStrobe_O[2] ;
 wire \Tile_X1Y1_FrameStrobe_O[3] ;
 wire \Tile_X1Y1_FrameStrobe_O[4] ;
 wire \Tile_X1Y1_FrameStrobe_O[5] ;
 wire \Tile_X1Y1_FrameStrobe_O[6] ;
 wire \Tile_X1Y1_FrameStrobe_O[7] ;
 wire \Tile_X1Y1_FrameStrobe_O[8] ;
 wire \Tile_X1Y1_FrameStrobe_O[9] ;
 wire \Tile_X1Y1_N1BEG[0] ;
 wire \Tile_X1Y1_N1BEG[1] ;
 wire \Tile_X1Y1_N1BEG[2] ;
 wire \Tile_X1Y1_N1BEG[3] ;
 wire \Tile_X1Y1_N2BEG[0] ;
 wire \Tile_X1Y1_N2BEG[1] ;
 wire \Tile_X1Y1_N2BEG[2] ;
 wire \Tile_X1Y1_N2BEG[3] ;
 wire \Tile_X1Y1_N2BEG[4] ;
 wire \Tile_X1Y1_N2BEG[5] ;
 wire \Tile_X1Y1_N2BEG[6] ;
 wire \Tile_X1Y1_N2BEG[7] ;
 wire \Tile_X1Y1_N2BEGb[0] ;
 wire \Tile_X1Y1_N2BEGb[1] ;
 wire \Tile_X1Y1_N2BEGb[2] ;
 wire \Tile_X1Y1_N2BEGb[3] ;
 wire \Tile_X1Y1_N2BEGb[4] ;
 wire \Tile_X1Y1_N2BEGb[5] ;
 wire \Tile_X1Y1_N2BEGb[6] ;
 wire \Tile_X1Y1_N2BEGb[7] ;
 wire \Tile_X1Y1_N4BEG[0] ;
 wire \Tile_X1Y1_N4BEG[10] ;
 wire \Tile_X1Y1_N4BEG[11] ;
 wire \Tile_X1Y1_N4BEG[12] ;
 wire \Tile_X1Y1_N4BEG[13] ;
 wire \Tile_X1Y1_N4BEG[14] ;
 wire \Tile_X1Y1_N4BEG[15] ;
 wire \Tile_X1Y1_N4BEG[1] ;
 wire \Tile_X1Y1_N4BEG[2] ;
 wire \Tile_X1Y1_N4BEG[3] ;
 wire \Tile_X1Y1_N4BEG[4] ;
 wire \Tile_X1Y1_N4BEG[5] ;
 wire \Tile_X1Y1_N4BEG[6] ;
 wire \Tile_X1Y1_N4BEG[7] ;
 wire \Tile_X1Y1_N4BEG[8] ;
 wire \Tile_X1Y1_N4BEG[9] ;
 wire \Tile_X1Y1_NN4BEG[0] ;
 wire \Tile_X1Y1_NN4BEG[10] ;
 wire \Tile_X1Y1_NN4BEG[11] ;
 wire \Tile_X1Y1_NN4BEG[12] ;
 wire \Tile_X1Y1_NN4BEG[13] ;
 wire \Tile_X1Y1_NN4BEG[14] ;
 wire \Tile_X1Y1_NN4BEG[15] ;
 wire \Tile_X1Y1_NN4BEG[1] ;
 wire \Tile_X1Y1_NN4BEG[2] ;
 wire \Tile_X1Y1_NN4BEG[3] ;
 wire \Tile_X1Y1_NN4BEG[4] ;
 wire \Tile_X1Y1_NN4BEG[5] ;
 wire \Tile_X1Y1_NN4BEG[6] ;
 wire \Tile_X1Y1_NN4BEG[7] ;
 wire \Tile_X1Y1_NN4BEG[8] ;
 wire \Tile_X1Y1_NN4BEG[9] ;
 wire \Tile_X1Y1_S1BEG[0] ;
 wire \Tile_X1Y1_S1BEG[1] ;
 wire \Tile_X1Y1_S1BEG[2] ;
 wire \Tile_X1Y1_S1BEG[3] ;
 wire \Tile_X1Y1_S2BEG[0] ;
 wire \Tile_X1Y1_S2BEG[1] ;
 wire \Tile_X1Y1_S2BEG[2] ;
 wire \Tile_X1Y1_S2BEG[3] ;
 wire \Tile_X1Y1_S2BEG[4] ;
 wire \Tile_X1Y1_S2BEG[5] ;
 wire \Tile_X1Y1_S2BEG[6] ;
 wire \Tile_X1Y1_S2BEG[7] ;
 wire \Tile_X1Y1_S2BEGb[0] ;
 wire \Tile_X1Y1_S2BEGb[1] ;
 wire \Tile_X1Y1_S2BEGb[2] ;
 wire \Tile_X1Y1_S2BEGb[3] ;
 wire \Tile_X1Y1_S2BEGb[4] ;
 wire \Tile_X1Y1_S2BEGb[5] ;
 wire \Tile_X1Y1_S2BEGb[6] ;
 wire \Tile_X1Y1_S2BEGb[7] ;
 wire \Tile_X1Y1_S4BEG[0] ;
 wire \Tile_X1Y1_S4BEG[10] ;
 wire \Tile_X1Y1_S4BEG[11] ;
 wire \Tile_X1Y1_S4BEG[12] ;
 wire \Tile_X1Y1_S4BEG[13] ;
 wire \Tile_X1Y1_S4BEG[14] ;
 wire \Tile_X1Y1_S4BEG[15] ;
 wire \Tile_X1Y1_S4BEG[1] ;
 wire \Tile_X1Y1_S4BEG[2] ;
 wire \Tile_X1Y1_S4BEG[3] ;
 wire \Tile_X1Y1_S4BEG[4] ;
 wire \Tile_X1Y1_S4BEG[5] ;
 wire \Tile_X1Y1_S4BEG[6] ;
 wire \Tile_X1Y1_S4BEG[7] ;
 wire \Tile_X1Y1_S4BEG[8] ;
 wire \Tile_X1Y1_S4BEG[9] ;
 wire \Tile_X1Y1_SS4BEG[0] ;
 wire \Tile_X1Y1_SS4BEG[10] ;
 wire \Tile_X1Y1_SS4BEG[11] ;
 wire \Tile_X1Y1_SS4BEG[12] ;
 wire \Tile_X1Y1_SS4BEG[13] ;
 wire \Tile_X1Y1_SS4BEG[14] ;
 wire \Tile_X1Y1_SS4BEG[15] ;
 wire \Tile_X1Y1_SS4BEG[1] ;
 wire \Tile_X1Y1_SS4BEG[2] ;
 wire \Tile_X1Y1_SS4BEG[3] ;
 wire \Tile_X1Y1_SS4BEG[4] ;
 wire \Tile_X1Y1_SS4BEG[5] ;
 wire \Tile_X1Y1_SS4BEG[6] ;
 wire \Tile_X1Y1_SS4BEG[7] ;
 wire \Tile_X1Y1_SS4BEG[8] ;
 wire \Tile_X1Y1_SS4BEG[9] ;
 wire Tile_X1Y1_UserCLKo;
 wire \Tile_X1Y1_W1BEG[0] ;
 wire \Tile_X1Y1_W1BEG[1] ;
 wire \Tile_X1Y1_W1BEG[2] ;
 wire \Tile_X1Y1_W1BEG[3] ;
 wire \Tile_X1Y1_W2BEG[0] ;
 wire \Tile_X1Y1_W2BEG[1] ;
 wire \Tile_X1Y1_W2BEG[2] ;
 wire \Tile_X1Y1_W2BEG[3] ;
 wire \Tile_X1Y1_W2BEG[4] ;
 wire \Tile_X1Y1_W2BEG[5] ;
 wire \Tile_X1Y1_W2BEG[6] ;
 wire \Tile_X1Y1_W2BEG[7] ;
 wire \Tile_X1Y1_W2BEGb[0] ;
 wire \Tile_X1Y1_W2BEGb[1] ;
 wire \Tile_X1Y1_W2BEGb[2] ;
 wire \Tile_X1Y1_W2BEGb[3] ;
 wire \Tile_X1Y1_W2BEGb[4] ;
 wire \Tile_X1Y1_W2BEGb[5] ;
 wire \Tile_X1Y1_W2BEGb[6] ;
 wire \Tile_X1Y1_W2BEGb[7] ;
 wire \Tile_X1Y1_W6BEG[0] ;
 wire \Tile_X1Y1_W6BEG[10] ;
 wire \Tile_X1Y1_W6BEG[11] ;
 wire \Tile_X1Y1_W6BEG[1] ;
 wire \Tile_X1Y1_W6BEG[2] ;
 wire \Tile_X1Y1_W6BEG[3] ;
 wire \Tile_X1Y1_W6BEG[4] ;
 wire \Tile_X1Y1_W6BEG[5] ;
 wire \Tile_X1Y1_W6BEG[6] ;
 wire \Tile_X1Y1_W6BEG[7] ;
 wire \Tile_X1Y1_W6BEG[8] ;
 wire \Tile_X1Y1_W6BEG[9] ;
 wire \Tile_X1Y1_WW4BEG[0] ;
 wire \Tile_X1Y1_WW4BEG[10] ;
 wire \Tile_X1Y1_WW4BEG[11] ;
 wire \Tile_X1Y1_WW4BEG[12] ;
 wire \Tile_X1Y1_WW4BEG[13] ;
 wire \Tile_X1Y1_WW4BEG[14] ;
 wire \Tile_X1Y1_WW4BEG[15] ;
 wire \Tile_X1Y1_WW4BEG[1] ;
 wire \Tile_X1Y1_WW4BEG[2] ;
 wire \Tile_X1Y1_WW4BEG[3] ;
 wire \Tile_X1Y1_WW4BEG[4] ;
 wire \Tile_X1Y1_WW4BEG[5] ;
 wire \Tile_X1Y1_WW4BEG[6] ;
 wire \Tile_X1Y1_WW4BEG[7] ;
 wire \Tile_X1Y1_WW4BEG[8] ;
 wire \Tile_X1Y1_WW4BEG[9] ;
 wire Tile_X1Y2_Co;
 wire \Tile_X1Y2_E1BEG[0] ;
 wire \Tile_X1Y2_E1BEG[1] ;
 wire \Tile_X1Y2_E1BEG[2] ;
 wire \Tile_X1Y2_E1BEG[3] ;
 wire \Tile_X1Y2_E2BEG[0] ;
 wire \Tile_X1Y2_E2BEG[1] ;
 wire \Tile_X1Y2_E2BEG[2] ;
 wire \Tile_X1Y2_E2BEG[3] ;
 wire \Tile_X1Y2_E2BEG[4] ;
 wire \Tile_X1Y2_E2BEG[5] ;
 wire \Tile_X1Y2_E2BEG[6] ;
 wire \Tile_X1Y2_E2BEG[7] ;
 wire \Tile_X1Y2_E2BEGb[0] ;
 wire \Tile_X1Y2_E2BEGb[1] ;
 wire \Tile_X1Y2_E2BEGb[2] ;
 wire \Tile_X1Y2_E2BEGb[3] ;
 wire \Tile_X1Y2_E2BEGb[4] ;
 wire \Tile_X1Y2_E2BEGb[5] ;
 wire \Tile_X1Y2_E2BEGb[6] ;
 wire \Tile_X1Y2_E2BEGb[7] ;
 wire \Tile_X1Y2_E6BEG[0] ;
 wire \Tile_X1Y2_E6BEG[10] ;
 wire \Tile_X1Y2_E6BEG[11] ;
 wire \Tile_X1Y2_E6BEG[1] ;
 wire \Tile_X1Y2_E6BEG[2] ;
 wire \Tile_X1Y2_E6BEG[3] ;
 wire \Tile_X1Y2_E6BEG[4] ;
 wire \Tile_X1Y2_E6BEG[5] ;
 wire \Tile_X1Y2_E6BEG[6] ;
 wire \Tile_X1Y2_E6BEG[7] ;
 wire \Tile_X1Y2_E6BEG[8] ;
 wire \Tile_X1Y2_E6BEG[9] ;
 wire \Tile_X1Y2_EE4BEG[0] ;
 wire \Tile_X1Y2_EE4BEG[10] ;
 wire \Tile_X1Y2_EE4BEG[11] ;
 wire \Tile_X1Y2_EE4BEG[12] ;
 wire \Tile_X1Y2_EE4BEG[13] ;
 wire \Tile_X1Y2_EE4BEG[14] ;
 wire \Tile_X1Y2_EE4BEG[15] ;
 wire \Tile_X1Y2_EE4BEG[1] ;
 wire \Tile_X1Y2_EE4BEG[2] ;
 wire \Tile_X1Y2_EE4BEG[3] ;
 wire \Tile_X1Y2_EE4BEG[4] ;
 wire \Tile_X1Y2_EE4BEG[5] ;
 wire \Tile_X1Y2_EE4BEG[6] ;
 wire \Tile_X1Y2_EE4BEG[7] ;
 wire \Tile_X1Y2_EE4BEG[8] ;
 wire \Tile_X1Y2_EE4BEG[9] ;
 wire \Tile_X1Y2_FrameData_O[0] ;
 wire \Tile_X1Y2_FrameData_O[10] ;
 wire \Tile_X1Y2_FrameData_O[11] ;
 wire \Tile_X1Y2_FrameData_O[12] ;
 wire \Tile_X1Y2_FrameData_O[13] ;
 wire \Tile_X1Y2_FrameData_O[14] ;
 wire \Tile_X1Y2_FrameData_O[15] ;
 wire \Tile_X1Y2_FrameData_O[16] ;
 wire \Tile_X1Y2_FrameData_O[17] ;
 wire \Tile_X1Y2_FrameData_O[18] ;
 wire \Tile_X1Y2_FrameData_O[19] ;
 wire \Tile_X1Y2_FrameData_O[1] ;
 wire \Tile_X1Y2_FrameData_O[20] ;
 wire \Tile_X1Y2_FrameData_O[21] ;
 wire \Tile_X1Y2_FrameData_O[22] ;
 wire \Tile_X1Y2_FrameData_O[23] ;
 wire \Tile_X1Y2_FrameData_O[24] ;
 wire \Tile_X1Y2_FrameData_O[25] ;
 wire \Tile_X1Y2_FrameData_O[26] ;
 wire \Tile_X1Y2_FrameData_O[27] ;
 wire \Tile_X1Y2_FrameData_O[28] ;
 wire \Tile_X1Y2_FrameData_O[29] ;
 wire \Tile_X1Y2_FrameData_O[2] ;
 wire \Tile_X1Y2_FrameData_O[30] ;
 wire \Tile_X1Y2_FrameData_O[31] ;
 wire \Tile_X1Y2_FrameData_O[3] ;
 wire \Tile_X1Y2_FrameData_O[4] ;
 wire \Tile_X1Y2_FrameData_O[5] ;
 wire \Tile_X1Y2_FrameData_O[6] ;
 wire \Tile_X1Y2_FrameData_O[7] ;
 wire \Tile_X1Y2_FrameData_O[8] ;
 wire \Tile_X1Y2_FrameData_O[9] ;
 wire \Tile_X1Y2_FrameStrobe_O[0] ;
 wire \Tile_X1Y2_FrameStrobe_O[10] ;
 wire \Tile_X1Y2_FrameStrobe_O[11] ;
 wire \Tile_X1Y2_FrameStrobe_O[12] ;
 wire \Tile_X1Y2_FrameStrobe_O[13] ;
 wire \Tile_X1Y2_FrameStrobe_O[14] ;
 wire \Tile_X1Y2_FrameStrobe_O[15] ;
 wire \Tile_X1Y2_FrameStrobe_O[16] ;
 wire \Tile_X1Y2_FrameStrobe_O[17] ;
 wire \Tile_X1Y2_FrameStrobe_O[18] ;
 wire \Tile_X1Y2_FrameStrobe_O[19] ;
 wire \Tile_X1Y2_FrameStrobe_O[1] ;
 wire \Tile_X1Y2_FrameStrobe_O[2] ;
 wire \Tile_X1Y2_FrameStrobe_O[3] ;
 wire \Tile_X1Y2_FrameStrobe_O[4] ;
 wire \Tile_X1Y2_FrameStrobe_O[5] ;
 wire \Tile_X1Y2_FrameStrobe_O[6] ;
 wire \Tile_X1Y2_FrameStrobe_O[7] ;
 wire \Tile_X1Y2_FrameStrobe_O[8] ;
 wire \Tile_X1Y2_FrameStrobe_O[9] ;
 wire \Tile_X1Y2_N1BEG[0] ;
 wire \Tile_X1Y2_N1BEG[1] ;
 wire \Tile_X1Y2_N1BEG[2] ;
 wire \Tile_X1Y2_N1BEG[3] ;
 wire \Tile_X1Y2_N2BEG[0] ;
 wire \Tile_X1Y2_N2BEG[1] ;
 wire \Tile_X1Y2_N2BEG[2] ;
 wire \Tile_X1Y2_N2BEG[3] ;
 wire \Tile_X1Y2_N2BEG[4] ;
 wire \Tile_X1Y2_N2BEG[5] ;
 wire \Tile_X1Y2_N2BEG[6] ;
 wire \Tile_X1Y2_N2BEG[7] ;
 wire \Tile_X1Y2_N2BEGb[0] ;
 wire \Tile_X1Y2_N2BEGb[1] ;
 wire \Tile_X1Y2_N2BEGb[2] ;
 wire \Tile_X1Y2_N2BEGb[3] ;
 wire \Tile_X1Y2_N2BEGb[4] ;
 wire \Tile_X1Y2_N2BEGb[5] ;
 wire \Tile_X1Y2_N2BEGb[6] ;
 wire \Tile_X1Y2_N2BEGb[7] ;
 wire \Tile_X1Y2_N4BEG[0] ;
 wire \Tile_X1Y2_N4BEG[10] ;
 wire \Tile_X1Y2_N4BEG[11] ;
 wire \Tile_X1Y2_N4BEG[12] ;
 wire \Tile_X1Y2_N4BEG[13] ;
 wire \Tile_X1Y2_N4BEG[14] ;
 wire \Tile_X1Y2_N4BEG[15] ;
 wire \Tile_X1Y2_N4BEG[1] ;
 wire \Tile_X1Y2_N4BEG[2] ;
 wire \Tile_X1Y2_N4BEG[3] ;
 wire \Tile_X1Y2_N4BEG[4] ;
 wire \Tile_X1Y2_N4BEG[5] ;
 wire \Tile_X1Y2_N4BEG[6] ;
 wire \Tile_X1Y2_N4BEG[7] ;
 wire \Tile_X1Y2_N4BEG[8] ;
 wire \Tile_X1Y2_N4BEG[9] ;
 wire \Tile_X1Y2_NN4BEG[0] ;
 wire \Tile_X1Y2_NN4BEG[10] ;
 wire \Tile_X1Y2_NN4BEG[11] ;
 wire \Tile_X1Y2_NN4BEG[12] ;
 wire \Tile_X1Y2_NN4BEG[13] ;
 wire \Tile_X1Y2_NN4BEG[14] ;
 wire \Tile_X1Y2_NN4BEG[15] ;
 wire \Tile_X1Y2_NN4BEG[1] ;
 wire \Tile_X1Y2_NN4BEG[2] ;
 wire \Tile_X1Y2_NN4BEG[3] ;
 wire \Tile_X1Y2_NN4BEG[4] ;
 wire \Tile_X1Y2_NN4BEG[5] ;
 wire \Tile_X1Y2_NN4BEG[6] ;
 wire \Tile_X1Y2_NN4BEG[7] ;
 wire \Tile_X1Y2_NN4BEG[8] ;
 wire \Tile_X1Y2_NN4BEG[9] ;
 wire \Tile_X1Y2_S1BEG[0] ;
 wire \Tile_X1Y2_S1BEG[1] ;
 wire \Tile_X1Y2_S1BEG[2] ;
 wire \Tile_X1Y2_S1BEG[3] ;
 wire \Tile_X1Y2_S2BEG[0] ;
 wire \Tile_X1Y2_S2BEG[1] ;
 wire \Tile_X1Y2_S2BEG[2] ;
 wire \Tile_X1Y2_S2BEG[3] ;
 wire \Tile_X1Y2_S2BEG[4] ;
 wire \Tile_X1Y2_S2BEG[5] ;
 wire \Tile_X1Y2_S2BEG[6] ;
 wire \Tile_X1Y2_S2BEG[7] ;
 wire \Tile_X1Y2_S2BEGb[0] ;
 wire \Tile_X1Y2_S2BEGb[1] ;
 wire \Tile_X1Y2_S2BEGb[2] ;
 wire \Tile_X1Y2_S2BEGb[3] ;
 wire \Tile_X1Y2_S2BEGb[4] ;
 wire \Tile_X1Y2_S2BEGb[5] ;
 wire \Tile_X1Y2_S2BEGb[6] ;
 wire \Tile_X1Y2_S2BEGb[7] ;
 wire \Tile_X1Y2_S4BEG[0] ;
 wire \Tile_X1Y2_S4BEG[10] ;
 wire \Tile_X1Y2_S4BEG[11] ;
 wire \Tile_X1Y2_S4BEG[12] ;
 wire \Tile_X1Y2_S4BEG[13] ;
 wire \Tile_X1Y2_S4BEG[14] ;
 wire \Tile_X1Y2_S4BEG[15] ;
 wire \Tile_X1Y2_S4BEG[1] ;
 wire \Tile_X1Y2_S4BEG[2] ;
 wire \Tile_X1Y2_S4BEG[3] ;
 wire \Tile_X1Y2_S4BEG[4] ;
 wire \Tile_X1Y2_S4BEG[5] ;
 wire \Tile_X1Y2_S4BEG[6] ;
 wire \Tile_X1Y2_S4BEG[7] ;
 wire \Tile_X1Y2_S4BEG[8] ;
 wire \Tile_X1Y2_S4BEG[9] ;
 wire \Tile_X1Y2_SS4BEG[0] ;
 wire \Tile_X1Y2_SS4BEG[10] ;
 wire \Tile_X1Y2_SS4BEG[11] ;
 wire \Tile_X1Y2_SS4BEG[12] ;
 wire \Tile_X1Y2_SS4BEG[13] ;
 wire \Tile_X1Y2_SS4BEG[14] ;
 wire \Tile_X1Y2_SS4BEG[15] ;
 wire \Tile_X1Y2_SS4BEG[1] ;
 wire \Tile_X1Y2_SS4BEG[2] ;
 wire \Tile_X1Y2_SS4BEG[3] ;
 wire \Tile_X1Y2_SS4BEG[4] ;
 wire \Tile_X1Y2_SS4BEG[5] ;
 wire \Tile_X1Y2_SS4BEG[6] ;
 wire \Tile_X1Y2_SS4BEG[7] ;
 wire \Tile_X1Y2_SS4BEG[8] ;
 wire \Tile_X1Y2_SS4BEG[9] ;
 wire Tile_X1Y2_UserCLKo;
 wire \Tile_X1Y2_W1BEG[0] ;
 wire \Tile_X1Y2_W1BEG[1] ;
 wire \Tile_X1Y2_W1BEG[2] ;
 wire \Tile_X1Y2_W1BEG[3] ;
 wire \Tile_X1Y2_W2BEG[0] ;
 wire \Tile_X1Y2_W2BEG[1] ;
 wire \Tile_X1Y2_W2BEG[2] ;
 wire \Tile_X1Y2_W2BEG[3] ;
 wire \Tile_X1Y2_W2BEG[4] ;
 wire \Tile_X1Y2_W2BEG[5] ;
 wire \Tile_X1Y2_W2BEG[6] ;
 wire \Tile_X1Y2_W2BEG[7] ;
 wire \Tile_X1Y2_W2BEGb[0] ;
 wire \Tile_X1Y2_W2BEGb[1] ;
 wire \Tile_X1Y2_W2BEGb[2] ;
 wire \Tile_X1Y2_W2BEGb[3] ;
 wire \Tile_X1Y2_W2BEGb[4] ;
 wire \Tile_X1Y2_W2BEGb[5] ;
 wire \Tile_X1Y2_W2BEGb[6] ;
 wire \Tile_X1Y2_W2BEGb[7] ;
 wire \Tile_X1Y2_W6BEG[0] ;
 wire \Tile_X1Y2_W6BEG[10] ;
 wire \Tile_X1Y2_W6BEG[11] ;
 wire \Tile_X1Y2_W6BEG[1] ;
 wire \Tile_X1Y2_W6BEG[2] ;
 wire \Tile_X1Y2_W6BEG[3] ;
 wire \Tile_X1Y2_W6BEG[4] ;
 wire \Tile_X1Y2_W6BEG[5] ;
 wire \Tile_X1Y2_W6BEG[6] ;
 wire \Tile_X1Y2_W6BEG[7] ;
 wire \Tile_X1Y2_W6BEG[8] ;
 wire \Tile_X1Y2_W6BEG[9] ;
 wire \Tile_X1Y2_WW4BEG[0] ;
 wire \Tile_X1Y2_WW4BEG[10] ;
 wire \Tile_X1Y2_WW4BEG[11] ;
 wire \Tile_X1Y2_WW4BEG[12] ;
 wire \Tile_X1Y2_WW4BEG[13] ;
 wire \Tile_X1Y2_WW4BEG[14] ;
 wire \Tile_X1Y2_WW4BEG[15] ;
 wire \Tile_X1Y2_WW4BEG[1] ;
 wire \Tile_X1Y2_WW4BEG[2] ;
 wire \Tile_X1Y2_WW4BEG[3] ;
 wire \Tile_X1Y2_WW4BEG[4] ;
 wire \Tile_X1Y2_WW4BEG[5] ;
 wire \Tile_X1Y2_WW4BEG[6] ;
 wire \Tile_X1Y2_WW4BEG[7] ;
 wire \Tile_X1Y2_WW4BEG[8] ;
 wire \Tile_X1Y2_WW4BEG[9] ;
 wire Tile_X1Y3_Co;
 wire \Tile_X1Y3_E1BEG[0] ;
 wire \Tile_X1Y3_E1BEG[1] ;
 wire \Tile_X1Y3_E1BEG[2] ;
 wire \Tile_X1Y3_E1BEG[3] ;
 wire \Tile_X1Y3_E2BEG[0] ;
 wire \Tile_X1Y3_E2BEG[1] ;
 wire \Tile_X1Y3_E2BEG[2] ;
 wire \Tile_X1Y3_E2BEG[3] ;
 wire \Tile_X1Y3_E2BEG[4] ;
 wire \Tile_X1Y3_E2BEG[5] ;
 wire \Tile_X1Y3_E2BEG[6] ;
 wire \Tile_X1Y3_E2BEG[7] ;
 wire \Tile_X1Y3_E2BEGb[0] ;
 wire \Tile_X1Y3_E2BEGb[1] ;
 wire \Tile_X1Y3_E2BEGb[2] ;
 wire \Tile_X1Y3_E2BEGb[3] ;
 wire \Tile_X1Y3_E2BEGb[4] ;
 wire \Tile_X1Y3_E2BEGb[5] ;
 wire \Tile_X1Y3_E2BEGb[6] ;
 wire \Tile_X1Y3_E2BEGb[7] ;
 wire \Tile_X1Y3_E6BEG[0] ;
 wire \Tile_X1Y3_E6BEG[10] ;
 wire \Tile_X1Y3_E6BEG[11] ;
 wire \Tile_X1Y3_E6BEG[1] ;
 wire \Tile_X1Y3_E6BEG[2] ;
 wire \Tile_X1Y3_E6BEG[3] ;
 wire \Tile_X1Y3_E6BEG[4] ;
 wire \Tile_X1Y3_E6BEG[5] ;
 wire \Tile_X1Y3_E6BEG[6] ;
 wire \Tile_X1Y3_E6BEG[7] ;
 wire \Tile_X1Y3_E6BEG[8] ;
 wire \Tile_X1Y3_E6BEG[9] ;
 wire \Tile_X1Y3_EE4BEG[0] ;
 wire \Tile_X1Y3_EE4BEG[10] ;
 wire \Tile_X1Y3_EE4BEG[11] ;
 wire \Tile_X1Y3_EE4BEG[12] ;
 wire \Tile_X1Y3_EE4BEG[13] ;
 wire \Tile_X1Y3_EE4BEG[14] ;
 wire \Tile_X1Y3_EE4BEG[15] ;
 wire \Tile_X1Y3_EE4BEG[1] ;
 wire \Tile_X1Y3_EE4BEG[2] ;
 wire \Tile_X1Y3_EE4BEG[3] ;
 wire \Tile_X1Y3_EE4BEG[4] ;
 wire \Tile_X1Y3_EE4BEG[5] ;
 wire \Tile_X1Y3_EE4BEG[6] ;
 wire \Tile_X1Y3_EE4BEG[7] ;
 wire \Tile_X1Y3_EE4BEG[8] ;
 wire \Tile_X1Y3_EE4BEG[9] ;
 wire \Tile_X1Y3_FrameData_O[0] ;
 wire \Tile_X1Y3_FrameData_O[10] ;
 wire \Tile_X1Y3_FrameData_O[11] ;
 wire \Tile_X1Y3_FrameData_O[12] ;
 wire \Tile_X1Y3_FrameData_O[13] ;
 wire \Tile_X1Y3_FrameData_O[14] ;
 wire \Tile_X1Y3_FrameData_O[15] ;
 wire \Tile_X1Y3_FrameData_O[16] ;
 wire \Tile_X1Y3_FrameData_O[17] ;
 wire \Tile_X1Y3_FrameData_O[18] ;
 wire \Tile_X1Y3_FrameData_O[19] ;
 wire \Tile_X1Y3_FrameData_O[1] ;
 wire \Tile_X1Y3_FrameData_O[20] ;
 wire \Tile_X1Y3_FrameData_O[21] ;
 wire \Tile_X1Y3_FrameData_O[22] ;
 wire \Tile_X1Y3_FrameData_O[23] ;
 wire \Tile_X1Y3_FrameData_O[24] ;
 wire \Tile_X1Y3_FrameData_O[25] ;
 wire \Tile_X1Y3_FrameData_O[26] ;
 wire \Tile_X1Y3_FrameData_O[27] ;
 wire \Tile_X1Y3_FrameData_O[28] ;
 wire \Tile_X1Y3_FrameData_O[29] ;
 wire \Tile_X1Y3_FrameData_O[2] ;
 wire \Tile_X1Y3_FrameData_O[30] ;
 wire \Tile_X1Y3_FrameData_O[31] ;
 wire \Tile_X1Y3_FrameData_O[3] ;
 wire \Tile_X1Y3_FrameData_O[4] ;
 wire \Tile_X1Y3_FrameData_O[5] ;
 wire \Tile_X1Y3_FrameData_O[6] ;
 wire \Tile_X1Y3_FrameData_O[7] ;
 wire \Tile_X1Y3_FrameData_O[8] ;
 wire \Tile_X1Y3_FrameData_O[9] ;
 wire \Tile_X1Y3_FrameStrobe_O[0] ;
 wire \Tile_X1Y3_FrameStrobe_O[10] ;
 wire \Tile_X1Y3_FrameStrobe_O[11] ;
 wire \Tile_X1Y3_FrameStrobe_O[12] ;
 wire \Tile_X1Y3_FrameStrobe_O[13] ;
 wire \Tile_X1Y3_FrameStrobe_O[14] ;
 wire \Tile_X1Y3_FrameStrobe_O[15] ;
 wire \Tile_X1Y3_FrameStrobe_O[16] ;
 wire \Tile_X1Y3_FrameStrobe_O[17] ;
 wire \Tile_X1Y3_FrameStrobe_O[18] ;
 wire \Tile_X1Y3_FrameStrobe_O[19] ;
 wire \Tile_X1Y3_FrameStrobe_O[1] ;
 wire \Tile_X1Y3_FrameStrobe_O[2] ;
 wire \Tile_X1Y3_FrameStrobe_O[3] ;
 wire \Tile_X1Y3_FrameStrobe_O[4] ;
 wire \Tile_X1Y3_FrameStrobe_O[5] ;
 wire \Tile_X1Y3_FrameStrobe_O[6] ;
 wire \Tile_X1Y3_FrameStrobe_O[7] ;
 wire \Tile_X1Y3_FrameStrobe_O[8] ;
 wire \Tile_X1Y3_FrameStrobe_O[9] ;
 wire \Tile_X1Y3_N1BEG[0] ;
 wire \Tile_X1Y3_N1BEG[1] ;
 wire \Tile_X1Y3_N1BEG[2] ;
 wire \Tile_X1Y3_N1BEG[3] ;
 wire \Tile_X1Y3_N2BEG[0] ;
 wire \Tile_X1Y3_N2BEG[1] ;
 wire \Tile_X1Y3_N2BEG[2] ;
 wire \Tile_X1Y3_N2BEG[3] ;
 wire \Tile_X1Y3_N2BEG[4] ;
 wire \Tile_X1Y3_N2BEG[5] ;
 wire \Tile_X1Y3_N2BEG[6] ;
 wire \Tile_X1Y3_N2BEG[7] ;
 wire \Tile_X1Y3_N2BEGb[0] ;
 wire \Tile_X1Y3_N2BEGb[1] ;
 wire \Tile_X1Y3_N2BEGb[2] ;
 wire \Tile_X1Y3_N2BEGb[3] ;
 wire \Tile_X1Y3_N2BEGb[4] ;
 wire \Tile_X1Y3_N2BEGb[5] ;
 wire \Tile_X1Y3_N2BEGb[6] ;
 wire \Tile_X1Y3_N2BEGb[7] ;
 wire \Tile_X1Y3_N4BEG[0] ;
 wire \Tile_X1Y3_N4BEG[10] ;
 wire \Tile_X1Y3_N4BEG[11] ;
 wire \Tile_X1Y3_N4BEG[12] ;
 wire \Tile_X1Y3_N4BEG[13] ;
 wire \Tile_X1Y3_N4BEG[14] ;
 wire \Tile_X1Y3_N4BEG[15] ;
 wire \Tile_X1Y3_N4BEG[1] ;
 wire \Tile_X1Y3_N4BEG[2] ;
 wire \Tile_X1Y3_N4BEG[3] ;
 wire \Tile_X1Y3_N4BEG[4] ;
 wire \Tile_X1Y3_N4BEG[5] ;
 wire \Tile_X1Y3_N4BEG[6] ;
 wire \Tile_X1Y3_N4BEG[7] ;
 wire \Tile_X1Y3_N4BEG[8] ;
 wire \Tile_X1Y3_N4BEG[9] ;
 wire \Tile_X1Y3_NN4BEG[0] ;
 wire \Tile_X1Y3_NN4BEG[10] ;
 wire \Tile_X1Y3_NN4BEG[11] ;
 wire \Tile_X1Y3_NN4BEG[12] ;
 wire \Tile_X1Y3_NN4BEG[13] ;
 wire \Tile_X1Y3_NN4BEG[14] ;
 wire \Tile_X1Y3_NN4BEG[15] ;
 wire \Tile_X1Y3_NN4BEG[1] ;
 wire \Tile_X1Y3_NN4BEG[2] ;
 wire \Tile_X1Y3_NN4BEG[3] ;
 wire \Tile_X1Y3_NN4BEG[4] ;
 wire \Tile_X1Y3_NN4BEG[5] ;
 wire \Tile_X1Y3_NN4BEG[6] ;
 wire \Tile_X1Y3_NN4BEG[7] ;
 wire \Tile_X1Y3_NN4BEG[8] ;
 wire \Tile_X1Y3_NN4BEG[9] ;
 wire \Tile_X1Y3_S1BEG[0] ;
 wire \Tile_X1Y3_S1BEG[1] ;
 wire \Tile_X1Y3_S1BEG[2] ;
 wire \Tile_X1Y3_S1BEG[3] ;
 wire \Tile_X1Y3_S2BEG[0] ;
 wire \Tile_X1Y3_S2BEG[1] ;
 wire \Tile_X1Y3_S2BEG[2] ;
 wire \Tile_X1Y3_S2BEG[3] ;
 wire \Tile_X1Y3_S2BEG[4] ;
 wire \Tile_X1Y3_S2BEG[5] ;
 wire \Tile_X1Y3_S2BEG[6] ;
 wire \Tile_X1Y3_S2BEG[7] ;
 wire \Tile_X1Y3_S2BEGb[0] ;
 wire \Tile_X1Y3_S2BEGb[1] ;
 wire \Tile_X1Y3_S2BEGb[2] ;
 wire \Tile_X1Y3_S2BEGb[3] ;
 wire \Tile_X1Y3_S2BEGb[4] ;
 wire \Tile_X1Y3_S2BEGb[5] ;
 wire \Tile_X1Y3_S2BEGb[6] ;
 wire \Tile_X1Y3_S2BEGb[7] ;
 wire \Tile_X1Y3_S4BEG[0] ;
 wire \Tile_X1Y3_S4BEG[10] ;
 wire \Tile_X1Y3_S4BEG[11] ;
 wire \Tile_X1Y3_S4BEG[12] ;
 wire \Tile_X1Y3_S4BEG[13] ;
 wire \Tile_X1Y3_S4BEG[14] ;
 wire \Tile_X1Y3_S4BEG[15] ;
 wire \Tile_X1Y3_S4BEG[1] ;
 wire \Tile_X1Y3_S4BEG[2] ;
 wire \Tile_X1Y3_S4BEG[3] ;
 wire \Tile_X1Y3_S4BEG[4] ;
 wire \Tile_X1Y3_S4BEG[5] ;
 wire \Tile_X1Y3_S4BEG[6] ;
 wire \Tile_X1Y3_S4BEG[7] ;
 wire \Tile_X1Y3_S4BEG[8] ;
 wire \Tile_X1Y3_S4BEG[9] ;
 wire \Tile_X1Y3_SS4BEG[0] ;
 wire \Tile_X1Y3_SS4BEG[10] ;
 wire \Tile_X1Y3_SS4BEG[11] ;
 wire \Tile_X1Y3_SS4BEG[12] ;
 wire \Tile_X1Y3_SS4BEG[13] ;
 wire \Tile_X1Y3_SS4BEG[14] ;
 wire \Tile_X1Y3_SS4BEG[15] ;
 wire \Tile_X1Y3_SS4BEG[1] ;
 wire \Tile_X1Y3_SS4BEG[2] ;
 wire \Tile_X1Y3_SS4BEG[3] ;
 wire \Tile_X1Y3_SS4BEG[4] ;
 wire \Tile_X1Y3_SS4BEG[5] ;
 wire \Tile_X1Y3_SS4BEG[6] ;
 wire \Tile_X1Y3_SS4BEG[7] ;
 wire \Tile_X1Y3_SS4BEG[8] ;
 wire \Tile_X1Y3_SS4BEG[9] ;
 wire Tile_X1Y3_UserCLKo;
 wire \Tile_X1Y3_W1BEG[0] ;
 wire \Tile_X1Y3_W1BEG[1] ;
 wire \Tile_X1Y3_W1BEG[2] ;
 wire \Tile_X1Y3_W1BEG[3] ;
 wire \Tile_X1Y3_W2BEG[0] ;
 wire \Tile_X1Y3_W2BEG[1] ;
 wire \Tile_X1Y3_W2BEG[2] ;
 wire \Tile_X1Y3_W2BEG[3] ;
 wire \Tile_X1Y3_W2BEG[4] ;
 wire \Tile_X1Y3_W2BEG[5] ;
 wire \Tile_X1Y3_W2BEG[6] ;
 wire \Tile_X1Y3_W2BEG[7] ;
 wire \Tile_X1Y3_W2BEGb[0] ;
 wire \Tile_X1Y3_W2BEGb[1] ;
 wire \Tile_X1Y3_W2BEGb[2] ;
 wire \Tile_X1Y3_W2BEGb[3] ;
 wire \Tile_X1Y3_W2BEGb[4] ;
 wire \Tile_X1Y3_W2BEGb[5] ;
 wire \Tile_X1Y3_W2BEGb[6] ;
 wire \Tile_X1Y3_W2BEGb[7] ;
 wire \Tile_X1Y3_W6BEG[0] ;
 wire \Tile_X1Y3_W6BEG[10] ;
 wire \Tile_X1Y3_W6BEG[11] ;
 wire \Tile_X1Y3_W6BEG[1] ;
 wire \Tile_X1Y3_W6BEG[2] ;
 wire \Tile_X1Y3_W6BEG[3] ;
 wire \Tile_X1Y3_W6BEG[4] ;
 wire \Tile_X1Y3_W6BEG[5] ;
 wire \Tile_X1Y3_W6BEG[6] ;
 wire \Tile_X1Y3_W6BEG[7] ;
 wire \Tile_X1Y3_W6BEG[8] ;
 wire \Tile_X1Y3_W6BEG[9] ;
 wire \Tile_X1Y3_WW4BEG[0] ;
 wire \Tile_X1Y3_WW4BEG[10] ;
 wire \Tile_X1Y3_WW4BEG[11] ;
 wire \Tile_X1Y3_WW4BEG[12] ;
 wire \Tile_X1Y3_WW4BEG[13] ;
 wire \Tile_X1Y3_WW4BEG[14] ;
 wire \Tile_X1Y3_WW4BEG[15] ;
 wire \Tile_X1Y3_WW4BEG[1] ;
 wire \Tile_X1Y3_WW4BEG[2] ;
 wire \Tile_X1Y3_WW4BEG[3] ;
 wire \Tile_X1Y3_WW4BEG[4] ;
 wire \Tile_X1Y3_WW4BEG[5] ;
 wire \Tile_X1Y3_WW4BEG[6] ;
 wire \Tile_X1Y3_WW4BEG[7] ;
 wire \Tile_X1Y3_WW4BEG[8] ;
 wire \Tile_X1Y3_WW4BEG[9] ;
 wire Tile_X1Y4_Co;
 wire \Tile_X1Y4_E1BEG[0] ;
 wire \Tile_X1Y4_E1BEG[1] ;
 wire \Tile_X1Y4_E1BEG[2] ;
 wire \Tile_X1Y4_E1BEG[3] ;
 wire \Tile_X1Y4_E2BEG[0] ;
 wire \Tile_X1Y4_E2BEG[1] ;
 wire \Tile_X1Y4_E2BEG[2] ;
 wire \Tile_X1Y4_E2BEG[3] ;
 wire \Tile_X1Y4_E2BEG[4] ;
 wire \Tile_X1Y4_E2BEG[5] ;
 wire \Tile_X1Y4_E2BEG[6] ;
 wire \Tile_X1Y4_E2BEG[7] ;
 wire \Tile_X1Y4_E2BEGb[0] ;
 wire \Tile_X1Y4_E2BEGb[1] ;
 wire \Tile_X1Y4_E2BEGb[2] ;
 wire \Tile_X1Y4_E2BEGb[3] ;
 wire \Tile_X1Y4_E2BEGb[4] ;
 wire \Tile_X1Y4_E2BEGb[5] ;
 wire \Tile_X1Y4_E2BEGb[6] ;
 wire \Tile_X1Y4_E2BEGb[7] ;
 wire \Tile_X1Y4_E6BEG[0] ;
 wire \Tile_X1Y4_E6BEG[10] ;
 wire \Tile_X1Y4_E6BEG[11] ;
 wire \Tile_X1Y4_E6BEG[1] ;
 wire \Tile_X1Y4_E6BEG[2] ;
 wire \Tile_X1Y4_E6BEG[3] ;
 wire \Tile_X1Y4_E6BEG[4] ;
 wire \Tile_X1Y4_E6BEG[5] ;
 wire \Tile_X1Y4_E6BEG[6] ;
 wire \Tile_X1Y4_E6BEG[7] ;
 wire \Tile_X1Y4_E6BEG[8] ;
 wire \Tile_X1Y4_E6BEG[9] ;
 wire \Tile_X1Y4_EE4BEG[0] ;
 wire \Tile_X1Y4_EE4BEG[10] ;
 wire \Tile_X1Y4_EE4BEG[11] ;
 wire \Tile_X1Y4_EE4BEG[12] ;
 wire \Tile_X1Y4_EE4BEG[13] ;
 wire \Tile_X1Y4_EE4BEG[14] ;
 wire \Tile_X1Y4_EE4BEG[15] ;
 wire \Tile_X1Y4_EE4BEG[1] ;
 wire \Tile_X1Y4_EE4BEG[2] ;
 wire \Tile_X1Y4_EE4BEG[3] ;
 wire \Tile_X1Y4_EE4BEG[4] ;
 wire \Tile_X1Y4_EE4BEG[5] ;
 wire \Tile_X1Y4_EE4BEG[6] ;
 wire \Tile_X1Y4_EE4BEG[7] ;
 wire \Tile_X1Y4_EE4BEG[8] ;
 wire \Tile_X1Y4_EE4BEG[9] ;
 wire \Tile_X1Y4_FrameData_O[0] ;
 wire \Tile_X1Y4_FrameData_O[10] ;
 wire \Tile_X1Y4_FrameData_O[11] ;
 wire \Tile_X1Y4_FrameData_O[12] ;
 wire \Tile_X1Y4_FrameData_O[13] ;
 wire \Tile_X1Y4_FrameData_O[14] ;
 wire \Tile_X1Y4_FrameData_O[15] ;
 wire \Tile_X1Y4_FrameData_O[16] ;
 wire \Tile_X1Y4_FrameData_O[17] ;
 wire \Tile_X1Y4_FrameData_O[18] ;
 wire \Tile_X1Y4_FrameData_O[19] ;
 wire \Tile_X1Y4_FrameData_O[1] ;
 wire \Tile_X1Y4_FrameData_O[20] ;
 wire \Tile_X1Y4_FrameData_O[21] ;
 wire \Tile_X1Y4_FrameData_O[22] ;
 wire \Tile_X1Y4_FrameData_O[23] ;
 wire \Tile_X1Y4_FrameData_O[24] ;
 wire \Tile_X1Y4_FrameData_O[25] ;
 wire \Tile_X1Y4_FrameData_O[26] ;
 wire \Tile_X1Y4_FrameData_O[27] ;
 wire \Tile_X1Y4_FrameData_O[28] ;
 wire \Tile_X1Y4_FrameData_O[29] ;
 wire \Tile_X1Y4_FrameData_O[2] ;
 wire \Tile_X1Y4_FrameData_O[30] ;
 wire \Tile_X1Y4_FrameData_O[31] ;
 wire \Tile_X1Y4_FrameData_O[3] ;
 wire \Tile_X1Y4_FrameData_O[4] ;
 wire \Tile_X1Y4_FrameData_O[5] ;
 wire \Tile_X1Y4_FrameData_O[6] ;
 wire \Tile_X1Y4_FrameData_O[7] ;
 wire \Tile_X1Y4_FrameData_O[8] ;
 wire \Tile_X1Y4_FrameData_O[9] ;
 wire \Tile_X1Y4_FrameStrobe_O[0] ;
 wire \Tile_X1Y4_FrameStrobe_O[10] ;
 wire \Tile_X1Y4_FrameStrobe_O[11] ;
 wire \Tile_X1Y4_FrameStrobe_O[12] ;
 wire \Tile_X1Y4_FrameStrobe_O[13] ;
 wire \Tile_X1Y4_FrameStrobe_O[14] ;
 wire \Tile_X1Y4_FrameStrobe_O[15] ;
 wire \Tile_X1Y4_FrameStrobe_O[16] ;
 wire \Tile_X1Y4_FrameStrobe_O[17] ;
 wire \Tile_X1Y4_FrameStrobe_O[18] ;
 wire \Tile_X1Y4_FrameStrobe_O[19] ;
 wire \Tile_X1Y4_FrameStrobe_O[1] ;
 wire \Tile_X1Y4_FrameStrobe_O[2] ;
 wire \Tile_X1Y4_FrameStrobe_O[3] ;
 wire \Tile_X1Y4_FrameStrobe_O[4] ;
 wire \Tile_X1Y4_FrameStrobe_O[5] ;
 wire \Tile_X1Y4_FrameStrobe_O[6] ;
 wire \Tile_X1Y4_FrameStrobe_O[7] ;
 wire \Tile_X1Y4_FrameStrobe_O[8] ;
 wire \Tile_X1Y4_FrameStrobe_O[9] ;
 wire \Tile_X1Y4_N1BEG[0] ;
 wire \Tile_X1Y4_N1BEG[1] ;
 wire \Tile_X1Y4_N1BEG[2] ;
 wire \Tile_X1Y4_N1BEG[3] ;
 wire \Tile_X1Y4_N2BEG[0] ;
 wire \Tile_X1Y4_N2BEG[1] ;
 wire \Tile_X1Y4_N2BEG[2] ;
 wire \Tile_X1Y4_N2BEG[3] ;
 wire \Tile_X1Y4_N2BEG[4] ;
 wire \Tile_X1Y4_N2BEG[5] ;
 wire \Tile_X1Y4_N2BEG[6] ;
 wire \Tile_X1Y4_N2BEG[7] ;
 wire \Tile_X1Y4_N2BEGb[0] ;
 wire \Tile_X1Y4_N2BEGb[1] ;
 wire \Tile_X1Y4_N2BEGb[2] ;
 wire \Tile_X1Y4_N2BEGb[3] ;
 wire \Tile_X1Y4_N2BEGb[4] ;
 wire \Tile_X1Y4_N2BEGb[5] ;
 wire \Tile_X1Y4_N2BEGb[6] ;
 wire \Tile_X1Y4_N2BEGb[7] ;
 wire \Tile_X1Y4_N4BEG[0] ;
 wire \Tile_X1Y4_N4BEG[10] ;
 wire \Tile_X1Y4_N4BEG[11] ;
 wire \Tile_X1Y4_N4BEG[12] ;
 wire \Tile_X1Y4_N4BEG[13] ;
 wire \Tile_X1Y4_N4BEG[14] ;
 wire \Tile_X1Y4_N4BEG[15] ;
 wire \Tile_X1Y4_N4BEG[1] ;
 wire \Tile_X1Y4_N4BEG[2] ;
 wire \Tile_X1Y4_N4BEG[3] ;
 wire \Tile_X1Y4_N4BEG[4] ;
 wire \Tile_X1Y4_N4BEG[5] ;
 wire \Tile_X1Y4_N4BEG[6] ;
 wire \Tile_X1Y4_N4BEG[7] ;
 wire \Tile_X1Y4_N4BEG[8] ;
 wire \Tile_X1Y4_N4BEG[9] ;
 wire \Tile_X1Y4_NN4BEG[0] ;
 wire \Tile_X1Y4_NN4BEG[10] ;
 wire \Tile_X1Y4_NN4BEG[11] ;
 wire \Tile_X1Y4_NN4BEG[12] ;
 wire \Tile_X1Y4_NN4BEG[13] ;
 wire \Tile_X1Y4_NN4BEG[14] ;
 wire \Tile_X1Y4_NN4BEG[15] ;
 wire \Tile_X1Y4_NN4BEG[1] ;
 wire \Tile_X1Y4_NN4BEG[2] ;
 wire \Tile_X1Y4_NN4BEG[3] ;
 wire \Tile_X1Y4_NN4BEG[4] ;
 wire \Tile_X1Y4_NN4BEG[5] ;
 wire \Tile_X1Y4_NN4BEG[6] ;
 wire \Tile_X1Y4_NN4BEG[7] ;
 wire \Tile_X1Y4_NN4BEG[8] ;
 wire \Tile_X1Y4_NN4BEG[9] ;
 wire \Tile_X1Y4_S1BEG[0] ;
 wire \Tile_X1Y4_S1BEG[1] ;
 wire \Tile_X1Y4_S1BEG[2] ;
 wire \Tile_X1Y4_S1BEG[3] ;
 wire \Tile_X1Y4_S2BEG[0] ;
 wire \Tile_X1Y4_S2BEG[1] ;
 wire \Tile_X1Y4_S2BEG[2] ;
 wire \Tile_X1Y4_S2BEG[3] ;
 wire \Tile_X1Y4_S2BEG[4] ;
 wire \Tile_X1Y4_S2BEG[5] ;
 wire \Tile_X1Y4_S2BEG[6] ;
 wire \Tile_X1Y4_S2BEG[7] ;
 wire \Tile_X1Y4_S2BEGb[0] ;
 wire \Tile_X1Y4_S2BEGb[1] ;
 wire \Tile_X1Y4_S2BEGb[2] ;
 wire \Tile_X1Y4_S2BEGb[3] ;
 wire \Tile_X1Y4_S2BEGb[4] ;
 wire \Tile_X1Y4_S2BEGb[5] ;
 wire \Tile_X1Y4_S2BEGb[6] ;
 wire \Tile_X1Y4_S2BEGb[7] ;
 wire \Tile_X1Y4_S4BEG[0] ;
 wire \Tile_X1Y4_S4BEG[10] ;
 wire \Tile_X1Y4_S4BEG[11] ;
 wire \Tile_X1Y4_S4BEG[12] ;
 wire \Tile_X1Y4_S4BEG[13] ;
 wire \Tile_X1Y4_S4BEG[14] ;
 wire \Tile_X1Y4_S4BEG[15] ;
 wire \Tile_X1Y4_S4BEG[1] ;
 wire \Tile_X1Y4_S4BEG[2] ;
 wire \Tile_X1Y4_S4BEG[3] ;
 wire \Tile_X1Y4_S4BEG[4] ;
 wire \Tile_X1Y4_S4BEG[5] ;
 wire \Tile_X1Y4_S4BEG[6] ;
 wire \Tile_X1Y4_S4BEG[7] ;
 wire \Tile_X1Y4_S4BEG[8] ;
 wire \Tile_X1Y4_S4BEG[9] ;
 wire \Tile_X1Y4_SS4BEG[0] ;
 wire \Tile_X1Y4_SS4BEG[10] ;
 wire \Tile_X1Y4_SS4BEG[11] ;
 wire \Tile_X1Y4_SS4BEG[12] ;
 wire \Tile_X1Y4_SS4BEG[13] ;
 wire \Tile_X1Y4_SS4BEG[14] ;
 wire \Tile_X1Y4_SS4BEG[15] ;
 wire \Tile_X1Y4_SS4BEG[1] ;
 wire \Tile_X1Y4_SS4BEG[2] ;
 wire \Tile_X1Y4_SS4BEG[3] ;
 wire \Tile_X1Y4_SS4BEG[4] ;
 wire \Tile_X1Y4_SS4BEG[5] ;
 wire \Tile_X1Y4_SS4BEG[6] ;
 wire \Tile_X1Y4_SS4BEG[7] ;
 wire \Tile_X1Y4_SS4BEG[8] ;
 wire \Tile_X1Y4_SS4BEG[9] ;
 wire Tile_X1Y4_UserCLKo;
 wire \Tile_X1Y4_W1BEG[0] ;
 wire \Tile_X1Y4_W1BEG[1] ;
 wire \Tile_X1Y4_W1BEG[2] ;
 wire \Tile_X1Y4_W1BEG[3] ;
 wire \Tile_X1Y4_W2BEG[0] ;
 wire \Tile_X1Y4_W2BEG[1] ;
 wire \Tile_X1Y4_W2BEG[2] ;
 wire \Tile_X1Y4_W2BEG[3] ;
 wire \Tile_X1Y4_W2BEG[4] ;
 wire \Tile_X1Y4_W2BEG[5] ;
 wire \Tile_X1Y4_W2BEG[6] ;
 wire \Tile_X1Y4_W2BEG[7] ;
 wire \Tile_X1Y4_W2BEGb[0] ;
 wire \Tile_X1Y4_W2BEGb[1] ;
 wire \Tile_X1Y4_W2BEGb[2] ;
 wire \Tile_X1Y4_W2BEGb[3] ;
 wire \Tile_X1Y4_W2BEGb[4] ;
 wire \Tile_X1Y4_W2BEGb[5] ;
 wire \Tile_X1Y4_W2BEGb[6] ;
 wire \Tile_X1Y4_W2BEGb[7] ;
 wire \Tile_X1Y4_W6BEG[0] ;
 wire \Tile_X1Y4_W6BEG[10] ;
 wire \Tile_X1Y4_W6BEG[11] ;
 wire \Tile_X1Y4_W6BEG[1] ;
 wire \Tile_X1Y4_W6BEG[2] ;
 wire \Tile_X1Y4_W6BEG[3] ;
 wire \Tile_X1Y4_W6BEG[4] ;
 wire \Tile_X1Y4_W6BEG[5] ;
 wire \Tile_X1Y4_W6BEG[6] ;
 wire \Tile_X1Y4_W6BEG[7] ;
 wire \Tile_X1Y4_W6BEG[8] ;
 wire \Tile_X1Y4_W6BEG[9] ;
 wire \Tile_X1Y4_WW4BEG[0] ;
 wire \Tile_X1Y4_WW4BEG[10] ;
 wire \Tile_X1Y4_WW4BEG[11] ;
 wire \Tile_X1Y4_WW4BEG[12] ;
 wire \Tile_X1Y4_WW4BEG[13] ;
 wire \Tile_X1Y4_WW4BEG[14] ;
 wire \Tile_X1Y4_WW4BEG[15] ;
 wire \Tile_X1Y4_WW4BEG[1] ;
 wire \Tile_X1Y4_WW4BEG[2] ;
 wire \Tile_X1Y4_WW4BEG[3] ;
 wire \Tile_X1Y4_WW4BEG[4] ;
 wire \Tile_X1Y4_WW4BEG[5] ;
 wire \Tile_X1Y4_WW4BEG[6] ;
 wire \Tile_X1Y4_WW4BEG[7] ;
 wire \Tile_X1Y4_WW4BEG[8] ;
 wire \Tile_X1Y4_WW4BEG[9] ;
 wire Tile_X1Y5_Co;
 wire \Tile_X1Y5_E1BEG[0] ;
 wire \Tile_X1Y5_E1BEG[1] ;
 wire \Tile_X1Y5_E1BEG[2] ;
 wire \Tile_X1Y5_E1BEG[3] ;
 wire \Tile_X1Y5_E2BEG[0] ;
 wire \Tile_X1Y5_E2BEG[1] ;
 wire \Tile_X1Y5_E2BEG[2] ;
 wire \Tile_X1Y5_E2BEG[3] ;
 wire \Tile_X1Y5_E2BEG[4] ;
 wire \Tile_X1Y5_E2BEG[5] ;
 wire \Tile_X1Y5_E2BEG[6] ;
 wire \Tile_X1Y5_E2BEG[7] ;
 wire \Tile_X1Y5_E2BEGb[0] ;
 wire \Tile_X1Y5_E2BEGb[1] ;
 wire \Tile_X1Y5_E2BEGb[2] ;
 wire \Tile_X1Y5_E2BEGb[3] ;
 wire \Tile_X1Y5_E2BEGb[4] ;
 wire \Tile_X1Y5_E2BEGb[5] ;
 wire \Tile_X1Y5_E2BEGb[6] ;
 wire \Tile_X1Y5_E2BEGb[7] ;
 wire \Tile_X1Y5_E6BEG[0] ;
 wire \Tile_X1Y5_E6BEG[10] ;
 wire \Tile_X1Y5_E6BEG[11] ;
 wire \Tile_X1Y5_E6BEG[1] ;
 wire \Tile_X1Y5_E6BEG[2] ;
 wire \Tile_X1Y5_E6BEG[3] ;
 wire \Tile_X1Y5_E6BEG[4] ;
 wire \Tile_X1Y5_E6BEG[5] ;
 wire \Tile_X1Y5_E6BEG[6] ;
 wire \Tile_X1Y5_E6BEG[7] ;
 wire \Tile_X1Y5_E6BEG[8] ;
 wire \Tile_X1Y5_E6BEG[9] ;
 wire \Tile_X1Y5_EE4BEG[0] ;
 wire \Tile_X1Y5_EE4BEG[10] ;
 wire \Tile_X1Y5_EE4BEG[11] ;
 wire \Tile_X1Y5_EE4BEG[12] ;
 wire \Tile_X1Y5_EE4BEG[13] ;
 wire \Tile_X1Y5_EE4BEG[14] ;
 wire \Tile_X1Y5_EE4BEG[15] ;
 wire \Tile_X1Y5_EE4BEG[1] ;
 wire \Tile_X1Y5_EE4BEG[2] ;
 wire \Tile_X1Y5_EE4BEG[3] ;
 wire \Tile_X1Y5_EE4BEG[4] ;
 wire \Tile_X1Y5_EE4BEG[5] ;
 wire \Tile_X1Y5_EE4BEG[6] ;
 wire \Tile_X1Y5_EE4BEG[7] ;
 wire \Tile_X1Y5_EE4BEG[8] ;
 wire \Tile_X1Y5_EE4BEG[9] ;
 wire \Tile_X1Y5_FrameData_O[0] ;
 wire \Tile_X1Y5_FrameData_O[10] ;
 wire \Tile_X1Y5_FrameData_O[11] ;
 wire \Tile_X1Y5_FrameData_O[12] ;
 wire \Tile_X1Y5_FrameData_O[13] ;
 wire \Tile_X1Y5_FrameData_O[14] ;
 wire \Tile_X1Y5_FrameData_O[15] ;
 wire \Tile_X1Y5_FrameData_O[16] ;
 wire \Tile_X1Y5_FrameData_O[17] ;
 wire \Tile_X1Y5_FrameData_O[18] ;
 wire \Tile_X1Y5_FrameData_O[19] ;
 wire \Tile_X1Y5_FrameData_O[1] ;
 wire \Tile_X1Y5_FrameData_O[20] ;
 wire \Tile_X1Y5_FrameData_O[21] ;
 wire \Tile_X1Y5_FrameData_O[22] ;
 wire \Tile_X1Y5_FrameData_O[23] ;
 wire \Tile_X1Y5_FrameData_O[24] ;
 wire \Tile_X1Y5_FrameData_O[25] ;
 wire \Tile_X1Y5_FrameData_O[26] ;
 wire \Tile_X1Y5_FrameData_O[27] ;
 wire \Tile_X1Y5_FrameData_O[28] ;
 wire \Tile_X1Y5_FrameData_O[29] ;
 wire \Tile_X1Y5_FrameData_O[2] ;
 wire \Tile_X1Y5_FrameData_O[30] ;
 wire \Tile_X1Y5_FrameData_O[31] ;
 wire \Tile_X1Y5_FrameData_O[3] ;
 wire \Tile_X1Y5_FrameData_O[4] ;
 wire \Tile_X1Y5_FrameData_O[5] ;
 wire \Tile_X1Y5_FrameData_O[6] ;
 wire \Tile_X1Y5_FrameData_O[7] ;
 wire \Tile_X1Y5_FrameData_O[8] ;
 wire \Tile_X1Y5_FrameData_O[9] ;
 wire \Tile_X1Y5_FrameStrobe_O[0] ;
 wire \Tile_X1Y5_FrameStrobe_O[10] ;
 wire \Tile_X1Y5_FrameStrobe_O[11] ;
 wire \Tile_X1Y5_FrameStrobe_O[12] ;
 wire \Tile_X1Y5_FrameStrobe_O[13] ;
 wire \Tile_X1Y5_FrameStrobe_O[14] ;
 wire \Tile_X1Y5_FrameStrobe_O[15] ;
 wire \Tile_X1Y5_FrameStrobe_O[16] ;
 wire \Tile_X1Y5_FrameStrobe_O[17] ;
 wire \Tile_X1Y5_FrameStrobe_O[18] ;
 wire \Tile_X1Y5_FrameStrobe_O[19] ;
 wire \Tile_X1Y5_FrameStrobe_O[1] ;
 wire \Tile_X1Y5_FrameStrobe_O[2] ;
 wire \Tile_X1Y5_FrameStrobe_O[3] ;
 wire \Tile_X1Y5_FrameStrobe_O[4] ;
 wire \Tile_X1Y5_FrameStrobe_O[5] ;
 wire \Tile_X1Y5_FrameStrobe_O[6] ;
 wire \Tile_X1Y5_FrameStrobe_O[7] ;
 wire \Tile_X1Y5_FrameStrobe_O[8] ;
 wire \Tile_X1Y5_FrameStrobe_O[9] ;
 wire \Tile_X1Y5_N1BEG[0] ;
 wire \Tile_X1Y5_N1BEG[1] ;
 wire \Tile_X1Y5_N1BEG[2] ;
 wire \Tile_X1Y5_N1BEG[3] ;
 wire \Tile_X1Y5_N2BEG[0] ;
 wire \Tile_X1Y5_N2BEG[1] ;
 wire \Tile_X1Y5_N2BEG[2] ;
 wire \Tile_X1Y5_N2BEG[3] ;
 wire \Tile_X1Y5_N2BEG[4] ;
 wire \Tile_X1Y5_N2BEG[5] ;
 wire \Tile_X1Y5_N2BEG[6] ;
 wire \Tile_X1Y5_N2BEG[7] ;
 wire \Tile_X1Y5_N2BEGb[0] ;
 wire \Tile_X1Y5_N2BEGb[1] ;
 wire \Tile_X1Y5_N2BEGb[2] ;
 wire \Tile_X1Y5_N2BEGb[3] ;
 wire \Tile_X1Y5_N2BEGb[4] ;
 wire \Tile_X1Y5_N2BEGb[5] ;
 wire \Tile_X1Y5_N2BEGb[6] ;
 wire \Tile_X1Y5_N2BEGb[7] ;
 wire \Tile_X1Y5_N4BEG[0] ;
 wire \Tile_X1Y5_N4BEG[10] ;
 wire \Tile_X1Y5_N4BEG[11] ;
 wire \Tile_X1Y5_N4BEG[12] ;
 wire \Tile_X1Y5_N4BEG[13] ;
 wire \Tile_X1Y5_N4BEG[14] ;
 wire \Tile_X1Y5_N4BEG[15] ;
 wire \Tile_X1Y5_N4BEG[1] ;
 wire \Tile_X1Y5_N4BEG[2] ;
 wire \Tile_X1Y5_N4BEG[3] ;
 wire \Tile_X1Y5_N4BEG[4] ;
 wire \Tile_X1Y5_N4BEG[5] ;
 wire \Tile_X1Y5_N4BEG[6] ;
 wire \Tile_X1Y5_N4BEG[7] ;
 wire \Tile_X1Y5_N4BEG[8] ;
 wire \Tile_X1Y5_N4BEG[9] ;
 wire \Tile_X1Y5_NN4BEG[0] ;
 wire \Tile_X1Y5_NN4BEG[10] ;
 wire \Tile_X1Y5_NN4BEG[11] ;
 wire \Tile_X1Y5_NN4BEG[12] ;
 wire \Tile_X1Y5_NN4BEG[13] ;
 wire \Tile_X1Y5_NN4BEG[14] ;
 wire \Tile_X1Y5_NN4BEG[15] ;
 wire \Tile_X1Y5_NN4BEG[1] ;
 wire \Tile_X1Y5_NN4BEG[2] ;
 wire \Tile_X1Y5_NN4BEG[3] ;
 wire \Tile_X1Y5_NN4BEG[4] ;
 wire \Tile_X1Y5_NN4BEG[5] ;
 wire \Tile_X1Y5_NN4BEG[6] ;
 wire \Tile_X1Y5_NN4BEG[7] ;
 wire \Tile_X1Y5_NN4BEG[8] ;
 wire \Tile_X1Y5_NN4BEG[9] ;
 wire \Tile_X1Y5_S1BEG[0] ;
 wire \Tile_X1Y5_S1BEG[1] ;
 wire \Tile_X1Y5_S1BEG[2] ;
 wire \Tile_X1Y5_S1BEG[3] ;
 wire \Tile_X1Y5_S2BEG[0] ;
 wire \Tile_X1Y5_S2BEG[1] ;
 wire \Tile_X1Y5_S2BEG[2] ;
 wire \Tile_X1Y5_S2BEG[3] ;
 wire \Tile_X1Y5_S2BEG[4] ;
 wire \Tile_X1Y5_S2BEG[5] ;
 wire \Tile_X1Y5_S2BEG[6] ;
 wire \Tile_X1Y5_S2BEG[7] ;
 wire \Tile_X1Y5_S2BEGb[0] ;
 wire \Tile_X1Y5_S2BEGb[1] ;
 wire \Tile_X1Y5_S2BEGb[2] ;
 wire \Tile_X1Y5_S2BEGb[3] ;
 wire \Tile_X1Y5_S2BEGb[4] ;
 wire \Tile_X1Y5_S2BEGb[5] ;
 wire \Tile_X1Y5_S2BEGb[6] ;
 wire \Tile_X1Y5_S2BEGb[7] ;
 wire \Tile_X1Y5_S4BEG[0] ;
 wire \Tile_X1Y5_S4BEG[10] ;
 wire \Tile_X1Y5_S4BEG[11] ;
 wire \Tile_X1Y5_S4BEG[12] ;
 wire \Tile_X1Y5_S4BEG[13] ;
 wire \Tile_X1Y5_S4BEG[14] ;
 wire \Tile_X1Y5_S4BEG[15] ;
 wire \Tile_X1Y5_S4BEG[1] ;
 wire \Tile_X1Y5_S4BEG[2] ;
 wire \Tile_X1Y5_S4BEG[3] ;
 wire \Tile_X1Y5_S4BEG[4] ;
 wire \Tile_X1Y5_S4BEG[5] ;
 wire \Tile_X1Y5_S4BEG[6] ;
 wire \Tile_X1Y5_S4BEG[7] ;
 wire \Tile_X1Y5_S4BEG[8] ;
 wire \Tile_X1Y5_S4BEG[9] ;
 wire \Tile_X1Y5_SS4BEG[0] ;
 wire \Tile_X1Y5_SS4BEG[10] ;
 wire \Tile_X1Y5_SS4BEG[11] ;
 wire \Tile_X1Y5_SS4BEG[12] ;
 wire \Tile_X1Y5_SS4BEG[13] ;
 wire \Tile_X1Y5_SS4BEG[14] ;
 wire \Tile_X1Y5_SS4BEG[15] ;
 wire \Tile_X1Y5_SS4BEG[1] ;
 wire \Tile_X1Y5_SS4BEG[2] ;
 wire \Tile_X1Y5_SS4BEG[3] ;
 wire \Tile_X1Y5_SS4BEG[4] ;
 wire \Tile_X1Y5_SS4BEG[5] ;
 wire \Tile_X1Y5_SS4BEG[6] ;
 wire \Tile_X1Y5_SS4BEG[7] ;
 wire \Tile_X1Y5_SS4BEG[8] ;
 wire \Tile_X1Y5_SS4BEG[9] ;
 wire Tile_X1Y5_UserCLKo;
 wire \Tile_X1Y5_W1BEG[0] ;
 wire \Tile_X1Y5_W1BEG[1] ;
 wire \Tile_X1Y5_W1BEG[2] ;
 wire \Tile_X1Y5_W1BEG[3] ;
 wire \Tile_X1Y5_W2BEG[0] ;
 wire \Tile_X1Y5_W2BEG[1] ;
 wire \Tile_X1Y5_W2BEG[2] ;
 wire \Tile_X1Y5_W2BEG[3] ;
 wire \Tile_X1Y5_W2BEG[4] ;
 wire \Tile_X1Y5_W2BEG[5] ;
 wire \Tile_X1Y5_W2BEG[6] ;
 wire \Tile_X1Y5_W2BEG[7] ;
 wire \Tile_X1Y5_W2BEGb[0] ;
 wire \Tile_X1Y5_W2BEGb[1] ;
 wire \Tile_X1Y5_W2BEGb[2] ;
 wire \Tile_X1Y5_W2BEGb[3] ;
 wire \Tile_X1Y5_W2BEGb[4] ;
 wire \Tile_X1Y5_W2BEGb[5] ;
 wire \Tile_X1Y5_W2BEGb[6] ;
 wire \Tile_X1Y5_W2BEGb[7] ;
 wire \Tile_X1Y5_W6BEG[0] ;
 wire \Tile_X1Y5_W6BEG[10] ;
 wire \Tile_X1Y5_W6BEG[11] ;
 wire \Tile_X1Y5_W6BEG[1] ;
 wire \Tile_X1Y5_W6BEG[2] ;
 wire \Tile_X1Y5_W6BEG[3] ;
 wire \Tile_X1Y5_W6BEG[4] ;
 wire \Tile_X1Y5_W6BEG[5] ;
 wire \Tile_X1Y5_W6BEG[6] ;
 wire \Tile_X1Y5_W6BEG[7] ;
 wire \Tile_X1Y5_W6BEG[8] ;
 wire \Tile_X1Y5_W6BEG[9] ;
 wire \Tile_X1Y5_WW4BEG[0] ;
 wire \Tile_X1Y5_WW4BEG[10] ;
 wire \Tile_X1Y5_WW4BEG[11] ;
 wire \Tile_X1Y5_WW4BEG[12] ;
 wire \Tile_X1Y5_WW4BEG[13] ;
 wire \Tile_X1Y5_WW4BEG[14] ;
 wire \Tile_X1Y5_WW4BEG[15] ;
 wire \Tile_X1Y5_WW4BEG[1] ;
 wire \Tile_X1Y5_WW4BEG[2] ;
 wire \Tile_X1Y5_WW4BEG[3] ;
 wire \Tile_X1Y5_WW4BEG[4] ;
 wire \Tile_X1Y5_WW4BEG[5] ;
 wire \Tile_X1Y5_WW4BEG[6] ;
 wire \Tile_X1Y5_WW4BEG[7] ;
 wire \Tile_X1Y5_WW4BEG[8] ;
 wire \Tile_X1Y5_WW4BEG[9] ;
 wire Tile_X1Y6_Co;
 wire \Tile_X1Y6_E1BEG[0] ;
 wire \Tile_X1Y6_E1BEG[1] ;
 wire \Tile_X1Y6_E1BEG[2] ;
 wire \Tile_X1Y6_E1BEG[3] ;
 wire \Tile_X1Y6_E2BEG[0] ;
 wire \Tile_X1Y6_E2BEG[1] ;
 wire \Tile_X1Y6_E2BEG[2] ;
 wire \Tile_X1Y6_E2BEG[3] ;
 wire \Tile_X1Y6_E2BEG[4] ;
 wire \Tile_X1Y6_E2BEG[5] ;
 wire \Tile_X1Y6_E2BEG[6] ;
 wire \Tile_X1Y6_E2BEG[7] ;
 wire \Tile_X1Y6_E2BEGb[0] ;
 wire \Tile_X1Y6_E2BEGb[1] ;
 wire \Tile_X1Y6_E2BEGb[2] ;
 wire \Tile_X1Y6_E2BEGb[3] ;
 wire \Tile_X1Y6_E2BEGb[4] ;
 wire \Tile_X1Y6_E2BEGb[5] ;
 wire \Tile_X1Y6_E2BEGb[6] ;
 wire \Tile_X1Y6_E2BEGb[7] ;
 wire \Tile_X1Y6_E6BEG[0] ;
 wire \Tile_X1Y6_E6BEG[10] ;
 wire \Tile_X1Y6_E6BEG[11] ;
 wire \Tile_X1Y6_E6BEG[1] ;
 wire \Tile_X1Y6_E6BEG[2] ;
 wire \Tile_X1Y6_E6BEG[3] ;
 wire \Tile_X1Y6_E6BEG[4] ;
 wire \Tile_X1Y6_E6BEG[5] ;
 wire \Tile_X1Y6_E6BEG[6] ;
 wire \Tile_X1Y6_E6BEG[7] ;
 wire \Tile_X1Y6_E6BEG[8] ;
 wire \Tile_X1Y6_E6BEG[9] ;
 wire \Tile_X1Y6_EE4BEG[0] ;
 wire \Tile_X1Y6_EE4BEG[10] ;
 wire \Tile_X1Y6_EE4BEG[11] ;
 wire \Tile_X1Y6_EE4BEG[12] ;
 wire \Tile_X1Y6_EE4BEG[13] ;
 wire \Tile_X1Y6_EE4BEG[14] ;
 wire \Tile_X1Y6_EE4BEG[15] ;
 wire \Tile_X1Y6_EE4BEG[1] ;
 wire \Tile_X1Y6_EE4BEG[2] ;
 wire \Tile_X1Y6_EE4BEG[3] ;
 wire \Tile_X1Y6_EE4BEG[4] ;
 wire \Tile_X1Y6_EE4BEG[5] ;
 wire \Tile_X1Y6_EE4BEG[6] ;
 wire \Tile_X1Y6_EE4BEG[7] ;
 wire \Tile_X1Y6_EE4BEG[8] ;
 wire \Tile_X1Y6_EE4BEG[9] ;
 wire \Tile_X1Y6_FrameData_O[0] ;
 wire \Tile_X1Y6_FrameData_O[10] ;
 wire \Tile_X1Y6_FrameData_O[11] ;
 wire \Tile_X1Y6_FrameData_O[12] ;
 wire \Tile_X1Y6_FrameData_O[13] ;
 wire \Tile_X1Y6_FrameData_O[14] ;
 wire \Tile_X1Y6_FrameData_O[15] ;
 wire \Tile_X1Y6_FrameData_O[16] ;
 wire \Tile_X1Y6_FrameData_O[17] ;
 wire \Tile_X1Y6_FrameData_O[18] ;
 wire \Tile_X1Y6_FrameData_O[19] ;
 wire \Tile_X1Y6_FrameData_O[1] ;
 wire \Tile_X1Y6_FrameData_O[20] ;
 wire \Tile_X1Y6_FrameData_O[21] ;
 wire \Tile_X1Y6_FrameData_O[22] ;
 wire \Tile_X1Y6_FrameData_O[23] ;
 wire \Tile_X1Y6_FrameData_O[24] ;
 wire \Tile_X1Y6_FrameData_O[25] ;
 wire \Tile_X1Y6_FrameData_O[26] ;
 wire \Tile_X1Y6_FrameData_O[27] ;
 wire \Tile_X1Y6_FrameData_O[28] ;
 wire \Tile_X1Y6_FrameData_O[29] ;
 wire \Tile_X1Y6_FrameData_O[2] ;
 wire \Tile_X1Y6_FrameData_O[30] ;
 wire \Tile_X1Y6_FrameData_O[31] ;
 wire \Tile_X1Y6_FrameData_O[3] ;
 wire \Tile_X1Y6_FrameData_O[4] ;
 wire \Tile_X1Y6_FrameData_O[5] ;
 wire \Tile_X1Y6_FrameData_O[6] ;
 wire \Tile_X1Y6_FrameData_O[7] ;
 wire \Tile_X1Y6_FrameData_O[8] ;
 wire \Tile_X1Y6_FrameData_O[9] ;
 wire \Tile_X1Y6_FrameStrobe_O[0] ;
 wire \Tile_X1Y6_FrameStrobe_O[10] ;
 wire \Tile_X1Y6_FrameStrobe_O[11] ;
 wire \Tile_X1Y6_FrameStrobe_O[12] ;
 wire \Tile_X1Y6_FrameStrobe_O[13] ;
 wire \Tile_X1Y6_FrameStrobe_O[14] ;
 wire \Tile_X1Y6_FrameStrobe_O[15] ;
 wire \Tile_X1Y6_FrameStrobe_O[16] ;
 wire \Tile_X1Y6_FrameStrobe_O[17] ;
 wire \Tile_X1Y6_FrameStrobe_O[18] ;
 wire \Tile_X1Y6_FrameStrobe_O[19] ;
 wire \Tile_X1Y6_FrameStrobe_O[1] ;
 wire \Tile_X1Y6_FrameStrobe_O[2] ;
 wire \Tile_X1Y6_FrameStrobe_O[3] ;
 wire \Tile_X1Y6_FrameStrobe_O[4] ;
 wire \Tile_X1Y6_FrameStrobe_O[5] ;
 wire \Tile_X1Y6_FrameStrobe_O[6] ;
 wire \Tile_X1Y6_FrameStrobe_O[7] ;
 wire \Tile_X1Y6_FrameStrobe_O[8] ;
 wire \Tile_X1Y6_FrameStrobe_O[9] ;
 wire \Tile_X1Y6_N1BEG[0] ;
 wire \Tile_X1Y6_N1BEG[1] ;
 wire \Tile_X1Y6_N1BEG[2] ;
 wire \Tile_X1Y6_N1BEG[3] ;
 wire \Tile_X1Y6_N2BEG[0] ;
 wire \Tile_X1Y6_N2BEG[1] ;
 wire \Tile_X1Y6_N2BEG[2] ;
 wire \Tile_X1Y6_N2BEG[3] ;
 wire \Tile_X1Y6_N2BEG[4] ;
 wire \Tile_X1Y6_N2BEG[5] ;
 wire \Tile_X1Y6_N2BEG[6] ;
 wire \Tile_X1Y6_N2BEG[7] ;
 wire \Tile_X1Y6_N2BEGb[0] ;
 wire \Tile_X1Y6_N2BEGb[1] ;
 wire \Tile_X1Y6_N2BEGb[2] ;
 wire \Tile_X1Y6_N2BEGb[3] ;
 wire \Tile_X1Y6_N2BEGb[4] ;
 wire \Tile_X1Y6_N2BEGb[5] ;
 wire \Tile_X1Y6_N2BEGb[6] ;
 wire \Tile_X1Y6_N2BEGb[7] ;
 wire \Tile_X1Y6_N4BEG[0] ;
 wire \Tile_X1Y6_N4BEG[10] ;
 wire \Tile_X1Y6_N4BEG[11] ;
 wire \Tile_X1Y6_N4BEG[12] ;
 wire \Tile_X1Y6_N4BEG[13] ;
 wire \Tile_X1Y6_N4BEG[14] ;
 wire \Tile_X1Y6_N4BEG[15] ;
 wire \Tile_X1Y6_N4BEG[1] ;
 wire \Tile_X1Y6_N4BEG[2] ;
 wire \Tile_X1Y6_N4BEG[3] ;
 wire \Tile_X1Y6_N4BEG[4] ;
 wire \Tile_X1Y6_N4BEG[5] ;
 wire \Tile_X1Y6_N4BEG[6] ;
 wire \Tile_X1Y6_N4BEG[7] ;
 wire \Tile_X1Y6_N4BEG[8] ;
 wire \Tile_X1Y6_N4BEG[9] ;
 wire \Tile_X1Y6_NN4BEG[0] ;
 wire \Tile_X1Y6_NN4BEG[10] ;
 wire \Tile_X1Y6_NN4BEG[11] ;
 wire \Tile_X1Y6_NN4BEG[12] ;
 wire \Tile_X1Y6_NN4BEG[13] ;
 wire \Tile_X1Y6_NN4BEG[14] ;
 wire \Tile_X1Y6_NN4BEG[15] ;
 wire \Tile_X1Y6_NN4BEG[1] ;
 wire \Tile_X1Y6_NN4BEG[2] ;
 wire \Tile_X1Y6_NN4BEG[3] ;
 wire \Tile_X1Y6_NN4BEG[4] ;
 wire \Tile_X1Y6_NN4BEG[5] ;
 wire \Tile_X1Y6_NN4BEG[6] ;
 wire \Tile_X1Y6_NN4BEG[7] ;
 wire \Tile_X1Y6_NN4BEG[8] ;
 wire \Tile_X1Y6_NN4BEG[9] ;
 wire \Tile_X1Y6_S1BEG[0] ;
 wire \Tile_X1Y6_S1BEG[1] ;
 wire \Tile_X1Y6_S1BEG[2] ;
 wire \Tile_X1Y6_S1BEG[3] ;
 wire \Tile_X1Y6_S2BEG[0] ;
 wire \Tile_X1Y6_S2BEG[1] ;
 wire \Tile_X1Y6_S2BEG[2] ;
 wire \Tile_X1Y6_S2BEG[3] ;
 wire \Tile_X1Y6_S2BEG[4] ;
 wire \Tile_X1Y6_S2BEG[5] ;
 wire \Tile_X1Y6_S2BEG[6] ;
 wire \Tile_X1Y6_S2BEG[7] ;
 wire \Tile_X1Y6_S2BEGb[0] ;
 wire \Tile_X1Y6_S2BEGb[1] ;
 wire \Tile_X1Y6_S2BEGb[2] ;
 wire \Tile_X1Y6_S2BEGb[3] ;
 wire \Tile_X1Y6_S2BEGb[4] ;
 wire \Tile_X1Y6_S2BEGb[5] ;
 wire \Tile_X1Y6_S2BEGb[6] ;
 wire \Tile_X1Y6_S2BEGb[7] ;
 wire \Tile_X1Y6_S4BEG[0] ;
 wire \Tile_X1Y6_S4BEG[10] ;
 wire \Tile_X1Y6_S4BEG[11] ;
 wire \Tile_X1Y6_S4BEG[12] ;
 wire \Tile_X1Y6_S4BEG[13] ;
 wire \Tile_X1Y6_S4BEG[14] ;
 wire \Tile_X1Y6_S4BEG[15] ;
 wire \Tile_X1Y6_S4BEG[1] ;
 wire \Tile_X1Y6_S4BEG[2] ;
 wire \Tile_X1Y6_S4BEG[3] ;
 wire \Tile_X1Y6_S4BEG[4] ;
 wire \Tile_X1Y6_S4BEG[5] ;
 wire \Tile_X1Y6_S4BEG[6] ;
 wire \Tile_X1Y6_S4BEG[7] ;
 wire \Tile_X1Y6_S4BEG[8] ;
 wire \Tile_X1Y6_S4BEG[9] ;
 wire \Tile_X1Y6_SS4BEG[0] ;
 wire \Tile_X1Y6_SS4BEG[10] ;
 wire \Tile_X1Y6_SS4BEG[11] ;
 wire \Tile_X1Y6_SS4BEG[12] ;
 wire \Tile_X1Y6_SS4BEG[13] ;
 wire \Tile_X1Y6_SS4BEG[14] ;
 wire \Tile_X1Y6_SS4BEG[15] ;
 wire \Tile_X1Y6_SS4BEG[1] ;
 wire \Tile_X1Y6_SS4BEG[2] ;
 wire \Tile_X1Y6_SS4BEG[3] ;
 wire \Tile_X1Y6_SS4BEG[4] ;
 wire \Tile_X1Y6_SS4BEG[5] ;
 wire \Tile_X1Y6_SS4BEG[6] ;
 wire \Tile_X1Y6_SS4BEG[7] ;
 wire \Tile_X1Y6_SS4BEG[8] ;
 wire \Tile_X1Y6_SS4BEG[9] ;
 wire Tile_X1Y6_UserCLKo;
 wire \Tile_X1Y6_W1BEG[0] ;
 wire \Tile_X1Y6_W1BEG[1] ;
 wire \Tile_X1Y6_W1BEG[2] ;
 wire \Tile_X1Y6_W1BEG[3] ;
 wire \Tile_X1Y6_W2BEG[0] ;
 wire \Tile_X1Y6_W2BEG[1] ;
 wire \Tile_X1Y6_W2BEG[2] ;
 wire \Tile_X1Y6_W2BEG[3] ;
 wire \Tile_X1Y6_W2BEG[4] ;
 wire \Tile_X1Y6_W2BEG[5] ;
 wire \Tile_X1Y6_W2BEG[6] ;
 wire \Tile_X1Y6_W2BEG[7] ;
 wire \Tile_X1Y6_W2BEGb[0] ;
 wire \Tile_X1Y6_W2BEGb[1] ;
 wire \Tile_X1Y6_W2BEGb[2] ;
 wire \Tile_X1Y6_W2BEGb[3] ;
 wire \Tile_X1Y6_W2BEGb[4] ;
 wire \Tile_X1Y6_W2BEGb[5] ;
 wire \Tile_X1Y6_W2BEGb[6] ;
 wire \Tile_X1Y6_W2BEGb[7] ;
 wire \Tile_X1Y6_W6BEG[0] ;
 wire \Tile_X1Y6_W6BEG[10] ;
 wire \Tile_X1Y6_W6BEG[11] ;
 wire \Tile_X1Y6_W6BEG[1] ;
 wire \Tile_X1Y6_W6BEG[2] ;
 wire \Tile_X1Y6_W6BEG[3] ;
 wire \Tile_X1Y6_W6BEG[4] ;
 wire \Tile_X1Y6_W6BEG[5] ;
 wire \Tile_X1Y6_W6BEG[6] ;
 wire \Tile_X1Y6_W6BEG[7] ;
 wire \Tile_X1Y6_W6BEG[8] ;
 wire \Tile_X1Y6_W6BEG[9] ;
 wire \Tile_X1Y6_WW4BEG[0] ;
 wire \Tile_X1Y6_WW4BEG[10] ;
 wire \Tile_X1Y6_WW4BEG[11] ;
 wire \Tile_X1Y6_WW4BEG[12] ;
 wire \Tile_X1Y6_WW4BEG[13] ;
 wire \Tile_X1Y6_WW4BEG[14] ;
 wire \Tile_X1Y6_WW4BEG[15] ;
 wire \Tile_X1Y6_WW4BEG[1] ;
 wire \Tile_X1Y6_WW4BEG[2] ;
 wire \Tile_X1Y6_WW4BEG[3] ;
 wire \Tile_X1Y6_WW4BEG[4] ;
 wire \Tile_X1Y6_WW4BEG[5] ;
 wire \Tile_X1Y6_WW4BEG[6] ;
 wire \Tile_X1Y6_WW4BEG[7] ;
 wire \Tile_X1Y6_WW4BEG[8] ;
 wire \Tile_X1Y6_WW4BEG[9] ;
 wire Tile_X1Y7_Co;
 wire \Tile_X1Y7_E1BEG[0] ;
 wire \Tile_X1Y7_E1BEG[1] ;
 wire \Tile_X1Y7_E1BEG[2] ;
 wire \Tile_X1Y7_E1BEG[3] ;
 wire \Tile_X1Y7_E2BEG[0] ;
 wire \Tile_X1Y7_E2BEG[1] ;
 wire \Tile_X1Y7_E2BEG[2] ;
 wire \Tile_X1Y7_E2BEG[3] ;
 wire \Tile_X1Y7_E2BEG[4] ;
 wire \Tile_X1Y7_E2BEG[5] ;
 wire \Tile_X1Y7_E2BEG[6] ;
 wire \Tile_X1Y7_E2BEG[7] ;
 wire \Tile_X1Y7_E2BEGb[0] ;
 wire \Tile_X1Y7_E2BEGb[1] ;
 wire \Tile_X1Y7_E2BEGb[2] ;
 wire \Tile_X1Y7_E2BEGb[3] ;
 wire \Tile_X1Y7_E2BEGb[4] ;
 wire \Tile_X1Y7_E2BEGb[5] ;
 wire \Tile_X1Y7_E2BEGb[6] ;
 wire \Tile_X1Y7_E2BEGb[7] ;
 wire \Tile_X1Y7_E6BEG[0] ;
 wire \Tile_X1Y7_E6BEG[10] ;
 wire \Tile_X1Y7_E6BEG[11] ;
 wire \Tile_X1Y7_E6BEG[1] ;
 wire \Tile_X1Y7_E6BEG[2] ;
 wire \Tile_X1Y7_E6BEG[3] ;
 wire \Tile_X1Y7_E6BEG[4] ;
 wire \Tile_X1Y7_E6BEG[5] ;
 wire \Tile_X1Y7_E6BEG[6] ;
 wire \Tile_X1Y7_E6BEG[7] ;
 wire \Tile_X1Y7_E6BEG[8] ;
 wire \Tile_X1Y7_E6BEG[9] ;
 wire \Tile_X1Y7_EE4BEG[0] ;
 wire \Tile_X1Y7_EE4BEG[10] ;
 wire \Tile_X1Y7_EE4BEG[11] ;
 wire \Tile_X1Y7_EE4BEG[12] ;
 wire \Tile_X1Y7_EE4BEG[13] ;
 wire \Tile_X1Y7_EE4BEG[14] ;
 wire \Tile_X1Y7_EE4BEG[15] ;
 wire \Tile_X1Y7_EE4BEG[1] ;
 wire \Tile_X1Y7_EE4BEG[2] ;
 wire \Tile_X1Y7_EE4BEG[3] ;
 wire \Tile_X1Y7_EE4BEG[4] ;
 wire \Tile_X1Y7_EE4BEG[5] ;
 wire \Tile_X1Y7_EE4BEG[6] ;
 wire \Tile_X1Y7_EE4BEG[7] ;
 wire \Tile_X1Y7_EE4BEG[8] ;
 wire \Tile_X1Y7_EE4BEG[9] ;
 wire \Tile_X1Y7_FrameData_O[0] ;
 wire \Tile_X1Y7_FrameData_O[10] ;
 wire \Tile_X1Y7_FrameData_O[11] ;
 wire \Tile_X1Y7_FrameData_O[12] ;
 wire \Tile_X1Y7_FrameData_O[13] ;
 wire \Tile_X1Y7_FrameData_O[14] ;
 wire \Tile_X1Y7_FrameData_O[15] ;
 wire \Tile_X1Y7_FrameData_O[16] ;
 wire \Tile_X1Y7_FrameData_O[17] ;
 wire \Tile_X1Y7_FrameData_O[18] ;
 wire \Tile_X1Y7_FrameData_O[19] ;
 wire \Tile_X1Y7_FrameData_O[1] ;
 wire \Tile_X1Y7_FrameData_O[20] ;
 wire \Tile_X1Y7_FrameData_O[21] ;
 wire \Tile_X1Y7_FrameData_O[22] ;
 wire \Tile_X1Y7_FrameData_O[23] ;
 wire \Tile_X1Y7_FrameData_O[24] ;
 wire \Tile_X1Y7_FrameData_O[25] ;
 wire \Tile_X1Y7_FrameData_O[26] ;
 wire \Tile_X1Y7_FrameData_O[27] ;
 wire \Tile_X1Y7_FrameData_O[28] ;
 wire \Tile_X1Y7_FrameData_O[29] ;
 wire \Tile_X1Y7_FrameData_O[2] ;
 wire \Tile_X1Y7_FrameData_O[30] ;
 wire \Tile_X1Y7_FrameData_O[31] ;
 wire \Tile_X1Y7_FrameData_O[3] ;
 wire \Tile_X1Y7_FrameData_O[4] ;
 wire \Tile_X1Y7_FrameData_O[5] ;
 wire \Tile_X1Y7_FrameData_O[6] ;
 wire \Tile_X1Y7_FrameData_O[7] ;
 wire \Tile_X1Y7_FrameData_O[8] ;
 wire \Tile_X1Y7_FrameData_O[9] ;
 wire \Tile_X1Y7_FrameStrobe_O[0] ;
 wire \Tile_X1Y7_FrameStrobe_O[10] ;
 wire \Tile_X1Y7_FrameStrobe_O[11] ;
 wire \Tile_X1Y7_FrameStrobe_O[12] ;
 wire \Tile_X1Y7_FrameStrobe_O[13] ;
 wire \Tile_X1Y7_FrameStrobe_O[14] ;
 wire \Tile_X1Y7_FrameStrobe_O[15] ;
 wire \Tile_X1Y7_FrameStrobe_O[16] ;
 wire \Tile_X1Y7_FrameStrobe_O[17] ;
 wire \Tile_X1Y7_FrameStrobe_O[18] ;
 wire \Tile_X1Y7_FrameStrobe_O[19] ;
 wire \Tile_X1Y7_FrameStrobe_O[1] ;
 wire \Tile_X1Y7_FrameStrobe_O[2] ;
 wire \Tile_X1Y7_FrameStrobe_O[3] ;
 wire \Tile_X1Y7_FrameStrobe_O[4] ;
 wire \Tile_X1Y7_FrameStrobe_O[5] ;
 wire \Tile_X1Y7_FrameStrobe_O[6] ;
 wire \Tile_X1Y7_FrameStrobe_O[7] ;
 wire \Tile_X1Y7_FrameStrobe_O[8] ;
 wire \Tile_X1Y7_FrameStrobe_O[9] ;
 wire \Tile_X1Y7_N1BEG[0] ;
 wire \Tile_X1Y7_N1BEG[1] ;
 wire \Tile_X1Y7_N1BEG[2] ;
 wire \Tile_X1Y7_N1BEG[3] ;
 wire \Tile_X1Y7_N2BEG[0] ;
 wire \Tile_X1Y7_N2BEG[1] ;
 wire \Tile_X1Y7_N2BEG[2] ;
 wire \Tile_X1Y7_N2BEG[3] ;
 wire \Tile_X1Y7_N2BEG[4] ;
 wire \Tile_X1Y7_N2BEG[5] ;
 wire \Tile_X1Y7_N2BEG[6] ;
 wire \Tile_X1Y7_N2BEG[7] ;
 wire \Tile_X1Y7_N2BEGb[0] ;
 wire \Tile_X1Y7_N2BEGb[1] ;
 wire \Tile_X1Y7_N2BEGb[2] ;
 wire \Tile_X1Y7_N2BEGb[3] ;
 wire \Tile_X1Y7_N2BEGb[4] ;
 wire \Tile_X1Y7_N2BEGb[5] ;
 wire \Tile_X1Y7_N2BEGb[6] ;
 wire \Tile_X1Y7_N2BEGb[7] ;
 wire \Tile_X1Y7_N4BEG[0] ;
 wire \Tile_X1Y7_N4BEG[10] ;
 wire \Tile_X1Y7_N4BEG[11] ;
 wire \Tile_X1Y7_N4BEG[12] ;
 wire \Tile_X1Y7_N4BEG[13] ;
 wire \Tile_X1Y7_N4BEG[14] ;
 wire \Tile_X1Y7_N4BEG[15] ;
 wire \Tile_X1Y7_N4BEG[1] ;
 wire \Tile_X1Y7_N4BEG[2] ;
 wire \Tile_X1Y7_N4BEG[3] ;
 wire \Tile_X1Y7_N4BEG[4] ;
 wire \Tile_X1Y7_N4BEG[5] ;
 wire \Tile_X1Y7_N4BEG[6] ;
 wire \Tile_X1Y7_N4BEG[7] ;
 wire \Tile_X1Y7_N4BEG[8] ;
 wire \Tile_X1Y7_N4BEG[9] ;
 wire \Tile_X1Y7_NN4BEG[0] ;
 wire \Tile_X1Y7_NN4BEG[10] ;
 wire \Tile_X1Y7_NN4BEG[11] ;
 wire \Tile_X1Y7_NN4BEG[12] ;
 wire \Tile_X1Y7_NN4BEG[13] ;
 wire \Tile_X1Y7_NN4BEG[14] ;
 wire \Tile_X1Y7_NN4BEG[15] ;
 wire \Tile_X1Y7_NN4BEG[1] ;
 wire \Tile_X1Y7_NN4BEG[2] ;
 wire \Tile_X1Y7_NN4BEG[3] ;
 wire \Tile_X1Y7_NN4BEG[4] ;
 wire \Tile_X1Y7_NN4BEG[5] ;
 wire \Tile_X1Y7_NN4BEG[6] ;
 wire \Tile_X1Y7_NN4BEG[7] ;
 wire \Tile_X1Y7_NN4BEG[8] ;
 wire \Tile_X1Y7_NN4BEG[9] ;
 wire \Tile_X1Y7_S1BEG[0] ;
 wire \Tile_X1Y7_S1BEG[1] ;
 wire \Tile_X1Y7_S1BEG[2] ;
 wire \Tile_X1Y7_S1BEG[3] ;
 wire \Tile_X1Y7_S2BEG[0] ;
 wire \Tile_X1Y7_S2BEG[1] ;
 wire \Tile_X1Y7_S2BEG[2] ;
 wire \Tile_X1Y7_S2BEG[3] ;
 wire \Tile_X1Y7_S2BEG[4] ;
 wire \Tile_X1Y7_S2BEG[5] ;
 wire \Tile_X1Y7_S2BEG[6] ;
 wire \Tile_X1Y7_S2BEG[7] ;
 wire \Tile_X1Y7_S2BEGb[0] ;
 wire \Tile_X1Y7_S2BEGb[1] ;
 wire \Tile_X1Y7_S2BEGb[2] ;
 wire \Tile_X1Y7_S2BEGb[3] ;
 wire \Tile_X1Y7_S2BEGb[4] ;
 wire \Tile_X1Y7_S2BEGb[5] ;
 wire \Tile_X1Y7_S2BEGb[6] ;
 wire \Tile_X1Y7_S2BEGb[7] ;
 wire \Tile_X1Y7_S4BEG[0] ;
 wire \Tile_X1Y7_S4BEG[10] ;
 wire \Tile_X1Y7_S4BEG[11] ;
 wire \Tile_X1Y7_S4BEG[12] ;
 wire \Tile_X1Y7_S4BEG[13] ;
 wire \Tile_X1Y7_S4BEG[14] ;
 wire \Tile_X1Y7_S4BEG[15] ;
 wire \Tile_X1Y7_S4BEG[1] ;
 wire \Tile_X1Y7_S4BEG[2] ;
 wire \Tile_X1Y7_S4BEG[3] ;
 wire \Tile_X1Y7_S4BEG[4] ;
 wire \Tile_X1Y7_S4BEG[5] ;
 wire \Tile_X1Y7_S4BEG[6] ;
 wire \Tile_X1Y7_S4BEG[7] ;
 wire \Tile_X1Y7_S4BEG[8] ;
 wire \Tile_X1Y7_S4BEG[9] ;
 wire \Tile_X1Y7_SS4BEG[0] ;
 wire \Tile_X1Y7_SS4BEG[10] ;
 wire \Tile_X1Y7_SS4BEG[11] ;
 wire \Tile_X1Y7_SS4BEG[12] ;
 wire \Tile_X1Y7_SS4BEG[13] ;
 wire \Tile_X1Y7_SS4BEG[14] ;
 wire \Tile_X1Y7_SS4BEG[15] ;
 wire \Tile_X1Y7_SS4BEG[1] ;
 wire \Tile_X1Y7_SS4BEG[2] ;
 wire \Tile_X1Y7_SS4BEG[3] ;
 wire \Tile_X1Y7_SS4BEG[4] ;
 wire \Tile_X1Y7_SS4BEG[5] ;
 wire \Tile_X1Y7_SS4BEG[6] ;
 wire \Tile_X1Y7_SS4BEG[7] ;
 wire \Tile_X1Y7_SS4BEG[8] ;
 wire \Tile_X1Y7_SS4BEG[9] ;
 wire Tile_X1Y7_UserCLKo;
 wire \Tile_X1Y7_W1BEG[0] ;
 wire \Tile_X1Y7_W1BEG[1] ;
 wire \Tile_X1Y7_W1BEG[2] ;
 wire \Tile_X1Y7_W1BEG[3] ;
 wire \Tile_X1Y7_W2BEG[0] ;
 wire \Tile_X1Y7_W2BEG[1] ;
 wire \Tile_X1Y7_W2BEG[2] ;
 wire \Tile_X1Y7_W2BEG[3] ;
 wire \Tile_X1Y7_W2BEG[4] ;
 wire \Tile_X1Y7_W2BEG[5] ;
 wire \Tile_X1Y7_W2BEG[6] ;
 wire \Tile_X1Y7_W2BEG[7] ;
 wire \Tile_X1Y7_W2BEGb[0] ;
 wire \Tile_X1Y7_W2BEGb[1] ;
 wire \Tile_X1Y7_W2BEGb[2] ;
 wire \Tile_X1Y7_W2BEGb[3] ;
 wire \Tile_X1Y7_W2BEGb[4] ;
 wire \Tile_X1Y7_W2BEGb[5] ;
 wire \Tile_X1Y7_W2BEGb[6] ;
 wire \Tile_X1Y7_W2BEGb[7] ;
 wire \Tile_X1Y7_W6BEG[0] ;
 wire \Tile_X1Y7_W6BEG[10] ;
 wire \Tile_X1Y7_W6BEG[11] ;
 wire \Tile_X1Y7_W6BEG[1] ;
 wire \Tile_X1Y7_W6BEG[2] ;
 wire \Tile_X1Y7_W6BEG[3] ;
 wire \Tile_X1Y7_W6BEG[4] ;
 wire \Tile_X1Y7_W6BEG[5] ;
 wire \Tile_X1Y7_W6BEG[6] ;
 wire \Tile_X1Y7_W6BEG[7] ;
 wire \Tile_X1Y7_W6BEG[8] ;
 wire \Tile_X1Y7_W6BEG[9] ;
 wire \Tile_X1Y7_WW4BEG[0] ;
 wire \Tile_X1Y7_WW4BEG[10] ;
 wire \Tile_X1Y7_WW4BEG[11] ;
 wire \Tile_X1Y7_WW4BEG[12] ;
 wire \Tile_X1Y7_WW4BEG[13] ;
 wire \Tile_X1Y7_WW4BEG[14] ;
 wire \Tile_X1Y7_WW4BEG[15] ;
 wire \Tile_X1Y7_WW4BEG[1] ;
 wire \Tile_X1Y7_WW4BEG[2] ;
 wire \Tile_X1Y7_WW4BEG[3] ;
 wire \Tile_X1Y7_WW4BEG[4] ;
 wire \Tile_X1Y7_WW4BEG[5] ;
 wire \Tile_X1Y7_WW4BEG[6] ;
 wire \Tile_X1Y7_WW4BEG[7] ;
 wire \Tile_X1Y7_WW4BEG[8] ;
 wire \Tile_X1Y7_WW4BEG[9] ;
 wire Tile_X1Y8_Co;
 wire \Tile_X1Y8_E1BEG[0] ;
 wire \Tile_X1Y8_E1BEG[1] ;
 wire \Tile_X1Y8_E1BEG[2] ;
 wire \Tile_X1Y8_E1BEG[3] ;
 wire \Tile_X1Y8_E2BEG[0] ;
 wire \Tile_X1Y8_E2BEG[1] ;
 wire \Tile_X1Y8_E2BEG[2] ;
 wire \Tile_X1Y8_E2BEG[3] ;
 wire \Tile_X1Y8_E2BEG[4] ;
 wire \Tile_X1Y8_E2BEG[5] ;
 wire \Tile_X1Y8_E2BEG[6] ;
 wire \Tile_X1Y8_E2BEG[7] ;
 wire \Tile_X1Y8_E2BEGb[0] ;
 wire \Tile_X1Y8_E2BEGb[1] ;
 wire \Tile_X1Y8_E2BEGb[2] ;
 wire \Tile_X1Y8_E2BEGb[3] ;
 wire \Tile_X1Y8_E2BEGb[4] ;
 wire \Tile_X1Y8_E2BEGb[5] ;
 wire \Tile_X1Y8_E2BEGb[6] ;
 wire \Tile_X1Y8_E2BEGb[7] ;
 wire \Tile_X1Y8_E6BEG[0] ;
 wire \Tile_X1Y8_E6BEG[10] ;
 wire \Tile_X1Y8_E6BEG[11] ;
 wire \Tile_X1Y8_E6BEG[1] ;
 wire \Tile_X1Y8_E6BEG[2] ;
 wire \Tile_X1Y8_E6BEG[3] ;
 wire \Tile_X1Y8_E6BEG[4] ;
 wire \Tile_X1Y8_E6BEG[5] ;
 wire \Tile_X1Y8_E6BEG[6] ;
 wire \Tile_X1Y8_E6BEG[7] ;
 wire \Tile_X1Y8_E6BEG[8] ;
 wire \Tile_X1Y8_E6BEG[9] ;
 wire \Tile_X1Y8_EE4BEG[0] ;
 wire \Tile_X1Y8_EE4BEG[10] ;
 wire \Tile_X1Y8_EE4BEG[11] ;
 wire \Tile_X1Y8_EE4BEG[12] ;
 wire \Tile_X1Y8_EE4BEG[13] ;
 wire \Tile_X1Y8_EE4BEG[14] ;
 wire \Tile_X1Y8_EE4BEG[15] ;
 wire \Tile_X1Y8_EE4BEG[1] ;
 wire \Tile_X1Y8_EE4BEG[2] ;
 wire \Tile_X1Y8_EE4BEG[3] ;
 wire \Tile_X1Y8_EE4BEG[4] ;
 wire \Tile_X1Y8_EE4BEG[5] ;
 wire \Tile_X1Y8_EE4BEG[6] ;
 wire \Tile_X1Y8_EE4BEG[7] ;
 wire \Tile_X1Y8_EE4BEG[8] ;
 wire \Tile_X1Y8_EE4BEG[9] ;
 wire \Tile_X1Y8_FrameData_O[0] ;
 wire \Tile_X1Y8_FrameData_O[10] ;
 wire \Tile_X1Y8_FrameData_O[11] ;
 wire \Tile_X1Y8_FrameData_O[12] ;
 wire \Tile_X1Y8_FrameData_O[13] ;
 wire \Tile_X1Y8_FrameData_O[14] ;
 wire \Tile_X1Y8_FrameData_O[15] ;
 wire \Tile_X1Y8_FrameData_O[16] ;
 wire \Tile_X1Y8_FrameData_O[17] ;
 wire \Tile_X1Y8_FrameData_O[18] ;
 wire \Tile_X1Y8_FrameData_O[19] ;
 wire \Tile_X1Y8_FrameData_O[1] ;
 wire \Tile_X1Y8_FrameData_O[20] ;
 wire \Tile_X1Y8_FrameData_O[21] ;
 wire \Tile_X1Y8_FrameData_O[22] ;
 wire \Tile_X1Y8_FrameData_O[23] ;
 wire \Tile_X1Y8_FrameData_O[24] ;
 wire \Tile_X1Y8_FrameData_O[25] ;
 wire \Tile_X1Y8_FrameData_O[26] ;
 wire \Tile_X1Y8_FrameData_O[27] ;
 wire \Tile_X1Y8_FrameData_O[28] ;
 wire \Tile_X1Y8_FrameData_O[29] ;
 wire \Tile_X1Y8_FrameData_O[2] ;
 wire \Tile_X1Y8_FrameData_O[30] ;
 wire \Tile_X1Y8_FrameData_O[31] ;
 wire \Tile_X1Y8_FrameData_O[3] ;
 wire \Tile_X1Y8_FrameData_O[4] ;
 wire \Tile_X1Y8_FrameData_O[5] ;
 wire \Tile_X1Y8_FrameData_O[6] ;
 wire \Tile_X1Y8_FrameData_O[7] ;
 wire \Tile_X1Y8_FrameData_O[8] ;
 wire \Tile_X1Y8_FrameData_O[9] ;
 wire \Tile_X1Y8_FrameStrobe_O[0] ;
 wire \Tile_X1Y8_FrameStrobe_O[10] ;
 wire \Tile_X1Y8_FrameStrobe_O[11] ;
 wire \Tile_X1Y8_FrameStrobe_O[12] ;
 wire \Tile_X1Y8_FrameStrobe_O[13] ;
 wire \Tile_X1Y8_FrameStrobe_O[14] ;
 wire \Tile_X1Y8_FrameStrobe_O[15] ;
 wire \Tile_X1Y8_FrameStrobe_O[16] ;
 wire \Tile_X1Y8_FrameStrobe_O[17] ;
 wire \Tile_X1Y8_FrameStrobe_O[18] ;
 wire \Tile_X1Y8_FrameStrobe_O[19] ;
 wire \Tile_X1Y8_FrameStrobe_O[1] ;
 wire \Tile_X1Y8_FrameStrobe_O[2] ;
 wire \Tile_X1Y8_FrameStrobe_O[3] ;
 wire \Tile_X1Y8_FrameStrobe_O[4] ;
 wire \Tile_X1Y8_FrameStrobe_O[5] ;
 wire \Tile_X1Y8_FrameStrobe_O[6] ;
 wire \Tile_X1Y8_FrameStrobe_O[7] ;
 wire \Tile_X1Y8_FrameStrobe_O[8] ;
 wire \Tile_X1Y8_FrameStrobe_O[9] ;
 wire \Tile_X1Y8_N1BEG[0] ;
 wire \Tile_X1Y8_N1BEG[1] ;
 wire \Tile_X1Y8_N1BEG[2] ;
 wire \Tile_X1Y8_N1BEG[3] ;
 wire \Tile_X1Y8_N2BEG[0] ;
 wire \Tile_X1Y8_N2BEG[1] ;
 wire \Tile_X1Y8_N2BEG[2] ;
 wire \Tile_X1Y8_N2BEG[3] ;
 wire \Tile_X1Y8_N2BEG[4] ;
 wire \Tile_X1Y8_N2BEG[5] ;
 wire \Tile_X1Y8_N2BEG[6] ;
 wire \Tile_X1Y8_N2BEG[7] ;
 wire \Tile_X1Y8_N2BEGb[0] ;
 wire \Tile_X1Y8_N2BEGb[1] ;
 wire \Tile_X1Y8_N2BEGb[2] ;
 wire \Tile_X1Y8_N2BEGb[3] ;
 wire \Tile_X1Y8_N2BEGb[4] ;
 wire \Tile_X1Y8_N2BEGb[5] ;
 wire \Tile_X1Y8_N2BEGb[6] ;
 wire \Tile_X1Y8_N2BEGb[7] ;
 wire \Tile_X1Y8_N4BEG[0] ;
 wire \Tile_X1Y8_N4BEG[10] ;
 wire \Tile_X1Y8_N4BEG[11] ;
 wire \Tile_X1Y8_N4BEG[12] ;
 wire \Tile_X1Y8_N4BEG[13] ;
 wire \Tile_X1Y8_N4BEG[14] ;
 wire \Tile_X1Y8_N4BEG[15] ;
 wire \Tile_X1Y8_N4BEG[1] ;
 wire \Tile_X1Y8_N4BEG[2] ;
 wire \Tile_X1Y8_N4BEG[3] ;
 wire \Tile_X1Y8_N4BEG[4] ;
 wire \Tile_X1Y8_N4BEG[5] ;
 wire \Tile_X1Y8_N4BEG[6] ;
 wire \Tile_X1Y8_N4BEG[7] ;
 wire \Tile_X1Y8_N4BEG[8] ;
 wire \Tile_X1Y8_N4BEG[9] ;
 wire \Tile_X1Y8_NN4BEG[0] ;
 wire \Tile_X1Y8_NN4BEG[10] ;
 wire \Tile_X1Y8_NN4BEG[11] ;
 wire \Tile_X1Y8_NN4BEG[12] ;
 wire \Tile_X1Y8_NN4BEG[13] ;
 wire \Tile_X1Y8_NN4BEG[14] ;
 wire \Tile_X1Y8_NN4BEG[15] ;
 wire \Tile_X1Y8_NN4BEG[1] ;
 wire \Tile_X1Y8_NN4BEG[2] ;
 wire \Tile_X1Y8_NN4BEG[3] ;
 wire \Tile_X1Y8_NN4BEG[4] ;
 wire \Tile_X1Y8_NN4BEG[5] ;
 wire \Tile_X1Y8_NN4BEG[6] ;
 wire \Tile_X1Y8_NN4BEG[7] ;
 wire \Tile_X1Y8_NN4BEG[8] ;
 wire \Tile_X1Y8_NN4BEG[9] ;
 wire \Tile_X1Y8_S1BEG[0] ;
 wire \Tile_X1Y8_S1BEG[1] ;
 wire \Tile_X1Y8_S1BEG[2] ;
 wire \Tile_X1Y8_S1BEG[3] ;
 wire \Tile_X1Y8_S2BEG[0] ;
 wire \Tile_X1Y8_S2BEG[1] ;
 wire \Tile_X1Y8_S2BEG[2] ;
 wire \Tile_X1Y8_S2BEG[3] ;
 wire \Tile_X1Y8_S2BEG[4] ;
 wire \Tile_X1Y8_S2BEG[5] ;
 wire \Tile_X1Y8_S2BEG[6] ;
 wire \Tile_X1Y8_S2BEG[7] ;
 wire \Tile_X1Y8_S2BEGb[0] ;
 wire \Tile_X1Y8_S2BEGb[1] ;
 wire \Tile_X1Y8_S2BEGb[2] ;
 wire \Tile_X1Y8_S2BEGb[3] ;
 wire \Tile_X1Y8_S2BEGb[4] ;
 wire \Tile_X1Y8_S2BEGb[5] ;
 wire \Tile_X1Y8_S2BEGb[6] ;
 wire \Tile_X1Y8_S2BEGb[7] ;
 wire \Tile_X1Y8_S4BEG[0] ;
 wire \Tile_X1Y8_S4BEG[10] ;
 wire \Tile_X1Y8_S4BEG[11] ;
 wire \Tile_X1Y8_S4BEG[12] ;
 wire \Tile_X1Y8_S4BEG[13] ;
 wire \Tile_X1Y8_S4BEG[14] ;
 wire \Tile_X1Y8_S4BEG[15] ;
 wire \Tile_X1Y8_S4BEG[1] ;
 wire \Tile_X1Y8_S4BEG[2] ;
 wire \Tile_X1Y8_S4BEG[3] ;
 wire \Tile_X1Y8_S4BEG[4] ;
 wire \Tile_X1Y8_S4BEG[5] ;
 wire \Tile_X1Y8_S4BEG[6] ;
 wire \Tile_X1Y8_S4BEG[7] ;
 wire \Tile_X1Y8_S4BEG[8] ;
 wire \Tile_X1Y8_S4BEG[9] ;
 wire \Tile_X1Y8_SS4BEG[0] ;
 wire \Tile_X1Y8_SS4BEG[10] ;
 wire \Tile_X1Y8_SS4BEG[11] ;
 wire \Tile_X1Y8_SS4BEG[12] ;
 wire \Tile_X1Y8_SS4BEG[13] ;
 wire \Tile_X1Y8_SS4BEG[14] ;
 wire \Tile_X1Y8_SS4BEG[15] ;
 wire \Tile_X1Y8_SS4BEG[1] ;
 wire \Tile_X1Y8_SS4BEG[2] ;
 wire \Tile_X1Y8_SS4BEG[3] ;
 wire \Tile_X1Y8_SS4BEG[4] ;
 wire \Tile_X1Y8_SS4BEG[5] ;
 wire \Tile_X1Y8_SS4BEG[6] ;
 wire \Tile_X1Y8_SS4BEG[7] ;
 wire \Tile_X1Y8_SS4BEG[8] ;
 wire \Tile_X1Y8_SS4BEG[9] ;
 wire Tile_X1Y8_UserCLKo;
 wire \Tile_X1Y8_W1BEG[0] ;
 wire \Tile_X1Y8_W1BEG[1] ;
 wire \Tile_X1Y8_W1BEG[2] ;
 wire \Tile_X1Y8_W1BEG[3] ;
 wire \Tile_X1Y8_W2BEG[0] ;
 wire \Tile_X1Y8_W2BEG[1] ;
 wire \Tile_X1Y8_W2BEG[2] ;
 wire \Tile_X1Y8_W2BEG[3] ;
 wire \Tile_X1Y8_W2BEG[4] ;
 wire \Tile_X1Y8_W2BEG[5] ;
 wire \Tile_X1Y8_W2BEG[6] ;
 wire \Tile_X1Y8_W2BEG[7] ;
 wire \Tile_X1Y8_W2BEGb[0] ;
 wire \Tile_X1Y8_W2BEGb[1] ;
 wire \Tile_X1Y8_W2BEGb[2] ;
 wire \Tile_X1Y8_W2BEGb[3] ;
 wire \Tile_X1Y8_W2BEGb[4] ;
 wire \Tile_X1Y8_W2BEGb[5] ;
 wire \Tile_X1Y8_W2BEGb[6] ;
 wire \Tile_X1Y8_W2BEGb[7] ;
 wire \Tile_X1Y8_W6BEG[0] ;
 wire \Tile_X1Y8_W6BEG[10] ;
 wire \Tile_X1Y8_W6BEG[11] ;
 wire \Tile_X1Y8_W6BEG[1] ;
 wire \Tile_X1Y8_W6BEG[2] ;
 wire \Tile_X1Y8_W6BEG[3] ;
 wire \Tile_X1Y8_W6BEG[4] ;
 wire \Tile_X1Y8_W6BEG[5] ;
 wire \Tile_X1Y8_W6BEG[6] ;
 wire \Tile_X1Y8_W6BEG[7] ;
 wire \Tile_X1Y8_W6BEG[8] ;
 wire \Tile_X1Y8_W6BEG[9] ;
 wire \Tile_X1Y8_WW4BEG[0] ;
 wire \Tile_X1Y8_WW4BEG[10] ;
 wire \Tile_X1Y8_WW4BEG[11] ;
 wire \Tile_X1Y8_WW4BEG[12] ;
 wire \Tile_X1Y8_WW4BEG[13] ;
 wire \Tile_X1Y8_WW4BEG[14] ;
 wire \Tile_X1Y8_WW4BEG[15] ;
 wire \Tile_X1Y8_WW4BEG[1] ;
 wire \Tile_X1Y8_WW4BEG[2] ;
 wire \Tile_X1Y8_WW4BEG[3] ;
 wire \Tile_X1Y8_WW4BEG[4] ;
 wire \Tile_X1Y8_WW4BEG[5] ;
 wire \Tile_X1Y8_WW4BEG[6] ;
 wire \Tile_X1Y8_WW4BEG[7] ;
 wire \Tile_X1Y8_WW4BEG[8] ;
 wire \Tile_X1Y8_WW4BEG[9] ;
 wire Tile_X1Y9_Co;
 wire \Tile_X1Y9_E1BEG[0] ;
 wire \Tile_X1Y9_E1BEG[1] ;
 wire \Tile_X1Y9_E1BEG[2] ;
 wire \Tile_X1Y9_E1BEG[3] ;
 wire \Tile_X1Y9_E2BEG[0] ;
 wire \Tile_X1Y9_E2BEG[1] ;
 wire \Tile_X1Y9_E2BEG[2] ;
 wire \Tile_X1Y9_E2BEG[3] ;
 wire \Tile_X1Y9_E2BEG[4] ;
 wire \Tile_X1Y9_E2BEG[5] ;
 wire \Tile_X1Y9_E2BEG[6] ;
 wire \Tile_X1Y9_E2BEG[7] ;
 wire \Tile_X1Y9_E2BEGb[0] ;
 wire \Tile_X1Y9_E2BEGb[1] ;
 wire \Tile_X1Y9_E2BEGb[2] ;
 wire \Tile_X1Y9_E2BEGb[3] ;
 wire \Tile_X1Y9_E2BEGb[4] ;
 wire \Tile_X1Y9_E2BEGb[5] ;
 wire \Tile_X1Y9_E2BEGb[6] ;
 wire \Tile_X1Y9_E2BEGb[7] ;
 wire \Tile_X1Y9_E6BEG[0] ;
 wire \Tile_X1Y9_E6BEG[10] ;
 wire \Tile_X1Y9_E6BEG[11] ;
 wire \Tile_X1Y9_E6BEG[1] ;
 wire \Tile_X1Y9_E6BEG[2] ;
 wire \Tile_X1Y9_E6BEG[3] ;
 wire \Tile_X1Y9_E6BEG[4] ;
 wire \Tile_X1Y9_E6BEG[5] ;
 wire \Tile_X1Y9_E6BEG[6] ;
 wire \Tile_X1Y9_E6BEG[7] ;
 wire \Tile_X1Y9_E6BEG[8] ;
 wire \Tile_X1Y9_E6BEG[9] ;
 wire \Tile_X1Y9_EE4BEG[0] ;
 wire \Tile_X1Y9_EE4BEG[10] ;
 wire \Tile_X1Y9_EE4BEG[11] ;
 wire \Tile_X1Y9_EE4BEG[12] ;
 wire \Tile_X1Y9_EE4BEG[13] ;
 wire \Tile_X1Y9_EE4BEG[14] ;
 wire \Tile_X1Y9_EE4BEG[15] ;
 wire \Tile_X1Y9_EE4BEG[1] ;
 wire \Tile_X1Y9_EE4BEG[2] ;
 wire \Tile_X1Y9_EE4BEG[3] ;
 wire \Tile_X1Y9_EE4BEG[4] ;
 wire \Tile_X1Y9_EE4BEG[5] ;
 wire \Tile_X1Y9_EE4BEG[6] ;
 wire \Tile_X1Y9_EE4BEG[7] ;
 wire \Tile_X1Y9_EE4BEG[8] ;
 wire \Tile_X1Y9_EE4BEG[9] ;
 wire \Tile_X1Y9_FrameData_O[0] ;
 wire \Tile_X1Y9_FrameData_O[10] ;
 wire \Tile_X1Y9_FrameData_O[11] ;
 wire \Tile_X1Y9_FrameData_O[12] ;
 wire \Tile_X1Y9_FrameData_O[13] ;
 wire \Tile_X1Y9_FrameData_O[14] ;
 wire \Tile_X1Y9_FrameData_O[15] ;
 wire \Tile_X1Y9_FrameData_O[16] ;
 wire \Tile_X1Y9_FrameData_O[17] ;
 wire \Tile_X1Y9_FrameData_O[18] ;
 wire \Tile_X1Y9_FrameData_O[19] ;
 wire \Tile_X1Y9_FrameData_O[1] ;
 wire \Tile_X1Y9_FrameData_O[20] ;
 wire \Tile_X1Y9_FrameData_O[21] ;
 wire \Tile_X1Y9_FrameData_O[22] ;
 wire \Tile_X1Y9_FrameData_O[23] ;
 wire \Tile_X1Y9_FrameData_O[24] ;
 wire \Tile_X1Y9_FrameData_O[25] ;
 wire \Tile_X1Y9_FrameData_O[26] ;
 wire \Tile_X1Y9_FrameData_O[27] ;
 wire \Tile_X1Y9_FrameData_O[28] ;
 wire \Tile_X1Y9_FrameData_O[29] ;
 wire \Tile_X1Y9_FrameData_O[2] ;
 wire \Tile_X1Y9_FrameData_O[30] ;
 wire \Tile_X1Y9_FrameData_O[31] ;
 wire \Tile_X1Y9_FrameData_O[3] ;
 wire \Tile_X1Y9_FrameData_O[4] ;
 wire \Tile_X1Y9_FrameData_O[5] ;
 wire \Tile_X1Y9_FrameData_O[6] ;
 wire \Tile_X1Y9_FrameData_O[7] ;
 wire \Tile_X1Y9_FrameData_O[8] ;
 wire \Tile_X1Y9_FrameData_O[9] ;
 wire \Tile_X1Y9_FrameStrobe_O[0] ;
 wire \Tile_X1Y9_FrameStrobe_O[10] ;
 wire \Tile_X1Y9_FrameStrobe_O[11] ;
 wire \Tile_X1Y9_FrameStrobe_O[12] ;
 wire \Tile_X1Y9_FrameStrobe_O[13] ;
 wire \Tile_X1Y9_FrameStrobe_O[14] ;
 wire \Tile_X1Y9_FrameStrobe_O[15] ;
 wire \Tile_X1Y9_FrameStrobe_O[16] ;
 wire \Tile_X1Y9_FrameStrobe_O[17] ;
 wire \Tile_X1Y9_FrameStrobe_O[18] ;
 wire \Tile_X1Y9_FrameStrobe_O[19] ;
 wire \Tile_X1Y9_FrameStrobe_O[1] ;
 wire \Tile_X1Y9_FrameStrobe_O[2] ;
 wire \Tile_X1Y9_FrameStrobe_O[3] ;
 wire \Tile_X1Y9_FrameStrobe_O[4] ;
 wire \Tile_X1Y9_FrameStrobe_O[5] ;
 wire \Tile_X1Y9_FrameStrobe_O[6] ;
 wire \Tile_X1Y9_FrameStrobe_O[7] ;
 wire \Tile_X1Y9_FrameStrobe_O[8] ;
 wire \Tile_X1Y9_FrameStrobe_O[9] ;
 wire \Tile_X1Y9_N1BEG[0] ;
 wire \Tile_X1Y9_N1BEG[1] ;
 wire \Tile_X1Y9_N1BEG[2] ;
 wire \Tile_X1Y9_N1BEG[3] ;
 wire \Tile_X1Y9_N2BEG[0] ;
 wire \Tile_X1Y9_N2BEG[1] ;
 wire \Tile_X1Y9_N2BEG[2] ;
 wire \Tile_X1Y9_N2BEG[3] ;
 wire \Tile_X1Y9_N2BEG[4] ;
 wire \Tile_X1Y9_N2BEG[5] ;
 wire \Tile_X1Y9_N2BEG[6] ;
 wire \Tile_X1Y9_N2BEG[7] ;
 wire \Tile_X1Y9_N2BEGb[0] ;
 wire \Tile_X1Y9_N2BEGb[1] ;
 wire \Tile_X1Y9_N2BEGb[2] ;
 wire \Tile_X1Y9_N2BEGb[3] ;
 wire \Tile_X1Y9_N2BEGb[4] ;
 wire \Tile_X1Y9_N2BEGb[5] ;
 wire \Tile_X1Y9_N2BEGb[6] ;
 wire \Tile_X1Y9_N2BEGb[7] ;
 wire \Tile_X1Y9_N4BEG[0] ;
 wire \Tile_X1Y9_N4BEG[10] ;
 wire \Tile_X1Y9_N4BEG[11] ;
 wire \Tile_X1Y9_N4BEG[12] ;
 wire \Tile_X1Y9_N4BEG[13] ;
 wire \Tile_X1Y9_N4BEG[14] ;
 wire \Tile_X1Y9_N4BEG[15] ;
 wire \Tile_X1Y9_N4BEG[1] ;
 wire \Tile_X1Y9_N4BEG[2] ;
 wire \Tile_X1Y9_N4BEG[3] ;
 wire \Tile_X1Y9_N4BEG[4] ;
 wire \Tile_X1Y9_N4BEG[5] ;
 wire \Tile_X1Y9_N4BEG[6] ;
 wire \Tile_X1Y9_N4BEG[7] ;
 wire \Tile_X1Y9_N4BEG[8] ;
 wire \Tile_X1Y9_N4BEG[9] ;
 wire \Tile_X1Y9_NN4BEG[0] ;
 wire \Tile_X1Y9_NN4BEG[10] ;
 wire \Tile_X1Y9_NN4BEG[11] ;
 wire \Tile_X1Y9_NN4BEG[12] ;
 wire \Tile_X1Y9_NN4BEG[13] ;
 wire \Tile_X1Y9_NN4BEG[14] ;
 wire \Tile_X1Y9_NN4BEG[15] ;
 wire \Tile_X1Y9_NN4BEG[1] ;
 wire \Tile_X1Y9_NN4BEG[2] ;
 wire \Tile_X1Y9_NN4BEG[3] ;
 wire \Tile_X1Y9_NN4BEG[4] ;
 wire \Tile_X1Y9_NN4BEG[5] ;
 wire \Tile_X1Y9_NN4BEG[6] ;
 wire \Tile_X1Y9_NN4BEG[7] ;
 wire \Tile_X1Y9_NN4BEG[8] ;
 wire \Tile_X1Y9_NN4BEG[9] ;
 wire \Tile_X1Y9_S1BEG[0] ;
 wire \Tile_X1Y9_S1BEG[1] ;
 wire \Tile_X1Y9_S1BEG[2] ;
 wire \Tile_X1Y9_S1BEG[3] ;
 wire \Tile_X1Y9_S2BEG[0] ;
 wire \Tile_X1Y9_S2BEG[1] ;
 wire \Tile_X1Y9_S2BEG[2] ;
 wire \Tile_X1Y9_S2BEG[3] ;
 wire \Tile_X1Y9_S2BEG[4] ;
 wire \Tile_X1Y9_S2BEG[5] ;
 wire \Tile_X1Y9_S2BEG[6] ;
 wire \Tile_X1Y9_S2BEG[7] ;
 wire \Tile_X1Y9_S2BEGb[0] ;
 wire \Tile_X1Y9_S2BEGb[1] ;
 wire \Tile_X1Y9_S2BEGb[2] ;
 wire \Tile_X1Y9_S2BEGb[3] ;
 wire \Tile_X1Y9_S2BEGb[4] ;
 wire \Tile_X1Y9_S2BEGb[5] ;
 wire \Tile_X1Y9_S2BEGb[6] ;
 wire \Tile_X1Y9_S2BEGb[7] ;
 wire \Tile_X1Y9_S4BEG[0] ;
 wire \Tile_X1Y9_S4BEG[10] ;
 wire \Tile_X1Y9_S4BEG[11] ;
 wire \Tile_X1Y9_S4BEG[12] ;
 wire \Tile_X1Y9_S4BEG[13] ;
 wire \Tile_X1Y9_S4BEG[14] ;
 wire \Tile_X1Y9_S4BEG[15] ;
 wire \Tile_X1Y9_S4BEG[1] ;
 wire \Tile_X1Y9_S4BEG[2] ;
 wire \Tile_X1Y9_S4BEG[3] ;
 wire \Tile_X1Y9_S4BEG[4] ;
 wire \Tile_X1Y9_S4BEG[5] ;
 wire \Tile_X1Y9_S4BEG[6] ;
 wire \Tile_X1Y9_S4BEG[7] ;
 wire \Tile_X1Y9_S4BEG[8] ;
 wire \Tile_X1Y9_S4BEG[9] ;
 wire \Tile_X1Y9_SS4BEG[0] ;
 wire \Tile_X1Y9_SS4BEG[10] ;
 wire \Tile_X1Y9_SS4BEG[11] ;
 wire \Tile_X1Y9_SS4BEG[12] ;
 wire \Tile_X1Y9_SS4BEG[13] ;
 wire \Tile_X1Y9_SS4BEG[14] ;
 wire \Tile_X1Y9_SS4BEG[15] ;
 wire \Tile_X1Y9_SS4BEG[1] ;
 wire \Tile_X1Y9_SS4BEG[2] ;
 wire \Tile_X1Y9_SS4BEG[3] ;
 wire \Tile_X1Y9_SS4BEG[4] ;
 wire \Tile_X1Y9_SS4BEG[5] ;
 wire \Tile_X1Y9_SS4BEG[6] ;
 wire \Tile_X1Y9_SS4BEG[7] ;
 wire \Tile_X1Y9_SS4BEG[8] ;
 wire \Tile_X1Y9_SS4BEG[9] ;
 wire Tile_X1Y9_UserCLKo;
 wire \Tile_X1Y9_W1BEG[0] ;
 wire \Tile_X1Y9_W1BEG[1] ;
 wire \Tile_X1Y9_W1BEG[2] ;
 wire \Tile_X1Y9_W1BEG[3] ;
 wire \Tile_X1Y9_W2BEG[0] ;
 wire \Tile_X1Y9_W2BEG[1] ;
 wire \Tile_X1Y9_W2BEG[2] ;
 wire \Tile_X1Y9_W2BEG[3] ;
 wire \Tile_X1Y9_W2BEG[4] ;
 wire \Tile_X1Y9_W2BEG[5] ;
 wire \Tile_X1Y9_W2BEG[6] ;
 wire \Tile_X1Y9_W2BEG[7] ;
 wire \Tile_X1Y9_W2BEGb[0] ;
 wire \Tile_X1Y9_W2BEGb[1] ;
 wire \Tile_X1Y9_W2BEGb[2] ;
 wire \Tile_X1Y9_W2BEGb[3] ;
 wire \Tile_X1Y9_W2BEGb[4] ;
 wire \Tile_X1Y9_W2BEGb[5] ;
 wire \Tile_X1Y9_W2BEGb[6] ;
 wire \Tile_X1Y9_W2BEGb[7] ;
 wire \Tile_X1Y9_W6BEG[0] ;
 wire \Tile_X1Y9_W6BEG[10] ;
 wire \Tile_X1Y9_W6BEG[11] ;
 wire \Tile_X1Y9_W6BEG[1] ;
 wire \Tile_X1Y9_W6BEG[2] ;
 wire \Tile_X1Y9_W6BEG[3] ;
 wire \Tile_X1Y9_W6BEG[4] ;
 wire \Tile_X1Y9_W6BEG[5] ;
 wire \Tile_X1Y9_W6BEG[6] ;
 wire \Tile_X1Y9_W6BEG[7] ;
 wire \Tile_X1Y9_W6BEG[8] ;
 wire \Tile_X1Y9_W6BEG[9] ;
 wire \Tile_X1Y9_WW4BEG[0] ;
 wire \Tile_X1Y9_WW4BEG[10] ;
 wire \Tile_X1Y9_WW4BEG[11] ;
 wire \Tile_X1Y9_WW4BEG[12] ;
 wire \Tile_X1Y9_WW4BEG[13] ;
 wire \Tile_X1Y9_WW4BEG[14] ;
 wire \Tile_X1Y9_WW4BEG[15] ;
 wire \Tile_X1Y9_WW4BEG[1] ;
 wire \Tile_X1Y9_WW4BEG[2] ;
 wire \Tile_X1Y9_WW4BEG[3] ;
 wire \Tile_X1Y9_WW4BEG[4] ;
 wire \Tile_X1Y9_WW4BEG[5] ;
 wire \Tile_X1Y9_WW4BEG[6] ;
 wire \Tile_X1Y9_WW4BEG[7] ;
 wire \Tile_X1Y9_WW4BEG[8] ;
 wire \Tile_X1Y9_WW4BEG[9] ;
 wire \Tile_X2Y0_FrameData_O[0] ;
 wire \Tile_X2Y0_FrameData_O[10] ;
 wire \Tile_X2Y0_FrameData_O[11] ;
 wire \Tile_X2Y0_FrameData_O[12] ;
 wire \Tile_X2Y0_FrameData_O[13] ;
 wire \Tile_X2Y0_FrameData_O[14] ;
 wire \Tile_X2Y0_FrameData_O[15] ;
 wire \Tile_X2Y0_FrameData_O[16] ;
 wire \Tile_X2Y0_FrameData_O[17] ;
 wire \Tile_X2Y0_FrameData_O[18] ;
 wire \Tile_X2Y0_FrameData_O[19] ;
 wire \Tile_X2Y0_FrameData_O[1] ;
 wire \Tile_X2Y0_FrameData_O[20] ;
 wire \Tile_X2Y0_FrameData_O[21] ;
 wire \Tile_X2Y0_FrameData_O[22] ;
 wire \Tile_X2Y0_FrameData_O[23] ;
 wire \Tile_X2Y0_FrameData_O[24] ;
 wire \Tile_X2Y0_FrameData_O[25] ;
 wire \Tile_X2Y0_FrameData_O[26] ;
 wire \Tile_X2Y0_FrameData_O[27] ;
 wire \Tile_X2Y0_FrameData_O[28] ;
 wire \Tile_X2Y0_FrameData_O[29] ;
 wire \Tile_X2Y0_FrameData_O[2] ;
 wire \Tile_X2Y0_FrameData_O[30] ;
 wire \Tile_X2Y0_FrameData_O[31] ;
 wire \Tile_X2Y0_FrameData_O[3] ;
 wire \Tile_X2Y0_FrameData_O[4] ;
 wire \Tile_X2Y0_FrameData_O[5] ;
 wire \Tile_X2Y0_FrameData_O[6] ;
 wire \Tile_X2Y0_FrameData_O[7] ;
 wire \Tile_X2Y0_FrameData_O[8] ;
 wire \Tile_X2Y0_FrameData_O[9] ;
 wire \Tile_X2Y0_FrameStrobe_O[0] ;
 wire \Tile_X2Y0_FrameStrobe_O[10] ;
 wire \Tile_X2Y0_FrameStrobe_O[11] ;
 wire \Tile_X2Y0_FrameStrobe_O[12] ;
 wire \Tile_X2Y0_FrameStrobe_O[13] ;
 wire \Tile_X2Y0_FrameStrobe_O[14] ;
 wire \Tile_X2Y0_FrameStrobe_O[15] ;
 wire \Tile_X2Y0_FrameStrobe_O[16] ;
 wire \Tile_X2Y0_FrameStrobe_O[17] ;
 wire \Tile_X2Y0_FrameStrobe_O[18] ;
 wire \Tile_X2Y0_FrameStrobe_O[19] ;
 wire \Tile_X2Y0_FrameStrobe_O[1] ;
 wire \Tile_X2Y0_FrameStrobe_O[2] ;
 wire \Tile_X2Y0_FrameStrobe_O[3] ;
 wire \Tile_X2Y0_FrameStrobe_O[4] ;
 wire \Tile_X2Y0_FrameStrobe_O[5] ;
 wire \Tile_X2Y0_FrameStrobe_O[6] ;
 wire \Tile_X2Y0_FrameStrobe_O[7] ;
 wire \Tile_X2Y0_FrameStrobe_O[8] ;
 wire \Tile_X2Y0_FrameStrobe_O[9] ;
 wire \Tile_X2Y0_S1BEG[0] ;
 wire \Tile_X2Y0_S1BEG[1] ;
 wire \Tile_X2Y0_S1BEG[2] ;
 wire \Tile_X2Y0_S1BEG[3] ;
 wire \Tile_X2Y0_S2BEG[0] ;
 wire \Tile_X2Y0_S2BEG[1] ;
 wire \Tile_X2Y0_S2BEG[2] ;
 wire \Tile_X2Y0_S2BEG[3] ;
 wire \Tile_X2Y0_S2BEG[4] ;
 wire \Tile_X2Y0_S2BEG[5] ;
 wire \Tile_X2Y0_S2BEG[6] ;
 wire \Tile_X2Y0_S2BEG[7] ;
 wire \Tile_X2Y0_S2BEGb[0] ;
 wire \Tile_X2Y0_S2BEGb[1] ;
 wire \Tile_X2Y0_S2BEGb[2] ;
 wire \Tile_X2Y0_S2BEGb[3] ;
 wire \Tile_X2Y0_S2BEGb[4] ;
 wire \Tile_X2Y0_S2BEGb[5] ;
 wire \Tile_X2Y0_S2BEGb[6] ;
 wire \Tile_X2Y0_S2BEGb[7] ;
 wire \Tile_X2Y0_S4BEG[0] ;
 wire \Tile_X2Y0_S4BEG[10] ;
 wire \Tile_X2Y0_S4BEG[11] ;
 wire \Tile_X2Y0_S4BEG[12] ;
 wire \Tile_X2Y0_S4BEG[13] ;
 wire \Tile_X2Y0_S4BEG[14] ;
 wire \Tile_X2Y0_S4BEG[15] ;
 wire \Tile_X2Y0_S4BEG[1] ;
 wire \Tile_X2Y0_S4BEG[2] ;
 wire \Tile_X2Y0_S4BEG[3] ;
 wire \Tile_X2Y0_S4BEG[4] ;
 wire \Tile_X2Y0_S4BEG[5] ;
 wire \Tile_X2Y0_S4BEG[6] ;
 wire \Tile_X2Y0_S4BEG[7] ;
 wire \Tile_X2Y0_S4BEG[8] ;
 wire \Tile_X2Y0_S4BEG[9] ;
 wire \Tile_X2Y0_SS4BEG[0] ;
 wire \Tile_X2Y0_SS4BEG[10] ;
 wire \Tile_X2Y0_SS4BEG[11] ;
 wire \Tile_X2Y0_SS4BEG[12] ;
 wire \Tile_X2Y0_SS4BEG[13] ;
 wire \Tile_X2Y0_SS4BEG[14] ;
 wire \Tile_X2Y0_SS4BEG[15] ;
 wire \Tile_X2Y0_SS4BEG[1] ;
 wire \Tile_X2Y0_SS4BEG[2] ;
 wire \Tile_X2Y0_SS4BEG[3] ;
 wire \Tile_X2Y0_SS4BEG[4] ;
 wire \Tile_X2Y0_SS4BEG[5] ;
 wire \Tile_X2Y0_SS4BEG[6] ;
 wire \Tile_X2Y0_SS4BEG[7] ;
 wire \Tile_X2Y0_SS4BEG[8] ;
 wire \Tile_X2Y0_SS4BEG[9] ;
 wire Tile_X2Y0_UserCLKo;
 wire Tile_X2Y10_Co;
 wire \Tile_X2Y10_E1BEG[0] ;
 wire \Tile_X2Y10_E1BEG[1] ;
 wire \Tile_X2Y10_E1BEG[2] ;
 wire \Tile_X2Y10_E1BEG[3] ;
 wire \Tile_X2Y10_E2BEG[0] ;
 wire \Tile_X2Y10_E2BEG[1] ;
 wire \Tile_X2Y10_E2BEG[2] ;
 wire \Tile_X2Y10_E2BEG[3] ;
 wire \Tile_X2Y10_E2BEG[4] ;
 wire \Tile_X2Y10_E2BEG[5] ;
 wire \Tile_X2Y10_E2BEG[6] ;
 wire \Tile_X2Y10_E2BEG[7] ;
 wire \Tile_X2Y10_E2BEGb[0] ;
 wire \Tile_X2Y10_E2BEGb[1] ;
 wire \Tile_X2Y10_E2BEGb[2] ;
 wire \Tile_X2Y10_E2BEGb[3] ;
 wire \Tile_X2Y10_E2BEGb[4] ;
 wire \Tile_X2Y10_E2BEGb[5] ;
 wire \Tile_X2Y10_E2BEGb[6] ;
 wire \Tile_X2Y10_E2BEGb[7] ;
 wire \Tile_X2Y10_E6BEG[0] ;
 wire \Tile_X2Y10_E6BEG[10] ;
 wire \Tile_X2Y10_E6BEG[11] ;
 wire \Tile_X2Y10_E6BEG[1] ;
 wire \Tile_X2Y10_E6BEG[2] ;
 wire \Tile_X2Y10_E6BEG[3] ;
 wire \Tile_X2Y10_E6BEG[4] ;
 wire \Tile_X2Y10_E6BEG[5] ;
 wire \Tile_X2Y10_E6BEG[6] ;
 wire \Tile_X2Y10_E6BEG[7] ;
 wire \Tile_X2Y10_E6BEG[8] ;
 wire \Tile_X2Y10_E6BEG[9] ;
 wire \Tile_X2Y10_EE4BEG[0] ;
 wire \Tile_X2Y10_EE4BEG[10] ;
 wire \Tile_X2Y10_EE4BEG[11] ;
 wire \Tile_X2Y10_EE4BEG[12] ;
 wire \Tile_X2Y10_EE4BEG[13] ;
 wire \Tile_X2Y10_EE4BEG[14] ;
 wire \Tile_X2Y10_EE4BEG[15] ;
 wire \Tile_X2Y10_EE4BEG[1] ;
 wire \Tile_X2Y10_EE4BEG[2] ;
 wire \Tile_X2Y10_EE4BEG[3] ;
 wire \Tile_X2Y10_EE4BEG[4] ;
 wire \Tile_X2Y10_EE4BEG[5] ;
 wire \Tile_X2Y10_EE4BEG[6] ;
 wire \Tile_X2Y10_EE4BEG[7] ;
 wire \Tile_X2Y10_EE4BEG[8] ;
 wire \Tile_X2Y10_EE4BEG[9] ;
 wire \Tile_X2Y10_FrameData_O[0] ;
 wire \Tile_X2Y10_FrameData_O[10] ;
 wire \Tile_X2Y10_FrameData_O[11] ;
 wire \Tile_X2Y10_FrameData_O[12] ;
 wire \Tile_X2Y10_FrameData_O[13] ;
 wire \Tile_X2Y10_FrameData_O[14] ;
 wire \Tile_X2Y10_FrameData_O[15] ;
 wire \Tile_X2Y10_FrameData_O[16] ;
 wire \Tile_X2Y10_FrameData_O[17] ;
 wire \Tile_X2Y10_FrameData_O[18] ;
 wire \Tile_X2Y10_FrameData_O[19] ;
 wire \Tile_X2Y10_FrameData_O[1] ;
 wire \Tile_X2Y10_FrameData_O[20] ;
 wire \Tile_X2Y10_FrameData_O[21] ;
 wire \Tile_X2Y10_FrameData_O[22] ;
 wire \Tile_X2Y10_FrameData_O[23] ;
 wire \Tile_X2Y10_FrameData_O[24] ;
 wire \Tile_X2Y10_FrameData_O[25] ;
 wire \Tile_X2Y10_FrameData_O[26] ;
 wire \Tile_X2Y10_FrameData_O[27] ;
 wire \Tile_X2Y10_FrameData_O[28] ;
 wire \Tile_X2Y10_FrameData_O[29] ;
 wire \Tile_X2Y10_FrameData_O[2] ;
 wire \Tile_X2Y10_FrameData_O[30] ;
 wire \Tile_X2Y10_FrameData_O[31] ;
 wire \Tile_X2Y10_FrameData_O[3] ;
 wire \Tile_X2Y10_FrameData_O[4] ;
 wire \Tile_X2Y10_FrameData_O[5] ;
 wire \Tile_X2Y10_FrameData_O[6] ;
 wire \Tile_X2Y10_FrameData_O[7] ;
 wire \Tile_X2Y10_FrameData_O[8] ;
 wire \Tile_X2Y10_FrameData_O[9] ;
 wire \Tile_X2Y10_FrameStrobe_O[0] ;
 wire \Tile_X2Y10_FrameStrobe_O[10] ;
 wire \Tile_X2Y10_FrameStrobe_O[11] ;
 wire \Tile_X2Y10_FrameStrobe_O[12] ;
 wire \Tile_X2Y10_FrameStrobe_O[13] ;
 wire \Tile_X2Y10_FrameStrobe_O[14] ;
 wire \Tile_X2Y10_FrameStrobe_O[15] ;
 wire \Tile_X2Y10_FrameStrobe_O[16] ;
 wire \Tile_X2Y10_FrameStrobe_O[17] ;
 wire \Tile_X2Y10_FrameStrobe_O[18] ;
 wire \Tile_X2Y10_FrameStrobe_O[19] ;
 wire \Tile_X2Y10_FrameStrobe_O[1] ;
 wire \Tile_X2Y10_FrameStrobe_O[2] ;
 wire \Tile_X2Y10_FrameStrobe_O[3] ;
 wire \Tile_X2Y10_FrameStrobe_O[4] ;
 wire \Tile_X2Y10_FrameStrobe_O[5] ;
 wire \Tile_X2Y10_FrameStrobe_O[6] ;
 wire \Tile_X2Y10_FrameStrobe_O[7] ;
 wire \Tile_X2Y10_FrameStrobe_O[8] ;
 wire \Tile_X2Y10_FrameStrobe_O[9] ;
 wire \Tile_X2Y10_N1BEG[0] ;
 wire \Tile_X2Y10_N1BEG[1] ;
 wire \Tile_X2Y10_N1BEG[2] ;
 wire \Tile_X2Y10_N1BEG[3] ;
 wire \Tile_X2Y10_N2BEG[0] ;
 wire \Tile_X2Y10_N2BEG[1] ;
 wire \Tile_X2Y10_N2BEG[2] ;
 wire \Tile_X2Y10_N2BEG[3] ;
 wire \Tile_X2Y10_N2BEG[4] ;
 wire \Tile_X2Y10_N2BEG[5] ;
 wire \Tile_X2Y10_N2BEG[6] ;
 wire \Tile_X2Y10_N2BEG[7] ;
 wire \Tile_X2Y10_N2BEGb[0] ;
 wire \Tile_X2Y10_N2BEGb[1] ;
 wire \Tile_X2Y10_N2BEGb[2] ;
 wire \Tile_X2Y10_N2BEGb[3] ;
 wire \Tile_X2Y10_N2BEGb[4] ;
 wire \Tile_X2Y10_N2BEGb[5] ;
 wire \Tile_X2Y10_N2BEGb[6] ;
 wire \Tile_X2Y10_N2BEGb[7] ;
 wire \Tile_X2Y10_N4BEG[0] ;
 wire \Tile_X2Y10_N4BEG[10] ;
 wire \Tile_X2Y10_N4BEG[11] ;
 wire \Tile_X2Y10_N4BEG[12] ;
 wire \Tile_X2Y10_N4BEG[13] ;
 wire \Tile_X2Y10_N4BEG[14] ;
 wire \Tile_X2Y10_N4BEG[15] ;
 wire \Tile_X2Y10_N4BEG[1] ;
 wire \Tile_X2Y10_N4BEG[2] ;
 wire \Tile_X2Y10_N4BEG[3] ;
 wire \Tile_X2Y10_N4BEG[4] ;
 wire \Tile_X2Y10_N4BEG[5] ;
 wire \Tile_X2Y10_N4BEG[6] ;
 wire \Tile_X2Y10_N4BEG[7] ;
 wire \Tile_X2Y10_N4BEG[8] ;
 wire \Tile_X2Y10_N4BEG[9] ;
 wire \Tile_X2Y10_NN4BEG[0] ;
 wire \Tile_X2Y10_NN4BEG[10] ;
 wire \Tile_X2Y10_NN4BEG[11] ;
 wire \Tile_X2Y10_NN4BEG[12] ;
 wire \Tile_X2Y10_NN4BEG[13] ;
 wire \Tile_X2Y10_NN4BEG[14] ;
 wire \Tile_X2Y10_NN4BEG[15] ;
 wire \Tile_X2Y10_NN4BEG[1] ;
 wire \Tile_X2Y10_NN4BEG[2] ;
 wire \Tile_X2Y10_NN4BEG[3] ;
 wire \Tile_X2Y10_NN4BEG[4] ;
 wire \Tile_X2Y10_NN4BEG[5] ;
 wire \Tile_X2Y10_NN4BEG[6] ;
 wire \Tile_X2Y10_NN4BEG[7] ;
 wire \Tile_X2Y10_NN4BEG[8] ;
 wire \Tile_X2Y10_NN4BEG[9] ;
 wire \Tile_X2Y10_S1BEG[0] ;
 wire \Tile_X2Y10_S1BEG[1] ;
 wire \Tile_X2Y10_S1BEG[2] ;
 wire \Tile_X2Y10_S1BEG[3] ;
 wire \Tile_X2Y10_S2BEG[0] ;
 wire \Tile_X2Y10_S2BEG[1] ;
 wire \Tile_X2Y10_S2BEG[2] ;
 wire \Tile_X2Y10_S2BEG[3] ;
 wire \Tile_X2Y10_S2BEG[4] ;
 wire \Tile_X2Y10_S2BEG[5] ;
 wire \Tile_X2Y10_S2BEG[6] ;
 wire \Tile_X2Y10_S2BEG[7] ;
 wire \Tile_X2Y10_S2BEGb[0] ;
 wire \Tile_X2Y10_S2BEGb[1] ;
 wire \Tile_X2Y10_S2BEGb[2] ;
 wire \Tile_X2Y10_S2BEGb[3] ;
 wire \Tile_X2Y10_S2BEGb[4] ;
 wire \Tile_X2Y10_S2BEGb[5] ;
 wire \Tile_X2Y10_S2BEGb[6] ;
 wire \Tile_X2Y10_S2BEGb[7] ;
 wire \Tile_X2Y10_S4BEG[0] ;
 wire \Tile_X2Y10_S4BEG[10] ;
 wire \Tile_X2Y10_S4BEG[11] ;
 wire \Tile_X2Y10_S4BEG[12] ;
 wire \Tile_X2Y10_S4BEG[13] ;
 wire \Tile_X2Y10_S4BEG[14] ;
 wire \Tile_X2Y10_S4BEG[15] ;
 wire \Tile_X2Y10_S4BEG[1] ;
 wire \Tile_X2Y10_S4BEG[2] ;
 wire \Tile_X2Y10_S4BEG[3] ;
 wire \Tile_X2Y10_S4BEG[4] ;
 wire \Tile_X2Y10_S4BEG[5] ;
 wire \Tile_X2Y10_S4BEG[6] ;
 wire \Tile_X2Y10_S4BEG[7] ;
 wire \Tile_X2Y10_S4BEG[8] ;
 wire \Tile_X2Y10_S4BEG[9] ;
 wire \Tile_X2Y10_SS4BEG[0] ;
 wire \Tile_X2Y10_SS4BEG[10] ;
 wire \Tile_X2Y10_SS4BEG[11] ;
 wire \Tile_X2Y10_SS4BEG[12] ;
 wire \Tile_X2Y10_SS4BEG[13] ;
 wire \Tile_X2Y10_SS4BEG[14] ;
 wire \Tile_X2Y10_SS4BEG[15] ;
 wire \Tile_X2Y10_SS4BEG[1] ;
 wire \Tile_X2Y10_SS4BEG[2] ;
 wire \Tile_X2Y10_SS4BEG[3] ;
 wire \Tile_X2Y10_SS4BEG[4] ;
 wire \Tile_X2Y10_SS4BEG[5] ;
 wire \Tile_X2Y10_SS4BEG[6] ;
 wire \Tile_X2Y10_SS4BEG[7] ;
 wire \Tile_X2Y10_SS4BEG[8] ;
 wire \Tile_X2Y10_SS4BEG[9] ;
 wire Tile_X2Y10_UserCLKo;
 wire \Tile_X2Y10_W1BEG[0] ;
 wire \Tile_X2Y10_W1BEG[1] ;
 wire \Tile_X2Y10_W1BEG[2] ;
 wire \Tile_X2Y10_W1BEG[3] ;
 wire \Tile_X2Y10_W2BEG[0] ;
 wire \Tile_X2Y10_W2BEG[1] ;
 wire \Tile_X2Y10_W2BEG[2] ;
 wire \Tile_X2Y10_W2BEG[3] ;
 wire \Tile_X2Y10_W2BEG[4] ;
 wire \Tile_X2Y10_W2BEG[5] ;
 wire \Tile_X2Y10_W2BEG[6] ;
 wire \Tile_X2Y10_W2BEG[7] ;
 wire \Tile_X2Y10_W2BEGb[0] ;
 wire \Tile_X2Y10_W2BEGb[1] ;
 wire \Tile_X2Y10_W2BEGb[2] ;
 wire \Tile_X2Y10_W2BEGb[3] ;
 wire \Tile_X2Y10_W2BEGb[4] ;
 wire \Tile_X2Y10_W2BEGb[5] ;
 wire \Tile_X2Y10_W2BEGb[6] ;
 wire \Tile_X2Y10_W2BEGb[7] ;
 wire \Tile_X2Y10_W6BEG[0] ;
 wire \Tile_X2Y10_W6BEG[10] ;
 wire \Tile_X2Y10_W6BEG[11] ;
 wire \Tile_X2Y10_W6BEG[1] ;
 wire \Tile_X2Y10_W6BEG[2] ;
 wire \Tile_X2Y10_W6BEG[3] ;
 wire \Tile_X2Y10_W6BEG[4] ;
 wire \Tile_X2Y10_W6BEG[5] ;
 wire \Tile_X2Y10_W6BEG[6] ;
 wire \Tile_X2Y10_W6BEG[7] ;
 wire \Tile_X2Y10_W6BEG[8] ;
 wire \Tile_X2Y10_W6BEG[9] ;
 wire \Tile_X2Y10_WW4BEG[0] ;
 wire \Tile_X2Y10_WW4BEG[10] ;
 wire \Tile_X2Y10_WW4BEG[11] ;
 wire \Tile_X2Y10_WW4BEG[12] ;
 wire \Tile_X2Y10_WW4BEG[13] ;
 wire \Tile_X2Y10_WW4BEG[14] ;
 wire \Tile_X2Y10_WW4BEG[15] ;
 wire \Tile_X2Y10_WW4BEG[1] ;
 wire \Tile_X2Y10_WW4BEG[2] ;
 wire \Tile_X2Y10_WW4BEG[3] ;
 wire \Tile_X2Y10_WW4BEG[4] ;
 wire \Tile_X2Y10_WW4BEG[5] ;
 wire \Tile_X2Y10_WW4BEG[6] ;
 wire \Tile_X2Y10_WW4BEG[7] ;
 wire \Tile_X2Y10_WW4BEG[8] ;
 wire \Tile_X2Y10_WW4BEG[9] ;
 wire Tile_X2Y11_Co;
 wire \Tile_X2Y11_E1BEG[0] ;
 wire \Tile_X2Y11_E1BEG[1] ;
 wire \Tile_X2Y11_E1BEG[2] ;
 wire \Tile_X2Y11_E1BEG[3] ;
 wire \Tile_X2Y11_E2BEG[0] ;
 wire \Tile_X2Y11_E2BEG[1] ;
 wire \Tile_X2Y11_E2BEG[2] ;
 wire \Tile_X2Y11_E2BEG[3] ;
 wire \Tile_X2Y11_E2BEG[4] ;
 wire \Tile_X2Y11_E2BEG[5] ;
 wire \Tile_X2Y11_E2BEG[6] ;
 wire \Tile_X2Y11_E2BEG[7] ;
 wire \Tile_X2Y11_E2BEGb[0] ;
 wire \Tile_X2Y11_E2BEGb[1] ;
 wire \Tile_X2Y11_E2BEGb[2] ;
 wire \Tile_X2Y11_E2BEGb[3] ;
 wire \Tile_X2Y11_E2BEGb[4] ;
 wire \Tile_X2Y11_E2BEGb[5] ;
 wire \Tile_X2Y11_E2BEGb[6] ;
 wire \Tile_X2Y11_E2BEGb[7] ;
 wire \Tile_X2Y11_E6BEG[0] ;
 wire \Tile_X2Y11_E6BEG[10] ;
 wire \Tile_X2Y11_E6BEG[11] ;
 wire \Tile_X2Y11_E6BEG[1] ;
 wire \Tile_X2Y11_E6BEG[2] ;
 wire \Tile_X2Y11_E6BEG[3] ;
 wire \Tile_X2Y11_E6BEG[4] ;
 wire \Tile_X2Y11_E6BEG[5] ;
 wire \Tile_X2Y11_E6BEG[6] ;
 wire \Tile_X2Y11_E6BEG[7] ;
 wire \Tile_X2Y11_E6BEG[8] ;
 wire \Tile_X2Y11_E6BEG[9] ;
 wire \Tile_X2Y11_EE4BEG[0] ;
 wire \Tile_X2Y11_EE4BEG[10] ;
 wire \Tile_X2Y11_EE4BEG[11] ;
 wire \Tile_X2Y11_EE4BEG[12] ;
 wire \Tile_X2Y11_EE4BEG[13] ;
 wire \Tile_X2Y11_EE4BEG[14] ;
 wire \Tile_X2Y11_EE4BEG[15] ;
 wire \Tile_X2Y11_EE4BEG[1] ;
 wire \Tile_X2Y11_EE4BEG[2] ;
 wire \Tile_X2Y11_EE4BEG[3] ;
 wire \Tile_X2Y11_EE4BEG[4] ;
 wire \Tile_X2Y11_EE4BEG[5] ;
 wire \Tile_X2Y11_EE4BEG[6] ;
 wire \Tile_X2Y11_EE4BEG[7] ;
 wire \Tile_X2Y11_EE4BEG[8] ;
 wire \Tile_X2Y11_EE4BEG[9] ;
 wire \Tile_X2Y11_FrameData_O[0] ;
 wire \Tile_X2Y11_FrameData_O[10] ;
 wire \Tile_X2Y11_FrameData_O[11] ;
 wire \Tile_X2Y11_FrameData_O[12] ;
 wire \Tile_X2Y11_FrameData_O[13] ;
 wire \Tile_X2Y11_FrameData_O[14] ;
 wire \Tile_X2Y11_FrameData_O[15] ;
 wire \Tile_X2Y11_FrameData_O[16] ;
 wire \Tile_X2Y11_FrameData_O[17] ;
 wire \Tile_X2Y11_FrameData_O[18] ;
 wire \Tile_X2Y11_FrameData_O[19] ;
 wire \Tile_X2Y11_FrameData_O[1] ;
 wire \Tile_X2Y11_FrameData_O[20] ;
 wire \Tile_X2Y11_FrameData_O[21] ;
 wire \Tile_X2Y11_FrameData_O[22] ;
 wire \Tile_X2Y11_FrameData_O[23] ;
 wire \Tile_X2Y11_FrameData_O[24] ;
 wire \Tile_X2Y11_FrameData_O[25] ;
 wire \Tile_X2Y11_FrameData_O[26] ;
 wire \Tile_X2Y11_FrameData_O[27] ;
 wire \Tile_X2Y11_FrameData_O[28] ;
 wire \Tile_X2Y11_FrameData_O[29] ;
 wire \Tile_X2Y11_FrameData_O[2] ;
 wire \Tile_X2Y11_FrameData_O[30] ;
 wire \Tile_X2Y11_FrameData_O[31] ;
 wire \Tile_X2Y11_FrameData_O[3] ;
 wire \Tile_X2Y11_FrameData_O[4] ;
 wire \Tile_X2Y11_FrameData_O[5] ;
 wire \Tile_X2Y11_FrameData_O[6] ;
 wire \Tile_X2Y11_FrameData_O[7] ;
 wire \Tile_X2Y11_FrameData_O[8] ;
 wire \Tile_X2Y11_FrameData_O[9] ;
 wire \Tile_X2Y11_FrameStrobe_O[0] ;
 wire \Tile_X2Y11_FrameStrobe_O[10] ;
 wire \Tile_X2Y11_FrameStrobe_O[11] ;
 wire \Tile_X2Y11_FrameStrobe_O[12] ;
 wire \Tile_X2Y11_FrameStrobe_O[13] ;
 wire \Tile_X2Y11_FrameStrobe_O[14] ;
 wire \Tile_X2Y11_FrameStrobe_O[15] ;
 wire \Tile_X2Y11_FrameStrobe_O[16] ;
 wire \Tile_X2Y11_FrameStrobe_O[17] ;
 wire \Tile_X2Y11_FrameStrobe_O[18] ;
 wire \Tile_X2Y11_FrameStrobe_O[19] ;
 wire \Tile_X2Y11_FrameStrobe_O[1] ;
 wire \Tile_X2Y11_FrameStrobe_O[2] ;
 wire \Tile_X2Y11_FrameStrobe_O[3] ;
 wire \Tile_X2Y11_FrameStrobe_O[4] ;
 wire \Tile_X2Y11_FrameStrobe_O[5] ;
 wire \Tile_X2Y11_FrameStrobe_O[6] ;
 wire \Tile_X2Y11_FrameStrobe_O[7] ;
 wire \Tile_X2Y11_FrameStrobe_O[8] ;
 wire \Tile_X2Y11_FrameStrobe_O[9] ;
 wire \Tile_X2Y11_N1BEG[0] ;
 wire \Tile_X2Y11_N1BEG[1] ;
 wire \Tile_X2Y11_N1BEG[2] ;
 wire \Tile_X2Y11_N1BEG[3] ;
 wire \Tile_X2Y11_N2BEG[0] ;
 wire \Tile_X2Y11_N2BEG[1] ;
 wire \Tile_X2Y11_N2BEG[2] ;
 wire \Tile_X2Y11_N2BEG[3] ;
 wire \Tile_X2Y11_N2BEG[4] ;
 wire \Tile_X2Y11_N2BEG[5] ;
 wire \Tile_X2Y11_N2BEG[6] ;
 wire \Tile_X2Y11_N2BEG[7] ;
 wire \Tile_X2Y11_N2BEGb[0] ;
 wire \Tile_X2Y11_N2BEGb[1] ;
 wire \Tile_X2Y11_N2BEGb[2] ;
 wire \Tile_X2Y11_N2BEGb[3] ;
 wire \Tile_X2Y11_N2BEGb[4] ;
 wire \Tile_X2Y11_N2BEGb[5] ;
 wire \Tile_X2Y11_N2BEGb[6] ;
 wire \Tile_X2Y11_N2BEGb[7] ;
 wire \Tile_X2Y11_N4BEG[0] ;
 wire \Tile_X2Y11_N4BEG[10] ;
 wire \Tile_X2Y11_N4BEG[11] ;
 wire \Tile_X2Y11_N4BEG[12] ;
 wire \Tile_X2Y11_N4BEG[13] ;
 wire \Tile_X2Y11_N4BEG[14] ;
 wire \Tile_X2Y11_N4BEG[15] ;
 wire \Tile_X2Y11_N4BEG[1] ;
 wire \Tile_X2Y11_N4BEG[2] ;
 wire \Tile_X2Y11_N4BEG[3] ;
 wire \Tile_X2Y11_N4BEG[4] ;
 wire \Tile_X2Y11_N4BEG[5] ;
 wire \Tile_X2Y11_N4BEG[6] ;
 wire \Tile_X2Y11_N4BEG[7] ;
 wire \Tile_X2Y11_N4BEG[8] ;
 wire \Tile_X2Y11_N4BEG[9] ;
 wire \Tile_X2Y11_NN4BEG[0] ;
 wire \Tile_X2Y11_NN4BEG[10] ;
 wire \Tile_X2Y11_NN4BEG[11] ;
 wire \Tile_X2Y11_NN4BEG[12] ;
 wire \Tile_X2Y11_NN4BEG[13] ;
 wire \Tile_X2Y11_NN4BEG[14] ;
 wire \Tile_X2Y11_NN4BEG[15] ;
 wire \Tile_X2Y11_NN4BEG[1] ;
 wire \Tile_X2Y11_NN4BEG[2] ;
 wire \Tile_X2Y11_NN4BEG[3] ;
 wire \Tile_X2Y11_NN4BEG[4] ;
 wire \Tile_X2Y11_NN4BEG[5] ;
 wire \Tile_X2Y11_NN4BEG[6] ;
 wire \Tile_X2Y11_NN4BEG[7] ;
 wire \Tile_X2Y11_NN4BEG[8] ;
 wire \Tile_X2Y11_NN4BEG[9] ;
 wire \Tile_X2Y11_S1BEG[0] ;
 wire \Tile_X2Y11_S1BEG[1] ;
 wire \Tile_X2Y11_S1BEG[2] ;
 wire \Tile_X2Y11_S1BEG[3] ;
 wire \Tile_X2Y11_S2BEG[0] ;
 wire \Tile_X2Y11_S2BEG[1] ;
 wire \Tile_X2Y11_S2BEG[2] ;
 wire \Tile_X2Y11_S2BEG[3] ;
 wire \Tile_X2Y11_S2BEG[4] ;
 wire \Tile_X2Y11_S2BEG[5] ;
 wire \Tile_X2Y11_S2BEG[6] ;
 wire \Tile_X2Y11_S2BEG[7] ;
 wire \Tile_X2Y11_S2BEGb[0] ;
 wire \Tile_X2Y11_S2BEGb[1] ;
 wire \Tile_X2Y11_S2BEGb[2] ;
 wire \Tile_X2Y11_S2BEGb[3] ;
 wire \Tile_X2Y11_S2BEGb[4] ;
 wire \Tile_X2Y11_S2BEGb[5] ;
 wire \Tile_X2Y11_S2BEGb[6] ;
 wire \Tile_X2Y11_S2BEGb[7] ;
 wire \Tile_X2Y11_S4BEG[0] ;
 wire \Tile_X2Y11_S4BEG[10] ;
 wire \Tile_X2Y11_S4BEG[11] ;
 wire \Tile_X2Y11_S4BEG[12] ;
 wire \Tile_X2Y11_S4BEG[13] ;
 wire \Tile_X2Y11_S4BEG[14] ;
 wire \Tile_X2Y11_S4BEG[15] ;
 wire \Tile_X2Y11_S4BEG[1] ;
 wire \Tile_X2Y11_S4BEG[2] ;
 wire \Tile_X2Y11_S4BEG[3] ;
 wire \Tile_X2Y11_S4BEG[4] ;
 wire \Tile_X2Y11_S4BEG[5] ;
 wire \Tile_X2Y11_S4BEG[6] ;
 wire \Tile_X2Y11_S4BEG[7] ;
 wire \Tile_X2Y11_S4BEG[8] ;
 wire \Tile_X2Y11_S4BEG[9] ;
 wire \Tile_X2Y11_SS4BEG[0] ;
 wire \Tile_X2Y11_SS4BEG[10] ;
 wire \Tile_X2Y11_SS4BEG[11] ;
 wire \Tile_X2Y11_SS4BEG[12] ;
 wire \Tile_X2Y11_SS4BEG[13] ;
 wire \Tile_X2Y11_SS4BEG[14] ;
 wire \Tile_X2Y11_SS4BEG[15] ;
 wire \Tile_X2Y11_SS4BEG[1] ;
 wire \Tile_X2Y11_SS4BEG[2] ;
 wire \Tile_X2Y11_SS4BEG[3] ;
 wire \Tile_X2Y11_SS4BEG[4] ;
 wire \Tile_X2Y11_SS4BEG[5] ;
 wire \Tile_X2Y11_SS4BEG[6] ;
 wire \Tile_X2Y11_SS4BEG[7] ;
 wire \Tile_X2Y11_SS4BEG[8] ;
 wire \Tile_X2Y11_SS4BEG[9] ;
 wire Tile_X2Y11_UserCLKo;
 wire \Tile_X2Y11_W1BEG[0] ;
 wire \Tile_X2Y11_W1BEG[1] ;
 wire \Tile_X2Y11_W1BEG[2] ;
 wire \Tile_X2Y11_W1BEG[3] ;
 wire \Tile_X2Y11_W2BEG[0] ;
 wire \Tile_X2Y11_W2BEG[1] ;
 wire \Tile_X2Y11_W2BEG[2] ;
 wire \Tile_X2Y11_W2BEG[3] ;
 wire \Tile_X2Y11_W2BEG[4] ;
 wire \Tile_X2Y11_W2BEG[5] ;
 wire \Tile_X2Y11_W2BEG[6] ;
 wire \Tile_X2Y11_W2BEG[7] ;
 wire \Tile_X2Y11_W2BEGb[0] ;
 wire \Tile_X2Y11_W2BEGb[1] ;
 wire \Tile_X2Y11_W2BEGb[2] ;
 wire \Tile_X2Y11_W2BEGb[3] ;
 wire \Tile_X2Y11_W2BEGb[4] ;
 wire \Tile_X2Y11_W2BEGb[5] ;
 wire \Tile_X2Y11_W2BEGb[6] ;
 wire \Tile_X2Y11_W2BEGb[7] ;
 wire \Tile_X2Y11_W6BEG[0] ;
 wire \Tile_X2Y11_W6BEG[10] ;
 wire \Tile_X2Y11_W6BEG[11] ;
 wire \Tile_X2Y11_W6BEG[1] ;
 wire \Tile_X2Y11_W6BEG[2] ;
 wire \Tile_X2Y11_W6BEG[3] ;
 wire \Tile_X2Y11_W6BEG[4] ;
 wire \Tile_X2Y11_W6BEG[5] ;
 wire \Tile_X2Y11_W6BEG[6] ;
 wire \Tile_X2Y11_W6BEG[7] ;
 wire \Tile_X2Y11_W6BEG[8] ;
 wire \Tile_X2Y11_W6BEG[9] ;
 wire \Tile_X2Y11_WW4BEG[0] ;
 wire \Tile_X2Y11_WW4BEG[10] ;
 wire \Tile_X2Y11_WW4BEG[11] ;
 wire \Tile_X2Y11_WW4BEG[12] ;
 wire \Tile_X2Y11_WW4BEG[13] ;
 wire \Tile_X2Y11_WW4BEG[14] ;
 wire \Tile_X2Y11_WW4BEG[15] ;
 wire \Tile_X2Y11_WW4BEG[1] ;
 wire \Tile_X2Y11_WW4BEG[2] ;
 wire \Tile_X2Y11_WW4BEG[3] ;
 wire \Tile_X2Y11_WW4BEG[4] ;
 wire \Tile_X2Y11_WW4BEG[5] ;
 wire \Tile_X2Y11_WW4BEG[6] ;
 wire \Tile_X2Y11_WW4BEG[7] ;
 wire \Tile_X2Y11_WW4BEG[8] ;
 wire \Tile_X2Y11_WW4BEG[9] ;
 wire Tile_X2Y12_Co;
 wire \Tile_X2Y12_E1BEG[0] ;
 wire \Tile_X2Y12_E1BEG[1] ;
 wire \Tile_X2Y12_E1BEG[2] ;
 wire \Tile_X2Y12_E1BEG[3] ;
 wire \Tile_X2Y12_E2BEG[0] ;
 wire \Tile_X2Y12_E2BEG[1] ;
 wire \Tile_X2Y12_E2BEG[2] ;
 wire \Tile_X2Y12_E2BEG[3] ;
 wire \Tile_X2Y12_E2BEG[4] ;
 wire \Tile_X2Y12_E2BEG[5] ;
 wire \Tile_X2Y12_E2BEG[6] ;
 wire \Tile_X2Y12_E2BEG[7] ;
 wire \Tile_X2Y12_E2BEGb[0] ;
 wire \Tile_X2Y12_E2BEGb[1] ;
 wire \Tile_X2Y12_E2BEGb[2] ;
 wire \Tile_X2Y12_E2BEGb[3] ;
 wire \Tile_X2Y12_E2BEGb[4] ;
 wire \Tile_X2Y12_E2BEGb[5] ;
 wire \Tile_X2Y12_E2BEGb[6] ;
 wire \Tile_X2Y12_E2BEGb[7] ;
 wire \Tile_X2Y12_E6BEG[0] ;
 wire \Tile_X2Y12_E6BEG[10] ;
 wire \Tile_X2Y12_E6BEG[11] ;
 wire \Tile_X2Y12_E6BEG[1] ;
 wire \Tile_X2Y12_E6BEG[2] ;
 wire \Tile_X2Y12_E6BEG[3] ;
 wire \Tile_X2Y12_E6BEG[4] ;
 wire \Tile_X2Y12_E6BEG[5] ;
 wire \Tile_X2Y12_E6BEG[6] ;
 wire \Tile_X2Y12_E6BEG[7] ;
 wire \Tile_X2Y12_E6BEG[8] ;
 wire \Tile_X2Y12_E6BEG[9] ;
 wire \Tile_X2Y12_EE4BEG[0] ;
 wire \Tile_X2Y12_EE4BEG[10] ;
 wire \Tile_X2Y12_EE4BEG[11] ;
 wire \Tile_X2Y12_EE4BEG[12] ;
 wire \Tile_X2Y12_EE4BEG[13] ;
 wire \Tile_X2Y12_EE4BEG[14] ;
 wire \Tile_X2Y12_EE4BEG[15] ;
 wire \Tile_X2Y12_EE4BEG[1] ;
 wire \Tile_X2Y12_EE4BEG[2] ;
 wire \Tile_X2Y12_EE4BEG[3] ;
 wire \Tile_X2Y12_EE4BEG[4] ;
 wire \Tile_X2Y12_EE4BEG[5] ;
 wire \Tile_X2Y12_EE4BEG[6] ;
 wire \Tile_X2Y12_EE4BEG[7] ;
 wire \Tile_X2Y12_EE4BEG[8] ;
 wire \Tile_X2Y12_EE4BEG[9] ;
 wire \Tile_X2Y12_FrameData_O[0] ;
 wire \Tile_X2Y12_FrameData_O[10] ;
 wire \Tile_X2Y12_FrameData_O[11] ;
 wire \Tile_X2Y12_FrameData_O[12] ;
 wire \Tile_X2Y12_FrameData_O[13] ;
 wire \Tile_X2Y12_FrameData_O[14] ;
 wire \Tile_X2Y12_FrameData_O[15] ;
 wire \Tile_X2Y12_FrameData_O[16] ;
 wire \Tile_X2Y12_FrameData_O[17] ;
 wire \Tile_X2Y12_FrameData_O[18] ;
 wire \Tile_X2Y12_FrameData_O[19] ;
 wire \Tile_X2Y12_FrameData_O[1] ;
 wire \Tile_X2Y12_FrameData_O[20] ;
 wire \Tile_X2Y12_FrameData_O[21] ;
 wire \Tile_X2Y12_FrameData_O[22] ;
 wire \Tile_X2Y12_FrameData_O[23] ;
 wire \Tile_X2Y12_FrameData_O[24] ;
 wire \Tile_X2Y12_FrameData_O[25] ;
 wire \Tile_X2Y12_FrameData_O[26] ;
 wire \Tile_X2Y12_FrameData_O[27] ;
 wire \Tile_X2Y12_FrameData_O[28] ;
 wire \Tile_X2Y12_FrameData_O[29] ;
 wire \Tile_X2Y12_FrameData_O[2] ;
 wire \Tile_X2Y12_FrameData_O[30] ;
 wire \Tile_X2Y12_FrameData_O[31] ;
 wire \Tile_X2Y12_FrameData_O[3] ;
 wire \Tile_X2Y12_FrameData_O[4] ;
 wire \Tile_X2Y12_FrameData_O[5] ;
 wire \Tile_X2Y12_FrameData_O[6] ;
 wire \Tile_X2Y12_FrameData_O[7] ;
 wire \Tile_X2Y12_FrameData_O[8] ;
 wire \Tile_X2Y12_FrameData_O[9] ;
 wire \Tile_X2Y12_FrameStrobe_O[0] ;
 wire \Tile_X2Y12_FrameStrobe_O[10] ;
 wire \Tile_X2Y12_FrameStrobe_O[11] ;
 wire \Tile_X2Y12_FrameStrobe_O[12] ;
 wire \Tile_X2Y12_FrameStrobe_O[13] ;
 wire \Tile_X2Y12_FrameStrobe_O[14] ;
 wire \Tile_X2Y12_FrameStrobe_O[15] ;
 wire \Tile_X2Y12_FrameStrobe_O[16] ;
 wire \Tile_X2Y12_FrameStrobe_O[17] ;
 wire \Tile_X2Y12_FrameStrobe_O[18] ;
 wire \Tile_X2Y12_FrameStrobe_O[19] ;
 wire \Tile_X2Y12_FrameStrobe_O[1] ;
 wire \Tile_X2Y12_FrameStrobe_O[2] ;
 wire \Tile_X2Y12_FrameStrobe_O[3] ;
 wire \Tile_X2Y12_FrameStrobe_O[4] ;
 wire \Tile_X2Y12_FrameStrobe_O[5] ;
 wire \Tile_X2Y12_FrameStrobe_O[6] ;
 wire \Tile_X2Y12_FrameStrobe_O[7] ;
 wire \Tile_X2Y12_FrameStrobe_O[8] ;
 wire \Tile_X2Y12_FrameStrobe_O[9] ;
 wire \Tile_X2Y12_N1BEG[0] ;
 wire \Tile_X2Y12_N1BEG[1] ;
 wire \Tile_X2Y12_N1BEG[2] ;
 wire \Tile_X2Y12_N1BEG[3] ;
 wire \Tile_X2Y12_N2BEG[0] ;
 wire \Tile_X2Y12_N2BEG[1] ;
 wire \Tile_X2Y12_N2BEG[2] ;
 wire \Tile_X2Y12_N2BEG[3] ;
 wire \Tile_X2Y12_N2BEG[4] ;
 wire \Tile_X2Y12_N2BEG[5] ;
 wire \Tile_X2Y12_N2BEG[6] ;
 wire \Tile_X2Y12_N2BEG[7] ;
 wire \Tile_X2Y12_N2BEGb[0] ;
 wire \Tile_X2Y12_N2BEGb[1] ;
 wire \Tile_X2Y12_N2BEGb[2] ;
 wire \Tile_X2Y12_N2BEGb[3] ;
 wire \Tile_X2Y12_N2BEGb[4] ;
 wire \Tile_X2Y12_N2BEGb[5] ;
 wire \Tile_X2Y12_N2BEGb[6] ;
 wire \Tile_X2Y12_N2BEGb[7] ;
 wire \Tile_X2Y12_N4BEG[0] ;
 wire \Tile_X2Y12_N4BEG[10] ;
 wire \Tile_X2Y12_N4BEG[11] ;
 wire \Tile_X2Y12_N4BEG[12] ;
 wire \Tile_X2Y12_N4BEG[13] ;
 wire \Tile_X2Y12_N4BEG[14] ;
 wire \Tile_X2Y12_N4BEG[15] ;
 wire \Tile_X2Y12_N4BEG[1] ;
 wire \Tile_X2Y12_N4BEG[2] ;
 wire \Tile_X2Y12_N4BEG[3] ;
 wire \Tile_X2Y12_N4BEG[4] ;
 wire \Tile_X2Y12_N4BEG[5] ;
 wire \Tile_X2Y12_N4BEG[6] ;
 wire \Tile_X2Y12_N4BEG[7] ;
 wire \Tile_X2Y12_N4BEG[8] ;
 wire \Tile_X2Y12_N4BEG[9] ;
 wire \Tile_X2Y12_NN4BEG[0] ;
 wire \Tile_X2Y12_NN4BEG[10] ;
 wire \Tile_X2Y12_NN4BEG[11] ;
 wire \Tile_X2Y12_NN4BEG[12] ;
 wire \Tile_X2Y12_NN4BEG[13] ;
 wire \Tile_X2Y12_NN4BEG[14] ;
 wire \Tile_X2Y12_NN4BEG[15] ;
 wire \Tile_X2Y12_NN4BEG[1] ;
 wire \Tile_X2Y12_NN4BEG[2] ;
 wire \Tile_X2Y12_NN4BEG[3] ;
 wire \Tile_X2Y12_NN4BEG[4] ;
 wire \Tile_X2Y12_NN4BEG[5] ;
 wire \Tile_X2Y12_NN4BEG[6] ;
 wire \Tile_X2Y12_NN4BEG[7] ;
 wire \Tile_X2Y12_NN4BEG[8] ;
 wire \Tile_X2Y12_NN4BEG[9] ;
 wire \Tile_X2Y12_S1BEG[0] ;
 wire \Tile_X2Y12_S1BEG[1] ;
 wire \Tile_X2Y12_S1BEG[2] ;
 wire \Tile_X2Y12_S1BEG[3] ;
 wire \Tile_X2Y12_S2BEG[0] ;
 wire \Tile_X2Y12_S2BEG[1] ;
 wire \Tile_X2Y12_S2BEG[2] ;
 wire \Tile_X2Y12_S2BEG[3] ;
 wire \Tile_X2Y12_S2BEG[4] ;
 wire \Tile_X2Y12_S2BEG[5] ;
 wire \Tile_X2Y12_S2BEG[6] ;
 wire \Tile_X2Y12_S2BEG[7] ;
 wire \Tile_X2Y12_S2BEGb[0] ;
 wire \Tile_X2Y12_S2BEGb[1] ;
 wire \Tile_X2Y12_S2BEGb[2] ;
 wire \Tile_X2Y12_S2BEGb[3] ;
 wire \Tile_X2Y12_S2BEGb[4] ;
 wire \Tile_X2Y12_S2BEGb[5] ;
 wire \Tile_X2Y12_S2BEGb[6] ;
 wire \Tile_X2Y12_S2BEGb[7] ;
 wire \Tile_X2Y12_S4BEG[0] ;
 wire \Tile_X2Y12_S4BEG[10] ;
 wire \Tile_X2Y12_S4BEG[11] ;
 wire \Tile_X2Y12_S4BEG[12] ;
 wire \Tile_X2Y12_S4BEG[13] ;
 wire \Tile_X2Y12_S4BEG[14] ;
 wire \Tile_X2Y12_S4BEG[15] ;
 wire \Tile_X2Y12_S4BEG[1] ;
 wire \Tile_X2Y12_S4BEG[2] ;
 wire \Tile_X2Y12_S4BEG[3] ;
 wire \Tile_X2Y12_S4BEG[4] ;
 wire \Tile_X2Y12_S4BEG[5] ;
 wire \Tile_X2Y12_S4BEG[6] ;
 wire \Tile_X2Y12_S4BEG[7] ;
 wire \Tile_X2Y12_S4BEG[8] ;
 wire \Tile_X2Y12_S4BEG[9] ;
 wire \Tile_X2Y12_SS4BEG[0] ;
 wire \Tile_X2Y12_SS4BEG[10] ;
 wire \Tile_X2Y12_SS4BEG[11] ;
 wire \Tile_X2Y12_SS4BEG[12] ;
 wire \Tile_X2Y12_SS4BEG[13] ;
 wire \Tile_X2Y12_SS4BEG[14] ;
 wire \Tile_X2Y12_SS4BEG[15] ;
 wire \Tile_X2Y12_SS4BEG[1] ;
 wire \Tile_X2Y12_SS4BEG[2] ;
 wire \Tile_X2Y12_SS4BEG[3] ;
 wire \Tile_X2Y12_SS4BEG[4] ;
 wire \Tile_X2Y12_SS4BEG[5] ;
 wire \Tile_X2Y12_SS4BEG[6] ;
 wire \Tile_X2Y12_SS4BEG[7] ;
 wire \Tile_X2Y12_SS4BEG[8] ;
 wire \Tile_X2Y12_SS4BEG[9] ;
 wire Tile_X2Y12_UserCLKo;
 wire \Tile_X2Y12_W1BEG[0] ;
 wire \Tile_X2Y12_W1BEG[1] ;
 wire \Tile_X2Y12_W1BEG[2] ;
 wire \Tile_X2Y12_W1BEG[3] ;
 wire \Tile_X2Y12_W2BEG[0] ;
 wire \Tile_X2Y12_W2BEG[1] ;
 wire \Tile_X2Y12_W2BEG[2] ;
 wire \Tile_X2Y12_W2BEG[3] ;
 wire \Tile_X2Y12_W2BEG[4] ;
 wire \Tile_X2Y12_W2BEG[5] ;
 wire \Tile_X2Y12_W2BEG[6] ;
 wire \Tile_X2Y12_W2BEG[7] ;
 wire \Tile_X2Y12_W2BEGb[0] ;
 wire \Tile_X2Y12_W2BEGb[1] ;
 wire \Tile_X2Y12_W2BEGb[2] ;
 wire \Tile_X2Y12_W2BEGb[3] ;
 wire \Tile_X2Y12_W2BEGb[4] ;
 wire \Tile_X2Y12_W2BEGb[5] ;
 wire \Tile_X2Y12_W2BEGb[6] ;
 wire \Tile_X2Y12_W2BEGb[7] ;
 wire \Tile_X2Y12_W6BEG[0] ;
 wire \Tile_X2Y12_W6BEG[10] ;
 wire \Tile_X2Y12_W6BEG[11] ;
 wire \Tile_X2Y12_W6BEG[1] ;
 wire \Tile_X2Y12_W6BEG[2] ;
 wire \Tile_X2Y12_W6BEG[3] ;
 wire \Tile_X2Y12_W6BEG[4] ;
 wire \Tile_X2Y12_W6BEG[5] ;
 wire \Tile_X2Y12_W6BEG[6] ;
 wire \Tile_X2Y12_W6BEG[7] ;
 wire \Tile_X2Y12_W6BEG[8] ;
 wire \Tile_X2Y12_W6BEG[9] ;
 wire \Tile_X2Y12_WW4BEG[0] ;
 wire \Tile_X2Y12_WW4BEG[10] ;
 wire \Tile_X2Y12_WW4BEG[11] ;
 wire \Tile_X2Y12_WW4BEG[12] ;
 wire \Tile_X2Y12_WW4BEG[13] ;
 wire \Tile_X2Y12_WW4BEG[14] ;
 wire \Tile_X2Y12_WW4BEG[15] ;
 wire \Tile_X2Y12_WW4BEG[1] ;
 wire \Tile_X2Y12_WW4BEG[2] ;
 wire \Tile_X2Y12_WW4BEG[3] ;
 wire \Tile_X2Y12_WW4BEG[4] ;
 wire \Tile_X2Y12_WW4BEG[5] ;
 wire \Tile_X2Y12_WW4BEG[6] ;
 wire \Tile_X2Y12_WW4BEG[7] ;
 wire \Tile_X2Y12_WW4BEG[8] ;
 wire \Tile_X2Y12_WW4BEG[9] ;
 wire Tile_X2Y13_Co;
 wire \Tile_X2Y13_E1BEG[0] ;
 wire \Tile_X2Y13_E1BEG[1] ;
 wire \Tile_X2Y13_E1BEG[2] ;
 wire \Tile_X2Y13_E1BEG[3] ;
 wire \Tile_X2Y13_E2BEG[0] ;
 wire \Tile_X2Y13_E2BEG[1] ;
 wire \Tile_X2Y13_E2BEG[2] ;
 wire \Tile_X2Y13_E2BEG[3] ;
 wire \Tile_X2Y13_E2BEG[4] ;
 wire \Tile_X2Y13_E2BEG[5] ;
 wire \Tile_X2Y13_E2BEG[6] ;
 wire \Tile_X2Y13_E2BEG[7] ;
 wire \Tile_X2Y13_E2BEGb[0] ;
 wire \Tile_X2Y13_E2BEGb[1] ;
 wire \Tile_X2Y13_E2BEGb[2] ;
 wire \Tile_X2Y13_E2BEGb[3] ;
 wire \Tile_X2Y13_E2BEGb[4] ;
 wire \Tile_X2Y13_E2BEGb[5] ;
 wire \Tile_X2Y13_E2BEGb[6] ;
 wire \Tile_X2Y13_E2BEGb[7] ;
 wire \Tile_X2Y13_E6BEG[0] ;
 wire \Tile_X2Y13_E6BEG[10] ;
 wire \Tile_X2Y13_E6BEG[11] ;
 wire \Tile_X2Y13_E6BEG[1] ;
 wire \Tile_X2Y13_E6BEG[2] ;
 wire \Tile_X2Y13_E6BEG[3] ;
 wire \Tile_X2Y13_E6BEG[4] ;
 wire \Tile_X2Y13_E6BEG[5] ;
 wire \Tile_X2Y13_E6BEG[6] ;
 wire \Tile_X2Y13_E6BEG[7] ;
 wire \Tile_X2Y13_E6BEG[8] ;
 wire \Tile_X2Y13_E6BEG[9] ;
 wire \Tile_X2Y13_EE4BEG[0] ;
 wire \Tile_X2Y13_EE4BEG[10] ;
 wire \Tile_X2Y13_EE4BEG[11] ;
 wire \Tile_X2Y13_EE4BEG[12] ;
 wire \Tile_X2Y13_EE4BEG[13] ;
 wire \Tile_X2Y13_EE4BEG[14] ;
 wire \Tile_X2Y13_EE4BEG[15] ;
 wire \Tile_X2Y13_EE4BEG[1] ;
 wire \Tile_X2Y13_EE4BEG[2] ;
 wire \Tile_X2Y13_EE4BEG[3] ;
 wire \Tile_X2Y13_EE4BEG[4] ;
 wire \Tile_X2Y13_EE4BEG[5] ;
 wire \Tile_X2Y13_EE4BEG[6] ;
 wire \Tile_X2Y13_EE4BEG[7] ;
 wire \Tile_X2Y13_EE4BEG[8] ;
 wire \Tile_X2Y13_EE4BEG[9] ;
 wire \Tile_X2Y13_FrameData_O[0] ;
 wire \Tile_X2Y13_FrameData_O[10] ;
 wire \Tile_X2Y13_FrameData_O[11] ;
 wire \Tile_X2Y13_FrameData_O[12] ;
 wire \Tile_X2Y13_FrameData_O[13] ;
 wire \Tile_X2Y13_FrameData_O[14] ;
 wire \Tile_X2Y13_FrameData_O[15] ;
 wire \Tile_X2Y13_FrameData_O[16] ;
 wire \Tile_X2Y13_FrameData_O[17] ;
 wire \Tile_X2Y13_FrameData_O[18] ;
 wire \Tile_X2Y13_FrameData_O[19] ;
 wire \Tile_X2Y13_FrameData_O[1] ;
 wire \Tile_X2Y13_FrameData_O[20] ;
 wire \Tile_X2Y13_FrameData_O[21] ;
 wire \Tile_X2Y13_FrameData_O[22] ;
 wire \Tile_X2Y13_FrameData_O[23] ;
 wire \Tile_X2Y13_FrameData_O[24] ;
 wire \Tile_X2Y13_FrameData_O[25] ;
 wire \Tile_X2Y13_FrameData_O[26] ;
 wire \Tile_X2Y13_FrameData_O[27] ;
 wire \Tile_X2Y13_FrameData_O[28] ;
 wire \Tile_X2Y13_FrameData_O[29] ;
 wire \Tile_X2Y13_FrameData_O[2] ;
 wire \Tile_X2Y13_FrameData_O[30] ;
 wire \Tile_X2Y13_FrameData_O[31] ;
 wire \Tile_X2Y13_FrameData_O[3] ;
 wire \Tile_X2Y13_FrameData_O[4] ;
 wire \Tile_X2Y13_FrameData_O[5] ;
 wire \Tile_X2Y13_FrameData_O[6] ;
 wire \Tile_X2Y13_FrameData_O[7] ;
 wire \Tile_X2Y13_FrameData_O[8] ;
 wire \Tile_X2Y13_FrameData_O[9] ;
 wire \Tile_X2Y13_FrameStrobe_O[0] ;
 wire \Tile_X2Y13_FrameStrobe_O[10] ;
 wire \Tile_X2Y13_FrameStrobe_O[11] ;
 wire \Tile_X2Y13_FrameStrobe_O[12] ;
 wire \Tile_X2Y13_FrameStrobe_O[13] ;
 wire \Tile_X2Y13_FrameStrobe_O[14] ;
 wire \Tile_X2Y13_FrameStrobe_O[15] ;
 wire \Tile_X2Y13_FrameStrobe_O[16] ;
 wire \Tile_X2Y13_FrameStrobe_O[17] ;
 wire \Tile_X2Y13_FrameStrobe_O[18] ;
 wire \Tile_X2Y13_FrameStrobe_O[19] ;
 wire \Tile_X2Y13_FrameStrobe_O[1] ;
 wire \Tile_X2Y13_FrameStrobe_O[2] ;
 wire \Tile_X2Y13_FrameStrobe_O[3] ;
 wire \Tile_X2Y13_FrameStrobe_O[4] ;
 wire \Tile_X2Y13_FrameStrobe_O[5] ;
 wire \Tile_X2Y13_FrameStrobe_O[6] ;
 wire \Tile_X2Y13_FrameStrobe_O[7] ;
 wire \Tile_X2Y13_FrameStrobe_O[8] ;
 wire \Tile_X2Y13_FrameStrobe_O[9] ;
 wire \Tile_X2Y13_N1BEG[0] ;
 wire \Tile_X2Y13_N1BEG[1] ;
 wire \Tile_X2Y13_N1BEG[2] ;
 wire \Tile_X2Y13_N1BEG[3] ;
 wire \Tile_X2Y13_N2BEG[0] ;
 wire \Tile_X2Y13_N2BEG[1] ;
 wire \Tile_X2Y13_N2BEG[2] ;
 wire \Tile_X2Y13_N2BEG[3] ;
 wire \Tile_X2Y13_N2BEG[4] ;
 wire \Tile_X2Y13_N2BEG[5] ;
 wire \Tile_X2Y13_N2BEG[6] ;
 wire \Tile_X2Y13_N2BEG[7] ;
 wire \Tile_X2Y13_N2BEGb[0] ;
 wire \Tile_X2Y13_N2BEGb[1] ;
 wire \Tile_X2Y13_N2BEGb[2] ;
 wire \Tile_X2Y13_N2BEGb[3] ;
 wire \Tile_X2Y13_N2BEGb[4] ;
 wire \Tile_X2Y13_N2BEGb[5] ;
 wire \Tile_X2Y13_N2BEGb[6] ;
 wire \Tile_X2Y13_N2BEGb[7] ;
 wire \Tile_X2Y13_N4BEG[0] ;
 wire \Tile_X2Y13_N4BEG[10] ;
 wire \Tile_X2Y13_N4BEG[11] ;
 wire \Tile_X2Y13_N4BEG[12] ;
 wire \Tile_X2Y13_N4BEG[13] ;
 wire \Tile_X2Y13_N4BEG[14] ;
 wire \Tile_X2Y13_N4BEG[15] ;
 wire \Tile_X2Y13_N4BEG[1] ;
 wire \Tile_X2Y13_N4BEG[2] ;
 wire \Tile_X2Y13_N4BEG[3] ;
 wire \Tile_X2Y13_N4BEG[4] ;
 wire \Tile_X2Y13_N4BEG[5] ;
 wire \Tile_X2Y13_N4BEG[6] ;
 wire \Tile_X2Y13_N4BEG[7] ;
 wire \Tile_X2Y13_N4BEG[8] ;
 wire \Tile_X2Y13_N4BEG[9] ;
 wire \Tile_X2Y13_NN4BEG[0] ;
 wire \Tile_X2Y13_NN4BEG[10] ;
 wire \Tile_X2Y13_NN4BEG[11] ;
 wire \Tile_X2Y13_NN4BEG[12] ;
 wire \Tile_X2Y13_NN4BEG[13] ;
 wire \Tile_X2Y13_NN4BEG[14] ;
 wire \Tile_X2Y13_NN4BEG[15] ;
 wire \Tile_X2Y13_NN4BEG[1] ;
 wire \Tile_X2Y13_NN4BEG[2] ;
 wire \Tile_X2Y13_NN4BEG[3] ;
 wire \Tile_X2Y13_NN4BEG[4] ;
 wire \Tile_X2Y13_NN4BEG[5] ;
 wire \Tile_X2Y13_NN4BEG[6] ;
 wire \Tile_X2Y13_NN4BEG[7] ;
 wire \Tile_X2Y13_NN4BEG[8] ;
 wire \Tile_X2Y13_NN4BEG[9] ;
 wire \Tile_X2Y13_S1BEG[0] ;
 wire \Tile_X2Y13_S1BEG[1] ;
 wire \Tile_X2Y13_S1BEG[2] ;
 wire \Tile_X2Y13_S1BEG[3] ;
 wire \Tile_X2Y13_S2BEG[0] ;
 wire \Tile_X2Y13_S2BEG[1] ;
 wire \Tile_X2Y13_S2BEG[2] ;
 wire \Tile_X2Y13_S2BEG[3] ;
 wire \Tile_X2Y13_S2BEG[4] ;
 wire \Tile_X2Y13_S2BEG[5] ;
 wire \Tile_X2Y13_S2BEG[6] ;
 wire \Tile_X2Y13_S2BEG[7] ;
 wire \Tile_X2Y13_S2BEGb[0] ;
 wire \Tile_X2Y13_S2BEGb[1] ;
 wire \Tile_X2Y13_S2BEGb[2] ;
 wire \Tile_X2Y13_S2BEGb[3] ;
 wire \Tile_X2Y13_S2BEGb[4] ;
 wire \Tile_X2Y13_S2BEGb[5] ;
 wire \Tile_X2Y13_S2BEGb[6] ;
 wire \Tile_X2Y13_S2BEGb[7] ;
 wire \Tile_X2Y13_S4BEG[0] ;
 wire \Tile_X2Y13_S4BEG[10] ;
 wire \Tile_X2Y13_S4BEG[11] ;
 wire \Tile_X2Y13_S4BEG[12] ;
 wire \Tile_X2Y13_S4BEG[13] ;
 wire \Tile_X2Y13_S4BEG[14] ;
 wire \Tile_X2Y13_S4BEG[15] ;
 wire \Tile_X2Y13_S4BEG[1] ;
 wire \Tile_X2Y13_S4BEG[2] ;
 wire \Tile_X2Y13_S4BEG[3] ;
 wire \Tile_X2Y13_S4BEG[4] ;
 wire \Tile_X2Y13_S4BEG[5] ;
 wire \Tile_X2Y13_S4BEG[6] ;
 wire \Tile_X2Y13_S4BEG[7] ;
 wire \Tile_X2Y13_S4BEG[8] ;
 wire \Tile_X2Y13_S4BEG[9] ;
 wire \Tile_X2Y13_SS4BEG[0] ;
 wire \Tile_X2Y13_SS4BEG[10] ;
 wire \Tile_X2Y13_SS4BEG[11] ;
 wire \Tile_X2Y13_SS4BEG[12] ;
 wire \Tile_X2Y13_SS4BEG[13] ;
 wire \Tile_X2Y13_SS4BEG[14] ;
 wire \Tile_X2Y13_SS4BEG[15] ;
 wire \Tile_X2Y13_SS4BEG[1] ;
 wire \Tile_X2Y13_SS4BEG[2] ;
 wire \Tile_X2Y13_SS4BEG[3] ;
 wire \Tile_X2Y13_SS4BEG[4] ;
 wire \Tile_X2Y13_SS4BEG[5] ;
 wire \Tile_X2Y13_SS4BEG[6] ;
 wire \Tile_X2Y13_SS4BEG[7] ;
 wire \Tile_X2Y13_SS4BEG[8] ;
 wire \Tile_X2Y13_SS4BEG[9] ;
 wire Tile_X2Y13_UserCLKo;
 wire \Tile_X2Y13_W1BEG[0] ;
 wire \Tile_X2Y13_W1BEG[1] ;
 wire \Tile_X2Y13_W1BEG[2] ;
 wire \Tile_X2Y13_W1BEG[3] ;
 wire \Tile_X2Y13_W2BEG[0] ;
 wire \Tile_X2Y13_W2BEG[1] ;
 wire \Tile_X2Y13_W2BEG[2] ;
 wire \Tile_X2Y13_W2BEG[3] ;
 wire \Tile_X2Y13_W2BEG[4] ;
 wire \Tile_X2Y13_W2BEG[5] ;
 wire \Tile_X2Y13_W2BEG[6] ;
 wire \Tile_X2Y13_W2BEG[7] ;
 wire \Tile_X2Y13_W2BEGb[0] ;
 wire \Tile_X2Y13_W2BEGb[1] ;
 wire \Tile_X2Y13_W2BEGb[2] ;
 wire \Tile_X2Y13_W2BEGb[3] ;
 wire \Tile_X2Y13_W2BEGb[4] ;
 wire \Tile_X2Y13_W2BEGb[5] ;
 wire \Tile_X2Y13_W2BEGb[6] ;
 wire \Tile_X2Y13_W2BEGb[7] ;
 wire \Tile_X2Y13_W6BEG[0] ;
 wire \Tile_X2Y13_W6BEG[10] ;
 wire \Tile_X2Y13_W6BEG[11] ;
 wire \Tile_X2Y13_W6BEG[1] ;
 wire \Tile_X2Y13_W6BEG[2] ;
 wire \Tile_X2Y13_W6BEG[3] ;
 wire \Tile_X2Y13_W6BEG[4] ;
 wire \Tile_X2Y13_W6BEG[5] ;
 wire \Tile_X2Y13_W6BEG[6] ;
 wire \Tile_X2Y13_W6BEG[7] ;
 wire \Tile_X2Y13_W6BEG[8] ;
 wire \Tile_X2Y13_W6BEG[9] ;
 wire \Tile_X2Y13_WW4BEG[0] ;
 wire \Tile_X2Y13_WW4BEG[10] ;
 wire \Tile_X2Y13_WW4BEG[11] ;
 wire \Tile_X2Y13_WW4BEG[12] ;
 wire \Tile_X2Y13_WW4BEG[13] ;
 wire \Tile_X2Y13_WW4BEG[14] ;
 wire \Tile_X2Y13_WW4BEG[15] ;
 wire \Tile_X2Y13_WW4BEG[1] ;
 wire \Tile_X2Y13_WW4BEG[2] ;
 wire \Tile_X2Y13_WW4BEG[3] ;
 wire \Tile_X2Y13_WW4BEG[4] ;
 wire \Tile_X2Y13_WW4BEG[5] ;
 wire \Tile_X2Y13_WW4BEG[6] ;
 wire \Tile_X2Y13_WW4BEG[7] ;
 wire \Tile_X2Y13_WW4BEG[8] ;
 wire \Tile_X2Y13_WW4BEG[9] ;
 wire Tile_X2Y14_Co;
 wire \Tile_X2Y14_E1BEG[0] ;
 wire \Tile_X2Y14_E1BEG[1] ;
 wire \Tile_X2Y14_E1BEG[2] ;
 wire \Tile_X2Y14_E1BEG[3] ;
 wire \Tile_X2Y14_E2BEG[0] ;
 wire \Tile_X2Y14_E2BEG[1] ;
 wire \Tile_X2Y14_E2BEG[2] ;
 wire \Tile_X2Y14_E2BEG[3] ;
 wire \Tile_X2Y14_E2BEG[4] ;
 wire \Tile_X2Y14_E2BEG[5] ;
 wire \Tile_X2Y14_E2BEG[6] ;
 wire \Tile_X2Y14_E2BEG[7] ;
 wire \Tile_X2Y14_E2BEGb[0] ;
 wire \Tile_X2Y14_E2BEGb[1] ;
 wire \Tile_X2Y14_E2BEGb[2] ;
 wire \Tile_X2Y14_E2BEGb[3] ;
 wire \Tile_X2Y14_E2BEGb[4] ;
 wire \Tile_X2Y14_E2BEGb[5] ;
 wire \Tile_X2Y14_E2BEGb[6] ;
 wire \Tile_X2Y14_E2BEGb[7] ;
 wire \Tile_X2Y14_E6BEG[0] ;
 wire \Tile_X2Y14_E6BEG[10] ;
 wire \Tile_X2Y14_E6BEG[11] ;
 wire \Tile_X2Y14_E6BEG[1] ;
 wire \Tile_X2Y14_E6BEG[2] ;
 wire \Tile_X2Y14_E6BEG[3] ;
 wire \Tile_X2Y14_E6BEG[4] ;
 wire \Tile_X2Y14_E6BEG[5] ;
 wire \Tile_X2Y14_E6BEG[6] ;
 wire \Tile_X2Y14_E6BEG[7] ;
 wire \Tile_X2Y14_E6BEG[8] ;
 wire \Tile_X2Y14_E6BEG[9] ;
 wire \Tile_X2Y14_EE4BEG[0] ;
 wire \Tile_X2Y14_EE4BEG[10] ;
 wire \Tile_X2Y14_EE4BEG[11] ;
 wire \Tile_X2Y14_EE4BEG[12] ;
 wire \Tile_X2Y14_EE4BEG[13] ;
 wire \Tile_X2Y14_EE4BEG[14] ;
 wire \Tile_X2Y14_EE4BEG[15] ;
 wire \Tile_X2Y14_EE4BEG[1] ;
 wire \Tile_X2Y14_EE4BEG[2] ;
 wire \Tile_X2Y14_EE4BEG[3] ;
 wire \Tile_X2Y14_EE4BEG[4] ;
 wire \Tile_X2Y14_EE4BEG[5] ;
 wire \Tile_X2Y14_EE4BEG[6] ;
 wire \Tile_X2Y14_EE4BEG[7] ;
 wire \Tile_X2Y14_EE4BEG[8] ;
 wire \Tile_X2Y14_EE4BEG[9] ;
 wire \Tile_X2Y14_FrameData_O[0] ;
 wire \Tile_X2Y14_FrameData_O[10] ;
 wire \Tile_X2Y14_FrameData_O[11] ;
 wire \Tile_X2Y14_FrameData_O[12] ;
 wire \Tile_X2Y14_FrameData_O[13] ;
 wire \Tile_X2Y14_FrameData_O[14] ;
 wire \Tile_X2Y14_FrameData_O[15] ;
 wire \Tile_X2Y14_FrameData_O[16] ;
 wire \Tile_X2Y14_FrameData_O[17] ;
 wire \Tile_X2Y14_FrameData_O[18] ;
 wire \Tile_X2Y14_FrameData_O[19] ;
 wire \Tile_X2Y14_FrameData_O[1] ;
 wire \Tile_X2Y14_FrameData_O[20] ;
 wire \Tile_X2Y14_FrameData_O[21] ;
 wire \Tile_X2Y14_FrameData_O[22] ;
 wire \Tile_X2Y14_FrameData_O[23] ;
 wire \Tile_X2Y14_FrameData_O[24] ;
 wire \Tile_X2Y14_FrameData_O[25] ;
 wire \Tile_X2Y14_FrameData_O[26] ;
 wire \Tile_X2Y14_FrameData_O[27] ;
 wire \Tile_X2Y14_FrameData_O[28] ;
 wire \Tile_X2Y14_FrameData_O[29] ;
 wire \Tile_X2Y14_FrameData_O[2] ;
 wire \Tile_X2Y14_FrameData_O[30] ;
 wire \Tile_X2Y14_FrameData_O[31] ;
 wire \Tile_X2Y14_FrameData_O[3] ;
 wire \Tile_X2Y14_FrameData_O[4] ;
 wire \Tile_X2Y14_FrameData_O[5] ;
 wire \Tile_X2Y14_FrameData_O[6] ;
 wire \Tile_X2Y14_FrameData_O[7] ;
 wire \Tile_X2Y14_FrameData_O[8] ;
 wire \Tile_X2Y14_FrameData_O[9] ;
 wire \Tile_X2Y14_FrameStrobe_O[0] ;
 wire \Tile_X2Y14_FrameStrobe_O[10] ;
 wire \Tile_X2Y14_FrameStrobe_O[11] ;
 wire \Tile_X2Y14_FrameStrobe_O[12] ;
 wire \Tile_X2Y14_FrameStrobe_O[13] ;
 wire \Tile_X2Y14_FrameStrobe_O[14] ;
 wire \Tile_X2Y14_FrameStrobe_O[15] ;
 wire \Tile_X2Y14_FrameStrobe_O[16] ;
 wire \Tile_X2Y14_FrameStrobe_O[17] ;
 wire \Tile_X2Y14_FrameStrobe_O[18] ;
 wire \Tile_X2Y14_FrameStrobe_O[19] ;
 wire \Tile_X2Y14_FrameStrobe_O[1] ;
 wire \Tile_X2Y14_FrameStrobe_O[2] ;
 wire \Tile_X2Y14_FrameStrobe_O[3] ;
 wire \Tile_X2Y14_FrameStrobe_O[4] ;
 wire \Tile_X2Y14_FrameStrobe_O[5] ;
 wire \Tile_X2Y14_FrameStrobe_O[6] ;
 wire \Tile_X2Y14_FrameStrobe_O[7] ;
 wire \Tile_X2Y14_FrameStrobe_O[8] ;
 wire \Tile_X2Y14_FrameStrobe_O[9] ;
 wire \Tile_X2Y14_N1BEG[0] ;
 wire \Tile_X2Y14_N1BEG[1] ;
 wire \Tile_X2Y14_N1BEG[2] ;
 wire \Tile_X2Y14_N1BEG[3] ;
 wire \Tile_X2Y14_N2BEG[0] ;
 wire \Tile_X2Y14_N2BEG[1] ;
 wire \Tile_X2Y14_N2BEG[2] ;
 wire \Tile_X2Y14_N2BEG[3] ;
 wire \Tile_X2Y14_N2BEG[4] ;
 wire \Tile_X2Y14_N2BEG[5] ;
 wire \Tile_X2Y14_N2BEG[6] ;
 wire \Tile_X2Y14_N2BEG[7] ;
 wire \Tile_X2Y14_N2BEGb[0] ;
 wire \Tile_X2Y14_N2BEGb[1] ;
 wire \Tile_X2Y14_N2BEGb[2] ;
 wire \Tile_X2Y14_N2BEGb[3] ;
 wire \Tile_X2Y14_N2BEGb[4] ;
 wire \Tile_X2Y14_N2BEGb[5] ;
 wire \Tile_X2Y14_N2BEGb[6] ;
 wire \Tile_X2Y14_N2BEGb[7] ;
 wire \Tile_X2Y14_N4BEG[0] ;
 wire \Tile_X2Y14_N4BEG[10] ;
 wire \Tile_X2Y14_N4BEG[11] ;
 wire \Tile_X2Y14_N4BEG[12] ;
 wire \Tile_X2Y14_N4BEG[13] ;
 wire \Tile_X2Y14_N4BEG[14] ;
 wire \Tile_X2Y14_N4BEG[15] ;
 wire \Tile_X2Y14_N4BEG[1] ;
 wire \Tile_X2Y14_N4BEG[2] ;
 wire \Tile_X2Y14_N4BEG[3] ;
 wire \Tile_X2Y14_N4BEG[4] ;
 wire \Tile_X2Y14_N4BEG[5] ;
 wire \Tile_X2Y14_N4BEG[6] ;
 wire \Tile_X2Y14_N4BEG[7] ;
 wire \Tile_X2Y14_N4BEG[8] ;
 wire \Tile_X2Y14_N4BEG[9] ;
 wire \Tile_X2Y14_NN4BEG[0] ;
 wire \Tile_X2Y14_NN4BEG[10] ;
 wire \Tile_X2Y14_NN4BEG[11] ;
 wire \Tile_X2Y14_NN4BEG[12] ;
 wire \Tile_X2Y14_NN4BEG[13] ;
 wire \Tile_X2Y14_NN4BEG[14] ;
 wire \Tile_X2Y14_NN4BEG[15] ;
 wire \Tile_X2Y14_NN4BEG[1] ;
 wire \Tile_X2Y14_NN4BEG[2] ;
 wire \Tile_X2Y14_NN4BEG[3] ;
 wire \Tile_X2Y14_NN4BEG[4] ;
 wire \Tile_X2Y14_NN4BEG[5] ;
 wire \Tile_X2Y14_NN4BEG[6] ;
 wire \Tile_X2Y14_NN4BEG[7] ;
 wire \Tile_X2Y14_NN4BEG[8] ;
 wire \Tile_X2Y14_NN4BEG[9] ;
 wire \Tile_X2Y14_S1BEG[0] ;
 wire \Tile_X2Y14_S1BEG[1] ;
 wire \Tile_X2Y14_S1BEG[2] ;
 wire \Tile_X2Y14_S1BEG[3] ;
 wire \Tile_X2Y14_S2BEG[0] ;
 wire \Tile_X2Y14_S2BEG[1] ;
 wire \Tile_X2Y14_S2BEG[2] ;
 wire \Tile_X2Y14_S2BEG[3] ;
 wire \Tile_X2Y14_S2BEG[4] ;
 wire \Tile_X2Y14_S2BEG[5] ;
 wire \Tile_X2Y14_S2BEG[6] ;
 wire \Tile_X2Y14_S2BEG[7] ;
 wire \Tile_X2Y14_S2BEGb[0] ;
 wire \Tile_X2Y14_S2BEGb[1] ;
 wire \Tile_X2Y14_S2BEGb[2] ;
 wire \Tile_X2Y14_S2BEGb[3] ;
 wire \Tile_X2Y14_S2BEGb[4] ;
 wire \Tile_X2Y14_S2BEGb[5] ;
 wire \Tile_X2Y14_S2BEGb[6] ;
 wire \Tile_X2Y14_S2BEGb[7] ;
 wire \Tile_X2Y14_S4BEG[0] ;
 wire \Tile_X2Y14_S4BEG[10] ;
 wire \Tile_X2Y14_S4BEG[11] ;
 wire \Tile_X2Y14_S4BEG[12] ;
 wire \Tile_X2Y14_S4BEG[13] ;
 wire \Tile_X2Y14_S4BEG[14] ;
 wire \Tile_X2Y14_S4BEG[15] ;
 wire \Tile_X2Y14_S4BEG[1] ;
 wire \Tile_X2Y14_S4BEG[2] ;
 wire \Tile_X2Y14_S4BEG[3] ;
 wire \Tile_X2Y14_S4BEG[4] ;
 wire \Tile_X2Y14_S4BEG[5] ;
 wire \Tile_X2Y14_S4BEG[6] ;
 wire \Tile_X2Y14_S4BEG[7] ;
 wire \Tile_X2Y14_S4BEG[8] ;
 wire \Tile_X2Y14_S4BEG[9] ;
 wire \Tile_X2Y14_SS4BEG[0] ;
 wire \Tile_X2Y14_SS4BEG[10] ;
 wire \Tile_X2Y14_SS4BEG[11] ;
 wire \Tile_X2Y14_SS4BEG[12] ;
 wire \Tile_X2Y14_SS4BEG[13] ;
 wire \Tile_X2Y14_SS4BEG[14] ;
 wire \Tile_X2Y14_SS4BEG[15] ;
 wire \Tile_X2Y14_SS4BEG[1] ;
 wire \Tile_X2Y14_SS4BEG[2] ;
 wire \Tile_X2Y14_SS4BEG[3] ;
 wire \Tile_X2Y14_SS4BEG[4] ;
 wire \Tile_X2Y14_SS4BEG[5] ;
 wire \Tile_X2Y14_SS4BEG[6] ;
 wire \Tile_X2Y14_SS4BEG[7] ;
 wire \Tile_X2Y14_SS4BEG[8] ;
 wire \Tile_X2Y14_SS4BEG[9] ;
 wire Tile_X2Y14_UserCLKo;
 wire \Tile_X2Y14_W1BEG[0] ;
 wire \Tile_X2Y14_W1BEG[1] ;
 wire \Tile_X2Y14_W1BEG[2] ;
 wire \Tile_X2Y14_W1BEG[3] ;
 wire \Tile_X2Y14_W2BEG[0] ;
 wire \Tile_X2Y14_W2BEG[1] ;
 wire \Tile_X2Y14_W2BEG[2] ;
 wire \Tile_X2Y14_W2BEG[3] ;
 wire \Tile_X2Y14_W2BEG[4] ;
 wire \Tile_X2Y14_W2BEG[5] ;
 wire \Tile_X2Y14_W2BEG[6] ;
 wire \Tile_X2Y14_W2BEG[7] ;
 wire \Tile_X2Y14_W2BEGb[0] ;
 wire \Tile_X2Y14_W2BEGb[1] ;
 wire \Tile_X2Y14_W2BEGb[2] ;
 wire \Tile_X2Y14_W2BEGb[3] ;
 wire \Tile_X2Y14_W2BEGb[4] ;
 wire \Tile_X2Y14_W2BEGb[5] ;
 wire \Tile_X2Y14_W2BEGb[6] ;
 wire \Tile_X2Y14_W2BEGb[7] ;
 wire \Tile_X2Y14_W6BEG[0] ;
 wire \Tile_X2Y14_W6BEG[10] ;
 wire \Tile_X2Y14_W6BEG[11] ;
 wire \Tile_X2Y14_W6BEG[1] ;
 wire \Tile_X2Y14_W6BEG[2] ;
 wire \Tile_X2Y14_W6BEG[3] ;
 wire \Tile_X2Y14_W6BEG[4] ;
 wire \Tile_X2Y14_W6BEG[5] ;
 wire \Tile_X2Y14_W6BEG[6] ;
 wire \Tile_X2Y14_W6BEG[7] ;
 wire \Tile_X2Y14_W6BEG[8] ;
 wire \Tile_X2Y14_W6BEG[9] ;
 wire \Tile_X2Y14_WW4BEG[0] ;
 wire \Tile_X2Y14_WW4BEG[10] ;
 wire \Tile_X2Y14_WW4BEG[11] ;
 wire \Tile_X2Y14_WW4BEG[12] ;
 wire \Tile_X2Y14_WW4BEG[13] ;
 wire \Tile_X2Y14_WW4BEG[14] ;
 wire \Tile_X2Y14_WW4BEG[15] ;
 wire \Tile_X2Y14_WW4BEG[1] ;
 wire \Tile_X2Y14_WW4BEG[2] ;
 wire \Tile_X2Y14_WW4BEG[3] ;
 wire \Tile_X2Y14_WW4BEG[4] ;
 wire \Tile_X2Y14_WW4BEG[5] ;
 wire \Tile_X2Y14_WW4BEG[6] ;
 wire \Tile_X2Y14_WW4BEG[7] ;
 wire \Tile_X2Y14_WW4BEG[8] ;
 wire \Tile_X2Y14_WW4BEG[9] ;
 wire Tile_X2Y15_Co;
 wire \Tile_X2Y15_FrameData_O[0] ;
 wire \Tile_X2Y15_FrameData_O[10] ;
 wire \Tile_X2Y15_FrameData_O[11] ;
 wire \Tile_X2Y15_FrameData_O[12] ;
 wire \Tile_X2Y15_FrameData_O[13] ;
 wire \Tile_X2Y15_FrameData_O[14] ;
 wire \Tile_X2Y15_FrameData_O[15] ;
 wire \Tile_X2Y15_FrameData_O[16] ;
 wire \Tile_X2Y15_FrameData_O[17] ;
 wire \Tile_X2Y15_FrameData_O[18] ;
 wire \Tile_X2Y15_FrameData_O[19] ;
 wire \Tile_X2Y15_FrameData_O[1] ;
 wire \Tile_X2Y15_FrameData_O[20] ;
 wire \Tile_X2Y15_FrameData_O[21] ;
 wire \Tile_X2Y15_FrameData_O[22] ;
 wire \Tile_X2Y15_FrameData_O[23] ;
 wire \Tile_X2Y15_FrameData_O[24] ;
 wire \Tile_X2Y15_FrameData_O[25] ;
 wire \Tile_X2Y15_FrameData_O[26] ;
 wire \Tile_X2Y15_FrameData_O[27] ;
 wire \Tile_X2Y15_FrameData_O[28] ;
 wire \Tile_X2Y15_FrameData_O[29] ;
 wire \Tile_X2Y15_FrameData_O[2] ;
 wire \Tile_X2Y15_FrameData_O[30] ;
 wire \Tile_X2Y15_FrameData_O[31] ;
 wire \Tile_X2Y15_FrameData_O[3] ;
 wire \Tile_X2Y15_FrameData_O[4] ;
 wire \Tile_X2Y15_FrameData_O[5] ;
 wire \Tile_X2Y15_FrameData_O[6] ;
 wire \Tile_X2Y15_FrameData_O[7] ;
 wire \Tile_X2Y15_FrameData_O[8] ;
 wire \Tile_X2Y15_FrameData_O[9] ;
 wire \Tile_X2Y15_FrameStrobe_O[0] ;
 wire \Tile_X2Y15_FrameStrobe_O[10] ;
 wire \Tile_X2Y15_FrameStrobe_O[11] ;
 wire \Tile_X2Y15_FrameStrobe_O[12] ;
 wire \Tile_X2Y15_FrameStrobe_O[13] ;
 wire \Tile_X2Y15_FrameStrobe_O[14] ;
 wire \Tile_X2Y15_FrameStrobe_O[15] ;
 wire \Tile_X2Y15_FrameStrobe_O[16] ;
 wire \Tile_X2Y15_FrameStrobe_O[17] ;
 wire \Tile_X2Y15_FrameStrobe_O[18] ;
 wire \Tile_X2Y15_FrameStrobe_O[19] ;
 wire \Tile_X2Y15_FrameStrobe_O[1] ;
 wire \Tile_X2Y15_FrameStrobe_O[2] ;
 wire \Tile_X2Y15_FrameStrobe_O[3] ;
 wire \Tile_X2Y15_FrameStrobe_O[4] ;
 wire \Tile_X2Y15_FrameStrobe_O[5] ;
 wire \Tile_X2Y15_FrameStrobe_O[6] ;
 wire \Tile_X2Y15_FrameStrobe_O[7] ;
 wire \Tile_X2Y15_FrameStrobe_O[8] ;
 wire \Tile_X2Y15_FrameStrobe_O[9] ;
 wire \Tile_X2Y15_N1BEG[0] ;
 wire \Tile_X2Y15_N1BEG[1] ;
 wire \Tile_X2Y15_N1BEG[2] ;
 wire \Tile_X2Y15_N1BEG[3] ;
 wire \Tile_X2Y15_N2BEG[0] ;
 wire \Tile_X2Y15_N2BEG[1] ;
 wire \Tile_X2Y15_N2BEG[2] ;
 wire \Tile_X2Y15_N2BEG[3] ;
 wire \Tile_X2Y15_N2BEG[4] ;
 wire \Tile_X2Y15_N2BEG[5] ;
 wire \Tile_X2Y15_N2BEG[6] ;
 wire \Tile_X2Y15_N2BEG[7] ;
 wire \Tile_X2Y15_N2BEGb[0] ;
 wire \Tile_X2Y15_N2BEGb[1] ;
 wire \Tile_X2Y15_N2BEGb[2] ;
 wire \Tile_X2Y15_N2BEGb[3] ;
 wire \Tile_X2Y15_N2BEGb[4] ;
 wire \Tile_X2Y15_N2BEGb[5] ;
 wire \Tile_X2Y15_N2BEGb[6] ;
 wire \Tile_X2Y15_N2BEGb[7] ;
 wire \Tile_X2Y15_N4BEG[0] ;
 wire \Tile_X2Y15_N4BEG[10] ;
 wire \Tile_X2Y15_N4BEG[11] ;
 wire \Tile_X2Y15_N4BEG[12] ;
 wire \Tile_X2Y15_N4BEG[13] ;
 wire \Tile_X2Y15_N4BEG[14] ;
 wire \Tile_X2Y15_N4BEG[15] ;
 wire \Tile_X2Y15_N4BEG[1] ;
 wire \Tile_X2Y15_N4BEG[2] ;
 wire \Tile_X2Y15_N4BEG[3] ;
 wire \Tile_X2Y15_N4BEG[4] ;
 wire \Tile_X2Y15_N4BEG[5] ;
 wire \Tile_X2Y15_N4BEG[6] ;
 wire \Tile_X2Y15_N4BEG[7] ;
 wire \Tile_X2Y15_N4BEG[8] ;
 wire \Tile_X2Y15_N4BEG[9] ;
 wire \Tile_X2Y15_NN4BEG[0] ;
 wire \Tile_X2Y15_NN4BEG[10] ;
 wire \Tile_X2Y15_NN4BEG[11] ;
 wire \Tile_X2Y15_NN4BEG[12] ;
 wire \Tile_X2Y15_NN4BEG[13] ;
 wire \Tile_X2Y15_NN4BEG[14] ;
 wire \Tile_X2Y15_NN4BEG[15] ;
 wire \Tile_X2Y15_NN4BEG[1] ;
 wire \Tile_X2Y15_NN4BEG[2] ;
 wire \Tile_X2Y15_NN4BEG[3] ;
 wire \Tile_X2Y15_NN4BEG[4] ;
 wire \Tile_X2Y15_NN4BEG[5] ;
 wire \Tile_X2Y15_NN4BEG[6] ;
 wire \Tile_X2Y15_NN4BEG[7] ;
 wire \Tile_X2Y15_NN4BEG[8] ;
 wire \Tile_X2Y15_NN4BEG[9] ;
 wire Tile_X2Y15_UserCLKo;
 wire Tile_X2Y1_Co;
 wire \Tile_X2Y1_E1BEG[0] ;
 wire \Tile_X2Y1_E1BEG[1] ;
 wire \Tile_X2Y1_E1BEG[2] ;
 wire \Tile_X2Y1_E1BEG[3] ;
 wire \Tile_X2Y1_E2BEG[0] ;
 wire \Tile_X2Y1_E2BEG[1] ;
 wire \Tile_X2Y1_E2BEG[2] ;
 wire \Tile_X2Y1_E2BEG[3] ;
 wire \Tile_X2Y1_E2BEG[4] ;
 wire \Tile_X2Y1_E2BEG[5] ;
 wire \Tile_X2Y1_E2BEG[6] ;
 wire \Tile_X2Y1_E2BEG[7] ;
 wire \Tile_X2Y1_E2BEGb[0] ;
 wire \Tile_X2Y1_E2BEGb[1] ;
 wire \Tile_X2Y1_E2BEGb[2] ;
 wire \Tile_X2Y1_E2BEGb[3] ;
 wire \Tile_X2Y1_E2BEGb[4] ;
 wire \Tile_X2Y1_E2BEGb[5] ;
 wire \Tile_X2Y1_E2BEGb[6] ;
 wire \Tile_X2Y1_E2BEGb[7] ;
 wire \Tile_X2Y1_E6BEG[0] ;
 wire \Tile_X2Y1_E6BEG[10] ;
 wire \Tile_X2Y1_E6BEG[11] ;
 wire \Tile_X2Y1_E6BEG[1] ;
 wire \Tile_X2Y1_E6BEG[2] ;
 wire \Tile_X2Y1_E6BEG[3] ;
 wire \Tile_X2Y1_E6BEG[4] ;
 wire \Tile_X2Y1_E6BEG[5] ;
 wire \Tile_X2Y1_E6BEG[6] ;
 wire \Tile_X2Y1_E6BEG[7] ;
 wire \Tile_X2Y1_E6BEG[8] ;
 wire \Tile_X2Y1_E6BEG[9] ;
 wire \Tile_X2Y1_EE4BEG[0] ;
 wire \Tile_X2Y1_EE4BEG[10] ;
 wire \Tile_X2Y1_EE4BEG[11] ;
 wire \Tile_X2Y1_EE4BEG[12] ;
 wire \Tile_X2Y1_EE4BEG[13] ;
 wire \Tile_X2Y1_EE4BEG[14] ;
 wire \Tile_X2Y1_EE4BEG[15] ;
 wire \Tile_X2Y1_EE4BEG[1] ;
 wire \Tile_X2Y1_EE4BEG[2] ;
 wire \Tile_X2Y1_EE4BEG[3] ;
 wire \Tile_X2Y1_EE4BEG[4] ;
 wire \Tile_X2Y1_EE4BEG[5] ;
 wire \Tile_X2Y1_EE4BEG[6] ;
 wire \Tile_X2Y1_EE4BEG[7] ;
 wire \Tile_X2Y1_EE4BEG[8] ;
 wire \Tile_X2Y1_EE4BEG[9] ;
 wire \Tile_X2Y1_FrameData_O[0] ;
 wire \Tile_X2Y1_FrameData_O[10] ;
 wire \Tile_X2Y1_FrameData_O[11] ;
 wire \Tile_X2Y1_FrameData_O[12] ;
 wire \Tile_X2Y1_FrameData_O[13] ;
 wire \Tile_X2Y1_FrameData_O[14] ;
 wire \Tile_X2Y1_FrameData_O[15] ;
 wire \Tile_X2Y1_FrameData_O[16] ;
 wire \Tile_X2Y1_FrameData_O[17] ;
 wire \Tile_X2Y1_FrameData_O[18] ;
 wire \Tile_X2Y1_FrameData_O[19] ;
 wire \Tile_X2Y1_FrameData_O[1] ;
 wire \Tile_X2Y1_FrameData_O[20] ;
 wire \Tile_X2Y1_FrameData_O[21] ;
 wire \Tile_X2Y1_FrameData_O[22] ;
 wire \Tile_X2Y1_FrameData_O[23] ;
 wire \Tile_X2Y1_FrameData_O[24] ;
 wire \Tile_X2Y1_FrameData_O[25] ;
 wire \Tile_X2Y1_FrameData_O[26] ;
 wire \Tile_X2Y1_FrameData_O[27] ;
 wire \Tile_X2Y1_FrameData_O[28] ;
 wire \Tile_X2Y1_FrameData_O[29] ;
 wire \Tile_X2Y1_FrameData_O[2] ;
 wire \Tile_X2Y1_FrameData_O[30] ;
 wire \Tile_X2Y1_FrameData_O[31] ;
 wire \Tile_X2Y1_FrameData_O[3] ;
 wire \Tile_X2Y1_FrameData_O[4] ;
 wire \Tile_X2Y1_FrameData_O[5] ;
 wire \Tile_X2Y1_FrameData_O[6] ;
 wire \Tile_X2Y1_FrameData_O[7] ;
 wire \Tile_X2Y1_FrameData_O[8] ;
 wire \Tile_X2Y1_FrameData_O[9] ;
 wire \Tile_X2Y1_FrameStrobe_O[0] ;
 wire \Tile_X2Y1_FrameStrobe_O[10] ;
 wire \Tile_X2Y1_FrameStrobe_O[11] ;
 wire \Tile_X2Y1_FrameStrobe_O[12] ;
 wire \Tile_X2Y1_FrameStrobe_O[13] ;
 wire \Tile_X2Y1_FrameStrobe_O[14] ;
 wire \Tile_X2Y1_FrameStrobe_O[15] ;
 wire \Tile_X2Y1_FrameStrobe_O[16] ;
 wire \Tile_X2Y1_FrameStrobe_O[17] ;
 wire \Tile_X2Y1_FrameStrobe_O[18] ;
 wire \Tile_X2Y1_FrameStrobe_O[19] ;
 wire \Tile_X2Y1_FrameStrobe_O[1] ;
 wire \Tile_X2Y1_FrameStrobe_O[2] ;
 wire \Tile_X2Y1_FrameStrobe_O[3] ;
 wire \Tile_X2Y1_FrameStrobe_O[4] ;
 wire \Tile_X2Y1_FrameStrobe_O[5] ;
 wire \Tile_X2Y1_FrameStrobe_O[6] ;
 wire \Tile_X2Y1_FrameStrobe_O[7] ;
 wire \Tile_X2Y1_FrameStrobe_O[8] ;
 wire \Tile_X2Y1_FrameStrobe_O[9] ;
 wire \Tile_X2Y1_N1BEG[0] ;
 wire \Tile_X2Y1_N1BEG[1] ;
 wire \Tile_X2Y1_N1BEG[2] ;
 wire \Tile_X2Y1_N1BEG[3] ;
 wire \Tile_X2Y1_N2BEG[0] ;
 wire \Tile_X2Y1_N2BEG[1] ;
 wire \Tile_X2Y1_N2BEG[2] ;
 wire \Tile_X2Y1_N2BEG[3] ;
 wire \Tile_X2Y1_N2BEG[4] ;
 wire \Tile_X2Y1_N2BEG[5] ;
 wire \Tile_X2Y1_N2BEG[6] ;
 wire \Tile_X2Y1_N2BEG[7] ;
 wire \Tile_X2Y1_N2BEGb[0] ;
 wire \Tile_X2Y1_N2BEGb[1] ;
 wire \Tile_X2Y1_N2BEGb[2] ;
 wire \Tile_X2Y1_N2BEGb[3] ;
 wire \Tile_X2Y1_N2BEGb[4] ;
 wire \Tile_X2Y1_N2BEGb[5] ;
 wire \Tile_X2Y1_N2BEGb[6] ;
 wire \Tile_X2Y1_N2BEGb[7] ;
 wire \Tile_X2Y1_N4BEG[0] ;
 wire \Tile_X2Y1_N4BEG[10] ;
 wire \Tile_X2Y1_N4BEG[11] ;
 wire \Tile_X2Y1_N4BEG[12] ;
 wire \Tile_X2Y1_N4BEG[13] ;
 wire \Tile_X2Y1_N4BEG[14] ;
 wire \Tile_X2Y1_N4BEG[15] ;
 wire \Tile_X2Y1_N4BEG[1] ;
 wire \Tile_X2Y1_N4BEG[2] ;
 wire \Tile_X2Y1_N4BEG[3] ;
 wire \Tile_X2Y1_N4BEG[4] ;
 wire \Tile_X2Y1_N4BEG[5] ;
 wire \Tile_X2Y1_N4BEG[6] ;
 wire \Tile_X2Y1_N4BEG[7] ;
 wire \Tile_X2Y1_N4BEG[8] ;
 wire \Tile_X2Y1_N4BEG[9] ;
 wire \Tile_X2Y1_NN4BEG[0] ;
 wire \Tile_X2Y1_NN4BEG[10] ;
 wire \Tile_X2Y1_NN4BEG[11] ;
 wire \Tile_X2Y1_NN4BEG[12] ;
 wire \Tile_X2Y1_NN4BEG[13] ;
 wire \Tile_X2Y1_NN4BEG[14] ;
 wire \Tile_X2Y1_NN4BEG[15] ;
 wire \Tile_X2Y1_NN4BEG[1] ;
 wire \Tile_X2Y1_NN4BEG[2] ;
 wire \Tile_X2Y1_NN4BEG[3] ;
 wire \Tile_X2Y1_NN4BEG[4] ;
 wire \Tile_X2Y1_NN4BEG[5] ;
 wire \Tile_X2Y1_NN4BEG[6] ;
 wire \Tile_X2Y1_NN4BEG[7] ;
 wire \Tile_X2Y1_NN4BEG[8] ;
 wire \Tile_X2Y1_NN4BEG[9] ;
 wire \Tile_X2Y1_S1BEG[0] ;
 wire \Tile_X2Y1_S1BEG[1] ;
 wire \Tile_X2Y1_S1BEG[2] ;
 wire \Tile_X2Y1_S1BEG[3] ;
 wire \Tile_X2Y1_S2BEG[0] ;
 wire \Tile_X2Y1_S2BEG[1] ;
 wire \Tile_X2Y1_S2BEG[2] ;
 wire \Tile_X2Y1_S2BEG[3] ;
 wire \Tile_X2Y1_S2BEG[4] ;
 wire \Tile_X2Y1_S2BEG[5] ;
 wire \Tile_X2Y1_S2BEG[6] ;
 wire \Tile_X2Y1_S2BEG[7] ;
 wire \Tile_X2Y1_S2BEGb[0] ;
 wire \Tile_X2Y1_S2BEGb[1] ;
 wire \Tile_X2Y1_S2BEGb[2] ;
 wire \Tile_X2Y1_S2BEGb[3] ;
 wire \Tile_X2Y1_S2BEGb[4] ;
 wire \Tile_X2Y1_S2BEGb[5] ;
 wire \Tile_X2Y1_S2BEGb[6] ;
 wire \Tile_X2Y1_S2BEGb[7] ;
 wire \Tile_X2Y1_S4BEG[0] ;
 wire \Tile_X2Y1_S4BEG[10] ;
 wire \Tile_X2Y1_S4BEG[11] ;
 wire \Tile_X2Y1_S4BEG[12] ;
 wire \Tile_X2Y1_S4BEG[13] ;
 wire \Tile_X2Y1_S4BEG[14] ;
 wire \Tile_X2Y1_S4BEG[15] ;
 wire \Tile_X2Y1_S4BEG[1] ;
 wire \Tile_X2Y1_S4BEG[2] ;
 wire \Tile_X2Y1_S4BEG[3] ;
 wire \Tile_X2Y1_S4BEG[4] ;
 wire \Tile_X2Y1_S4BEG[5] ;
 wire \Tile_X2Y1_S4BEG[6] ;
 wire \Tile_X2Y1_S4BEG[7] ;
 wire \Tile_X2Y1_S4BEG[8] ;
 wire \Tile_X2Y1_S4BEG[9] ;
 wire \Tile_X2Y1_SS4BEG[0] ;
 wire \Tile_X2Y1_SS4BEG[10] ;
 wire \Tile_X2Y1_SS4BEG[11] ;
 wire \Tile_X2Y1_SS4BEG[12] ;
 wire \Tile_X2Y1_SS4BEG[13] ;
 wire \Tile_X2Y1_SS4BEG[14] ;
 wire \Tile_X2Y1_SS4BEG[15] ;
 wire \Tile_X2Y1_SS4BEG[1] ;
 wire \Tile_X2Y1_SS4BEG[2] ;
 wire \Tile_X2Y1_SS4BEG[3] ;
 wire \Tile_X2Y1_SS4BEG[4] ;
 wire \Tile_X2Y1_SS4BEG[5] ;
 wire \Tile_X2Y1_SS4BEG[6] ;
 wire \Tile_X2Y1_SS4BEG[7] ;
 wire \Tile_X2Y1_SS4BEG[8] ;
 wire \Tile_X2Y1_SS4BEG[9] ;
 wire Tile_X2Y1_UserCLKo;
 wire \Tile_X2Y1_W1BEG[0] ;
 wire \Tile_X2Y1_W1BEG[1] ;
 wire \Tile_X2Y1_W1BEG[2] ;
 wire \Tile_X2Y1_W1BEG[3] ;
 wire \Tile_X2Y1_W2BEG[0] ;
 wire \Tile_X2Y1_W2BEG[1] ;
 wire \Tile_X2Y1_W2BEG[2] ;
 wire \Tile_X2Y1_W2BEG[3] ;
 wire \Tile_X2Y1_W2BEG[4] ;
 wire \Tile_X2Y1_W2BEG[5] ;
 wire \Tile_X2Y1_W2BEG[6] ;
 wire \Tile_X2Y1_W2BEG[7] ;
 wire \Tile_X2Y1_W2BEGb[0] ;
 wire \Tile_X2Y1_W2BEGb[1] ;
 wire \Tile_X2Y1_W2BEGb[2] ;
 wire \Tile_X2Y1_W2BEGb[3] ;
 wire \Tile_X2Y1_W2BEGb[4] ;
 wire \Tile_X2Y1_W2BEGb[5] ;
 wire \Tile_X2Y1_W2BEGb[6] ;
 wire \Tile_X2Y1_W2BEGb[7] ;
 wire \Tile_X2Y1_W6BEG[0] ;
 wire \Tile_X2Y1_W6BEG[10] ;
 wire \Tile_X2Y1_W6BEG[11] ;
 wire \Tile_X2Y1_W6BEG[1] ;
 wire \Tile_X2Y1_W6BEG[2] ;
 wire \Tile_X2Y1_W6BEG[3] ;
 wire \Tile_X2Y1_W6BEG[4] ;
 wire \Tile_X2Y1_W6BEG[5] ;
 wire \Tile_X2Y1_W6BEG[6] ;
 wire \Tile_X2Y1_W6BEG[7] ;
 wire \Tile_X2Y1_W6BEG[8] ;
 wire \Tile_X2Y1_W6BEG[9] ;
 wire \Tile_X2Y1_WW4BEG[0] ;
 wire \Tile_X2Y1_WW4BEG[10] ;
 wire \Tile_X2Y1_WW4BEG[11] ;
 wire \Tile_X2Y1_WW4BEG[12] ;
 wire \Tile_X2Y1_WW4BEG[13] ;
 wire \Tile_X2Y1_WW4BEG[14] ;
 wire \Tile_X2Y1_WW4BEG[15] ;
 wire \Tile_X2Y1_WW4BEG[1] ;
 wire \Tile_X2Y1_WW4BEG[2] ;
 wire \Tile_X2Y1_WW4BEG[3] ;
 wire \Tile_X2Y1_WW4BEG[4] ;
 wire \Tile_X2Y1_WW4BEG[5] ;
 wire \Tile_X2Y1_WW4BEG[6] ;
 wire \Tile_X2Y1_WW4BEG[7] ;
 wire \Tile_X2Y1_WW4BEG[8] ;
 wire \Tile_X2Y1_WW4BEG[9] ;
 wire Tile_X2Y2_Co;
 wire \Tile_X2Y2_E1BEG[0] ;
 wire \Tile_X2Y2_E1BEG[1] ;
 wire \Tile_X2Y2_E1BEG[2] ;
 wire \Tile_X2Y2_E1BEG[3] ;
 wire \Tile_X2Y2_E2BEG[0] ;
 wire \Tile_X2Y2_E2BEG[1] ;
 wire \Tile_X2Y2_E2BEG[2] ;
 wire \Tile_X2Y2_E2BEG[3] ;
 wire \Tile_X2Y2_E2BEG[4] ;
 wire \Tile_X2Y2_E2BEG[5] ;
 wire \Tile_X2Y2_E2BEG[6] ;
 wire \Tile_X2Y2_E2BEG[7] ;
 wire \Tile_X2Y2_E2BEGb[0] ;
 wire \Tile_X2Y2_E2BEGb[1] ;
 wire \Tile_X2Y2_E2BEGb[2] ;
 wire \Tile_X2Y2_E2BEGb[3] ;
 wire \Tile_X2Y2_E2BEGb[4] ;
 wire \Tile_X2Y2_E2BEGb[5] ;
 wire \Tile_X2Y2_E2BEGb[6] ;
 wire \Tile_X2Y2_E2BEGb[7] ;
 wire \Tile_X2Y2_E6BEG[0] ;
 wire \Tile_X2Y2_E6BEG[10] ;
 wire \Tile_X2Y2_E6BEG[11] ;
 wire \Tile_X2Y2_E6BEG[1] ;
 wire \Tile_X2Y2_E6BEG[2] ;
 wire \Tile_X2Y2_E6BEG[3] ;
 wire \Tile_X2Y2_E6BEG[4] ;
 wire \Tile_X2Y2_E6BEG[5] ;
 wire \Tile_X2Y2_E6BEG[6] ;
 wire \Tile_X2Y2_E6BEG[7] ;
 wire \Tile_X2Y2_E6BEG[8] ;
 wire \Tile_X2Y2_E6BEG[9] ;
 wire \Tile_X2Y2_EE4BEG[0] ;
 wire \Tile_X2Y2_EE4BEG[10] ;
 wire \Tile_X2Y2_EE4BEG[11] ;
 wire \Tile_X2Y2_EE4BEG[12] ;
 wire \Tile_X2Y2_EE4BEG[13] ;
 wire \Tile_X2Y2_EE4BEG[14] ;
 wire \Tile_X2Y2_EE4BEG[15] ;
 wire \Tile_X2Y2_EE4BEG[1] ;
 wire \Tile_X2Y2_EE4BEG[2] ;
 wire \Tile_X2Y2_EE4BEG[3] ;
 wire \Tile_X2Y2_EE4BEG[4] ;
 wire \Tile_X2Y2_EE4BEG[5] ;
 wire \Tile_X2Y2_EE4BEG[6] ;
 wire \Tile_X2Y2_EE4BEG[7] ;
 wire \Tile_X2Y2_EE4BEG[8] ;
 wire \Tile_X2Y2_EE4BEG[9] ;
 wire \Tile_X2Y2_FrameData_O[0] ;
 wire \Tile_X2Y2_FrameData_O[10] ;
 wire \Tile_X2Y2_FrameData_O[11] ;
 wire \Tile_X2Y2_FrameData_O[12] ;
 wire \Tile_X2Y2_FrameData_O[13] ;
 wire \Tile_X2Y2_FrameData_O[14] ;
 wire \Tile_X2Y2_FrameData_O[15] ;
 wire \Tile_X2Y2_FrameData_O[16] ;
 wire \Tile_X2Y2_FrameData_O[17] ;
 wire \Tile_X2Y2_FrameData_O[18] ;
 wire \Tile_X2Y2_FrameData_O[19] ;
 wire \Tile_X2Y2_FrameData_O[1] ;
 wire \Tile_X2Y2_FrameData_O[20] ;
 wire \Tile_X2Y2_FrameData_O[21] ;
 wire \Tile_X2Y2_FrameData_O[22] ;
 wire \Tile_X2Y2_FrameData_O[23] ;
 wire \Tile_X2Y2_FrameData_O[24] ;
 wire \Tile_X2Y2_FrameData_O[25] ;
 wire \Tile_X2Y2_FrameData_O[26] ;
 wire \Tile_X2Y2_FrameData_O[27] ;
 wire \Tile_X2Y2_FrameData_O[28] ;
 wire \Tile_X2Y2_FrameData_O[29] ;
 wire \Tile_X2Y2_FrameData_O[2] ;
 wire \Tile_X2Y2_FrameData_O[30] ;
 wire \Tile_X2Y2_FrameData_O[31] ;
 wire \Tile_X2Y2_FrameData_O[3] ;
 wire \Tile_X2Y2_FrameData_O[4] ;
 wire \Tile_X2Y2_FrameData_O[5] ;
 wire \Tile_X2Y2_FrameData_O[6] ;
 wire \Tile_X2Y2_FrameData_O[7] ;
 wire \Tile_X2Y2_FrameData_O[8] ;
 wire \Tile_X2Y2_FrameData_O[9] ;
 wire \Tile_X2Y2_FrameStrobe_O[0] ;
 wire \Tile_X2Y2_FrameStrobe_O[10] ;
 wire \Tile_X2Y2_FrameStrobe_O[11] ;
 wire \Tile_X2Y2_FrameStrobe_O[12] ;
 wire \Tile_X2Y2_FrameStrobe_O[13] ;
 wire \Tile_X2Y2_FrameStrobe_O[14] ;
 wire \Tile_X2Y2_FrameStrobe_O[15] ;
 wire \Tile_X2Y2_FrameStrobe_O[16] ;
 wire \Tile_X2Y2_FrameStrobe_O[17] ;
 wire \Tile_X2Y2_FrameStrobe_O[18] ;
 wire \Tile_X2Y2_FrameStrobe_O[19] ;
 wire \Tile_X2Y2_FrameStrobe_O[1] ;
 wire \Tile_X2Y2_FrameStrobe_O[2] ;
 wire \Tile_X2Y2_FrameStrobe_O[3] ;
 wire \Tile_X2Y2_FrameStrobe_O[4] ;
 wire \Tile_X2Y2_FrameStrobe_O[5] ;
 wire \Tile_X2Y2_FrameStrobe_O[6] ;
 wire \Tile_X2Y2_FrameStrobe_O[7] ;
 wire \Tile_X2Y2_FrameStrobe_O[8] ;
 wire \Tile_X2Y2_FrameStrobe_O[9] ;
 wire \Tile_X2Y2_N1BEG[0] ;
 wire \Tile_X2Y2_N1BEG[1] ;
 wire \Tile_X2Y2_N1BEG[2] ;
 wire \Tile_X2Y2_N1BEG[3] ;
 wire \Tile_X2Y2_N2BEG[0] ;
 wire \Tile_X2Y2_N2BEG[1] ;
 wire \Tile_X2Y2_N2BEG[2] ;
 wire \Tile_X2Y2_N2BEG[3] ;
 wire \Tile_X2Y2_N2BEG[4] ;
 wire \Tile_X2Y2_N2BEG[5] ;
 wire \Tile_X2Y2_N2BEG[6] ;
 wire \Tile_X2Y2_N2BEG[7] ;
 wire \Tile_X2Y2_N2BEGb[0] ;
 wire \Tile_X2Y2_N2BEGb[1] ;
 wire \Tile_X2Y2_N2BEGb[2] ;
 wire \Tile_X2Y2_N2BEGb[3] ;
 wire \Tile_X2Y2_N2BEGb[4] ;
 wire \Tile_X2Y2_N2BEGb[5] ;
 wire \Tile_X2Y2_N2BEGb[6] ;
 wire \Tile_X2Y2_N2BEGb[7] ;
 wire \Tile_X2Y2_N4BEG[0] ;
 wire \Tile_X2Y2_N4BEG[10] ;
 wire \Tile_X2Y2_N4BEG[11] ;
 wire \Tile_X2Y2_N4BEG[12] ;
 wire \Tile_X2Y2_N4BEG[13] ;
 wire \Tile_X2Y2_N4BEG[14] ;
 wire \Tile_X2Y2_N4BEG[15] ;
 wire \Tile_X2Y2_N4BEG[1] ;
 wire \Tile_X2Y2_N4BEG[2] ;
 wire \Tile_X2Y2_N4BEG[3] ;
 wire \Tile_X2Y2_N4BEG[4] ;
 wire \Tile_X2Y2_N4BEG[5] ;
 wire \Tile_X2Y2_N4BEG[6] ;
 wire \Tile_X2Y2_N4BEG[7] ;
 wire \Tile_X2Y2_N4BEG[8] ;
 wire \Tile_X2Y2_N4BEG[9] ;
 wire \Tile_X2Y2_NN4BEG[0] ;
 wire \Tile_X2Y2_NN4BEG[10] ;
 wire \Tile_X2Y2_NN4BEG[11] ;
 wire \Tile_X2Y2_NN4BEG[12] ;
 wire \Tile_X2Y2_NN4BEG[13] ;
 wire \Tile_X2Y2_NN4BEG[14] ;
 wire \Tile_X2Y2_NN4BEG[15] ;
 wire \Tile_X2Y2_NN4BEG[1] ;
 wire \Tile_X2Y2_NN4BEG[2] ;
 wire \Tile_X2Y2_NN4BEG[3] ;
 wire \Tile_X2Y2_NN4BEG[4] ;
 wire \Tile_X2Y2_NN4BEG[5] ;
 wire \Tile_X2Y2_NN4BEG[6] ;
 wire \Tile_X2Y2_NN4BEG[7] ;
 wire \Tile_X2Y2_NN4BEG[8] ;
 wire \Tile_X2Y2_NN4BEG[9] ;
 wire \Tile_X2Y2_S1BEG[0] ;
 wire \Tile_X2Y2_S1BEG[1] ;
 wire \Tile_X2Y2_S1BEG[2] ;
 wire \Tile_X2Y2_S1BEG[3] ;
 wire \Tile_X2Y2_S2BEG[0] ;
 wire \Tile_X2Y2_S2BEG[1] ;
 wire \Tile_X2Y2_S2BEG[2] ;
 wire \Tile_X2Y2_S2BEG[3] ;
 wire \Tile_X2Y2_S2BEG[4] ;
 wire \Tile_X2Y2_S2BEG[5] ;
 wire \Tile_X2Y2_S2BEG[6] ;
 wire \Tile_X2Y2_S2BEG[7] ;
 wire \Tile_X2Y2_S2BEGb[0] ;
 wire \Tile_X2Y2_S2BEGb[1] ;
 wire \Tile_X2Y2_S2BEGb[2] ;
 wire \Tile_X2Y2_S2BEGb[3] ;
 wire \Tile_X2Y2_S2BEGb[4] ;
 wire \Tile_X2Y2_S2BEGb[5] ;
 wire \Tile_X2Y2_S2BEGb[6] ;
 wire \Tile_X2Y2_S2BEGb[7] ;
 wire \Tile_X2Y2_S4BEG[0] ;
 wire \Tile_X2Y2_S4BEG[10] ;
 wire \Tile_X2Y2_S4BEG[11] ;
 wire \Tile_X2Y2_S4BEG[12] ;
 wire \Tile_X2Y2_S4BEG[13] ;
 wire \Tile_X2Y2_S4BEG[14] ;
 wire \Tile_X2Y2_S4BEG[15] ;
 wire \Tile_X2Y2_S4BEG[1] ;
 wire \Tile_X2Y2_S4BEG[2] ;
 wire \Tile_X2Y2_S4BEG[3] ;
 wire \Tile_X2Y2_S4BEG[4] ;
 wire \Tile_X2Y2_S4BEG[5] ;
 wire \Tile_X2Y2_S4BEG[6] ;
 wire \Tile_X2Y2_S4BEG[7] ;
 wire \Tile_X2Y2_S4BEG[8] ;
 wire \Tile_X2Y2_S4BEG[9] ;
 wire \Tile_X2Y2_SS4BEG[0] ;
 wire \Tile_X2Y2_SS4BEG[10] ;
 wire \Tile_X2Y2_SS4BEG[11] ;
 wire \Tile_X2Y2_SS4BEG[12] ;
 wire \Tile_X2Y2_SS4BEG[13] ;
 wire \Tile_X2Y2_SS4BEG[14] ;
 wire \Tile_X2Y2_SS4BEG[15] ;
 wire \Tile_X2Y2_SS4BEG[1] ;
 wire \Tile_X2Y2_SS4BEG[2] ;
 wire \Tile_X2Y2_SS4BEG[3] ;
 wire \Tile_X2Y2_SS4BEG[4] ;
 wire \Tile_X2Y2_SS4BEG[5] ;
 wire \Tile_X2Y2_SS4BEG[6] ;
 wire \Tile_X2Y2_SS4BEG[7] ;
 wire \Tile_X2Y2_SS4BEG[8] ;
 wire \Tile_X2Y2_SS4BEG[9] ;
 wire Tile_X2Y2_UserCLKo;
 wire \Tile_X2Y2_W1BEG[0] ;
 wire \Tile_X2Y2_W1BEG[1] ;
 wire \Tile_X2Y2_W1BEG[2] ;
 wire \Tile_X2Y2_W1BEG[3] ;
 wire \Tile_X2Y2_W2BEG[0] ;
 wire \Tile_X2Y2_W2BEG[1] ;
 wire \Tile_X2Y2_W2BEG[2] ;
 wire \Tile_X2Y2_W2BEG[3] ;
 wire \Tile_X2Y2_W2BEG[4] ;
 wire \Tile_X2Y2_W2BEG[5] ;
 wire \Tile_X2Y2_W2BEG[6] ;
 wire \Tile_X2Y2_W2BEG[7] ;
 wire \Tile_X2Y2_W2BEGb[0] ;
 wire \Tile_X2Y2_W2BEGb[1] ;
 wire \Tile_X2Y2_W2BEGb[2] ;
 wire \Tile_X2Y2_W2BEGb[3] ;
 wire \Tile_X2Y2_W2BEGb[4] ;
 wire \Tile_X2Y2_W2BEGb[5] ;
 wire \Tile_X2Y2_W2BEGb[6] ;
 wire \Tile_X2Y2_W2BEGb[7] ;
 wire \Tile_X2Y2_W6BEG[0] ;
 wire \Tile_X2Y2_W6BEG[10] ;
 wire \Tile_X2Y2_W6BEG[11] ;
 wire \Tile_X2Y2_W6BEG[1] ;
 wire \Tile_X2Y2_W6BEG[2] ;
 wire \Tile_X2Y2_W6BEG[3] ;
 wire \Tile_X2Y2_W6BEG[4] ;
 wire \Tile_X2Y2_W6BEG[5] ;
 wire \Tile_X2Y2_W6BEG[6] ;
 wire \Tile_X2Y2_W6BEG[7] ;
 wire \Tile_X2Y2_W6BEG[8] ;
 wire \Tile_X2Y2_W6BEG[9] ;
 wire \Tile_X2Y2_WW4BEG[0] ;
 wire \Tile_X2Y2_WW4BEG[10] ;
 wire \Tile_X2Y2_WW4BEG[11] ;
 wire \Tile_X2Y2_WW4BEG[12] ;
 wire \Tile_X2Y2_WW4BEG[13] ;
 wire \Tile_X2Y2_WW4BEG[14] ;
 wire \Tile_X2Y2_WW4BEG[15] ;
 wire \Tile_X2Y2_WW4BEG[1] ;
 wire \Tile_X2Y2_WW4BEG[2] ;
 wire \Tile_X2Y2_WW4BEG[3] ;
 wire \Tile_X2Y2_WW4BEG[4] ;
 wire \Tile_X2Y2_WW4BEG[5] ;
 wire \Tile_X2Y2_WW4BEG[6] ;
 wire \Tile_X2Y2_WW4BEG[7] ;
 wire \Tile_X2Y2_WW4BEG[8] ;
 wire \Tile_X2Y2_WW4BEG[9] ;
 wire Tile_X2Y3_Co;
 wire \Tile_X2Y3_E1BEG[0] ;
 wire \Tile_X2Y3_E1BEG[1] ;
 wire \Tile_X2Y3_E1BEG[2] ;
 wire \Tile_X2Y3_E1BEG[3] ;
 wire \Tile_X2Y3_E2BEG[0] ;
 wire \Tile_X2Y3_E2BEG[1] ;
 wire \Tile_X2Y3_E2BEG[2] ;
 wire \Tile_X2Y3_E2BEG[3] ;
 wire \Tile_X2Y3_E2BEG[4] ;
 wire \Tile_X2Y3_E2BEG[5] ;
 wire \Tile_X2Y3_E2BEG[6] ;
 wire \Tile_X2Y3_E2BEG[7] ;
 wire \Tile_X2Y3_E2BEGb[0] ;
 wire \Tile_X2Y3_E2BEGb[1] ;
 wire \Tile_X2Y3_E2BEGb[2] ;
 wire \Tile_X2Y3_E2BEGb[3] ;
 wire \Tile_X2Y3_E2BEGb[4] ;
 wire \Tile_X2Y3_E2BEGb[5] ;
 wire \Tile_X2Y3_E2BEGb[6] ;
 wire \Tile_X2Y3_E2BEGb[7] ;
 wire \Tile_X2Y3_E6BEG[0] ;
 wire \Tile_X2Y3_E6BEG[10] ;
 wire \Tile_X2Y3_E6BEG[11] ;
 wire \Tile_X2Y3_E6BEG[1] ;
 wire \Tile_X2Y3_E6BEG[2] ;
 wire \Tile_X2Y3_E6BEG[3] ;
 wire \Tile_X2Y3_E6BEG[4] ;
 wire \Tile_X2Y3_E6BEG[5] ;
 wire \Tile_X2Y3_E6BEG[6] ;
 wire \Tile_X2Y3_E6BEG[7] ;
 wire \Tile_X2Y3_E6BEG[8] ;
 wire \Tile_X2Y3_E6BEG[9] ;
 wire \Tile_X2Y3_EE4BEG[0] ;
 wire \Tile_X2Y3_EE4BEG[10] ;
 wire \Tile_X2Y3_EE4BEG[11] ;
 wire \Tile_X2Y3_EE4BEG[12] ;
 wire \Tile_X2Y3_EE4BEG[13] ;
 wire \Tile_X2Y3_EE4BEG[14] ;
 wire \Tile_X2Y3_EE4BEG[15] ;
 wire \Tile_X2Y3_EE4BEG[1] ;
 wire \Tile_X2Y3_EE4BEG[2] ;
 wire \Tile_X2Y3_EE4BEG[3] ;
 wire \Tile_X2Y3_EE4BEG[4] ;
 wire \Tile_X2Y3_EE4BEG[5] ;
 wire \Tile_X2Y3_EE4BEG[6] ;
 wire \Tile_X2Y3_EE4BEG[7] ;
 wire \Tile_X2Y3_EE4BEG[8] ;
 wire \Tile_X2Y3_EE4BEG[9] ;
 wire \Tile_X2Y3_FrameData_O[0] ;
 wire \Tile_X2Y3_FrameData_O[10] ;
 wire \Tile_X2Y3_FrameData_O[11] ;
 wire \Tile_X2Y3_FrameData_O[12] ;
 wire \Tile_X2Y3_FrameData_O[13] ;
 wire \Tile_X2Y3_FrameData_O[14] ;
 wire \Tile_X2Y3_FrameData_O[15] ;
 wire \Tile_X2Y3_FrameData_O[16] ;
 wire \Tile_X2Y3_FrameData_O[17] ;
 wire \Tile_X2Y3_FrameData_O[18] ;
 wire \Tile_X2Y3_FrameData_O[19] ;
 wire \Tile_X2Y3_FrameData_O[1] ;
 wire \Tile_X2Y3_FrameData_O[20] ;
 wire \Tile_X2Y3_FrameData_O[21] ;
 wire \Tile_X2Y3_FrameData_O[22] ;
 wire \Tile_X2Y3_FrameData_O[23] ;
 wire \Tile_X2Y3_FrameData_O[24] ;
 wire \Tile_X2Y3_FrameData_O[25] ;
 wire \Tile_X2Y3_FrameData_O[26] ;
 wire \Tile_X2Y3_FrameData_O[27] ;
 wire \Tile_X2Y3_FrameData_O[28] ;
 wire \Tile_X2Y3_FrameData_O[29] ;
 wire \Tile_X2Y3_FrameData_O[2] ;
 wire \Tile_X2Y3_FrameData_O[30] ;
 wire \Tile_X2Y3_FrameData_O[31] ;
 wire \Tile_X2Y3_FrameData_O[3] ;
 wire \Tile_X2Y3_FrameData_O[4] ;
 wire \Tile_X2Y3_FrameData_O[5] ;
 wire \Tile_X2Y3_FrameData_O[6] ;
 wire \Tile_X2Y3_FrameData_O[7] ;
 wire \Tile_X2Y3_FrameData_O[8] ;
 wire \Tile_X2Y3_FrameData_O[9] ;
 wire \Tile_X2Y3_FrameStrobe_O[0] ;
 wire \Tile_X2Y3_FrameStrobe_O[10] ;
 wire \Tile_X2Y3_FrameStrobe_O[11] ;
 wire \Tile_X2Y3_FrameStrobe_O[12] ;
 wire \Tile_X2Y3_FrameStrobe_O[13] ;
 wire \Tile_X2Y3_FrameStrobe_O[14] ;
 wire \Tile_X2Y3_FrameStrobe_O[15] ;
 wire \Tile_X2Y3_FrameStrobe_O[16] ;
 wire \Tile_X2Y3_FrameStrobe_O[17] ;
 wire \Tile_X2Y3_FrameStrobe_O[18] ;
 wire \Tile_X2Y3_FrameStrobe_O[19] ;
 wire \Tile_X2Y3_FrameStrobe_O[1] ;
 wire \Tile_X2Y3_FrameStrobe_O[2] ;
 wire \Tile_X2Y3_FrameStrobe_O[3] ;
 wire \Tile_X2Y3_FrameStrobe_O[4] ;
 wire \Tile_X2Y3_FrameStrobe_O[5] ;
 wire \Tile_X2Y3_FrameStrobe_O[6] ;
 wire \Tile_X2Y3_FrameStrobe_O[7] ;
 wire \Tile_X2Y3_FrameStrobe_O[8] ;
 wire \Tile_X2Y3_FrameStrobe_O[9] ;
 wire \Tile_X2Y3_N1BEG[0] ;
 wire \Tile_X2Y3_N1BEG[1] ;
 wire \Tile_X2Y3_N1BEG[2] ;
 wire \Tile_X2Y3_N1BEG[3] ;
 wire \Tile_X2Y3_N2BEG[0] ;
 wire \Tile_X2Y3_N2BEG[1] ;
 wire \Tile_X2Y3_N2BEG[2] ;
 wire \Tile_X2Y3_N2BEG[3] ;
 wire \Tile_X2Y3_N2BEG[4] ;
 wire \Tile_X2Y3_N2BEG[5] ;
 wire \Tile_X2Y3_N2BEG[6] ;
 wire \Tile_X2Y3_N2BEG[7] ;
 wire \Tile_X2Y3_N2BEGb[0] ;
 wire \Tile_X2Y3_N2BEGb[1] ;
 wire \Tile_X2Y3_N2BEGb[2] ;
 wire \Tile_X2Y3_N2BEGb[3] ;
 wire \Tile_X2Y3_N2BEGb[4] ;
 wire \Tile_X2Y3_N2BEGb[5] ;
 wire \Tile_X2Y3_N2BEGb[6] ;
 wire \Tile_X2Y3_N2BEGb[7] ;
 wire \Tile_X2Y3_N4BEG[0] ;
 wire \Tile_X2Y3_N4BEG[10] ;
 wire \Tile_X2Y3_N4BEG[11] ;
 wire \Tile_X2Y3_N4BEG[12] ;
 wire \Tile_X2Y3_N4BEG[13] ;
 wire \Tile_X2Y3_N4BEG[14] ;
 wire \Tile_X2Y3_N4BEG[15] ;
 wire \Tile_X2Y3_N4BEG[1] ;
 wire \Tile_X2Y3_N4BEG[2] ;
 wire \Tile_X2Y3_N4BEG[3] ;
 wire \Tile_X2Y3_N4BEG[4] ;
 wire \Tile_X2Y3_N4BEG[5] ;
 wire \Tile_X2Y3_N4BEG[6] ;
 wire \Tile_X2Y3_N4BEG[7] ;
 wire \Tile_X2Y3_N4BEG[8] ;
 wire \Tile_X2Y3_N4BEG[9] ;
 wire \Tile_X2Y3_NN4BEG[0] ;
 wire \Tile_X2Y3_NN4BEG[10] ;
 wire \Tile_X2Y3_NN4BEG[11] ;
 wire \Tile_X2Y3_NN4BEG[12] ;
 wire \Tile_X2Y3_NN4BEG[13] ;
 wire \Tile_X2Y3_NN4BEG[14] ;
 wire \Tile_X2Y3_NN4BEG[15] ;
 wire \Tile_X2Y3_NN4BEG[1] ;
 wire \Tile_X2Y3_NN4BEG[2] ;
 wire \Tile_X2Y3_NN4BEG[3] ;
 wire \Tile_X2Y3_NN4BEG[4] ;
 wire \Tile_X2Y3_NN4BEG[5] ;
 wire \Tile_X2Y3_NN4BEG[6] ;
 wire \Tile_X2Y3_NN4BEG[7] ;
 wire \Tile_X2Y3_NN4BEG[8] ;
 wire \Tile_X2Y3_NN4BEG[9] ;
 wire \Tile_X2Y3_S1BEG[0] ;
 wire \Tile_X2Y3_S1BEG[1] ;
 wire \Tile_X2Y3_S1BEG[2] ;
 wire \Tile_X2Y3_S1BEG[3] ;
 wire \Tile_X2Y3_S2BEG[0] ;
 wire \Tile_X2Y3_S2BEG[1] ;
 wire \Tile_X2Y3_S2BEG[2] ;
 wire \Tile_X2Y3_S2BEG[3] ;
 wire \Tile_X2Y3_S2BEG[4] ;
 wire \Tile_X2Y3_S2BEG[5] ;
 wire \Tile_X2Y3_S2BEG[6] ;
 wire \Tile_X2Y3_S2BEG[7] ;
 wire \Tile_X2Y3_S2BEGb[0] ;
 wire \Tile_X2Y3_S2BEGb[1] ;
 wire \Tile_X2Y3_S2BEGb[2] ;
 wire \Tile_X2Y3_S2BEGb[3] ;
 wire \Tile_X2Y3_S2BEGb[4] ;
 wire \Tile_X2Y3_S2BEGb[5] ;
 wire \Tile_X2Y3_S2BEGb[6] ;
 wire \Tile_X2Y3_S2BEGb[7] ;
 wire \Tile_X2Y3_S4BEG[0] ;
 wire \Tile_X2Y3_S4BEG[10] ;
 wire \Tile_X2Y3_S4BEG[11] ;
 wire \Tile_X2Y3_S4BEG[12] ;
 wire \Tile_X2Y3_S4BEG[13] ;
 wire \Tile_X2Y3_S4BEG[14] ;
 wire \Tile_X2Y3_S4BEG[15] ;
 wire \Tile_X2Y3_S4BEG[1] ;
 wire \Tile_X2Y3_S4BEG[2] ;
 wire \Tile_X2Y3_S4BEG[3] ;
 wire \Tile_X2Y3_S4BEG[4] ;
 wire \Tile_X2Y3_S4BEG[5] ;
 wire \Tile_X2Y3_S4BEG[6] ;
 wire \Tile_X2Y3_S4BEG[7] ;
 wire \Tile_X2Y3_S4BEG[8] ;
 wire \Tile_X2Y3_S4BEG[9] ;
 wire \Tile_X2Y3_SS4BEG[0] ;
 wire \Tile_X2Y3_SS4BEG[10] ;
 wire \Tile_X2Y3_SS4BEG[11] ;
 wire \Tile_X2Y3_SS4BEG[12] ;
 wire \Tile_X2Y3_SS4BEG[13] ;
 wire \Tile_X2Y3_SS4BEG[14] ;
 wire \Tile_X2Y3_SS4BEG[15] ;
 wire \Tile_X2Y3_SS4BEG[1] ;
 wire \Tile_X2Y3_SS4BEG[2] ;
 wire \Tile_X2Y3_SS4BEG[3] ;
 wire \Tile_X2Y3_SS4BEG[4] ;
 wire \Tile_X2Y3_SS4BEG[5] ;
 wire \Tile_X2Y3_SS4BEG[6] ;
 wire \Tile_X2Y3_SS4BEG[7] ;
 wire \Tile_X2Y3_SS4BEG[8] ;
 wire \Tile_X2Y3_SS4BEG[9] ;
 wire Tile_X2Y3_UserCLKo;
 wire \Tile_X2Y3_W1BEG[0] ;
 wire \Tile_X2Y3_W1BEG[1] ;
 wire \Tile_X2Y3_W1BEG[2] ;
 wire \Tile_X2Y3_W1BEG[3] ;
 wire \Tile_X2Y3_W2BEG[0] ;
 wire \Tile_X2Y3_W2BEG[1] ;
 wire \Tile_X2Y3_W2BEG[2] ;
 wire \Tile_X2Y3_W2BEG[3] ;
 wire \Tile_X2Y3_W2BEG[4] ;
 wire \Tile_X2Y3_W2BEG[5] ;
 wire \Tile_X2Y3_W2BEG[6] ;
 wire \Tile_X2Y3_W2BEG[7] ;
 wire \Tile_X2Y3_W2BEGb[0] ;
 wire \Tile_X2Y3_W2BEGb[1] ;
 wire \Tile_X2Y3_W2BEGb[2] ;
 wire \Tile_X2Y3_W2BEGb[3] ;
 wire \Tile_X2Y3_W2BEGb[4] ;
 wire \Tile_X2Y3_W2BEGb[5] ;
 wire \Tile_X2Y3_W2BEGb[6] ;
 wire \Tile_X2Y3_W2BEGb[7] ;
 wire \Tile_X2Y3_W6BEG[0] ;
 wire \Tile_X2Y3_W6BEG[10] ;
 wire \Tile_X2Y3_W6BEG[11] ;
 wire \Tile_X2Y3_W6BEG[1] ;
 wire \Tile_X2Y3_W6BEG[2] ;
 wire \Tile_X2Y3_W6BEG[3] ;
 wire \Tile_X2Y3_W6BEG[4] ;
 wire \Tile_X2Y3_W6BEG[5] ;
 wire \Tile_X2Y3_W6BEG[6] ;
 wire \Tile_X2Y3_W6BEG[7] ;
 wire \Tile_X2Y3_W6BEG[8] ;
 wire \Tile_X2Y3_W6BEG[9] ;
 wire \Tile_X2Y3_WW4BEG[0] ;
 wire \Tile_X2Y3_WW4BEG[10] ;
 wire \Tile_X2Y3_WW4BEG[11] ;
 wire \Tile_X2Y3_WW4BEG[12] ;
 wire \Tile_X2Y3_WW4BEG[13] ;
 wire \Tile_X2Y3_WW4BEG[14] ;
 wire \Tile_X2Y3_WW4BEG[15] ;
 wire \Tile_X2Y3_WW4BEG[1] ;
 wire \Tile_X2Y3_WW4BEG[2] ;
 wire \Tile_X2Y3_WW4BEG[3] ;
 wire \Tile_X2Y3_WW4BEG[4] ;
 wire \Tile_X2Y3_WW4BEG[5] ;
 wire \Tile_X2Y3_WW4BEG[6] ;
 wire \Tile_X2Y3_WW4BEG[7] ;
 wire \Tile_X2Y3_WW4BEG[8] ;
 wire \Tile_X2Y3_WW4BEG[9] ;
 wire Tile_X2Y4_Co;
 wire \Tile_X2Y4_E1BEG[0] ;
 wire \Tile_X2Y4_E1BEG[1] ;
 wire \Tile_X2Y4_E1BEG[2] ;
 wire \Tile_X2Y4_E1BEG[3] ;
 wire \Tile_X2Y4_E2BEG[0] ;
 wire \Tile_X2Y4_E2BEG[1] ;
 wire \Tile_X2Y4_E2BEG[2] ;
 wire \Tile_X2Y4_E2BEG[3] ;
 wire \Tile_X2Y4_E2BEG[4] ;
 wire \Tile_X2Y4_E2BEG[5] ;
 wire \Tile_X2Y4_E2BEG[6] ;
 wire \Tile_X2Y4_E2BEG[7] ;
 wire \Tile_X2Y4_E2BEGb[0] ;
 wire \Tile_X2Y4_E2BEGb[1] ;
 wire \Tile_X2Y4_E2BEGb[2] ;
 wire \Tile_X2Y4_E2BEGb[3] ;
 wire \Tile_X2Y4_E2BEGb[4] ;
 wire \Tile_X2Y4_E2BEGb[5] ;
 wire \Tile_X2Y4_E2BEGb[6] ;
 wire \Tile_X2Y4_E2BEGb[7] ;
 wire \Tile_X2Y4_E6BEG[0] ;
 wire \Tile_X2Y4_E6BEG[10] ;
 wire \Tile_X2Y4_E6BEG[11] ;
 wire \Tile_X2Y4_E6BEG[1] ;
 wire \Tile_X2Y4_E6BEG[2] ;
 wire \Tile_X2Y4_E6BEG[3] ;
 wire \Tile_X2Y4_E6BEG[4] ;
 wire \Tile_X2Y4_E6BEG[5] ;
 wire \Tile_X2Y4_E6BEG[6] ;
 wire \Tile_X2Y4_E6BEG[7] ;
 wire \Tile_X2Y4_E6BEG[8] ;
 wire \Tile_X2Y4_E6BEG[9] ;
 wire \Tile_X2Y4_EE4BEG[0] ;
 wire \Tile_X2Y4_EE4BEG[10] ;
 wire \Tile_X2Y4_EE4BEG[11] ;
 wire \Tile_X2Y4_EE4BEG[12] ;
 wire \Tile_X2Y4_EE4BEG[13] ;
 wire \Tile_X2Y4_EE4BEG[14] ;
 wire \Tile_X2Y4_EE4BEG[15] ;
 wire \Tile_X2Y4_EE4BEG[1] ;
 wire \Tile_X2Y4_EE4BEG[2] ;
 wire \Tile_X2Y4_EE4BEG[3] ;
 wire \Tile_X2Y4_EE4BEG[4] ;
 wire \Tile_X2Y4_EE4BEG[5] ;
 wire \Tile_X2Y4_EE4BEG[6] ;
 wire \Tile_X2Y4_EE4BEG[7] ;
 wire \Tile_X2Y4_EE4BEG[8] ;
 wire \Tile_X2Y4_EE4BEG[9] ;
 wire \Tile_X2Y4_FrameData_O[0] ;
 wire \Tile_X2Y4_FrameData_O[10] ;
 wire \Tile_X2Y4_FrameData_O[11] ;
 wire \Tile_X2Y4_FrameData_O[12] ;
 wire \Tile_X2Y4_FrameData_O[13] ;
 wire \Tile_X2Y4_FrameData_O[14] ;
 wire \Tile_X2Y4_FrameData_O[15] ;
 wire \Tile_X2Y4_FrameData_O[16] ;
 wire \Tile_X2Y4_FrameData_O[17] ;
 wire \Tile_X2Y4_FrameData_O[18] ;
 wire \Tile_X2Y4_FrameData_O[19] ;
 wire \Tile_X2Y4_FrameData_O[1] ;
 wire \Tile_X2Y4_FrameData_O[20] ;
 wire \Tile_X2Y4_FrameData_O[21] ;
 wire \Tile_X2Y4_FrameData_O[22] ;
 wire \Tile_X2Y4_FrameData_O[23] ;
 wire \Tile_X2Y4_FrameData_O[24] ;
 wire \Tile_X2Y4_FrameData_O[25] ;
 wire \Tile_X2Y4_FrameData_O[26] ;
 wire \Tile_X2Y4_FrameData_O[27] ;
 wire \Tile_X2Y4_FrameData_O[28] ;
 wire \Tile_X2Y4_FrameData_O[29] ;
 wire \Tile_X2Y4_FrameData_O[2] ;
 wire \Tile_X2Y4_FrameData_O[30] ;
 wire \Tile_X2Y4_FrameData_O[31] ;
 wire \Tile_X2Y4_FrameData_O[3] ;
 wire \Tile_X2Y4_FrameData_O[4] ;
 wire \Tile_X2Y4_FrameData_O[5] ;
 wire \Tile_X2Y4_FrameData_O[6] ;
 wire \Tile_X2Y4_FrameData_O[7] ;
 wire \Tile_X2Y4_FrameData_O[8] ;
 wire \Tile_X2Y4_FrameData_O[9] ;
 wire \Tile_X2Y4_FrameStrobe_O[0] ;
 wire \Tile_X2Y4_FrameStrobe_O[10] ;
 wire \Tile_X2Y4_FrameStrobe_O[11] ;
 wire \Tile_X2Y4_FrameStrobe_O[12] ;
 wire \Tile_X2Y4_FrameStrobe_O[13] ;
 wire \Tile_X2Y4_FrameStrobe_O[14] ;
 wire \Tile_X2Y4_FrameStrobe_O[15] ;
 wire \Tile_X2Y4_FrameStrobe_O[16] ;
 wire \Tile_X2Y4_FrameStrobe_O[17] ;
 wire \Tile_X2Y4_FrameStrobe_O[18] ;
 wire \Tile_X2Y4_FrameStrobe_O[19] ;
 wire \Tile_X2Y4_FrameStrobe_O[1] ;
 wire \Tile_X2Y4_FrameStrobe_O[2] ;
 wire \Tile_X2Y4_FrameStrobe_O[3] ;
 wire \Tile_X2Y4_FrameStrobe_O[4] ;
 wire \Tile_X2Y4_FrameStrobe_O[5] ;
 wire \Tile_X2Y4_FrameStrobe_O[6] ;
 wire \Tile_X2Y4_FrameStrobe_O[7] ;
 wire \Tile_X2Y4_FrameStrobe_O[8] ;
 wire \Tile_X2Y4_FrameStrobe_O[9] ;
 wire \Tile_X2Y4_N1BEG[0] ;
 wire \Tile_X2Y4_N1BEG[1] ;
 wire \Tile_X2Y4_N1BEG[2] ;
 wire \Tile_X2Y4_N1BEG[3] ;
 wire \Tile_X2Y4_N2BEG[0] ;
 wire \Tile_X2Y4_N2BEG[1] ;
 wire \Tile_X2Y4_N2BEG[2] ;
 wire \Tile_X2Y4_N2BEG[3] ;
 wire \Tile_X2Y4_N2BEG[4] ;
 wire \Tile_X2Y4_N2BEG[5] ;
 wire \Tile_X2Y4_N2BEG[6] ;
 wire \Tile_X2Y4_N2BEG[7] ;
 wire \Tile_X2Y4_N2BEGb[0] ;
 wire \Tile_X2Y4_N2BEGb[1] ;
 wire \Tile_X2Y4_N2BEGb[2] ;
 wire \Tile_X2Y4_N2BEGb[3] ;
 wire \Tile_X2Y4_N2BEGb[4] ;
 wire \Tile_X2Y4_N2BEGb[5] ;
 wire \Tile_X2Y4_N2BEGb[6] ;
 wire \Tile_X2Y4_N2BEGb[7] ;
 wire \Tile_X2Y4_N4BEG[0] ;
 wire \Tile_X2Y4_N4BEG[10] ;
 wire \Tile_X2Y4_N4BEG[11] ;
 wire \Tile_X2Y4_N4BEG[12] ;
 wire \Tile_X2Y4_N4BEG[13] ;
 wire \Tile_X2Y4_N4BEG[14] ;
 wire \Tile_X2Y4_N4BEG[15] ;
 wire \Tile_X2Y4_N4BEG[1] ;
 wire \Tile_X2Y4_N4BEG[2] ;
 wire \Tile_X2Y4_N4BEG[3] ;
 wire \Tile_X2Y4_N4BEG[4] ;
 wire \Tile_X2Y4_N4BEG[5] ;
 wire \Tile_X2Y4_N4BEG[6] ;
 wire \Tile_X2Y4_N4BEG[7] ;
 wire \Tile_X2Y4_N4BEG[8] ;
 wire \Tile_X2Y4_N4BEG[9] ;
 wire \Tile_X2Y4_NN4BEG[0] ;
 wire \Tile_X2Y4_NN4BEG[10] ;
 wire \Tile_X2Y4_NN4BEG[11] ;
 wire \Tile_X2Y4_NN4BEG[12] ;
 wire \Tile_X2Y4_NN4BEG[13] ;
 wire \Tile_X2Y4_NN4BEG[14] ;
 wire \Tile_X2Y4_NN4BEG[15] ;
 wire \Tile_X2Y4_NN4BEG[1] ;
 wire \Tile_X2Y4_NN4BEG[2] ;
 wire \Tile_X2Y4_NN4BEG[3] ;
 wire \Tile_X2Y4_NN4BEG[4] ;
 wire \Tile_X2Y4_NN4BEG[5] ;
 wire \Tile_X2Y4_NN4BEG[6] ;
 wire \Tile_X2Y4_NN4BEG[7] ;
 wire \Tile_X2Y4_NN4BEG[8] ;
 wire \Tile_X2Y4_NN4BEG[9] ;
 wire \Tile_X2Y4_S1BEG[0] ;
 wire \Tile_X2Y4_S1BEG[1] ;
 wire \Tile_X2Y4_S1BEG[2] ;
 wire \Tile_X2Y4_S1BEG[3] ;
 wire \Tile_X2Y4_S2BEG[0] ;
 wire \Tile_X2Y4_S2BEG[1] ;
 wire \Tile_X2Y4_S2BEG[2] ;
 wire \Tile_X2Y4_S2BEG[3] ;
 wire \Tile_X2Y4_S2BEG[4] ;
 wire \Tile_X2Y4_S2BEG[5] ;
 wire \Tile_X2Y4_S2BEG[6] ;
 wire \Tile_X2Y4_S2BEG[7] ;
 wire \Tile_X2Y4_S2BEGb[0] ;
 wire \Tile_X2Y4_S2BEGb[1] ;
 wire \Tile_X2Y4_S2BEGb[2] ;
 wire \Tile_X2Y4_S2BEGb[3] ;
 wire \Tile_X2Y4_S2BEGb[4] ;
 wire \Tile_X2Y4_S2BEGb[5] ;
 wire \Tile_X2Y4_S2BEGb[6] ;
 wire \Tile_X2Y4_S2BEGb[7] ;
 wire \Tile_X2Y4_S4BEG[0] ;
 wire \Tile_X2Y4_S4BEG[10] ;
 wire \Tile_X2Y4_S4BEG[11] ;
 wire \Tile_X2Y4_S4BEG[12] ;
 wire \Tile_X2Y4_S4BEG[13] ;
 wire \Tile_X2Y4_S4BEG[14] ;
 wire \Tile_X2Y4_S4BEG[15] ;
 wire \Tile_X2Y4_S4BEG[1] ;
 wire \Tile_X2Y4_S4BEG[2] ;
 wire \Tile_X2Y4_S4BEG[3] ;
 wire \Tile_X2Y4_S4BEG[4] ;
 wire \Tile_X2Y4_S4BEG[5] ;
 wire \Tile_X2Y4_S4BEG[6] ;
 wire \Tile_X2Y4_S4BEG[7] ;
 wire \Tile_X2Y4_S4BEG[8] ;
 wire \Tile_X2Y4_S4BEG[9] ;
 wire \Tile_X2Y4_SS4BEG[0] ;
 wire \Tile_X2Y4_SS4BEG[10] ;
 wire \Tile_X2Y4_SS4BEG[11] ;
 wire \Tile_X2Y4_SS4BEG[12] ;
 wire \Tile_X2Y4_SS4BEG[13] ;
 wire \Tile_X2Y4_SS4BEG[14] ;
 wire \Tile_X2Y4_SS4BEG[15] ;
 wire \Tile_X2Y4_SS4BEG[1] ;
 wire \Tile_X2Y4_SS4BEG[2] ;
 wire \Tile_X2Y4_SS4BEG[3] ;
 wire \Tile_X2Y4_SS4BEG[4] ;
 wire \Tile_X2Y4_SS4BEG[5] ;
 wire \Tile_X2Y4_SS4BEG[6] ;
 wire \Tile_X2Y4_SS4BEG[7] ;
 wire \Tile_X2Y4_SS4BEG[8] ;
 wire \Tile_X2Y4_SS4BEG[9] ;
 wire Tile_X2Y4_UserCLKo;
 wire \Tile_X2Y4_W1BEG[0] ;
 wire \Tile_X2Y4_W1BEG[1] ;
 wire \Tile_X2Y4_W1BEG[2] ;
 wire \Tile_X2Y4_W1BEG[3] ;
 wire \Tile_X2Y4_W2BEG[0] ;
 wire \Tile_X2Y4_W2BEG[1] ;
 wire \Tile_X2Y4_W2BEG[2] ;
 wire \Tile_X2Y4_W2BEG[3] ;
 wire \Tile_X2Y4_W2BEG[4] ;
 wire \Tile_X2Y4_W2BEG[5] ;
 wire \Tile_X2Y4_W2BEG[6] ;
 wire \Tile_X2Y4_W2BEG[7] ;
 wire \Tile_X2Y4_W2BEGb[0] ;
 wire \Tile_X2Y4_W2BEGb[1] ;
 wire \Tile_X2Y4_W2BEGb[2] ;
 wire \Tile_X2Y4_W2BEGb[3] ;
 wire \Tile_X2Y4_W2BEGb[4] ;
 wire \Tile_X2Y4_W2BEGb[5] ;
 wire \Tile_X2Y4_W2BEGb[6] ;
 wire \Tile_X2Y4_W2BEGb[7] ;
 wire \Tile_X2Y4_W6BEG[0] ;
 wire \Tile_X2Y4_W6BEG[10] ;
 wire \Tile_X2Y4_W6BEG[11] ;
 wire \Tile_X2Y4_W6BEG[1] ;
 wire \Tile_X2Y4_W6BEG[2] ;
 wire \Tile_X2Y4_W6BEG[3] ;
 wire \Tile_X2Y4_W6BEG[4] ;
 wire \Tile_X2Y4_W6BEG[5] ;
 wire \Tile_X2Y4_W6BEG[6] ;
 wire \Tile_X2Y4_W6BEG[7] ;
 wire \Tile_X2Y4_W6BEG[8] ;
 wire \Tile_X2Y4_W6BEG[9] ;
 wire \Tile_X2Y4_WW4BEG[0] ;
 wire \Tile_X2Y4_WW4BEG[10] ;
 wire \Tile_X2Y4_WW4BEG[11] ;
 wire \Tile_X2Y4_WW4BEG[12] ;
 wire \Tile_X2Y4_WW4BEG[13] ;
 wire \Tile_X2Y4_WW4BEG[14] ;
 wire \Tile_X2Y4_WW4BEG[15] ;
 wire \Tile_X2Y4_WW4BEG[1] ;
 wire \Tile_X2Y4_WW4BEG[2] ;
 wire \Tile_X2Y4_WW4BEG[3] ;
 wire \Tile_X2Y4_WW4BEG[4] ;
 wire \Tile_X2Y4_WW4BEG[5] ;
 wire \Tile_X2Y4_WW4BEG[6] ;
 wire \Tile_X2Y4_WW4BEG[7] ;
 wire \Tile_X2Y4_WW4BEG[8] ;
 wire \Tile_X2Y4_WW4BEG[9] ;
 wire Tile_X2Y5_Co;
 wire \Tile_X2Y5_E1BEG[0] ;
 wire \Tile_X2Y5_E1BEG[1] ;
 wire \Tile_X2Y5_E1BEG[2] ;
 wire \Tile_X2Y5_E1BEG[3] ;
 wire \Tile_X2Y5_E2BEG[0] ;
 wire \Tile_X2Y5_E2BEG[1] ;
 wire \Tile_X2Y5_E2BEG[2] ;
 wire \Tile_X2Y5_E2BEG[3] ;
 wire \Tile_X2Y5_E2BEG[4] ;
 wire \Tile_X2Y5_E2BEG[5] ;
 wire \Tile_X2Y5_E2BEG[6] ;
 wire \Tile_X2Y5_E2BEG[7] ;
 wire \Tile_X2Y5_E2BEGb[0] ;
 wire \Tile_X2Y5_E2BEGb[1] ;
 wire \Tile_X2Y5_E2BEGb[2] ;
 wire \Tile_X2Y5_E2BEGb[3] ;
 wire \Tile_X2Y5_E2BEGb[4] ;
 wire \Tile_X2Y5_E2BEGb[5] ;
 wire \Tile_X2Y5_E2BEGb[6] ;
 wire \Tile_X2Y5_E2BEGb[7] ;
 wire \Tile_X2Y5_E6BEG[0] ;
 wire \Tile_X2Y5_E6BEG[10] ;
 wire \Tile_X2Y5_E6BEG[11] ;
 wire \Tile_X2Y5_E6BEG[1] ;
 wire \Tile_X2Y5_E6BEG[2] ;
 wire \Tile_X2Y5_E6BEG[3] ;
 wire \Tile_X2Y5_E6BEG[4] ;
 wire \Tile_X2Y5_E6BEG[5] ;
 wire \Tile_X2Y5_E6BEG[6] ;
 wire \Tile_X2Y5_E6BEG[7] ;
 wire \Tile_X2Y5_E6BEG[8] ;
 wire \Tile_X2Y5_E6BEG[9] ;
 wire \Tile_X2Y5_EE4BEG[0] ;
 wire \Tile_X2Y5_EE4BEG[10] ;
 wire \Tile_X2Y5_EE4BEG[11] ;
 wire \Tile_X2Y5_EE4BEG[12] ;
 wire \Tile_X2Y5_EE4BEG[13] ;
 wire \Tile_X2Y5_EE4BEG[14] ;
 wire \Tile_X2Y5_EE4BEG[15] ;
 wire \Tile_X2Y5_EE4BEG[1] ;
 wire \Tile_X2Y5_EE4BEG[2] ;
 wire \Tile_X2Y5_EE4BEG[3] ;
 wire \Tile_X2Y5_EE4BEG[4] ;
 wire \Tile_X2Y5_EE4BEG[5] ;
 wire \Tile_X2Y5_EE4BEG[6] ;
 wire \Tile_X2Y5_EE4BEG[7] ;
 wire \Tile_X2Y5_EE4BEG[8] ;
 wire \Tile_X2Y5_EE4BEG[9] ;
 wire \Tile_X2Y5_FrameData_O[0] ;
 wire \Tile_X2Y5_FrameData_O[10] ;
 wire \Tile_X2Y5_FrameData_O[11] ;
 wire \Tile_X2Y5_FrameData_O[12] ;
 wire \Tile_X2Y5_FrameData_O[13] ;
 wire \Tile_X2Y5_FrameData_O[14] ;
 wire \Tile_X2Y5_FrameData_O[15] ;
 wire \Tile_X2Y5_FrameData_O[16] ;
 wire \Tile_X2Y5_FrameData_O[17] ;
 wire \Tile_X2Y5_FrameData_O[18] ;
 wire \Tile_X2Y5_FrameData_O[19] ;
 wire \Tile_X2Y5_FrameData_O[1] ;
 wire \Tile_X2Y5_FrameData_O[20] ;
 wire \Tile_X2Y5_FrameData_O[21] ;
 wire \Tile_X2Y5_FrameData_O[22] ;
 wire \Tile_X2Y5_FrameData_O[23] ;
 wire \Tile_X2Y5_FrameData_O[24] ;
 wire \Tile_X2Y5_FrameData_O[25] ;
 wire \Tile_X2Y5_FrameData_O[26] ;
 wire \Tile_X2Y5_FrameData_O[27] ;
 wire \Tile_X2Y5_FrameData_O[28] ;
 wire \Tile_X2Y5_FrameData_O[29] ;
 wire \Tile_X2Y5_FrameData_O[2] ;
 wire \Tile_X2Y5_FrameData_O[30] ;
 wire \Tile_X2Y5_FrameData_O[31] ;
 wire \Tile_X2Y5_FrameData_O[3] ;
 wire \Tile_X2Y5_FrameData_O[4] ;
 wire \Tile_X2Y5_FrameData_O[5] ;
 wire \Tile_X2Y5_FrameData_O[6] ;
 wire \Tile_X2Y5_FrameData_O[7] ;
 wire \Tile_X2Y5_FrameData_O[8] ;
 wire \Tile_X2Y5_FrameData_O[9] ;
 wire \Tile_X2Y5_FrameStrobe_O[0] ;
 wire \Tile_X2Y5_FrameStrobe_O[10] ;
 wire \Tile_X2Y5_FrameStrobe_O[11] ;
 wire \Tile_X2Y5_FrameStrobe_O[12] ;
 wire \Tile_X2Y5_FrameStrobe_O[13] ;
 wire \Tile_X2Y5_FrameStrobe_O[14] ;
 wire \Tile_X2Y5_FrameStrobe_O[15] ;
 wire \Tile_X2Y5_FrameStrobe_O[16] ;
 wire \Tile_X2Y5_FrameStrobe_O[17] ;
 wire \Tile_X2Y5_FrameStrobe_O[18] ;
 wire \Tile_X2Y5_FrameStrobe_O[19] ;
 wire \Tile_X2Y5_FrameStrobe_O[1] ;
 wire \Tile_X2Y5_FrameStrobe_O[2] ;
 wire \Tile_X2Y5_FrameStrobe_O[3] ;
 wire \Tile_X2Y5_FrameStrobe_O[4] ;
 wire \Tile_X2Y5_FrameStrobe_O[5] ;
 wire \Tile_X2Y5_FrameStrobe_O[6] ;
 wire \Tile_X2Y5_FrameStrobe_O[7] ;
 wire \Tile_X2Y5_FrameStrobe_O[8] ;
 wire \Tile_X2Y5_FrameStrobe_O[9] ;
 wire \Tile_X2Y5_N1BEG[0] ;
 wire \Tile_X2Y5_N1BEG[1] ;
 wire \Tile_X2Y5_N1BEG[2] ;
 wire \Tile_X2Y5_N1BEG[3] ;
 wire \Tile_X2Y5_N2BEG[0] ;
 wire \Tile_X2Y5_N2BEG[1] ;
 wire \Tile_X2Y5_N2BEG[2] ;
 wire \Tile_X2Y5_N2BEG[3] ;
 wire \Tile_X2Y5_N2BEG[4] ;
 wire \Tile_X2Y5_N2BEG[5] ;
 wire \Tile_X2Y5_N2BEG[6] ;
 wire \Tile_X2Y5_N2BEG[7] ;
 wire \Tile_X2Y5_N2BEGb[0] ;
 wire \Tile_X2Y5_N2BEGb[1] ;
 wire \Tile_X2Y5_N2BEGb[2] ;
 wire \Tile_X2Y5_N2BEGb[3] ;
 wire \Tile_X2Y5_N2BEGb[4] ;
 wire \Tile_X2Y5_N2BEGb[5] ;
 wire \Tile_X2Y5_N2BEGb[6] ;
 wire \Tile_X2Y5_N2BEGb[7] ;
 wire \Tile_X2Y5_N4BEG[0] ;
 wire \Tile_X2Y5_N4BEG[10] ;
 wire \Tile_X2Y5_N4BEG[11] ;
 wire \Tile_X2Y5_N4BEG[12] ;
 wire \Tile_X2Y5_N4BEG[13] ;
 wire \Tile_X2Y5_N4BEG[14] ;
 wire \Tile_X2Y5_N4BEG[15] ;
 wire \Tile_X2Y5_N4BEG[1] ;
 wire \Tile_X2Y5_N4BEG[2] ;
 wire \Tile_X2Y5_N4BEG[3] ;
 wire \Tile_X2Y5_N4BEG[4] ;
 wire \Tile_X2Y5_N4BEG[5] ;
 wire \Tile_X2Y5_N4BEG[6] ;
 wire \Tile_X2Y5_N4BEG[7] ;
 wire \Tile_X2Y5_N4BEG[8] ;
 wire \Tile_X2Y5_N4BEG[9] ;
 wire \Tile_X2Y5_NN4BEG[0] ;
 wire \Tile_X2Y5_NN4BEG[10] ;
 wire \Tile_X2Y5_NN4BEG[11] ;
 wire \Tile_X2Y5_NN4BEG[12] ;
 wire \Tile_X2Y5_NN4BEG[13] ;
 wire \Tile_X2Y5_NN4BEG[14] ;
 wire \Tile_X2Y5_NN4BEG[15] ;
 wire \Tile_X2Y5_NN4BEG[1] ;
 wire \Tile_X2Y5_NN4BEG[2] ;
 wire \Tile_X2Y5_NN4BEG[3] ;
 wire \Tile_X2Y5_NN4BEG[4] ;
 wire \Tile_X2Y5_NN4BEG[5] ;
 wire \Tile_X2Y5_NN4BEG[6] ;
 wire \Tile_X2Y5_NN4BEG[7] ;
 wire \Tile_X2Y5_NN4BEG[8] ;
 wire \Tile_X2Y5_NN4BEG[9] ;
 wire \Tile_X2Y5_S1BEG[0] ;
 wire \Tile_X2Y5_S1BEG[1] ;
 wire \Tile_X2Y5_S1BEG[2] ;
 wire \Tile_X2Y5_S1BEG[3] ;
 wire \Tile_X2Y5_S2BEG[0] ;
 wire \Tile_X2Y5_S2BEG[1] ;
 wire \Tile_X2Y5_S2BEG[2] ;
 wire \Tile_X2Y5_S2BEG[3] ;
 wire \Tile_X2Y5_S2BEG[4] ;
 wire \Tile_X2Y5_S2BEG[5] ;
 wire \Tile_X2Y5_S2BEG[6] ;
 wire \Tile_X2Y5_S2BEG[7] ;
 wire \Tile_X2Y5_S2BEGb[0] ;
 wire \Tile_X2Y5_S2BEGb[1] ;
 wire \Tile_X2Y5_S2BEGb[2] ;
 wire \Tile_X2Y5_S2BEGb[3] ;
 wire \Tile_X2Y5_S2BEGb[4] ;
 wire \Tile_X2Y5_S2BEGb[5] ;
 wire \Tile_X2Y5_S2BEGb[6] ;
 wire \Tile_X2Y5_S2BEGb[7] ;
 wire \Tile_X2Y5_S4BEG[0] ;
 wire \Tile_X2Y5_S4BEG[10] ;
 wire \Tile_X2Y5_S4BEG[11] ;
 wire \Tile_X2Y5_S4BEG[12] ;
 wire \Tile_X2Y5_S4BEG[13] ;
 wire \Tile_X2Y5_S4BEG[14] ;
 wire \Tile_X2Y5_S4BEG[15] ;
 wire \Tile_X2Y5_S4BEG[1] ;
 wire \Tile_X2Y5_S4BEG[2] ;
 wire \Tile_X2Y5_S4BEG[3] ;
 wire \Tile_X2Y5_S4BEG[4] ;
 wire \Tile_X2Y5_S4BEG[5] ;
 wire \Tile_X2Y5_S4BEG[6] ;
 wire \Tile_X2Y5_S4BEG[7] ;
 wire \Tile_X2Y5_S4BEG[8] ;
 wire \Tile_X2Y5_S4BEG[9] ;
 wire \Tile_X2Y5_SS4BEG[0] ;
 wire \Tile_X2Y5_SS4BEG[10] ;
 wire \Tile_X2Y5_SS4BEG[11] ;
 wire \Tile_X2Y5_SS4BEG[12] ;
 wire \Tile_X2Y5_SS4BEG[13] ;
 wire \Tile_X2Y5_SS4BEG[14] ;
 wire \Tile_X2Y5_SS4BEG[15] ;
 wire \Tile_X2Y5_SS4BEG[1] ;
 wire \Tile_X2Y5_SS4BEG[2] ;
 wire \Tile_X2Y5_SS4BEG[3] ;
 wire \Tile_X2Y5_SS4BEG[4] ;
 wire \Tile_X2Y5_SS4BEG[5] ;
 wire \Tile_X2Y5_SS4BEG[6] ;
 wire \Tile_X2Y5_SS4BEG[7] ;
 wire \Tile_X2Y5_SS4BEG[8] ;
 wire \Tile_X2Y5_SS4BEG[9] ;
 wire Tile_X2Y5_UserCLKo;
 wire \Tile_X2Y5_W1BEG[0] ;
 wire \Tile_X2Y5_W1BEG[1] ;
 wire \Tile_X2Y5_W1BEG[2] ;
 wire \Tile_X2Y5_W1BEG[3] ;
 wire \Tile_X2Y5_W2BEG[0] ;
 wire \Tile_X2Y5_W2BEG[1] ;
 wire \Tile_X2Y5_W2BEG[2] ;
 wire \Tile_X2Y5_W2BEG[3] ;
 wire \Tile_X2Y5_W2BEG[4] ;
 wire \Tile_X2Y5_W2BEG[5] ;
 wire \Tile_X2Y5_W2BEG[6] ;
 wire \Tile_X2Y5_W2BEG[7] ;
 wire \Tile_X2Y5_W2BEGb[0] ;
 wire \Tile_X2Y5_W2BEGb[1] ;
 wire \Tile_X2Y5_W2BEGb[2] ;
 wire \Tile_X2Y5_W2BEGb[3] ;
 wire \Tile_X2Y5_W2BEGb[4] ;
 wire \Tile_X2Y5_W2BEGb[5] ;
 wire \Tile_X2Y5_W2BEGb[6] ;
 wire \Tile_X2Y5_W2BEGb[7] ;
 wire \Tile_X2Y5_W6BEG[0] ;
 wire \Tile_X2Y5_W6BEG[10] ;
 wire \Tile_X2Y5_W6BEG[11] ;
 wire \Tile_X2Y5_W6BEG[1] ;
 wire \Tile_X2Y5_W6BEG[2] ;
 wire \Tile_X2Y5_W6BEG[3] ;
 wire \Tile_X2Y5_W6BEG[4] ;
 wire \Tile_X2Y5_W6BEG[5] ;
 wire \Tile_X2Y5_W6BEG[6] ;
 wire \Tile_X2Y5_W6BEG[7] ;
 wire \Tile_X2Y5_W6BEG[8] ;
 wire \Tile_X2Y5_W6BEG[9] ;
 wire \Tile_X2Y5_WW4BEG[0] ;
 wire \Tile_X2Y5_WW4BEG[10] ;
 wire \Tile_X2Y5_WW4BEG[11] ;
 wire \Tile_X2Y5_WW4BEG[12] ;
 wire \Tile_X2Y5_WW4BEG[13] ;
 wire \Tile_X2Y5_WW4BEG[14] ;
 wire \Tile_X2Y5_WW4BEG[15] ;
 wire \Tile_X2Y5_WW4BEG[1] ;
 wire \Tile_X2Y5_WW4BEG[2] ;
 wire \Tile_X2Y5_WW4BEG[3] ;
 wire \Tile_X2Y5_WW4BEG[4] ;
 wire \Tile_X2Y5_WW4BEG[5] ;
 wire \Tile_X2Y5_WW4BEG[6] ;
 wire \Tile_X2Y5_WW4BEG[7] ;
 wire \Tile_X2Y5_WW4BEG[8] ;
 wire \Tile_X2Y5_WW4BEG[9] ;
 wire Tile_X2Y6_Co;
 wire \Tile_X2Y6_E1BEG[0] ;
 wire \Tile_X2Y6_E1BEG[1] ;
 wire \Tile_X2Y6_E1BEG[2] ;
 wire \Tile_X2Y6_E1BEG[3] ;
 wire \Tile_X2Y6_E2BEG[0] ;
 wire \Tile_X2Y6_E2BEG[1] ;
 wire \Tile_X2Y6_E2BEG[2] ;
 wire \Tile_X2Y6_E2BEG[3] ;
 wire \Tile_X2Y6_E2BEG[4] ;
 wire \Tile_X2Y6_E2BEG[5] ;
 wire \Tile_X2Y6_E2BEG[6] ;
 wire \Tile_X2Y6_E2BEG[7] ;
 wire \Tile_X2Y6_E2BEGb[0] ;
 wire \Tile_X2Y6_E2BEGb[1] ;
 wire \Tile_X2Y6_E2BEGb[2] ;
 wire \Tile_X2Y6_E2BEGb[3] ;
 wire \Tile_X2Y6_E2BEGb[4] ;
 wire \Tile_X2Y6_E2BEGb[5] ;
 wire \Tile_X2Y6_E2BEGb[6] ;
 wire \Tile_X2Y6_E2BEGb[7] ;
 wire \Tile_X2Y6_E6BEG[0] ;
 wire \Tile_X2Y6_E6BEG[10] ;
 wire \Tile_X2Y6_E6BEG[11] ;
 wire \Tile_X2Y6_E6BEG[1] ;
 wire \Tile_X2Y6_E6BEG[2] ;
 wire \Tile_X2Y6_E6BEG[3] ;
 wire \Tile_X2Y6_E6BEG[4] ;
 wire \Tile_X2Y6_E6BEG[5] ;
 wire \Tile_X2Y6_E6BEG[6] ;
 wire \Tile_X2Y6_E6BEG[7] ;
 wire \Tile_X2Y6_E6BEG[8] ;
 wire \Tile_X2Y6_E6BEG[9] ;
 wire \Tile_X2Y6_EE4BEG[0] ;
 wire \Tile_X2Y6_EE4BEG[10] ;
 wire \Tile_X2Y6_EE4BEG[11] ;
 wire \Tile_X2Y6_EE4BEG[12] ;
 wire \Tile_X2Y6_EE4BEG[13] ;
 wire \Tile_X2Y6_EE4BEG[14] ;
 wire \Tile_X2Y6_EE4BEG[15] ;
 wire \Tile_X2Y6_EE4BEG[1] ;
 wire \Tile_X2Y6_EE4BEG[2] ;
 wire \Tile_X2Y6_EE4BEG[3] ;
 wire \Tile_X2Y6_EE4BEG[4] ;
 wire \Tile_X2Y6_EE4BEG[5] ;
 wire \Tile_X2Y6_EE4BEG[6] ;
 wire \Tile_X2Y6_EE4BEG[7] ;
 wire \Tile_X2Y6_EE4BEG[8] ;
 wire \Tile_X2Y6_EE4BEG[9] ;
 wire \Tile_X2Y6_FrameData_O[0] ;
 wire \Tile_X2Y6_FrameData_O[10] ;
 wire \Tile_X2Y6_FrameData_O[11] ;
 wire \Tile_X2Y6_FrameData_O[12] ;
 wire \Tile_X2Y6_FrameData_O[13] ;
 wire \Tile_X2Y6_FrameData_O[14] ;
 wire \Tile_X2Y6_FrameData_O[15] ;
 wire \Tile_X2Y6_FrameData_O[16] ;
 wire \Tile_X2Y6_FrameData_O[17] ;
 wire \Tile_X2Y6_FrameData_O[18] ;
 wire \Tile_X2Y6_FrameData_O[19] ;
 wire \Tile_X2Y6_FrameData_O[1] ;
 wire \Tile_X2Y6_FrameData_O[20] ;
 wire \Tile_X2Y6_FrameData_O[21] ;
 wire \Tile_X2Y6_FrameData_O[22] ;
 wire \Tile_X2Y6_FrameData_O[23] ;
 wire \Tile_X2Y6_FrameData_O[24] ;
 wire \Tile_X2Y6_FrameData_O[25] ;
 wire \Tile_X2Y6_FrameData_O[26] ;
 wire \Tile_X2Y6_FrameData_O[27] ;
 wire \Tile_X2Y6_FrameData_O[28] ;
 wire \Tile_X2Y6_FrameData_O[29] ;
 wire \Tile_X2Y6_FrameData_O[2] ;
 wire \Tile_X2Y6_FrameData_O[30] ;
 wire \Tile_X2Y6_FrameData_O[31] ;
 wire \Tile_X2Y6_FrameData_O[3] ;
 wire \Tile_X2Y6_FrameData_O[4] ;
 wire \Tile_X2Y6_FrameData_O[5] ;
 wire \Tile_X2Y6_FrameData_O[6] ;
 wire \Tile_X2Y6_FrameData_O[7] ;
 wire \Tile_X2Y6_FrameData_O[8] ;
 wire \Tile_X2Y6_FrameData_O[9] ;
 wire \Tile_X2Y6_FrameStrobe_O[0] ;
 wire \Tile_X2Y6_FrameStrobe_O[10] ;
 wire \Tile_X2Y6_FrameStrobe_O[11] ;
 wire \Tile_X2Y6_FrameStrobe_O[12] ;
 wire \Tile_X2Y6_FrameStrobe_O[13] ;
 wire \Tile_X2Y6_FrameStrobe_O[14] ;
 wire \Tile_X2Y6_FrameStrobe_O[15] ;
 wire \Tile_X2Y6_FrameStrobe_O[16] ;
 wire \Tile_X2Y6_FrameStrobe_O[17] ;
 wire \Tile_X2Y6_FrameStrobe_O[18] ;
 wire \Tile_X2Y6_FrameStrobe_O[19] ;
 wire \Tile_X2Y6_FrameStrobe_O[1] ;
 wire \Tile_X2Y6_FrameStrobe_O[2] ;
 wire \Tile_X2Y6_FrameStrobe_O[3] ;
 wire \Tile_X2Y6_FrameStrobe_O[4] ;
 wire \Tile_X2Y6_FrameStrobe_O[5] ;
 wire \Tile_X2Y6_FrameStrobe_O[6] ;
 wire \Tile_X2Y6_FrameStrobe_O[7] ;
 wire \Tile_X2Y6_FrameStrobe_O[8] ;
 wire \Tile_X2Y6_FrameStrobe_O[9] ;
 wire \Tile_X2Y6_N1BEG[0] ;
 wire \Tile_X2Y6_N1BEG[1] ;
 wire \Tile_X2Y6_N1BEG[2] ;
 wire \Tile_X2Y6_N1BEG[3] ;
 wire \Tile_X2Y6_N2BEG[0] ;
 wire \Tile_X2Y6_N2BEG[1] ;
 wire \Tile_X2Y6_N2BEG[2] ;
 wire \Tile_X2Y6_N2BEG[3] ;
 wire \Tile_X2Y6_N2BEG[4] ;
 wire \Tile_X2Y6_N2BEG[5] ;
 wire \Tile_X2Y6_N2BEG[6] ;
 wire \Tile_X2Y6_N2BEG[7] ;
 wire \Tile_X2Y6_N2BEGb[0] ;
 wire \Tile_X2Y6_N2BEGb[1] ;
 wire \Tile_X2Y6_N2BEGb[2] ;
 wire \Tile_X2Y6_N2BEGb[3] ;
 wire \Tile_X2Y6_N2BEGb[4] ;
 wire \Tile_X2Y6_N2BEGb[5] ;
 wire \Tile_X2Y6_N2BEGb[6] ;
 wire \Tile_X2Y6_N2BEGb[7] ;
 wire \Tile_X2Y6_N4BEG[0] ;
 wire \Tile_X2Y6_N4BEG[10] ;
 wire \Tile_X2Y6_N4BEG[11] ;
 wire \Tile_X2Y6_N4BEG[12] ;
 wire \Tile_X2Y6_N4BEG[13] ;
 wire \Tile_X2Y6_N4BEG[14] ;
 wire \Tile_X2Y6_N4BEG[15] ;
 wire \Tile_X2Y6_N4BEG[1] ;
 wire \Tile_X2Y6_N4BEG[2] ;
 wire \Tile_X2Y6_N4BEG[3] ;
 wire \Tile_X2Y6_N4BEG[4] ;
 wire \Tile_X2Y6_N4BEG[5] ;
 wire \Tile_X2Y6_N4BEG[6] ;
 wire \Tile_X2Y6_N4BEG[7] ;
 wire \Tile_X2Y6_N4BEG[8] ;
 wire \Tile_X2Y6_N4BEG[9] ;
 wire \Tile_X2Y6_NN4BEG[0] ;
 wire \Tile_X2Y6_NN4BEG[10] ;
 wire \Tile_X2Y6_NN4BEG[11] ;
 wire \Tile_X2Y6_NN4BEG[12] ;
 wire \Tile_X2Y6_NN4BEG[13] ;
 wire \Tile_X2Y6_NN4BEG[14] ;
 wire \Tile_X2Y6_NN4BEG[15] ;
 wire \Tile_X2Y6_NN4BEG[1] ;
 wire \Tile_X2Y6_NN4BEG[2] ;
 wire \Tile_X2Y6_NN4BEG[3] ;
 wire \Tile_X2Y6_NN4BEG[4] ;
 wire \Tile_X2Y6_NN4BEG[5] ;
 wire \Tile_X2Y6_NN4BEG[6] ;
 wire \Tile_X2Y6_NN4BEG[7] ;
 wire \Tile_X2Y6_NN4BEG[8] ;
 wire \Tile_X2Y6_NN4BEG[9] ;
 wire \Tile_X2Y6_S1BEG[0] ;
 wire \Tile_X2Y6_S1BEG[1] ;
 wire \Tile_X2Y6_S1BEG[2] ;
 wire \Tile_X2Y6_S1BEG[3] ;
 wire \Tile_X2Y6_S2BEG[0] ;
 wire \Tile_X2Y6_S2BEG[1] ;
 wire \Tile_X2Y6_S2BEG[2] ;
 wire \Tile_X2Y6_S2BEG[3] ;
 wire \Tile_X2Y6_S2BEG[4] ;
 wire \Tile_X2Y6_S2BEG[5] ;
 wire \Tile_X2Y6_S2BEG[6] ;
 wire \Tile_X2Y6_S2BEG[7] ;
 wire \Tile_X2Y6_S2BEGb[0] ;
 wire \Tile_X2Y6_S2BEGb[1] ;
 wire \Tile_X2Y6_S2BEGb[2] ;
 wire \Tile_X2Y6_S2BEGb[3] ;
 wire \Tile_X2Y6_S2BEGb[4] ;
 wire \Tile_X2Y6_S2BEGb[5] ;
 wire \Tile_X2Y6_S2BEGb[6] ;
 wire \Tile_X2Y6_S2BEGb[7] ;
 wire \Tile_X2Y6_S4BEG[0] ;
 wire \Tile_X2Y6_S4BEG[10] ;
 wire \Tile_X2Y6_S4BEG[11] ;
 wire \Tile_X2Y6_S4BEG[12] ;
 wire \Tile_X2Y6_S4BEG[13] ;
 wire \Tile_X2Y6_S4BEG[14] ;
 wire \Tile_X2Y6_S4BEG[15] ;
 wire \Tile_X2Y6_S4BEG[1] ;
 wire \Tile_X2Y6_S4BEG[2] ;
 wire \Tile_X2Y6_S4BEG[3] ;
 wire \Tile_X2Y6_S4BEG[4] ;
 wire \Tile_X2Y6_S4BEG[5] ;
 wire \Tile_X2Y6_S4BEG[6] ;
 wire \Tile_X2Y6_S4BEG[7] ;
 wire \Tile_X2Y6_S4BEG[8] ;
 wire \Tile_X2Y6_S4BEG[9] ;
 wire \Tile_X2Y6_SS4BEG[0] ;
 wire \Tile_X2Y6_SS4BEG[10] ;
 wire \Tile_X2Y6_SS4BEG[11] ;
 wire \Tile_X2Y6_SS4BEG[12] ;
 wire \Tile_X2Y6_SS4BEG[13] ;
 wire \Tile_X2Y6_SS4BEG[14] ;
 wire \Tile_X2Y6_SS4BEG[15] ;
 wire \Tile_X2Y6_SS4BEG[1] ;
 wire \Tile_X2Y6_SS4BEG[2] ;
 wire \Tile_X2Y6_SS4BEG[3] ;
 wire \Tile_X2Y6_SS4BEG[4] ;
 wire \Tile_X2Y6_SS4BEG[5] ;
 wire \Tile_X2Y6_SS4BEG[6] ;
 wire \Tile_X2Y6_SS4BEG[7] ;
 wire \Tile_X2Y6_SS4BEG[8] ;
 wire \Tile_X2Y6_SS4BEG[9] ;
 wire Tile_X2Y6_UserCLKo;
 wire \Tile_X2Y6_W1BEG[0] ;
 wire \Tile_X2Y6_W1BEG[1] ;
 wire \Tile_X2Y6_W1BEG[2] ;
 wire \Tile_X2Y6_W1BEG[3] ;
 wire \Tile_X2Y6_W2BEG[0] ;
 wire \Tile_X2Y6_W2BEG[1] ;
 wire \Tile_X2Y6_W2BEG[2] ;
 wire \Tile_X2Y6_W2BEG[3] ;
 wire \Tile_X2Y6_W2BEG[4] ;
 wire \Tile_X2Y6_W2BEG[5] ;
 wire \Tile_X2Y6_W2BEG[6] ;
 wire \Tile_X2Y6_W2BEG[7] ;
 wire \Tile_X2Y6_W2BEGb[0] ;
 wire \Tile_X2Y6_W2BEGb[1] ;
 wire \Tile_X2Y6_W2BEGb[2] ;
 wire \Tile_X2Y6_W2BEGb[3] ;
 wire \Tile_X2Y6_W2BEGb[4] ;
 wire \Tile_X2Y6_W2BEGb[5] ;
 wire \Tile_X2Y6_W2BEGb[6] ;
 wire \Tile_X2Y6_W2BEGb[7] ;
 wire \Tile_X2Y6_W6BEG[0] ;
 wire \Tile_X2Y6_W6BEG[10] ;
 wire \Tile_X2Y6_W6BEG[11] ;
 wire \Tile_X2Y6_W6BEG[1] ;
 wire \Tile_X2Y6_W6BEG[2] ;
 wire \Tile_X2Y6_W6BEG[3] ;
 wire \Tile_X2Y6_W6BEG[4] ;
 wire \Tile_X2Y6_W6BEG[5] ;
 wire \Tile_X2Y6_W6BEG[6] ;
 wire \Tile_X2Y6_W6BEG[7] ;
 wire \Tile_X2Y6_W6BEG[8] ;
 wire \Tile_X2Y6_W6BEG[9] ;
 wire \Tile_X2Y6_WW4BEG[0] ;
 wire \Tile_X2Y6_WW4BEG[10] ;
 wire \Tile_X2Y6_WW4BEG[11] ;
 wire \Tile_X2Y6_WW4BEG[12] ;
 wire \Tile_X2Y6_WW4BEG[13] ;
 wire \Tile_X2Y6_WW4BEG[14] ;
 wire \Tile_X2Y6_WW4BEG[15] ;
 wire \Tile_X2Y6_WW4BEG[1] ;
 wire \Tile_X2Y6_WW4BEG[2] ;
 wire \Tile_X2Y6_WW4BEG[3] ;
 wire \Tile_X2Y6_WW4BEG[4] ;
 wire \Tile_X2Y6_WW4BEG[5] ;
 wire \Tile_X2Y6_WW4BEG[6] ;
 wire \Tile_X2Y6_WW4BEG[7] ;
 wire \Tile_X2Y6_WW4BEG[8] ;
 wire \Tile_X2Y6_WW4BEG[9] ;
 wire Tile_X2Y7_Co;
 wire \Tile_X2Y7_E1BEG[0] ;
 wire \Tile_X2Y7_E1BEG[1] ;
 wire \Tile_X2Y7_E1BEG[2] ;
 wire \Tile_X2Y7_E1BEG[3] ;
 wire \Tile_X2Y7_E2BEG[0] ;
 wire \Tile_X2Y7_E2BEG[1] ;
 wire \Tile_X2Y7_E2BEG[2] ;
 wire \Tile_X2Y7_E2BEG[3] ;
 wire \Tile_X2Y7_E2BEG[4] ;
 wire \Tile_X2Y7_E2BEG[5] ;
 wire \Tile_X2Y7_E2BEG[6] ;
 wire \Tile_X2Y7_E2BEG[7] ;
 wire \Tile_X2Y7_E2BEGb[0] ;
 wire \Tile_X2Y7_E2BEGb[1] ;
 wire \Tile_X2Y7_E2BEGb[2] ;
 wire \Tile_X2Y7_E2BEGb[3] ;
 wire \Tile_X2Y7_E2BEGb[4] ;
 wire \Tile_X2Y7_E2BEGb[5] ;
 wire \Tile_X2Y7_E2BEGb[6] ;
 wire \Tile_X2Y7_E2BEGb[7] ;
 wire \Tile_X2Y7_E6BEG[0] ;
 wire \Tile_X2Y7_E6BEG[10] ;
 wire \Tile_X2Y7_E6BEG[11] ;
 wire \Tile_X2Y7_E6BEG[1] ;
 wire \Tile_X2Y7_E6BEG[2] ;
 wire \Tile_X2Y7_E6BEG[3] ;
 wire \Tile_X2Y7_E6BEG[4] ;
 wire \Tile_X2Y7_E6BEG[5] ;
 wire \Tile_X2Y7_E6BEG[6] ;
 wire \Tile_X2Y7_E6BEG[7] ;
 wire \Tile_X2Y7_E6BEG[8] ;
 wire \Tile_X2Y7_E6BEG[9] ;
 wire \Tile_X2Y7_EE4BEG[0] ;
 wire \Tile_X2Y7_EE4BEG[10] ;
 wire \Tile_X2Y7_EE4BEG[11] ;
 wire \Tile_X2Y7_EE4BEG[12] ;
 wire \Tile_X2Y7_EE4BEG[13] ;
 wire \Tile_X2Y7_EE4BEG[14] ;
 wire \Tile_X2Y7_EE4BEG[15] ;
 wire \Tile_X2Y7_EE4BEG[1] ;
 wire \Tile_X2Y7_EE4BEG[2] ;
 wire \Tile_X2Y7_EE4BEG[3] ;
 wire \Tile_X2Y7_EE4BEG[4] ;
 wire \Tile_X2Y7_EE4BEG[5] ;
 wire \Tile_X2Y7_EE4BEG[6] ;
 wire \Tile_X2Y7_EE4BEG[7] ;
 wire \Tile_X2Y7_EE4BEG[8] ;
 wire \Tile_X2Y7_EE4BEG[9] ;
 wire \Tile_X2Y7_FrameData_O[0] ;
 wire \Tile_X2Y7_FrameData_O[10] ;
 wire \Tile_X2Y7_FrameData_O[11] ;
 wire \Tile_X2Y7_FrameData_O[12] ;
 wire \Tile_X2Y7_FrameData_O[13] ;
 wire \Tile_X2Y7_FrameData_O[14] ;
 wire \Tile_X2Y7_FrameData_O[15] ;
 wire \Tile_X2Y7_FrameData_O[16] ;
 wire \Tile_X2Y7_FrameData_O[17] ;
 wire \Tile_X2Y7_FrameData_O[18] ;
 wire \Tile_X2Y7_FrameData_O[19] ;
 wire \Tile_X2Y7_FrameData_O[1] ;
 wire \Tile_X2Y7_FrameData_O[20] ;
 wire \Tile_X2Y7_FrameData_O[21] ;
 wire \Tile_X2Y7_FrameData_O[22] ;
 wire \Tile_X2Y7_FrameData_O[23] ;
 wire \Tile_X2Y7_FrameData_O[24] ;
 wire \Tile_X2Y7_FrameData_O[25] ;
 wire \Tile_X2Y7_FrameData_O[26] ;
 wire \Tile_X2Y7_FrameData_O[27] ;
 wire \Tile_X2Y7_FrameData_O[28] ;
 wire \Tile_X2Y7_FrameData_O[29] ;
 wire \Tile_X2Y7_FrameData_O[2] ;
 wire \Tile_X2Y7_FrameData_O[30] ;
 wire \Tile_X2Y7_FrameData_O[31] ;
 wire \Tile_X2Y7_FrameData_O[3] ;
 wire \Tile_X2Y7_FrameData_O[4] ;
 wire \Tile_X2Y7_FrameData_O[5] ;
 wire \Tile_X2Y7_FrameData_O[6] ;
 wire \Tile_X2Y7_FrameData_O[7] ;
 wire \Tile_X2Y7_FrameData_O[8] ;
 wire \Tile_X2Y7_FrameData_O[9] ;
 wire \Tile_X2Y7_FrameStrobe_O[0] ;
 wire \Tile_X2Y7_FrameStrobe_O[10] ;
 wire \Tile_X2Y7_FrameStrobe_O[11] ;
 wire \Tile_X2Y7_FrameStrobe_O[12] ;
 wire \Tile_X2Y7_FrameStrobe_O[13] ;
 wire \Tile_X2Y7_FrameStrobe_O[14] ;
 wire \Tile_X2Y7_FrameStrobe_O[15] ;
 wire \Tile_X2Y7_FrameStrobe_O[16] ;
 wire \Tile_X2Y7_FrameStrobe_O[17] ;
 wire \Tile_X2Y7_FrameStrobe_O[18] ;
 wire \Tile_X2Y7_FrameStrobe_O[19] ;
 wire \Tile_X2Y7_FrameStrobe_O[1] ;
 wire \Tile_X2Y7_FrameStrobe_O[2] ;
 wire \Tile_X2Y7_FrameStrobe_O[3] ;
 wire \Tile_X2Y7_FrameStrobe_O[4] ;
 wire \Tile_X2Y7_FrameStrobe_O[5] ;
 wire \Tile_X2Y7_FrameStrobe_O[6] ;
 wire \Tile_X2Y7_FrameStrobe_O[7] ;
 wire \Tile_X2Y7_FrameStrobe_O[8] ;
 wire \Tile_X2Y7_FrameStrobe_O[9] ;
 wire \Tile_X2Y7_N1BEG[0] ;
 wire \Tile_X2Y7_N1BEG[1] ;
 wire \Tile_X2Y7_N1BEG[2] ;
 wire \Tile_X2Y7_N1BEG[3] ;
 wire \Tile_X2Y7_N2BEG[0] ;
 wire \Tile_X2Y7_N2BEG[1] ;
 wire \Tile_X2Y7_N2BEG[2] ;
 wire \Tile_X2Y7_N2BEG[3] ;
 wire \Tile_X2Y7_N2BEG[4] ;
 wire \Tile_X2Y7_N2BEG[5] ;
 wire \Tile_X2Y7_N2BEG[6] ;
 wire \Tile_X2Y7_N2BEG[7] ;
 wire \Tile_X2Y7_N2BEGb[0] ;
 wire \Tile_X2Y7_N2BEGb[1] ;
 wire \Tile_X2Y7_N2BEGb[2] ;
 wire \Tile_X2Y7_N2BEGb[3] ;
 wire \Tile_X2Y7_N2BEGb[4] ;
 wire \Tile_X2Y7_N2BEGb[5] ;
 wire \Tile_X2Y7_N2BEGb[6] ;
 wire \Tile_X2Y7_N2BEGb[7] ;
 wire \Tile_X2Y7_N4BEG[0] ;
 wire \Tile_X2Y7_N4BEG[10] ;
 wire \Tile_X2Y7_N4BEG[11] ;
 wire \Tile_X2Y7_N4BEG[12] ;
 wire \Tile_X2Y7_N4BEG[13] ;
 wire \Tile_X2Y7_N4BEG[14] ;
 wire \Tile_X2Y7_N4BEG[15] ;
 wire \Tile_X2Y7_N4BEG[1] ;
 wire \Tile_X2Y7_N4BEG[2] ;
 wire \Tile_X2Y7_N4BEG[3] ;
 wire \Tile_X2Y7_N4BEG[4] ;
 wire \Tile_X2Y7_N4BEG[5] ;
 wire \Tile_X2Y7_N4BEG[6] ;
 wire \Tile_X2Y7_N4BEG[7] ;
 wire \Tile_X2Y7_N4BEG[8] ;
 wire \Tile_X2Y7_N4BEG[9] ;
 wire \Tile_X2Y7_NN4BEG[0] ;
 wire \Tile_X2Y7_NN4BEG[10] ;
 wire \Tile_X2Y7_NN4BEG[11] ;
 wire \Tile_X2Y7_NN4BEG[12] ;
 wire \Tile_X2Y7_NN4BEG[13] ;
 wire \Tile_X2Y7_NN4BEG[14] ;
 wire \Tile_X2Y7_NN4BEG[15] ;
 wire \Tile_X2Y7_NN4BEG[1] ;
 wire \Tile_X2Y7_NN4BEG[2] ;
 wire \Tile_X2Y7_NN4BEG[3] ;
 wire \Tile_X2Y7_NN4BEG[4] ;
 wire \Tile_X2Y7_NN4BEG[5] ;
 wire \Tile_X2Y7_NN4BEG[6] ;
 wire \Tile_X2Y7_NN4BEG[7] ;
 wire \Tile_X2Y7_NN4BEG[8] ;
 wire \Tile_X2Y7_NN4BEG[9] ;
 wire \Tile_X2Y7_S1BEG[0] ;
 wire \Tile_X2Y7_S1BEG[1] ;
 wire \Tile_X2Y7_S1BEG[2] ;
 wire \Tile_X2Y7_S1BEG[3] ;
 wire \Tile_X2Y7_S2BEG[0] ;
 wire \Tile_X2Y7_S2BEG[1] ;
 wire \Tile_X2Y7_S2BEG[2] ;
 wire \Tile_X2Y7_S2BEG[3] ;
 wire \Tile_X2Y7_S2BEG[4] ;
 wire \Tile_X2Y7_S2BEG[5] ;
 wire \Tile_X2Y7_S2BEG[6] ;
 wire \Tile_X2Y7_S2BEG[7] ;
 wire \Tile_X2Y7_S2BEGb[0] ;
 wire \Tile_X2Y7_S2BEGb[1] ;
 wire \Tile_X2Y7_S2BEGb[2] ;
 wire \Tile_X2Y7_S2BEGb[3] ;
 wire \Tile_X2Y7_S2BEGb[4] ;
 wire \Tile_X2Y7_S2BEGb[5] ;
 wire \Tile_X2Y7_S2BEGb[6] ;
 wire \Tile_X2Y7_S2BEGb[7] ;
 wire \Tile_X2Y7_S4BEG[0] ;
 wire \Tile_X2Y7_S4BEG[10] ;
 wire \Tile_X2Y7_S4BEG[11] ;
 wire \Tile_X2Y7_S4BEG[12] ;
 wire \Tile_X2Y7_S4BEG[13] ;
 wire \Tile_X2Y7_S4BEG[14] ;
 wire \Tile_X2Y7_S4BEG[15] ;
 wire \Tile_X2Y7_S4BEG[1] ;
 wire \Tile_X2Y7_S4BEG[2] ;
 wire \Tile_X2Y7_S4BEG[3] ;
 wire \Tile_X2Y7_S4BEG[4] ;
 wire \Tile_X2Y7_S4BEG[5] ;
 wire \Tile_X2Y7_S4BEG[6] ;
 wire \Tile_X2Y7_S4BEG[7] ;
 wire \Tile_X2Y7_S4BEG[8] ;
 wire \Tile_X2Y7_S4BEG[9] ;
 wire \Tile_X2Y7_SS4BEG[0] ;
 wire \Tile_X2Y7_SS4BEG[10] ;
 wire \Tile_X2Y7_SS4BEG[11] ;
 wire \Tile_X2Y7_SS4BEG[12] ;
 wire \Tile_X2Y7_SS4BEG[13] ;
 wire \Tile_X2Y7_SS4BEG[14] ;
 wire \Tile_X2Y7_SS4BEG[15] ;
 wire \Tile_X2Y7_SS4BEG[1] ;
 wire \Tile_X2Y7_SS4BEG[2] ;
 wire \Tile_X2Y7_SS4BEG[3] ;
 wire \Tile_X2Y7_SS4BEG[4] ;
 wire \Tile_X2Y7_SS4BEG[5] ;
 wire \Tile_X2Y7_SS4BEG[6] ;
 wire \Tile_X2Y7_SS4BEG[7] ;
 wire \Tile_X2Y7_SS4BEG[8] ;
 wire \Tile_X2Y7_SS4BEG[9] ;
 wire Tile_X2Y7_UserCLKo;
 wire \Tile_X2Y7_W1BEG[0] ;
 wire \Tile_X2Y7_W1BEG[1] ;
 wire \Tile_X2Y7_W1BEG[2] ;
 wire \Tile_X2Y7_W1BEG[3] ;
 wire \Tile_X2Y7_W2BEG[0] ;
 wire \Tile_X2Y7_W2BEG[1] ;
 wire \Tile_X2Y7_W2BEG[2] ;
 wire \Tile_X2Y7_W2BEG[3] ;
 wire \Tile_X2Y7_W2BEG[4] ;
 wire \Tile_X2Y7_W2BEG[5] ;
 wire \Tile_X2Y7_W2BEG[6] ;
 wire \Tile_X2Y7_W2BEG[7] ;
 wire \Tile_X2Y7_W2BEGb[0] ;
 wire \Tile_X2Y7_W2BEGb[1] ;
 wire \Tile_X2Y7_W2BEGb[2] ;
 wire \Tile_X2Y7_W2BEGb[3] ;
 wire \Tile_X2Y7_W2BEGb[4] ;
 wire \Tile_X2Y7_W2BEGb[5] ;
 wire \Tile_X2Y7_W2BEGb[6] ;
 wire \Tile_X2Y7_W2BEGb[7] ;
 wire \Tile_X2Y7_W6BEG[0] ;
 wire \Tile_X2Y7_W6BEG[10] ;
 wire \Tile_X2Y7_W6BEG[11] ;
 wire \Tile_X2Y7_W6BEG[1] ;
 wire \Tile_X2Y7_W6BEG[2] ;
 wire \Tile_X2Y7_W6BEG[3] ;
 wire \Tile_X2Y7_W6BEG[4] ;
 wire \Tile_X2Y7_W6BEG[5] ;
 wire \Tile_X2Y7_W6BEG[6] ;
 wire \Tile_X2Y7_W6BEG[7] ;
 wire \Tile_X2Y7_W6BEG[8] ;
 wire \Tile_X2Y7_W6BEG[9] ;
 wire \Tile_X2Y7_WW4BEG[0] ;
 wire \Tile_X2Y7_WW4BEG[10] ;
 wire \Tile_X2Y7_WW4BEG[11] ;
 wire \Tile_X2Y7_WW4BEG[12] ;
 wire \Tile_X2Y7_WW4BEG[13] ;
 wire \Tile_X2Y7_WW4BEG[14] ;
 wire \Tile_X2Y7_WW4BEG[15] ;
 wire \Tile_X2Y7_WW4BEG[1] ;
 wire \Tile_X2Y7_WW4BEG[2] ;
 wire \Tile_X2Y7_WW4BEG[3] ;
 wire \Tile_X2Y7_WW4BEG[4] ;
 wire \Tile_X2Y7_WW4BEG[5] ;
 wire \Tile_X2Y7_WW4BEG[6] ;
 wire \Tile_X2Y7_WW4BEG[7] ;
 wire \Tile_X2Y7_WW4BEG[8] ;
 wire \Tile_X2Y7_WW4BEG[9] ;
 wire Tile_X2Y8_Co;
 wire \Tile_X2Y8_E1BEG[0] ;
 wire \Tile_X2Y8_E1BEG[1] ;
 wire \Tile_X2Y8_E1BEG[2] ;
 wire \Tile_X2Y8_E1BEG[3] ;
 wire \Tile_X2Y8_E2BEG[0] ;
 wire \Tile_X2Y8_E2BEG[1] ;
 wire \Tile_X2Y8_E2BEG[2] ;
 wire \Tile_X2Y8_E2BEG[3] ;
 wire \Tile_X2Y8_E2BEG[4] ;
 wire \Tile_X2Y8_E2BEG[5] ;
 wire \Tile_X2Y8_E2BEG[6] ;
 wire \Tile_X2Y8_E2BEG[7] ;
 wire \Tile_X2Y8_E2BEGb[0] ;
 wire \Tile_X2Y8_E2BEGb[1] ;
 wire \Tile_X2Y8_E2BEGb[2] ;
 wire \Tile_X2Y8_E2BEGb[3] ;
 wire \Tile_X2Y8_E2BEGb[4] ;
 wire \Tile_X2Y8_E2BEGb[5] ;
 wire \Tile_X2Y8_E2BEGb[6] ;
 wire \Tile_X2Y8_E2BEGb[7] ;
 wire \Tile_X2Y8_E6BEG[0] ;
 wire \Tile_X2Y8_E6BEG[10] ;
 wire \Tile_X2Y8_E6BEG[11] ;
 wire \Tile_X2Y8_E6BEG[1] ;
 wire \Tile_X2Y8_E6BEG[2] ;
 wire \Tile_X2Y8_E6BEG[3] ;
 wire \Tile_X2Y8_E6BEG[4] ;
 wire \Tile_X2Y8_E6BEG[5] ;
 wire \Tile_X2Y8_E6BEG[6] ;
 wire \Tile_X2Y8_E6BEG[7] ;
 wire \Tile_X2Y8_E6BEG[8] ;
 wire \Tile_X2Y8_E6BEG[9] ;
 wire \Tile_X2Y8_EE4BEG[0] ;
 wire \Tile_X2Y8_EE4BEG[10] ;
 wire \Tile_X2Y8_EE4BEG[11] ;
 wire \Tile_X2Y8_EE4BEG[12] ;
 wire \Tile_X2Y8_EE4BEG[13] ;
 wire \Tile_X2Y8_EE4BEG[14] ;
 wire \Tile_X2Y8_EE4BEG[15] ;
 wire \Tile_X2Y8_EE4BEG[1] ;
 wire \Tile_X2Y8_EE4BEG[2] ;
 wire \Tile_X2Y8_EE4BEG[3] ;
 wire \Tile_X2Y8_EE4BEG[4] ;
 wire \Tile_X2Y8_EE4BEG[5] ;
 wire \Tile_X2Y8_EE4BEG[6] ;
 wire \Tile_X2Y8_EE4BEG[7] ;
 wire \Tile_X2Y8_EE4BEG[8] ;
 wire \Tile_X2Y8_EE4BEG[9] ;
 wire \Tile_X2Y8_FrameData_O[0] ;
 wire \Tile_X2Y8_FrameData_O[10] ;
 wire \Tile_X2Y8_FrameData_O[11] ;
 wire \Tile_X2Y8_FrameData_O[12] ;
 wire \Tile_X2Y8_FrameData_O[13] ;
 wire \Tile_X2Y8_FrameData_O[14] ;
 wire \Tile_X2Y8_FrameData_O[15] ;
 wire \Tile_X2Y8_FrameData_O[16] ;
 wire \Tile_X2Y8_FrameData_O[17] ;
 wire \Tile_X2Y8_FrameData_O[18] ;
 wire \Tile_X2Y8_FrameData_O[19] ;
 wire \Tile_X2Y8_FrameData_O[1] ;
 wire \Tile_X2Y8_FrameData_O[20] ;
 wire \Tile_X2Y8_FrameData_O[21] ;
 wire \Tile_X2Y8_FrameData_O[22] ;
 wire \Tile_X2Y8_FrameData_O[23] ;
 wire \Tile_X2Y8_FrameData_O[24] ;
 wire \Tile_X2Y8_FrameData_O[25] ;
 wire \Tile_X2Y8_FrameData_O[26] ;
 wire \Tile_X2Y8_FrameData_O[27] ;
 wire \Tile_X2Y8_FrameData_O[28] ;
 wire \Tile_X2Y8_FrameData_O[29] ;
 wire \Tile_X2Y8_FrameData_O[2] ;
 wire \Tile_X2Y8_FrameData_O[30] ;
 wire \Tile_X2Y8_FrameData_O[31] ;
 wire \Tile_X2Y8_FrameData_O[3] ;
 wire \Tile_X2Y8_FrameData_O[4] ;
 wire \Tile_X2Y8_FrameData_O[5] ;
 wire \Tile_X2Y8_FrameData_O[6] ;
 wire \Tile_X2Y8_FrameData_O[7] ;
 wire \Tile_X2Y8_FrameData_O[8] ;
 wire \Tile_X2Y8_FrameData_O[9] ;
 wire \Tile_X2Y8_FrameStrobe_O[0] ;
 wire \Tile_X2Y8_FrameStrobe_O[10] ;
 wire \Tile_X2Y8_FrameStrobe_O[11] ;
 wire \Tile_X2Y8_FrameStrobe_O[12] ;
 wire \Tile_X2Y8_FrameStrobe_O[13] ;
 wire \Tile_X2Y8_FrameStrobe_O[14] ;
 wire \Tile_X2Y8_FrameStrobe_O[15] ;
 wire \Tile_X2Y8_FrameStrobe_O[16] ;
 wire \Tile_X2Y8_FrameStrobe_O[17] ;
 wire \Tile_X2Y8_FrameStrobe_O[18] ;
 wire \Tile_X2Y8_FrameStrobe_O[19] ;
 wire \Tile_X2Y8_FrameStrobe_O[1] ;
 wire \Tile_X2Y8_FrameStrobe_O[2] ;
 wire \Tile_X2Y8_FrameStrobe_O[3] ;
 wire \Tile_X2Y8_FrameStrobe_O[4] ;
 wire \Tile_X2Y8_FrameStrobe_O[5] ;
 wire \Tile_X2Y8_FrameStrobe_O[6] ;
 wire \Tile_X2Y8_FrameStrobe_O[7] ;
 wire \Tile_X2Y8_FrameStrobe_O[8] ;
 wire \Tile_X2Y8_FrameStrobe_O[9] ;
 wire \Tile_X2Y8_N1BEG[0] ;
 wire \Tile_X2Y8_N1BEG[1] ;
 wire \Tile_X2Y8_N1BEG[2] ;
 wire \Tile_X2Y8_N1BEG[3] ;
 wire \Tile_X2Y8_N2BEG[0] ;
 wire \Tile_X2Y8_N2BEG[1] ;
 wire \Tile_X2Y8_N2BEG[2] ;
 wire \Tile_X2Y8_N2BEG[3] ;
 wire \Tile_X2Y8_N2BEG[4] ;
 wire \Tile_X2Y8_N2BEG[5] ;
 wire \Tile_X2Y8_N2BEG[6] ;
 wire \Tile_X2Y8_N2BEG[7] ;
 wire \Tile_X2Y8_N2BEGb[0] ;
 wire \Tile_X2Y8_N2BEGb[1] ;
 wire \Tile_X2Y8_N2BEGb[2] ;
 wire \Tile_X2Y8_N2BEGb[3] ;
 wire \Tile_X2Y8_N2BEGb[4] ;
 wire \Tile_X2Y8_N2BEGb[5] ;
 wire \Tile_X2Y8_N2BEGb[6] ;
 wire \Tile_X2Y8_N2BEGb[7] ;
 wire \Tile_X2Y8_N4BEG[0] ;
 wire \Tile_X2Y8_N4BEG[10] ;
 wire \Tile_X2Y8_N4BEG[11] ;
 wire \Tile_X2Y8_N4BEG[12] ;
 wire \Tile_X2Y8_N4BEG[13] ;
 wire \Tile_X2Y8_N4BEG[14] ;
 wire \Tile_X2Y8_N4BEG[15] ;
 wire \Tile_X2Y8_N4BEG[1] ;
 wire \Tile_X2Y8_N4BEG[2] ;
 wire \Tile_X2Y8_N4BEG[3] ;
 wire \Tile_X2Y8_N4BEG[4] ;
 wire \Tile_X2Y8_N4BEG[5] ;
 wire \Tile_X2Y8_N4BEG[6] ;
 wire \Tile_X2Y8_N4BEG[7] ;
 wire \Tile_X2Y8_N4BEG[8] ;
 wire \Tile_X2Y8_N4BEG[9] ;
 wire \Tile_X2Y8_NN4BEG[0] ;
 wire \Tile_X2Y8_NN4BEG[10] ;
 wire \Tile_X2Y8_NN4BEG[11] ;
 wire \Tile_X2Y8_NN4BEG[12] ;
 wire \Tile_X2Y8_NN4BEG[13] ;
 wire \Tile_X2Y8_NN4BEG[14] ;
 wire \Tile_X2Y8_NN4BEG[15] ;
 wire \Tile_X2Y8_NN4BEG[1] ;
 wire \Tile_X2Y8_NN4BEG[2] ;
 wire \Tile_X2Y8_NN4BEG[3] ;
 wire \Tile_X2Y8_NN4BEG[4] ;
 wire \Tile_X2Y8_NN4BEG[5] ;
 wire \Tile_X2Y8_NN4BEG[6] ;
 wire \Tile_X2Y8_NN4BEG[7] ;
 wire \Tile_X2Y8_NN4BEG[8] ;
 wire \Tile_X2Y8_NN4BEG[9] ;
 wire \Tile_X2Y8_S1BEG[0] ;
 wire \Tile_X2Y8_S1BEG[1] ;
 wire \Tile_X2Y8_S1BEG[2] ;
 wire \Tile_X2Y8_S1BEG[3] ;
 wire \Tile_X2Y8_S2BEG[0] ;
 wire \Tile_X2Y8_S2BEG[1] ;
 wire \Tile_X2Y8_S2BEG[2] ;
 wire \Tile_X2Y8_S2BEG[3] ;
 wire \Tile_X2Y8_S2BEG[4] ;
 wire \Tile_X2Y8_S2BEG[5] ;
 wire \Tile_X2Y8_S2BEG[6] ;
 wire \Tile_X2Y8_S2BEG[7] ;
 wire \Tile_X2Y8_S2BEGb[0] ;
 wire \Tile_X2Y8_S2BEGb[1] ;
 wire \Tile_X2Y8_S2BEGb[2] ;
 wire \Tile_X2Y8_S2BEGb[3] ;
 wire \Tile_X2Y8_S2BEGb[4] ;
 wire \Tile_X2Y8_S2BEGb[5] ;
 wire \Tile_X2Y8_S2BEGb[6] ;
 wire \Tile_X2Y8_S2BEGb[7] ;
 wire \Tile_X2Y8_S4BEG[0] ;
 wire \Tile_X2Y8_S4BEG[10] ;
 wire \Tile_X2Y8_S4BEG[11] ;
 wire \Tile_X2Y8_S4BEG[12] ;
 wire \Tile_X2Y8_S4BEG[13] ;
 wire \Tile_X2Y8_S4BEG[14] ;
 wire \Tile_X2Y8_S4BEG[15] ;
 wire \Tile_X2Y8_S4BEG[1] ;
 wire \Tile_X2Y8_S4BEG[2] ;
 wire \Tile_X2Y8_S4BEG[3] ;
 wire \Tile_X2Y8_S4BEG[4] ;
 wire \Tile_X2Y8_S4BEG[5] ;
 wire \Tile_X2Y8_S4BEG[6] ;
 wire \Tile_X2Y8_S4BEG[7] ;
 wire \Tile_X2Y8_S4BEG[8] ;
 wire \Tile_X2Y8_S4BEG[9] ;
 wire \Tile_X2Y8_SS4BEG[0] ;
 wire \Tile_X2Y8_SS4BEG[10] ;
 wire \Tile_X2Y8_SS4BEG[11] ;
 wire \Tile_X2Y8_SS4BEG[12] ;
 wire \Tile_X2Y8_SS4BEG[13] ;
 wire \Tile_X2Y8_SS4BEG[14] ;
 wire \Tile_X2Y8_SS4BEG[15] ;
 wire \Tile_X2Y8_SS4BEG[1] ;
 wire \Tile_X2Y8_SS4BEG[2] ;
 wire \Tile_X2Y8_SS4BEG[3] ;
 wire \Tile_X2Y8_SS4BEG[4] ;
 wire \Tile_X2Y8_SS4BEG[5] ;
 wire \Tile_X2Y8_SS4BEG[6] ;
 wire \Tile_X2Y8_SS4BEG[7] ;
 wire \Tile_X2Y8_SS4BEG[8] ;
 wire \Tile_X2Y8_SS4BEG[9] ;
 wire Tile_X2Y8_UserCLKo;
 wire \Tile_X2Y8_W1BEG[0] ;
 wire \Tile_X2Y8_W1BEG[1] ;
 wire \Tile_X2Y8_W1BEG[2] ;
 wire \Tile_X2Y8_W1BEG[3] ;
 wire \Tile_X2Y8_W2BEG[0] ;
 wire \Tile_X2Y8_W2BEG[1] ;
 wire \Tile_X2Y8_W2BEG[2] ;
 wire \Tile_X2Y8_W2BEG[3] ;
 wire \Tile_X2Y8_W2BEG[4] ;
 wire \Tile_X2Y8_W2BEG[5] ;
 wire \Tile_X2Y8_W2BEG[6] ;
 wire \Tile_X2Y8_W2BEG[7] ;
 wire \Tile_X2Y8_W2BEGb[0] ;
 wire \Tile_X2Y8_W2BEGb[1] ;
 wire \Tile_X2Y8_W2BEGb[2] ;
 wire \Tile_X2Y8_W2BEGb[3] ;
 wire \Tile_X2Y8_W2BEGb[4] ;
 wire \Tile_X2Y8_W2BEGb[5] ;
 wire \Tile_X2Y8_W2BEGb[6] ;
 wire \Tile_X2Y8_W2BEGb[7] ;
 wire \Tile_X2Y8_W6BEG[0] ;
 wire \Tile_X2Y8_W6BEG[10] ;
 wire \Tile_X2Y8_W6BEG[11] ;
 wire \Tile_X2Y8_W6BEG[1] ;
 wire \Tile_X2Y8_W6BEG[2] ;
 wire \Tile_X2Y8_W6BEG[3] ;
 wire \Tile_X2Y8_W6BEG[4] ;
 wire \Tile_X2Y8_W6BEG[5] ;
 wire \Tile_X2Y8_W6BEG[6] ;
 wire \Tile_X2Y8_W6BEG[7] ;
 wire \Tile_X2Y8_W6BEG[8] ;
 wire \Tile_X2Y8_W6BEG[9] ;
 wire \Tile_X2Y8_WW4BEG[0] ;
 wire \Tile_X2Y8_WW4BEG[10] ;
 wire \Tile_X2Y8_WW4BEG[11] ;
 wire \Tile_X2Y8_WW4BEG[12] ;
 wire \Tile_X2Y8_WW4BEG[13] ;
 wire \Tile_X2Y8_WW4BEG[14] ;
 wire \Tile_X2Y8_WW4BEG[15] ;
 wire \Tile_X2Y8_WW4BEG[1] ;
 wire \Tile_X2Y8_WW4BEG[2] ;
 wire \Tile_X2Y8_WW4BEG[3] ;
 wire \Tile_X2Y8_WW4BEG[4] ;
 wire \Tile_X2Y8_WW4BEG[5] ;
 wire \Tile_X2Y8_WW4BEG[6] ;
 wire \Tile_X2Y8_WW4BEG[7] ;
 wire \Tile_X2Y8_WW4BEG[8] ;
 wire \Tile_X2Y8_WW4BEG[9] ;
 wire Tile_X2Y9_Co;
 wire \Tile_X2Y9_E1BEG[0] ;
 wire \Tile_X2Y9_E1BEG[1] ;
 wire \Tile_X2Y9_E1BEG[2] ;
 wire \Tile_X2Y9_E1BEG[3] ;
 wire \Tile_X2Y9_E2BEG[0] ;
 wire \Tile_X2Y9_E2BEG[1] ;
 wire \Tile_X2Y9_E2BEG[2] ;
 wire \Tile_X2Y9_E2BEG[3] ;
 wire \Tile_X2Y9_E2BEG[4] ;
 wire \Tile_X2Y9_E2BEG[5] ;
 wire \Tile_X2Y9_E2BEG[6] ;
 wire \Tile_X2Y9_E2BEG[7] ;
 wire \Tile_X2Y9_E2BEGb[0] ;
 wire \Tile_X2Y9_E2BEGb[1] ;
 wire \Tile_X2Y9_E2BEGb[2] ;
 wire \Tile_X2Y9_E2BEGb[3] ;
 wire \Tile_X2Y9_E2BEGb[4] ;
 wire \Tile_X2Y9_E2BEGb[5] ;
 wire \Tile_X2Y9_E2BEGb[6] ;
 wire \Tile_X2Y9_E2BEGb[7] ;
 wire \Tile_X2Y9_E6BEG[0] ;
 wire \Tile_X2Y9_E6BEG[10] ;
 wire \Tile_X2Y9_E6BEG[11] ;
 wire \Tile_X2Y9_E6BEG[1] ;
 wire \Tile_X2Y9_E6BEG[2] ;
 wire \Tile_X2Y9_E6BEG[3] ;
 wire \Tile_X2Y9_E6BEG[4] ;
 wire \Tile_X2Y9_E6BEG[5] ;
 wire \Tile_X2Y9_E6BEG[6] ;
 wire \Tile_X2Y9_E6BEG[7] ;
 wire \Tile_X2Y9_E6BEG[8] ;
 wire \Tile_X2Y9_E6BEG[9] ;
 wire \Tile_X2Y9_EE4BEG[0] ;
 wire \Tile_X2Y9_EE4BEG[10] ;
 wire \Tile_X2Y9_EE4BEG[11] ;
 wire \Tile_X2Y9_EE4BEG[12] ;
 wire \Tile_X2Y9_EE4BEG[13] ;
 wire \Tile_X2Y9_EE4BEG[14] ;
 wire \Tile_X2Y9_EE4BEG[15] ;
 wire \Tile_X2Y9_EE4BEG[1] ;
 wire \Tile_X2Y9_EE4BEG[2] ;
 wire \Tile_X2Y9_EE4BEG[3] ;
 wire \Tile_X2Y9_EE4BEG[4] ;
 wire \Tile_X2Y9_EE4BEG[5] ;
 wire \Tile_X2Y9_EE4BEG[6] ;
 wire \Tile_X2Y9_EE4BEG[7] ;
 wire \Tile_X2Y9_EE4BEG[8] ;
 wire \Tile_X2Y9_EE4BEG[9] ;
 wire \Tile_X2Y9_FrameData_O[0] ;
 wire \Tile_X2Y9_FrameData_O[10] ;
 wire \Tile_X2Y9_FrameData_O[11] ;
 wire \Tile_X2Y9_FrameData_O[12] ;
 wire \Tile_X2Y9_FrameData_O[13] ;
 wire \Tile_X2Y9_FrameData_O[14] ;
 wire \Tile_X2Y9_FrameData_O[15] ;
 wire \Tile_X2Y9_FrameData_O[16] ;
 wire \Tile_X2Y9_FrameData_O[17] ;
 wire \Tile_X2Y9_FrameData_O[18] ;
 wire \Tile_X2Y9_FrameData_O[19] ;
 wire \Tile_X2Y9_FrameData_O[1] ;
 wire \Tile_X2Y9_FrameData_O[20] ;
 wire \Tile_X2Y9_FrameData_O[21] ;
 wire \Tile_X2Y9_FrameData_O[22] ;
 wire \Tile_X2Y9_FrameData_O[23] ;
 wire \Tile_X2Y9_FrameData_O[24] ;
 wire \Tile_X2Y9_FrameData_O[25] ;
 wire \Tile_X2Y9_FrameData_O[26] ;
 wire \Tile_X2Y9_FrameData_O[27] ;
 wire \Tile_X2Y9_FrameData_O[28] ;
 wire \Tile_X2Y9_FrameData_O[29] ;
 wire \Tile_X2Y9_FrameData_O[2] ;
 wire \Tile_X2Y9_FrameData_O[30] ;
 wire \Tile_X2Y9_FrameData_O[31] ;
 wire \Tile_X2Y9_FrameData_O[3] ;
 wire \Tile_X2Y9_FrameData_O[4] ;
 wire \Tile_X2Y9_FrameData_O[5] ;
 wire \Tile_X2Y9_FrameData_O[6] ;
 wire \Tile_X2Y9_FrameData_O[7] ;
 wire \Tile_X2Y9_FrameData_O[8] ;
 wire \Tile_X2Y9_FrameData_O[9] ;
 wire \Tile_X2Y9_FrameStrobe_O[0] ;
 wire \Tile_X2Y9_FrameStrobe_O[10] ;
 wire \Tile_X2Y9_FrameStrobe_O[11] ;
 wire \Tile_X2Y9_FrameStrobe_O[12] ;
 wire \Tile_X2Y9_FrameStrobe_O[13] ;
 wire \Tile_X2Y9_FrameStrobe_O[14] ;
 wire \Tile_X2Y9_FrameStrobe_O[15] ;
 wire \Tile_X2Y9_FrameStrobe_O[16] ;
 wire \Tile_X2Y9_FrameStrobe_O[17] ;
 wire \Tile_X2Y9_FrameStrobe_O[18] ;
 wire \Tile_X2Y9_FrameStrobe_O[19] ;
 wire \Tile_X2Y9_FrameStrobe_O[1] ;
 wire \Tile_X2Y9_FrameStrobe_O[2] ;
 wire \Tile_X2Y9_FrameStrobe_O[3] ;
 wire \Tile_X2Y9_FrameStrobe_O[4] ;
 wire \Tile_X2Y9_FrameStrobe_O[5] ;
 wire \Tile_X2Y9_FrameStrobe_O[6] ;
 wire \Tile_X2Y9_FrameStrobe_O[7] ;
 wire \Tile_X2Y9_FrameStrobe_O[8] ;
 wire \Tile_X2Y9_FrameStrobe_O[9] ;
 wire \Tile_X2Y9_N1BEG[0] ;
 wire \Tile_X2Y9_N1BEG[1] ;
 wire \Tile_X2Y9_N1BEG[2] ;
 wire \Tile_X2Y9_N1BEG[3] ;
 wire \Tile_X2Y9_N2BEG[0] ;
 wire \Tile_X2Y9_N2BEG[1] ;
 wire \Tile_X2Y9_N2BEG[2] ;
 wire \Tile_X2Y9_N2BEG[3] ;
 wire \Tile_X2Y9_N2BEG[4] ;
 wire \Tile_X2Y9_N2BEG[5] ;
 wire \Tile_X2Y9_N2BEG[6] ;
 wire \Tile_X2Y9_N2BEG[7] ;
 wire \Tile_X2Y9_N2BEGb[0] ;
 wire \Tile_X2Y9_N2BEGb[1] ;
 wire \Tile_X2Y9_N2BEGb[2] ;
 wire \Tile_X2Y9_N2BEGb[3] ;
 wire \Tile_X2Y9_N2BEGb[4] ;
 wire \Tile_X2Y9_N2BEGb[5] ;
 wire \Tile_X2Y9_N2BEGb[6] ;
 wire \Tile_X2Y9_N2BEGb[7] ;
 wire \Tile_X2Y9_N4BEG[0] ;
 wire \Tile_X2Y9_N4BEG[10] ;
 wire \Tile_X2Y9_N4BEG[11] ;
 wire \Tile_X2Y9_N4BEG[12] ;
 wire \Tile_X2Y9_N4BEG[13] ;
 wire \Tile_X2Y9_N4BEG[14] ;
 wire \Tile_X2Y9_N4BEG[15] ;
 wire \Tile_X2Y9_N4BEG[1] ;
 wire \Tile_X2Y9_N4BEG[2] ;
 wire \Tile_X2Y9_N4BEG[3] ;
 wire \Tile_X2Y9_N4BEG[4] ;
 wire \Tile_X2Y9_N4BEG[5] ;
 wire \Tile_X2Y9_N4BEG[6] ;
 wire \Tile_X2Y9_N4BEG[7] ;
 wire \Tile_X2Y9_N4BEG[8] ;
 wire \Tile_X2Y9_N4BEG[9] ;
 wire \Tile_X2Y9_NN4BEG[0] ;
 wire \Tile_X2Y9_NN4BEG[10] ;
 wire \Tile_X2Y9_NN4BEG[11] ;
 wire \Tile_X2Y9_NN4BEG[12] ;
 wire \Tile_X2Y9_NN4BEG[13] ;
 wire \Tile_X2Y9_NN4BEG[14] ;
 wire \Tile_X2Y9_NN4BEG[15] ;
 wire \Tile_X2Y9_NN4BEG[1] ;
 wire \Tile_X2Y9_NN4BEG[2] ;
 wire \Tile_X2Y9_NN4BEG[3] ;
 wire \Tile_X2Y9_NN4BEG[4] ;
 wire \Tile_X2Y9_NN4BEG[5] ;
 wire \Tile_X2Y9_NN4BEG[6] ;
 wire \Tile_X2Y9_NN4BEG[7] ;
 wire \Tile_X2Y9_NN4BEG[8] ;
 wire \Tile_X2Y9_NN4BEG[9] ;
 wire \Tile_X2Y9_S1BEG[0] ;
 wire \Tile_X2Y9_S1BEG[1] ;
 wire \Tile_X2Y9_S1BEG[2] ;
 wire \Tile_X2Y9_S1BEG[3] ;
 wire \Tile_X2Y9_S2BEG[0] ;
 wire \Tile_X2Y9_S2BEG[1] ;
 wire \Tile_X2Y9_S2BEG[2] ;
 wire \Tile_X2Y9_S2BEG[3] ;
 wire \Tile_X2Y9_S2BEG[4] ;
 wire \Tile_X2Y9_S2BEG[5] ;
 wire \Tile_X2Y9_S2BEG[6] ;
 wire \Tile_X2Y9_S2BEG[7] ;
 wire \Tile_X2Y9_S2BEGb[0] ;
 wire \Tile_X2Y9_S2BEGb[1] ;
 wire \Tile_X2Y9_S2BEGb[2] ;
 wire \Tile_X2Y9_S2BEGb[3] ;
 wire \Tile_X2Y9_S2BEGb[4] ;
 wire \Tile_X2Y9_S2BEGb[5] ;
 wire \Tile_X2Y9_S2BEGb[6] ;
 wire \Tile_X2Y9_S2BEGb[7] ;
 wire \Tile_X2Y9_S4BEG[0] ;
 wire \Tile_X2Y9_S4BEG[10] ;
 wire \Tile_X2Y9_S4BEG[11] ;
 wire \Tile_X2Y9_S4BEG[12] ;
 wire \Tile_X2Y9_S4BEG[13] ;
 wire \Tile_X2Y9_S4BEG[14] ;
 wire \Tile_X2Y9_S4BEG[15] ;
 wire \Tile_X2Y9_S4BEG[1] ;
 wire \Tile_X2Y9_S4BEG[2] ;
 wire \Tile_X2Y9_S4BEG[3] ;
 wire \Tile_X2Y9_S4BEG[4] ;
 wire \Tile_X2Y9_S4BEG[5] ;
 wire \Tile_X2Y9_S4BEG[6] ;
 wire \Tile_X2Y9_S4BEG[7] ;
 wire \Tile_X2Y9_S4BEG[8] ;
 wire \Tile_X2Y9_S4BEG[9] ;
 wire \Tile_X2Y9_SS4BEG[0] ;
 wire \Tile_X2Y9_SS4BEG[10] ;
 wire \Tile_X2Y9_SS4BEG[11] ;
 wire \Tile_X2Y9_SS4BEG[12] ;
 wire \Tile_X2Y9_SS4BEG[13] ;
 wire \Tile_X2Y9_SS4BEG[14] ;
 wire \Tile_X2Y9_SS4BEG[15] ;
 wire \Tile_X2Y9_SS4BEG[1] ;
 wire \Tile_X2Y9_SS4BEG[2] ;
 wire \Tile_X2Y9_SS4BEG[3] ;
 wire \Tile_X2Y9_SS4BEG[4] ;
 wire \Tile_X2Y9_SS4BEG[5] ;
 wire \Tile_X2Y9_SS4BEG[6] ;
 wire \Tile_X2Y9_SS4BEG[7] ;
 wire \Tile_X2Y9_SS4BEG[8] ;
 wire \Tile_X2Y9_SS4BEG[9] ;
 wire Tile_X2Y9_UserCLKo;
 wire \Tile_X2Y9_W1BEG[0] ;
 wire \Tile_X2Y9_W1BEG[1] ;
 wire \Tile_X2Y9_W1BEG[2] ;
 wire \Tile_X2Y9_W1BEG[3] ;
 wire \Tile_X2Y9_W2BEG[0] ;
 wire \Tile_X2Y9_W2BEG[1] ;
 wire \Tile_X2Y9_W2BEG[2] ;
 wire \Tile_X2Y9_W2BEG[3] ;
 wire \Tile_X2Y9_W2BEG[4] ;
 wire \Tile_X2Y9_W2BEG[5] ;
 wire \Tile_X2Y9_W2BEG[6] ;
 wire \Tile_X2Y9_W2BEG[7] ;
 wire \Tile_X2Y9_W2BEGb[0] ;
 wire \Tile_X2Y9_W2BEGb[1] ;
 wire \Tile_X2Y9_W2BEGb[2] ;
 wire \Tile_X2Y9_W2BEGb[3] ;
 wire \Tile_X2Y9_W2BEGb[4] ;
 wire \Tile_X2Y9_W2BEGb[5] ;
 wire \Tile_X2Y9_W2BEGb[6] ;
 wire \Tile_X2Y9_W2BEGb[7] ;
 wire \Tile_X2Y9_W6BEG[0] ;
 wire \Tile_X2Y9_W6BEG[10] ;
 wire \Tile_X2Y9_W6BEG[11] ;
 wire \Tile_X2Y9_W6BEG[1] ;
 wire \Tile_X2Y9_W6BEG[2] ;
 wire \Tile_X2Y9_W6BEG[3] ;
 wire \Tile_X2Y9_W6BEG[4] ;
 wire \Tile_X2Y9_W6BEG[5] ;
 wire \Tile_X2Y9_W6BEG[6] ;
 wire \Tile_X2Y9_W6BEG[7] ;
 wire \Tile_X2Y9_W6BEG[8] ;
 wire \Tile_X2Y9_W6BEG[9] ;
 wire \Tile_X2Y9_WW4BEG[0] ;
 wire \Tile_X2Y9_WW4BEG[10] ;
 wire \Tile_X2Y9_WW4BEG[11] ;
 wire \Tile_X2Y9_WW4BEG[12] ;
 wire \Tile_X2Y9_WW4BEG[13] ;
 wire \Tile_X2Y9_WW4BEG[14] ;
 wire \Tile_X2Y9_WW4BEG[15] ;
 wire \Tile_X2Y9_WW4BEG[1] ;
 wire \Tile_X2Y9_WW4BEG[2] ;
 wire \Tile_X2Y9_WW4BEG[3] ;
 wire \Tile_X2Y9_WW4BEG[4] ;
 wire \Tile_X2Y9_WW4BEG[5] ;
 wire \Tile_X2Y9_WW4BEG[6] ;
 wire \Tile_X2Y9_WW4BEG[7] ;
 wire \Tile_X2Y9_WW4BEG[8] ;
 wire \Tile_X2Y9_WW4BEG[9] ;
 wire \Tile_X3Y0_FrameData_O[0] ;
 wire \Tile_X3Y0_FrameData_O[10] ;
 wire \Tile_X3Y0_FrameData_O[11] ;
 wire \Tile_X3Y0_FrameData_O[12] ;
 wire \Tile_X3Y0_FrameData_O[13] ;
 wire \Tile_X3Y0_FrameData_O[14] ;
 wire \Tile_X3Y0_FrameData_O[15] ;
 wire \Tile_X3Y0_FrameData_O[16] ;
 wire \Tile_X3Y0_FrameData_O[17] ;
 wire \Tile_X3Y0_FrameData_O[18] ;
 wire \Tile_X3Y0_FrameData_O[19] ;
 wire \Tile_X3Y0_FrameData_O[1] ;
 wire \Tile_X3Y0_FrameData_O[20] ;
 wire \Tile_X3Y0_FrameData_O[21] ;
 wire \Tile_X3Y0_FrameData_O[22] ;
 wire \Tile_X3Y0_FrameData_O[23] ;
 wire \Tile_X3Y0_FrameData_O[24] ;
 wire \Tile_X3Y0_FrameData_O[25] ;
 wire \Tile_X3Y0_FrameData_O[26] ;
 wire \Tile_X3Y0_FrameData_O[27] ;
 wire \Tile_X3Y0_FrameData_O[28] ;
 wire \Tile_X3Y0_FrameData_O[29] ;
 wire \Tile_X3Y0_FrameData_O[2] ;
 wire \Tile_X3Y0_FrameData_O[30] ;
 wire \Tile_X3Y0_FrameData_O[31] ;
 wire \Tile_X3Y0_FrameData_O[3] ;
 wire \Tile_X3Y0_FrameData_O[4] ;
 wire \Tile_X3Y0_FrameData_O[5] ;
 wire \Tile_X3Y0_FrameData_O[6] ;
 wire \Tile_X3Y0_FrameData_O[7] ;
 wire \Tile_X3Y0_FrameData_O[8] ;
 wire \Tile_X3Y0_FrameData_O[9] ;
 wire \Tile_X3Y0_FrameStrobe_O[0] ;
 wire \Tile_X3Y0_FrameStrobe_O[10] ;
 wire \Tile_X3Y0_FrameStrobe_O[11] ;
 wire \Tile_X3Y0_FrameStrobe_O[12] ;
 wire \Tile_X3Y0_FrameStrobe_O[13] ;
 wire \Tile_X3Y0_FrameStrobe_O[14] ;
 wire \Tile_X3Y0_FrameStrobe_O[15] ;
 wire \Tile_X3Y0_FrameStrobe_O[16] ;
 wire \Tile_X3Y0_FrameStrobe_O[17] ;
 wire \Tile_X3Y0_FrameStrobe_O[18] ;
 wire \Tile_X3Y0_FrameStrobe_O[19] ;
 wire \Tile_X3Y0_FrameStrobe_O[1] ;
 wire \Tile_X3Y0_FrameStrobe_O[2] ;
 wire \Tile_X3Y0_FrameStrobe_O[3] ;
 wire \Tile_X3Y0_FrameStrobe_O[4] ;
 wire \Tile_X3Y0_FrameStrobe_O[5] ;
 wire \Tile_X3Y0_FrameStrobe_O[6] ;
 wire \Tile_X3Y0_FrameStrobe_O[7] ;
 wire \Tile_X3Y0_FrameStrobe_O[8] ;
 wire \Tile_X3Y0_FrameStrobe_O[9] ;
 wire \Tile_X3Y0_S1BEG[0] ;
 wire \Tile_X3Y0_S1BEG[1] ;
 wire \Tile_X3Y0_S1BEG[2] ;
 wire \Tile_X3Y0_S1BEG[3] ;
 wire \Tile_X3Y0_S2BEG[0] ;
 wire \Tile_X3Y0_S2BEG[1] ;
 wire \Tile_X3Y0_S2BEG[2] ;
 wire \Tile_X3Y0_S2BEG[3] ;
 wire \Tile_X3Y0_S2BEG[4] ;
 wire \Tile_X3Y0_S2BEG[5] ;
 wire \Tile_X3Y0_S2BEG[6] ;
 wire \Tile_X3Y0_S2BEG[7] ;
 wire \Tile_X3Y0_S2BEGb[0] ;
 wire \Tile_X3Y0_S2BEGb[1] ;
 wire \Tile_X3Y0_S2BEGb[2] ;
 wire \Tile_X3Y0_S2BEGb[3] ;
 wire \Tile_X3Y0_S2BEGb[4] ;
 wire \Tile_X3Y0_S2BEGb[5] ;
 wire \Tile_X3Y0_S2BEGb[6] ;
 wire \Tile_X3Y0_S2BEGb[7] ;
 wire \Tile_X3Y0_S4BEG[0] ;
 wire \Tile_X3Y0_S4BEG[10] ;
 wire \Tile_X3Y0_S4BEG[11] ;
 wire \Tile_X3Y0_S4BEG[12] ;
 wire \Tile_X3Y0_S4BEG[13] ;
 wire \Tile_X3Y0_S4BEG[14] ;
 wire \Tile_X3Y0_S4BEG[15] ;
 wire \Tile_X3Y0_S4BEG[1] ;
 wire \Tile_X3Y0_S4BEG[2] ;
 wire \Tile_X3Y0_S4BEG[3] ;
 wire \Tile_X3Y0_S4BEG[4] ;
 wire \Tile_X3Y0_S4BEG[5] ;
 wire \Tile_X3Y0_S4BEG[6] ;
 wire \Tile_X3Y0_S4BEG[7] ;
 wire \Tile_X3Y0_S4BEG[8] ;
 wire \Tile_X3Y0_S4BEG[9] ;
 wire \Tile_X3Y0_SS4BEG[0] ;
 wire \Tile_X3Y0_SS4BEG[10] ;
 wire \Tile_X3Y0_SS4BEG[11] ;
 wire \Tile_X3Y0_SS4BEG[12] ;
 wire \Tile_X3Y0_SS4BEG[13] ;
 wire \Tile_X3Y0_SS4BEG[14] ;
 wire \Tile_X3Y0_SS4BEG[15] ;
 wire \Tile_X3Y0_SS4BEG[1] ;
 wire \Tile_X3Y0_SS4BEG[2] ;
 wire \Tile_X3Y0_SS4BEG[3] ;
 wire \Tile_X3Y0_SS4BEG[4] ;
 wire \Tile_X3Y0_SS4BEG[5] ;
 wire \Tile_X3Y0_SS4BEG[6] ;
 wire \Tile_X3Y0_SS4BEG[7] ;
 wire \Tile_X3Y0_SS4BEG[8] ;
 wire \Tile_X3Y0_SS4BEG[9] ;
 wire Tile_X3Y0_UserCLKo;
 wire Tile_X3Y10_Co;
 wire \Tile_X3Y10_E1BEG[0] ;
 wire \Tile_X3Y10_E1BEG[1] ;
 wire \Tile_X3Y10_E1BEG[2] ;
 wire \Tile_X3Y10_E1BEG[3] ;
 wire \Tile_X3Y10_E2BEG[0] ;
 wire \Tile_X3Y10_E2BEG[1] ;
 wire \Tile_X3Y10_E2BEG[2] ;
 wire \Tile_X3Y10_E2BEG[3] ;
 wire \Tile_X3Y10_E2BEG[4] ;
 wire \Tile_X3Y10_E2BEG[5] ;
 wire \Tile_X3Y10_E2BEG[6] ;
 wire \Tile_X3Y10_E2BEG[7] ;
 wire \Tile_X3Y10_E2BEGb[0] ;
 wire \Tile_X3Y10_E2BEGb[1] ;
 wire \Tile_X3Y10_E2BEGb[2] ;
 wire \Tile_X3Y10_E2BEGb[3] ;
 wire \Tile_X3Y10_E2BEGb[4] ;
 wire \Tile_X3Y10_E2BEGb[5] ;
 wire \Tile_X3Y10_E2BEGb[6] ;
 wire \Tile_X3Y10_E2BEGb[7] ;
 wire \Tile_X3Y10_E6BEG[0] ;
 wire \Tile_X3Y10_E6BEG[10] ;
 wire \Tile_X3Y10_E6BEG[11] ;
 wire \Tile_X3Y10_E6BEG[1] ;
 wire \Tile_X3Y10_E6BEG[2] ;
 wire \Tile_X3Y10_E6BEG[3] ;
 wire \Tile_X3Y10_E6BEG[4] ;
 wire \Tile_X3Y10_E6BEG[5] ;
 wire \Tile_X3Y10_E6BEG[6] ;
 wire \Tile_X3Y10_E6BEG[7] ;
 wire \Tile_X3Y10_E6BEG[8] ;
 wire \Tile_X3Y10_E6BEG[9] ;
 wire \Tile_X3Y10_EE4BEG[0] ;
 wire \Tile_X3Y10_EE4BEG[10] ;
 wire \Tile_X3Y10_EE4BEG[11] ;
 wire \Tile_X3Y10_EE4BEG[12] ;
 wire \Tile_X3Y10_EE4BEG[13] ;
 wire \Tile_X3Y10_EE4BEG[14] ;
 wire \Tile_X3Y10_EE4BEG[15] ;
 wire \Tile_X3Y10_EE4BEG[1] ;
 wire \Tile_X3Y10_EE4BEG[2] ;
 wire \Tile_X3Y10_EE4BEG[3] ;
 wire \Tile_X3Y10_EE4BEG[4] ;
 wire \Tile_X3Y10_EE4BEG[5] ;
 wire \Tile_X3Y10_EE4BEG[6] ;
 wire \Tile_X3Y10_EE4BEG[7] ;
 wire \Tile_X3Y10_EE4BEG[8] ;
 wire \Tile_X3Y10_EE4BEG[9] ;
 wire \Tile_X3Y10_FrameData_O[0] ;
 wire \Tile_X3Y10_FrameData_O[10] ;
 wire \Tile_X3Y10_FrameData_O[11] ;
 wire \Tile_X3Y10_FrameData_O[12] ;
 wire \Tile_X3Y10_FrameData_O[13] ;
 wire \Tile_X3Y10_FrameData_O[14] ;
 wire \Tile_X3Y10_FrameData_O[15] ;
 wire \Tile_X3Y10_FrameData_O[16] ;
 wire \Tile_X3Y10_FrameData_O[17] ;
 wire \Tile_X3Y10_FrameData_O[18] ;
 wire \Tile_X3Y10_FrameData_O[19] ;
 wire \Tile_X3Y10_FrameData_O[1] ;
 wire \Tile_X3Y10_FrameData_O[20] ;
 wire \Tile_X3Y10_FrameData_O[21] ;
 wire \Tile_X3Y10_FrameData_O[22] ;
 wire \Tile_X3Y10_FrameData_O[23] ;
 wire \Tile_X3Y10_FrameData_O[24] ;
 wire \Tile_X3Y10_FrameData_O[25] ;
 wire \Tile_X3Y10_FrameData_O[26] ;
 wire \Tile_X3Y10_FrameData_O[27] ;
 wire \Tile_X3Y10_FrameData_O[28] ;
 wire \Tile_X3Y10_FrameData_O[29] ;
 wire \Tile_X3Y10_FrameData_O[2] ;
 wire \Tile_X3Y10_FrameData_O[30] ;
 wire \Tile_X3Y10_FrameData_O[31] ;
 wire \Tile_X3Y10_FrameData_O[3] ;
 wire \Tile_X3Y10_FrameData_O[4] ;
 wire \Tile_X3Y10_FrameData_O[5] ;
 wire \Tile_X3Y10_FrameData_O[6] ;
 wire \Tile_X3Y10_FrameData_O[7] ;
 wire \Tile_X3Y10_FrameData_O[8] ;
 wire \Tile_X3Y10_FrameData_O[9] ;
 wire \Tile_X3Y10_FrameStrobe_O[0] ;
 wire \Tile_X3Y10_FrameStrobe_O[10] ;
 wire \Tile_X3Y10_FrameStrobe_O[11] ;
 wire \Tile_X3Y10_FrameStrobe_O[12] ;
 wire \Tile_X3Y10_FrameStrobe_O[13] ;
 wire \Tile_X3Y10_FrameStrobe_O[14] ;
 wire \Tile_X3Y10_FrameStrobe_O[15] ;
 wire \Tile_X3Y10_FrameStrobe_O[16] ;
 wire \Tile_X3Y10_FrameStrobe_O[17] ;
 wire \Tile_X3Y10_FrameStrobe_O[18] ;
 wire \Tile_X3Y10_FrameStrobe_O[19] ;
 wire \Tile_X3Y10_FrameStrobe_O[1] ;
 wire \Tile_X3Y10_FrameStrobe_O[2] ;
 wire \Tile_X3Y10_FrameStrobe_O[3] ;
 wire \Tile_X3Y10_FrameStrobe_O[4] ;
 wire \Tile_X3Y10_FrameStrobe_O[5] ;
 wire \Tile_X3Y10_FrameStrobe_O[6] ;
 wire \Tile_X3Y10_FrameStrobe_O[7] ;
 wire \Tile_X3Y10_FrameStrobe_O[8] ;
 wire \Tile_X3Y10_FrameStrobe_O[9] ;
 wire \Tile_X3Y10_N1BEG[0] ;
 wire \Tile_X3Y10_N1BEG[1] ;
 wire \Tile_X3Y10_N1BEG[2] ;
 wire \Tile_X3Y10_N1BEG[3] ;
 wire \Tile_X3Y10_N2BEG[0] ;
 wire \Tile_X3Y10_N2BEG[1] ;
 wire \Tile_X3Y10_N2BEG[2] ;
 wire \Tile_X3Y10_N2BEG[3] ;
 wire \Tile_X3Y10_N2BEG[4] ;
 wire \Tile_X3Y10_N2BEG[5] ;
 wire \Tile_X3Y10_N2BEG[6] ;
 wire \Tile_X3Y10_N2BEG[7] ;
 wire \Tile_X3Y10_N2BEGb[0] ;
 wire \Tile_X3Y10_N2BEGb[1] ;
 wire \Tile_X3Y10_N2BEGb[2] ;
 wire \Tile_X3Y10_N2BEGb[3] ;
 wire \Tile_X3Y10_N2BEGb[4] ;
 wire \Tile_X3Y10_N2BEGb[5] ;
 wire \Tile_X3Y10_N2BEGb[6] ;
 wire \Tile_X3Y10_N2BEGb[7] ;
 wire \Tile_X3Y10_N4BEG[0] ;
 wire \Tile_X3Y10_N4BEG[10] ;
 wire \Tile_X3Y10_N4BEG[11] ;
 wire \Tile_X3Y10_N4BEG[12] ;
 wire \Tile_X3Y10_N4BEG[13] ;
 wire \Tile_X3Y10_N4BEG[14] ;
 wire \Tile_X3Y10_N4BEG[15] ;
 wire \Tile_X3Y10_N4BEG[1] ;
 wire \Tile_X3Y10_N4BEG[2] ;
 wire \Tile_X3Y10_N4BEG[3] ;
 wire \Tile_X3Y10_N4BEG[4] ;
 wire \Tile_X3Y10_N4BEG[5] ;
 wire \Tile_X3Y10_N4BEG[6] ;
 wire \Tile_X3Y10_N4BEG[7] ;
 wire \Tile_X3Y10_N4BEG[8] ;
 wire \Tile_X3Y10_N4BEG[9] ;
 wire \Tile_X3Y10_NN4BEG[0] ;
 wire \Tile_X3Y10_NN4BEG[10] ;
 wire \Tile_X3Y10_NN4BEG[11] ;
 wire \Tile_X3Y10_NN4BEG[12] ;
 wire \Tile_X3Y10_NN4BEG[13] ;
 wire \Tile_X3Y10_NN4BEG[14] ;
 wire \Tile_X3Y10_NN4BEG[15] ;
 wire \Tile_X3Y10_NN4BEG[1] ;
 wire \Tile_X3Y10_NN4BEG[2] ;
 wire \Tile_X3Y10_NN4BEG[3] ;
 wire \Tile_X3Y10_NN4BEG[4] ;
 wire \Tile_X3Y10_NN4BEG[5] ;
 wire \Tile_X3Y10_NN4BEG[6] ;
 wire \Tile_X3Y10_NN4BEG[7] ;
 wire \Tile_X3Y10_NN4BEG[8] ;
 wire \Tile_X3Y10_NN4BEG[9] ;
 wire \Tile_X3Y10_S1BEG[0] ;
 wire \Tile_X3Y10_S1BEG[1] ;
 wire \Tile_X3Y10_S1BEG[2] ;
 wire \Tile_X3Y10_S1BEG[3] ;
 wire \Tile_X3Y10_S2BEG[0] ;
 wire \Tile_X3Y10_S2BEG[1] ;
 wire \Tile_X3Y10_S2BEG[2] ;
 wire \Tile_X3Y10_S2BEG[3] ;
 wire \Tile_X3Y10_S2BEG[4] ;
 wire \Tile_X3Y10_S2BEG[5] ;
 wire \Tile_X3Y10_S2BEG[6] ;
 wire \Tile_X3Y10_S2BEG[7] ;
 wire \Tile_X3Y10_S2BEGb[0] ;
 wire \Tile_X3Y10_S2BEGb[1] ;
 wire \Tile_X3Y10_S2BEGb[2] ;
 wire \Tile_X3Y10_S2BEGb[3] ;
 wire \Tile_X3Y10_S2BEGb[4] ;
 wire \Tile_X3Y10_S2BEGb[5] ;
 wire \Tile_X3Y10_S2BEGb[6] ;
 wire \Tile_X3Y10_S2BEGb[7] ;
 wire \Tile_X3Y10_S4BEG[0] ;
 wire \Tile_X3Y10_S4BEG[10] ;
 wire \Tile_X3Y10_S4BEG[11] ;
 wire \Tile_X3Y10_S4BEG[12] ;
 wire \Tile_X3Y10_S4BEG[13] ;
 wire \Tile_X3Y10_S4BEG[14] ;
 wire \Tile_X3Y10_S4BEG[15] ;
 wire \Tile_X3Y10_S4BEG[1] ;
 wire \Tile_X3Y10_S4BEG[2] ;
 wire \Tile_X3Y10_S4BEG[3] ;
 wire \Tile_X3Y10_S4BEG[4] ;
 wire \Tile_X3Y10_S4BEG[5] ;
 wire \Tile_X3Y10_S4BEG[6] ;
 wire \Tile_X3Y10_S4BEG[7] ;
 wire \Tile_X3Y10_S4BEG[8] ;
 wire \Tile_X3Y10_S4BEG[9] ;
 wire \Tile_X3Y10_SS4BEG[0] ;
 wire \Tile_X3Y10_SS4BEG[10] ;
 wire \Tile_X3Y10_SS4BEG[11] ;
 wire \Tile_X3Y10_SS4BEG[12] ;
 wire \Tile_X3Y10_SS4BEG[13] ;
 wire \Tile_X3Y10_SS4BEG[14] ;
 wire \Tile_X3Y10_SS4BEG[15] ;
 wire \Tile_X3Y10_SS4BEG[1] ;
 wire \Tile_X3Y10_SS4BEG[2] ;
 wire \Tile_X3Y10_SS4BEG[3] ;
 wire \Tile_X3Y10_SS4BEG[4] ;
 wire \Tile_X3Y10_SS4BEG[5] ;
 wire \Tile_X3Y10_SS4BEG[6] ;
 wire \Tile_X3Y10_SS4BEG[7] ;
 wire \Tile_X3Y10_SS4BEG[8] ;
 wire \Tile_X3Y10_SS4BEG[9] ;
 wire Tile_X3Y10_UserCLKo;
 wire \Tile_X3Y10_W1BEG[0] ;
 wire \Tile_X3Y10_W1BEG[1] ;
 wire \Tile_X3Y10_W1BEG[2] ;
 wire \Tile_X3Y10_W1BEG[3] ;
 wire \Tile_X3Y10_W2BEG[0] ;
 wire \Tile_X3Y10_W2BEG[1] ;
 wire \Tile_X3Y10_W2BEG[2] ;
 wire \Tile_X3Y10_W2BEG[3] ;
 wire \Tile_X3Y10_W2BEG[4] ;
 wire \Tile_X3Y10_W2BEG[5] ;
 wire \Tile_X3Y10_W2BEG[6] ;
 wire \Tile_X3Y10_W2BEG[7] ;
 wire \Tile_X3Y10_W2BEGb[0] ;
 wire \Tile_X3Y10_W2BEGb[1] ;
 wire \Tile_X3Y10_W2BEGb[2] ;
 wire \Tile_X3Y10_W2BEGb[3] ;
 wire \Tile_X3Y10_W2BEGb[4] ;
 wire \Tile_X3Y10_W2BEGb[5] ;
 wire \Tile_X3Y10_W2BEGb[6] ;
 wire \Tile_X3Y10_W2BEGb[7] ;
 wire \Tile_X3Y10_W6BEG[0] ;
 wire \Tile_X3Y10_W6BEG[10] ;
 wire \Tile_X3Y10_W6BEG[11] ;
 wire \Tile_X3Y10_W6BEG[1] ;
 wire \Tile_X3Y10_W6BEG[2] ;
 wire \Tile_X3Y10_W6BEG[3] ;
 wire \Tile_X3Y10_W6BEG[4] ;
 wire \Tile_X3Y10_W6BEG[5] ;
 wire \Tile_X3Y10_W6BEG[6] ;
 wire \Tile_X3Y10_W6BEG[7] ;
 wire \Tile_X3Y10_W6BEG[8] ;
 wire \Tile_X3Y10_W6BEG[9] ;
 wire \Tile_X3Y10_WW4BEG[0] ;
 wire \Tile_X3Y10_WW4BEG[10] ;
 wire \Tile_X3Y10_WW4BEG[11] ;
 wire \Tile_X3Y10_WW4BEG[12] ;
 wire \Tile_X3Y10_WW4BEG[13] ;
 wire \Tile_X3Y10_WW4BEG[14] ;
 wire \Tile_X3Y10_WW4BEG[15] ;
 wire \Tile_X3Y10_WW4BEG[1] ;
 wire \Tile_X3Y10_WW4BEG[2] ;
 wire \Tile_X3Y10_WW4BEG[3] ;
 wire \Tile_X3Y10_WW4BEG[4] ;
 wire \Tile_X3Y10_WW4BEG[5] ;
 wire \Tile_X3Y10_WW4BEG[6] ;
 wire \Tile_X3Y10_WW4BEG[7] ;
 wire \Tile_X3Y10_WW4BEG[8] ;
 wire \Tile_X3Y10_WW4BEG[9] ;
 wire Tile_X3Y11_Co;
 wire \Tile_X3Y11_E1BEG[0] ;
 wire \Tile_X3Y11_E1BEG[1] ;
 wire \Tile_X3Y11_E1BEG[2] ;
 wire \Tile_X3Y11_E1BEG[3] ;
 wire \Tile_X3Y11_E2BEG[0] ;
 wire \Tile_X3Y11_E2BEG[1] ;
 wire \Tile_X3Y11_E2BEG[2] ;
 wire \Tile_X3Y11_E2BEG[3] ;
 wire \Tile_X3Y11_E2BEG[4] ;
 wire \Tile_X3Y11_E2BEG[5] ;
 wire \Tile_X3Y11_E2BEG[6] ;
 wire \Tile_X3Y11_E2BEG[7] ;
 wire \Tile_X3Y11_E2BEGb[0] ;
 wire \Tile_X3Y11_E2BEGb[1] ;
 wire \Tile_X3Y11_E2BEGb[2] ;
 wire \Tile_X3Y11_E2BEGb[3] ;
 wire \Tile_X3Y11_E2BEGb[4] ;
 wire \Tile_X3Y11_E2BEGb[5] ;
 wire \Tile_X3Y11_E2BEGb[6] ;
 wire \Tile_X3Y11_E2BEGb[7] ;
 wire \Tile_X3Y11_E6BEG[0] ;
 wire \Tile_X3Y11_E6BEG[10] ;
 wire \Tile_X3Y11_E6BEG[11] ;
 wire \Tile_X3Y11_E6BEG[1] ;
 wire \Tile_X3Y11_E6BEG[2] ;
 wire \Tile_X3Y11_E6BEG[3] ;
 wire \Tile_X3Y11_E6BEG[4] ;
 wire \Tile_X3Y11_E6BEG[5] ;
 wire \Tile_X3Y11_E6BEG[6] ;
 wire \Tile_X3Y11_E6BEG[7] ;
 wire \Tile_X3Y11_E6BEG[8] ;
 wire \Tile_X3Y11_E6BEG[9] ;
 wire \Tile_X3Y11_EE4BEG[0] ;
 wire \Tile_X3Y11_EE4BEG[10] ;
 wire \Tile_X3Y11_EE4BEG[11] ;
 wire \Tile_X3Y11_EE4BEG[12] ;
 wire \Tile_X3Y11_EE4BEG[13] ;
 wire \Tile_X3Y11_EE4BEG[14] ;
 wire \Tile_X3Y11_EE4BEG[15] ;
 wire \Tile_X3Y11_EE4BEG[1] ;
 wire \Tile_X3Y11_EE4BEG[2] ;
 wire \Tile_X3Y11_EE4BEG[3] ;
 wire \Tile_X3Y11_EE4BEG[4] ;
 wire \Tile_X3Y11_EE4BEG[5] ;
 wire \Tile_X3Y11_EE4BEG[6] ;
 wire \Tile_X3Y11_EE4BEG[7] ;
 wire \Tile_X3Y11_EE4BEG[8] ;
 wire \Tile_X3Y11_EE4BEG[9] ;
 wire \Tile_X3Y11_FrameData_O[0] ;
 wire \Tile_X3Y11_FrameData_O[10] ;
 wire \Tile_X3Y11_FrameData_O[11] ;
 wire \Tile_X3Y11_FrameData_O[12] ;
 wire \Tile_X3Y11_FrameData_O[13] ;
 wire \Tile_X3Y11_FrameData_O[14] ;
 wire \Tile_X3Y11_FrameData_O[15] ;
 wire \Tile_X3Y11_FrameData_O[16] ;
 wire \Tile_X3Y11_FrameData_O[17] ;
 wire \Tile_X3Y11_FrameData_O[18] ;
 wire \Tile_X3Y11_FrameData_O[19] ;
 wire \Tile_X3Y11_FrameData_O[1] ;
 wire \Tile_X3Y11_FrameData_O[20] ;
 wire \Tile_X3Y11_FrameData_O[21] ;
 wire \Tile_X3Y11_FrameData_O[22] ;
 wire \Tile_X3Y11_FrameData_O[23] ;
 wire \Tile_X3Y11_FrameData_O[24] ;
 wire \Tile_X3Y11_FrameData_O[25] ;
 wire \Tile_X3Y11_FrameData_O[26] ;
 wire \Tile_X3Y11_FrameData_O[27] ;
 wire \Tile_X3Y11_FrameData_O[28] ;
 wire \Tile_X3Y11_FrameData_O[29] ;
 wire \Tile_X3Y11_FrameData_O[2] ;
 wire \Tile_X3Y11_FrameData_O[30] ;
 wire \Tile_X3Y11_FrameData_O[31] ;
 wire \Tile_X3Y11_FrameData_O[3] ;
 wire \Tile_X3Y11_FrameData_O[4] ;
 wire \Tile_X3Y11_FrameData_O[5] ;
 wire \Tile_X3Y11_FrameData_O[6] ;
 wire \Tile_X3Y11_FrameData_O[7] ;
 wire \Tile_X3Y11_FrameData_O[8] ;
 wire \Tile_X3Y11_FrameData_O[9] ;
 wire \Tile_X3Y11_FrameStrobe_O[0] ;
 wire \Tile_X3Y11_FrameStrobe_O[10] ;
 wire \Tile_X3Y11_FrameStrobe_O[11] ;
 wire \Tile_X3Y11_FrameStrobe_O[12] ;
 wire \Tile_X3Y11_FrameStrobe_O[13] ;
 wire \Tile_X3Y11_FrameStrobe_O[14] ;
 wire \Tile_X3Y11_FrameStrobe_O[15] ;
 wire \Tile_X3Y11_FrameStrobe_O[16] ;
 wire \Tile_X3Y11_FrameStrobe_O[17] ;
 wire \Tile_X3Y11_FrameStrobe_O[18] ;
 wire \Tile_X3Y11_FrameStrobe_O[19] ;
 wire \Tile_X3Y11_FrameStrobe_O[1] ;
 wire \Tile_X3Y11_FrameStrobe_O[2] ;
 wire \Tile_X3Y11_FrameStrobe_O[3] ;
 wire \Tile_X3Y11_FrameStrobe_O[4] ;
 wire \Tile_X3Y11_FrameStrobe_O[5] ;
 wire \Tile_X3Y11_FrameStrobe_O[6] ;
 wire \Tile_X3Y11_FrameStrobe_O[7] ;
 wire \Tile_X3Y11_FrameStrobe_O[8] ;
 wire \Tile_X3Y11_FrameStrobe_O[9] ;
 wire \Tile_X3Y11_N1BEG[0] ;
 wire \Tile_X3Y11_N1BEG[1] ;
 wire \Tile_X3Y11_N1BEG[2] ;
 wire \Tile_X3Y11_N1BEG[3] ;
 wire \Tile_X3Y11_N2BEG[0] ;
 wire \Tile_X3Y11_N2BEG[1] ;
 wire \Tile_X3Y11_N2BEG[2] ;
 wire \Tile_X3Y11_N2BEG[3] ;
 wire \Tile_X3Y11_N2BEG[4] ;
 wire \Tile_X3Y11_N2BEG[5] ;
 wire \Tile_X3Y11_N2BEG[6] ;
 wire \Tile_X3Y11_N2BEG[7] ;
 wire \Tile_X3Y11_N2BEGb[0] ;
 wire \Tile_X3Y11_N2BEGb[1] ;
 wire \Tile_X3Y11_N2BEGb[2] ;
 wire \Tile_X3Y11_N2BEGb[3] ;
 wire \Tile_X3Y11_N2BEGb[4] ;
 wire \Tile_X3Y11_N2BEGb[5] ;
 wire \Tile_X3Y11_N2BEGb[6] ;
 wire \Tile_X3Y11_N2BEGb[7] ;
 wire \Tile_X3Y11_N4BEG[0] ;
 wire \Tile_X3Y11_N4BEG[10] ;
 wire \Tile_X3Y11_N4BEG[11] ;
 wire \Tile_X3Y11_N4BEG[12] ;
 wire \Tile_X3Y11_N4BEG[13] ;
 wire \Tile_X3Y11_N4BEG[14] ;
 wire \Tile_X3Y11_N4BEG[15] ;
 wire \Tile_X3Y11_N4BEG[1] ;
 wire \Tile_X3Y11_N4BEG[2] ;
 wire \Tile_X3Y11_N4BEG[3] ;
 wire \Tile_X3Y11_N4BEG[4] ;
 wire \Tile_X3Y11_N4BEG[5] ;
 wire \Tile_X3Y11_N4BEG[6] ;
 wire \Tile_X3Y11_N4BEG[7] ;
 wire \Tile_X3Y11_N4BEG[8] ;
 wire \Tile_X3Y11_N4BEG[9] ;
 wire \Tile_X3Y11_NN4BEG[0] ;
 wire \Tile_X3Y11_NN4BEG[10] ;
 wire \Tile_X3Y11_NN4BEG[11] ;
 wire \Tile_X3Y11_NN4BEG[12] ;
 wire \Tile_X3Y11_NN4BEG[13] ;
 wire \Tile_X3Y11_NN4BEG[14] ;
 wire \Tile_X3Y11_NN4BEG[15] ;
 wire \Tile_X3Y11_NN4BEG[1] ;
 wire \Tile_X3Y11_NN4BEG[2] ;
 wire \Tile_X3Y11_NN4BEG[3] ;
 wire \Tile_X3Y11_NN4BEG[4] ;
 wire \Tile_X3Y11_NN4BEG[5] ;
 wire \Tile_X3Y11_NN4BEG[6] ;
 wire \Tile_X3Y11_NN4BEG[7] ;
 wire \Tile_X3Y11_NN4BEG[8] ;
 wire \Tile_X3Y11_NN4BEG[9] ;
 wire \Tile_X3Y11_S1BEG[0] ;
 wire \Tile_X3Y11_S1BEG[1] ;
 wire \Tile_X3Y11_S1BEG[2] ;
 wire \Tile_X3Y11_S1BEG[3] ;
 wire \Tile_X3Y11_S2BEG[0] ;
 wire \Tile_X3Y11_S2BEG[1] ;
 wire \Tile_X3Y11_S2BEG[2] ;
 wire \Tile_X3Y11_S2BEG[3] ;
 wire \Tile_X3Y11_S2BEG[4] ;
 wire \Tile_X3Y11_S2BEG[5] ;
 wire \Tile_X3Y11_S2BEG[6] ;
 wire \Tile_X3Y11_S2BEG[7] ;
 wire \Tile_X3Y11_S2BEGb[0] ;
 wire \Tile_X3Y11_S2BEGb[1] ;
 wire \Tile_X3Y11_S2BEGb[2] ;
 wire \Tile_X3Y11_S2BEGb[3] ;
 wire \Tile_X3Y11_S2BEGb[4] ;
 wire \Tile_X3Y11_S2BEGb[5] ;
 wire \Tile_X3Y11_S2BEGb[6] ;
 wire \Tile_X3Y11_S2BEGb[7] ;
 wire \Tile_X3Y11_S4BEG[0] ;
 wire \Tile_X3Y11_S4BEG[10] ;
 wire \Tile_X3Y11_S4BEG[11] ;
 wire \Tile_X3Y11_S4BEG[12] ;
 wire \Tile_X3Y11_S4BEG[13] ;
 wire \Tile_X3Y11_S4BEG[14] ;
 wire \Tile_X3Y11_S4BEG[15] ;
 wire \Tile_X3Y11_S4BEG[1] ;
 wire \Tile_X3Y11_S4BEG[2] ;
 wire \Tile_X3Y11_S4BEG[3] ;
 wire \Tile_X3Y11_S4BEG[4] ;
 wire \Tile_X3Y11_S4BEG[5] ;
 wire \Tile_X3Y11_S4BEG[6] ;
 wire \Tile_X3Y11_S4BEG[7] ;
 wire \Tile_X3Y11_S4BEG[8] ;
 wire \Tile_X3Y11_S4BEG[9] ;
 wire \Tile_X3Y11_SS4BEG[0] ;
 wire \Tile_X3Y11_SS4BEG[10] ;
 wire \Tile_X3Y11_SS4BEG[11] ;
 wire \Tile_X3Y11_SS4BEG[12] ;
 wire \Tile_X3Y11_SS4BEG[13] ;
 wire \Tile_X3Y11_SS4BEG[14] ;
 wire \Tile_X3Y11_SS4BEG[15] ;
 wire \Tile_X3Y11_SS4BEG[1] ;
 wire \Tile_X3Y11_SS4BEG[2] ;
 wire \Tile_X3Y11_SS4BEG[3] ;
 wire \Tile_X3Y11_SS4BEG[4] ;
 wire \Tile_X3Y11_SS4BEG[5] ;
 wire \Tile_X3Y11_SS4BEG[6] ;
 wire \Tile_X3Y11_SS4BEG[7] ;
 wire \Tile_X3Y11_SS4BEG[8] ;
 wire \Tile_X3Y11_SS4BEG[9] ;
 wire Tile_X3Y11_UserCLKo;
 wire \Tile_X3Y11_W1BEG[0] ;
 wire \Tile_X3Y11_W1BEG[1] ;
 wire \Tile_X3Y11_W1BEG[2] ;
 wire \Tile_X3Y11_W1BEG[3] ;
 wire \Tile_X3Y11_W2BEG[0] ;
 wire \Tile_X3Y11_W2BEG[1] ;
 wire \Tile_X3Y11_W2BEG[2] ;
 wire \Tile_X3Y11_W2BEG[3] ;
 wire \Tile_X3Y11_W2BEG[4] ;
 wire \Tile_X3Y11_W2BEG[5] ;
 wire \Tile_X3Y11_W2BEG[6] ;
 wire \Tile_X3Y11_W2BEG[7] ;
 wire \Tile_X3Y11_W2BEGb[0] ;
 wire \Tile_X3Y11_W2BEGb[1] ;
 wire \Tile_X3Y11_W2BEGb[2] ;
 wire \Tile_X3Y11_W2BEGb[3] ;
 wire \Tile_X3Y11_W2BEGb[4] ;
 wire \Tile_X3Y11_W2BEGb[5] ;
 wire \Tile_X3Y11_W2BEGb[6] ;
 wire \Tile_X3Y11_W2BEGb[7] ;
 wire \Tile_X3Y11_W6BEG[0] ;
 wire \Tile_X3Y11_W6BEG[10] ;
 wire \Tile_X3Y11_W6BEG[11] ;
 wire \Tile_X3Y11_W6BEG[1] ;
 wire \Tile_X3Y11_W6BEG[2] ;
 wire \Tile_X3Y11_W6BEG[3] ;
 wire \Tile_X3Y11_W6BEG[4] ;
 wire \Tile_X3Y11_W6BEG[5] ;
 wire \Tile_X3Y11_W6BEG[6] ;
 wire \Tile_X3Y11_W6BEG[7] ;
 wire \Tile_X3Y11_W6BEG[8] ;
 wire \Tile_X3Y11_W6BEG[9] ;
 wire \Tile_X3Y11_WW4BEG[0] ;
 wire \Tile_X3Y11_WW4BEG[10] ;
 wire \Tile_X3Y11_WW4BEG[11] ;
 wire \Tile_X3Y11_WW4BEG[12] ;
 wire \Tile_X3Y11_WW4BEG[13] ;
 wire \Tile_X3Y11_WW4BEG[14] ;
 wire \Tile_X3Y11_WW4BEG[15] ;
 wire \Tile_X3Y11_WW4BEG[1] ;
 wire \Tile_X3Y11_WW4BEG[2] ;
 wire \Tile_X3Y11_WW4BEG[3] ;
 wire \Tile_X3Y11_WW4BEG[4] ;
 wire \Tile_X3Y11_WW4BEG[5] ;
 wire \Tile_X3Y11_WW4BEG[6] ;
 wire \Tile_X3Y11_WW4BEG[7] ;
 wire \Tile_X3Y11_WW4BEG[8] ;
 wire \Tile_X3Y11_WW4BEG[9] ;
 wire Tile_X3Y12_Co;
 wire \Tile_X3Y12_E1BEG[0] ;
 wire \Tile_X3Y12_E1BEG[1] ;
 wire \Tile_X3Y12_E1BEG[2] ;
 wire \Tile_X3Y12_E1BEG[3] ;
 wire \Tile_X3Y12_E2BEG[0] ;
 wire \Tile_X3Y12_E2BEG[1] ;
 wire \Tile_X3Y12_E2BEG[2] ;
 wire \Tile_X3Y12_E2BEG[3] ;
 wire \Tile_X3Y12_E2BEG[4] ;
 wire \Tile_X3Y12_E2BEG[5] ;
 wire \Tile_X3Y12_E2BEG[6] ;
 wire \Tile_X3Y12_E2BEG[7] ;
 wire \Tile_X3Y12_E2BEGb[0] ;
 wire \Tile_X3Y12_E2BEGb[1] ;
 wire \Tile_X3Y12_E2BEGb[2] ;
 wire \Tile_X3Y12_E2BEGb[3] ;
 wire \Tile_X3Y12_E2BEGb[4] ;
 wire \Tile_X3Y12_E2BEGb[5] ;
 wire \Tile_X3Y12_E2BEGb[6] ;
 wire \Tile_X3Y12_E2BEGb[7] ;
 wire \Tile_X3Y12_E6BEG[0] ;
 wire \Tile_X3Y12_E6BEG[10] ;
 wire \Tile_X3Y12_E6BEG[11] ;
 wire \Tile_X3Y12_E6BEG[1] ;
 wire \Tile_X3Y12_E6BEG[2] ;
 wire \Tile_X3Y12_E6BEG[3] ;
 wire \Tile_X3Y12_E6BEG[4] ;
 wire \Tile_X3Y12_E6BEG[5] ;
 wire \Tile_X3Y12_E6BEG[6] ;
 wire \Tile_X3Y12_E6BEG[7] ;
 wire \Tile_X3Y12_E6BEG[8] ;
 wire \Tile_X3Y12_E6BEG[9] ;
 wire \Tile_X3Y12_EE4BEG[0] ;
 wire \Tile_X3Y12_EE4BEG[10] ;
 wire \Tile_X3Y12_EE4BEG[11] ;
 wire \Tile_X3Y12_EE4BEG[12] ;
 wire \Tile_X3Y12_EE4BEG[13] ;
 wire \Tile_X3Y12_EE4BEG[14] ;
 wire \Tile_X3Y12_EE4BEG[15] ;
 wire \Tile_X3Y12_EE4BEG[1] ;
 wire \Tile_X3Y12_EE4BEG[2] ;
 wire \Tile_X3Y12_EE4BEG[3] ;
 wire \Tile_X3Y12_EE4BEG[4] ;
 wire \Tile_X3Y12_EE4BEG[5] ;
 wire \Tile_X3Y12_EE4BEG[6] ;
 wire \Tile_X3Y12_EE4BEG[7] ;
 wire \Tile_X3Y12_EE4BEG[8] ;
 wire \Tile_X3Y12_EE4BEG[9] ;
 wire \Tile_X3Y12_FrameData_O[0] ;
 wire \Tile_X3Y12_FrameData_O[10] ;
 wire \Tile_X3Y12_FrameData_O[11] ;
 wire \Tile_X3Y12_FrameData_O[12] ;
 wire \Tile_X3Y12_FrameData_O[13] ;
 wire \Tile_X3Y12_FrameData_O[14] ;
 wire \Tile_X3Y12_FrameData_O[15] ;
 wire \Tile_X3Y12_FrameData_O[16] ;
 wire \Tile_X3Y12_FrameData_O[17] ;
 wire \Tile_X3Y12_FrameData_O[18] ;
 wire \Tile_X3Y12_FrameData_O[19] ;
 wire \Tile_X3Y12_FrameData_O[1] ;
 wire \Tile_X3Y12_FrameData_O[20] ;
 wire \Tile_X3Y12_FrameData_O[21] ;
 wire \Tile_X3Y12_FrameData_O[22] ;
 wire \Tile_X3Y12_FrameData_O[23] ;
 wire \Tile_X3Y12_FrameData_O[24] ;
 wire \Tile_X3Y12_FrameData_O[25] ;
 wire \Tile_X3Y12_FrameData_O[26] ;
 wire \Tile_X3Y12_FrameData_O[27] ;
 wire \Tile_X3Y12_FrameData_O[28] ;
 wire \Tile_X3Y12_FrameData_O[29] ;
 wire \Tile_X3Y12_FrameData_O[2] ;
 wire \Tile_X3Y12_FrameData_O[30] ;
 wire \Tile_X3Y12_FrameData_O[31] ;
 wire \Tile_X3Y12_FrameData_O[3] ;
 wire \Tile_X3Y12_FrameData_O[4] ;
 wire \Tile_X3Y12_FrameData_O[5] ;
 wire \Tile_X3Y12_FrameData_O[6] ;
 wire \Tile_X3Y12_FrameData_O[7] ;
 wire \Tile_X3Y12_FrameData_O[8] ;
 wire \Tile_X3Y12_FrameData_O[9] ;
 wire \Tile_X3Y12_FrameStrobe_O[0] ;
 wire \Tile_X3Y12_FrameStrobe_O[10] ;
 wire \Tile_X3Y12_FrameStrobe_O[11] ;
 wire \Tile_X3Y12_FrameStrobe_O[12] ;
 wire \Tile_X3Y12_FrameStrobe_O[13] ;
 wire \Tile_X3Y12_FrameStrobe_O[14] ;
 wire \Tile_X3Y12_FrameStrobe_O[15] ;
 wire \Tile_X3Y12_FrameStrobe_O[16] ;
 wire \Tile_X3Y12_FrameStrobe_O[17] ;
 wire \Tile_X3Y12_FrameStrobe_O[18] ;
 wire \Tile_X3Y12_FrameStrobe_O[19] ;
 wire \Tile_X3Y12_FrameStrobe_O[1] ;
 wire \Tile_X3Y12_FrameStrobe_O[2] ;
 wire \Tile_X3Y12_FrameStrobe_O[3] ;
 wire \Tile_X3Y12_FrameStrobe_O[4] ;
 wire \Tile_X3Y12_FrameStrobe_O[5] ;
 wire \Tile_X3Y12_FrameStrobe_O[6] ;
 wire \Tile_X3Y12_FrameStrobe_O[7] ;
 wire \Tile_X3Y12_FrameStrobe_O[8] ;
 wire \Tile_X3Y12_FrameStrobe_O[9] ;
 wire \Tile_X3Y12_N1BEG[0] ;
 wire \Tile_X3Y12_N1BEG[1] ;
 wire \Tile_X3Y12_N1BEG[2] ;
 wire \Tile_X3Y12_N1BEG[3] ;
 wire \Tile_X3Y12_N2BEG[0] ;
 wire \Tile_X3Y12_N2BEG[1] ;
 wire \Tile_X3Y12_N2BEG[2] ;
 wire \Tile_X3Y12_N2BEG[3] ;
 wire \Tile_X3Y12_N2BEG[4] ;
 wire \Tile_X3Y12_N2BEG[5] ;
 wire \Tile_X3Y12_N2BEG[6] ;
 wire \Tile_X3Y12_N2BEG[7] ;
 wire \Tile_X3Y12_N2BEGb[0] ;
 wire \Tile_X3Y12_N2BEGb[1] ;
 wire \Tile_X3Y12_N2BEGb[2] ;
 wire \Tile_X3Y12_N2BEGb[3] ;
 wire \Tile_X3Y12_N2BEGb[4] ;
 wire \Tile_X3Y12_N2BEGb[5] ;
 wire \Tile_X3Y12_N2BEGb[6] ;
 wire \Tile_X3Y12_N2BEGb[7] ;
 wire \Tile_X3Y12_N4BEG[0] ;
 wire \Tile_X3Y12_N4BEG[10] ;
 wire \Tile_X3Y12_N4BEG[11] ;
 wire \Tile_X3Y12_N4BEG[12] ;
 wire \Tile_X3Y12_N4BEG[13] ;
 wire \Tile_X3Y12_N4BEG[14] ;
 wire \Tile_X3Y12_N4BEG[15] ;
 wire \Tile_X3Y12_N4BEG[1] ;
 wire \Tile_X3Y12_N4BEG[2] ;
 wire \Tile_X3Y12_N4BEG[3] ;
 wire \Tile_X3Y12_N4BEG[4] ;
 wire \Tile_X3Y12_N4BEG[5] ;
 wire \Tile_X3Y12_N4BEG[6] ;
 wire \Tile_X3Y12_N4BEG[7] ;
 wire \Tile_X3Y12_N4BEG[8] ;
 wire \Tile_X3Y12_N4BEG[9] ;
 wire \Tile_X3Y12_NN4BEG[0] ;
 wire \Tile_X3Y12_NN4BEG[10] ;
 wire \Tile_X3Y12_NN4BEG[11] ;
 wire \Tile_X3Y12_NN4BEG[12] ;
 wire \Tile_X3Y12_NN4BEG[13] ;
 wire \Tile_X3Y12_NN4BEG[14] ;
 wire \Tile_X3Y12_NN4BEG[15] ;
 wire \Tile_X3Y12_NN4BEG[1] ;
 wire \Tile_X3Y12_NN4BEG[2] ;
 wire \Tile_X3Y12_NN4BEG[3] ;
 wire \Tile_X3Y12_NN4BEG[4] ;
 wire \Tile_X3Y12_NN4BEG[5] ;
 wire \Tile_X3Y12_NN4BEG[6] ;
 wire \Tile_X3Y12_NN4BEG[7] ;
 wire \Tile_X3Y12_NN4BEG[8] ;
 wire \Tile_X3Y12_NN4BEG[9] ;
 wire \Tile_X3Y12_S1BEG[0] ;
 wire \Tile_X3Y12_S1BEG[1] ;
 wire \Tile_X3Y12_S1BEG[2] ;
 wire \Tile_X3Y12_S1BEG[3] ;
 wire \Tile_X3Y12_S2BEG[0] ;
 wire \Tile_X3Y12_S2BEG[1] ;
 wire \Tile_X3Y12_S2BEG[2] ;
 wire \Tile_X3Y12_S2BEG[3] ;
 wire \Tile_X3Y12_S2BEG[4] ;
 wire \Tile_X3Y12_S2BEG[5] ;
 wire \Tile_X3Y12_S2BEG[6] ;
 wire \Tile_X3Y12_S2BEG[7] ;
 wire \Tile_X3Y12_S2BEGb[0] ;
 wire \Tile_X3Y12_S2BEGb[1] ;
 wire \Tile_X3Y12_S2BEGb[2] ;
 wire \Tile_X3Y12_S2BEGb[3] ;
 wire \Tile_X3Y12_S2BEGb[4] ;
 wire \Tile_X3Y12_S2BEGb[5] ;
 wire \Tile_X3Y12_S2BEGb[6] ;
 wire \Tile_X3Y12_S2BEGb[7] ;
 wire \Tile_X3Y12_S4BEG[0] ;
 wire \Tile_X3Y12_S4BEG[10] ;
 wire \Tile_X3Y12_S4BEG[11] ;
 wire \Tile_X3Y12_S4BEG[12] ;
 wire \Tile_X3Y12_S4BEG[13] ;
 wire \Tile_X3Y12_S4BEG[14] ;
 wire \Tile_X3Y12_S4BEG[15] ;
 wire \Tile_X3Y12_S4BEG[1] ;
 wire \Tile_X3Y12_S4BEG[2] ;
 wire \Tile_X3Y12_S4BEG[3] ;
 wire \Tile_X3Y12_S4BEG[4] ;
 wire \Tile_X3Y12_S4BEG[5] ;
 wire \Tile_X3Y12_S4BEG[6] ;
 wire \Tile_X3Y12_S4BEG[7] ;
 wire \Tile_X3Y12_S4BEG[8] ;
 wire \Tile_X3Y12_S4BEG[9] ;
 wire \Tile_X3Y12_SS4BEG[0] ;
 wire \Tile_X3Y12_SS4BEG[10] ;
 wire \Tile_X3Y12_SS4BEG[11] ;
 wire \Tile_X3Y12_SS4BEG[12] ;
 wire \Tile_X3Y12_SS4BEG[13] ;
 wire \Tile_X3Y12_SS4BEG[14] ;
 wire \Tile_X3Y12_SS4BEG[15] ;
 wire \Tile_X3Y12_SS4BEG[1] ;
 wire \Tile_X3Y12_SS4BEG[2] ;
 wire \Tile_X3Y12_SS4BEG[3] ;
 wire \Tile_X3Y12_SS4BEG[4] ;
 wire \Tile_X3Y12_SS4BEG[5] ;
 wire \Tile_X3Y12_SS4BEG[6] ;
 wire \Tile_X3Y12_SS4BEG[7] ;
 wire \Tile_X3Y12_SS4BEG[8] ;
 wire \Tile_X3Y12_SS4BEG[9] ;
 wire Tile_X3Y12_UserCLKo;
 wire \Tile_X3Y12_W1BEG[0] ;
 wire \Tile_X3Y12_W1BEG[1] ;
 wire \Tile_X3Y12_W1BEG[2] ;
 wire \Tile_X3Y12_W1BEG[3] ;
 wire \Tile_X3Y12_W2BEG[0] ;
 wire \Tile_X3Y12_W2BEG[1] ;
 wire \Tile_X3Y12_W2BEG[2] ;
 wire \Tile_X3Y12_W2BEG[3] ;
 wire \Tile_X3Y12_W2BEG[4] ;
 wire \Tile_X3Y12_W2BEG[5] ;
 wire \Tile_X3Y12_W2BEG[6] ;
 wire \Tile_X3Y12_W2BEG[7] ;
 wire \Tile_X3Y12_W2BEGb[0] ;
 wire \Tile_X3Y12_W2BEGb[1] ;
 wire \Tile_X3Y12_W2BEGb[2] ;
 wire \Tile_X3Y12_W2BEGb[3] ;
 wire \Tile_X3Y12_W2BEGb[4] ;
 wire \Tile_X3Y12_W2BEGb[5] ;
 wire \Tile_X3Y12_W2BEGb[6] ;
 wire \Tile_X3Y12_W2BEGb[7] ;
 wire \Tile_X3Y12_W6BEG[0] ;
 wire \Tile_X3Y12_W6BEG[10] ;
 wire \Tile_X3Y12_W6BEG[11] ;
 wire \Tile_X3Y12_W6BEG[1] ;
 wire \Tile_X3Y12_W6BEG[2] ;
 wire \Tile_X3Y12_W6BEG[3] ;
 wire \Tile_X3Y12_W6BEG[4] ;
 wire \Tile_X3Y12_W6BEG[5] ;
 wire \Tile_X3Y12_W6BEG[6] ;
 wire \Tile_X3Y12_W6BEG[7] ;
 wire \Tile_X3Y12_W6BEG[8] ;
 wire \Tile_X3Y12_W6BEG[9] ;
 wire \Tile_X3Y12_WW4BEG[0] ;
 wire \Tile_X3Y12_WW4BEG[10] ;
 wire \Tile_X3Y12_WW4BEG[11] ;
 wire \Tile_X3Y12_WW4BEG[12] ;
 wire \Tile_X3Y12_WW4BEG[13] ;
 wire \Tile_X3Y12_WW4BEG[14] ;
 wire \Tile_X3Y12_WW4BEG[15] ;
 wire \Tile_X3Y12_WW4BEG[1] ;
 wire \Tile_X3Y12_WW4BEG[2] ;
 wire \Tile_X3Y12_WW4BEG[3] ;
 wire \Tile_X3Y12_WW4BEG[4] ;
 wire \Tile_X3Y12_WW4BEG[5] ;
 wire \Tile_X3Y12_WW4BEG[6] ;
 wire \Tile_X3Y12_WW4BEG[7] ;
 wire \Tile_X3Y12_WW4BEG[8] ;
 wire \Tile_X3Y12_WW4BEG[9] ;
 wire Tile_X3Y13_Co;
 wire \Tile_X3Y13_E1BEG[0] ;
 wire \Tile_X3Y13_E1BEG[1] ;
 wire \Tile_X3Y13_E1BEG[2] ;
 wire \Tile_X3Y13_E1BEG[3] ;
 wire \Tile_X3Y13_E2BEG[0] ;
 wire \Tile_X3Y13_E2BEG[1] ;
 wire \Tile_X3Y13_E2BEG[2] ;
 wire \Tile_X3Y13_E2BEG[3] ;
 wire \Tile_X3Y13_E2BEG[4] ;
 wire \Tile_X3Y13_E2BEG[5] ;
 wire \Tile_X3Y13_E2BEG[6] ;
 wire \Tile_X3Y13_E2BEG[7] ;
 wire \Tile_X3Y13_E2BEGb[0] ;
 wire \Tile_X3Y13_E2BEGb[1] ;
 wire \Tile_X3Y13_E2BEGb[2] ;
 wire \Tile_X3Y13_E2BEGb[3] ;
 wire \Tile_X3Y13_E2BEGb[4] ;
 wire \Tile_X3Y13_E2BEGb[5] ;
 wire \Tile_X3Y13_E2BEGb[6] ;
 wire \Tile_X3Y13_E2BEGb[7] ;
 wire \Tile_X3Y13_E6BEG[0] ;
 wire \Tile_X3Y13_E6BEG[10] ;
 wire \Tile_X3Y13_E6BEG[11] ;
 wire \Tile_X3Y13_E6BEG[1] ;
 wire \Tile_X3Y13_E6BEG[2] ;
 wire \Tile_X3Y13_E6BEG[3] ;
 wire \Tile_X3Y13_E6BEG[4] ;
 wire \Tile_X3Y13_E6BEG[5] ;
 wire \Tile_X3Y13_E6BEG[6] ;
 wire \Tile_X3Y13_E6BEG[7] ;
 wire \Tile_X3Y13_E6BEG[8] ;
 wire \Tile_X3Y13_E6BEG[9] ;
 wire \Tile_X3Y13_EE4BEG[0] ;
 wire \Tile_X3Y13_EE4BEG[10] ;
 wire \Tile_X3Y13_EE4BEG[11] ;
 wire \Tile_X3Y13_EE4BEG[12] ;
 wire \Tile_X3Y13_EE4BEG[13] ;
 wire \Tile_X3Y13_EE4BEG[14] ;
 wire \Tile_X3Y13_EE4BEG[15] ;
 wire \Tile_X3Y13_EE4BEG[1] ;
 wire \Tile_X3Y13_EE4BEG[2] ;
 wire \Tile_X3Y13_EE4BEG[3] ;
 wire \Tile_X3Y13_EE4BEG[4] ;
 wire \Tile_X3Y13_EE4BEG[5] ;
 wire \Tile_X3Y13_EE4BEG[6] ;
 wire \Tile_X3Y13_EE4BEG[7] ;
 wire \Tile_X3Y13_EE4BEG[8] ;
 wire \Tile_X3Y13_EE4BEG[9] ;
 wire \Tile_X3Y13_FrameData_O[0] ;
 wire \Tile_X3Y13_FrameData_O[10] ;
 wire \Tile_X3Y13_FrameData_O[11] ;
 wire \Tile_X3Y13_FrameData_O[12] ;
 wire \Tile_X3Y13_FrameData_O[13] ;
 wire \Tile_X3Y13_FrameData_O[14] ;
 wire \Tile_X3Y13_FrameData_O[15] ;
 wire \Tile_X3Y13_FrameData_O[16] ;
 wire \Tile_X3Y13_FrameData_O[17] ;
 wire \Tile_X3Y13_FrameData_O[18] ;
 wire \Tile_X3Y13_FrameData_O[19] ;
 wire \Tile_X3Y13_FrameData_O[1] ;
 wire \Tile_X3Y13_FrameData_O[20] ;
 wire \Tile_X3Y13_FrameData_O[21] ;
 wire \Tile_X3Y13_FrameData_O[22] ;
 wire \Tile_X3Y13_FrameData_O[23] ;
 wire \Tile_X3Y13_FrameData_O[24] ;
 wire \Tile_X3Y13_FrameData_O[25] ;
 wire \Tile_X3Y13_FrameData_O[26] ;
 wire \Tile_X3Y13_FrameData_O[27] ;
 wire \Tile_X3Y13_FrameData_O[28] ;
 wire \Tile_X3Y13_FrameData_O[29] ;
 wire \Tile_X3Y13_FrameData_O[2] ;
 wire \Tile_X3Y13_FrameData_O[30] ;
 wire \Tile_X3Y13_FrameData_O[31] ;
 wire \Tile_X3Y13_FrameData_O[3] ;
 wire \Tile_X3Y13_FrameData_O[4] ;
 wire \Tile_X3Y13_FrameData_O[5] ;
 wire \Tile_X3Y13_FrameData_O[6] ;
 wire \Tile_X3Y13_FrameData_O[7] ;
 wire \Tile_X3Y13_FrameData_O[8] ;
 wire \Tile_X3Y13_FrameData_O[9] ;
 wire \Tile_X3Y13_FrameStrobe_O[0] ;
 wire \Tile_X3Y13_FrameStrobe_O[10] ;
 wire \Tile_X3Y13_FrameStrobe_O[11] ;
 wire \Tile_X3Y13_FrameStrobe_O[12] ;
 wire \Tile_X3Y13_FrameStrobe_O[13] ;
 wire \Tile_X3Y13_FrameStrobe_O[14] ;
 wire \Tile_X3Y13_FrameStrobe_O[15] ;
 wire \Tile_X3Y13_FrameStrobe_O[16] ;
 wire \Tile_X3Y13_FrameStrobe_O[17] ;
 wire \Tile_X3Y13_FrameStrobe_O[18] ;
 wire \Tile_X3Y13_FrameStrobe_O[19] ;
 wire \Tile_X3Y13_FrameStrobe_O[1] ;
 wire \Tile_X3Y13_FrameStrobe_O[2] ;
 wire \Tile_X3Y13_FrameStrobe_O[3] ;
 wire \Tile_X3Y13_FrameStrobe_O[4] ;
 wire \Tile_X3Y13_FrameStrobe_O[5] ;
 wire \Tile_X3Y13_FrameStrobe_O[6] ;
 wire \Tile_X3Y13_FrameStrobe_O[7] ;
 wire \Tile_X3Y13_FrameStrobe_O[8] ;
 wire \Tile_X3Y13_FrameStrobe_O[9] ;
 wire \Tile_X3Y13_N1BEG[0] ;
 wire \Tile_X3Y13_N1BEG[1] ;
 wire \Tile_X3Y13_N1BEG[2] ;
 wire \Tile_X3Y13_N1BEG[3] ;
 wire \Tile_X3Y13_N2BEG[0] ;
 wire \Tile_X3Y13_N2BEG[1] ;
 wire \Tile_X3Y13_N2BEG[2] ;
 wire \Tile_X3Y13_N2BEG[3] ;
 wire \Tile_X3Y13_N2BEG[4] ;
 wire \Tile_X3Y13_N2BEG[5] ;
 wire \Tile_X3Y13_N2BEG[6] ;
 wire \Tile_X3Y13_N2BEG[7] ;
 wire \Tile_X3Y13_N2BEGb[0] ;
 wire \Tile_X3Y13_N2BEGb[1] ;
 wire \Tile_X3Y13_N2BEGb[2] ;
 wire \Tile_X3Y13_N2BEGb[3] ;
 wire \Tile_X3Y13_N2BEGb[4] ;
 wire \Tile_X3Y13_N2BEGb[5] ;
 wire \Tile_X3Y13_N2BEGb[6] ;
 wire \Tile_X3Y13_N2BEGb[7] ;
 wire \Tile_X3Y13_N4BEG[0] ;
 wire \Tile_X3Y13_N4BEG[10] ;
 wire \Tile_X3Y13_N4BEG[11] ;
 wire \Tile_X3Y13_N4BEG[12] ;
 wire \Tile_X3Y13_N4BEG[13] ;
 wire \Tile_X3Y13_N4BEG[14] ;
 wire \Tile_X3Y13_N4BEG[15] ;
 wire \Tile_X3Y13_N4BEG[1] ;
 wire \Tile_X3Y13_N4BEG[2] ;
 wire \Tile_X3Y13_N4BEG[3] ;
 wire \Tile_X3Y13_N4BEG[4] ;
 wire \Tile_X3Y13_N4BEG[5] ;
 wire \Tile_X3Y13_N4BEG[6] ;
 wire \Tile_X3Y13_N4BEG[7] ;
 wire \Tile_X3Y13_N4BEG[8] ;
 wire \Tile_X3Y13_N4BEG[9] ;
 wire \Tile_X3Y13_NN4BEG[0] ;
 wire \Tile_X3Y13_NN4BEG[10] ;
 wire \Tile_X3Y13_NN4BEG[11] ;
 wire \Tile_X3Y13_NN4BEG[12] ;
 wire \Tile_X3Y13_NN4BEG[13] ;
 wire \Tile_X3Y13_NN4BEG[14] ;
 wire \Tile_X3Y13_NN4BEG[15] ;
 wire \Tile_X3Y13_NN4BEG[1] ;
 wire \Tile_X3Y13_NN4BEG[2] ;
 wire \Tile_X3Y13_NN4BEG[3] ;
 wire \Tile_X3Y13_NN4BEG[4] ;
 wire \Tile_X3Y13_NN4BEG[5] ;
 wire \Tile_X3Y13_NN4BEG[6] ;
 wire \Tile_X3Y13_NN4BEG[7] ;
 wire \Tile_X3Y13_NN4BEG[8] ;
 wire \Tile_X3Y13_NN4BEG[9] ;
 wire \Tile_X3Y13_S1BEG[0] ;
 wire \Tile_X3Y13_S1BEG[1] ;
 wire \Tile_X3Y13_S1BEG[2] ;
 wire \Tile_X3Y13_S1BEG[3] ;
 wire \Tile_X3Y13_S2BEG[0] ;
 wire \Tile_X3Y13_S2BEG[1] ;
 wire \Tile_X3Y13_S2BEG[2] ;
 wire \Tile_X3Y13_S2BEG[3] ;
 wire \Tile_X3Y13_S2BEG[4] ;
 wire \Tile_X3Y13_S2BEG[5] ;
 wire \Tile_X3Y13_S2BEG[6] ;
 wire \Tile_X3Y13_S2BEG[7] ;
 wire \Tile_X3Y13_S2BEGb[0] ;
 wire \Tile_X3Y13_S2BEGb[1] ;
 wire \Tile_X3Y13_S2BEGb[2] ;
 wire \Tile_X3Y13_S2BEGb[3] ;
 wire \Tile_X3Y13_S2BEGb[4] ;
 wire \Tile_X3Y13_S2BEGb[5] ;
 wire \Tile_X3Y13_S2BEGb[6] ;
 wire \Tile_X3Y13_S2BEGb[7] ;
 wire \Tile_X3Y13_S4BEG[0] ;
 wire \Tile_X3Y13_S4BEG[10] ;
 wire \Tile_X3Y13_S4BEG[11] ;
 wire \Tile_X3Y13_S4BEG[12] ;
 wire \Tile_X3Y13_S4BEG[13] ;
 wire \Tile_X3Y13_S4BEG[14] ;
 wire \Tile_X3Y13_S4BEG[15] ;
 wire \Tile_X3Y13_S4BEG[1] ;
 wire \Tile_X3Y13_S4BEG[2] ;
 wire \Tile_X3Y13_S4BEG[3] ;
 wire \Tile_X3Y13_S4BEG[4] ;
 wire \Tile_X3Y13_S4BEG[5] ;
 wire \Tile_X3Y13_S4BEG[6] ;
 wire \Tile_X3Y13_S4BEG[7] ;
 wire \Tile_X3Y13_S4BEG[8] ;
 wire \Tile_X3Y13_S4BEG[9] ;
 wire \Tile_X3Y13_SS4BEG[0] ;
 wire \Tile_X3Y13_SS4BEG[10] ;
 wire \Tile_X3Y13_SS4BEG[11] ;
 wire \Tile_X3Y13_SS4BEG[12] ;
 wire \Tile_X3Y13_SS4BEG[13] ;
 wire \Tile_X3Y13_SS4BEG[14] ;
 wire \Tile_X3Y13_SS4BEG[15] ;
 wire \Tile_X3Y13_SS4BEG[1] ;
 wire \Tile_X3Y13_SS4BEG[2] ;
 wire \Tile_X3Y13_SS4BEG[3] ;
 wire \Tile_X3Y13_SS4BEG[4] ;
 wire \Tile_X3Y13_SS4BEG[5] ;
 wire \Tile_X3Y13_SS4BEG[6] ;
 wire \Tile_X3Y13_SS4BEG[7] ;
 wire \Tile_X3Y13_SS4BEG[8] ;
 wire \Tile_X3Y13_SS4BEG[9] ;
 wire Tile_X3Y13_UserCLKo;
 wire \Tile_X3Y13_W1BEG[0] ;
 wire \Tile_X3Y13_W1BEG[1] ;
 wire \Tile_X3Y13_W1BEG[2] ;
 wire \Tile_X3Y13_W1BEG[3] ;
 wire \Tile_X3Y13_W2BEG[0] ;
 wire \Tile_X3Y13_W2BEG[1] ;
 wire \Tile_X3Y13_W2BEG[2] ;
 wire \Tile_X3Y13_W2BEG[3] ;
 wire \Tile_X3Y13_W2BEG[4] ;
 wire \Tile_X3Y13_W2BEG[5] ;
 wire \Tile_X3Y13_W2BEG[6] ;
 wire \Tile_X3Y13_W2BEG[7] ;
 wire \Tile_X3Y13_W2BEGb[0] ;
 wire \Tile_X3Y13_W2BEGb[1] ;
 wire \Tile_X3Y13_W2BEGb[2] ;
 wire \Tile_X3Y13_W2BEGb[3] ;
 wire \Tile_X3Y13_W2BEGb[4] ;
 wire \Tile_X3Y13_W2BEGb[5] ;
 wire \Tile_X3Y13_W2BEGb[6] ;
 wire \Tile_X3Y13_W2BEGb[7] ;
 wire \Tile_X3Y13_W6BEG[0] ;
 wire \Tile_X3Y13_W6BEG[10] ;
 wire \Tile_X3Y13_W6BEG[11] ;
 wire \Tile_X3Y13_W6BEG[1] ;
 wire \Tile_X3Y13_W6BEG[2] ;
 wire \Tile_X3Y13_W6BEG[3] ;
 wire \Tile_X3Y13_W6BEG[4] ;
 wire \Tile_X3Y13_W6BEG[5] ;
 wire \Tile_X3Y13_W6BEG[6] ;
 wire \Tile_X3Y13_W6BEG[7] ;
 wire \Tile_X3Y13_W6BEG[8] ;
 wire \Tile_X3Y13_W6BEG[9] ;
 wire \Tile_X3Y13_WW4BEG[0] ;
 wire \Tile_X3Y13_WW4BEG[10] ;
 wire \Tile_X3Y13_WW4BEG[11] ;
 wire \Tile_X3Y13_WW4BEG[12] ;
 wire \Tile_X3Y13_WW4BEG[13] ;
 wire \Tile_X3Y13_WW4BEG[14] ;
 wire \Tile_X3Y13_WW4BEG[15] ;
 wire \Tile_X3Y13_WW4BEG[1] ;
 wire \Tile_X3Y13_WW4BEG[2] ;
 wire \Tile_X3Y13_WW4BEG[3] ;
 wire \Tile_X3Y13_WW4BEG[4] ;
 wire \Tile_X3Y13_WW4BEG[5] ;
 wire \Tile_X3Y13_WW4BEG[6] ;
 wire \Tile_X3Y13_WW4BEG[7] ;
 wire \Tile_X3Y13_WW4BEG[8] ;
 wire \Tile_X3Y13_WW4BEG[9] ;
 wire Tile_X3Y14_Co;
 wire \Tile_X3Y14_E1BEG[0] ;
 wire \Tile_X3Y14_E1BEG[1] ;
 wire \Tile_X3Y14_E1BEG[2] ;
 wire \Tile_X3Y14_E1BEG[3] ;
 wire \Tile_X3Y14_E2BEG[0] ;
 wire \Tile_X3Y14_E2BEG[1] ;
 wire \Tile_X3Y14_E2BEG[2] ;
 wire \Tile_X3Y14_E2BEG[3] ;
 wire \Tile_X3Y14_E2BEG[4] ;
 wire \Tile_X3Y14_E2BEG[5] ;
 wire \Tile_X3Y14_E2BEG[6] ;
 wire \Tile_X3Y14_E2BEG[7] ;
 wire \Tile_X3Y14_E2BEGb[0] ;
 wire \Tile_X3Y14_E2BEGb[1] ;
 wire \Tile_X3Y14_E2BEGb[2] ;
 wire \Tile_X3Y14_E2BEGb[3] ;
 wire \Tile_X3Y14_E2BEGb[4] ;
 wire \Tile_X3Y14_E2BEGb[5] ;
 wire \Tile_X3Y14_E2BEGb[6] ;
 wire \Tile_X3Y14_E2BEGb[7] ;
 wire \Tile_X3Y14_E6BEG[0] ;
 wire \Tile_X3Y14_E6BEG[10] ;
 wire \Tile_X3Y14_E6BEG[11] ;
 wire \Tile_X3Y14_E6BEG[1] ;
 wire \Tile_X3Y14_E6BEG[2] ;
 wire \Tile_X3Y14_E6BEG[3] ;
 wire \Tile_X3Y14_E6BEG[4] ;
 wire \Tile_X3Y14_E6BEG[5] ;
 wire \Tile_X3Y14_E6BEG[6] ;
 wire \Tile_X3Y14_E6BEG[7] ;
 wire \Tile_X3Y14_E6BEG[8] ;
 wire \Tile_X3Y14_E6BEG[9] ;
 wire \Tile_X3Y14_EE4BEG[0] ;
 wire \Tile_X3Y14_EE4BEG[10] ;
 wire \Tile_X3Y14_EE4BEG[11] ;
 wire \Tile_X3Y14_EE4BEG[12] ;
 wire \Tile_X3Y14_EE4BEG[13] ;
 wire \Tile_X3Y14_EE4BEG[14] ;
 wire \Tile_X3Y14_EE4BEG[15] ;
 wire \Tile_X3Y14_EE4BEG[1] ;
 wire \Tile_X3Y14_EE4BEG[2] ;
 wire \Tile_X3Y14_EE4BEG[3] ;
 wire \Tile_X3Y14_EE4BEG[4] ;
 wire \Tile_X3Y14_EE4BEG[5] ;
 wire \Tile_X3Y14_EE4BEG[6] ;
 wire \Tile_X3Y14_EE4BEG[7] ;
 wire \Tile_X3Y14_EE4BEG[8] ;
 wire \Tile_X3Y14_EE4BEG[9] ;
 wire \Tile_X3Y14_FrameData_O[0] ;
 wire \Tile_X3Y14_FrameData_O[10] ;
 wire \Tile_X3Y14_FrameData_O[11] ;
 wire \Tile_X3Y14_FrameData_O[12] ;
 wire \Tile_X3Y14_FrameData_O[13] ;
 wire \Tile_X3Y14_FrameData_O[14] ;
 wire \Tile_X3Y14_FrameData_O[15] ;
 wire \Tile_X3Y14_FrameData_O[16] ;
 wire \Tile_X3Y14_FrameData_O[17] ;
 wire \Tile_X3Y14_FrameData_O[18] ;
 wire \Tile_X3Y14_FrameData_O[19] ;
 wire \Tile_X3Y14_FrameData_O[1] ;
 wire \Tile_X3Y14_FrameData_O[20] ;
 wire \Tile_X3Y14_FrameData_O[21] ;
 wire \Tile_X3Y14_FrameData_O[22] ;
 wire \Tile_X3Y14_FrameData_O[23] ;
 wire \Tile_X3Y14_FrameData_O[24] ;
 wire \Tile_X3Y14_FrameData_O[25] ;
 wire \Tile_X3Y14_FrameData_O[26] ;
 wire \Tile_X3Y14_FrameData_O[27] ;
 wire \Tile_X3Y14_FrameData_O[28] ;
 wire \Tile_X3Y14_FrameData_O[29] ;
 wire \Tile_X3Y14_FrameData_O[2] ;
 wire \Tile_X3Y14_FrameData_O[30] ;
 wire \Tile_X3Y14_FrameData_O[31] ;
 wire \Tile_X3Y14_FrameData_O[3] ;
 wire \Tile_X3Y14_FrameData_O[4] ;
 wire \Tile_X3Y14_FrameData_O[5] ;
 wire \Tile_X3Y14_FrameData_O[6] ;
 wire \Tile_X3Y14_FrameData_O[7] ;
 wire \Tile_X3Y14_FrameData_O[8] ;
 wire \Tile_X3Y14_FrameData_O[9] ;
 wire \Tile_X3Y14_FrameStrobe_O[0] ;
 wire \Tile_X3Y14_FrameStrobe_O[10] ;
 wire \Tile_X3Y14_FrameStrobe_O[11] ;
 wire \Tile_X3Y14_FrameStrobe_O[12] ;
 wire \Tile_X3Y14_FrameStrobe_O[13] ;
 wire \Tile_X3Y14_FrameStrobe_O[14] ;
 wire \Tile_X3Y14_FrameStrobe_O[15] ;
 wire \Tile_X3Y14_FrameStrobe_O[16] ;
 wire \Tile_X3Y14_FrameStrobe_O[17] ;
 wire \Tile_X3Y14_FrameStrobe_O[18] ;
 wire \Tile_X3Y14_FrameStrobe_O[19] ;
 wire \Tile_X3Y14_FrameStrobe_O[1] ;
 wire \Tile_X3Y14_FrameStrobe_O[2] ;
 wire \Tile_X3Y14_FrameStrobe_O[3] ;
 wire \Tile_X3Y14_FrameStrobe_O[4] ;
 wire \Tile_X3Y14_FrameStrobe_O[5] ;
 wire \Tile_X3Y14_FrameStrobe_O[6] ;
 wire \Tile_X3Y14_FrameStrobe_O[7] ;
 wire \Tile_X3Y14_FrameStrobe_O[8] ;
 wire \Tile_X3Y14_FrameStrobe_O[9] ;
 wire \Tile_X3Y14_N1BEG[0] ;
 wire \Tile_X3Y14_N1BEG[1] ;
 wire \Tile_X3Y14_N1BEG[2] ;
 wire \Tile_X3Y14_N1BEG[3] ;
 wire \Tile_X3Y14_N2BEG[0] ;
 wire \Tile_X3Y14_N2BEG[1] ;
 wire \Tile_X3Y14_N2BEG[2] ;
 wire \Tile_X3Y14_N2BEG[3] ;
 wire \Tile_X3Y14_N2BEG[4] ;
 wire \Tile_X3Y14_N2BEG[5] ;
 wire \Tile_X3Y14_N2BEG[6] ;
 wire \Tile_X3Y14_N2BEG[7] ;
 wire \Tile_X3Y14_N2BEGb[0] ;
 wire \Tile_X3Y14_N2BEGb[1] ;
 wire \Tile_X3Y14_N2BEGb[2] ;
 wire \Tile_X3Y14_N2BEGb[3] ;
 wire \Tile_X3Y14_N2BEGb[4] ;
 wire \Tile_X3Y14_N2BEGb[5] ;
 wire \Tile_X3Y14_N2BEGb[6] ;
 wire \Tile_X3Y14_N2BEGb[7] ;
 wire \Tile_X3Y14_N4BEG[0] ;
 wire \Tile_X3Y14_N4BEG[10] ;
 wire \Tile_X3Y14_N4BEG[11] ;
 wire \Tile_X3Y14_N4BEG[12] ;
 wire \Tile_X3Y14_N4BEG[13] ;
 wire \Tile_X3Y14_N4BEG[14] ;
 wire \Tile_X3Y14_N4BEG[15] ;
 wire \Tile_X3Y14_N4BEG[1] ;
 wire \Tile_X3Y14_N4BEG[2] ;
 wire \Tile_X3Y14_N4BEG[3] ;
 wire \Tile_X3Y14_N4BEG[4] ;
 wire \Tile_X3Y14_N4BEG[5] ;
 wire \Tile_X3Y14_N4BEG[6] ;
 wire \Tile_X3Y14_N4BEG[7] ;
 wire \Tile_X3Y14_N4BEG[8] ;
 wire \Tile_X3Y14_N4BEG[9] ;
 wire \Tile_X3Y14_NN4BEG[0] ;
 wire \Tile_X3Y14_NN4BEG[10] ;
 wire \Tile_X3Y14_NN4BEG[11] ;
 wire \Tile_X3Y14_NN4BEG[12] ;
 wire \Tile_X3Y14_NN4BEG[13] ;
 wire \Tile_X3Y14_NN4BEG[14] ;
 wire \Tile_X3Y14_NN4BEG[15] ;
 wire \Tile_X3Y14_NN4BEG[1] ;
 wire \Tile_X3Y14_NN4BEG[2] ;
 wire \Tile_X3Y14_NN4BEG[3] ;
 wire \Tile_X3Y14_NN4BEG[4] ;
 wire \Tile_X3Y14_NN4BEG[5] ;
 wire \Tile_X3Y14_NN4BEG[6] ;
 wire \Tile_X3Y14_NN4BEG[7] ;
 wire \Tile_X3Y14_NN4BEG[8] ;
 wire \Tile_X3Y14_NN4BEG[9] ;
 wire \Tile_X3Y14_S1BEG[0] ;
 wire \Tile_X3Y14_S1BEG[1] ;
 wire \Tile_X3Y14_S1BEG[2] ;
 wire \Tile_X3Y14_S1BEG[3] ;
 wire \Tile_X3Y14_S2BEG[0] ;
 wire \Tile_X3Y14_S2BEG[1] ;
 wire \Tile_X3Y14_S2BEG[2] ;
 wire \Tile_X3Y14_S2BEG[3] ;
 wire \Tile_X3Y14_S2BEG[4] ;
 wire \Tile_X3Y14_S2BEG[5] ;
 wire \Tile_X3Y14_S2BEG[6] ;
 wire \Tile_X3Y14_S2BEG[7] ;
 wire \Tile_X3Y14_S2BEGb[0] ;
 wire \Tile_X3Y14_S2BEGb[1] ;
 wire \Tile_X3Y14_S2BEGb[2] ;
 wire \Tile_X3Y14_S2BEGb[3] ;
 wire \Tile_X3Y14_S2BEGb[4] ;
 wire \Tile_X3Y14_S2BEGb[5] ;
 wire \Tile_X3Y14_S2BEGb[6] ;
 wire \Tile_X3Y14_S2BEGb[7] ;
 wire \Tile_X3Y14_S4BEG[0] ;
 wire \Tile_X3Y14_S4BEG[10] ;
 wire \Tile_X3Y14_S4BEG[11] ;
 wire \Tile_X3Y14_S4BEG[12] ;
 wire \Tile_X3Y14_S4BEG[13] ;
 wire \Tile_X3Y14_S4BEG[14] ;
 wire \Tile_X3Y14_S4BEG[15] ;
 wire \Tile_X3Y14_S4BEG[1] ;
 wire \Tile_X3Y14_S4BEG[2] ;
 wire \Tile_X3Y14_S4BEG[3] ;
 wire \Tile_X3Y14_S4BEG[4] ;
 wire \Tile_X3Y14_S4BEG[5] ;
 wire \Tile_X3Y14_S4BEG[6] ;
 wire \Tile_X3Y14_S4BEG[7] ;
 wire \Tile_X3Y14_S4BEG[8] ;
 wire \Tile_X3Y14_S4BEG[9] ;
 wire \Tile_X3Y14_SS4BEG[0] ;
 wire \Tile_X3Y14_SS4BEG[10] ;
 wire \Tile_X3Y14_SS4BEG[11] ;
 wire \Tile_X3Y14_SS4BEG[12] ;
 wire \Tile_X3Y14_SS4BEG[13] ;
 wire \Tile_X3Y14_SS4BEG[14] ;
 wire \Tile_X3Y14_SS4BEG[15] ;
 wire \Tile_X3Y14_SS4BEG[1] ;
 wire \Tile_X3Y14_SS4BEG[2] ;
 wire \Tile_X3Y14_SS4BEG[3] ;
 wire \Tile_X3Y14_SS4BEG[4] ;
 wire \Tile_X3Y14_SS4BEG[5] ;
 wire \Tile_X3Y14_SS4BEG[6] ;
 wire \Tile_X3Y14_SS4BEG[7] ;
 wire \Tile_X3Y14_SS4BEG[8] ;
 wire \Tile_X3Y14_SS4BEG[9] ;
 wire Tile_X3Y14_UserCLKo;
 wire \Tile_X3Y14_W1BEG[0] ;
 wire \Tile_X3Y14_W1BEG[1] ;
 wire \Tile_X3Y14_W1BEG[2] ;
 wire \Tile_X3Y14_W1BEG[3] ;
 wire \Tile_X3Y14_W2BEG[0] ;
 wire \Tile_X3Y14_W2BEG[1] ;
 wire \Tile_X3Y14_W2BEG[2] ;
 wire \Tile_X3Y14_W2BEG[3] ;
 wire \Tile_X3Y14_W2BEG[4] ;
 wire \Tile_X3Y14_W2BEG[5] ;
 wire \Tile_X3Y14_W2BEG[6] ;
 wire \Tile_X3Y14_W2BEG[7] ;
 wire \Tile_X3Y14_W2BEGb[0] ;
 wire \Tile_X3Y14_W2BEGb[1] ;
 wire \Tile_X3Y14_W2BEGb[2] ;
 wire \Tile_X3Y14_W2BEGb[3] ;
 wire \Tile_X3Y14_W2BEGb[4] ;
 wire \Tile_X3Y14_W2BEGb[5] ;
 wire \Tile_X3Y14_W2BEGb[6] ;
 wire \Tile_X3Y14_W2BEGb[7] ;
 wire \Tile_X3Y14_W6BEG[0] ;
 wire \Tile_X3Y14_W6BEG[10] ;
 wire \Tile_X3Y14_W6BEG[11] ;
 wire \Tile_X3Y14_W6BEG[1] ;
 wire \Tile_X3Y14_W6BEG[2] ;
 wire \Tile_X3Y14_W6BEG[3] ;
 wire \Tile_X3Y14_W6BEG[4] ;
 wire \Tile_X3Y14_W6BEG[5] ;
 wire \Tile_X3Y14_W6BEG[6] ;
 wire \Tile_X3Y14_W6BEG[7] ;
 wire \Tile_X3Y14_W6BEG[8] ;
 wire \Tile_X3Y14_W6BEG[9] ;
 wire \Tile_X3Y14_WW4BEG[0] ;
 wire \Tile_X3Y14_WW4BEG[10] ;
 wire \Tile_X3Y14_WW4BEG[11] ;
 wire \Tile_X3Y14_WW4BEG[12] ;
 wire \Tile_X3Y14_WW4BEG[13] ;
 wire \Tile_X3Y14_WW4BEG[14] ;
 wire \Tile_X3Y14_WW4BEG[15] ;
 wire \Tile_X3Y14_WW4BEG[1] ;
 wire \Tile_X3Y14_WW4BEG[2] ;
 wire \Tile_X3Y14_WW4BEG[3] ;
 wire \Tile_X3Y14_WW4BEG[4] ;
 wire \Tile_X3Y14_WW4BEG[5] ;
 wire \Tile_X3Y14_WW4BEG[6] ;
 wire \Tile_X3Y14_WW4BEG[7] ;
 wire \Tile_X3Y14_WW4BEG[8] ;
 wire \Tile_X3Y14_WW4BEG[9] ;
 wire Tile_X3Y15_Co;
 wire \Tile_X3Y15_FrameData_O[0] ;
 wire \Tile_X3Y15_FrameData_O[10] ;
 wire \Tile_X3Y15_FrameData_O[11] ;
 wire \Tile_X3Y15_FrameData_O[12] ;
 wire \Tile_X3Y15_FrameData_O[13] ;
 wire \Tile_X3Y15_FrameData_O[14] ;
 wire \Tile_X3Y15_FrameData_O[15] ;
 wire \Tile_X3Y15_FrameData_O[16] ;
 wire \Tile_X3Y15_FrameData_O[17] ;
 wire \Tile_X3Y15_FrameData_O[18] ;
 wire \Tile_X3Y15_FrameData_O[19] ;
 wire \Tile_X3Y15_FrameData_O[1] ;
 wire \Tile_X3Y15_FrameData_O[20] ;
 wire \Tile_X3Y15_FrameData_O[21] ;
 wire \Tile_X3Y15_FrameData_O[22] ;
 wire \Tile_X3Y15_FrameData_O[23] ;
 wire \Tile_X3Y15_FrameData_O[24] ;
 wire \Tile_X3Y15_FrameData_O[25] ;
 wire \Tile_X3Y15_FrameData_O[26] ;
 wire \Tile_X3Y15_FrameData_O[27] ;
 wire \Tile_X3Y15_FrameData_O[28] ;
 wire \Tile_X3Y15_FrameData_O[29] ;
 wire \Tile_X3Y15_FrameData_O[2] ;
 wire \Tile_X3Y15_FrameData_O[30] ;
 wire \Tile_X3Y15_FrameData_O[31] ;
 wire \Tile_X3Y15_FrameData_O[3] ;
 wire \Tile_X3Y15_FrameData_O[4] ;
 wire \Tile_X3Y15_FrameData_O[5] ;
 wire \Tile_X3Y15_FrameData_O[6] ;
 wire \Tile_X3Y15_FrameData_O[7] ;
 wire \Tile_X3Y15_FrameData_O[8] ;
 wire \Tile_X3Y15_FrameData_O[9] ;
 wire \Tile_X3Y15_FrameStrobe_O[0] ;
 wire \Tile_X3Y15_FrameStrobe_O[10] ;
 wire \Tile_X3Y15_FrameStrobe_O[11] ;
 wire \Tile_X3Y15_FrameStrobe_O[12] ;
 wire \Tile_X3Y15_FrameStrobe_O[13] ;
 wire \Tile_X3Y15_FrameStrobe_O[14] ;
 wire \Tile_X3Y15_FrameStrobe_O[15] ;
 wire \Tile_X3Y15_FrameStrobe_O[16] ;
 wire \Tile_X3Y15_FrameStrobe_O[17] ;
 wire \Tile_X3Y15_FrameStrobe_O[18] ;
 wire \Tile_X3Y15_FrameStrobe_O[19] ;
 wire \Tile_X3Y15_FrameStrobe_O[1] ;
 wire \Tile_X3Y15_FrameStrobe_O[2] ;
 wire \Tile_X3Y15_FrameStrobe_O[3] ;
 wire \Tile_X3Y15_FrameStrobe_O[4] ;
 wire \Tile_X3Y15_FrameStrobe_O[5] ;
 wire \Tile_X3Y15_FrameStrobe_O[6] ;
 wire \Tile_X3Y15_FrameStrobe_O[7] ;
 wire \Tile_X3Y15_FrameStrobe_O[8] ;
 wire \Tile_X3Y15_FrameStrobe_O[9] ;
 wire \Tile_X3Y15_N1BEG[0] ;
 wire \Tile_X3Y15_N1BEG[1] ;
 wire \Tile_X3Y15_N1BEG[2] ;
 wire \Tile_X3Y15_N1BEG[3] ;
 wire \Tile_X3Y15_N2BEG[0] ;
 wire \Tile_X3Y15_N2BEG[1] ;
 wire \Tile_X3Y15_N2BEG[2] ;
 wire \Tile_X3Y15_N2BEG[3] ;
 wire \Tile_X3Y15_N2BEG[4] ;
 wire \Tile_X3Y15_N2BEG[5] ;
 wire \Tile_X3Y15_N2BEG[6] ;
 wire \Tile_X3Y15_N2BEG[7] ;
 wire \Tile_X3Y15_N2BEGb[0] ;
 wire \Tile_X3Y15_N2BEGb[1] ;
 wire \Tile_X3Y15_N2BEGb[2] ;
 wire \Tile_X3Y15_N2BEGb[3] ;
 wire \Tile_X3Y15_N2BEGb[4] ;
 wire \Tile_X3Y15_N2BEGb[5] ;
 wire \Tile_X3Y15_N2BEGb[6] ;
 wire \Tile_X3Y15_N2BEGb[7] ;
 wire \Tile_X3Y15_N4BEG[0] ;
 wire \Tile_X3Y15_N4BEG[10] ;
 wire \Tile_X3Y15_N4BEG[11] ;
 wire \Tile_X3Y15_N4BEG[12] ;
 wire \Tile_X3Y15_N4BEG[13] ;
 wire \Tile_X3Y15_N4BEG[14] ;
 wire \Tile_X3Y15_N4BEG[15] ;
 wire \Tile_X3Y15_N4BEG[1] ;
 wire \Tile_X3Y15_N4BEG[2] ;
 wire \Tile_X3Y15_N4BEG[3] ;
 wire \Tile_X3Y15_N4BEG[4] ;
 wire \Tile_X3Y15_N4BEG[5] ;
 wire \Tile_X3Y15_N4BEG[6] ;
 wire \Tile_X3Y15_N4BEG[7] ;
 wire \Tile_X3Y15_N4BEG[8] ;
 wire \Tile_X3Y15_N4BEG[9] ;
 wire \Tile_X3Y15_NN4BEG[0] ;
 wire \Tile_X3Y15_NN4BEG[10] ;
 wire \Tile_X3Y15_NN4BEG[11] ;
 wire \Tile_X3Y15_NN4BEG[12] ;
 wire \Tile_X3Y15_NN4BEG[13] ;
 wire \Tile_X3Y15_NN4BEG[14] ;
 wire \Tile_X3Y15_NN4BEG[15] ;
 wire \Tile_X3Y15_NN4BEG[1] ;
 wire \Tile_X3Y15_NN4BEG[2] ;
 wire \Tile_X3Y15_NN4BEG[3] ;
 wire \Tile_X3Y15_NN4BEG[4] ;
 wire \Tile_X3Y15_NN4BEG[5] ;
 wire \Tile_X3Y15_NN4BEG[6] ;
 wire \Tile_X3Y15_NN4BEG[7] ;
 wire \Tile_X3Y15_NN4BEG[8] ;
 wire \Tile_X3Y15_NN4BEG[9] ;
 wire Tile_X3Y15_UserCLKo;
 wire Tile_X3Y1_Co;
 wire \Tile_X3Y1_E1BEG[0] ;
 wire \Tile_X3Y1_E1BEG[1] ;
 wire \Tile_X3Y1_E1BEG[2] ;
 wire \Tile_X3Y1_E1BEG[3] ;
 wire \Tile_X3Y1_E2BEG[0] ;
 wire \Tile_X3Y1_E2BEG[1] ;
 wire \Tile_X3Y1_E2BEG[2] ;
 wire \Tile_X3Y1_E2BEG[3] ;
 wire \Tile_X3Y1_E2BEG[4] ;
 wire \Tile_X3Y1_E2BEG[5] ;
 wire \Tile_X3Y1_E2BEG[6] ;
 wire \Tile_X3Y1_E2BEG[7] ;
 wire \Tile_X3Y1_E2BEGb[0] ;
 wire \Tile_X3Y1_E2BEGb[1] ;
 wire \Tile_X3Y1_E2BEGb[2] ;
 wire \Tile_X3Y1_E2BEGb[3] ;
 wire \Tile_X3Y1_E2BEGb[4] ;
 wire \Tile_X3Y1_E2BEGb[5] ;
 wire \Tile_X3Y1_E2BEGb[6] ;
 wire \Tile_X3Y1_E2BEGb[7] ;
 wire \Tile_X3Y1_E6BEG[0] ;
 wire \Tile_X3Y1_E6BEG[10] ;
 wire \Tile_X3Y1_E6BEG[11] ;
 wire \Tile_X3Y1_E6BEG[1] ;
 wire \Tile_X3Y1_E6BEG[2] ;
 wire \Tile_X3Y1_E6BEG[3] ;
 wire \Tile_X3Y1_E6BEG[4] ;
 wire \Tile_X3Y1_E6BEG[5] ;
 wire \Tile_X3Y1_E6BEG[6] ;
 wire \Tile_X3Y1_E6BEG[7] ;
 wire \Tile_X3Y1_E6BEG[8] ;
 wire \Tile_X3Y1_E6BEG[9] ;
 wire \Tile_X3Y1_EE4BEG[0] ;
 wire \Tile_X3Y1_EE4BEG[10] ;
 wire \Tile_X3Y1_EE4BEG[11] ;
 wire \Tile_X3Y1_EE4BEG[12] ;
 wire \Tile_X3Y1_EE4BEG[13] ;
 wire \Tile_X3Y1_EE4BEG[14] ;
 wire \Tile_X3Y1_EE4BEG[15] ;
 wire \Tile_X3Y1_EE4BEG[1] ;
 wire \Tile_X3Y1_EE4BEG[2] ;
 wire \Tile_X3Y1_EE4BEG[3] ;
 wire \Tile_X3Y1_EE4BEG[4] ;
 wire \Tile_X3Y1_EE4BEG[5] ;
 wire \Tile_X3Y1_EE4BEG[6] ;
 wire \Tile_X3Y1_EE4BEG[7] ;
 wire \Tile_X3Y1_EE4BEG[8] ;
 wire \Tile_X3Y1_EE4BEG[9] ;
 wire \Tile_X3Y1_FrameData_O[0] ;
 wire \Tile_X3Y1_FrameData_O[10] ;
 wire \Tile_X3Y1_FrameData_O[11] ;
 wire \Tile_X3Y1_FrameData_O[12] ;
 wire \Tile_X3Y1_FrameData_O[13] ;
 wire \Tile_X3Y1_FrameData_O[14] ;
 wire \Tile_X3Y1_FrameData_O[15] ;
 wire \Tile_X3Y1_FrameData_O[16] ;
 wire \Tile_X3Y1_FrameData_O[17] ;
 wire \Tile_X3Y1_FrameData_O[18] ;
 wire \Tile_X3Y1_FrameData_O[19] ;
 wire \Tile_X3Y1_FrameData_O[1] ;
 wire \Tile_X3Y1_FrameData_O[20] ;
 wire \Tile_X3Y1_FrameData_O[21] ;
 wire \Tile_X3Y1_FrameData_O[22] ;
 wire \Tile_X3Y1_FrameData_O[23] ;
 wire \Tile_X3Y1_FrameData_O[24] ;
 wire \Tile_X3Y1_FrameData_O[25] ;
 wire \Tile_X3Y1_FrameData_O[26] ;
 wire \Tile_X3Y1_FrameData_O[27] ;
 wire \Tile_X3Y1_FrameData_O[28] ;
 wire \Tile_X3Y1_FrameData_O[29] ;
 wire \Tile_X3Y1_FrameData_O[2] ;
 wire \Tile_X3Y1_FrameData_O[30] ;
 wire \Tile_X3Y1_FrameData_O[31] ;
 wire \Tile_X3Y1_FrameData_O[3] ;
 wire \Tile_X3Y1_FrameData_O[4] ;
 wire \Tile_X3Y1_FrameData_O[5] ;
 wire \Tile_X3Y1_FrameData_O[6] ;
 wire \Tile_X3Y1_FrameData_O[7] ;
 wire \Tile_X3Y1_FrameData_O[8] ;
 wire \Tile_X3Y1_FrameData_O[9] ;
 wire \Tile_X3Y1_FrameStrobe_O[0] ;
 wire \Tile_X3Y1_FrameStrobe_O[10] ;
 wire \Tile_X3Y1_FrameStrobe_O[11] ;
 wire \Tile_X3Y1_FrameStrobe_O[12] ;
 wire \Tile_X3Y1_FrameStrobe_O[13] ;
 wire \Tile_X3Y1_FrameStrobe_O[14] ;
 wire \Tile_X3Y1_FrameStrobe_O[15] ;
 wire \Tile_X3Y1_FrameStrobe_O[16] ;
 wire \Tile_X3Y1_FrameStrobe_O[17] ;
 wire \Tile_X3Y1_FrameStrobe_O[18] ;
 wire \Tile_X3Y1_FrameStrobe_O[19] ;
 wire \Tile_X3Y1_FrameStrobe_O[1] ;
 wire \Tile_X3Y1_FrameStrobe_O[2] ;
 wire \Tile_X3Y1_FrameStrobe_O[3] ;
 wire \Tile_X3Y1_FrameStrobe_O[4] ;
 wire \Tile_X3Y1_FrameStrobe_O[5] ;
 wire \Tile_X3Y1_FrameStrobe_O[6] ;
 wire \Tile_X3Y1_FrameStrobe_O[7] ;
 wire \Tile_X3Y1_FrameStrobe_O[8] ;
 wire \Tile_X3Y1_FrameStrobe_O[9] ;
 wire \Tile_X3Y1_N1BEG[0] ;
 wire \Tile_X3Y1_N1BEG[1] ;
 wire \Tile_X3Y1_N1BEG[2] ;
 wire \Tile_X3Y1_N1BEG[3] ;
 wire \Tile_X3Y1_N2BEG[0] ;
 wire \Tile_X3Y1_N2BEG[1] ;
 wire \Tile_X3Y1_N2BEG[2] ;
 wire \Tile_X3Y1_N2BEG[3] ;
 wire \Tile_X3Y1_N2BEG[4] ;
 wire \Tile_X3Y1_N2BEG[5] ;
 wire \Tile_X3Y1_N2BEG[6] ;
 wire \Tile_X3Y1_N2BEG[7] ;
 wire \Tile_X3Y1_N2BEGb[0] ;
 wire \Tile_X3Y1_N2BEGb[1] ;
 wire \Tile_X3Y1_N2BEGb[2] ;
 wire \Tile_X3Y1_N2BEGb[3] ;
 wire \Tile_X3Y1_N2BEGb[4] ;
 wire \Tile_X3Y1_N2BEGb[5] ;
 wire \Tile_X3Y1_N2BEGb[6] ;
 wire \Tile_X3Y1_N2BEGb[7] ;
 wire \Tile_X3Y1_N4BEG[0] ;
 wire \Tile_X3Y1_N4BEG[10] ;
 wire \Tile_X3Y1_N4BEG[11] ;
 wire \Tile_X3Y1_N4BEG[12] ;
 wire \Tile_X3Y1_N4BEG[13] ;
 wire \Tile_X3Y1_N4BEG[14] ;
 wire \Tile_X3Y1_N4BEG[15] ;
 wire \Tile_X3Y1_N4BEG[1] ;
 wire \Tile_X3Y1_N4BEG[2] ;
 wire \Tile_X3Y1_N4BEG[3] ;
 wire \Tile_X3Y1_N4BEG[4] ;
 wire \Tile_X3Y1_N4BEG[5] ;
 wire \Tile_X3Y1_N4BEG[6] ;
 wire \Tile_X3Y1_N4BEG[7] ;
 wire \Tile_X3Y1_N4BEG[8] ;
 wire \Tile_X3Y1_N4BEG[9] ;
 wire \Tile_X3Y1_NN4BEG[0] ;
 wire \Tile_X3Y1_NN4BEG[10] ;
 wire \Tile_X3Y1_NN4BEG[11] ;
 wire \Tile_X3Y1_NN4BEG[12] ;
 wire \Tile_X3Y1_NN4BEG[13] ;
 wire \Tile_X3Y1_NN4BEG[14] ;
 wire \Tile_X3Y1_NN4BEG[15] ;
 wire \Tile_X3Y1_NN4BEG[1] ;
 wire \Tile_X3Y1_NN4BEG[2] ;
 wire \Tile_X3Y1_NN4BEG[3] ;
 wire \Tile_X3Y1_NN4BEG[4] ;
 wire \Tile_X3Y1_NN4BEG[5] ;
 wire \Tile_X3Y1_NN4BEG[6] ;
 wire \Tile_X3Y1_NN4BEG[7] ;
 wire \Tile_X3Y1_NN4BEG[8] ;
 wire \Tile_X3Y1_NN4BEG[9] ;
 wire \Tile_X3Y1_S1BEG[0] ;
 wire \Tile_X3Y1_S1BEG[1] ;
 wire \Tile_X3Y1_S1BEG[2] ;
 wire \Tile_X3Y1_S1BEG[3] ;
 wire \Tile_X3Y1_S2BEG[0] ;
 wire \Tile_X3Y1_S2BEG[1] ;
 wire \Tile_X3Y1_S2BEG[2] ;
 wire \Tile_X3Y1_S2BEG[3] ;
 wire \Tile_X3Y1_S2BEG[4] ;
 wire \Tile_X3Y1_S2BEG[5] ;
 wire \Tile_X3Y1_S2BEG[6] ;
 wire \Tile_X3Y1_S2BEG[7] ;
 wire \Tile_X3Y1_S2BEGb[0] ;
 wire \Tile_X3Y1_S2BEGb[1] ;
 wire \Tile_X3Y1_S2BEGb[2] ;
 wire \Tile_X3Y1_S2BEGb[3] ;
 wire \Tile_X3Y1_S2BEGb[4] ;
 wire \Tile_X3Y1_S2BEGb[5] ;
 wire \Tile_X3Y1_S2BEGb[6] ;
 wire \Tile_X3Y1_S2BEGb[7] ;
 wire \Tile_X3Y1_S4BEG[0] ;
 wire \Tile_X3Y1_S4BEG[10] ;
 wire \Tile_X3Y1_S4BEG[11] ;
 wire \Tile_X3Y1_S4BEG[12] ;
 wire \Tile_X3Y1_S4BEG[13] ;
 wire \Tile_X3Y1_S4BEG[14] ;
 wire \Tile_X3Y1_S4BEG[15] ;
 wire \Tile_X3Y1_S4BEG[1] ;
 wire \Tile_X3Y1_S4BEG[2] ;
 wire \Tile_X3Y1_S4BEG[3] ;
 wire \Tile_X3Y1_S4BEG[4] ;
 wire \Tile_X3Y1_S4BEG[5] ;
 wire \Tile_X3Y1_S4BEG[6] ;
 wire \Tile_X3Y1_S4BEG[7] ;
 wire \Tile_X3Y1_S4BEG[8] ;
 wire \Tile_X3Y1_S4BEG[9] ;
 wire \Tile_X3Y1_SS4BEG[0] ;
 wire \Tile_X3Y1_SS4BEG[10] ;
 wire \Tile_X3Y1_SS4BEG[11] ;
 wire \Tile_X3Y1_SS4BEG[12] ;
 wire \Tile_X3Y1_SS4BEG[13] ;
 wire \Tile_X3Y1_SS4BEG[14] ;
 wire \Tile_X3Y1_SS4BEG[15] ;
 wire \Tile_X3Y1_SS4BEG[1] ;
 wire \Tile_X3Y1_SS4BEG[2] ;
 wire \Tile_X3Y1_SS4BEG[3] ;
 wire \Tile_X3Y1_SS4BEG[4] ;
 wire \Tile_X3Y1_SS4BEG[5] ;
 wire \Tile_X3Y1_SS4BEG[6] ;
 wire \Tile_X3Y1_SS4BEG[7] ;
 wire \Tile_X3Y1_SS4BEG[8] ;
 wire \Tile_X3Y1_SS4BEG[9] ;
 wire Tile_X3Y1_UserCLKo;
 wire \Tile_X3Y1_W1BEG[0] ;
 wire \Tile_X3Y1_W1BEG[1] ;
 wire \Tile_X3Y1_W1BEG[2] ;
 wire \Tile_X3Y1_W1BEG[3] ;
 wire \Tile_X3Y1_W2BEG[0] ;
 wire \Tile_X3Y1_W2BEG[1] ;
 wire \Tile_X3Y1_W2BEG[2] ;
 wire \Tile_X3Y1_W2BEG[3] ;
 wire \Tile_X3Y1_W2BEG[4] ;
 wire \Tile_X3Y1_W2BEG[5] ;
 wire \Tile_X3Y1_W2BEG[6] ;
 wire \Tile_X3Y1_W2BEG[7] ;
 wire \Tile_X3Y1_W2BEGb[0] ;
 wire \Tile_X3Y1_W2BEGb[1] ;
 wire \Tile_X3Y1_W2BEGb[2] ;
 wire \Tile_X3Y1_W2BEGb[3] ;
 wire \Tile_X3Y1_W2BEGb[4] ;
 wire \Tile_X3Y1_W2BEGb[5] ;
 wire \Tile_X3Y1_W2BEGb[6] ;
 wire \Tile_X3Y1_W2BEGb[7] ;
 wire \Tile_X3Y1_W6BEG[0] ;
 wire \Tile_X3Y1_W6BEG[10] ;
 wire \Tile_X3Y1_W6BEG[11] ;
 wire \Tile_X3Y1_W6BEG[1] ;
 wire \Tile_X3Y1_W6BEG[2] ;
 wire \Tile_X3Y1_W6BEG[3] ;
 wire \Tile_X3Y1_W6BEG[4] ;
 wire \Tile_X3Y1_W6BEG[5] ;
 wire \Tile_X3Y1_W6BEG[6] ;
 wire \Tile_X3Y1_W6BEG[7] ;
 wire \Tile_X3Y1_W6BEG[8] ;
 wire \Tile_X3Y1_W6BEG[9] ;
 wire \Tile_X3Y1_WW4BEG[0] ;
 wire \Tile_X3Y1_WW4BEG[10] ;
 wire \Tile_X3Y1_WW4BEG[11] ;
 wire \Tile_X3Y1_WW4BEG[12] ;
 wire \Tile_X3Y1_WW4BEG[13] ;
 wire \Tile_X3Y1_WW4BEG[14] ;
 wire \Tile_X3Y1_WW4BEG[15] ;
 wire \Tile_X3Y1_WW4BEG[1] ;
 wire \Tile_X3Y1_WW4BEG[2] ;
 wire \Tile_X3Y1_WW4BEG[3] ;
 wire \Tile_X3Y1_WW4BEG[4] ;
 wire \Tile_X3Y1_WW4BEG[5] ;
 wire \Tile_X3Y1_WW4BEG[6] ;
 wire \Tile_X3Y1_WW4BEG[7] ;
 wire \Tile_X3Y1_WW4BEG[8] ;
 wire \Tile_X3Y1_WW4BEG[9] ;
 wire Tile_X3Y2_Co;
 wire \Tile_X3Y2_E1BEG[0] ;
 wire \Tile_X3Y2_E1BEG[1] ;
 wire \Tile_X3Y2_E1BEG[2] ;
 wire \Tile_X3Y2_E1BEG[3] ;
 wire \Tile_X3Y2_E2BEG[0] ;
 wire \Tile_X3Y2_E2BEG[1] ;
 wire \Tile_X3Y2_E2BEG[2] ;
 wire \Tile_X3Y2_E2BEG[3] ;
 wire \Tile_X3Y2_E2BEG[4] ;
 wire \Tile_X3Y2_E2BEG[5] ;
 wire \Tile_X3Y2_E2BEG[6] ;
 wire \Tile_X3Y2_E2BEG[7] ;
 wire \Tile_X3Y2_E2BEGb[0] ;
 wire \Tile_X3Y2_E2BEGb[1] ;
 wire \Tile_X3Y2_E2BEGb[2] ;
 wire \Tile_X3Y2_E2BEGb[3] ;
 wire \Tile_X3Y2_E2BEGb[4] ;
 wire \Tile_X3Y2_E2BEGb[5] ;
 wire \Tile_X3Y2_E2BEGb[6] ;
 wire \Tile_X3Y2_E2BEGb[7] ;
 wire \Tile_X3Y2_E6BEG[0] ;
 wire \Tile_X3Y2_E6BEG[10] ;
 wire \Tile_X3Y2_E6BEG[11] ;
 wire \Tile_X3Y2_E6BEG[1] ;
 wire \Tile_X3Y2_E6BEG[2] ;
 wire \Tile_X3Y2_E6BEG[3] ;
 wire \Tile_X3Y2_E6BEG[4] ;
 wire \Tile_X3Y2_E6BEG[5] ;
 wire \Tile_X3Y2_E6BEG[6] ;
 wire \Tile_X3Y2_E6BEG[7] ;
 wire \Tile_X3Y2_E6BEG[8] ;
 wire \Tile_X3Y2_E6BEG[9] ;
 wire \Tile_X3Y2_EE4BEG[0] ;
 wire \Tile_X3Y2_EE4BEG[10] ;
 wire \Tile_X3Y2_EE4BEG[11] ;
 wire \Tile_X3Y2_EE4BEG[12] ;
 wire \Tile_X3Y2_EE4BEG[13] ;
 wire \Tile_X3Y2_EE4BEG[14] ;
 wire \Tile_X3Y2_EE4BEG[15] ;
 wire \Tile_X3Y2_EE4BEG[1] ;
 wire \Tile_X3Y2_EE4BEG[2] ;
 wire \Tile_X3Y2_EE4BEG[3] ;
 wire \Tile_X3Y2_EE4BEG[4] ;
 wire \Tile_X3Y2_EE4BEG[5] ;
 wire \Tile_X3Y2_EE4BEG[6] ;
 wire \Tile_X3Y2_EE4BEG[7] ;
 wire \Tile_X3Y2_EE4BEG[8] ;
 wire \Tile_X3Y2_EE4BEG[9] ;
 wire \Tile_X3Y2_FrameData_O[0] ;
 wire \Tile_X3Y2_FrameData_O[10] ;
 wire \Tile_X3Y2_FrameData_O[11] ;
 wire \Tile_X3Y2_FrameData_O[12] ;
 wire \Tile_X3Y2_FrameData_O[13] ;
 wire \Tile_X3Y2_FrameData_O[14] ;
 wire \Tile_X3Y2_FrameData_O[15] ;
 wire \Tile_X3Y2_FrameData_O[16] ;
 wire \Tile_X3Y2_FrameData_O[17] ;
 wire \Tile_X3Y2_FrameData_O[18] ;
 wire \Tile_X3Y2_FrameData_O[19] ;
 wire \Tile_X3Y2_FrameData_O[1] ;
 wire \Tile_X3Y2_FrameData_O[20] ;
 wire \Tile_X3Y2_FrameData_O[21] ;
 wire \Tile_X3Y2_FrameData_O[22] ;
 wire \Tile_X3Y2_FrameData_O[23] ;
 wire \Tile_X3Y2_FrameData_O[24] ;
 wire \Tile_X3Y2_FrameData_O[25] ;
 wire \Tile_X3Y2_FrameData_O[26] ;
 wire \Tile_X3Y2_FrameData_O[27] ;
 wire \Tile_X3Y2_FrameData_O[28] ;
 wire \Tile_X3Y2_FrameData_O[29] ;
 wire \Tile_X3Y2_FrameData_O[2] ;
 wire \Tile_X3Y2_FrameData_O[30] ;
 wire \Tile_X3Y2_FrameData_O[31] ;
 wire \Tile_X3Y2_FrameData_O[3] ;
 wire \Tile_X3Y2_FrameData_O[4] ;
 wire \Tile_X3Y2_FrameData_O[5] ;
 wire \Tile_X3Y2_FrameData_O[6] ;
 wire \Tile_X3Y2_FrameData_O[7] ;
 wire \Tile_X3Y2_FrameData_O[8] ;
 wire \Tile_X3Y2_FrameData_O[9] ;
 wire \Tile_X3Y2_FrameStrobe_O[0] ;
 wire \Tile_X3Y2_FrameStrobe_O[10] ;
 wire \Tile_X3Y2_FrameStrobe_O[11] ;
 wire \Tile_X3Y2_FrameStrobe_O[12] ;
 wire \Tile_X3Y2_FrameStrobe_O[13] ;
 wire \Tile_X3Y2_FrameStrobe_O[14] ;
 wire \Tile_X3Y2_FrameStrobe_O[15] ;
 wire \Tile_X3Y2_FrameStrobe_O[16] ;
 wire \Tile_X3Y2_FrameStrobe_O[17] ;
 wire \Tile_X3Y2_FrameStrobe_O[18] ;
 wire \Tile_X3Y2_FrameStrobe_O[19] ;
 wire \Tile_X3Y2_FrameStrobe_O[1] ;
 wire \Tile_X3Y2_FrameStrobe_O[2] ;
 wire \Tile_X3Y2_FrameStrobe_O[3] ;
 wire \Tile_X3Y2_FrameStrobe_O[4] ;
 wire \Tile_X3Y2_FrameStrobe_O[5] ;
 wire \Tile_X3Y2_FrameStrobe_O[6] ;
 wire \Tile_X3Y2_FrameStrobe_O[7] ;
 wire \Tile_X3Y2_FrameStrobe_O[8] ;
 wire \Tile_X3Y2_FrameStrobe_O[9] ;
 wire \Tile_X3Y2_N1BEG[0] ;
 wire \Tile_X3Y2_N1BEG[1] ;
 wire \Tile_X3Y2_N1BEG[2] ;
 wire \Tile_X3Y2_N1BEG[3] ;
 wire \Tile_X3Y2_N2BEG[0] ;
 wire \Tile_X3Y2_N2BEG[1] ;
 wire \Tile_X3Y2_N2BEG[2] ;
 wire \Tile_X3Y2_N2BEG[3] ;
 wire \Tile_X3Y2_N2BEG[4] ;
 wire \Tile_X3Y2_N2BEG[5] ;
 wire \Tile_X3Y2_N2BEG[6] ;
 wire \Tile_X3Y2_N2BEG[7] ;
 wire \Tile_X3Y2_N2BEGb[0] ;
 wire \Tile_X3Y2_N2BEGb[1] ;
 wire \Tile_X3Y2_N2BEGb[2] ;
 wire \Tile_X3Y2_N2BEGb[3] ;
 wire \Tile_X3Y2_N2BEGb[4] ;
 wire \Tile_X3Y2_N2BEGb[5] ;
 wire \Tile_X3Y2_N2BEGb[6] ;
 wire \Tile_X3Y2_N2BEGb[7] ;
 wire \Tile_X3Y2_N4BEG[0] ;
 wire \Tile_X3Y2_N4BEG[10] ;
 wire \Tile_X3Y2_N4BEG[11] ;
 wire \Tile_X3Y2_N4BEG[12] ;
 wire \Tile_X3Y2_N4BEG[13] ;
 wire \Tile_X3Y2_N4BEG[14] ;
 wire \Tile_X3Y2_N4BEG[15] ;
 wire \Tile_X3Y2_N4BEG[1] ;
 wire \Tile_X3Y2_N4BEG[2] ;
 wire \Tile_X3Y2_N4BEG[3] ;
 wire \Tile_X3Y2_N4BEG[4] ;
 wire \Tile_X3Y2_N4BEG[5] ;
 wire \Tile_X3Y2_N4BEG[6] ;
 wire \Tile_X3Y2_N4BEG[7] ;
 wire \Tile_X3Y2_N4BEG[8] ;
 wire \Tile_X3Y2_N4BEG[9] ;
 wire \Tile_X3Y2_NN4BEG[0] ;
 wire \Tile_X3Y2_NN4BEG[10] ;
 wire \Tile_X3Y2_NN4BEG[11] ;
 wire \Tile_X3Y2_NN4BEG[12] ;
 wire \Tile_X3Y2_NN4BEG[13] ;
 wire \Tile_X3Y2_NN4BEG[14] ;
 wire \Tile_X3Y2_NN4BEG[15] ;
 wire \Tile_X3Y2_NN4BEG[1] ;
 wire \Tile_X3Y2_NN4BEG[2] ;
 wire \Tile_X3Y2_NN4BEG[3] ;
 wire \Tile_X3Y2_NN4BEG[4] ;
 wire \Tile_X3Y2_NN4BEG[5] ;
 wire \Tile_X3Y2_NN4BEG[6] ;
 wire \Tile_X3Y2_NN4BEG[7] ;
 wire \Tile_X3Y2_NN4BEG[8] ;
 wire \Tile_X3Y2_NN4BEG[9] ;
 wire \Tile_X3Y2_S1BEG[0] ;
 wire \Tile_X3Y2_S1BEG[1] ;
 wire \Tile_X3Y2_S1BEG[2] ;
 wire \Tile_X3Y2_S1BEG[3] ;
 wire \Tile_X3Y2_S2BEG[0] ;
 wire \Tile_X3Y2_S2BEG[1] ;
 wire \Tile_X3Y2_S2BEG[2] ;
 wire \Tile_X3Y2_S2BEG[3] ;
 wire \Tile_X3Y2_S2BEG[4] ;
 wire \Tile_X3Y2_S2BEG[5] ;
 wire \Tile_X3Y2_S2BEG[6] ;
 wire \Tile_X3Y2_S2BEG[7] ;
 wire \Tile_X3Y2_S2BEGb[0] ;
 wire \Tile_X3Y2_S2BEGb[1] ;
 wire \Tile_X3Y2_S2BEGb[2] ;
 wire \Tile_X3Y2_S2BEGb[3] ;
 wire \Tile_X3Y2_S2BEGb[4] ;
 wire \Tile_X3Y2_S2BEGb[5] ;
 wire \Tile_X3Y2_S2BEGb[6] ;
 wire \Tile_X3Y2_S2BEGb[7] ;
 wire \Tile_X3Y2_S4BEG[0] ;
 wire \Tile_X3Y2_S4BEG[10] ;
 wire \Tile_X3Y2_S4BEG[11] ;
 wire \Tile_X3Y2_S4BEG[12] ;
 wire \Tile_X3Y2_S4BEG[13] ;
 wire \Tile_X3Y2_S4BEG[14] ;
 wire \Tile_X3Y2_S4BEG[15] ;
 wire \Tile_X3Y2_S4BEG[1] ;
 wire \Tile_X3Y2_S4BEG[2] ;
 wire \Tile_X3Y2_S4BEG[3] ;
 wire \Tile_X3Y2_S4BEG[4] ;
 wire \Tile_X3Y2_S4BEG[5] ;
 wire \Tile_X3Y2_S4BEG[6] ;
 wire \Tile_X3Y2_S4BEG[7] ;
 wire \Tile_X3Y2_S4BEG[8] ;
 wire \Tile_X3Y2_S4BEG[9] ;
 wire \Tile_X3Y2_SS4BEG[0] ;
 wire \Tile_X3Y2_SS4BEG[10] ;
 wire \Tile_X3Y2_SS4BEG[11] ;
 wire \Tile_X3Y2_SS4BEG[12] ;
 wire \Tile_X3Y2_SS4BEG[13] ;
 wire \Tile_X3Y2_SS4BEG[14] ;
 wire \Tile_X3Y2_SS4BEG[15] ;
 wire \Tile_X3Y2_SS4BEG[1] ;
 wire \Tile_X3Y2_SS4BEG[2] ;
 wire \Tile_X3Y2_SS4BEG[3] ;
 wire \Tile_X3Y2_SS4BEG[4] ;
 wire \Tile_X3Y2_SS4BEG[5] ;
 wire \Tile_X3Y2_SS4BEG[6] ;
 wire \Tile_X3Y2_SS4BEG[7] ;
 wire \Tile_X3Y2_SS4BEG[8] ;
 wire \Tile_X3Y2_SS4BEG[9] ;
 wire Tile_X3Y2_UserCLKo;
 wire \Tile_X3Y2_W1BEG[0] ;
 wire \Tile_X3Y2_W1BEG[1] ;
 wire \Tile_X3Y2_W1BEG[2] ;
 wire \Tile_X3Y2_W1BEG[3] ;
 wire \Tile_X3Y2_W2BEG[0] ;
 wire \Tile_X3Y2_W2BEG[1] ;
 wire \Tile_X3Y2_W2BEG[2] ;
 wire \Tile_X3Y2_W2BEG[3] ;
 wire \Tile_X3Y2_W2BEG[4] ;
 wire \Tile_X3Y2_W2BEG[5] ;
 wire \Tile_X3Y2_W2BEG[6] ;
 wire \Tile_X3Y2_W2BEG[7] ;
 wire \Tile_X3Y2_W2BEGb[0] ;
 wire \Tile_X3Y2_W2BEGb[1] ;
 wire \Tile_X3Y2_W2BEGb[2] ;
 wire \Tile_X3Y2_W2BEGb[3] ;
 wire \Tile_X3Y2_W2BEGb[4] ;
 wire \Tile_X3Y2_W2BEGb[5] ;
 wire \Tile_X3Y2_W2BEGb[6] ;
 wire \Tile_X3Y2_W2BEGb[7] ;
 wire \Tile_X3Y2_W6BEG[0] ;
 wire \Tile_X3Y2_W6BEG[10] ;
 wire \Tile_X3Y2_W6BEG[11] ;
 wire \Tile_X3Y2_W6BEG[1] ;
 wire \Tile_X3Y2_W6BEG[2] ;
 wire \Tile_X3Y2_W6BEG[3] ;
 wire \Tile_X3Y2_W6BEG[4] ;
 wire \Tile_X3Y2_W6BEG[5] ;
 wire \Tile_X3Y2_W6BEG[6] ;
 wire \Tile_X3Y2_W6BEG[7] ;
 wire \Tile_X3Y2_W6BEG[8] ;
 wire \Tile_X3Y2_W6BEG[9] ;
 wire \Tile_X3Y2_WW4BEG[0] ;
 wire \Tile_X3Y2_WW4BEG[10] ;
 wire \Tile_X3Y2_WW4BEG[11] ;
 wire \Tile_X3Y2_WW4BEG[12] ;
 wire \Tile_X3Y2_WW4BEG[13] ;
 wire \Tile_X3Y2_WW4BEG[14] ;
 wire \Tile_X3Y2_WW4BEG[15] ;
 wire \Tile_X3Y2_WW4BEG[1] ;
 wire \Tile_X3Y2_WW4BEG[2] ;
 wire \Tile_X3Y2_WW4BEG[3] ;
 wire \Tile_X3Y2_WW4BEG[4] ;
 wire \Tile_X3Y2_WW4BEG[5] ;
 wire \Tile_X3Y2_WW4BEG[6] ;
 wire \Tile_X3Y2_WW4BEG[7] ;
 wire \Tile_X3Y2_WW4BEG[8] ;
 wire \Tile_X3Y2_WW4BEG[9] ;
 wire Tile_X3Y3_Co;
 wire \Tile_X3Y3_E1BEG[0] ;
 wire \Tile_X3Y3_E1BEG[1] ;
 wire \Tile_X3Y3_E1BEG[2] ;
 wire \Tile_X3Y3_E1BEG[3] ;
 wire \Tile_X3Y3_E2BEG[0] ;
 wire \Tile_X3Y3_E2BEG[1] ;
 wire \Tile_X3Y3_E2BEG[2] ;
 wire \Tile_X3Y3_E2BEG[3] ;
 wire \Tile_X3Y3_E2BEG[4] ;
 wire \Tile_X3Y3_E2BEG[5] ;
 wire \Tile_X3Y3_E2BEG[6] ;
 wire \Tile_X3Y3_E2BEG[7] ;
 wire \Tile_X3Y3_E2BEGb[0] ;
 wire \Tile_X3Y3_E2BEGb[1] ;
 wire \Tile_X3Y3_E2BEGb[2] ;
 wire \Tile_X3Y3_E2BEGb[3] ;
 wire \Tile_X3Y3_E2BEGb[4] ;
 wire \Tile_X3Y3_E2BEGb[5] ;
 wire \Tile_X3Y3_E2BEGb[6] ;
 wire \Tile_X3Y3_E2BEGb[7] ;
 wire \Tile_X3Y3_E6BEG[0] ;
 wire \Tile_X3Y3_E6BEG[10] ;
 wire \Tile_X3Y3_E6BEG[11] ;
 wire \Tile_X3Y3_E6BEG[1] ;
 wire \Tile_X3Y3_E6BEG[2] ;
 wire \Tile_X3Y3_E6BEG[3] ;
 wire \Tile_X3Y3_E6BEG[4] ;
 wire \Tile_X3Y3_E6BEG[5] ;
 wire \Tile_X3Y3_E6BEG[6] ;
 wire \Tile_X3Y3_E6BEG[7] ;
 wire \Tile_X3Y3_E6BEG[8] ;
 wire \Tile_X3Y3_E6BEG[9] ;
 wire \Tile_X3Y3_EE4BEG[0] ;
 wire \Tile_X3Y3_EE4BEG[10] ;
 wire \Tile_X3Y3_EE4BEG[11] ;
 wire \Tile_X3Y3_EE4BEG[12] ;
 wire \Tile_X3Y3_EE4BEG[13] ;
 wire \Tile_X3Y3_EE4BEG[14] ;
 wire \Tile_X3Y3_EE4BEG[15] ;
 wire \Tile_X3Y3_EE4BEG[1] ;
 wire \Tile_X3Y3_EE4BEG[2] ;
 wire \Tile_X3Y3_EE4BEG[3] ;
 wire \Tile_X3Y3_EE4BEG[4] ;
 wire \Tile_X3Y3_EE4BEG[5] ;
 wire \Tile_X3Y3_EE4BEG[6] ;
 wire \Tile_X3Y3_EE4BEG[7] ;
 wire \Tile_X3Y3_EE4BEG[8] ;
 wire \Tile_X3Y3_EE4BEG[9] ;
 wire \Tile_X3Y3_FrameData_O[0] ;
 wire \Tile_X3Y3_FrameData_O[10] ;
 wire \Tile_X3Y3_FrameData_O[11] ;
 wire \Tile_X3Y3_FrameData_O[12] ;
 wire \Tile_X3Y3_FrameData_O[13] ;
 wire \Tile_X3Y3_FrameData_O[14] ;
 wire \Tile_X3Y3_FrameData_O[15] ;
 wire \Tile_X3Y3_FrameData_O[16] ;
 wire \Tile_X3Y3_FrameData_O[17] ;
 wire \Tile_X3Y3_FrameData_O[18] ;
 wire \Tile_X3Y3_FrameData_O[19] ;
 wire \Tile_X3Y3_FrameData_O[1] ;
 wire \Tile_X3Y3_FrameData_O[20] ;
 wire \Tile_X3Y3_FrameData_O[21] ;
 wire \Tile_X3Y3_FrameData_O[22] ;
 wire \Tile_X3Y3_FrameData_O[23] ;
 wire \Tile_X3Y3_FrameData_O[24] ;
 wire \Tile_X3Y3_FrameData_O[25] ;
 wire \Tile_X3Y3_FrameData_O[26] ;
 wire \Tile_X3Y3_FrameData_O[27] ;
 wire \Tile_X3Y3_FrameData_O[28] ;
 wire \Tile_X3Y3_FrameData_O[29] ;
 wire \Tile_X3Y3_FrameData_O[2] ;
 wire \Tile_X3Y3_FrameData_O[30] ;
 wire \Tile_X3Y3_FrameData_O[31] ;
 wire \Tile_X3Y3_FrameData_O[3] ;
 wire \Tile_X3Y3_FrameData_O[4] ;
 wire \Tile_X3Y3_FrameData_O[5] ;
 wire \Tile_X3Y3_FrameData_O[6] ;
 wire \Tile_X3Y3_FrameData_O[7] ;
 wire \Tile_X3Y3_FrameData_O[8] ;
 wire \Tile_X3Y3_FrameData_O[9] ;
 wire \Tile_X3Y3_FrameStrobe_O[0] ;
 wire \Tile_X3Y3_FrameStrobe_O[10] ;
 wire \Tile_X3Y3_FrameStrobe_O[11] ;
 wire \Tile_X3Y3_FrameStrobe_O[12] ;
 wire \Tile_X3Y3_FrameStrobe_O[13] ;
 wire \Tile_X3Y3_FrameStrobe_O[14] ;
 wire \Tile_X3Y3_FrameStrobe_O[15] ;
 wire \Tile_X3Y3_FrameStrobe_O[16] ;
 wire \Tile_X3Y3_FrameStrobe_O[17] ;
 wire \Tile_X3Y3_FrameStrobe_O[18] ;
 wire \Tile_X3Y3_FrameStrobe_O[19] ;
 wire \Tile_X3Y3_FrameStrobe_O[1] ;
 wire \Tile_X3Y3_FrameStrobe_O[2] ;
 wire \Tile_X3Y3_FrameStrobe_O[3] ;
 wire \Tile_X3Y3_FrameStrobe_O[4] ;
 wire \Tile_X3Y3_FrameStrobe_O[5] ;
 wire \Tile_X3Y3_FrameStrobe_O[6] ;
 wire \Tile_X3Y3_FrameStrobe_O[7] ;
 wire \Tile_X3Y3_FrameStrobe_O[8] ;
 wire \Tile_X3Y3_FrameStrobe_O[9] ;
 wire \Tile_X3Y3_N1BEG[0] ;
 wire \Tile_X3Y3_N1BEG[1] ;
 wire \Tile_X3Y3_N1BEG[2] ;
 wire \Tile_X3Y3_N1BEG[3] ;
 wire \Tile_X3Y3_N2BEG[0] ;
 wire \Tile_X3Y3_N2BEG[1] ;
 wire \Tile_X3Y3_N2BEG[2] ;
 wire \Tile_X3Y3_N2BEG[3] ;
 wire \Tile_X3Y3_N2BEG[4] ;
 wire \Tile_X3Y3_N2BEG[5] ;
 wire \Tile_X3Y3_N2BEG[6] ;
 wire \Tile_X3Y3_N2BEG[7] ;
 wire \Tile_X3Y3_N2BEGb[0] ;
 wire \Tile_X3Y3_N2BEGb[1] ;
 wire \Tile_X3Y3_N2BEGb[2] ;
 wire \Tile_X3Y3_N2BEGb[3] ;
 wire \Tile_X3Y3_N2BEGb[4] ;
 wire \Tile_X3Y3_N2BEGb[5] ;
 wire \Tile_X3Y3_N2BEGb[6] ;
 wire \Tile_X3Y3_N2BEGb[7] ;
 wire \Tile_X3Y3_N4BEG[0] ;
 wire \Tile_X3Y3_N4BEG[10] ;
 wire \Tile_X3Y3_N4BEG[11] ;
 wire \Tile_X3Y3_N4BEG[12] ;
 wire \Tile_X3Y3_N4BEG[13] ;
 wire \Tile_X3Y3_N4BEG[14] ;
 wire \Tile_X3Y3_N4BEG[15] ;
 wire \Tile_X3Y3_N4BEG[1] ;
 wire \Tile_X3Y3_N4BEG[2] ;
 wire \Tile_X3Y3_N4BEG[3] ;
 wire \Tile_X3Y3_N4BEG[4] ;
 wire \Tile_X3Y3_N4BEG[5] ;
 wire \Tile_X3Y3_N4BEG[6] ;
 wire \Tile_X3Y3_N4BEG[7] ;
 wire \Tile_X3Y3_N4BEG[8] ;
 wire \Tile_X3Y3_N4BEG[9] ;
 wire \Tile_X3Y3_NN4BEG[0] ;
 wire \Tile_X3Y3_NN4BEG[10] ;
 wire \Tile_X3Y3_NN4BEG[11] ;
 wire \Tile_X3Y3_NN4BEG[12] ;
 wire \Tile_X3Y3_NN4BEG[13] ;
 wire \Tile_X3Y3_NN4BEG[14] ;
 wire \Tile_X3Y3_NN4BEG[15] ;
 wire \Tile_X3Y3_NN4BEG[1] ;
 wire \Tile_X3Y3_NN4BEG[2] ;
 wire \Tile_X3Y3_NN4BEG[3] ;
 wire \Tile_X3Y3_NN4BEG[4] ;
 wire \Tile_X3Y3_NN4BEG[5] ;
 wire \Tile_X3Y3_NN4BEG[6] ;
 wire \Tile_X3Y3_NN4BEG[7] ;
 wire \Tile_X3Y3_NN4BEG[8] ;
 wire \Tile_X3Y3_NN4BEG[9] ;
 wire \Tile_X3Y3_S1BEG[0] ;
 wire \Tile_X3Y3_S1BEG[1] ;
 wire \Tile_X3Y3_S1BEG[2] ;
 wire \Tile_X3Y3_S1BEG[3] ;
 wire \Tile_X3Y3_S2BEG[0] ;
 wire \Tile_X3Y3_S2BEG[1] ;
 wire \Tile_X3Y3_S2BEG[2] ;
 wire \Tile_X3Y3_S2BEG[3] ;
 wire \Tile_X3Y3_S2BEG[4] ;
 wire \Tile_X3Y3_S2BEG[5] ;
 wire \Tile_X3Y3_S2BEG[6] ;
 wire \Tile_X3Y3_S2BEG[7] ;
 wire \Tile_X3Y3_S2BEGb[0] ;
 wire \Tile_X3Y3_S2BEGb[1] ;
 wire \Tile_X3Y3_S2BEGb[2] ;
 wire \Tile_X3Y3_S2BEGb[3] ;
 wire \Tile_X3Y3_S2BEGb[4] ;
 wire \Tile_X3Y3_S2BEGb[5] ;
 wire \Tile_X3Y3_S2BEGb[6] ;
 wire \Tile_X3Y3_S2BEGb[7] ;
 wire \Tile_X3Y3_S4BEG[0] ;
 wire \Tile_X3Y3_S4BEG[10] ;
 wire \Tile_X3Y3_S4BEG[11] ;
 wire \Tile_X3Y3_S4BEG[12] ;
 wire \Tile_X3Y3_S4BEG[13] ;
 wire \Tile_X3Y3_S4BEG[14] ;
 wire \Tile_X3Y3_S4BEG[15] ;
 wire \Tile_X3Y3_S4BEG[1] ;
 wire \Tile_X3Y3_S4BEG[2] ;
 wire \Tile_X3Y3_S4BEG[3] ;
 wire \Tile_X3Y3_S4BEG[4] ;
 wire \Tile_X3Y3_S4BEG[5] ;
 wire \Tile_X3Y3_S4BEG[6] ;
 wire \Tile_X3Y3_S4BEG[7] ;
 wire \Tile_X3Y3_S4BEG[8] ;
 wire \Tile_X3Y3_S4BEG[9] ;
 wire \Tile_X3Y3_SS4BEG[0] ;
 wire \Tile_X3Y3_SS4BEG[10] ;
 wire \Tile_X3Y3_SS4BEG[11] ;
 wire \Tile_X3Y3_SS4BEG[12] ;
 wire \Tile_X3Y3_SS4BEG[13] ;
 wire \Tile_X3Y3_SS4BEG[14] ;
 wire \Tile_X3Y3_SS4BEG[15] ;
 wire \Tile_X3Y3_SS4BEG[1] ;
 wire \Tile_X3Y3_SS4BEG[2] ;
 wire \Tile_X3Y3_SS4BEG[3] ;
 wire \Tile_X3Y3_SS4BEG[4] ;
 wire \Tile_X3Y3_SS4BEG[5] ;
 wire \Tile_X3Y3_SS4BEG[6] ;
 wire \Tile_X3Y3_SS4BEG[7] ;
 wire \Tile_X3Y3_SS4BEG[8] ;
 wire \Tile_X3Y3_SS4BEG[9] ;
 wire Tile_X3Y3_UserCLKo;
 wire \Tile_X3Y3_W1BEG[0] ;
 wire \Tile_X3Y3_W1BEG[1] ;
 wire \Tile_X3Y3_W1BEG[2] ;
 wire \Tile_X3Y3_W1BEG[3] ;
 wire \Tile_X3Y3_W2BEG[0] ;
 wire \Tile_X3Y3_W2BEG[1] ;
 wire \Tile_X3Y3_W2BEG[2] ;
 wire \Tile_X3Y3_W2BEG[3] ;
 wire \Tile_X3Y3_W2BEG[4] ;
 wire \Tile_X3Y3_W2BEG[5] ;
 wire \Tile_X3Y3_W2BEG[6] ;
 wire \Tile_X3Y3_W2BEG[7] ;
 wire \Tile_X3Y3_W2BEGb[0] ;
 wire \Tile_X3Y3_W2BEGb[1] ;
 wire \Tile_X3Y3_W2BEGb[2] ;
 wire \Tile_X3Y3_W2BEGb[3] ;
 wire \Tile_X3Y3_W2BEGb[4] ;
 wire \Tile_X3Y3_W2BEGb[5] ;
 wire \Tile_X3Y3_W2BEGb[6] ;
 wire \Tile_X3Y3_W2BEGb[7] ;
 wire \Tile_X3Y3_W6BEG[0] ;
 wire \Tile_X3Y3_W6BEG[10] ;
 wire \Tile_X3Y3_W6BEG[11] ;
 wire \Tile_X3Y3_W6BEG[1] ;
 wire \Tile_X3Y3_W6BEG[2] ;
 wire \Tile_X3Y3_W6BEG[3] ;
 wire \Tile_X3Y3_W6BEG[4] ;
 wire \Tile_X3Y3_W6BEG[5] ;
 wire \Tile_X3Y3_W6BEG[6] ;
 wire \Tile_X3Y3_W6BEG[7] ;
 wire \Tile_X3Y3_W6BEG[8] ;
 wire \Tile_X3Y3_W6BEG[9] ;
 wire \Tile_X3Y3_WW4BEG[0] ;
 wire \Tile_X3Y3_WW4BEG[10] ;
 wire \Tile_X3Y3_WW4BEG[11] ;
 wire \Tile_X3Y3_WW4BEG[12] ;
 wire \Tile_X3Y3_WW4BEG[13] ;
 wire \Tile_X3Y3_WW4BEG[14] ;
 wire \Tile_X3Y3_WW4BEG[15] ;
 wire \Tile_X3Y3_WW4BEG[1] ;
 wire \Tile_X3Y3_WW4BEG[2] ;
 wire \Tile_X3Y3_WW4BEG[3] ;
 wire \Tile_X3Y3_WW4BEG[4] ;
 wire \Tile_X3Y3_WW4BEG[5] ;
 wire \Tile_X3Y3_WW4BEG[6] ;
 wire \Tile_X3Y3_WW4BEG[7] ;
 wire \Tile_X3Y3_WW4BEG[8] ;
 wire \Tile_X3Y3_WW4BEG[9] ;
 wire Tile_X3Y4_Co;
 wire \Tile_X3Y4_E1BEG[0] ;
 wire \Tile_X3Y4_E1BEG[1] ;
 wire \Tile_X3Y4_E1BEG[2] ;
 wire \Tile_X3Y4_E1BEG[3] ;
 wire \Tile_X3Y4_E2BEG[0] ;
 wire \Tile_X3Y4_E2BEG[1] ;
 wire \Tile_X3Y4_E2BEG[2] ;
 wire \Tile_X3Y4_E2BEG[3] ;
 wire \Tile_X3Y4_E2BEG[4] ;
 wire \Tile_X3Y4_E2BEG[5] ;
 wire \Tile_X3Y4_E2BEG[6] ;
 wire \Tile_X3Y4_E2BEG[7] ;
 wire \Tile_X3Y4_E2BEGb[0] ;
 wire \Tile_X3Y4_E2BEGb[1] ;
 wire \Tile_X3Y4_E2BEGb[2] ;
 wire \Tile_X3Y4_E2BEGb[3] ;
 wire \Tile_X3Y4_E2BEGb[4] ;
 wire \Tile_X3Y4_E2BEGb[5] ;
 wire \Tile_X3Y4_E2BEGb[6] ;
 wire \Tile_X3Y4_E2BEGb[7] ;
 wire \Tile_X3Y4_E6BEG[0] ;
 wire \Tile_X3Y4_E6BEG[10] ;
 wire \Tile_X3Y4_E6BEG[11] ;
 wire \Tile_X3Y4_E6BEG[1] ;
 wire \Tile_X3Y4_E6BEG[2] ;
 wire \Tile_X3Y4_E6BEG[3] ;
 wire \Tile_X3Y4_E6BEG[4] ;
 wire \Tile_X3Y4_E6BEG[5] ;
 wire \Tile_X3Y4_E6BEG[6] ;
 wire \Tile_X3Y4_E6BEG[7] ;
 wire \Tile_X3Y4_E6BEG[8] ;
 wire \Tile_X3Y4_E6BEG[9] ;
 wire \Tile_X3Y4_EE4BEG[0] ;
 wire \Tile_X3Y4_EE4BEG[10] ;
 wire \Tile_X3Y4_EE4BEG[11] ;
 wire \Tile_X3Y4_EE4BEG[12] ;
 wire \Tile_X3Y4_EE4BEG[13] ;
 wire \Tile_X3Y4_EE4BEG[14] ;
 wire \Tile_X3Y4_EE4BEG[15] ;
 wire \Tile_X3Y4_EE4BEG[1] ;
 wire \Tile_X3Y4_EE4BEG[2] ;
 wire \Tile_X3Y4_EE4BEG[3] ;
 wire \Tile_X3Y4_EE4BEG[4] ;
 wire \Tile_X3Y4_EE4BEG[5] ;
 wire \Tile_X3Y4_EE4BEG[6] ;
 wire \Tile_X3Y4_EE4BEG[7] ;
 wire \Tile_X3Y4_EE4BEG[8] ;
 wire \Tile_X3Y4_EE4BEG[9] ;
 wire \Tile_X3Y4_FrameData_O[0] ;
 wire \Tile_X3Y4_FrameData_O[10] ;
 wire \Tile_X3Y4_FrameData_O[11] ;
 wire \Tile_X3Y4_FrameData_O[12] ;
 wire \Tile_X3Y4_FrameData_O[13] ;
 wire \Tile_X3Y4_FrameData_O[14] ;
 wire \Tile_X3Y4_FrameData_O[15] ;
 wire \Tile_X3Y4_FrameData_O[16] ;
 wire \Tile_X3Y4_FrameData_O[17] ;
 wire \Tile_X3Y4_FrameData_O[18] ;
 wire \Tile_X3Y4_FrameData_O[19] ;
 wire \Tile_X3Y4_FrameData_O[1] ;
 wire \Tile_X3Y4_FrameData_O[20] ;
 wire \Tile_X3Y4_FrameData_O[21] ;
 wire \Tile_X3Y4_FrameData_O[22] ;
 wire \Tile_X3Y4_FrameData_O[23] ;
 wire \Tile_X3Y4_FrameData_O[24] ;
 wire \Tile_X3Y4_FrameData_O[25] ;
 wire \Tile_X3Y4_FrameData_O[26] ;
 wire \Tile_X3Y4_FrameData_O[27] ;
 wire \Tile_X3Y4_FrameData_O[28] ;
 wire \Tile_X3Y4_FrameData_O[29] ;
 wire \Tile_X3Y4_FrameData_O[2] ;
 wire \Tile_X3Y4_FrameData_O[30] ;
 wire \Tile_X3Y4_FrameData_O[31] ;
 wire \Tile_X3Y4_FrameData_O[3] ;
 wire \Tile_X3Y4_FrameData_O[4] ;
 wire \Tile_X3Y4_FrameData_O[5] ;
 wire \Tile_X3Y4_FrameData_O[6] ;
 wire \Tile_X3Y4_FrameData_O[7] ;
 wire \Tile_X3Y4_FrameData_O[8] ;
 wire \Tile_X3Y4_FrameData_O[9] ;
 wire \Tile_X3Y4_FrameStrobe_O[0] ;
 wire \Tile_X3Y4_FrameStrobe_O[10] ;
 wire \Tile_X3Y4_FrameStrobe_O[11] ;
 wire \Tile_X3Y4_FrameStrobe_O[12] ;
 wire \Tile_X3Y4_FrameStrobe_O[13] ;
 wire \Tile_X3Y4_FrameStrobe_O[14] ;
 wire \Tile_X3Y4_FrameStrobe_O[15] ;
 wire \Tile_X3Y4_FrameStrobe_O[16] ;
 wire \Tile_X3Y4_FrameStrobe_O[17] ;
 wire \Tile_X3Y4_FrameStrobe_O[18] ;
 wire \Tile_X3Y4_FrameStrobe_O[19] ;
 wire \Tile_X3Y4_FrameStrobe_O[1] ;
 wire \Tile_X3Y4_FrameStrobe_O[2] ;
 wire \Tile_X3Y4_FrameStrobe_O[3] ;
 wire \Tile_X3Y4_FrameStrobe_O[4] ;
 wire \Tile_X3Y4_FrameStrobe_O[5] ;
 wire \Tile_X3Y4_FrameStrobe_O[6] ;
 wire \Tile_X3Y4_FrameStrobe_O[7] ;
 wire \Tile_X3Y4_FrameStrobe_O[8] ;
 wire \Tile_X3Y4_FrameStrobe_O[9] ;
 wire \Tile_X3Y4_N1BEG[0] ;
 wire \Tile_X3Y4_N1BEG[1] ;
 wire \Tile_X3Y4_N1BEG[2] ;
 wire \Tile_X3Y4_N1BEG[3] ;
 wire \Tile_X3Y4_N2BEG[0] ;
 wire \Tile_X3Y4_N2BEG[1] ;
 wire \Tile_X3Y4_N2BEG[2] ;
 wire \Tile_X3Y4_N2BEG[3] ;
 wire \Tile_X3Y4_N2BEG[4] ;
 wire \Tile_X3Y4_N2BEG[5] ;
 wire \Tile_X3Y4_N2BEG[6] ;
 wire \Tile_X3Y4_N2BEG[7] ;
 wire \Tile_X3Y4_N2BEGb[0] ;
 wire \Tile_X3Y4_N2BEGb[1] ;
 wire \Tile_X3Y4_N2BEGb[2] ;
 wire \Tile_X3Y4_N2BEGb[3] ;
 wire \Tile_X3Y4_N2BEGb[4] ;
 wire \Tile_X3Y4_N2BEGb[5] ;
 wire \Tile_X3Y4_N2BEGb[6] ;
 wire \Tile_X3Y4_N2BEGb[7] ;
 wire \Tile_X3Y4_N4BEG[0] ;
 wire \Tile_X3Y4_N4BEG[10] ;
 wire \Tile_X3Y4_N4BEG[11] ;
 wire \Tile_X3Y4_N4BEG[12] ;
 wire \Tile_X3Y4_N4BEG[13] ;
 wire \Tile_X3Y4_N4BEG[14] ;
 wire \Tile_X3Y4_N4BEG[15] ;
 wire \Tile_X3Y4_N4BEG[1] ;
 wire \Tile_X3Y4_N4BEG[2] ;
 wire \Tile_X3Y4_N4BEG[3] ;
 wire \Tile_X3Y4_N4BEG[4] ;
 wire \Tile_X3Y4_N4BEG[5] ;
 wire \Tile_X3Y4_N4BEG[6] ;
 wire \Tile_X3Y4_N4BEG[7] ;
 wire \Tile_X3Y4_N4BEG[8] ;
 wire \Tile_X3Y4_N4BEG[9] ;
 wire \Tile_X3Y4_NN4BEG[0] ;
 wire \Tile_X3Y4_NN4BEG[10] ;
 wire \Tile_X3Y4_NN4BEG[11] ;
 wire \Tile_X3Y4_NN4BEG[12] ;
 wire \Tile_X3Y4_NN4BEG[13] ;
 wire \Tile_X3Y4_NN4BEG[14] ;
 wire \Tile_X3Y4_NN4BEG[15] ;
 wire \Tile_X3Y4_NN4BEG[1] ;
 wire \Tile_X3Y4_NN4BEG[2] ;
 wire \Tile_X3Y4_NN4BEG[3] ;
 wire \Tile_X3Y4_NN4BEG[4] ;
 wire \Tile_X3Y4_NN4BEG[5] ;
 wire \Tile_X3Y4_NN4BEG[6] ;
 wire \Tile_X3Y4_NN4BEG[7] ;
 wire \Tile_X3Y4_NN4BEG[8] ;
 wire \Tile_X3Y4_NN4BEG[9] ;
 wire \Tile_X3Y4_S1BEG[0] ;
 wire \Tile_X3Y4_S1BEG[1] ;
 wire \Tile_X3Y4_S1BEG[2] ;
 wire \Tile_X3Y4_S1BEG[3] ;
 wire \Tile_X3Y4_S2BEG[0] ;
 wire \Tile_X3Y4_S2BEG[1] ;
 wire \Tile_X3Y4_S2BEG[2] ;
 wire \Tile_X3Y4_S2BEG[3] ;
 wire \Tile_X3Y4_S2BEG[4] ;
 wire \Tile_X3Y4_S2BEG[5] ;
 wire \Tile_X3Y4_S2BEG[6] ;
 wire \Tile_X3Y4_S2BEG[7] ;
 wire \Tile_X3Y4_S2BEGb[0] ;
 wire \Tile_X3Y4_S2BEGb[1] ;
 wire \Tile_X3Y4_S2BEGb[2] ;
 wire \Tile_X3Y4_S2BEGb[3] ;
 wire \Tile_X3Y4_S2BEGb[4] ;
 wire \Tile_X3Y4_S2BEGb[5] ;
 wire \Tile_X3Y4_S2BEGb[6] ;
 wire \Tile_X3Y4_S2BEGb[7] ;
 wire \Tile_X3Y4_S4BEG[0] ;
 wire \Tile_X3Y4_S4BEG[10] ;
 wire \Tile_X3Y4_S4BEG[11] ;
 wire \Tile_X3Y4_S4BEG[12] ;
 wire \Tile_X3Y4_S4BEG[13] ;
 wire \Tile_X3Y4_S4BEG[14] ;
 wire \Tile_X3Y4_S4BEG[15] ;
 wire \Tile_X3Y4_S4BEG[1] ;
 wire \Tile_X3Y4_S4BEG[2] ;
 wire \Tile_X3Y4_S4BEG[3] ;
 wire \Tile_X3Y4_S4BEG[4] ;
 wire \Tile_X3Y4_S4BEG[5] ;
 wire \Tile_X3Y4_S4BEG[6] ;
 wire \Tile_X3Y4_S4BEG[7] ;
 wire \Tile_X3Y4_S4BEG[8] ;
 wire \Tile_X3Y4_S4BEG[9] ;
 wire \Tile_X3Y4_SS4BEG[0] ;
 wire \Tile_X3Y4_SS4BEG[10] ;
 wire \Tile_X3Y4_SS4BEG[11] ;
 wire \Tile_X3Y4_SS4BEG[12] ;
 wire \Tile_X3Y4_SS4BEG[13] ;
 wire \Tile_X3Y4_SS4BEG[14] ;
 wire \Tile_X3Y4_SS4BEG[15] ;
 wire \Tile_X3Y4_SS4BEG[1] ;
 wire \Tile_X3Y4_SS4BEG[2] ;
 wire \Tile_X3Y4_SS4BEG[3] ;
 wire \Tile_X3Y4_SS4BEG[4] ;
 wire \Tile_X3Y4_SS4BEG[5] ;
 wire \Tile_X3Y4_SS4BEG[6] ;
 wire \Tile_X3Y4_SS4BEG[7] ;
 wire \Tile_X3Y4_SS4BEG[8] ;
 wire \Tile_X3Y4_SS4BEG[9] ;
 wire Tile_X3Y4_UserCLKo;
 wire \Tile_X3Y4_W1BEG[0] ;
 wire \Tile_X3Y4_W1BEG[1] ;
 wire \Tile_X3Y4_W1BEG[2] ;
 wire \Tile_X3Y4_W1BEG[3] ;
 wire \Tile_X3Y4_W2BEG[0] ;
 wire \Tile_X3Y4_W2BEG[1] ;
 wire \Tile_X3Y4_W2BEG[2] ;
 wire \Tile_X3Y4_W2BEG[3] ;
 wire \Tile_X3Y4_W2BEG[4] ;
 wire \Tile_X3Y4_W2BEG[5] ;
 wire \Tile_X3Y4_W2BEG[6] ;
 wire \Tile_X3Y4_W2BEG[7] ;
 wire \Tile_X3Y4_W2BEGb[0] ;
 wire \Tile_X3Y4_W2BEGb[1] ;
 wire \Tile_X3Y4_W2BEGb[2] ;
 wire \Tile_X3Y4_W2BEGb[3] ;
 wire \Tile_X3Y4_W2BEGb[4] ;
 wire \Tile_X3Y4_W2BEGb[5] ;
 wire \Tile_X3Y4_W2BEGb[6] ;
 wire \Tile_X3Y4_W2BEGb[7] ;
 wire \Tile_X3Y4_W6BEG[0] ;
 wire \Tile_X3Y4_W6BEG[10] ;
 wire \Tile_X3Y4_W6BEG[11] ;
 wire \Tile_X3Y4_W6BEG[1] ;
 wire \Tile_X3Y4_W6BEG[2] ;
 wire \Tile_X3Y4_W6BEG[3] ;
 wire \Tile_X3Y4_W6BEG[4] ;
 wire \Tile_X3Y4_W6BEG[5] ;
 wire \Tile_X3Y4_W6BEG[6] ;
 wire \Tile_X3Y4_W6BEG[7] ;
 wire \Tile_X3Y4_W6BEG[8] ;
 wire \Tile_X3Y4_W6BEG[9] ;
 wire \Tile_X3Y4_WW4BEG[0] ;
 wire \Tile_X3Y4_WW4BEG[10] ;
 wire \Tile_X3Y4_WW4BEG[11] ;
 wire \Tile_X3Y4_WW4BEG[12] ;
 wire \Tile_X3Y4_WW4BEG[13] ;
 wire \Tile_X3Y4_WW4BEG[14] ;
 wire \Tile_X3Y4_WW4BEG[15] ;
 wire \Tile_X3Y4_WW4BEG[1] ;
 wire \Tile_X3Y4_WW4BEG[2] ;
 wire \Tile_X3Y4_WW4BEG[3] ;
 wire \Tile_X3Y4_WW4BEG[4] ;
 wire \Tile_X3Y4_WW4BEG[5] ;
 wire \Tile_X3Y4_WW4BEG[6] ;
 wire \Tile_X3Y4_WW4BEG[7] ;
 wire \Tile_X3Y4_WW4BEG[8] ;
 wire \Tile_X3Y4_WW4BEG[9] ;
 wire Tile_X3Y5_Co;
 wire \Tile_X3Y5_E1BEG[0] ;
 wire \Tile_X3Y5_E1BEG[1] ;
 wire \Tile_X3Y5_E1BEG[2] ;
 wire \Tile_X3Y5_E1BEG[3] ;
 wire \Tile_X3Y5_E2BEG[0] ;
 wire \Tile_X3Y5_E2BEG[1] ;
 wire \Tile_X3Y5_E2BEG[2] ;
 wire \Tile_X3Y5_E2BEG[3] ;
 wire \Tile_X3Y5_E2BEG[4] ;
 wire \Tile_X3Y5_E2BEG[5] ;
 wire \Tile_X3Y5_E2BEG[6] ;
 wire \Tile_X3Y5_E2BEG[7] ;
 wire \Tile_X3Y5_E2BEGb[0] ;
 wire \Tile_X3Y5_E2BEGb[1] ;
 wire \Tile_X3Y5_E2BEGb[2] ;
 wire \Tile_X3Y5_E2BEGb[3] ;
 wire \Tile_X3Y5_E2BEGb[4] ;
 wire \Tile_X3Y5_E2BEGb[5] ;
 wire \Tile_X3Y5_E2BEGb[6] ;
 wire \Tile_X3Y5_E2BEGb[7] ;
 wire \Tile_X3Y5_E6BEG[0] ;
 wire \Tile_X3Y5_E6BEG[10] ;
 wire \Tile_X3Y5_E6BEG[11] ;
 wire \Tile_X3Y5_E6BEG[1] ;
 wire \Tile_X3Y5_E6BEG[2] ;
 wire \Tile_X3Y5_E6BEG[3] ;
 wire \Tile_X3Y5_E6BEG[4] ;
 wire \Tile_X3Y5_E6BEG[5] ;
 wire \Tile_X3Y5_E6BEG[6] ;
 wire \Tile_X3Y5_E6BEG[7] ;
 wire \Tile_X3Y5_E6BEG[8] ;
 wire \Tile_X3Y5_E6BEG[9] ;
 wire \Tile_X3Y5_EE4BEG[0] ;
 wire \Tile_X3Y5_EE4BEG[10] ;
 wire \Tile_X3Y5_EE4BEG[11] ;
 wire \Tile_X3Y5_EE4BEG[12] ;
 wire \Tile_X3Y5_EE4BEG[13] ;
 wire \Tile_X3Y5_EE4BEG[14] ;
 wire \Tile_X3Y5_EE4BEG[15] ;
 wire \Tile_X3Y5_EE4BEG[1] ;
 wire \Tile_X3Y5_EE4BEG[2] ;
 wire \Tile_X3Y5_EE4BEG[3] ;
 wire \Tile_X3Y5_EE4BEG[4] ;
 wire \Tile_X3Y5_EE4BEG[5] ;
 wire \Tile_X3Y5_EE4BEG[6] ;
 wire \Tile_X3Y5_EE4BEG[7] ;
 wire \Tile_X3Y5_EE4BEG[8] ;
 wire \Tile_X3Y5_EE4BEG[9] ;
 wire \Tile_X3Y5_FrameData_O[0] ;
 wire \Tile_X3Y5_FrameData_O[10] ;
 wire \Tile_X3Y5_FrameData_O[11] ;
 wire \Tile_X3Y5_FrameData_O[12] ;
 wire \Tile_X3Y5_FrameData_O[13] ;
 wire \Tile_X3Y5_FrameData_O[14] ;
 wire \Tile_X3Y5_FrameData_O[15] ;
 wire \Tile_X3Y5_FrameData_O[16] ;
 wire \Tile_X3Y5_FrameData_O[17] ;
 wire \Tile_X3Y5_FrameData_O[18] ;
 wire \Tile_X3Y5_FrameData_O[19] ;
 wire \Tile_X3Y5_FrameData_O[1] ;
 wire \Tile_X3Y5_FrameData_O[20] ;
 wire \Tile_X3Y5_FrameData_O[21] ;
 wire \Tile_X3Y5_FrameData_O[22] ;
 wire \Tile_X3Y5_FrameData_O[23] ;
 wire \Tile_X3Y5_FrameData_O[24] ;
 wire \Tile_X3Y5_FrameData_O[25] ;
 wire \Tile_X3Y5_FrameData_O[26] ;
 wire \Tile_X3Y5_FrameData_O[27] ;
 wire \Tile_X3Y5_FrameData_O[28] ;
 wire \Tile_X3Y5_FrameData_O[29] ;
 wire \Tile_X3Y5_FrameData_O[2] ;
 wire \Tile_X3Y5_FrameData_O[30] ;
 wire \Tile_X3Y5_FrameData_O[31] ;
 wire \Tile_X3Y5_FrameData_O[3] ;
 wire \Tile_X3Y5_FrameData_O[4] ;
 wire \Tile_X3Y5_FrameData_O[5] ;
 wire \Tile_X3Y5_FrameData_O[6] ;
 wire \Tile_X3Y5_FrameData_O[7] ;
 wire \Tile_X3Y5_FrameData_O[8] ;
 wire \Tile_X3Y5_FrameData_O[9] ;
 wire \Tile_X3Y5_FrameStrobe_O[0] ;
 wire \Tile_X3Y5_FrameStrobe_O[10] ;
 wire \Tile_X3Y5_FrameStrobe_O[11] ;
 wire \Tile_X3Y5_FrameStrobe_O[12] ;
 wire \Tile_X3Y5_FrameStrobe_O[13] ;
 wire \Tile_X3Y5_FrameStrobe_O[14] ;
 wire \Tile_X3Y5_FrameStrobe_O[15] ;
 wire \Tile_X3Y5_FrameStrobe_O[16] ;
 wire \Tile_X3Y5_FrameStrobe_O[17] ;
 wire \Tile_X3Y5_FrameStrobe_O[18] ;
 wire \Tile_X3Y5_FrameStrobe_O[19] ;
 wire \Tile_X3Y5_FrameStrobe_O[1] ;
 wire \Tile_X3Y5_FrameStrobe_O[2] ;
 wire \Tile_X3Y5_FrameStrobe_O[3] ;
 wire \Tile_X3Y5_FrameStrobe_O[4] ;
 wire \Tile_X3Y5_FrameStrobe_O[5] ;
 wire \Tile_X3Y5_FrameStrobe_O[6] ;
 wire \Tile_X3Y5_FrameStrobe_O[7] ;
 wire \Tile_X3Y5_FrameStrobe_O[8] ;
 wire \Tile_X3Y5_FrameStrobe_O[9] ;
 wire \Tile_X3Y5_N1BEG[0] ;
 wire \Tile_X3Y5_N1BEG[1] ;
 wire \Tile_X3Y5_N1BEG[2] ;
 wire \Tile_X3Y5_N1BEG[3] ;
 wire \Tile_X3Y5_N2BEG[0] ;
 wire \Tile_X3Y5_N2BEG[1] ;
 wire \Tile_X3Y5_N2BEG[2] ;
 wire \Tile_X3Y5_N2BEG[3] ;
 wire \Tile_X3Y5_N2BEG[4] ;
 wire \Tile_X3Y5_N2BEG[5] ;
 wire \Tile_X3Y5_N2BEG[6] ;
 wire \Tile_X3Y5_N2BEG[7] ;
 wire \Tile_X3Y5_N2BEGb[0] ;
 wire \Tile_X3Y5_N2BEGb[1] ;
 wire \Tile_X3Y5_N2BEGb[2] ;
 wire \Tile_X3Y5_N2BEGb[3] ;
 wire \Tile_X3Y5_N2BEGb[4] ;
 wire \Tile_X3Y5_N2BEGb[5] ;
 wire \Tile_X3Y5_N2BEGb[6] ;
 wire \Tile_X3Y5_N2BEGb[7] ;
 wire \Tile_X3Y5_N4BEG[0] ;
 wire \Tile_X3Y5_N4BEG[10] ;
 wire \Tile_X3Y5_N4BEG[11] ;
 wire \Tile_X3Y5_N4BEG[12] ;
 wire \Tile_X3Y5_N4BEG[13] ;
 wire \Tile_X3Y5_N4BEG[14] ;
 wire \Tile_X3Y5_N4BEG[15] ;
 wire \Tile_X3Y5_N4BEG[1] ;
 wire \Tile_X3Y5_N4BEG[2] ;
 wire \Tile_X3Y5_N4BEG[3] ;
 wire \Tile_X3Y5_N4BEG[4] ;
 wire \Tile_X3Y5_N4BEG[5] ;
 wire \Tile_X3Y5_N4BEG[6] ;
 wire \Tile_X3Y5_N4BEG[7] ;
 wire \Tile_X3Y5_N4BEG[8] ;
 wire \Tile_X3Y5_N4BEG[9] ;
 wire \Tile_X3Y5_NN4BEG[0] ;
 wire \Tile_X3Y5_NN4BEG[10] ;
 wire \Tile_X3Y5_NN4BEG[11] ;
 wire \Tile_X3Y5_NN4BEG[12] ;
 wire \Tile_X3Y5_NN4BEG[13] ;
 wire \Tile_X3Y5_NN4BEG[14] ;
 wire \Tile_X3Y5_NN4BEG[15] ;
 wire \Tile_X3Y5_NN4BEG[1] ;
 wire \Tile_X3Y5_NN4BEG[2] ;
 wire \Tile_X3Y5_NN4BEG[3] ;
 wire \Tile_X3Y5_NN4BEG[4] ;
 wire \Tile_X3Y5_NN4BEG[5] ;
 wire \Tile_X3Y5_NN4BEG[6] ;
 wire \Tile_X3Y5_NN4BEG[7] ;
 wire \Tile_X3Y5_NN4BEG[8] ;
 wire \Tile_X3Y5_NN4BEG[9] ;
 wire \Tile_X3Y5_S1BEG[0] ;
 wire \Tile_X3Y5_S1BEG[1] ;
 wire \Tile_X3Y5_S1BEG[2] ;
 wire \Tile_X3Y5_S1BEG[3] ;
 wire \Tile_X3Y5_S2BEG[0] ;
 wire \Tile_X3Y5_S2BEG[1] ;
 wire \Tile_X3Y5_S2BEG[2] ;
 wire \Tile_X3Y5_S2BEG[3] ;
 wire \Tile_X3Y5_S2BEG[4] ;
 wire \Tile_X3Y5_S2BEG[5] ;
 wire \Tile_X3Y5_S2BEG[6] ;
 wire \Tile_X3Y5_S2BEG[7] ;
 wire \Tile_X3Y5_S2BEGb[0] ;
 wire \Tile_X3Y5_S2BEGb[1] ;
 wire \Tile_X3Y5_S2BEGb[2] ;
 wire \Tile_X3Y5_S2BEGb[3] ;
 wire \Tile_X3Y5_S2BEGb[4] ;
 wire \Tile_X3Y5_S2BEGb[5] ;
 wire \Tile_X3Y5_S2BEGb[6] ;
 wire \Tile_X3Y5_S2BEGb[7] ;
 wire \Tile_X3Y5_S4BEG[0] ;
 wire \Tile_X3Y5_S4BEG[10] ;
 wire \Tile_X3Y5_S4BEG[11] ;
 wire \Tile_X3Y5_S4BEG[12] ;
 wire \Tile_X3Y5_S4BEG[13] ;
 wire \Tile_X3Y5_S4BEG[14] ;
 wire \Tile_X3Y5_S4BEG[15] ;
 wire \Tile_X3Y5_S4BEG[1] ;
 wire \Tile_X3Y5_S4BEG[2] ;
 wire \Tile_X3Y5_S4BEG[3] ;
 wire \Tile_X3Y5_S4BEG[4] ;
 wire \Tile_X3Y5_S4BEG[5] ;
 wire \Tile_X3Y5_S4BEG[6] ;
 wire \Tile_X3Y5_S4BEG[7] ;
 wire \Tile_X3Y5_S4BEG[8] ;
 wire \Tile_X3Y5_S4BEG[9] ;
 wire \Tile_X3Y5_SS4BEG[0] ;
 wire \Tile_X3Y5_SS4BEG[10] ;
 wire \Tile_X3Y5_SS4BEG[11] ;
 wire \Tile_X3Y5_SS4BEG[12] ;
 wire \Tile_X3Y5_SS4BEG[13] ;
 wire \Tile_X3Y5_SS4BEG[14] ;
 wire \Tile_X3Y5_SS4BEG[15] ;
 wire \Tile_X3Y5_SS4BEG[1] ;
 wire \Tile_X3Y5_SS4BEG[2] ;
 wire \Tile_X3Y5_SS4BEG[3] ;
 wire \Tile_X3Y5_SS4BEG[4] ;
 wire \Tile_X3Y5_SS4BEG[5] ;
 wire \Tile_X3Y5_SS4BEG[6] ;
 wire \Tile_X3Y5_SS4BEG[7] ;
 wire \Tile_X3Y5_SS4BEG[8] ;
 wire \Tile_X3Y5_SS4BEG[9] ;
 wire Tile_X3Y5_UserCLKo;
 wire \Tile_X3Y5_W1BEG[0] ;
 wire \Tile_X3Y5_W1BEG[1] ;
 wire \Tile_X3Y5_W1BEG[2] ;
 wire \Tile_X3Y5_W1BEG[3] ;
 wire \Tile_X3Y5_W2BEG[0] ;
 wire \Tile_X3Y5_W2BEG[1] ;
 wire \Tile_X3Y5_W2BEG[2] ;
 wire \Tile_X3Y5_W2BEG[3] ;
 wire \Tile_X3Y5_W2BEG[4] ;
 wire \Tile_X3Y5_W2BEG[5] ;
 wire \Tile_X3Y5_W2BEG[6] ;
 wire \Tile_X3Y5_W2BEG[7] ;
 wire \Tile_X3Y5_W2BEGb[0] ;
 wire \Tile_X3Y5_W2BEGb[1] ;
 wire \Tile_X3Y5_W2BEGb[2] ;
 wire \Tile_X3Y5_W2BEGb[3] ;
 wire \Tile_X3Y5_W2BEGb[4] ;
 wire \Tile_X3Y5_W2BEGb[5] ;
 wire \Tile_X3Y5_W2BEGb[6] ;
 wire \Tile_X3Y5_W2BEGb[7] ;
 wire \Tile_X3Y5_W6BEG[0] ;
 wire \Tile_X3Y5_W6BEG[10] ;
 wire \Tile_X3Y5_W6BEG[11] ;
 wire \Tile_X3Y5_W6BEG[1] ;
 wire \Tile_X3Y5_W6BEG[2] ;
 wire \Tile_X3Y5_W6BEG[3] ;
 wire \Tile_X3Y5_W6BEG[4] ;
 wire \Tile_X3Y5_W6BEG[5] ;
 wire \Tile_X3Y5_W6BEG[6] ;
 wire \Tile_X3Y5_W6BEG[7] ;
 wire \Tile_X3Y5_W6BEG[8] ;
 wire \Tile_X3Y5_W6BEG[9] ;
 wire \Tile_X3Y5_WW4BEG[0] ;
 wire \Tile_X3Y5_WW4BEG[10] ;
 wire \Tile_X3Y5_WW4BEG[11] ;
 wire \Tile_X3Y5_WW4BEG[12] ;
 wire \Tile_X3Y5_WW4BEG[13] ;
 wire \Tile_X3Y5_WW4BEG[14] ;
 wire \Tile_X3Y5_WW4BEG[15] ;
 wire \Tile_X3Y5_WW4BEG[1] ;
 wire \Tile_X3Y5_WW4BEG[2] ;
 wire \Tile_X3Y5_WW4BEG[3] ;
 wire \Tile_X3Y5_WW4BEG[4] ;
 wire \Tile_X3Y5_WW4BEG[5] ;
 wire \Tile_X3Y5_WW4BEG[6] ;
 wire \Tile_X3Y5_WW4BEG[7] ;
 wire \Tile_X3Y5_WW4BEG[8] ;
 wire \Tile_X3Y5_WW4BEG[9] ;
 wire Tile_X3Y6_Co;
 wire \Tile_X3Y6_E1BEG[0] ;
 wire \Tile_X3Y6_E1BEG[1] ;
 wire \Tile_X3Y6_E1BEG[2] ;
 wire \Tile_X3Y6_E1BEG[3] ;
 wire \Tile_X3Y6_E2BEG[0] ;
 wire \Tile_X3Y6_E2BEG[1] ;
 wire \Tile_X3Y6_E2BEG[2] ;
 wire \Tile_X3Y6_E2BEG[3] ;
 wire \Tile_X3Y6_E2BEG[4] ;
 wire \Tile_X3Y6_E2BEG[5] ;
 wire \Tile_X3Y6_E2BEG[6] ;
 wire \Tile_X3Y6_E2BEG[7] ;
 wire \Tile_X3Y6_E2BEGb[0] ;
 wire \Tile_X3Y6_E2BEGb[1] ;
 wire \Tile_X3Y6_E2BEGb[2] ;
 wire \Tile_X3Y6_E2BEGb[3] ;
 wire \Tile_X3Y6_E2BEGb[4] ;
 wire \Tile_X3Y6_E2BEGb[5] ;
 wire \Tile_X3Y6_E2BEGb[6] ;
 wire \Tile_X3Y6_E2BEGb[7] ;
 wire \Tile_X3Y6_E6BEG[0] ;
 wire \Tile_X3Y6_E6BEG[10] ;
 wire \Tile_X3Y6_E6BEG[11] ;
 wire \Tile_X3Y6_E6BEG[1] ;
 wire \Tile_X3Y6_E6BEG[2] ;
 wire \Tile_X3Y6_E6BEG[3] ;
 wire \Tile_X3Y6_E6BEG[4] ;
 wire \Tile_X3Y6_E6BEG[5] ;
 wire \Tile_X3Y6_E6BEG[6] ;
 wire \Tile_X3Y6_E6BEG[7] ;
 wire \Tile_X3Y6_E6BEG[8] ;
 wire \Tile_X3Y6_E6BEG[9] ;
 wire \Tile_X3Y6_EE4BEG[0] ;
 wire \Tile_X3Y6_EE4BEG[10] ;
 wire \Tile_X3Y6_EE4BEG[11] ;
 wire \Tile_X3Y6_EE4BEG[12] ;
 wire \Tile_X3Y6_EE4BEG[13] ;
 wire \Tile_X3Y6_EE4BEG[14] ;
 wire \Tile_X3Y6_EE4BEG[15] ;
 wire \Tile_X3Y6_EE4BEG[1] ;
 wire \Tile_X3Y6_EE4BEG[2] ;
 wire \Tile_X3Y6_EE4BEG[3] ;
 wire \Tile_X3Y6_EE4BEG[4] ;
 wire \Tile_X3Y6_EE4BEG[5] ;
 wire \Tile_X3Y6_EE4BEG[6] ;
 wire \Tile_X3Y6_EE4BEG[7] ;
 wire \Tile_X3Y6_EE4BEG[8] ;
 wire \Tile_X3Y6_EE4BEG[9] ;
 wire \Tile_X3Y6_FrameData_O[0] ;
 wire \Tile_X3Y6_FrameData_O[10] ;
 wire \Tile_X3Y6_FrameData_O[11] ;
 wire \Tile_X3Y6_FrameData_O[12] ;
 wire \Tile_X3Y6_FrameData_O[13] ;
 wire \Tile_X3Y6_FrameData_O[14] ;
 wire \Tile_X3Y6_FrameData_O[15] ;
 wire \Tile_X3Y6_FrameData_O[16] ;
 wire \Tile_X3Y6_FrameData_O[17] ;
 wire \Tile_X3Y6_FrameData_O[18] ;
 wire \Tile_X3Y6_FrameData_O[19] ;
 wire \Tile_X3Y6_FrameData_O[1] ;
 wire \Tile_X3Y6_FrameData_O[20] ;
 wire \Tile_X3Y6_FrameData_O[21] ;
 wire \Tile_X3Y6_FrameData_O[22] ;
 wire \Tile_X3Y6_FrameData_O[23] ;
 wire \Tile_X3Y6_FrameData_O[24] ;
 wire \Tile_X3Y6_FrameData_O[25] ;
 wire \Tile_X3Y6_FrameData_O[26] ;
 wire \Tile_X3Y6_FrameData_O[27] ;
 wire \Tile_X3Y6_FrameData_O[28] ;
 wire \Tile_X3Y6_FrameData_O[29] ;
 wire \Tile_X3Y6_FrameData_O[2] ;
 wire \Tile_X3Y6_FrameData_O[30] ;
 wire \Tile_X3Y6_FrameData_O[31] ;
 wire \Tile_X3Y6_FrameData_O[3] ;
 wire \Tile_X3Y6_FrameData_O[4] ;
 wire \Tile_X3Y6_FrameData_O[5] ;
 wire \Tile_X3Y6_FrameData_O[6] ;
 wire \Tile_X3Y6_FrameData_O[7] ;
 wire \Tile_X3Y6_FrameData_O[8] ;
 wire \Tile_X3Y6_FrameData_O[9] ;
 wire \Tile_X3Y6_FrameStrobe_O[0] ;
 wire \Tile_X3Y6_FrameStrobe_O[10] ;
 wire \Tile_X3Y6_FrameStrobe_O[11] ;
 wire \Tile_X3Y6_FrameStrobe_O[12] ;
 wire \Tile_X3Y6_FrameStrobe_O[13] ;
 wire \Tile_X3Y6_FrameStrobe_O[14] ;
 wire \Tile_X3Y6_FrameStrobe_O[15] ;
 wire \Tile_X3Y6_FrameStrobe_O[16] ;
 wire \Tile_X3Y6_FrameStrobe_O[17] ;
 wire \Tile_X3Y6_FrameStrobe_O[18] ;
 wire \Tile_X3Y6_FrameStrobe_O[19] ;
 wire \Tile_X3Y6_FrameStrobe_O[1] ;
 wire \Tile_X3Y6_FrameStrobe_O[2] ;
 wire \Tile_X3Y6_FrameStrobe_O[3] ;
 wire \Tile_X3Y6_FrameStrobe_O[4] ;
 wire \Tile_X3Y6_FrameStrobe_O[5] ;
 wire \Tile_X3Y6_FrameStrobe_O[6] ;
 wire \Tile_X3Y6_FrameStrobe_O[7] ;
 wire \Tile_X3Y6_FrameStrobe_O[8] ;
 wire \Tile_X3Y6_FrameStrobe_O[9] ;
 wire \Tile_X3Y6_N1BEG[0] ;
 wire \Tile_X3Y6_N1BEG[1] ;
 wire \Tile_X3Y6_N1BEG[2] ;
 wire \Tile_X3Y6_N1BEG[3] ;
 wire \Tile_X3Y6_N2BEG[0] ;
 wire \Tile_X3Y6_N2BEG[1] ;
 wire \Tile_X3Y6_N2BEG[2] ;
 wire \Tile_X3Y6_N2BEG[3] ;
 wire \Tile_X3Y6_N2BEG[4] ;
 wire \Tile_X3Y6_N2BEG[5] ;
 wire \Tile_X3Y6_N2BEG[6] ;
 wire \Tile_X3Y6_N2BEG[7] ;
 wire \Tile_X3Y6_N2BEGb[0] ;
 wire \Tile_X3Y6_N2BEGb[1] ;
 wire \Tile_X3Y6_N2BEGb[2] ;
 wire \Tile_X3Y6_N2BEGb[3] ;
 wire \Tile_X3Y6_N2BEGb[4] ;
 wire \Tile_X3Y6_N2BEGb[5] ;
 wire \Tile_X3Y6_N2BEGb[6] ;
 wire \Tile_X3Y6_N2BEGb[7] ;
 wire \Tile_X3Y6_N4BEG[0] ;
 wire \Tile_X3Y6_N4BEG[10] ;
 wire \Tile_X3Y6_N4BEG[11] ;
 wire \Tile_X3Y6_N4BEG[12] ;
 wire \Tile_X3Y6_N4BEG[13] ;
 wire \Tile_X3Y6_N4BEG[14] ;
 wire \Tile_X3Y6_N4BEG[15] ;
 wire \Tile_X3Y6_N4BEG[1] ;
 wire \Tile_X3Y6_N4BEG[2] ;
 wire \Tile_X3Y6_N4BEG[3] ;
 wire \Tile_X3Y6_N4BEG[4] ;
 wire \Tile_X3Y6_N4BEG[5] ;
 wire \Tile_X3Y6_N4BEG[6] ;
 wire \Tile_X3Y6_N4BEG[7] ;
 wire \Tile_X3Y6_N4BEG[8] ;
 wire \Tile_X3Y6_N4BEG[9] ;
 wire \Tile_X3Y6_NN4BEG[0] ;
 wire \Tile_X3Y6_NN4BEG[10] ;
 wire \Tile_X3Y6_NN4BEG[11] ;
 wire \Tile_X3Y6_NN4BEG[12] ;
 wire \Tile_X3Y6_NN4BEG[13] ;
 wire \Tile_X3Y6_NN4BEG[14] ;
 wire \Tile_X3Y6_NN4BEG[15] ;
 wire \Tile_X3Y6_NN4BEG[1] ;
 wire \Tile_X3Y6_NN4BEG[2] ;
 wire \Tile_X3Y6_NN4BEG[3] ;
 wire \Tile_X3Y6_NN4BEG[4] ;
 wire \Tile_X3Y6_NN4BEG[5] ;
 wire \Tile_X3Y6_NN4BEG[6] ;
 wire \Tile_X3Y6_NN4BEG[7] ;
 wire \Tile_X3Y6_NN4BEG[8] ;
 wire \Tile_X3Y6_NN4BEG[9] ;
 wire \Tile_X3Y6_S1BEG[0] ;
 wire \Tile_X3Y6_S1BEG[1] ;
 wire \Tile_X3Y6_S1BEG[2] ;
 wire \Tile_X3Y6_S1BEG[3] ;
 wire \Tile_X3Y6_S2BEG[0] ;
 wire \Tile_X3Y6_S2BEG[1] ;
 wire \Tile_X3Y6_S2BEG[2] ;
 wire \Tile_X3Y6_S2BEG[3] ;
 wire \Tile_X3Y6_S2BEG[4] ;
 wire \Tile_X3Y6_S2BEG[5] ;
 wire \Tile_X3Y6_S2BEG[6] ;
 wire \Tile_X3Y6_S2BEG[7] ;
 wire \Tile_X3Y6_S2BEGb[0] ;
 wire \Tile_X3Y6_S2BEGb[1] ;
 wire \Tile_X3Y6_S2BEGb[2] ;
 wire \Tile_X3Y6_S2BEGb[3] ;
 wire \Tile_X3Y6_S2BEGb[4] ;
 wire \Tile_X3Y6_S2BEGb[5] ;
 wire \Tile_X3Y6_S2BEGb[6] ;
 wire \Tile_X3Y6_S2BEGb[7] ;
 wire \Tile_X3Y6_S4BEG[0] ;
 wire \Tile_X3Y6_S4BEG[10] ;
 wire \Tile_X3Y6_S4BEG[11] ;
 wire \Tile_X3Y6_S4BEG[12] ;
 wire \Tile_X3Y6_S4BEG[13] ;
 wire \Tile_X3Y6_S4BEG[14] ;
 wire \Tile_X3Y6_S4BEG[15] ;
 wire \Tile_X3Y6_S4BEG[1] ;
 wire \Tile_X3Y6_S4BEG[2] ;
 wire \Tile_X3Y6_S4BEG[3] ;
 wire \Tile_X3Y6_S4BEG[4] ;
 wire \Tile_X3Y6_S4BEG[5] ;
 wire \Tile_X3Y6_S4BEG[6] ;
 wire \Tile_X3Y6_S4BEG[7] ;
 wire \Tile_X3Y6_S4BEG[8] ;
 wire \Tile_X3Y6_S4BEG[9] ;
 wire \Tile_X3Y6_SS4BEG[0] ;
 wire \Tile_X3Y6_SS4BEG[10] ;
 wire \Tile_X3Y6_SS4BEG[11] ;
 wire \Tile_X3Y6_SS4BEG[12] ;
 wire \Tile_X3Y6_SS4BEG[13] ;
 wire \Tile_X3Y6_SS4BEG[14] ;
 wire \Tile_X3Y6_SS4BEG[15] ;
 wire \Tile_X3Y6_SS4BEG[1] ;
 wire \Tile_X3Y6_SS4BEG[2] ;
 wire \Tile_X3Y6_SS4BEG[3] ;
 wire \Tile_X3Y6_SS4BEG[4] ;
 wire \Tile_X3Y6_SS4BEG[5] ;
 wire \Tile_X3Y6_SS4BEG[6] ;
 wire \Tile_X3Y6_SS4BEG[7] ;
 wire \Tile_X3Y6_SS4BEG[8] ;
 wire \Tile_X3Y6_SS4BEG[9] ;
 wire Tile_X3Y6_UserCLKo;
 wire \Tile_X3Y6_W1BEG[0] ;
 wire \Tile_X3Y6_W1BEG[1] ;
 wire \Tile_X3Y6_W1BEG[2] ;
 wire \Tile_X3Y6_W1BEG[3] ;
 wire \Tile_X3Y6_W2BEG[0] ;
 wire \Tile_X3Y6_W2BEG[1] ;
 wire \Tile_X3Y6_W2BEG[2] ;
 wire \Tile_X3Y6_W2BEG[3] ;
 wire \Tile_X3Y6_W2BEG[4] ;
 wire \Tile_X3Y6_W2BEG[5] ;
 wire \Tile_X3Y6_W2BEG[6] ;
 wire \Tile_X3Y6_W2BEG[7] ;
 wire \Tile_X3Y6_W2BEGb[0] ;
 wire \Tile_X3Y6_W2BEGb[1] ;
 wire \Tile_X3Y6_W2BEGb[2] ;
 wire \Tile_X3Y6_W2BEGb[3] ;
 wire \Tile_X3Y6_W2BEGb[4] ;
 wire \Tile_X3Y6_W2BEGb[5] ;
 wire \Tile_X3Y6_W2BEGb[6] ;
 wire \Tile_X3Y6_W2BEGb[7] ;
 wire \Tile_X3Y6_W6BEG[0] ;
 wire \Tile_X3Y6_W6BEG[10] ;
 wire \Tile_X3Y6_W6BEG[11] ;
 wire \Tile_X3Y6_W6BEG[1] ;
 wire \Tile_X3Y6_W6BEG[2] ;
 wire \Tile_X3Y6_W6BEG[3] ;
 wire \Tile_X3Y6_W6BEG[4] ;
 wire \Tile_X3Y6_W6BEG[5] ;
 wire \Tile_X3Y6_W6BEG[6] ;
 wire \Tile_X3Y6_W6BEG[7] ;
 wire \Tile_X3Y6_W6BEG[8] ;
 wire \Tile_X3Y6_W6BEG[9] ;
 wire \Tile_X3Y6_WW4BEG[0] ;
 wire \Tile_X3Y6_WW4BEG[10] ;
 wire \Tile_X3Y6_WW4BEG[11] ;
 wire \Tile_X3Y6_WW4BEG[12] ;
 wire \Tile_X3Y6_WW4BEG[13] ;
 wire \Tile_X3Y6_WW4BEG[14] ;
 wire \Tile_X3Y6_WW4BEG[15] ;
 wire \Tile_X3Y6_WW4BEG[1] ;
 wire \Tile_X3Y6_WW4BEG[2] ;
 wire \Tile_X3Y6_WW4BEG[3] ;
 wire \Tile_X3Y6_WW4BEG[4] ;
 wire \Tile_X3Y6_WW4BEG[5] ;
 wire \Tile_X3Y6_WW4BEG[6] ;
 wire \Tile_X3Y6_WW4BEG[7] ;
 wire \Tile_X3Y6_WW4BEG[8] ;
 wire \Tile_X3Y6_WW4BEG[9] ;
 wire Tile_X3Y7_Co;
 wire \Tile_X3Y7_E1BEG[0] ;
 wire \Tile_X3Y7_E1BEG[1] ;
 wire \Tile_X3Y7_E1BEG[2] ;
 wire \Tile_X3Y7_E1BEG[3] ;
 wire \Tile_X3Y7_E2BEG[0] ;
 wire \Tile_X3Y7_E2BEG[1] ;
 wire \Tile_X3Y7_E2BEG[2] ;
 wire \Tile_X3Y7_E2BEG[3] ;
 wire \Tile_X3Y7_E2BEG[4] ;
 wire \Tile_X3Y7_E2BEG[5] ;
 wire \Tile_X3Y7_E2BEG[6] ;
 wire \Tile_X3Y7_E2BEG[7] ;
 wire \Tile_X3Y7_E2BEGb[0] ;
 wire \Tile_X3Y7_E2BEGb[1] ;
 wire \Tile_X3Y7_E2BEGb[2] ;
 wire \Tile_X3Y7_E2BEGb[3] ;
 wire \Tile_X3Y7_E2BEGb[4] ;
 wire \Tile_X3Y7_E2BEGb[5] ;
 wire \Tile_X3Y7_E2BEGb[6] ;
 wire \Tile_X3Y7_E2BEGb[7] ;
 wire \Tile_X3Y7_E6BEG[0] ;
 wire \Tile_X3Y7_E6BEG[10] ;
 wire \Tile_X3Y7_E6BEG[11] ;
 wire \Tile_X3Y7_E6BEG[1] ;
 wire \Tile_X3Y7_E6BEG[2] ;
 wire \Tile_X3Y7_E6BEG[3] ;
 wire \Tile_X3Y7_E6BEG[4] ;
 wire \Tile_X3Y7_E6BEG[5] ;
 wire \Tile_X3Y7_E6BEG[6] ;
 wire \Tile_X3Y7_E6BEG[7] ;
 wire \Tile_X3Y7_E6BEG[8] ;
 wire \Tile_X3Y7_E6BEG[9] ;
 wire \Tile_X3Y7_EE4BEG[0] ;
 wire \Tile_X3Y7_EE4BEG[10] ;
 wire \Tile_X3Y7_EE4BEG[11] ;
 wire \Tile_X3Y7_EE4BEG[12] ;
 wire \Tile_X3Y7_EE4BEG[13] ;
 wire \Tile_X3Y7_EE4BEG[14] ;
 wire \Tile_X3Y7_EE4BEG[15] ;
 wire \Tile_X3Y7_EE4BEG[1] ;
 wire \Tile_X3Y7_EE4BEG[2] ;
 wire \Tile_X3Y7_EE4BEG[3] ;
 wire \Tile_X3Y7_EE4BEG[4] ;
 wire \Tile_X3Y7_EE4BEG[5] ;
 wire \Tile_X3Y7_EE4BEG[6] ;
 wire \Tile_X3Y7_EE4BEG[7] ;
 wire \Tile_X3Y7_EE4BEG[8] ;
 wire \Tile_X3Y7_EE4BEG[9] ;
 wire \Tile_X3Y7_FrameData_O[0] ;
 wire \Tile_X3Y7_FrameData_O[10] ;
 wire \Tile_X3Y7_FrameData_O[11] ;
 wire \Tile_X3Y7_FrameData_O[12] ;
 wire \Tile_X3Y7_FrameData_O[13] ;
 wire \Tile_X3Y7_FrameData_O[14] ;
 wire \Tile_X3Y7_FrameData_O[15] ;
 wire \Tile_X3Y7_FrameData_O[16] ;
 wire \Tile_X3Y7_FrameData_O[17] ;
 wire \Tile_X3Y7_FrameData_O[18] ;
 wire \Tile_X3Y7_FrameData_O[19] ;
 wire \Tile_X3Y7_FrameData_O[1] ;
 wire \Tile_X3Y7_FrameData_O[20] ;
 wire \Tile_X3Y7_FrameData_O[21] ;
 wire \Tile_X3Y7_FrameData_O[22] ;
 wire \Tile_X3Y7_FrameData_O[23] ;
 wire \Tile_X3Y7_FrameData_O[24] ;
 wire \Tile_X3Y7_FrameData_O[25] ;
 wire \Tile_X3Y7_FrameData_O[26] ;
 wire \Tile_X3Y7_FrameData_O[27] ;
 wire \Tile_X3Y7_FrameData_O[28] ;
 wire \Tile_X3Y7_FrameData_O[29] ;
 wire \Tile_X3Y7_FrameData_O[2] ;
 wire \Tile_X3Y7_FrameData_O[30] ;
 wire \Tile_X3Y7_FrameData_O[31] ;
 wire \Tile_X3Y7_FrameData_O[3] ;
 wire \Tile_X3Y7_FrameData_O[4] ;
 wire \Tile_X3Y7_FrameData_O[5] ;
 wire \Tile_X3Y7_FrameData_O[6] ;
 wire \Tile_X3Y7_FrameData_O[7] ;
 wire \Tile_X3Y7_FrameData_O[8] ;
 wire \Tile_X3Y7_FrameData_O[9] ;
 wire \Tile_X3Y7_FrameStrobe_O[0] ;
 wire \Tile_X3Y7_FrameStrobe_O[10] ;
 wire \Tile_X3Y7_FrameStrobe_O[11] ;
 wire \Tile_X3Y7_FrameStrobe_O[12] ;
 wire \Tile_X3Y7_FrameStrobe_O[13] ;
 wire \Tile_X3Y7_FrameStrobe_O[14] ;
 wire \Tile_X3Y7_FrameStrobe_O[15] ;
 wire \Tile_X3Y7_FrameStrobe_O[16] ;
 wire \Tile_X3Y7_FrameStrobe_O[17] ;
 wire \Tile_X3Y7_FrameStrobe_O[18] ;
 wire \Tile_X3Y7_FrameStrobe_O[19] ;
 wire \Tile_X3Y7_FrameStrobe_O[1] ;
 wire \Tile_X3Y7_FrameStrobe_O[2] ;
 wire \Tile_X3Y7_FrameStrobe_O[3] ;
 wire \Tile_X3Y7_FrameStrobe_O[4] ;
 wire \Tile_X3Y7_FrameStrobe_O[5] ;
 wire \Tile_X3Y7_FrameStrobe_O[6] ;
 wire \Tile_X3Y7_FrameStrobe_O[7] ;
 wire \Tile_X3Y7_FrameStrobe_O[8] ;
 wire \Tile_X3Y7_FrameStrobe_O[9] ;
 wire \Tile_X3Y7_N1BEG[0] ;
 wire \Tile_X3Y7_N1BEG[1] ;
 wire \Tile_X3Y7_N1BEG[2] ;
 wire \Tile_X3Y7_N1BEG[3] ;
 wire \Tile_X3Y7_N2BEG[0] ;
 wire \Tile_X3Y7_N2BEG[1] ;
 wire \Tile_X3Y7_N2BEG[2] ;
 wire \Tile_X3Y7_N2BEG[3] ;
 wire \Tile_X3Y7_N2BEG[4] ;
 wire \Tile_X3Y7_N2BEG[5] ;
 wire \Tile_X3Y7_N2BEG[6] ;
 wire \Tile_X3Y7_N2BEG[7] ;
 wire \Tile_X3Y7_N2BEGb[0] ;
 wire \Tile_X3Y7_N2BEGb[1] ;
 wire \Tile_X3Y7_N2BEGb[2] ;
 wire \Tile_X3Y7_N2BEGb[3] ;
 wire \Tile_X3Y7_N2BEGb[4] ;
 wire \Tile_X3Y7_N2BEGb[5] ;
 wire \Tile_X3Y7_N2BEGb[6] ;
 wire \Tile_X3Y7_N2BEGb[7] ;
 wire \Tile_X3Y7_N4BEG[0] ;
 wire \Tile_X3Y7_N4BEG[10] ;
 wire \Tile_X3Y7_N4BEG[11] ;
 wire \Tile_X3Y7_N4BEG[12] ;
 wire \Tile_X3Y7_N4BEG[13] ;
 wire \Tile_X3Y7_N4BEG[14] ;
 wire \Tile_X3Y7_N4BEG[15] ;
 wire \Tile_X3Y7_N4BEG[1] ;
 wire \Tile_X3Y7_N4BEG[2] ;
 wire \Tile_X3Y7_N4BEG[3] ;
 wire \Tile_X3Y7_N4BEG[4] ;
 wire \Tile_X3Y7_N4BEG[5] ;
 wire \Tile_X3Y7_N4BEG[6] ;
 wire \Tile_X3Y7_N4BEG[7] ;
 wire \Tile_X3Y7_N4BEG[8] ;
 wire \Tile_X3Y7_N4BEG[9] ;
 wire \Tile_X3Y7_NN4BEG[0] ;
 wire \Tile_X3Y7_NN4BEG[10] ;
 wire \Tile_X3Y7_NN4BEG[11] ;
 wire \Tile_X3Y7_NN4BEG[12] ;
 wire \Tile_X3Y7_NN4BEG[13] ;
 wire \Tile_X3Y7_NN4BEG[14] ;
 wire \Tile_X3Y7_NN4BEG[15] ;
 wire \Tile_X3Y7_NN4BEG[1] ;
 wire \Tile_X3Y7_NN4BEG[2] ;
 wire \Tile_X3Y7_NN4BEG[3] ;
 wire \Tile_X3Y7_NN4BEG[4] ;
 wire \Tile_X3Y7_NN4BEG[5] ;
 wire \Tile_X3Y7_NN4BEG[6] ;
 wire \Tile_X3Y7_NN4BEG[7] ;
 wire \Tile_X3Y7_NN4BEG[8] ;
 wire \Tile_X3Y7_NN4BEG[9] ;
 wire \Tile_X3Y7_S1BEG[0] ;
 wire \Tile_X3Y7_S1BEG[1] ;
 wire \Tile_X3Y7_S1BEG[2] ;
 wire \Tile_X3Y7_S1BEG[3] ;
 wire \Tile_X3Y7_S2BEG[0] ;
 wire \Tile_X3Y7_S2BEG[1] ;
 wire \Tile_X3Y7_S2BEG[2] ;
 wire \Tile_X3Y7_S2BEG[3] ;
 wire \Tile_X3Y7_S2BEG[4] ;
 wire \Tile_X3Y7_S2BEG[5] ;
 wire \Tile_X3Y7_S2BEG[6] ;
 wire \Tile_X3Y7_S2BEG[7] ;
 wire \Tile_X3Y7_S2BEGb[0] ;
 wire \Tile_X3Y7_S2BEGb[1] ;
 wire \Tile_X3Y7_S2BEGb[2] ;
 wire \Tile_X3Y7_S2BEGb[3] ;
 wire \Tile_X3Y7_S2BEGb[4] ;
 wire \Tile_X3Y7_S2BEGb[5] ;
 wire \Tile_X3Y7_S2BEGb[6] ;
 wire \Tile_X3Y7_S2BEGb[7] ;
 wire \Tile_X3Y7_S4BEG[0] ;
 wire \Tile_X3Y7_S4BEG[10] ;
 wire \Tile_X3Y7_S4BEG[11] ;
 wire \Tile_X3Y7_S4BEG[12] ;
 wire \Tile_X3Y7_S4BEG[13] ;
 wire \Tile_X3Y7_S4BEG[14] ;
 wire \Tile_X3Y7_S4BEG[15] ;
 wire \Tile_X3Y7_S4BEG[1] ;
 wire \Tile_X3Y7_S4BEG[2] ;
 wire \Tile_X3Y7_S4BEG[3] ;
 wire \Tile_X3Y7_S4BEG[4] ;
 wire \Tile_X3Y7_S4BEG[5] ;
 wire \Tile_X3Y7_S4BEG[6] ;
 wire \Tile_X3Y7_S4BEG[7] ;
 wire \Tile_X3Y7_S4BEG[8] ;
 wire \Tile_X3Y7_S4BEG[9] ;
 wire \Tile_X3Y7_SS4BEG[0] ;
 wire \Tile_X3Y7_SS4BEG[10] ;
 wire \Tile_X3Y7_SS4BEG[11] ;
 wire \Tile_X3Y7_SS4BEG[12] ;
 wire \Tile_X3Y7_SS4BEG[13] ;
 wire \Tile_X3Y7_SS4BEG[14] ;
 wire \Tile_X3Y7_SS4BEG[15] ;
 wire \Tile_X3Y7_SS4BEG[1] ;
 wire \Tile_X3Y7_SS4BEG[2] ;
 wire \Tile_X3Y7_SS4BEG[3] ;
 wire \Tile_X3Y7_SS4BEG[4] ;
 wire \Tile_X3Y7_SS4BEG[5] ;
 wire \Tile_X3Y7_SS4BEG[6] ;
 wire \Tile_X3Y7_SS4BEG[7] ;
 wire \Tile_X3Y7_SS4BEG[8] ;
 wire \Tile_X3Y7_SS4BEG[9] ;
 wire Tile_X3Y7_UserCLKo;
 wire \Tile_X3Y7_W1BEG[0] ;
 wire \Tile_X3Y7_W1BEG[1] ;
 wire \Tile_X3Y7_W1BEG[2] ;
 wire \Tile_X3Y7_W1BEG[3] ;
 wire \Tile_X3Y7_W2BEG[0] ;
 wire \Tile_X3Y7_W2BEG[1] ;
 wire \Tile_X3Y7_W2BEG[2] ;
 wire \Tile_X3Y7_W2BEG[3] ;
 wire \Tile_X3Y7_W2BEG[4] ;
 wire \Tile_X3Y7_W2BEG[5] ;
 wire \Tile_X3Y7_W2BEG[6] ;
 wire \Tile_X3Y7_W2BEG[7] ;
 wire \Tile_X3Y7_W2BEGb[0] ;
 wire \Tile_X3Y7_W2BEGb[1] ;
 wire \Tile_X3Y7_W2BEGb[2] ;
 wire \Tile_X3Y7_W2BEGb[3] ;
 wire \Tile_X3Y7_W2BEGb[4] ;
 wire \Tile_X3Y7_W2BEGb[5] ;
 wire \Tile_X3Y7_W2BEGb[6] ;
 wire \Tile_X3Y7_W2BEGb[7] ;
 wire \Tile_X3Y7_W6BEG[0] ;
 wire \Tile_X3Y7_W6BEG[10] ;
 wire \Tile_X3Y7_W6BEG[11] ;
 wire \Tile_X3Y7_W6BEG[1] ;
 wire \Tile_X3Y7_W6BEG[2] ;
 wire \Tile_X3Y7_W6BEG[3] ;
 wire \Tile_X3Y7_W6BEG[4] ;
 wire \Tile_X3Y7_W6BEG[5] ;
 wire \Tile_X3Y7_W6BEG[6] ;
 wire \Tile_X3Y7_W6BEG[7] ;
 wire \Tile_X3Y7_W6BEG[8] ;
 wire \Tile_X3Y7_W6BEG[9] ;
 wire \Tile_X3Y7_WW4BEG[0] ;
 wire \Tile_X3Y7_WW4BEG[10] ;
 wire \Tile_X3Y7_WW4BEG[11] ;
 wire \Tile_X3Y7_WW4BEG[12] ;
 wire \Tile_X3Y7_WW4BEG[13] ;
 wire \Tile_X3Y7_WW4BEG[14] ;
 wire \Tile_X3Y7_WW4BEG[15] ;
 wire \Tile_X3Y7_WW4BEG[1] ;
 wire \Tile_X3Y7_WW4BEG[2] ;
 wire \Tile_X3Y7_WW4BEG[3] ;
 wire \Tile_X3Y7_WW4BEG[4] ;
 wire \Tile_X3Y7_WW4BEG[5] ;
 wire \Tile_X3Y7_WW4BEG[6] ;
 wire \Tile_X3Y7_WW4BEG[7] ;
 wire \Tile_X3Y7_WW4BEG[8] ;
 wire \Tile_X3Y7_WW4BEG[9] ;
 wire Tile_X3Y8_Co;
 wire \Tile_X3Y8_E1BEG[0] ;
 wire \Tile_X3Y8_E1BEG[1] ;
 wire \Tile_X3Y8_E1BEG[2] ;
 wire \Tile_X3Y8_E1BEG[3] ;
 wire \Tile_X3Y8_E2BEG[0] ;
 wire \Tile_X3Y8_E2BEG[1] ;
 wire \Tile_X3Y8_E2BEG[2] ;
 wire \Tile_X3Y8_E2BEG[3] ;
 wire \Tile_X3Y8_E2BEG[4] ;
 wire \Tile_X3Y8_E2BEG[5] ;
 wire \Tile_X3Y8_E2BEG[6] ;
 wire \Tile_X3Y8_E2BEG[7] ;
 wire \Tile_X3Y8_E2BEGb[0] ;
 wire \Tile_X3Y8_E2BEGb[1] ;
 wire \Tile_X3Y8_E2BEGb[2] ;
 wire \Tile_X3Y8_E2BEGb[3] ;
 wire \Tile_X3Y8_E2BEGb[4] ;
 wire \Tile_X3Y8_E2BEGb[5] ;
 wire \Tile_X3Y8_E2BEGb[6] ;
 wire \Tile_X3Y8_E2BEGb[7] ;
 wire \Tile_X3Y8_E6BEG[0] ;
 wire \Tile_X3Y8_E6BEG[10] ;
 wire \Tile_X3Y8_E6BEG[11] ;
 wire \Tile_X3Y8_E6BEG[1] ;
 wire \Tile_X3Y8_E6BEG[2] ;
 wire \Tile_X3Y8_E6BEG[3] ;
 wire \Tile_X3Y8_E6BEG[4] ;
 wire \Tile_X3Y8_E6BEG[5] ;
 wire \Tile_X3Y8_E6BEG[6] ;
 wire \Tile_X3Y8_E6BEG[7] ;
 wire \Tile_X3Y8_E6BEG[8] ;
 wire \Tile_X3Y8_E6BEG[9] ;
 wire \Tile_X3Y8_EE4BEG[0] ;
 wire \Tile_X3Y8_EE4BEG[10] ;
 wire \Tile_X3Y8_EE4BEG[11] ;
 wire \Tile_X3Y8_EE4BEG[12] ;
 wire \Tile_X3Y8_EE4BEG[13] ;
 wire \Tile_X3Y8_EE4BEG[14] ;
 wire \Tile_X3Y8_EE4BEG[15] ;
 wire \Tile_X3Y8_EE4BEG[1] ;
 wire \Tile_X3Y8_EE4BEG[2] ;
 wire \Tile_X3Y8_EE4BEG[3] ;
 wire \Tile_X3Y8_EE4BEG[4] ;
 wire \Tile_X3Y8_EE4BEG[5] ;
 wire \Tile_X3Y8_EE4BEG[6] ;
 wire \Tile_X3Y8_EE4BEG[7] ;
 wire \Tile_X3Y8_EE4BEG[8] ;
 wire \Tile_X3Y8_EE4BEG[9] ;
 wire \Tile_X3Y8_FrameData_O[0] ;
 wire \Tile_X3Y8_FrameData_O[10] ;
 wire \Tile_X3Y8_FrameData_O[11] ;
 wire \Tile_X3Y8_FrameData_O[12] ;
 wire \Tile_X3Y8_FrameData_O[13] ;
 wire \Tile_X3Y8_FrameData_O[14] ;
 wire \Tile_X3Y8_FrameData_O[15] ;
 wire \Tile_X3Y8_FrameData_O[16] ;
 wire \Tile_X3Y8_FrameData_O[17] ;
 wire \Tile_X3Y8_FrameData_O[18] ;
 wire \Tile_X3Y8_FrameData_O[19] ;
 wire \Tile_X3Y8_FrameData_O[1] ;
 wire \Tile_X3Y8_FrameData_O[20] ;
 wire \Tile_X3Y8_FrameData_O[21] ;
 wire \Tile_X3Y8_FrameData_O[22] ;
 wire \Tile_X3Y8_FrameData_O[23] ;
 wire \Tile_X3Y8_FrameData_O[24] ;
 wire \Tile_X3Y8_FrameData_O[25] ;
 wire \Tile_X3Y8_FrameData_O[26] ;
 wire \Tile_X3Y8_FrameData_O[27] ;
 wire \Tile_X3Y8_FrameData_O[28] ;
 wire \Tile_X3Y8_FrameData_O[29] ;
 wire \Tile_X3Y8_FrameData_O[2] ;
 wire \Tile_X3Y8_FrameData_O[30] ;
 wire \Tile_X3Y8_FrameData_O[31] ;
 wire \Tile_X3Y8_FrameData_O[3] ;
 wire \Tile_X3Y8_FrameData_O[4] ;
 wire \Tile_X3Y8_FrameData_O[5] ;
 wire \Tile_X3Y8_FrameData_O[6] ;
 wire \Tile_X3Y8_FrameData_O[7] ;
 wire \Tile_X3Y8_FrameData_O[8] ;
 wire \Tile_X3Y8_FrameData_O[9] ;
 wire \Tile_X3Y8_FrameStrobe_O[0] ;
 wire \Tile_X3Y8_FrameStrobe_O[10] ;
 wire \Tile_X3Y8_FrameStrobe_O[11] ;
 wire \Tile_X3Y8_FrameStrobe_O[12] ;
 wire \Tile_X3Y8_FrameStrobe_O[13] ;
 wire \Tile_X3Y8_FrameStrobe_O[14] ;
 wire \Tile_X3Y8_FrameStrobe_O[15] ;
 wire \Tile_X3Y8_FrameStrobe_O[16] ;
 wire \Tile_X3Y8_FrameStrobe_O[17] ;
 wire \Tile_X3Y8_FrameStrobe_O[18] ;
 wire \Tile_X3Y8_FrameStrobe_O[19] ;
 wire \Tile_X3Y8_FrameStrobe_O[1] ;
 wire \Tile_X3Y8_FrameStrobe_O[2] ;
 wire \Tile_X3Y8_FrameStrobe_O[3] ;
 wire \Tile_X3Y8_FrameStrobe_O[4] ;
 wire \Tile_X3Y8_FrameStrobe_O[5] ;
 wire \Tile_X3Y8_FrameStrobe_O[6] ;
 wire \Tile_X3Y8_FrameStrobe_O[7] ;
 wire \Tile_X3Y8_FrameStrobe_O[8] ;
 wire \Tile_X3Y8_FrameStrobe_O[9] ;
 wire \Tile_X3Y8_N1BEG[0] ;
 wire \Tile_X3Y8_N1BEG[1] ;
 wire \Tile_X3Y8_N1BEG[2] ;
 wire \Tile_X3Y8_N1BEG[3] ;
 wire \Tile_X3Y8_N2BEG[0] ;
 wire \Tile_X3Y8_N2BEG[1] ;
 wire \Tile_X3Y8_N2BEG[2] ;
 wire \Tile_X3Y8_N2BEG[3] ;
 wire \Tile_X3Y8_N2BEG[4] ;
 wire \Tile_X3Y8_N2BEG[5] ;
 wire \Tile_X3Y8_N2BEG[6] ;
 wire \Tile_X3Y8_N2BEG[7] ;
 wire \Tile_X3Y8_N2BEGb[0] ;
 wire \Tile_X3Y8_N2BEGb[1] ;
 wire \Tile_X3Y8_N2BEGb[2] ;
 wire \Tile_X3Y8_N2BEGb[3] ;
 wire \Tile_X3Y8_N2BEGb[4] ;
 wire \Tile_X3Y8_N2BEGb[5] ;
 wire \Tile_X3Y8_N2BEGb[6] ;
 wire \Tile_X3Y8_N2BEGb[7] ;
 wire \Tile_X3Y8_N4BEG[0] ;
 wire \Tile_X3Y8_N4BEG[10] ;
 wire \Tile_X3Y8_N4BEG[11] ;
 wire \Tile_X3Y8_N4BEG[12] ;
 wire \Tile_X3Y8_N4BEG[13] ;
 wire \Tile_X3Y8_N4BEG[14] ;
 wire \Tile_X3Y8_N4BEG[15] ;
 wire \Tile_X3Y8_N4BEG[1] ;
 wire \Tile_X3Y8_N4BEG[2] ;
 wire \Tile_X3Y8_N4BEG[3] ;
 wire \Tile_X3Y8_N4BEG[4] ;
 wire \Tile_X3Y8_N4BEG[5] ;
 wire \Tile_X3Y8_N4BEG[6] ;
 wire \Tile_X3Y8_N4BEG[7] ;
 wire \Tile_X3Y8_N4BEG[8] ;
 wire \Tile_X3Y8_N4BEG[9] ;
 wire \Tile_X3Y8_NN4BEG[0] ;
 wire \Tile_X3Y8_NN4BEG[10] ;
 wire \Tile_X3Y8_NN4BEG[11] ;
 wire \Tile_X3Y8_NN4BEG[12] ;
 wire \Tile_X3Y8_NN4BEG[13] ;
 wire \Tile_X3Y8_NN4BEG[14] ;
 wire \Tile_X3Y8_NN4BEG[15] ;
 wire \Tile_X3Y8_NN4BEG[1] ;
 wire \Tile_X3Y8_NN4BEG[2] ;
 wire \Tile_X3Y8_NN4BEG[3] ;
 wire \Tile_X3Y8_NN4BEG[4] ;
 wire \Tile_X3Y8_NN4BEG[5] ;
 wire \Tile_X3Y8_NN4BEG[6] ;
 wire \Tile_X3Y8_NN4BEG[7] ;
 wire \Tile_X3Y8_NN4BEG[8] ;
 wire \Tile_X3Y8_NN4BEG[9] ;
 wire \Tile_X3Y8_S1BEG[0] ;
 wire \Tile_X3Y8_S1BEG[1] ;
 wire \Tile_X3Y8_S1BEG[2] ;
 wire \Tile_X3Y8_S1BEG[3] ;
 wire \Tile_X3Y8_S2BEG[0] ;
 wire \Tile_X3Y8_S2BEG[1] ;
 wire \Tile_X3Y8_S2BEG[2] ;
 wire \Tile_X3Y8_S2BEG[3] ;
 wire \Tile_X3Y8_S2BEG[4] ;
 wire \Tile_X3Y8_S2BEG[5] ;
 wire \Tile_X3Y8_S2BEG[6] ;
 wire \Tile_X3Y8_S2BEG[7] ;
 wire \Tile_X3Y8_S2BEGb[0] ;
 wire \Tile_X3Y8_S2BEGb[1] ;
 wire \Tile_X3Y8_S2BEGb[2] ;
 wire \Tile_X3Y8_S2BEGb[3] ;
 wire \Tile_X3Y8_S2BEGb[4] ;
 wire \Tile_X3Y8_S2BEGb[5] ;
 wire \Tile_X3Y8_S2BEGb[6] ;
 wire \Tile_X3Y8_S2BEGb[7] ;
 wire \Tile_X3Y8_S4BEG[0] ;
 wire \Tile_X3Y8_S4BEG[10] ;
 wire \Tile_X3Y8_S4BEG[11] ;
 wire \Tile_X3Y8_S4BEG[12] ;
 wire \Tile_X3Y8_S4BEG[13] ;
 wire \Tile_X3Y8_S4BEG[14] ;
 wire \Tile_X3Y8_S4BEG[15] ;
 wire \Tile_X3Y8_S4BEG[1] ;
 wire \Tile_X3Y8_S4BEG[2] ;
 wire \Tile_X3Y8_S4BEG[3] ;
 wire \Tile_X3Y8_S4BEG[4] ;
 wire \Tile_X3Y8_S4BEG[5] ;
 wire \Tile_X3Y8_S4BEG[6] ;
 wire \Tile_X3Y8_S4BEG[7] ;
 wire \Tile_X3Y8_S4BEG[8] ;
 wire \Tile_X3Y8_S4BEG[9] ;
 wire \Tile_X3Y8_SS4BEG[0] ;
 wire \Tile_X3Y8_SS4BEG[10] ;
 wire \Tile_X3Y8_SS4BEG[11] ;
 wire \Tile_X3Y8_SS4BEG[12] ;
 wire \Tile_X3Y8_SS4BEG[13] ;
 wire \Tile_X3Y8_SS4BEG[14] ;
 wire \Tile_X3Y8_SS4BEG[15] ;
 wire \Tile_X3Y8_SS4BEG[1] ;
 wire \Tile_X3Y8_SS4BEG[2] ;
 wire \Tile_X3Y8_SS4BEG[3] ;
 wire \Tile_X3Y8_SS4BEG[4] ;
 wire \Tile_X3Y8_SS4BEG[5] ;
 wire \Tile_X3Y8_SS4BEG[6] ;
 wire \Tile_X3Y8_SS4BEG[7] ;
 wire \Tile_X3Y8_SS4BEG[8] ;
 wire \Tile_X3Y8_SS4BEG[9] ;
 wire Tile_X3Y8_UserCLKo;
 wire \Tile_X3Y8_W1BEG[0] ;
 wire \Tile_X3Y8_W1BEG[1] ;
 wire \Tile_X3Y8_W1BEG[2] ;
 wire \Tile_X3Y8_W1BEG[3] ;
 wire \Tile_X3Y8_W2BEG[0] ;
 wire \Tile_X3Y8_W2BEG[1] ;
 wire \Tile_X3Y8_W2BEG[2] ;
 wire \Tile_X3Y8_W2BEG[3] ;
 wire \Tile_X3Y8_W2BEG[4] ;
 wire \Tile_X3Y8_W2BEG[5] ;
 wire \Tile_X3Y8_W2BEG[6] ;
 wire \Tile_X3Y8_W2BEG[7] ;
 wire \Tile_X3Y8_W2BEGb[0] ;
 wire \Tile_X3Y8_W2BEGb[1] ;
 wire \Tile_X3Y8_W2BEGb[2] ;
 wire \Tile_X3Y8_W2BEGb[3] ;
 wire \Tile_X3Y8_W2BEGb[4] ;
 wire \Tile_X3Y8_W2BEGb[5] ;
 wire \Tile_X3Y8_W2BEGb[6] ;
 wire \Tile_X3Y8_W2BEGb[7] ;
 wire \Tile_X3Y8_W6BEG[0] ;
 wire \Tile_X3Y8_W6BEG[10] ;
 wire \Tile_X3Y8_W6BEG[11] ;
 wire \Tile_X3Y8_W6BEG[1] ;
 wire \Tile_X3Y8_W6BEG[2] ;
 wire \Tile_X3Y8_W6BEG[3] ;
 wire \Tile_X3Y8_W6BEG[4] ;
 wire \Tile_X3Y8_W6BEG[5] ;
 wire \Tile_X3Y8_W6BEG[6] ;
 wire \Tile_X3Y8_W6BEG[7] ;
 wire \Tile_X3Y8_W6BEG[8] ;
 wire \Tile_X3Y8_W6BEG[9] ;
 wire \Tile_X3Y8_WW4BEG[0] ;
 wire \Tile_X3Y8_WW4BEG[10] ;
 wire \Tile_X3Y8_WW4BEG[11] ;
 wire \Tile_X3Y8_WW4BEG[12] ;
 wire \Tile_X3Y8_WW4BEG[13] ;
 wire \Tile_X3Y8_WW4BEG[14] ;
 wire \Tile_X3Y8_WW4BEG[15] ;
 wire \Tile_X3Y8_WW4BEG[1] ;
 wire \Tile_X3Y8_WW4BEG[2] ;
 wire \Tile_X3Y8_WW4BEG[3] ;
 wire \Tile_X3Y8_WW4BEG[4] ;
 wire \Tile_X3Y8_WW4BEG[5] ;
 wire \Tile_X3Y8_WW4BEG[6] ;
 wire \Tile_X3Y8_WW4BEG[7] ;
 wire \Tile_X3Y8_WW4BEG[8] ;
 wire \Tile_X3Y8_WW4BEG[9] ;
 wire Tile_X3Y9_Co;
 wire \Tile_X3Y9_E1BEG[0] ;
 wire \Tile_X3Y9_E1BEG[1] ;
 wire \Tile_X3Y9_E1BEG[2] ;
 wire \Tile_X3Y9_E1BEG[3] ;
 wire \Tile_X3Y9_E2BEG[0] ;
 wire \Tile_X3Y9_E2BEG[1] ;
 wire \Tile_X3Y9_E2BEG[2] ;
 wire \Tile_X3Y9_E2BEG[3] ;
 wire \Tile_X3Y9_E2BEG[4] ;
 wire \Tile_X3Y9_E2BEG[5] ;
 wire \Tile_X3Y9_E2BEG[6] ;
 wire \Tile_X3Y9_E2BEG[7] ;
 wire \Tile_X3Y9_E2BEGb[0] ;
 wire \Tile_X3Y9_E2BEGb[1] ;
 wire \Tile_X3Y9_E2BEGb[2] ;
 wire \Tile_X3Y9_E2BEGb[3] ;
 wire \Tile_X3Y9_E2BEGb[4] ;
 wire \Tile_X3Y9_E2BEGb[5] ;
 wire \Tile_X3Y9_E2BEGb[6] ;
 wire \Tile_X3Y9_E2BEGb[7] ;
 wire \Tile_X3Y9_E6BEG[0] ;
 wire \Tile_X3Y9_E6BEG[10] ;
 wire \Tile_X3Y9_E6BEG[11] ;
 wire \Tile_X3Y9_E6BEG[1] ;
 wire \Tile_X3Y9_E6BEG[2] ;
 wire \Tile_X3Y9_E6BEG[3] ;
 wire \Tile_X3Y9_E6BEG[4] ;
 wire \Tile_X3Y9_E6BEG[5] ;
 wire \Tile_X3Y9_E6BEG[6] ;
 wire \Tile_X3Y9_E6BEG[7] ;
 wire \Tile_X3Y9_E6BEG[8] ;
 wire \Tile_X3Y9_E6BEG[9] ;
 wire \Tile_X3Y9_EE4BEG[0] ;
 wire \Tile_X3Y9_EE4BEG[10] ;
 wire \Tile_X3Y9_EE4BEG[11] ;
 wire \Tile_X3Y9_EE4BEG[12] ;
 wire \Tile_X3Y9_EE4BEG[13] ;
 wire \Tile_X3Y9_EE4BEG[14] ;
 wire \Tile_X3Y9_EE4BEG[15] ;
 wire \Tile_X3Y9_EE4BEG[1] ;
 wire \Tile_X3Y9_EE4BEG[2] ;
 wire \Tile_X3Y9_EE4BEG[3] ;
 wire \Tile_X3Y9_EE4BEG[4] ;
 wire \Tile_X3Y9_EE4BEG[5] ;
 wire \Tile_X3Y9_EE4BEG[6] ;
 wire \Tile_X3Y9_EE4BEG[7] ;
 wire \Tile_X3Y9_EE4BEG[8] ;
 wire \Tile_X3Y9_EE4BEG[9] ;
 wire \Tile_X3Y9_FrameData_O[0] ;
 wire \Tile_X3Y9_FrameData_O[10] ;
 wire \Tile_X3Y9_FrameData_O[11] ;
 wire \Tile_X3Y9_FrameData_O[12] ;
 wire \Tile_X3Y9_FrameData_O[13] ;
 wire \Tile_X3Y9_FrameData_O[14] ;
 wire \Tile_X3Y9_FrameData_O[15] ;
 wire \Tile_X3Y9_FrameData_O[16] ;
 wire \Tile_X3Y9_FrameData_O[17] ;
 wire \Tile_X3Y9_FrameData_O[18] ;
 wire \Tile_X3Y9_FrameData_O[19] ;
 wire \Tile_X3Y9_FrameData_O[1] ;
 wire \Tile_X3Y9_FrameData_O[20] ;
 wire \Tile_X3Y9_FrameData_O[21] ;
 wire \Tile_X3Y9_FrameData_O[22] ;
 wire \Tile_X3Y9_FrameData_O[23] ;
 wire \Tile_X3Y9_FrameData_O[24] ;
 wire \Tile_X3Y9_FrameData_O[25] ;
 wire \Tile_X3Y9_FrameData_O[26] ;
 wire \Tile_X3Y9_FrameData_O[27] ;
 wire \Tile_X3Y9_FrameData_O[28] ;
 wire \Tile_X3Y9_FrameData_O[29] ;
 wire \Tile_X3Y9_FrameData_O[2] ;
 wire \Tile_X3Y9_FrameData_O[30] ;
 wire \Tile_X3Y9_FrameData_O[31] ;
 wire \Tile_X3Y9_FrameData_O[3] ;
 wire \Tile_X3Y9_FrameData_O[4] ;
 wire \Tile_X3Y9_FrameData_O[5] ;
 wire \Tile_X3Y9_FrameData_O[6] ;
 wire \Tile_X3Y9_FrameData_O[7] ;
 wire \Tile_X3Y9_FrameData_O[8] ;
 wire \Tile_X3Y9_FrameData_O[9] ;
 wire \Tile_X3Y9_FrameStrobe_O[0] ;
 wire \Tile_X3Y9_FrameStrobe_O[10] ;
 wire \Tile_X3Y9_FrameStrobe_O[11] ;
 wire \Tile_X3Y9_FrameStrobe_O[12] ;
 wire \Tile_X3Y9_FrameStrobe_O[13] ;
 wire \Tile_X3Y9_FrameStrobe_O[14] ;
 wire \Tile_X3Y9_FrameStrobe_O[15] ;
 wire \Tile_X3Y9_FrameStrobe_O[16] ;
 wire \Tile_X3Y9_FrameStrobe_O[17] ;
 wire \Tile_X3Y9_FrameStrobe_O[18] ;
 wire \Tile_X3Y9_FrameStrobe_O[19] ;
 wire \Tile_X3Y9_FrameStrobe_O[1] ;
 wire \Tile_X3Y9_FrameStrobe_O[2] ;
 wire \Tile_X3Y9_FrameStrobe_O[3] ;
 wire \Tile_X3Y9_FrameStrobe_O[4] ;
 wire \Tile_X3Y9_FrameStrobe_O[5] ;
 wire \Tile_X3Y9_FrameStrobe_O[6] ;
 wire \Tile_X3Y9_FrameStrobe_O[7] ;
 wire \Tile_X3Y9_FrameStrobe_O[8] ;
 wire \Tile_X3Y9_FrameStrobe_O[9] ;
 wire \Tile_X3Y9_N1BEG[0] ;
 wire \Tile_X3Y9_N1BEG[1] ;
 wire \Tile_X3Y9_N1BEG[2] ;
 wire \Tile_X3Y9_N1BEG[3] ;
 wire \Tile_X3Y9_N2BEG[0] ;
 wire \Tile_X3Y9_N2BEG[1] ;
 wire \Tile_X3Y9_N2BEG[2] ;
 wire \Tile_X3Y9_N2BEG[3] ;
 wire \Tile_X3Y9_N2BEG[4] ;
 wire \Tile_X3Y9_N2BEG[5] ;
 wire \Tile_X3Y9_N2BEG[6] ;
 wire \Tile_X3Y9_N2BEG[7] ;
 wire \Tile_X3Y9_N2BEGb[0] ;
 wire \Tile_X3Y9_N2BEGb[1] ;
 wire \Tile_X3Y9_N2BEGb[2] ;
 wire \Tile_X3Y9_N2BEGb[3] ;
 wire \Tile_X3Y9_N2BEGb[4] ;
 wire \Tile_X3Y9_N2BEGb[5] ;
 wire \Tile_X3Y9_N2BEGb[6] ;
 wire \Tile_X3Y9_N2BEGb[7] ;
 wire \Tile_X3Y9_N4BEG[0] ;
 wire \Tile_X3Y9_N4BEG[10] ;
 wire \Tile_X3Y9_N4BEG[11] ;
 wire \Tile_X3Y9_N4BEG[12] ;
 wire \Tile_X3Y9_N4BEG[13] ;
 wire \Tile_X3Y9_N4BEG[14] ;
 wire \Tile_X3Y9_N4BEG[15] ;
 wire \Tile_X3Y9_N4BEG[1] ;
 wire \Tile_X3Y9_N4BEG[2] ;
 wire \Tile_X3Y9_N4BEG[3] ;
 wire \Tile_X3Y9_N4BEG[4] ;
 wire \Tile_X3Y9_N4BEG[5] ;
 wire \Tile_X3Y9_N4BEG[6] ;
 wire \Tile_X3Y9_N4BEG[7] ;
 wire \Tile_X3Y9_N4BEG[8] ;
 wire \Tile_X3Y9_N4BEG[9] ;
 wire \Tile_X3Y9_NN4BEG[0] ;
 wire \Tile_X3Y9_NN4BEG[10] ;
 wire \Tile_X3Y9_NN4BEG[11] ;
 wire \Tile_X3Y9_NN4BEG[12] ;
 wire \Tile_X3Y9_NN4BEG[13] ;
 wire \Tile_X3Y9_NN4BEG[14] ;
 wire \Tile_X3Y9_NN4BEG[15] ;
 wire \Tile_X3Y9_NN4BEG[1] ;
 wire \Tile_X3Y9_NN4BEG[2] ;
 wire \Tile_X3Y9_NN4BEG[3] ;
 wire \Tile_X3Y9_NN4BEG[4] ;
 wire \Tile_X3Y9_NN4BEG[5] ;
 wire \Tile_X3Y9_NN4BEG[6] ;
 wire \Tile_X3Y9_NN4BEG[7] ;
 wire \Tile_X3Y9_NN4BEG[8] ;
 wire \Tile_X3Y9_NN4BEG[9] ;
 wire \Tile_X3Y9_S1BEG[0] ;
 wire \Tile_X3Y9_S1BEG[1] ;
 wire \Tile_X3Y9_S1BEG[2] ;
 wire \Tile_X3Y9_S1BEG[3] ;
 wire \Tile_X3Y9_S2BEG[0] ;
 wire \Tile_X3Y9_S2BEG[1] ;
 wire \Tile_X3Y9_S2BEG[2] ;
 wire \Tile_X3Y9_S2BEG[3] ;
 wire \Tile_X3Y9_S2BEG[4] ;
 wire \Tile_X3Y9_S2BEG[5] ;
 wire \Tile_X3Y9_S2BEG[6] ;
 wire \Tile_X3Y9_S2BEG[7] ;
 wire \Tile_X3Y9_S2BEGb[0] ;
 wire \Tile_X3Y9_S2BEGb[1] ;
 wire \Tile_X3Y9_S2BEGb[2] ;
 wire \Tile_X3Y9_S2BEGb[3] ;
 wire \Tile_X3Y9_S2BEGb[4] ;
 wire \Tile_X3Y9_S2BEGb[5] ;
 wire \Tile_X3Y9_S2BEGb[6] ;
 wire \Tile_X3Y9_S2BEGb[7] ;
 wire \Tile_X3Y9_S4BEG[0] ;
 wire \Tile_X3Y9_S4BEG[10] ;
 wire \Tile_X3Y9_S4BEG[11] ;
 wire \Tile_X3Y9_S4BEG[12] ;
 wire \Tile_X3Y9_S4BEG[13] ;
 wire \Tile_X3Y9_S4BEG[14] ;
 wire \Tile_X3Y9_S4BEG[15] ;
 wire \Tile_X3Y9_S4BEG[1] ;
 wire \Tile_X3Y9_S4BEG[2] ;
 wire \Tile_X3Y9_S4BEG[3] ;
 wire \Tile_X3Y9_S4BEG[4] ;
 wire \Tile_X3Y9_S4BEG[5] ;
 wire \Tile_X3Y9_S4BEG[6] ;
 wire \Tile_X3Y9_S4BEG[7] ;
 wire \Tile_X3Y9_S4BEG[8] ;
 wire \Tile_X3Y9_S4BEG[9] ;
 wire \Tile_X3Y9_SS4BEG[0] ;
 wire \Tile_X3Y9_SS4BEG[10] ;
 wire \Tile_X3Y9_SS4BEG[11] ;
 wire \Tile_X3Y9_SS4BEG[12] ;
 wire \Tile_X3Y9_SS4BEG[13] ;
 wire \Tile_X3Y9_SS4BEG[14] ;
 wire \Tile_X3Y9_SS4BEG[15] ;
 wire \Tile_X3Y9_SS4BEG[1] ;
 wire \Tile_X3Y9_SS4BEG[2] ;
 wire \Tile_X3Y9_SS4BEG[3] ;
 wire \Tile_X3Y9_SS4BEG[4] ;
 wire \Tile_X3Y9_SS4BEG[5] ;
 wire \Tile_X3Y9_SS4BEG[6] ;
 wire \Tile_X3Y9_SS4BEG[7] ;
 wire \Tile_X3Y9_SS4BEG[8] ;
 wire \Tile_X3Y9_SS4BEG[9] ;
 wire Tile_X3Y9_UserCLKo;
 wire \Tile_X3Y9_W1BEG[0] ;
 wire \Tile_X3Y9_W1BEG[1] ;
 wire \Tile_X3Y9_W1BEG[2] ;
 wire \Tile_X3Y9_W1BEG[3] ;
 wire \Tile_X3Y9_W2BEG[0] ;
 wire \Tile_X3Y9_W2BEG[1] ;
 wire \Tile_X3Y9_W2BEG[2] ;
 wire \Tile_X3Y9_W2BEG[3] ;
 wire \Tile_X3Y9_W2BEG[4] ;
 wire \Tile_X3Y9_W2BEG[5] ;
 wire \Tile_X3Y9_W2BEG[6] ;
 wire \Tile_X3Y9_W2BEG[7] ;
 wire \Tile_X3Y9_W2BEGb[0] ;
 wire \Tile_X3Y9_W2BEGb[1] ;
 wire \Tile_X3Y9_W2BEGb[2] ;
 wire \Tile_X3Y9_W2BEGb[3] ;
 wire \Tile_X3Y9_W2BEGb[4] ;
 wire \Tile_X3Y9_W2BEGb[5] ;
 wire \Tile_X3Y9_W2BEGb[6] ;
 wire \Tile_X3Y9_W2BEGb[7] ;
 wire \Tile_X3Y9_W6BEG[0] ;
 wire \Tile_X3Y9_W6BEG[10] ;
 wire \Tile_X3Y9_W6BEG[11] ;
 wire \Tile_X3Y9_W6BEG[1] ;
 wire \Tile_X3Y9_W6BEG[2] ;
 wire \Tile_X3Y9_W6BEG[3] ;
 wire \Tile_X3Y9_W6BEG[4] ;
 wire \Tile_X3Y9_W6BEG[5] ;
 wire \Tile_X3Y9_W6BEG[6] ;
 wire \Tile_X3Y9_W6BEG[7] ;
 wire \Tile_X3Y9_W6BEG[8] ;
 wire \Tile_X3Y9_W6BEG[9] ;
 wire \Tile_X3Y9_WW4BEG[0] ;
 wire \Tile_X3Y9_WW4BEG[10] ;
 wire \Tile_X3Y9_WW4BEG[11] ;
 wire \Tile_X3Y9_WW4BEG[12] ;
 wire \Tile_X3Y9_WW4BEG[13] ;
 wire \Tile_X3Y9_WW4BEG[14] ;
 wire \Tile_X3Y9_WW4BEG[15] ;
 wire \Tile_X3Y9_WW4BEG[1] ;
 wire \Tile_X3Y9_WW4BEG[2] ;
 wire \Tile_X3Y9_WW4BEG[3] ;
 wire \Tile_X3Y9_WW4BEG[4] ;
 wire \Tile_X3Y9_WW4BEG[5] ;
 wire \Tile_X3Y9_WW4BEG[6] ;
 wire \Tile_X3Y9_WW4BEG[7] ;
 wire \Tile_X3Y9_WW4BEG[8] ;
 wire \Tile_X3Y9_WW4BEG[9] ;
 wire \Tile_X4Y0_FrameData_O[0] ;
 wire \Tile_X4Y0_FrameData_O[10] ;
 wire \Tile_X4Y0_FrameData_O[11] ;
 wire \Tile_X4Y0_FrameData_O[12] ;
 wire \Tile_X4Y0_FrameData_O[13] ;
 wire \Tile_X4Y0_FrameData_O[14] ;
 wire \Tile_X4Y0_FrameData_O[15] ;
 wire \Tile_X4Y0_FrameData_O[16] ;
 wire \Tile_X4Y0_FrameData_O[17] ;
 wire \Tile_X4Y0_FrameData_O[18] ;
 wire \Tile_X4Y0_FrameData_O[19] ;
 wire \Tile_X4Y0_FrameData_O[1] ;
 wire \Tile_X4Y0_FrameData_O[20] ;
 wire \Tile_X4Y0_FrameData_O[21] ;
 wire \Tile_X4Y0_FrameData_O[22] ;
 wire \Tile_X4Y0_FrameData_O[23] ;
 wire \Tile_X4Y0_FrameData_O[24] ;
 wire \Tile_X4Y0_FrameData_O[25] ;
 wire \Tile_X4Y0_FrameData_O[26] ;
 wire \Tile_X4Y0_FrameData_O[27] ;
 wire \Tile_X4Y0_FrameData_O[28] ;
 wire \Tile_X4Y0_FrameData_O[29] ;
 wire \Tile_X4Y0_FrameData_O[2] ;
 wire \Tile_X4Y0_FrameData_O[30] ;
 wire \Tile_X4Y0_FrameData_O[31] ;
 wire \Tile_X4Y0_FrameData_O[3] ;
 wire \Tile_X4Y0_FrameData_O[4] ;
 wire \Tile_X4Y0_FrameData_O[5] ;
 wire \Tile_X4Y0_FrameData_O[6] ;
 wire \Tile_X4Y0_FrameData_O[7] ;
 wire \Tile_X4Y0_FrameData_O[8] ;
 wire \Tile_X4Y0_FrameData_O[9] ;
 wire \Tile_X4Y0_FrameStrobe_O[0] ;
 wire \Tile_X4Y0_FrameStrobe_O[10] ;
 wire \Tile_X4Y0_FrameStrobe_O[11] ;
 wire \Tile_X4Y0_FrameStrobe_O[12] ;
 wire \Tile_X4Y0_FrameStrobe_O[13] ;
 wire \Tile_X4Y0_FrameStrobe_O[14] ;
 wire \Tile_X4Y0_FrameStrobe_O[15] ;
 wire \Tile_X4Y0_FrameStrobe_O[16] ;
 wire \Tile_X4Y0_FrameStrobe_O[17] ;
 wire \Tile_X4Y0_FrameStrobe_O[18] ;
 wire \Tile_X4Y0_FrameStrobe_O[19] ;
 wire \Tile_X4Y0_FrameStrobe_O[1] ;
 wire \Tile_X4Y0_FrameStrobe_O[2] ;
 wire \Tile_X4Y0_FrameStrobe_O[3] ;
 wire \Tile_X4Y0_FrameStrobe_O[4] ;
 wire \Tile_X4Y0_FrameStrobe_O[5] ;
 wire \Tile_X4Y0_FrameStrobe_O[6] ;
 wire \Tile_X4Y0_FrameStrobe_O[7] ;
 wire \Tile_X4Y0_FrameStrobe_O[8] ;
 wire \Tile_X4Y0_FrameStrobe_O[9] ;
 wire \Tile_X4Y0_S1BEG[0] ;
 wire \Tile_X4Y0_S1BEG[1] ;
 wire \Tile_X4Y0_S1BEG[2] ;
 wire \Tile_X4Y0_S1BEG[3] ;
 wire \Tile_X4Y0_S2BEG[0] ;
 wire \Tile_X4Y0_S2BEG[1] ;
 wire \Tile_X4Y0_S2BEG[2] ;
 wire \Tile_X4Y0_S2BEG[3] ;
 wire \Tile_X4Y0_S2BEG[4] ;
 wire \Tile_X4Y0_S2BEG[5] ;
 wire \Tile_X4Y0_S2BEG[6] ;
 wire \Tile_X4Y0_S2BEG[7] ;
 wire \Tile_X4Y0_S2BEGb[0] ;
 wire \Tile_X4Y0_S2BEGb[1] ;
 wire \Tile_X4Y0_S2BEGb[2] ;
 wire \Tile_X4Y0_S2BEGb[3] ;
 wire \Tile_X4Y0_S2BEGb[4] ;
 wire \Tile_X4Y0_S2BEGb[5] ;
 wire \Tile_X4Y0_S2BEGb[6] ;
 wire \Tile_X4Y0_S2BEGb[7] ;
 wire \Tile_X4Y0_S4BEG[0] ;
 wire \Tile_X4Y0_S4BEG[10] ;
 wire \Tile_X4Y0_S4BEG[11] ;
 wire \Tile_X4Y0_S4BEG[12] ;
 wire \Tile_X4Y0_S4BEG[13] ;
 wire \Tile_X4Y0_S4BEG[14] ;
 wire \Tile_X4Y0_S4BEG[15] ;
 wire \Tile_X4Y0_S4BEG[1] ;
 wire \Tile_X4Y0_S4BEG[2] ;
 wire \Tile_X4Y0_S4BEG[3] ;
 wire \Tile_X4Y0_S4BEG[4] ;
 wire \Tile_X4Y0_S4BEG[5] ;
 wire \Tile_X4Y0_S4BEG[6] ;
 wire \Tile_X4Y0_S4BEG[7] ;
 wire \Tile_X4Y0_S4BEG[8] ;
 wire \Tile_X4Y0_S4BEG[9] ;
 wire \Tile_X4Y0_SS4BEG[0] ;
 wire \Tile_X4Y0_SS4BEG[10] ;
 wire \Tile_X4Y0_SS4BEG[11] ;
 wire \Tile_X4Y0_SS4BEG[12] ;
 wire \Tile_X4Y0_SS4BEG[13] ;
 wire \Tile_X4Y0_SS4BEG[14] ;
 wire \Tile_X4Y0_SS4BEG[15] ;
 wire \Tile_X4Y0_SS4BEG[1] ;
 wire \Tile_X4Y0_SS4BEG[2] ;
 wire \Tile_X4Y0_SS4BEG[3] ;
 wire \Tile_X4Y0_SS4BEG[4] ;
 wire \Tile_X4Y0_SS4BEG[5] ;
 wire \Tile_X4Y0_SS4BEG[6] ;
 wire \Tile_X4Y0_SS4BEG[7] ;
 wire \Tile_X4Y0_SS4BEG[8] ;
 wire \Tile_X4Y0_SS4BEG[9] ;
 wire Tile_X4Y0_UserCLKo;
 wire \Tile_X4Y10_E1BEG[0] ;
 wire \Tile_X4Y10_E1BEG[1] ;
 wire \Tile_X4Y10_E1BEG[2] ;
 wire \Tile_X4Y10_E1BEG[3] ;
 wire \Tile_X4Y10_E2BEG[0] ;
 wire \Tile_X4Y10_E2BEG[1] ;
 wire \Tile_X4Y10_E2BEG[2] ;
 wire \Tile_X4Y10_E2BEG[3] ;
 wire \Tile_X4Y10_E2BEG[4] ;
 wire \Tile_X4Y10_E2BEG[5] ;
 wire \Tile_X4Y10_E2BEG[6] ;
 wire \Tile_X4Y10_E2BEG[7] ;
 wire \Tile_X4Y10_E2BEGb[0] ;
 wire \Tile_X4Y10_E2BEGb[1] ;
 wire \Tile_X4Y10_E2BEGb[2] ;
 wire \Tile_X4Y10_E2BEGb[3] ;
 wire \Tile_X4Y10_E2BEGb[4] ;
 wire \Tile_X4Y10_E2BEGb[5] ;
 wire \Tile_X4Y10_E2BEGb[6] ;
 wire \Tile_X4Y10_E2BEGb[7] ;
 wire \Tile_X4Y10_E6BEG[0] ;
 wire \Tile_X4Y10_E6BEG[10] ;
 wire \Tile_X4Y10_E6BEG[11] ;
 wire \Tile_X4Y10_E6BEG[1] ;
 wire \Tile_X4Y10_E6BEG[2] ;
 wire \Tile_X4Y10_E6BEG[3] ;
 wire \Tile_X4Y10_E6BEG[4] ;
 wire \Tile_X4Y10_E6BEG[5] ;
 wire \Tile_X4Y10_E6BEG[6] ;
 wire \Tile_X4Y10_E6BEG[7] ;
 wire \Tile_X4Y10_E6BEG[8] ;
 wire \Tile_X4Y10_E6BEG[9] ;
 wire \Tile_X4Y10_EE4BEG[0] ;
 wire \Tile_X4Y10_EE4BEG[10] ;
 wire \Tile_X4Y10_EE4BEG[11] ;
 wire \Tile_X4Y10_EE4BEG[12] ;
 wire \Tile_X4Y10_EE4BEG[13] ;
 wire \Tile_X4Y10_EE4BEG[14] ;
 wire \Tile_X4Y10_EE4BEG[15] ;
 wire \Tile_X4Y10_EE4BEG[1] ;
 wire \Tile_X4Y10_EE4BEG[2] ;
 wire \Tile_X4Y10_EE4BEG[3] ;
 wire \Tile_X4Y10_EE4BEG[4] ;
 wire \Tile_X4Y10_EE4BEG[5] ;
 wire \Tile_X4Y10_EE4BEG[6] ;
 wire \Tile_X4Y10_EE4BEG[7] ;
 wire \Tile_X4Y10_EE4BEG[8] ;
 wire \Tile_X4Y10_EE4BEG[9] ;
 wire \Tile_X4Y10_FrameData_O[0] ;
 wire \Tile_X4Y10_FrameData_O[10] ;
 wire \Tile_X4Y10_FrameData_O[11] ;
 wire \Tile_X4Y10_FrameData_O[12] ;
 wire \Tile_X4Y10_FrameData_O[13] ;
 wire \Tile_X4Y10_FrameData_O[14] ;
 wire \Tile_X4Y10_FrameData_O[15] ;
 wire \Tile_X4Y10_FrameData_O[16] ;
 wire \Tile_X4Y10_FrameData_O[17] ;
 wire \Tile_X4Y10_FrameData_O[18] ;
 wire \Tile_X4Y10_FrameData_O[19] ;
 wire \Tile_X4Y10_FrameData_O[1] ;
 wire \Tile_X4Y10_FrameData_O[20] ;
 wire \Tile_X4Y10_FrameData_O[21] ;
 wire \Tile_X4Y10_FrameData_O[22] ;
 wire \Tile_X4Y10_FrameData_O[23] ;
 wire \Tile_X4Y10_FrameData_O[24] ;
 wire \Tile_X4Y10_FrameData_O[25] ;
 wire \Tile_X4Y10_FrameData_O[26] ;
 wire \Tile_X4Y10_FrameData_O[27] ;
 wire \Tile_X4Y10_FrameData_O[28] ;
 wire \Tile_X4Y10_FrameData_O[29] ;
 wire \Tile_X4Y10_FrameData_O[2] ;
 wire \Tile_X4Y10_FrameData_O[30] ;
 wire \Tile_X4Y10_FrameData_O[31] ;
 wire \Tile_X4Y10_FrameData_O[3] ;
 wire \Tile_X4Y10_FrameData_O[4] ;
 wire \Tile_X4Y10_FrameData_O[5] ;
 wire \Tile_X4Y10_FrameData_O[6] ;
 wire \Tile_X4Y10_FrameData_O[7] ;
 wire \Tile_X4Y10_FrameData_O[8] ;
 wire \Tile_X4Y10_FrameData_O[9] ;
 wire \Tile_X4Y10_FrameStrobe_O[0] ;
 wire \Tile_X4Y10_FrameStrobe_O[10] ;
 wire \Tile_X4Y10_FrameStrobe_O[11] ;
 wire \Tile_X4Y10_FrameStrobe_O[12] ;
 wire \Tile_X4Y10_FrameStrobe_O[13] ;
 wire \Tile_X4Y10_FrameStrobe_O[14] ;
 wire \Tile_X4Y10_FrameStrobe_O[15] ;
 wire \Tile_X4Y10_FrameStrobe_O[16] ;
 wire \Tile_X4Y10_FrameStrobe_O[17] ;
 wire \Tile_X4Y10_FrameStrobe_O[18] ;
 wire \Tile_X4Y10_FrameStrobe_O[19] ;
 wire \Tile_X4Y10_FrameStrobe_O[1] ;
 wire \Tile_X4Y10_FrameStrobe_O[2] ;
 wire \Tile_X4Y10_FrameStrobe_O[3] ;
 wire \Tile_X4Y10_FrameStrobe_O[4] ;
 wire \Tile_X4Y10_FrameStrobe_O[5] ;
 wire \Tile_X4Y10_FrameStrobe_O[6] ;
 wire \Tile_X4Y10_FrameStrobe_O[7] ;
 wire \Tile_X4Y10_FrameStrobe_O[8] ;
 wire \Tile_X4Y10_FrameStrobe_O[9] ;
 wire \Tile_X4Y10_N1BEG[0] ;
 wire \Tile_X4Y10_N1BEG[1] ;
 wire \Tile_X4Y10_N1BEG[2] ;
 wire \Tile_X4Y10_N1BEG[3] ;
 wire \Tile_X4Y10_N2BEG[0] ;
 wire \Tile_X4Y10_N2BEG[1] ;
 wire \Tile_X4Y10_N2BEG[2] ;
 wire \Tile_X4Y10_N2BEG[3] ;
 wire \Tile_X4Y10_N2BEG[4] ;
 wire \Tile_X4Y10_N2BEG[5] ;
 wire \Tile_X4Y10_N2BEG[6] ;
 wire \Tile_X4Y10_N2BEG[7] ;
 wire \Tile_X4Y10_N2BEGb[0] ;
 wire \Tile_X4Y10_N2BEGb[1] ;
 wire \Tile_X4Y10_N2BEGb[2] ;
 wire \Tile_X4Y10_N2BEGb[3] ;
 wire \Tile_X4Y10_N2BEGb[4] ;
 wire \Tile_X4Y10_N2BEGb[5] ;
 wire \Tile_X4Y10_N2BEGb[6] ;
 wire \Tile_X4Y10_N2BEGb[7] ;
 wire \Tile_X4Y10_N4BEG[0] ;
 wire \Tile_X4Y10_N4BEG[10] ;
 wire \Tile_X4Y10_N4BEG[11] ;
 wire \Tile_X4Y10_N4BEG[12] ;
 wire \Tile_X4Y10_N4BEG[13] ;
 wire \Tile_X4Y10_N4BEG[14] ;
 wire \Tile_X4Y10_N4BEG[15] ;
 wire \Tile_X4Y10_N4BEG[1] ;
 wire \Tile_X4Y10_N4BEG[2] ;
 wire \Tile_X4Y10_N4BEG[3] ;
 wire \Tile_X4Y10_N4BEG[4] ;
 wire \Tile_X4Y10_N4BEG[5] ;
 wire \Tile_X4Y10_N4BEG[6] ;
 wire \Tile_X4Y10_N4BEG[7] ;
 wire \Tile_X4Y10_N4BEG[8] ;
 wire \Tile_X4Y10_N4BEG[9] ;
 wire \Tile_X4Y10_NN4BEG[0] ;
 wire \Tile_X4Y10_NN4BEG[10] ;
 wire \Tile_X4Y10_NN4BEG[11] ;
 wire \Tile_X4Y10_NN4BEG[12] ;
 wire \Tile_X4Y10_NN4BEG[13] ;
 wire \Tile_X4Y10_NN4BEG[14] ;
 wire \Tile_X4Y10_NN4BEG[15] ;
 wire \Tile_X4Y10_NN4BEG[1] ;
 wire \Tile_X4Y10_NN4BEG[2] ;
 wire \Tile_X4Y10_NN4BEG[3] ;
 wire \Tile_X4Y10_NN4BEG[4] ;
 wire \Tile_X4Y10_NN4BEG[5] ;
 wire \Tile_X4Y10_NN4BEG[6] ;
 wire \Tile_X4Y10_NN4BEG[7] ;
 wire \Tile_X4Y10_NN4BEG[8] ;
 wire \Tile_X4Y10_NN4BEG[9] ;
 wire \Tile_X4Y10_S1BEG[0] ;
 wire \Tile_X4Y10_S1BEG[1] ;
 wire \Tile_X4Y10_S1BEG[2] ;
 wire \Tile_X4Y10_S1BEG[3] ;
 wire \Tile_X4Y10_S2BEG[0] ;
 wire \Tile_X4Y10_S2BEG[1] ;
 wire \Tile_X4Y10_S2BEG[2] ;
 wire \Tile_X4Y10_S2BEG[3] ;
 wire \Tile_X4Y10_S2BEG[4] ;
 wire \Tile_X4Y10_S2BEG[5] ;
 wire \Tile_X4Y10_S2BEG[6] ;
 wire \Tile_X4Y10_S2BEG[7] ;
 wire \Tile_X4Y10_S2BEGb[0] ;
 wire \Tile_X4Y10_S2BEGb[1] ;
 wire \Tile_X4Y10_S2BEGb[2] ;
 wire \Tile_X4Y10_S2BEGb[3] ;
 wire \Tile_X4Y10_S2BEGb[4] ;
 wire \Tile_X4Y10_S2BEGb[5] ;
 wire \Tile_X4Y10_S2BEGb[6] ;
 wire \Tile_X4Y10_S2BEGb[7] ;
 wire \Tile_X4Y10_S4BEG[0] ;
 wire \Tile_X4Y10_S4BEG[10] ;
 wire \Tile_X4Y10_S4BEG[11] ;
 wire \Tile_X4Y10_S4BEG[12] ;
 wire \Tile_X4Y10_S4BEG[13] ;
 wire \Tile_X4Y10_S4BEG[14] ;
 wire \Tile_X4Y10_S4BEG[15] ;
 wire \Tile_X4Y10_S4BEG[1] ;
 wire \Tile_X4Y10_S4BEG[2] ;
 wire \Tile_X4Y10_S4BEG[3] ;
 wire \Tile_X4Y10_S4BEG[4] ;
 wire \Tile_X4Y10_S4BEG[5] ;
 wire \Tile_X4Y10_S4BEG[6] ;
 wire \Tile_X4Y10_S4BEG[7] ;
 wire \Tile_X4Y10_S4BEG[8] ;
 wire \Tile_X4Y10_S4BEG[9] ;
 wire \Tile_X4Y10_SS4BEG[0] ;
 wire \Tile_X4Y10_SS4BEG[10] ;
 wire \Tile_X4Y10_SS4BEG[11] ;
 wire \Tile_X4Y10_SS4BEG[12] ;
 wire \Tile_X4Y10_SS4BEG[13] ;
 wire \Tile_X4Y10_SS4BEG[14] ;
 wire \Tile_X4Y10_SS4BEG[15] ;
 wire \Tile_X4Y10_SS4BEG[1] ;
 wire \Tile_X4Y10_SS4BEG[2] ;
 wire \Tile_X4Y10_SS4BEG[3] ;
 wire \Tile_X4Y10_SS4BEG[4] ;
 wire \Tile_X4Y10_SS4BEG[5] ;
 wire \Tile_X4Y10_SS4BEG[6] ;
 wire \Tile_X4Y10_SS4BEG[7] ;
 wire \Tile_X4Y10_SS4BEG[8] ;
 wire \Tile_X4Y10_SS4BEG[9] ;
 wire Tile_X4Y10_UserCLKo;
 wire \Tile_X4Y10_W1BEG[0] ;
 wire \Tile_X4Y10_W1BEG[1] ;
 wire \Tile_X4Y10_W1BEG[2] ;
 wire \Tile_X4Y10_W1BEG[3] ;
 wire \Tile_X4Y10_W2BEG[0] ;
 wire \Tile_X4Y10_W2BEG[1] ;
 wire \Tile_X4Y10_W2BEG[2] ;
 wire \Tile_X4Y10_W2BEG[3] ;
 wire \Tile_X4Y10_W2BEG[4] ;
 wire \Tile_X4Y10_W2BEG[5] ;
 wire \Tile_X4Y10_W2BEG[6] ;
 wire \Tile_X4Y10_W2BEG[7] ;
 wire \Tile_X4Y10_W2BEGb[0] ;
 wire \Tile_X4Y10_W2BEGb[1] ;
 wire \Tile_X4Y10_W2BEGb[2] ;
 wire \Tile_X4Y10_W2BEGb[3] ;
 wire \Tile_X4Y10_W2BEGb[4] ;
 wire \Tile_X4Y10_W2BEGb[5] ;
 wire \Tile_X4Y10_W2BEGb[6] ;
 wire \Tile_X4Y10_W2BEGb[7] ;
 wire \Tile_X4Y10_W6BEG[0] ;
 wire \Tile_X4Y10_W6BEG[10] ;
 wire \Tile_X4Y10_W6BEG[11] ;
 wire \Tile_X4Y10_W6BEG[1] ;
 wire \Tile_X4Y10_W6BEG[2] ;
 wire \Tile_X4Y10_W6BEG[3] ;
 wire \Tile_X4Y10_W6BEG[4] ;
 wire \Tile_X4Y10_W6BEG[5] ;
 wire \Tile_X4Y10_W6BEG[6] ;
 wire \Tile_X4Y10_W6BEG[7] ;
 wire \Tile_X4Y10_W6BEG[8] ;
 wire \Tile_X4Y10_W6BEG[9] ;
 wire \Tile_X4Y10_WW4BEG[0] ;
 wire \Tile_X4Y10_WW4BEG[10] ;
 wire \Tile_X4Y10_WW4BEG[11] ;
 wire \Tile_X4Y10_WW4BEG[12] ;
 wire \Tile_X4Y10_WW4BEG[13] ;
 wire \Tile_X4Y10_WW4BEG[14] ;
 wire \Tile_X4Y10_WW4BEG[15] ;
 wire \Tile_X4Y10_WW4BEG[1] ;
 wire \Tile_X4Y10_WW4BEG[2] ;
 wire \Tile_X4Y10_WW4BEG[3] ;
 wire \Tile_X4Y10_WW4BEG[4] ;
 wire \Tile_X4Y10_WW4BEG[5] ;
 wire \Tile_X4Y10_WW4BEG[6] ;
 wire \Tile_X4Y10_WW4BEG[7] ;
 wire \Tile_X4Y10_WW4BEG[8] ;
 wire \Tile_X4Y10_WW4BEG[9] ;
 wire \Tile_X4Y11_E1BEG[0] ;
 wire \Tile_X4Y11_E1BEG[1] ;
 wire \Tile_X4Y11_E1BEG[2] ;
 wire \Tile_X4Y11_E1BEG[3] ;
 wire \Tile_X4Y11_E2BEG[0] ;
 wire \Tile_X4Y11_E2BEG[1] ;
 wire \Tile_X4Y11_E2BEG[2] ;
 wire \Tile_X4Y11_E2BEG[3] ;
 wire \Tile_X4Y11_E2BEG[4] ;
 wire \Tile_X4Y11_E2BEG[5] ;
 wire \Tile_X4Y11_E2BEG[6] ;
 wire \Tile_X4Y11_E2BEG[7] ;
 wire \Tile_X4Y11_E2BEGb[0] ;
 wire \Tile_X4Y11_E2BEGb[1] ;
 wire \Tile_X4Y11_E2BEGb[2] ;
 wire \Tile_X4Y11_E2BEGb[3] ;
 wire \Tile_X4Y11_E2BEGb[4] ;
 wire \Tile_X4Y11_E2BEGb[5] ;
 wire \Tile_X4Y11_E2BEGb[6] ;
 wire \Tile_X4Y11_E2BEGb[7] ;
 wire \Tile_X4Y11_E6BEG[0] ;
 wire \Tile_X4Y11_E6BEG[10] ;
 wire \Tile_X4Y11_E6BEG[11] ;
 wire \Tile_X4Y11_E6BEG[1] ;
 wire \Tile_X4Y11_E6BEG[2] ;
 wire \Tile_X4Y11_E6BEG[3] ;
 wire \Tile_X4Y11_E6BEG[4] ;
 wire \Tile_X4Y11_E6BEG[5] ;
 wire \Tile_X4Y11_E6BEG[6] ;
 wire \Tile_X4Y11_E6BEG[7] ;
 wire \Tile_X4Y11_E6BEG[8] ;
 wire \Tile_X4Y11_E6BEG[9] ;
 wire \Tile_X4Y11_EE4BEG[0] ;
 wire \Tile_X4Y11_EE4BEG[10] ;
 wire \Tile_X4Y11_EE4BEG[11] ;
 wire \Tile_X4Y11_EE4BEG[12] ;
 wire \Tile_X4Y11_EE4BEG[13] ;
 wire \Tile_X4Y11_EE4BEG[14] ;
 wire \Tile_X4Y11_EE4BEG[15] ;
 wire \Tile_X4Y11_EE4BEG[1] ;
 wire \Tile_X4Y11_EE4BEG[2] ;
 wire \Tile_X4Y11_EE4BEG[3] ;
 wire \Tile_X4Y11_EE4BEG[4] ;
 wire \Tile_X4Y11_EE4BEG[5] ;
 wire \Tile_X4Y11_EE4BEG[6] ;
 wire \Tile_X4Y11_EE4BEG[7] ;
 wire \Tile_X4Y11_EE4BEG[8] ;
 wire \Tile_X4Y11_EE4BEG[9] ;
 wire \Tile_X4Y11_FrameData_O[0] ;
 wire \Tile_X4Y11_FrameData_O[10] ;
 wire \Tile_X4Y11_FrameData_O[11] ;
 wire \Tile_X4Y11_FrameData_O[12] ;
 wire \Tile_X4Y11_FrameData_O[13] ;
 wire \Tile_X4Y11_FrameData_O[14] ;
 wire \Tile_X4Y11_FrameData_O[15] ;
 wire \Tile_X4Y11_FrameData_O[16] ;
 wire \Tile_X4Y11_FrameData_O[17] ;
 wire \Tile_X4Y11_FrameData_O[18] ;
 wire \Tile_X4Y11_FrameData_O[19] ;
 wire \Tile_X4Y11_FrameData_O[1] ;
 wire \Tile_X4Y11_FrameData_O[20] ;
 wire \Tile_X4Y11_FrameData_O[21] ;
 wire \Tile_X4Y11_FrameData_O[22] ;
 wire \Tile_X4Y11_FrameData_O[23] ;
 wire \Tile_X4Y11_FrameData_O[24] ;
 wire \Tile_X4Y11_FrameData_O[25] ;
 wire \Tile_X4Y11_FrameData_O[26] ;
 wire \Tile_X4Y11_FrameData_O[27] ;
 wire \Tile_X4Y11_FrameData_O[28] ;
 wire \Tile_X4Y11_FrameData_O[29] ;
 wire \Tile_X4Y11_FrameData_O[2] ;
 wire \Tile_X4Y11_FrameData_O[30] ;
 wire \Tile_X4Y11_FrameData_O[31] ;
 wire \Tile_X4Y11_FrameData_O[3] ;
 wire \Tile_X4Y11_FrameData_O[4] ;
 wire \Tile_X4Y11_FrameData_O[5] ;
 wire \Tile_X4Y11_FrameData_O[6] ;
 wire \Tile_X4Y11_FrameData_O[7] ;
 wire \Tile_X4Y11_FrameData_O[8] ;
 wire \Tile_X4Y11_FrameData_O[9] ;
 wire \Tile_X4Y11_FrameStrobe_O[0] ;
 wire \Tile_X4Y11_FrameStrobe_O[10] ;
 wire \Tile_X4Y11_FrameStrobe_O[11] ;
 wire \Tile_X4Y11_FrameStrobe_O[12] ;
 wire \Tile_X4Y11_FrameStrobe_O[13] ;
 wire \Tile_X4Y11_FrameStrobe_O[14] ;
 wire \Tile_X4Y11_FrameStrobe_O[15] ;
 wire \Tile_X4Y11_FrameStrobe_O[16] ;
 wire \Tile_X4Y11_FrameStrobe_O[17] ;
 wire \Tile_X4Y11_FrameStrobe_O[18] ;
 wire \Tile_X4Y11_FrameStrobe_O[19] ;
 wire \Tile_X4Y11_FrameStrobe_O[1] ;
 wire \Tile_X4Y11_FrameStrobe_O[2] ;
 wire \Tile_X4Y11_FrameStrobe_O[3] ;
 wire \Tile_X4Y11_FrameStrobe_O[4] ;
 wire \Tile_X4Y11_FrameStrobe_O[5] ;
 wire \Tile_X4Y11_FrameStrobe_O[6] ;
 wire \Tile_X4Y11_FrameStrobe_O[7] ;
 wire \Tile_X4Y11_FrameStrobe_O[8] ;
 wire \Tile_X4Y11_FrameStrobe_O[9] ;
 wire \Tile_X4Y11_N1BEG[0] ;
 wire \Tile_X4Y11_N1BEG[1] ;
 wire \Tile_X4Y11_N1BEG[2] ;
 wire \Tile_X4Y11_N1BEG[3] ;
 wire \Tile_X4Y11_N2BEG[0] ;
 wire \Tile_X4Y11_N2BEG[1] ;
 wire \Tile_X4Y11_N2BEG[2] ;
 wire \Tile_X4Y11_N2BEG[3] ;
 wire \Tile_X4Y11_N2BEG[4] ;
 wire \Tile_X4Y11_N2BEG[5] ;
 wire \Tile_X4Y11_N2BEG[6] ;
 wire \Tile_X4Y11_N2BEG[7] ;
 wire \Tile_X4Y11_N2BEGb[0] ;
 wire \Tile_X4Y11_N2BEGb[1] ;
 wire \Tile_X4Y11_N2BEGb[2] ;
 wire \Tile_X4Y11_N2BEGb[3] ;
 wire \Tile_X4Y11_N2BEGb[4] ;
 wire \Tile_X4Y11_N2BEGb[5] ;
 wire \Tile_X4Y11_N2BEGb[6] ;
 wire \Tile_X4Y11_N2BEGb[7] ;
 wire \Tile_X4Y11_N4BEG[0] ;
 wire \Tile_X4Y11_N4BEG[10] ;
 wire \Tile_X4Y11_N4BEG[11] ;
 wire \Tile_X4Y11_N4BEG[12] ;
 wire \Tile_X4Y11_N4BEG[13] ;
 wire \Tile_X4Y11_N4BEG[14] ;
 wire \Tile_X4Y11_N4BEG[15] ;
 wire \Tile_X4Y11_N4BEG[1] ;
 wire \Tile_X4Y11_N4BEG[2] ;
 wire \Tile_X4Y11_N4BEG[3] ;
 wire \Tile_X4Y11_N4BEG[4] ;
 wire \Tile_X4Y11_N4BEG[5] ;
 wire \Tile_X4Y11_N4BEG[6] ;
 wire \Tile_X4Y11_N4BEG[7] ;
 wire \Tile_X4Y11_N4BEG[8] ;
 wire \Tile_X4Y11_N4BEG[9] ;
 wire \Tile_X4Y11_NN4BEG[0] ;
 wire \Tile_X4Y11_NN4BEG[10] ;
 wire \Tile_X4Y11_NN4BEG[11] ;
 wire \Tile_X4Y11_NN4BEG[12] ;
 wire \Tile_X4Y11_NN4BEG[13] ;
 wire \Tile_X4Y11_NN4BEG[14] ;
 wire \Tile_X4Y11_NN4BEG[15] ;
 wire \Tile_X4Y11_NN4BEG[1] ;
 wire \Tile_X4Y11_NN4BEG[2] ;
 wire \Tile_X4Y11_NN4BEG[3] ;
 wire \Tile_X4Y11_NN4BEG[4] ;
 wire \Tile_X4Y11_NN4BEG[5] ;
 wire \Tile_X4Y11_NN4BEG[6] ;
 wire \Tile_X4Y11_NN4BEG[7] ;
 wire \Tile_X4Y11_NN4BEG[8] ;
 wire \Tile_X4Y11_NN4BEG[9] ;
 wire \Tile_X4Y11_S1BEG[0] ;
 wire \Tile_X4Y11_S1BEG[1] ;
 wire \Tile_X4Y11_S1BEG[2] ;
 wire \Tile_X4Y11_S1BEG[3] ;
 wire \Tile_X4Y11_S2BEG[0] ;
 wire \Tile_X4Y11_S2BEG[1] ;
 wire \Tile_X4Y11_S2BEG[2] ;
 wire \Tile_X4Y11_S2BEG[3] ;
 wire \Tile_X4Y11_S2BEG[4] ;
 wire \Tile_X4Y11_S2BEG[5] ;
 wire \Tile_X4Y11_S2BEG[6] ;
 wire \Tile_X4Y11_S2BEG[7] ;
 wire \Tile_X4Y11_S2BEGb[0] ;
 wire \Tile_X4Y11_S2BEGb[1] ;
 wire \Tile_X4Y11_S2BEGb[2] ;
 wire \Tile_X4Y11_S2BEGb[3] ;
 wire \Tile_X4Y11_S2BEGb[4] ;
 wire \Tile_X4Y11_S2BEGb[5] ;
 wire \Tile_X4Y11_S2BEGb[6] ;
 wire \Tile_X4Y11_S2BEGb[7] ;
 wire \Tile_X4Y11_S4BEG[0] ;
 wire \Tile_X4Y11_S4BEG[10] ;
 wire \Tile_X4Y11_S4BEG[11] ;
 wire \Tile_X4Y11_S4BEG[12] ;
 wire \Tile_X4Y11_S4BEG[13] ;
 wire \Tile_X4Y11_S4BEG[14] ;
 wire \Tile_X4Y11_S4BEG[15] ;
 wire \Tile_X4Y11_S4BEG[1] ;
 wire \Tile_X4Y11_S4BEG[2] ;
 wire \Tile_X4Y11_S4BEG[3] ;
 wire \Tile_X4Y11_S4BEG[4] ;
 wire \Tile_X4Y11_S4BEG[5] ;
 wire \Tile_X4Y11_S4BEG[6] ;
 wire \Tile_X4Y11_S4BEG[7] ;
 wire \Tile_X4Y11_S4BEG[8] ;
 wire \Tile_X4Y11_S4BEG[9] ;
 wire \Tile_X4Y11_SS4BEG[0] ;
 wire \Tile_X4Y11_SS4BEG[10] ;
 wire \Tile_X4Y11_SS4BEG[11] ;
 wire \Tile_X4Y11_SS4BEG[12] ;
 wire \Tile_X4Y11_SS4BEG[13] ;
 wire \Tile_X4Y11_SS4BEG[14] ;
 wire \Tile_X4Y11_SS4BEG[15] ;
 wire \Tile_X4Y11_SS4BEG[1] ;
 wire \Tile_X4Y11_SS4BEG[2] ;
 wire \Tile_X4Y11_SS4BEG[3] ;
 wire \Tile_X4Y11_SS4BEG[4] ;
 wire \Tile_X4Y11_SS4BEG[5] ;
 wire \Tile_X4Y11_SS4BEG[6] ;
 wire \Tile_X4Y11_SS4BEG[7] ;
 wire \Tile_X4Y11_SS4BEG[8] ;
 wire \Tile_X4Y11_SS4BEG[9] ;
 wire Tile_X4Y11_UserCLKo;
 wire \Tile_X4Y11_W1BEG[0] ;
 wire \Tile_X4Y11_W1BEG[1] ;
 wire \Tile_X4Y11_W1BEG[2] ;
 wire \Tile_X4Y11_W1BEG[3] ;
 wire \Tile_X4Y11_W2BEG[0] ;
 wire \Tile_X4Y11_W2BEG[1] ;
 wire \Tile_X4Y11_W2BEG[2] ;
 wire \Tile_X4Y11_W2BEG[3] ;
 wire \Tile_X4Y11_W2BEG[4] ;
 wire \Tile_X4Y11_W2BEG[5] ;
 wire \Tile_X4Y11_W2BEG[6] ;
 wire \Tile_X4Y11_W2BEG[7] ;
 wire \Tile_X4Y11_W2BEGb[0] ;
 wire \Tile_X4Y11_W2BEGb[1] ;
 wire \Tile_X4Y11_W2BEGb[2] ;
 wire \Tile_X4Y11_W2BEGb[3] ;
 wire \Tile_X4Y11_W2BEGb[4] ;
 wire \Tile_X4Y11_W2BEGb[5] ;
 wire \Tile_X4Y11_W2BEGb[6] ;
 wire \Tile_X4Y11_W2BEGb[7] ;
 wire \Tile_X4Y11_W6BEG[0] ;
 wire \Tile_X4Y11_W6BEG[10] ;
 wire \Tile_X4Y11_W6BEG[11] ;
 wire \Tile_X4Y11_W6BEG[1] ;
 wire \Tile_X4Y11_W6BEG[2] ;
 wire \Tile_X4Y11_W6BEG[3] ;
 wire \Tile_X4Y11_W6BEG[4] ;
 wire \Tile_X4Y11_W6BEG[5] ;
 wire \Tile_X4Y11_W6BEG[6] ;
 wire \Tile_X4Y11_W6BEG[7] ;
 wire \Tile_X4Y11_W6BEG[8] ;
 wire \Tile_X4Y11_W6BEG[9] ;
 wire \Tile_X4Y11_WW4BEG[0] ;
 wire \Tile_X4Y11_WW4BEG[10] ;
 wire \Tile_X4Y11_WW4BEG[11] ;
 wire \Tile_X4Y11_WW4BEG[12] ;
 wire \Tile_X4Y11_WW4BEG[13] ;
 wire \Tile_X4Y11_WW4BEG[14] ;
 wire \Tile_X4Y11_WW4BEG[15] ;
 wire \Tile_X4Y11_WW4BEG[1] ;
 wire \Tile_X4Y11_WW4BEG[2] ;
 wire \Tile_X4Y11_WW4BEG[3] ;
 wire \Tile_X4Y11_WW4BEG[4] ;
 wire \Tile_X4Y11_WW4BEG[5] ;
 wire \Tile_X4Y11_WW4BEG[6] ;
 wire \Tile_X4Y11_WW4BEG[7] ;
 wire \Tile_X4Y11_WW4BEG[8] ;
 wire \Tile_X4Y11_WW4BEG[9] ;
 wire \Tile_X4Y12_E1BEG[0] ;
 wire \Tile_X4Y12_E1BEG[1] ;
 wire \Tile_X4Y12_E1BEG[2] ;
 wire \Tile_X4Y12_E1BEG[3] ;
 wire \Tile_X4Y12_E2BEG[0] ;
 wire \Tile_X4Y12_E2BEG[1] ;
 wire \Tile_X4Y12_E2BEG[2] ;
 wire \Tile_X4Y12_E2BEG[3] ;
 wire \Tile_X4Y12_E2BEG[4] ;
 wire \Tile_X4Y12_E2BEG[5] ;
 wire \Tile_X4Y12_E2BEG[6] ;
 wire \Tile_X4Y12_E2BEG[7] ;
 wire \Tile_X4Y12_E2BEGb[0] ;
 wire \Tile_X4Y12_E2BEGb[1] ;
 wire \Tile_X4Y12_E2BEGb[2] ;
 wire \Tile_X4Y12_E2BEGb[3] ;
 wire \Tile_X4Y12_E2BEGb[4] ;
 wire \Tile_X4Y12_E2BEGb[5] ;
 wire \Tile_X4Y12_E2BEGb[6] ;
 wire \Tile_X4Y12_E2BEGb[7] ;
 wire \Tile_X4Y12_E6BEG[0] ;
 wire \Tile_X4Y12_E6BEG[10] ;
 wire \Tile_X4Y12_E6BEG[11] ;
 wire \Tile_X4Y12_E6BEG[1] ;
 wire \Tile_X4Y12_E6BEG[2] ;
 wire \Tile_X4Y12_E6BEG[3] ;
 wire \Tile_X4Y12_E6BEG[4] ;
 wire \Tile_X4Y12_E6BEG[5] ;
 wire \Tile_X4Y12_E6BEG[6] ;
 wire \Tile_X4Y12_E6BEG[7] ;
 wire \Tile_X4Y12_E6BEG[8] ;
 wire \Tile_X4Y12_E6BEG[9] ;
 wire \Tile_X4Y12_EE4BEG[0] ;
 wire \Tile_X4Y12_EE4BEG[10] ;
 wire \Tile_X4Y12_EE4BEG[11] ;
 wire \Tile_X4Y12_EE4BEG[12] ;
 wire \Tile_X4Y12_EE4BEG[13] ;
 wire \Tile_X4Y12_EE4BEG[14] ;
 wire \Tile_X4Y12_EE4BEG[15] ;
 wire \Tile_X4Y12_EE4BEG[1] ;
 wire \Tile_X4Y12_EE4BEG[2] ;
 wire \Tile_X4Y12_EE4BEG[3] ;
 wire \Tile_X4Y12_EE4BEG[4] ;
 wire \Tile_X4Y12_EE4BEG[5] ;
 wire \Tile_X4Y12_EE4BEG[6] ;
 wire \Tile_X4Y12_EE4BEG[7] ;
 wire \Tile_X4Y12_EE4BEG[8] ;
 wire \Tile_X4Y12_EE4BEG[9] ;
 wire \Tile_X4Y12_FrameData_O[0] ;
 wire \Tile_X4Y12_FrameData_O[10] ;
 wire \Tile_X4Y12_FrameData_O[11] ;
 wire \Tile_X4Y12_FrameData_O[12] ;
 wire \Tile_X4Y12_FrameData_O[13] ;
 wire \Tile_X4Y12_FrameData_O[14] ;
 wire \Tile_X4Y12_FrameData_O[15] ;
 wire \Tile_X4Y12_FrameData_O[16] ;
 wire \Tile_X4Y12_FrameData_O[17] ;
 wire \Tile_X4Y12_FrameData_O[18] ;
 wire \Tile_X4Y12_FrameData_O[19] ;
 wire \Tile_X4Y12_FrameData_O[1] ;
 wire \Tile_X4Y12_FrameData_O[20] ;
 wire \Tile_X4Y12_FrameData_O[21] ;
 wire \Tile_X4Y12_FrameData_O[22] ;
 wire \Tile_X4Y12_FrameData_O[23] ;
 wire \Tile_X4Y12_FrameData_O[24] ;
 wire \Tile_X4Y12_FrameData_O[25] ;
 wire \Tile_X4Y12_FrameData_O[26] ;
 wire \Tile_X4Y12_FrameData_O[27] ;
 wire \Tile_X4Y12_FrameData_O[28] ;
 wire \Tile_X4Y12_FrameData_O[29] ;
 wire \Tile_X4Y12_FrameData_O[2] ;
 wire \Tile_X4Y12_FrameData_O[30] ;
 wire \Tile_X4Y12_FrameData_O[31] ;
 wire \Tile_X4Y12_FrameData_O[3] ;
 wire \Tile_X4Y12_FrameData_O[4] ;
 wire \Tile_X4Y12_FrameData_O[5] ;
 wire \Tile_X4Y12_FrameData_O[6] ;
 wire \Tile_X4Y12_FrameData_O[7] ;
 wire \Tile_X4Y12_FrameData_O[8] ;
 wire \Tile_X4Y12_FrameData_O[9] ;
 wire \Tile_X4Y12_FrameStrobe_O[0] ;
 wire \Tile_X4Y12_FrameStrobe_O[10] ;
 wire \Tile_X4Y12_FrameStrobe_O[11] ;
 wire \Tile_X4Y12_FrameStrobe_O[12] ;
 wire \Tile_X4Y12_FrameStrobe_O[13] ;
 wire \Tile_X4Y12_FrameStrobe_O[14] ;
 wire \Tile_X4Y12_FrameStrobe_O[15] ;
 wire \Tile_X4Y12_FrameStrobe_O[16] ;
 wire \Tile_X4Y12_FrameStrobe_O[17] ;
 wire \Tile_X4Y12_FrameStrobe_O[18] ;
 wire \Tile_X4Y12_FrameStrobe_O[19] ;
 wire \Tile_X4Y12_FrameStrobe_O[1] ;
 wire \Tile_X4Y12_FrameStrobe_O[2] ;
 wire \Tile_X4Y12_FrameStrobe_O[3] ;
 wire \Tile_X4Y12_FrameStrobe_O[4] ;
 wire \Tile_X4Y12_FrameStrobe_O[5] ;
 wire \Tile_X4Y12_FrameStrobe_O[6] ;
 wire \Tile_X4Y12_FrameStrobe_O[7] ;
 wire \Tile_X4Y12_FrameStrobe_O[8] ;
 wire \Tile_X4Y12_FrameStrobe_O[9] ;
 wire \Tile_X4Y12_N1BEG[0] ;
 wire \Tile_X4Y12_N1BEG[1] ;
 wire \Tile_X4Y12_N1BEG[2] ;
 wire \Tile_X4Y12_N1BEG[3] ;
 wire \Tile_X4Y12_N2BEG[0] ;
 wire \Tile_X4Y12_N2BEG[1] ;
 wire \Tile_X4Y12_N2BEG[2] ;
 wire \Tile_X4Y12_N2BEG[3] ;
 wire \Tile_X4Y12_N2BEG[4] ;
 wire \Tile_X4Y12_N2BEG[5] ;
 wire \Tile_X4Y12_N2BEG[6] ;
 wire \Tile_X4Y12_N2BEG[7] ;
 wire \Tile_X4Y12_N2BEGb[0] ;
 wire \Tile_X4Y12_N2BEGb[1] ;
 wire \Tile_X4Y12_N2BEGb[2] ;
 wire \Tile_X4Y12_N2BEGb[3] ;
 wire \Tile_X4Y12_N2BEGb[4] ;
 wire \Tile_X4Y12_N2BEGb[5] ;
 wire \Tile_X4Y12_N2BEGb[6] ;
 wire \Tile_X4Y12_N2BEGb[7] ;
 wire \Tile_X4Y12_N4BEG[0] ;
 wire \Tile_X4Y12_N4BEG[10] ;
 wire \Tile_X4Y12_N4BEG[11] ;
 wire \Tile_X4Y12_N4BEG[12] ;
 wire \Tile_X4Y12_N4BEG[13] ;
 wire \Tile_X4Y12_N4BEG[14] ;
 wire \Tile_X4Y12_N4BEG[15] ;
 wire \Tile_X4Y12_N4BEG[1] ;
 wire \Tile_X4Y12_N4BEG[2] ;
 wire \Tile_X4Y12_N4BEG[3] ;
 wire \Tile_X4Y12_N4BEG[4] ;
 wire \Tile_X4Y12_N4BEG[5] ;
 wire \Tile_X4Y12_N4BEG[6] ;
 wire \Tile_X4Y12_N4BEG[7] ;
 wire \Tile_X4Y12_N4BEG[8] ;
 wire \Tile_X4Y12_N4BEG[9] ;
 wire \Tile_X4Y12_NN4BEG[0] ;
 wire \Tile_X4Y12_NN4BEG[10] ;
 wire \Tile_X4Y12_NN4BEG[11] ;
 wire \Tile_X4Y12_NN4BEG[12] ;
 wire \Tile_X4Y12_NN4BEG[13] ;
 wire \Tile_X4Y12_NN4BEG[14] ;
 wire \Tile_X4Y12_NN4BEG[15] ;
 wire \Tile_X4Y12_NN4BEG[1] ;
 wire \Tile_X4Y12_NN4BEG[2] ;
 wire \Tile_X4Y12_NN4BEG[3] ;
 wire \Tile_X4Y12_NN4BEG[4] ;
 wire \Tile_X4Y12_NN4BEG[5] ;
 wire \Tile_X4Y12_NN4BEG[6] ;
 wire \Tile_X4Y12_NN4BEG[7] ;
 wire \Tile_X4Y12_NN4BEG[8] ;
 wire \Tile_X4Y12_NN4BEG[9] ;
 wire \Tile_X4Y12_S1BEG[0] ;
 wire \Tile_X4Y12_S1BEG[1] ;
 wire \Tile_X4Y12_S1BEG[2] ;
 wire \Tile_X4Y12_S1BEG[3] ;
 wire \Tile_X4Y12_S2BEG[0] ;
 wire \Tile_X4Y12_S2BEG[1] ;
 wire \Tile_X4Y12_S2BEG[2] ;
 wire \Tile_X4Y12_S2BEG[3] ;
 wire \Tile_X4Y12_S2BEG[4] ;
 wire \Tile_X4Y12_S2BEG[5] ;
 wire \Tile_X4Y12_S2BEG[6] ;
 wire \Tile_X4Y12_S2BEG[7] ;
 wire \Tile_X4Y12_S2BEGb[0] ;
 wire \Tile_X4Y12_S2BEGb[1] ;
 wire \Tile_X4Y12_S2BEGb[2] ;
 wire \Tile_X4Y12_S2BEGb[3] ;
 wire \Tile_X4Y12_S2BEGb[4] ;
 wire \Tile_X4Y12_S2BEGb[5] ;
 wire \Tile_X4Y12_S2BEGb[6] ;
 wire \Tile_X4Y12_S2BEGb[7] ;
 wire \Tile_X4Y12_S4BEG[0] ;
 wire \Tile_X4Y12_S4BEG[10] ;
 wire \Tile_X4Y12_S4BEG[11] ;
 wire \Tile_X4Y12_S4BEG[12] ;
 wire \Tile_X4Y12_S4BEG[13] ;
 wire \Tile_X4Y12_S4BEG[14] ;
 wire \Tile_X4Y12_S4BEG[15] ;
 wire \Tile_X4Y12_S4BEG[1] ;
 wire \Tile_X4Y12_S4BEG[2] ;
 wire \Tile_X4Y12_S4BEG[3] ;
 wire \Tile_X4Y12_S4BEG[4] ;
 wire \Tile_X4Y12_S4BEG[5] ;
 wire \Tile_X4Y12_S4BEG[6] ;
 wire \Tile_X4Y12_S4BEG[7] ;
 wire \Tile_X4Y12_S4BEG[8] ;
 wire \Tile_X4Y12_S4BEG[9] ;
 wire \Tile_X4Y12_SS4BEG[0] ;
 wire \Tile_X4Y12_SS4BEG[10] ;
 wire \Tile_X4Y12_SS4BEG[11] ;
 wire \Tile_X4Y12_SS4BEG[12] ;
 wire \Tile_X4Y12_SS4BEG[13] ;
 wire \Tile_X4Y12_SS4BEG[14] ;
 wire \Tile_X4Y12_SS4BEG[15] ;
 wire \Tile_X4Y12_SS4BEG[1] ;
 wire \Tile_X4Y12_SS4BEG[2] ;
 wire \Tile_X4Y12_SS4BEG[3] ;
 wire \Tile_X4Y12_SS4BEG[4] ;
 wire \Tile_X4Y12_SS4BEG[5] ;
 wire \Tile_X4Y12_SS4BEG[6] ;
 wire \Tile_X4Y12_SS4BEG[7] ;
 wire \Tile_X4Y12_SS4BEG[8] ;
 wire \Tile_X4Y12_SS4BEG[9] ;
 wire Tile_X4Y12_UserCLKo;
 wire \Tile_X4Y12_W1BEG[0] ;
 wire \Tile_X4Y12_W1BEG[1] ;
 wire \Tile_X4Y12_W1BEG[2] ;
 wire \Tile_X4Y12_W1BEG[3] ;
 wire \Tile_X4Y12_W2BEG[0] ;
 wire \Tile_X4Y12_W2BEG[1] ;
 wire \Tile_X4Y12_W2BEG[2] ;
 wire \Tile_X4Y12_W2BEG[3] ;
 wire \Tile_X4Y12_W2BEG[4] ;
 wire \Tile_X4Y12_W2BEG[5] ;
 wire \Tile_X4Y12_W2BEG[6] ;
 wire \Tile_X4Y12_W2BEG[7] ;
 wire \Tile_X4Y12_W2BEGb[0] ;
 wire \Tile_X4Y12_W2BEGb[1] ;
 wire \Tile_X4Y12_W2BEGb[2] ;
 wire \Tile_X4Y12_W2BEGb[3] ;
 wire \Tile_X4Y12_W2BEGb[4] ;
 wire \Tile_X4Y12_W2BEGb[5] ;
 wire \Tile_X4Y12_W2BEGb[6] ;
 wire \Tile_X4Y12_W2BEGb[7] ;
 wire \Tile_X4Y12_W6BEG[0] ;
 wire \Tile_X4Y12_W6BEG[10] ;
 wire \Tile_X4Y12_W6BEG[11] ;
 wire \Tile_X4Y12_W6BEG[1] ;
 wire \Tile_X4Y12_W6BEG[2] ;
 wire \Tile_X4Y12_W6BEG[3] ;
 wire \Tile_X4Y12_W6BEG[4] ;
 wire \Tile_X4Y12_W6BEG[5] ;
 wire \Tile_X4Y12_W6BEG[6] ;
 wire \Tile_X4Y12_W6BEG[7] ;
 wire \Tile_X4Y12_W6BEG[8] ;
 wire \Tile_X4Y12_W6BEG[9] ;
 wire \Tile_X4Y12_WW4BEG[0] ;
 wire \Tile_X4Y12_WW4BEG[10] ;
 wire \Tile_X4Y12_WW4BEG[11] ;
 wire \Tile_X4Y12_WW4BEG[12] ;
 wire \Tile_X4Y12_WW4BEG[13] ;
 wire \Tile_X4Y12_WW4BEG[14] ;
 wire \Tile_X4Y12_WW4BEG[15] ;
 wire \Tile_X4Y12_WW4BEG[1] ;
 wire \Tile_X4Y12_WW4BEG[2] ;
 wire \Tile_X4Y12_WW4BEG[3] ;
 wire \Tile_X4Y12_WW4BEG[4] ;
 wire \Tile_X4Y12_WW4BEG[5] ;
 wire \Tile_X4Y12_WW4BEG[6] ;
 wire \Tile_X4Y12_WW4BEG[7] ;
 wire \Tile_X4Y12_WW4BEG[8] ;
 wire \Tile_X4Y12_WW4BEG[9] ;
 wire \Tile_X4Y13_E1BEG[0] ;
 wire \Tile_X4Y13_E1BEG[1] ;
 wire \Tile_X4Y13_E1BEG[2] ;
 wire \Tile_X4Y13_E1BEG[3] ;
 wire \Tile_X4Y13_E2BEG[0] ;
 wire \Tile_X4Y13_E2BEG[1] ;
 wire \Tile_X4Y13_E2BEG[2] ;
 wire \Tile_X4Y13_E2BEG[3] ;
 wire \Tile_X4Y13_E2BEG[4] ;
 wire \Tile_X4Y13_E2BEG[5] ;
 wire \Tile_X4Y13_E2BEG[6] ;
 wire \Tile_X4Y13_E2BEG[7] ;
 wire \Tile_X4Y13_E2BEGb[0] ;
 wire \Tile_X4Y13_E2BEGb[1] ;
 wire \Tile_X4Y13_E2BEGb[2] ;
 wire \Tile_X4Y13_E2BEGb[3] ;
 wire \Tile_X4Y13_E2BEGb[4] ;
 wire \Tile_X4Y13_E2BEGb[5] ;
 wire \Tile_X4Y13_E2BEGb[6] ;
 wire \Tile_X4Y13_E2BEGb[7] ;
 wire \Tile_X4Y13_E6BEG[0] ;
 wire \Tile_X4Y13_E6BEG[10] ;
 wire \Tile_X4Y13_E6BEG[11] ;
 wire \Tile_X4Y13_E6BEG[1] ;
 wire \Tile_X4Y13_E6BEG[2] ;
 wire \Tile_X4Y13_E6BEG[3] ;
 wire \Tile_X4Y13_E6BEG[4] ;
 wire \Tile_X4Y13_E6BEG[5] ;
 wire \Tile_X4Y13_E6BEG[6] ;
 wire \Tile_X4Y13_E6BEG[7] ;
 wire \Tile_X4Y13_E6BEG[8] ;
 wire \Tile_X4Y13_E6BEG[9] ;
 wire \Tile_X4Y13_EE4BEG[0] ;
 wire \Tile_X4Y13_EE4BEG[10] ;
 wire \Tile_X4Y13_EE4BEG[11] ;
 wire \Tile_X4Y13_EE4BEG[12] ;
 wire \Tile_X4Y13_EE4BEG[13] ;
 wire \Tile_X4Y13_EE4BEG[14] ;
 wire \Tile_X4Y13_EE4BEG[15] ;
 wire \Tile_X4Y13_EE4BEG[1] ;
 wire \Tile_X4Y13_EE4BEG[2] ;
 wire \Tile_X4Y13_EE4BEG[3] ;
 wire \Tile_X4Y13_EE4BEG[4] ;
 wire \Tile_X4Y13_EE4BEG[5] ;
 wire \Tile_X4Y13_EE4BEG[6] ;
 wire \Tile_X4Y13_EE4BEG[7] ;
 wire \Tile_X4Y13_EE4BEG[8] ;
 wire \Tile_X4Y13_EE4BEG[9] ;
 wire \Tile_X4Y13_FrameData_O[0] ;
 wire \Tile_X4Y13_FrameData_O[10] ;
 wire \Tile_X4Y13_FrameData_O[11] ;
 wire \Tile_X4Y13_FrameData_O[12] ;
 wire \Tile_X4Y13_FrameData_O[13] ;
 wire \Tile_X4Y13_FrameData_O[14] ;
 wire \Tile_X4Y13_FrameData_O[15] ;
 wire \Tile_X4Y13_FrameData_O[16] ;
 wire \Tile_X4Y13_FrameData_O[17] ;
 wire \Tile_X4Y13_FrameData_O[18] ;
 wire \Tile_X4Y13_FrameData_O[19] ;
 wire \Tile_X4Y13_FrameData_O[1] ;
 wire \Tile_X4Y13_FrameData_O[20] ;
 wire \Tile_X4Y13_FrameData_O[21] ;
 wire \Tile_X4Y13_FrameData_O[22] ;
 wire \Tile_X4Y13_FrameData_O[23] ;
 wire \Tile_X4Y13_FrameData_O[24] ;
 wire \Tile_X4Y13_FrameData_O[25] ;
 wire \Tile_X4Y13_FrameData_O[26] ;
 wire \Tile_X4Y13_FrameData_O[27] ;
 wire \Tile_X4Y13_FrameData_O[28] ;
 wire \Tile_X4Y13_FrameData_O[29] ;
 wire \Tile_X4Y13_FrameData_O[2] ;
 wire \Tile_X4Y13_FrameData_O[30] ;
 wire \Tile_X4Y13_FrameData_O[31] ;
 wire \Tile_X4Y13_FrameData_O[3] ;
 wire \Tile_X4Y13_FrameData_O[4] ;
 wire \Tile_X4Y13_FrameData_O[5] ;
 wire \Tile_X4Y13_FrameData_O[6] ;
 wire \Tile_X4Y13_FrameData_O[7] ;
 wire \Tile_X4Y13_FrameData_O[8] ;
 wire \Tile_X4Y13_FrameData_O[9] ;
 wire \Tile_X4Y13_FrameStrobe_O[0] ;
 wire \Tile_X4Y13_FrameStrobe_O[10] ;
 wire \Tile_X4Y13_FrameStrobe_O[11] ;
 wire \Tile_X4Y13_FrameStrobe_O[12] ;
 wire \Tile_X4Y13_FrameStrobe_O[13] ;
 wire \Tile_X4Y13_FrameStrobe_O[14] ;
 wire \Tile_X4Y13_FrameStrobe_O[15] ;
 wire \Tile_X4Y13_FrameStrobe_O[16] ;
 wire \Tile_X4Y13_FrameStrobe_O[17] ;
 wire \Tile_X4Y13_FrameStrobe_O[18] ;
 wire \Tile_X4Y13_FrameStrobe_O[19] ;
 wire \Tile_X4Y13_FrameStrobe_O[1] ;
 wire \Tile_X4Y13_FrameStrobe_O[2] ;
 wire \Tile_X4Y13_FrameStrobe_O[3] ;
 wire \Tile_X4Y13_FrameStrobe_O[4] ;
 wire \Tile_X4Y13_FrameStrobe_O[5] ;
 wire \Tile_X4Y13_FrameStrobe_O[6] ;
 wire \Tile_X4Y13_FrameStrobe_O[7] ;
 wire \Tile_X4Y13_FrameStrobe_O[8] ;
 wire \Tile_X4Y13_FrameStrobe_O[9] ;
 wire \Tile_X4Y13_N1BEG[0] ;
 wire \Tile_X4Y13_N1BEG[1] ;
 wire \Tile_X4Y13_N1BEG[2] ;
 wire \Tile_X4Y13_N1BEG[3] ;
 wire \Tile_X4Y13_N2BEG[0] ;
 wire \Tile_X4Y13_N2BEG[1] ;
 wire \Tile_X4Y13_N2BEG[2] ;
 wire \Tile_X4Y13_N2BEG[3] ;
 wire \Tile_X4Y13_N2BEG[4] ;
 wire \Tile_X4Y13_N2BEG[5] ;
 wire \Tile_X4Y13_N2BEG[6] ;
 wire \Tile_X4Y13_N2BEG[7] ;
 wire \Tile_X4Y13_N2BEGb[0] ;
 wire \Tile_X4Y13_N2BEGb[1] ;
 wire \Tile_X4Y13_N2BEGb[2] ;
 wire \Tile_X4Y13_N2BEGb[3] ;
 wire \Tile_X4Y13_N2BEGb[4] ;
 wire \Tile_X4Y13_N2BEGb[5] ;
 wire \Tile_X4Y13_N2BEGb[6] ;
 wire \Tile_X4Y13_N2BEGb[7] ;
 wire \Tile_X4Y13_N4BEG[0] ;
 wire \Tile_X4Y13_N4BEG[10] ;
 wire \Tile_X4Y13_N4BEG[11] ;
 wire \Tile_X4Y13_N4BEG[12] ;
 wire \Tile_X4Y13_N4BEG[13] ;
 wire \Tile_X4Y13_N4BEG[14] ;
 wire \Tile_X4Y13_N4BEG[15] ;
 wire \Tile_X4Y13_N4BEG[1] ;
 wire \Tile_X4Y13_N4BEG[2] ;
 wire \Tile_X4Y13_N4BEG[3] ;
 wire \Tile_X4Y13_N4BEG[4] ;
 wire \Tile_X4Y13_N4BEG[5] ;
 wire \Tile_X4Y13_N4BEG[6] ;
 wire \Tile_X4Y13_N4BEG[7] ;
 wire \Tile_X4Y13_N4BEG[8] ;
 wire \Tile_X4Y13_N4BEG[9] ;
 wire \Tile_X4Y13_NN4BEG[0] ;
 wire \Tile_X4Y13_NN4BEG[10] ;
 wire \Tile_X4Y13_NN4BEG[11] ;
 wire \Tile_X4Y13_NN4BEG[12] ;
 wire \Tile_X4Y13_NN4BEG[13] ;
 wire \Tile_X4Y13_NN4BEG[14] ;
 wire \Tile_X4Y13_NN4BEG[15] ;
 wire \Tile_X4Y13_NN4BEG[1] ;
 wire \Tile_X4Y13_NN4BEG[2] ;
 wire \Tile_X4Y13_NN4BEG[3] ;
 wire \Tile_X4Y13_NN4BEG[4] ;
 wire \Tile_X4Y13_NN4BEG[5] ;
 wire \Tile_X4Y13_NN4BEG[6] ;
 wire \Tile_X4Y13_NN4BEG[7] ;
 wire \Tile_X4Y13_NN4BEG[8] ;
 wire \Tile_X4Y13_NN4BEG[9] ;
 wire \Tile_X4Y13_S1BEG[0] ;
 wire \Tile_X4Y13_S1BEG[1] ;
 wire \Tile_X4Y13_S1BEG[2] ;
 wire \Tile_X4Y13_S1BEG[3] ;
 wire \Tile_X4Y13_S2BEG[0] ;
 wire \Tile_X4Y13_S2BEG[1] ;
 wire \Tile_X4Y13_S2BEG[2] ;
 wire \Tile_X4Y13_S2BEG[3] ;
 wire \Tile_X4Y13_S2BEG[4] ;
 wire \Tile_X4Y13_S2BEG[5] ;
 wire \Tile_X4Y13_S2BEG[6] ;
 wire \Tile_X4Y13_S2BEG[7] ;
 wire \Tile_X4Y13_S2BEGb[0] ;
 wire \Tile_X4Y13_S2BEGb[1] ;
 wire \Tile_X4Y13_S2BEGb[2] ;
 wire \Tile_X4Y13_S2BEGb[3] ;
 wire \Tile_X4Y13_S2BEGb[4] ;
 wire \Tile_X4Y13_S2BEGb[5] ;
 wire \Tile_X4Y13_S2BEGb[6] ;
 wire \Tile_X4Y13_S2BEGb[7] ;
 wire \Tile_X4Y13_S4BEG[0] ;
 wire \Tile_X4Y13_S4BEG[10] ;
 wire \Tile_X4Y13_S4BEG[11] ;
 wire \Tile_X4Y13_S4BEG[12] ;
 wire \Tile_X4Y13_S4BEG[13] ;
 wire \Tile_X4Y13_S4BEG[14] ;
 wire \Tile_X4Y13_S4BEG[15] ;
 wire \Tile_X4Y13_S4BEG[1] ;
 wire \Tile_X4Y13_S4BEG[2] ;
 wire \Tile_X4Y13_S4BEG[3] ;
 wire \Tile_X4Y13_S4BEG[4] ;
 wire \Tile_X4Y13_S4BEG[5] ;
 wire \Tile_X4Y13_S4BEG[6] ;
 wire \Tile_X4Y13_S4BEG[7] ;
 wire \Tile_X4Y13_S4BEG[8] ;
 wire \Tile_X4Y13_S4BEG[9] ;
 wire \Tile_X4Y13_SS4BEG[0] ;
 wire \Tile_X4Y13_SS4BEG[10] ;
 wire \Tile_X4Y13_SS4BEG[11] ;
 wire \Tile_X4Y13_SS4BEG[12] ;
 wire \Tile_X4Y13_SS4BEG[13] ;
 wire \Tile_X4Y13_SS4BEG[14] ;
 wire \Tile_X4Y13_SS4BEG[15] ;
 wire \Tile_X4Y13_SS4BEG[1] ;
 wire \Tile_X4Y13_SS4BEG[2] ;
 wire \Tile_X4Y13_SS4BEG[3] ;
 wire \Tile_X4Y13_SS4BEG[4] ;
 wire \Tile_X4Y13_SS4BEG[5] ;
 wire \Tile_X4Y13_SS4BEG[6] ;
 wire \Tile_X4Y13_SS4BEG[7] ;
 wire \Tile_X4Y13_SS4BEG[8] ;
 wire \Tile_X4Y13_SS4BEG[9] ;
 wire Tile_X4Y13_UserCLKo;
 wire \Tile_X4Y13_W1BEG[0] ;
 wire \Tile_X4Y13_W1BEG[1] ;
 wire \Tile_X4Y13_W1BEG[2] ;
 wire \Tile_X4Y13_W1BEG[3] ;
 wire \Tile_X4Y13_W2BEG[0] ;
 wire \Tile_X4Y13_W2BEG[1] ;
 wire \Tile_X4Y13_W2BEG[2] ;
 wire \Tile_X4Y13_W2BEG[3] ;
 wire \Tile_X4Y13_W2BEG[4] ;
 wire \Tile_X4Y13_W2BEG[5] ;
 wire \Tile_X4Y13_W2BEG[6] ;
 wire \Tile_X4Y13_W2BEG[7] ;
 wire \Tile_X4Y13_W2BEGb[0] ;
 wire \Tile_X4Y13_W2BEGb[1] ;
 wire \Tile_X4Y13_W2BEGb[2] ;
 wire \Tile_X4Y13_W2BEGb[3] ;
 wire \Tile_X4Y13_W2BEGb[4] ;
 wire \Tile_X4Y13_W2BEGb[5] ;
 wire \Tile_X4Y13_W2BEGb[6] ;
 wire \Tile_X4Y13_W2BEGb[7] ;
 wire \Tile_X4Y13_W6BEG[0] ;
 wire \Tile_X4Y13_W6BEG[10] ;
 wire \Tile_X4Y13_W6BEG[11] ;
 wire \Tile_X4Y13_W6BEG[1] ;
 wire \Tile_X4Y13_W6BEG[2] ;
 wire \Tile_X4Y13_W6BEG[3] ;
 wire \Tile_X4Y13_W6BEG[4] ;
 wire \Tile_X4Y13_W6BEG[5] ;
 wire \Tile_X4Y13_W6BEG[6] ;
 wire \Tile_X4Y13_W6BEG[7] ;
 wire \Tile_X4Y13_W6BEG[8] ;
 wire \Tile_X4Y13_W6BEG[9] ;
 wire \Tile_X4Y13_WW4BEG[0] ;
 wire \Tile_X4Y13_WW4BEG[10] ;
 wire \Tile_X4Y13_WW4BEG[11] ;
 wire \Tile_X4Y13_WW4BEG[12] ;
 wire \Tile_X4Y13_WW4BEG[13] ;
 wire \Tile_X4Y13_WW4BEG[14] ;
 wire \Tile_X4Y13_WW4BEG[15] ;
 wire \Tile_X4Y13_WW4BEG[1] ;
 wire \Tile_X4Y13_WW4BEG[2] ;
 wire \Tile_X4Y13_WW4BEG[3] ;
 wire \Tile_X4Y13_WW4BEG[4] ;
 wire \Tile_X4Y13_WW4BEG[5] ;
 wire \Tile_X4Y13_WW4BEG[6] ;
 wire \Tile_X4Y13_WW4BEG[7] ;
 wire \Tile_X4Y13_WW4BEG[8] ;
 wire \Tile_X4Y13_WW4BEG[9] ;
 wire \Tile_X4Y14_E1BEG[0] ;
 wire \Tile_X4Y14_E1BEG[1] ;
 wire \Tile_X4Y14_E1BEG[2] ;
 wire \Tile_X4Y14_E1BEG[3] ;
 wire \Tile_X4Y14_E2BEG[0] ;
 wire \Tile_X4Y14_E2BEG[1] ;
 wire \Tile_X4Y14_E2BEG[2] ;
 wire \Tile_X4Y14_E2BEG[3] ;
 wire \Tile_X4Y14_E2BEG[4] ;
 wire \Tile_X4Y14_E2BEG[5] ;
 wire \Tile_X4Y14_E2BEG[6] ;
 wire \Tile_X4Y14_E2BEG[7] ;
 wire \Tile_X4Y14_E2BEGb[0] ;
 wire \Tile_X4Y14_E2BEGb[1] ;
 wire \Tile_X4Y14_E2BEGb[2] ;
 wire \Tile_X4Y14_E2BEGb[3] ;
 wire \Tile_X4Y14_E2BEGb[4] ;
 wire \Tile_X4Y14_E2BEGb[5] ;
 wire \Tile_X4Y14_E2BEGb[6] ;
 wire \Tile_X4Y14_E2BEGb[7] ;
 wire \Tile_X4Y14_E6BEG[0] ;
 wire \Tile_X4Y14_E6BEG[10] ;
 wire \Tile_X4Y14_E6BEG[11] ;
 wire \Tile_X4Y14_E6BEG[1] ;
 wire \Tile_X4Y14_E6BEG[2] ;
 wire \Tile_X4Y14_E6BEG[3] ;
 wire \Tile_X4Y14_E6BEG[4] ;
 wire \Tile_X4Y14_E6BEG[5] ;
 wire \Tile_X4Y14_E6BEG[6] ;
 wire \Tile_X4Y14_E6BEG[7] ;
 wire \Tile_X4Y14_E6BEG[8] ;
 wire \Tile_X4Y14_E6BEG[9] ;
 wire \Tile_X4Y14_EE4BEG[0] ;
 wire \Tile_X4Y14_EE4BEG[10] ;
 wire \Tile_X4Y14_EE4BEG[11] ;
 wire \Tile_X4Y14_EE4BEG[12] ;
 wire \Tile_X4Y14_EE4BEG[13] ;
 wire \Tile_X4Y14_EE4BEG[14] ;
 wire \Tile_X4Y14_EE4BEG[15] ;
 wire \Tile_X4Y14_EE4BEG[1] ;
 wire \Tile_X4Y14_EE4BEG[2] ;
 wire \Tile_X4Y14_EE4BEG[3] ;
 wire \Tile_X4Y14_EE4BEG[4] ;
 wire \Tile_X4Y14_EE4BEG[5] ;
 wire \Tile_X4Y14_EE4BEG[6] ;
 wire \Tile_X4Y14_EE4BEG[7] ;
 wire \Tile_X4Y14_EE4BEG[8] ;
 wire \Tile_X4Y14_EE4BEG[9] ;
 wire \Tile_X4Y14_FrameData_O[0] ;
 wire \Tile_X4Y14_FrameData_O[10] ;
 wire \Tile_X4Y14_FrameData_O[11] ;
 wire \Tile_X4Y14_FrameData_O[12] ;
 wire \Tile_X4Y14_FrameData_O[13] ;
 wire \Tile_X4Y14_FrameData_O[14] ;
 wire \Tile_X4Y14_FrameData_O[15] ;
 wire \Tile_X4Y14_FrameData_O[16] ;
 wire \Tile_X4Y14_FrameData_O[17] ;
 wire \Tile_X4Y14_FrameData_O[18] ;
 wire \Tile_X4Y14_FrameData_O[19] ;
 wire \Tile_X4Y14_FrameData_O[1] ;
 wire \Tile_X4Y14_FrameData_O[20] ;
 wire \Tile_X4Y14_FrameData_O[21] ;
 wire \Tile_X4Y14_FrameData_O[22] ;
 wire \Tile_X4Y14_FrameData_O[23] ;
 wire \Tile_X4Y14_FrameData_O[24] ;
 wire \Tile_X4Y14_FrameData_O[25] ;
 wire \Tile_X4Y14_FrameData_O[26] ;
 wire \Tile_X4Y14_FrameData_O[27] ;
 wire \Tile_X4Y14_FrameData_O[28] ;
 wire \Tile_X4Y14_FrameData_O[29] ;
 wire \Tile_X4Y14_FrameData_O[2] ;
 wire \Tile_X4Y14_FrameData_O[30] ;
 wire \Tile_X4Y14_FrameData_O[31] ;
 wire \Tile_X4Y14_FrameData_O[3] ;
 wire \Tile_X4Y14_FrameData_O[4] ;
 wire \Tile_X4Y14_FrameData_O[5] ;
 wire \Tile_X4Y14_FrameData_O[6] ;
 wire \Tile_X4Y14_FrameData_O[7] ;
 wire \Tile_X4Y14_FrameData_O[8] ;
 wire \Tile_X4Y14_FrameData_O[9] ;
 wire \Tile_X4Y14_FrameStrobe_O[0] ;
 wire \Tile_X4Y14_FrameStrobe_O[10] ;
 wire \Tile_X4Y14_FrameStrobe_O[11] ;
 wire \Tile_X4Y14_FrameStrobe_O[12] ;
 wire \Tile_X4Y14_FrameStrobe_O[13] ;
 wire \Tile_X4Y14_FrameStrobe_O[14] ;
 wire \Tile_X4Y14_FrameStrobe_O[15] ;
 wire \Tile_X4Y14_FrameStrobe_O[16] ;
 wire \Tile_X4Y14_FrameStrobe_O[17] ;
 wire \Tile_X4Y14_FrameStrobe_O[18] ;
 wire \Tile_X4Y14_FrameStrobe_O[19] ;
 wire \Tile_X4Y14_FrameStrobe_O[1] ;
 wire \Tile_X4Y14_FrameStrobe_O[2] ;
 wire \Tile_X4Y14_FrameStrobe_O[3] ;
 wire \Tile_X4Y14_FrameStrobe_O[4] ;
 wire \Tile_X4Y14_FrameStrobe_O[5] ;
 wire \Tile_X4Y14_FrameStrobe_O[6] ;
 wire \Tile_X4Y14_FrameStrobe_O[7] ;
 wire \Tile_X4Y14_FrameStrobe_O[8] ;
 wire \Tile_X4Y14_FrameStrobe_O[9] ;
 wire \Tile_X4Y14_N1BEG[0] ;
 wire \Tile_X4Y14_N1BEG[1] ;
 wire \Tile_X4Y14_N1BEG[2] ;
 wire \Tile_X4Y14_N1BEG[3] ;
 wire \Tile_X4Y14_N2BEG[0] ;
 wire \Tile_X4Y14_N2BEG[1] ;
 wire \Tile_X4Y14_N2BEG[2] ;
 wire \Tile_X4Y14_N2BEG[3] ;
 wire \Tile_X4Y14_N2BEG[4] ;
 wire \Tile_X4Y14_N2BEG[5] ;
 wire \Tile_X4Y14_N2BEG[6] ;
 wire \Tile_X4Y14_N2BEG[7] ;
 wire \Tile_X4Y14_N2BEGb[0] ;
 wire \Tile_X4Y14_N2BEGb[1] ;
 wire \Tile_X4Y14_N2BEGb[2] ;
 wire \Tile_X4Y14_N2BEGb[3] ;
 wire \Tile_X4Y14_N2BEGb[4] ;
 wire \Tile_X4Y14_N2BEGb[5] ;
 wire \Tile_X4Y14_N2BEGb[6] ;
 wire \Tile_X4Y14_N2BEGb[7] ;
 wire \Tile_X4Y14_N4BEG[0] ;
 wire \Tile_X4Y14_N4BEG[10] ;
 wire \Tile_X4Y14_N4BEG[11] ;
 wire \Tile_X4Y14_N4BEG[12] ;
 wire \Tile_X4Y14_N4BEG[13] ;
 wire \Tile_X4Y14_N4BEG[14] ;
 wire \Tile_X4Y14_N4BEG[15] ;
 wire \Tile_X4Y14_N4BEG[1] ;
 wire \Tile_X4Y14_N4BEG[2] ;
 wire \Tile_X4Y14_N4BEG[3] ;
 wire \Tile_X4Y14_N4BEG[4] ;
 wire \Tile_X4Y14_N4BEG[5] ;
 wire \Tile_X4Y14_N4BEG[6] ;
 wire \Tile_X4Y14_N4BEG[7] ;
 wire \Tile_X4Y14_N4BEG[8] ;
 wire \Tile_X4Y14_N4BEG[9] ;
 wire \Tile_X4Y14_NN4BEG[0] ;
 wire \Tile_X4Y14_NN4BEG[10] ;
 wire \Tile_X4Y14_NN4BEG[11] ;
 wire \Tile_X4Y14_NN4BEG[12] ;
 wire \Tile_X4Y14_NN4BEG[13] ;
 wire \Tile_X4Y14_NN4BEG[14] ;
 wire \Tile_X4Y14_NN4BEG[15] ;
 wire \Tile_X4Y14_NN4BEG[1] ;
 wire \Tile_X4Y14_NN4BEG[2] ;
 wire \Tile_X4Y14_NN4BEG[3] ;
 wire \Tile_X4Y14_NN4BEG[4] ;
 wire \Tile_X4Y14_NN4BEG[5] ;
 wire \Tile_X4Y14_NN4BEG[6] ;
 wire \Tile_X4Y14_NN4BEG[7] ;
 wire \Tile_X4Y14_NN4BEG[8] ;
 wire \Tile_X4Y14_NN4BEG[9] ;
 wire \Tile_X4Y14_S1BEG[0] ;
 wire \Tile_X4Y14_S1BEG[1] ;
 wire \Tile_X4Y14_S1BEG[2] ;
 wire \Tile_X4Y14_S1BEG[3] ;
 wire \Tile_X4Y14_S2BEG[0] ;
 wire \Tile_X4Y14_S2BEG[1] ;
 wire \Tile_X4Y14_S2BEG[2] ;
 wire \Tile_X4Y14_S2BEG[3] ;
 wire \Tile_X4Y14_S2BEG[4] ;
 wire \Tile_X4Y14_S2BEG[5] ;
 wire \Tile_X4Y14_S2BEG[6] ;
 wire \Tile_X4Y14_S2BEG[7] ;
 wire \Tile_X4Y14_S2BEGb[0] ;
 wire \Tile_X4Y14_S2BEGb[1] ;
 wire \Tile_X4Y14_S2BEGb[2] ;
 wire \Tile_X4Y14_S2BEGb[3] ;
 wire \Tile_X4Y14_S2BEGb[4] ;
 wire \Tile_X4Y14_S2BEGb[5] ;
 wire \Tile_X4Y14_S2BEGb[6] ;
 wire \Tile_X4Y14_S2BEGb[7] ;
 wire \Tile_X4Y14_S4BEG[0] ;
 wire \Tile_X4Y14_S4BEG[10] ;
 wire \Tile_X4Y14_S4BEG[11] ;
 wire \Tile_X4Y14_S4BEG[12] ;
 wire \Tile_X4Y14_S4BEG[13] ;
 wire \Tile_X4Y14_S4BEG[14] ;
 wire \Tile_X4Y14_S4BEG[15] ;
 wire \Tile_X4Y14_S4BEG[1] ;
 wire \Tile_X4Y14_S4BEG[2] ;
 wire \Tile_X4Y14_S4BEG[3] ;
 wire \Tile_X4Y14_S4BEG[4] ;
 wire \Tile_X4Y14_S4BEG[5] ;
 wire \Tile_X4Y14_S4BEG[6] ;
 wire \Tile_X4Y14_S4BEG[7] ;
 wire \Tile_X4Y14_S4BEG[8] ;
 wire \Tile_X4Y14_S4BEG[9] ;
 wire \Tile_X4Y14_SS4BEG[0] ;
 wire \Tile_X4Y14_SS4BEG[10] ;
 wire \Tile_X4Y14_SS4BEG[11] ;
 wire \Tile_X4Y14_SS4BEG[12] ;
 wire \Tile_X4Y14_SS4BEG[13] ;
 wire \Tile_X4Y14_SS4BEG[14] ;
 wire \Tile_X4Y14_SS4BEG[15] ;
 wire \Tile_X4Y14_SS4BEG[1] ;
 wire \Tile_X4Y14_SS4BEG[2] ;
 wire \Tile_X4Y14_SS4BEG[3] ;
 wire \Tile_X4Y14_SS4BEG[4] ;
 wire \Tile_X4Y14_SS4BEG[5] ;
 wire \Tile_X4Y14_SS4BEG[6] ;
 wire \Tile_X4Y14_SS4BEG[7] ;
 wire \Tile_X4Y14_SS4BEG[8] ;
 wire \Tile_X4Y14_SS4BEG[9] ;
 wire Tile_X4Y14_UserCLKo;
 wire \Tile_X4Y14_W1BEG[0] ;
 wire \Tile_X4Y14_W1BEG[1] ;
 wire \Tile_X4Y14_W1BEG[2] ;
 wire \Tile_X4Y14_W1BEG[3] ;
 wire \Tile_X4Y14_W2BEG[0] ;
 wire \Tile_X4Y14_W2BEG[1] ;
 wire \Tile_X4Y14_W2BEG[2] ;
 wire \Tile_X4Y14_W2BEG[3] ;
 wire \Tile_X4Y14_W2BEG[4] ;
 wire \Tile_X4Y14_W2BEG[5] ;
 wire \Tile_X4Y14_W2BEG[6] ;
 wire \Tile_X4Y14_W2BEG[7] ;
 wire \Tile_X4Y14_W2BEGb[0] ;
 wire \Tile_X4Y14_W2BEGb[1] ;
 wire \Tile_X4Y14_W2BEGb[2] ;
 wire \Tile_X4Y14_W2BEGb[3] ;
 wire \Tile_X4Y14_W2BEGb[4] ;
 wire \Tile_X4Y14_W2BEGb[5] ;
 wire \Tile_X4Y14_W2BEGb[6] ;
 wire \Tile_X4Y14_W2BEGb[7] ;
 wire \Tile_X4Y14_W6BEG[0] ;
 wire \Tile_X4Y14_W6BEG[10] ;
 wire \Tile_X4Y14_W6BEG[11] ;
 wire \Tile_X4Y14_W6BEG[1] ;
 wire \Tile_X4Y14_W6BEG[2] ;
 wire \Tile_X4Y14_W6BEG[3] ;
 wire \Tile_X4Y14_W6BEG[4] ;
 wire \Tile_X4Y14_W6BEG[5] ;
 wire \Tile_X4Y14_W6BEG[6] ;
 wire \Tile_X4Y14_W6BEG[7] ;
 wire \Tile_X4Y14_W6BEG[8] ;
 wire \Tile_X4Y14_W6BEG[9] ;
 wire \Tile_X4Y14_WW4BEG[0] ;
 wire \Tile_X4Y14_WW4BEG[10] ;
 wire \Tile_X4Y14_WW4BEG[11] ;
 wire \Tile_X4Y14_WW4BEG[12] ;
 wire \Tile_X4Y14_WW4BEG[13] ;
 wire \Tile_X4Y14_WW4BEG[14] ;
 wire \Tile_X4Y14_WW4BEG[15] ;
 wire \Tile_X4Y14_WW4BEG[1] ;
 wire \Tile_X4Y14_WW4BEG[2] ;
 wire \Tile_X4Y14_WW4BEG[3] ;
 wire \Tile_X4Y14_WW4BEG[4] ;
 wire \Tile_X4Y14_WW4BEG[5] ;
 wire \Tile_X4Y14_WW4BEG[6] ;
 wire \Tile_X4Y14_WW4BEG[7] ;
 wire \Tile_X4Y14_WW4BEG[8] ;
 wire \Tile_X4Y14_WW4BEG[9] ;
 wire \Tile_X4Y15_FrameData_O[0] ;
 wire \Tile_X4Y15_FrameData_O[10] ;
 wire \Tile_X4Y15_FrameData_O[11] ;
 wire \Tile_X4Y15_FrameData_O[12] ;
 wire \Tile_X4Y15_FrameData_O[13] ;
 wire \Tile_X4Y15_FrameData_O[14] ;
 wire \Tile_X4Y15_FrameData_O[15] ;
 wire \Tile_X4Y15_FrameData_O[16] ;
 wire \Tile_X4Y15_FrameData_O[17] ;
 wire \Tile_X4Y15_FrameData_O[18] ;
 wire \Tile_X4Y15_FrameData_O[19] ;
 wire \Tile_X4Y15_FrameData_O[1] ;
 wire \Tile_X4Y15_FrameData_O[20] ;
 wire \Tile_X4Y15_FrameData_O[21] ;
 wire \Tile_X4Y15_FrameData_O[22] ;
 wire \Tile_X4Y15_FrameData_O[23] ;
 wire \Tile_X4Y15_FrameData_O[24] ;
 wire \Tile_X4Y15_FrameData_O[25] ;
 wire \Tile_X4Y15_FrameData_O[26] ;
 wire \Tile_X4Y15_FrameData_O[27] ;
 wire \Tile_X4Y15_FrameData_O[28] ;
 wire \Tile_X4Y15_FrameData_O[29] ;
 wire \Tile_X4Y15_FrameData_O[2] ;
 wire \Tile_X4Y15_FrameData_O[30] ;
 wire \Tile_X4Y15_FrameData_O[31] ;
 wire \Tile_X4Y15_FrameData_O[3] ;
 wire \Tile_X4Y15_FrameData_O[4] ;
 wire \Tile_X4Y15_FrameData_O[5] ;
 wire \Tile_X4Y15_FrameData_O[6] ;
 wire \Tile_X4Y15_FrameData_O[7] ;
 wire \Tile_X4Y15_FrameData_O[8] ;
 wire \Tile_X4Y15_FrameData_O[9] ;
 wire \Tile_X4Y15_FrameStrobe_O[0] ;
 wire \Tile_X4Y15_FrameStrobe_O[10] ;
 wire \Tile_X4Y15_FrameStrobe_O[11] ;
 wire \Tile_X4Y15_FrameStrobe_O[12] ;
 wire \Tile_X4Y15_FrameStrobe_O[13] ;
 wire \Tile_X4Y15_FrameStrobe_O[14] ;
 wire \Tile_X4Y15_FrameStrobe_O[15] ;
 wire \Tile_X4Y15_FrameStrobe_O[16] ;
 wire \Tile_X4Y15_FrameStrobe_O[17] ;
 wire \Tile_X4Y15_FrameStrobe_O[18] ;
 wire \Tile_X4Y15_FrameStrobe_O[19] ;
 wire \Tile_X4Y15_FrameStrobe_O[1] ;
 wire \Tile_X4Y15_FrameStrobe_O[2] ;
 wire \Tile_X4Y15_FrameStrobe_O[3] ;
 wire \Tile_X4Y15_FrameStrobe_O[4] ;
 wire \Tile_X4Y15_FrameStrobe_O[5] ;
 wire \Tile_X4Y15_FrameStrobe_O[6] ;
 wire \Tile_X4Y15_FrameStrobe_O[7] ;
 wire \Tile_X4Y15_FrameStrobe_O[8] ;
 wire \Tile_X4Y15_FrameStrobe_O[9] ;
 wire \Tile_X4Y15_N1BEG[0] ;
 wire \Tile_X4Y15_N1BEG[1] ;
 wire \Tile_X4Y15_N1BEG[2] ;
 wire \Tile_X4Y15_N1BEG[3] ;
 wire \Tile_X4Y15_N2BEG[0] ;
 wire \Tile_X4Y15_N2BEG[1] ;
 wire \Tile_X4Y15_N2BEG[2] ;
 wire \Tile_X4Y15_N2BEG[3] ;
 wire \Tile_X4Y15_N2BEG[4] ;
 wire \Tile_X4Y15_N2BEG[5] ;
 wire \Tile_X4Y15_N2BEG[6] ;
 wire \Tile_X4Y15_N2BEG[7] ;
 wire \Tile_X4Y15_N2BEGb[0] ;
 wire \Tile_X4Y15_N2BEGb[1] ;
 wire \Tile_X4Y15_N2BEGb[2] ;
 wire \Tile_X4Y15_N2BEGb[3] ;
 wire \Tile_X4Y15_N2BEGb[4] ;
 wire \Tile_X4Y15_N2BEGb[5] ;
 wire \Tile_X4Y15_N2BEGb[6] ;
 wire \Tile_X4Y15_N2BEGb[7] ;
 wire \Tile_X4Y15_N4BEG[0] ;
 wire \Tile_X4Y15_N4BEG[10] ;
 wire \Tile_X4Y15_N4BEG[11] ;
 wire \Tile_X4Y15_N4BEG[12] ;
 wire \Tile_X4Y15_N4BEG[13] ;
 wire \Tile_X4Y15_N4BEG[14] ;
 wire \Tile_X4Y15_N4BEG[15] ;
 wire \Tile_X4Y15_N4BEG[1] ;
 wire \Tile_X4Y15_N4BEG[2] ;
 wire \Tile_X4Y15_N4BEG[3] ;
 wire \Tile_X4Y15_N4BEG[4] ;
 wire \Tile_X4Y15_N4BEG[5] ;
 wire \Tile_X4Y15_N4BEG[6] ;
 wire \Tile_X4Y15_N4BEG[7] ;
 wire \Tile_X4Y15_N4BEG[8] ;
 wire \Tile_X4Y15_N4BEG[9] ;
 wire \Tile_X4Y15_NN4BEG[0] ;
 wire \Tile_X4Y15_NN4BEG[10] ;
 wire \Tile_X4Y15_NN4BEG[11] ;
 wire \Tile_X4Y15_NN4BEG[12] ;
 wire \Tile_X4Y15_NN4BEG[13] ;
 wire \Tile_X4Y15_NN4BEG[14] ;
 wire \Tile_X4Y15_NN4BEG[15] ;
 wire \Tile_X4Y15_NN4BEG[1] ;
 wire \Tile_X4Y15_NN4BEG[2] ;
 wire \Tile_X4Y15_NN4BEG[3] ;
 wire \Tile_X4Y15_NN4BEG[4] ;
 wire \Tile_X4Y15_NN4BEG[5] ;
 wire \Tile_X4Y15_NN4BEG[6] ;
 wire \Tile_X4Y15_NN4BEG[7] ;
 wire \Tile_X4Y15_NN4BEG[8] ;
 wire \Tile_X4Y15_NN4BEG[9] ;
 wire Tile_X4Y15_UserCLKo;
 wire \Tile_X4Y1_E1BEG[0] ;
 wire \Tile_X4Y1_E1BEG[1] ;
 wire \Tile_X4Y1_E1BEG[2] ;
 wire \Tile_X4Y1_E1BEG[3] ;
 wire \Tile_X4Y1_E2BEG[0] ;
 wire \Tile_X4Y1_E2BEG[1] ;
 wire \Tile_X4Y1_E2BEG[2] ;
 wire \Tile_X4Y1_E2BEG[3] ;
 wire \Tile_X4Y1_E2BEG[4] ;
 wire \Tile_X4Y1_E2BEG[5] ;
 wire \Tile_X4Y1_E2BEG[6] ;
 wire \Tile_X4Y1_E2BEG[7] ;
 wire \Tile_X4Y1_E2BEGb[0] ;
 wire \Tile_X4Y1_E2BEGb[1] ;
 wire \Tile_X4Y1_E2BEGb[2] ;
 wire \Tile_X4Y1_E2BEGb[3] ;
 wire \Tile_X4Y1_E2BEGb[4] ;
 wire \Tile_X4Y1_E2BEGb[5] ;
 wire \Tile_X4Y1_E2BEGb[6] ;
 wire \Tile_X4Y1_E2BEGb[7] ;
 wire \Tile_X4Y1_E6BEG[0] ;
 wire \Tile_X4Y1_E6BEG[10] ;
 wire \Tile_X4Y1_E6BEG[11] ;
 wire \Tile_X4Y1_E6BEG[1] ;
 wire \Tile_X4Y1_E6BEG[2] ;
 wire \Tile_X4Y1_E6BEG[3] ;
 wire \Tile_X4Y1_E6BEG[4] ;
 wire \Tile_X4Y1_E6BEG[5] ;
 wire \Tile_X4Y1_E6BEG[6] ;
 wire \Tile_X4Y1_E6BEG[7] ;
 wire \Tile_X4Y1_E6BEG[8] ;
 wire \Tile_X4Y1_E6BEG[9] ;
 wire \Tile_X4Y1_EE4BEG[0] ;
 wire \Tile_X4Y1_EE4BEG[10] ;
 wire \Tile_X4Y1_EE4BEG[11] ;
 wire \Tile_X4Y1_EE4BEG[12] ;
 wire \Tile_X4Y1_EE4BEG[13] ;
 wire \Tile_X4Y1_EE4BEG[14] ;
 wire \Tile_X4Y1_EE4BEG[15] ;
 wire \Tile_X4Y1_EE4BEG[1] ;
 wire \Tile_X4Y1_EE4BEG[2] ;
 wire \Tile_X4Y1_EE4BEG[3] ;
 wire \Tile_X4Y1_EE4BEG[4] ;
 wire \Tile_X4Y1_EE4BEG[5] ;
 wire \Tile_X4Y1_EE4BEG[6] ;
 wire \Tile_X4Y1_EE4BEG[7] ;
 wire \Tile_X4Y1_EE4BEG[8] ;
 wire \Tile_X4Y1_EE4BEG[9] ;
 wire \Tile_X4Y1_FrameData_O[0] ;
 wire \Tile_X4Y1_FrameData_O[10] ;
 wire \Tile_X4Y1_FrameData_O[11] ;
 wire \Tile_X4Y1_FrameData_O[12] ;
 wire \Tile_X4Y1_FrameData_O[13] ;
 wire \Tile_X4Y1_FrameData_O[14] ;
 wire \Tile_X4Y1_FrameData_O[15] ;
 wire \Tile_X4Y1_FrameData_O[16] ;
 wire \Tile_X4Y1_FrameData_O[17] ;
 wire \Tile_X4Y1_FrameData_O[18] ;
 wire \Tile_X4Y1_FrameData_O[19] ;
 wire \Tile_X4Y1_FrameData_O[1] ;
 wire \Tile_X4Y1_FrameData_O[20] ;
 wire \Tile_X4Y1_FrameData_O[21] ;
 wire \Tile_X4Y1_FrameData_O[22] ;
 wire \Tile_X4Y1_FrameData_O[23] ;
 wire \Tile_X4Y1_FrameData_O[24] ;
 wire \Tile_X4Y1_FrameData_O[25] ;
 wire \Tile_X4Y1_FrameData_O[26] ;
 wire \Tile_X4Y1_FrameData_O[27] ;
 wire \Tile_X4Y1_FrameData_O[28] ;
 wire \Tile_X4Y1_FrameData_O[29] ;
 wire \Tile_X4Y1_FrameData_O[2] ;
 wire \Tile_X4Y1_FrameData_O[30] ;
 wire \Tile_X4Y1_FrameData_O[31] ;
 wire \Tile_X4Y1_FrameData_O[3] ;
 wire \Tile_X4Y1_FrameData_O[4] ;
 wire \Tile_X4Y1_FrameData_O[5] ;
 wire \Tile_X4Y1_FrameData_O[6] ;
 wire \Tile_X4Y1_FrameData_O[7] ;
 wire \Tile_X4Y1_FrameData_O[8] ;
 wire \Tile_X4Y1_FrameData_O[9] ;
 wire \Tile_X4Y1_FrameStrobe_O[0] ;
 wire \Tile_X4Y1_FrameStrobe_O[10] ;
 wire \Tile_X4Y1_FrameStrobe_O[11] ;
 wire \Tile_X4Y1_FrameStrobe_O[12] ;
 wire \Tile_X4Y1_FrameStrobe_O[13] ;
 wire \Tile_X4Y1_FrameStrobe_O[14] ;
 wire \Tile_X4Y1_FrameStrobe_O[15] ;
 wire \Tile_X4Y1_FrameStrobe_O[16] ;
 wire \Tile_X4Y1_FrameStrobe_O[17] ;
 wire \Tile_X4Y1_FrameStrobe_O[18] ;
 wire \Tile_X4Y1_FrameStrobe_O[19] ;
 wire \Tile_X4Y1_FrameStrobe_O[1] ;
 wire \Tile_X4Y1_FrameStrobe_O[2] ;
 wire \Tile_X4Y1_FrameStrobe_O[3] ;
 wire \Tile_X4Y1_FrameStrobe_O[4] ;
 wire \Tile_X4Y1_FrameStrobe_O[5] ;
 wire \Tile_X4Y1_FrameStrobe_O[6] ;
 wire \Tile_X4Y1_FrameStrobe_O[7] ;
 wire \Tile_X4Y1_FrameStrobe_O[8] ;
 wire \Tile_X4Y1_FrameStrobe_O[9] ;
 wire \Tile_X4Y1_N1BEG[0] ;
 wire \Tile_X4Y1_N1BEG[1] ;
 wire \Tile_X4Y1_N1BEG[2] ;
 wire \Tile_X4Y1_N1BEG[3] ;
 wire \Tile_X4Y1_N2BEG[0] ;
 wire \Tile_X4Y1_N2BEG[1] ;
 wire \Tile_X4Y1_N2BEG[2] ;
 wire \Tile_X4Y1_N2BEG[3] ;
 wire \Tile_X4Y1_N2BEG[4] ;
 wire \Tile_X4Y1_N2BEG[5] ;
 wire \Tile_X4Y1_N2BEG[6] ;
 wire \Tile_X4Y1_N2BEG[7] ;
 wire \Tile_X4Y1_N2BEGb[0] ;
 wire \Tile_X4Y1_N2BEGb[1] ;
 wire \Tile_X4Y1_N2BEGb[2] ;
 wire \Tile_X4Y1_N2BEGb[3] ;
 wire \Tile_X4Y1_N2BEGb[4] ;
 wire \Tile_X4Y1_N2BEGb[5] ;
 wire \Tile_X4Y1_N2BEGb[6] ;
 wire \Tile_X4Y1_N2BEGb[7] ;
 wire \Tile_X4Y1_N4BEG[0] ;
 wire \Tile_X4Y1_N4BEG[10] ;
 wire \Tile_X4Y1_N4BEG[11] ;
 wire \Tile_X4Y1_N4BEG[12] ;
 wire \Tile_X4Y1_N4BEG[13] ;
 wire \Tile_X4Y1_N4BEG[14] ;
 wire \Tile_X4Y1_N4BEG[15] ;
 wire \Tile_X4Y1_N4BEG[1] ;
 wire \Tile_X4Y1_N4BEG[2] ;
 wire \Tile_X4Y1_N4BEG[3] ;
 wire \Tile_X4Y1_N4BEG[4] ;
 wire \Tile_X4Y1_N4BEG[5] ;
 wire \Tile_X4Y1_N4BEG[6] ;
 wire \Tile_X4Y1_N4BEG[7] ;
 wire \Tile_X4Y1_N4BEG[8] ;
 wire \Tile_X4Y1_N4BEG[9] ;
 wire \Tile_X4Y1_NN4BEG[0] ;
 wire \Tile_X4Y1_NN4BEG[10] ;
 wire \Tile_X4Y1_NN4BEG[11] ;
 wire \Tile_X4Y1_NN4BEG[12] ;
 wire \Tile_X4Y1_NN4BEG[13] ;
 wire \Tile_X4Y1_NN4BEG[14] ;
 wire \Tile_X4Y1_NN4BEG[15] ;
 wire \Tile_X4Y1_NN4BEG[1] ;
 wire \Tile_X4Y1_NN4BEG[2] ;
 wire \Tile_X4Y1_NN4BEG[3] ;
 wire \Tile_X4Y1_NN4BEG[4] ;
 wire \Tile_X4Y1_NN4BEG[5] ;
 wire \Tile_X4Y1_NN4BEG[6] ;
 wire \Tile_X4Y1_NN4BEG[7] ;
 wire \Tile_X4Y1_NN4BEG[8] ;
 wire \Tile_X4Y1_NN4BEG[9] ;
 wire \Tile_X4Y1_S1BEG[0] ;
 wire \Tile_X4Y1_S1BEG[1] ;
 wire \Tile_X4Y1_S1BEG[2] ;
 wire \Tile_X4Y1_S1BEG[3] ;
 wire \Tile_X4Y1_S2BEG[0] ;
 wire \Tile_X4Y1_S2BEG[1] ;
 wire \Tile_X4Y1_S2BEG[2] ;
 wire \Tile_X4Y1_S2BEG[3] ;
 wire \Tile_X4Y1_S2BEG[4] ;
 wire \Tile_X4Y1_S2BEG[5] ;
 wire \Tile_X4Y1_S2BEG[6] ;
 wire \Tile_X4Y1_S2BEG[7] ;
 wire \Tile_X4Y1_S2BEGb[0] ;
 wire \Tile_X4Y1_S2BEGb[1] ;
 wire \Tile_X4Y1_S2BEGb[2] ;
 wire \Tile_X4Y1_S2BEGb[3] ;
 wire \Tile_X4Y1_S2BEGb[4] ;
 wire \Tile_X4Y1_S2BEGb[5] ;
 wire \Tile_X4Y1_S2BEGb[6] ;
 wire \Tile_X4Y1_S2BEGb[7] ;
 wire \Tile_X4Y1_S4BEG[0] ;
 wire \Tile_X4Y1_S4BEG[10] ;
 wire \Tile_X4Y1_S4BEG[11] ;
 wire \Tile_X4Y1_S4BEG[12] ;
 wire \Tile_X4Y1_S4BEG[13] ;
 wire \Tile_X4Y1_S4BEG[14] ;
 wire \Tile_X4Y1_S4BEG[15] ;
 wire \Tile_X4Y1_S4BEG[1] ;
 wire \Tile_X4Y1_S4BEG[2] ;
 wire \Tile_X4Y1_S4BEG[3] ;
 wire \Tile_X4Y1_S4BEG[4] ;
 wire \Tile_X4Y1_S4BEG[5] ;
 wire \Tile_X4Y1_S4BEG[6] ;
 wire \Tile_X4Y1_S4BEG[7] ;
 wire \Tile_X4Y1_S4BEG[8] ;
 wire \Tile_X4Y1_S4BEG[9] ;
 wire \Tile_X4Y1_SS4BEG[0] ;
 wire \Tile_X4Y1_SS4BEG[10] ;
 wire \Tile_X4Y1_SS4BEG[11] ;
 wire \Tile_X4Y1_SS4BEG[12] ;
 wire \Tile_X4Y1_SS4BEG[13] ;
 wire \Tile_X4Y1_SS4BEG[14] ;
 wire \Tile_X4Y1_SS4BEG[15] ;
 wire \Tile_X4Y1_SS4BEG[1] ;
 wire \Tile_X4Y1_SS4BEG[2] ;
 wire \Tile_X4Y1_SS4BEG[3] ;
 wire \Tile_X4Y1_SS4BEG[4] ;
 wire \Tile_X4Y1_SS4BEG[5] ;
 wire \Tile_X4Y1_SS4BEG[6] ;
 wire \Tile_X4Y1_SS4BEG[7] ;
 wire \Tile_X4Y1_SS4BEG[8] ;
 wire \Tile_X4Y1_SS4BEG[9] ;
 wire Tile_X4Y1_UserCLKo;
 wire \Tile_X4Y1_W1BEG[0] ;
 wire \Tile_X4Y1_W1BEG[1] ;
 wire \Tile_X4Y1_W1BEG[2] ;
 wire \Tile_X4Y1_W1BEG[3] ;
 wire \Tile_X4Y1_W2BEG[0] ;
 wire \Tile_X4Y1_W2BEG[1] ;
 wire \Tile_X4Y1_W2BEG[2] ;
 wire \Tile_X4Y1_W2BEG[3] ;
 wire \Tile_X4Y1_W2BEG[4] ;
 wire \Tile_X4Y1_W2BEG[5] ;
 wire \Tile_X4Y1_W2BEG[6] ;
 wire \Tile_X4Y1_W2BEG[7] ;
 wire \Tile_X4Y1_W2BEGb[0] ;
 wire \Tile_X4Y1_W2BEGb[1] ;
 wire \Tile_X4Y1_W2BEGb[2] ;
 wire \Tile_X4Y1_W2BEGb[3] ;
 wire \Tile_X4Y1_W2BEGb[4] ;
 wire \Tile_X4Y1_W2BEGb[5] ;
 wire \Tile_X4Y1_W2BEGb[6] ;
 wire \Tile_X4Y1_W2BEGb[7] ;
 wire \Tile_X4Y1_W6BEG[0] ;
 wire \Tile_X4Y1_W6BEG[10] ;
 wire \Tile_X4Y1_W6BEG[11] ;
 wire \Tile_X4Y1_W6BEG[1] ;
 wire \Tile_X4Y1_W6BEG[2] ;
 wire \Tile_X4Y1_W6BEG[3] ;
 wire \Tile_X4Y1_W6BEG[4] ;
 wire \Tile_X4Y1_W6BEG[5] ;
 wire \Tile_X4Y1_W6BEG[6] ;
 wire \Tile_X4Y1_W6BEG[7] ;
 wire \Tile_X4Y1_W6BEG[8] ;
 wire \Tile_X4Y1_W6BEG[9] ;
 wire \Tile_X4Y1_WW4BEG[0] ;
 wire \Tile_X4Y1_WW4BEG[10] ;
 wire \Tile_X4Y1_WW4BEG[11] ;
 wire \Tile_X4Y1_WW4BEG[12] ;
 wire \Tile_X4Y1_WW4BEG[13] ;
 wire \Tile_X4Y1_WW4BEG[14] ;
 wire \Tile_X4Y1_WW4BEG[15] ;
 wire \Tile_X4Y1_WW4BEG[1] ;
 wire \Tile_X4Y1_WW4BEG[2] ;
 wire \Tile_X4Y1_WW4BEG[3] ;
 wire \Tile_X4Y1_WW4BEG[4] ;
 wire \Tile_X4Y1_WW4BEG[5] ;
 wire \Tile_X4Y1_WW4BEG[6] ;
 wire \Tile_X4Y1_WW4BEG[7] ;
 wire \Tile_X4Y1_WW4BEG[8] ;
 wire \Tile_X4Y1_WW4BEG[9] ;
 wire \Tile_X4Y2_E1BEG[0] ;
 wire \Tile_X4Y2_E1BEG[1] ;
 wire \Tile_X4Y2_E1BEG[2] ;
 wire \Tile_X4Y2_E1BEG[3] ;
 wire \Tile_X4Y2_E2BEG[0] ;
 wire \Tile_X4Y2_E2BEG[1] ;
 wire \Tile_X4Y2_E2BEG[2] ;
 wire \Tile_X4Y2_E2BEG[3] ;
 wire \Tile_X4Y2_E2BEG[4] ;
 wire \Tile_X4Y2_E2BEG[5] ;
 wire \Tile_X4Y2_E2BEG[6] ;
 wire \Tile_X4Y2_E2BEG[7] ;
 wire \Tile_X4Y2_E2BEGb[0] ;
 wire \Tile_X4Y2_E2BEGb[1] ;
 wire \Tile_X4Y2_E2BEGb[2] ;
 wire \Tile_X4Y2_E2BEGb[3] ;
 wire \Tile_X4Y2_E2BEGb[4] ;
 wire \Tile_X4Y2_E2BEGb[5] ;
 wire \Tile_X4Y2_E2BEGb[6] ;
 wire \Tile_X4Y2_E2BEGb[7] ;
 wire \Tile_X4Y2_E6BEG[0] ;
 wire \Tile_X4Y2_E6BEG[10] ;
 wire \Tile_X4Y2_E6BEG[11] ;
 wire \Tile_X4Y2_E6BEG[1] ;
 wire \Tile_X4Y2_E6BEG[2] ;
 wire \Tile_X4Y2_E6BEG[3] ;
 wire \Tile_X4Y2_E6BEG[4] ;
 wire \Tile_X4Y2_E6BEG[5] ;
 wire \Tile_X4Y2_E6BEG[6] ;
 wire \Tile_X4Y2_E6BEG[7] ;
 wire \Tile_X4Y2_E6BEG[8] ;
 wire \Tile_X4Y2_E6BEG[9] ;
 wire \Tile_X4Y2_EE4BEG[0] ;
 wire \Tile_X4Y2_EE4BEG[10] ;
 wire \Tile_X4Y2_EE4BEG[11] ;
 wire \Tile_X4Y2_EE4BEG[12] ;
 wire \Tile_X4Y2_EE4BEG[13] ;
 wire \Tile_X4Y2_EE4BEG[14] ;
 wire \Tile_X4Y2_EE4BEG[15] ;
 wire \Tile_X4Y2_EE4BEG[1] ;
 wire \Tile_X4Y2_EE4BEG[2] ;
 wire \Tile_X4Y2_EE4BEG[3] ;
 wire \Tile_X4Y2_EE4BEG[4] ;
 wire \Tile_X4Y2_EE4BEG[5] ;
 wire \Tile_X4Y2_EE4BEG[6] ;
 wire \Tile_X4Y2_EE4BEG[7] ;
 wire \Tile_X4Y2_EE4BEG[8] ;
 wire \Tile_X4Y2_EE4BEG[9] ;
 wire \Tile_X4Y2_FrameData_O[0] ;
 wire \Tile_X4Y2_FrameData_O[10] ;
 wire \Tile_X4Y2_FrameData_O[11] ;
 wire \Tile_X4Y2_FrameData_O[12] ;
 wire \Tile_X4Y2_FrameData_O[13] ;
 wire \Tile_X4Y2_FrameData_O[14] ;
 wire \Tile_X4Y2_FrameData_O[15] ;
 wire \Tile_X4Y2_FrameData_O[16] ;
 wire \Tile_X4Y2_FrameData_O[17] ;
 wire \Tile_X4Y2_FrameData_O[18] ;
 wire \Tile_X4Y2_FrameData_O[19] ;
 wire \Tile_X4Y2_FrameData_O[1] ;
 wire \Tile_X4Y2_FrameData_O[20] ;
 wire \Tile_X4Y2_FrameData_O[21] ;
 wire \Tile_X4Y2_FrameData_O[22] ;
 wire \Tile_X4Y2_FrameData_O[23] ;
 wire \Tile_X4Y2_FrameData_O[24] ;
 wire \Tile_X4Y2_FrameData_O[25] ;
 wire \Tile_X4Y2_FrameData_O[26] ;
 wire \Tile_X4Y2_FrameData_O[27] ;
 wire \Tile_X4Y2_FrameData_O[28] ;
 wire \Tile_X4Y2_FrameData_O[29] ;
 wire \Tile_X4Y2_FrameData_O[2] ;
 wire \Tile_X4Y2_FrameData_O[30] ;
 wire \Tile_X4Y2_FrameData_O[31] ;
 wire \Tile_X4Y2_FrameData_O[3] ;
 wire \Tile_X4Y2_FrameData_O[4] ;
 wire \Tile_X4Y2_FrameData_O[5] ;
 wire \Tile_X4Y2_FrameData_O[6] ;
 wire \Tile_X4Y2_FrameData_O[7] ;
 wire \Tile_X4Y2_FrameData_O[8] ;
 wire \Tile_X4Y2_FrameData_O[9] ;
 wire \Tile_X4Y2_FrameStrobe_O[0] ;
 wire \Tile_X4Y2_FrameStrobe_O[10] ;
 wire \Tile_X4Y2_FrameStrobe_O[11] ;
 wire \Tile_X4Y2_FrameStrobe_O[12] ;
 wire \Tile_X4Y2_FrameStrobe_O[13] ;
 wire \Tile_X4Y2_FrameStrobe_O[14] ;
 wire \Tile_X4Y2_FrameStrobe_O[15] ;
 wire \Tile_X4Y2_FrameStrobe_O[16] ;
 wire \Tile_X4Y2_FrameStrobe_O[17] ;
 wire \Tile_X4Y2_FrameStrobe_O[18] ;
 wire \Tile_X4Y2_FrameStrobe_O[19] ;
 wire \Tile_X4Y2_FrameStrobe_O[1] ;
 wire \Tile_X4Y2_FrameStrobe_O[2] ;
 wire \Tile_X4Y2_FrameStrobe_O[3] ;
 wire \Tile_X4Y2_FrameStrobe_O[4] ;
 wire \Tile_X4Y2_FrameStrobe_O[5] ;
 wire \Tile_X4Y2_FrameStrobe_O[6] ;
 wire \Tile_X4Y2_FrameStrobe_O[7] ;
 wire \Tile_X4Y2_FrameStrobe_O[8] ;
 wire \Tile_X4Y2_FrameStrobe_O[9] ;
 wire \Tile_X4Y2_N1BEG[0] ;
 wire \Tile_X4Y2_N1BEG[1] ;
 wire \Tile_X4Y2_N1BEG[2] ;
 wire \Tile_X4Y2_N1BEG[3] ;
 wire \Tile_X4Y2_N2BEG[0] ;
 wire \Tile_X4Y2_N2BEG[1] ;
 wire \Tile_X4Y2_N2BEG[2] ;
 wire \Tile_X4Y2_N2BEG[3] ;
 wire \Tile_X4Y2_N2BEG[4] ;
 wire \Tile_X4Y2_N2BEG[5] ;
 wire \Tile_X4Y2_N2BEG[6] ;
 wire \Tile_X4Y2_N2BEG[7] ;
 wire \Tile_X4Y2_N2BEGb[0] ;
 wire \Tile_X4Y2_N2BEGb[1] ;
 wire \Tile_X4Y2_N2BEGb[2] ;
 wire \Tile_X4Y2_N2BEGb[3] ;
 wire \Tile_X4Y2_N2BEGb[4] ;
 wire \Tile_X4Y2_N2BEGb[5] ;
 wire \Tile_X4Y2_N2BEGb[6] ;
 wire \Tile_X4Y2_N2BEGb[7] ;
 wire \Tile_X4Y2_N4BEG[0] ;
 wire \Tile_X4Y2_N4BEG[10] ;
 wire \Tile_X4Y2_N4BEG[11] ;
 wire \Tile_X4Y2_N4BEG[12] ;
 wire \Tile_X4Y2_N4BEG[13] ;
 wire \Tile_X4Y2_N4BEG[14] ;
 wire \Tile_X4Y2_N4BEG[15] ;
 wire \Tile_X4Y2_N4BEG[1] ;
 wire \Tile_X4Y2_N4BEG[2] ;
 wire \Tile_X4Y2_N4BEG[3] ;
 wire \Tile_X4Y2_N4BEG[4] ;
 wire \Tile_X4Y2_N4BEG[5] ;
 wire \Tile_X4Y2_N4BEG[6] ;
 wire \Tile_X4Y2_N4BEG[7] ;
 wire \Tile_X4Y2_N4BEG[8] ;
 wire \Tile_X4Y2_N4BEG[9] ;
 wire \Tile_X4Y2_NN4BEG[0] ;
 wire \Tile_X4Y2_NN4BEG[10] ;
 wire \Tile_X4Y2_NN4BEG[11] ;
 wire \Tile_X4Y2_NN4BEG[12] ;
 wire \Tile_X4Y2_NN4BEG[13] ;
 wire \Tile_X4Y2_NN4BEG[14] ;
 wire \Tile_X4Y2_NN4BEG[15] ;
 wire \Tile_X4Y2_NN4BEG[1] ;
 wire \Tile_X4Y2_NN4BEG[2] ;
 wire \Tile_X4Y2_NN4BEG[3] ;
 wire \Tile_X4Y2_NN4BEG[4] ;
 wire \Tile_X4Y2_NN4BEG[5] ;
 wire \Tile_X4Y2_NN4BEG[6] ;
 wire \Tile_X4Y2_NN4BEG[7] ;
 wire \Tile_X4Y2_NN4BEG[8] ;
 wire \Tile_X4Y2_NN4BEG[9] ;
 wire \Tile_X4Y2_S1BEG[0] ;
 wire \Tile_X4Y2_S1BEG[1] ;
 wire \Tile_X4Y2_S1BEG[2] ;
 wire \Tile_X4Y2_S1BEG[3] ;
 wire \Tile_X4Y2_S2BEG[0] ;
 wire \Tile_X4Y2_S2BEG[1] ;
 wire \Tile_X4Y2_S2BEG[2] ;
 wire \Tile_X4Y2_S2BEG[3] ;
 wire \Tile_X4Y2_S2BEG[4] ;
 wire \Tile_X4Y2_S2BEG[5] ;
 wire \Tile_X4Y2_S2BEG[6] ;
 wire \Tile_X4Y2_S2BEG[7] ;
 wire \Tile_X4Y2_S2BEGb[0] ;
 wire \Tile_X4Y2_S2BEGb[1] ;
 wire \Tile_X4Y2_S2BEGb[2] ;
 wire \Tile_X4Y2_S2BEGb[3] ;
 wire \Tile_X4Y2_S2BEGb[4] ;
 wire \Tile_X4Y2_S2BEGb[5] ;
 wire \Tile_X4Y2_S2BEGb[6] ;
 wire \Tile_X4Y2_S2BEGb[7] ;
 wire \Tile_X4Y2_S4BEG[0] ;
 wire \Tile_X4Y2_S4BEG[10] ;
 wire \Tile_X4Y2_S4BEG[11] ;
 wire \Tile_X4Y2_S4BEG[12] ;
 wire \Tile_X4Y2_S4BEG[13] ;
 wire \Tile_X4Y2_S4BEG[14] ;
 wire \Tile_X4Y2_S4BEG[15] ;
 wire \Tile_X4Y2_S4BEG[1] ;
 wire \Tile_X4Y2_S4BEG[2] ;
 wire \Tile_X4Y2_S4BEG[3] ;
 wire \Tile_X4Y2_S4BEG[4] ;
 wire \Tile_X4Y2_S4BEG[5] ;
 wire \Tile_X4Y2_S4BEG[6] ;
 wire \Tile_X4Y2_S4BEG[7] ;
 wire \Tile_X4Y2_S4BEG[8] ;
 wire \Tile_X4Y2_S4BEG[9] ;
 wire \Tile_X4Y2_SS4BEG[0] ;
 wire \Tile_X4Y2_SS4BEG[10] ;
 wire \Tile_X4Y2_SS4BEG[11] ;
 wire \Tile_X4Y2_SS4BEG[12] ;
 wire \Tile_X4Y2_SS4BEG[13] ;
 wire \Tile_X4Y2_SS4BEG[14] ;
 wire \Tile_X4Y2_SS4BEG[15] ;
 wire \Tile_X4Y2_SS4BEG[1] ;
 wire \Tile_X4Y2_SS4BEG[2] ;
 wire \Tile_X4Y2_SS4BEG[3] ;
 wire \Tile_X4Y2_SS4BEG[4] ;
 wire \Tile_X4Y2_SS4BEG[5] ;
 wire \Tile_X4Y2_SS4BEG[6] ;
 wire \Tile_X4Y2_SS4BEG[7] ;
 wire \Tile_X4Y2_SS4BEG[8] ;
 wire \Tile_X4Y2_SS4BEG[9] ;
 wire Tile_X4Y2_UserCLKo;
 wire \Tile_X4Y2_W1BEG[0] ;
 wire \Tile_X4Y2_W1BEG[1] ;
 wire \Tile_X4Y2_W1BEG[2] ;
 wire \Tile_X4Y2_W1BEG[3] ;
 wire \Tile_X4Y2_W2BEG[0] ;
 wire \Tile_X4Y2_W2BEG[1] ;
 wire \Tile_X4Y2_W2BEG[2] ;
 wire \Tile_X4Y2_W2BEG[3] ;
 wire \Tile_X4Y2_W2BEG[4] ;
 wire \Tile_X4Y2_W2BEG[5] ;
 wire \Tile_X4Y2_W2BEG[6] ;
 wire \Tile_X4Y2_W2BEG[7] ;
 wire \Tile_X4Y2_W2BEGb[0] ;
 wire \Tile_X4Y2_W2BEGb[1] ;
 wire \Tile_X4Y2_W2BEGb[2] ;
 wire \Tile_X4Y2_W2BEGb[3] ;
 wire \Tile_X4Y2_W2BEGb[4] ;
 wire \Tile_X4Y2_W2BEGb[5] ;
 wire \Tile_X4Y2_W2BEGb[6] ;
 wire \Tile_X4Y2_W2BEGb[7] ;
 wire \Tile_X4Y2_W6BEG[0] ;
 wire \Tile_X4Y2_W6BEG[10] ;
 wire \Tile_X4Y2_W6BEG[11] ;
 wire \Tile_X4Y2_W6BEG[1] ;
 wire \Tile_X4Y2_W6BEG[2] ;
 wire \Tile_X4Y2_W6BEG[3] ;
 wire \Tile_X4Y2_W6BEG[4] ;
 wire \Tile_X4Y2_W6BEG[5] ;
 wire \Tile_X4Y2_W6BEG[6] ;
 wire \Tile_X4Y2_W6BEG[7] ;
 wire \Tile_X4Y2_W6BEG[8] ;
 wire \Tile_X4Y2_W6BEG[9] ;
 wire \Tile_X4Y2_WW4BEG[0] ;
 wire \Tile_X4Y2_WW4BEG[10] ;
 wire \Tile_X4Y2_WW4BEG[11] ;
 wire \Tile_X4Y2_WW4BEG[12] ;
 wire \Tile_X4Y2_WW4BEG[13] ;
 wire \Tile_X4Y2_WW4BEG[14] ;
 wire \Tile_X4Y2_WW4BEG[15] ;
 wire \Tile_X4Y2_WW4BEG[1] ;
 wire \Tile_X4Y2_WW4BEG[2] ;
 wire \Tile_X4Y2_WW4BEG[3] ;
 wire \Tile_X4Y2_WW4BEG[4] ;
 wire \Tile_X4Y2_WW4BEG[5] ;
 wire \Tile_X4Y2_WW4BEG[6] ;
 wire \Tile_X4Y2_WW4BEG[7] ;
 wire \Tile_X4Y2_WW4BEG[8] ;
 wire \Tile_X4Y2_WW4BEG[9] ;
 wire \Tile_X4Y3_E1BEG[0] ;
 wire \Tile_X4Y3_E1BEG[1] ;
 wire \Tile_X4Y3_E1BEG[2] ;
 wire \Tile_X4Y3_E1BEG[3] ;
 wire \Tile_X4Y3_E2BEG[0] ;
 wire \Tile_X4Y3_E2BEG[1] ;
 wire \Tile_X4Y3_E2BEG[2] ;
 wire \Tile_X4Y3_E2BEG[3] ;
 wire \Tile_X4Y3_E2BEG[4] ;
 wire \Tile_X4Y3_E2BEG[5] ;
 wire \Tile_X4Y3_E2BEG[6] ;
 wire \Tile_X4Y3_E2BEG[7] ;
 wire \Tile_X4Y3_E2BEGb[0] ;
 wire \Tile_X4Y3_E2BEGb[1] ;
 wire \Tile_X4Y3_E2BEGb[2] ;
 wire \Tile_X4Y3_E2BEGb[3] ;
 wire \Tile_X4Y3_E2BEGb[4] ;
 wire \Tile_X4Y3_E2BEGb[5] ;
 wire \Tile_X4Y3_E2BEGb[6] ;
 wire \Tile_X4Y3_E2BEGb[7] ;
 wire \Tile_X4Y3_E6BEG[0] ;
 wire \Tile_X4Y3_E6BEG[10] ;
 wire \Tile_X4Y3_E6BEG[11] ;
 wire \Tile_X4Y3_E6BEG[1] ;
 wire \Tile_X4Y3_E6BEG[2] ;
 wire \Tile_X4Y3_E6BEG[3] ;
 wire \Tile_X4Y3_E6BEG[4] ;
 wire \Tile_X4Y3_E6BEG[5] ;
 wire \Tile_X4Y3_E6BEG[6] ;
 wire \Tile_X4Y3_E6BEG[7] ;
 wire \Tile_X4Y3_E6BEG[8] ;
 wire \Tile_X4Y3_E6BEG[9] ;
 wire \Tile_X4Y3_EE4BEG[0] ;
 wire \Tile_X4Y3_EE4BEG[10] ;
 wire \Tile_X4Y3_EE4BEG[11] ;
 wire \Tile_X4Y3_EE4BEG[12] ;
 wire \Tile_X4Y3_EE4BEG[13] ;
 wire \Tile_X4Y3_EE4BEG[14] ;
 wire \Tile_X4Y3_EE4BEG[15] ;
 wire \Tile_X4Y3_EE4BEG[1] ;
 wire \Tile_X4Y3_EE4BEG[2] ;
 wire \Tile_X4Y3_EE4BEG[3] ;
 wire \Tile_X4Y3_EE4BEG[4] ;
 wire \Tile_X4Y3_EE4BEG[5] ;
 wire \Tile_X4Y3_EE4BEG[6] ;
 wire \Tile_X4Y3_EE4BEG[7] ;
 wire \Tile_X4Y3_EE4BEG[8] ;
 wire \Tile_X4Y3_EE4BEG[9] ;
 wire \Tile_X4Y3_FrameData_O[0] ;
 wire \Tile_X4Y3_FrameData_O[10] ;
 wire \Tile_X4Y3_FrameData_O[11] ;
 wire \Tile_X4Y3_FrameData_O[12] ;
 wire \Tile_X4Y3_FrameData_O[13] ;
 wire \Tile_X4Y3_FrameData_O[14] ;
 wire \Tile_X4Y3_FrameData_O[15] ;
 wire \Tile_X4Y3_FrameData_O[16] ;
 wire \Tile_X4Y3_FrameData_O[17] ;
 wire \Tile_X4Y3_FrameData_O[18] ;
 wire \Tile_X4Y3_FrameData_O[19] ;
 wire \Tile_X4Y3_FrameData_O[1] ;
 wire \Tile_X4Y3_FrameData_O[20] ;
 wire \Tile_X4Y3_FrameData_O[21] ;
 wire \Tile_X4Y3_FrameData_O[22] ;
 wire \Tile_X4Y3_FrameData_O[23] ;
 wire \Tile_X4Y3_FrameData_O[24] ;
 wire \Tile_X4Y3_FrameData_O[25] ;
 wire \Tile_X4Y3_FrameData_O[26] ;
 wire \Tile_X4Y3_FrameData_O[27] ;
 wire \Tile_X4Y3_FrameData_O[28] ;
 wire \Tile_X4Y3_FrameData_O[29] ;
 wire \Tile_X4Y3_FrameData_O[2] ;
 wire \Tile_X4Y3_FrameData_O[30] ;
 wire \Tile_X4Y3_FrameData_O[31] ;
 wire \Tile_X4Y3_FrameData_O[3] ;
 wire \Tile_X4Y3_FrameData_O[4] ;
 wire \Tile_X4Y3_FrameData_O[5] ;
 wire \Tile_X4Y3_FrameData_O[6] ;
 wire \Tile_X4Y3_FrameData_O[7] ;
 wire \Tile_X4Y3_FrameData_O[8] ;
 wire \Tile_X4Y3_FrameData_O[9] ;
 wire \Tile_X4Y3_FrameStrobe_O[0] ;
 wire \Tile_X4Y3_FrameStrobe_O[10] ;
 wire \Tile_X4Y3_FrameStrobe_O[11] ;
 wire \Tile_X4Y3_FrameStrobe_O[12] ;
 wire \Tile_X4Y3_FrameStrobe_O[13] ;
 wire \Tile_X4Y3_FrameStrobe_O[14] ;
 wire \Tile_X4Y3_FrameStrobe_O[15] ;
 wire \Tile_X4Y3_FrameStrobe_O[16] ;
 wire \Tile_X4Y3_FrameStrobe_O[17] ;
 wire \Tile_X4Y3_FrameStrobe_O[18] ;
 wire \Tile_X4Y3_FrameStrobe_O[19] ;
 wire \Tile_X4Y3_FrameStrobe_O[1] ;
 wire \Tile_X4Y3_FrameStrobe_O[2] ;
 wire \Tile_X4Y3_FrameStrobe_O[3] ;
 wire \Tile_X4Y3_FrameStrobe_O[4] ;
 wire \Tile_X4Y3_FrameStrobe_O[5] ;
 wire \Tile_X4Y3_FrameStrobe_O[6] ;
 wire \Tile_X4Y3_FrameStrobe_O[7] ;
 wire \Tile_X4Y3_FrameStrobe_O[8] ;
 wire \Tile_X4Y3_FrameStrobe_O[9] ;
 wire \Tile_X4Y3_N1BEG[0] ;
 wire \Tile_X4Y3_N1BEG[1] ;
 wire \Tile_X4Y3_N1BEG[2] ;
 wire \Tile_X4Y3_N1BEG[3] ;
 wire \Tile_X4Y3_N2BEG[0] ;
 wire \Tile_X4Y3_N2BEG[1] ;
 wire \Tile_X4Y3_N2BEG[2] ;
 wire \Tile_X4Y3_N2BEG[3] ;
 wire \Tile_X4Y3_N2BEG[4] ;
 wire \Tile_X4Y3_N2BEG[5] ;
 wire \Tile_X4Y3_N2BEG[6] ;
 wire \Tile_X4Y3_N2BEG[7] ;
 wire \Tile_X4Y3_N2BEGb[0] ;
 wire \Tile_X4Y3_N2BEGb[1] ;
 wire \Tile_X4Y3_N2BEGb[2] ;
 wire \Tile_X4Y3_N2BEGb[3] ;
 wire \Tile_X4Y3_N2BEGb[4] ;
 wire \Tile_X4Y3_N2BEGb[5] ;
 wire \Tile_X4Y3_N2BEGb[6] ;
 wire \Tile_X4Y3_N2BEGb[7] ;
 wire \Tile_X4Y3_N4BEG[0] ;
 wire \Tile_X4Y3_N4BEG[10] ;
 wire \Tile_X4Y3_N4BEG[11] ;
 wire \Tile_X4Y3_N4BEG[12] ;
 wire \Tile_X4Y3_N4BEG[13] ;
 wire \Tile_X4Y3_N4BEG[14] ;
 wire \Tile_X4Y3_N4BEG[15] ;
 wire \Tile_X4Y3_N4BEG[1] ;
 wire \Tile_X4Y3_N4BEG[2] ;
 wire \Tile_X4Y3_N4BEG[3] ;
 wire \Tile_X4Y3_N4BEG[4] ;
 wire \Tile_X4Y3_N4BEG[5] ;
 wire \Tile_X4Y3_N4BEG[6] ;
 wire \Tile_X4Y3_N4BEG[7] ;
 wire \Tile_X4Y3_N4BEG[8] ;
 wire \Tile_X4Y3_N4BEG[9] ;
 wire \Tile_X4Y3_NN4BEG[0] ;
 wire \Tile_X4Y3_NN4BEG[10] ;
 wire \Tile_X4Y3_NN4BEG[11] ;
 wire \Tile_X4Y3_NN4BEG[12] ;
 wire \Tile_X4Y3_NN4BEG[13] ;
 wire \Tile_X4Y3_NN4BEG[14] ;
 wire \Tile_X4Y3_NN4BEG[15] ;
 wire \Tile_X4Y3_NN4BEG[1] ;
 wire \Tile_X4Y3_NN4BEG[2] ;
 wire \Tile_X4Y3_NN4BEG[3] ;
 wire \Tile_X4Y3_NN4BEG[4] ;
 wire \Tile_X4Y3_NN4BEG[5] ;
 wire \Tile_X4Y3_NN4BEG[6] ;
 wire \Tile_X4Y3_NN4BEG[7] ;
 wire \Tile_X4Y3_NN4BEG[8] ;
 wire \Tile_X4Y3_NN4BEG[9] ;
 wire \Tile_X4Y3_S1BEG[0] ;
 wire \Tile_X4Y3_S1BEG[1] ;
 wire \Tile_X4Y3_S1BEG[2] ;
 wire \Tile_X4Y3_S1BEG[3] ;
 wire \Tile_X4Y3_S2BEG[0] ;
 wire \Tile_X4Y3_S2BEG[1] ;
 wire \Tile_X4Y3_S2BEG[2] ;
 wire \Tile_X4Y3_S2BEG[3] ;
 wire \Tile_X4Y3_S2BEG[4] ;
 wire \Tile_X4Y3_S2BEG[5] ;
 wire \Tile_X4Y3_S2BEG[6] ;
 wire \Tile_X4Y3_S2BEG[7] ;
 wire \Tile_X4Y3_S2BEGb[0] ;
 wire \Tile_X4Y3_S2BEGb[1] ;
 wire \Tile_X4Y3_S2BEGb[2] ;
 wire \Tile_X4Y3_S2BEGb[3] ;
 wire \Tile_X4Y3_S2BEGb[4] ;
 wire \Tile_X4Y3_S2BEGb[5] ;
 wire \Tile_X4Y3_S2BEGb[6] ;
 wire \Tile_X4Y3_S2BEGb[7] ;
 wire \Tile_X4Y3_S4BEG[0] ;
 wire \Tile_X4Y3_S4BEG[10] ;
 wire \Tile_X4Y3_S4BEG[11] ;
 wire \Tile_X4Y3_S4BEG[12] ;
 wire \Tile_X4Y3_S4BEG[13] ;
 wire \Tile_X4Y3_S4BEG[14] ;
 wire \Tile_X4Y3_S4BEG[15] ;
 wire \Tile_X4Y3_S4BEG[1] ;
 wire \Tile_X4Y3_S4BEG[2] ;
 wire \Tile_X4Y3_S4BEG[3] ;
 wire \Tile_X4Y3_S4BEG[4] ;
 wire \Tile_X4Y3_S4BEG[5] ;
 wire \Tile_X4Y3_S4BEG[6] ;
 wire \Tile_X4Y3_S4BEG[7] ;
 wire \Tile_X4Y3_S4BEG[8] ;
 wire \Tile_X4Y3_S4BEG[9] ;
 wire \Tile_X4Y3_SS4BEG[0] ;
 wire \Tile_X4Y3_SS4BEG[10] ;
 wire \Tile_X4Y3_SS4BEG[11] ;
 wire \Tile_X4Y3_SS4BEG[12] ;
 wire \Tile_X4Y3_SS4BEG[13] ;
 wire \Tile_X4Y3_SS4BEG[14] ;
 wire \Tile_X4Y3_SS4BEG[15] ;
 wire \Tile_X4Y3_SS4BEG[1] ;
 wire \Tile_X4Y3_SS4BEG[2] ;
 wire \Tile_X4Y3_SS4BEG[3] ;
 wire \Tile_X4Y3_SS4BEG[4] ;
 wire \Tile_X4Y3_SS4BEG[5] ;
 wire \Tile_X4Y3_SS4BEG[6] ;
 wire \Tile_X4Y3_SS4BEG[7] ;
 wire \Tile_X4Y3_SS4BEG[8] ;
 wire \Tile_X4Y3_SS4BEG[9] ;
 wire Tile_X4Y3_UserCLKo;
 wire \Tile_X4Y3_W1BEG[0] ;
 wire \Tile_X4Y3_W1BEG[1] ;
 wire \Tile_X4Y3_W1BEG[2] ;
 wire \Tile_X4Y3_W1BEG[3] ;
 wire \Tile_X4Y3_W2BEG[0] ;
 wire \Tile_X4Y3_W2BEG[1] ;
 wire \Tile_X4Y3_W2BEG[2] ;
 wire \Tile_X4Y3_W2BEG[3] ;
 wire \Tile_X4Y3_W2BEG[4] ;
 wire \Tile_X4Y3_W2BEG[5] ;
 wire \Tile_X4Y3_W2BEG[6] ;
 wire \Tile_X4Y3_W2BEG[7] ;
 wire \Tile_X4Y3_W2BEGb[0] ;
 wire \Tile_X4Y3_W2BEGb[1] ;
 wire \Tile_X4Y3_W2BEGb[2] ;
 wire \Tile_X4Y3_W2BEGb[3] ;
 wire \Tile_X4Y3_W2BEGb[4] ;
 wire \Tile_X4Y3_W2BEGb[5] ;
 wire \Tile_X4Y3_W2BEGb[6] ;
 wire \Tile_X4Y3_W2BEGb[7] ;
 wire \Tile_X4Y3_W6BEG[0] ;
 wire \Tile_X4Y3_W6BEG[10] ;
 wire \Tile_X4Y3_W6BEG[11] ;
 wire \Tile_X4Y3_W6BEG[1] ;
 wire \Tile_X4Y3_W6BEG[2] ;
 wire \Tile_X4Y3_W6BEG[3] ;
 wire \Tile_X4Y3_W6BEG[4] ;
 wire \Tile_X4Y3_W6BEG[5] ;
 wire \Tile_X4Y3_W6BEG[6] ;
 wire \Tile_X4Y3_W6BEG[7] ;
 wire \Tile_X4Y3_W6BEG[8] ;
 wire \Tile_X4Y3_W6BEG[9] ;
 wire \Tile_X4Y3_WW4BEG[0] ;
 wire \Tile_X4Y3_WW4BEG[10] ;
 wire \Tile_X4Y3_WW4BEG[11] ;
 wire \Tile_X4Y3_WW4BEG[12] ;
 wire \Tile_X4Y3_WW4BEG[13] ;
 wire \Tile_X4Y3_WW4BEG[14] ;
 wire \Tile_X4Y3_WW4BEG[15] ;
 wire \Tile_X4Y3_WW4BEG[1] ;
 wire \Tile_X4Y3_WW4BEG[2] ;
 wire \Tile_X4Y3_WW4BEG[3] ;
 wire \Tile_X4Y3_WW4BEG[4] ;
 wire \Tile_X4Y3_WW4BEG[5] ;
 wire \Tile_X4Y3_WW4BEG[6] ;
 wire \Tile_X4Y3_WW4BEG[7] ;
 wire \Tile_X4Y3_WW4BEG[8] ;
 wire \Tile_X4Y3_WW4BEG[9] ;
 wire \Tile_X4Y4_E1BEG[0] ;
 wire \Tile_X4Y4_E1BEG[1] ;
 wire \Tile_X4Y4_E1BEG[2] ;
 wire \Tile_X4Y4_E1BEG[3] ;
 wire \Tile_X4Y4_E2BEG[0] ;
 wire \Tile_X4Y4_E2BEG[1] ;
 wire \Tile_X4Y4_E2BEG[2] ;
 wire \Tile_X4Y4_E2BEG[3] ;
 wire \Tile_X4Y4_E2BEG[4] ;
 wire \Tile_X4Y4_E2BEG[5] ;
 wire \Tile_X4Y4_E2BEG[6] ;
 wire \Tile_X4Y4_E2BEG[7] ;
 wire \Tile_X4Y4_E2BEGb[0] ;
 wire \Tile_X4Y4_E2BEGb[1] ;
 wire \Tile_X4Y4_E2BEGb[2] ;
 wire \Tile_X4Y4_E2BEGb[3] ;
 wire \Tile_X4Y4_E2BEGb[4] ;
 wire \Tile_X4Y4_E2BEGb[5] ;
 wire \Tile_X4Y4_E2BEGb[6] ;
 wire \Tile_X4Y4_E2BEGb[7] ;
 wire \Tile_X4Y4_E6BEG[0] ;
 wire \Tile_X4Y4_E6BEG[10] ;
 wire \Tile_X4Y4_E6BEG[11] ;
 wire \Tile_X4Y4_E6BEG[1] ;
 wire \Tile_X4Y4_E6BEG[2] ;
 wire \Tile_X4Y4_E6BEG[3] ;
 wire \Tile_X4Y4_E6BEG[4] ;
 wire \Tile_X4Y4_E6BEG[5] ;
 wire \Tile_X4Y4_E6BEG[6] ;
 wire \Tile_X4Y4_E6BEG[7] ;
 wire \Tile_X4Y4_E6BEG[8] ;
 wire \Tile_X4Y4_E6BEG[9] ;
 wire \Tile_X4Y4_EE4BEG[0] ;
 wire \Tile_X4Y4_EE4BEG[10] ;
 wire \Tile_X4Y4_EE4BEG[11] ;
 wire \Tile_X4Y4_EE4BEG[12] ;
 wire \Tile_X4Y4_EE4BEG[13] ;
 wire \Tile_X4Y4_EE4BEG[14] ;
 wire \Tile_X4Y4_EE4BEG[15] ;
 wire \Tile_X4Y4_EE4BEG[1] ;
 wire \Tile_X4Y4_EE4BEG[2] ;
 wire \Tile_X4Y4_EE4BEG[3] ;
 wire \Tile_X4Y4_EE4BEG[4] ;
 wire \Tile_X4Y4_EE4BEG[5] ;
 wire \Tile_X4Y4_EE4BEG[6] ;
 wire \Tile_X4Y4_EE4BEG[7] ;
 wire \Tile_X4Y4_EE4BEG[8] ;
 wire \Tile_X4Y4_EE4BEG[9] ;
 wire \Tile_X4Y4_FrameData_O[0] ;
 wire \Tile_X4Y4_FrameData_O[10] ;
 wire \Tile_X4Y4_FrameData_O[11] ;
 wire \Tile_X4Y4_FrameData_O[12] ;
 wire \Tile_X4Y4_FrameData_O[13] ;
 wire \Tile_X4Y4_FrameData_O[14] ;
 wire \Tile_X4Y4_FrameData_O[15] ;
 wire \Tile_X4Y4_FrameData_O[16] ;
 wire \Tile_X4Y4_FrameData_O[17] ;
 wire \Tile_X4Y4_FrameData_O[18] ;
 wire \Tile_X4Y4_FrameData_O[19] ;
 wire \Tile_X4Y4_FrameData_O[1] ;
 wire \Tile_X4Y4_FrameData_O[20] ;
 wire \Tile_X4Y4_FrameData_O[21] ;
 wire \Tile_X4Y4_FrameData_O[22] ;
 wire \Tile_X4Y4_FrameData_O[23] ;
 wire \Tile_X4Y4_FrameData_O[24] ;
 wire \Tile_X4Y4_FrameData_O[25] ;
 wire \Tile_X4Y4_FrameData_O[26] ;
 wire \Tile_X4Y4_FrameData_O[27] ;
 wire \Tile_X4Y4_FrameData_O[28] ;
 wire \Tile_X4Y4_FrameData_O[29] ;
 wire \Tile_X4Y4_FrameData_O[2] ;
 wire \Tile_X4Y4_FrameData_O[30] ;
 wire \Tile_X4Y4_FrameData_O[31] ;
 wire \Tile_X4Y4_FrameData_O[3] ;
 wire \Tile_X4Y4_FrameData_O[4] ;
 wire \Tile_X4Y4_FrameData_O[5] ;
 wire \Tile_X4Y4_FrameData_O[6] ;
 wire \Tile_X4Y4_FrameData_O[7] ;
 wire \Tile_X4Y4_FrameData_O[8] ;
 wire \Tile_X4Y4_FrameData_O[9] ;
 wire \Tile_X4Y4_FrameStrobe_O[0] ;
 wire \Tile_X4Y4_FrameStrobe_O[10] ;
 wire \Tile_X4Y4_FrameStrobe_O[11] ;
 wire \Tile_X4Y4_FrameStrobe_O[12] ;
 wire \Tile_X4Y4_FrameStrobe_O[13] ;
 wire \Tile_X4Y4_FrameStrobe_O[14] ;
 wire \Tile_X4Y4_FrameStrobe_O[15] ;
 wire \Tile_X4Y4_FrameStrobe_O[16] ;
 wire \Tile_X4Y4_FrameStrobe_O[17] ;
 wire \Tile_X4Y4_FrameStrobe_O[18] ;
 wire \Tile_X4Y4_FrameStrobe_O[19] ;
 wire \Tile_X4Y4_FrameStrobe_O[1] ;
 wire \Tile_X4Y4_FrameStrobe_O[2] ;
 wire \Tile_X4Y4_FrameStrobe_O[3] ;
 wire \Tile_X4Y4_FrameStrobe_O[4] ;
 wire \Tile_X4Y4_FrameStrobe_O[5] ;
 wire \Tile_X4Y4_FrameStrobe_O[6] ;
 wire \Tile_X4Y4_FrameStrobe_O[7] ;
 wire \Tile_X4Y4_FrameStrobe_O[8] ;
 wire \Tile_X4Y4_FrameStrobe_O[9] ;
 wire \Tile_X4Y4_N1BEG[0] ;
 wire \Tile_X4Y4_N1BEG[1] ;
 wire \Tile_X4Y4_N1BEG[2] ;
 wire \Tile_X4Y4_N1BEG[3] ;
 wire \Tile_X4Y4_N2BEG[0] ;
 wire \Tile_X4Y4_N2BEG[1] ;
 wire \Tile_X4Y4_N2BEG[2] ;
 wire \Tile_X4Y4_N2BEG[3] ;
 wire \Tile_X4Y4_N2BEG[4] ;
 wire \Tile_X4Y4_N2BEG[5] ;
 wire \Tile_X4Y4_N2BEG[6] ;
 wire \Tile_X4Y4_N2BEG[7] ;
 wire \Tile_X4Y4_N2BEGb[0] ;
 wire \Tile_X4Y4_N2BEGb[1] ;
 wire \Tile_X4Y4_N2BEGb[2] ;
 wire \Tile_X4Y4_N2BEGb[3] ;
 wire \Tile_X4Y4_N2BEGb[4] ;
 wire \Tile_X4Y4_N2BEGb[5] ;
 wire \Tile_X4Y4_N2BEGb[6] ;
 wire \Tile_X4Y4_N2BEGb[7] ;
 wire \Tile_X4Y4_N4BEG[0] ;
 wire \Tile_X4Y4_N4BEG[10] ;
 wire \Tile_X4Y4_N4BEG[11] ;
 wire \Tile_X4Y4_N4BEG[12] ;
 wire \Tile_X4Y4_N4BEG[13] ;
 wire \Tile_X4Y4_N4BEG[14] ;
 wire \Tile_X4Y4_N4BEG[15] ;
 wire \Tile_X4Y4_N4BEG[1] ;
 wire \Tile_X4Y4_N4BEG[2] ;
 wire \Tile_X4Y4_N4BEG[3] ;
 wire \Tile_X4Y4_N4BEG[4] ;
 wire \Tile_X4Y4_N4BEG[5] ;
 wire \Tile_X4Y4_N4BEG[6] ;
 wire \Tile_X4Y4_N4BEG[7] ;
 wire \Tile_X4Y4_N4BEG[8] ;
 wire \Tile_X4Y4_N4BEG[9] ;
 wire \Tile_X4Y4_NN4BEG[0] ;
 wire \Tile_X4Y4_NN4BEG[10] ;
 wire \Tile_X4Y4_NN4BEG[11] ;
 wire \Tile_X4Y4_NN4BEG[12] ;
 wire \Tile_X4Y4_NN4BEG[13] ;
 wire \Tile_X4Y4_NN4BEG[14] ;
 wire \Tile_X4Y4_NN4BEG[15] ;
 wire \Tile_X4Y4_NN4BEG[1] ;
 wire \Tile_X4Y4_NN4BEG[2] ;
 wire \Tile_X4Y4_NN4BEG[3] ;
 wire \Tile_X4Y4_NN4BEG[4] ;
 wire \Tile_X4Y4_NN4BEG[5] ;
 wire \Tile_X4Y4_NN4BEG[6] ;
 wire \Tile_X4Y4_NN4BEG[7] ;
 wire \Tile_X4Y4_NN4BEG[8] ;
 wire \Tile_X4Y4_NN4BEG[9] ;
 wire \Tile_X4Y4_S1BEG[0] ;
 wire \Tile_X4Y4_S1BEG[1] ;
 wire \Tile_X4Y4_S1BEG[2] ;
 wire \Tile_X4Y4_S1BEG[3] ;
 wire \Tile_X4Y4_S2BEG[0] ;
 wire \Tile_X4Y4_S2BEG[1] ;
 wire \Tile_X4Y4_S2BEG[2] ;
 wire \Tile_X4Y4_S2BEG[3] ;
 wire \Tile_X4Y4_S2BEG[4] ;
 wire \Tile_X4Y4_S2BEG[5] ;
 wire \Tile_X4Y4_S2BEG[6] ;
 wire \Tile_X4Y4_S2BEG[7] ;
 wire \Tile_X4Y4_S2BEGb[0] ;
 wire \Tile_X4Y4_S2BEGb[1] ;
 wire \Tile_X4Y4_S2BEGb[2] ;
 wire \Tile_X4Y4_S2BEGb[3] ;
 wire \Tile_X4Y4_S2BEGb[4] ;
 wire \Tile_X4Y4_S2BEGb[5] ;
 wire \Tile_X4Y4_S2BEGb[6] ;
 wire \Tile_X4Y4_S2BEGb[7] ;
 wire \Tile_X4Y4_S4BEG[0] ;
 wire \Tile_X4Y4_S4BEG[10] ;
 wire \Tile_X4Y4_S4BEG[11] ;
 wire \Tile_X4Y4_S4BEG[12] ;
 wire \Tile_X4Y4_S4BEG[13] ;
 wire \Tile_X4Y4_S4BEG[14] ;
 wire \Tile_X4Y4_S4BEG[15] ;
 wire \Tile_X4Y4_S4BEG[1] ;
 wire \Tile_X4Y4_S4BEG[2] ;
 wire \Tile_X4Y4_S4BEG[3] ;
 wire \Tile_X4Y4_S4BEG[4] ;
 wire \Tile_X4Y4_S4BEG[5] ;
 wire \Tile_X4Y4_S4BEG[6] ;
 wire \Tile_X4Y4_S4BEG[7] ;
 wire \Tile_X4Y4_S4BEG[8] ;
 wire \Tile_X4Y4_S4BEG[9] ;
 wire \Tile_X4Y4_SS4BEG[0] ;
 wire \Tile_X4Y4_SS4BEG[10] ;
 wire \Tile_X4Y4_SS4BEG[11] ;
 wire \Tile_X4Y4_SS4BEG[12] ;
 wire \Tile_X4Y4_SS4BEG[13] ;
 wire \Tile_X4Y4_SS4BEG[14] ;
 wire \Tile_X4Y4_SS4BEG[15] ;
 wire \Tile_X4Y4_SS4BEG[1] ;
 wire \Tile_X4Y4_SS4BEG[2] ;
 wire \Tile_X4Y4_SS4BEG[3] ;
 wire \Tile_X4Y4_SS4BEG[4] ;
 wire \Tile_X4Y4_SS4BEG[5] ;
 wire \Tile_X4Y4_SS4BEG[6] ;
 wire \Tile_X4Y4_SS4BEG[7] ;
 wire \Tile_X4Y4_SS4BEG[8] ;
 wire \Tile_X4Y4_SS4BEG[9] ;
 wire Tile_X4Y4_UserCLKo;
 wire \Tile_X4Y4_W1BEG[0] ;
 wire \Tile_X4Y4_W1BEG[1] ;
 wire \Tile_X4Y4_W1BEG[2] ;
 wire \Tile_X4Y4_W1BEG[3] ;
 wire \Tile_X4Y4_W2BEG[0] ;
 wire \Tile_X4Y4_W2BEG[1] ;
 wire \Tile_X4Y4_W2BEG[2] ;
 wire \Tile_X4Y4_W2BEG[3] ;
 wire \Tile_X4Y4_W2BEG[4] ;
 wire \Tile_X4Y4_W2BEG[5] ;
 wire \Tile_X4Y4_W2BEG[6] ;
 wire \Tile_X4Y4_W2BEG[7] ;
 wire \Tile_X4Y4_W2BEGb[0] ;
 wire \Tile_X4Y4_W2BEGb[1] ;
 wire \Tile_X4Y4_W2BEGb[2] ;
 wire \Tile_X4Y4_W2BEGb[3] ;
 wire \Tile_X4Y4_W2BEGb[4] ;
 wire \Tile_X4Y4_W2BEGb[5] ;
 wire \Tile_X4Y4_W2BEGb[6] ;
 wire \Tile_X4Y4_W2BEGb[7] ;
 wire \Tile_X4Y4_W6BEG[0] ;
 wire \Tile_X4Y4_W6BEG[10] ;
 wire \Tile_X4Y4_W6BEG[11] ;
 wire \Tile_X4Y4_W6BEG[1] ;
 wire \Tile_X4Y4_W6BEG[2] ;
 wire \Tile_X4Y4_W6BEG[3] ;
 wire \Tile_X4Y4_W6BEG[4] ;
 wire \Tile_X4Y4_W6BEG[5] ;
 wire \Tile_X4Y4_W6BEG[6] ;
 wire \Tile_X4Y4_W6BEG[7] ;
 wire \Tile_X4Y4_W6BEG[8] ;
 wire \Tile_X4Y4_W6BEG[9] ;
 wire \Tile_X4Y4_WW4BEG[0] ;
 wire \Tile_X4Y4_WW4BEG[10] ;
 wire \Tile_X4Y4_WW4BEG[11] ;
 wire \Tile_X4Y4_WW4BEG[12] ;
 wire \Tile_X4Y4_WW4BEG[13] ;
 wire \Tile_X4Y4_WW4BEG[14] ;
 wire \Tile_X4Y4_WW4BEG[15] ;
 wire \Tile_X4Y4_WW4BEG[1] ;
 wire \Tile_X4Y4_WW4BEG[2] ;
 wire \Tile_X4Y4_WW4BEG[3] ;
 wire \Tile_X4Y4_WW4BEG[4] ;
 wire \Tile_X4Y4_WW4BEG[5] ;
 wire \Tile_X4Y4_WW4BEG[6] ;
 wire \Tile_X4Y4_WW4BEG[7] ;
 wire \Tile_X4Y4_WW4BEG[8] ;
 wire \Tile_X4Y4_WW4BEG[9] ;
 wire \Tile_X4Y5_E1BEG[0] ;
 wire \Tile_X4Y5_E1BEG[1] ;
 wire \Tile_X4Y5_E1BEG[2] ;
 wire \Tile_X4Y5_E1BEG[3] ;
 wire \Tile_X4Y5_E2BEG[0] ;
 wire \Tile_X4Y5_E2BEG[1] ;
 wire \Tile_X4Y5_E2BEG[2] ;
 wire \Tile_X4Y5_E2BEG[3] ;
 wire \Tile_X4Y5_E2BEG[4] ;
 wire \Tile_X4Y5_E2BEG[5] ;
 wire \Tile_X4Y5_E2BEG[6] ;
 wire \Tile_X4Y5_E2BEG[7] ;
 wire \Tile_X4Y5_E2BEGb[0] ;
 wire \Tile_X4Y5_E2BEGb[1] ;
 wire \Tile_X4Y5_E2BEGb[2] ;
 wire \Tile_X4Y5_E2BEGb[3] ;
 wire \Tile_X4Y5_E2BEGb[4] ;
 wire \Tile_X4Y5_E2BEGb[5] ;
 wire \Tile_X4Y5_E2BEGb[6] ;
 wire \Tile_X4Y5_E2BEGb[7] ;
 wire \Tile_X4Y5_E6BEG[0] ;
 wire \Tile_X4Y5_E6BEG[10] ;
 wire \Tile_X4Y5_E6BEG[11] ;
 wire \Tile_X4Y5_E6BEG[1] ;
 wire \Tile_X4Y5_E6BEG[2] ;
 wire \Tile_X4Y5_E6BEG[3] ;
 wire \Tile_X4Y5_E6BEG[4] ;
 wire \Tile_X4Y5_E6BEG[5] ;
 wire \Tile_X4Y5_E6BEG[6] ;
 wire \Tile_X4Y5_E6BEG[7] ;
 wire \Tile_X4Y5_E6BEG[8] ;
 wire \Tile_X4Y5_E6BEG[9] ;
 wire \Tile_X4Y5_EE4BEG[0] ;
 wire \Tile_X4Y5_EE4BEG[10] ;
 wire \Tile_X4Y5_EE4BEG[11] ;
 wire \Tile_X4Y5_EE4BEG[12] ;
 wire \Tile_X4Y5_EE4BEG[13] ;
 wire \Tile_X4Y5_EE4BEG[14] ;
 wire \Tile_X4Y5_EE4BEG[15] ;
 wire \Tile_X4Y5_EE4BEG[1] ;
 wire \Tile_X4Y5_EE4BEG[2] ;
 wire \Tile_X4Y5_EE4BEG[3] ;
 wire \Tile_X4Y5_EE4BEG[4] ;
 wire \Tile_X4Y5_EE4BEG[5] ;
 wire \Tile_X4Y5_EE4BEG[6] ;
 wire \Tile_X4Y5_EE4BEG[7] ;
 wire \Tile_X4Y5_EE4BEG[8] ;
 wire \Tile_X4Y5_EE4BEG[9] ;
 wire \Tile_X4Y5_FrameData_O[0] ;
 wire \Tile_X4Y5_FrameData_O[10] ;
 wire \Tile_X4Y5_FrameData_O[11] ;
 wire \Tile_X4Y5_FrameData_O[12] ;
 wire \Tile_X4Y5_FrameData_O[13] ;
 wire \Tile_X4Y5_FrameData_O[14] ;
 wire \Tile_X4Y5_FrameData_O[15] ;
 wire \Tile_X4Y5_FrameData_O[16] ;
 wire \Tile_X4Y5_FrameData_O[17] ;
 wire \Tile_X4Y5_FrameData_O[18] ;
 wire \Tile_X4Y5_FrameData_O[19] ;
 wire \Tile_X4Y5_FrameData_O[1] ;
 wire \Tile_X4Y5_FrameData_O[20] ;
 wire \Tile_X4Y5_FrameData_O[21] ;
 wire \Tile_X4Y5_FrameData_O[22] ;
 wire \Tile_X4Y5_FrameData_O[23] ;
 wire \Tile_X4Y5_FrameData_O[24] ;
 wire \Tile_X4Y5_FrameData_O[25] ;
 wire \Tile_X4Y5_FrameData_O[26] ;
 wire \Tile_X4Y5_FrameData_O[27] ;
 wire \Tile_X4Y5_FrameData_O[28] ;
 wire \Tile_X4Y5_FrameData_O[29] ;
 wire \Tile_X4Y5_FrameData_O[2] ;
 wire \Tile_X4Y5_FrameData_O[30] ;
 wire \Tile_X4Y5_FrameData_O[31] ;
 wire \Tile_X4Y5_FrameData_O[3] ;
 wire \Tile_X4Y5_FrameData_O[4] ;
 wire \Tile_X4Y5_FrameData_O[5] ;
 wire \Tile_X4Y5_FrameData_O[6] ;
 wire \Tile_X4Y5_FrameData_O[7] ;
 wire \Tile_X4Y5_FrameData_O[8] ;
 wire \Tile_X4Y5_FrameData_O[9] ;
 wire \Tile_X4Y5_FrameStrobe_O[0] ;
 wire \Tile_X4Y5_FrameStrobe_O[10] ;
 wire \Tile_X4Y5_FrameStrobe_O[11] ;
 wire \Tile_X4Y5_FrameStrobe_O[12] ;
 wire \Tile_X4Y5_FrameStrobe_O[13] ;
 wire \Tile_X4Y5_FrameStrobe_O[14] ;
 wire \Tile_X4Y5_FrameStrobe_O[15] ;
 wire \Tile_X4Y5_FrameStrobe_O[16] ;
 wire \Tile_X4Y5_FrameStrobe_O[17] ;
 wire \Tile_X4Y5_FrameStrobe_O[18] ;
 wire \Tile_X4Y5_FrameStrobe_O[19] ;
 wire \Tile_X4Y5_FrameStrobe_O[1] ;
 wire \Tile_X4Y5_FrameStrobe_O[2] ;
 wire \Tile_X4Y5_FrameStrobe_O[3] ;
 wire \Tile_X4Y5_FrameStrobe_O[4] ;
 wire \Tile_X4Y5_FrameStrobe_O[5] ;
 wire \Tile_X4Y5_FrameStrobe_O[6] ;
 wire \Tile_X4Y5_FrameStrobe_O[7] ;
 wire \Tile_X4Y5_FrameStrobe_O[8] ;
 wire \Tile_X4Y5_FrameStrobe_O[9] ;
 wire \Tile_X4Y5_N1BEG[0] ;
 wire \Tile_X4Y5_N1BEG[1] ;
 wire \Tile_X4Y5_N1BEG[2] ;
 wire \Tile_X4Y5_N1BEG[3] ;
 wire \Tile_X4Y5_N2BEG[0] ;
 wire \Tile_X4Y5_N2BEG[1] ;
 wire \Tile_X4Y5_N2BEG[2] ;
 wire \Tile_X4Y5_N2BEG[3] ;
 wire \Tile_X4Y5_N2BEG[4] ;
 wire \Tile_X4Y5_N2BEG[5] ;
 wire \Tile_X4Y5_N2BEG[6] ;
 wire \Tile_X4Y5_N2BEG[7] ;
 wire \Tile_X4Y5_N2BEGb[0] ;
 wire \Tile_X4Y5_N2BEGb[1] ;
 wire \Tile_X4Y5_N2BEGb[2] ;
 wire \Tile_X4Y5_N2BEGb[3] ;
 wire \Tile_X4Y5_N2BEGb[4] ;
 wire \Tile_X4Y5_N2BEGb[5] ;
 wire \Tile_X4Y5_N2BEGb[6] ;
 wire \Tile_X4Y5_N2BEGb[7] ;
 wire \Tile_X4Y5_N4BEG[0] ;
 wire \Tile_X4Y5_N4BEG[10] ;
 wire \Tile_X4Y5_N4BEG[11] ;
 wire \Tile_X4Y5_N4BEG[12] ;
 wire \Tile_X4Y5_N4BEG[13] ;
 wire \Tile_X4Y5_N4BEG[14] ;
 wire \Tile_X4Y5_N4BEG[15] ;
 wire \Tile_X4Y5_N4BEG[1] ;
 wire \Tile_X4Y5_N4BEG[2] ;
 wire \Tile_X4Y5_N4BEG[3] ;
 wire \Tile_X4Y5_N4BEG[4] ;
 wire \Tile_X4Y5_N4BEG[5] ;
 wire \Tile_X4Y5_N4BEG[6] ;
 wire \Tile_X4Y5_N4BEG[7] ;
 wire \Tile_X4Y5_N4BEG[8] ;
 wire \Tile_X4Y5_N4BEG[9] ;
 wire \Tile_X4Y5_NN4BEG[0] ;
 wire \Tile_X4Y5_NN4BEG[10] ;
 wire \Tile_X4Y5_NN4BEG[11] ;
 wire \Tile_X4Y5_NN4BEG[12] ;
 wire \Tile_X4Y5_NN4BEG[13] ;
 wire \Tile_X4Y5_NN4BEG[14] ;
 wire \Tile_X4Y5_NN4BEG[15] ;
 wire \Tile_X4Y5_NN4BEG[1] ;
 wire \Tile_X4Y5_NN4BEG[2] ;
 wire \Tile_X4Y5_NN4BEG[3] ;
 wire \Tile_X4Y5_NN4BEG[4] ;
 wire \Tile_X4Y5_NN4BEG[5] ;
 wire \Tile_X4Y5_NN4BEG[6] ;
 wire \Tile_X4Y5_NN4BEG[7] ;
 wire \Tile_X4Y5_NN4BEG[8] ;
 wire \Tile_X4Y5_NN4BEG[9] ;
 wire \Tile_X4Y5_S1BEG[0] ;
 wire \Tile_X4Y5_S1BEG[1] ;
 wire \Tile_X4Y5_S1BEG[2] ;
 wire \Tile_X4Y5_S1BEG[3] ;
 wire \Tile_X4Y5_S2BEG[0] ;
 wire \Tile_X4Y5_S2BEG[1] ;
 wire \Tile_X4Y5_S2BEG[2] ;
 wire \Tile_X4Y5_S2BEG[3] ;
 wire \Tile_X4Y5_S2BEG[4] ;
 wire \Tile_X4Y5_S2BEG[5] ;
 wire \Tile_X4Y5_S2BEG[6] ;
 wire \Tile_X4Y5_S2BEG[7] ;
 wire \Tile_X4Y5_S2BEGb[0] ;
 wire \Tile_X4Y5_S2BEGb[1] ;
 wire \Tile_X4Y5_S2BEGb[2] ;
 wire \Tile_X4Y5_S2BEGb[3] ;
 wire \Tile_X4Y5_S2BEGb[4] ;
 wire \Tile_X4Y5_S2BEGb[5] ;
 wire \Tile_X4Y5_S2BEGb[6] ;
 wire \Tile_X4Y5_S2BEGb[7] ;
 wire \Tile_X4Y5_S4BEG[0] ;
 wire \Tile_X4Y5_S4BEG[10] ;
 wire \Tile_X4Y5_S4BEG[11] ;
 wire \Tile_X4Y5_S4BEG[12] ;
 wire \Tile_X4Y5_S4BEG[13] ;
 wire \Tile_X4Y5_S4BEG[14] ;
 wire \Tile_X4Y5_S4BEG[15] ;
 wire \Tile_X4Y5_S4BEG[1] ;
 wire \Tile_X4Y5_S4BEG[2] ;
 wire \Tile_X4Y5_S4BEG[3] ;
 wire \Tile_X4Y5_S4BEG[4] ;
 wire \Tile_X4Y5_S4BEG[5] ;
 wire \Tile_X4Y5_S4BEG[6] ;
 wire \Tile_X4Y5_S4BEG[7] ;
 wire \Tile_X4Y5_S4BEG[8] ;
 wire \Tile_X4Y5_S4BEG[9] ;
 wire \Tile_X4Y5_SS4BEG[0] ;
 wire \Tile_X4Y5_SS4BEG[10] ;
 wire \Tile_X4Y5_SS4BEG[11] ;
 wire \Tile_X4Y5_SS4BEG[12] ;
 wire \Tile_X4Y5_SS4BEG[13] ;
 wire \Tile_X4Y5_SS4BEG[14] ;
 wire \Tile_X4Y5_SS4BEG[15] ;
 wire \Tile_X4Y5_SS4BEG[1] ;
 wire \Tile_X4Y5_SS4BEG[2] ;
 wire \Tile_X4Y5_SS4BEG[3] ;
 wire \Tile_X4Y5_SS4BEG[4] ;
 wire \Tile_X4Y5_SS4BEG[5] ;
 wire \Tile_X4Y5_SS4BEG[6] ;
 wire \Tile_X4Y5_SS4BEG[7] ;
 wire \Tile_X4Y5_SS4BEG[8] ;
 wire \Tile_X4Y5_SS4BEG[9] ;
 wire Tile_X4Y5_UserCLKo;
 wire \Tile_X4Y5_W1BEG[0] ;
 wire \Tile_X4Y5_W1BEG[1] ;
 wire \Tile_X4Y5_W1BEG[2] ;
 wire \Tile_X4Y5_W1BEG[3] ;
 wire \Tile_X4Y5_W2BEG[0] ;
 wire \Tile_X4Y5_W2BEG[1] ;
 wire \Tile_X4Y5_W2BEG[2] ;
 wire \Tile_X4Y5_W2BEG[3] ;
 wire \Tile_X4Y5_W2BEG[4] ;
 wire \Tile_X4Y5_W2BEG[5] ;
 wire \Tile_X4Y5_W2BEG[6] ;
 wire \Tile_X4Y5_W2BEG[7] ;
 wire \Tile_X4Y5_W2BEGb[0] ;
 wire \Tile_X4Y5_W2BEGb[1] ;
 wire \Tile_X4Y5_W2BEGb[2] ;
 wire \Tile_X4Y5_W2BEGb[3] ;
 wire \Tile_X4Y5_W2BEGb[4] ;
 wire \Tile_X4Y5_W2BEGb[5] ;
 wire \Tile_X4Y5_W2BEGb[6] ;
 wire \Tile_X4Y5_W2BEGb[7] ;
 wire \Tile_X4Y5_W6BEG[0] ;
 wire \Tile_X4Y5_W6BEG[10] ;
 wire \Tile_X4Y5_W6BEG[11] ;
 wire \Tile_X4Y5_W6BEG[1] ;
 wire \Tile_X4Y5_W6BEG[2] ;
 wire \Tile_X4Y5_W6BEG[3] ;
 wire \Tile_X4Y5_W6BEG[4] ;
 wire \Tile_X4Y5_W6BEG[5] ;
 wire \Tile_X4Y5_W6BEG[6] ;
 wire \Tile_X4Y5_W6BEG[7] ;
 wire \Tile_X4Y5_W6BEG[8] ;
 wire \Tile_X4Y5_W6BEG[9] ;
 wire \Tile_X4Y5_WW4BEG[0] ;
 wire \Tile_X4Y5_WW4BEG[10] ;
 wire \Tile_X4Y5_WW4BEG[11] ;
 wire \Tile_X4Y5_WW4BEG[12] ;
 wire \Tile_X4Y5_WW4BEG[13] ;
 wire \Tile_X4Y5_WW4BEG[14] ;
 wire \Tile_X4Y5_WW4BEG[15] ;
 wire \Tile_X4Y5_WW4BEG[1] ;
 wire \Tile_X4Y5_WW4BEG[2] ;
 wire \Tile_X4Y5_WW4BEG[3] ;
 wire \Tile_X4Y5_WW4BEG[4] ;
 wire \Tile_X4Y5_WW4BEG[5] ;
 wire \Tile_X4Y5_WW4BEG[6] ;
 wire \Tile_X4Y5_WW4BEG[7] ;
 wire \Tile_X4Y5_WW4BEG[8] ;
 wire \Tile_X4Y5_WW4BEG[9] ;
 wire \Tile_X4Y6_E1BEG[0] ;
 wire \Tile_X4Y6_E1BEG[1] ;
 wire \Tile_X4Y6_E1BEG[2] ;
 wire \Tile_X4Y6_E1BEG[3] ;
 wire \Tile_X4Y6_E2BEG[0] ;
 wire \Tile_X4Y6_E2BEG[1] ;
 wire \Tile_X4Y6_E2BEG[2] ;
 wire \Tile_X4Y6_E2BEG[3] ;
 wire \Tile_X4Y6_E2BEG[4] ;
 wire \Tile_X4Y6_E2BEG[5] ;
 wire \Tile_X4Y6_E2BEG[6] ;
 wire \Tile_X4Y6_E2BEG[7] ;
 wire \Tile_X4Y6_E2BEGb[0] ;
 wire \Tile_X4Y6_E2BEGb[1] ;
 wire \Tile_X4Y6_E2BEGb[2] ;
 wire \Tile_X4Y6_E2BEGb[3] ;
 wire \Tile_X4Y6_E2BEGb[4] ;
 wire \Tile_X4Y6_E2BEGb[5] ;
 wire \Tile_X4Y6_E2BEGb[6] ;
 wire \Tile_X4Y6_E2BEGb[7] ;
 wire \Tile_X4Y6_E6BEG[0] ;
 wire \Tile_X4Y6_E6BEG[10] ;
 wire \Tile_X4Y6_E6BEG[11] ;
 wire \Tile_X4Y6_E6BEG[1] ;
 wire \Tile_X4Y6_E6BEG[2] ;
 wire \Tile_X4Y6_E6BEG[3] ;
 wire \Tile_X4Y6_E6BEG[4] ;
 wire \Tile_X4Y6_E6BEG[5] ;
 wire \Tile_X4Y6_E6BEG[6] ;
 wire \Tile_X4Y6_E6BEG[7] ;
 wire \Tile_X4Y6_E6BEG[8] ;
 wire \Tile_X4Y6_E6BEG[9] ;
 wire \Tile_X4Y6_EE4BEG[0] ;
 wire \Tile_X4Y6_EE4BEG[10] ;
 wire \Tile_X4Y6_EE4BEG[11] ;
 wire \Tile_X4Y6_EE4BEG[12] ;
 wire \Tile_X4Y6_EE4BEG[13] ;
 wire \Tile_X4Y6_EE4BEG[14] ;
 wire \Tile_X4Y6_EE4BEG[15] ;
 wire \Tile_X4Y6_EE4BEG[1] ;
 wire \Tile_X4Y6_EE4BEG[2] ;
 wire \Tile_X4Y6_EE4BEG[3] ;
 wire \Tile_X4Y6_EE4BEG[4] ;
 wire \Tile_X4Y6_EE4BEG[5] ;
 wire \Tile_X4Y6_EE4BEG[6] ;
 wire \Tile_X4Y6_EE4BEG[7] ;
 wire \Tile_X4Y6_EE4BEG[8] ;
 wire \Tile_X4Y6_EE4BEG[9] ;
 wire \Tile_X4Y6_FrameData_O[0] ;
 wire \Tile_X4Y6_FrameData_O[10] ;
 wire \Tile_X4Y6_FrameData_O[11] ;
 wire \Tile_X4Y6_FrameData_O[12] ;
 wire \Tile_X4Y6_FrameData_O[13] ;
 wire \Tile_X4Y6_FrameData_O[14] ;
 wire \Tile_X4Y6_FrameData_O[15] ;
 wire \Tile_X4Y6_FrameData_O[16] ;
 wire \Tile_X4Y6_FrameData_O[17] ;
 wire \Tile_X4Y6_FrameData_O[18] ;
 wire \Tile_X4Y6_FrameData_O[19] ;
 wire \Tile_X4Y6_FrameData_O[1] ;
 wire \Tile_X4Y6_FrameData_O[20] ;
 wire \Tile_X4Y6_FrameData_O[21] ;
 wire \Tile_X4Y6_FrameData_O[22] ;
 wire \Tile_X4Y6_FrameData_O[23] ;
 wire \Tile_X4Y6_FrameData_O[24] ;
 wire \Tile_X4Y6_FrameData_O[25] ;
 wire \Tile_X4Y6_FrameData_O[26] ;
 wire \Tile_X4Y6_FrameData_O[27] ;
 wire \Tile_X4Y6_FrameData_O[28] ;
 wire \Tile_X4Y6_FrameData_O[29] ;
 wire \Tile_X4Y6_FrameData_O[2] ;
 wire \Tile_X4Y6_FrameData_O[30] ;
 wire \Tile_X4Y6_FrameData_O[31] ;
 wire \Tile_X4Y6_FrameData_O[3] ;
 wire \Tile_X4Y6_FrameData_O[4] ;
 wire \Tile_X4Y6_FrameData_O[5] ;
 wire \Tile_X4Y6_FrameData_O[6] ;
 wire \Tile_X4Y6_FrameData_O[7] ;
 wire \Tile_X4Y6_FrameData_O[8] ;
 wire \Tile_X4Y6_FrameData_O[9] ;
 wire \Tile_X4Y6_FrameStrobe_O[0] ;
 wire \Tile_X4Y6_FrameStrobe_O[10] ;
 wire \Tile_X4Y6_FrameStrobe_O[11] ;
 wire \Tile_X4Y6_FrameStrobe_O[12] ;
 wire \Tile_X4Y6_FrameStrobe_O[13] ;
 wire \Tile_X4Y6_FrameStrobe_O[14] ;
 wire \Tile_X4Y6_FrameStrobe_O[15] ;
 wire \Tile_X4Y6_FrameStrobe_O[16] ;
 wire \Tile_X4Y6_FrameStrobe_O[17] ;
 wire \Tile_X4Y6_FrameStrobe_O[18] ;
 wire \Tile_X4Y6_FrameStrobe_O[19] ;
 wire \Tile_X4Y6_FrameStrobe_O[1] ;
 wire \Tile_X4Y6_FrameStrobe_O[2] ;
 wire \Tile_X4Y6_FrameStrobe_O[3] ;
 wire \Tile_X4Y6_FrameStrobe_O[4] ;
 wire \Tile_X4Y6_FrameStrobe_O[5] ;
 wire \Tile_X4Y6_FrameStrobe_O[6] ;
 wire \Tile_X4Y6_FrameStrobe_O[7] ;
 wire \Tile_X4Y6_FrameStrobe_O[8] ;
 wire \Tile_X4Y6_FrameStrobe_O[9] ;
 wire \Tile_X4Y6_N1BEG[0] ;
 wire \Tile_X4Y6_N1BEG[1] ;
 wire \Tile_X4Y6_N1BEG[2] ;
 wire \Tile_X4Y6_N1BEG[3] ;
 wire \Tile_X4Y6_N2BEG[0] ;
 wire \Tile_X4Y6_N2BEG[1] ;
 wire \Tile_X4Y6_N2BEG[2] ;
 wire \Tile_X4Y6_N2BEG[3] ;
 wire \Tile_X4Y6_N2BEG[4] ;
 wire \Tile_X4Y6_N2BEG[5] ;
 wire \Tile_X4Y6_N2BEG[6] ;
 wire \Tile_X4Y6_N2BEG[7] ;
 wire \Tile_X4Y6_N2BEGb[0] ;
 wire \Tile_X4Y6_N2BEGb[1] ;
 wire \Tile_X4Y6_N2BEGb[2] ;
 wire \Tile_X4Y6_N2BEGb[3] ;
 wire \Tile_X4Y6_N2BEGb[4] ;
 wire \Tile_X4Y6_N2BEGb[5] ;
 wire \Tile_X4Y6_N2BEGb[6] ;
 wire \Tile_X4Y6_N2BEGb[7] ;
 wire \Tile_X4Y6_N4BEG[0] ;
 wire \Tile_X4Y6_N4BEG[10] ;
 wire \Tile_X4Y6_N4BEG[11] ;
 wire \Tile_X4Y6_N4BEG[12] ;
 wire \Tile_X4Y6_N4BEG[13] ;
 wire \Tile_X4Y6_N4BEG[14] ;
 wire \Tile_X4Y6_N4BEG[15] ;
 wire \Tile_X4Y6_N4BEG[1] ;
 wire \Tile_X4Y6_N4BEG[2] ;
 wire \Tile_X4Y6_N4BEG[3] ;
 wire \Tile_X4Y6_N4BEG[4] ;
 wire \Tile_X4Y6_N4BEG[5] ;
 wire \Tile_X4Y6_N4BEG[6] ;
 wire \Tile_X4Y6_N4BEG[7] ;
 wire \Tile_X4Y6_N4BEG[8] ;
 wire \Tile_X4Y6_N4BEG[9] ;
 wire \Tile_X4Y6_NN4BEG[0] ;
 wire \Tile_X4Y6_NN4BEG[10] ;
 wire \Tile_X4Y6_NN4BEG[11] ;
 wire \Tile_X4Y6_NN4BEG[12] ;
 wire \Tile_X4Y6_NN4BEG[13] ;
 wire \Tile_X4Y6_NN4BEG[14] ;
 wire \Tile_X4Y6_NN4BEG[15] ;
 wire \Tile_X4Y6_NN4BEG[1] ;
 wire \Tile_X4Y6_NN4BEG[2] ;
 wire \Tile_X4Y6_NN4BEG[3] ;
 wire \Tile_X4Y6_NN4BEG[4] ;
 wire \Tile_X4Y6_NN4BEG[5] ;
 wire \Tile_X4Y6_NN4BEG[6] ;
 wire \Tile_X4Y6_NN4BEG[7] ;
 wire \Tile_X4Y6_NN4BEG[8] ;
 wire \Tile_X4Y6_NN4BEG[9] ;
 wire \Tile_X4Y6_S1BEG[0] ;
 wire \Tile_X4Y6_S1BEG[1] ;
 wire \Tile_X4Y6_S1BEG[2] ;
 wire \Tile_X4Y6_S1BEG[3] ;
 wire \Tile_X4Y6_S2BEG[0] ;
 wire \Tile_X4Y6_S2BEG[1] ;
 wire \Tile_X4Y6_S2BEG[2] ;
 wire \Tile_X4Y6_S2BEG[3] ;
 wire \Tile_X4Y6_S2BEG[4] ;
 wire \Tile_X4Y6_S2BEG[5] ;
 wire \Tile_X4Y6_S2BEG[6] ;
 wire \Tile_X4Y6_S2BEG[7] ;
 wire \Tile_X4Y6_S2BEGb[0] ;
 wire \Tile_X4Y6_S2BEGb[1] ;
 wire \Tile_X4Y6_S2BEGb[2] ;
 wire \Tile_X4Y6_S2BEGb[3] ;
 wire \Tile_X4Y6_S2BEGb[4] ;
 wire \Tile_X4Y6_S2BEGb[5] ;
 wire \Tile_X4Y6_S2BEGb[6] ;
 wire \Tile_X4Y6_S2BEGb[7] ;
 wire \Tile_X4Y6_S4BEG[0] ;
 wire \Tile_X4Y6_S4BEG[10] ;
 wire \Tile_X4Y6_S4BEG[11] ;
 wire \Tile_X4Y6_S4BEG[12] ;
 wire \Tile_X4Y6_S4BEG[13] ;
 wire \Tile_X4Y6_S4BEG[14] ;
 wire \Tile_X4Y6_S4BEG[15] ;
 wire \Tile_X4Y6_S4BEG[1] ;
 wire \Tile_X4Y6_S4BEG[2] ;
 wire \Tile_X4Y6_S4BEG[3] ;
 wire \Tile_X4Y6_S4BEG[4] ;
 wire \Tile_X4Y6_S4BEG[5] ;
 wire \Tile_X4Y6_S4BEG[6] ;
 wire \Tile_X4Y6_S4BEG[7] ;
 wire \Tile_X4Y6_S4BEG[8] ;
 wire \Tile_X4Y6_S4BEG[9] ;
 wire \Tile_X4Y6_SS4BEG[0] ;
 wire \Tile_X4Y6_SS4BEG[10] ;
 wire \Tile_X4Y6_SS4BEG[11] ;
 wire \Tile_X4Y6_SS4BEG[12] ;
 wire \Tile_X4Y6_SS4BEG[13] ;
 wire \Tile_X4Y6_SS4BEG[14] ;
 wire \Tile_X4Y6_SS4BEG[15] ;
 wire \Tile_X4Y6_SS4BEG[1] ;
 wire \Tile_X4Y6_SS4BEG[2] ;
 wire \Tile_X4Y6_SS4BEG[3] ;
 wire \Tile_X4Y6_SS4BEG[4] ;
 wire \Tile_X4Y6_SS4BEG[5] ;
 wire \Tile_X4Y6_SS4BEG[6] ;
 wire \Tile_X4Y6_SS4BEG[7] ;
 wire \Tile_X4Y6_SS4BEG[8] ;
 wire \Tile_X4Y6_SS4BEG[9] ;
 wire Tile_X4Y6_UserCLKo;
 wire \Tile_X4Y6_W1BEG[0] ;
 wire \Tile_X4Y6_W1BEG[1] ;
 wire \Tile_X4Y6_W1BEG[2] ;
 wire \Tile_X4Y6_W1BEG[3] ;
 wire \Tile_X4Y6_W2BEG[0] ;
 wire \Tile_X4Y6_W2BEG[1] ;
 wire \Tile_X4Y6_W2BEG[2] ;
 wire \Tile_X4Y6_W2BEG[3] ;
 wire \Tile_X4Y6_W2BEG[4] ;
 wire \Tile_X4Y6_W2BEG[5] ;
 wire \Tile_X4Y6_W2BEG[6] ;
 wire \Tile_X4Y6_W2BEG[7] ;
 wire \Tile_X4Y6_W2BEGb[0] ;
 wire \Tile_X4Y6_W2BEGb[1] ;
 wire \Tile_X4Y6_W2BEGb[2] ;
 wire \Tile_X4Y6_W2BEGb[3] ;
 wire \Tile_X4Y6_W2BEGb[4] ;
 wire \Tile_X4Y6_W2BEGb[5] ;
 wire \Tile_X4Y6_W2BEGb[6] ;
 wire \Tile_X4Y6_W2BEGb[7] ;
 wire \Tile_X4Y6_W6BEG[0] ;
 wire \Tile_X4Y6_W6BEG[10] ;
 wire \Tile_X4Y6_W6BEG[11] ;
 wire \Tile_X4Y6_W6BEG[1] ;
 wire \Tile_X4Y6_W6BEG[2] ;
 wire \Tile_X4Y6_W6BEG[3] ;
 wire \Tile_X4Y6_W6BEG[4] ;
 wire \Tile_X4Y6_W6BEG[5] ;
 wire \Tile_X4Y6_W6BEG[6] ;
 wire \Tile_X4Y6_W6BEG[7] ;
 wire \Tile_X4Y6_W6BEG[8] ;
 wire \Tile_X4Y6_W6BEG[9] ;
 wire \Tile_X4Y6_WW4BEG[0] ;
 wire \Tile_X4Y6_WW4BEG[10] ;
 wire \Tile_X4Y6_WW4BEG[11] ;
 wire \Tile_X4Y6_WW4BEG[12] ;
 wire \Tile_X4Y6_WW4BEG[13] ;
 wire \Tile_X4Y6_WW4BEG[14] ;
 wire \Tile_X4Y6_WW4BEG[15] ;
 wire \Tile_X4Y6_WW4BEG[1] ;
 wire \Tile_X4Y6_WW4BEG[2] ;
 wire \Tile_X4Y6_WW4BEG[3] ;
 wire \Tile_X4Y6_WW4BEG[4] ;
 wire \Tile_X4Y6_WW4BEG[5] ;
 wire \Tile_X4Y6_WW4BEG[6] ;
 wire \Tile_X4Y6_WW4BEG[7] ;
 wire \Tile_X4Y6_WW4BEG[8] ;
 wire \Tile_X4Y6_WW4BEG[9] ;
 wire \Tile_X4Y7_E1BEG[0] ;
 wire \Tile_X4Y7_E1BEG[1] ;
 wire \Tile_X4Y7_E1BEG[2] ;
 wire \Tile_X4Y7_E1BEG[3] ;
 wire \Tile_X4Y7_E2BEG[0] ;
 wire \Tile_X4Y7_E2BEG[1] ;
 wire \Tile_X4Y7_E2BEG[2] ;
 wire \Tile_X4Y7_E2BEG[3] ;
 wire \Tile_X4Y7_E2BEG[4] ;
 wire \Tile_X4Y7_E2BEG[5] ;
 wire \Tile_X4Y7_E2BEG[6] ;
 wire \Tile_X4Y7_E2BEG[7] ;
 wire \Tile_X4Y7_E2BEGb[0] ;
 wire \Tile_X4Y7_E2BEGb[1] ;
 wire \Tile_X4Y7_E2BEGb[2] ;
 wire \Tile_X4Y7_E2BEGb[3] ;
 wire \Tile_X4Y7_E2BEGb[4] ;
 wire \Tile_X4Y7_E2BEGb[5] ;
 wire \Tile_X4Y7_E2BEGb[6] ;
 wire \Tile_X4Y7_E2BEGb[7] ;
 wire \Tile_X4Y7_E6BEG[0] ;
 wire \Tile_X4Y7_E6BEG[10] ;
 wire \Tile_X4Y7_E6BEG[11] ;
 wire \Tile_X4Y7_E6BEG[1] ;
 wire \Tile_X4Y7_E6BEG[2] ;
 wire \Tile_X4Y7_E6BEG[3] ;
 wire \Tile_X4Y7_E6BEG[4] ;
 wire \Tile_X4Y7_E6BEG[5] ;
 wire \Tile_X4Y7_E6BEG[6] ;
 wire \Tile_X4Y7_E6BEG[7] ;
 wire \Tile_X4Y7_E6BEG[8] ;
 wire \Tile_X4Y7_E6BEG[9] ;
 wire \Tile_X4Y7_EE4BEG[0] ;
 wire \Tile_X4Y7_EE4BEG[10] ;
 wire \Tile_X4Y7_EE4BEG[11] ;
 wire \Tile_X4Y7_EE4BEG[12] ;
 wire \Tile_X4Y7_EE4BEG[13] ;
 wire \Tile_X4Y7_EE4BEG[14] ;
 wire \Tile_X4Y7_EE4BEG[15] ;
 wire \Tile_X4Y7_EE4BEG[1] ;
 wire \Tile_X4Y7_EE4BEG[2] ;
 wire \Tile_X4Y7_EE4BEG[3] ;
 wire \Tile_X4Y7_EE4BEG[4] ;
 wire \Tile_X4Y7_EE4BEG[5] ;
 wire \Tile_X4Y7_EE4BEG[6] ;
 wire \Tile_X4Y7_EE4BEG[7] ;
 wire \Tile_X4Y7_EE4BEG[8] ;
 wire \Tile_X4Y7_EE4BEG[9] ;
 wire \Tile_X4Y7_FrameData_O[0] ;
 wire \Tile_X4Y7_FrameData_O[10] ;
 wire \Tile_X4Y7_FrameData_O[11] ;
 wire \Tile_X4Y7_FrameData_O[12] ;
 wire \Tile_X4Y7_FrameData_O[13] ;
 wire \Tile_X4Y7_FrameData_O[14] ;
 wire \Tile_X4Y7_FrameData_O[15] ;
 wire \Tile_X4Y7_FrameData_O[16] ;
 wire \Tile_X4Y7_FrameData_O[17] ;
 wire \Tile_X4Y7_FrameData_O[18] ;
 wire \Tile_X4Y7_FrameData_O[19] ;
 wire \Tile_X4Y7_FrameData_O[1] ;
 wire \Tile_X4Y7_FrameData_O[20] ;
 wire \Tile_X4Y7_FrameData_O[21] ;
 wire \Tile_X4Y7_FrameData_O[22] ;
 wire \Tile_X4Y7_FrameData_O[23] ;
 wire \Tile_X4Y7_FrameData_O[24] ;
 wire \Tile_X4Y7_FrameData_O[25] ;
 wire \Tile_X4Y7_FrameData_O[26] ;
 wire \Tile_X4Y7_FrameData_O[27] ;
 wire \Tile_X4Y7_FrameData_O[28] ;
 wire \Tile_X4Y7_FrameData_O[29] ;
 wire \Tile_X4Y7_FrameData_O[2] ;
 wire \Tile_X4Y7_FrameData_O[30] ;
 wire \Tile_X4Y7_FrameData_O[31] ;
 wire \Tile_X4Y7_FrameData_O[3] ;
 wire \Tile_X4Y7_FrameData_O[4] ;
 wire \Tile_X4Y7_FrameData_O[5] ;
 wire \Tile_X4Y7_FrameData_O[6] ;
 wire \Tile_X4Y7_FrameData_O[7] ;
 wire \Tile_X4Y7_FrameData_O[8] ;
 wire \Tile_X4Y7_FrameData_O[9] ;
 wire \Tile_X4Y7_FrameStrobe_O[0] ;
 wire \Tile_X4Y7_FrameStrobe_O[10] ;
 wire \Tile_X4Y7_FrameStrobe_O[11] ;
 wire \Tile_X4Y7_FrameStrobe_O[12] ;
 wire \Tile_X4Y7_FrameStrobe_O[13] ;
 wire \Tile_X4Y7_FrameStrobe_O[14] ;
 wire \Tile_X4Y7_FrameStrobe_O[15] ;
 wire \Tile_X4Y7_FrameStrobe_O[16] ;
 wire \Tile_X4Y7_FrameStrobe_O[17] ;
 wire \Tile_X4Y7_FrameStrobe_O[18] ;
 wire \Tile_X4Y7_FrameStrobe_O[19] ;
 wire \Tile_X4Y7_FrameStrobe_O[1] ;
 wire \Tile_X4Y7_FrameStrobe_O[2] ;
 wire \Tile_X4Y7_FrameStrobe_O[3] ;
 wire \Tile_X4Y7_FrameStrobe_O[4] ;
 wire \Tile_X4Y7_FrameStrobe_O[5] ;
 wire \Tile_X4Y7_FrameStrobe_O[6] ;
 wire \Tile_X4Y7_FrameStrobe_O[7] ;
 wire \Tile_X4Y7_FrameStrobe_O[8] ;
 wire \Tile_X4Y7_FrameStrobe_O[9] ;
 wire \Tile_X4Y7_N1BEG[0] ;
 wire \Tile_X4Y7_N1BEG[1] ;
 wire \Tile_X4Y7_N1BEG[2] ;
 wire \Tile_X4Y7_N1BEG[3] ;
 wire \Tile_X4Y7_N2BEG[0] ;
 wire \Tile_X4Y7_N2BEG[1] ;
 wire \Tile_X4Y7_N2BEG[2] ;
 wire \Tile_X4Y7_N2BEG[3] ;
 wire \Tile_X4Y7_N2BEG[4] ;
 wire \Tile_X4Y7_N2BEG[5] ;
 wire \Tile_X4Y7_N2BEG[6] ;
 wire \Tile_X4Y7_N2BEG[7] ;
 wire \Tile_X4Y7_N2BEGb[0] ;
 wire \Tile_X4Y7_N2BEGb[1] ;
 wire \Tile_X4Y7_N2BEGb[2] ;
 wire \Tile_X4Y7_N2BEGb[3] ;
 wire \Tile_X4Y7_N2BEGb[4] ;
 wire \Tile_X4Y7_N2BEGb[5] ;
 wire \Tile_X4Y7_N2BEGb[6] ;
 wire \Tile_X4Y7_N2BEGb[7] ;
 wire \Tile_X4Y7_N4BEG[0] ;
 wire \Tile_X4Y7_N4BEG[10] ;
 wire \Tile_X4Y7_N4BEG[11] ;
 wire \Tile_X4Y7_N4BEG[12] ;
 wire \Tile_X4Y7_N4BEG[13] ;
 wire \Tile_X4Y7_N4BEG[14] ;
 wire \Tile_X4Y7_N4BEG[15] ;
 wire \Tile_X4Y7_N4BEG[1] ;
 wire \Tile_X4Y7_N4BEG[2] ;
 wire \Tile_X4Y7_N4BEG[3] ;
 wire \Tile_X4Y7_N4BEG[4] ;
 wire \Tile_X4Y7_N4BEG[5] ;
 wire \Tile_X4Y7_N4BEG[6] ;
 wire \Tile_X4Y7_N4BEG[7] ;
 wire \Tile_X4Y7_N4BEG[8] ;
 wire \Tile_X4Y7_N4BEG[9] ;
 wire \Tile_X4Y7_NN4BEG[0] ;
 wire \Tile_X4Y7_NN4BEG[10] ;
 wire \Tile_X4Y7_NN4BEG[11] ;
 wire \Tile_X4Y7_NN4BEG[12] ;
 wire \Tile_X4Y7_NN4BEG[13] ;
 wire \Tile_X4Y7_NN4BEG[14] ;
 wire \Tile_X4Y7_NN4BEG[15] ;
 wire \Tile_X4Y7_NN4BEG[1] ;
 wire \Tile_X4Y7_NN4BEG[2] ;
 wire \Tile_X4Y7_NN4BEG[3] ;
 wire \Tile_X4Y7_NN4BEG[4] ;
 wire \Tile_X4Y7_NN4BEG[5] ;
 wire \Tile_X4Y7_NN4BEG[6] ;
 wire \Tile_X4Y7_NN4BEG[7] ;
 wire \Tile_X4Y7_NN4BEG[8] ;
 wire \Tile_X4Y7_NN4BEG[9] ;
 wire \Tile_X4Y7_S1BEG[0] ;
 wire \Tile_X4Y7_S1BEG[1] ;
 wire \Tile_X4Y7_S1BEG[2] ;
 wire \Tile_X4Y7_S1BEG[3] ;
 wire \Tile_X4Y7_S2BEG[0] ;
 wire \Tile_X4Y7_S2BEG[1] ;
 wire \Tile_X4Y7_S2BEG[2] ;
 wire \Tile_X4Y7_S2BEG[3] ;
 wire \Tile_X4Y7_S2BEG[4] ;
 wire \Tile_X4Y7_S2BEG[5] ;
 wire \Tile_X4Y7_S2BEG[6] ;
 wire \Tile_X4Y7_S2BEG[7] ;
 wire \Tile_X4Y7_S2BEGb[0] ;
 wire \Tile_X4Y7_S2BEGb[1] ;
 wire \Tile_X4Y7_S2BEGb[2] ;
 wire \Tile_X4Y7_S2BEGb[3] ;
 wire \Tile_X4Y7_S2BEGb[4] ;
 wire \Tile_X4Y7_S2BEGb[5] ;
 wire \Tile_X4Y7_S2BEGb[6] ;
 wire \Tile_X4Y7_S2BEGb[7] ;
 wire \Tile_X4Y7_S4BEG[0] ;
 wire \Tile_X4Y7_S4BEG[10] ;
 wire \Tile_X4Y7_S4BEG[11] ;
 wire \Tile_X4Y7_S4BEG[12] ;
 wire \Tile_X4Y7_S4BEG[13] ;
 wire \Tile_X4Y7_S4BEG[14] ;
 wire \Tile_X4Y7_S4BEG[15] ;
 wire \Tile_X4Y7_S4BEG[1] ;
 wire \Tile_X4Y7_S4BEG[2] ;
 wire \Tile_X4Y7_S4BEG[3] ;
 wire \Tile_X4Y7_S4BEG[4] ;
 wire \Tile_X4Y7_S4BEG[5] ;
 wire \Tile_X4Y7_S4BEG[6] ;
 wire \Tile_X4Y7_S4BEG[7] ;
 wire \Tile_X4Y7_S4BEG[8] ;
 wire \Tile_X4Y7_S4BEG[9] ;
 wire \Tile_X4Y7_SS4BEG[0] ;
 wire \Tile_X4Y7_SS4BEG[10] ;
 wire \Tile_X4Y7_SS4BEG[11] ;
 wire \Tile_X4Y7_SS4BEG[12] ;
 wire \Tile_X4Y7_SS4BEG[13] ;
 wire \Tile_X4Y7_SS4BEG[14] ;
 wire \Tile_X4Y7_SS4BEG[15] ;
 wire \Tile_X4Y7_SS4BEG[1] ;
 wire \Tile_X4Y7_SS4BEG[2] ;
 wire \Tile_X4Y7_SS4BEG[3] ;
 wire \Tile_X4Y7_SS4BEG[4] ;
 wire \Tile_X4Y7_SS4BEG[5] ;
 wire \Tile_X4Y7_SS4BEG[6] ;
 wire \Tile_X4Y7_SS4BEG[7] ;
 wire \Tile_X4Y7_SS4BEG[8] ;
 wire \Tile_X4Y7_SS4BEG[9] ;
 wire Tile_X4Y7_UserCLKo;
 wire \Tile_X4Y7_W1BEG[0] ;
 wire \Tile_X4Y7_W1BEG[1] ;
 wire \Tile_X4Y7_W1BEG[2] ;
 wire \Tile_X4Y7_W1BEG[3] ;
 wire \Tile_X4Y7_W2BEG[0] ;
 wire \Tile_X4Y7_W2BEG[1] ;
 wire \Tile_X4Y7_W2BEG[2] ;
 wire \Tile_X4Y7_W2BEG[3] ;
 wire \Tile_X4Y7_W2BEG[4] ;
 wire \Tile_X4Y7_W2BEG[5] ;
 wire \Tile_X4Y7_W2BEG[6] ;
 wire \Tile_X4Y7_W2BEG[7] ;
 wire \Tile_X4Y7_W2BEGb[0] ;
 wire \Tile_X4Y7_W2BEGb[1] ;
 wire \Tile_X4Y7_W2BEGb[2] ;
 wire \Tile_X4Y7_W2BEGb[3] ;
 wire \Tile_X4Y7_W2BEGb[4] ;
 wire \Tile_X4Y7_W2BEGb[5] ;
 wire \Tile_X4Y7_W2BEGb[6] ;
 wire \Tile_X4Y7_W2BEGb[7] ;
 wire \Tile_X4Y7_W6BEG[0] ;
 wire \Tile_X4Y7_W6BEG[10] ;
 wire \Tile_X4Y7_W6BEG[11] ;
 wire \Tile_X4Y7_W6BEG[1] ;
 wire \Tile_X4Y7_W6BEG[2] ;
 wire \Tile_X4Y7_W6BEG[3] ;
 wire \Tile_X4Y7_W6BEG[4] ;
 wire \Tile_X4Y7_W6BEG[5] ;
 wire \Tile_X4Y7_W6BEG[6] ;
 wire \Tile_X4Y7_W6BEG[7] ;
 wire \Tile_X4Y7_W6BEG[8] ;
 wire \Tile_X4Y7_W6BEG[9] ;
 wire \Tile_X4Y7_WW4BEG[0] ;
 wire \Tile_X4Y7_WW4BEG[10] ;
 wire \Tile_X4Y7_WW4BEG[11] ;
 wire \Tile_X4Y7_WW4BEG[12] ;
 wire \Tile_X4Y7_WW4BEG[13] ;
 wire \Tile_X4Y7_WW4BEG[14] ;
 wire \Tile_X4Y7_WW4BEG[15] ;
 wire \Tile_X4Y7_WW4BEG[1] ;
 wire \Tile_X4Y7_WW4BEG[2] ;
 wire \Tile_X4Y7_WW4BEG[3] ;
 wire \Tile_X4Y7_WW4BEG[4] ;
 wire \Tile_X4Y7_WW4BEG[5] ;
 wire \Tile_X4Y7_WW4BEG[6] ;
 wire \Tile_X4Y7_WW4BEG[7] ;
 wire \Tile_X4Y7_WW4BEG[8] ;
 wire \Tile_X4Y7_WW4BEG[9] ;
 wire \Tile_X4Y8_E1BEG[0] ;
 wire \Tile_X4Y8_E1BEG[1] ;
 wire \Tile_X4Y8_E1BEG[2] ;
 wire \Tile_X4Y8_E1BEG[3] ;
 wire \Tile_X4Y8_E2BEG[0] ;
 wire \Tile_X4Y8_E2BEG[1] ;
 wire \Tile_X4Y8_E2BEG[2] ;
 wire \Tile_X4Y8_E2BEG[3] ;
 wire \Tile_X4Y8_E2BEG[4] ;
 wire \Tile_X4Y8_E2BEG[5] ;
 wire \Tile_X4Y8_E2BEG[6] ;
 wire \Tile_X4Y8_E2BEG[7] ;
 wire \Tile_X4Y8_E2BEGb[0] ;
 wire \Tile_X4Y8_E2BEGb[1] ;
 wire \Tile_X4Y8_E2BEGb[2] ;
 wire \Tile_X4Y8_E2BEGb[3] ;
 wire \Tile_X4Y8_E2BEGb[4] ;
 wire \Tile_X4Y8_E2BEGb[5] ;
 wire \Tile_X4Y8_E2BEGb[6] ;
 wire \Tile_X4Y8_E2BEGb[7] ;
 wire \Tile_X4Y8_E6BEG[0] ;
 wire \Tile_X4Y8_E6BEG[10] ;
 wire \Tile_X4Y8_E6BEG[11] ;
 wire \Tile_X4Y8_E6BEG[1] ;
 wire \Tile_X4Y8_E6BEG[2] ;
 wire \Tile_X4Y8_E6BEG[3] ;
 wire \Tile_X4Y8_E6BEG[4] ;
 wire \Tile_X4Y8_E6BEG[5] ;
 wire \Tile_X4Y8_E6BEG[6] ;
 wire \Tile_X4Y8_E6BEG[7] ;
 wire \Tile_X4Y8_E6BEG[8] ;
 wire \Tile_X4Y8_E6BEG[9] ;
 wire \Tile_X4Y8_EE4BEG[0] ;
 wire \Tile_X4Y8_EE4BEG[10] ;
 wire \Tile_X4Y8_EE4BEG[11] ;
 wire \Tile_X4Y8_EE4BEG[12] ;
 wire \Tile_X4Y8_EE4BEG[13] ;
 wire \Tile_X4Y8_EE4BEG[14] ;
 wire \Tile_X4Y8_EE4BEG[15] ;
 wire \Tile_X4Y8_EE4BEG[1] ;
 wire \Tile_X4Y8_EE4BEG[2] ;
 wire \Tile_X4Y8_EE4BEG[3] ;
 wire \Tile_X4Y8_EE4BEG[4] ;
 wire \Tile_X4Y8_EE4BEG[5] ;
 wire \Tile_X4Y8_EE4BEG[6] ;
 wire \Tile_X4Y8_EE4BEG[7] ;
 wire \Tile_X4Y8_EE4BEG[8] ;
 wire \Tile_X4Y8_EE4BEG[9] ;
 wire \Tile_X4Y8_FrameData_O[0] ;
 wire \Tile_X4Y8_FrameData_O[10] ;
 wire \Tile_X4Y8_FrameData_O[11] ;
 wire \Tile_X4Y8_FrameData_O[12] ;
 wire \Tile_X4Y8_FrameData_O[13] ;
 wire \Tile_X4Y8_FrameData_O[14] ;
 wire \Tile_X4Y8_FrameData_O[15] ;
 wire \Tile_X4Y8_FrameData_O[16] ;
 wire \Tile_X4Y8_FrameData_O[17] ;
 wire \Tile_X4Y8_FrameData_O[18] ;
 wire \Tile_X4Y8_FrameData_O[19] ;
 wire \Tile_X4Y8_FrameData_O[1] ;
 wire \Tile_X4Y8_FrameData_O[20] ;
 wire \Tile_X4Y8_FrameData_O[21] ;
 wire \Tile_X4Y8_FrameData_O[22] ;
 wire \Tile_X4Y8_FrameData_O[23] ;
 wire \Tile_X4Y8_FrameData_O[24] ;
 wire \Tile_X4Y8_FrameData_O[25] ;
 wire \Tile_X4Y8_FrameData_O[26] ;
 wire \Tile_X4Y8_FrameData_O[27] ;
 wire \Tile_X4Y8_FrameData_O[28] ;
 wire \Tile_X4Y8_FrameData_O[29] ;
 wire \Tile_X4Y8_FrameData_O[2] ;
 wire \Tile_X4Y8_FrameData_O[30] ;
 wire \Tile_X4Y8_FrameData_O[31] ;
 wire \Tile_X4Y8_FrameData_O[3] ;
 wire \Tile_X4Y8_FrameData_O[4] ;
 wire \Tile_X4Y8_FrameData_O[5] ;
 wire \Tile_X4Y8_FrameData_O[6] ;
 wire \Tile_X4Y8_FrameData_O[7] ;
 wire \Tile_X4Y8_FrameData_O[8] ;
 wire \Tile_X4Y8_FrameData_O[9] ;
 wire \Tile_X4Y8_FrameStrobe_O[0] ;
 wire \Tile_X4Y8_FrameStrobe_O[10] ;
 wire \Tile_X4Y8_FrameStrobe_O[11] ;
 wire \Tile_X4Y8_FrameStrobe_O[12] ;
 wire \Tile_X4Y8_FrameStrobe_O[13] ;
 wire \Tile_X4Y8_FrameStrobe_O[14] ;
 wire \Tile_X4Y8_FrameStrobe_O[15] ;
 wire \Tile_X4Y8_FrameStrobe_O[16] ;
 wire \Tile_X4Y8_FrameStrobe_O[17] ;
 wire \Tile_X4Y8_FrameStrobe_O[18] ;
 wire \Tile_X4Y8_FrameStrobe_O[19] ;
 wire \Tile_X4Y8_FrameStrobe_O[1] ;
 wire \Tile_X4Y8_FrameStrobe_O[2] ;
 wire \Tile_X4Y8_FrameStrobe_O[3] ;
 wire \Tile_X4Y8_FrameStrobe_O[4] ;
 wire \Tile_X4Y8_FrameStrobe_O[5] ;
 wire \Tile_X4Y8_FrameStrobe_O[6] ;
 wire \Tile_X4Y8_FrameStrobe_O[7] ;
 wire \Tile_X4Y8_FrameStrobe_O[8] ;
 wire \Tile_X4Y8_FrameStrobe_O[9] ;
 wire \Tile_X4Y8_N1BEG[0] ;
 wire \Tile_X4Y8_N1BEG[1] ;
 wire \Tile_X4Y8_N1BEG[2] ;
 wire \Tile_X4Y8_N1BEG[3] ;
 wire \Tile_X4Y8_N2BEG[0] ;
 wire \Tile_X4Y8_N2BEG[1] ;
 wire \Tile_X4Y8_N2BEG[2] ;
 wire \Tile_X4Y8_N2BEG[3] ;
 wire \Tile_X4Y8_N2BEG[4] ;
 wire \Tile_X4Y8_N2BEG[5] ;
 wire \Tile_X4Y8_N2BEG[6] ;
 wire \Tile_X4Y8_N2BEG[7] ;
 wire \Tile_X4Y8_N2BEGb[0] ;
 wire \Tile_X4Y8_N2BEGb[1] ;
 wire \Tile_X4Y8_N2BEGb[2] ;
 wire \Tile_X4Y8_N2BEGb[3] ;
 wire \Tile_X4Y8_N2BEGb[4] ;
 wire \Tile_X4Y8_N2BEGb[5] ;
 wire \Tile_X4Y8_N2BEGb[6] ;
 wire \Tile_X4Y8_N2BEGb[7] ;
 wire \Tile_X4Y8_N4BEG[0] ;
 wire \Tile_X4Y8_N4BEG[10] ;
 wire \Tile_X4Y8_N4BEG[11] ;
 wire \Tile_X4Y8_N4BEG[12] ;
 wire \Tile_X4Y8_N4BEG[13] ;
 wire \Tile_X4Y8_N4BEG[14] ;
 wire \Tile_X4Y8_N4BEG[15] ;
 wire \Tile_X4Y8_N4BEG[1] ;
 wire \Tile_X4Y8_N4BEG[2] ;
 wire \Tile_X4Y8_N4BEG[3] ;
 wire \Tile_X4Y8_N4BEG[4] ;
 wire \Tile_X4Y8_N4BEG[5] ;
 wire \Tile_X4Y8_N4BEG[6] ;
 wire \Tile_X4Y8_N4BEG[7] ;
 wire \Tile_X4Y8_N4BEG[8] ;
 wire \Tile_X4Y8_N4BEG[9] ;
 wire \Tile_X4Y8_NN4BEG[0] ;
 wire \Tile_X4Y8_NN4BEG[10] ;
 wire \Tile_X4Y8_NN4BEG[11] ;
 wire \Tile_X4Y8_NN4BEG[12] ;
 wire \Tile_X4Y8_NN4BEG[13] ;
 wire \Tile_X4Y8_NN4BEG[14] ;
 wire \Tile_X4Y8_NN4BEG[15] ;
 wire \Tile_X4Y8_NN4BEG[1] ;
 wire \Tile_X4Y8_NN4BEG[2] ;
 wire \Tile_X4Y8_NN4BEG[3] ;
 wire \Tile_X4Y8_NN4BEG[4] ;
 wire \Tile_X4Y8_NN4BEG[5] ;
 wire \Tile_X4Y8_NN4BEG[6] ;
 wire \Tile_X4Y8_NN4BEG[7] ;
 wire \Tile_X4Y8_NN4BEG[8] ;
 wire \Tile_X4Y8_NN4BEG[9] ;
 wire \Tile_X4Y8_S1BEG[0] ;
 wire \Tile_X4Y8_S1BEG[1] ;
 wire \Tile_X4Y8_S1BEG[2] ;
 wire \Tile_X4Y8_S1BEG[3] ;
 wire \Tile_X4Y8_S2BEG[0] ;
 wire \Tile_X4Y8_S2BEG[1] ;
 wire \Tile_X4Y8_S2BEG[2] ;
 wire \Tile_X4Y8_S2BEG[3] ;
 wire \Tile_X4Y8_S2BEG[4] ;
 wire \Tile_X4Y8_S2BEG[5] ;
 wire \Tile_X4Y8_S2BEG[6] ;
 wire \Tile_X4Y8_S2BEG[7] ;
 wire \Tile_X4Y8_S2BEGb[0] ;
 wire \Tile_X4Y8_S2BEGb[1] ;
 wire \Tile_X4Y8_S2BEGb[2] ;
 wire \Tile_X4Y8_S2BEGb[3] ;
 wire \Tile_X4Y8_S2BEGb[4] ;
 wire \Tile_X4Y8_S2BEGb[5] ;
 wire \Tile_X4Y8_S2BEGb[6] ;
 wire \Tile_X4Y8_S2BEGb[7] ;
 wire \Tile_X4Y8_S4BEG[0] ;
 wire \Tile_X4Y8_S4BEG[10] ;
 wire \Tile_X4Y8_S4BEG[11] ;
 wire \Tile_X4Y8_S4BEG[12] ;
 wire \Tile_X4Y8_S4BEG[13] ;
 wire \Tile_X4Y8_S4BEG[14] ;
 wire \Tile_X4Y8_S4BEG[15] ;
 wire \Tile_X4Y8_S4BEG[1] ;
 wire \Tile_X4Y8_S4BEG[2] ;
 wire \Tile_X4Y8_S4BEG[3] ;
 wire \Tile_X4Y8_S4BEG[4] ;
 wire \Tile_X4Y8_S4BEG[5] ;
 wire \Tile_X4Y8_S4BEG[6] ;
 wire \Tile_X4Y8_S4BEG[7] ;
 wire \Tile_X4Y8_S4BEG[8] ;
 wire \Tile_X4Y8_S4BEG[9] ;
 wire \Tile_X4Y8_SS4BEG[0] ;
 wire \Tile_X4Y8_SS4BEG[10] ;
 wire \Tile_X4Y8_SS4BEG[11] ;
 wire \Tile_X4Y8_SS4BEG[12] ;
 wire \Tile_X4Y8_SS4BEG[13] ;
 wire \Tile_X4Y8_SS4BEG[14] ;
 wire \Tile_X4Y8_SS4BEG[15] ;
 wire \Tile_X4Y8_SS4BEG[1] ;
 wire \Tile_X4Y8_SS4BEG[2] ;
 wire \Tile_X4Y8_SS4BEG[3] ;
 wire \Tile_X4Y8_SS4BEG[4] ;
 wire \Tile_X4Y8_SS4BEG[5] ;
 wire \Tile_X4Y8_SS4BEG[6] ;
 wire \Tile_X4Y8_SS4BEG[7] ;
 wire \Tile_X4Y8_SS4BEG[8] ;
 wire \Tile_X4Y8_SS4BEG[9] ;
 wire Tile_X4Y8_UserCLKo;
 wire \Tile_X4Y8_W1BEG[0] ;
 wire \Tile_X4Y8_W1BEG[1] ;
 wire \Tile_X4Y8_W1BEG[2] ;
 wire \Tile_X4Y8_W1BEG[3] ;
 wire \Tile_X4Y8_W2BEG[0] ;
 wire \Tile_X4Y8_W2BEG[1] ;
 wire \Tile_X4Y8_W2BEG[2] ;
 wire \Tile_X4Y8_W2BEG[3] ;
 wire \Tile_X4Y8_W2BEG[4] ;
 wire \Tile_X4Y8_W2BEG[5] ;
 wire \Tile_X4Y8_W2BEG[6] ;
 wire \Tile_X4Y8_W2BEG[7] ;
 wire \Tile_X4Y8_W2BEGb[0] ;
 wire \Tile_X4Y8_W2BEGb[1] ;
 wire \Tile_X4Y8_W2BEGb[2] ;
 wire \Tile_X4Y8_W2BEGb[3] ;
 wire \Tile_X4Y8_W2BEGb[4] ;
 wire \Tile_X4Y8_W2BEGb[5] ;
 wire \Tile_X4Y8_W2BEGb[6] ;
 wire \Tile_X4Y8_W2BEGb[7] ;
 wire \Tile_X4Y8_W6BEG[0] ;
 wire \Tile_X4Y8_W6BEG[10] ;
 wire \Tile_X4Y8_W6BEG[11] ;
 wire \Tile_X4Y8_W6BEG[1] ;
 wire \Tile_X4Y8_W6BEG[2] ;
 wire \Tile_X4Y8_W6BEG[3] ;
 wire \Tile_X4Y8_W6BEG[4] ;
 wire \Tile_X4Y8_W6BEG[5] ;
 wire \Tile_X4Y8_W6BEG[6] ;
 wire \Tile_X4Y8_W6BEG[7] ;
 wire \Tile_X4Y8_W6BEG[8] ;
 wire \Tile_X4Y8_W6BEG[9] ;
 wire \Tile_X4Y8_WW4BEG[0] ;
 wire \Tile_X4Y8_WW4BEG[10] ;
 wire \Tile_X4Y8_WW4BEG[11] ;
 wire \Tile_X4Y8_WW4BEG[12] ;
 wire \Tile_X4Y8_WW4BEG[13] ;
 wire \Tile_X4Y8_WW4BEG[14] ;
 wire \Tile_X4Y8_WW4BEG[15] ;
 wire \Tile_X4Y8_WW4BEG[1] ;
 wire \Tile_X4Y8_WW4BEG[2] ;
 wire \Tile_X4Y8_WW4BEG[3] ;
 wire \Tile_X4Y8_WW4BEG[4] ;
 wire \Tile_X4Y8_WW4BEG[5] ;
 wire \Tile_X4Y8_WW4BEG[6] ;
 wire \Tile_X4Y8_WW4BEG[7] ;
 wire \Tile_X4Y8_WW4BEG[8] ;
 wire \Tile_X4Y8_WW4BEG[9] ;
 wire \Tile_X4Y9_E1BEG[0] ;
 wire \Tile_X4Y9_E1BEG[1] ;
 wire \Tile_X4Y9_E1BEG[2] ;
 wire \Tile_X4Y9_E1BEG[3] ;
 wire \Tile_X4Y9_E2BEG[0] ;
 wire \Tile_X4Y9_E2BEG[1] ;
 wire \Tile_X4Y9_E2BEG[2] ;
 wire \Tile_X4Y9_E2BEG[3] ;
 wire \Tile_X4Y9_E2BEG[4] ;
 wire \Tile_X4Y9_E2BEG[5] ;
 wire \Tile_X4Y9_E2BEG[6] ;
 wire \Tile_X4Y9_E2BEG[7] ;
 wire \Tile_X4Y9_E2BEGb[0] ;
 wire \Tile_X4Y9_E2BEGb[1] ;
 wire \Tile_X4Y9_E2BEGb[2] ;
 wire \Tile_X4Y9_E2BEGb[3] ;
 wire \Tile_X4Y9_E2BEGb[4] ;
 wire \Tile_X4Y9_E2BEGb[5] ;
 wire \Tile_X4Y9_E2BEGb[6] ;
 wire \Tile_X4Y9_E2BEGb[7] ;
 wire \Tile_X4Y9_E6BEG[0] ;
 wire \Tile_X4Y9_E6BEG[10] ;
 wire \Tile_X4Y9_E6BEG[11] ;
 wire \Tile_X4Y9_E6BEG[1] ;
 wire \Tile_X4Y9_E6BEG[2] ;
 wire \Tile_X4Y9_E6BEG[3] ;
 wire \Tile_X4Y9_E6BEG[4] ;
 wire \Tile_X4Y9_E6BEG[5] ;
 wire \Tile_X4Y9_E6BEG[6] ;
 wire \Tile_X4Y9_E6BEG[7] ;
 wire \Tile_X4Y9_E6BEG[8] ;
 wire \Tile_X4Y9_E6BEG[9] ;
 wire \Tile_X4Y9_EE4BEG[0] ;
 wire \Tile_X4Y9_EE4BEG[10] ;
 wire \Tile_X4Y9_EE4BEG[11] ;
 wire \Tile_X4Y9_EE4BEG[12] ;
 wire \Tile_X4Y9_EE4BEG[13] ;
 wire \Tile_X4Y9_EE4BEG[14] ;
 wire \Tile_X4Y9_EE4BEG[15] ;
 wire \Tile_X4Y9_EE4BEG[1] ;
 wire \Tile_X4Y9_EE4BEG[2] ;
 wire \Tile_X4Y9_EE4BEG[3] ;
 wire \Tile_X4Y9_EE4BEG[4] ;
 wire \Tile_X4Y9_EE4BEG[5] ;
 wire \Tile_X4Y9_EE4BEG[6] ;
 wire \Tile_X4Y9_EE4BEG[7] ;
 wire \Tile_X4Y9_EE4BEG[8] ;
 wire \Tile_X4Y9_EE4BEG[9] ;
 wire \Tile_X4Y9_FrameData_O[0] ;
 wire \Tile_X4Y9_FrameData_O[10] ;
 wire \Tile_X4Y9_FrameData_O[11] ;
 wire \Tile_X4Y9_FrameData_O[12] ;
 wire \Tile_X4Y9_FrameData_O[13] ;
 wire \Tile_X4Y9_FrameData_O[14] ;
 wire \Tile_X4Y9_FrameData_O[15] ;
 wire \Tile_X4Y9_FrameData_O[16] ;
 wire \Tile_X4Y9_FrameData_O[17] ;
 wire \Tile_X4Y9_FrameData_O[18] ;
 wire \Tile_X4Y9_FrameData_O[19] ;
 wire \Tile_X4Y9_FrameData_O[1] ;
 wire \Tile_X4Y9_FrameData_O[20] ;
 wire \Tile_X4Y9_FrameData_O[21] ;
 wire \Tile_X4Y9_FrameData_O[22] ;
 wire \Tile_X4Y9_FrameData_O[23] ;
 wire \Tile_X4Y9_FrameData_O[24] ;
 wire \Tile_X4Y9_FrameData_O[25] ;
 wire \Tile_X4Y9_FrameData_O[26] ;
 wire \Tile_X4Y9_FrameData_O[27] ;
 wire \Tile_X4Y9_FrameData_O[28] ;
 wire \Tile_X4Y9_FrameData_O[29] ;
 wire \Tile_X4Y9_FrameData_O[2] ;
 wire \Tile_X4Y9_FrameData_O[30] ;
 wire \Tile_X4Y9_FrameData_O[31] ;
 wire \Tile_X4Y9_FrameData_O[3] ;
 wire \Tile_X4Y9_FrameData_O[4] ;
 wire \Tile_X4Y9_FrameData_O[5] ;
 wire \Tile_X4Y9_FrameData_O[6] ;
 wire \Tile_X4Y9_FrameData_O[7] ;
 wire \Tile_X4Y9_FrameData_O[8] ;
 wire \Tile_X4Y9_FrameData_O[9] ;
 wire \Tile_X4Y9_FrameStrobe_O[0] ;
 wire \Tile_X4Y9_FrameStrobe_O[10] ;
 wire \Tile_X4Y9_FrameStrobe_O[11] ;
 wire \Tile_X4Y9_FrameStrobe_O[12] ;
 wire \Tile_X4Y9_FrameStrobe_O[13] ;
 wire \Tile_X4Y9_FrameStrobe_O[14] ;
 wire \Tile_X4Y9_FrameStrobe_O[15] ;
 wire \Tile_X4Y9_FrameStrobe_O[16] ;
 wire \Tile_X4Y9_FrameStrobe_O[17] ;
 wire \Tile_X4Y9_FrameStrobe_O[18] ;
 wire \Tile_X4Y9_FrameStrobe_O[19] ;
 wire \Tile_X4Y9_FrameStrobe_O[1] ;
 wire \Tile_X4Y9_FrameStrobe_O[2] ;
 wire \Tile_X4Y9_FrameStrobe_O[3] ;
 wire \Tile_X4Y9_FrameStrobe_O[4] ;
 wire \Tile_X4Y9_FrameStrobe_O[5] ;
 wire \Tile_X4Y9_FrameStrobe_O[6] ;
 wire \Tile_X4Y9_FrameStrobe_O[7] ;
 wire \Tile_X4Y9_FrameStrobe_O[8] ;
 wire \Tile_X4Y9_FrameStrobe_O[9] ;
 wire \Tile_X4Y9_N1BEG[0] ;
 wire \Tile_X4Y9_N1BEG[1] ;
 wire \Tile_X4Y9_N1BEG[2] ;
 wire \Tile_X4Y9_N1BEG[3] ;
 wire \Tile_X4Y9_N2BEG[0] ;
 wire \Tile_X4Y9_N2BEG[1] ;
 wire \Tile_X4Y9_N2BEG[2] ;
 wire \Tile_X4Y9_N2BEG[3] ;
 wire \Tile_X4Y9_N2BEG[4] ;
 wire \Tile_X4Y9_N2BEG[5] ;
 wire \Tile_X4Y9_N2BEG[6] ;
 wire \Tile_X4Y9_N2BEG[7] ;
 wire \Tile_X4Y9_N2BEGb[0] ;
 wire \Tile_X4Y9_N2BEGb[1] ;
 wire \Tile_X4Y9_N2BEGb[2] ;
 wire \Tile_X4Y9_N2BEGb[3] ;
 wire \Tile_X4Y9_N2BEGb[4] ;
 wire \Tile_X4Y9_N2BEGb[5] ;
 wire \Tile_X4Y9_N2BEGb[6] ;
 wire \Tile_X4Y9_N2BEGb[7] ;
 wire \Tile_X4Y9_N4BEG[0] ;
 wire \Tile_X4Y9_N4BEG[10] ;
 wire \Tile_X4Y9_N4BEG[11] ;
 wire \Tile_X4Y9_N4BEG[12] ;
 wire \Tile_X4Y9_N4BEG[13] ;
 wire \Tile_X4Y9_N4BEG[14] ;
 wire \Tile_X4Y9_N4BEG[15] ;
 wire \Tile_X4Y9_N4BEG[1] ;
 wire \Tile_X4Y9_N4BEG[2] ;
 wire \Tile_X4Y9_N4BEG[3] ;
 wire \Tile_X4Y9_N4BEG[4] ;
 wire \Tile_X4Y9_N4BEG[5] ;
 wire \Tile_X4Y9_N4BEG[6] ;
 wire \Tile_X4Y9_N4BEG[7] ;
 wire \Tile_X4Y9_N4BEG[8] ;
 wire \Tile_X4Y9_N4BEG[9] ;
 wire \Tile_X4Y9_NN4BEG[0] ;
 wire \Tile_X4Y9_NN4BEG[10] ;
 wire \Tile_X4Y9_NN4BEG[11] ;
 wire \Tile_X4Y9_NN4BEG[12] ;
 wire \Tile_X4Y9_NN4BEG[13] ;
 wire \Tile_X4Y9_NN4BEG[14] ;
 wire \Tile_X4Y9_NN4BEG[15] ;
 wire \Tile_X4Y9_NN4BEG[1] ;
 wire \Tile_X4Y9_NN4BEG[2] ;
 wire \Tile_X4Y9_NN4BEG[3] ;
 wire \Tile_X4Y9_NN4BEG[4] ;
 wire \Tile_X4Y9_NN4BEG[5] ;
 wire \Tile_X4Y9_NN4BEG[6] ;
 wire \Tile_X4Y9_NN4BEG[7] ;
 wire \Tile_X4Y9_NN4BEG[8] ;
 wire \Tile_X4Y9_NN4BEG[9] ;
 wire \Tile_X4Y9_S1BEG[0] ;
 wire \Tile_X4Y9_S1BEG[1] ;
 wire \Tile_X4Y9_S1BEG[2] ;
 wire \Tile_X4Y9_S1BEG[3] ;
 wire \Tile_X4Y9_S2BEG[0] ;
 wire \Tile_X4Y9_S2BEG[1] ;
 wire \Tile_X4Y9_S2BEG[2] ;
 wire \Tile_X4Y9_S2BEG[3] ;
 wire \Tile_X4Y9_S2BEG[4] ;
 wire \Tile_X4Y9_S2BEG[5] ;
 wire \Tile_X4Y9_S2BEG[6] ;
 wire \Tile_X4Y9_S2BEG[7] ;
 wire \Tile_X4Y9_S2BEGb[0] ;
 wire \Tile_X4Y9_S2BEGb[1] ;
 wire \Tile_X4Y9_S2BEGb[2] ;
 wire \Tile_X4Y9_S2BEGb[3] ;
 wire \Tile_X4Y9_S2BEGb[4] ;
 wire \Tile_X4Y9_S2BEGb[5] ;
 wire \Tile_X4Y9_S2BEGb[6] ;
 wire \Tile_X4Y9_S2BEGb[7] ;
 wire \Tile_X4Y9_S4BEG[0] ;
 wire \Tile_X4Y9_S4BEG[10] ;
 wire \Tile_X4Y9_S4BEG[11] ;
 wire \Tile_X4Y9_S4BEG[12] ;
 wire \Tile_X4Y9_S4BEG[13] ;
 wire \Tile_X4Y9_S4BEG[14] ;
 wire \Tile_X4Y9_S4BEG[15] ;
 wire \Tile_X4Y9_S4BEG[1] ;
 wire \Tile_X4Y9_S4BEG[2] ;
 wire \Tile_X4Y9_S4BEG[3] ;
 wire \Tile_X4Y9_S4BEG[4] ;
 wire \Tile_X4Y9_S4BEG[5] ;
 wire \Tile_X4Y9_S4BEG[6] ;
 wire \Tile_X4Y9_S4BEG[7] ;
 wire \Tile_X4Y9_S4BEG[8] ;
 wire \Tile_X4Y9_S4BEG[9] ;
 wire \Tile_X4Y9_SS4BEG[0] ;
 wire \Tile_X4Y9_SS4BEG[10] ;
 wire \Tile_X4Y9_SS4BEG[11] ;
 wire \Tile_X4Y9_SS4BEG[12] ;
 wire \Tile_X4Y9_SS4BEG[13] ;
 wire \Tile_X4Y9_SS4BEG[14] ;
 wire \Tile_X4Y9_SS4BEG[15] ;
 wire \Tile_X4Y9_SS4BEG[1] ;
 wire \Tile_X4Y9_SS4BEG[2] ;
 wire \Tile_X4Y9_SS4BEG[3] ;
 wire \Tile_X4Y9_SS4BEG[4] ;
 wire \Tile_X4Y9_SS4BEG[5] ;
 wire \Tile_X4Y9_SS4BEG[6] ;
 wire \Tile_X4Y9_SS4BEG[7] ;
 wire \Tile_X4Y9_SS4BEG[8] ;
 wire \Tile_X4Y9_SS4BEG[9] ;
 wire Tile_X4Y9_UserCLKo;
 wire \Tile_X4Y9_W1BEG[0] ;
 wire \Tile_X4Y9_W1BEG[1] ;
 wire \Tile_X4Y9_W1BEG[2] ;
 wire \Tile_X4Y9_W1BEG[3] ;
 wire \Tile_X4Y9_W2BEG[0] ;
 wire \Tile_X4Y9_W2BEG[1] ;
 wire \Tile_X4Y9_W2BEG[2] ;
 wire \Tile_X4Y9_W2BEG[3] ;
 wire \Tile_X4Y9_W2BEG[4] ;
 wire \Tile_X4Y9_W2BEG[5] ;
 wire \Tile_X4Y9_W2BEG[6] ;
 wire \Tile_X4Y9_W2BEG[7] ;
 wire \Tile_X4Y9_W2BEGb[0] ;
 wire \Tile_X4Y9_W2BEGb[1] ;
 wire \Tile_X4Y9_W2BEGb[2] ;
 wire \Tile_X4Y9_W2BEGb[3] ;
 wire \Tile_X4Y9_W2BEGb[4] ;
 wire \Tile_X4Y9_W2BEGb[5] ;
 wire \Tile_X4Y9_W2BEGb[6] ;
 wire \Tile_X4Y9_W2BEGb[7] ;
 wire \Tile_X4Y9_W6BEG[0] ;
 wire \Tile_X4Y9_W6BEG[10] ;
 wire \Tile_X4Y9_W6BEG[11] ;
 wire \Tile_X4Y9_W6BEG[1] ;
 wire \Tile_X4Y9_W6BEG[2] ;
 wire \Tile_X4Y9_W6BEG[3] ;
 wire \Tile_X4Y9_W6BEG[4] ;
 wire \Tile_X4Y9_W6BEG[5] ;
 wire \Tile_X4Y9_W6BEG[6] ;
 wire \Tile_X4Y9_W6BEG[7] ;
 wire \Tile_X4Y9_W6BEG[8] ;
 wire \Tile_X4Y9_W6BEG[9] ;
 wire \Tile_X4Y9_WW4BEG[0] ;
 wire \Tile_X4Y9_WW4BEG[10] ;
 wire \Tile_X4Y9_WW4BEG[11] ;
 wire \Tile_X4Y9_WW4BEG[12] ;
 wire \Tile_X4Y9_WW4BEG[13] ;
 wire \Tile_X4Y9_WW4BEG[14] ;
 wire \Tile_X4Y9_WW4BEG[15] ;
 wire \Tile_X4Y9_WW4BEG[1] ;
 wire \Tile_X4Y9_WW4BEG[2] ;
 wire \Tile_X4Y9_WW4BEG[3] ;
 wire \Tile_X4Y9_WW4BEG[4] ;
 wire \Tile_X4Y9_WW4BEG[5] ;
 wire \Tile_X4Y9_WW4BEG[6] ;
 wire \Tile_X4Y9_WW4BEG[7] ;
 wire \Tile_X4Y9_WW4BEG[8] ;
 wire \Tile_X4Y9_WW4BEG[9] ;
 wire \Tile_X5Y0_FrameData_O[0] ;
 wire \Tile_X5Y0_FrameData_O[10] ;
 wire \Tile_X5Y0_FrameData_O[11] ;
 wire \Tile_X5Y0_FrameData_O[12] ;
 wire \Tile_X5Y0_FrameData_O[13] ;
 wire \Tile_X5Y0_FrameData_O[14] ;
 wire \Tile_X5Y0_FrameData_O[15] ;
 wire \Tile_X5Y0_FrameData_O[16] ;
 wire \Tile_X5Y0_FrameData_O[17] ;
 wire \Tile_X5Y0_FrameData_O[18] ;
 wire \Tile_X5Y0_FrameData_O[19] ;
 wire \Tile_X5Y0_FrameData_O[1] ;
 wire \Tile_X5Y0_FrameData_O[20] ;
 wire \Tile_X5Y0_FrameData_O[21] ;
 wire \Tile_X5Y0_FrameData_O[22] ;
 wire \Tile_X5Y0_FrameData_O[23] ;
 wire \Tile_X5Y0_FrameData_O[24] ;
 wire \Tile_X5Y0_FrameData_O[25] ;
 wire \Tile_X5Y0_FrameData_O[26] ;
 wire \Tile_X5Y0_FrameData_O[27] ;
 wire \Tile_X5Y0_FrameData_O[28] ;
 wire \Tile_X5Y0_FrameData_O[29] ;
 wire \Tile_X5Y0_FrameData_O[2] ;
 wire \Tile_X5Y0_FrameData_O[30] ;
 wire \Tile_X5Y0_FrameData_O[31] ;
 wire \Tile_X5Y0_FrameData_O[3] ;
 wire \Tile_X5Y0_FrameData_O[4] ;
 wire \Tile_X5Y0_FrameData_O[5] ;
 wire \Tile_X5Y0_FrameData_O[6] ;
 wire \Tile_X5Y0_FrameData_O[7] ;
 wire \Tile_X5Y0_FrameData_O[8] ;
 wire \Tile_X5Y0_FrameData_O[9] ;
 wire \Tile_X5Y0_FrameStrobe_O[0] ;
 wire \Tile_X5Y0_FrameStrobe_O[10] ;
 wire \Tile_X5Y0_FrameStrobe_O[11] ;
 wire \Tile_X5Y0_FrameStrobe_O[12] ;
 wire \Tile_X5Y0_FrameStrobe_O[13] ;
 wire \Tile_X5Y0_FrameStrobe_O[14] ;
 wire \Tile_X5Y0_FrameStrobe_O[15] ;
 wire \Tile_X5Y0_FrameStrobe_O[16] ;
 wire \Tile_X5Y0_FrameStrobe_O[17] ;
 wire \Tile_X5Y0_FrameStrobe_O[18] ;
 wire \Tile_X5Y0_FrameStrobe_O[19] ;
 wire \Tile_X5Y0_FrameStrobe_O[1] ;
 wire \Tile_X5Y0_FrameStrobe_O[2] ;
 wire \Tile_X5Y0_FrameStrobe_O[3] ;
 wire \Tile_X5Y0_FrameStrobe_O[4] ;
 wire \Tile_X5Y0_FrameStrobe_O[5] ;
 wire \Tile_X5Y0_FrameStrobe_O[6] ;
 wire \Tile_X5Y0_FrameStrobe_O[7] ;
 wire \Tile_X5Y0_FrameStrobe_O[8] ;
 wire \Tile_X5Y0_FrameStrobe_O[9] ;
 wire \Tile_X5Y0_S1BEG[0] ;
 wire \Tile_X5Y0_S1BEG[1] ;
 wire \Tile_X5Y0_S1BEG[2] ;
 wire \Tile_X5Y0_S1BEG[3] ;
 wire \Tile_X5Y0_S2BEG[0] ;
 wire \Tile_X5Y0_S2BEG[1] ;
 wire \Tile_X5Y0_S2BEG[2] ;
 wire \Tile_X5Y0_S2BEG[3] ;
 wire \Tile_X5Y0_S2BEG[4] ;
 wire \Tile_X5Y0_S2BEG[5] ;
 wire \Tile_X5Y0_S2BEG[6] ;
 wire \Tile_X5Y0_S2BEG[7] ;
 wire \Tile_X5Y0_S2BEGb[0] ;
 wire \Tile_X5Y0_S2BEGb[1] ;
 wire \Tile_X5Y0_S2BEGb[2] ;
 wire \Tile_X5Y0_S2BEGb[3] ;
 wire \Tile_X5Y0_S2BEGb[4] ;
 wire \Tile_X5Y0_S2BEGb[5] ;
 wire \Tile_X5Y0_S2BEGb[6] ;
 wire \Tile_X5Y0_S2BEGb[7] ;
 wire \Tile_X5Y0_S4BEG[0] ;
 wire \Tile_X5Y0_S4BEG[10] ;
 wire \Tile_X5Y0_S4BEG[11] ;
 wire \Tile_X5Y0_S4BEG[12] ;
 wire \Tile_X5Y0_S4BEG[13] ;
 wire \Tile_X5Y0_S4BEG[14] ;
 wire \Tile_X5Y0_S4BEG[15] ;
 wire \Tile_X5Y0_S4BEG[1] ;
 wire \Tile_X5Y0_S4BEG[2] ;
 wire \Tile_X5Y0_S4BEG[3] ;
 wire \Tile_X5Y0_S4BEG[4] ;
 wire \Tile_X5Y0_S4BEG[5] ;
 wire \Tile_X5Y0_S4BEG[6] ;
 wire \Tile_X5Y0_S4BEG[7] ;
 wire \Tile_X5Y0_S4BEG[8] ;
 wire \Tile_X5Y0_S4BEG[9] ;
 wire \Tile_X5Y0_SS4BEG[0] ;
 wire \Tile_X5Y0_SS4BEG[10] ;
 wire \Tile_X5Y0_SS4BEG[11] ;
 wire \Tile_X5Y0_SS4BEG[12] ;
 wire \Tile_X5Y0_SS4BEG[13] ;
 wire \Tile_X5Y0_SS4BEG[14] ;
 wire \Tile_X5Y0_SS4BEG[15] ;
 wire \Tile_X5Y0_SS4BEG[1] ;
 wire \Tile_X5Y0_SS4BEG[2] ;
 wire \Tile_X5Y0_SS4BEG[3] ;
 wire \Tile_X5Y0_SS4BEG[4] ;
 wire \Tile_X5Y0_SS4BEG[5] ;
 wire \Tile_X5Y0_SS4BEG[6] ;
 wire \Tile_X5Y0_SS4BEG[7] ;
 wire \Tile_X5Y0_SS4BEG[8] ;
 wire \Tile_X5Y0_SS4BEG[9] ;
 wire Tile_X5Y0_UserCLKo;
 wire Tile_X5Y10_Co;
 wire \Tile_X5Y10_E1BEG[0] ;
 wire \Tile_X5Y10_E1BEG[1] ;
 wire \Tile_X5Y10_E1BEG[2] ;
 wire \Tile_X5Y10_E1BEG[3] ;
 wire \Tile_X5Y10_E2BEG[0] ;
 wire \Tile_X5Y10_E2BEG[1] ;
 wire \Tile_X5Y10_E2BEG[2] ;
 wire \Tile_X5Y10_E2BEG[3] ;
 wire \Tile_X5Y10_E2BEG[4] ;
 wire \Tile_X5Y10_E2BEG[5] ;
 wire \Tile_X5Y10_E2BEG[6] ;
 wire \Tile_X5Y10_E2BEG[7] ;
 wire \Tile_X5Y10_E2BEGb[0] ;
 wire \Tile_X5Y10_E2BEGb[1] ;
 wire \Tile_X5Y10_E2BEGb[2] ;
 wire \Tile_X5Y10_E2BEGb[3] ;
 wire \Tile_X5Y10_E2BEGb[4] ;
 wire \Tile_X5Y10_E2BEGb[5] ;
 wire \Tile_X5Y10_E2BEGb[6] ;
 wire \Tile_X5Y10_E2BEGb[7] ;
 wire \Tile_X5Y10_E6BEG[0] ;
 wire \Tile_X5Y10_E6BEG[10] ;
 wire \Tile_X5Y10_E6BEG[11] ;
 wire \Tile_X5Y10_E6BEG[1] ;
 wire \Tile_X5Y10_E6BEG[2] ;
 wire \Tile_X5Y10_E6BEG[3] ;
 wire \Tile_X5Y10_E6BEG[4] ;
 wire \Tile_X5Y10_E6BEG[5] ;
 wire \Tile_X5Y10_E6BEG[6] ;
 wire \Tile_X5Y10_E6BEG[7] ;
 wire \Tile_X5Y10_E6BEG[8] ;
 wire \Tile_X5Y10_E6BEG[9] ;
 wire \Tile_X5Y10_EE4BEG[0] ;
 wire \Tile_X5Y10_EE4BEG[10] ;
 wire \Tile_X5Y10_EE4BEG[11] ;
 wire \Tile_X5Y10_EE4BEG[12] ;
 wire \Tile_X5Y10_EE4BEG[13] ;
 wire \Tile_X5Y10_EE4BEG[14] ;
 wire \Tile_X5Y10_EE4BEG[15] ;
 wire \Tile_X5Y10_EE4BEG[1] ;
 wire \Tile_X5Y10_EE4BEG[2] ;
 wire \Tile_X5Y10_EE4BEG[3] ;
 wire \Tile_X5Y10_EE4BEG[4] ;
 wire \Tile_X5Y10_EE4BEG[5] ;
 wire \Tile_X5Y10_EE4BEG[6] ;
 wire \Tile_X5Y10_EE4BEG[7] ;
 wire \Tile_X5Y10_EE4BEG[8] ;
 wire \Tile_X5Y10_EE4BEG[9] ;
 wire \Tile_X5Y10_FrameData_O[0] ;
 wire \Tile_X5Y10_FrameData_O[10] ;
 wire \Tile_X5Y10_FrameData_O[11] ;
 wire \Tile_X5Y10_FrameData_O[12] ;
 wire \Tile_X5Y10_FrameData_O[13] ;
 wire \Tile_X5Y10_FrameData_O[14] ;
 wire \Tile_X5Y10_FrameData_O[15] ;
 wire \Tile_X5Y10_FrameData_O[16] ;
 wire \Tile_X5Y10_FrameData_O[17] ;
 wire \Tile_X5Y10_FrameData_O[18] ;
 wire \Tile_X5Y10_FrameData_O[19] ;
 wire \Tile_X5Y10_FrameData_O[1] ;
 wire \Tile_X5Y10_FrameData_O[20] ;
 wire \Tile_X5Y10_FrameData_O[21] ;
 wire \Tile_X5Y10_FrameData_O[22] ;
 wire \Tile_X5Y10_FrameData_O[23] ;
 wire \Tile_X5Y10_FrameData_O[24] ;
 wire \Tile_X5Y10_FrameData_O[25] ;
 wire \Tile_X5Y10_FrameData_O[26] ;
 wire \Tile_X5Y10_FrameData_O[27] ;
 wire \Tile_X5Y10_FrameData_O[28] ;
 wire \Tile_X5Y10_FrameData_O[29] ;
 wire \Tile_X5Y10_FrameData_O[2] ;
 wire \Tile_X5Y10_FrameData_O[30] ;
 wire \Tile_X5Y10_FrameData_O[31] ;
 wire \Tile_X5Y10_FrameData_O[3] ;
 wire \Tile_X5Y10_FrameData_O[4] ;
 wire \Tile_X5Y10_FrameData_O[5] ;
 wire \Tile_X5Y10_FrameData_O[6] ;
 wire \Tile_X5Y10_FrameData_O[7] ;
 wire \Tile_X5Y10_FrameData_O[8] ;
 wire \Tile_X5Y10_FrameData_O[9] ;
 wire \Tile_X5Y10_FrameStrobe_O[0] ;
 wire \Tile_X5Y10_FrameStrobe_O[10] ;
 wire \Tile_X5Y10_FrameStrobe_O[11] ;
 wire \Tile_X5Y10_FrameStrobe_O[12] ;
 wire \Tile_X5Y10_FrameStrobe_O[13] ;
 wire \Tile_X5Y10_FrameStrobe_O[14] ;
 wire \Tile_X5Y10_FrameStrobe_O[15] ;
 wire \Tile_X5Y10_FrameStrobe_O[16] ;
 wire \Tile_X5Y10_FrameStrobe_O[17] ;
 wire \Tile_X5Y10_FrameStrobe_O[18] ;
 wire \Tile_X5Y10_FrameStrobe_O[19] ;
 wire \Tile_X5Y10_FrameStrobe_O[1] ;
 wire \Tile_X5Y10_FrameStrobe_O[2] ;
 wire \Tile_X5Y10_FrameStrobe_O[3] ;
 wire \Tile_X5Y10_FrameStrobe_O[4] ;
 wire \Tile_X5Y10_FrameStrobe_O[5] ;
 wire \Tile_X5Y10_FrameStrobe_O[6] ;
 wire \Tile_X5Y10_FrameStrobe_O[7] ;
 wire \Tile_X5Y10_FrameStrobe_O[8] ;
 wire \Tile_X5Y10_FrameStrobe_O[9] ;
 wire \Tile_X5Y10_N1BEG[0] ;
 wire \Tile_X5Y10_N1BEG[1] ;
 wire \Tile_X5Y10_N1BEG[2] ;
 wire \Tile_X5Y10_N1BEG[3] ;
 wire \Tile_X5Y10_N2BEG[0] ;
 wire \Tile_X5Y10_N2BEG[1] ;
 wire \Tile_X5Y10_N2BEG[2] ;
 wire \Tile_X5Y10_N2BEG[3] ;
 wire \Tile_X5Y10_N2BEG[4] ;
 wire \Tile_X5Y10_N2BEG[5] ;
 wire \Tile_X5Y10_N2BEG[6] ;
 wire \Tile_X5Y10_N2BEG[7] ;
 wire \Tile_X5Y10_N2BEGb[0] ;
 wire \Tile_X5Y10_N2BEGb[1] ;
 wire \Tile_X5Y10_N2BEGb[2] ;
 wire \Tile_X5Y10_N2BEGb[3] ;
 wire \Tile_X5Y10_N2BEGb[4] ;
 wire \Tile_X5Y10_N2BEGb[5] ;
 wire \Tile_X5Y10_N2BEGb[6] ;
 wire \Tile_X5Y10_N2BEGb[7] ;
 wire \Tile_X5Y10_N4BEG[0] ;
 wire \Tile_X5Y10_N4BEG[10] ;
 wire \Tile_X5Y10_N4BEG[11] ;
 wire \Tile_X5Y10_N4BEG[12] ;
 wire \Tile_X5Y10_N4BEG[13] ;
 wire \Tile_X5Y10_N4BEG[14] ;
 wire \Tile_X5Y10_N4BEG[15] ;
 wire \Tile_X5Y10_N4BEG[1] ;
 wire \Tile_X5Y10_N4BEG[2] ;
 wire \Tile_X5Y10_N4BEG[3] ;
 wire \Tile_X5Y10_N4BEG[4] ;
 wire \Tile_X5Y10_N4BEG[5] ;
 wire \Tile_X5Y10_N4BEG[6] ;
 wire \Tile_X5Y10_N4BEG[7] ;
 wire \Tile_X5Y10_N4BEG[8] ;
 wire \Tile_X5Y10_N4BEG[9] ;
 wire \Tile_X5Y10_NN4BEG[0] ;
 wire \Tile_X5Y10_NN4BEG[10] ;
 wire \Tile_X5Y10_NN4BEG[11] ;
 wire \Tile_X5Y10_NN4BEG[12] ;
 wire \Tile_X5Y10_NN4BEG[13] ;
 wire \Tile_X5Y10_NN4BEG[14] ;
 wire \Tile_X5Y10_NN4BEG[15] ;
 wire \Tile_X5Y10_NN4BEG[1] ;
 wire \Tile_X5Y10_NN4BEG[2] ;
 wire \Tile_X5Y10_NN4BEG[3] ;
 wire \Tile_X5Y10_NN4BEG[4] ;
 wire \Tile_X5Y10_NN4BEG[5] ;
 wire \Tile_X5Y10_NN4BEG[6] ;
 wire \Tile_X5Y10_NN4BEG[7] ;
 wire \Tile_X5Y10_NN4BEG[8] ;
 wire \Tile_X5Y10_NN4BEG[9] ;
 wire \Tile_X5Y10_S1BEG[0] ;
 wire \Tile_X5Y10_S1BEG[1] ;
 wire \Tile_X5Y10_S1BEG[2] ;
 wire \Tile_X5Y10_S1BEG[3] ;
 wire \Tile_X5Y10_S2BEG[0] ;
 wire \Tile_X5Y10_S2BEG[1] ;
 wire \Tile_X5Y10_S2BEG[2] ;
 wire \Tile_X5Y10_S2BEG[3] ;
 wire \Tile_X5Y10_S2BEG[4] ;
 wire \Tile_X5Y10_S2BEG[5] ;
 wire \Tile_X5Y10_S2BEG[6] ;
 wire \Tile_X5Y10_S2BEG[7] ;
 wire \Tile_X5Y10_S2BEGb[0] ;
 wire \Tile_X5Y10_S2BEGb[1] ;
 wire \Tile_X5Y10_S2BEGb[2] ;
 wire \Tile_X5Y10_S2BEGb[3] ;
 wire \Tile_X5Y10_S2BEGb[4] ;
 wire \Tile_X5Y10_S2BEGb[5] ;
 wire \Tile_X5Y10_S2BEGb[6] ;
 wire \Tile_X5Y10_S2BEGb[7] ;
 wire \Tile_X5Y10_S4BEG[0] ;
 wire \Tile_X5Y10_S4BEG[10] ;
 wire \Tile_X5Y10_S4BEG[11] ;
 wire \Tile_X5Y10_S4BEG[12] ;
 wire \Tile_X5Y10_S4BEG[13] ;
 wire \Tile_X5Y10_S4BEG[14] ;
 wire \Tile_X5Y10_S4BEG[15] ;
 wire \Tile_X5Y10_S4BEG[1] ;
 wire \Tile_X5Y10_S4BEG[2] ;
 wire \Tile_X5Y10_S4BEG[3] ;
 wire \Tile_X5Y10_S4BEG[4] ;
 wire \Tile_X5Y10_S4BEG[5] ;
 wire \Tile_X5Y10_S4BEG[6] ;
 wire \Tile_X5Y10_S4BEG[7] ;
 wire \Tile_X5Y10_S4BEG[8] ;
 wire \Tile_X5Y10_S4BEG[9] ;
 wire \Tile_X5Y10_SS4BEG[0] ;
 wire \Tile_X5Y10_SS4BEG[10] ;
 wire \Tile_X5Y10_SS4BEG[11] ;
 wire \Tile_X5Y10_SS4BEG[12] ;
 wire \Tile_X5Y10_SS4BEG[13] ;
 wire \Tile_X5Y10_SS4BEG[14] ;
 wire \Tile_X5Y10_SS4BEG[15] ;
 wire \Tile_X5Y10_SS4BEG[1] ;
 wire \Tile_X5Y10_SS4BEG[2] ;
 wire \Tile_X5Y10_SS4BEG[3] ;
 wire \Tile_X5Y10_SS4BEG[4] ;
 wire \Tile_X5Y10_SS4BEG[5] ;
 wire \Tile_X5Y10_SS4BEG[6] ;
 wire \Tile_X5Y10_SS4BEG[7] ;
 wire \Tile_X5Y10_SS4BEG[8] ;
 wire \Tile_X5Y10_SS4BEG[9] ;
 wire Tile_X5Y10_UserCLKo;
 wire \Tile_X5Y10_W1BEG[0] ;
 wire \Tile_X5Y10_W1BEG[1] ;
 wire \Tile_X5Y10_W1BEG[2] ;
 wire \Tile_X5Y10_W1BEG[3] ;
 wire \Tile_X5Y10_W2BEG[0] ;
 wire \Tile_X5Y10_W2BEG[1] ;
 wire \Tile_X5Y10_W2BEG[2] ;
 wire \Tile_X5Y10_W2BEG[3] ;
 wire \Tile_X5Y10_W2BEG[4] ;
 wire \Tile_X5Y10_W2BEG[5] ;
 wire \Tile_X5Y10_W2BEG[6] ;
 wire \Tile_X5Y10_W2BEG[7] ;
 wire \Tile_X5Y10_W2BEGb[0] ;
 wire \Tile_X5Y10_W2BEGb[1] ;
 wire \Tile_X5Y10_W2BEGb[2] ;
 wire \Tile_X5Y10_W2BEGb[3] ;
 wire \Tile_X5Y10_W2BEGb[4] ;
 wire \Tile_X5Y10_W2BEGb[5] ;
 wire \Tile_X5Y10_W2BEGb[6] ;
 wire \Tile_X5Y10_W2BEGb[7] ;
 wire \Tile_X5Y10_W6BEG[0] ;
 wire \Tile_X5Y10_W6BEG[10] ;
 wire \Tile_X5Y10_W6BEG[11] ;
 wire \Tile_X5Y10_W6BEG[1] ;
 wire \Tile_X5Y10_W6BEG[2] ;
 wire \Tile_X5Y10_W6BEG[3] ;
 wire \Tile_X5Y10_W6BEG[4] ;
 wire \Tile_X5Y10_W6BEG[5] ;
 wire \Tile_X5Y10_W6BEG[6] ;
 wire \Tile_X5Y10_W6BEG[7] ;
 wire \Tile_X5Y10_W6BEG[8] ;
 wire \Tile_X5Y10_W6BEG[9] ;
 wire \Tile_X5Y10_WW4BEG[0] ;
 wire \Tile_X5Y10_WW4BEG[10] ;
 wire \Tile_X5Y10_WW4BEG[11] ;
 wire \Tile_X5Y10_WW4BEG[12] ;
 wire \Tile_X5Y10_WW4BEG[13] ;
 wire \Tile_X5Y10_WW4BEG[14] ;
 wire \Tile_X5Y10_WW4BEG[15] ;
 wire \Tile_X5Y10_WW4BEG[1] ;
 wire \Tile_X5Y10_WW4BEG[2] ;
 wire \Tile_X5Y10_WW4BEG[3] ;
 wire \Tile_X5Y10_WW4BEG[4] ;
 wire \Tile_X5Y10_WW4BEG[5] ;
 wire \Tile_X5Y10_WW4BEG[6] ;
 wire \Tile_X5Y10_WW4BEG[7] ;
 wire \Tile_X5Y10_WW4BEG[8] ;
 wire \Tile_X5Y10_WW4BEG[9] ;
 wire Tile_X5Y11_Co;
 wire \Tile_X5Y11_E1BEG[0] ;
 wire \Tile_X5Y11_E1BEG[1] ;
 wire \Tile_X5Y11_E1BEG[2] ;
 wire \Tile_X5Y11_E1BEG[3] ;
 wire \Tile_X5Y11_E2BEG[0] ;
 wire \Tile_X5Y11_E2BEG[1] ;
 wire \Tile_X5Y11_E2BEG[2] ;
 wire \Tile_X5Y11_E2BEG[3] ;
 wire \Tile_X5Y11_E2BEG[4] ;
 wire \Tile_X5Y11_E2BEG[5] ;
 wire \Tile_X5Y11_E2BEG[6] ;
 wire \Tile_X5Y11_E2BEG[7] ;
 wire \Tile_X5Y11_E2BEGb[0] ;
 wire \Tile_X5Y11_E2BEGb[1] ;
 wire \Tile_X5Y11_E2BEGb[2] ;
 wire \Tile_X5Y11_E2BEGb[3] ;
 wire \Tile_X5Y11_E2BEGb[4] ;
 wire \Tile_X5Y11_E2BEGb[5] ;
 wire \Tile_X5Y11_E2BEGb[6] ;
 wire \Tile_X5Y11_E2BEGb[7] ;
 wire \Tile_X5Y11_E6BEG[0] ;
 wire \Tile_X5Y11_E6BEG[10] ;
 wire \Tile_X5Y11_E6BEG[11] ;
 wire \Tile_X5Y11_E6BEG[1] ;
 wire \Tile_X5Y11_E6BEG[2] ;
 wire \Tile_X5Y11_E6BEG[3] ;
 wire \Tile_X5Y11_E6BEG[4] ;
 wire \Tile_X5Y11_E6BEG[5] ;
 wire \Tile_X5Y11_E6BEG[6] ;
 wire \Tile_X5Y11_E6BEG[7] ;
 wire \Tile_X5Y11_E6BEG[8] ;
 wire \Tile_X5Y11_E6BEG[9] ;
 wire \Tile_X5Y11_EE4BEG[0] ;
 wire \Tile_X5Y11_EE4BEG[10] ;
 wire \Tile_X5Y11_EE4BEG[11] ;
 wire \Tile_X5Y11_EE4BEG[12] ;
 wire \Tile_X5Y11_EE4BEG[13] ;
 wire \Tile_X5Y11_EE4BEG[14] ;
 wire \Tile_X5Y11_EE4BEG[15] ;
 wire \Tile_X5Y11_EE4BEG[1] ;
 wire \Tile_X5Y11_EE4BEG[2] ;
 wire \Tile_X5Y11_EE4BEG[3] ;
 wire \Tile_X5Y11_EE4BEG[4] ;
 wire \Tile_X5Y11_EE4BEG[5] ;
 wire \Tile_X5Y11_EE4BEG[6] ;
 wire \Tile_X5Y11_EE4BEG[7] ;
 wire \Tile_X5Y11_EE4BEG[8] ;
 wire \Tile_X5Y11_EE4BEG[9] ;
 wire \Tile_X5Y11_FrameData_O[0] ;
 wire \Tile_X5Y11_FrameData_O[10] ;
 wire \Tile_X5Y11_FrameData_O[11] ;
 wire \Tile_X5Y11_FrameData_O[12] ;
 wire \Tile_X5Y11_FrameData_O[13] ;
 wire \Tile_X5Y11_FrameData_O[14] ;
 wire \Tile_X5Y11_FrameData_O[15] ;
 wire \Tile_X5Y11_FrameData_O[16] ;
 wire \Tile_X5Y11_FrameData_O[17] ;
 wire \Tile_X5Y11_FrameData_O[18] ;
 wire \Tile_X5Y11_FrameData_O[19] ;
 wire \Tile_X5Y11_FrameData_O[1] ;
 wire \Tile_X5Y11_FrameData_O[20] ;
 wire \Tile_X5Y11_FrameData_O[21] ;
 wire \Tile_X5Y11_FrameData_O[22] ;
 wire \Tile_X5Y11_FrameData_O[23] ;
 wire \Tile_X5Y11_FrameData_O[24] ;
 wire \Tile_X5Y11_FrameData_O[25] ;
 wire \Tile_X5Y11_FrameData_O[26] ;
 wire \Tile_X5Y11_FrameData_O[27] ;
 wire \Tile_X5Y11_FrameData_O[28] ;
 wire \Tile_X5Y11_FrameData_O[29] ;
 wire \Tile_X5Y11_FrameData_O[2] ;
 wire \Tile_X5Y11_FrameData_O[30] ;
 wire \Tile_X5Y11_FrameData_O[31] ;
 wire \Tile_X5Y11_FrameData_O[3] ;
 wire \Tile_X5Y11_FrameData_O[4] ;
 wire \Tile_X5Y11_FrameData_O[5] ;
 wire \Tile_X5Y11_FrameData_O[6] ;
 wire \Tile_X5Y11_FrameData_O[7] ;
 wire \Tile_X5Y11_FrameData_O[8] ;
 wire \Tile_X5Y11_FrameData_O[9] ;
 wire \Tile_X5Y11_FrameStrobe_O[0] ;
 wire \Tile_X5Y11_FrameStrobe_O[10] ;
 wire \Tile_X5Y11_FrameStrobe_O[11] ;
 wire \Tile_X5Y11_FrameStrobe_O[12] ;
 wire \Tile_X5Y11_FrameStrobe_O[13] ;
 wire \Tile_X5Y11_FrameStrobe_O[14] ;
 wire \Tile_X5Y11_FrameStrobe_O[15] ;
 wire \Tile_X5Y11_FrameStrobe_O[16] ;
 wire \Tile_X5Y11_FrameStrobe_O[17] ;
 wire \Tile_X5Y11_FrameStrobe_O[18] ;
 wire \Tile_X5Y11_FrameStrobe_O[19] ;
 wire \Tile_X5Y11_FrameStrobe_O[1] ;
 wire \Tile_X5Y11_FrameStrobe_O[2] ;
 wire \Tile_X5Y11_FrameStrobe_O[3] ;
 wire \Tile_X5Y11_FrameStrobe_O[4] ;
 wire \Tile_X5Y11_FrameStrobe_O[5] ;
 wire \Tile_X5Y11_FrameStrobe_O[6] ;
 wire \Tile_X5Y11_FrameStrobe_O[7] ;
 wire \Tile_X5Y11_FrameStrobe_O[8] ;
 wire \Tile_X5Y11_FrameStrobe_O[9] ;
 wire \Tile_X5Y11_N1BEG[0] ;
 wire \Tile_X5Y11_N1BEG[1] ;
 wire \Tile_X5Y11_N1BEG[2] ;
 wire \Tile_X5Y11_N1BEG[3] ;
 wire \Tile_X5Y11_N2BEG[0] ;
 wire \Tile_X5Y11_N2BEG[1] ;
 wire \Tile_X5Y11_N2BEG[2] ;
 wire \Tile_X5Y11_N2BEG[3] ;
 wire \Tile_X5Y11_N2BEG[4] ;
 wire \Tile_X5Y11_N2BEG[5] ;
 wire \Tile_X5Y11_N2BEG[6] ;
 wire \Tile_X5Y11_N2BEG[7] ;
 wire \Tile_X5Y11_N2BEGb[0] ;
 wire \Tile_X5Y11_N2BEGb[1] ;
 wire \Tile_X5Y11_N2BEGb[2] ;
 wire \Tile_X5Y11_N2BEGb[3] ;
 wire \Tile_X5Y11_N2BEGb[4] ;
 wire \Tile_X5Y11_N2BEGb[5] ;
 wire \Tile_X5Y11_N2BEGb[6] ;
 wire \Tile_X5Y11_N2BEGb[7] ;
 wire \Tile_X5Y11_N4BEG[0] ;
 wire \Tile_X5Y11_N4BEG[10] ;
 wire \Tile_X5Y11_N4BEG[11] ;
 wire \Tile_X5Y11_N4BEG[12] ;
 wire \Tile_X5Y11_N4BEG[13] ;
 wire \Tile_X5Y11_N4BEG[14] ;
 wire \Tile_X5Y11_N4BEG[15] ;
 wire \Tile_X5Y11_N4BEG[1] ;
 wire \Tile_X5Y11_N4BEG[2] ;
 wire \Tile_X5Y11_N4BEG[3] ;
 wire \Tile_X5Y11_N4BEG[4] ;
 wire \Tile_X5Y11_N4BEG[5] ;
 wire \Tile_X5Y11_N4BEG[6] ;
 wire \Tile_X5Y11_N4BEG[7] ;
 wire \Tile_X5Y11_N4BEG[8] ;
 wire \Tile_X5Y11_N4BEG[9] ;
 wire \Tile_X5Y11_NN4BEG[0] ;
 wire \Tile_X5Y11_NN4BEG[10] ;
 wire \Tile_X5Y11_NN4BEG[11] ;
 wire \Tile_X5Y11_NN4BEG[12] ;
 wire \Tile_X5Y11_NN4BEG[13] ;
 wire \Tile_X5Y11_NN4BEG[14] ;
 wire \Tile_X5Y11_NN4BEG[15] ;
 wire \Tile_X5Y11_NN4BEG[1] ;
 wire \Tile_X5Y11_NN4BEG[2] ;
 wire \Tile_X5Y11_NN4BEG[3] ;
 wire \Tile_X5Y11_NN4BEG[4] ;
 wire \Tile_X5Y11_NN4BEG[5] ;
 wire \Tile_X5Y11_NN4BEG[6] ;
 wire \Tile_X5Y11_NN4BEG[7] ;
 wire \Tile_X5Y11_NN4BEG[8] ;
 wire \Tile_X5Y11_NN4BEG[9] ;
 wire \Tile_X5Y11_S1BEG[0] ;
 wire \Tile_X5Y11_S1BEG[1] ;
 wire \Tile_X5Y11_S1BEG[2] ;
 wire \Tile_X5Y11_S1BEG[3] ;
 wire \Tile_X5Y11_S2BEG[0] ;
 wire \Tile_X5Y11_S2BEG[1] ;
 wire \Tile_X5Y11_S2BEG[2] ;
 wire \Tile_X5Y11_S2BEG[3] ;
 wire \Tile_X5Y11_S2BEG[4] ;
 wire \Tile_X5Y11_S2BEG[5] ;
 wire \Tile_X5Y11_S2BEG[6] ;
 wire \Tile_X5Y11_S2BEG[7] ;
 wire \Tile_X5Y11_S2BEGb[0] ;
 wire \Tile_X5Y11_S2BEGb[1] ;
 wire \Tile_X5Y11_S2BEGb[2] ;
 wire \Tile_X5Y11_S2BEGb[3] ;
 wire \Tile_X5Y11_S2BEGb[4] ;
 wire \Tile_X5Y11_S2BEGb[5] ;
 wire \Tile_X5Y11_S2BEGb[6] ;
 wire \Tile_X5Y11_S2BEGb[7] ;
 wire \Tile_X5Y11_S4BEG[0] ;
 wire \Tile_X5Y11_S4BEG[10] ;
 wire \Tile_X5Y11_S4BEG[11] ;
 wire \Tile_X5Y11_S4BEG[12] ;
 wire \Tile_X5Y11_S4BEG[13] ;
 wire \Tile_X5Y11_S4BEG[14] ;
 wire \Tile_X5Y11_S4BEG[15] ;
 wire \Tile_X5Y11_S4BEG[1] ;
 wire \Tile_X5Y11_S4BEG[2] ;
 wire \Tile_X5Y11_S4BEG[3] ;
 wire \Tile_X5Y11_S4BEG[4] ;
 wire \Tile_X5Y11_S4BEG[5] ;
 wire \Tile_X5Y11_S4BEG[6] ;
 wire \Tile_X5Y11_S4BEG[7] ;
 wire \Tile_X5Y11_S4BEG[8] ;
 wire \Tile_X5Y11_S4BEG[9] ;
 wire \Tile_X5Y11_SS4BEG[0] ;
 wire \Tile_X5Y11_SS4BEG[10] ;
 wire \Tile_X5Y11_SS4BEG[11] ;
 wire \Tile_X5Y11_SS4BEG[12] ;
 wire \Tile_X5Y11_SS4BEG[13] ;
 wire \Tile_X5Y11_SS4BEG[14] ;
 wire \Tile_X5Y11_SS4BEG[15] ;
 wire \Tile_X5Y11_SS4BEG[1] ;
 wire \Tile_X5Y11_SS4BEG[2] ;
 wire \Tile_X5Y11_SS4BEG[3] ;
 wire \Tile_X5Y11_SS4BEG[4] ;
 wire \Tile_X5Y11_SS4BEG[5] ;
 wire \Tile_X5Y11_SS4BEG[6] ;
 wire \Tile_X5Y11_SS4BEG[7] ;
 wire \Tile_X5Y11_SS4BEG[8] ;
 wire \Tile_X5Y11_SS4BEG[9] ;
 wire Tile_X5Y11_UserCLKo;
 wire \Tile_X5Y11_W1BEG[0] ;
 wire \Tile_X5Y11_W1BEG[1] ;
 wire \Tile_X5Y11_W1BEG[2] ;
 wire \Tile_X5Y11_W1BEG[3] ;
 wire \Tile_X5Y11_W2BEG[0] ;
 wire \Tile_X5Y11_W2BEG[1] ;
 wire \Tile_X5Y11_W2BEG[2] ;
 wire \Tile_X5Y11_W2BEG[3] ;
 wire \Tile_X5Y11_W2BEG[4] ;
 wire \Tile_X5Y11_W2BEG[5] ;
 wire \Tile_X5Y11_W2BEG[6] ;
 wire \Tile_X5Y11_W2BEG[7] ;
 wire \Tile_X5Y11_W2BEGb[0] ;
 wire \Tile_X5Y11_W2BEGb[1] ;
 wire \Tile_X5Y11_W2BEGb[2] ;
 wire \Tile_X5Y11_W2BEGb[3] ;
 wire \Tile_X5Y11_W2BEGb[4] ;
 wire \Tile_X5Y11_W2BEGb[5] ;
 wire \Tile_X5Y11_W2BEGb[6] ;
 wire \Tile_X5Y11_W2BEGb[7] ;
 wire \Tile_X5Y11_W6BEG[0] ;
 wire \Tile_X5Y11_W6BEG[10] ;
 wire \Tile_X5Y11_W6BEG[11] ;
 wire \Tile_X5Y11_W6BEG[1] ;
 wire \Tile_X5Y11_W6BEG[2] ;
 wire \Tile_X5Y11_W6BEG[3] ;
 wire \Tile_X5Y11_W6BEG[4] ;
 wire \Tile_X5Y11_W6BEG[5] ;
 wire \Tile_X5Y11_W6BEG[6] ;
 wire \Tile_X5Y11_W6BEG[7] ;
 wire \Tile_X5Y11_W6BEG[8] ;
 wire \Tile_X5Y11_W6BEG[9] ;
 wire \Tile_X5Y11_WW4BEG[0] ;
 wire \Tile_X5Y11_WW4BEG[10] ;
 wire \Tile_X5Y11_WW4BEG[11] ;
 wire \Tile_X5Y11_WW4BEG[12] ;
 wire \Tile_X5Y11_WW4BEG[13] ;
 wire \Tile_X5Y11_WW4BEG[14] ;
 wire \Tile_X5Y11_WW4BEG[15] ;
 wire \Tile_X5Y11_WW4BEG[1] ;
 wire \Tile_X5Y11_WW4BEG[2] ;
 wire \Tile_X5Y11_WW4BEG[3] ;
 wire \Tile_X5Y11_WW4BEG[4] ;
 wire \Tile_X5Y11_WW4BEG[5] ;
 wire \Tile_X5Y11_WW4BEG[6] ;
 wire \Tile_X5Y11_WW4BEG[7] ;
 wire \Tile_X5Y11_WW4BEG[8] ;
 wire \Tile_X5Y11_WW4BEG[9] ;
 wire Tile_X5Y12_Co;
 wire \Tile_X5Y12_E1BEG[0] ;
 wire \Tile_X5Y12_E1BEG[1] ;
 wire \Tile_X5Y12_E1BEG[2] ;
 wire \Tile_X5Y12_E1BEG[3] ;
 wire \Tile_X5Y12_E2BEG[0] ;
 wire \Tile_X5Y12_E2BEG[1] ;
 wire \Tile_X5Y12_E2BEG[2] ;
 wire \Tile_X5Y12_E2BEG[3] ;
 wire \Tile_X5Y12_E2BEG[4] ;
 wire \Tile_X5Y12_E2BEG[5] ;
 wire \Tile_X5Y12_E2BEG[6] ;
 wire \Tile_X5Y12_E2BEG[7] ;
 wire \Tile_X5Y12_E2BEGb[0] ;
 wire \Tile_X5Y12_E2BEGb[1] ;
 wire \Tile_X5Y12_E2BEGb[2] ;
 wire \Tile_X5Y12_E2BEGb[3] ;
 wire \Tile_X5Y12_E2BEGb[4] ;
 wire \Tile_X5Y12_E2BEGb[5] ;
 wire \Tile_X5Y12_E2BEGb[6] ;
 wire \Tile_X5Y12_E2BEGb[7] ;
 wire \Tile_X5Y12_E6BEG[0] ;
 wire \Tile_X5Y12_E6BEG[10] ;
 wire \Tile_X5Y12_E6BEG[11] ;
 wire \Tile_X5Y12_E6BEG[1] ;
 wire \Tile_X5Y12_E6BEG[2] ;
 wire \Tile_X5Y12_E6BEG[3] ;
 wire \Tile_X5Y12_E6BEG[4] ;
 wire \Tile_X5Y12_E6BEG[5] ;
 wire \Tile_X5Y12_E6BEG[6] ;
 wire \Tile_X5Y12_E6BEG[7] ;
 wire \Tile_X5Y12_E6BEG[8] ;
 wire \Tile_X5Y12_E6BEG[9] ;
 wire \Tile_X5Y12_EE4BEG[0] ;
 wire \Tile_X5Y12_EE4BEG[10] ;
 wire \Tile_X5Y12_EE4BEG[11] ;
 wire \Tile_X5Y12_EE4BEG[12] ;
 wire \Tile_X5Y12_EE4BEG[13] ;
 wire \Tile_X5Y12_EE4BEG[14] ;
 wire \Tile_X5Y12_EE4BEG[15] ;
 wire \Tile_X5Y12_EE4BEG[1] ;
 wire \Tile_X5Y12_EE4BEG[2] ;
 wire \Tile_X5Y12_EE4BEG[3] ;
 wire \Tile_X5Y12_EE4BEG[4] ;
 wire \Tile_X5Y12_EE4BEG[5] ;
 wire \Tile_X5Y12_EE4BEG[6] ;
 wire \Tile_X5Y12_EE4BEG[7] ;
 wire \Tile_X5Y12_EE4BEG[8] ;
 wire \Tile_X5Y12_EE4BEG[9] ;
 wire \Tile_X5Y12_FrameData_O[0] ;
 wire \Tile_X5Y12_FrameData_O[10] ;
 wire \Tile_X5Y12_FrameData_O[11] ;
 wire \Tile_X5Y12_FrameData_O[12] ;
 wire \Tile_X5Y12_FrameData_O[13] ;
 wire \Tile_X5Y12_FrameData_O[14] ;
 wire \Tile_X5Y12_FrameData_O[15] ;
 wire \Tile_X5Y12_FrameData_O[16] ;
 wire \Tile_X5Y12_FrameData_O[17] ;
 wire \Tile_X5Y12_FrameData_O[18] ;
 wire \Tile_X5Y12_FrameData_O[19] ;
 wire \Tile_X5Y12_FrameData_O[1] ;
 wire \Tile_X5Y12_FrameData_O[20] ;
 wire \Tile_X5Y12_FrameData_O[21] ;
 wire \Tile_X5Y12_FrameData_O[22] ;
 wire \Tile_X5Y12_FrameData_O[23] ;
 wire \Tile_X5Y12_FrameData_O[24] ;
 wire \Tile_X5Y12_FrameData_O[25] ;
 wire \Tile_X5Y12_FrameData_O[26] ;
 wire \Tile_X5Y12_FrameData_O[27] ;
 wire \Tile_X5Y12_FrameData_O[28] ;
 wire \Tile_X5Y12_FrameData_O[29] ;
 wire \Tile_X5Y12_FrameData_O[2] ;
 wire \Tile_X5Y12_FrameData_O[30] ;
 wire \Tile_X5Y12_FrameData_O[31] ;
 wire \Tile_X5Y12_FrameData_O[3] ;
 wire \Tile_X5Y12_FrameData_O[4] ;
 wire \Tile_X5Y12_FrameData_O[5] ;
 wire \Tile_X5Y12_FrameData_O[6] ;
 wire \Tile_X5Y12_FrameData_O[7] ;
 wire \Tile_X5Y12_FrameData_O[8] ;
 wire \Tile_X5Y12_FrameData_O[9] ;
 wire \Tile_X5Y12_FrameStrobe_O[0] ;
 wire \Tile_X5Y12_FrameStrobe_O[10] ;
 wire \Tile_X5Y12_FrameStrobe_O[11] ;
 wire \Tile_X5Y12_FrameStrobe_O[12] ;
 wire \Tile_X5Y12_FrameStrobe_O[13] ;
 wire \Tile_X5Y12_FrameStrobe_O[14] ;
 wire \Tile_X5Y12_FrameStrobe_O[15] ;
 wire \Tile_X5Y12_FrameStrobe_O[16] ;
 wire \Tile_X5Y12_FrameStrobe_O[17] ;
 wire \Tile_X5Y12_FrameStrobe_O[18] ;
 wire \Tile_X5Y12_FrameStrobe_O[19] ;
 wire \Tile_X5Y12_FrameStrobe_O[1] ;
 wire \Tile_X5Y12_FrameStrobe_O[2] ;
 wire \Tile_X5Y12_FrameStrobe_O[3] ;
 wire \Tile_X5Y12_FrameStrobe_O[4] ;
 wire \Tile_X5Y12_FrameStrobe_O[5] ;
 wire \Tile_X5Y12_FrameStrobe_O[6] ;
 wire \Tile_X5Y12_FrameStrobe_O[7] ;
 wire \Tile_X5Y12_FrameStrobe_O[8] ;
 wire \Tile_X5Y12_FrameStrobe_O[9] ;
 wire \Tile_X5Y12_N1BEG[0] ;
 wire \Tile_X5Y12_N1BEG[1] ;
 wire \Tile_X5Y12_N1BEG[2] ;
 wire \Tile_X5Y12_N1BEG[3] ;
 wire \Tile_X5Y12_N2BEG[0] ;
 wire \Tile_X5Y12_N2BEG[1] ;
 wire \Tile_X5Y12_N2BEG[2] ;
 wire \Tile_X5Y12_N2BEG[3] ;
 wire \Tile_X5Y12_N2BEG[4] ;
 wire \Tile_X5Y12_N2BEG[5] ;
 wire \Tile_X5Y12_N2BEG[6] ;
 wire \Tile_X5Y12_N2BEG[7] ;
 wire \Tile_X5Y12_N2BEGb[0] ;
 wire \Tile_X5Y12_N2BEGb[1] ;
 wire \Tile_X5Y12_N2BEGb[2] ;
 wire \Tile_X5Y12_N2BEGb[3] ;
 wire \Tile_X5Y12_N2BEGb[4] ;
 wire \Tile_X5Y12_N2BEGb[5] ;
 wire \Tile_X5Y12_N2BEGb[6] ;
 wire \Tile_X5Y12_N2BEGb[7] ;
 wire \Tile_X5Y12_N4BEG[0] ;
 wire \Tile_X5Y12_N4BEG[10] ;
 wire \Tile_X5Y12_N4BEG[11] ;
 wire \Tile_X5Y12_N4BEG[12] ;
 wire \Tile_X5Y12_N4BEG[13] ;
 wire \Tile_X5Y12_N4BEG[14] ;
 wire \Tile_X5Y12_N4BEG[15] ;
 wire \Tile_X5Y12_N4BEG[1] ;
 wire \Tile_X5Y12_N4BEG[2] ;
 wire \Tile_X5Y12_N4BEG[3] ;
 wire \Tile_X5Y12_N4BEG[4] ;
 wire \Tile_X5Y12_N4BEG[5] ;
 wire \Tile_X5Y12_N4BEG[6] ;
 wire \Tile_X5Y12_N4BEG[7] ;
 wire \Tile_X5Y12_N4BEG[8] ;
 wire \Tile_X5Y12_N4BEG[9] ;
 wire \Tile_X5Y12_NN4BEG[0] ;
 wire \Tile_X5Y12_NN4BEG[10] ;
 wire \Tile_X5Y12_NN4BEG[11] ;
 wire \Tile_X5Y12_NN4BEG[12] ;
 wire \Tile_X5Y12_NN4BEG[13] ;
 wire \Tile_X5Y12_NN4BEG[14] ;
 wire \Tile_X5Y12_NN4BEG[15] ;
 wire \Tile_X5Y12_NN4BEG[1] ;
 wire \Tile_X5Y12_NN4BEG[2] ;
 wire \Tile_X5Y12_NN4BEG[3] ;
 wire \Tile_X5Y12_NN4BEG[4] ;
 wire \Tile_X5Y12_NN4BEG[5] ;
 wire \Tile_X5Y12_NN4BEG[6] ;
 wire \Tile_X5Y12_NN4BEG[7] ;
 wire \Tile_X5Y12_NN4BEG[8] ;
 wire \Tile_X5Y12_NN4BEG[9] ;
 wire \Tile_X5Y12_S1BEG[0] ;
 wire \Tile_X5Y12_S1BEG[1] ;
 wire \Tile_X5Y12_S1BEG[2] ;
 wire \Tile_X5Y12_S1BEG[3] ;
 wire \Tile_X5Y12_S2BEG[0] ;
 wire \Tile_X5Y12_S2BEG[1] ;
 wire \Tile_X5Y12_S2BEG[2] ;
 wire \Tile_X5Y12_S2BEG[3] ;
 wire \Tile_X5Y12_S2BEG[4] ;
 wire \Tile_X5Y12_S2BEG[5] ;
 wire \Tile_X5Y12_S2BEG[6] ;
 wire \Tile_X5Y12_S2BEG[7] ;
 wire \Tile_X5Y12_S2BEGb[0] ;
 wire \Tile_X5Y12_S2BEGb[1] ;
 wire \Tile_X5Y12_S2BEGb[2] ;
 wire \Tile_X5Y12_S2BEGb[3] ;
 wire \Tile_X5Y12_S2BEGb[4] ;
 wire \Tile_X5Y12_S2BEGb[5] ;
 wire \Tile_X5Y12_S2BEGb[6] ;
 wire \Tile_X5Y12_S2BEGb[7] ;
 wire \Tile_X5Y12_S4BEG[0] ;
 wire \Tile_X5Y12_S4BEG[10] ;
 wire \Tile_X5Y12_S4BEG[11] ;
 wire \Tile_X5Y12_S4BEG[12] ;
 wire \Tile_X5Y12_S4BEG[13] ;
 wire \Tile_X5Y12_S4BEG[14] ;
 wire \Tile_X5Y12_S4BEG[15] ;
 wire \Tile_X5Y12_S4BEG[1] ;
 wire \Tile_X5Y12_S4BEG[2] ;
 wire \Tile_X5Y12_S4BEG[3] ;
 wire \Tile_X5Y12_S4BEG[4] ;
 wire \Tile_X5Y12_S4BEG[5] ;
 wire \Tile_X5Y12_S4BEG[6] ;
 wire \Tile_X5Y12_S4BEG[7] ;
 wire \Tile_X5Y12_S4BEG[8] ;
 wire \Tile_X5Y12_S4BEG[9] ;
 wire \Tile_X5Y12_SS4BEG[0] ;
 wire \Tile_X5Y12_SS4BEG[10] ;
 wire \Tile_X5Y12_SS4BEG[11] ;
 wire \Tile_X5Y12_SS4BEG[12] ;
 wire \Tile_X5Y12_SS4BEG[13] ;
 wire \Tile_X5Y12_SS4BEG[14] ;
 wire \Tile_X5Y12_SS4BEG[15] ;
 wire \Tile_X5Y12_SS4BEG[1] ;
 wire \Tile_X5Y12_SS4BEG[2] ;
 wire \Tile_X5Y12_SS4BEG[3] ;
 wire \Tile_X5Y12_SS4BEG[4] ;
 wire \Tile_X5Y12_SS4BEG[5] ;
 wire \Tile_X5Y12_SS4BEG[6] ;
 wire \Tile_X5Y12_SS4BEG[7] ;
 wire \Tile_X5Y12_SS4BEG[8] ;
 wire \Tile_X5Y12_SS4BEG[9] ;
 wire Tile_X5Y12_UserCLKo;
 wire \Tile_X5Y12_W1BEG[0] ;
 wire \Tile_X5Y12_W1BEG[1] ;
 wire \Tile_X5Y12_W1BEG[2] ;
 wire \Tile_X5Y12_W1BEG[3] ;
 wire \Tile_X5Y12_W2BEG[0] ;
 wire \Tile_X5Y12_W2BEG[1] ;
 wire \Tile_X5Y12_W2BEG[2] ;
 wire \Tile_X5Y12_W2BEG[3] ;
 wire \Tile_X5Y12_W2BEG[4] ;
 wire \Tile_X5Y12_W2BEG[5] ;
 wire \Tile_X5Y12_W2BEG[6] ;
 wire \Tile_X5Y12_W2BEG[7] ;
 wire \Tile_X5Y12_W2BEGb[0] ;
 wire \Tile_X5Y12_W2BEGb[1] ;
 wire \Tile_X5Y12_W2BEGb[2] ;
 wire \Tile_X5Y12_W2BEGb[3] ;
 wire \Tile_X5Y12_W2BEGb[4] ;
 wire \Tile_X5Y12_W2BEGb[5] ;
 wire \Tile_X5Y12_W2BEGb[6] ;
 wire \Tile_X5Y12_W2BEGb[7] ;
 wire \Tile_X5Y12_W6BEG[0] ;
 wire \Tile_X5Y12_W6BEG[10] ;
 wire \Tile_X5Y12_W6BEG[11] ;
 wire \Tile_X5Y12_W6BEG[1] ;
 wire \Tile_X5Y12_W6BEG[2] ;
 wire \Tile_X5Y12_W6BEG[3] ;
 wire \Tile_X5Y12_W6BEG[4] ;
 wire \Tile_X5Y12_W6BEG[5] ;
 wire \Tile_X5Y12_W6BEG[6] ;
 wire \Tile_X5Y12_W6BEG[7] ;
 wire \Tile_X5Y12_W6BEG[8] ;
 wire \Tile_X5Y12_W6BEG[9] ;
 wire \Tile_X5Y12_WW4BEG[0] ;
 wire \Tile_X5Y12_WW4BEG[10] ;
 wire \Tile_X5Y12_WW4BEG[11] ;
 wire \Tile_X5Y12_WW4BEG[12] ;
 wire \Tile_X5Y12_WW4BEG[13] ;
 wire \Tile_X5Y12_WW4BEG[14] ;
 wire \Tile_X5Y12_WW4BEG[15] ;
 wire \Tile_X5Y12_WW4BEG[1] ;
 wire \Tile_X5Y12_WW4BEG[2] ;
 wire \Tile_X5Y12_WW4BEG[3] ;
 wire \Tile_X5Y12_WW4BEG[4] ;
 wire \Tile_X5Y12_WW4BEG[5] ;
 wire \Tile_X5Y12_WW4BEG[6] ;
 wire \Tile_X5Y12_WW4BEG[7] ;
 wire \Tile_X5Y12_WW4BEG[8] ;
 wire \Tile_X5Y12_WW4BEG[9] ;
 wire Tile_X5Y13_Co;
 wire \Tile_X5Y13_E1BEG[0] ;
 wire \Tile_X5Y13_E1BEG[1] ;
 wire \Tile_X5Y13_E1BEG[2] ;
 wire \Tile_X5Y13_E1BEG[3] ;
 wire \Tile_X5Y13_E2BEG[0] ;
 wire \Tile_X5Y13_E2BEG[1] ;
 wire \Tile_X5Y13_E2BEG[2] ;
 wire \Tile_X5Y13_E2BEG[3] ;
 wire \Tile_X5Y13_E2BEG[4] ;
 wire \Tile_X5Y13_E2BEG[5] ;
 wire \Tile_X5Y13_E2BEG[6] ;
 wire \Tile_X5Y13_E2BEG[7] ;
 wire \Tile_X5Y13_E2BEGb[0] ;
 wire \Tile_X5Y13_E2BEGb[1] ;
 wire \Tile_X5Y13_E2BEGb[2] ;
 wire \Tile_X5Y13_E2BEGb[3] ;
 wire \Tile_X5Y13_E2BEGb[4] ;
 wire \Tile_X5Y13_E2BEGb[5] ;
 wire \Tile_X5Y13_E2BEGb[6] ;
 wire \Tile_X5Y13_E2BEGb[7] ;
 wire \Tile_X5Y13_E6BEG[0] ;
 wire \Tile_X5Y13_E6BEG[10] ;
 wire \Tile_X5Y13_E6BEG[11] ;
 wire \Tile_X5Y13_E6BEG[1] ;
 wire \Tile_X5Y13_E6BEG[2] ;
 wire \Tile_X5Y13_E6BEG[3] ;
 wire \Tile_X5Y13_E6BEG[4] ;
 wire \Tile_X5Y13_E6BEG[5] ;
 wire \Tile_X5Y13_E6BEG[6] ;
 wire \Tile_X5Y13_E6BEG[7] ;
 wire \Tile_X5Y13_E6BEG[8] ;
 wire \Tile_X5Y13_E6BEG[9] ;
 wire \Tile_X5Y13_EE4BEG[0] ;
 wire \Tile_X5Y13_EE4BEG[10] ;
 wire \Tile_X5Y13_EE4BEG[11] ;
 wire \Tile_X5Y13_EE4BEG[12] ;
 wire \Tile_X5Y13_EE4BEG[13] ;
 wire \Tile_X5Y13_EE4BEG[14] ;
 wire \Tile_X5Y13_EE4BEG[15] ;
 wire \Tile_X5Y13_EE4BEG[1] ;
 wire \Tile_X5Y13_EE4BEG[2] ;
 wire \Tile_X5Y13_EE4BEG[3] ;
 wire \Tile_X5Y13_EE4BEG[4] ;
 wire \Tile_X5Y13_EE4BEG[5] ;
 wire \Tile_X5Y13_EE4BEG[6] ;
 wire \Tile_X5Y13_EE4BEG[7] ;
 wire \Tile_X5Y13_EE4BEG[8] ;
 wire \Tile_X5Y13_EE4BEG[9] ;
 wire \Tile_X5Y13_FrameData_O[0] ;
 wire \Tile_X5Y13_FrameData_O[10] ;
 wire \Tile_X5Y13_FrameData_O[11] ;
 wire \Tile_X5Y13_FrameData_O[12] ;
 wire \Tile_X5Y13_FrameData_O[13] ;
 wire \Tile_X5Y13_FrameData_O[14] ;
 wire \Tile_X5Y13_FrameData_O[15] ;
 wire \Tile_X5Y13_FrameData_O[16] ;
 wire \Tile_X5Y13_FrameData_O[17] ;
 wire \Tile_X5Y13_FrameData_O[18] ;
 wire \Tile_X5Y13_FrameData_O[19] ;
 wire \Tile_X5Y13_FrameData_O[1] ;
 wire \Tile_X5Y13_FrameData_O[20] ;
 wire \Tile_X5Y13_FrameData_O[21] ;
 wire \Tile_X5Y13_FrameData_O[22] ;
 wire \Tile_X5Y13_FrameData_O[23] ;
 wire \Tile_X5Y13_FrameData_O[24] ;
 wire \Tile_X5Y13_FrameData_O[25] ;
 wire \Tile_X5Y13_FrameData_O[26] ;
 wire \Tile_X5Y13_FrameData_O[27] ;
 wire \Tile_X5Y13_FrameData_O[28] ;
 wire \Tile_X5Y13_FrameData_O[29] ;
 wire \Tile_X5Y13_FrameData_O[2] ;
 wire \Tile_X5Y13_FrameData_O[30] ;
 wire \Tile_X5Y13_FrameData_O[31] ;
 wire \Tile_X5Y13_FrameData_O[3] ;
 wire \Tile_X5Y13_FrameData_O[4] ;
 wire \Tile_X5Y13_FrameData_O[5] ;
 wire \Tile_X5Y13_FrameData_O[6] ;
 wire \Tile_X5Y13_FrameData_O[7] ;
 wire \Tile_X5Y13_FrameData_O[8] ;
 wire \Tile_X5Y13_FrameData_O[9] ;
 wire \Tile_X5Y13_FrameStrobe_O[0] ;
 wire \Tile_X5Y13_FrameStrobe_O[10] ;
 wire \Tile_X5Y13_FrameStrobe_O[11] ;
 wire \Tile_X5Y13_FrameStrobe_O[12] ;
 wire \Tile_X5Y13_FrameStrobe_O[13] ;
 wire \Tile_X5Y13_FrameStrobe_O[14] ;
 wire \Tile_X5Y13_FrameStrobe_O[15] ;
 wire \Tile_X5Y13_FrameStrobe_O[16] ;
 wire \Tile_X5Y13_FrameStrobe_O[17] ;
 wire \Tile_X5Y13_FrameStrobe_O[18] ;
 wire \Tile_X5Y13_FrameStrobe_O[19] ;
 wire \Tile_X5Y13_FrameStrobe_O[1] ;
 wire \Tile_X5Y13_FrameStrobe_O[2] ;
 wire \Tile_X5Y13_FrameStrobe_O[3] ;
 wire \Tile_X5Y13_FrameStrobe_O[4] ;
 wire \Tile_X5Y13_FrameStrobe_O[5] ;
 wire \Tile_X5Y13_FrameStrobe_O[6] ;
 wire \Tile_X5Y13_FrameStrobe_O[7] ;
 wire \Tile_X5Y13_FrameStrobe_O[8] ;
 wire \Tile_X5Y13_FrameStrobe_O[9] ;
 wire \Tile_X5Y13_N1BEG[0] ;
 wire \Tile_X5Y13_N1BEG[1] ;
 wire \Tile_X5Y13_N1BEG[2] ;
 wire \Tile_X5Y13_N1BEG[3] ;
 wire \Tile_X5Y13_N2BEG[0] ;
 wire \Tile_X5Y13_N2BEG[1] ;
 wire \Tile_X5Y13_N2BEG[2] ;
 wire \Tile_X5Y13_N2BEG[3] ;
 wire \Tile_X5Y13_N2BEG[4] ;
 wire \Tile_X5Y13_N2BEG[5] ;
 wire \Tile_X5Y13_N2BEG[6] ;
 wire \Tile_X5Y13_N2BEG[7] ;
 wire \Tile_X5Y13_N2BEGb[0] ;
 wire \Tile_X5Y13_N2BEGb[1] ;
 wire \Tile_X5Y13_N2BEGb[2] ;
 wire \Tile_X5Y13_N2BEGb[3] ;
 wire \Tile_X5Y13_N2BEGb[4] ;
 wire \Tile_X5Y13_N2BEGb[5] ;
 wire \Tile_X5Y13_N2BEGb[6] ;
 wire \Tile_X5Y13_N2BEGb[7] ;
 wire \Tile_X5Y13_N4BEG[0] ;
 wire \Tile_X5Y13_N4BEG[10] ;
 wire \Tile_X5Y13_N4BEG[11] ;
 wire \Tile_X5Y13_N4BEG[12] ;
 wire \Tile_X5Y13_N4BEG[13] ;
 wire \Tile_X5Y13_N4BEG[14] ;
 wire \Tile_X5Y13_N4BEG[15] ;
 wire \Tile_X5Y13_N4BEG[1] ;
 wire \Tile_X5Y13_N4BEG[2] ;
 wire \Tile_X5Y13_N4BEG[3] ;
 wire \Tile_X5Y13_N4BEG[4] ;
 wire \Tile_X5Y13_N4BEG[5] ;
 wire \Tile_X5Y13_N4BEG[6] ;
 wire \Tile_X5Y13_N4BEG[7] ;
 wire \Tile_X5Y13_N4BEG[8] ;
 wire \Tile_X5Y13_N4BEG[9] ;
 wire \Tile_X5Y13_NN4BEG[0] ;
 wire \Tile_X5Y13_NN4BEG[10] ;
 wire \Tile_X5Y13_NN4BEG[11] ;
 wire \Tile_X5Y13_NN4BEG[12] ;
 wire \Tile_X5Y13_NN4BEG[13] ;
 wire \Tile_X5Y13_NN4BEG[14] ;
 wire \Tile_X5Y13_NN4BEG[15] ;
 wire \Tile_X5Y13_NN4BEG[1] ;
 wire \Tile_X5Y13_NN4BEG[2] ;
 wire \Tile_X5Y13_NN4BEG[3] ;
 wire \Tile_X5Y13_NN4BEG[4] ;
 wire \Tile_X5Y13_NN4BEG[5] ;
 wire \Tile_X5Y13_NN4BEG[6] ;
 wire \Tile_X5Y13_NN4BEG[7] ;
 wire \Tile_X5Y13_NN4BEG[8] ;
 wire \Tile_X5Y13_NN4BEG[9] ;
 wire \Tile_X5Y13_S1BEG[0] ;
 wire \Tile_X5Y13_S1BEG[1] ;
 wire \Tile_X5Y13_S1BEG[2] ;
 wire \Tile_X5Y13_S1BEG[3] ;
 wire \Tile_X5Y13_S2BEG[0] ;
 wire \Tile_X5Y13_S2BEG[1] ;
 wire \Tile_X5Y13_S2BEG[2] ;
 wire \Tile_X5Y13_S2BEG[3] ;
 wire \Tile_X5Y13_S2BEG[4] ;
 wire \Tile_X5Y13_S2BEG[5] ;
 wire \Tile_X5Y13_S2BEG[6] ;
 wire \Tile_X5Y13_S2BEG[7] ;
 wire \Tile_X5Y13_S2BEGb[0] ;
 wire \Tile_X5Y13_S2BEGb[1] ;
 wire \Tile_X5Y13_S2BEGb[2] ;
 wire \Tile_X5Y13_S2BEGb[3] ;
 wire \Tile_X5Y13_S2BEGb[4] ;
 wire \Tile_X5Y13_S2BEGb[5] ;
 wire \Tile_X5Y13_S2BEGb[6] ;
 wire \Tile_X5Y13_S2BEGb[7] ;
 wire \Tile_X5Y13_S4BEG[0] ;
 wire \Tile_X5Y13_S4BEG[10] ;
 wire \Tile_X5Y13_S4BEG[11] ;
 wire \Tile_X5Y13_S4BEG[12] ;
 wire \Tile_X5Y13_S4BEG[13] ;
 wire \Tile_X5Y13_S4BEG[14] ;
 wire \Tile_X5Y13_S4BEG[15] ;
 wire \Tile_X5Y13_S4BEG[1] ;
 wire \Tile_X5Y13_S4BEG[2] ;
 wire \Tile_X5Y13_S4BEG[3] ;
 wire \Tile_X5Y13_S4BEG[4] ;
 wire \Tile_X5Y13_S4BEG[5] ;
 wire \Tile_X5Y13_S4BEG[6] ;
 wire \Tile_X5Y13_S4BEG[7] ;
 wire \Tile_X5Y13_S4BEG[8] ;
 wire \Tile_X5Y13_S4BEG[9] ;
 wire \Tile_X5Y13_SS4BEG[0] ;
 wire \Tile_X5Y13_SS4BEG[10] ;
 wire \Tile_X5Y13_SS4BEG[11] ;
 wire \Tile_X5Y13_SS4BEG[12] ;
 wire \Tile_X5Y13_SS4BEG[13] ;
 wire \Tile_X5Y13_SS4BEG[14] ;
 wire \Tile_X5Y13_SS4BEG[15] ;
 wire \Tile_X5Y13_SS4BEG[1] ;
 wire \Tile_X5Y13_SS4BEG[2] ;
 wire \Tile_X5Y13_SS4BEG[3] ;
 wire \Tile_X5Y13_SS4BEG[4] ;
 wire \Tile_X5Y13_SS4BEG[5] ;
 wire \Tile_X5Y13_SS4BEG[6] ;
 wire \Tile_X5Y13_SS4BEG[7] ;
 wire \Tile_X5Y13_SS4BEG[8] ;
 wire \Tile_X5Y13_SS4BEG[9] ;
 wire Tile_X5Y13_UserCLKo;
 wire \Tile_X5Y13_W1BEG[0] ;
 wire \Tile_X5Y13_W1BEG[1] ;
 wire \Tile_X5Y13_W1BEG[2] ;
 wire \Tile_X5Y13_W1BEG[3] ;
 wire \Tile_X5Y13_W2BEG[0] ;
 wire \Tile_X5Y13_W2BEG[1] ;
 wire \Tile_X5Y13_W2BEG[2] ;
 wire \Tile_X5Y13_W2BEG[3] ;
 wire \Tile_X5Y13_W2BEG[4] ;
 wire \Tile_X5Y13_W2BEG[5] ;
 wire \Tile_X5Y13_W2BEG[6] ;
 wire \Tile_X5Y13_W2BEG[7] ;
 wire \Tile_X5Y13_W2BEGb[0] ;
 wire \Tile_X5Y13_W2BEGb[1] ;
 wire \Tile_X5Y13_W2BEGb[2] ;
 wire \Tile_X5Y13_W2BEGb[3] ;
 wire \Tile_X5Y13_W2BEGb[4] ;
 wire \Tile_X5Y13_W2BEGb[5] ;
 wire \Tile_X5Y13_W2BEGb[6] ;
 wire \Tile_X5Y13_W2BEGb[7] ;
 wire \Tile_X5Y13_W6BEG[0] ;
 wire \Tile_X5Y13_W6BEG[10] ;
 wire \Tile_X5Y13_W6BEG[11] ;
 wire \Tile_X5Y13_W6BEG[1] ;
 wire \Tile_X5Y13_W6BEG[2] ;
 wire \Tile_X5Y13_W6BEG[3] ;
 wire \Tile_X5Y13_W6BEG[4] ;
 wire \Tile_X5Y13_W6BEG[5] ;
 wire \Tile_X5Y13_W6BEG[6] ;
 wire \Tile_X5Y13_W6BEG[7] ;
 wire \Tile_X5Y13_W6BEG[8] ;
 wire \Tile_X5Y13_W6BEG[9] ;
 wire \Tile_X5Y13_WW4BEG[0] ;
 wire \Tile_X5Y13_WW4BEG[10] ;
 wire \Tile_X5Y13_WW4BEG[11] ;
 wire \Tile_X5Y13_WW4BEG[12] ;
 wire \Tile_X5Y13_WW4BEG[13] ;
 wire \Tile_X5Y13_WW4BEG[14] ;
 wire \Tile_X5Y13_WW4BEG[15] ;
 wire \Tile_X5Y13_WW4BEG[1] ;
 wire \Tile_X5Y13_WW4BEG[2] ;
 wire \Tile_X5Y13_WW4BEG[3] ;
 wire \Tile_X5Y13_WW4BEG[4] ;
 wire \Tile_X5Y13_WW4BEG[5] ;
 wire \Tile_X5Y13_WW4BEG[6] ;
 wire \Tile_X5Y13_WW4BEG[7] ;
 wire \Tile_X5Y13_WW4BEG[8] ;
 wire \Tile_X5Y13_WW4BEG[9] ;
 wire Tile_X5Y14_Co;
 wire \Tile_X5Y14_E1BEG[0] ;
 wire \Tile_X5Y14_E1BEG[1] ;
 wire \Tile_X5Y14_E1BEG[2] ;
 wire \Tile_X5Y14_E1BEG[3] ;
 wire \Tile_X5Y14_E2BEG[0] ;
 wire \Tile_X5Y14_E2BEG[1] ;
 wire \Tile_X5Y14_E2BEG[2] ;
 wire \Tile_X5Y14_E2BEG[3] ;
 wire \Tile_X5Y14_E2BEG[4] ;
 wire \Tile_X5Y14_E2BEG[5] ;
 wire \Tile_X5Y14_E2BEG[6] ;
 wire \Tile_X5Y14_E2BEG[7] ;
 wire \Tile_X5Y14_E2BEGb[0] ;
 wire \Tile_X5Y14_E2BEGb[1] ;
 wire \Tile_X5Y14_E2BEGb[2] ;
 wire \Tile_X5Y14_E2BEGb[3] ;
 wire \Tile_X5Y14_E2BEGb[4] ;
 wire \Tile_X5Y14_E2BEGb[5] ;
 wire \Tile_X5Y14_E2BEGb[6] ;
 wire \Tile_X5Y14_E2BEGb[7] ;
 wire \Tile_X5Y14_E6BEG[0] ;
 wire \Tile_X5Y14_E6BEG[10] ;
 wire \Tile_X5Y14_E6BEG[11] ;
 wire \Tile_X5Y14_E6BEG[1] ;
 wire \Tile_X5Y14_E6BEG[2] ;
 wire \Tile_X5Y14_E6BEG[3] ;
 wire \Tile_X5Y14_E6BEG[4] ;
 wire \Tile_X5Y14_E6BEG[5] ;
 wire \Tile_X5Y14_E6BEG[6] ;
 wire \Tile_X5Y14_E6BEG[7] ;
 wire \Tile_X5Y14_E6BEG[8] ;
 wire \Tile_X5Y14_E6BEG[9] ;
 wire \Tile_X5Y14_EE4BEG[0] ;
 wire \Tile_X5Y14_EE4BEG[10] ;
 wire \Tile_X5Y14_EE4BEG[11] ;
 wire \Tile_X5Y14_EE4BEG[12] ;
 wire \Tile_X5Y14_EE4BEG[13] ;
 wire \Tile_X5Y14_EE4BEG[14] ;
 wire \Tile_X5Y14_EE4BEG[15] ;
 wire \Tile_X5Y14_EE4BEG[1] ;
 wire \Tile_X5Y14_EE4BEG[2] ;
 wire \Tile_X5Y14_EE4BEG[3] ;
 wire \Tile_X5Y14_EE4BEG[4] ;
 wire \Tile_X5Y14_EE4BEG[5] ;
 wire \Tile_X5Y14_EE4BEG[6] ;
 wire \Tile_X5Y14_EE4BEG[7] ;
 wire \Tile_X5Y14_EE4BEG[8] ;
 wire \Tile_X5Y14_EE4BEG[9] ;
 wire \Tile_X5Y14_FrameData_O[0] ;
 wire \Tile_X5Y14_FrameData_O[10] ;
 wire \Tile_X5Y14_FrameData_O[11] ;
 wire \Tile_X5Y14_FrameData_O[12] ;
 wire \Tile_X5Y14_FrameData_O[13] ;
 wire \Tile_X5Y14_FrameData_O[14] ;
 wire \Tile_X5Y14_FrameData_O[15] ;
 wire \Tile_X5Y14_FrameData_O[16] ;
 wire \Tile_X5Y14_FrameData_O[17] ;
 wire \Tile_X5Y14_FrameData_O[18] ;
 wire \Tile_X5Y14_FrameData_O[19] ;
 wire \Tile_X5Y14_FrameData_O[1] ;
 wire \Tile_X5Y14_FrameData_O[20] ;
 wire \Tile_X5Y14_FrameData_O[21] ;
 wire \Tile_X5Y14_FrameData_O[22] ;
 wire \Tile_X5Y14_FrameData_O[23] ;
 wire \Tile_X5Y14_FrameData_O[24] ;
 wire \Tile_X5Y14_FrameData_O[25] ;
 wire \Tile_X5Y14_FrameData_O[26] ;
 wire \Tile_X5Y14_FrameData_O[27] ;
 wire \Tile_X5Y14_FrameData_O[28] ;
 wire \Tile_X5Y14_FrameData_O[29] ;
 wire \Tile_X5Y14_FrameData_O[2] ;
 wire \Tile_X5Y14_FrameData_O[30] ;
 wire \Tile_X5Y14_FrameData_O[31] ;
 wire \Tile_X5Y14_FrameData_O[3] ;
 wire \Tile_X5Y14_FrameData_O[4] ;
 wire \Tile_X5Y14_FrameData_O[5] ;
 wire \Tile_X5Y14_FrameData_O[6] ;
 wire \Tile_X5Y14_FrameData_O[7] ;
 wire \Tile_X5Y14_FrameData_O[8] ;
 wire \Tile_X5Y14_FrameData_O[9] ;
 wire \Tile_X5Y14_FrameStrobe_O[0] ;
 wire \Tile_X5Y14_FrameStrobe_O[10] ;
 wire \Tile_X5Y14_FrameStrobe_O[11] ;
 wire \Tile_X5Y14_FrameStrobe_O[12] ;
 wire \Tile_X5Y14_FrameStrobe_O[13] ;
 wire \Tile_X5Y14_FrameStrobe_O[14] ;
 wire \Tile_X5Y14_FrameStrobe_O[15] ;
 wire \Tile_X5Y14_FrameStrobe_O[16] ;
 wire \Tile_X5Y14_FrameStrobe_O[17] ;
 wire \Tile_X5Y14_FrameStrobe_O[18] ;
 wire \Tile_X5Y14_FrameStrobe_O[19] ;
 wire \Tile_X5Y14_FrameStrobe_O[1] ;
 wire \Tile_X5Y14_FrameStrobe_O[2] ;
 wire \Tile_X5Y14_FrameStrobe_O[3] ;
 wire \Tile_X5Y14_FrameStrobe_O[4] ;
 wire \Tile_X5Y14_FrameStrobe_O[5] ;
 wire \Tile_X5Y14_FrameStrobe_O[6] ;
 wire \Tile_X5Y14_FrameStrobe_O[7] ;
 wire \Tile_X5Y14_FrameStrobe_O[8] ;
 wire \Tile_X5Y14_FrameStrobe_O[9] ;
 wire \Tile_X5Y14_N1BEG[0] ;
 wire \Tile_X5Y14_N1BEG[1] ;
 wire \Tile_X5Y14_N1BEG[2] ;
 wire \Tile_X5Y14_N1BEG[3] ;
 wire \Tile_X5Y14_N2BEG[0] ;
 wire \Tile_X5Y14_N2BEG[1] ;
 wire \Tile_X5Y14_N2BEG[2] ;
 wire \Tile_X5Y14_N2BEG[3] ;
 wire \Tile_X5Y14_N2BEG[4] ;
 wire \Tile_X5Y14_N2BEG[5] ;
 wire \Tile_X5Y14_N2BEG[6] ;
 wire \Tile_X5Y14_N2BEG[7] ;
 wire \Tile_X5Y14_N2BEGb[0] ;
 wire \Tile_X5Y14_N2BEGb[1] ;
 wire \Tile_X5Y14_N2BEGb[2] ;
 wire \Tile_X5Y14_N2BEGb[3] ;
 wire \Tile_X5Y14_N2BEGb[4] ;
 wire \Tile_X5Y14_N2BEGb[5] ;
 wire \Tile_X5Y14_N2BEGb[6] ;
 wire \Tile_X5Y14_N2BEGb[7] ;
 wire \Tile_X5Y14_N4BEG[0] ;
 wire \Tile_X5Y14_N4BEG[10] ;
 wire \Tile_X5Y14_N4BEG[11] ;
 wire \Tile_X5Y14_N4BEG[12] ;
 wire \Tile_X5Y14_N4BEG[13] ;
 wire \Tile_X5Y14_N4BEG[14] ;
 wire \Tile_X5Y14_N4BEG[15] ;
 wire \Tile_X5Y14_N4BEG[1] ;
 wire \Tile_X5Y14_N4BEG[2] ;
 wire \Tile_X5Y14_N4BEG[3] ;
 wire \Tile_X5Y14_N4BEG[4] ;
 wire \Tile_X5Y14_N4BEG[5] ;
 wire \Tile_X5Y14_N4BEG[6] ;
 wire \Tile_X5Y14_N4BEG[7] ;
 wire \Tile_X5Y14_N4BEG[8] ;
 wire \Tile_X5Y14_N4BEG[9] ;
 wire \Tile_X5Y14_NN4BEG[0] ;
 wire \Tile_X5Y14_NN4BEG[10] ;
 wire \Tile_X5Y14_NN4BEG[11] ;
 wire \Tile_X5Y14_NN4BEG[12] ;
 wire \Tile_X5Y14_NN4BEG[13] ;
 wire \Tile_X5Y14_NN4BEG[14] ;
 wire \Tile_X5Y14_NN4BEG[15] ;
 wire \Tile_X5Y14_NN4BEG[1] ;
 wire \Tile_X5Y14_NN4BEG[2] ;
 wire \Tile_X5Y14_NN4BEG[3] ;
 wire \Tile_X5Y14_NN4BEG[4] ;
 wire \Tile_X5Y14_NN4BEG[5] ;
 wire \Tile_X5Y14_NN4BEG[6] ;
 wire \Tile_X5Y14_NN4BEG[7] ;
 wire \Tile_X5Y14_NN4BEG[8] ;
 wire \Tile_X5Y14_NN4BEG[9] ;
 wire \Tile_X5Y14_S1BEG[0] ;
 wire \Tile_X5Y14_S1BEG[1] ;
 wire \Tile_X5Y14_S1BEG[2] ;
 wire \Tile_X5Y14_S1BEG[3] ;
 wire \Tile_X5Y14_S2BEG[0] ;
 wire \Tile_X5Y14_S2BEG[1] ;
 wire \Tile_X5Y14_S2BEG[2] ;
 wire \Tile_X5Y14_S2BEG[3] ;
 wire \Tile_X5Y14_S2BEG[4] ;
 wire \Tile_X5Y14_S2BEG[5] ;
 wire \Tile_X5Y14_S2BEG[6] ;
 wire \Tile_X5Y14_S2BEG[7] ;
 wire \Tile_X5Y14_S2BEGb[0] ;
 wire \Tile_X5Y14_S2BEGb[1] ;
 wire \Tile_X5Y14_S2BEGb[2] ;
 wire \Tile_X5Y14_S2BEGb[3] ;
 wire \Tile_X5Y14_S2BEGb[4] ;
 wire \Tile_X5Y14_S2BEGb[5] ;
 wire \Tile_X5Y14_S2BEGb[6] ;
 wire \Tile_X5Y14_S2BEGb[7] ;
 wire \Tile_X5Y14_S4BEG[0] ;
 wire \Tile_X5Y14_S4BEG[10] ;
 wire \Tile_X5Y14_S4BEG[11] ;
 wire \Tile_X5Y14_S4BEG[12] ;
 wire \Tile_X5Y14_S4BEG[13] ;
 wire \Tile_X5Y14_S4BEG[14] ;
 wire \Tile_X5Y14_S4BEG[15] ;
 wire \Tile_X5Y14_S4BEG[1] ;
 wire \Tile_X5Y14_S4BEG[2] ;
 wire \Tile_X5Y14_S4BEG[3] ;
 wire \Tile_X5Y14_S4BEG[4] ;
 wire \Tile_X5Y14_S4BEG[5] ;
 wire \Tile_X5Y14_S4BEG[6] ;
 wire \Tile_X5Y14_S4BEG[7] ;
 wire \Tile_X5Y14_S4BEG[8] ;
 wire \Tile_X5Y14_S4BEG[9] ;
 wire \Tile_X5Y14_SS4BEG[0] ;
 wire \Tile_X5Y14_SS4BEG[10] ;
 wire \Tile_X5Y14_SS4BEG[11] ;
 wire \Tile_X5Y14_SS4BEG[12] ;
 wire \Tile_X5Y14_SS4BEG[13] ;
 wire \Tile_X5Y14_SS4BEG[14] ;
 wire \Tile_X5Y14_SS4BEG[15] ;
 wire \Tile_X5Y14_SS4BEG[1] ;
 wire \Tile_X5Y14_SS4BEG[2] ;
 wire \Tile_X5Y14_SS4BEG[3] ;
 wire \Tile_X5Y14_SS4BEG[4] ;
 wire \Tile_X5Y14_SS4BEG[5] ;
 wire \Tile_X5Y14_SS4BEG[6] ;
 wire \Tile_X5Y14_SS4BEG[7] ;
 wire \Tile_X5Y14_SS4BEG[8] ;
 wire \Tile_X5Y14_SS4BEG[9] ;
 wire Tile_X5Y14_UserCLKo;
 wire \Tile_X5Y14_W1BEG[0] ;
 wire \Tile_X5Y14_W1BEG[1] ;
 wire \Tile_X5Y14_W1BEG[2] ;
 wire \Tile_X5Y14_W1BEG[3] ;
 wire \Tile_X5Y14_W2BEG[0] ;
 wire \Tile_X5Y14_W2BEG[1] ;
 wire \Tile_X5Y14_W2BEG[2] ;
 wire \Tile_X5Y14_W2BEG[3] ;
 wire \Tile_X5Y14_W2BEG[4] ;
 wire \Tile_X5Y14_W2BEG[5] ;
 wire \Tile_X5Y14_W2BEG[6] ;
 wire \Tile_X5Y14_W2BEG[7] ;
 wire \Tile_X5Y14_W2BEGb[0] ;
 wire \Tile_X5Y14_W2BEGb[1] ;
 wire \Tile_X5Y14_W2BEGb[2] ;
 wire \Tile_X5Y14_W2BEGb[3] ;
 wire \Tile_X5Y14_W2BEGb[4] ;
 wire \Tile_X5Y14_W2BEGb[5] ;
 wire \Tile_X5Y14_W2BEGb[6] ;
 wire \Tile_X5Y14_W2BEGb[7] ;
 wire \Tile_X5Y14_W6BEG[0] ;
 wire \Tile_X5Y14_W6BEG[10] ;
 wire \Tile_X5Y14_W6BEG[11] ;
 wire \Tile_X5Y14_W6BEG[1] ;
 wire \Tile_X5Y14_W6BEG[2] ;
 wire \Tile_X5Y14_W6BEG[3] ;
 wire \Tile_X5Y14_W6BEG[4] ;
 wire \Tile_X5Y14_W6BEG[5] ;
 wire \Tile_X5Y14_W6BEG[6] ;
 wire \Tile_X5Y14_W6BEG[7] ;
 wire \Tile_X5Y14_W6BEG[8] ;
 wire \Tile_X5Y14_W6BEG[9] ;
 wire \Tile_X5Y14_WW4BEG[0] ;
 wire \Tile_X5Y14_WW4BEG[10] ;
 wire \Tile_X5Y14_WW4BEG[11] ;
 wire \Tile_X5Y14_WW4BEG[12] ;
 wire \Tile_X5Y14_WW4BEG[13] ;
 wire \Tile_X5Y14_WW4BEG[14] ;
 wire \Tile_X5Y14_WW4BEG[15] ;
 wire \Tile_X5Y14_WW4BEG[1] ;
 wire \Tile_X5Y14_WW4BEG[2] ;
 wire \Tile_X5Y14_WW4BEG[3] ;
 wire \Tile_X5Y14_WW4BEG[4] ;
 wire \Tile_X5Y14_WW4BEG[5] ;
 wire \Tile_X5Y14_WW4BEG[6] ;
 wire \Tile_X5Y14_WW4BEG[7] ;
 wire \Tile_X5Y14_WW4BEG[8] ;
 wire \Tile_X5Y14_WW4BEG[9] ;
 wire Tile_X5Y15_Co;
 wire \Tile_X5Y15_FrameData_O[0] ;
 wire \Tile_X5Y15_FrameData_O[10] ;
 wire \Tile_X5Y15_FrameData_O[11] ;
 wire \Tile_X5Y15_FrameData_O[12] ;
 wire \Tile_X5Y15_FrameData_O[13] ;
 wire \Tile_X5Y15_FrameData_O[14] ;
 wire \Tile_X5Y15_FrameData_O[15] ;
 wire \Tile_X5Y15_FrameData_O[16] ;
 wire \Tile_X5Y15_FrameData_O[17] ;
 wire \Tile_X5Y15_FrameData_O[18] ;
 wire \Tile_X5Y15_FrameData_O[19] ;
 wire \Tile_X5Y15_FrameData_O[1] ;
 wire \Tile_X5Y15_FrameData_O[20] ;
 wire \Tile_X5Y15_FrameData_O[21] ;
 wire \Tile_X5Y15_FrameData_O[22] ;
 wire \Tile_X5Y15_FrameData_O[23] ;
 wire \Tile_X5Y15_FrameData_O[24] ;
 wire \Tile_X5Y15_FrameData_O[25] ;
 wire \Tile_X5Y15_FrameData_O[26] ;
 wire \Tile_X5Y15_FrameData_O[27] ;
 wire \Tile_X5Y15_FrameData_O[28] ;
 wire \Tile_X5Y15_FrameData_O[29] ;
 wire \Tile_X5Y15_FrameData_O[2] ;
 wire \Tile_X5Y15_FrameData_O[30] ;
 wire \Tile_X5Y15_FrameData_O[31] ;
 wire \Tile_X5Y15_FrameData_O[3] ;
 wire \Tile_X5Y15_FrameData_O[4] ;
 wire \Tile_X5Y15_FrameData_O[5] ;
 wire \Tile_X5Y15_FrameData_O[6] ;
 wire \Tile_X5Y15_FrameData_O[7] ;
 wire \Tile_X5Y15_FrameData_O[8] ;
 wire \Tile_X5Y15_FrameData_O[9] ;
 wire \Tile_X5Y15_FrameStrobe_O[0] ;
 wire \Tile_X5Y15_FrameStrobe_O[10] ;
 wire \Tile_X5Y15_FrameStrobe_O[11] ;
 wire \Tile_X5Y15_FrameStrobe_O[12] ;
 wire \Tile_X5Y15_FrameStrobe_O[13] ;
 wire \Tile_X5Y15_FrameStrobe_O[14] ;
 wire \Tile_X5Y15_FrameStrobe_O[15] ;
 wire \Tile_X5Y15_FrameStrobe_O[16] ;
 wire \Tile_X5Y15_FrameStrobe_O[17] ;
 wire \Tile_X5Y15_FrameStrobe_O[18] ;
 wire \Tile_X5Y15_FrameStrobe_O[19] ;
 wire \Tile_X5Y15_FrameStrobe_O[1] ;
 wire \Tile_X5Y15_FrameStrobe_O[2] ;
 wire \Tile_X5Y15_FrameStrobe_O[3] ;
 wire \Tile_X5Y15_FrameStrobe_O[4] ;
 wire \Tile_X5Y15_FrameStrobe_O[5] ;
 wire \Tile_X5Y15_FrameStrobe_O[6] ;
 wire \Tile_X5Y15_FrameStrobe_O[7] ;
 wire \Tile_X5Y15_FrameStrobe_O[8] ;
 wire \Tile_X5Y15_FrameStrobe_O[9] ;
 wire \Tile_X5Y15_N1BEG[0] ;
 wire \Tile_X5Y15_N1BEG[1] ;
 wire \Tile_X5Y15_N1BEG[2] ;
 wire \Tile_X5Y15_N1BEG[3] ;
 wire \Tile_X5Y15_N2BEG[0] ;
 wire \Tile_X5Y15_N2BEG[1] ;
 wire \Tile_X5Y15_N2BEG[2] ;
 wire \Tile_X5Y15_N2BEG[3] ;
 wire \Tile_X5Y15_N2BEG[4] ;
 wire \Tile_X5Y15_N2BEG[5] ;
 wire \Tile_X5Y15_N2BEG[6] ;
 wire \Tile_X5Y15_N2BEG[7] ;
 wire \Tile_X5Y15_N2BEGb[0] ;
 wire \Tile_X5Y15_N2BEGb[1] ;
 wire \Tile_X5Y15_N2BEGb[2] ;
 wire \Tile_X5Y15_N2BEGb[3] ;
 wire \Tile_X5Y15_N2BEGb[4] ;
 wire \Tile_X5Y15_N2BEGb[5] ;
 wire \Tile_X5Y15_N2BEGb[6] ;
 wire \Tile_X5Y15_N2BEGb[7] ;
 wire \Tile_X5Y15_N4BEG[0] ;
 wire \Tile_X5Y15_N4BEG[10] ;
 wire \Tile_X5Y15_N4BEG[11] ;
 wire \Tile_X5Y15_N4BEG[12] ;
 wire \Tile_X5Y15_N4BEG[13] ;
 wire \Tile_X5Y15_N4BEG[14] ;
 wire \Tile_X5Y15_N4BEG[15] ;
 wire \Tile_X5Y15_N4BEG[1] ;
 wire \Tile_X5Y15_N4BEG[2] ;
 wire \Tile_X5Y15_N4BEG[3] ;
 wire \Tile_X5Y15_N4BEG[4] ;
 wire \Tile_X5Y15_N4BEG[5] ;
 wire \Tile_X5Y15_N4BEG[6] ;
 wire \Tile_X5Y15_N4BEG[7] ;
 wire \Tile_X5Y15_N4BEG[8] ;
 wire \Tile_X5Y15_N4BEG[9] ;
 wire \Tile_X5Y15_NN4BEG[0] ;
 wire \Tile_X5Y15_NN4BEG[10] ;
 wire \Tile_X5Y15_NN4BEG[11] ;
 wire \Tile_X5Y15_NN4BEG[12] ;
 wire \Tile_X5Y15_NN4BEG[13] ;
 wire \Tile_X5Y15_NN4BEG[14] ;
 wire \Tile_X5Y15_NN4BEG[15] ;
 wire \Tile_X5Y15_NN4BEG[1] ;
 wire \Tile_X5Y15_NN4BEG[2] ;
 wire \Tile_X5Y15_NN4BEG[3] ;
 wire \Tile_X5Y15_NN4BEG[4] ;
 wire \Tile_X5Y15_NN4BEG[5] ;
 wire \Tile_X5Y15_NN4BEG[6] ;
 wire \Tile_X5Y15_NN4BEG[7] ;
 wire \Tile_X5Y15_NN4BEG[8] ;
 wire \Tile_X5Y15_NN4BEG[9] ;
 wire Tile_X5Y15_UserCLKo;
 wire Tile_X5Y1_Co;
 wire \Tile_X5Y1_E1BEG[0] ;
 wire \Tile_X5Y1_E1BEG[1] ;
 wire \Tile_X5Y1_E1BEG[2] ;
 wire \Tile_X5Y1_E1BEG[3] ;
 wire \Tile_X5Y1_E2BEG[0] ;
 wire \Tile_X5Y1_E2BEG[1] ;
 wire \Tile_X5Y1_E2BEG[2] ;
 wire \Tile_X5Y1_E2BEG[3] ;
 wire \Tile_X5Y1_E2BEG[4] ;
 wire \Tile_X5Y1_E2BEG[5] ;
 wire \Tile_X5Y1_E2BEG[6] ;
 wire \Tile_X5Y1_E2BEG[7] ;
 wire \Tile_X5Y1_E2BEGb[0] ;
 wire \Tile_X5Y1_E2BEGb[1] ;
 wire \Tile_X5Y1_E2BEGb[2] ;
 wire \Tile_X5Y1_E2BEGb[3] ;
 wire \Tile_X5Y1_E2BEGb[4] ;
 wire \Tile_X5Y1_E2BEGb[5] ;
 wire \Tile_X5Y1_E2BEGb[6] ;
 wire \Tile_X5Y1_E2BEGb[7] ;
 wire \Tile_X5Y1_E6BEG[0] ;
 wire \Tile_X5Y1_E6BEG[10] ;
 wire \Tile_X5Y1_E6BEG[11] ;
 wire \Tile_X5Y1_E6BEG[1] ;
 wire \Tile_X5Y1_E6BEG[2] ;
 wire \Tile_X5Y1_E6BEG[3] ;
 wire \Tile_X5Y1_E6BEG[4] ;
 wire \Tile_X5Y1_E6BEG[5] ;
 wire \Tile_X5Y1_E6BEG[6] ;
 wire \Tile_X5Y1_E6BEG[7] ;
 wire \Tile_X5Y1_E6BEG[8] ;
 wire \Tile_X5Y1_E6BEG[9] ;
 wire \Tile_X5Y1_EE4BEG[0] ;
 wire \Tile_X5Y1_EE4BEG[10] ;
 wire \Tile_X5Y1_EE4BEG[11] ;
 wire \Tile_X5Y1_EE4BEG[12] ;
 wire \Tile_X5Y1_EE4BEG[13] ;
 wire \Tile_X5Y1_EE4BEG[14] ;
 wire \Tile_X5Y1_EE4BEG[15] ;
 wire \Tile_X5Y1_EE4BEG[1] ;
 wire \Tile_X5Y1_EE4BEG[2] ;
 wire \Tile_X5Y1_EE4BEG[3] ;
 wire \Tile_X5Y1_EE4BEG[4] ;
 wire \Tile_X5Y1_EE4BEG[5] ;
 wire \Tile_X5Y1_EE4BEG[6] ;
 wire \Tile_X5Y1_EE4BEG[7] ;
 wire \Tile_X5Y1_EE4BEG[8] ;
 wire \Tile_X5Y1_EE4BEG[9] ;
 wire \Tile_X5Y1_FrameData_O[0] ;
 wire \Tile_X5Y1_FrameData_O[10] ;
 wire \Tile_X5Y1_FrameData_O[11] ;
 wire \Tile_X5Y1_FrameData_O[12] ;
 wire \Tile_X5Y1_FrameData_O[13] ;
 wire \Tile_X5Y1_FrameData_O[14] ;
 wire \Tile_X5Y1_FrameData_O[15] ;
 wire \Tile_X5Y1_FrameData_O[16] ;
 wire \Tile_X5Y1_FrameData_O[17] ;
 wire \Tile_X5Y1_FrameData_O[18] ;
 wire \Tile_X5Y1_FrameData_O[19] ;
 wire \Tile_X5Y1_FrameData_O[1] ;
 wire \Tile_X5Y1_FrameData_O[20] ;
 wire \Tile_X5Y1_FrameData_O[21] ;
 wire \Tile_X5Y1_FrameData_O[22] ;
 wire \Tile_X5Y1_FrameData_O[23] ;
 wire \Tile_X5Y1_FrameData_O[24] ;
 wire \Tile_X5Y1_FrameData_O[25] ;
 wire \Tile_X5Y1_FrameData_O[26] ;
 wire \Tile_X5Y1_FrameData_O[27] ;
 wire \Tile_X5Y1_FrameData_O[28] ;
 wire \Tile_X5Y1_FrameData_O[29] ;
 wire \Tile_X5Y1_FrameData_O[2] ;
 wire \Tile_X5Y1_FrameData_O[30] ;
 wire \Tile_X5Y1_FrameData_O[31] ;
 wire \Tile_X5Y1_FrameData_O[3] ;
 wire \Tile_X5Y1_FrameData_O[4] ;
 wire \Tile_X5Y1_FrameData_O[5] ;
 wire \Tile_X5Y1_FrameData_O[6] ;
 wire \Tile_X5Y1_FrameData_O[7] ;
 wire \Tile_X5Y1_FrameData_O[8] ;
 wire \Tile_X5Y1_FrameData_O[9] ;
 wire \Tile_X5Y1_FrameStrobe_O[0] ;
 wire \Tile_X5Y1_FrameStrobe_O[10] ;
 wire \Tile_X5Y1_FrameStrobe_O[11] ;
 wire \Tile_X5Y1_FrameStrobe_O[12] ;
 wire \Tile_X5Y1_FrameStrobe_O[13] ;
 wire \Tile_X5Y1_FrameStrobe_O[14] ;
 wire \Tile_X5Y1_FrameStrobe_O[15] ;
 wire \Tile_X5Y1_FrameStrobe_O[16] ;
 wire \Tile_X5Y1_FrameStrobe_O[17] ;
 wire \Tile_X5Y1_FrameStrobe_O[18] ;
 wire \Tile_X5Y1_FrameStrobe_O[19] ;
 wire \Tile_X5Y1_FrameStrobe_O[1] ;
 wire \Tile_X5Y1_FrameStrobe_O[2] ;
 wire \Tile_X5Y1_FrameStrobe_O[3] ;
 wire \Tile_X5Y1_FrameStrobe_O[4] ;
 wire \Tile_X5Y1_FrameStrobe_O[5] ;
 wire \Tile_X5Y1_FrameStrobe_O[6] ;
 wire \Tile_X5Y1_FrameStrobe_O[7] ;
 wire \Tile_X5Y1_FrameStrobe_O[8] ;
 wire \Tile_X5Y1_FrameStrobe_O[9] ;
 wire \Tile_X5Y1_N1BEG[0] ;
 wire \Tile_X5Y1_N1BEG[1] ;
 wire \Tile_X5Y1_N1BEG[2] ;
 wire \Tile_X5Y1_N1BEG[3] ;
 wire \Tile_X5Y1_N2BEG[0] ;
 wire \Tile_X5Y1_N2BEG[1] ;
 wire \Tile_X5Y1_N2BEG[2] ;
 wire \Tile_X5Y1_N2BEG[3] ;
 wire \Tile_X5Y1_N2BEG[4] ;
 wire \Tile_X5Y1_N2BEG[5] ;
 wire \Tile_X5Y1_N2BEG[6] ;
 wire \Tile_X5Y1_N2BEG[7] ;
 wire \Tile_X5Y1_N2BEGb[0] ;
 wire \Tile_X5Y1_N2BEGb[1] ;
 wire \Tile_X5Y1_N2BEGb[2] ;
 wire \Tile_X5Y1_N2BEGb[3] ;
 wire \Tile_X5Y1_N2BEGb[4] ;
 wire \Tile_X5Y1_N2BEGb[5] ;
 wire \Tile_X5Y1_N2BEGb[6] ;
 wire \Tile_X5Y1_N2BEGb[7] ;
 wire \Tile_X5Y1_N4BEG[0] ;
 wire \Tile_X5Y1_N4BEG[10] ;
 wire \Tile_X5Y1_N4BEG[11] ;
 wire \Tile_X5Y1_N4BEG[12] ;
 wire \Tile_X5Y1_N4BEG[13] ;
 wire \Tile_X5Y1_N4BEG[14] ;
 wire \Tile_X5Y1_N4BEG[15] ;
 wire \Tile_X5Y1_N4BEG[1] ;
 wire \Tile_X5Y1_N4BEG[2] ;
 wire \Tile_X5Y1_N4BEG[3] ;
 wire \Tile_X5Y1_N4BEG[4] ;
 wire \Tile_X5Y1_N4BEG[5] ;
 wire \Tile_X5Y1_N4BEG[6] ;
 wire \Tile_X5Y1_N4BEG[7] ;
 wire \Tile_X5Y1_N4BEG[8] ;
 wire \Tile_X5Y1_N4BEG[9] ;
 wire \Tile_X5Y1_NN4BEG[0] ;
 wire \Tile_X5Y1_NN4BEG[10] ;
 wire \Tile_X5Y1_NN4BEG[11] ;
 wire \Tile_X5Y1_NN4BEG[12] ;
 wire \Tile_X5Y1_NN4BEG[13] ;
 wire \Tile_X5Y1_NN4BEG[14] ;
 wire \Tile_X5Y1_NN4BEG[15] ;
 wire \Tile_X5Y1_NN4BEG[1] ;
 wire \Tile_X5Y1_NN4BEG[2] ;
 wire \Tile_X5Y1_NN4BEG[3] ;
 wire \Tile_X5Y1_NN4BEG[4] ;
 wire \Tile_X5Y1_NN4BEG[5] ;
 wire \Tile_X5Y1_NN4BEG[6] ;
 wire \Tile_X5Y1_NN4BEG[7] ;
 wire \Tile_X5Y1_NN4BEG[8] ;
 wire \Tile_X5Y1_NN4BEG[9] ;
 wire \Tile_X5Y1_S1BEG[0] ;
 wire \Tile_X5Y1_S1BEG[1] ;
 wire \Tile_X5Y1_S1BEG[2] ;
 wire \Tile_X5Y1_S1BEG[3] ;
 wire \Tile_X5Y1_S2BEG[0] ;
 wire \Tile_X5Y1_S2BEG[1] ;
 wire \Tile_X5Y1_S2BEG[2] ;
 wire \Tile_X5Y1_S2BEG[3] ;
 wire \Tile_X5Y1_S2BEG[4] ;
 wire \Tile_X5Y1_S2BEG[5] ;
 wire \Tile_X5Y1_S2BEG[6] ;
 wire \Tile_X5Y1_S2BEG[7] ;
 wire \Tile_X5Y1_S2BEGb[0] ;
 wire \Tile_X5Y1_S2BEGb[1] ;
 wire \Tile_X5Y1_S2BEGb[2] ;
 wire \Tile_X5Y1_S2BEGb[3] ;
 wire \Tile_X5Y1_S2BEGb[4] ;
 wire \Tile_X5Y1_S2BEGb[5] ;
 wire \Tile_X5Y1_S2BEGb[6] ;
 wire \Tile_X5Y1_S2BEGb[7] ;
 wire \Tile_X5Y1_S4BEG[0] ;
 wire \Tile_X5Y1_S4BEG[10] ;
 wire \Tile_X5Y1_S4BEG[11] ;
 wire \Tile_X5Y1_S4BEG[12] ;
 wire \Tile_X5Y1_S4BEG[13] ;
 wire \Tile_X5Y1_S4BEG[14] ;
 wire \Tile_X5Y1_S4BEG[15] ;
 wire \Tile_X5Y1_S4BEG[1] ;
 wire \Tile_X5Y1_S4BEG[2] ;
 wire \Tile_X5Y1_S4BEG[3] ;
 wire \Tile_X5Y1_S4BEG[4] ;
 wire \Tile_X5Y1_S4BEG[5] ;
 wire \Tile_X5Y1_S4BEG[6] ;
 wire \Tile_X5Y1_S4BEG[7] ;
 wire \Tile_X5Y1_S4BEG[8] ;
 wire \Tile_X5Y1_S4BEG[9] ;
 wire \Tile_X5Y1_SS4BEG[0] ;
 wire \Tile_X5Y1_SS4BEG[10] ;
 wire \Tile_X5Y1_SS4BEG[11] ;
 wire \Tile_X5Y1_SS4BEG[12] ;
 wire \Tile_X5Y1_SS4BEG[13] ;
 wire \Tile_X5Y1_SS4BEG[14] ;
 wire \Tile_X5Y1_SS4BEG[15] ;
 wire \Tile_X5Y1_SS4BEG[1] ;
 wire \Tile_X5Y1_SS4BEG[2] ;
 wire \Tile_X5Y1_SS4BEG[3] ;
 wire \Tile_X5Y1_SS4BEG[4] ;
 wire \Tile_X5Y1_SS4BEG[5] ;
 wire \Tile_X5Y1_SS4BEG[6] ;
 wire \Tile_X5Y1_SS4BEG[7] ;
 wire \Tile_X5Y1_SS4BEG[8] ;
 wire \Tile_X5Y1_SS4BEG[9] ;
 wire Tile_X5Y1_UserCLKo;
 wire \Tile_X5Y1_W1BEG[0] ;
 wire \Tile_X5Y1_W1BEG[1] ;
 wire \Tile_X5Y1_W1BEG[2] ;
 wire \Tile_X5Y1_W1BEG[3] ;
 wire \Tile_X5Y1_W2BEG[0] ;
 wire \Tile_X5Y1_W2BEG[1] ;
 wire \Tile_X5Y1_W2BEG[2] ;
 wire \Tile_X5Y1_W2BEG[3] ;
 wire \Tile_X5Y1_W2BEG[4] ;
 wire \Tile_X5Y1_W2BEG[5] ;
 wire \Tile_X5Y1_W2BEG[6] ;
 wire \Tile_X5Y1_W2BEG[7] ;
 wire \Tile_X5Y1_W2BEGb[0] ;
 wire \Tile_X5Y1_W2BEGb[1] ;
 wire \Tile_X5Y1_W2BEGb[2] ;
 wire \Tile_X5Y1_W2BEGb[3] ;
 wire \Tile_X5Y1_W2BEGb[4] ;
 wire \Tile_X5Y1_W2BEGb[5] ;
 wire \Tile_X5Y1_W2BEGb[6] ;
 wire \Tile_X5Y1_W2BEGb[7] ;
 wire \Tile_X5Y1_W6BEG[0] ;
 wire \Tile_X5Y1_W6BEG[10] ;
 wire \Tile_X5Y1_W6BEG[11] ;
 wire \Tile_X5Y1_W6BEG[1] ;
 wire \Tile_X5Y1_W6BEG[2] ;
 wire \Tile_X5Y1_W6BEG[3] ;
 wire \Tile_X5Y1_W6BEG[4] ;
 wire \Tile_X5Y1_W6BEG[5] ;
 wire \Tile_X5Y1_W6BEG[6] ;
 wire \Tile_X5Y1_W6BEG[7] ;
 wire \Tile_X5Y1_W6BEG[8] ;
 wire \Tile_X5Y1_W6BEG[9] ;
 wire \Tile_X5Y1_WW4BEG[0] ;
 wire \Tile_X5Y1_WW4BEG[10] ;
 wire \Tile_X5Y1_WW4BEG[11] ;
 wire \Tile_X5Y1_WW4BEG[12] ;
 wire \Tile_X5Y1_WW4BEG[13] ;
 wire \Tile_X5Y1_WW4BEG[14] ;
 wire \Tile_X5Y1_WW4BEG[15] ;
 wire \Tile_X5Y1_WW4BEG[1] ;
 wire \Tile_X5Y1_WW4BEG[2] ;
 wire \Tile_X5Y1_WW4BEG[3] ;
 wire \Tile_X5Y1_WW4BEG[4] ;
 wire \Tile_X5Y1_WW4BEG[5] ;
 wire \Tile_X5Y1_WW4BEG[6] ;
 wire \Tile_X5Y1_WW4BEG[7] ;
 wire \Tile_X5Y1_WW4BEG[8] ;
 wire \Tile_X5Y1_WW4BEG[9] ;
 wire Tile_X5Y2_Co;
 wire \Tile_X5Y2_E1BEG[0] ;
 wire \Tile_X5Y2_E1BEG[1] ;
 wire \Tile_X5Y2_E1BEG[2] ;
 wire \Tile_X5Y2_E1BEG[3] ;
 wire \Tile_X5Y2_E2BEG[0] ;
 wire \Tile_X5Y2_E2BEG[1] ;
 wire \Tile_X5Y2_E2BEG[2] ;
 wire \Tile_X5Y2_E2BEG[3] ;
 wire \Tile_X5Y2_E2BEG[4] ;
 wire \Tile_X5Y2_E2BEG[5] ;
 wire \Tile_X5Y2_E2BEG[6] ;
 wire \Tile_X5Y2_E2BEG[7] ;
 wire \Tile_X5Y2_E2BEGb[0] ;
 wire \Tile_X5Y2_E2BEGb[1] ;
 wire \Tile_X5Y2_E2BEGb[2] ;
 wire \Tile_X5Y2_E2BEGb[3] ;
 wire \Tile_X5Y2_E2BEGb[4] ;
 wire \Tile_X5Y2_E2BEGb[5] ;
 wire \Tile_X5Y2_E2BEGb[6] ;
 wire \Tile_X5Y2_E2BEGb[7] ;
 wire \Tile_X5Y2_E6BEG[0] ;
 wire \Tile_X5Y2_E6BEG[10] ;
 wire \Tile_X5Y2_E6BEG[11] ;
 wire \Tile_X5Y2_E6BEG[1] ;
 wire \Tile_X5Y2_E6BEG[2] ;
 wire \Tile_X5Y2_E6BEG[3] ;
 wire \Tile_X5Y2_E6BEG[4] ;
 wire \Tile_X5Y2_E6BEG[5] ;
 wire \Tile_X5Y2_E6BEG[6] ;
 wire \Tile_X5Y2_E6BEG[7] ;
 wire \Tile_X5Y2_E6BEG[8] ;
 wire \Tile_X5Y2_E6BEG[9] ;
 wire \Tile_X5Y2_EE4BEG[0] ;
 wire \Tile_X5Y2_EE4BEG[10] ;
 wire \Tile_X5Y2_EE4BEG[11] ;
 wire \Tile_X5Y2_EE4BEG[12] ;
 wire \Tile_X5Y2_EE4BEG[13] ;
 wire \Tile_X5Y2_EE4BEG[14] ;
 wire \Tile_X5Y2_EE4BEG[15] ;
 wire \Tile_X5Y2_EE4BEG[1] ;
 wire \Tile_X5Y2_EE4BEG[2] ;
 wire \Tile_X5Y2_EE4BEG[3] ;
 wire \Tile_X5Y2_EE4BEG[4] ;
 wire \Tile_X5Y2_EE4BEG[5] ;
 wire \Tile_X5Y2_EE4BEG[6] ;
 wire \Tile_X5Y2_EE4BEG[7] ;
 wire \Tile_X5Y2_EE4BEG[8] ;
 wire \Tile_X5Y2_EE4BEG[9] ;
 wire \Tile_X5Y2_FrameData_O[0] ;
 wire \Tile_X5Y2_FrameData_O[10] ;
 wire \Tile_X5Y2_FrameData_O[11] ;
 wire \Tile_X5Y2_FrameData_O[12] ;
 wire \Tile_X5Y2_FrameData_O[13] ;
 wire \Tile_X5Y2_FrameData_O[14] ;
 wire \Tile_X5Y2_FrameData_O[15] ;
 wire \Tile_X5Y2_FrameData_O[16] ;
 wire \Tile_X5Y2_FrameData_O[17] ;
 wire \Tile_X5Y2_FrameData_O[18] ;
 wire \Tile_X5Y2_FrameData_O[19] ;
 wire \Tile_X5Y2_FrameData_O[1] ;
 wire \Tile_X5Y2_FrameData_O[20] ;
 wire \Tile_X5Y2_FrameData_O[21] ;
 wire \Tile_X5Y2_FrameData_O[22] ;
 wire \Tile_X5Y2_FrameData_O[23] ;
 wire \Tile_X5Y2_FrameData_O[24] ;
 wire \Tile_X5Y2_FrameData_O[25] ;
 wire \Tile_X5Y2_FrameData_O[26] ;
 wire \Tile_X5Y2_FrameData_O[27] ;
 wire \Tile_X5Y2_FrameData_O[28] ;
 wire \Tile_X5Y2_FrameData_O[29] ;
 wire \Tile_X5Y2_FrameData_O[2] ;
 wire \Tile_X5Y2_FrameData_O[30] ;
 wire \Tile_X5Y2_FrameData_O[31] ;
 wire \Tile_X5Y2_FrameData_O[3] ;
 wire \Tile_X5Y2_FrameData_O[4] ;
 wire \Tile_X5Y2_FrameData_O[5] ;
 wire \Tile_X5Y2_FrameData_O[6] ;
 wire \Tile_X5Y2_FrameData_O[7] ;
 wire \Tile_X5Y2_FrameData_O[8] ;
 wire \Tile_X5Y2_FrameData_O[9] ;
 wire \Tile_X5Y2_FrameStrobe_O[0] ;
 wire \Tile_X5Y2_FrameStrobe_O[10] ;
 wire \Tile_X5Y2_FrameStrobe_O[11] ;
 wire \Tile_X5Y2_FrameStrobe_O[12] ;
 wire \Tile_X5Y2_FrameStrobe_O[13] ;
 wire \Tile_X5Y2_FrameStrobe_O[14] ;
 wire \Tile_X5Y2_FrameStrobe_O[15] ;
 wire \Tile_X5Y2_FrameStrobe_O[16] ;
 wire \Tile_X5Y2_FrameStrobe_O[17] ;
 wire \Tile_X5Y2_FrameStrobe_O[18] ;
 wire \Tile_X5Y2_FrameStrobe_O[19] ;
 wire \Tile_X5Y2_FrameStrobe_O[1] ;
 wire \Tile_X5Y2_FrameStrobe_O[2] ;
 wire \Tile_X5Y2_FrameStrobe_O[3] ;
 wire \Tile_X5Y2_FrameStrobe_O[4] ;
 wire \Tile_X5Y2_FrameStrobe_O[5] ;
 wire \Tile_X5Y2_FrameStrobe_O[6] ;
 wire \Tile_X5Y2_FrameStrobe_O[7] ;
 wire \Tile_X5Y2_FrameStrobe_O[8] ;
 wire \Tile_X5Y2_FrameStrobe_O[9] ;
 wire \Tile_X5Y2_N1BEG[0] ;
 wire \Tile_X5Y2_N1BEG[1] ;
 wire \Tile_X5Y2_N1BEG[2] ;
 wire \Tile_X5Y2_N1BEG[3] ;
 wire \Tile_X5Y2_N2BEG[0] ;
 wire \Tile_X5Y2_N2BEG[1] ;
 wire \Tile_X5Y2_N2BEG[2] ;
 wire \Tile_X5Y2_N2BEG[3] ;
 wire \Tile_X5Y2_N2BEG[4] ;
 wire \Tile_X5Y2_N2BEG[5] ;
 wire \Tile_X5Y2_N2BEG[6] ;
 wire \Tile_X5Y2_N2BEG[7] ;
 wire \Tile_X5Y2_N2BEGb[0] ;
 wire \Tile_X5Y2_N2BEGb[1] ;
 wire \Tile_X5Y2_N2BEGb[2] ;
 wire \Tile_X5Y2_N2BEGb[3] ;
 wire \Tile_X5Y2_N2BEGb[4] ;
 wire \Tile_X5Y2_N2BEGb[5] ;
 wire \Tile_X5Y2_N2BEGb[6] ;
 wire \Tile_X5Y2_N2BEGb[7] ;
 wire \Tile_X5Y2_N4BEG[0] ;
 wire \Tile_X5Y2_N4BEG[10] ;
 wire \Tile_X5Y2_N4BEG[11] ;
 wire \Tile_X5Y2_N4BEG[12] ;
 wire \Tile_X5Y2_N4BEG[13] ;
 wire \Tile_X5Y2_N4BEG[14] ;
 wire \Tile_X5Y2_N4BEG[15] ;
 wire \Tile_X5Y2_N4BEG[1] ;
 wire \Tile_X5Y2_N4BEG[2] ;
 wire \Tile_X5Y2_N4BEG[3] ;
 wire \Tile_X5Y2_N4BEG[4] ;
 wire \Tile_X5Y2_N4BEG[5] ;
 wire \Tile_X5Y2_N4BEG[6] ;
 wire \Tile_X5Y2_N4BEG[7] ;
 wire \Tile_X5Y2_N4BEG[8] ;
 wire \Tile_X5Y2_N4BEG[9] ;
 wire \Tile_X5Y2_NN4BEG[0] ;
 wire \Tile_X5Y2_NN4BEG[10] ;
 wire \Tile_X5Y2_NN4BEG[11] ;
 wire \Tile_X5Y2_NN4BEG[12] ;
 wire \Tile_X5Y2_NN4BEG[13] ;
 wire \Tile_X5Y2_NN4BEG[14] ;
 wire \Tile_X5Y2_NN4BEG[15] ;
 wire \Tile_X5Y2_NN4BEG[1] ;
 wire \Tile_X5Y2_NN4BEG[2] ;
 wire \Tile_X5Y2_NN4BEG[3] ;
 wire \Tile_X5Y2_NN4BEG[4] ;
 wire \Tile_X5Y2_NN4BEG[5] ;
 wire \Tile_X5Y2_NN4BEG[6] ;
 wire \Tile_X5Y2_NN4BEG[7] ;
 wire \Tile_X5Y2_NN4BEG[8] ;
 wire \Tile_X5Y2_NN4BEG[9] ;
 wire \Tile_X5Y2_S1BEG[0] ;
 wire \Tile_X5Y2_S1BEG[1] ;
 wire \Tile_X5Y2_S1BEG[2] ;
 wire \Tile_X5Y2_S1BEG[3] ;
 wire \Tile_X5Y2_S2BEG[0] ;
 wire \Tile_X5Y2_S2BEG[1] ;
 wire \Tile_X5Y2_S2BEG[2] ;
 wire \Tile_X5Y2_S2BEG[3] ;
 wire \Tile_X5Y2_S2BEG[4] ;
 wire \Tile_X5Y2_S2BEG[5] ;
 wire \Tile_X5Y2_S2BEG[6] ;
 wire \Tile_X5Y2_S2BEG[7] ;
 wire \Tile_X5Y2_S2BEGb[0] ;
 wire \Tile_X5Y2_S2BEGb[1] ;
 wire \Tile_X5Y2_S2BEGb[2] ;
 wire \Tile_X5Y2_S2BEGb[3] ;
 wire \Tile_X5Y2_S2BEGb[4] ;
 wire \Tile_X5Y2_S2BEGb[5] ;
 wire \Tile_X5Y2_S2BEGb[6] ;
 wire \Tile_X5Y2_S2BEGb[7] ;
 wire \Tile_X5Y2_S4BEG[0] ;
 wire \Tile_X5Y2_S4BEG[10] ;
 wire \Tile_X5Y2_S4BEG[11] ;
 wire \Tile_X5Y2_S4BEG[12] ;
 wire \Tile_X5Y2_S4BEG[13] ;
 wire \Tile_X5Y2_S4BEG[14] ;
 wire \Tile_X5Y2_S4BEG[15] ;
 wire \Tile_X5Y2_S4BEG[1] ;
 wire \Tile_X5Y2_S4BEG[2] ;
 wire \Tile_X5Y2_S4BEG[3] ;
 wire \Tile_X5Y2_S4BEG[4] ;
 wire \Tile_X5Y2_S4BEG[5] ;
 wire \Tile_X5Y2_S4BEG[6] ;
 wire \Tile_X5Y2_S4BEG[7] ;
 wire \Tile_X5Y2_S4BEG[8] ;
 wire \Tile_X5Y2_S4BEG[9] ;
 wire \Tile_X5Y2_SS4BEG[0] ;
 wire \Tile_X5Y2_SS4BEG[10] ;
 wire \Tile_X5Y2_SS4BEG[11] ;
 wire \Tile_X5Y2_SS4BEG[12] ;
 wire \Tile_X5Y2_SS4BEG[13] ;
 wire \Tile_X5Y2_SS4BEG[14] ;
 wire \Tile_X5Y2_SS4BEG[15] ;
 wire \Tile_X5Y2_SS4BEG[1] ;
 wire \Tile_X5Y2_SS4BEG[2] ;
 wire \Tile_X5Y2_SS4BEG[3] ;
 wire \Tile_X5Y2_SS4BEG[4] ;
 wire \Tile_X5Y2_SS4BEG[5] ;
 wire \Tile_X5Y2_SS4BEG[6] ;
 wire \Tile_X5Y2_SS4BEG[7] ;
 wire \Tile_X5Y2_SS4BEG[8] ;
 wire \Tile_X5Y2_SS4BEG[9] ;
 wire Tile_X5Y2_UserCLKo;
 wire \Tile_X5Y2_W1BEG[0] ;
 wire \Tile_X5Y2_W1BEG[1] ;
 wire \Tile_X5Y2_W1BEG[2] ;
 wire \Tile_X5Y2_W1BEG[3] ;
 wire \Tile_X5Y2_W2BEG[0] ;
 wire \Tile_X5Y2_W2BEG[1] ;
 wire \Tile_X5Y2_W2BEG[2] ;
 wire \Tile_X5Y2_W2BEG[3] ;
 wire \Tile_X5Y2_W2BEG[4] ;
 wire \Tile_X5Y2_W2BEG[5] ;
 wire \Tile_X5Y2_W2BEG[6] ;
 wire \Tile_X5Y2_W2BEG[7] ;
 wire \Tile_X5Y2_W2BEGb[0] ;
 wire \Tile_X5Y2_W2BEGb[1] ;
 wire \Tile_X5Y2_W2BEGb[2] ;
 wire \Tile_X5Y2_W2BEGb[3] ;
 wire \Tile_X5Y2_W2BEGb[4] ;
 wire \Tile_X5Y2_W2BEGb[5] ;
 wire \Tile_X5Y2_W2BEGb[6] ;
 wire \Tile_X5Y2_W2BEGb[7] ;
 wire \Tile_X5Y2_W6BEG[0] ;
 wire \Tile_X5Y2_W6BEG[10] ;
 wire \Tile_X5Y2_W6BEG[11] ;
 wire \Tile_X5Y2_W6BEG[1] ;
 wire \Tile_X5Y2_W6BEG[2] ;
 wire \Tile_X5Y2_W6BEG[3] ;
 wire \Tile_X5Y2_W6BEG[4] ;
 wire \Tile_X5Y2_W6BEG[5] ;
 wire \Tile_X5Y2_W6BEG[6] ;
 wire \Tile_X5Y2_W6BEG[7] ;
 wire \Tile_X5Y2_W6BEG[8] ;
 wire \Tile_X5Y2_W6BEG[9] ;
 wire \Tile_X5Y2_WW4BEG[0] ;
 wire \Tile_X5Y2_WW4BEG[10] ;
 wire \Tile_X5Y2_WW4BEG[11] ;
 wire \Tile_X5Y2_WW4BEG[12] ;
 wire \Tile_X5Y2_WW4BEG[13] ;
 wire \Tile_X5Y2_WW4BEG[14] ;
 wire \Tile_X5Y2_WW4BEG[15] ;
 wire \Tile_X5Y2_WW4BEG[1] ;
 wire \Tile_X5Y2_WW4BEG[2] ;
 wire \Tile_X5Y2_WW4BEG[3] ;
 wire \Tile_X5Y2_WW4BEG[4] ;
 wire \Tile_X5Y2_WW4BEG[5] ;
 wire \Tile_X5Y2_WW4BEG[6] ;
 wire \Tile_X5Y2_WW4BEG[7] ;
 wire \Tile_X5Y2_WW4BEG[8] ;
 wire \Tile_X5Y2_WW4BEG[9] ;
 wire Tile_X5Y3_Co;
 wire \Tile_X5Y3_E1BEG[0] ;
 wire \Tile_X5Y3_E1BEG[1] ;
 wire \Tile_X5Y3_E1BEG[2] ;
 wire \Tile_X5Y3_E1BEG[3] ;
 wire \Tile_X5Y3_E2BEG[0] ;
 wire \Tile_X5Y3_E2BEG[1] ;
 wire \Tile_X5Y3_E2BEG[2] ;
 wire \Tile_X5Y3_E2BEG[3] ;
 wire \Tile_X5Y3_E2BEG[4] ;
 wire \Tile_X5Y3_E2BEG[5] ;
 wire \Tile_X5Y3_E2BEG[6] ;
 wire \Tile_X5Y3_E2BEG[7] ;
 wire \Tile_X5Y3_E2BEGb[0] ;
 wire \Tile_X5Y3_E2BEGb[1] ;
 wire \Tile_X5Y3_E2BEGb[2] ;
 wire \Tile_X5Y3_E2BEGb[3] ;
 wire \Tile_X5Y3_E2BEGb[4] ;
 wire \Tile_X5Y3_E2BEGb[5] ;
 wire \Tile_X5Y3_E2BEGb[6] ;
 wire \Tile_X5Y3_E2BEGb[7] ;
 wire \Tile_X5Y3_E6BEG[0] ;
 wire \Tile_X5Y3_E6BEG[10] ;
 wire \Tile_X5Y3_E6BEG[11] ;
 wire \Tile_X5Y3_E6BEG[1] ;
 wire \Tile_X5Y3_E6BEG[2] ;
 wire \Tile_X5Y3_E6BEG[3] ;
 wire \Tile_X5Y3_E6BEG[4] ;
 wire \Tile_X5Y3_E6BEG[5] ;
 wire \Tile_X5Y3_E6BEG[6] ;
 wire \Tile_X5Y3_E6BEG[7] ;
 wire \Tile_X5Y3_E6BEG[8] ;
 wire \Tile_X5Y3_E6BEG[9] ;
 wire \Tile_X5Y3_EE4BEG[0] ;
 wire \Tile_X5Y3_EE4BEG[10] ;
 wire \Tile_X5Y3_EE4BEG[11] ;
 wire \Tile_X5Y3_EE4BEG[12] ;
 wire \Tile_X5Y3_EE4BEG[13] ;
 wire \Tile_X5Y3_EE4BEG[14] ;
 wire \Tile_X5Y3_EE4BEG[15] ;
 wire \Tile_X5Y3_EE4BEG[1] ;
 wire \Tile_X5Y3_EE4BEG[2] ;
 wire \Tile_X5Y3_EE4BEG[3] ;
 wire \Tile_X5Y3_EE4BEG[4] ;
 wire \Tile_X5Y3_EE4BEG[5] ;
 wire \Tile_X5Y3_EE4BEG[6] ;
 wire \Tile_X5Y3_EE4BEG[7] ;
 wire \Tile_X5Y3_EE4BEG[8] ;
 wire \Tile_X5Y3_EE4BEG[9] ;
 wire \Tile_X5Y3_FrameData_O[0] ;
 wire \Tile_X5Y3_FrameData_O[10] ;
 wire \Tile_X5Y3_FrameData_O[11] ;
 wire \Tile_X5Y3_FrameData_O[12] ;
 wire \Tile_X5Y3_FrameData_O[13] ;
 wire \Tile_X5Y3_FrameData_O[14] ;
 wire \Tile_X5Y3_FrameData_O[15] ;
 wire \Tile_X5Y3_FrameData_O[16] ;
 wire \Tile_X5Y3_FrameData_O[17] ;
 wire \Tile_X5Y3_FrameData_O[18] ;
 wire \Tile_X5Y3_FrameData_O[19] ;
 wire \Tile_X5Y3_FrameData_O[1] ;
 wire \Tile_X5Y3_FrameData_O[20] ;
 wire \Tile_X5Y3_FrameData_O[21] ;
 wire \Tile_X5Y3_FrameData_O[22] ;
 wire \Tile_X5Y3_FrameData_O[23] ;
 wire \Tile_X5Y3_FrameData_O[24] ;
 wire \Tile_X5Y3_FrameData_O[25] ;
 wire \Tile_X5Y3_FrameData_O[26] ;
 wire \Tile_X5Y3_FrameData_O[27] ;
 wire \Tile_X5Y3_FrameData_O[28] ;
 wire \Tile_X5Y3_FrameData_O[29] ;
 wire \Tile_X5Y3_FrameData_O[2] ;
 wire \Tile_X5Y3_FrameData_O[30] ;
 wire \Tile_X5Y3_FrameData_O[31] ;
 wire \Tile_X5Y3_FrameData_O[3] ;
 wire \Tile_X5Y3_FrameData_O[4] ;
 wire \Tile_X5Y3_FrameData_O[5] ;
 wire \Tile_X5Y3_FrameData_O[6] ;
 wire \Tile_X5Y3_FrameData_O[7] ;
 wire \Tile_X5Y3_FrameData_O[8] ;
 wire \Tile_X5Y3_FrameData_O[9] ;
 wire \Tile_X5Y3_FrameStrobe_O[0] ;
 wire \Tile_X5Y3_FrameStrobe_O[10] ;
 wire \Tile_X5Y3_FrameStrobe_O[11] ;
 wire \Tile_X5Y3_FrameStrobe_O[12] ;
 wire \Tile_X5Y3_FrameStrobe_O[13] ;
 wire \Tile_X5Y3_FrameStrobe_O[14] ;
 wire \Tile_X5Y3_FrameStrobe_O[15] ;
 wire \Tile_X5Y3_FrameStrobe_O[16] ;
 wire \Tile_X5Y3_FrameStrobe_O[17] ;
 wire \Tile_X5Y3_FrameStrobe_O[18] ;
 wire \Tile_X5Y3_FrameStrobe_O[19] ;
 wire \Tile_X5Y3_FrameStrobe_O[1] ;
 wire \Tile_X5Y3_FrameStrobe_O[2] ;
 wire \Tile_X5Y3_FrameStrobe_O[3] ;
 wire \Tile_X5Y3_FrameStrobe_O[4] ;
 wire \Tile_X5Y3_FrameStrobe_O[5] ;
 wire \Tile_X5Y3_FrameStrobe_O[6] ;
 wire \Tile_X5Y3_FrameStrobe_O[7] ;
 wire \Tile_X5Y3_FrameStrobe_O[8] ;
 wire \Tile_X5Y3_FrameStrobe_O[9] ;
 wire \Tile_X5Y3_N1BEG[0] ;
 wire \Tile_X5Y3_N1BEG[1] ;
 wire \Tile_X5Y3_N1BEG[2] ;
 wire \Tile_X5Y3_N1BEG[3] ;
 wire \Tile_X5Y3_N2BEG[0] ;
 wire \Tile_X5Y3_N2BEG[1] ;
 wire \Tile_X5Y3_N2BEG[2] ;
 wire \Tile_X5Y3_N2BEG[3] ;
 wire \Tile_X5Y3_N2BEG[4] ;
 wire \Tile_X5Y3_N2BEG[5] ;
 wire \Tile_X5Y3_N2BEG[6] ;
 wire \Tile_X5Y3_N2BEG[7] ;
 wire \Tile_X5Y3_N2BEGb[0] ;
 wire \Tile_X5Y3_N2BEGb[1] ;
 wire \Tile_X5Y3_N2BEGb[2] ;
 wire \Tile_X5Y3_N2BEGb[3] ;
 wire \Tile_X5Y3_N2BEGb[4] ;
 wire \Tile_X5Y3_N2BEGb[5] ;
 wire \Tile_X5Y3_N2BEGb[6] ;
 wire \Tile_X5Y3_N2BEGb[7] ;
 wire \Tile_X5Y3_N4BEG[0] ;
 wire \Tile_X5Y3_N4BEG[10] ;
 wire \Tile_X5Y3_N4BEG[11] ;
 wire \Tile_X5Y3_N4BEG[12] ;
 wire \Tile_X5Y3_N4BEG[13] ;
 wire \Tile_X5Y3_N4BEG[14] ;
 wire \Tile_X5Y3_N4BEG[15] ;
 wire \Tile_X5Y3_N4BEG[1] ;
 wire \Tile_X5Y3_N4BEG[2] ;
 wire \Tile_X5Y3_N4BEG[3] ;
 wire \Tile_X5Y3_N4BEG[4] ;
 wire \Tile_X5Y3_N4BEG[5] ;
 wire \Tile_X5Y3_N4BEG[6] ;
 wire \Tile_X5Y3_N4BEG[7] ;
 wire \Tile_X5Y3_N4BEG[8] ;
 wire \Tile_X5Y3_N4BEG[9] ;
 wire \Tile_X5Y3_NN4BEG[0] ;
 wire \Tile_X5Y3_NN4BEG[10] ;
 wire \Tile_X5Y3_NN4BEG[11] ;
 wire \Tile_X5Y3_NN4BEG[12] ;
 wire \Tile_X5Y3_NN4BEG[13] ;
 wire \Tile_X5Y3_NN4BEG[14] ;
 wire \Tile_X5Y3_NN4BEG[15] ;
 wire \Tile_X5Y3_NN4BEG[1] ;
 wire \Tile_X5Y3_NN4BEG[2] ;
 wire \Tile_X5Y3_NN4BEG[3] ;
 wire \Tile_X5Y3_NN4BEG[4] ;
 wire \Tile_X5Y3_NN4BEG[5] ;
 wire \Tile_X5Y3_NN4BEG[6] ;
 wire \Tile_X5Y3_NN4BEG[7] ;
 wire \Tile_X5Y3_NN4BEG[8] ;
 wire \Tile_X5Y3_NN4BEG[9] ;
 wire \Tile_X5Y3_S1BEG[0] ;
 wire \Tile_X5Y3_S1BEG[1] ;
 wire \Tile_X5Y3_S1BEG[2] ;
 wire \Tile_X5Y3_S1BEG[3] ;
 wire \Tile_X5Y3_S2BEG[0] ;
 wire \Tile_X5Y3_S2BEG[1] ;
 wire \Tile_X5Y3_S2BEG[2] ;
 wire \Tile_X5Y3_S2BEG[3] ;
 wire \Tile_X5Y3_S2BEG[4] ;
 wire \Tile_X5Y3_S2BEG[5] ;
 wire \Tile_X5Y3_S2BEG[6] ;
 wire \Tile_X5Y3_S2BEG[7] ;
 wire \Tile_X5Y3_S2BEGb[0] ;
 wire \Tile_X5Y3_S2BEGb[1] ;
 wire \Tile_X5Y3_S2BEGb[2] ;
 wire \Tile_X5Y3_S2BEGb[3] ;
 wire \Tile_X5Y3_S2BEGb[4] ;
 wire \Tile_X5Y3_S2BEGb[5] ;
 wire \Tile_X5Y3_S2BEGb[6] ;
 wire \Tile_X5Y3_S2BEGb[7] ;
 wire \Tile_X5Y3_S4BEG[0] ;
 wire \Tile_X5Y3_S4BEG[10] ;
 wire \Tile_X5Y3_S4BEG[11] ;
 wire \Tile_X5Y3_S4BEG[12] ;
 wire \Tile_X5Y3_S4BEG[13] ;
 wire \Tile_X5Y3_S4BEG[14] ;
 wire \Tile_X5Y3_S4BEG[15] ;
 wire \Tile_X5Y3_S4BEG[1] ;
 wire \Tile_X5Y3_S4BEG[2] ;
 wire \Tile_X5Y3_S4BEG[3] ;
 wire \Tile_X5Y3_S4BEG[4] ;
 wire \Tile_X5Y3_S4BEG[5] ;
 wire \Tile_X5Y3_S4BEG[6] ;
 wire \Tile_X5Y3_S4BEG[7] ;
 wire \Tile_X5Y3_S4BEG[8] ;
 wire \Tile_X5Y3_S4BEG[9] ;
 wire \Tile_X5Y3_SS4BEG[0] ;
 wire \Tile_X5Y3_SS4BEG[10] ;
 wire \Tile_X5Y3_SS4BEG[11] ;
 wire \Tile_X5Y3_SS4BEG[12] ;
 wire \Tile_X5Y3_SS4BEG[13] ;
 wire \Tile_X5Y3_SS4BEG[14] ;
 wire \Tile_X5Y3_SS4BEG[15] ;
 wire \Tile_X5Y3_SS4BEG[1] ;
 wire \Tile_X5Y3_SS4BEG[2] ;
 wire \Tile_X5Y3_SS4BEG[3] ;
 wire \Tile_X5Y3_SS4BEG[4] ;
 wire \Tile_X5Y3_SS4BEG[5] ;
 wire \Tile_X5Y3_SS4BEG[6] ;
 wire \Tile_X5Y3_SS4BEG[7] ;
 wire \Tile_X5Y3_SS4BEG[8] ;
 wire \Tile_X5Y3_SS4BEG[9] ;
 wire Tile_X5Y3_UserCLKo;
 wire \Tile_X5Y3_W1BEG[0] ;
 wire \Tile_X5Y3_W1BEG[1] ;
 wire \Tile_X5Y3_W1BEG[2] ;
 wire \Tile_X5Y3_W1BEG[3] ;
 wire \Tile_X5Y3_W2BEG[0] ;
 wire \Tile_X5Y3_W2BEG[1] ;
 wire \Tile_X5Y3_W2BEG[2] ;
 wire \Tile_X5Y3_W2BEG[3] ;
 wire \Tile_X5Y3_W2BEG[4] ;
 wire \Tile_X5Y3_W2BEG[5] ;
 wire \Tile_X5Y3_W2BEG[6] ;
 wire \Tile_X5Y3_W2BEG[7] ;
 wire \Tile_X5Y3_W2BEGb[0] ;
 wire \Tile_X5Y3_W2BEGb[1] ;
 wire \Tile_X5Y3_W2BEGb[2] ;
 wire \Tile_X5Y3_W2BEGb[3] ;
 wire \Tile_X5Y3_W2BEGb[4] ;
 wire \Tile_X5Y3_W2BEGb[5] ;
 wire \Tile_X5Y3_W2BEGb[6] ;
 wire \Tile_X5Y3_W2BEGb[7] ;
 wire \Tile_X5Y3_W6BEG[0] ;
 wire \Tile_X5Y3_W6BEG[10] ;
 wire \Tile_X5Y3_W6BEG[11] ;
 wire \Tile_X5Y3_W6BEG[1] ;
 wire \Tile_X5Y3_W6BEG[2] ;
 wire \Tile_X5Y3_W6BEG[3] ;
 wire \Tile_X5Y3_W6BEG[4] ;
 wire \Tile_X5Y3_W6BEG[5] ;
 wire \Tile_X5Y3_W6BEG[6] ;
 wire \Tile_X5Y3_W6BEG[7] ;
 wire \Tile_X5Y3_W6BEG[8] ;
 wire \Tile_X5Y3_W6BEG[9] ;
 wire \Tile_X5Y3_WW4BEG[0] ;
 wire \Tile_X5Y3_WW4BEG[10] ;
 wire \Tile_X5Y3_WW4BEG[11] ;
 wire \Tile_X5Y3_WW4BEG[12] ;
 wire \Tile_X5Y3_WW4BEG[13] ;
 wire \Tile_X5Y3_WW4BEG[14] ;
 wire \Tile_X5Y3_WW4BEG[15] ;
 wire \Tile_X5Y3_WW4BEG[1] ;
 wire \Tile_X5Y3_WW4BEG[2] ;
 wire \Tile_X5Y3_WW4BEG[3] ;
 wire \Tile_X5Y3_WW4BEG[4] ;
 wire \Tile_X5Y3_WW4BEG[5] ;
 wire \Tile_X5Y3_WW4BEG[6] ;
 wire \Tile_X5Y3_WW4BEG[7] ;
 wire \Tile_X5Y3_WW4BEG[8] ;
 wire \Tile_X5Y3_WW4BEG[9] ;
 wire Tile_X5Y4_Co;
 wire \Tile_X5Y4_E1BEG[0] ;
 wire \Tile_X5Y4_E1BEG[1] ;
 wire \Tile_X5Y4_E1BEG[2] ;
 wire \Tile_X5Y4_E1BEG[3] ;
 wire \Tile_X5Y4_E2BEG[0] ;
 wire \Tile_X5Y4_E2BEG[1] ;
 wire \Tile_X5Y4_E2BEG[2] ;
 wire \Tile_X5Y4_E2BEG[3] ;
 wire \Tile_X5Y4_E2BEG[4] ;
 wire \Tile_X5Y4_E2BEG[5] ;
 wire \Tile_X5Y4_E2BEG[6] ;
 wire \Tile_X5Y4_E2BEG[7] ;
 wire \Tile_X5Y4_E2BEGb[0] ;
 wire \Tile_X5Y4_E2BEGb[1] ;
 wire \Tile_X5Y4_E2BEGb[2] ;
 wire \Tile_X5Y4_E2BEGb[3] ;
 wire \Tile_X5Y4_E2BEGb[4] ;
 wire \Tile_X5Y4_E2BEGb[5] ;
 wire \Tile_X5Y4_E2BEGb[6] ;
 wire \Tile_X5Y4_E2BEGb[7] ;
 wire \Tile_X5Y4_E6BEG[0] ;
 wire \Tile_X5Y4_E6BEG[10] ;
 wire \Tile_X5Y4_E6BEG[11] ;
 wire \Tile_X5Y4_E6BEG[1] ;
 wire \Tile_X5Y4_E6BEG[2] ;
 wire \Tile_X5Y4_E6BEG[3] ;
 wire \Tile_X5Y4_E6BEG[4] ;
 wire \Tile_X5Y4_E6BEG[5] ;
 wire \Tile_X5Y4_E6BEG[6] ;
 wire \Tile_X5Y4_E6BEG[7] ;
 wire \Tile_X5Y4_E6BEG[8] ;
 wire \Tile_X5Y4_E6BEG[9] ;
 wire \Tile_X5Y4_EE4BEG[0] ;
 wire \Tile_X5Y4_EE4BEG[10] ;
 wire \Tile_X5Y4_EE4BEG[11] ;
 wire \Tile_X5Y4_EE4BEG[12] ;
 wire \Tile_X5Y4_EE4BEG[13] ;
 wire \Tile_X5Y4_EE4BEG[14] ;
 wire \Tile_X5Y4_EE4BEG[15] ;
 wire \Tile_X5Y4_EE4BEG[1] ;
 wire \Tile_X5Y4_EE4BEG[2] ;
 wire \Tile_X5Y4_EE4BEG[3] ;
 wire \Tile_X5Y4_EE4BEG[4] ;
 wire \Tile_X5Y4_EE4BEG[5] ;
 wire \Tile_X5Y4_EE4BEG[6] ;
 wire \Tile_X5Y4_EE4BEG[7] ;
 wire \Tile_X5Y4_EE4BEG[8] ;
 wire \Tile_X5Y4_EE4BEG[9] ;
 wire \Tile_X5Y4_FrameData_O[0] ;
 wire \Tile_X5Y4_FrameData_O[10] ;
 wire \Tile_X5Y4_FrameData_O[11] ;
 wire \Tile_X5Y4_FrameData_O[12] ;
 wire \Tile_X5Y4_FrameData_O[13] ;
 wire \Tile_X5Y4_FrameData_O[14] ;
 wire \Tile_X5Y4_FrameData_O[15] ;
 wire \Tile_X5Y4_FrameData_O[16] ;
 wire \Tile_X5Y4_FrameData_O[17] ;
 wire \Tile_X5Y4_FrameData_O[18] ;
 wire \Tile_X5Y4_FrameData_O[19] ;
 wire \Tile_X5Y4_FrameData_O[1] ;
 wire \Tile_X5Y4_FrameData_O[20] ;
 wire \Tile_X5Y4_FrameData_O[21] ;
 wire \Tile_X5Y4_FrameData_O[22] ;
 wire \Tile_X5Y4_FrameData_O[23] ;
 wire \Tile_X5Y4_FrameData_O[24] ;
 wire \Tile_X5Y4_FrameData_O[25] ;
 wire \Tile_X5Y4_FrameData_O[26] ;
 wire \Tile_X5Y4_FrameData_O[27] ;
 wire \Tile_X5Y4_FrameData_O[28] ;
 wire \Tile_X5Y4_FrameData_O[29] ;
 wire \Tile_X5Y4_FrameData_O[2] ;
 wire \Tile_X5Y4_FrameData_O[30] ;
 wire \Tile_X5Y4_FrameData_O[31] ;
 wire \Tile_X5Y4_FrameData_O[3] ;
 wire \Tile_X5Y4_FrameData_O[4] ;
 wire \Tile_X5Y4_FrameData_O[5] ;
 wire \Tile_X5Y4_FrameData_O[6] ;
 wire \Tile_X5Y4_FrameData_O[7] ;
 wire \Tile_X5Y4_FrameData_O[8] ;
 wire \Tile_X5Y4_FrameData_O[9] ;
 wire \Tile_X5Y4_FrameStrobe_O[0] ;
 wire \Tile_X5Y4_FrameStrobe_O[10] ;
 wire \Tile_X5Y4_FrameStrobe_O[11] ;
 wire \Tile_X5Y4_FrameStrobe_O[12] ;
 wire \Tile_X5Y4_FrameStrobe_O[13] ;
 wire \Tile_X5Y4_FrameStrobe_O[14] ;
 wire \Tile_X5Y4_FrameStrobe_O[15] ;
 wire \Tile_X5Y4_FrameStrobe_O[16] ;
 wire \Tile_X5Y4_FrameStrobe_O[17] ;
 wire \Tile_X5Y4_FrameStrobe_O[18] ;
 wire \Tile_X5Y4_FrameStrobe_O[19] ;
 wire \Tile_X5Y4_FrameStrobe_O[1] ;
 wire \Tile_X5Y4_FrameStrobe_O[2] ;
 wire \Tile_X5Y4_FrameStrobe_O[3] ;
 wire \Tile_X5Y4_FrameStrobe_O[4] ;
 wire \Tile_X5Y4_FrameStrobe_O[5] ;
 wire \Tile_X5Y4_FrameStrobe_O[6] ;
 wire \Tile_X5Y4_FrameStrobe_O[7] ;
 wire \Tile_X5Y4_FrameStrobe_O[8] ;
 wire \Tile_X5Y4_FrameStrobe_O[9] ;
 wire \Tile_X5Y4_N1BEG[0] ;
 wire \Tile_X5Y4_N1BEG[1] ;
 wire \Tile_X5Y4_N1BEG[2] ;
 wire \Tile_X5Y4_N1BEG[3] ;
 wire \Tile_X5Y4_N2BEG[0] ;
 wire \Tile_X5Y4_N2BEG[1] ;
 wire \Tile_X5Y4_N2BEG[2] ;
 wire \Tile_X5Y4_N2BEG[3] ;
 wire \Tile_X5Y4_N2BEG[4] ;
 wire \Tile_X5Y4_N2BEG[5] ;
 wire \Tile_X5Y4_N2BEG[6] ;
 wire \Tile_X5Y4_N2BEG[7] ;
 wire \Tile_X5Y4_N2BEGb[0] ;
 wire \Tile_X5Y4_N2BEGb[1] ;
 wire \Tile_X5Y4_N2BEGb[2] ;
 wire \Tile_X5Y4_N2BEGb[3] ;
 wire \Tile_X5Y4_N2BEGb[4] ;
 wire \Tile_X5Y4_N2BEGb[5] ;
 wire \Tile_X5Y4_N2BEGb[6] ;
 wire \Tile_X5Y4_N2BEGb[7] ;
 wire \Tile_X5Y4_N4BEG[0] ;
 wire \Tile_X5Y4_N4BEG[10] ;
 wire \Tile_X5Y4_N4BEG[11] ;
 wire \Tile_X5Y4_N4BEG[12] ;
 wire \Tile_X5Y4_N4BEG[13] ;
 wire \Tile_X5Y4_N4BEG[14] ;
 wire \Tile_X5Y4_N4BEG[15] ;
 wire \Tile_X5Y4_N4BEG[1] ;
 wire \Tile_X5Y4_N4BEG[2] ;
 wire \Tile_X5Y4_N4BEG[3] ;
 wire \Tile_X5Y4_N4BEG[4] ;
 wire \Tile_X5Y4_N4BEG[5] ;
 wire \Tile_X5Y4_N4BEG[6] ;
 wire \Tile_X5Y4_N4BEG[7] ;
 wire \Tile_X5Y4_N4BEG[8] ;
 wire \Tile_X5Y4_N4BEG[9] ;
 wire \Tile_X5Y4_NN4BEG[0] ;
 wire \Tile_X5Y4_NN4BEG[10] ;
 wire \Tile_X5Y4_NN4BEG[11] ;
 wire \Tile_X5Y4_NN4BEG[12] ;
 wire \Tile_X5Y4_NN4BEG[13] ;
 wire \Tile_X5Y4_NN4BEG[14] ;
 wire \Tile_X5Y4_NN4BEG[15] ;
 wire \Tile_X5Y4_NN4BEG[1] ;
 wire \Tile_X5Y4_NN4BEG[2] ;
 wire \Tile_X5Y4_NN4BEG[3] ;
 wire \Tile_X5Y4_NN4BEG[4] ;
 wire \Tile_X5Y4_NN4BEG[5] ;
 wire \Tile_X5Y4_NN4BEG[6] ;
 wire \Tile_X5Y4_NN4BEG[7] ;
 wire \Tile_X5Y4_NN4BEG[8] ;
 wire \Tile_X5Y4_NN4BEG[9] ;
 wire \Tile_X5Y4_S1BEG[0] ;
 wire \Tile_X5Y4_S1BEG[1] ;
 wire \Tile_X5Y4_S1BEG[2] ;
 wire \Tile_X5Y4_S1BEG[3] ;
 wire \Tile_X5Y4_S2BEG[0] ;
 wire \Tile_X5Y4_S2BEG[1] ;
 wire \Tile_X5Y4_S2BEG[2] ;
 wire \Tile_X5Y4_S2BEG[3] ;
 wire \Tile_X5Y4_S2BEG[4] ;
 wire \Tile_X5Y4_S2BEG[5] ;
 wire \Tile_X5Y4_S2BEG[6] ;
 wire \Tile_X5Y4_S2BEG[7] ;
 wire \Tile_X5Y4_S2BEGb[0] ;
 wire \Tile_X5Y4_S2BEGb[1] ;
 wire \Tile_X5Y4_S2BEGb[2] ;
 wire \Tile_X5Y4_S2BEGb[3] ;
 wire \Tile_X5Y4_S2BEGb[4] ;
 wire \Tile_X5Y4_S2BEGb[5] ;
 wire \Tile_X5Y4_S2BEGb[6] ;
 wire \Tile_X5Y4_S2BEGb[7] ;
 wire \Tile_X5Y4_S4BEG[0] ;
 wire \Tile_X5Y4_S4BEG[10] ;
 wire \Tile_X5Y4_S4BEG[11] ;
 wire \Tile_X5Y4_S4BEG[12] ;
 wire \Tile_X5Y4_S4BEG[13] ;
 wire \Tile_X5Y4_S4BEG[14] ;
 wire \Tile_X5Y4_S4BEG[15] ;
 wire \Tile_X5Y4_S4BEG[1] ;
 wire \Tile_X5Y4_S4BEG[2] ;
 wire \Tile_X5Y4_S4BEG[3] ;
 wire \Tile_X5Y4_S4BEG[4] ;
 wire \Tile_X5Y4_S4BEG[5] ;
 wire \Tile_X5Y4_S4BEG[6] ;
 wire \Tile_X5Y4_S4BEG[7] ;
 wire \Tile_X5Y4_S4BEG[8] ;
 wire \Tile_X5Y4_S4BEG[9] ;
 wire \Tile_X5Y4_SS4BEG[0] ;
 wire \Tile_X5Y4_SS4BEG[10] ;
 wire \Tile_X5Y4_SS4BEG[11] ;
 wire \Tile_X5Y4_SS4BEG[12] ;
 wire \Tile_X5Y4_SS4BEG[13] ;
 wire \Tile_X5Y4_SS4BEG[14] ;
 wire \Tile_X5Y4_SS4BEG[15] ;
 wire \Tile_X5Y4_SS4BEG[1] ;
 wire \Tile_X5Y4_SS4BEG[2] ;
 wire \Tile_X5Y4_SS4BEG[3] ;
 wire \Tile_X5Y4_SS4BEG[4] ;
 wire \Tile_X5Y4_SS4BEG[5] ;
 wire \Tile_X5Y4_SS4BEG[6] ;
 wire \Tile_X5Y4_SS4BEG[7] ;
 wire \Tile_X5Y4_SS4BEG[8] ;
 wire \Tile_X5Y4_SS4BEG[9] ;
 wire Tile_X5Y4_UserCLKo;
 wire \Tile_X5Y4_W1BEG[0] ;
 wire \Tile_X5Y4_W1BEG[1] ;
 wire \Tile_X5Y4_W1BEG[2] ;
 wire \Tile_X5Y4_W1BEG[3] ;
 wire \Tile_X5Y4_W2BEG[0] ;
 wire \Tile_X5Y4_W2BEG[1] ;
 wire \Tile_X5Y4_W2BEG[2] ;
 wire \Tile_X5Y4_W2BEG[3] ;
 wire \Tile_X5Y4_W2BEG[4] ;
 wire \Tile_X5Y4_W2BEG[5] ;
 wire \Tile_X5Y4_W2BEG[6] ;
 wire \Tile_X5Y4_W2BEG[7] ;
 wire \Tile_X5Y4_W2BEGb[0] ;
 wire \Tile_X5Y4_W2BEGb[1] ;
 wire \Tile_X5Y4_W2BEGb[2] ;
 wire \Tile_X5Y4_W2BEGb[3] ;
 wire \Tile_X5Y4_W2BEGb[4] ;
 wire \Tile_X5Y4_W2BEGb[5] ;
 wire \Tile_X5Y4_W2BEGb[6] ;
 wire \Tile_X5Y4_W2BEGb[7] ;
 wire \Tile_X5Y4_W6BEG[0] ;
 wire \Tile_X5Y4_W6BEG[10] ;
 wire \Tile_X5Y4_W6BEG[11] ;
 wire \Tile_X5Y4_W6BEG[1] ;
 wire \Tile_X5Y4_W6BEG[2] ;
 wire \Tile_X5Y4_W6BEG[3] ;
 wire \Tile_X5Y4_W6BEG[4] ;
 wire \Tile_X5Y4_W6BEG[5] ;
 wire \Tile_X5Y4_W6BEG[6] ;
 wire \Tile_X5Y4_W6BEG[7] ;
 wire \Tile_X5Y4_W6BEG[8] ;
 wire \Tile_X5Y4_W6BEG[9] ;
 wire \Tile_X5Y4_WW4BEG[0] ;
 wire \Tile_X5Y4_WW4BEG[10] ;
 wire \Tile_X5Y4_WW4BEG[11] ;
 wire \Tile_X5Y4_WW4BEG[12] ;
 wire \Tile_X5Y4_WW4BEG[13] ;
 wire \Tile_X5Y4_WW4BEG[14] ;
 wire \Tile_X5Y4_WW4BEG[15] ;
 wire \Tile_X5Y4_WW4BEG[1] ;
 wire \Tile_X5Y4_WW4BEG[2] ;
 wire \Tile_X5Y4_WW4BEG[3] ;
 wire \Tile_X5Y4_WW4BEG[4] ;
 wire \Tile_X5Y4_WW4BEG[5] ;
 wire \Tile_X5Y4_WW4BEG[6] ;
 wire \Tile_X5Y4_WW4BEG[7] ;
 wire \Tile_X5Y4_WW4BEG[8] ;
 wire \Tile_X5Y4_WW4BEG[9] ;
 wire Tile_X5Y5_Co;
 wire \Tile_X5Y5_E1BEG[0] ;
 wire \Tile_X5Y5_E1BEG[1] ;
 wire \Tile_X5Y5_E1BEG[2] ;
 wire \Tile_X5Y5_E1BEG[3] ;
 wire \Tile_X5Y5_E2BEG[0] ;
 wire \Tile_X5Y5_E2BEG[1] ;
 wire \Tile_X5Y5_E2BEG[2] ;
 wire \Tile_X5Y5_E2BEG[3] ;
 wire \Tile_X5Y5_E2BEG[4] ;
 wire \Tile_X5Y5_E2BEG[5] ;
 wire \Tile_X5Y5_E2BEG[6] ;
 wire \Tile_X5Y5_E2BEG[7] ;
 wire \Tile_X5Y5_E2BEGb[0] ;
 wire \Tile_X5Y5_E2BEGb[1] ;
 wire \Tile_X5Y5_E2BEGb[2] ;
 wire \Tile_X5Y5_E2BEGb[3] ;
 wire \Tile_X5Y5_E2BEGb[4] ;
 wire \Tile_X5Y5_E2BEGb[5] ;
 wire \Tile_X5Y5_E2BEGb[6] ;
 wire \Tile_X5Y5_E2BEGb[7] ;
 wire \Tile_X5Y5_E6BEG[0] ;
 wire \Tile_X5Y5_E6BEG[10] ;
 wire \Tile_X5Y5_E6BEG[11] ;
 wire \Tile_X5Y5_E6BEG[1] ;
 wire \Tile_X5Y5_E6BEG[2] ;
 wire \Tile_X5Y5_E6BEG[3] ;
 wire \Tile_X5Y5_E6BEG[4] ;
 wire \Tile_X5Y5_E6BEG[5] ;
 wire \Tile_X5Y5_E6BEG[6] ;
 wire \Tile_X5Y5_E6BEG[7] ;
 wire \Tile_X5Y5_E6BEG[8] ;
 wire \Tile_X5Y5_E6BEG[9] ;
 wire \Tile_X5Y5_EE4BEG[0] ;
 wire \Tile_X5Y5_EE4BEG[10] ;
 wire \Tile_X5Y5_EE4BEG[11] ;
 wire \Tile_X5Y5_EE4BEG[12] ;
 wire \Tile_X5Y5_EE4BEG[13] ;
 wire \Tile_X5Y5_EE4BEG[14] ;
 wire \Tile_X5Y5_EE4BEG[15] ;
 wire \Tile_X5Y5_EE4BEG[1] ;
 wire \Tile_X5Y5_EE4BEG[2] ;
 wire \Tile_X5Y5_EE4BEG[3] ;
 wire \Tile_X5Y5_EE4BEG[4] ;
 wire \Tile_X5Y5_EE4BEG[5] ;
 wire \Tile_X5Y5_EE4BEG[6] ;
 wire \Tile_X5Y5_EE4BEG[7] ;
 wire \Tile_X5Y5_EE4BEG[8] ;
 wire \Tile_X5Y5_EE4BEG[9] ;
 wire \Tile_X5Y5_FrameData_O[0] ;
 wire \Tile_X5Y5_FrameData_O[10] ;
 wire \Tile_X5Y5_FrameData_O[11] ;
 wire \Tile_X5Y5_FrameData_O[12] ;
 wire \Tile_X5Y5_FrameData_O[13] ;
 wire \Tile_X5Y5_FrameData_O[14] ;
 wire \Tile_X5Y5_FrameData_O[15] ;
 wire \Tile_X5Y5_FrameData_O[16] ;
 wire \Tile_X5Y5_FrameData_O[17] ;
 wire \Tile_X5Y5_FrameData_O[18] ;
 wire \Tile_X5Y5_FrameData_O[19] ;
 wire \Tile_X5Y5_FrameData_O[1] ;
 wire \Tile_X5Y5_FrameData_O[20] ;
 wire \Tile_X5Y5_FrameData_O[21] ;
 wire \Tile_X5Y5_FrameData_O[22] ;
 wire \Tile_X5Y5_FrameData_O[23] ;
 wire \Tile_X5Y5_FrameData_O[24] ;
 wire \Tile_X5Y5_FrameData_O[25] ;
 wire \Tile_X5Y5_FrameData_O[26] ;
 wire \Tile_X5Y5_FrameData_O[27] ;
 wire \Tile_X5Y5_FrameData_O[28] ;
 wire \Tile_X5Y5_FrameData_O[29] ;
 wire \Tile_X5Y5_FrameData_O[2] ;
 wire \Tile_X5Y5_FrameData_O[30] ;
 wire \Tile_X5Y5_FrameData_O[31] ;
 wire \Tile_X5Y5_FrameData_O[3] ;
 wire \Tile_X5Y5_FrameData_O[4] ;
 wire \Tile_X5Y5_FrameData_O[5] ;
 wire \Tile_X5Y5_FrameData_O[6] ;
 wire \Tile_X5Y5_FrameData_O[7] ;
 wire \Tile_X5Y5_FrameData_O[8] ;
 wire \Tile_X5Y5_FrameData_O[9] ;
 wire \Tile_X5Y5_FrameStrobe_O[0] ;
 wire \Tile_X5Y5_FrameStrobe_O[10] ;
 wire \Tile_X5Y5_FrameStrobe_O[11] ;
 wire \Tile_X5Y5_FrameStrobe_O[12] ;
 wire \Tile_X5Y5_FrameStrobe_O[13] ;
 wire \Tile_X5Y5_FrameStrobe_O[14] ;
 wire \Tile_X5Y5_FrameStrobe_O[15] ;
 wire \Tile_X5Y5_FrameStrobe_O[16] ;
 wire \Tile_X5Y5_FrameStrobe_O[17] ;
 wire \Tile_X5Y5_FrameStrobe_O[18] ;
 wire \Tile_X5Y5_FrameStrobe_O[19] ;
 wire \Tile_X5Y5_FrameStrobe_O[1] ;
 wire \Tile_X5Y5_FrameStrobe_O[2] ;
 wire \Tile_X5Y5_FrameStrobe_O[3] ;
 wire \Tile_X5Y5_FrameStrobe_O[4] ;
 wire \Tile_X5Y5_FrameStrobe_O[5] ;
 wire \Tile_X5Y5_FrameStrobe_O[6] ;
 wire \Tile_X5Y5_FrameStrobe_O[7] ;
 wire \Tile_X5Y5_FrameStrobe_O[8] ;
 wire \Tile_X5Y5_FrameStrobe_O[9] ;
 wire \Tile_X5Y5_N1BEG[0] ;
 wire \Tile_X5Y5_N1BEG[1] ;
 wire \Tile_X5Y5_N1BEG[2] ;
 wire \Tile_X5Y5_N1BEG[3] ;
 wire \Tile_X5Y5_N2BEG[0] ;
 wire \Tile_X5Y5_N2BEG[1] ;
 wire \Tile_X5Y5_N2BEG[2] ;
 wire \Tile_X5Y5_N2BEG[3] ;
 wire \Tile_X5Y5_N2BEG[4] ;
 wire \Tile_X5Y5_N2BEG[5] ;
 wire \Tile_X5Y5_N2BEG[6] ;
 wire \Tile_X5Y5_N2BEG[7] ;
 wire \Tile_X5Y5_N2BEGb[0] ;
 wire \Tile_X5Y5_N2BEGb[1] ;
 wire \Tile_X5Y5_N2BEGb[2] ;
 wire \Tile_X5Y5_N2BEGb[3] ;
 wire \Tile_X5Y5_N2BEGb[4] ;
 wire \Tile_X5Y5_N2BEGb[5] ;
 wire \Tile_X5Y5_N2BEGb[6] ;
 wire \Tile_X5Y5_N2BEGb[7] ;
 wire \Tile_X5Y5_N4BEG[0] ;
 wire \Tile_X5Y5_N4BEG[10] ;
 wire \Tile_X5Y5_N4BEG[11] ;
 wire \Tile_X5Y5_N4BEG[12] ;
 wire \Tile_X5Y5_N4BEG[13] ;
 wire \Tile_X5Y5_N4BEG[14] ;
 wire \Tile_X5Y5_N4BEG[15] ;
 wire \Tile_X5Y5_N4BEG[1] ;
 wire \Tile_X5Y5_N4BEG[2] ;
 wire \Tile_X5Y5_N4BEG[3] ;
 wire \Tile_X5Y5_N4BEG[4] ;
 wire \Tile_X5Y5_N4BEG[5] ;
 wire \Tile_X5Y5_N4BEG[6] ;
 wire \Tile_X5Y5_N4BEG[7] ;
 wire \Tile_X5Y5_N4BEG[8] ;
 wire \Tile_X5Y5_N4BEG[9] ;
 wire \Tile_X5Y5_NN4BEG[0] ;
 wire \Tile_X5Y5_NN4BEG[10] ;
 wire \Tile_X5Y5_NN4BEG[11] ;
 wire \Tile_X5Y5_NN4BEG[12] ;
 wire \Tile_X5Y5_NN4BEG[13] ;
 wire \Tile_X5Y5_NN4BEG[14] ;
 wire \Tile_X5Y5_NN4BEG[15] ;
 wire \Tile_X5Y5_NN4BEG[1] ;
 wire \Tile_X5Y5_NN4BEG[2] ;
 wire \Tile_X5Y5_NN4BEG[3] ;
 wire \Tile_X5Y5_NN4BEG[4] ;
 wire \Tile_X5Y5_NN4BEG[5] ;
 wire \Tile_X5Y5_NN4BEG[6] ;
 wire \Tile_X5Y5_NN4BEG[7] ;
 wire \Tile_X5Y5_NN4BEG[8] ;
 wire \Tile_X5Y5_NN4BEG[9] ;
 wire \Tile_X5Y5_S1BEG[0] ;
 wire \Tile_X5Y5_S1BEG[1] ;
 wire \Tile_X5Y5_S1BEG[2] ;
 wire \Tile_X5Y5_S1BEG[3] ;
 wire \Tile_X5Y5_S2BEG[0] ;
 wire \Tile_X5Y5_S2BEG[1] ;
 wire \Tile_X5Y5_S2BEG[2] ;
 wire \Tile_X5Y5_S2BEG[3] ;
 wire \Tile_X5Y5_S2BEG[4] ;
 wire \Tile_X5Y5_S2BEG[5] ;
 wire \Tile_X5Y5_S2BEG[6] ;
 wire \Tile_X5Y5_S2BEG[7] ;
 wire \Tile_X5Y5_S2BEGb[0] ;
 wire \Tile_X5Y5_S2BEGb[1] ;
 wire \Tile_X5Y5_S2BEGb[2] ;
 wire \Tile_X5Y5_S2BEGb[3] ;
 wire \Tile_X5Y5_S2BEGb[4] ;
 wire \Tile_X5Y5_S2BEGb[5] ;
 wire \Tile_X5Y5_S2BEGb[6] ;
 wire \Tile_X5Y5_S2BEGb[7] ;
 wire \Tile_X5Y5_S4BEG[0] ;
 wire \Tile_X5Y5_S4BEG[10] ;
 wire \Tile_X5Y5_S4BEG[11] ;
 wire \Tile_X5Y5_S4BEG[12] ;
 wire \Tile_X5Y5_S4BEG[13] ;
 wire \Tile_X5Y5_S4BEG[14] ;
 wire \Tile_X5Y5_S4BEG[15] ;
 wire \Tile_X5Y5_S4BEG[1] ;
 wire \Tile_X5Y5_S4BEG[2] ;
 wire \Tile_X5Y5_S4BEG[3] ;
 wire \Tile_X5Y5_S4BEG[4] ;
 wire \Tile_X5Y5_S4BEG[5] ;
 wire \Tile_X5Y5_S4BEG[6] ;
 wire \Tile_X5Y5_S4BEG[7] ;
 wire \Tile_X5Y5_S4BEG[8] ;
 wire \Tile_X5Y5_S4BEG[9] ;
 wire \Tile_X5Y5_SS4BEG[0] ;
 wire \Tile_X5Y5_SS4BEG[10] ;
 wire \Tile_X5Y5_SS4BEG[11] ;
 wire \Tile_X5Y5_SS4BEG[12] ;
 wire \Tile_X5Y5_SS4BEG[13] ;
 wire \Tile_X5Y5_SS4BEG[14] ;
 wire \Tile_X5Y5_SS4BEG[15] ;
 wire \Tile_X5Y5_SS4BEG[1] ;
 wire \Tile_X5Y5_SS4BEG[2] ;
 wire \Tile_X5Y5_SS4BEG[3] ;
 wire \Tile_X5Y5_SS4BEG[4] ;
 wire \Tile_X5Y5_SS4BEG[5] ;
 wire \Tile_X5Y5_SS4BEG[6] ;
 wire \Tile_X5Y5_SS4BEG[7] ;
 wire \Tile_X5Y5_SS4BEG[8] ;
 wire \Tile_X5Y5_SS4BEG[9] ;
 wire Tile_X5Y5_UserCLKo;
 wire \Tile_X5Y5_W1BEG[0] ;
 wire \Tile_X5Y5_W1BEG[1] ;
 wire \Tile_X5Y5_W1BEG[2] ;
 wire \Tile_X5Y5_W1BEG[3] ;
 wire \Tile_X5Y5_W2BEG[0] ;
 wire \Tile_X5Y5_W2BEG[1] ;
 wire \Tile_X5Y5_W2BEG[2] ;
 wire \Tile_X5Y5_W2BEG[3] ;
 wire \Tile_X5Y5_W2BEG[4] ;
 wire \Tile_X5Y5_W2BEG[5] ;
 wire \Tile_X5Y5_W2BEG[6] ;
 wire \Tile_X5Y5_W2BEG[7] ;
 wire \Tile_X5Y5_W2BEGb[0] ;
 wire \Tile_X5Y5_W2BEGb[1] ;
 wire \Tile_X5Y5_W2BEGb[2] ;
 wire \Tile_X5Y5_W2BEGb[3] ;
 wire \Tile_X5Y5_W2BEGb[4] ;
 wire \Tile_X5Y5_W2BEGb[5] ;
 wire \Tile_X5Y5_W2BEGb[6] ;
 wire \Tile_X5Y5_W2BEGb[7] ;
 wire \Tile_X5Y5_W6BEG[0] ;
 wire \Tile_X5Y5_W6BEG[10] ;
 wire \Tile_X5Y5_W6BEG[11] ;
 wire \Tile_X5Y5_W6BEG[1] ;
 wire \Tile_X5Y5_W6BEG[2] ;
 wire \Tile_X5Y5_W6BEG[3] ;
 wire \Tile_X5Y5_W6BEG[4] ;
 wire \Tile_X5Y5_W6BEG[5] ;
 wire \Tile_X5Y5_W6BEG[6] ;
 wire \Tile_X5Y5_W6BEG[7] ;
 wire \Tile_X5Y5_W6BEG[8] ;
 wire \Tile_X5Y5_W6BEG[9] ;
 wire \Tile_X5Y5_WW4BEG[0] ;
 wire \Tile_X5Y5_WW4BEG[10] ;
 wire \Tile_X5Y5_WW4BEG[11] ;
 wire \Tile_X5Y5_WW4BEG[12] ;
 wire \Tile_X5Y5_WW4BEG[13] ;
 wire \Tile_X5Y5_WW4BEG[14] ;
 wire \Tile_X5Y5_WW4BEG[15] ;
 wire \Tile_X5Y5_WW4BEG[1] ;
 wire \Tile_X5Y5_WW4BEG[2] ;
 wire \Tile_X5Y5_WW4BEG[3] ;
 wire \Tile_X5Y5_WW4BEG[4] ;
 wire \Tile_X5Y5_WW4BEG[5] ;
 wire \Tile_X5Y5_WW4BEG[6] ;
 wire \Tile_X5Y5_WW4BEG[7] ;
 wire \Tile_X5Y5_WW4BEG[8] ;
 wire \Tile_X5Y5_WW4BEG[9] ;
 wire Tile_X5Y6_Co;
 wire \Tile_X5Y6_E1BEG[0] ;
 wire \Tile_X5Y6_E1BEG[1] ;
 wire \Tile_X5Y6_E1BEG[2] ;
 wire \Tile_X5Y6_E1BEG[3] ;
 wire \Tile_X5Y6_E2BEG[0] ;
 wire \Tile_X5Y6_E2BEG[1] ;
 wire \Tile_X5Y6_E2BEG[2] ;
 wire \Tile_X5Y6_E2BEG[3] ;
 wire \Tile_X5Y6_E2BEG[4] ;
 wire \Tile_X5Y6_E2BEG[5] ;
 wire \Tile_X5Y6_E2BEG[6] ;
 wire \Tile_X5Y6_E2BEG[7] ;
 wire \Tile_X5Y6_E2BEGb[0] ;
 wire \Tile_X5Y6_E2BEGb[1] ;
 wire \Tile_X5Y6_E2BEGb[2] ;
 wire \Tile_X5Y6_E2BEGb[3] ;
 wire \Tile_X5Y6_E2BEGb[4] ;
 wire \Tile_X5Y6_E2BEGb[5] ;
 wire \Tile_X5Y6_E2BEGb[6] ;
 wire \Tile_X5Y6_E2BEGb[7] ;
 wire \Tile_X5Y6_E6BEG[0] ;
 wire \Tile_X5Y6_E6BEG[10] ;
 wire \Tile_X5Y6_E6BEG[11] ;
 wire \Tile_X5Y6_E6BEG[1] ;
 wire \Tile_X5Y6_E6BEG[2] ;
 wire \Tile_X5Y6_E6BEG[3] ;
 wire \Tile_X5Y6_E6BEG[4] ;
 wire \Tile_X5Y6_E6BEG[5] ;
 wire \Tile_X5Y6_E6BEG[6] ;
 wire \Tile_X5Y6_E6BEG[7] ;
 wire \Tile_X5Y6_E6BEG[8] ;
 wire \Tile_X5Y6_E6BEG[9] ;
 wire \Tile_X5Y6_EE4BEG[0] ;
 wire \Tile_X5Y6_EE4BEG[10] ;
 wire \Tile_X5Y6_EE4BEG[11] ;
 wire \Tile_X5Y6_EE4BEG[12] ;
 wire \Tile_X5Y6_EE4BEG[13] ;
 wire \Tile_X5Y6_EE4BEG[14] ;
 wire \Tile_X5Y6_EE4BEG[15] ;
 wire \Tile_X5Y6_EE4BEG[1] ;
 wire \Tile_X5Y6_EE4BEG[2] ;
 wire \Tile_X5Y6_EE4BEG[3] ;
 wire \Tile_X5Y6_EE4BEG[4] ;
 wire \Tile_X5Y6_EE4BEG[5] ;
 wire \Tile_X5Y6_EE4BEG[6] ;
 wire \Tile_X5Y6_EE4BEG[7] ;
 wire \Tile_X5Y6_EE4BEG[8] ;
 wire \Tile_X5Y6_EE4BEG[9] ;
 wire \Tile_X5Y6_FrameData_O[0] ;
 wire \Tile_X5Y6_FrameData_O[10] ;
 wire \Tile_X5Y6_FrameData_O[11] ;
 wire \Tile_X5Y6_FrameData_O[12] ;
 wire \Tile_X5Y6_FrameData_O[13] ;
 wire \Tile_X5Y6_FrameData_O[14] ;
 wire \Tile_X5Y6_FrameData_O[15] ;
 wire \Tile_X5Y6_FrameData_O[16] ;
 wire \Tile_X5Y6_FrameData_O[17] ;
 wire \Tile_X5Y6_FrameData_O[18] ;
 wire \Tile_X5Y6_FrameData_O[19] ;
 wire \Tile_X5Y6_FrameData_O[1] ;
 wire \Tile_X5Y6_FrameData_O[20] ;
 wire \Tile_X5Y6_FrameData_O[21] ;
 wire \Tile_X5Y6_FrameData_O[22] ;
 wire \Tile_X5Y6_FrameData_O[23] ;
 wire \Tile_X5Y6_FrameData_O[24] ;
 wire \Tile_X5Y6_FrameData_O[25] ;
 wire \Tile_X5Y6_FrameData_O[26] ;
 wire \Tile_X5Y6_FrameData_O[27] ;
 wire \Tile_X5Y6_FrameData_O[28] ;
 wire \Tile_X5Y6_FrameData_O[29] ;
 wire \Tile_X5Y6_FrameData_O[2] ;
 wire \Tile_X5Y6_FrameData_O[30] ;
 wire \Tile_X5Y6_FrameData_O[31] ;
 wire \Tile_X5Y6_FrameData_O[3] ;
 wire \Tile_X5Y6_FrameData_O[4] ;
 wire \Tile_X5Y6_FrameData_O[5] ;
 wire \Tile_X5Y6_FrameData_O[6] ;
 wire \Tile_X5Y6_FrameData_O[7] ;
 wire \Tile_X5Y6_FrameData_O[8] ;
 wire \Tile_X5Y6_FrameData_O[9] ;
 wire \Tile_X5Y6_FrameStrobe_O[0] ;
 wire \Tile_X5Y6_FrameStrobe_O[10] ;
 wire \Tile_X5Y6_FrameStrobe_O[11] ;
 wire \Tile_X5Y6_FrameStrobe_O[12] ;
 wire \Tile_X5Y6_FrameStrobe_O[13] ;
 wire \Tile_X5Y6_FrameStrobe_O[14] ;
 wire \Tile_X5Y6_FrameStrobe_O[15] ;
 wire \Tile_X5Y6_FrameStrobe_O[16] ;
 wire \Tile_X5Y6_FrameStrobe_O[17] ;
 wire \Tile_X5Y6_FrameStrobe_O[18] ;
 wire \Tile_X5Y6_FrameStrobe_O[19] ;
 wire \Tile_X5Y6_FrameStrobe_O[1] ;
 wire \Tile_X5Y6_FrameStrobe_O[2] ;
 wire \Tile_X5Y6_FrameStrobe_O[3] ;
 wire \Tile_X5Y6_FrameStrobe_O[4] ;
 wire \Tile_X5Y6_FrameStrobe_O[5] ;
 wire \Tile_X5Y6_FrameStrobe_O[6] ;
 wire \Tile_X5Y6_FrameStrobe_O[7] ;
 wire \Tile_X5Y6_FrameStrobe_O[8] ;
 wire \Tile_X5Y6_FrameStrobe_O[9] ;
 wire \Tile_X5Y6_N1BEG[0] ;
 wire \Tile_X5Y6_N1BEG[1] ;
 wire \Tile_X5Y6_N1BEG[2] ;
 wire \Tile_X5Y6_N1BEG[3] ;
 wire \Tile_X5Y6_N2BEG[0] ;
 wire \Tile_X5Y6_N2BEG[1] ;
 wire \Tile_X5Y6_N2BEG[2] ;
 wire \Tile_X5Y6_N2BEG[3] ;
 wire \Tile_X5Y6_N2BEG[4] ;
 wire \Tile_X5Y6_N2BEG[5] ;
 wire \Tile_X5Y6_N2BEG[6] ;
 wire \Tile_X5Y6_N2BEG[7] ;
 wire \Tile_X5Y6_N2BEGb[0] ;
 wire \Tile_X5Y6_N2BEGb[1] ;
 wire \Tile_X5Y6_N2BEGb[2] ;
 wire \Tile_X5Y6_N2BEGb[3] ;
 wire \Tile_X5Y6_N2BEGb[4] ;
 wire \Tile_X5Y6_N2BEGb[5] ;
 wire \Tile_X5Y6_N2BEGb[6] ;
 wire \Tile_X5Y6_N2BEGb[7] ;
 wire \Tile_X5Y6_N4BEG[0] ;
 wire \Tile_X5Y6_N4BEG[10] ;
 wire \Tile_X5Y6_N4BEG[11] ;
 wire \Tile_X5Y6_N4BEG[12] ;
 wire \Tile_X5Y6_N4BEG[13] ;
 wire \Tile_X5Y6_N4BEG[14] ;
 wire \Tile_X5Y6_N4BEG[15] ;
 wire \Tile_X5Y6_N4BEG[1] ;
 wire \Tile_X5Y6_N4BEG[2] ;
 wire \Tile_X5Y6_N4BEG[3] ;
 wire \Tile_X5Y6_N4BEG[4] ;
 wire \Tile_X5Y6_N4BEG[5] ;
 wire \Tile_X5Y6_N4BEG[6] ;
 wire \Tile_X5Y6_N4BEG[7] ;
 wire \Tile_X5Y6_N4BEG[8] ;
 wire \Tile_X5Y6_N4BEG[9] ;
 wire \Tile_X5Y6_NN4BEG[0] ;
 wire \Tile_X5Y6_NN4BEG[10] ;
 wire \Tile_X5Y6_NN4BEG[11] ;
 wire \Tile_X5Y6_NN4BEG[12] ;
 wire \Tile_X5Y6_NN4BEG[13] ;
 wire \Tile_X5Y6_NN4BEG[14] ;
 wire \Tile_X5Y6_NN4BEG[15] ;
 wire \Tile_X5Y6_NN4BEG[1] ;
 wire \Tile_X5Y6_NN4BEG[2] ;
 wire \Tile_X5Y6_NN4BEG[3] ;
 wire \Tile_X5Y6_NN4BEG[4] ;
 wire \Tile_X5Y6_NN4BEG[5] ;
 wire \Tile_X5Y6_NN4BEG[6] ;
 wire \Tile_X5Y6_NN4BEG[7] ;
 wire \Tile_X5Y6_NN4BEG[8] ;
 wire \Tile_X5Y6_NN4BEG[9] ;
 wire \Tile_X5Y6_S1BEG[0] ;
 wire \Tile_X5Y6_S1BEG[1] ;
 wire \Tile_X5Y6_S1BEG[2] ;
 wire \Tile_X5Y6_S1BEG[3] ;
 wire \Tile_X5Y6_S2BEG[0] ;
 wire \Tile_X5Y6_S2BEG[1] ;
 wire \Tile_X5Y6_S2BEG[2] ;
 wire \Tile_X5Y6_S2BEG[3] ;
 wire \Tile_X5Y6_S2BEG[4] ;
 wire \Tile_X5Y6_S2BEG[5] ;
 wire \Tile_X5Y6_S2BEG[6] ;
 wire \Tile_X5Y6_S2BEG[7] ;
 wire \Tile_X5Y6_S2BEGb[0] ;
 wire \Tile_X5Y6_S2BEGb[1] ;
 wire \Tile_X5Y6_S2BEGb[2] ;
 wire \Tile_X5Y6_S2BEGb[3] ;
 wire \Tile_X5Y6_S2BEGb[4] ;
 wire \Tile_X5Y6_S2BEGb[5] ;
 wire \Tile_X5Y6_S2BEGb[6] ;
 wire \Tile_X5Y6_S2BEGb[7] ;
 wire \Tile_X5Y6_S4BEG[0] ;
 wire \Tile_X5Y6_S4BEG[10] ;
 wire \Tile_X5Y6_S4BEG[11] ;
 wire \Tile_X5Y6_S4BEG[12] ;
 wire \Tile_X5Y6_S4BEG[13] ;
 wire \Tile_X5Y6_S4BEG[14] ;
 wire \Tile_X5Y6_S4BEG[15] ;
 wire \Tile_X5Y6_S4BEG[1] ;
 wire \Tile_X5Y6_S4BEG[2] ;
 wire \Tile_X5Y6_S4BEG[3] ;
 wire \Tile_X5Y6_S4BEG[4] ;
 wire \Tile_X5Y6_S4BEG[5] ;
 wire \Tile_X5Y6_S4BEG[6] ;
 wire \Tile_X5Y6_S4BEG[7] ;
 wire \Tile_X5Y6_S4BEG[8] ;
 wire \Tile_X5Y6_S4BEG[9] ;
 wire \Tile_X5Y6_SS4BEG[0] ;
 wire \Tile_X5Y6_SS4BEG[10] ;
 wire \Tile_X5Y6_SS4BEG[11] ;
 wire \Tile_X5Y6_SS4BEG[12] ;
 wire \Tile_X5Y6_SS4BEG[13] ;
 wire \Tile_X5Y6_SS4BEG[14] ;
 wire \Tile_X5Y6_SS4BEG[15] ;
 wire \Tile_X5Y6_SS4BEG[1] ;
 wire \Tile_X5Y6_SS4BEG[2] ;
 wire \Tile_X5Y6_SS4BEG[3] ;
 wire \Tile_X5Y6_SS4BEG[4] ;
 wire \Tile_X5Y6_SS4BEG[5] ;
 wire \Tile_X5Y6_SS4BEG[6] ;
 wire \Tile_X5Y6_SS4BEG[7] ;
 wire \Tile_X5Y6_SS4BEG[8] ;
 wire \Tile_X5Y6_SS4BEG[9] ;
 wire Tile_X5Y6_UserCLKo;
 wire \Tile_X5Y6_W1BEG[0] ;
 wire \Tile_X5Y6_W1BEG[1] ;
 wire \Tile_X5Y6_W1BEG[2] ;
 wire \Tile_X5Y6_W1BEG[3] ;
 wire \Tile_X5Y6_W2BEG[0] ;
 wire \Tile_X5Y6_W2BEG[1] ;
 wire \Tile_X5Y6_W2BEG[2] ;
 wire \Tile_X5Y6_W2BEG[3] ;
 wire \Tile_X5Y6_W2BEG[4] ;
 wire \Tile_X5Y6_W2BEG[5] ;
 wire \Tile_X5Y6_W2BEG[6] ;
 wire \Tile_X5Y6_W2BEG[7] ;
 wire \Tile_X5Y6_W2BEGb[0] ;
 wire \Tile_X5Y6_W2BEGb[1] ;
 wire \Tile_X5Y6_W2BEGb[2] ;
 wire \Tile_X5Y6_W2BEGb[3] ;
 wire \Tile_X5Y6_W2BEGb[4] ;
 wire \Tile_X5Y6_W2BEGb[5] ;
 wire \Tile_X5Y6_W2BEGb[6] ;
 wire \Tile_X5Y6_W2BEGb[7] ;
 wire \Tile_X5Y6_W6BEG[0] ;
 wire \Tile_X5Y6_W6BEG[10] ;
 wire \Tile_X5Y6_W6BEG[11] ;
 wire \Tile_X5Y6_W6BEG[1] ;
 wire \Tile_X5Y6_W6BEG[2] ;
 wire \Tile_X5Y6_W6BEG[3] ;
 wire \Tile_X5Y6_W6BEG[4] ;
 wire \Tile_X5Y6_W6BEG[5] ;
 wire \Tile_X5Y6_W6BEG[6] ;
 wire \Tile_X5Y6_W6BEG[7] ;
 wire \Tile_X5Y6_W6BEG[8] ;
 wire \Tile_X5Y6_W6BEG[9] ;
 wire \Tile_X5Y6_WW4BEG[0] ;
 wire \Tile_X5Y6_WW4BEG[10] ;
 wire \Tile_X5Y6_WW4BEG[11] ;
 wire \Tile_X5Y6_WW4BEG[12] ;
 wire \Tile_X5Y6_WW4BEG[13] ;
 wire \Tile_X5Y6_WW4BEG[14] ;
 wire \Tile_X5Y6_WW4BEG[15] ;
 wire \Tile_X5Y6_WW4BEG[1] ;
 wire \Tile_X5Y6_WW4BEG[2] ;
 wire \Tile_X5Y6_WW4BEG[3] ;
 wire \Tile_X5Y6_WW4BEG[4] ;
 wire \Tile_X5Y6_WW4BEG[5] ;
 wire \Tile_X5Y6_WW4BEG[6] ;
 wire \Tile_X5Y6_WW4BEG[7] ;
 wire \Tile_X5Y6_WW4BEG[8] ;
 wire \Tile_X5Y6_WW4BEG[9] ;
 wire Tile_X5Y7_Co;
 wire \Tile_X5Y7_E1BEG[0] ;
 wire \Tile_X5Y7_E1BEG[1] ;
 wire \Tile_X5Y7_E1BEG[2] ;
 wire \Tile_X5Y7_E1BEG[3] ;
 wire \Tile_X5Y7_E2BEG[0] ;
 wire \Tile_X5Y7_E2BEG[1] ;
 wire \Tile_X5Y7_E2BEG[2] ;
 wire \Tile_X5Y7_E2BEG[3] ;
 wire \Tile_X5Y7_E2BEG[4] ;
 wire \Tile_X5Y7_E2BEG[5] ;
 wire \Tile_X5Y7_E2BEG[6] ;
 wire \Tile_X5Y7_E2BEG[7] ;
 wire \Tile_X5Y7_E2BEGb[0] ;
 wire \Tile_X5Y7_E2BEGb[1] ;
 wire \Tile_X5Y7_E2BEGb[2] ;
 wire \Tile_X5Y7_E2BEGb[3] ;
 wire \Tile_X5Y7_E2BEGb[4] ;
 wire \Tile_X5Y7_E2BEGb[5] ;
 wire \Tile_X5Y7_E2BEGb[6] ;
 wire \Tile_X5Y7_E2BEGb[7] ;
 wire \Tile_X5Y7_E6BEG[0] ;
 wire \Tile_X5Y7_E6BEG[10] ;
 wire \Tile_X5Y7_E6BEG[11] ;
 wire \Tile_X5Y7_E6BEG[1] ;
 wire \Tile_X5Y7_E6BEG[2] ;
 wire \Tile_X5Y7_E6BEG[3] ;
 wire \Tile_X5Y7_E6BEG[4] ;
 wire \Tile_X5Y7_E6BEG[5] ;
 wire \Tile_X5Y7_E6BEG[6] ;
 wire \Tile_X5Y7_E6BEG[7] ;
 wire \Tile_X5Y7_E6BEG[8] ;
 wire \Tile_X5Y7_E6BEG[9] ;
 wire \Tile_X5Y7_EE4BEG[0] ;
 wire \Tile_X5Y7_EE4BEG[10] ;
 wire \Tile_X5Y7_EE4BEG[11] ;
 wire \Tile_X5Y7_EE4BEG[12] ;
 wire \Tile_X5Y7_EE4BEG[13] ;
 wire \Tile_X5Y7_EE4BEG[14] ;
 wire \Tile_X5Y7_EE4BEG[15] ;
 wire \Tile_X5Y7_EE4BEG[1] ;
 wire \Tile_X5Y7_EE4BEG[2] ;
 wire \Tile_X5Y7_EE4BEG[3] ;
 wire \Tile_X5Y7_EE4BEG[4] ;
 wire \Tile_X5Y7_EE4BEG[5] ;
 wire \Tile_X5Y7_EE4BEG[6] ;
 wire \Tile_X5Y7_EE4BEG[7] ;
 wire \Tile_X5Y7_EE4BEG[8] ;
 wire \Tile_X5Y7_EE4BEG[9] ;
 wire \Tile_X5Y7_FrameData_O[0] ;
 wire \Tile_X5Y7_FrameData_O[10] ;
 wire \Tile_X5Y7_FrameData_O[11] ;
 wire \Tile_X5Y7_FrameData_O[12] ;
 wire \Tile_X5Y7_FrameData_O[13] ;
 wire \Tile_X5Y7_FrameData_O[14] ;
 wire \Tile_X5Y7_FrameData_O[15] ;
 wire \Tile_X5Y7_FrameData_O[16] ;
 wire \Tile_X5Y7_FrameData_O[17] ;
 wire \Tile_X5Y7_FrameData_O[18] ;
 wire \Tile_X5Y7_FrameData_O[19] ;
 wire \Tile_X5Y7_FrameData_O[1] ;
 wire \Tile_X5Y7_FrameData_O[20] ;
 wire \Tile_X5Y7_FrameData_O[21] ;
 wire \Tile_X5Y7_FrameData_O[22] ;
 wire \Tile_X5Y7_FrameData_O[23] ;
 wire \Tile_X5Y7_FrameData_O[24] ;
 wire \Tile_X5Y7_FrameData_O[25] ;
 wire \Tile_X5Y7_FrameData_O[26] ;
 wire \Tile_X5Y7_FrameData_O[27] ;
 wire \Tile_X5Y7_FrameData_O[28] ;
 wire \Tile_X5Y7_FrameData_O[29] ;
 wire \Tile_X5Y7_FrameData_O[2] ;
 wire \Tile_X5Y7_FrameData_O[30] ;
 wire \Tile_X5Y7_FrameData_O[31] ;
 wire \Tile_X5Y7_FrameData_O[3] ;
 wire \Tile_X5Y7_FrameData_O[4] ;
 wire \Tile_X5Y7_FrameData_O[5] ;
 wire \Tile_X5Y7_FrameData_O[6] ;
 wire \Tile_X5Y7_FrameData_O[7] ;
 wire \Tile_X5Y7_FrameData_O[8] ;
 wire \Tile_X5Y7_FrameData_O[9] ;
 wire \Tile_X5Y7_FrameStrobe_O[0] ;
 wire \Tile_X5Y7_FrameStrobe_O[10] ;
 wire \Tile_X5Y7_FrameStrobe_O[11] ;
 wire \Tile_X5Y7_FrameStrobe_O[12] ;
 wire \Tile_X5Y7_FrameStrobe_O[13] ;
 wire \Tile_X5Y7_FrameStrobe_O[14] ;
 wire \Tile_X5Y7_FrameStrobe_O[15] ;
 wire \Tile_X5Y7_FrameStrobe_O[16] ;
 wire \Tile_X5Y7_FrameStrobe_O[17] ;
 wire \Tile_X5Y7_FrameStrobe_O[18] ;
 wire \Tile_X5Y7_FrameStrobe_O[19] ;
 wire \Tile_X5Y7_FrameStrobe_O[1] ;
 wire \Tile_X5Y7_FrameStrobe_O[2] ;
 wire \Tile_X5Y7_FrameStrobe_O[3] ;
 wire \Tile_X5Y7_FrameStrobe_O[4] ;
 wire \Tile_X5Y7_FrameStrobe_O[5] ;
 wire \Tile_X5Y7_FrameStrobe_O[6] ;
 wire \Tile_X5Y7_FrameStrobe_O[7] ;
 wire \Tile_X5Y7_FrameStrobe_O[8] ;
 wire \Tile_X5Y7_FrameStrobe_O[9] ;
 wire \Tile_X5Y7_N1BEG[0] ;
 wire \Tile_X5Y7_N1BEG[1] ;
 wire \Tile_X5Y7_N1BEG[2] ;
 wire \Tile_X5Y7_N1BEG[3] ;
 wire \Tile_X5Y7_N2BEG[0] ;
 wire \Tile_X5Y7_N2BEG[1] ;
 wire \Tile_X5Y7_N2BEG[2] ;
 wire \Tile_X5Y7_N2BEG[3] ;
 wire \Tile_X5Y7_N2BEG[4] ;
 wire \Tile_X5Y7_N2BEG[5] ;
 wire \Tile_X5Y7_N2BEG[6] ;
 wire \Tile_X5Y7_N2BEG[7] ;
 wire \Tile_X5Y7_N2BEGb[0] ;
 wire \Tile_X5Y7_N2BEGb[1] ;
 wire \Tile_X5Y7_N2BEGb[2] ;
 wire \Tile_X5Y7_N2BEGb[3] ;
 wire \Tile_X5Y7_N2BEGb[4] ;
 wire \Tile_X5Y7_N2BEGb[5] ;
 wire \Tile_X5Y7_N2BEGb[6] ;
 wire \Tile_X5Y7_N2BEGb[7] ;
 wire \Tile_X5Y7_N4BEG[0] ;
 wire \Tile_X5Y7_N4BEG[10] ;
 wire \Tile_X5Y7_N4BEG[11] ;
 wire \Tile_X5Y7_N4BEG[12] ;
 wire \Tile_X5Y7_N4BEG[13] ;
 wire \Tile_X5Y7_N4BEG[14] ;
 wire \Tile_X5Y7_N4BEG[15] ;
 wire \Tile_X5Y7_N4BEG[1] ;
 wire \Tile_X5Y7_N4BEG[2] ;
 wire \Tile_X5Y7_N4BEG[3] ;
 wire \Tile_X5Y7_N4BEG[4] ;
 wire \Tile_X5Y7_N4BEG[5] ;
 wire \Tile_X5Y7_N4BEG[6] ;
 wire \Tile_X5Y7_N4BEG[7] ;
 wire \Tile_X5Y7_N4BEG[8] ;
 wire \Tile_X5Y7_N4BEG[9] ;
 wire \Tile_X5Y7_NN4BEG[0] ;
 wire \Tile_X5Y7_NN4BEG[10] ;
 wire \Tile_X5Y7_NN4BEG[11] ;
 wire \Tile_X5Y7_NN4BEG[12] ;
 wire \Tile_X5Y7_NN4BEG[13] ;
 wire \Tile_X5Y7_NN4BEG[14] ;
 wire \Tile_X5Y7_NN4BEG[15] ;
 wire \Tile_X5Y7_NN4BEG[1] ;
 wire \Tile_X5Y7_NN4BEG[2] ;
 wire \Tile_X5Y7_NN4BEG[3] ;
 wire \Tile_X5Y7_NN4BEG[4] ;
 wire \Tile_X5Y7_NN4BEG[5] ;
 wire \Tile_X5Y7_NN4BEG[6] ;
 wire \Tile_X5Y7_NN4BEG[7] ;
 wire \Tile_X5Y7_NN4BEG[8] ;
 wire \Tile_X5Y7_NN4BEG[9] ;
 wire \Tile_X5Y7_S1BEG[0] ;
 wire \Tile_X5Y7_S1BEG[1] ;
 wire \Tile_X5Y7_S1BEG[2] ;
 wire \Tile_X5Y7_S1BEG[3] ;
 wire \Tile_X5Y7_S2BEG[0] ;
 wire \Tile_X5Y7_S2BEG[1] ;
 wire \Tile_X5Y7_S2BEG[2] ;
 wire \Tile_X5Y7_S2BEG[3] ;
 wire \Tile_X5Y7_S2BEG[4] ;
 wire \Tile_X5Y7_S2BEG[5] ;
 wire \Tile_X5Y7_S2BEG[6] ;
 wire \Tile_X5Y7_S2BEG[7] ;
 wire \Tile_X5Y7_S2BEGb[0] ;
 wire \Tile_X5Y7_S2BEGb[1] ;
 wire \Tile_X5Y7_S2BEGb[2] ;
 wire \Tile_X5Y7_S2BEGb[3] ;
 wire \Tile_X5Y7_S2BEGb[4] ;
 wire \Tile_X5Y7_S2BEGb[5] ;
 wire \Tile_X5Y7_S2BEGb[6] ;
 wire \Tile_X5Y7_S2BEGb[7] ;
 wire \Tile_X5Y7_S4BEG[0] ;
 wire \Tile_X5Y7_S4BEG[10] ;
 wire \Tile_X5Y7_S4BEG[11] ;
 wire \Tile_X5Y7_S4BEG[12] ;
 wire \Tile_X5Y7_S4BEG[13] ;
 wire \Tile_X5Y7_S4BEG[14] ;
 wire \Tile_X5Y7_S4BEG[15] ;
 wire \Tile_X5Y7_S4BEG[1] ;
 wire \Tile_X5Y7_S4BEG[2] ;
 wire \Tile_X5Y7_S4BEG[3] ;
 wire \Tile_X5Y7_S4BEG[4] ;
 wire \Tile_X5Y7_S4BEG[5] ;
 wire \Tile_X5Y7_S4BEG[6] ;
 wire \Tile_X5Y7_S4BEG[7] ;
 wire \Tile_X5Y7_S4BEG[8] ;
 wire \Tile_X5Y7_S4BEG[9] ;
 wire \Tile_X5Y7_SS4BEG[0] ;
 wire \Tile_X5Y7_SS4BEG[10] ;
 wire \Tile_X5Y7_SS4BEG[11] ;
 wire \Tile_X5Y7_SS4BEG[12] ;
 wire \Tile_X5Y7_SS4BEG[13] ;
 wire \Tile_X5Y7_SS4BEG[14] ;
 wire \Tile_X5Y7_SS4BEG[15] ;
 wire \Tile_X5Y7_SS4BEG[1] ;
 wire \Tile_X5Y7_SS4BEG[2] ;
 wire \Tile_X5Y7_SS4BEG[3] ;
 wire \Tile_X5Y7_SS4BEG[4] ;
 wire \Tile_X5Y7_SS4BEG[5] ;
 wire \Tile_X5Y7_SS4BEG[6] ;
 wire \Tile_X5Y7_SS4BEG[7] ;
 wire \Tile_X5Y7_SS4BEG[8] ;
 wire \Tile_X5Y7_SS4BEG[9] ;
 wire Tile_X5Y7_UserCLKo;
 wire \Tile_X5Y7_W1BEG[0] ;
 wire \Tile_X5Y7_W1BEG[1] ;
 wire \Tile_X5Y7_W1BEG[2] ;
 wire \Tile_X5Y7_W1BEG[3] ;
 wire \Tile_X5Y7_W2BEG[0] ;
 wire \Tile_X5Y7_W2BEG[1] ;
 wire \Tile_X5Y7_W2BEG[2] ;
 wire \Tile_X5Y7_W2BEG[3] ;
 wire \Tile_X5Y7_W2BEG[4] ;
 wire \Tile_X5Y7_W2BEG[5] ;
 wire \Tile_X5Y7_W2BEG[6] ;
 wire \Tile_X5Y7_W2BEG[7] ;
 wire \Tile_X5Y7_W2BEGb[0] ;
 wire \Tile_X5Y7_W2BEGb[1] ;
 wire \Tile_X5Y7_W2BEGb[2] ;
 wire \Tile_X5Y7_W2BEGb[3] ;
 wire \Tile_X5Y7_W2BEGb[4] ;
 wire \Tile_X5Y7_W2BEGb[5] ;
 wire \Tile_X5Y7_W2BEGb[6] ;
 wire \Tile_X5Y7_W2BEGb[7] ;
 wire \Tile_X5Y7_W6BEG[0] ;
 wire \Tile_X5Y7_W6BEG[10] ;
 wire \Tile_X5Y7_W6BEG[11] ;
 wire \Tile_X5Y7_W6BEG[1] ;
 wire \Tile_X5Y7_W6BEG[2] ;
 wire \Tile_X5Y7_W6BEG[3] ;
 wire \Tile_X5Y7_W6BEG[4] ;
 wire \Tile_X5Y7_W6BEG[5] ;
 wire \Tile_X5Y7_W6BEG[6] ;
 wire \Tile_X5Y7_W6BEG[7] ;
 wire \Tile_X5Y7_W6BEG[8] ;
 wire \Tile_X5Y7_W6BEG[9] ;
 wire \Tile_X5Y7_WW4BEG[0] ;
 wire \Tile_X5Y7_WW4BEG[10] ;
 wire \Tile_X5Y7_WW4BEG[11] ;
 wire \Tile_X5Y7_WW4BEG[12] ;
 wire \Tile_X5Y7_WW4BEG[13] ;
 wire \Tile_X5Y7_WW4BEG[14] ;
 wire \Tile_X5Y7_WW4BEG[15] ;
 wire \Tile_X5Y7_WW4BEG[1] ;
 wire \Tile_X5Y7_WW4BEG[2] ;
 wire \Tile_X5Y7_WW4BEG[3] ;
 wire \Tile_X5Y7_WW4BEG[4] ;
 wire \Tile_X5Y7_WW4BEG[5] ;
 wire \Tile_X5Y7_WW4BEG[6] ;
 wire \Tile_X5Y7_WW4BEG[7] ;
 wire \Tile_X5Y7_WW4BEG[8] ;
 wire \Tile_X5Y7_WW4BEG[9] ;
 wire Tile_X5Y8_Co;
 wire \Tile_X5Y8_E1BEG[0] ;
 wire \Tile_X5Y8_E1BEG[1] ;
 wire \Tile_X5Y8_E1BEG[2] ;
 wire \Tile_X5Y8_E1BEG[3] ;
 wire \Tile_X5Y8_E2BEG[0] ;
 wire \Tile_X5Y8_E2BEG[1] ;
 wire \Tile_X5Y8_E2BEG[2] ;
 wire \Tile_X5Y8_E2BEG[3] ;
 wire \Tile_X5Y8_E2BEG[4] ;
 wire \Tile_X5Y8_E2BEG[5] ;
 wire \Tile_X5Y8_E2BEG[6] ;
 wire \Tile_X5Y8_E2BEG[7] ;
 wire \Tile_X5Y8_E2BEGb[0] ;
 wire \Tile_X5Y8_E2BEGb[1] ;
 wire \Tile_X5Y8_E2BEGb[2] ;
 wire \Tile_X5Y8_E2BEGb[3] ;
 wire \Tile_X5Y8_E2BEGb[4] ;
 wire \Tile_X5Y8_E2BEGb[5] ;
 wire \Tile_X5Y8_E2BEGb[6] ;
 wire \Tile_X5Y8_E2BEGb[7] ;
 wire \Tile_X5Y8_E6BEG[0] ;
 wire \Tile_X5Y8_E6BEG[10] ;
 wire \Tile_X5Y8_E6BEG[11] ;
 wire \Tile_X5Y8_E6BEG[1] ;
 wire \Tile_X5Y8_E6BEG[2] ;
 wire \Tile_X5Y8_E6BEG[3] ;
 wire \Tile_X5Y8_E6BEG[4] ;
 wire \Tile_X5Y8_E6BEG[5] ;
 wire \Tile_X5Y8_E6BEG[6] ;
 wire \Tile_X5Y8_E6BEG[7] ;
 wire \Tile_X5Y8_E6BEG[8] ;
 wire \Tile_X5Y8_E6BEG[9] ;
 wire \Tile_X5Y8_EE4BEG[0] ;
 wire \Tile_X5Y8_EE4BEG[10] ;
 wire \Tile_X5Y8_EE4BEG[11] ;
 wire \Tile_X5Y8_EE4BEG[12] ;
 wire \Tile_X5Y8_EE4BEG[13] ;
 wire \Tile_X5Y8_EE4BEG[14] ;
 wire \Tile_X5Y8_EE4BEG[15] ;
 wire \Tile_X5Y8_EE4BEG[1] ;
 wire \Tile_X5Y8_EE4BEG[2] ;
 wire \Tile_X5Y8_EE4BEG[3] ;
 wire \Tile_X5Y8_EE4BEG[4] ;
 wire \Tile_X5Y8_EE4BEG[5] ;
 wire \Tile_X5Y8_EE4BEG[6] ;
 wire \Tile_X5Y8_EE4BEG[7] ;
 wire \Tile_X5Y8_EE4BEG[8] ;
 wire \Tile_X5Y8_EE4BEG[9] ;
 wire \Tile_X5Y8_FrameData_O[0] ;
 wire \Tile_X5Y8_FrameData_O[10] ;
 wire \Tile_X5Y8_FrameData_O[11] ;
 wire \Tile_X5Y8_FrameData_O[12] ;
 wire \Tile_X5Y8_FrameData_O[13] ;
 wire \Tile_X5Y8_FrameData_O[14] ;
 wire \Tile_X5Y8_FrameData_O[15] ;
 wire \Tile_X5Y8_FrameData_O[16] ;
 wire \Tile_X5Y8_FrameData_O[17] ;
 wire \Tile_X5Y8_FrameData_O[18] ;
 wire \Tile_X5Y8_FrameData_O[19] ;
 wire \Tile_X5Y8_FrameData_O[1] ;
 wire \Tile_X5Y8_FrameData_O[20] ;
 wire \Tile_X5Y8_FrameData_O[21] ;
 wire \Tile_X5Y8_FrameData_O[22] ;
 wire \Tile_X5Y8_FrameData_O[23] ;
 wire \Tile_X5Y8_FrameData_O[24] ;
 wire \Tile_X5Y8_FrameData_O[25] ;
 wire \Tile_X5Y8_FrameData_O[26] ;
 wire \Tile_X5Y8_FrameData_O[27] ;
 wire \Tile_X5Y8_FrameData_O[28] ;
 wire \Tile_X5Y8_FrameData_O[29] ;
 wire \Tile_X5Y8_FrameData_O[2] ;
 wire \Tile_X5Y8_FrameData_O[30] ;
 wire \Tile_X5Y8_FrameData_O[31] ;
 wire \Tile_X5Y8_FrameData_O[3] ;
 wire \Tile_X5Y8_FrameData_O[4] ;
 wire \Tile_X5Y8_FrameData_O[5] ;
 wire \Tile_X5Y8_FrameData_O[6] ;
 wire \Tile_X5Y8_FrameData_O[7] ;
 wire \Tile_X5Y8_FrameData_O[8] ;
 wire \Tile_X5Y8_FrameData_O[9] ;
 wire \Tile_X5Y8_FrameStrobe_O[0] ;
 wire \Tile_X5Y8_FrameStrobe_O[10] ;
 wire \Tile_X5Y8_FrameStrobe_O[11] ;
 wire \Tile_X5Y8_FrameStrobe_O[12] ;
 wire \Tile_X5Y8_FrameStrobe_O[13] ;
 wire \Tile_X5Y8_FrameStrobe_O[14] ;
 wire \Tile_X5Y8_FrameStrobe_O[15] ;
 wire \Tile_X5Y8_FrameStrobe_O[16] ;
 wire \Tile_X5Y8_FrameStrobe_O[17] ;
 wire \Tile_X5Y8_FrameStrobe_O[18] ;
 wire \Tile_X5Y8_FrameStrobe_O[19] ;
 wire \Tile_X5Y8_FrameStrobe_O[1] ;
 wire \Tile_X5Y8_FrameStrobe_O[2] ;
 wire \Tile_X5Y8_FrameStrobe_O[3] ;
 wire \Tile_X5Y8_FrameStrobe_O[4] ;
 wire \Tile_X5Y8_FrameStrobe_O[5] ;
 wire \Tile_X5Y8_FrameStrobe_O[6] ;
 wire \Tile_X5Y8_FrameStrobe_O[7] ;
 wire \Tile_X5Y8_FrameStrobe_O[8] ;
 wire \Tile_X5Y8_FrameStrobe_O[9] ;
 wire \Tile_X5Y8_N1BEG[0] ;
 wire \Tile_X5Y8_N1BEG[1] ;
 wire \Tile_X5Y8_N1BEG[2] ;
 wire \Tile_X5Y8_N1BEG[3] ;
 wire \Tile_X5Y8_N2BEG[0] ;
 wire \Tile_X5Y8_N2BEG[1] ;
 wire \Tile_X5Y8_N2BEG[2] ;
 wire \Tile_X5Y8_N2BEG[3] ;
 wire \Tile_X5Y8_N2BEG[4] ;
 wire \Tile_X5Y8_N2BEG[5] ;
 wire \Tile_X5Y8_N2BEG[6] ;
 wire \Tile_X5Y8_N2BEG[7] ;
 wire \Tile_X5Y8_N2BEGb[0] ;
 wire \Tile_X5Y8_N2BEGb[1] ;
 wire \Tile_X5Y8_N2BEGb[2] ;
 wire \Tile_X5Y8_N2BEGb[3] ;
 wire \Tile_X5Y8_N2BEGb[4] ;
 wire \Tile_X5Y8_N2BEGb[5] ;
 wire \Tile_X5Y8_N2BEGb[6] ;
 wire \Tile_X5Y8_N2BEGb[7] ;
 wire \Tile_X5Y8_N4BEG[0] ;
 wire \Tile_X5Y8_N4BEG[10] ;
 wire \Tile_X5Y8_N4BEG[11] ;
 wire \Tile_X5Y8_N4BEG[12] ;
 wire \Tile_X5Y8_N4BEG[13] ;
 wire \Tile_X5Y8_N4BEG[14] ;
 wire \Tile_X5Y8_N4BEG[15] ;
 wire \Tile_X5Y8_N4BEG[1] ;
 wire \Tile_X5Y8_N4BEG[2] ;
 wire \Tile_X5Y8_N4BEG[3] ;
 wire \Tile_X5Y8_N4BEG[4] ;
 wire \Tile_X5Y8_N4BEG[5] ;
 wire \Tile_X5Y8_N4BEG[6] ;
 wire \Tile_X5Y8_N4BEG[7] ;
 wire \Tile_X5Y8_N4BEG[8] ;
 wire \Tile_X5Y8_N4BEG[9] ;
 wire \Tile_X5Y8_NN4BEG[0] ;
 wire \Tile_X5Y8_NN4BEG[10] ;
 wire \Tile_X5Y8_NN4BEG[11] ;
 wire \Tile_X5Y8_NN4BEG[12] ;
 wire \Tile_X5Y8_NN4BEG[13] ;
 wire \Tile_X5Y8_NN4BEG[14] ;
 wire \Tile_X5Y8_NN4BEG[15] ;
 wire \Tile_X5Y8_NN4BEG[1] ;
 wire \Tile_X5Y8_NN4BEG[2] ;
 wire \Tile_X5Y8_NN4BEG[3] ;
 wire \Tile_X5Y8_NN4BEG[4] ;
 wire \Tile_X5Y8_NN4BEG[5] ;
 wire \Tile_X5Y8_NN4BEG[6] ;
 wire \Tile_X5Y8_NN4BEG[7] ;
 wire \Tile_X5Y8_NN4BEG[8] ;
 wire \Tile_X5Y8_NN4BEG[9] ;
 wire \Tile_X5Y8_S1BEG[0] ;
 wire \Tile_X5Y8_S1BEG[1] ;
 wire \Tile_X5Y8_S1BEG[2] ;
 wire \Tile_X5Y8_S1BEG[3] ;
 wire \Tile_X5Y8_S2BEG[0] ;
 wire \Tile_X5Y8_S2BEG[1] ;
 wire \Tile_X5Y8_S2BEG[2] ;
 wire \Tile_X5Y8_S2BEG[3] ;
 wire \Tile_X5Y8_S2BEG[4] ;
 wire \Tile_X5Y8_S2BEG[5] ;
 wire \Tile_X5Y8_S2BEG[6] ;
 wire \Tile_X5Y8_S2BEG[7] ;
 wire \Tile_X5Y8_S2BEGb[0] ;
 wire \Tile_X5Y8_S2BEGb[1] ;
 wire \Tile_X5Y8_S2BEGb[2] ;
 wire \Tile_X5Y8_S2BEGb[3] ;
 wire \Tile_X5Y8_S2BEGb[4] ;
 wire \Tile_X5Y8_S2BEGb[5] ;
 wire \Tile_X5Y8_S2BEGb[6] ;
 wire \Tile_X5Y8_S2BEGb[7] ;
 wire \Tile_X5Y8_S4BEG[0] ;
 wire \Tile_X5Y8_S4BEG[10] ;
 wire \Tile_X5Y8_S4BEG[11] ;
 wire \Tile_X5Y8_S4BEG[12] ;
 wire \Tile_X5Y8_S4BEG[13] ;
 wire \Tile_X5Y8_S4BEG[14] ;
 wire \Tile_X5Y8_S4BEG[15] ;
 wire \Tile_X5Y8_S4BEG[1] ;
 wire \Tile_X5Y8_S4BEG[2] ;
 wire \Tile_X5Y8_S4BEG[3] ;
 wire \Tile_X5Y8_S4BEG[4] ;
 wire \Tile_X5Y8_S4BEG[5] ;
 wire \Tile_X5Y8_S4BEG[6] ;
 wire \Tile_X5Y8_S4BEG[7] ;
 wire \Tile_X5Y8_S4BEG[8] ;
 wire \Tile_X5Y8_S4BEG[9] ;
 wire \Tile_X5Y8_SS4BEG[0] ;
 wire \Tile_X5Y8_SS4BEG[10] ;
 wire \Tile_X5Y8_SS4BEG[11] ;
 wire \Tile_X5Y8_SS4BEG[12] ;
 wire \Tile_X5Y8_SS4BEG[13] ;
 wire \Tile_X5Y8_SS4BEG[14] ;
 wire \Tile_X5Y8_SS4BEG[15] ;
 wire \Tile_X5Y8_SS4BEG[1] ;
 wire \Tile_X5Y8_SS4BEG[2] ;
 wire \Tile_X5Y8_SS4BEG[3] ;
 wire \Tile_X5Y8_SS4BEG[4] ;
 wire \Tile_X5Y8_SS4BEG[5] ;
 wire \Tile_X5Y8_SS4BEG[6] ;
 wire \Tile_X5Y8_SS4BEG[7] ;
 wire \Tile_X5Y8_SS4BEG[8] ;
 wire \Tile_X5Y8_SS4BEG[9] ;
 wire Tile_X5Y8_UserCLKo;
 wire \Tile_X5Y8_W1BEG[0] ;
 wire \Tile_X5Y8_W1BEG[1] ;
 wire \Tile_X5Y8_W1BEG[2] ;
 wire \Tile_X5Y8_W1BEG[3] ;
 wire \Tile_X5Y8_W2BEG[0] ;
 wire \Tile_X5Y8_W2BEG[1] ;
 wire \Tile_X5Y8_W2BEG[2] ;
 wire \Tile_X5Y8_W2BEG[3] ;
 wire \Tile_X5Y8_W2BEG[4] ;
 wire \Tile_X5Y8_W2BEG[5] ;
 wire \Tile_X5Y8_W2BEG[6] ;
 wire \Tile_X5Y8_W2BEG[7] ;
 wire \Tile_X5Y8_W2BEGb[0] ;
 wire \Tile_X5Y8_W2BEGb[1] ;
 wire \Tile_X5Y8_W2BEGb[2] ;
 wire \Tile_X5Y8_W2BEGb[3] ;
 wire \Tile_X5Y8_W2BEGb[4] ;
 wire \Tile_X5Y8_W2BEGb[5] ;
 wire \Tile_X5Y8_W2BEGb[6] ;
 wire \Tile_X5Y8_W2BEGb[7] ;
 wire \Tile_X5Y8_W6BEG[0] ;
 wire \Tile_X5Y8_W6BEG[10] ;
 wire \Tile_X5Y8_W6BEG[11] ;
 wire \Tile_X5Y8_W6BEG[1] ;
 wire \Tile_X5Y8_W6BEG[2] ;
 wire \Tile_X5Y8_W6BEG[3] ;
 wire \Tile_X5Y8_W6BEG[4] ;
 wire \Tile_X5Y8_W6BEG[5] ;
 wire \Tile_X5Y8_W6BEG[6] ;
 wire \Tile_X5Y8_W6BEG[7] ;
 wire \Tile_X5Y8_W6BEG[8] ;
 wire \Tile_X5Y8_W6BEG[9] ;
 wire \Tile_X5Y8_WW4BEG[0] ;
 wire \Tile_X5Y8_WW4BEG[10] ;
 wire \Tile_X5Y8_WW4BEG[11] ;
 wire \Tile_X5Y8_WW4BEG[12] ;
 wire \Tile_X5Y8_WW4BEG[13] ;
 wire \Tile_X5Y8_WW4BEG[14] ;
 wire \Tile_X5Y8_WW4BEG[15] ;
 wire \Tile_X5Y8_WW4BEG[1] ;
 wire \Tile_X5Y8_WW4BEG[2] ;
 wire \Tile_X5Y8_WW4BEG[3] ;
 wire \Tile_X5Y8_WW4BEG[4] ;
 wire \Tile_X5Y8_WW4BEG[5] ;
 wire \Tile_X5Y8_WW4BEG[6] ;
 wire \Tile_X5Y8_WW4BEG[7] ;
 wire \Tile_X5Y8_WW4BEG[8] ;
 wire \Tile_X5Y8_WW4BEG[9] ;
 wire Tile_X5Y9_Co;
 wire \Tile_X5Y9_E1BEG[0] ;
 wire \Tile_X5Y9_E1BEG[1] ;
 wire \Tile_X5Y9_E1BEG[2] ;
 wire \Tile_X5Y9_E1BEG[3] ;
 wire \Tile_X5Y9_E2BEG[0] ;
 wire \Tile_X5Y9_E2BEG[1] ;
 wire \Tile_X5Y9_E2BEG[2] ;
 wire \Tile_X5Y9_E2BEG[3] ;
 wire \Tile_X5Y9_E2BEG[4] ;
 wire \Tile_X5Y9_E2BEG[5] ;
 wire \Tile_X5Y9_E2BEG[6] ;
 wire \Tile_X5Y9_E2BEG[7] ;
 wire \Tile_X5Y9_E2BEGb[0] ;
 wire \Tile_X5Y9_E2BEGb[1] ;
 wire \Tile_X5Y9_E2BEGb[2] ;
 wire \Tile_X5Y9_E2BEGb[3] ;
 wire \Tile_X5Y9_E2BEGb[4] ;
 wire \Tile_X5Y9_E2BEGb[5] ;
 wire \Tile_X5Y9_E2BEGb[6] ;
 wire \Tile_X5Y9_E2BEGb[7] ;
 wire \Tile_X5Y9_E6BEG[0] ;
 wire \Tile_X5Y9_E6BEG[10] ;
 wire \Tile_X5Y9_E6BEG[11] ;
 wire \Tile_X5Y9_E6BEG[1] ;
 wire \Tile_X5Y9_E6BEG[2] ;
 wire \Tile_X5Y9_E6BEG[3] ;
 wire \Tile_X5Y9_E6BEG[4] ;
 wire \Tile_X5Y9_E6BEG[5] ;
 wire \Tile_X5Y9_E6BEG[6] ;
 wire \Tile_X5Y9_E6BEG[7] ;
 wire \Tile_X5Y9_E6BEG[8] ;
 wire \Tile_X5Y9_E6BEG[9] ;
 wire \Tile_X5Y9_EE4BEG[0] ;
 wire \Tile_X5Y9_EE4BEG[10] ;
 wire \Tile_X5Y9_EE4BEG[11] ;
 wire \Tile_X5Y9_EE4BEG[12] ;
 wire \Tile_X5Y9_EE4BEG[13] ;
 wire \Tile_X5Y9_EE4BEG[14] ;
 wire \Tile_X5Y9_EE4BEG[15] ;
 wire \Tile_X5Y9_EE4BEG[1] ;
 wire \Tile_X5Y9_EE4BEG[2] ;
 wire \Tile_X5Y9_EE4BEG[3] ;
 wire \Tile_X5Y9_EE4BEG[4] ;
 wire \Tile_X5Y9_EE4BEG[5] ;
 wire \Tile_X5Y9_EE4BEG[6] ;
 wire \Tile_X5Y9_EE4BEG[7] ;
 wire \Tile_X5Y9_EE4BEG[8] ;
 wire \Tile_X5Y9_EE4BEG[9] ;
 wire \Tile_X5Y9_FrameData_O[0] ;
 wire \Tile_X5Y9_FrameData_O[10] ;
 wire \Tile_X5Y9_FrameData_O[11] ;
 wire \Tile_X5Y9_FrameData_O[12] ;
 wire \Tile_X5Y9_FrameData_O[13] ;
 wire \Tile_X5Y9_FrameData_O[14] ;
 wire \Tile_X5Y9_FrameData_O[15] ;
 wire \Tile_X5Y9_FrameData_O[16] ;
 wire \Tile_X5Y9_FrameData_O[17] ;
 wire \Tile_X5Y9_FrameData_O[18] ;
 wire \Tile_X5Y9_FrameData_O[19] ;
 wire \Tile_X5Y9_FrameData_O[1] ;
 wire \Tile_X5Y9_FrameData_O[20] ;
 wire \Tile_X5Y9_FrameData_O[21] ;
 wire \Tile_X5Y9_FrameData_O[22] ;
 wire \Tile_X5Y9_FrameData_O[23] ;
 wire \Tile_X5Y9_FrameData_O[24] ;
 wire \Tile_X5Y9_FrameData_O[25] ;
 wire \Tile_X5Y9_FrameData_O[26] ;
 wire \Tile_X5Y9_FrameData_O[27] ;
 wire \Tile_X5Y9_FrameData_O[28] ;
 wire \Tile_X5Y9_FrameData_O[29] ;
 wire \Tile_X5Y9_FrameData_O[2] ;
 wire \Tile_X5Y9_FrameData_O[30] ;
 wire \Tile_X5Y9_FrameData_O[31] ;
 wire \Tile_X5Y9_FrameData_O[3] ;
 wire \Tile_X5Y9_FrameData_O[4] ;
 wire \Tile_X5Y9_FrameData_O[5] ;
 wire \Tile_X5Y9_FrameData_O[6] ;
 wire \Tile_X5Y9_FrameData_O[7] ;
 wire \Tile_X5Y9_FrameData_O[8] ;
 wire \Tile_X5Y9_FrameData_O[9] ;
 wire \Tile_X5Y9_FrameStrobe_O[0] ;
 wire \Tile_X5Y9_FrameStrobe_O[10] ;
 wire \Tile_X5Y9_FrameStrobe_O[11] ;
 wire \Tile_X5Y9_FrameStrobe_O[12] ;
 wire \Tile_X5Y9_FrameStrobe_O[13] ;
 wire \Tile_X5Y9_FrameStrobe_O[14] ;
 wire \Tile_X5Y9_FrameStrobe_O[15] ;
 wire \Tile_X5Y9_FrameStrobe_O[16] ;
 wire \Tile_X5Y9_FrameStrobe_O[17] ;
 wire \Tile_X5Y9_FrameStrobe_O[18] ;
 wire \Tile_X5Y9_FrameStrobe_O[19] ;
 wire \Tile_X5Y9_FrameStrobe_O[1] ;
 wire \Tile_X5Y9_FrameStrobe_O[2] ;
 wire \Tile_X5Y9_FrameStrobe_O[3] ;
 wire \Tile_X5Y9_FrameStrobe_O[4] ;
 wire \Tile_X5Y9_FrameStrobe_O[5] ;
 wire \Tile_X5Y9_FrameStrobe_O[6] ;
 wire \Tile_X5Y9_FrameStrobe_O[7] ;
 wire \Tile_X5Y9_FrameStrobe_O[8] ;
 wire \Tile_X5Y9_FrameStrobe_O[9] ;
 wire \Tile_X5Y9_N1BEG[0] ;
 wire \Tile_X5Y9_N1BEG[1] ;
 wire \Tile_X5Y9_N1BEG[2] ;
 wire \Tile_X5Y9_N1BEG[3] ;
 wire \Tile_X5Y9_N2BEG[0] ;
 wire \Tile_X5Y9_N2BEG[1] ;
 wire \Tile_X5Y9_N2BEG[2] ;
 wire \Tile_X5Y9_N2BEG[3] ;
 wire \Tile_X5Y9_N2BEG[4] ;
 wire \Tile_X5Y9_N2BEG[5] ;
 wire \Tile_X5Y9_N2BEG[6] ;
 wire \Tile_X5Y9_N2BEG[7] ;
 wire \Tile_X5Y9_N2BEGb[0] ;
 wire \Tile_X5Y9_N2BEGb[1] ;
 wire \Tile_X5Y9_N2BEGb[2] ;
 wire \Tile_X5Y9_N2BEGb[3] ;
 wire \Tile_X5Y9_N2BEGb[4] ;
 wire \Tile_X5Y9_N2BEGb[5] ;
 wire \Tile_X5Y9_N2BEGb[6] ;
 wire \Tile_X5Y9_N2BEGb[7] ;
 wire \Tile_X5Y9_N4BEG[0] ;
 wire \Tile_X5Y9_N4BEG[10] ;
 wire \Tile_X5Y9_N4BEG[11] ;
 wire \Tile_X5Y9_N4BEG[12] ;
 wire \Tile_X5Y9_N4BEG[13] ;
 wire \Tile_X5Y9_N4BEG[14] ;
 wire \Tile_X5Y9_N4BEG[15] ;
 wire \Tile_X5Y9_N4BEG[1] ;
 wire \Tile_X5Y9_N4BEG[2] ;
 wire \Tile_X5Y9_N4BEG[3] ;
 wire \Tile_X5Y9_N4BEG[4] ;
 wire \Tile_X5Y9_N4BEG[5] ;
 wire \Tile_X5Y9_N4BEG[6] ;
 wire \Tile_X5Y9_N4BEG[7] ;
 wire \Tile_X5Y9_N4BEG[8] ;
 wire \Tile_X5Y9_N4BEG[9] ;
 wire \Tile_X5Y9_NN4BEG[0] ;
 wire \Tile_X5Y9_NN4BEG[10] ;
 wire \Tile_X5Y9_NN4BEG[11] ;
 wire \Tile_X5Y9_NN4BEG[12] ;
 wire \Tile_X5Y9_NN4BEG[13] ;
 wire \Tile_X5Y9_NN4BEG[14] ;
 wire \Tile_X5Y9_NN4BEG[15] ;
 wire \Tile_X5Y9_NN4BEG[1] ;
 wire \Tile_X5Y9_NN4BEG[2] ;
 wire \Tile_X5Y9_NN4BEG[3] ;
 wire \Tile_X5Y9_NN4BEG[4] ;
 wire \Tile_X5Y9_NN4BEG[5] ;
 wire \Tile_X5Y9_NN4BEG[6] ;
 wire \Tile_X5Y9_NN4BEG[7] ;
 wire \Tile_X5Y9_NN4BEG[8] ;
 wire \Tile_X5Y9_NN4BEG[9] ;
 wire \Tile_X5Y9_S1BEG[0] ;
 wire \Tile_X5Y9_S1BEG[1] ;
 wire \Tile_X5Y9_S1BEG[2] ;
 wire \Tile_X5Y9_S1BEG[3] ;
 wire \Tile_X5Y9_S2BEG[0] ;
 wire \Tile_X5Y9_S2BEG[1] ;
 wire \Tile_X5Y9_S2BEG[2] ;
 wire \Tile_X5Y9_S2BEG[3] ;
 wire \Tile_X5Y9_S2BEG[4] ;
 wire \Tile_X5Y9_S2BEG[5] ;
 wire \Tile_X5Y9_S2BEG[6] ;
 wire \Tile_X5Y9_S2BEG[7] ;
 wire \Tile_X5Y9_S2BEGb[0] ;
 wire \Tile_X5Y9_S2BEGb[1] ;
 wire \Tile_X5Y9_S2BEGb[2] ;
 wire \Tile_X5Y9_S2BEGb[3] ;
 wire \Tile_X5Y9_S2BEGb[4] ;
 wire \Tile_X5Y9_S2BEGb[5] ;
 wire \Tile_X5Y9_S2BEGb[6] ;
 wire \Tile_X5Y9_S2BEGb[7] ;
 wire \Tile_X5Y9_S4BEG[0] ;
 wire \Tile_X5Y9_S4BEG[10] ;
 wire \Tile_X5Y9_S4BEG[11] ;
 wire \Tile_X5Y9_S4BEG[12] ;
 wire \Tile_X5Y9_S4BEG[13] ;
 wire \Tile_X5Y9_S4BEG[14] ;
 wire \Tile_X5Y9_S4BEG[15] ;
 wire \Tile_X5Y9_S4BEG[1] ;
 wire \Tile_X5Y9_S4BEG[2] ;
 wire \Tile_X5Y9_S4BEG[3] ;
 wire \Tile_X5Y9_S4BEG[4] ;
 wire \Tile_X5Y9_S4BEG[5] ;
 wire \Tile_X5Y9_S4BEG[6] ;
 wire \Tile_X5Y9_S4BEG[7] ;
 wire \Tile_X5Y9_S4BEG[8] ;
 wire \Tile_X5Y9_S4BEG[9] ;
 wire \Tile_X5Y9_SS4BEG[0] ;
 wire \Tile_X5Y9_SS4BEG[10] ;
 wire \Tile_X5Y9_SS4BEG[11] ;
 wire \Tile_X5Y9_SS4BEG[12] ;
 wire \Tile_X5Y9_SS4BEG[13] ;
 wire \Tile_X5Y9_SS4BEG[14] ;
 wire \Tile_X5Y9_SS4BEG[15] ;
 wire \Tile_X5Y9_SS4BEG[1] ;
 wire \Tile_X5Y9_SS4BEG[2] ;
 wire \Tile_X5Y9_SS4BEG[3] ;
 wire \Tile_X5Y9_SS4BEG[4] ;
 wire \Tile_X5Y9_SS4BEG[5] ;
 wire \Tile_X5Y9_SS4BEG[6] ;
 wire \Tile_X5Y9_SS4BEG[7] ;
 wire \Tile_X5Y9_SS4BEG[8] ;
 wire \Tile_X5Y9_SS4BEG[9] ;
 wire Tile_X5Y9_UserCLKo;
 wire \Tile_X5Y9_W1BEG[0] ;
 wire \Tile_X5Y9_W1BEG[1] ;
 wire \Tile_X5Y9_W1BEG[2] ;
 wire \Tile_X5Y9_W1BEG[3] ;
 wire \Tile_X5Y9_W2BEG[0] ;
 wire \Tile_X5Y9_W2BEG[1] ;
 wire \Tile_X5Y9_W2BEG[2] ;
 wire \Tile_X5Y9_W2BEG[3] ;
 wire \Tile_X5Y9_W2BEG[4] ;
 wire \Tile_X5Y9_W2BEG[5] ;
 wire \Tile_X5Y9_W2BEG[6] ;
 wire \Tile_X5Y9_W2BEG[7] ;
 wire \Tile_X5Y9_W2BEGb[0] ;
 wire \Tile_X5Y9_W2BEGb[1] ;
 wire \Tile_X5Y9_W2BEGb[2] ;
 wire \Tile_X5Y9_W2BEGb[3] ;
 wire \Tile_X5Y9_W2BEGb[4] ;
 wire \Tile_X5Y9_W2BEGb[5] ;
 wire \Tile_X5Y9_W2BEGb[6] ;
 wire \Tile_X5Y9_W2BEGb[7] ;
 wire \Tile_X5Y9_W6BEG[0] ;
 wire \Tile_X5Y9_W6BEG[10] ;
 wire \Tile_X5Y9_W6BEG[11] ;
 wire \Tile_X5Y9_W6BEG[1] ;
 wire \Tile_X5Y9_W6BEG[2] ;
 wire \Tile_X5Y9_W6BEG[3] ;
 wire \Tile_X5Y9_W6BEG[4] ;
 wire \Tile_X5Y9_W6BEG[5] ;
 wire \Tile_X5Y9_W6BEG[6] ;
 wire \Tile_X5Y9_W6BEG[7] ;
 wire \Tile_X5Y9_W6BEG[8] ;
 wire \Tile_X5Y9_W6BEG[9] ;
 wire \Tile_X5Y9_WW4BEG[0] ;
 wire \Tile_X5Y9_WW4BEG[10] ;
 wire \Tile_X5Y9_WW4BEG[11] ;
 wire \Tile_X5Y9_WW4BEG[12] ;
 wire \Tile_X5Y9_WW4BEG[13] ;
 wire \Tile_X5Y9_WW4BEG[14] ;
 wire \Tile_X5Y9_WW4BEG[15] ;
 wire \Tile_X5Y9_WW4BEG[1] ;
 wire \Tile_X5Y9_WW4BEG[2] ;
 wire \Tile_X5Y9_WW4BEG[3] ;
 wire \Tile_X5Y9_WW4BEG[4] ;
 wire \Tile_X5Y9_WW4BEG[5] ;
 wire \Tile_X5Y9_WW4BEG[6] ;
 wire \Tile_X5Y9_WW4BEG[7] ;
 wire \Tile_X5Y9_WW4BEG[8] ;
 wire \Tile_X5Y9_WW4BEG[9] ;
 wire \Tile_X6Y0_FrameData_O[0] ;
 wire \Tile_X6Y0_FrameData_O[10] ;
 wire \Tile_X6Y0_FrameData_O[11] ;
 wire \Tile_X6Y0_FrameData_O[12] ;
 wire \Tile_X6Y0_FrameData_O[13] ;
 wire \Tile_X6Y0_FrameData_O[14] ;
 wire \Tile_X6Y0_FrameData_O[15] ;
 wire \Tile_X6Y0_FrameData_O[16] ;
 wire \Tile_X6Y0_FrameData_O[17] ;
 wire \Tile_X6Y0_FrameData_O[18] ;
 wire \Tile_X6Y0_FrameData_O[19] ;
 wire \Tile_X6Y0_FrameData_O[1] ;
 wire \Tile_X6Y0_FrameData_O[20] ;
 wire \Tile_X6Y0_FrameData_O[21] ;
 wire \Tile_X6Y0_FrameData_O[22] ;
 wire \Tile_X6Y0_FrameData_O[23] ;
 wire \Tile_X6Y0_FrameData_O[24] ;
 wire \Tile_X6Y0_FrameData_O[25] ;
 wire \Tile_X6Y0_FrameData_O[26] ;
 wire \Tile_X6Y0_FrameData_O[27] ;
 wire \Tile_X6Y0_FrameData_O[28] ;
 wire \Tile_X6Y0_FrameData_O[29] ;
 wire \Tile_X6Y0_FrameData_O[2] ;
 wire \Tile_X6Y0_FrameData_O[30] ;
 wire \Tile_X6Y0_FrameData_O[31] ;
 wire \Tile_X6Y0_FrameData_O[3] ;
 wire \Tile_X6Y0_FrameData_O[4] ;
 wire \Tile_X6Y0_FrameData_O[5] ;
 wire \Tile_X6Y0_FrameData_O[6] ;
 wire \Tile_X6Y0_FrameData_O[7] ;
 wire \Tile_X6Y0_FrameData_O[8] ;
 wire \Tile_X6Y0_FrameData_O[9] ;
 wire \Tile_X6Y0_FrameStrobe_O[0] ;
 wire \Tile_X6Y0_FrameStrobe_O[10] ;
 wire \Tile_X6Y0_FrameStrobe_O[11] ;
 wire \Tile_X6Y0_FrameStrobe_O[12] ;
 wire \Tile_X6Y0_FrameStrobe_O[13] ;
 wire \Tile_X6Y0_FrameStrobe_O[14] ;
 wire \Tile_X6Y0_FrameStrobe_O[15] ;
 wire \Tile_X6Y0_FrameStrobe_O[16] ;
 wire \Tile_X6Y0_FrameStrobe_O[17] ;
 wire \Tile_X6Y0_FrameStrobe_O[18] ;
 wire \Tile_X6Y0_FrameStrobe_O[19] ;
 wire \Tile_X6Y0_FrameStrobe_O[1] ;
 wire \Tile_X6Y0_FrameStrobe_O[2] ;
 wire \Tile_X6Y0_FrameStrobe_O[3] ;
 wire \Tile_X6Y0_FrameStrobe_O[4] ;
 wire \Tile_X6Y0_FrameStrobe_O[5] ;
 wire \Tile_X6Y0_FrameStrobe_O[6] ;
 wire \Tile_X6Y0_FrameStrobe_O[7] ;
 wire \Tile_X6Y0_FrameStrobe_O[8] ;
 wire \Tile_X6Y0_FrameStrobe_O[9] ;
 wire \Tile_X6Y0_S1BEG[0] ;
 wire \Tile_X6Y0_S1BEG[1] ;
 wire \Tile_X6Y0_S1BEG[2] ;
 wire \Tile_X6Y0_S1BEG[3] ;
 wire \Tile_X6Y0_S2BEG[0] ;
 wire \Tile_X6Y0_S2BEG[1] ;
 wire \Tile_X6Y0_S2BEG[2] ;
 wire \Tile_X6Y0_S2BEG[3] ;
 wire \Tile_X6Y0_S2BEG[4] ;
 wire \Tile_X6Y0_S2BEG[5] ;
 wire \Tile_X6Y0_S2BEG[6] ;
 wire \Tile_X6Y0_S2BEG[7] ;
 wire \Tile_X6Y0_S2BEGb[0] ;
 wire \Tile_X6Y0_S2BEGb[1] ;
 wire \Tile_X6Y0_S2BEGb[2] ;
 wire \Tile_X6Y0_S2BEGb[3] ;
 wire \Tile_X6Y0_S2BEGb[4] ;
 wire \Tile_X6Y0_S2BEGb[5] ;
 wire \Tile_X6Y0_S2BEGb[6] ;
 wire \Tile_X6Y0_S2BEGb[7] ;
 wire \Tile_X6Y0_S4BEG[0] ;
 wire \Tile_X6Y0_S4BEG[10] ;
 wire \Tile_X6Y0_S4BEG[11] ;
 wire \Tile_X6Y0_S4BEG[12] ;
 wire \Tile_X6Y0_S4BEG[13] ;
 wire \Tile_X6Y0_S4BEG[14] ;
 wire \Tile_X6Y0_S4BEG[15] ;
 wire \Tile_X6Y0_S4BEG[1] ;
 wire \Tile_X6Y0_S4BEG[2] ;
 wire \Tile_X6Y0_S4BEG[3] ;
 wire \Tile_X6Y0_S4BEG[4] ;
 wire \Tile_X6Y0_S4BEG[5] ;
 wire \Tile_X6Y0_S4BEG[6] ;
 wire \Tile_X6Y0_S4BEG[7] ;
 wire \Tile_X6Y0_S4BEG[8] ;
 wire \Tile_X6Y0_S4BEG[9] ;
 wire \Tile_X6Y0_SS4BEG[0] ;
 wire \Tile_X6Y0_SS4BEG[10] ;
 wire \Tile_X6Y0_SS4BEG[11] ;
 wire \Tile_X6Y0_SS4BEG[12] ;
 wire \Tile_X6Y0_SS4BEG[13] ;
 wire \Tile_X6Y0_SS4BEG[14] ;
 wire \Tile_X6Y0_SS4BEG[15] ;
 wire \Tile_X6Y0_SS4BEG[1] ;
 wire \Tile_X6Y0_SS4BEG[2] ;
 wire \Tile_X6Y0_SS4BEG[3] ;
 wire \Tile_X6Y0_SS4BEG[4] ;
 wire \Tile_X6Y0_SS4BEG[5] ;
 wire \Tile_X6Y0_SS4BEG[6] ;
 wire \Tile_X6Y0_SS4BEG[7] ;
 wire \Tile_X6Y0_SS4BEG[8] ;
 wire \Tile_X6Y0_SS4BEG[9] ;
 wire Tile_X6Y0_UserCLKo;
 wire Tile_X6Y10_Co;
 wire \Tile_X6Y10_E1BEG[0] ;
 wire \Tile_X6Y10_E1BEG[1] ;
 wire \Tile_X6Y10_E1BEG[2] ;
 wire \Tile_X6Y10_E1BEG[3] ;
 wire \Tile_X6Y10_E2BEG[0] ;
 wire \Tile_X6Y10_E2BEG[1] ;
 wire \Tile_X6Y10_E2BEG[2] ;
 wire \Tile_X6Y10_E2BEG[3] ;
 wire \Tile_X6Y10_E2BEG[4] ;
 wire \Tile_X6Y10_E2BEG[5] ;
 wire \Tile_X6Y10_E2BEG[6] ;
 wire \Tile_X6Y10_E2BEG[7] ;
 wire \Tile_X6Y10_E2BEGb[0] ;
 wire \Tile_X6Y10_E2BEGb[1] ;
 wire \Tile_X6Y10_E2BEGb[2] ;
 wire \Tile_X6Y10_E2BEGb[3] ;
 wire \Tile_X6Y10_E2BEGb[4] ;
 wire \Tile_X6Y10_E2BEGb[5] ;
 wire \Tile_X6Y10_E2BEGb[6] ;
 wire \Tile_X6Y10_E2BEGb[7] ;
 wire \Tile_X6Y10_E6BEG[0] ;
 wire \Tile_X6Y10_E6BEG[10] ;
 wire \Tile_X6Y10_E6BEG[11] ;
 wire \Tile_X6Y10_E6BEG[1] ;
 wire \Tile_X6Y10_E6BEG[2] ;
 wire \Tile_X6Y10_E6BEG[3] ;
 wire \Tile_X6Y10_E6BEG[4] ;
 wire \Tile_X6Y10_E6BEG[5] ;
 wire \Tile_X6Y10_E6BEG[6] ;
 wire \Tile_X6Y10_E6BEG[7] ;
 wire \Tile_X6Y10_E6BEG[8] ;
 wire \Tile_X6Y10_E6BEG[9] ;
 wire \Tile_X6Y10_EE4BEG[0] ;
 wire \Tile_X6Y10_EE4BEG[10] ;
 wire \Tile_X6Y10_EE4BEG[11] ;
 wire \Tile_X6Y10_EE4BEG[12] ;
 wire \Tile_X6Y10_EE4BEG[13] ;
 wire \Tile_X6Y10_EE4BEG[14] ;
 wire \Tile_X6Y10_EE4BEG[15] ;
 wire \Tile_X6Y10_EE4BEG[1] ;
 wire \Tile_X6Y10_EE4BEG[2] ;
 wire \Tile_X6Y10_EE4BEG[3] ;
 wire \Tile_X6Y10_EE4BEG[4] ;
 wire \Tile_X6Y10_EE4BEG[5] ;
 wire \Tile_X6Y10_EE4BEG[6] ;
 wire \Tile_X6Y10_EE4BEG[7] ;
 wire \Tile_X6Y10_EE4BEG[8] ;
 wire \Tile_X6Y10_EE4BEG[9] ;
 wire \Tile_X6Y10_FrameData_O[0] ;
 wire \Tile_X6Y10_FrameData_O[10] ;
 wire \Tile_X6Y10_FrameData_O[11] ;
 wire \Tile_X6Y10_FrameData_O[12] ;
 wire \Tile_X6Y10_FrameData_O[13] ;
 wire \Tile_X6Y10_FrameData_O[14] ;
 wire \Tile_X6Y10_FrameData_O[15] ;
 wire \Tile_X6Y10_FrameData_O[16] ;
 wire \Tile_X6Y10_FrameData_O[17] ;
 wire \Tile_X6Y10_FrameData_O[18] ;
 wire \Tile_X6Y10_FrameData_O[19] ;
 wire \Tile_X6Y10_FrameData_O[1] ;
 wire \Tile_X6Y10_FrameData_O[20] ;
 wire \Tile_X6Y10_FrameData_O[21] ;
 wire \Tile_X6Y10_FrameData_O[22] ;
 wire \Tile_X6Y10_FrameData_O[23] ;
 wire \Tile_X6Y10_FrameData_O[24] ;
 wire \Tile_X6Y10_FrameData_O[25] ;
 wire \Tile_X6Y10_FrameData_O[26] ;
 wire \Tile_X6Y10_FrameData_O[27] ;
 wire \Tile_X6Y10_FrameData_O[28] ;
 wire \Tile_X6Y10_FrameData_O[29] ;
 wire \Tile_X6Y10_FrameData_O[2] ;
 wire \Tile_X6Y10_FrameData_O[30] ;
 wire \Tile_X6Y10_FrameData_O[31] ;
 wire \Tile_X6Y10_FrameData_O[3] ;
 wire \Tile_X6Y10_FrameData_O[4] ;
 wire \Tile_X6Y10_FrameData_O[5] ;
 wire \Tile_X6Y10_FrameData_O[6] ;
 wire \Tile_X6Y10_FrameData_O[7] ;
 wire \Tile_X6Y10_FrameData_O[8] ;
 wire \Tile_X6Y10_FrameData_O[9] ;
 wire \Tile_X6Y10_FrameStrobe_O[0] ;
 wire \Tile_X6Y10_FrameStrobe_O[10] ;
 wire \Tile_X6Y10_FrameStrobe_O[11] ;
 wire \Tile_X6Y10_FrameStrobe_O[12] ;
 wire \Tile_X6Y10_FrameStrobe_O[13] ;
 wire \Tile_X6Y10_FrameStrobe_O[14] ;
 wire \Tile_X6Y10_FrameStrobe_O[15] ;
 wire \Tile_X6Y10_FrameStrobe_O[16] ;
 wire \Tile_X6Y10_FrameStrobe_O[17] ;
 wire \Tile_X6Y10_FrameStrobe_O[18] ;
 wire \Tile_X6Y10_FrameStrobe_O[19] ;
 wire \Tile_X6Y10_FrameStrobe_O[1] ;
 wire \Tile_X6Y10_FrameStrobe_O[2] ;
 wire \Tile_X6Y10_FrameStrobe_O[3] ;
 wire \Tile_X6Y10_FrameStrobe_O[4] ;
 wire \Tile_X6Y10_FrameStrobe_O[5] ;
 wire \Tile_X6Y10_FrameStrobe_O[6] ;
 wire \Tile_X6Y10_FrameStrobe_O[7] ;
 wire \Tile_X6Y10_FrameStrobe_O[8] ;
 wire \Tile_X6Y10_FrameStrobe_O[9] ;
 wire \Tile_X6Y10_N1BEG[0] ;
 wire \Tile_X6Y10_N1BEG[1] ;
 wire \Tile_X6Y10_N1BEG[2] ;
 wire \Tile_X6Y10_N1BEG[3] ;
 wire \Tile_X6Y10_N2BEG[0] ;
 wire \Tile_X6Y10_N2BEG[1] ;
 wire \Tile_X6Y10_N2BEG[2] ;
 wire \Tile_X6Y10_N2BEG[3] ;
 wire \Tile_X6Y10_N2BEG[4] ;
 wire \Tile_X6Y10_N2BEG[5] ;
 wire \Tile_X6Y10_N2BEG[6] ;
 wire \Tile_X6Y10_N2BEG[7] ;
 wire \Tile_X6Y10_N2BEGb[0] ;
 wire \Tile_X6Y10_N2BEGb[1] ;
 wire \Tile_X6Y10_N2BEGb[2] ;
 wire \Tile_X6Y10_N2BEGb[3] ;
 wire \Tile_X6Y10_N2BEGb[4] ;
 wire \Tile_X6Y10_N2BEGb[5] ;
 wire \Tile_X6Y10_N2BEGb[6] ;
 wire \Tile_X6Y10_N2BEGb[7] ;
 wire \Tile_X6Y10_N4BEG[0] ;
 wire \Tile_X6Y10_N4BEG[10] ;
 wire \Tile_X6Y10_N4BEG[11] ;
 wire \Tile_X6Y10_N4BEG[12] ;
 wire \Tile_X6Y10_N4BEG[13] ;
 wire \Tile_X6Y10_N4BEG[14] ;
 wire \Tile_X6Y10_N4BEG[15] ;
 wire \Tile_X6Y10_N4BEG[1] ;
 wire \Tile_X6Y10_N4BEG[2] ;
 wire \Tile_X6Y10_N4BEG[3] ;
 wire \Tile_X6Y10_N4BEG[4] ;
 wire \Tile_X6Y10_N4BEG[5] ;
 wire \Tile_X6Y10_N4BEG[6] ;
 wire \Tile_X6Y10_N4BEG[7] ;
 wire \Tile_X6Y10_N4BEG[8] ;
 wire \Tile_X6Y10_N4BEG[9] ;
 wire \Tile_X6Y10_NN4BEG[0] ;
 wire \Tile_X6Y10_NN4BEG[10] ;
 wire \Tile_X6Y10_NN4BEG[11] ;
 wire \Tile_X6Y10_NN4BEG[12] ;
 wire \Tile_X6Y10_NN4BEG[13] ;
 wire \Tile_X6Y10_NN4BEG[14] ;
 wire \Tile_X6Y10_NN4BEG[15] ;
 wire \Tile_X6Y10_NN4BEG[1] ;
 wire \Tile_X6Y10_NN4BEG[2] ;
 wire \Tile_X6Y10_NN4BEG[3] ;
 wire \Tile_X6Y10_NN4BEG[4] ;
 wire \Tile_X6Y10_NN4BEG[5] ;
 wire \Tile_X6Y10_NN4BEG[6] ;
 wire \Tile_X6Y10_NN4BEG[7] ;
 wire \Tile_X6Y10_NN4BEG[8] ;
 wire \Tile_X6Y10_NN4BEG[9] ;
 wire \Tile_X6Y10_S1BEG[0] ;
 wire \Tile_X6Y10_S1BEG[1] ;
 wire \Tile_X6Y10_S1BEG[2] ;
 wire \Tile_X6Y10_S1BEG[3] ;
 wire \Tile_X6Y10_S2BEG[0] ;
 wire \Tile_X6Y10_S2BEG[1] ;
 wire \Tile_X6Y10_S2BEG[2] ;
 wire \Tile_X6Y10_S2BEG[3] ;
 wire \Tile_X6Y10_S2BEG[4] ;
 wire \Tile_X6Y10_S2BEG[5] ;
 wire \Tile_X6Y10_S2BEG[6] ;
 wire \Tile_X6Y10_S2BEG[7] ;
 wire \Tile_X6Y10_S2BEGb[0] ;
 wire \Tile_X6Y10_S2BEGb[1] ;
 wire \Tile_X6Y10_S2BEGb[2] ;
 wire \Tile_X6Y10_S2BEGb[3] ;
 wire \Tile_X6Y10_S2BEGb[4] ;
 wire \Tile_X6Y10_S2BEGb[5] ;
 wire \Tile_X6Y10_S2BEGb[6] ;
 wire \Tile_X6Y10_S2BEGb[7] ;
 wire \Tile_X6Y10_S4BEG[0] ;
 wire \Tile_X6Y10_S4BEG[10] ;
 wire \Tile_X6Y10_S4BEG[11] ;
 wire \Tile_X6Y10_S4BEG[12] ;
 wire \Tile_X6Y10_S4BEG[13] ;
 wire \Tile_X6Y10_S4BEG[14] ;
 wire \Tile_X6Y10_S4BEG[15] ;
 wire \Tile_X6Y10_S4BEG[1] ;
 wire \Tile_X6Y10_S4BEG[2] ;
 wire \Tile_X6Y10_S4BEG[3] ;
 wire \Tile_X6Y10_S4BEG[4] ;
 wire \Tile_X6Y10_S4BEG[5] ;
 wire \Tile_X6Y10_S4BEG[6] ;
 wire \Tile_X6Y10_S4BEG[7] ;
 wire \Tile_X6Y10_S4BEG[8] ;
 wire \Tile_X6Y10_S4BEG[9] ;
 wire \Tile_X6Y10_SS4BEG[0] ;
 wire \Tile_X6Y10_SS4BEG[10] ;
 wire \Tile_X6Y10_SS4BEG[11] ;
 wire \Tile_X6Y10_SS4BEG[12] ;
 wire \Tile_X6Y10_SS4BEG[13] ;
 wire \Tile_X6Y10_SS4BEG[14] ;
 wire \Tile_X6Y10_SS4BEG[15] ;
 wire \Tile_X6Y10_SS4BEG[1] ;
 wire \Tile_X6Y10_SS4BEG[2] ;
 wire \Tile_X6Y10_SS4BEG[3] ;
 wire \Tile_X6Y10_SS4BEG[4] ;
 wire \Tile_X6Y10_SS4BEG[5] ;
 wire \Tile_X6Y10_SS4BEG[6] ;
 wire \Tile_X6Y10_SS4BEG[7] ;
 wire \Tile_X6Y10_SS4BEG[8] ;
 wire \Tile_X6Y10_SS4BEG[9] ;
 wire Tile_X6Y10_UserCLKo;
 wire \Tile_X6Y10_W1BEG[0] ;
 wire \Tile_X6Y10_W1BEG[1] ;
 wire \Tile_X6Y10_W1BEG[2] ;
 wire \Tile_X6Y10_W1BEG[3] ;
 wire \Tile_X6Y10_W2BEG[0] ;
 wire \Tile_X6Y10_W2BEG[1] ;
 wire \Tile_X6Y10_W2BEG[2] ;
 wire \Tile_X6Y10_W2BEG[3] ;
 wire \Tile_X6Y10_W2BEG[4] ;
 wire \Tile_X6Y10_W2BEG[5] ;
 wire \Tile_X6Y10_W2BEG[6] ;
 wire \Tile_X6Y10_W2BEG[7] ;
 wire \Tile_X6Y10_W2BEGb[0] ;
 wire \Tile_X6Y10_W2BEGb[1] ;
 wire \Tile_X6Y10_W2BEGb[2] ;
 wire \Tile_X6Y10_W2BEGb[3] ;
 wire \Tile_X6Y10_W2BEGb[4] ;
 wire \Tile_X6Y10_W2BEGb[5] ;
 wire \Tile_X6Y10_W2BEGb[6] ;
 wire \Tile_X6Y10_W2BEGb[7] ;
 wire \Tile_X6Y10_W6BEG[0] ;
 wire \Tile_X6Y10_W6BEG[10] ;
 wire \Tile_X6Y10_W6BEG[11] ;
 wire \Tile_X6Y10_W6BEG[1] ;
 wire \Tile_X6Y10_W6BEG[2] ;
 wire \Tile_X6Y10_W6BEG[3] ;
 wire \Tile_X6Y10_W6BEG[4] ;
 wire \Tile_X6Y10_W6BEG[5] ;
 wire \Tile_X6Y10_W6BEG[6] ;
 wire \Tile_X6Y10_W6BEG[7] ;
 wire \Tile_X6Y10_W6BEG[8] ;
 wire \Tile_X6Y10_W6BEG[9] ;
 wire \Tile_X6Y10_WW4BEG[0] ;
 wire \Tile_X6Y10_WW4BEG[10] ;
 wire \Tile_X6Y10_WW4BEG[11] ;
 wire \Tile_X6Y10_WW4BEG[12] ;
 wire \Tile_X6Y10_WW4BEG[13] ;
 wire \Tile_X6Y10_WW4BEG[14] ;
 wire \Tile_X6Y10_WW4BEG[15] ;
 wire \Tile_X6Y10_WW4BEG[1] ;
 wire \Tile_X6Y10_WW4BEG[2] ;
 wire \Tile_X6Y10_WW4BEG[3] ;
 wire \Tile_X6Y10_WW4BEG[4] ;
 wire \Tile_X6Y10_WW4BEG[5] ;
 wire \Tile_X6Y10_WW4BEG[6] ;
 wire \Tile_X6Y10_WW4BEG[7] ;
 wire \Tile_X6Y10_WW4BEG[8] ;
 wire \Tile_X6Y10_WW4BEG[9] ;
 wire Tile_X6Y11_Co;
 wire \Tile_X6Y11_E1BEG[0] ;
 wire \Tile_X6Y11_E1BEG[1] ;
 wire \Tile_X6Y11_E1BEG[2] ;
 wire \Tile_X6Y11_E1BEG[3] ;
 wire \Tile_X6Y11_E2BEG[0] ;
 wire \Tile_X6Y11_E2BEG[1] ;
 wire \Tile_X6Y11_E2BEG[2] ;
 wire \Tile_X6Y11_E2BEG[3] ;
 wire \Tile_X6Y11_E2BEG[4] ;
 wire \Tile_X6Y11_E2BEG[5] ;
 wire \Tile_X6Y11_E2BEG[6] ;
 wire \Tile_X6Y11_E2BEG[7] ;
 wire \Tile_X6Y11_E2BEGb[0] ;
 wire \Tile_X6Y11_E2BEGb[1] ;
 wire \Tile_X6Y11_E2BEGb[2] ;
 wire \Tile_X6Y11_E2BEGb[3] ;
 wire \Tile_X6Y11_E2BEGb[4] ;
 wire \Tile_X6Y11_E2BEGb[5] ;
 wire \Tile_X6Y11_E2BEGb[6] ;
 wire \Tile_X6Y11_E2BEGb[7] ;
 wire \Tile_X6Y11_E6BEG[0] ;
 wire \Tile_X6Y11_E6BEG[10] ;
 wire \Tile_X6Y11_E6BEG[11] ;
 wire \Tile_X6Y11_E6BEG[1] ;
 wire \Tile_X6Y11_E6BEG[2] ;
 wire \Tile_X6Y11_E6BEG[3] ;
 wire \Tile_X6Y11_E6BEG[4] ;
 wire \Tile_X6Y11_E6BEG[5] ;
 wire \Tile_X6Y11_E6BEG[6] ;
 wire \Tile_X6Y11_E6BEG[7] ;
 wire \Tile_X6Y11_E6BEG[8] ;
 wire \Tile_X6Y11_E6BEG[9] ;
 wire \Tile_X6Y11_EE4BEG[0] ;
 wire \Tile_X6Y11_EE4BEG[10] ;
 wire \Tile_X6Y11_EE4BEG[11] ;
 wire \Tile_X6Y11_EE4BEG[12] ;
 wire \Tile_X6Y11_EE4BEG[13] ;
 wire \Tile_X6Y11_EE4BEG[14] ;
 wire \Tile_X6Y11_EE4BEG[15] ;
 wire \Tile_X6Y11_EE4BEG[1] ;
 wire \Tile_X6Y11_EE4BEG[2] ;
 wire \Tile_X6Y11_EE4BEG[3] ;
 wire \Tile_X6Y11_EE4BEG[4] ;
 wire \Tile_X6Y11_EE4BEG[5] ;
 wire \Tile_X6Y11_EE4BEG[6] ;
 wire \Tile_X6Y11_EE4BEG[7] ;
 wire \Tile_X6Y11_EE4BEG[8] ;
 wire \Tile_X6Y11_EE4BEG[9] ;
 wire \Tile_X6Y11_FrameData_O[0] ;
 wire \Tile_X6Y11_FrameData_O[10] ;
 wire \Tile_X6Y11_FrameData_O[11] ;
 wire \Tile_X6Y11_FrameData_O[12] ;
 wire \Tile_X6Y11_FrameData_O[13] ;
 wire \Tile_X6Y11_FrameData_O[14] ;
 wire \Tile_X6Y11_FrameData_O[15] ;
 wire \Tile_X6Y11_FrameData_O[16] ;
 wire \Tile_X6Y11_FrameData_O[17] ;
 wire \Tile_X6Y11_FrameData_O[18] ;
 wire \Tile_X6Y11_FrameData_O[19] ;
 wire \Tile_X6Y11_FrameData_O[1] ;
 wire \Tile_X6Y11_FrameData_O[20] ;
 wire \Tile_X6Y11_FrameData_O[21] ;
 wire \Tile_X6Y11_FrameData_O[22] ;
 wire \Tile_X6Y11_FrameData_O[23] ;
 wire \Tile_X6Y11_FrameData_O[24] ;
 wire \Tile_X6Y11_FrameData_O[25] ;
 wire \Tile_X6Y11_FrameData_O[26] ;
 wire \Tile_X6Y11_FrameData_O[27] ;
 wire \Tile_X6Y11_FrameData_O[28] ;
 wire \Tile_X6Y11_FrameData_O[29] ;
 wire \Tile_X6Y11_FrameData_O[2] ;
 wire \Tile_X6Y11_FrameData_O[30] ;
 wire \Tile_X6Y11_FrameData_O[31] ;
 wire \Tile_X6Y11_FrameData_O[3] ;
 wire \Tile_X6Y11_FrameData_O[4] ;
 wire \Tile_X6Y11_FrameData_O[5] ;
 wire \Tile_X6Y11_FrameData_O[6] ;
 wire \Tile_X6Y11_FrameData_O[7] ;
 wire \Tile_X6Y11_FrameData_O[8] ;
 wire \Tile_X6Y11_FrameData_O[9] ;
 wire \Tile_X6Y11_FrameStrobe_O[0] ;
 wire \Tile_X6Y11_FrameStrobe_O[10] ;
 wire \Tile_X6Y11_FrameStrobe_O[11] ;
 wire \Tile_X6Y11_FrameStrobe_O[12] ;
 wire \Tile_X6Y11_FrameStrobe_O[13] ;
 wire \Tile_X6Y11_FrameStrobe_O[14] ;
 wire \Tile_X6Y11_FrameStrobe_O[15] ;
 wire \Tile_X6Y11_FrameStrobe_O[16] ;
 wire \Tile_X6Y11_FrameStrobe_O[17] ;
 wire \Tile_X6Y11_FrameStrobe_O[18] ;
 wire \Tile_X6Y11_FrameStrobe_O[19] ;
 wire \Tile_X6Y11_FrameStrobe_O[1] ;
 wire \Tile_X6Y11_FrameStrobe_O[2] ;
 wire \Tile_X6Y11_FrameStrobe_O[3] ;
 wire \Tile_X6Y11_FrameStrobe_O[4] ;
 wire \Tile_X6Y11_FrameStrobe_O[5] ;
 wire \Tile_X6Y11_FrameStrobe_O[6] ;
 wire \Tile_X6Y11_FrameStrobe_O[7] ;
 wire \Tile_X6Y11_FrameStrobe_O[8] ;
 wire \Tile_X6Y11_FrameStrobe_O[9] ;
 wire \Tile_X6Y11_N1BEG[0] ;
 wire \Tile_X6Y11_N1BEG[1] ;
 wire \Tile_X6Y11_N1BEG[2] ;
 wire \Tile_X6Y11_N1BEG[3] ;
 wire \Tile_X6Y11_N2BEG[0] ;
 wire \Tile_X6Y11_N2BEG[1] ;
 wire \Tile_X6Y11_N2BEG[2] ;
 wire \Tile_X6Y11_N2BEG[3] ;
 wire \Tile_X6Y11_N2BEG[4] ;
 wire \Tile_X6Y11_N2BEG[5] ;
 wire \Tile_X6Y11_N2BEG[6] ;
 wire \Tile_X6Y11_N2BEG[7] ;
 wire \Tile_X6Y11_N2BEGb[0] ;
 wire \Tile_X6Y11_N2BEGb[1] ;
 wire \Tile_X6Y11_N2BEGb[2] ;
 wire \Tile_X6Y11_N2BEGb[3] ;
 wire \Tile_X6Y11_N2BEGb[4] ;
 wire \Tile_X6Y11_N2BEGb[5] ;
 wire \Tile_X6Y11_N2BEGb[6] ;
 wire \Tile_X6Y11_N2BEGb[7] ;
 wire \Tile_X6Y11_N4BEG[0] ;
 wire \Tile_X6Y11_N4BEG[10] ;
 wire \Tile_X6Y11_N4BEG[11] ;
 wire \Tile_X6Y11_N4BEG[12] ;
 wire \Tile_X6Y11_N4BEG[13] ;
 wire \Tile_X6Y11_N4BEG[14] ;
 wire \Tile_X6Y11_N4BEG[15] ;
 wire \Tile_X6Y11_N4BEG[1] ;
 wire \Tile_X6Y11_N4BEG[2] ;
 wire \Tile_X6Y11_N4BEG[3] ;
 wire \Tile_X6Y11_N4BEG[4] ;
 wire \Tile_X6Y11_N4BEG[5] ;
 wire \Tile_X6Y11_N4BEG[6] ;
 wire \Tile_X6Y11_N4BEG[7] ;
 wire \Tile_X6Y11_N4BEG[8] ;
 wire \Tile_X6Y11_N4BEG[9] ;
 wire \Tile_X6Y11_NN4BEG[0] ;
 wire \Tile_X6Y11_NN4BEG[10] ;
 wire \Tile_X6Y11_NN4BEG[11] ;
 wire \Tile_X6Y11_NN4BEG[12] ;
 wire \Tile_X6Y11_NN4BEG[13] ;
 wire \Tile_X6Y11_NN4BEG[14] ;
 wire \Tile_X6Y11_NN4BEG[15] ;
 wire \Tile_X6Y11_NN4BEG[1] ;
 wire \Tile_X6Y11_NN4BEG[2] ;
 wire \Tile_X6Y11_NN4BEG[3] ;
 wire \Tile_X6Y11_NN4BEG[4] ;
 wire \Tile_X6Y11_NN4BEG[5] ;
 wire \Tile_X6Y11_NN4BEG[6] ;
 wire \Tile_X6Y11_NN4BEG[7] ;
 wire \Tile_X6Y11_NN4BEG[8] ;
 wire \Tile_X6Y11_NN4BEG[9] ;
 wire \Tile_X6Y11_S1BEG[0] ;
 wire \Tile_X6Y11_S1BEG[1] ;
 wire \Tile_X6Y11_S1BEG[2] ;
 wire \Tile_X6Y11_S1BEG[3] ;
 wire \Tile_X6Y11_S2BEG[0] ;
 wire \Tile_X6Y11_S2BEG[1] ;
 wire \Tile_X6Y11_S2BEG[2] ;
 wire \Tile_X6Y11_S2BEG[3] ;
 wire \Tile_X6Y11_S2BEG[4] ;
 wire \Tile_X6Y11_S2BEG[5] ;
 wire \Tile_X6Y11_S2BEG[6] ;
 wire \Tile_X6Y11_S2BEG[7] ;
 wire \Tile_X6Y11_S2BEGb[0] ;
 wire \Tile_X6Y11_S2BEGb[1] ;
 wire \Tile_X6Y11_S2BEGb[2] ;
 wire \Tile_X6Y11_S2BEGb[3] ;
 wire \Tile_X6Y11_S2BEGb[4] ;
 wire \Tile_X6Y11_S2BEGb[5] ;
 wire \Tile_X6Y11_S2BEGb[6] ;
 wire \Tile_X6Y11_S2BEGb[7] ;
 wire \Tile_X6Y11_S4BEG[0] ;
 wire \Tile_X6Y11_S4BEG[10] ;
 wire \Tile_X6Y11_S4BEG[11] ;
 wire \Tile_X6Y11_S4BEG[12] ;
 wire \Tile_X6Y11_S4BEG[13] ;
 wire \Tile_X6Y11_S4BEG[14] ;
 wire \Tile_X6Y11_S4BEG[15] ;
 wire \Tile_X6Y11_S4BEG[1] ;
 wire \Tile_X6Y11_S4BEG[2] ;
 wire \Tile_X6Y11_S4BEG[3] ;
 wire \Tile_X6Y11_S4BEG[4] ;
 wire \Tile_X6Y11_S4BEG[5] ;
 wire \Tile_X6Y11_S4BEG[6] ;
 wire \Tile_X6Y11_S4BEG[7] ;
 wire \Tile_X6Y11_S4BEG[8] ;
 wire \Tile_X6Y11_S4BEG[9] ;
 wire \Tile_X6Y11_SS4BEG[0] ;
 wire \Tile_X6Y11_SS4BEG[10] ;
 wire \Tile_X6Y11_SS4BEG[11] ;
 wire \Tile_X6Y11_SS4BEG[12] ;
 wire \Tile_X6Y11_SS4BEG[13] ;
 wire \Tile_X6Y11_SS4BEG[14] ;
 wire \Tile_X6Y11_SS4BEG[15] ;
 wire \Tile_X6Y11_SS4BEG[1] ;
 wire \Tile_X6Y11_SS4BEG[2] ;
 wire \Tile_X6Y11_SS4BEG[3] ;
 wire \Tile_X6Y11_SS4BEG[4] ;
 wire \Tile_X6Y11_SS4BEG[5] ;
 wire \Tile_X6Y11_SS4BEG[6] ;
 wire \Tile_X6Y11_SS4BEG[7] ;
 wire \Tile_X6Y11_SS4BEG[8] ;
 wire \Tile_X6Y11_SS4BEG[9] ;
 wire Tile_X6Y11_UserCLKo;
 wire \Tile_X6Y11_W1BEG[0] ;
 wire \Tile_X6Y11_W1BEG[1] ;
 wire \Tile_X6Y11_W1BEG[2] ;
 wire \Tile_X6Y11_W1BEG[3] ;
 wire \Tile_X6Y11_W2BEG[0] ;
 wire \Tile_X6Y11_W2BEG[1] ;
 wire \Tile_X6Y11_W2BEG[2] ;
 wire \Tile_X6Y11_W2BEG[3] ;
 wire \Tile_X6Y11_W2BEG[4] ;
 wire \Tile_X6Y11_W2BEG[5] ;
 wire \Tile_X6Y11_W2BEG[6] ;
 wire \Tile_X6Y11_W2BEG[7] ;
 wire \Tile_X6Y11_W2BEGb[0] ;
 wire \Tile_X6Y11_W2BEGb[1] ;
 wire \Tile_X6Y11_W2BEGb[2] ;
 wire \Tile_X6Y11_W2BEGb[3] ;
 wire \Tile_X6Y11_W2BEGb[4] ;
 wire \Tile_X6Y11_W2BEGb[5] ;
 wire \Tile_X6Y11_W2BEGb[6] ;
 wire \Tile_X6Y11_W2BEGb[7] ;
 wire \Tile_X6Y11_W6BEG[0] ;
 wire \Tile_X6Y11_W6BEG[10] ;
 wire \Tile_X6Y11_W6BEG[11] ;
 wire \Tile_X6Y11_W6BEG[1] ;
 wire \Tile_X6Y11_W6BEG[2] ;
 wire \Tile_X6Y11_W6BEG[3] ;
 wire \Tile_X6Y11_W6BEG[4] ;
 wire \Tile_X6Y11_W6BEG[5] ;
 wire \Tile_X6Y11_W6BEG[6] ;
 wire \Tile_X6Y11_W6BEG[7] ;
 wire \Tile_X6Y11_W6BEG[8] ;
 wire \Tile_X6Y11_W6BEG[9] ;
 wire \Tile_X6Y11_WW4BEG[0] ;
 wire \Tile_X6Y11_WW4BEG[10] ;
 wire \Tile_X6Y11_WW4BEG[11] ;
 wire \Tile_X6Y11_WW4BEG[12] ;
 wire \Tile_X6Y11_WW4BEG[13] ;
 wire \Tile_X6Y11_WW4BEG[14] ;
 wire \Tile_X6Y11_WW4BEG[15] ;
 wire \Tile_X6Y11_WW4BEG[1] ;
 wire \Tile_X6Y11_WW4BEG[2] ;
 wire \Tile_X6Y11_WW4BEG[3] ;
 wire \Tile_X6Y11_WW4BEG[4] ;
 wire \Tile_X6Y11_WW4BEG[5] ;
 wire \Tile_X6Y11_WW4BEG[6] ;
 wire \Tile_X6Y11_WW4BEG[7] ;
 wire \Tile_X6Y11_WW4BEG[8] ;
 wire \Tile_X6Y11_WW4BEG[9] ;
 wire Tile_X6Y12_Co;
 wire \Tile_X6Y12_E1BEG[0] ;
 wire \Tile_X6Y12_E1BEG[1] ;
 wire \Tile_X6Y12_E1BEG[2] ;
 wire \Tile_X6Y12_E1BEG[3] ;
 wire \Tile_X6Y12_E2BEG[0] ;
 wire \Tile_X6Y12_E2BEG[1] ;
 wire \Tile_X6Y12_E2BEG[2] ;
 wire \Tile_X6Y12_E2BEG[3] ;
 wire \Tile_X6Y12_E2BEG[4] ;
 wire \Tile_X6Y12_E2BEG[5] ;
 wire \Tile_X6Y12_E2BEG[6] ;
 wire \Tile_X6Y12_E2BEG[7] ;
 wire \Tile_X6Y12_E2BEGb[0] ;
 wire \Tile_X6Y12_E2BEGb[1] ;
 wire \Tile_X6Y12_E2BEGb[2] ;
 wire \Tile_X6Y12_E2BEGb[3] ;
 wire \Tile_X6Y12_E2BEGb[4] ;
 wire \Tile_X6Y12_E2BEGb[5] ;
 wire \Tile_X6Y12_E2BEGb[6] ;
 wire \Tile_X6Y12_E2BEGb[7] ;
 wire \Tile_X6Y12_E6BEG[0] ;
 wire \Tile_X6Y12_E6BEG[10] ;
 wire \Tile_X6Y12_E6BEG[11] ;
 wire \Tile_X6Y12_E6BEG[1] ;
 wire \Tile_X6Y12_E6BEG[2] ;
 wire \Tile_X6Y12_E6BEG[3] ;
 wire \Tile_X6Y12_E6BEG[4] ;
 wire \Tile_X6Y12_E6BEG[5] ;
 wire \Tile_X6Y12_E6BEG[6] ;
 wire \Tile_X6Y12_E6BEG[7] ;
 wire \Tile_X6Y12_E6BEG[8] ;
 wire \Tile_X6Y12_E6BEG[9] ;
 wire \Tile_X6Y12_EE4BEG[0] ;
 wire \Tile_X6Y12_EE4BEG[10] ;
 wire \Tile_X6Y12_EE4BEG[11] ;
 wire \Tile_X6Y12_EE4BEG[12] ;
 wire \Tile_X6Y12_EE4BEG[13] ;
 wire \Tile_X6Y12_EE4BEG[14] ;
 wire \Tile_X6Y12_EE4BEG[15] ;
 wire \Tile_X6Y12_EE4BEG[1] ;
 wire \Tile_X6Y12_EE4BEG[2] ;
 wire \Tile_X6Y12_EE4BEG[3] ;
 wire \Tile_X6Y12_EE4BEG[4] ;
 wire \Tile_X6Y12_EE4BEG[5] ;
 wire \Tile_X6Y12_EE4BEG[6] ;
 wire \Tile_X6Y12_EE4BEG[7] ;
 wire \Tile_X6Y12_EE4BEG[8] ;
 wire \Tile_X6Y12_EE4BEG[9] ;
 wire \Tile_X6Y12_FrameData_O[0] ;
 wire \Tile_X6Y12_FrameData_O[10] ;
 wire \Tile_X6Y12_FrameData_O[11] ;
 wire \Tile_X6Y12_FrameData_O[12] ;
 wire \Tile_X6Y12_FrameData_O[13] ;
 wire \Tile_X6Y12_FrameData_O[14] ;
 wire \Tile_X6Y12_FrameData_O[15] ;
 wire \Tile_X6Y12_FrameData_O[16] ;
 wire \Tile_X6Y12_FrameData_O[17] ;
 wire \Tile_X6Y12_FrameData_O[18] ;
 wire \Tile_X6Y12_FrameData_O[19] ;
 wire \Tile_X6Y12_FrameData_O[1] ;
 wire \Tile_X6Y12_FrameData_O[20] ;
 wire \Tile_X6Y12_FrameData_O[21] ;
 wire \Tile_X6Y12_FrameData_O[22] ;
 wire \Tile_X6Y12_FrameData_O[23] ;
 wire \Tile_X6Y12_FrameData_O[24] ;
 wire \Tile_X6Y12_FrameData_O[25] ;
 wire \Tile_X6Y12_FrameData_O[26] ;
 wire \Tile_X6Y12_FrameData_O[27] ;
 wire \Tile_X6Y12_FrameData_O[28] ;
 wire \Tile_X6Y12_FrameData_O[29] ;
 wire \Tile_X6Y12_FrameData_O[2] ;
 wire \Tile_X6Y12_FrameData_O[30] ;
 wire \Tile_X6Y12_FrameData_O[31] ;
 wire \Tile_X6Y12_FrameData_O[3] ;
 wire \Tile_X6Y12_FrameData_O[4] ;
 wire \Tile_X6Y12_FrameData_O[5] ;
 wire \Tile_X6Y12_FrameData_O[6] ;
 wire \Tile_X6Y12_FrameData_O[7] ;
 wire \Tile_X6Y12_FrameData_O[8] ;
 wire \Tile_X6Y12_FrameData_O[9] ;
 wire \Tile_X6Y12_FrameStrobe_O[0] ;
 wire \Tile_X6Y12_FrameStrobe_O[10] ;
 wire \Tile_X6Y12_FrameStrobe_O[11] ;
 wire \Tile_X6Y12_FrameStrobe_O[12] ;
 wire \Tile_X6Y12_FrameStrobe_O[13] ;
 wire \Tile_X6Y12_FrameStrobe_O[14] ;
 wire \Tile_X6Y12_FrameStrobe_O[15] ;
 wire \Tile_X6Y12_FrameStrobe_O[16] ;
 wire \Tile_X6Y12_FrameStrobe_O[17] ;
 wire \Tile_X6Y12_FrameStrobe_O[18] ;
 wire \Tile_X6Y12_FrameStrobe_O[19] ;
 wire \Tile_X6Y12_FrameStrobe_O[1] ;
 wire \Tile_X6Y12_FrameStrobe_O[2] ;
 wire \Tile_X6Y12_FrameStrobe_O[3] ;
 wire \Tile_X6Y12_FrameStrobe_O[4] ;
 wire \Tile_X6Y12_FrameStrobe_O[5] ;
 wire \Tile_X6Y12_FrameStrobe_O[6] ;
 wire \Tile_X6Y12_FrameStrobe_O[7] ;
 wire \Tile_X6Y12_FrameStrobe_O[8] ;
 wire \Tile_X6Y12_FrameStrobe_O[9] ;
 wire \Tile_X6Y12_N1BEG[0] ;
 wire \Tile_X6Y12_N1BEG[1] ;
 wire \Tile_X6Y12_N1BEG[2] ;
 wire \Tile_X6Y12_N1BEG[3] ;
 wire \Tile_X6Y12_N2BEG[0] ;
 wire \Tile_X6Y12_N2BEG[1] ;
 wire \Tile_X6Y12_N2BEG[2] ;
 wire \Tile_X6Y12_N2BEG[3] ;
 wire \Tile_X6Y12_N2BEG[4] ;
 wire \Tile_X6Y12_N2BEG[5] ;
 wire \Tile_X6Y12_N2BEG[6] ;
 wire \Tile_X6Y12_N2BEG[7] ;
 wire \Tile_X6Y12_N2BEGb[0] ;
 wire \Tile_X6Y12_N2BEGb[1] ;
 wire \Tile_X6Y12_N2BEGb[2] ;
 wire \Tile_X6Y12_N2BEGb[3] ;
 wire \Tile_X6Y12_N2BEGb[4] ;
 wire \Tile_X6Y12_N2BEGb[5] ;
 wire \Tile_X6Y12_N2BEGb[6] ;
 wire \Tile_X6Y12_N2BEGb[7] ;
 wire \Tile_X6Y12_N4BEG[0] ;
 wire \Tile_X6Y12_N4BEG[10] ;
 wire \Tile_X6Y12_N4BEG[11] ;
 wire \Tile_X6Y12_N4BEG[12] ;
 wire \Tile_X6Y12_N4BEG[13] ;
 wire \Tile_X6Y12_N4BEG[14] ;
 wire \Tile_X6Y12_N4BEG[15] ;
 wire \Tile_X6Y12_N4BEG[1] ;
 wire \Tile_X6Y12_N4BEG[2] ;
 wire \Tile_X6Y12_N4BEG[3] ;
 wire \Tile_X6Y12_N4BEG[4] ;
 wire \Tile_X6Y12_N4BEG[5] ;
 wire \Tile_X6Y12_N4BEG[6] ;
 wire \Tile_X6Y12_N4BEG[7] ;
 wire \Tile_X6Y12_N4BEG[8] ;
 wire \Tile_X6Y12_N4BEG[9] ;
 wire \Tile_X6Y12_NN4BEG[0] ;
 wire \Tile_X6Y12_NN4BEG[10] ;
 wire \Tile_X6Y12_NN4BEG[11] ;
 wire \Tile_X6Y12_NN4BEG[12] ;
 wire \Tile_X6Y12_NN4BEG[13] ;
 wire \Tile_X6Y12_NN4BEG[14] ;
 wire \Tile_X6Y12_NN4BEG[15] ;
 wire \Tile_X6Y12_NN4BEG[1] ;
 wire \Tile_X6Y12_NN4BEG[2] ;
 wire \Tile_X6Y12_NN4BEG[3] ;
 wire \Tile_X6Y12_NN4BEG[4] ;
 wire \Tile_X6Y12_NN4BEG[5] ;
 wire \Tile_X6Y12_NN4BEG[6] ;
 wire \Tile_X6Y12_NN4BEG[7] ;
 wire \Tile_X6Y12_NN4BEG[8] ;
 wire \Tile_X6Y12_NN4BEG[9] ;
 wire \Tile_X6Y12_S1BEG[0] ;
 wire \Tile_X6Y12_S1BEG[1] ;
 wire \Tile_X6Y12_S1BEG[2] ;
 wire \Tile_X6Y12_S1BEG[3] ;
 wire \Tile_X6Y12_S2BEG[0] ;
 wire \Tile_X6Y12_S2BEG[1] ;
 wire \Tile_X6Y12_S2BEG[2] ;
 wire \Tile_X6Y12_S2BEG[3] ;
 wire \Tile_X6Y12_S2BEG[4] ;
 wire \Tile_X6Y12_S2BEG[5] ;
 wire \Tile_X6Y12_S2BEG[6] ;
 wire \Tile_X6Y12_S2BEG[7] ;
 wire \Tile_X6Y12_S2BEGb[0] ;
 wire \Tile_X6Y12_S2BEGb[1] ;
 wire \Tile_X6Y12_S2BEGb[2] ;
 wire \Tile_X6Y12_S2BEGb[3] ;
 wire \Tile_X6Y12_S2BEGb[4] ;
 wire \Tile_X6Y12_S2BEGb[5] ;
 wire \Tile_X6Y12_S2BEGb[6] ;
 wire \Tile_X6Y12_S2BEGb[7] ;
 wire \Tile_X6Y12_S4BEG[0] ;
 wire \Tile_X6Y12_S4BEG[10] ;
 wire \Tile_X6Y12_S4BEG[11] ;
 wire \Tile_X6Y12_S4BEG[12] ;
 wire \Tile_X6Y12_S4BEG[13] ;
 wire \Tile_X6Y12_S4BEG[14] ;
 wire \Tile_X6Y12_S4BEG[15] ;
 wire \Tile_X6Y12_S4BEG[1] ;
 wire \Tile_X6Y12_S4BEG[2] ;
 wire \Tile_X6Y12_S4BEG[3] ;
 wire \Tile_X6Y12_S4BEG[4] ;
 wire \Tile_X6Y12_S4BEG[5] ;
 wire \Tile_X6Y12_S4BEG[6] ;
 wire \Tile_X6Y12_S4BEG[7] ;
 wire \Tile_X6Y12_S4BEG[8] ;
 wire \Tile_X6Y12_S4BEG[9] ;
 wire \Tile_X6Y12_SS4BEG[0] ;
 wire \Tile_X6Y12_SS4BEG[10] ;
 wire \Tile_X6Y12_SS4BEG[11] ;
 wire \Tile_X6Y12_SS4BEG[12] ;
 wire \Tile_X6Y12_SS4BEG[13] ;
 wire \Tile_X6Y12_SS4BEG[14] ;
 wire \Tile_X6Y12_SS4BEG[15] ;
 wire \Tile_X6Y12_SS4BEG[1] ;
 wire \Tile_X6Y12_SS4BEG[2] ;
 wire \Tile_X6Y12_SS4BEG[3] ;
 wire \Tile_X6Y12_SS4BEG[4] ;
 wire \Tile_X6Y12_SS4BEG[5] ;
 wire \Tile_X6Y12_SS4BEG[6] ;
 wire \Tile_X6Y12_SS4BEG[7] ;
 wire \Tile_X6Y12_SS4BEG[8] ;
 wire \Tile_X6Y12_SS4BEG[9] ;
 wire Tile_X6Y12_UserCLKo;
 wire \Tile_X6Y12_W1BEG[0] ;
 wire \Tile_X6Y12_W1BEG[1] ;
 wire \Tile_X6Y12_W1BEG[2] ;
 wire \Tile_X6Y12_W1BEG[3] ;
 wire \Tile_X6Y12_W2BEG[0] ;
 wire \Tile_X6Y12_W2BEG[1] ;
 wire \Tile_X6Y12_W2BEG[2] ;
 wire \Tile_X6Y12_W2BEG[3] ;
 wire \Tile_X6Y12_W2BEG[4] ;
 wire \Tile_X6Y12_W2BEG[5] ;
 wire \Tile_X6Y12_W2BEG[6] ;
 wire \Tile_X6Y12_W2BEG[7] ;
 wire \Tile_X6Y12_W2BEGb[0] ;
 wire \Tile_X6Y12_W2BEGb[1] ;
 wire \Tile_X6Y12_W2BEGb[2] ;
 wire \Tile_X6Y12_W2BEGb[3] ;
 wire \Tile_X6Y12_W2BEGb[4] ;
 wire \Tile_X6Y12_W2BEGb[5] ;
 wire \Tile_X6Y12_W2BEGb[6] ;
 wire \Tile_X6Y12_W2BEGb[7] ;
 wire \Tile_X6Y12_W6BEG[0] ;
 wire \Tile_X6Y12_W6BEG[10] ;
 wire \Tile_X6Y12_W6BEG[11] ;
 wire \Tile_X6Y12_W6BEG[1] ;
 wire \Tile_X6Y12_W6BEG[2] ;
 wire \Tile_X6Y12_W6BEG[3] ;
 wire \Tile_X6Y12_W6BEG[4] ;
 wire \Tile_X6Y12_W6BEG[5] ;
 wire \Tile_X6Y12_W6BEG[6] ;
 wire \Tile_X6Y12_W6BEG[7] ;
 wire \Tile_X6Y12_W6BEG[8] ;
 wire \Tile_X6Y12_W6BEG[9] ;
 wire \Tile_X6Y12_WW4BEG[0] ;
 wire \Tile_X6Y12_WW4BEG[10] ;
 wire \Tile_X6Y12_WW4BEG[11] ;
 wire \Tile_X6Y12_WW4BEG[12] ;
 wire \Tile_X6Y12_WW4BEG[13] ;
 wire \Tile_X6Y12_WW4BEG[14] ;
 wire \Tile_X6Y12_WW4BEG[15] ;
 wire \Tile_X6Y12_WW4BEG[1] ;
 wire \Tile_X6Y12_WW4BEG[2] ;
 wire \Tile_X6Y12_WW4BEG[3] ;
 wire \Tile_X6Y12_WW4BEG[4] ;
 wire \Tile_X6Y12_WW4BEG[5] ;
 wire \Tile_X6Y12_WW4BEG[6] ;
 wire \Tile_X6Y12_WW4BEG[7] ;
 wire \Tile_X6Y12_WW4BEG[8] ;
 wire \Tile_X6Y12_WW4BEG[9] ;
 wire Tile_X6Y13_Co;
 wire \Tile_X6Y13_E1BEG[0] ;
 wire \Tile_X6Y13_E1BEG[1] ;
 wire \Tile_X6Y13_E1BEG[2] ;
 wire \Tile_X6Y13_E1BEG[3] ;
 wire \Tile_X6Y13_E2BEG[0] ;
 wire \Tile_X6Y13_E2BEG[1] ;
 wire \Tile_X6Y13_E2BEG[2] ;
 wire \Tile_X6Y13_E2BEG[3] ;
 wire \Tile_X6Y13_E2BEG[4] ;
 wire \Tile_X6Y13_E2BEG[5] ;
 wire \Tile_X6Y13_E2BEG[6] ;
 wire \Tile_X6Y13_E2BEG[7] ;
 wire \Tile_X6Y13_E2BEGb[0] ;
 wire \Tile_X6Y13_E2BEGb[1] ;
 wire \Tile_X6Y13_E2BEGb[2] ;
 wire \Tile_X6Y13_E2BEGb[3] ;
 wire \Tile_X6Y13_E2BEGb[4] ;
 wire \Tile_X6Y13_E2BEGb[5] ;
 wire \Tile_X6Y13_E2BEGb[6] ;
 wire \Tile_X6Y13_E2BEGb[7] ;
 wire \Tile_X6Y13_E6BEG[0] ;
 wire \Tile_X6Y13_E6BEG[10] ;
 wire \Tile_X6Y13_E6BEG[11] ;
 wire \Tile_X6Y13_E6BEG[1] ;
 wire \Tile_X6Y13_E6BEG[2] ;
 wire \Tile_X6Y13_E6BEG[3] ;
 wire \Tile_X6Y13_E6BEG[4] ;
 wire \Tile_X6Y13_E6BEG[5] ;
 wire \Tile_X6Y13_E6BEG[6] ;
 wire \Tile_X6Y13_E6BEG[7] ;
 wire \Tile_X6Y13_E6BEG[8] ;
 wire \Tile_X6Y13_E6BEG[9] ;
 wire \Tile_X6Y13_EE4BEG[0] ;
 wire \Tile_X6Y13_EE4BEG[10] ;
 wire \Tile_X6Y13_EE4BEG[11] ;
 wire \Tile_X6Y13_EE4BEG[12] ;
 wire \Tile_X6Y13_EE4BEG[13] ;
 wire \Tile_X6Y13_EE4BEG[14] ;
 wire \Tile_X6Y13_EE4BEG[15] ;
 wire \Tile_X6Y13_EE4BEG[1] ;
 wire \Tile_X6Y13_EE4BEG[2] ;
 wire \Tile_X6Y13_EE4BEG[3] ;
 wire \Tile_X6Y13_EE4BEG[4] ;
 wire \Tile_X6Y13_EE4BEG[5] ;
 wire \Tile_X6Y13_EE4BEG[6] ;
 wire \Tile_X6Y13_EE4BEG[7] ;
 wire \Tile_X6Y13_EE4BEG[8] ;
 wire \Tile_X6Y13_EE4BEG[9] ;
 wire \Tile_X6Y13_FrameData_O[0] ;
 wire \Tile_X6Y13_FrameData_O[10] ;
 wire \Tile_X6Y13_FrameData_O[11] ;
 wire \Tile_X6Y13_FrameData_O[12] ;
 wire \Tile_X6Y13_FrameData_O[13] ;
 wire \Tile_X6Y13_FrameData_O[14] ;
 wire \Tile_X6Y13_FrameData_O[15] ;
 wire \Tile_X6Y13_FrameData_O[16] ;
 wire \Tile_X6Y13_FrameData_O[17] ;
 wire \Tile_X6Y13_FrameData_O[18] ;
 wire \Tile_X6Y13_FrameData_O[19] ;
 wire \Tile_X6Y13_FrameData_O[1] ;
 wire \Tile_X6Y13_FrameData_O[20] ;
 wire \Tile_X6Y13_FrameData_O[21] ;
 wire \Tile_X6Y13_FrameData_O[22] ;
 wire \Tile_X6Y13_FrameData_O[23] ;
 wire \Tile_X6Y13_FrameData_O[24] ;
 wire \Tile_X6Y13_FrameData_O[25] ;
 wire \Tile_X6Y13_FrameData_O[26] ;
 wire \Tile_X6Y13_FrameData_O[27] ;
 wire \Tile_X6Y13_FrameData_O[28] ;
 wire \Tile_X6Y13_FrameData_O[29] ;
 wire \Tile_X6Y13_FrameData_O[2] ;
 wire \Tile_X6Y13_FrameData_O[30] ;
 wire \Tile_X6Y13_FrameData_O[31] ;
 wire \Tile_X6Y13_FrameData_O[3] ;
 wire \Tile_X6Y13_FrameData_O[4] ;
 wire \Tile_X6Y13_FrameData_O[5] ;
 wire \Tile_X6Y13_FrameData_O[6] ;
 wire \Tile_X6Y13_FrameData_O[7] ;
 wire \Tile_X6Y13_FrameData_O[8] ;
 wire \Tile_X6Y13_FrameData_O[9] ;
 wire \Tile_X6Y13_FrameStrobe_O[0] ;
 wire \Tile_X6Y13_FrameStrobe_O[10] ;
 wire \Tile_X6Y13_FrameStrobe_O[11] ;
 wire \Tile_X6Y13_FrameStrobe_O[12] ;
 wire \Tile_X6Y13_FrameStrobe_O[13] ;
 wire \Tile_X6Y13_FrameStrobe_O[14] ;
 wire \Tile_X6Y13_FrameStrobe_O[15] ;
 wire \Tile_X6Y13_FrameStrobe_O[16] ;
 wire \Tile_X6Y13_FrameStrobe_O[17] ;
 wire \Tile_X6Y13_FrameStrobe_O[18] ;
 wire \Tile_X6Y13_FrameStrobe_O[19] ;
 wire \Tile_X6Y13_FrameStrobe_O[1] ;
 wire \Tile_X6Y13_FrameStrobe_O[2] ;
 wire \Tile_X6Y13_FrameStrobe_O[3] ;
 wire \Tile_X6Y13_FrameStrobe_O[4] ;
 wire \Tile_X6Y13_FrameStrobe_O[5] ;
 wire \Tile_X6Y13_FrameStrobe_O[6] ;
 wire \Tile_X6Y13_FrameStrobe_O[7] ;
 wire \Tile_X6Y13_FrameStrobe_O[8] ;
 wire \Tile_X6Y13_FrameStrobe_O[9] ;
 wire \Tile_X6Y13_N1BEG[0] ;
 wire \Tile_X6Y13_N1BEG[1] ;
 wire \Tile_X6Y13_N1BEG[2] ;
 wire \Tile_X6Y13_N1BEG[3] ;
 wire \Tile_X6Y13_N2BEG[0] ;
 wire \Tile_X6Y13_N2BEG[1] ;
 wire \Tile_X6Y13_N2BEG[2] ;
 wire \Tile_X6Y13_N2BEG[3] ;
 wire \Tile_X6Y13_N2BEG[4] ;
 wire \Tile_X6Y13_N2BEG[5] ;
 wire \Tile_X6Y13_N2BEG[6] ;
 wire \Tile_X6Y13_N2BEG[7] ;
 wire \Tile_X6Y13_N2BEGb[0] ;
 wire \Tile_X6Y13_N2BEGb[1] ;
 wire \Tile_X6Y13_N2BEGb[2] ;
 wire \Tile_X6Y13_N2BEGb[3] ;
 wire \Tile_X6Y13_N2BEGb[4] ;
 wire \Tile_X6Y13_N2BEGb[5] ;
 wire \Tile_X6Y13_N2BEGb[6] ;
 wire \Tile_X6Y13_N2BEGb[7] ;
 wire \Tile_X6Y13_N4BEG[0] ;
 wire \Tile_X6Y13_N4BEG[10] ;
 wire \Tile_X6Y13_N4BEG[11] ;
 wire \Tile_X6Y13_N4BEG[12] ;
 wire \Tile_X6Y13_N4BEG[13] ;
 wire \Tile_X6Y13_N4BEG[14] ;
 wire \Tile_X6Y13_N4BEG[15] ;
 wire \Tile_X6Y13_N4BEG[1] ;
 wire \Tile_X6Y13_N4BEG[2] ;
 wire \Tile_X6Y13_N4BEG[3] ;
 wire \Tile_X6Y13_N4BEG[4] ;
 wire \Tile_X6Y13_N4BEG[5] ;
 wire \Tile_X6Y13_N4BEG[6] ;
 wire \Tile_X6Y13_N4BEG[7] ;
 wire \Tile_X6Y13_N4BEG[8] ;
 wire \Tile_X6Y13_N4BEG[9] ;
 wire \Tile_X6Y13_NN4BEG[0] ;
 wire \Tile_X6Y13_NN4BEG[10] ;
 wire \Tile_X6Y13_NN4BEG[11] ;
 wire \Tile_X6Y13_NN4BEG[12] ;
 wire \Tile_X6Y13_NN4BEG[13] ;
 wire \Tile_X6Y13_NN4BEG[14] ;
 wire \Tile_X6Y13_NN4BEG[15] ;
 wire \Tile_X6Y13_NN4BEG[1] ;
 wire \Tile_X6Y13_NN4BEG[2] ;
 wire \Tile_X6Y13_NN4BEG[3] ;
 wire \Tile_X6Y13_NN4BEG[4] ;
 wire \Tile_X6Y13_NN4BEG[5] ;
 wire \Tile_X6Y13_NN4BEG[6] ;
 wire \Tile_X6Y13_NN4BEG[7] ;
 wire \Tile_X6Y13_NN4BEG[8] ;
 wire \Tile_X6Y13_NN4BEG[9] ;
 wire \Tile_X6Y13_S1BEG[0] ;
 wire \Tile_X6Y13_S1BEG[1] ;
 wire \Tile_X6Y13_S1BEG[2] ;
 wire \Tile_X6Y13_S1BEG[3] ;
 wire \Tile_X6Y13_S2BEG[0] ;
 wire \Tile_X6Y13_S2BEG[1] ;
 wire \Tile_X6Y13_S2BEG[2] ;
 wire \Tile_X6Y13_S2BEG[3] ;
 wire \Tile_X6Y13_S2BEG[4] ;
 wire \Tile_X6Y13_S2BEG[5] ;
 wire \Tile_X6Y13_S2BEG[6] ;
 wire \Tile_X6Y13_S2BEG[7] ;
 wire \Tile_X6Y13_S2BEGb[0] ;
 wire \Tile_X6Y13_S2BEGb[1] ;
 wire \Tile_X6Y13_S2BEGb[2] ;
 wire \Tile_X6Y13_S2BEGb[3] ;
 wire \Tile_X6Y13_S2BEGb[4] ;
 wire \Tile_X6Y13_S2BEGb[5] ;
 wire \Tile_X6Y13_S2BEGb[6] ;
 wire \Tile_X6Y13_S2BEGb[7] ;
 wire \Tile_X6Y13_S4BEG[0] ;
 wire \Tile_X6Y13_S4BEG[10] ;
 wire \Tile_X6Y13_S4BEG[11] ;
 wire \Tile_X6Y13_S4BEG[12] ;
 wire \Tile_X6Y13_S4BEG[13] ;
 wire \Tile_X6Y13_S4BEG[14] ;
 wire \Tile_X6Y13_S4BEG[15] ;
 wire \Tile_X6Y13_S4BEG[1] ;
 wire \Tile_X6Y13_S4BEG[2] ;
 wire \Tile_X6Y13_S4BEG[3] ;
 wire \Tile_X6Y13_S4BEG[4] ;
 wire \Tile_X6Y13_S4BEG[5] ;
 wire \Tile_X6Y13_S4BEG[6] ;
 wire \Tile_X6Y13_S4BEG[7] ;
 wire \Tile_X6Y13_S4BEG[8] ;
 wire \Tile_X6Y13_S4BEG[9] ;
 wire \Tile_X6Y13_SS4BEG[0] ;
 wire \Tile_X6Y13_SS4BEG[10] ;
 wire \Tile_X6Y13_SS4BEG[11] ;
 wire \Tile_X6Y13_SS4BEG[12] ;
 wire \Tile_X6Y13_SS4BEG[13] ;
 wire \Tile_X6Y13_SS4BEG[14] ;
 wire \Tile_X6Y13_SS4BEG[15] ;
 wire \Tile_X6Y13_SS4BEG[1] ;
 wire \Tile_X6Y13_SS4BEG[2] ;
 wire \Tile_X6Y13_SS4BEG[3] ;
 wire \Tile_X6Y13_SS4BEG[4] ;
 wire \Tile_X6Y13_SS4BEG[5] ;
 wire \Tile_X6Y13_SS4BEG[6] ;
 wire \Tile_X6Y13_SS4BEG[7] ;
 wire \Tile_X6Y13_SS4BEG[8] ;
 wire \Tile_X6Y13_SS4BEG[9] ;
 wire Tile_X6Y13_UserCLKo;
 wire \Tile_X6Y13_W1BEG[0] ;
 wire \Tile_X6Y13_W1BEG[1] ;
 wire \Tile_X6Y13_W1BEG[2] ;
 wire \Tile_X6Y13_W1BEG[3] ;
 wire \Tile_X6Y13_W2BEG[0] ;
 wire \Tile_X6Y13_W2BEG[1] ;
 wire \Tile_X6Y13_W2BEG[2] ;
 wire \Tile_X6Y13_W2BEG[3] ;
 wire \Tile_X6Y13_W2BEG[4] ;
 wire \Tile_X6Y13_W2BEG[5] ;
 wire \Tile_X6Y13_W2BEG[6] ;
 wire \Tile_X6Y13_W2BEG[7] ;
 wire \Tile_X6Y13_W2BEGb[0] ;
 wire \Tile_X6Y13_W2BEGb[1] ;
 wire \Tile_X6Y13_W2BEGb[2] ;
 wire \Tile_X6Y13_W2BEGb[3] ;
 wire \Tile_X6Y13_W2BEGb[4] ;
 wire \Tile_X6Y13_W2BEGb[5] ;
 wire \Tile_X6Y13_W2BEGb[6] ;
 wire \Tile_X6Y13_W2BEGb[7] ;
 wire \Tile_X6Y13_W6BEG[0] ;
 wire \Tile_X6Y13_W6BEG[10] ;
 wire \Tile_X6Y13_W6BEG[11] ;
 wire \Tile_X6Y13_W6BEG[1] ;
 wire \Tile_X6Y13_W6BEG[2] ;
 wire \Tile_X6Y13_W6BEG[3] ;
 wire \Tile_X6Y13_W6BEG[4] ;
 wire \Tile_X6Y13_W6BEG[5] ;
 wire \Tile_X6Y13_W6BEG[6] ;
 wire \Tile_X6Y13_W6BEG[7] ;
 wire \Tile_X6Y13_W6BEG[8] ;
 wire \Tile_X6Y13_W6BEG[9] ;
 wire \Tile_X6Y13_WW4BEG[0] ;
 wire \Tile_X6Y13_WW4BEG[10] ;
 wire \Tile_X6Y13_WW4BEG[11] ;
 wire \Tile_X6Y13_WW4BEG[12] ;
 wire \Tile_X6Y13_WW4BEG[13] ;
 wire \Tile_X6Y13_WW4BEG[14] ;
 wire \Tile_X6Y13_WW4BEG[15] ;
 wire \Tile_X6Y13_WW4BEG[1] ;
 wire \Tile_X6Y13_WW4BEG[2] ;
 wire \Tile_X6Y13_WW4BEG[3] ;
 wire \Tile_X6Y13_WW4BEG[4] ;
 wire \Tile_X6Y13_WW4BEG[5] ;
 wire \Tile_X6Y13_WW4BEG[6] ;
 wire \Tile_X6Y13_WW4BEG[7] ;
 wire \Tile_X6Y13_WW4BEG[8] ;
 wire \Tile_X6Y13_WW4BEG[9] ;
 wire Tile_X6Y14_Co;
 wire \Tile_X6Y14_E1BEG[0] ;
 wire \Tile_X6Y14_E1BEG[1] ;
 wire \Tile_X6Y14_E1BEG[2] ;
 wire \Tile_X6Y14_E1BEG[3] ;
 wire \Tile_X6Y14_E2BEG[0] ;
 wire \Tile_X6Y14_E2BEG[1] ;
 wire \Tile_X6Y14_E2BEG[2] ;
 wire \Tile_X6Y14_E2BEG[3] ;
 wire \Tile_X6Y14_E2BEG[4] ;
 wire \Tile_X6Y14_E2BEG[5] ;
 wire \Tile_X6Y14_E2BEG[6] ;
 wire \Tile_X6Y14_E2BEG[7] ;
 wire \Tile_X6Y14_E2BEGb[0] ;
 wire \Tile_X6Y14_E2BEGb[1] ;
 wire \Tile_X6Y14_E2BEGb[2] ;
 wire \Tile_X6Y14_E2BEGb[3] ;
 wire \Tile_X6Y14_E2BEGb[4] ;
 wire \Tile_X6Y14_E2BEGb[5] ;
 wire \Tile_X6Y14_E2BEGb[6] ;
 wire \Tile_X6Y14_E2BEGb[7] ;
 wire \Tile_X6Y14_E6BEG[0] ;
 wire \Tile_X6Y14_E6BEG[10] ;
 wire \Tile_X6Y14_E6BEG[11] ;
 wire \Tile_X6Y14_E6BEG[1] ;
 wire \Tile_X6Y14_E6BEG[2] ;
 wire \Tile_X6Y14_E6BEG[3] ;
 wire \Tile_X6Y14_E6BEG[4] ;
 wire \Tile_X6Y14_E6BEG[5] ;
 wire \Tile_X6Y14_E6BEG[6] ;
 wire \Tile_X6Y14_E6BEG[7] ;
 wire \Tile_X6Y14_E6BEG[8] ;
 wire \Tile_X6Y14_E6BEG[9] ;
 wire \Tile_X6Y14_EE4BEG[0] ;
 wire \Tile_X6Y14_EE4BEG[10] ;
 wire \Tile_X6Y14_EE4BEG[11] ;
 wire \Tile_X6Y14_EE4BEG[12] ;
 wire \Tile_X6Y14_EE4BEG[13] ;
 wire \Tile_X6Y14_EE4BEG[14] ;
 wire \Tile_X6Y14_EE4BEG[15] ;
 wire \Tile_X6Y14_EE4BEG[1] ;
 wire \Tile_X6Y14_EE4BEG[2] ;
 wire \Tile_X6Y14_EE4BEG[3] ;
 wire \Tile_X6Y14_EE4BEG[4] ;
 wire \Tile_X6Y14_EE4BEG[5] ;
 wire \Tile_X6Y14_EE4BEG[6] ;
 wire \Tile_X6Y14_EE4BEG[7] ;
 wire \Tile_X6Y14_EE4BEG[8] ;
 wire \Tile_X6Y14_EE4BEG[9] ;
 wire \Tile_X6Y14_FrameData_O[0] ;
 wire \Tile_X6Y14_FrameData_O[10] ;
 wire \Tile_X6Y14_FrameData_O[11] ;
 wire \Tile_X6Y14_FrameData_O[12] ;
 wire \Tile_X6Y14_FrameData_O[13] ;
 wire \Tile_X6Y14_FrameData_O[14] ;
 wire \Tile_X6Y14_FrameData_O[15] ;
 wire \Tile_X6Y14_FrameData_O[16] ;
 wire \Tile_X6Y14_FrameData_O[17] ;
 wire \Tile_X6Y14_FrameData_O[18] ;
 wire \Tile_X6Y14_FrameData_O[19] ;
 wire \Tile_X6Y14_FrameData_O[1] ;
 wire \Tile_X6Y14_FrameData_O[20] ;
 wire \Tile_X6Y14_FrameData_O[21] ;
 wire \Tile_X6Y14_FrameData_O[22] ;
 wire \Tile_X6Y14_FrameData_O[23] ;
 wire \Tile_X6Y14_FrameData_O[24] ;
 wire \Tile_X6Y14_FrameData_O[25] ;
 wire \Tile_X6Y14_FrameData_O[26] ;
 wire \Tile_X6Y14_FrameData_O[27] ;
 wire \Tile_X6Y14_FrameData_O[28] ;
 wire \Tile_X6Y14_FrameData_O[29] ;
 wire \Tile_X6Y14_FrameData_O[2] ;
 wire \Tile_X6Y14_FrameData_O[30] ;
 wire \Tile_X6Y14_FrameData_O[31] ;
 wire \Tile_X6Y14_FrameData_O[3] ;
 wire \Tile_X6Y14_FrameData_O[4] ;
 wire \Tile_X6Y14_FrameData_O[5] ;
 wire \Tile_X6Y14_FrameData_O[6] ;
 wire \Tile_X6Y14_FrameData_O[7] ;
 wire \Tile_X6Y14_FrameData_O[8] ;
 wire \Tile_X6Y14_FrameData_O[9] ;
 wire \Tile_X6Y14_FrameStrobe_O[0] ;
 wire \Tile_X6Y14_FrameStrobe_O[10] ;
 wire \Tile_X6Y14_FrameStrobe_O[11] ;
 wire \Tile_X6Y14_FrameStrobe_O[12] ;
 wire \Tile_X6Y14_FrameStrobe_O[13] ;
 wire \Tile_X6Y14_FrameStrobe_O[14] ;
 wire \Tile_X6Y14_FrameStrobe_O[15] ;
 wire \Tile_X6Y14_FrameStrobe_O[16] ;
 wire \Tile_X6Y14_FrameStrobe_O[17] ;
 wire \Tile_X6Y14_FrameStrobe_O[18] ;
 wire \Tile_X6Y14_FrameStrobe_O[19] ;
 wire \Tile_X6Y14_FrameStrobe_O[1] ;
 wire \Tile_X6Y14_FrameStrobe_O[2] ;
 wire \Tile_X6Y14_FrameStrobe_O[3] ;
 wire \Tile_X6Y14_FrameStrobe_O[4] ;
 wire \Tile_X6Y14_FrameStrobe_O[5] ;
 wire \Tile_X6Y14_FrameStrobe_O[6] ;
 wire \Tile_X6Y14_FrameStrobe_O[7] ;
 wire \Tile_X6Y14_FrameStrobe_O[8] ;
 wire \Tile_X6Y14_FrameStrobe_O[9] ;
 wire \Tile_X6Y14_N1BEG[0] ;
 wire \Tile_X6Y14_N1BEG[1] ;
 wire \Tile_X6Y14_N1BEG[2] ;
 wire \Tile_X6Y14_N1BEG[3] ;
 wire \Tile_X6Y14_N2BEG[0] ;
 wire \Tile_X6Y14_N2BEG[1] ;
 wire \Tile_X6Y14_N2BEG[2] ;
 wire \Tile_X6Y14_N2BEG[3] ;
 wire \Tile_X6Y14_N2BEG[4] ;
 wire \Tile_X6Y14_N2BEG[5] ;
 wire \Tile_X6Y14_N2BEG[6] ;
 wire \Tile_X6Y14_N2BEG[7] ;
 wire \Tile_X6Y14_N2BEGb[0] ;
 wire \Tile_X6Y14_N2BEGb[1] ;
 wire \Tile_X6Y14_N2BEGb[2] ;
 wire \Tile_X6Y14_N2BEGb[3] ;
 wire \Tile_X6Y14_N2BEGb[4] ;
 wire \Tile_X6Y14_N2BEGb[5] ;
 wire \Tile_X6Y14_N2BEGb[6] ;
 wire \Tile_X6Y14_N2BEGb[7] ;
 wire \Tile_X6Y14_N4BEG[0] ;
 wire \Tile_X6Y14_N4BEG[10] ;
 wire \Tile_X6Y14_N4BEG[11] ;
 wire \Tile_X6Y14_N4BEG[12] ;
 wire \Tile_X6Y14_N4BEG[13] ;
 wire \Tile_X6Y14_N4BEG[14] ;
 wire \Tile_X6Y14_N4BEG[15] ;
 wire \Tile_X6Y14_N4BEG[1] ;
 wire \Tile_X6Y14_N4BEG[2] ;
 wire \Tile_X6Y14_N4BEG[3] ;
 wire \Tile_X6Y14_N4BEG[4] ;
 wire \Tile_X6Y14_N4BEG[5] ;
 wire \Tile_X6Y14_N4BEG[6] ;
 wire \Tile_X6Y14_N4BEG[7] ;
 wire \Tile_X6Y14_N4BEG[8] ;
 wire \Tile_X6Y14_N4BEG[9] ;
 wire \Tile_X6Y14_NN4BEG[0] ;
 wire \Tile_X6Y14_NN4BEG[10] ;
 wire \Tile_X6Y14_NN4BEG[11] ;
 wire \Tile_X6Y14_NN4BEG[12] ;
 wire \Tile_X6Y14_NN4BEG[13] ;
 wire \Tile_X6Y14_NN4BEG[14] ;
 wire \Tile_X6Y14_NN4BEG[15] ;
 wire \Tile_X6Y14_NN4BEG[1] ;
 wire \Tile_X6Y14_NN4BEG[2] ;
 wire \Tile_X6Y14_NN4BEG[3] ;
 wire \Tile_X6Y14_NN4BEG[4] ;
 wire \Tile_X6Y14_NN4BEG[5] ;
 wire \Tile_X6Y14_NN4BEG[6] ;
 wire \Tile_X6Y14_NN4BEG[7] ;
 wire \Tile_X6Y14_NN4BEG[8] ;
 wire \Tile_X6Y14_NN4BEG[9] ;
 wire \Tile_X6Y14_S1BEG[0] ;
 wire \Tile_X6Y14_S1BEG[1] ;
 wire \Tile_X6Y14_S1BEG[2] ;
 wire \Tile_X6Y14_S1BEG[3] ;
 wire \Tile_X6Y14_S2BEG[0] ;
 wire \Tile_X6Y14_S2BEG[1] ;
 wire \Tile_X6Y14_S2BEG[2] ;
 wire \Tile_X6Y14_S2BEG[3] ;
 wire \Tile_X6Y14_S2BEG[4] ;
 wire \Tile_X6Y14_S2BEG[5] ;
 wire \Tile_X6Y14_S2BEG[6] ;
 wire \Tile_X6Y14_S2BEG[7] ;
 wire \Tile_X6Y14_S2BEGb[0] ;
 wire \Tile_X6Y14_S2BEGb[1] ;
 wire \Tile_X6Y14_S2BEGb[2] ;
 wire \Tile_X6Y14_S2BEGb[3] ;
 wire \Tile_X6Y14_S2BEGb[4] ;
 wire \Tile_X6Y14_S2BEGb[5] ;
 wire \Tile_X6Y14_S2BEGb[6] ;
 wire \Tile_X6Y14_S2BEGb[7] ;
 wire \Tile_X6Y14_S4BEG[0] ;
 wire \Tile_X6Y14_S4BEG[10] ;
 wire \Tile_X6Y14_S4BEG[11] ;
 wire \Tile_X6Y14_S4BEG[12] ;
 wire \Tile_X6Y14_S4BEG[13] ;
 wire \Tile_X6Y14_S4BEG[14] ;
 wire \Tile_X6Y14_S4BEG[15] ;
 wire \Tile_X6Y14_S4BEG[1] ;
 wire \Tile_X6Y14_S4BEG[2] ;
 wire \Tile_X6Y14_S4BEG[3] ;
 wire \Tile_X6Y14_S4BEG[4] ;
 wire \Tile_X6Y14_S4BEG[5] ;
 wire \Tile_X6Y14_S4BEG[6] ;
 wire \Tile_X6Y14_S4BEG[7] ;
 wire \Tile_X6Y14_S4BEG[8] ;
 wire \Tile_X6Y14_S4BEG[9] ;
 wire \Tile_X6Y14_SS4BEG[0] ;
 wire \Tile_X6Y14_SS4BEG[10] ;
 wire \Tile_X6Y14_SS4BEG[11] ;
 wire \Tile_X6Y14_SS4BEG[12] ;
 wire \Tile_X6Y14_SS4BEG[13] ;
 wire \Tile_X6Y14_SS4BEG[14] ;
 wire \Tile_X6Y14_SS4BEG[15] ;
 wire \Tile_X6Y14_SS4BEG[1] ;
 wire \Tile_X6Y14_SS4BEG[2] ;
 wire \Tile_X6Y14_SS4BEG[3] ;
 wire \Tile_X6Y14_SS4BEG[4] ;
 wire \Tile_X6Y14_SS4BEG[5] ;
 wire \Tile_X6Y14_SS4BEG[6] ;
 wire \Tile_X6Y14_SS4BEG[7] ;
 wire \Tile_X6Y14_SS4BEG[8] ;
 wire \Tile_X6Y14_SS4BEG[9] ;
 wire Tile_X6Y14_UserCLKo;
 wire \Tile_X6Y14_W1BEG[0] ;
 wire \Tile_X6Y14_W1BEG[1] ;
 wire \Tile_X6Y14_W1BEG[2] ;
 wire \Tile_X6Y14_W1BEG[3] ;
 wire \Tile_X6Y14_W2BEG[0] ;
 wire \Tile_X6Y14_W2BEG[1] ;
 wire \Tile_X6Y14_W2BEG[2] ;
 wire \Tile_X6Y14_W2BEG[3] ;
 wire \Tile_X6Y14_W2BEG[4] ;
 wire \Tile_X6Y14_W2BEG[5] ;
 wire \Tile_X6Y14_W2BEG[6] ;
 wire \Tile_X6Y14_W2BEG[7] ;
 wire \Tile_X6Y14_W2BEGb[0] ;
 wire \Tile_X6Y14_W2BEGb[1] ;
 wire \Tile_X6Y14_W2BEGb[2] ;
 wire \Tile_X6Y14_W2BEGb[3] ;
 wire \Tile_X6Y14_W2BEGb[4] ;
 wire \Tile_X6Y14_W2BEGb[5] ;
 wire \Tile_X6Y14_W2BEGb[6] ;
 wire \Tile_X6Y14_W2BEGb[7] ;
 wire \Tile_X6Y14_W6BEG[0] ;
 wire \Tile_X6Y14_W6BEG[10] ;
 wire \Tile_X6Y14_W6BEG[11] ;
 wire \Tile_X6Y14_W6BEG[1] ;
 wire \Tile_X6Y14_W6BEG[2] ;
 wire \Tile_X6Y14_W6BEG[3] ;
 wire \Tile_X6Y14_W6BEG[4] ;
 wire \Tile_X6Y14_W6BEG[5] ;
 wire \Tile_X6Y14_W6BEG[6] ;
 wire \Tile_X6Y14_W6BEG[7] ;
 wire \Tile_X6Y14_W6BEG[8] ;
 wire \Tile_X6Y14_W6BEG[9] ;
 wire \Tile_X6Y14_WW4BEG[0] ;
 wire \Tile_X6Y14_WW4BEG[10] ;
 wire \Tile_X6Y14_WW4BEG[11] ;
 wire \Tile_X6Y14_WW4BEG[12] ;
 wire \Tile_X6Y14_WW4BEG[13] ;
 wire \Tile_X6Y14_WW4BEG[14] ;
 wire \Tile_X6Y14_WW4BEG[15] ;
 wire \Tile_X6Y14_WW4BEG[1] ;
 wire \Tile_X6Y14_WW4BEG[2] ;
 wire \Tile_X6Y14_WW4BEG[3] ;
 wire \Tile_X6Y14_WW4BEG[4] ;
 wire \Tile_X6Y14_WW4BEG[5] ;
 wire \Tile_X6Y14_WW4BEG[6] ;
 wire \Tile_X6Y14_WW4BEG[7] ;
 wire \Tile_X6Y14_WW4BEG[8] ;
 wire \Tile_X6Y14_WW4BEG[9] ;
 wire Tile_X6Y15_Co;
 wire \Tile_X6Y15_FrameData_O[0] ;
 wire \Tile_X6Y15_FrameData_O[10] ;
 wire \Tile_X6Y15_FrameData_O[11] ;
 wire \Tile_X6Y15_FrameData_O[12] ;
 wire \Tile_X6Y15_FrameData_O[13] ;
 wire \Tile_X6Y15_FrameData_O[14] ;
 wire \Tile_X6Y15_FrameData_O[15] ;
 wire \Tile_X6Y15_FrameData_O[16] ;
 wire \Tile_X6Y15_FrameData_O[17] ;
 wire \Tile_X6Y15_FrameData_O[18] ;
 wire \Tile_X6Y15_FrameData_O[19] ;
 wire \Tile_X6Y15_FrameData_O[1] ;
 wire \Tile_X6Y15_FrameData_O[20] ;
 wire \Tile_X6Y15_FrameData_O[21] ;
 wire \Tile_X6Y15_FrameData_O[22] ;
 wire \Tile_X6Y15_FrameData_O[23] ;
 wire \Tile_X6Y15_FrameData_O[24] ;
 wire \Tile_X6Y15_FrameData_O[25] ;
 wire \Tile_X6Y15_FrameData_O[26] ;
 wire \Tile_X6Y15_FrameData_O[27] ;
 wire \Tile_X6Y15_FrameData_O[28] ;
 wire \Tile_X6Y15_FrameData_O[29] ;
 wire \Tile_X6Y15_FrameData_O[2] ;
 wire \Tile_X6Y15_FrameData_O[30] ;
 wire \Tile_X6Y15_FrameData_O[31] ;
 wire \Tile_X6Y15_FrameData_O[3] ;
 wire \Tile_X6Y15_FrameData_O[4] ;
 wire \Tile_X6Y15_FrameData_O[5] ;
 wire \Tile_X6Y15_FrameData_O[6] ;
 wire \Tile_X6Y15_FrameData_O[7] ;
 wire \Tile_X6Y15_FrameData_O[8] ;
 wire \Tile_X6Y15_FrameData_O[9] ;
 wire \Tile_X6Y15_FrameStrobe_O[0] ;
 wire \Tile_X6Y15_FrameStrobe_O[10] ;
 wire \Tile_X6Y15_FrameStrobe_O[11] ;
 wire \Tile_X6Y15_FrameStrobe_O[12] ;
 wire \Tile_X6Y15_FrameStrobe_O[13] ;
 wire \Tile_X6Y15_FrameStrobe_O[14] ;
 wire \Tile_X6Y15_FrameStrobe_O[15] ;
 wire \Tile_X6Y15_FrameStrobe_O[16] ;
 wire \Tile_X6Y15_FrameStrobe_O[17] ;
 wire \Tile_X6Y15_FrameStrobe_O[18] ;
 wire \Tile_X6Y15_FrameStrobe_O[19] ;
 wire \Tile_X6Y15_FrameStrobe_O[1] ;
 wire \Tile_X6Y15_FrameStrobe_O[2] ;
 wire \Tile_X6Y15_FrameStrobe_O[3] ;
 wire \Tile_X6Y15_FrameStrobe_O[4] ;
 wire \Tile_X6Y15_FrameStrobe_O[5] ;
 wire \Tile_X6Y15_FrameStrobe_O[6] ;
 wire \Tile_X6Y15_FrameStrobe_O[7] ;
 wire \Tile_X6Y15_FrameStrobe_O[8] ;
 wire \Tile_X6Y15_FrameStrobe_O[9] ;
 wire \Tile_X6Y15_N1BEG[0] ;
 wire \Tile_X6Y15_N1BEG[1] ;
 wire \Tile_X6Y15_N1BEG[2] ;
 wire \Tile_X6Y15_N1BEG[3] ;
 wire \Tile_X6Y15_N2BEG[0] ;
 wire \Tile_X6Y15_N2BEG[1] ;
 wire \Tile_X6Y15_N2BEG[2] ;
 wire \Tile_X6Y15_N2BEG[3] ;
 wire \Tile_X6Y15_N2BEG[4] ;
 wire \Tile_X6Y15_N2BEG[5] ;
 wire \Tile_X6Y15_N2BEG[6] ;
 wire \Tile_X6Y15_N2BEG[7] ;
 wire \Tile_X6Y15_N2BEGb[0] ;
 wire \Tile_X6Y15_N2BEGb[1] ;
 wire \Tile_X6Y15_N2BEGb[2] ;
 wire \Tile_X6Y15_N2BEGb[3] ;
 wire \Tile_X6Y15_N2BEGb[4] ;
 wire \Tile_X6Y15_N2BEGb[5] ;
 wire \Tile_X6Y15_N2BEGb[6] ;
 wire \Tile_X6Y15_N2BEGb[7] ;
 wire \Tile_X6Y15_N4BEG[0] ;
 wire \Tile_X6Y15_N4BEG[10] ;
 wire \Tile_X6Y15_N4BEG[11] ;
 wire \Tile_X6Y15_N4BEG[12] ;
 wire \Tile_X6Y15_N4BEG[13] ;
 wire \Tile_X6Y15_N4BEG[14] ;
 wire \Tile_X6Y15_N4BEG[15] ;
 wire \Tile_X6Y15_N4BEG[1] ;
 wire \Tile_X6Y15_N4BEG[2] ;
 wire \Tile_X6Y15_N4BEG[3] ;
 wire \Tile_X6Y15_N4BEG[4] ;
 wire \Tile_X6Y15_N4BEG[5] ;
 wire \Tile_X6Y15_N4BEG[6] ;
 wire \Tile_X6Y15_N4BEG[7] ;
 wire \Tile_X6Y15_N4BEG[8] ;
 wire \Tile_X6Y15_N4BEG[9] ;
 wire \Tile_X6Y15_NN4BEG[0] ;
 wire \Tile_X6Y15_NN4BEG[10] ;
 wire \Tile_X6Y15_NN4BEG[11] ;
 wire \Tile_X6Y15_NN4BEG[12] ;
 wire \Tile_X6Y15_NN4BEG[13] ;
 wire \Tile_X6Y15_NN4BEG[14] ;
 wire \Tile_X6Y15_NN4BEG[15] ;
 wire \Tile_X6Y15_NN4BEG[1] ;
 wire \Tile_X6Y15_NN4BEG[2] ;
 wire \Tile_X6Y15_NN4BEG[3] ;
 wire \Tile_X6Y15_NN4BEG[4] ;
 wire \Tile_X6Y15_NN4BEG[5] ;
 wire \Tile_X6Y15_NN4BEG[6] ;
 wire \Tile_X6Y15_NN4BEG[7] ;
 wire \Tile_X6Y15_NN4BEG[8] ;
 wire \Tile_X6Y15_NN4BEG[9] ;
 wire Tile_X6Y15_UserCLKo;
 wire Tile_X6Y1_Co;
 wire \Tile_X6Y1_E1BEG[0] ;
 wire \Tile_X6Y1_E1BEG[1] ;
 wire \Tile_X6Y1_E1BEG[2] ;
 wire \Tile_X6Y1_E1BEG[3] ;
 wire \Tile_X6Y1_E2BEG[0] ;
 wire \Tile_X6Y1_E2BEG[1] ;
 wire \Tile_X6Y1_E2BEG[2] ;
 wire \Tile_X6Y1_E2BEG[3] ;
 wire \Tile_X6Y1_E2BEG[4] ;
 wire \Tile_X6Y1_E2BEG[5] ;
 wire \Tile_X6Y1_E2BEG[6] ;
 wire \Tile_X6Y1_E2BEG[7] ;
 wire \Tile_X6Y1_E2BEGb[0] ;
 wire \Tile_X6Y1_E2BEGb[1] ;
 wire \Tile_X6Y1_E2BEGb[2] ;
 wire \Tile_X6Y1_E2BEGb[3] ;
 wire \Tile_X6Y1_E2BEGb[4] ;
 wire \Tile_X6Y1_E2BEGb[5] ;
 wire \Tile_X6Y1_E2BEGb[6] ;
 wire \Tile_X6Y1_E2BEGb[7] ;
 wire \Tile_X6Y1_E6BEG[0] ;
 wire \Tile_X6Y1_E6BEG[10] ;
 wire \Tile_X6Y1_E6BEG[11] ;
 wire \Tile_X6Y1_E6BEG[1] ;
 wire \Tile_X6Y1_E6BEG[2] ;
 wire \Tile_X6Y1_E6BEG[3] ;
 wire \Tile_X6Y1_E6BEG[4] ;
 wire \Tile_X6Y1_E6BEG[5] ;
 wire \Tile_X6Y1_E6BEG[6] ;
 wire \Tile_X6Y1_E6BEG[7] ;
 wire \Tile_X6Y1_E6BEG[8] ;
 wire \Tile_X6Y1_E6BEG[9] ;
 wire \Tile_X6Y1_EE4BEG[0] ;
 wire \Tile_X6Y1_EE4BEG[10] ;
 wire \Tile_X6Y1_EE4BEG[11] ;
 wire \Tile_X6Y1_EE4BEG[12] ;
 wire \Tile_X6Y1_EE4BEG[13] ;
 wire \Tile_X6Y1_EE4BEG[14] ;
 wire \Tile_X6Y1_EE4BEG[15] ;
 wire \Tile_X6Y1_EE4BEG[1] ;
 wire \Tile_X6Y1_EE4BEG[2] ;
 wire \Tile_X6Y1_EE4BEG[3] ;
 wire \Tile_X6Y1_EE4BEG[4] ;
 wire \Tile_X6Y1_EE4BEG[5] ;
 wire \Tile_X6Y1_EE4BEG[6] ;
 wire \Tile_X6Y1_EE4BEG[7] ;
 wire \Tile_X6Y1_EE4BEG[8] ;
 wire \Tile_X6Y1_EE4BEG[9] ;
 wire \Tile_X6Y1_FrameData_O[0] ;
 wire \Tile_X6Y1_FrameData_O[10] ;
 wire \Tile_X6Y1_FrameData_O[11] ;
 wire \Tile_X6Y1_FrameData_O[12] ;
 wire \Tile_X6Y1_FrameData_O[13] ;
 wire \Tile_X6Y1_FrameData_O[14] ;
 wire \Tile_X6Y1_FrameData_O[15] ;
 wire \Tile_X6Y1_FrameData_O[16] ;
 wire \Tile_X6Y1_FrameData_O[17] ;
 wire \Tile_X6Y1_FrameData_O[18] ;
 wire \Tile_X6Y1_FrameData_O[19] ;
 wire \Tile_X6Y1_FrameData_O[1] ;
 wire \Tile_X6Y1_FrameData_O[20] ;
 wire \Tile_X6Y1_FrameData_O[21] ;
 wire \Tile_X6Y1_FrameData_O[22] ;
 wire \Tile_X6Y1_FrameData_O[23] ;
 wire \Tile_X6Y1_FrameData_O[24] ;
 wire \Tile_X6Y1_FrameData_O[25] ;
 wire \Tile_X6Y1_FrameData_O[26] ;
 wire \Tile_X6Y1_FrameData_O[27] ;
 wire \Tile_X6Y1_FrameData_O[28] ;
 wire \Tile_X6Y1_FrameData_O[29] ;
 wire \Tile_X6Y1_FrameData_O[2] ;
 wire \Tile_X6Y1_FrameData_O[30] ;
 wire \Tile_X6Y1_FrameData_O[31] ;
 wire \Tile_X6Y1_FrameData_O[3] ;
 wire \Tile_X6Y1_FrameData_O[4] ;
 wire \Tile_X6Y1_FrameData_O[5] ;
 wire \Tile_X6Y1_FrameData_O[6] ;
 wire \Tile_X6Y1_FrameData_O[7] ;
 wire \Tile_X6Y1_FrameData_O[8] ;
 wire \Tile_X6Y1_FrameData_O[9] ;
 wire \Tile_X6Y1_FrameStrobe_O[0] ;
 wire \Tile_X6Y1_FrameStrobe_O[10] ;
 wire \Tile_X6Y1_FrameStrobe_O[11] ;
 wire \Tile_X6Y1_FrameStrobe_O[12] ;
 wire \Tile_X6Y1_FrameStrobe_O[13] ;
 wire \Tile_X6Y1_FrameStrobe_O[14] ;
 wire \Tile_X6Y1_FrameStrobe_O[15] ;
 wire \Tile_X6Y1_FrameStrobe_O[16] ;
 wire \Tile_X6Y1_FrameStrobe_O[17] ;
 wire \Tile_X6Y1_FrameStrobe_O[18] ;
 wire \Tile_X6Y1_FrameStrobe_O[19] ;
 wire \Tile_X6Y1_FrameStrobe_O[1] ;
 wire \Tile_X6Y1_FrameStrobe_O[2] ;
 wire \Tile_X6Y1_FrameStrobe_O[3] ;
 wire \Tile_X6Y1_FrameStrobe_O[4] ;
 wire \Tile_X6Y1_FrameStrobe_O[5] ;
 wire \Tile_X6Y1_FrameStrobe_O[6] ;
 wire \Tile_X6Y1_FrameStrobe_O[7] ;
 wire \Tile_X6Y1_FrameStrobe_O[8] ;
 wire \Tile_X6Y1_FrameStrobe_O[9] ;
 wire \Tile_X6Y1_N1BEG[0] ;
 wire \Tile_X6Y1_N1BEG[1] ;
 wire \Tile_X6Y1_N1BEG[2] ;
 wire \Tile_X6Y1_N1BEG[3] ;
 wire \Tile_X6Y1_N2BEG[0] ;
 wire \Tile_X6Y1_N2BEG[1] ;
 wire \Tile_X6Y1_N2BEG[2] ;
 wire \Tile_X6Y1_N2BEG[3] ;
 wire \Tile_X6Y1_N2BEG[4] ;
 wire \Tile_X6Y1_N2BEG[5] ;
 wire \Tile_X6Y1_N2BEG[6] ;
 wire \Tile_X6Y1_N2BEG[7] ;
 wire \Tile_X6Y1_N2BEGb[0] ;
 wire \Tile_X6Y1_N2BEGb[1] ;
 wire \Tile_X6Y1_N2BEGb[2] ;
 wire \Tile_X6Y1_N2BEGb[3] ;
 wire \Tile_X6Y1_N2BEGb[4] ;
 wire \Tile_X6Y1_N2BEGb[5] ;
 wire \Tile_X6Y1_N2BEGb[6] ;
 wire \Tile_X6Y1_N2BEGb[7] ;
 wire \Tile_X6Y1_N4BEG[0] ;
 wire \Tile_X6Y1_N4BEG[10] ;
 wire \Tile_X6Y1_N4BEG[11] ;
 wire \Tile_X6Y1_N4BEG[12] ;
 wire \Tile_X6Y1_N4BEG[13] ;
 wire \Tile_X6Y1_N4BEG[14] ;
 wire \Tile_X6Y1_N4BEG[15] ;
 wire \Tile_X6Y1_N4BEG[1] ;
 wire \Tile_X6Y1_N4BEG[2] ;
 wire \Tile_X6Y1_N4BEG[3] ;
 wire \Tile_X6Y1_N4BEG[4] ;
 wire \Tile_X6Y1_N4BEG[5] ;
 wire \Tile_X6Y1_N4BEG[6] ;
 wire \Tile_X6Y1_N4BEG[7] ;
 wire \Tile_X6Y1_N4BEG[8] ;
 wire \Tile_X6Y1_N4BEG[9] ;
 wire \Tile_X6Y1_NN4BEG[0] ;
 wire \Tile_X6Y1_NN4BEG[10] ;
 wire \Tile_X6Y1_NN4BEG[11] ;
 wire \Tile_X6Y1_NN4BEG[12] ;
 wire \Tile_X6Y1_NN4BEG[13] ;
 wire \Tile_X6Y1_NN4BEG[14] ;
 wire \Tile_X6Y1_NN4BEG[15] ;
 wire \Tile_X6Y1_NN4BEG[1] ;
 wire \Tile_X6Y1_NN4BEG[2] ;
 wire \Tile_X6Y1_NN4BEG[3] ;
 wire \Tile_X6Y1_NN4BEG[4] ;
 wire \Tile_X6Y1_NN4BEG[5] ;
 wire \Tile_X6Y1_NN4BEG[6] ;
 wire \Tile_X6Y1_NN4BEG[7] ;
 wire \Tile_X6Y1_NN4BEG[8] ;
 wire \Tile_X6Y1_NN4BEG[9] ;
 wire \Tile_X6Y1_S1BEG[0] ;
 wire \Tile_X6Y1_S1BEG[1] ;
 wire \Tile_X6Y1_S1BEG[2] ;
 wire \Tile_X6Y1_S1BEG[3] ;
 wire \Tile_X6Y1_S2BEG[0] ;
 wire \Tile_X6Y1_S2BEG[1] ;
 wire \Tile_X6Y1_S2BEG[2] ;
 wire \Tile_X6Y1_S2BEG[3] ;
 wire \Tile_X6Y1_S2BEG[4] ;
 wire \Tile_X6Y1_S2BEG[5] ;
 wire \Tile_X6Y1_S2BEG[6] ;
 wire \Tile_X6Y1_S2BEG[7] ;
 wire \Tile_X6Y1_S2BEGb[0] ;
 wire \Tile_X6Y1_S2BEGb[1] ;
 wire \Tile_X6Y1_S2BEGb[2] ;
 wire \Tile_X6Y1_S2BEGb[3] ;
 wire \Tile_X6Y1_S2BEGb[4] ;
 wire \Tile_X6Y1_S2BEGb[5] ;
 wire \Tile_X6Y1_S2BEGb[6] ;
 wire \Tile_X6Y1_S2BEGb[7] ;
 wire \Tile_X6Y1_S4BEG[0] ;
 wire \Tile_X6Y1_S4BEG[10] ;
 wire \Tile_X6Y1_S4BEG[11] ;
 wire \Tile_X6Y1_S4BEG[12] ;
 wire \Tile_X6Y1_S4BEG[13] ;
 wire \Tile_X6Y1_S4BEG[14] ;
 wire \Tile_X6Y1_S4BEG[15] ;
 wire \Tile_X6Y1_S4BEG[1] ;
 wire \Tile_X6Y1_S4BEG[2] ;
 wire \Tile_X6Y1_S4BEG[3] ;
 wire \Tile_X6Y1_S4BEG[4] ;
 wire \Tile_X6Y1_S4BEG[5] ;
 wire \Tile_X6Y1_S4BEG[6] ;
 wire \Tile_X6Y1_S4BEG[7] ;
 wire \Tile_X6Y1_S4BEG[8] ;
 wire \Tile_X6Y1_S4BEG[9] ;
 wire \Tile_X6Y1_SS4BEG[0] ;
 wire \Tile_X6Y1_SS4BEG[10] ;
 wire \Tile_X6Y1_SS4BEG[11] ;
 wire \Tile_X6Y1_SS4BEG[12] ;
 wire \Tile_X6Y1_SS4BEG[13] ;
 wire \Tile_X6Y1_SS4BEG[14] ;
 wire \Tile_X6Y1_SS4BEG[15] ;
 wire \Tile_X6Y1_SS4BEG[1] ;
 wire \Tile_X6Y1_SS4BEG[2] ;
 wire \Tile_X6Y1_SS4BEG[3] ;
 wire \Tile_X6Y1_SS4BEG[4] ;
 wire \Tile_X6Y1_SS4BEG[5] ;
 wire \Tile_X6Y1_SS4BEG[6] ;
 wire \Tile_X6Y1_SS4BEG[7] ;
 wire \Tile_X6Y1_SS4BEG[8] ;
 wire \Tile_X6Y1_SS4BEG[9] ;
 wire Tile_X6Y1_UserCLKo;
 wire \Tile_X6Y1_W1BEG[0] ;
 wire \Tile_X6Y1_W1BEG[1] ;
 wire \Tile_X6Y1_W1BEG[2] ;
 wire \Tile_X6Y1_W1BEG[3] ;
 wire \Tile_X6Y1_W2BEG[0] ;
 wire \Tile_X6Y1_W2BEG[1] ;
 wire \Tile_X6Y1_W2BEG[2] ;
 wire \Tile_X6Y1_W2BEG[3] ;
 wire \Tile_X6Y1_W2BEG[4] ;
 wire \Tile_X6Y1_W2BEG[5] ;
 wire \Tile_X6Y1_W2BEG[6] ;
 wire \Tile_X6Y1_W2BEG[7] ;
 wire \Tile_X6Y1_W2BEGb[0] ;
 wire \Tile_X6Y1_W2BEGb[1] ;
 wire \Tile_X6Y1_W2BEGb[2] ;
 wire \Tile_X6Y1_W2BEGb[3] ;
 wire \Tile_X6Y1_W2BEGb[4] ;
 wire \Tile_X6Y1_W2BEGb[5] ;
 wire \Tile_X6Y1_W2BEGb[6] ;
 wire \Tile_X6Y1_W2BEGb[7] ;
 wire \Tile_X6Y1_W6BEG[0] ;
 wire \Tile_X6Y1_W6BEG[10] ;
 wire \Tile_X6Y1_W6BEG[11] ;
 wire \Tile_X6Y1_W6BEG[1] ;
 wire \Tile_X6Y1_W6BEG[2] ;
 wire \Tile_X6Y1_W6BEG[3] ;
 wire \Tile_X6Y1_W6BEG[4] ;
 wire \Tile_X6Y1_W6BEG[5] ;
 wire \Tile_X6Y1_W6BEG[6] ;
 wire \Tile_X6Y1_W6BEG[7] ;
 wire \Tile_X6Y1_W6BEG[8] ;
 wire \Tile_X6Y1_W6BEG[9] ;
 wire \Tile_X6Y1_WW4BEG[0] ;
 wire \Tile_X6Y1_WW4BEG[10] ;
 wire \Tile_X6Y1_WW4BEG[11] ;
 wire \Tile_X6Y1_WW4BEG[12] ;
 wire \Tile_X6Y1_WW4BEG[13] ;
 wire \Tile_X6Y1_WW4BEG[14] ;
 wire \Tile_X6Y1_WW4BEG[15] ;
 wire \Tile_X6Y1_WW4BEG[1] ;
 wire \Tile_X6Y1_WW4BEG[2] ;
 wire \Tile_X6Y1_WW4BEG[3] ;
 wire \Tile_X6Y1_WW4BEG[4] ;
 wire \Tile_X6Y1_WW4BEG[5] ;
 wire \Tile_X6Y1_WW4BEG[6] ;
 wire \Tile_X6Y1_WW4BEG[7] ;
 wire \Tile_X6Y1_WW4BEG[8] ;
 wire \Tile_X6Y1_WW4BEG[9] ;
 wire Tile_X6Y2_Co;
 wire \Tile_X6Y2_E1BEG[0] ;
 wire \Tile_X6Y2_E1BEG[1] ;
 wire \Tile_X6Y2_E1BEG[2] ;
 wire \Tile_X6Y2_E1BEG[3] ;
 wire \Tile_X6Y2_E2BEG[0] ;
 wire \Tile_X6Y2_E2BEG[1] ;
 wire \Tile_X6Y2_E2BEG[2] ;
 wire \Tile_X6Y2_E2BEG[3] ;
 wire \Tile_X6Y2_E2BEG[4] ;
 wire \Tile_X6Y2_E2BEG[5] ;
 wire \Tile_X6Y2_E2BEG[6] ;
 wire \Tile_X6Y2_E2BEG[7] ;
 wire \Tile_X6Y2_E2BEGb[0] ;
 wire \Tile_X6Y2_E2BEGb[1] ;
 wire \Tile_X6Y2_E2BEGb[2] ;
 wire \Tile_X6Y2_E2BEGb[3] ;
 wire \Tile_X6Y2_E2BEGb[4] ;
 wire \Tile_X6Y2_E2BEGb[5] ;
 wire \Tile_X6Y2_E2BEGb[6] ;
 wire \Tile_X6Y2_E2BEGb[7] ;
 wire \Tile_X6Y2_E6BEG[0] ;
 wire \Tile_X6Y2_E6BEG[10] ;
 wire \Tile_X6Y2_E6BEG[11] ;
 wire \Tile_X6Y2_E6BEG[1] ;
 wire \Tile_X6Y2_E6BEG[2] ;
 wire \Tile_X6Y2_E6BEG[3] ;
 wire \Tile_X6Y2_E6BEG[4] ;
 wire \Tile_X6Y2_E6BEG[5] ;
 wire \Tile_X6Y2_E6BEG[6] ;
 wire \Tile_X6Y2_E6BEG[7] ;
 wire \Tile_X6Y2_E6BEG[8] ;
 wire \Tile_X6Y2_E6BEG[9] ;
 wire \Tile_X6Y2_EE4BEG[0] ;
 wire \Tile_X6Y2_EE4BEG[10] ;
 wire \Tile_X6Y2_EE4BEG[11] ;
 wire \Tile_X6Y2_EE4BEG[12] ;
 wire \Tile_X6Y2_EE4BEG[13] ;
 wire \Tile_X6Y2_EE4BEG[14] ;
 wire \Tile_X6Y2_EE4BEG[15] ;
 wire \Tile_X6Y2_EE4BEG[1] ;
 wire \Tile_X6Y2_EE4BEG[2] ;
 wire \Tile_X6Y2_EE4BEG[3] ;
 wire \Tile_X6Y2_EE4BEG[4] ;
 wire \Tile_X6Y2_EE4BEG[5] ;
 wire \Tile_X6Y2_EE4BEG[6] ;
 wire \Tile_X6Y2_EE4BEG[7] ;
 wire \Tile_X6Y2_EE4BEG[8] ;
 wire \Tile_X6Y2_EE4BEG[9] ;
 wire \Tile_X6Y2_FrameData_O[0] ;
 wire \Tile_X6Y2_FrameData_O[10] ;
 wire \Tile_X6Y2_FrameData_O[11] ;
 wire \Tile_X6Y2_FrameData_O[12] ;
 wire \Tile_X6Y2_FrameData_O[13] ;
 wire \Tile_X6Y2_FrameData_O[14] ;
 wire \Tile_X6Y2_FrameData_O[15] ;
 wire \Tile_X6Y2_FrameData_O[16] ;
 wire \Tile_X6Y2_FrameData_O[17] ;
 wire \Tile_X6Y2_FrameData_O[18] ;
 wire \Tile_X6Y2_FrameData_O[19] ;
 wire \Tile_X6Y2_FrameData_O[1] ;
 wire \Tile_X6Y2_FrameData_O[20] ;
 wire \Tile_X6Y2_FrameData_O[21] ;
 wire \Tile_X6Y2_FrameData_O[22] ;
 wire \Tile_X6Y2_FrameData_O[23] ;
 wire \Tile_X6Y2_FrameData_O[24] ;
 wire \Tile_X6Y2_FrameData_O[25] ;
 wire \Tile_X6Y2_FrameData_O[26] ;
 wire \Tile_X6Y2_FrameData_O[27] ;
 wire \Tile_X6Y2_FrameData_O[28] ;
 wire \Tile_X6Y2_FrameData_O[29] ;
 wire \Tile_X6Y2_FrameData_O[2] ;
 wire \Tile_X6Y2_FrameData_O[30] ;
 wire \Tile_X6Y2_FrameData_O[31] ;
 wire \Tile_X6Y2_FrameData_O[3] ;
 wire \Tile_X6Y2_FrameData_O[4] ;
 wire \Tile_X6Y2_FrameData_O[5] ;
 wire \Tile_X6Y2_FrameData_O[6] ;
 wire \Tile_X6Y2_FrameData_O[7] ;
 wire \Tile_X6Y2_FrameData_O[8] ;
 wire \Tile_X6Y2_FrameData_O[9] ;
 wire \Tile_X6Y2_FrameStrobe_O[0] ;
 wire \Tile_X6Y2_FrameStrobe_O[10] ;
 wire \Tile_X6Y2_FrameStrobe_O[11] ;
 wire \Tile_X6Y2_FrameStrobe_O[12] ;
 wire \Tile_X6Y2_FrameStrobe_O[13] ;
 wire \Tile_X6Y2_FrameStrobe_O[14] ;
 wire \Tile_X6Y2_FrameStrobe_O[15] ;
 wire \Tile_X6Y2_FrameStrobe_O[16] ;
 wire \Tile_X6Y2_FrameStrobe_O[17] ;
 wire \Tile_X6Y2_FrameStrobe_O[18] ;
 wire \Tile_X6Y2_FrameStrobe_O[19] ;
 wire \Tile_X6Y2_FrameStrobe_O[1] ;
 wire \Tile_X6Y2_FrameStrobe_O[2] ;
 wire \Tile_X6Y2_FrameStrobe_O[3] ;
 wire \Tile_X6Y2_FrameStrobe_O[4] ;
 wire \Tile_X6Y2_FrameStrobe_O[5] ;
 wire \Tile_X6Y2_FrameStrobe_O[6] ;
 wire \Tile_X6Y2_FrameStrobe_O[7] ;
 wire \Tile_X6Y2_FrameStrobe_O[8] ;
 wire \Tile_X6Y2_FrameStrobe_O[9] ;
 wire \Tile_X6Y2_N1BEG[0] ;
 wire \Tile_X6Y2_N1BEG[1] ;
 wire \Tile_X6Y2_N1BEG[2] ;
 wire \Tile_X6Y2_N1BEG[3] ;
 wire \Tile_X6Y2_N2BEG[0] ;
 wire \Tile_X6Y2_N2BEG[1] ;
 wire \Tile_X6Y2_N2BEG[2] ;
 wire \Tile_X6Y2_N2BEG[3] ;
 wire \Tile_X6Y2_N2BEG[4] ;
 wire \Tile_X6Y2_N2BEG[5] ;
 wire \Tile_X6Y2_N2BEG[6] ;
 wire \Tile_X6Y2_N2BEG[7] ;
 wire \Tile_X6Y2_N2BEGb[0] ;
 wire \Tile_X6Y2_N2BEGb[1] ;
 wire \Tile_X6Y2_N2BEGb[2] ;
 wire \Tile_X6Y2_N2BEGb[3] ;
 wire \Tile_X6Y2_N2BEGb[4] ;
 wire \Tile_X6Y2_N2BEGb[5] ;
 wire \Tile_X6Y2_N2BEGb[6] ;
 wire \Tile_X6Y2_N2BEGb[7] ;
 wire \Tile_X6Y2_N4BEG[0] ;
 wire \Tile_X6Y2_N4BEG[10] ;
 wire \Tile_X6Y2_N4BEG[11] ;
 wire \Tile_X6Y2_N4BEG[12] ;
 wire \Tile_X6Y2_N4BEG[13] ;
 wire \Tile_X6Y2_N4BEG[14] ;
 wire \Tile_X6Y2_N4BEG[15] ;
 wire \Tile_X6Y2_N4BEG[1] ;
 wire \Tile_X6Y2_N4BEG[2] ;
 wire \Tile_X6Y2_N4BEG[3] ;
 wire \Tile_X6Y2_N4BEG[4] ;
 wire \Tile_X6Y2_N4BEG[5] ;
 wire \Tile_X6Y2_N4BEG[6] ;
 wire \Tile_X6Y2_N4BEG[7] ;
 wire \Tile_X6Y2_N4BEG[8] ;
 wire \Tile_X6Y2_N4BEG[9] ;
 wire \Tile_X6Y2_NN4BEG[0] ;
 wire \Tile_X6Y2_NN4BEG[10] ;
 wire \Tile_X6Y2_NN4BEG[11] ;
 wire \Tile_X6Y2_NN4BEG[12] ;
 wire \Tile_X6Y2_NN4BEG[13] ;
 wire \Tile_X6Y2_NN4BEG[14] ;
 wire \Tile_X6Y2_NN4BEG[15] ;
 wire \Tile_X6Y2_NN4BEG[1] ;
 wire \Tile_X6Y2_NN4BEG[2] ;
 wire \Tile_X6Y2_NN4BEG[3] ;
 wire \Tile_X6Y2_NN4BEG[4] ;
 wire \Tile_X6Y2_NN4BEG[5] ;
 wire \Tile_X6Y2_NN4BEG[6] ;
 wire \Tile_X6Y2_NN4BEG[7] ;
 wire \Tile_X6Y2_NN4BEG[8] ;
 wire \Tile_X6Y2_NN4BEG[9] ;
 wire \Tile_X6Y2_S1BEG[0] ;
 wire \Tile_X6Y2_S1BEG[1] ;
 wire \Tile_X6Y2_S1BEG[2] ;
 wire \Tile_X6Y2_S1BEG[3] ;
 wire \Tile_X6Y2_S2BEG[0] ;
 wire \Tile_X6Y2_S2BEG[1] ;
 wire \Tile_X6Y2_S2BEG[2] ;
 wire \Tile_X6Y2_S2BEG[3] ;
 wire \Tile_X6Y2_S2BEG[4] ;
 wire \Tile_X6Y2_S2BEG[5] ;
 wire \Tile_X6Y2_S2BEG[6] ;
 wire \Tile_X6Y2_S2BEG[7] ;
 wire \Tile_X6Y2_S2BEGb[0] ;
 wire \Tile_X6Y2_S2BEGb[1] ;
 wire \Tile_X6Y2_S2BEGb[2] ;
 wire \Tile_X6Y2_S2BEGb[3] ;
 wire \Tile_X6Y2_S2BEGb[4] ;
 wire \Tile_X6Y2_S2BEGb[5] ;
 wire \Tile_X6Y2_S2BEGb[6] ;
 wire \Tile_X6Y2_S2BEGb[7] ;
 wire \Tile_X6Y2_S4BEG[0] ;
 wire \Tile_X6Y2_S4BEG[10] ;
 wire \Tile_X6Y2_S4BEG[11] ;
 wire \Tile_X6Y2_S4BEG[12] ;
 wire \Tile_X6Y2_S4BEG[13] ;
 wire \Tile_X6Y2_S4BEG[14] ;
 wire \Tile_X6Y2_S4BEG[15] ;
 wire \Tile_X6Y2_S4BEG[1] ;
 wire \Tile_X6Y2_S4BEG[2] ;
 wire \Tile_X6Y2_S4BEG[3] ;
 wire \Tile_X6Y2_S4BEG[4] ;
 wire \Tile_X6Y2_S4BEG[5] ;
 wire \Tile_X6Y2_S4BEG[6] ;
 wire \Tile_X6Y2_S4BEG[7] ;
 wire \Tile_X6Y2_S4BEG[8] ;
 wire \Tile_X6Y2_S4BEG[9] ;
 wire \Tile_X6Y2_SS4BEG[0] ;
 wire \Tile_X6Y2_SS4BEG[10] ;
 wire \Tile_X6Y2_SS4BEG[11] ;
 wire \Tile_X6Y2_SS4BEG[12] ;
 wire \Tile_X6Y2_SS4BEG[13] ;
 wire \Tile_X6Y2_SS4BEG[14] ;
 wire \Tile_X6Y2_SS4BEG[15] ;
 wire \Tile_X6Y2_SS4BEG[1] ;
 wire \Tile_X6Y2_SS4BEG[2] ;
 wire \Tile_X6Y2_SS4BEG[3] ;
 wire \Tile_X6Y2_SS4BEG[4] ;
 wire \Tile_X6Y2_SS4BEG[5] ;
 wire \Tile_X6Y2_SS4BEG[6] ;
 wire \Tile_X6Y2_SS4BEG[7] ;
 wire \Tile_X6Y2_SS4BEG[8] ;
 wire \Tile_X6Y2_SS4BEG[9] ;
 wire Tile_X6Y2_UserCLKo;
 wire \Tile_X6Y2_W1BEG[0] ;
 wire \Tile_X6Y2_W1BEG[1] ;
 wire \Tile_X6Y2_W1BEG[2] ;
 wire \Tile_X6Y2_W1BEG[3] ;
 wire \Tile_X6Y2_W2BEG[0] ;
 wire \Tile_X6Y2_W2BEG[1] ;
 wire \Tile_X6Y2_W2BEG[2] ;
 wire \Tile_X6Y2_W2BEG[3] ;
 wire \Tile_X6Y2_W2BEG[4] ;
 wire \Tile_X6Y2_W2BEG[5] ;
 wire \Tile_X6Y2_W2BEG[6] ;
 wire \Tile_X6Y2_W2BEG[7] ;
 wire \Tile_X6Y2_W2BEGb[0] ;
 wire \Tile_X6Y2_W2BEGb[1] ;
 wire \Tile_X6Y2_W2BEGb[2] ;
 wire \Tile_X6Y2_W2BEGb[3] ;
 wire \Tile_X6Y2_W2BEGb[4] ;
 wire \Tile_X6Y2_W2BEGb[5] ;
 wire \Tile_X6Y2_W2BEGb[6] ;
 wire \Tile_X6Y2_W2BEGb[7] ;
 wire \Tile_X6Y2_W6BEG[0] ;
 wire \Tile_X6Y2_W6BEG[10] ;
 wire \Tile_X6Y2_W6BEG[11] ;
 wire \Tile_X6Y2_W6BEG[1] ;
 wire \Tile_X6Y2_W6BEG[2] ;
 wire \Tile_X6Y2_W6BEG[3] ;
 wire \Tile_X6Y2_W6BEG[4] ;
 wire \Tile_X6Y2_W6BEG[5] ;
 wire \Tile_X6Y2_W6BEG[6] ;
 wire \Tile_X6Y2_W6BEG[7] ;
 wire \Tile_X6Y2_W6BEG[8] ;
 wire \Tile_X6Y2_W6BEG[9] ;
 wire \Tile_X6Y2_WW4BEG[0] ;
 wire \Tile_X6Y2_WW4BEG[10] ;
 wire \Tile_X6Y2_WW4BEG[11] ;
 wire \Tile_X6Y2_WW4BEG[12] ;
 wire \Tile_X6Y2_WW4BEG[13] ;
 wire \Tile_X6Y2_WW4BEG[14] ;
 wire \Tile_X6Y2_WW4BEG[15] ;
 wire \Tile_X6Y2_WW4BEG[1] ;
 wire \Tile_X6Y2_WW4BEG[2] ;
 wire \Tile_X6Y2_WW4BEG[3] ;
 wire \Tile_X6Y2_WW4BEG[4] ;
 wire \Tile_X6Y2_WW4BEG[5] ;
 wire \Tile_X6Y2_WW4BEG[6] ;
 wire \Tile_X6Y2_WW4BEG[7] ;
 wire \Tile_X6Y2_WW4BEG[8] ;
 wire \Tile_X6Y2_WW4BEG[9] ;
 wire Tile_X6Y3_Co;
 wire \Tile_X6Y3_E1BEG[0] ;
 wire \Tile_X6Y3_E1BEG[1] ;
 wire \Tile_X6Y3_E1BEG[2] ;
 wire \Tile_X6Y3_E1BEG[3] ;
 wire \Tile_X6Y3_E2BEG[0] ;
 wire \Tile_X6Y3_E2BEG[1] ;
 wire \Tile_X6Y3_E2BEG[2] ;
 wire \Tile_X6Y3_E2BEG[3] ;
 wire \Tile_X6Y3_E2BEG[4] ;
 wire \Tile_X6Y3_E2BEG[5] ;
 wire \Tile_X6Y3_E2BEG[6] ;
 wire \Tile_X6Y3_E2BEG[7] ;
 wire \Tile_X6Y3_E2BEGb[0] ;
 wire \Tile_X6Y3_E2BEGb[1] ;
 wire \Tile_X6Y3_E2BEGb[2] ;
 wire \Tile_X6Y3_E2BEGb[3] ;
 wire \Tile_X6Y3_E2BEGb[4] ;
 wire \Tile_X6Y3_E2BEGb[5] ;
 wire \Tile_X6Y3_E2BEGb[6] ;
 wire \Tile_X6Y3_E2BEGb[7] ;
 wire \Tile_X6Y3_E6BEG[0] ;
 wire \Tile_X6Y3_E6BEG[10] ;
 wire \Tile_X6Y3_E6BEG[11] ;
 wire \Tile_X6Y3_E6BEG[1] ;
 wire \Tile_X6Y3_E6BEG[2] ;
 wire \Tile_X6Y3_E6BEG[3] ;
 wire \Tile_X6Y3_E6BEG[4] ;
 wire \Tile_X6Y3_E6BEG[5] ;
 wire \Tile_X6Y3_E6BEG[6] ;
 wire \Tile_X6Y3_E6BEG[7] ;
 wire \Tile_X6Y3_E6BEG[8] ;
 wire \Tile_X6Y3_E6BEG[9] ;
 wire \Tile_X6Y3_EE4BEG[0] ;
 wire \Tile_X6Y3_EE4BEG[10] ;
 wire \Tile_X6Y3_EE4BEG[11] ;
 wire \Tile_X6Y3_EE4BEG[12] ;
 wire \Tile_X6Y3_EE4BEG[13] ;
 wire \Tile_X6Y3_EE4BEG[14] ;
 wire \Tile_X6Y3_EE4BEG[15] ;
 wire \Tile_X6Y3_EE4BEG[1] ;
 wire \Tile_X6Y3_EE4BEG[2] ;
 wire \Tile_X6Y3_EE4BEG[3] ;
 wire \Tile_X6Y3_EE4BEG[4] ;
 wire \Tile_X6Y3_EE4BEG[5] ;
 wire \Tile_X6Y3_EE4BEG[6] ;
 wire \Tile_X6Y3_EE4BEG[7] ;
 wire \Tile_X6Y3_EE4BEG[8] ;
 wire \Tile_X6Y3_EE4BEG[9] ;
 wire \Tile_X6Y3_FrameData_O[0] ;
 wire \Tile_X6Y3_FrameData_O[10] ;
 wire \Tile_X6Y3_FrameData_O[11] ;
 wire \Tile_X6Y3_FrameData_O[12] ;
 wire \Tile_X6Y3_FrameData_O[13] ;
 wire \Tile_X6Y3_FrameData_O[14] ;
 wire \Tile_X6Y3_FrameData_O[15] ;
 wire \Tile_X6Y3_FrameData_O[16] ;
 wire \Tile_X6Y3_FrameData_O[17] ;
 wire \Tile_X6Y3_FrameData_O[18] ;
 wire \Tile_X6Y3_FrameData_O[19] ;
 wire \Tile_X6Y3_FrameData_O[1] ;
 wire \Tile_X6Y3_FrameData_O[20] ;
 wire \Tile_X6Y3_FrameData_O[21] ;
 wire \Tile_X6Y3_FrameData_O[22] ;
 wire \Tile_X6Y3_FrameData_O[23] ;
 wire \Tile_X6Y3_FrameData_O[24] ;
 wire \Tile_X6Y3_FrameData_O[25] ;
 wire \Tile_X6Y3_FrameData_O[26] ;
 wire \Tile_X6Y3_FrameData_O[27] ;
 wire \Tile_X6Y3_FrameData_O[28] ;
 wire \Tile_X6Y3_FrameData_O[29] ;
 wire \Tile_X6Y3_FrameData_O[2] ;
 wire \Tile_X6Y3_FrameData_O[30] ;
 wire \Tile_X6Y3_FrameData_O[31] ;
 wire \Tile_X6Y3_FrameData_O[3] ;
 wire \Tile_X6Y3_FrameData_O[4] ;
 wire \Tile_X6Y3_FrameData_O[5] ;
 wire \Tile_X6Y3_FrameData_O[6] ;
 wire \Tile_X6Y3_FrameData_O[7] ;
 wire \Tile_X6Y3_FrameData_O[8] ;
 wire \Tile_X6Y3_FrameData_O[9] ;
 wire \Tile_X6Y3_FrameStrobe_O[0] ;
 wire \Tile_X6Y3_FrameStrobe_O[10] ;
 wire \Tile_X6Y3_FrameStrobe_O[11] ;
 wire \Tile_X6Y3_FrameStrobe_O[12] ;
 wire \Tile_X6Y3_FrameStrobe_O[13] ;
 wire \Tile_X6Y3_FrameStrobe_O[14] ;
 wire \Tile_X6Y3_FrameStrobe_O[15] ;
 wire \Tile_X6Y3_FrameStrobe_O[16] ;
 wire \Tile_X6Y3_FrameStrobe_O[17] ;
 wire \Tile_X6Y3_FrameStrobe_O[18] ;
 wire \Tile_X6Y3_FrameStrobe_O[19] ;
 wire \Tile_X6Y3_FrameStrobe_O[1] ;
 wire \Tile_X6Y3_FrameStrobe_O[2] ;
 wire \Tile_X6Y3_FrameStrobe_O[3] ;
 wire \Tile_X6Y3_FrameStrobe_O[4] ;
 wire \Tile_X6Y3_FrameStrobe_O[5] ;
 wire \Tile_X6Y3_FrameStrobe_O[6] ;
 wire \Tile_X6Y3_FrameStrobe_O[7] ;
 wire \Tile_X6Y3_FrameStrobe_O[8] ;
 wire \Tile_X6Y3_FrameStrobe_O[9] ;
 wire \Tile_X6Y3_N1BEG[0] ;
 wire \Tile_X6Y3_N1BEG[1] ;
 wire \Tile_X6Y3_N1BEG[2] ;
 wire \Tile_X6Y3_N1BEG[3] ;
 wire \Tile_X6Y3_N2BEG[0] ;
 wire \Tile_X6Y3_N2BEG[1] ;
 wire \Tile_X6Y3_N2BEG[2] ;
 wire \Tile_X6Y3_N2BEG[3] ;
 wire \Tile_X6Y3_N2BEG[4] ;
 wire \Tile_X6Y3_N2BEG[5] ;
 wire \Tile_X6Y3_N2BEG[6] ;
 wire \Tile_X6Y3_N2BEG[7] ;
 wire \Tile_X6Y3_N2BEGb[0] ;
 wire \Tile_X6Y3_N2BEGb[1] ;
 wire \Tile_X6Y3_N2BEGb[2] ;
 wire \Tile_X6Y3_N2BEGb[3] ;
 wire \Tile_X6Y3_N2BEGb[4] ;
 wire \Tile_X6Y3_N2BEGb[5] ;
 wire \Tile_X6Y3_N2BEGb[6] ;
 wire \Tile_X6Y3_N2BEGb[7] ;
 wire \Tile_X6Y3_N4BEG[0] ;
 wire \Tile_X6Y3_N4BEG[10] ;
 wire \Tile_X6Y3_N4BEG[11] ;
 wire \Tile_X6Y3_N4BEG[12] ;
 wire \Tile_X6Y3_N4BEG[13] ;
 wire \Tile_X6Y3_N4BEG[14] ;
 wire \Tile_X6Y3_N4BEG[15] ;
 wire \Tile_X6Y3_N4BEG[1] ;
 wire \Tile_X6Y3_N4BEG[2] ;
 wire \Tile_X6Y3_N4BEG[3] ;
 wire \Tile_X6Y3_N4BEG[4] ;
 wire \Tile_X6Y3_N4BEG[5] ;
 wire \Tile_X6Y3_N4BEG[6] ;
 wire \Tile_X6Y3_N4BEG[7] ;
 wire \Tile_X6Y3_N4BEG[8] ;
 wire \Tile_X6Y3_N4BEG[9] ;
 wire \Tile_X6Y3_NN4BEG[0] ;
 wire \Tile_X6Y3_NN4BEG[10] ;
 wire \Tile_X6Y3_NN4BEG[11] ;
 wire \Tile_X6Y3_NN4BEG[12] ;
 wire \Tile_X6Y3_NN4BEG[13] ;
 wire \Tile_X6Y3_NN4BEG[14] ;
 wire \Tile_X6Y3_NN4BEG[15] ;
 wire \Tile_X6Y3_NN4BEG[1] ;
 wire \Tile_X6Y3_NN4BEG[2] ;
 wire \Tile_X6Y3_NN4BEG[3] ;
 wire \Tile_X6Y3_NN4BEG[4] ;
 wire \Tile_X6Y3_NN4BEG[5] ;
 wire \Tile_X6Y3_NN4BEG[6] ;
 wire \Tile_X6Y3_NN4BEG[7] ;
 wire \Tile_X6Y3_NN4BEG[8] ;
 wire \Tile_X6Y3_NN4BEG[9] ;
 wire \Tile_X6Y3_S1BEG[0] ;
 wire \Tile_X6Y3_S1BEG[1] ;
 wire \Tile_X6Y3_S1BEG[2] ;
 wire \Tile_X6Y3_S1BEG[3] ;
 wire \Tile_X6Y3_S2BEG[0] ;
 wire \Tile_X6Y3_S2BEG[1] ;
 wire \Tile_X6Y3_S2BEG[2] ;
 wire \Tile_X6Y3_S2BEG[3] ;
 wire \Tile_X6Y3_S2BEG[4] ;
 wire \Tile_X6Y3_S2BEG[5] ;
 wire \Tile_X6Y3_S2BEG[6] ;
 wire \Tile_X6Y3_S2BEG[7] ;
 wire \Tile_X6Y3_S2BEGb[0] ;
 wire \Tile_X6Y3_S2BEGb[1] ;
 wire \Tile_X6Y3_S2BEGb[2] ;
 wire \Tile_X6Y3_S2BEGb[3] ;
 wire \Tile_X6Y3_S2BEGb[4] ;
 wire \Tile_X6Y3_S2BEGb[5] ;
 wire \Tile_X6Y3_S2BEGb[6] ;
 wire \Tile_X6Y3_S2BEGb[7] ;
 wire \Tile_X6Y3_S4BEG[0] ;
 wire \Tile_X6Y3_S4BEG[10] ;
 wire \Tile_X6Y3_S4BEG[11] ;
 wire \Tile_X6Y3_S4BEG[12] ;
 wire \Tile_X6Y3_S4BEG[13] ;
 wire \Tile_X6Y3_S4BEG[14] ;
 wire \Tile_X6Y3_S4BEG[15] ;
 wire \Tile_X6Y3_S4BEG[1] ;
 wire \Tile_X6Y3_S4BEG[2] ;
 wire \Tile_X6Y3_S4BEG[3] ;
 wire \Tile_X6Y3_S4BEG[4] ;
 wire \Tile_X6Y3_S4BEG[5] ;
 wire \Tile_X6Y3_S4BEG[6] ;
 wire \Tile_X6Y3_S4BEG[7] ;
 wire \Tile_X6Y3_S4BEG[8] ;
 wire \Tile_X6Y3_S4BEG[9] ;
 wire \Tile_X6Y3_SS4BEG[0] ;
 wire \Tile_X6Y3_SS4BEG[10] ;
 wire \Tile_X6Y3_SS4BEG[11] ;
 wire \Tile_X6Y3_SS4BEG[12] ;
 wire \Tile_X6Y3_SS4BEG[13] ;
 wire \Tile_X6Y3_SS4BEG[14] ;
 wire \Tile_X6Y3_SS4BEG[15] ;
 wire \Tile_X6Y3_SS4BEG[1] ;
 wire \Tile_X6Y3_SS4BEG[2] ;
 wire \Tile_X6Y3_SS4BEG[3] ;
 wire \Tile_X6Y3_SS4BEG[4] ;
 wire \Tile_X6Y3_SS4BEG[5] ;
 wire \Tile_X6Y3_SS4BEG[6] ;
 wire \Tile_X6Y3_SS4BEG[7] ;
 wire \Tile_X6Y3_SS4BEG[8] ;
 wire \Tile_X6Y3_SS4BEG[9] ;
 wire Tile_X6Y3_UserCLKo;
 wire \Tile_X6Y3_W1BEG[0] ;
 wire \Tile_X6Y3_W1BEG[1] ;
 wire \Tile_X6Y3_W1BEG[2] ;
 wire \Tile_X6Y3_W1BEG[3] ;
 wire \Tile_X6Y3_W2BEG[0] ;
 wire \Tile_X6Y3_W2BEG[1] ;
 wire \Tile_X6Y3_W2BEG[2] ;
 wire \Tile_X6Y3_W2BEG[3] ;
 wire \Tile_X6Y3_W2BEG[4] ;
 wire \Tile_X6Y3_W2BEG[5] ;
 wire \Tile_X6Y3_W2BEG[6] ;
 wire \Tile_X6Y3_W2BEG[7] ;
 wire \Tile_X6Y3_W2BEGb[0] ;
 wire \Tile_X6Y3_W2BEGb[1] ;
 wire \Tile_X6Y3_W2BEGb[2] ;
 wire \Tile_X6Y3_W2BEGb[3] ;
 wire \Tile_X6Y3_W2BEGb[4] ;
 wire \Tile_X6Y3_W2BEGb[5] ;
 wire \Tile_X6Y3_W2BEGb[6] ;
 wire \Tile_X6Y3_W2BEGb[7] ;
 wire \Tile_X6Y3_W6BEG[0] ;
 wire \Tile_X6Y3_W6BEG[10] ;
 wire \Tile_X6Y3_W6BEG[11] ;
 wire \Tile_X6Y3_W6BEG[1] ;
 wire \Tile_X6Y3_W6BEG[2] ;
 wire \Tile_X6Y3_W6BEG[3] ;
 wire \Tile_X6Y3_W6BEG[4] ;
 wire \Tile_X6Y3_W6BEG[5] ;
 wire \Tile_X6Y3_W6BEG[6] ;
 wire \Tile_X6Y3_W6BEG[7] ;
 wire \Tile_X6Y3_W6BEG[8] ;
 wire \Tile_X6Y3_W6BEG[9] ;
 wire \Tile_X6Y3_WW4BEG[0] ;
 wire \Tile_X6Y3_WW4BEG[10] ;
 wire \Tile_X6Y3_WW4BEG[11] ;
 wire \Tile_X6Y3_WW4BEG[12] ;
 wire \Tile_X6Y3_WW4BEG[13] ;
 wire \Tile_X6Y3_WW4BEG[14] ;
 wire \Tile_X6Y3_WW4BEG[15] ;
 wire \Tile_X6Y3_WW4BEG[1] ;
 wire \Tile_X6Y3_WW4BEG[2] ;
 wire \Tile_X6Y3_WW4BEG[3] ;
 wire \Tile_X6Y3_WW4BEG[4] ;
 wire \Tile_X6Y3_WW4BEG[5] ;
 wire \Tile_X6Y3_WW4BEG[6] ;
 wire \Tile_X6Y3_WW4BEG[7] ;
 wire \Tile_X6Y3_WW4BEG[8] ;
 wire \Tile_X6Y3_WW4BEG[9] ;
 wire Tile_X6Y4_Co;
 wire \Tile_X6Y4_E1BEG[0] ;
 wire \Tile_X6Y4_E1BEG[1] ;
 wire \Tile_X6Y4_E1BEG[2] ;
 wire \Tile_X6Y4_E1BEG[3] ;
 wire \Tile_X6Y4_E2BEG[0] ;
 wire \Tile_X6Y4_E2BEG[1] ;
 wire \Tile_X6Y4_E2BEG[2] ;
 wire \Tile_X6Y4_E2BEG[3] ;
 wire \Tile_X6Y4_E2BEG[4] ;
 wire \Tile_X6Y4_E2BEG[5] ;
 wire \Tile_X6Y4_E2BEG[6] ;
 wire \Tile_X6Y4_E2BEG[7] ;
 wire \Tile_X6Y4_E2BEGb[0] ;
 wire \Tile_X6Y4_E2BEGb[1] ;
 wire \Tile_X6Y4_E2BEGb[2] ;
 wire \Tile_X6Y4_E2BEGb[3] ;
 wire \Tile_X6Y4_E2BEGb[4] ;
 wire \Tile_X6Y4_E2BEGb[5] ;
 wire \Tile_X6Y4_E2BEGb[6] ;
 wire \Tile_X6Y4_E2BEGb[7] ;
 wire \Tile_X6Y4_E6BEG[0] ;
 wire \Tile_X6Y4_E6BEG[10] ;
 wire \Tile_X6Y4_E6BEG[11] ;
 wire \Tile_X6Y4_E6BEG[1] ;
 wire \Tile_X6Y4_E6BEG[2] ;
 wire \Tile_X6Y4_E6BEG[3] ;
 wire \Tile_X6Y4_E6BEG[4] ;
 wire \Tile_X6Y4_E6BEG[5] ;
 wire \Tile_X6Y4_E6BEG[6] ;
 wire \Tile_X6Y4_E6BEG[7] ;
 wire \Tile_X6Y4_E6BEG[8] ;
 wire \Tile_X6Y4_E6BEG[9] ;
 wire \Tile_X6Y4_EE4BEG[0] ;
 wire \Tile_X6Y4_EE4BEG[10] ;
 wire \Tile_X6Y4_EE4BEG[11] ;
 wire \Tile_X6Y4_EE4BEG[12] ;
 wire \Tile_X6Y4_EE4BEG[13] ;
 wire \Tile_X6Y4_EE4BEG[14] ;
 wire \Tile_X6Y4_EE4BEG[15] ;
 wire \Tile_X6Y4_EE4BEG[1] ;
 wire \Tile_X6Y4_EE4BEG[2] ;
 wire \Tile_X6Y4_EE4BEG[3] ;
 wire \Tile_X6Y4_EE4BEG[4] ;
 wire \Tile_X6Y4_EE4BEG[5] ;
 wire \Tile_X6Y4_EE4BEG[6] ;
 wire \Tile_X6Y4_EE4BEG[7] ;
 wire \Tile_X6Y4_EE4BEG[8] ;
 wire \Tile_X6Y4_EE4BEG[9] ;
 wire \Tile_X6Y4_FrameData_O[0] ;
 wire \Tile_X6Y4_FrameData_O[10] ;
 wire \Tile_X6Y4_FrameData_O[11] ;
 wire \Tile_X6Y4_FrameData_O[12] ;
 wire \Tile_X6Y4_FrameData_O[13] ;
 wire \Tile_X6Y4_FrameData_O[14] ;
 wire \Tile_X6Y4_FrameData_O[15] ;
 wire \Tile_X6Y4_FrameData_O[16] ;
 wire \Tile_X6Y4_FrameData_O[17] ;
 wire \Tile_X6Y4_FrameData_O[18] ;
 wire \Tile_X6Y4_FrameData_O[19] ;
 wire \Tile_X6Y4_FrameData_O[1] ;
 wire \Tile_X6Y4_FrameData_O[20] ;
 wire \Tile_X6Y4_FrameData_O[21] ;
 wire \Tile_X6Y4_FrameData_O[22] ;
 wire \Tile_X6Y4_FrameData_O[23] ;
 wire \Tile_X6Y4_FrameData_O[24] ;
 wire \Tile_X6Y4_FrameData_O[25] ;
 wire \Tile_X6Y4_FrameData_O[26] ;
 wire \Tile_X6Y4_FrameData_O[27] ;
 wire \Tile_X6Y4_FrameData_O[28] ;
 wire \Tile_X6Y4_FrameData_O[29] ;
 wire \Tile_X6Y4_FrameData_O[2] ;
 wire \Tile_X6Y4_FrameData_O[30] ;
 wire \Tile_X6Y4_FrameData_O[31] ;
 wire \Tile_X6Y4_FrameData_O[3] ;
 wire \Tile_X6Y4_FrameData_O[4] ;
 wire \Tile_X6Y4_FrameData_O[5] ;
 wire \Tile_X6Y4_FrameData_O[6] ;
 wire \Tile_X6Y4_FrameData_O[7] ;
 wire \Tile_X6Y4_FrameData_O[8] ;
 wire \Tile_X6Y4_FrameData_O[9] ;
 wire \Tile_X6Y4_FrameStrobe_O[0] ;
 wire \Tile_X6Y4_FrameStrobe_O[10] ;
 wire \Tile_X6Y4_FrameStrobe_O[11] ;
 wire \Tile_X6Y4_FrameStrobe_O[12] ;
 wire \Tile_X6Y4_FrameStrobe_O[13] ;
 wire \Tile_X6Y4_FrameStrobe_O[14] ;
 wire \Tile_X6Y4_FrameStrobe_O[15] ;
 wire \Tile_X6Y4_FrameStrobe_O[16] ;
 wire \Tile_X6Y4_FrameStrobe_O[17] ;
 wire \Tile_X6Y4_FrameStrobe_O[18] ;
 wire \Tile_X6Y4_FrameStrobe_O[19] ;
 wire \Tile_X6Y4_FrameStrobe_O[1] ;
 wire \Tile_X6Y4_FrameStrobe_O[2] ;
 wire \Tile_X6Y4_FrameStrobe_O[3] ;
 wire \Tile_X6Y4_FrameStrobe_O[4] ;
 wire \Tile_X6Y4_FrameStrobe_O[5] ;
 wire \Tile_X6Y4_FrameStrobe_O[6] ;
 wire \Tile_X6Y4_FrameStrobe_O[7] ;
 wire \Tile_X6Y4_FrameStrobe_O[8] ;
 wire \Tile_X6Y4_FrameStrobe_O[9] ;
 wire \Tile_X6Y4_N1BEG[0] ;
 wire \Tile_X6Y4_N1BEG[1] ;
 wire \Tile_X6Y4_N1BEG[2] ;
 wire \Tile_X6Y4_N1BEG[3] ;
 wire \Tile_X6Y4_N2BEG[0] ;
 wire \Tile_X6Y4_N2BEG[1] ;
 wire \Tile_X6Y4_N2BEG[2] ;
 wire \Tile_X6Y4_N2BEG[3] ;
 wire \Tile_X6Y4_N2BEG[4] ;
 wire \Tile_X6Y4_N2BEG[5] ;
 wire \Tile_X6Y4_N2BEG[6] ;
 wire \Tile_X6Y4_N2BEG[7] ;
 wire \Tile_X6Y4_N2BEGb[0] ;
 wire \Tile_X6Y4_N2BEGb[1] ;
 wire \Tile_X6Y4_N2BEGb[2] ;
 wire \Tile_X6Y4_N2BEGb[3] ;
 wire \Tile_X6Y4_N2BEGb[4] ;
 wire \Tile_X6Y4_N2BEGb[5] ;
 wire \Tile_X6Y4_N2BEGb[6] ;
 wire \Tile_X6Y4_N2BEGb[7] ;
 wire \Tile_X6Y4_N4BEG[0] ;
 wire \Tile_X6Y4_N4BEG[10] ;
 wire \Tile_X6Y4_N4BEG[11] ;
 wire \Tile_X6Y4_N4BEG[12] ;
 wire \Tile_X6Y4_N4BEG[13] ;
 wire \Tile_X6Y4_N4BEG[14] ;
 wire \Tile_X6Y4_N4BEG[15] ;
 wire \Tile_X6Y4_N4BEG[1] ;
 wire \Tile_X6Y4_N4BEG[2] ;
 wire \Tile_X6Y4_N4BEG[3] ;
 wire \Tile_X6Y4_N4BEG[4] ;
 wire \Tile_X6Y4_N4BEG[5] ;
 wire \Tile_X6Y4_N4BEG[6] ;
 wire \Tile_X6Y4_N4BEG[7] ;
 wire \Tile_X6Y4_N4BEG[8] ;
 wire \Tile_X6Y4_N4BEG[9] ;
 wire \Tile_X6Y4_NN4BEG[0] ;
 wire \Tile_X6Y4_NN4BEG[10] ;
 wire \Tile_X6Y4_NN4BEG[11] ;
 wire \Tile_X6Y4_NN4BEG[12] ;
 wire \Tile_X6Y4_NN4BEG[13] ;
 wire \Tile_X6Y4_NN4BEG[14] ;
 wire \Tile_X6Y4_NN4BEG[15] ;
 wire \Tile_X6Y4_NN4BEG[1] ;
 wire \Tile_X6Y4_NN4BEG[2] ;
 wire \Tile_X6Y4_NN4BEG[3] ;
 wire \Tile_X6Y4_NN4BEG[4] ;
 wire \Tile_X6Y4_NN4BEG[5] ;
 wire \Tile_X6Y4_NN4BEG[6] ;
 wire \Tile_X6Y4_NN4BEG[7] ;
 wire \Tile_X6Y4_NN4BEG[8] ;
 wire \Tile_X6Y4_NN4BEG[9] ;
 wire \Tile_X6Y4_S1BEG[0] ;
 wire \Tile_X6Y4_S1BEG[1] ;
 wire \Tile_X6Y4_S1BEG[2] ;
 wire \Tile_X6Y4_S1BEG[3] ;
 wire \Tile_X6Y4_S2BEG[0] ;
 wire \Tile_X6Y4_S2BEG[1] ;
 wire \Tile_X6Y4_S2BEG[2] ;
 wire \Tile_X6Y4_S2BEG[3] ;
 wire \Tile_X6Y4_S2BEG[4] ;
 wire \Tile_X6Y4_S2BEG[5] ;
 wire \Tile_X6Y4_S2BEG[6] ;
 wire \Tile_X6Y4_S2BEG[7] ;
 wire \Tile_X6Y4_S2BEGb[0] ;
 wire \Tile_X6Y4_S2BEGb[1] ;
 wire \Tile_X6Y4_S2BEGb[2] ;
 wire \Tile_X6Y4_S2BEGb[3] ;
 wire \Tile_X6Y4_S2BEGb[4] ;
 wire \Tile_X6Y4_S2BEGb[5] ;
 wire \Tile_X6Y4_S2BEGb[6] ;
 wire \Tile_X6Y4_S2BEGb[7] ;
 wire \Tile_X6Y4_S4BEG[0] ;
 wire \Tile_X6Y4_S4BEG[10] ;
 wire \Tile_X6Y4_S4BEG[11] ;
 wire \Tile_X6Y4_S4BEG[12] ;
 wire \Tile_X6Y4_S4BEG[13] ;
 wire \Tile_X6Y4_S4BEG[14] ;
 wire \Tile_X6Y4_S4BEG[15] ;
 wire \Tile_X6Y4_S4BEG[1] ;
 wire \Tile_X6Y4_S4BEG[2] ;
 wire \Tile_X6Y4_S4BEG[3] ;
 wire \Tile_X6Y4_S4BEG[4] ;
 wire \Tile_X6Y4_S4BEG[5] ;
 wire \Tile_X6Y4_S4BEG[6] ;
 wire \Tile_X6Y4_S4BEG[7] ;
 wire \Tile_X6Y4_S4BEG[8] ;
 wire \Tile_X6Y4_S4BEG[9] ;
 wire \Tile_X6Y4_SS4BEG[0] ;
 wire \Tile_X6Y4_SS4BEG[10] ;
 wire \Tile_X6Y4_SS4BEG[11] ;
 wire \Tile_X6Y4_SS4BEG[12] ;
 wire \Tile_X6Y4_SS4BEG[13] ;
 wire \Tile_X6Y4_SS4BEG[14] ;
 wire \Tile_X6Y4_SS4BEG[15] ;
 wire \Tile_X6Y4_SS4BEG[1] ;
 wire \Tile_X6Y4_SS4BEG[2] ;
 wire \Tile_X6Y4_SS4BEG[3] ;
 wire \Tile_X6Y4_SS4BEG[4] ;
 wire \Tile_X6Y4_SS4BEG[5] ;
 wire \Tile_X6Y4_SS4BEG[6] ;
 wire \Tile_X6Y4_SS4BEG[7] ;
 wire \Tile_X6Y4_SS4BEG[8] ;
 wire \Tile_X6Y4_SS4BEG[9] ;
 wire Tile_X6Y4_UserCLKo;
 wire \Tile_X6Y4_W1BEG[0] ;
 wire \Tile_X6Y4_W1BEG[1] ;
 wire \Tile_X6Y4_W1BEG[2] ;
 wire \Tile_X6Y4_W1BEG[3] ;
 wire \Tile_X6Y4_W2BEG[0] ;
 wire \Tile_X6Y4_W2BEG[1] ;
 wire \Tile_X6Y4_W2BEG[2] ;
 wire \Tile_X6Y4_W2BEG[3] ;
 wire \Tile_X6Y4_W2BEG[4] ;
 wire \Tile_X6Y4_W2BEG[5] ;
 wire \Tile_X6Y4_W2BEG[6] ;
 wire \Tile_X6Y4_W2BEG[7] ;
 wire \Tile_X6Y4_W2BEGb[0] ;
 wire \Tile_X6Y4_W2BEGb[1] ;
 wire \Tile_X6Y4_W2BEGb[2] ;
 wire \Tile_X6Y4_W2BEGb[3] ;
 wire \Tile_X6Y4_W2BEGb[4] ;
 wire \Tile_X6Y4_W2BEGb[5] ;
 wire \Tile_X6Y4_W2BEGb[6] ;
 wire \Tile_X6Y4_W2BEGb[7] ;
 wire \Tile_X6Y4_W6BEG[0] ;
 wire \Tile_X6Y4_W6BEG[10] ;
 wire \Tile_X6Y4_W6BEG[11] ;
 wire \Tile_X6Y4_W6BEG[1] ;
 wire \Tile_X6Y4_W6BEG[2] ;
 wire \Tile_X6Y4_W6BEG[3] ;
 wire \Tile_X6Y4_W6BEG[4] ;
 wire \Tile_X6Y4_W6BEG[5] ;
 wire \Tile_X6Y4_W6BEG[6] ;
 wire \Tile_X6Y4_W6BEG[7] ;
 wire \Tile_X6Y4_W6BEG[8] ;
 wire \Tile_X6Y4_W6BEG[9] ;
 wire \Tile_X6Y4_WW4BEG[0] ;
 wire \Tile_X6Y4_WW4BEG[10] ;
 wire \Tile_X6Y4_WW4BEG[11] ;
 wire \Tile_X6Y4_WW4BEG[12] ;
 wire \Tile_X6Y4_WW4BEG[13] ;
 wire \Tile_X6Y4_WW4BEG[14] ;
 wire \Tile_X6Y4_WW4BEG[15] ;
 wire \Tile_X6Y4_WW4BEG[1] ;
 wire \Tile_X6Y4_WW4BEG[2] ;
 wire \Tile_X6Y4_WW4BEG[3] ;
 wire \Tile_X6Y4_WW4BEG[4] ;
 wire \Tile_X6Y4_WW4BEG[5] ;
 wire \Tile_X6Y4_WW4BEG[6] ;
 wire \Tile_X6Y4_WW4BEG[7] ;
 wire \Tile_X6Y4_WW4BEG[8] ;
 wire \Tile_X6Y4_WW4BEG[9] ;
 wire Tile_X6Y5_Co;
 wire \Tile_X6Y5_E1BEG[0] ;
 wire \Tile_X6Y5_E1BEG[1] ;
 wire \Tile_X6Y5_E1BEG[2] ;
 wire \Tile_X6Y5_E1BEG[3] ;
 wire \Tile_X6Y5_E2BEG[0] ;
 wire \Tile_X6Y5_E2BEG[1] ;
 wire \Tile_X6Y5_E2BEG[2] ;
 wire \Tile_X6Y5_E2BEG[3] ;
 wire \Tile_X6Y5_E2BEG[4] ;
 wire \Tile_X6Y5_E2BEG[5] ;
 wire \Tile_X6Y5_E2BEG[6] ;
 wire \Tile_X6Y5_E2BEG[7] ;
 wire \Tile_X6Y5_E2BEGb[0] ;
 wire \Tile_X6Y5_E2BEGb[1] ;
 wire \Tile_X6Y5_E2BEGb[2] ;
 wire \Tile_X6Y5_E2BEGb[3] ;
 wire \Tile_X6Y5_E2BEGb[4] ;
 wire \Tile_X6Y5_E2BEGb[5] ;
 wire \Tile_X6Y5_E2BEGb[6] ;
 wire \Tile_X6Y5_E2BEGb[7] ;
 wire \Tile_X6Y5_E6BEG[0] ;
 wire \Tile_X6Y5_E6BEG[10] ;
 wire \Tile_X6Y5_E6BEG[11] ;
 wire \Tile_X6Y5_E6BEG[1] ;
 wire \Tile_X6Y5_E6BEG[2] ;
 wire \Tile_X6Y5_E6BEG[3] ;
 wire \Tile_X6Y5_E6BEG[4] ;
 wire \Tile_X6Y5_E6BEG[5] ;
 wire \Tile_X6Y5_E6BEG[6] ;
 wire \Tile_X6Y5_E6BEG[7] ;
 wire \Tile_X6Y5_E6BEG[8] ;
 wire \Tile_X6Y5_E6BEG[9] ;
 wire \Tile_X6Y5_EE4BEG[0] ;
 wire \Tile_X6Y5_EE4BEG[10] ;
 wire \Tile_X6Y5_EE4BEG[11] ;
 wire \Tile_X6Y5_EE4BEG[12] ;
 wire \Tile_X6Y5_EE4BEG[13] ;
 wire \Tile_X6Y5_EE4BEG[14] ;
 wire \Tile_X6Y5_EE4BEG[15] ;
 wire \Tile_X6Y5_EE4BEG[1] ;
 wire \Tile_X6Y5_EE4BEG[2] ;
 wire \Tile_X6Y5_EE4BEG[3] ;
 wire \Tile_X6Y5_EE4BEG[4] ;
 wire \Tile_X6Y5_EE4BEG[5] ;
 wire \Tile_X6Y5_EE4BEG[6] ;
 wire \Tile_X6Y5_EE4BEG[7] ;
 wire \Tile_X6Y5_EE4BEG[8] ;
 wire \Tile_X6Y5_EE4BEG[9] ;
 wire \Tile_X6Y5_FrameData_O[0] ;
 wire \Tile_X6Y5_FrameData_O[10] ;
 wire \Tile_X6Y5_FrameData_O[11] ;
 wire \Tile_X6Y5_FrameData_O[12] ;
 wire \Tile_X6Y5_FrameData_O[13] ;
 wire \Tile_X6Y5_FrameData_O[14] ;
 wire \Tile_X6Y5_FrameData_O[15] ;
 wire \Tile_X6Y5_FrameData_O[16] ;
 wire \Tile_X6Y5_FrameData_O[17] ;
 wire \Tile_X6Y5_FrameData_O[18] ;
 wire \Tile_X6Y5_FrameData_O[19] ;
 wire \Tile_X6Y5_FrameData_O[1] ;
 wire \Tile_X6Y5_FrameData_O[20] ;
 wire \Tile_X6Y5_FrameData_O[21] ;
 wire \Tile_X6Y5_FrameData_O[22] ;
 wire \Tile_X6Y5_FrameData_O[23] ;
 wire \Tile_X6Y5_FrameData_O[24] ;
 wire \Tile_X6Y5_FrameData_O[25] ;
 wire \Tile_X6Y5_FrameData_O[26] ;
 wire \Tile_X6Y5_FrameData_O[27] ;
 wire \Tile_X6Y5_FrameData_O[28] ;
 wire \Tile_X6Y5_FrameData_O[29] ;
 wire \Tile_X6Y5_FrameData_O[2] ;
 wire \Tile_X6Y5_FrameData_O[30] ;
 wire \Tile_X6Y5_FrameData_O[31] ;
 wire \Tile_X6Y5_FrameData_O[3] ;
 wire \Tile_X6Y5_FrameData_O[4] ;
 wire \Tile_X6Y5_FrameData_O[5] ;
 wire \Tile_X6Y5_FrameData_O[6] ;
 wire \Tile_X6Y5_FrameData_O[7] ;
 wire \Tile_X6Y5_FrameData_O[8] ;
 wire \Tile_X6Y5_FrameData_O[9] ;
 wire \Tile_X6Y5_FrameStrobe_O[0] ;
 wire \Tile_X6Y5_FrameStrobe_O[10] ;
 wire \Tile_X6Y5_FrameStrobe_O[11] ;
 wire \Tile_X6Y5_FrameStrobe_O[12] ;
 wire \Tile_X6Y5_FrameStrobe_O[13] ;
 wire \Tile_X6Y5_FrameStrobe_O[14] ;
 wire \Tile_X6Y5_FrameStrobe_O[15] ;
 wire \Tile_X6Y5_FrameStrobe_O[16] ;
 wire \Tile_X6Y5_FrameStrobe_O[17] ;
 wire \Tile_X6Y5_FrameStrobe_O[18] ;
 wire \Tile_X6Y5_FrameStrobe_O[19] ;
 wire \Tile_X6Y5_FrameStrobe_O[1] ;
 wire \Tile_X6Y5_FrameStrobe_O[2] ;
 wire \Tile_X6Y5_FrameStrobe_O[3] ;
 wire \Tile_X6Y5_FrameStrobe_O[4] ;
 wire \Tile_X6Y5_FrameStrobe_O[5] ;
 wire \Tile_X6Y5_FrameStrobe_O[6] ;
 wire \Tile_X6Y5_FrameStrobe_O[7] ;
 wire \Tile_X6Y5_FrameStrobe_O[8] ;
 wire \Tile_X6Y5_FrameStrobe_O[9] ;
 wire \Tile_X6Y5_N1BEG[0] ;
 wire \Tile_X6Y5_N1BEG[1] ;
 wire \Tile_X6Y5_N1BEG[2] ;
 wire \Tile_X6Y5_N1BEG[3] ;
 wire \Tile_X6Y5_N2BEG[0] ;
 wire \Tile_X6Y5_N2BEG[1] ;
 wire \Tile_X6Y5_N2BEG[2] ;
 wire \Tile_X6Y5_N2BEG[3] ;
 wire \Tile_X6Y5_N2BEG[4] ;
 wire \Tile_X6Y5_N2BEG[5] ;
 wire \Tile_X6Y5_N2BEG[6] ;
 wire \Tile_X6Y5_N2BEG[7] ;
 wire \Tile_X6Y5_N2BEGb[0] ;
 wire \Tile_X6Y5_N2BEGb[1] ;
 wire \Tile_X6Y5_N2BEGb[2] ;
 wire \Tile_X6Y5_N2BEGb[3] ;
 wire \Tile_X6Y5_N2BEGb[4] ;
 wire \Tile_X6Y5_N2BEGb[5] ;
 wire \Tile_X6Y5_N2BEGb[6] ;
 wire \Tile_X6Y5_N2BEGb[7] ;
 wire \Tile_X6Y5_N4BEG[0] ;
 wire \Tile_X6Y5_N4BEG[10] ;
 wire \Tile_X6Y5_N4BEG[11] ;
 wire \Tile_X6Y5_N4BEG[12] ;
 wire \Tile_X6Y5_N4BEG[13] ;
 wire \Tile_X6Y5_N4BEG[14] ;
 wire \Tile_X6Y5_N4BEG[15] ;
 wire \Tile_X6Y5_N4BEG[1] ;
 wire \Tile_X6Y5_N4BEG[2] ;
 wire \Tile_X6Y5_N4BEG[3] ;
 wire \Tile_X6Y5_N4BEG[4] ;
 wire \Tile_X6Y5_N4BEG[5] ;
 wire \Tile_X6Y5_N4BEG[6] ;
 wire \Tile_X6Y5_N4BEG[7] ;
 wire \Tile_X6Y5_N4BEG[8] ;
 wire \Tile_X6Y5_N4BEG[9] ;
 wire \Tile_X6Y5_NN4BEG[0] ;
 wire \Tile_X6Y5_NN4BEG[10] ;
 wire \Tile_X6Y5_NN4BEG[11] ;
 wire \Tile_X6Y5_NN4BEG[12] ;
 wire \Tile_X6Y5_NN4BEG[13] ;
 wire \Tile_X6Y5_NN4BEG[14] ;
 wire \Tile_X6Y5_NN4BEG[15] ;
 wire \Tile_X6Y5_NN4BEG[1] ;
 wire \Tile_X6Y5_NN4BEG[2] ;
 wire \Tile_X6Y5_NN4BEG[3] ;
 wire \Tile_X6Y5_NN4BEG[4] ;
 wire \Tile_X6Y5_NN4BEG[5] ;
 wire \Tile_X6Y5_NN4BEG[6] ;
 wire \Tile_X6Y5_NN4BEG[7] ;
 wire \Tile_X6Y5_NN4BEG[8] ;
 wire \Tile_X6Y5_NN4BEG[9] ;
 wire \Tile_X6Y5_S1BEG[0] ;
 wire \Tile_X6Y5_S1BEG[1] ;
 wire \Tile_X6Y5_S1BEG[2] ;
 wire \Tile_X6Y5_S1BEG[3] ;
 wire \Tile_X6Y5_S2BEG[0] ;
 wire \Tile_X6Y5_S2BEG[1] ;
 wire \Tile_X6Y5_S2BEG[2] ;
 wire \Tile_X6Y5_S2BEG[3] ;
 wire \Tile_X6Y5_S2BEG[4] ;
 wire \Tile_X6Y5_S2BEG[5] ;
 wire \Tile_X6Y5_S2BEG[6] ;
 wire \Tile_X6Y5_S2BEG[7] ;
 wire \Tile_X6Y5_S2BEGb[0] ;
 wire \Tile_X6Y5_S2BEGb[1] ;
 wire \Tile_X6Y5_S2BEGb[2] ;
 wire \Tile_X6Y5_S2BEGb[3] ;
 wire \Tile_X6Y5_S2BEGb[4] ;
 wire \Tile_X6Y5_S2BEGb[5] ;
 wire \Tile_X6Y5_S2BEGb[6] ;
 wire \Tile_X6Y5_S2BEGb[7] ;
 wire \Tile_X6Y5_S4BEG[0] ;
 wire \Tile_X6Y5_S4BEG[10] ;
 wire \Tile_X6Y5_S4BEG[11] ;
 wire \Tile_X6Y5_S4BEG[12] ;
 wire \Tile_X6Y5_S4BEG[13] ;
 wire \Tile_X6Y5_S4BEG[14] ;
 wire \Tile_X6Y5_S4BEG[15] ;
 wire \Tile_X6Y5_S4BEG[1] ;
 wire \Tile_X6Y5_S4BEG[2] ;
 wire \Tile_X6Y5_S4BEG[3] ;
 wire \Tile_X6Y5_S4BEG[4] ;
 wire \Tile_X6Y5_S4BEG[5] ;
 wire \Tile_X6Y5_S4BEG[6] ;
 wire \Tile_X6Y5_S4BEG[7] ;
 wire \Tile_X6Y5_S4BEG[8] ;
 wire \Tile_X6Y5_S4BEG[9] ;
 wire \Tile_X6Y5_SS4BEG[0] ;
 wire \Tile_X6Y5_SS4BEG[10] ;
 wire \Tile_X6Y5_SS4BEG[11] ;
 wire \Tile_X6Y5_SS4BEG[12] ;
 wire \Tile_X6Y5_SS4BEG[13] ;
 wire \Tile_X6Y5_SS4BEG[14] ;
 wire \Tile_X6Y5_SS4BEG[15] ;
 wire \Tile_X6Y5_SS4BEG[1] ;
 wire \Tile_X6Y5_SS4BEG[2] ;
 wire \Tile_X6Y5_SS4BEG[3] ;
 wire \Tile_X6Y5_SS4BEG[4] ;
 wire \Tile_X6Y5_SS4BEG[5] ;
 wire \Tile_X6Y5_SS4BEG[6] ;
 wire \Tile_X6Y5_SS4BEG[7] ;
 wire \Tile_X6Y5_SS4BEG[8] ;
 wire \Tile_X6Y5_SS4BEG[9] ;
 wire Tile_X6Y5_UserCLKo;
 wire \Tile_X6Y5_W1BEG[0] ;
 wire \Tile_X6Y5_W1BEG[1] ;
 wire \Tile_X6Y5_W1BEG[2] ;
 wire \Tile_X6Y5_W1BEG[3] ;
 wire \Tile_X6Y5_W2BEG[0] ;
 wire \Tile_X6Y5_W2BEG[1] ;
 wire \Tile_X6Y5_W2BEG[2] ;
 wire \Tile_X6Y5_W2BEG[3] ;
 wire \Tile_X6Y5_W2BEG[4] ;
 wire \Tile_X6Y5_W2BEG[5] ;
 wire \Tile_X6Y5_W2BEG[6] ;
 wire \Tile_X6Y5_W2BEG[7] ;
 wire \Tile_X6Y5_W2BEGb[0] ;
 wire \Tile_X6Y5_W2BEGb[1] ;
 wire \Tile_X6Y5_W2BEGb[2] ;
 wire \Tile_X6Y5_W2BEGb[3] ;
 wire \Tile_X6Y5_W2BEGb[4] ;
 wire \Tile_X6Y5_W2BEGb[5] ;
 wire \Tile_X6Y5_W2BEGb[6] ;
 wire \Tile_X6Y5_W2BEGb[7] ;
 wire \Tile_X6Y5_W6BEG[0] ;
 wire \Tile_X6Y5_W6BEG[10] ;
 wire \Tile_X6Y5_W6BEG[11] ;
 wire \Tile_X6Y5_W6BEG[1] ;
 wire \Tile_X6Y5_W6BEG[2] ;
 wire \Tile_X6Y5_W6BEG[3] ;
 wire \Tile_X6Y5_W6BEG[4] ;
 wire \Tile_X6Y5_W6BEG[5] ;
 wire \Tile_X6Y5_W6BEG[6] ;
 wire \Tile_X6Y5_W6BEG[7] ;
 wire \Tile_X6Y5_W6BEG[8] ;
 wire \Tile_X6Y5_W6BEG[9] ;
 wire \Tile_X6Y5_WW4BEG[0] ;
 wire \Tile_X6Y5_WW4BEG[10] ;
 wire \Tile_X6Y5_WW4BEG[11] ;
 wire \Tile_X6Y5_WW4BEG[12] ;
 wire \Tile_X6Y5_WW4BEG[13] ;
 wire \Tile_X6Y5_WW4BEG[14] ;
 wire \Tile_X6Y5_WW4BEG[15] ;
 wire \Tile_X6Y5_WW4BEG[1] ;
 wire \Tile_X6Y5_WW4BEG[2] ;
 wire \Tile_X6Y5_WW4BEG[3] ;
 wire \Tile_X6Y5_WW4BEG[4] ;
 wire \Tile_X6Y5_WW4BEG[5] ;
 wire \Tile_X6Y5_WW4BEG[6] ;
 wire \Tile_X6Y5_WW4BEG[7] ;
 wire \Tile_X6Y5_WW4BEG[8] ;
 wire \Tile_X6Y5_WW4BEG[9] ;
 wire Tile_X6Y6_Co;
 wire \Tile_X6Y6_E1BEG[0] ;
 wire \Tile_X6Y6_E1BEG[1] ;
 wire \Tile_X6Y6_E1BEG[2] ;
 wire \Tile_X6Y6_E1BEG[3] ;
 wire \Tile_X6Y6_E2BEG[0] ;
 wire \Tile_X6Y6_E2BEG[1] ;
 wire \Tile_X6Y6_E2BEG[2] ;
 wire \Tile_X6Y6_E2BEG[3] ;
 wire \Tile_X6Y6_E2BEG[4] ;
 wire \Tile_X6Y6_E2BEG[5] ;
 wire \Tile_X6Y6_E2BEG[6] ;
 wire \Tile_X6Y6_E2BEG[7] ;
 wire \Tile_X6Y6_E2BEGb[0] ;
 wire \Tile_X6Y6_E2BEGb[1] ;
 wire \Tile_X6Y6_E2BEGb[2] ;
 wire \Tile_X6Y6_E2BEGb[3] ;
 wire \Tile_X6Y6_E2BEGb[4] ;
 wire \Tile_X6Y6_E2BEGb[5] ;
 wire \Tile_X6Y6_E2BEGb[6] ;
 wire \Tile_X6Y6_E2BEGb[7] ;
 wire \Tile_X6Y6_E6BEG[0] ;
 wire \Tile_X6Y6_E6BEG[10] ;
 wire \Tile_X6Y6_E6BEG[11] ;
 wire \Tile_X6Y6_E6BEG[1] ;
 wire \Tile_X6Y6_E6BEG[2] ;
 wire \Tile_X6Y6_E6BEG[3] ;
 wire \Tile_X6Y6_E6BEG[4] ;
 wire \Tile_X6Y6_E6BEG[5] ;
 wire \Tile_X6Y6_E6BEG[6] ;
 wire \Tile_X6Y6_E6BEG[7] ;
 wire \Tile_X6Y6_E6BEG[8] ;
 wire \Tile_X6Y6_E6BEG[9] ;
 wire \Tile_X6Y6_EE4BEG[0] ;
 wire \Tile_X6Y6_EE4BEG[10] ;
 wire \Tile_X6Y6_EE4BEG[11] ;
 wire \Tile_X6Y6_EE4BEG[12] ;
 wire \Tile_X6Y6_EE4BEG[13] ;
 wire \Tile_X6Y6_EE4BEG[14] ;
 wire \Tile_X6Y6_EE4BEG[15] ;
 wire \Tile_X6Y6_EE4BEG[1] ;
 wire \Tile_X6Y6_EE4BEG[2] ;
 wire \Tile_X6Y6_EE4BEG[3] ;
 wire \Tile_X6Y6_EE4BEG[4] ;
 wire \Tile_X6Y6_EE4BEG[5] ;
 wire \Tile_X6Y6_EE4BEG[6] ;
 wire \Tile_X6Y6_EE4BEG[7] ;
 wire \Tile_X6Y6_EE4BEG[8] ;
 wire \Tile_X6Y6_EE4BEG[9] ;
 wire \Tile_X6Y6_FrameData_O[0] ;
 wire \Tile_X6Y6_FrameData_O[10] ;
 wire \Tile_X6Y6_FrameData_O[11] ;
 wire \Tile_X6Y6_FrameData_O[12] ;
 wire \Tile_X6Y6_FrameData_O[13] ;
 wire \Tile_X6Y6_FrameData_O[14] ;
 wire \Tile_X6Y6_FrameData_O[15] ;
 wire \Tile_X6Y6_FrameData_O[16] ;
 wire \Tile_X6Y6_FrameData_O[17] ;
 wire \Tile_X6Y6_FrameData_O[18] ;
 wire \Tile_X6Y6_FrameData_O[19] ;
 wire \Tile_X6Y6_FrameData_O[1] ;
 wire \Tile_X6Y6_FrameData_O[20] ;
 wire \Tile_X6Y6_FrameData_O[21] ;
 wire \Tile_X6Y6_FrameData_O[22] ;
 wire \Tile_X6Y6_FrameData_O[23] ;
 wire \Tile_X6Y6_FrameData_O[24] ;
 wire \Tile_X6Y6_FrameData_O[25] ;
 wire \Tile_X6Y6_FrameData_O[26] ;
 wire \Tile_X6Y6_FrameData_O[27] ;
 wire \Tile_X6Y6_FrameData_O[28] ;
 wire \Tile_X6Y6_FrameData_O[29] ;
 wire \Tile_X6Y6_FrameData_O[2] ;
 wire \Tile_X6Y6_FrameData_O[30] ;
 wire \Tile_X6Y6_FrameData_O[31] ;
 wire \Tile_X6Y6_FrameData_O[3] ;
 wire \Tile_X6Y6_FrameData_O[4] ;
 wire \Tile_X6Y6_FrameData_O[5] ;
 wire \Tile_X6Y6_FrameData_O[6] ;
 wire \Tile_X6Y6_FrameData_O[7] ;
 wire \Tile_X6Y6_FrameData_O[8] ;
 wire \Tile_X6Y6_FrameData_O[9] ;
 wire \Tile_X6Y6_FrameStrobe_O[0] ;
 wire \Tile_X6Y6_FrameStrobe_O[10] ;
 wire \Tile_X6Y6_FrameStrobe_O[11] ;
 wire \Tile_X6Y6_FrameStrobe_O[12] ;
 wire \Tile_X6Y6_FrameStrobe_O[13] ;
 wire \Tile_X6Y6_FrameStrobe_O[14] ;
 wire \Tile_X6Y6_FrameStrobe_O[15] ;
 wire \Tile_X6Y6_FrameStrobe_O[16] ;
 wire \Tile_X6Y6_FrameStrobe_O[17] ;
 wire \Tile_X6Y6_FrameStrobe_O[18] ;
 wire \Tile_X6Y6_FrameStrobe_O[19] ;
 wire \Tile_X6Y6_FrameStrobe_O[1] ;
 wire \Tile_X6Y6_FrameStrobe_O[2] ;
 wire \Tile_X6Y6_FrameStrobe_O[3] ;
 wire \Tile_X6Y6_FrameStrobe_O[4] ;
 wire \Tile_X6Y6_FrameStrobe_O[5] ;
 wire \Tile_X6Y6_FrameStrobe_O[6] ;
 wire \Tile_X6Y6_FrameStrobe_O[7] ;
 wire \Tile_X6Y6_FrameStrobe_O[8] ;
 wire \Tile_X6Y6_FrameStrobe_O[9] ;
 wire \Tile_X6Y6_N1BEG[0] ;
 wire \Tile_X6Y6_N1BEG[1] ;
 wire \Tile_X6Y6_N1BEG[2] ;
 wire \Tile_X6Y6_N1BEG[3] ;
 wire \Tile_X6Y6_N2BEG[0] ;
 wire \Tile_X6Y6_N2BEG[1] ;
 wire \Tile_X6Y6_N2BEG[2] ;
 wire \Tile_X6Y6_N2BEG[3] ;
 wire \Tile_X6Y6_N2BEG[4] ;
 wire \Tile_X6Y6_N2BEG[5] ;
 wire \Tile_X6Y6_N2BEG[6] ;
 wire \Tile_X6Y6_N2BEG[7] ;
 wire \Tile_X6Y6_N2BEGb[0] ;
 wire \Tile_X6Y6_N2BEGb[1] ;
 wire \Tile_X6Y6_N2BEGb[2] ;
 wire \Tile_X6Y6_N2BEGb[3] ;
 wire \Tile_X6Y6_N2BEGb[4] ;
 wire \Tile_X6Y6_N2BEGb[5] ;
 wire \Tile_X6Y6_N2BEGb[6] ;
 wire \Tile_X6Y6_N2BEGb[7] ;
 wire \Tile_X6Y6_N4BEG[0] ;
 wire \Tile_X6Y6_N4BEG[10] ;
 wire \Tile_X6Y6_N4BEG[11] ;
 wire \Tile_X6Y6_N4BEG[12] ;
 wire \Tile_X6Y6_N4BEG[13] ;
 wire \Tile_X6Y6_N4BEG[14] ;
 wire \Tile_X6Y6_N4BEG[15] ;
 wire \Tile_X6Y6_N4BEG[1] ;
 wire \Tile_X6Y6_N4BEG[2] ;
 wire \Tile_X6Y6_N4BEG[3] ;
 wire \Tile_X6Y6_N4BEG[4] ;
 wire \Tile_X6Y6_N4BEG[5] ;
 wire \Tile_X6Y6_N4BEG[6] ;
 wire \Tile_X6Y6_N4BEG[7] ;
 wire \Tile_X6Y6_N4BEG[8] ;
 wire \Tile_X6Y6_N4BEG[9] ;
 wire \Tile_X6Y6_NN4BEG[0] ;
 wire \Tile_X6Y6_NN4BEG[10] ;
 wire \Tile_X6Y6_NN4BEG[11] ;
 wire \Tile_X6Y6_NN4BEG[12] ;
 wire \Tile_X6Y6_NN4BEG[13] ;
 wire \Tile_X6Y6_NN4BEG[14] ;
 wire \Tile_X6Y6_NN4BEG[15] ;
 wire \Tile_X6Y6_NN4BEG[1] ;
 wire \Tile_X6Y6_NN4BEG[2] ;
 wire \Tile_X6Y6_NN4BEG[3] ;
 wire \Tile_X6Y6_NN4BEG[4] ;
 wire \Tile_X6Y6_NN4BEG[5] ;
 wire \Tile_X6Y6_NN4BEG[6] ;
 wire \Tile_X6Y6_NN4BEG[7] ;
 wire \Tile_X6Y6_NN4BEG[8] ;
 wire \Tile_X6Y6_NN4BEG[9] ;
 wire \Tile_X6Y6_S1BEG[0] ;
 wire \Tile_X6Y6_S1BEG[1] ;
 wire \Tile_X6Y6_S1BEG[2] ;
 wire \Tile_X6Y6_S1BEG[3] ;
 wire \Tile_X6Y6_S2BEG[0] ;
 wire \Tile_X6Y6_S2BEG[1] ;
 wire \Tile_X6Y6_S2BEG[2] ;
 wire \Tile_X6Y6_S2BEG[3] ;
 wire \Tile_X6Y6_S2BEG[4] ;
 wire \Tile_X6Y6_S2BEG[5] ;
 wire \Tile_X6Y6_S2BEG[6] ;
 wire \Tile_X6Y6_S2BEG[7] ;
 wire \Tile_X6Y6_S2BEGb[0] ;
 wire \Tile_X6Y6_S2BEGb[1] ;
 wire \Tile_X6Y6_S2BEGb[2] ;
 wire \Tile_X6Y6_S2BEGb[3] ;
 wire \Tile_X6Y6_S2BEGb[4] ;
 wire \Tile_X6Y6_S2BEGb[5] ;
 wire \Tile_X6Y6_S2BEGb[6] ;
 wire \Tile_X6Y6_S2BEGb[7] ;
 wire \Tile_X6Y6_S4BEG[0] ;
 wire \Tile_X6Y6_S4BEG[10] ;
 wire \Tile_X6Y6_S4BEG[11] ;
 wire \Tile_X6Y6_S4BEG[12] ;
 wire \Tile_X6Y6_S4BEG[13] ;
 wire \Tile_X6Y6_S4BEG[14] ;
 wire \Tile_X6Y6_S4BEG[15] ;
 wire \Tile_X6Y6_S4BEG[1] ;
 wire \Tile_X6Y6_S4BEG[2] ;
 wire \Tile_X6Y6_S4BEG[3] ;
 wire \Tile_X6Y6_S4BEG[4] ;
 wire \Tile_X6Y6_S4BEG[5] ;
 wire \Tile_X6Y6_S4BEG[6] ;
 wire \Tile_X6Y6_S4BEG[7] ;
 wire \Tile_X6Y6_S4BEG[8] ;
 wire \Tile_X6Y6_S4BEG[9] ;
 wire \Tile_X6Y6_SS4BEG[0] ;
 wire \Tile_X6Y6_SS4BEG[10] ;
 wire \Tile_X6Y6_SS4BEG[11] ;
 wire \Tile_X6Y6_SS4BEG[12] ;
 wire \Tile_X6Y6_SS4BEG[13] ;
 wire \Tile_X6Y6_SS4BEG[14] ;
 wire \Tile_X6Y6_SS4BEG[15] ;
 wire \Tile_X6Y6_SS4BEG[1] ;
 wire \Tile_X6Y6_SS4BEG[2] ;
 wire \Tile_X6Y6_SS4BEG[3] ;
 wire \Tile_X6Y6_SS4BEG[4] ;
 wire \Tile_X6Y6_SS4BEG[5] ;
 wire \Tile_X6Y6_SS4BEG[6] ;
 wire \Tile_X6Y6_SS4BEG[7] ;
 wire \Tile_X6Y6_SS4BEG[8] ;
 wire \Tile_X6Y6_SS4BEG[9] ;
 wire Tile_X6Y6_UserCLKo;
 wire \Tile_X6Y6_W1BEG[0] ;
 wire \Tile_X6Y6_W1BEG[1] ;
 wire \Tile_X6Y6_W1BEG[2] ;
 wire \Tile_X6Y6_W1BEG[3] ;
 wire \Tile_X6Y6_W2BEG[0] ;
 wire \Tile_X6Y6_W2BEG[1] ;
 wire \Tile_X6Y6_W2BEG[2] ;
 wire \Tile_X6Y6_W2BEG[3] ;
 wire \Tile_X6Y6_W2BEG[4] ;
 wire \Tile_X6Y6_W2BEG[5] ;
 wire \Tile_X6Y6_W2BEG[6] ;
 wire \Tile_X6Y6_W2BEG[7] ;
 wire \Tile_X6Y6_W2BEGb[0] ;
 wire \Tile_X6Y6_W2BEGb[1] ;
 wire \Tile_X6Y6_W2BEGb[2] ;
 wire \Tile_X6Y6_W2BEGb[3] ;
 wire \Tile_X6Y6_W2BEGb[4] ;
 wire \Tile_X6Y6_W2BEGb[5] ;
 wire \Tile_X6Y6_W2BEGb[6] ;
 wire \Tile_X6Y6_W2BEGb[7] ;
 wire \Tile_X6Y6_W6BEG[0] ;
 wire \Tile_X6Y6_W6BEG[10] ;
 wire \Tile_X6Y6_W6BEG[11] ;
 wire \Tile_X6Y6_W6BEG[1] ;
 wire \Tile_X6Y6_W6BEG[2] ;
 wire \Tile_X6Y6_W6BEG[3] ;
 wire \Tile_X6Y6_W6BEG[4] ;
 wire \Tile_X6Y6_W6BEG[5] ;
 wire \Tile_X6Y6_W6BEG[6] ;
 wire \Tile_X6Y6_W6BEG[7] ;
 wire \Tile_X6Y6_W6BEG[8] ;
 wire \Tile_X6Y6_W6BEG[9] ;
 wire \Tile_X6Y6_WW4BEG[0] ;
 wire \Tile_X6Y6_WW4BEG[10] ;
 wire \Tile_X6Y6_WW4BEG[11] ;
 wire \Tile_X6Y6_WW4BEG[12] ;
 wire \Tile_X6Y6_WW4BEG[13] ;
 wire \Tile_X6Y6_WW4BEG[14] ;
 wire \Tile_X6Y6_WW4BEG[15] ;
 wire \Tile_X6Y6_WW4BEG[1] ;
 wire \Tile_X6Y6_WW4BEG[2] ;
 wire \Tile_X6Y6_WW4BEG[3] ;
 wire \Tile_X6Y6_WW4BEG[4] ;
 wire \Tile_X6Y6_WW4BEG[5] ;
 wire \Tile_X6Y6_WW4BEG[6] ;
 wire \Tile_X6Y6_WW4BEG[7] ;
 wire \Tile_X6Y6_WW4BEG[8] ;
 wire \Tile_X6Y6_WW4BEG[9] ;
 wire Tile_X6Y7_Co;
 wire \Tile_X6Y7_E1BEG[0] ;
 wire \Tile_X6Y7_E1BEG[1] ;
 wire \Tile_X6Y7_E1BEG[2] ;
 wire \Tile_X6Y7_E1BEG[3] ;
 wire \Tile_X6Y7_E2BEG[0] ;
 wire \Tile_X6Y7_E2BEG[1] ;
 wire \Tile_X6Y7_E2BEG[2] ;
 wire \Tile_X6Y7_E2BEG[3] ;
 wire \Tile_X6Y7_E2BEG[4] ;
 wire \Tile_X6Y7_E2BEG[5] ;
 wire \Tile_X6Y7_E2BEG[6] ;
 wire \Tile_X6Y7_E2BEG[7] ;
 wire \Tile_X6Y7_E2BEGb[0] ;
 wire \Tile_X6Y7_E2BEGb[1] ;
 wire \Tile_X6Y7_E2BEGb[2] ;
 wire \Tile_X6Y7_E2BEGb[3] ;
 wire \Tile_X6Y7_E2BEGb[4] ;
 wire \Tile_X6Y7_E2BEGb[5] ;
 wire \Tile_X6Y7_E2BEGb[6] ;
 wire \Tile_X6Y7_E2BEGb[7] ;
 wire \Tile_X6Y7_E6BEG[0] ;
 wire \Tile_X6Y7_E6BEG[10] ;
 wire \Tile_X6Y7_E6BEG[11] ;
 wire \Tile_X6Y7_E6BEG[1] ;
 wire \Tile_X6Y7_E6BEG[2] ;
 wire \Tile_X6Y7_E6BEG[3] ;
 wire \Tile_X6Y7_E6BEG[4] ;
 wire \Tile_X6Y7_E6BEG[5] ;
 wire \Tile_X6Y7_E6BEG[6] ;
 wire \Tile_X6Y7_E6BEG[7] ;
 wire \Tile_X6Y7_E6BEG[8] ;
 wire \Tile_X6Y7_E6BEG[9] ;
 wire \Tile_X6Y7_EE4BEG[0] ;
 wire \Tile_X6Y7_EE4BEG[10] ;
 wire \Tile_X6Y7_EE4BEG[11] ;
 wire \Tile_X6Y7_EE4BEG[12] ;
 wire \Tile_X6Y7_EE4BEG[13] ;
 wire \Tile_X6Y7_EE4BEG[14] ;
 wire \Tile_X6Y7_EE4BEG[15] ;
 wire \Tile_X6Y7_EE4BEG[1] ;
 wire \Tile_X6Y7_EE4BEG[2] ;
 wire \Tile_X6Y7_EE4BEG[3] ;
 wire \Tile_X6Y7_EE4BEG[4] ;
 wire \Tile_X6Y7_EE4BEG[5] ;
 wire \Tile_X6Y7_EE4BEG[6] ;
 wire \Tile_X6Y7_EE4BEG[7] ;
 wire \Tile_X6Y7_EE4BEG[8] ;
 wire \Tile_X6Y7_EE4BEG[9] ;
 wire \Tile_X6Y7_FrameData_O[0] ;
 wire \Tile_X6Y7_FrameData_O[10] ;
 wire \Tile_X6Y7_FrameData_O[11] ;
 wire \Tile_X6Y7_FrameData_O[12] ;
 wire \Tile_X6Y7_FrameData_O[13] ;
 wire \Tile_X6Y7_FrameData_O[14] ;
 wire \Tile_X6Y7_FrameData_O[15] ;
 wire \Tile_X6Y7_FrameData_O[16] ;
 wire \Tile_X6Y7_FrameData_O[17] ;
 wire \Tile_X6Y7_FrameData_O[18] ;
 wire \Tile_X6Y7_FrameData_O[19] ;
 wire \Tile_X6Y7_FrameData_O[1] ;
 wire \Tile_X6Y7_FrameData_O[20] ;
 wire \Tile_X6Y7_FrameData_O[21] ;
 wire \Tile_X6Y7_FrameData_O[22] ;
 wire \Tile_X6Y7_FrameData_O[23] ;
 wire \Tile_X6Y7_FrameData_O[24] ;
 wire \Tile_X6Y7_FrameData_O[25] ;
 wire \Tile_X6Y7_FrameData_O[26] ;
 wire \Tile_X6Y7_FrameData_O[27] ;
 wire \Tile_X6Y7_FrameData_O[28] ;
 wire \Tile_X6Y7_FrameData_O[29] ;
 wire \Tile_X6Y7_FrameData_O[2] ;
 wire \Tile_X6Y7_FrameData_O[30] ;
 wire \Tile_X6Y7_FrameData_O[31] ;
 wire \Tile_X6Y7_FrameData_O[3] ;
 wire \Tile_X6Y7_FrameData_O[4] ;
 wire \Tile_X6Y7_FrameData_O[5] ;
 wire \Tile_X6Y7_FrameData_O[6] ;
 wire \Tile_X6Y7_FrameData_O[7] ;
 wire \Tile_X6Y7_FrameData_O[8] ;
 wire \Tile_X6Y7_FrameData_O[9] ;
 wire \Tile_X6Y7_FrameStrobe_O[0] ;
 wire \Tile_X6Y7_FrameStrobe_O[10] ;
 wire \Tile_X6Y7_FrameStrobe_O[11] ;
 wire \Tile_X6Y7_FrameStrobe_O[12] ;
 wire \Tile_X6Y7_FrameStrobe_O[13] ;
 wire \Tile_X6Y7_FrameStrobe_O[14] ;
 wire \Tile_X6Y7_FrameStrobe_O[15] ;
 wire \Tile_X6Y7_FrameStrobe_O[16] ;
 wire \Tile_X6Y7_FrameStrobe_O[17] ;
 wire \Tile_X6Y7_FrameStrobe_O[18] ;
 wire \Tile_X6Y7_FrameStrobe_O[19] ;
 wire \Tile_X6Y7_FrameStrobe_O[1] ;
 wire \Tile_X6Y7_FrameStrobe_O[2] ;
 wire \Tile_X6Y7_FrameStrobe_O[3] ;
 wire \Tile_X6Y7_FrameStrobe_O[4] ;
 wire \Tile_X6Y7_FrameStrobe_O[5] ;
 wire \Tile_X6Y7_FrameStrobe_O[6] ;
 wire \Tile_X6Y7_FrameStrobe_O[7] ;
 wire \Tile_X6Y7_FrameStrobe_O[8] ;
 wire \Tile_X6Y7_FrameStrobe_O[9] ;
 wire \Tile_X6Y7_N1BEG[0] ;
 wire \Tile_X6Y7_N1BEG[1] ;
 wire \Tile_X6Y7_N1BEG[2] ;
 wire \Tile_X6Y7_N1BEG[3] ;
 wire \Tile_X6Y7_N2BEG[0] ;
 wire \Tile_X6Y7_N2BEG[1] ;
 wire \Tile_X6Y7_N2BEG[2] ;
 wire \Tile_X6Y7_N2BEG[3] ;
 wire \Tile_X6Y7_N2BEG[4] ;
 wire \Tile_X6Y7_N2BEG[5] ;
 wire \Tile_X6Y7_N2BEG[6] ;
 wire \Tile_X6Y7_N2BEG[7] ;
 wire \Tile_X6Y7_N2BEGb[0] ;
 wire \Tile_X6Y7_N2BEGb[1] ;
 wire \Tile_X6Y7_N2BEGb[2] ;
 wire \Tile_X6Y7_N2BEGb[3] ;
 wire \Tile_X6Y7_N2BEGb[4] ;
 wire \Tile_X6Y7_N2BEGb[5] ;
 wire \Tile_X6Y7_N2BEGb[6] ;
 wire \Tile_X6Y7_N2BEGb[7] ;
 wire \Tile_X6Y7_N4BEG[0] ;
 wire \Tile_X6Y7_N4BEG[10] ;
 wire \Tile_X6Y7_N4BEG[11] ;
 wire \Tile_X6Y7_N4BEG[12] ;
 wire \Tile_X6Y7_N4BEG[13] ;
 wire \Tile_X6Y7_N4BEG[14] ;
 wire \Tile_X6Y7_N4BEG[15] ;
 wire \Tile_X6Y7_N4BEG[1] ;
 wire \Tile_X6Y7_N4BEG[2] ;
 wire \Tile_X6Y7_N4BEG[3] ;
 wire \Tile_X6Y7_N4BEG[4] ;
 wire \Tile_X6Y7_N4BEG[5] ;
 wire \Tile_X6Y7_N4BEG[6] ;
 wire \Tile_X6Y7_N4BEG[7] ;
 wire \Tile_X6Y7_N4BEG[8] ;
 wire \Tile_X6Y7_N4BEG[9] ;
 wire \Tile_X6Y7_NN4BEG[0] ;
 wire \Tile_X6Y7_NN4BEG[10] ;
 wire \Tile_X6Y7_NN4BEG[11] ;
 wire \Tile_X6Y7_NN4BEG[12] ;
 wire \Tile_X6Y7_NN4BEG[13] ;
 wire \Tile_X6Y7_NN4BEG[14] ;
 wire \Tile_X6Y7_NN4BEG[15] ;
 wire \Tile_X6Y7_NN4BEG[1] ;
 wire \Tile_X6Y7_NN4BEG[2] ;
 wire \Tile_X6Y7_NN4BEG[3] ;
 wire \Tile_X6Y7_NN4BEG[4] ;
 wire \Tile_X6Y7_NN4BEG[5] ;
 wire \Tile_X6Y7_NN4BEG[6] ;
 wire \Tile_X6Y7_NN4BEG[7] ;
 wire \Tile_X6Y7_NN4BEG[8] ;
 wire \Tile_X6Y7_NN4BEG[9] ;
 wire \Tile_X6Y7_S1BEG[0] ;
 wire \Tile_X6Y7_S1BEG[1] ;
 wire \Tile_X6Y7_S1BEG[2] ;
 wire \Tile_X6Y7_S1BEG[3] ;
 wire \Tile_X6Y7_S2BEG[0] ;
 wire \Tile_X6Y7_S2BEG[1] ;
 wire \Tile_X6Y7_S2BEG[2] ;
 wire \Tile_X6Y7_S2BEG[3] ;
 wire \Tile_X6Y7_S2BEG[4] ;
 wire \Tile_X6Y7_S2BEG[5] ;
 wire \Tile_X6Y7_S2BEG[6] ;
 wire \Tile_X6Y7_S2BEG[7] ;
 wire \Tile_X6Y7_S2BEGb[0] ;
 wire \Tile_X6Y7_S2BEGb[1] ;
 wire \Tile_X6Y7_S2BEGb[2] ;
 wire \Tile_X6Y7_S2BEGb[3] ;
 wire \Tile_X6Y7_S2BEGb[4] ;
 wire \Tile_X6Y7_S2BEGb[5] ;
 wire \Tile_X6Y7_S2BEGb[6] ;
 wire \Tile_X6Y7_S2BEGb[7] ;
 wire \Tile_X6Y7_S4BEG[0] ;
 wire \Tile_X6Y7_S4BEG[10] ;
 wire \Tile_X6Y7_S4BEG[11] ;
 wire \Tile_X6Y7_S4BEG[12] ;
 wire \Tile_X6Y7_S4BEG[13] ;
 wire \Tile_X6Y7_S4BEG[14] ;
 wire \Tile_X6Y7_S4BEG[15] ;
 wire \Tile_X6Y7_S4BEG[1] ;
 wire \Tile_X6Y7_S4BEG[2] ;
 wire \Tile_X6Y7_S4BEG[3] ;
 wire \Tile_X6Y7_S4BEG[4] ;
 wire \Tile_X6Y7_S4BEG[5] ;
 wire \Tile_X6Y7_S4BEG[6] ;
 wire \Tile_X6Y7_S4BEG[7] ;
 wire \Tile_X6Y7_S4BEG[8] ;
 wire \Tile_X6Y7_S4BEG[9] ;
 wire \Tile_X6Y7_SS4BEG[0] ;
 wire \Tile_X6Y7_SS4BEG[10] ;
 wire \Tile_X6Y7_SS4BEG[11] ;
 wire \Tile_X6Y7_SS4BEG[12] ;
 wire \Tile_X6Y7_SS4BEG[13] ;
 wire \Tile_X6Y7_SS4BEG[14] ;
 wire \Tile_X6Y7_SS4BEG[15] ;
 wire \Tile_X6Y7_SS4BEG[1] ;
 wire \Tile_X6Y7_SS4BEG[2] ;
 wire \Tile_X6Y7_SS4BEG[3] ;
 wire \Tile_X6Y7_SS4BEG[4] ;
 wire \Tile_X6Y7_SS4BEG[5] ;
 wire \Tile_X6Y7_SS4BEG[6] ;
 wire \Tile_X6Y7_SS4BEG[7] ;
 wire \Tile_X6Y7_SS4BEG[8] ;
 wire \Tile_X6Y7_SS4BEG[9] ;
 wire Tile_X6Y7_UserCLKo;
 wire \Tile_X6Y7_W1BEG[0] ;
 wire \Tile_X6Y7_W1BEG[1] ;
 wire \Tile_X6Y7_W1BEG[2] ;
 wire \Tile_X6Y7_W1BEG[3] ;
 wire \Tile_X6Y7_W2BEG[0] ;
 wire \Tile_X6Y7_W2BEG[1] ;
 wire \Tile_X6Y7_W2BEG[2] ;
 wire \Tile_X6Y7_W2BEG[3] ;
 wire \Tile_X6Y7_W2BEG[4] ;
 wire \Tile_X6Y7_W2BEG[5] ;
 wire \Tile_X6Y7_W2BEG[6] ;
 wire \Tile_X6Y7_W2BEG[7] ;
 wire \Tile_X6Y7_W2BEGb[0] ;
 wire \Tile_X6Y7_W2BEGb[1] ;
 wire \Tile_X6Y7_W2BEGb[2] ;
 wire \Tile_X6Y7_W2BEGb[3] ;
 wire \Tile_X6Y7_W2BEGb[4] ;
 wire \Tile_X6Y7_W2BEGb[5] ;
 wire \Tile_X6Y7_W2BEGb[6] ;
 wire \Tile_X6Y7_W2BEGb[7] ;
 wire \Tile_X6Y7_W6BEG[0] ;
 wire \Tile_X6Y7_W6BEG[10] ;
 wire \Tile_X6Y7_W6BEG[11] ;
 wire \Tile_X6Y7_W6BEG[1] ;
 wire \Tile_X6Y7_W6BEG[2] ;
 wire \Tile_X6Y7_W6BEG[3] ;
 wire \Tile_X6Y7_W6BEG[4] ;
 wire \Tile_X6Y7_W6BEG[5] ;
 wire \Tile_X6Y7_W6BEG[6] ;
 wire \Tile_X6Y7_W6BEG[7] ;
 wire \Tile_X6Y7_W6BEG[8] ;
 wire \Tile_X6Y7_W6BEG[9] ;
 wire \Tile_X6Y7_WW4BEG[0] ;
 wire \Tile_X6Y7_WW4BEG[10] ;
 wire \Tile_X6Y7_WW4BEG[11] ;
 wire \Tile_X6Y7_WW4BEG[12] ;
 wire \Tile_X6Y7_WW4BEG[13] ;
 wire \Tile_X6Y7_WW4BEG[14] ;
 wire \Tile_X6Y7_WW4BEG[15] ;
 wire \Tile_X6Y7_WW4BEG[1] ;
 wire \Tile_X6Y7_WW4BEG[2] ;
 wire \Tile_X6Y7_WW4BEG[3] ;
 wire \Tile_X6Y7_WW4BEG[4] ;
 wire \Tile_X6Y7_WW4BEG[5] ;
 wire \Tile_X6Y7_WW4BEG[6] ;
 wire \Tile_X6Y7_WW4BEG[7] ;
 wire \Tile_X6Y7_WW4BEG[8] ;
 wire \Tile_X6Y7_WW4BEG[9] ;
 wire Tile_X6Y8_Co;
 wire \Tile_X6Y8_E1BEG[0] ;
 wire \Tile_X6Y8_E1BEG[1] ;
 wire \Tile_X6Y8_E1BEG[2] ;
 wire \Tile_X6Y8_E1BEG[3] ;
 wire \Tile_X6Y8_E2BEG[0] ;
 wire \Tile_X6Y8_E2BEG[1] ;
 wire \Tile_X6Y8_E2BEG[2] ;
 wire \Tile_X6Y8_E2BEG[3] ;
 wire \Tile_X6Y8_E2BEG[4] ;
 wire \Tile_X6Y8_E2BEG[5] ;
 wire \Tile_X6Y8_E2BEG[6] ;
 wire \Tile_X6Y8_E2BEG[7] ;
 wire \Tile_X6Y8_E2BEGb[0] ;
 wire \Tile_X6Y8_E2BEGb[1] ;
 wire \Tile_X6Y8_E2BEGb[2] ;
 wire \Tile_X6Y8_E2BEGb[3] ;
 wire \Tile_X6Y8_E2BEGb[4] ;
 wire \Tile_X6Y8_E2BEGb[5] ;
 wire \Tile_X6Y8_E2BEGb[6] ;
 wire \Tile_X6Y8_E2BEGb[7] ;
 wire \Tile_X6Y8_E6BEG[0] ;
 wire \Tile_X6Y8_E6BEG[10] ;
 wire \Tile_X6Y8_E6BEG[11] ;
 wire \Tile_X6Y8_E6BEG[1] ;
 wire \Tile_X6Y8_E6BEG[2] ;
 wire \Tile_X6Y8_E6BEG[3] ;
 wire \Tile_X6Y8_E6BEG[4] ;
 wire \Tile_X6Y8_E6BEG[5] ;
 wire \Tile_X6Y8_E6BEG[6] ;
 wire \Tile_X6Y8_E6BEG[7] ;
 wire \Tile_X6Y8_E6BEG[8] ;
 wire \Tile_X6Y8_E6BEG[9] ;
 wire \Tile_X6Y8_EE4BEG[0] ;
 wire \Tile_X6Y8_EE4BEG[10] ;
 wire \Tile_X6Y8_EE4BEG[11] ;
 wire \Tile_X6Y8_EE4BEG[12] ;
 wire \Tile_X6Y8_EE4BEG[13] ;
 wire \Tile_X6Y8_EE4BEG[14] ;
 wire \Tile_X6Y8_EE4BEG[15] ;
 wire \Tile_X6Y8_EE4BEG[1] ;
 wire \Tile_X6Y8_EE4BEG[2] ;
 wire \Tile_X6Y8_EE4BEG[3] ;
 wire \Tile_X6Y8_EE4BEG[4] ;
 wire \Tile_X6Y8_EE4BEG[5] ;
 wire \Tile_X6Y8_EE4BEG[6] ;
 wire \Tile_X6Y8_EE4BEG[7] ;
 wire \Tile_X6Y8_EE4BEG[8] ;
 wire \Tile_X6Y8_EE4BEG[9] ;
 wire \Tile_X6Y8_FrameData_O[0] ;
 wire \Tile_X6Y8_FrameData_O[10] ;
 wire \Tile_X6Y8_FrameData_O[11] ;
 wire \Tile_X6Y8_FrameData_O[12] ;
 wire \Tile_X6Y8_FrameData_O[13] ;
 wire \Tile_X6Y8_FrameData_O[14] ;
 wire \Tile_X6Y8_FrameData_O[15] ;
 wire \Tile_X6Y8_FrameData_O[16] ;
 wire \Tile_X6Y8_FrameData_O[17] ;
 wire \Tile_X6Y8_FrameData_O[18] ;
 wire \Tile_X6Y8_FrameData_O[19] ;
 wire \Tile_X6Y8_FrameData_O[1] ;
 wire \Tile_X6Y8_FrameData_O[20] ;
 wire \Tile_X6Y8_FrameData_O[21] ;
 wire \Tile_X6Y8_FrameData_O[22] ;
 wire \Tile_X6Y8_FrameData_O[23] ;
 wire \Tile_X6Y8_FrameData_O[24] ;
 wire \Tile_X6Y8_FrameData_O[25] ;
 wire \Tile_X6Y8_FrameData_O[26] ;
 wire \Tile_X6Y8_FrameData_O[27] ;
 wire \Tile_X6Y8_FrameData_O[28] ;
 wire \Tile_X6Y8_FrameData_O[29] ;
 wire \Tile_X6Y8_FrameData_O[2] ;
 wire \Tile_X6Y8_FrameData_O[30] ;
 wire \Tile_X6Y8_FrameData_O[31] ;
 wire \Tile_X6Y8_FrameData_O[3] ;
 wire \Tile_X6Y8_FrameData_O[4] ;
 wire \Tile_X6Y8_FrameData_O[5] ;
 wire \Tile_X6Y8_FrameData_O[6] ;
 wire \Tile_X6Y8_FrameData_O[7] ;
 wire \Tile_X6Y8_FrameData_O[8] ;
 wire \Tile_X6Y8_FrameData_O[9] ;
 wire \Tile_X6Y8_FrameStrobe_O[0] ;
 wire \Tile_X6Y8_FrameStrobe_O[10] ;
 wire \Tile_X6Y8_FrameStrobe_O[11] ;
 wire \Tile_X6Y8_FrameStrobe_O[12] ;
 wire \Tile_X6Y8_FrameStrobe_O[13] ;
 wire \Tile_X6Y8_FrameStrobe_O[14] ;
 wire \Tile_X6Y8_FrameStrobe_O[15] ;
 wire \Tile_X6Y8_FrameStrobe_O[16] ;
 wire \Tile_X6Y8_FrameStrobe_O[17] ;
 wire \Tile_X6Y8_FrameStrobe_O[18] ;
 wire \Tile_X6Y8_FrameStrobe_O[19] ;
 wire \Tile_X6Y8_FrameStrobe_O[1] ;
 wire \Tile_X6Y8_FrameStrobe_O[2] ;
 wire \Tile_X6Y8_FrameStrobe_O[3] ;
 wire \Tile_X6Y8_FrameStrobe_O[4] ;
 wire \Tile_X6Y8_FrameStrobe_O[5] ;
 wire \Tile_X6Y8_FrameStrobe_O[6] ;
 wire \Tile_X6Y8_FrameStrobe_O[7] ;
 wire \Tile_X6Y8_FrameStrobe_O[8] ;
 wire \Tile_X6Y8_FrameStrobe_O[9] ;
 wire \Tile_X6Y8_N1BEG[0] ;
 wire \Tile_X6Y8_N1BEG[1] ;
 wire \Tile_X6Y8_N1BEG[2] ;
 wire \Tile_X6Y8_N1BEG[3] ;
 wire \Tile_X6Y8_N2BEG[0] ;
 wire \Tile_X6Y8_N2BEG[1] ;
 wire \Tile_X6Y8_N2BEG[2] ;
 wire \Tile_X6Y8_N2BEG[3] ;
 wire \Tile_X6Y8_N2BEG[4] ;
 wire \Tile_X6Y8_N2BEG[5] ;
 wire \Tile_X6Y8_N2BEG[6] ;
 wire \Tile_X6Y8_N2BEG[7] ;
 wire \Tile_X6Y8_N2BEGb[0] ;
 wire \Tile_X6Y8_N2BEGb[1] ;
 wire \Tile_X6Y8_N2BEGb[2] ;
 wire \Tile_X6Y8_N2BEGb[3] ;
 wire \Tile_X6Y8_N2BEGb[4] ;
 wire \Tile_X6Y8_N2BEGb[5] ;
 wire \Tile_X6Y8_N2BEGb[6] ;
 wire \Tile_X6Y8_N2BEGb[7] ;
 wire \Tile_X6Y8_N4BEG[0] ;
 wire \Tile_X6Y8_N4BEG[10] ;
 wire \Tile_X6Y8_N4BEG[11] ;
 wire \Tile_X6Y8_N4BEG[12] ;
 wire \Tile_X6Y8_N4BEG[13] ;
 wire \Tile_X6Y8_N4BEG[14] ;
 wire \Tile_X6Y8_N4BEG[15] ;
 wire \Tile_X6Y8_N4BEG[1] ;
 wire \Tile_X6Y8_N4BEG[2] ;
 wire \Tile_X6Y8_N4BEG[3] ;
 wire \Tile_X6Y8_N4BEG[4] ;
 wire \Tile_X6Y8_N4BEG[5] ;
 wire \Tile_X6Y8_N4BEG[6] ;
 wire \Tile_X6Y8_N4BEG[7] ;
 wire \Tile_X6Y8_N4BEG[8] ;
 wire \Tile_X6Y8_N4BEG[9] ;
 wire \Tile_X6Y8_NN4BEG[0] ;
 wire \Tile_X6Y8_NN4BEG[10] ;
 wire \Tile_X6Y8_NN4BEG[11] ;
 wire \Tile_X6Y8_NN4BEG[12] ;
 wire \Tile_X6Y8_NN4BEG[13] ;
 wire \Tile_X6Y8_NN4BEG[14] ;
 wire \Tile_X6Y8_NN4BEG[15] ;
 wire \Tile_X6Y8_NN4BEG[1] ;
 wire \Tile_X6Y8_NN4BEG[2] ;
 wire \Tile_X6Y8_NN4BEG[3] ;
 wire \Tile_X6Y8_NN4BEG[4] ;
 wire \Tile_X6Y8_NN4BEG[5] ;
 wire \Tile_X6Y8_NN4BEG[6] ;
 wire \Tile_X6Y8_NN4BEG[7] ;
 wire \Tile_X6Y8_NN4BEG[8] ;
 wire \Tile_X6Y8_NN4BEG[9] ;
 wire \Tile_X6Y8_S1BEG[0] ;
 wire \Tile_X6Y8_S1BEG[1] ;
 wire \Tile_X6Y8_S1BEG[2] ;
 wire \Tile_X6Y8_S1BEG[3] ;
 wire \Tile_X6Y8_S2BEG[0] ;
 wire \Tile_X6Y8_S2BEG[1] ;
 wire \Tile_X6Y8_S2BEG[2] ;
 wire \Tile_X6Y8_S2BEG[3] ;
 wire \Tile_X6Y8_S2BEG[4] ;
 wire \Tile_X6Y8_S2BEG[5] ;
 wire \Tile_X6Y8_S2BEG[6] ;
 wire \Tile_X6Y8_S2BEG[7] ;
 wire \Tile_X6Y8_S2BEGb[0] ;
 wire \Tile_X6Y8_S2BEGb[1] ;
 wire \Tile_X6Y8_S2BEGb[2] ;
 wire \Tile_X6Y8_S2BEGb[3] ;
 wire \Tile_X6Y8_S2BEGb[4] ;
 wire \Tile_X6Y8_S2BEGb[5] ;
 wire \Tile_X6Y8_S2BEGb[6] ;
 wire \Tile_X6Y8_S2BEGb[7] ;
 wire \Tile_X6Y8_S4BEG[0] ;
 wire \Tile_X6Y8_S4BEG[10] ;
 wire \Tile_X6Y8_S4BEG[11] ;
 wire \Tile_X6Y8_S4BEG[12] ;
 wire \Tile_X6Y8_S4BEG[13] ;
 wire \Tile_X6Y8_S4BEG[14] ;
 wire \Tile_X6Y8_S4BEG[15] ;
 wire \Tile_X6Y8_S4BEG[1] ;
 wire \Tile_X6Y8_S4BEG[2] ;
 wire \Tile_X6Y8_S4BEG[3] ;
 wire \Tile_X6Y8_S4BEG[4] ;
 wire \Tile_X6Y8_S4BEG[5] ;
 wire \Tile_X6Y8_S4BEG[6] ;
 wire \Tile_X6Y8_S4BEG[7] ;
 wire \Tile_X6Y8_S4BEG[8] ;
 wire \Tile_X6Y8_S4BEG[9] ;
 wire \Tile_X6Y8_SS4BEG[0] ;
 wire \Tile_X6Y8_SS4BEG[10] ;
 wire \Tile_X6Y8_SS4BEG[11] ;
 wire \Tile_X6Y8_SS4BEG[12] ;
 wire \Tile_X6Y8_SS4BEG[13] ;
 wire \Tile_X6Y8_SS4BEG[14] ;
 wire \Tile_X6Y8_SS4BEG[15] ;
 wire \Tile_X6Y8_SS4BEG[1] ;
 wire \Tile_X6Y8_SS4BEG[2] ;
 wire \Tile_X6Y8_SS4BEG[3] ;
 wire \Tile_X6Y8_SS4BEG[4] ;
 wire \Tile_X6Y8_SS4BEG[5] ;
 wire \Tile_X6Y8_SS4BEG[6] ;
 wire \Tile_X6Y8_SS4BEG[7] ;
 wire \Tile_X6Y8_SS4BEG[8] ;
 wire \Tile_X6Y8_SS4BEG[9] ;
 wire Tile_X6Y8_UserCLKo;
 wire \Tile_X6Y8_W1BEG[0] ;
 wire \Tile_X6Y8_W1BEG[1] ;
 wire \Tile_X6Y8_W1BEG[2] ;
 wire \Tile_X6Y8_W1BEG[3] ;
 wire \Tile_X6Y8_W2BEG[0] ;
 wire \Tile_X6Y8_W2BEG[1] ;
 wire \Tile_X6Y8_W2BEG[2] ;
 wire \Tile_X6Y8_W2BEG[3] ;
 wire \Tile_X6Y8_W2BEG[4] ;
 wire \Tile_X6Y8_W2BEG[5] ;
 wire \Tile_X6Y8_W2BEG[6] ;
 wire \Tile_X6Y8_W2BEG[7] ;
 wire \Tile_X6Y8_W2BEGb[0] ;
 wire \Tile_X6Y8_W2BEGb[1] ;
 wire \Tile_X6Y8_W2BEGb[2] ;
 wire \Tile_X6Y8_W2BEGb[3] ;
 wire \Tile_X6Y8_W2BEGb[4] ;
 wire \Tile_X6Y8_W2BEGb[5] ;
 wire \Tile_X6Y8_W2BEGb[6] ;
 wire \Tile_X6Y8_W2BEGb[7] ;
 wire \Tile_X6Y8_W6BEG[0] ;
 wire \Tile_X6Y8_W6BEG[10] ;
 wire \Tile_X6Y8_W6BEG[11] ;
 wire \Tile_X6Y8_W6BEG[1] ;
 wire \Tile_X6Y8_W6BEG[2] ;
 wire \Tile_X6Y8_W6BEG[3] ;
 wire \Tile_X6Y8_W6BEG[4] ;
 wire \Tile_X6Y8_W6BEG[5] ;
 wire \Tile_X6Y8_W6BEG[6] ;
 wire \Tile_X6Y8_W6BEG[7] ;
 wire \Tile_X6Y8_W6BEG[8] ;
 wire \Tile_X6Y8_W6BEG[9] ;
 wire \Tile_X6Y8_WW4BEG[0] ;
 wire \Tile_X6Y8_WW4BEG[10] ;
 wire \Tile_X6Y8_WW4BEG[11] ;
 wire \Tile_X6Y8_WW4BEG[12] ;
 wire \Tile_X6Y8_WW4BEG[13] ;
 wire \Tile_X6Y8_WW4BEG[14] ;
 wire \Tile_X6Y8_WW4BEG[15] ;
 wire \Tile_X6Y8_WW4BEG[1] ;
 wire \Tile_X6Y8_WW4BEG[2] ;
 wire \Tile_X6Y8_WW4BEG[3] ;
 wire \Tile_X6Y8_WW4BEG[4] ;
 wire \Tile_X6Y8_WW4BEG[5] ;
 wire \Tile_X6Y8_WW4BEG[6] ;
 wire \Tile_X6Y8_WW4BEG[7] ;
 wire \Tile_X6Y8_WW4BEG[8] ;
 wire \Tile_X6Y8_WW4BEG[9] ;
 wire Tile_X6Y9_Co;
 wire \Tile_X6Y9_E1BEG[0] ;
 wire \Tile_X6Y9_E1BEG[1] ;
 wire \Tile_X6Y9_E1BEG[2] ;
 wire \Tile_X6Y9_E1BEG[3] ;
 wire \Tile_X6Y9_E2BEG[0] ;
 wire \Tile_X6Y9_E2BEG[1] ;
 wire \Tile_X6Y9_E2BEG[2] ;
 wire \Tile_X6Y9_E2BEG[3] ;
 wire \Tile_X6Y9_E2BEG[4] ;
 wire \Tile_X6Y9_E2BEG[5] ;
 wire \Tile_X6Y9_E2BEG[6] ;
 wire \Tile_X6Y9_E2BEG[7] ;
 wire \Tile_X6Y9_E2BEGb[0] ;
 wire \Tile_X6Y9_E2BEGb[1] ;
 wire \Tile_X6Y9_E2BEGb[2] ;
 wire \Tile_X6Y9_E2BEGb[3] ;
 wire \Tile_X6Y9_E2BEGb[4] ;
 wire \Tile_X6Y9_E2BEGb[5] ;
 wire \Tile_X6Y9_E2BEGb[6] ;
 wire \Tile_X6Y9_E2BEGb[7] ;
 wire \Tile_X6Y9_E6BEG[0] ;
 wire \Tile_X6Y9_E6BEG[10] ;
 wire \Tile_X6Y9_E6BEG[11] ;
 wire \Tile_X6Y9_E6BEG[1] ;
 wire \Tile_X6Y9_E6BEG[2] ;
 wire \Tile_X6Y9_E6BEG[3] ;
 wire \Tile_X6Y9_E6BEG[4] ;
 wire \Tile_X6Y9_E6BEG[5] ;
 wire \Tile_X6Y9_E6BEG[6] ;
 wire \Tile_X6Y9_E6BEG[7] ;
 wire \Tile_X6Y9_E6BEG[8] ;
 wire \Tile_X6Y9_E6BEG[9] ;
 wire \Tile_X6Y9_EE4BEG[0] ;
 wire \Tile_X6Y9_EE4BEG[10] ;
 wire \Tile_X6Y9_EE4BEG[11] ;
 wire \Tile_X6Y9_EE4BEG[12] ;
 wire \Tile_X6Y9_EE4BEG[13] ;
 wire \Tile_X6Y9_EE4BEG[14] ;
 wire \Tile_X6Y9_EE4BEG[15] ;
 wire \Tile_X6Y9_EE4BEG[1] ;
 wire \Tile_X6Y9_EE4BEG[2] ;
 wire \Tile_X6Y9_EE4BEG[3] ;
 wire \Tile_X6Y9_EE4BEG[4] ;
 wire \Tile_X6Y9_EE4BEG[5] ;
 wire \Tile_X6Y9_EE4BEG[6] ;
 wire \Tile_X6Y9_EE4BEG[7] ;
 wire \Tile_X6Y9_EE4BEG[8] ;
 wire \Tile_X6Y9_EE4BEG[9] ;
 wire \Tile_X6Y9_FrameData_O[0] ;
 wire \Tile_X6Y9_FrameData_O[10] ;
 wire \Tile_X6Y9_FrameData_O[11] ;
 wire \Tile_X6Y9_FrameData_O[12] ;
 wire \Tile_X6Y9_FrameData_O[13] ;
 wire \Tile_X6Y9_FrameData_O[14] ;
 wire \Tile_X6Y9_FrameData_O[15] ;
 wire \Tile_X6Y9_FrameData_O[16] ;
 wire \Tile_X6Y9_FrameData_O[17] ;
 wire \Tile_X6Y9_FrameData_O[18] ;
 wire \Tile_X6Y9_FrameData_O[19] ;
 wire \Tile_X6Y9_FrameData_O[1] ;
 wire \Tile_X6Y9_FrameData_O[20] ;
 wire \Tile_X6Y9_FrameData_O[21] ;
 wire \Tile_X6Y9_FrameData_O[22] ;
 wire \Tile_X6Y9_FrameData_O[23] ;
 wire \Tile_X6Y9_FrameData_O[24] ;
 wire \Tile_X6Y9_FrameData_O[25] ;
 wire \Tile_X6Y9_FrameData_O[26] ;
 wire \Tile_X6Y9_FrameData_O[27] ;
 wire \Tile_X6Y9_FrameData_O[28] ;
 wire \Tile_X6Y9_FrameData_O[29] ;
 wire \Tile_X6Y9_FrameData_O[2] ;
 wire \Tile_X6Y9_FrameData_O[30] ;
 wire \Tile_X6Y9_FrameData_O[31] ;
 wire \Tile_X6Y9_FrameData_O[3] ;
 wire \Tile_X6Y9_FrameData_O[4] ;
 wire \Tile_X6Y9_FrameData_O[5] ;
 wire \Tile_X6Y9_FrameData_O[6] ;
 wire \Tile_X6Y9_FrameData_O[7] ;
 wire \Tile_X6Y9_FrameData_O[8] ;
 wire \Tile_X6Y9_FrameData_O[9] ;
 wire \Tile_X6Y9_FrameStrobe_O[0] ;
 wire \Tile_X6Y9_FrameStrobe_O[10] ;
 wire \Tile_X6Y9_FrameStrobe_O[11] ;
 wire \Tile_X6Y9_FrameStrobe_O[12] ;
 wire \Tile_X6Y9_FrameStrobe_O[13] ;
 wire \Tile_X6Y9_FrameStrobe_O[14] ;
 wire \Tile_X6Y9_FrameStrobe_O[15] ;
 wire \Tile_X6Y9_FrameStrobe_O[16] ;
 wire \Tile_X6Y9_FrameStrobe_O[17] ;
 wire \Tile_X6Y9_FrameStrobe_O[18] ;
 wire \Tile_X6Y9_FrameStrobe_O[19] ;
 wire \Tile_X6Y9_FrameStrobe_O[1] ;
 wire \Tile_X6Y9_FrameStrobe_O[2] ;
 wire \Tile_X6Y9_FrameStrobe_O[3] ;
 wire \Tile_X6Y9_FrameStrobe_O[4] ;
 wire \Tile_X6Y9_FrameStrobe_O[5] ;
 wire \Tile_X6Y9_FrameStrobe_O[6] ;
 wire \Tile_X6Y9_FrameStrobe_O[7] ;
 wire \Tile_X6Y9_FrameStrobe_O[8] ;
 wire \Tile_X6Y9_FrameStrobe_O[9] ;
 wire \Tile_X6Y9_N1BEG[0] ;
 wire \Tile_X6Y9_N1BEG[1] ;
 wire \Tile_X6Y9_N1BEG[2] ;
 wire \Tile_X6Y9_N1BEG[3] ;
 wire \Tile_X6Y9_N2BEG[0] ;
 wire \Tile_X6Y9_N2BEG[1] ;
 wire \Tile_X6Y9_N2BEG[2] ;
 wire \Tile_X6Y9_N2BEG[3] ;
 wire \Tile_X6Y9_N2BEG[4] ;
 wire \Tile_X6Y9_N2BEG[5] ;
 wire \Tile_X6Y9_N2BEG[6] ;
 wire \Tile_X6Y9_N2BEG[7] ;
 wire \Tile_X6Y9_N2BEGb[0] ;
 wire \Tile_X6Y9_N2BEGb[1] ;
 wire \Tile_X6Y9_N2BEGb[2] ;
 wire \Tile_X6Y9_N2BEGb[3] ;
 wire \Tile_X6Y9_N2BEGb[4] ;
 wire \Tile_X6Y9_N2BEGb[5] ;
 wire \Tile_X6Y9_N2BEGb[6] ;
 wire \Tile_X6Y9_N2BEGb[7] ;
 wire \Tile_X6Y9_N4BEG[0] ;
 wire \Tile_X6Y9_N4BEG[10] ;
 wire \Tile_X6Y9_N4BEG[11] ;
 wire \Tile_X6Y9_N4BEG[12] ;
 wire \Tile_X6Y9_N4BEG[13] ;
 wire \Tile_X6Y9_N4BEG[14] ;
 wire \Tile_X6Y9_N4BEG[15] ;
 wire \Tile_X6Y9_N4BEG[1] ;
 wire \Tile_X6Y9_N4BEG[2] ;
 wire \Tile_X6Y9_N4BEG[3] ;
 wire \Tile_X6Y9_N4BEG[4] ;
 wire \Tile_X6Y9_N4BEG[5] ;
 wire \Tile_X6Y9_N4BEG[6] ;
 wire \Tile_X6Y9_N4BEG[7] ;
 wire \Tile_X6Y9_N4BEG[8] ;
 wire \Tile_X6Y9_N4BEG[9] ;
 wire \Tile_X6Y9_NN4BEG[0] ;
 wire \Tile_X6Y9_NN4BEG[10] ;
 wire \Tile_X6Y9_NN4BEG[11] ;
 wire \Tile_X6Y9_NN4BEG[12] ;
 wire \Tile_X6Y9_NN4BEG[13] ;
 wire \Tile_X6Y9_NN4BEG[14] ;
 wire \Tile_X6Y9_NN4BEG[15] ;
 wire \Tile_X6Y9_NN4BEG[1] ;
 wire \Tile_X6Y9_NN4BEG[2] ;
 wire \Tile_X6Y9_NN4BEG[3] ;
 wire \Tile_X6Y9_NN4BEG[4] ;
 wire \Tile_X6Y9_NN4BEG[5] ;
 wire \Tile_X6Y9_NN4BEG[6] ;
 wire \Tile_X6Y9_NN4BEG[7] ;
 wire \Tile_X6Y9_NN4BEG[8] ;
 wire \Tile_X6Y9_NN4BEG[9] ;
 wire \Tile_X6Y9_S1BEG[0] ;
 wire \Tile_X6Y9_S1BEG[1] ;
 wire \Tile_X6Y9_S1BEG[2] ;
 wire \Tile_X6Y9_S1BEG[3] ;
 wire \Tile_X6Y9_S2BEG[0] ;
 wire \Tile_X6Y9_S2BEG[1] ;
 wire \Tile_X6Y9_S2BEG[2] ;
 wire \Tile_X6Y9_S2BEG[3] ;
 wire \Tile_X6Y9_S2BEG[4] ;
 wire \Tile_X6Y9_S2BEG[5] ;
 wire \Tile_X6Y9_S2BEG[6] ;
 wire \Tile_X6Y9_S2BEG[7] ;
 wire \Tile_X6Y9_S2BEGb[0] ;
 wire \Tile_X6Y9_S2BEGb[1] ;
 wire \Tile_X6Y9_S2BEGb[2] ;
 wire \Tile_X6Y9_S2BEGb[3] ;
 wire \Tile_X6Y9_S2BEGb[4] ;
 wire \Tile_X6Y9_S2BEGb[5] ;
 wire \Tile_X6Y9_S2BEGb[6] ;
 wire \Tile_X6Y9_S2BEGb[7] ;
 wire \Tile_X6Y9_S4BEG[0] ;
 wire \Tile_X6Y9_S4BEG[10] ;
 wire \Tile_X6Y9_S4BEG[11] ;
 wire \Tile_X6Y9_S4BEG[12] ;
 wire \Tile_X6Y9_S4BEG[13] ;
 wire \Tile_X6Y9_S4BEG[14] ;
 wire \Tile_X6Y9_S4BEG[15] ;
 wire \Tile_X6Y9_S4BEG[1] ;
 wire \Tile_X6Y9_S4BEG[2] ;
 wire \Tile_X6Y9_S4BEG[3] ;
 wire \Tile_X6Y9_S4BEG[4] ;
 wire \Tile_X6Y9_S4BEG[5] ;
 wire \Tile_X6Y9_S4BEG[6] ;
 wire \Tile_X6Y9_S4BEG[7] ;
 wire \Tile_X6Y9_S4BEG[8] ;
 wire \Tile_X6Y9_S4BEG[9] ;
 wire \Tile_X6Y9_SS4BEG[0] ;
 wire \Tile_X6Y9_SS4BEG[10] ;
 wire \Tile_X6Y9_SS4BEG[11] ;
 wire \Tile_X6Y9_SS4BEG[12] ;
 wire \Tile_X6Y9_SS4BEG[13] ;
 wire \Tile_X6Y9_SS4BEG[14] ;
 wire \Tile_X6Y9_SS4BEG[15] ;
 wire \Tile_X6Y9_SS4BEG[1] ;
 wire \Tile_X6Y9_SS4BEG[2] ;
 wire \Tile_X6Y9_SS4BEG[3] ;
 wire \Tile_X6Y9_SS4BEG[4] ;
 wire \Tile_X6Y9_SS4BEG[5] ;
 wire \Tile_X6Y9_SS4BEG[6] ;
 wire \Tile_X6Y9_SS4BEG[7] ;
 wire \Tile_X6Y9_SS4BEG[8] ;
 wire \Tile_X6Y9_SS4BEG[9] ;
 wire Tile_X6Y9_UserCLKo;
 wire \Tile_X6Y9_W1BEG[0] ;
 wire \Tile_X6Y9_W1BEG[1] ;
 wire \Tile_X6Y9_W1BEG[2] ;
 wire \Tile_X6Y9_W1BEG[3] ;
 wire \Tile_X6Y9_W2BEG[0] ;
 wire \Tile_X6Y9_W2BEG[1] ;
 wire \Tile_X6Y9_W2BEG[2] ;
 wire \Tile_X6Y9_W2BEG[3] ;
 wire \Tile_X6Y9_W2BEG[4] ;
 wire \Tile_X6Y9_W2BEG[5] ;
 wire \Tile_X6Y9_W2BEG[6] ;
 wire \Tile_X6Y9_W2BEG[7] ;
 wire \Tile_X6Y9_W2BEGb[0] ;
 wire \Tile_X6Y9_W2BEGb[1] ;
 wire \Tile_X6Y9_W2BEGb[2] ;
 wire \Tile_X6Y9_W2BEGb[3] ;
 wire \Tile_X6Y9_W2BEGb[4] ;
 wire \Tile_X6Y9_W2BEGb[5] ;
 wire \Tile_X6Y9_W2BEGb[6] ;
 wire \Tile_X6Y9_W2BEGb[7] ;
 wire \Tile_X6Y9_W6BEG[0] ;
 wire \Tile_X6Y9_W6BEG[10] ;
 wire \Tile_X6Y9_W6BEG[11] ;
 wire \Tile_X6Y9_W6BEG[1] ;
 wire \Tile_X6Y9_W6BEG[2] ;
 wire \Tile_X6Y9_W6BEG[3] ;
 wire \Tile_X6Y9_W6BEG[4] ;
 wire \Tile_X6Y9_W6BEG[5] ;
 wire \Tile_X6Y9_W6BEG[6] ;
 wire \Tile_X6Y9_W6BEG[7] ;
 wire \Tile_X6Y9_W6BEG[8] ;
 wire \Tile_X6Y9_W6BEG[9] ;
 wire \Tile_X6Y9_WW4BEG[0] ;
 wire \Tile_X6Y9_WW4BEG[10] ;
 wire \Tile_X6Y9_WW4BEG[11] ;
 wire \Tile_X6Y9_WW4BEG[12] ;
 wire \Tile_X6Y9_WW4BEG[13] ;
 wire \Tile_X6Y9_WW4BEG[14] ;
 wire \Tile_X6Y9_WW4BEG[15] ;
 wire \Tile_X6Y9_WW4BEG[1] ;
 wire \Tile_X6Y9_WW4BEG[2] ;
 wire \Tile_X6Y9_WW4BEG[3] ;
 wire \Tile_X6Y9_WW4BEG[4] ;
 wire \Tile_X6Y9_WW4BEG[5] ;
 wire \Tile_X6Y9_WW4BEG[6] ;
 wire \Tile_X6Y9_WW4BEG[7] ;
 wire \Tile_X6Y9_WW4BEG[8] ;
 wire \Tile_X6Y9_WW4BEG[9] ;
 wire \Tile_X7Y0_FrameData_O[0] ;
 wire \Tile_X7Y0_FrameData_O[10] ;
 wire \Tile_X7Y0_FrameData_O[11] ;
 wire \Tile_X7Y0_FrameData_O[12] ;
 wire \Tile_X7Y0_FrameData_O[13] ;
 wire \Tile_X7Y0_FrameData_O[14] ;
 wire \Tile_X7Y0_FrameData_O[15] ;
 wire \Tile_X7Y0_FrameData_O[16] ;
 wire \Tile_X7Y0_FrameData_O[17] ;
 wire \Tile_X7Y0_FrameData_O[18] ;
 wire \Tile_X7Y0_FrameData_O[19] ;
 wire \Tile_X7Y0_FrameData_O[1] ;
 wire \Tile_X7Y0_FrameData_O[20] ;
 wire \Tile_X7Y0_FrameData_O[21] ;
 wire \Tile_X7Y0_FrameData_O[22] ;
 wire \Tile_X7Y0_FrameData_O[23] ;
 wire \Tile_X7Y0_FrameData_O[24] ;
 wire \Tile_X7Y0_FrameData_O[25] ;
 wire \Tile_X7Y0_FrameData_O[26] ;
 wire \Tile_X7Y0_FrameData_O[27] ;
 wire \Tile_X7Y0_FrameData_O[28] ;
 wire \Tile_X7Y0_FrameData_O[29] ;
 wire \Tile_X7Y0_FrameData_O[2] ;
 wire \Tile_X7Y0_FrameData_O[30] ;
 wire \Tile_X7Y0_FrameData_O[31] ;
 wire \Tile_X7Y0_FrameData_O[3] ;
 wire \Tile_X7Y0_FrameData_O[4] ;
 wire \Tile_X7Y0_FrameData_O[5] ;
 wire \Tile_X7Y0_FrameData_O[6] ;
 wire \Tile_X7Y0_FrameData_O[7] ;
 wire \Tile_X7Y0_FrameData_O[8] ;
 wire \Tile_X7Y0_FrameData_O[9] ;
 wire \Tile_X7Y0_FrameStrobe_O[0] ;
 wire \Tile_X7Y0_FrameStrobe_O[10] ;
 wire \Tile_X7Y0_FrameStrobe_O[11] ;
 wire \Tile_X7Y0_FrameStrobe_O[12] ;
 wire \Tile_X7Y0_FrameStrobe_O[13] ;
 wire \Tile_X7Y0_FrameStrobe_O[14] ;
 wire \Tile_X7Y0_FrameStrobe_O[15] ;
 wire \Tile_X7Y0_FrameStrobe_O[16] ;
 wire \Tile_X7Y0_FrameStrobe_O[17] ;
 wire \Tile_X7Y0_FrameStrobe_O[18] ;
 wire \Tile_X7Y0_FrameStrobe_O[19] ;
 wire \Tile_X7Y0_FrameStrobe_O[1] ;
 wire \Tile_X7Y0_FrameStrobe_O[2] ;
 wire \Tile_X7Y0_FrameStrobe_O[3] ;
 wire \Tile_X7Y0_FrameStrobe_O[4] ;
 wire \Tile_X7Y0_FrameStrobe_O[5] ;
 wire \Tile_X7Y0_FrameStrobe_O[6] ;
 wire \Tile_X7Y0_FrameStrobe_O[7] ;
 wire \Tile_X7Y0_FrameStrobe_O[8] ;
 wire \Tile_X7Y0_FrameStrobe_O[9] ;
 wire \Tile_X7Y0_S1BEG[0] ;
 wire \Tile_X7Y0_S1BEG[1] ;
 wire \Tile_X7Y0_S1BEG[2] ;
 wire \Tile_X7Y0_S1BEG[3] ;
 wire \Tile_X7Y0_S2BEG[0] ;
 wire \Tile_X7Y0_S2BEG[1] ;
 wire \Tile_X7Y0_S2BEG[2] ;
 wire \Tile_X7Y0_S2BEG[3] ;
 wire \Tile_X7Y0_S2BEG[4] ;
 wire \Tile_X7Y0_S2BEG[5] ;
 wire \Tile_X7Y0_S2BEG[6] ;
 wire \Tile_X7Y0_S2BEG[7] ;
 wire \Tile_X7Y0_S2BEGb[0] ;
 wire \Tile_X7Y0_S2BEGb[1] ;
 wire \Tile_X7Y0_S2BEGb[2] ;
 wire \Tile_X7Y0_S2BEGb[3] ;
 wire \Tile_X7Y0_S2BEGb[4] ;
 wire \Tile_X7Y0_S2BEGb[5] ;
 wire \Tile_X7Y0_S2BEGb[6] ;
 wire \Tile_X7Y0_S2BEGb[7] ;
 wire \Tile_X7Y0_S4BEG[0] ;
 wire \Tile_X7Y0_S4BEG[10] ;
 wire \Tile_X7Y0_S4BEG[11] ;
 wire \Tile_X7Y0_S4BEG[12] ;
 wire \Tile_X7Y0_S4BEG[13] ;
 wire \Tile_X7Y0_S4BEG[14] ;
 wire \Tile_X7Y0_S4BEG[15] ;
 wire \Tile_X7Y0_S4BEG[1] ;
 wire \Tile_X7Y0_S4BEG[2] ;
 wire \Tile_X7Y0_S4BEG[3] ;
 wire \Tile_X7Y0_S4BEG[4] ;
 wire \Tile_X7Y0_S4BEG[5] ;
 wire \Tile_X7Y0_S4BEG[6] ;
 wire \Tile_X7Y0_S4BEG[7] ;
 wire \Tile_X7Y0_S4BEG[8] ;
 wire \Tile_X7Y0_S4BEG[9] ;
 wire \Tile_X7Y0_SS4BEG[0] ;
 wire \Tile_X7Y0_SS4BEG[10] ;
 wire \Tile_X7Y0_SS4BEG[11] ;
 wire \Tile_X7Y0_SS4BEG[12] ;
 wire \Tile_X7Y0_SS4BEG[13] ;
 wire \Tile_X7Y0_SS4BEG[14] ;
 wire \Tile_X7Y0_SS4BEG[15] ;
 wire \Tile_X7Y0_SS4BEG[1] ;
 wire \Tile_X7Y0_SS4BEG[2] ;
 wire \Tile_X7Y0_SS4BEG[3] ;
 wire \Tile_X7Y0_SS4BEG[4] ;
 wire \Tile_X7Y0_SS4BEG[5] ;
 wire \Tile_X7Y0_SS4BEG[6] ;
 wire \Tile_X7Y0_SS4BEG[7] ;
 wire \Tile_X7Y0_SS4BEG[8] ;
 wire \Tile_X7Y0_SS4BEG[9] ;
 wire Tile_X7Y0_UserCLKo;
 wire \Tile_X7Y10_E1BEG[0] ;
 wire \Tile_X7Y10_E1BEG[1] ;
 wire \Tile_X7Y10_E1BEG[2] ;
 wire \Tile_X7Y10_E1BEG[3] ;
 wire \Tile_X7Y10_E2BEG[0] ;
 wire \Tile_X7Y10_E2BEG[1] ;
 wire \Tile_X7Y10_E2BEG[2] ;
 wire \Tile_X7Y10_E2BEG[3] ;
 wire \Tile_X7Y10_E2BEG[4] ;
 wire \Tile_X7Y10_E2BEG[5] ;
 wire \Tile_X7Y10_E2BEG[6] ;
 wire \Tile_X7Y10_E2BEG[7] ;
 wire \Tile_X7Y10_E2BEGb[0] ;
 wire \Tile_X7Y10_E2BEGb[1] ;
 wire \Tile_X7Y10_E2BEGb[2] ;
 wire \Tile_X7Y10_E2BEGb[3] ;
 wire \Tile_X7Y10_E2BEGb[4] ;
 wire \Tile_X7Y10_E2BEGb[5] ;
 wire \Tile_X7Y10_E2BEGb[6] ;
 wire \Tile_X7Y10_E2BEGb[7] ;
 wire \Tile_X7Y10_E6BEG[0] ;
 wire \Tile_X7Y10_E6BEG[10] ;
 wire \Tile_X7Y10_E6BEG[11] ;
 wire \Tile_X7Y10_E6BEG[1] ;
 wire \Tile_X7Y10_E6BEG[2] ;
 wire \Tile_X7Y10_E6BEG[3] ;
 wire \Tile_X7Y10_E6BEG[4] ;
 wire \Tile_X7Y10_E6BEG[5] ;
 wire \Tile_X7Y10_E6BEG[6] ;
 wire \Tile_X7Y10_E6BEG[7] ;
 wire \Tile_X7Y10_E6BEG[8] ;
 wire \Tile_X7Y10_E6BEG[9] ;
 wire \Tile_X7Y10_EE4BEG[0] ;
 wire \Tile_X7Y10_EE4BEG[10] ;
 wire \Tile_X7Y10_EE4BEG[11] ;
 wire \Tile_X7Y10_EE4BEG[12] ;
 wire \Tile_X7Y10_EE4BEG[13] ;
 wire \Tile_X7Y10_EE4BEG[14] ;
 wire \Tile_X7Y10_EE4BEG[15] ;
 wire \Tile_X7Y10_EE4BEG[1] ;
 wire \Tile_X7Y10_EE4BEG[2] ;
 wire \Tile_X7Y10_EE4BEG[3] ;
 wire \Tile_X7Y10_EE4BEG[4] ;
 wire \Tile_X7Y10_EE4BEG[5] ;
 wire \Tile_X7Y10_EE4BEG[6] ;
 wire \Tile_X7Y10_EE4BEG[7] ;
 wire \Tile_X7Y10_EE4BEG[8] ;
 wire \Tile_X7Y10_EE4BEG[9] ;
 wire \Tile_X7Y10_FrameData_O[0] ;
 wire \Tile_X7Y10_FrameData_O[10] ;
 wire \Tile_X7Y10_FrameData_O[11] ;
 wire \Tile_X7Y10_FrameData_O[12] ;
 wire \Tile_X7Y10_FrameData_O[13] ;
 wire \Tile_X7Y10_FrameData_O[14] ;
 wire \Tile_X7Y10_FrameData_O[15] ;
 wire \Tile_X7Y10_FrameData_O[16] ;
 wire \Tile_X7Y10_FrameData_O[17] ;
 wire \Tile_X7Y10_FrameData_O[18] ;
 wire \Tile_X7Y10_FrameData_O[19] ;
 wire \Tile_X7Y10_FrameData_O[1] ;
 wire \Tile_X7Y10_FrameData_O[20] ;
 wire \Tile_X7Y10_FrameData_O[21] ;
 wire \Tile_X7Y10_FrameData_O[22] ;
 wire \Tile_X7Y10_FrameData_O[23] ;
 wire \Tile_X7Y10_FrameData_O[24] ;
 wire \Tile_X7Y10_FrameData_O[25] ;
 wire \Tile_X7Y10_FrameData_O[26] ;
 wire \Tile_X7Y10_FrameData_O[27] ;
 wire \Tile_X7Y10_FrameData_O[28] ;
 wire \Tile_X7Y10_FrameData_O[29] ;
 wire \Tile_X7Y10_FrameData_O[2] ;
 wire \Tile_X7Y10_FrameData_O[30] ;
 wire \Tile_X7Y10_FrameData_O[31] ;
 wire \Tile_X7Y10_FrameData_O[3] ;
 wire \Tile_X7Y10_FrameData_O[4] ;
 wire \Tile_X7Y10_FrameData_O[5] ;
 wire \Tile_X7Y10_FrameData_O[6] ;
 wire \Tile_X7Y10_FrameData_O[7] ;
 wire \Tile_X7Y10_FrameData_O[8] ;
 wire \Tile_X7Y10_FrameData_O[9] ;
 wire \Tile_X7Y10_S1BEG[0] ;
 wire \Tile_X7Y10_S1BEG[1] ;
 wire \Tile_X7Y10_S1BEG[2] ;
 wire \Tile_X7Y10_S1BEG[3] ;
 wire \Tile_X7Y10_S2BEG[0] ;
 wire \Tile_X7Y10_S2BEG[1] ;
 wire \Tile_X7Y10_S2BEG[2] ;
 wire \Tile_X7Y10_S2BEG[3] ;
 wire \Tile_X7Y10_S2BEG[4] ;
 wire \Tile_X7Y10_S2BEG[5] ;
 wire \Tile_X7Y10_S2BEG[6] ;
 wire \Tile_X7Y10_S2BEG[7] ;
 wire \Tile_X7Y10_S2BEGb[0] ;
 wire \Tile_X7Y10_S2BEGb[1] ;
 wire \Tile_X7Y10_S2BEGb[2] ;
 wire \Tile_X7Y10_S2BEGb[3] ;
 wire \Tile_X7Y10_S2BEGb[4] ;
 wire \Tile_X7Y10_S2BEGb[5] ;
 wire \Tile_X7Y10_S2BEGb[6] ;
 wire \Tile_X7Y10_S2BEGb[7] ;
 wire \Tile_X7Y10_S4BEG[0] ;
 wire \Tile_X7Y10_S4BEG[10] ;
 wire \Tile_X7Y10_S4BEG[11] ;
 wire \Tile_X7Y10_S4BEG[12] ;
 wire \Tile_X7Y10_S4BEG[13] ;
 wire \Tile_X7Y10_S4BEG[14] ;
 wire \Tile_X7Y10_S4BEG[15] ;
 wire \Tile_X7Y10_S4BEG[1] ;
 wire \Tile_X7Y10_S4BEG[2] ;
 wire \Tile_X7Y10_S4BEG[3] ;
 wire \Tile_X7Y10_S4BEG[4] ;
 wire \Tile_X7Y10_S4BEG[5] ;
 wire \Tile_X7Y10_S4BEG[6] ;
 wire \Tile_X7Y10_S4BEG[7] ;
 wire \Tile_X7Y10_S4BEG[8] ;
 wire \Tile_X7Y10_S4BEG[9] ;
 wire \Tile_X7Y10_SS4BEG[0] ;
 wire \Tile_X7Y10_SS4BEG[10] ;
 wire \Tile_X7Y10_SS4BEG[11] ;
 wire \Tile_X7Y10_SS4BEG[12] ;
 wire \Tile_X7Y10_SS4BEG[13] ;
 wire \Tile_X7Y10_SS4BEG[14] ;
 wire \Tile_X7Y10_SS4BEG[15] ;
 wire \Tile_X7Y10_SS4BEG[1] ;
 wire \Tile_X7Y10_SS4BEG[2] ;
 wire \Tile_X7Y10_SS4BEG[3] ;
 wire \Tile_X7Y10_SS4BEG[4] ;
 wire \Tile_X7Y10_SS4BEG[5] ;
 wire \Tile_X7Y10_SS4BEG[6] ;
 wire \Tile_X7Y10_SS4BEG[7] ;
 wire \Tile_X7Y10_SS4BEG[8] ;
 wire \Tile_X7Y10_SS4BEG[9] ;
 wire \Tile_X7Y10_W1BEG[0] ;
 wire \Tile_X7Y10_W1BEG[1] ;
 wire \Tile_X7Y10_W1BEG[2] ;
 wire \Tile_X7Y10_W1BEG[3] ;
 wire \Tile_X7Y10_W2BEG[0] ;
 wire \Tile_X7Y10_W2BEG[1] ;
 wire \Tile_X7Y10_W2BEG[2] ;
 wire \Tile_X7Y10_W2BEG[3] ;
 wire \Tile_X7Y10_W2BEG[4] ;
 wire \Tile_X7Y10_W2BEG[5] ;
 wire \Tile_X7Y10_W2BEG[6] ;
 wire \Tile_X7Y10_W2BEG[7] ;
 wire \Tile_X7Y10_W2BEGb[0] ;
 wire \Tile_X7Y10_W2BEGb[1] ;
 wire \Tile_X7Y10_W2BEGb[2] ;
 wire \Tile_X7Y10_W2BEGb[3] ;
 wire \Tile_X7Y10_W2BEGb[4] ;
 wire \Tile_X7Y10_W2BEGb[5] ;
 wire \Tile_X7Y10_W2BEGb[6] ;
 wire \Tile_X7Y10_W2BEGb[7] ;
 wire \Tile_X7Y10_W6BEG[0] ;
 wire \Tile_X7Y10_W6BEG[10] ;
 wire \Tile_X7Y10_W6BEG[11] ;
 wire \Tile_X7Y10_W6BEG[1] ;
 wire \Tile_X7Y10_W6BEG[2] ;
 wire \Tile_X7Y10_W6BEG[3] ;
 wire \Tile_X7Y10_W6BEG[4] ;
 wire \Tile_X7Y10_W6BEG[5] ;
 wire \Tile_X7Y10_W6BEG[6] ;
 wire \Tile_X7Y10_W6BEG[7] ;
 wire \Tile_X7Y10_W6BEG[8] ;
 wire \Tile_X7Y10_W6BEG[9] ;
 wire \Tile_X7Y10_WW4BEG[0] ;
 wire \Tile_X7Y10_WW4BEG[10] ;
 wire \Tile_X7Y10_WW4BEG[11] ;
 wire \Tile_X7Y10_WW4BEG[12] ;
 wire \Tile_X7Y10_WW4BEG[13] ;
 wire \Tile_X7Y10_WW4BEG[14] ;
 wire \Tile_X7Y10_WW4BEG[15] ;
 wire \Tile_X7Y10_WW4BEG[1] ;
 wire \Tile_X7Y10_WW4BEG[2] ;
 wire \Tile_X7Y10_WW4BEG[3] ;
 wire \Tile_X7Y10_WW4BEG[4] ;
 wire \Tile_X7Y10_WW4BEG[5] ;
 wire \Tile_X7Y10_WW4BEG[6] ;
 wire \Tile_X7Y10_WW4BEG[7] ;
 wire \Tile_X7Y10_WW4BEG[8] ;
 wire \Tile_X7Y10_WW4BEG[9] ;
 wire \Tile_X7Y11_E1BEG[0] ;
 wire \Tile_X7Y11_E1BEG[1] ;
 wire \Tile_X7Y11_E1BEG[2] ;
 wire \Tile_X7Y11_E1BEG[3] ;
 wire \Tile_X7Y11_E2BEG[0] ;
 wire \Tile_X7Y11_E2BEG[1] ;
 wire \Tile_X7Y11_E2BEG[2] ;
 wire \Tile_X7Y11_E2BEG[3] ;
 wire \Tile_X7Y11_E2BEG[4] ;
 wire \Tile_X7Y11_E2BEG[5] ;
 wire \Tile_X7Y11_E2BEG[6] ;
 wire \Tile_X7Y11_E2BEG[7] ;
 wire \Tile_X7Y11_E2BEGb[0] ;
 wire \Tile_X7Y11_E2BEGb[1] ;
 wire \Tile_X7Y11_E2BEGb[2] ;
 wire \Tile_X7Y11_E2BEGb[3] ;
 wire \Tile_X7Y11_E2BEGb[4] ;
 wire \Tile_X7Y11_E2BEGb[5] ;
 wire \Tile_X7Y11_E2BEGb[6] ;
 wire \Tile_X7Y11_E2BEGb[7] ;
 wire \Tile_X7Y11_E6BEG[0] ;
 wire \Tile_X7Y11_E6BEG[10] ;
 wire \Tile_X7Y11_E6BEG[11] ;
 wire \Tile_X7Y11_E6BEG[1] ;
 wire \Tile_X7Y11_E6BEG[2] ;
 wire \Tile_X7Y11_E6BEG[3] ;
 wire \Tile_X7Y11_E6BEG[4] ;
 wire \Tile_X7Y11_E6BEG[5] ;
 wire \Tile_X7Y11_E6BEG[6] ;
 wire \Tile_X7Y11_E6BEG[7] ;
 wire \Tile_X7Y11_E6BEG[8] ;
 wire \Tile_X7Y11_E6BEG[9] ;
 wire \Tile_X7Y11_EE4BEG[0] ;
 wire \Tile_X7Y11_EE4BEG[10] ;
 wire \Tile_X7Y11_EE4BEG[11] ;
 wire \Tile_X7Y11_EE4BEG[12] ;
 wire \Tile_X7Y11_EE4BEG[13] ;
 wire \Tile_X7Y11_EE4BEG[14] ;
 wire \Tile_X7Y11_EE4BEG[15] ;
 wire \Tile_X7Y11_EE4BEG[1] ;
 wire \Tile_X7Y11_EE4BEG[2] ;
 wire \Tile_X7Y11_EE4BEG[3] ;
 wire \Tile_X7Y11_EE4BEG[4] ;
 wire \Tile_X7Y11_EE4BEG[5] ;
 wire \Tile_X7Y11_EE4BEG[6] ;
 wire \Tile_X7Y11_EE4BEG[7] ;
 wire \Tile_X7Y11_EE4BEG[8] ;
 wire \Tile_X7Y11_EE4BEG[9] ;
 wire \Tile_X7Y11_FrameData_O[0] ;
 wire \Tile_X7Y11_FrameData_O[10] ;
 wire \Tile_X7Y11_FrameData_O[11] ;
 wire \Tile_X7Y11_FrameData_O[12] ;
 wire \Tile_X7Y11_FrameData_O[13] ;
 wire \Tile_X7Y11_FrameData_O[14] ;
 wire \Tile_X7Y11_FrameData_O[15] ;
 wire \Tile_X7Y11_FrameData_O[16] ;
 wire \Tile_X7Y11_FrameData_O[17] ;
 wire \Tile_X7Y11_FrameData_O[18] ;
 wire \Tile_X7Y11_FrameData_O[19] ;
 wire \Tile_X7Y11_FrameData_O[1] ;
 wire \Tile_X7Y11_FrameData_O[20] ;
 wire \Tile_X7Y11_FrameData_O[21] ;
 wire \Tile_X7Y11_FrameData_O[22] ;
 wire \Tile_X7Y11_FrameData_O[23] ;
 wire \Tile_X7Y11_FrameData_O[24] ;
 wire \Tile_X7Y11_FrameData_O[25] ;
 wire \Tile_X7Y11_FrameData_O[26] ;
 wire \Tile_X7Y11_FrameData_O[27] ;
 wire \Tile_X7Y11_FrameData_O[28] ;
 wire \Tile_X7Y11_FrameData_O[29] ;
 wire \Tile_X7Y11_FrameData_O[2] ;
 wire \Tile_X7Y11_FrameData_O[30] ;
 wire \Tile_X7Y11_FrameData_O[31] ;
 wire \Tile_X7Y11_FrameData_O[3] ;
 wire \Tile_X7Y11_FrameData_O[4] ;
 wire \Tile_X7Y11_FrameData_O[5] ;
 wire \Tile_X7Y11_FrameData_O[6] ;
 wire \Tile_X7Y11_FrameData_O[7] ;
 wire \Tile_X7Y11_FrameData_O[8] ;
 wire \Tile_X7Y11_FrameData_O[9] ;
 wire \Tile_X7Y11_FrameStrobe_O[0] ;
 wire \Tile_X7Y11_FrameStrobe_O[10] ;
 wire \Tile_X7Y11_FrameStrobe_O[11] ;
 wire \Tile_X7Y11_FrameStrobe_O[12] ;
 wire \Tile_X7Y11_FrameStrobe_O[13] ;
 wire \Tile_X7Y11_FrameStrobe_O[14] ;
 wire \Tile_X7Y11_FrameStrobe_O[15] ;
 wire \Tile_X7Y11_FrameStrobe_O[16] ;
 wire \Tile_X7Y11_FrameStrobe_O[17] ;
 wire \Tile_X7Y11_FrameStrobe_O[18] ;
 wire \Tile_X7Y11_FrameStrobe_O[19] ;
 wire \Tile_X7Y11_FrameStrobe_O[1] ;
 wire \Tile_X7Y11_FrameStrobe_O[2] ;
 wire \Tile_X7Y11_FrameStrobe_O[3] ;
 wire \Tile_X7Y11_FrameStrobe_O[4] ;
 wire \Tile_X7Y11_FrameStrobe_O[5] ;
 wire \Tile_X7Y11_FrameStrobe_O[6] ;
 wire \Tile_X7Y11_FrameStrobe_O[7] ;
 wire \Tile_X7Y11_FrameStrobe_O[8] ;
 wire \Tile_X7Y11_FrameStrobe_O[9] ;
 wire \Tile_X7Y11_N1BEG[0] ;
 wire \Tile_X7Y11_N1BEG[1] ;
 wire \Tile_X7Y11_N1BEG[2] ;
 wire \Tile_X7Y11_N1BEG[3] ;
 wire \Tile_X7Y11_N2BEG[0] ;
 wire \Tile_X7Y11_N2BEG[1] ;
 wire \Tile_X7Y11_N2BEG[2] ;
 wire \Tile_X7Y11_N2BEG[3] ;
 wire \Tile_X7Y11_N2BEG[4] ;
 wire \Tile_X7Y11_N2BEG[5] ;
 wire \Tile_X7Y11_N2BEG[6] ;
 wire \Tile_X7Y11_N2BEG[7] ;
 wire \Tile_X7Y11_N2BEGb[0] ;
 wire \Tile_X7Y11_N2BEGb[1] ;
 wire \Tile_X7Y11_N2BEGb[2] ;
 wire \Tile_X7Y11_N2BEGb[3] ;
 wire \Tile_X7Y11_N2BEGb[4] ;
 wire \Tile_X7Y11_N2BEGb[5] ;
 wire \Tile_X7Y11_N2BEGb[6] ;
 wire \Tile_X7Y11_N2BEGb[7] ;
 wire \Tile_X7Y11_N4BEG[0] ;
 wire \Tile_X7Y11_N4BEG[10] ;
 wire \Tile_X7Y11_N4BEG[11] ;
 wire \Tile_X7Y11_N4BEG[12] ;
 wire \Tile_X7Y11_N4BEG[13] ;
 wire \Tile_X7Y11_N4BEG[14] ;
 wire \Tile_X7Y11_N4BEG[15] ;
 wire \Tile_X7Y11_N4BEG[1] ;
 wire \Tile_X7Y11_N4BEG[2] ;
 wire \Tile_X7Y11_N4BEG[3] ;
 wire \Tile_X7Y11_N4BEG[4] ;
 wire \Tile_X7Y11_N4BEG[5] ;
 wire \Tile_X7Y11_N4BEG[6] ;
 wire \Tile_X7Y11_N4BEG[7] ;
 wire \Tile_X7Y11_N4BEG[8] ;
 wire \Tile_X7Y11_N4BEG[9] ;
 wire \Tile_X7Y11_NN4BEG[0] ;
 wire \Tile_X7Y11_NN4BEG[10] ;
 wire \Tile_X7Y11_NN4BEG[11] ;
 wire \Tile_X7Y11_NN4BEG[12] ;
 wire \Tile_X7Y11_NN4BEG[13] ;
 wire \Tile_X7Y11_NN4BEG[14] ;
 wire \Tile_X7Y11_NN4BEG[15] ;
 wire \Tile_X7Y11_NN4BEG[1] ;
 wire \Tile_X7Y11_NN4BEG[2] ;
 wire \Tile_X7Y11_NN4BEG[3] ;
 wire \Tile_X7Y11_NN4BEG[4] ;
 wire \Tile_X7Y11_NN4BEG[5] ;
 wire \Tile_X7Y11_NN4BEG[6] ;
 wire \Tile_X7Y11_NN4BEG[7] ;
 wire \Tile_X7Y11_NN4BEG[8] ;
 wire \Tile_X7Y11_NN4BEG[9] ;
 wire Tile_X7Y11_UserCLKo;
 wire \Tile_X7Y11_W1BEG[0] ;
 wire \Tile_X7Y11_W1BEG[1] ;
 wire \Tile_X7Y11_W1BEG[2] ;
 wire \Tile_X7Y11_W1BEG[3] ;
 wire \Tile_X7Y11_W2BEG[0] ;
 wire \Tile_X7Y11_W2BEG[1] ;
 wire \Tile_X7Y11_W2BEG[2] ;
 wire \Tile_X7Y11_W2BEG[3] ;
 wire \Tile_X7Y11_W2BEG[4] ;
 wire \Tile_X7Y11_W2BEG[5] ;
 wire \Tile_X7Y11_W2BEG[6] ;
 wire \Tile_X7Y11_W2BEG[7] ;
 wire \Tile_X7Y11_W2BEGb[0] ;
 wire \Tile_X7Y11_W2BEGb[1] ;
 wire \Tile_X7Y11_W2BEGb[2] ;
 wire \Tile_X7Y11_W2BEGb[3] ;
 wire \Tile_X7Y11_W2BEGb[4] ;
 wire \Tile_X7Y11_W2BEGb[5] ;
 wire \Tile_X7Y11_W2BEGb[6] ;
 wire \Tile_X7Y11_W2BEGb[7] ;
 wire \Tile_X7Y11_W6BEG[0] ;
 wire \Tile_X7Y11_W6BEG[10] ;
 wire \Tile_X7Y11_W6BEG[11] ;
 wire \Tile_X7Y11_W6BEG[1] ;
 wire \Tile_X7Y11_W6BEG[2] ;
 wire \Tile_X7Y11_W6BEG[3] ;
 wire \Tile_X7Y11_W6BEG[4] ;
 wire \Tile_X7Y11_W6BEG[5] ;
 wire \Tile_X7Y11_W6BEG[6] ;
 wire \Tile_X7Y11_W6BEG[7] ;
 wire \Tile_X7Y11_W6BEG[8] ;
 wire \Tile_X7Y11_W6BEG[9] ;
 wire \Tile_X7Y11_WW4BEG[0] ;
 wire \Tile_X7Y11_WW4BEG[10] ;
 wire \Tile_X7Y11_WW4BEG[11] ;
 wire \Tile_X7Y11_WW4BEG[12] ;
 wire \Tile_X7Y11_WW4BEG[13] ;
 wire \Tile_X7Y11_WW4BEG[14] ;
 wire \Tile_X7Y11_WW4BEG[15] ;
 wire \Tile_X7Y11_WW4BEG[1] ;
 wire \Tile_X7Y11_WW4BEG[2] ;
 wire \Tile_X7Y11_WW4BEG[3] ;
 wire \Tile_X7Y11_WW4BEG[4] ;
 wire \Tile_X7Y11_WW4BEG[5] ;
 wire \Tile_X7Y11_WW4BEG[6] ;
 wire \Tile_X7Y11_WW4BEG[7] ;
 wire \Tile_X7Y11_WW4BEG[8] ;
 wire \Tile_X7Y11_WW4BEG[9] ;
 wire \Tile_X7Y12_E1BEG[0] ;
 wire \Tile_X7Y12_E1BEG[1] ;
 wire \Tile_X7Y12_E1BEG[2] ;
 wire \Tile_X7Y12_E1BEG[3] ;
 wire \Tile_X7Y12_E2BEG[0] ;
 wire \Tile_X7Y12_E2BEG[1] ;
 wire \Tile_X7Y12_E2BEG[2] ;
 wire \Tile_X7Y12_E2BEG[3] ;
 wire \Tile_X7Y12_E2BEG[4] ;
 wire \Tile_X7Y12_E2BEG[5] ;
 wire \Tile_X7Y12_E2BEG[6] ;
 wire \Tile_X7Y12_E2BEG[7] ;
 wire \Tile_X7Y12_E2BEGb[0] ;
 wire \Tile_X7Y12_E2BEGb[1] ;
 wire \Tile_X7Y12_E2BEGb[2] ;
 wire \Tile_X7Y12_E2BEGb[3] ;
 wire \Tile_X7Y12_E2BEGb[4] ;
 wire \Tile_X7Y12_E2BEGb[5] ;
 wire \Tile_X7Y12_E2BEGb[6] ;
 wire \Tile_X7Y12_E2BEGb[7] ;
 wire \Tile_X7Y12_E6BEG[0] ;
 wire \Tile_X7Y12_E6BEG[10] ;
 wire \Tile_X7Y12_E6BEG[11] ;
 wire \Tile_X7Y12_E6BEG[1] ;
 wire \Tile_X7Y12_E6BEG[2] ;
 wire \Tile_X7Y12_E6BEG[3] ;
 wire \Tile_X7Y12_E6BEG[4] ;
 wire \Tile_X7Y12_E6BEG[5] ;
 wire \Tile_X7Y12_E6BEG[6] ;
 wire \Tile_X7Y12_E6BEG[7] ;
 wire \Tile_X7Y12_E6BEG[8] ;
 wire \Tile_X7Y12_E6BEG[9] ;
 wire \Tile_X7Y12_EE4BEG[0] ;
 wire \Tile_X7Y12_EE4BEG[10] ;
 wire \Tile_X7Y12_EE4BEG[11] ;
 wire \Tile_X7Y12_EE4BEG[12] ;
 wire \Tile_X7Y12_EE4BEG[13] ;
 wire \Tile_X7Y12_EE4BEG[14] ;
 wire \Tile_X7Y12_EE4BEG[15] ;
 wire \Tile_X7Y12_EE4BEG[1] ;
 wire \Tile_X7Y12_EE4BEG[2] ;
 wire \Tile_X7Y12_EE4BEG[3] ;
 wire \Tile_X7Y12_EE4BEG[4] ;
 wire \Tile_X7Y12_EE4BEG[5] ;
 wire \Tile_X7Y12_EE4BEG[6] ;
 wire \Tile_X7Y12_EE4BEG[7] ;
 wire \Tile_X7Y12_EE4BEG[8] ;
 wire \Tile_X7Y12_EE4BEG[9] ;
 wire \Tile_X7Y12_FrameData_O[0] ;
 wire \Tile_X7Y12_FrameData_O[10] ;
 wire \Tile_X7Y12_FrameData_O[11] ;
 wire \Tile_X7Y12_FrameData_O[12] ;
 wire \Tile_X7Y12_FrameData_O[13] ;
 wire \Tile_X7Y12_FrameData_O[14] ;
 wire \Tile_X7Y12_FrameData_O[15] ;
 wire \Tile_X7Y12_FrameData_O[16] ;
 wire \Tile_X7Y12_FrameData_O[17] ;
 wire \Tile_X7Y12_FrameData_O[18] ;
 wire \Tile_X7Y12_FrameData_O[19] ;
 wire \Tile_X7Y12_FrameData_O[1] ;
 wire \Tile_X7Y12_FrameData_O[20] ;
 wire \Tile_X7Y12_FrameData_O[21] ;
 wire \Tile_X7Y12_FrameData_O[22] ;
 wire \Tile_X7Y12_FrameData_O[23] ;
 wire \Tile_X7Y12_FrameData_O[24] ;
 wire \Tile_X7Y12_FrameData_O[25] ;
 wire \Tile_X7Y12_FrameData_O[26] ;
 wire \Tile_X7Y12_FrameData_O[27] ;
 wire \Tile_X7Y12_FrameData_O[28] ;
 wire \Tile_X7Y12_FrameData_O[29] ;
 wire \Tile_X7Y12_FrameData_O[2] ;
 wire \Tile_X7Y12_FrameData_O[30] ;
 wire \Tile_X7Y12_FrameData_O[31] ;
 wire \Tile_X7Y12_FrameData_O[3] ;
 wire \Tile_X7Y12_FrameData_O[4] ;
 wire \Tile_X7Y12_FrameData_O[5] ;
 wire \Tile_X7Y12_FrameData_O[6] ;
 wire \Tile_X7Y12_FrameData_O[7] ;
 wire \Tile_X7Y12_FrameData_O[8] ;
 wire \Tile_X7Y12_FrameData_O[9] ;
 wire \Tile_X7Y12_S1BEG[0] ;
 wire \Tile_X7Y12_S1BEG[1] ;
 wire \Tile_X7Y12_S1BEG[2] ;
 wire \Tile_X7Y12_S1BEG[3] ;
 wire \Tile_X7Y12_S2BEG[0] ;
 wire \Tile_X7Y12_S2BEG[1] ;
 wire \Tile_X7Y12_S2BEG[2] ;
 wire \Tile_X7Y12_S2BEG[3] ;
 wire \Tile_X7Y12_S2BEG[4] ;
 wire \Tile_X7Y12_S2BEG[5] ;
 wire \Tile_X7Y12_S2BEG[6] ;
 wire \Tile_X7Y12_S2BEG[7] ;
 wire \Tile_X7Y12_S2BEGb[0] ;
 wire \Tile_X7Y12_S2BEGb[1] ;
 wire \Tile_X7Y12_S2BEGb[2] ;
 wire \Tile_X7Y12_S2BEGb[3] ;
 wire \Tile_X7Y12_S2BEGb[4] ;
 wire \Tile_X7Y12_S2BEGb[5] ;
 wire \Tile_X7Y12_S2BEGb[6] ;
 wire \Tile_X7Y12_S2BEGb[7] ;
 wire \Tile_X7Y12_S4BEG[0] ;
 wire \Tile_X7Y12_S4BEG[10] ;
 wire \Tile_X7Y12_S4BEG[11] ;
 wire \Tile_X7Y12_S4BEG[12] ;
 wire \Tile_X7Y12_S4BEG[13] ;
 wire \Tile_X7Y12_S4BEG[14] ;
 wire \Tile_X7Y12_S4BEG[15] ;
 wire \Tile_X7Y12_S4BEG[1] ;
 wire \Tile_X7Y12_S4BEG[2] ;
 wire \Tile_X7Y12_S4BEG[3] ;
 wire \Tile_X7Y12_S4BEG[4] ;
 wire \Tile_X7Y12_S4BEG[5] ;
 wire \Tile_X7Y12_S4BEG[6] ;
 wire \Tile_X7Y12_S4BEG[7] ;
 wire \Tile_X7Y12_S4BEG[8] ;
 wire \Tile_X7Y12_S4BEG[9] ;
 wire \Tile_X7Y12_SS4BEG[0] ;
 wire \Tile_X7Y12_SS4BEG[10] ;
 wire \Tile_X7Y12_SS4BEG[11] ;
 wire \Tile_X7Y12_SS4BEG[12] ;
 wire \Tile_X7Y12_SS4BEG[13] ;
 wire \Tile_X7Y12_SS4BEG[14] ;
 wire \Tile_X7Y12_SS4BEG[15] ;
 wire \Tile_X7Y12_SS4BEG[1] ;
 wire \Tile_X7Y12_SS4BEG[2] ;
 wire \Tile_X7Y12_SS4BEG[3] ;
 wire \Tile_X7Y12_SS4BEG[4] ;
 wire \Tile_X7Y12_SS4BEG[5] ;
 wire \Tile_X7Y12_SS4BEG[6] ;
 wire \Tile_X7Y12_SS4BEG[7] ;
 wire \Tile_X7Y12_SS4BEG[8] ;
 wire \Tile_X7Y12_SS4BEG[9] ;
 wire \Tile_X7Y12_W1BEG[0] ;
 wire \Tile_X7Y12_W1BEG[1] ;
 wire \Tile_X7Y12_W1BEG[2] ;
 wire \Tile_X7Y12_W1BEG[3] ;
 wire \Tile_X7Y12_W2BEG[0] ;
 wire \Tile_X7Y12_W2BEG[1] ;
 wire \Tile_X7Y12_W2BEG[2] ;
 wire \Tile_X7Y12_W2BEG[3] ;
 wire \Tile_X7Y12_W2BEG[4] ;
 wire \Tile_X7Y12_W2BEG[5] ;
 wire \Tile_X7Y12_W2BEG[6] ;
 wire \Tile_X7Y12_W2BEG[7] ;
 wire \Tile_X7Y12_W2BEGb[0] ;
 wire \Tile_X7Y12_W2BEGb[1] ;
 wire \Tile_X7Y12_W2BEGb[2] ;
 wire \Tile_X7Y12_W2BEGb[3] ;
 wire \Tile_X7Y12_W2BEGb[4] ;
 wire \Tile_X7Y12_W2BEGb[5] ;
 wire \Tile_X7Y12_W2BEGb[6] ;
 wire \Tile_X7Y12_W2BEGb[7] ;
 wire \Tile_X7Y12_W6BEG[0] ;
 wire \Tile_X7Y12_W6BEG[10] ;
 wire \Tile_X7Y12_W6BEG[11] ;
 wire \Tile_X7Y12_W6BEG[1] ;
 wire \Tile_X7Y12_W6BEG[2] ;
 wire \Tile_X7Y12_W6BEG[3] ;
 wire \Tile_X7Y12_W6BEG[4] ;
 wire \Tile_X7Y12_W6BEG[5] ;
 wire \Tile_X7Y12_W6BEG[6] ;
 wire \Tile_X7Y12_W6BEG[7] ;
 wire \Tile_X7Y12_W6BEG[8] ;
 wire \Tile_X7Y12_W6BEG[9] ;
 wire \Tile_X7Y12_WW4BEG[0] ;
 wire \Tile_X7Y12_WW4BEG[10] ;
 wire \Tile_X7Y12_WW4BEG[11] ;
 wire \Tile_X7Y12_WW4BEG[12] ;
 wire \Tile_X7Y12_WW4BEG[13] ;
 wire \Tile_X7Y12_WW4BEG[14] ;
 wire \Tile_X7Y12_WW4BEG[15] ;
 wire \Tile_X7Y12_WW4BEG[1] ;
 wire \Tile_X7Y12_WW4BEG[2] ;
 wire \Tile_X7Y12_WW4BEG[3] ;
 wire \Tile_X7Y12_WW4BEG[4] ;
 wire \Tile_X7Y12_WW4BEG[5] ;
 wire \Tile_X7Y12_WW4BEG[6] ;
 wire \Tile_X7Y12_WW4BEG[7] ;
 wire \Tile_X7Y12_WW4BEG[8] ;
 wire \Tile_X7Y12_WW4BEG[9] ;
 wire \Tile_X7Y13_E1BEG[0] ;
 wire \Tile_X7Y13_E1BEG[1] ;
 wire \Tile_X7Y13_E1BEG[2] ;
 wire \Tile_X7Y13_E1BEG[3] ;
 wire \Tile_X7Y13_E2BEG[0] ;
 wire \Tile_X7Y13_E2BEG[1] ;
 wire \Tile_X7Y13_E2BEG[2] ;
 wire \Tile_X7Y13_E2BEG[3] ;
 wire \Tile_X7Y13_E2BEG[4] ;
 wire \Tile_X7Y13_E2BEG[5] ;
 wire \Tile_X7Y13_E2BEG[6] ;
 wire \Tile_X7Y13_E2BEG[7] ;
 wire \Tile_X7Y13_E2BEGb[0] ;
 wire \Tile_X7Y13_E2BEGb[1] ;
 wire \Tile_X7Y13_E2BEGb[2] ;
 wire \Tile_X7Y13_E2BEGb[3] ;
 wire \Tile_X7Y13_E2BEGb[4] ;
 wire \Tile_X7Y13_E2BEGb[5] ;
 wire \Tile_X7Y13_E2BEGb[6] ;
 wire \Tile_X7Y13_E2BEGb[7] ;
 wire \Tile_X7Y13_E6BEG[0] ;
 wire \Tile_X7Y13_E6BEG[10] ;
 wire \Tile_X7Y13_E6BEG[11] ;
 wire \Tile_X7Y13_E6BEG[1] ;
 wire \Tile_X7Y13_E6BEG[2] ;
 wire \Tile_X7Y13_E6BEG[3] ;
 wire \Tile_X7Y13_E6BEG[4] ;
 wire \Tile_X7Y13_E6BEG[5] ;
 wire \Tile_X7Y13_E6BEG[6] ;
 wire \Tile_X7Y13_E6BEG[7] ;
 wire \Tile_X7Y13_E6BEG[8] ;
 wire \Tile_X7Y13_E6BEG[9] ;
 wire \Tile_X7Y13_EE4BEG[0] ;
 wire \Tile_X7Y13_EE4BEG[10] ;
 wire \Tile_X7Y13_EE4BEG[11] ;
 wire \Tile_X7Y13_EE4BEG[12] ;
 wire \Tile_X7Y13_EE4BEG[13] ;
 wire \Tile_X7Y13_EE4BEG[14] ;
 wire \Tile_X7Y13_EE4BEG[15] ;
 wire \Tile_X7Y13_EE4BEG[1] ;
 wire \Tile_X7Y13_EE4BEG[2] ;
 wire \Tile_X7Y13_EE4BEG[3] ;
 wire \Tile_X7Y13_EE4BEG[4] ;
 wire \Tile_X7Y13_EE4BEG[5] ;
 wire \Tile_X7Y13_EE4BEG[6] ;
 wire \Tile_X7Y13_EE4BEG[7] ;
 wire \Tile_X7Y13_EE4BEG[8] ;
 wire \Tile_X7Y13_EE4BEG[9] ;
 wire \Tile_X7Y13_FrameData_O[0] ;
 wire \Tile_X7Y13_FrameData_O[10] ;
 wire \Tile_X7Y13_FrameData_O[11] ;
 wire \Tile_X7Y13_FrameData_O[12] ;
 wire \Tile_X7Y13_FrameData_O[13] ;
 wire \Tile_X7Y13_FrameData_O[14] ;
 wire \Tile_X7Y13_FrameData_O[15] ;
 wire \Tile_X7Y13_FrameData_O[16] ;
 wire \Tile_X7Y13_FrameData_O[17] ;
 wire \Tile_X7Y13_FrameData_O[18] ;
 wire \Tile_X7Y13_FrameData_O[19] ;
 wire \Tile_X7Y13_FrameData_O[1] ;
 wire \Tile_X7Y13_FrameData_O[20] ;
 wire \Tile_X7Y13_FrameData_O[21] ;
 wire \Tile_X7Y13_FrameData_O[22] ;
 wire \Tile_X7Y13_FrameData_O[23] ;
 wire \Tile_X7Y13_FrameData_O[24] ;
 wire \Tile_X7Y13_FrameData_O[25] ;
 wire \Tile_X7Y13_FrameData_O[26] ;
 wire \Tile_X7Y13_FrameData_O[27] ;
 wire \Tile_X7Y13_FrameData_O[28] ;
 wire \Tile_X7Y13_FrameData_O[29] ;
 wire \Tile_X7Y13_FrameData_O[2] ;
 wire \Tile_X7Y13_FrameData_O[30] ;
 wire \Tile_X7Y13_FrameData_O[31] ;
 wire \Tile_X7Y13_FrameData_O[3] ;
 wire \Tile_X7Y13_FrameData_O[4] ;
 wire \Tile_X7Y13_FrameData_O[5] ;
 wire \Tile_X7Y13_FrameData_O[6] ;
 wire \Tile_X7Y13_FrameData_O[7] ;
 wire \Tile_X7Y13_FrameData_O[8] ;
 wire \Tile_X7Y13_FrameData_O[9] ;
 wire \Tile_X7Y13_FrameStrobe_O[0] ;
 wire \Tile_X7Y13_FrameStrobe_O[10] ;
 wire \Tile_X7Y13_FrameStrobe_O[11] ;
 wire \Tile_X7Y13_FrameStrobe_O[12] ;
 wire \Tile_X7Y13_FrameStrobe_O[13] ;
 wire \Tile_X7Y13_FrameStrobe_O[14] ;
 wire \Tile_X7Y13_FrameStrobe_O[15] ;
 wire \Tile_X7Y13_FrameStrobe_O[16] ;
 wire \Tile_X7Y13_FrameStrobe_O[17] ;
 wire \Tile_X7Y13_FrameStrobe_O[18] ;
 wire \Tile_X7Y13_FrameStrobe_O[19] ;
 wire \Tile_X7Y13_FrameStrobe_O[1] ;
 wire \Tile_X7Y13_FrameStrobe_O[2] ;
 wire \Tile_X7Y13_FrameStrobe_O[3] ;
 wire \Tile_X7Y13_FrameStrobe_O[4] ;
 wire \Tile_X7Y13_FrameStrobe_O[5] ;
 wire \Tile_X7Y13_FrameStrobe_O[6] ;
 wire \Tile_X7Y13_FrameStrobe_O[7] ;
 wire \Tile_X7Y13_FrameStrobe_O[8] ;
 wire \Tile_X7Y13_FrameStrobe_O[9] ;
 wire \Tile_X7Y13_N1BEG[0] ;
 wire \Tile_X7Y13_N1BEG[1] ;
 wire \Tile_X7Y13_N1BEG[2] ;
 wire \Tile_X7Y13_N1BEG[3] ;
 wire \Tile_X7Y13_N2BEG[0] ;
 wire \Tile_X7Y13_N2BEG[1] ;
 wire \Tile_X7Y13_N2BEG[2] ;
 wire \Tile_X7Y13_N2BEG[3] ;
 wire \Tile_X7Y13_N2BEG[4] ;
 wire \Tile_X7Y13_N2BEG[5] ;
 wire \Tile_X7Y13_N2BEG[6] ;
 wire \Tile_X7Y13_N2BEG[7] ;
 wire \Tile_X7Y13_N2BEGb[0] ;
 wire \Tile_X7Y13_N2BEGb[1] ;
 wire \Tile_X7Y13_N2BEGb[2] ;
 wire \Tile_X7Y13_N2BEGb[3] ;
 wire \Tile_X7Y13_N2BEGb[4] ;
 wire \Tile_X7Y13_N2BEGb[5] ;
 wire \Tile_X7Y13_N2BEGb[6] ;
 wire \Tile_X7Y13_N2BEGb[7] ;
 wire \Tile_X7Y13_N4BEG[0] ;
 wire \Tile_X7Y13_N4BEG[10] ;
 wire \Tile_X7Y13_N4BEG[11] ;
 wire \Tile_X7Y13_N4BEG[12] ;
 wire \Tile_X7Y13_N4BEG[13] ;
 wire \Tile_X7Y13_N4BEG[14] ;
 wire \Tile_X7Y13_N4BEG[15] ;
 wire \Tile_X7Y13_N4BEG[1] ;
 wire \Tile_X7Y13_N4BEG[2] ;
 wire \Tile_X7Y13_N4BEG[3] ;
 wire \Tile_X7Y13_N4BEG[4] ;
 wire \Tile_X7Y13_N4BEG[5] ;
 wire \Tile_X7Y13_N4BEG[6] ;
 wire \Tile_X7Y13_N4BEG[7] ;
 wire \Tile_X7Y13_N4BEG[8] ;
 wire \Tile_X7Y13_N4BEG[9] ;
 wire \Tile_X7Y13_NN4BEG[0] ;
 wire \Tile_X7Y13_NN4BEG[10] ;
 wire \Tile_X7Y13_NN4BEG[11] ;
 wire \Tile_X7Y13_NN4BEG[12] ;
 wire \Tile_X7Y13_NN4BEG[13] ;
 wire \Tile_X7Y13_NN4BEG[14] ;
 wire \Tile_X7Y13_NN4BEG[15] ;
 wire \Tile_X7Y13_NN4BEG[1] ;
 wire \Tile_X7Y13_NN4BEG[2] ;
 wire \Tile_X7Y13_NN4BEG[3] ;
 wire \Tile_X7Y13_NN4BEG[4] ;
 wire \Tile_X7Y13_NN4BEG[5] ;
 wire \Tile_X7Y13_NN4BEG[6] ;
 wire \Tile_X7Y13_NN4BEG[7] ;
 wire \Tile_X7Y13_NN4BEG[8] ;
 wire \Tile_X7Y13_NN4BEG[9] ;
 wire Tile_X7Y13_UserCLKo;
 wire \Tile_X7Y13_W1BEG[0] ;
 wire \Tile_X7Y13_W1BEG[1] ;
 wire \Tile_X7Y13_W1BEG[2] ;
 wire \Tile_X7Y13_W1BEG[3] ;
 wire \Tile_X7Y13_W2BEG[0] ;
 wire \Tile_X7Y13_W2BEG[1] ;
 wire \Tile_X7Y13_W2BEG[2] ;
 wire \Tile_X7Y13_W2BEG[3] ;
 wire \Tile_X7Y13_W2BEG[4] ;
 wire \Tile_X7Y13_W2BEG[5] ;
 wire \Tile_X7Y13_W2BEG[6] ;
 wire \Tile_X7Y13_W2BEG[7] ;
 wire \Tile_X7Y13_W2BEGb[0] ;
 wire \Tile_X7Y13_W2BEGb[1] ;
 wire \Tile_X7Y13_W2BEGb[2] ;
 wire \Tile_X7Y13_W2BEGb[3] ;
 wire \Tile_X7Y13_W2BEGb[4] ;
 wire \Tile_X7Y13_W2BEGb[5] ;
 wire \Tile_X7Y13_W2BEGb[6] ;
 wire \Tile_X7Y13_W2BEGb[7] ;
 wire \Tile_X7Y13_W6BEG[0] ;
 wire \Tile_X7Y13_W6BEG[10] ;
 wire \Tile_X7Y13_W6BEG[11] ;
 wire \Tile_X7Y13_W6BEG[1] ;
 wire \Tile_X7Y13_W6BEG[2] ;
 wire \Tile_X7Y13_W6BEG[3] ;
 wire \Tile_X7Y13_W6BEG[4] ;
 wire \Tile_X7Y13_W6BEG[5] ;
 wire \Tile_X7Y13_W6BEG[6] ;
 wire \Tile_X7Y13_W6BEG[7] ;
 wire \Tile_X7Y13_W6BEG[8] ;
 wire \Tile_X7Y13_W6BEG[9] ;
 wire \Tile_X7Y13_WW4BEG[0] ;
 wire \Tile_X7Y13_WW4BEG[10] ;
 wire \Tile_X7Y13_WW4BEG[11] ;
 wire \Tile_X7Y13_WW4BEG[12] ;
 wire \Tile_X7Y13_WW4BEG[13] ;
 wire \Tile_X7Y13_WW4BEG[14] ;
 wire \Tile_X7Y13_WW4BEG[15] ;
 wire \Tile_X7Y13_WW4BEG[1] ;
 wire \Tile_X7Y13_WW4BEG[2] ;
 wire \Tile_X7Y13_WW4BEG[3] ;
 wire \Tile_X7Y13_WW4BEG[4] ;
 wire \Tile_X7Y13_WW4BEG[5] ;
 wire \Tile_X7Y13_WW4BEG[6] ;
 wire \Tile_X7Y13_WW4BEG[7] ;
 wire \Tile_X7Y13_WW4BEG[8] ;
 wire \Tile_X7Y13_WW4BEG[9] ;
 wire \Tile_X7Y14_E1BEG[0] ;
 wire \Tile_X7Y14_E1BEG[1] ;
 wire \Tile_X7Y14_E1BEG[2] ;
 wire \Tile_X7Y14_E1BEG[3] ;
 wire \Tile_X7Y14_E2BEG[0] ;
 wire \Tile_X7Y14_E2BEG[1] ;
 wire \Tile_X7Y14_E2BEG[2] ;
 wire \Tile_X7Y14_E2BEG[3] ;
 wire \Tile_X7Y14_E2BEG[4] ;
 wire \Tile_X7Y14_E2BEG[5] ;
 wire \Tile_X7Y14_E2BEG[6] ;
 wire \Tile_X7Y14_E2BEG[7] ;
 wire \Tile_X7Y14_E2BEGb[0] ;
 wire \Tile_X7Y14_E2BEGb[1] ;
 wire \Tile_X7Y14_E2BEGb[2] ;
 wire \Tile_X7Y14_E2BEGb[3] ;
 wire \Tile_X7Y14_E2BEGb[4] ;
 wire \Tile_X7Y14_E2BEGb[5] ;
 wire \Tile_X7Y14_E2BEGb[6] ;
 wire \Tile_X7Y14_E2BEGb[7] ;
 wire \Tile_X7Y14_E6BEG[0] ;
 wire \Tile_X7Y14_E6BEG[10] ;
 wire \Tile_X7Y14_E6BEG[11] ;
 wire \Tile_X7Y14_E6BEG[1] ;
 wire \Tile_X7Y14_E6BEG[2] ;
 wire \Tile_X7Y14_E6BEG[3] ;
 wire \Tile_X7Y14_E6BEG[4] ;
 wire \Tile_X7Y14_E6BEG[5] ;
 wire \Tile_X7Y14_E6BEG[6] ;
 wire \Tile_X7Y14_E6BEG[7] ;
 wire \Tile_X7Y14_E6BEG[8] ;
 wire \Tile_X7Y14_E6BEG[9] ;
 wire \Tile_X7Y14_EE4BEG[0] ;
 wire \Tile_X7Y14_EE4BEG[10] ;
 wire \Tile_X7Y14_EE4BEG[11] ;
 wire \Tile_X7Y14_EE4BEG[12] ;
 wire \Tile_X7Y14_EE4BEG[13] ;
 wire \Tile_X7Y14_EE4BEG[14] ;
 wire \Tile_X7Y14_EE4BEG[15] ;
 wire \Tile_X7Y14_EE4BEG[1] ;
 wire \Tile_X7Y14_EE4BEG[2] ;
 wire \Tile_X7Y14_EE4BEG[3] ;
 wire \Tile_X7Y14_EE4BEG[4] ;
 wire \Tile_X7Y14_EE4BEG[5] ;
 wire \Tile_X7Y14_EE4BEG[6] ;
 wire \Tile_X7Y14_EE4BEG[7] ;
 wire \Tile_X7Y14_EE4BEG[8] ;
 wire \Tile_X7Y14_EE4BEG[9] ;
 wire \Tile_X7Y14_FrameData_O[0] ;
 wire \Tile_X7Y14_FrameData_O[10] ;
 wire \Tile_X7Y14_FrameData_O[11] ;
 wire \Tile_X7Y14_FrameData_O[12] ;
 wire \Tile_X7Y14_FrameData_O[13] ;
 wire \Tile_X7Y14_FrameData_O[14] ;
 wire \Tile_X7Y14_FrameData_O[15] ;
 wire \Tile_X7Y14_FrameData_O[16] ;
 wire \Tile_X7Y14_FrameData_O[17] ;
 wire \Tile_X7Y14_FrameData_O[18] ;
 wire \Tile_X7Y14_FrameData_O[19] ;
 wire \Tile_X7Y14_FrameData_O[1] ;
 wire \Tile_X7Y14_FrameData_O[20] ;
 wire \Tile_X7Y14_FrameData_O[21] ;
 wire \Tile_X7Y14_FrameData_O[22] ;
 wire \Tile_X7Y14_FrameData_O[23] ;
 wire \Tile_X7Y14_FrameData_O[24] ;
 wire \Tile_X7Y14_FrameData_O[25] ;
 wire \Tile_X7Y14_FrameData_O[26] ;
 wire \Tile_X7Y14_FrameData_O[27] ;
 wire \Tile_X7Y14_FrameData_O[28] ;
 wire \Tile_X7Y14_FrameData_O[29] ;
 wire \Tile_X7Y14_FrameData_O[2] ;
 wire \Tile_X7Y14_FrameData_O[30] ;
 wire \Tile_X7Y14_FrameData_O[31] ;
 wire \Tile_X7Y14_FrameData_O[3] ;
 wire \Tile_X7Y14_FrameData_O[4] ;
 wire \Tile_X7Y14_FrameData_O[5] ;
 wire \Tile_X7Y14_FrameData_O[6] ;
 wire \Tile_X7Y14_FrameData_O[7] ;
 wire \Tile_X7Y14_FrameData_O[8] ;
 wire \Tile_X7Y14_FrameData_O[9] ;
 wire \Tile_X7Y14_S1BEG[0] ;
 wire \Tile_X7Y14_S1BEG[1] ;
 wire \Tile_X7Y14_S1BEG[2] ;
 wire \Tile_X7Y14_S1BEG[3] ;
 wire \Tile_X7Y14_S2BEG[0] ;
 wire \Tile_X7Y14_S2BEG[1] ;
 wire \Tile_X7Y14_S2BEG[2] ;
 wire \Tile_X7Y14_S2BEG[3] ;
 wire \Tile_X7Y14_S2BEG[4] ;
 wire \Tile_X7Y14_S2BEG[5] ;
 wire \Tile_X7Y14_S2BEG[6] ;
 wire \Tile_X7Y14_S2BEG[7] ;
 wire \Tile_X7Y14_S2BEGb[0] ;
 wire \Tile_X7Y14_S2BEGb[1] ;
 wire \Tile_X7Y14_S2BEGb[2] ;
 wire \Tile_X7Y14_S2BEGb[3] ;
 wire \Tile_X7Y14_S2BEGb[4] ;
 wire \Tile_X7Y14_S2BEGb[5] ;
 wire \Tile_X7Y14_S2BEGb[6] ;
 wire \Tile_X7Y14_S2BEGb[7] ;
 wire \Tile_X7Y14_S4BEG[0] ;
 wire \Tile_X7Y14_S4BEG[10] ;
 wire \Tile_X7Y14_S4BEG[11] ;
 wire \Tile_X7Y14_S4BEG[12] ;
 wire \Tile_X7Y14_S4BEG[13] ;
 wire \Tile_X7Y14_S4BEG[14] ;
 wire \Tile_X7Y14_S4BEG[15] ;
 wire \Tile_X7Y14_S4BEG[1] ;
 wire \Tile_X7Y14_S4BEG[2] ;
 wire \Tile_X7Y14_S4BEG[3] ;
 wire \Tile_X7Y14_S4BEG[4] ;
 wire \Tile_X7Y14_S4BEG[5] ;
 wire \Tile_X7Y14_S4BEG[6] ;
 wire \Tile_X7Y14_S4BEG[7] ;
 wire \Tile_X7Y14_S4BEG[8] ;
 wire \Tile_X7Y14_S4BEG[9] ;
 wire \Tile_X7Y14_SS4BEG[0] ;
 wire \Tile_X7Y14_SS4BEG[10] ;
 wire \Tile_X7Y14_SS4BEG[11] ;
 wire \Tile_X7Y14_SS4BEG[12] ;
 wire \Tile_X7Y14_SS4BEG[13] ;
 wire \Tile_X7Y14_SS4BEG[14] ;
 wire \Tile_X7Y14_SS4BEG[15] ;
 wire \Tile_X7Y14_SS4BEG[1] ;
 wire \Tile_X7Y14_SS4BEG[2] ;
 wire \Tile_X7Y14_SS4BEG[3] ;
 wire \Tile_X7Y14_SS4BEG[4] ;
 wire \Tile_X7Y14_SS4BEG[5] ;
 wire \Tile_X7Y14_SS4BEG[6] ;
 wire \Tile_X7Y14_SS4BEG[7] ;
 wire \Tile_X7Y14_SS4BEG[8] ;
 wire \Tile_X7Y14_SS4BEG[9] ;
 wire \Tile_X7Y14_W1BEG[0] ;
 wire \Tile_X7Y14_W1BEG[1] ;
 wire \Tile_X7Y14_W1BEG[2] ;
 wire \Tile_X7Y14_W1BEG[3] ;
 wire \Tile_X7Y14_W2BEG[0] ;
 wire \Tile_X7Y14_W2BEG[1] ;
 wire \Tile_X7Y14_W2BEG[2] ;
 wire \Tile_X7Y14_W2BEG[3] ;
 wire \Tile_X7Y14_W2BEG[4] ;
 wire \Tile_X7Y14_W2BEG[5] ;
 wire \Tile_X7Y14_W2BEG[6] ;
 wire \Tile_X7Y14_W2BEG[7] ;
 wire \Tile_X7Y14_W2BEGb[0] ;
 wire \Tile_X7Y14_W2BEGb[1] ;
 wire \Tile_X7Y14_W2BEGb[2] ;
 wire \Tile_X7Y14_W2BEGb[3] ;
 wire \Tile_X7Y14_W2BEGb[4] ;
 wire \Tile_X7Y14_W2BEGb[5] ;
 wire \Tile_X7Y14_W2BEGb[6] ;
 wire \Tile_X7Y14_W2BEGb[7] ;
 wire \Tile_X7Y14_W6BEG[0] ;
 wire \Tile_X7Y14_W6BEG[10] ;
 wire \Tile_X7Y14_W6BEG[11] ;
 wire \Tile_X7Y14_W6BEG[1] ;
 wire \Tile_X7Y14_W6BEG[2] ;
 wire \Tile_X7Y14_W6BEG[3] ;
 wire \Tile_X7Y14_W6BEG[4] ;
 wire \Tile_X7Y14_W6BEG[5] ;
 wire \Tile_X7Y14_W6BEG[6] ;
 wire \Tile_X7Y14_W6BEG[7] ;
 wire \Tile_X7Y14_W6BEG[8] ;
 wire \Tile_X7Y14_W6BEG[9] ;
 wire \Tile_X7Y14_WW4BEG[0] ;
 wire \Tile_X7Y14_WW4BEG[10] ;
 wire \Tile_X7Y14_WW4BEG[11] ;
 wire \Tile_X7Y14_WW4BEG[12] ;
 wire \Tile_X7Y14_WW4BEG[13] ;
 wire \Tile_X7Y14_WW4BEG[14] ;
 wire \Tile_X7Y14_WW4BEG[15] ;
 wire \Tile_X7Y14_WW4BEG[1] ;
 wire \Tile_X7Y14_WW4BEG[2] ;
 wire \Tile_X7Y14_WW4BEG[3] ;
 wire \Tile_X7Y14_WW4BEG[4] ;
 wire \Tile_X7Y14_WW4BEG[5] ;
 wire \Tile_X7Y14_WW4BEG[6] ;
 wire \Tile_X7Y14_WW4BEG[7] ;
 wire \Tile_X7Y14_WW4BEG[8] ;
 wire \Tile_X7Y14_WW4BEG[9] ;
 wire \Tile_X7Y15_FrameData_O[0] ;
 wire \Tile_X7Y15_FrameData_O[10] ;
 wire \Tile_X7Y15_FrameData_O[11] ;
 wire \Tile_X7Y15_FrameData_O[12] ;
 wire \Tile_X7Y15_FrameData_O[13] ;
 wire \Tile_X7Y15_FrameData_O[14] ;
 wire \Tile_X7Y15_FrameData_O[15] ;
 wire \Tile_X7Y15_FrameData_O[16] ;
 wire \Tile_X7Y15_FrameData_O[17] ;
 wire \Tile_X7Y15_FrameData_O[18] ;
 wire \Tile_X7Y15_FrameData_O[19] ;
 wire \Tile_X7Y15_FrameData_O[1] ;
 wire \Tile_X7Y15_FrameData_O[20] ;
 wire \Tile_X7Y15_FrameData_O[21] ;
 wire \Tile_X7Y15_FrameData_O[22] ;
 wire \Tile_X7Y15_FrameData_O[23] ;
 wire \Tile_X7Y15_FrameData_O[24] ;
 wire \Tile_X7Y15_FrameData_O[25] ;
 wire \Tile_X7Y15_FrameData_O[26] ;
 wire \Tile_X7Y15_FrameData_O[27] ;
 wire \Tile_X7Y15_FrameData_O[28] ;
 wire \Tile_X7Y15_FrameData_O[29] ;
 wire \Tile_X7Y15_FrameData_O[2] ;
 wire \Tile_X7Y15_FrameData_O[30] ;
 wire \Tile_X7Y15_FrameData_O[31] ;
 wire \Tile_X7Y15_FrameData_O[3] ;
 wire \Tile_X7Y15_FrameData_O[4] ;
 wire \Tile_X7Y15_FrameData_O[5] ;
 wire \Tile_X7Y15_FrameData_O[6] ;
 wire \Tile_X7Y15_FrameData_O[7] ;
 wire \Tile_X7Y15_FrameData_O[8] ;
 wire \Tile_X7Y15_FrameData_O[9] ;
 wire \Tile_X7Y15_FrameStrobe_O[0] ;
 wire \Tile_X7Y15_FrameStrobe_O[10] ;
 wire \Tile_X7Y15_FrameStrobe_O[11] ;
 wire \Tile_X7Y15_FrameStrobe_O[12] ;
 wire \Tile_X7Y15_FrameStrobe_O[13] ;
 wire \Tile_X7Y15_FrameStrobe_O[14] ;
 wire \Tile_X7Y15_FrameStrobe_O[15] ;
 wire \Tile_X7Y15_FrameStrobe_O[16] ;
 wire \Tile_X7Y15_FrameStrobe_O[17] ;
 wire \Tile_X7Y15_FrameStrobe_O[18] ;
 wire \Tile_X7Y15_FrameStrobe_O[19] ;
 wire \Tile_X7Y15_FrameStrobe_O[1] ;
 wire \Tile_X7Y15_FrameStrobe_O[2] ;
 wire \Tile_X7Y15_FrameStrobe_O[3] ;
 wire \Tile_X7Y15_FrameStrobe_O[4] ;
 wire \Tile_X7Y15_FrameStrobe_O[5] ;
 wire \Tile_X7Y15_FrameStrobe_O[6] ;
 wire \Tile_X7Y15_FrameStrobe_O[7] ;
 wire \Tile_X7Y15_FrameStrobe_O[8] ;
 wire \Tile_X7Y15_FrameStrobe_O[9] ;
 wire \Tile_X7Y15_N1BEG[0] ;
 wire \Tile_X7Y15_N1BEG[1] ;
 wire \Tile_X7Y15_N1BEG[2] ;
 wire \Tile_X7Y15_N1BEG[3] ;
 wire \Tile_X7Y15_N2BEG[0] ;
 wire \Tile_X7Y15_N2BEG[1] ;
 wire \Tile_X7Y15_N2BEG[2] ;
 wire \Tile_X7Y15_N2BEG[3] ;
 wire \Tile_X7Y15_N2BEG[4] ;
 wire \Tile_X7Y15_N2BEG[5] ;
 wire \Tile_X7Y15_N2BEG[6] ;
 wire \Tile_X7Y15_N2BEG[7] ;
 wire \Tile_X7Y15_N2BEGb[0] ;
 wire \Tile_X7Y15_N2BEGb[1] ;
 wire \Tile_X7Y15_N2BEGb[2] ;
 wire \Tile_X7Y15_N2BEGb[3] ;
 wire \Tile_X7Y15_N2BEGb[4] ;
 wire \Tile_X7Y15_N2BEGb[5] ;
 wire \Tile_X7Y15_N2BEGb[6] ;
 wire \Tile_X7Y15_N2BEGb[7] ;
 wire \Tile_X7Y15_N4BEG[0] ;
 wire \Tile_X7Y15_N4BEG[10] ;
 wire \Tile_X7Y15_N4BEG[11] ;
 wire \Tile_X7Y15_N4BEG[12] ;
 wire \Tile_X7Y15_N4BEG[13] ;
 wire \Tile_X7Y15_N4BEG[14] ;
 wire \Tile_X7Y15_N4BEG[15] ;
 wire \Tile_X7Y15_N4BEG[1] ;
 wire \Tile_X7Y15_N4BEG[2] ;
 wire \Tile_X7Y15_N4BEG[3] ;
 wire \Tile_X7Y15_N4BEG[4] ;
 wire \Tile_X7Y15_N4BEG[5] ;
 wire \Tile_X7Y15_N4BEG[6] ;
 wire \Tile_X7Y15_N4BEG[7] ;
 wire \Tile_X7Y15_N4BEG[8] ;
 wire \Tile_X7Y15_N4BEG[9] ;
 wire \Tile_X7Y15_NN4BEG[0] ;
 wire \Tile_X7Y15_NN4BEG[10] ;
 wire \Tile_X7Y15_NN4BEG[11] ;
 wire \Tile_X7Y15_NN4BEG[12] ;
 wire \Tile_X7Y15_NN4BEG[13] ;
 wire \Tile_X7Y15_NN4BEG[14] ;
 wire \Tile_X7Y15_NN4BEG[15] ;
 wire \Tile_X7Y15_NN4BEG[1] ;
 wire \Tile_X7Y15_NN4BEG[2] ;
 wire \Tile_X7Y15_NN4BEG[3] ;
 wire \Tile_X7Y15_NN4BEG[4] ;
 wire \Tile_X7Y15_NN4BEG[5] ;
 wire \Tile_X7Y15_NN4BEG[6] ;
 wire \Tile_X7Y15_NN4BEG[7] ;
 wire \Tile_X7Y15_NN4BEG[8] ;
 wire \Tile_X7Y15_NN4BEG[9] ;
 wire Tile_X7Y15_UserCLKo;
 wire \Tile_X7Y1_E1BEG[0] ;
 wire \Tile_X7Y1_E1BEG[1] ;
 wire \Tile_X7Y1_E1BEG[2] ;
 wire \Tile_X7Y1_E1BEG[3] ;
 wire \Tile_X7Y1_E2BEG[0] ;
 wire \Tile_X7Y1_E2BEG[1] ;
 wire \Tile_X7Y1_E2BEG[2] ;
 wire \Tile_X7Y1_E2BEG[3] ;
 wire \Tile_X7Y1_E2BEG[4] ;
 wire \Tile_X7Y1_E2BEG[5] ;
 wire \Tile_X7Y1_E2BEG[6] ;
 wire \Tile_X7Y1_E2BEG[7] ;
 wire \Tile_X7Y1_E2BEGb[0] ;
 wire \Tile_X7Y1_E2BEGb[1] ;
 wire \Tile_X7Y1_E2BEGb[2] ;
 wire \Tile_X7Y1_E2BEGb[3] ;
 wire \Tile_X7Y1_E2BEGb[4] ;
 wire \Tile_X7Y1_E2BEGb[5] ;
 wire \Tile_X7Y1_E2BEGb[6] ;
 wire \Tile_X7Y1_E2BEGb[7] ;
 wire \Tile_X7Y1_E6BEG[0] ;
 wire \Tile_X7Y1_E6BEG[10] ;
 wire \Tile_X7Y1_E6BEG[11] ;
 wire \Tile_X7Y1_E6BEG[1] ;
 wire \Tile_X7Y1_E6BEG[2] ;
 wire \Tile_X7Y1_E6BEG[3] ;
 wire \Tile_X7Y1_E6BEG[4] ;
 wire \Tile_X7Y1_E6BEG[5] ;
 wire \Tile_X7Y1_E6BEG[6] ;
 wire \Tile_X7Y1_E6BEG[7] ;
 wire \Tile_X7Y1_E6BEG[8] ;
 wire \Tile_X7Y1_E6BEG[9] ;
 wire \Tile_X7Y1_EE4BEG[0] ;
 wire \Tile_X7Y1_EE4BEG[10] ;
 wire \Tile_X7Y1_EE4BEG[11] ;
 wire \Tile_X7Y1_EE4BEG[12] ;
 wire \Tile_X7Y1_EE4BEG[13] ;
 wire \Tile_X7Y1_EE4BEG[14] ;
 wire \Tile_X7Y1_EE4BEG[15] ;
 wire \Tile_X7Y1_EE4BEG[1] ;
 wire \Tile_X7Y1_EE4BEG[2] ;
 wire \Tile_X7Y1_EE4BEG[3] ;
 wire \Tile_X7Y1_EE4BEG[4] ;
 wire \Tile_X7Y1_EE4BEG[5] ;
 wire \Tile_X7Y1_EE4BEG[6] ;
 wire \Tile_X7Y1_EE4BEG[7] ;
 wire \Tile_X7Y1_EE4BEG[8] ;
 wire \Tile_X7Y1_EE4BEG[9] ;
 wire \Tile_X7Y1_FrameData_O[0] ;
 wire \Tile_X7Y1_FrameData_O[10] ;
 wire \Tile_X7Y1_FrameData_O[11] ;
 wire \Tile_X7Y1_FrameData_O[12] ;
 wire \Tile_X7Y1_FrameData_O[13] ;
 wire \Tile_X7Y1_FrameData_O[14] ;
 wire \Tile_X7Y1_FrameData_O[15] ;
 wire \Tile_X7Y1_FrameData_O[16] ;
 wire \Tile_X7Y1_FrameData_O[17] ;
 wire \Tile_X7Y1_FrameData_O[18] ;
 wire \Tile_X7Y1_FrameData_O[19] ;
 wire \Tile_X7Y1_FrameData_O[1] ;
 wire \Tile_X7Y1_FrameData_O[20] ;
 wire \Tile_X7Y1_FrameData_O[21] ;
 wire \Tile_X7Y1_FrameData_O[22] ;
 wire \Tile_X7Y1_FrameData_O[23] ;
 wire \Tile_X7Y1_FrameData_O[24] ;
 wire \Tile_X7Y1_FrameData_O[25] ;
 wire \Tile_X7Y1_FrameData_O[26] ;
 wire \Tile_X7Y1_FrameData_O[27] ;
 wire \Tile_X7Y1_FrameData_O[28] ;
 wire \Tile_X7Y1_FrameData_O[29] ;
 wire \Tile_X7Y1_FrameData_O[2] ;
 wire \Tile_X7Y1_FrameData_O[30] ;
 wire \Tile_X7Y1_FrameData_O[31] ;
 wire \Tile_X7Y1_FrameData_O[3] ;
 wire \Tile_X7Y1_FrameData_O[4] ;
 wire \Tile_X7Y1_FrameData_O[5] ;
 wire \Tile_X7Y1_FrameData_O[6] ;
 wire \Tile_X7Y1_FrameData_O[7] ;
 wire \Tile_X7Y1_FrameData_O[8] ;
 wire \Tile_X7Y1_FrameData_O[9] ;
 wire \Tile_X7Y1_FrameStrobe_O[0] ;
 wire \Tile_X7Y1_FrameStrobe_O[10] ;
 wire \Tile_X7Y1_FrameStrobe_O[11] ;
 wire \Tile_X7Y1_FrameStrobe_O[12] ;
 wire \Tile_X7Y1_FrameStrobe_O[13] ;
 wire \Tile_X7Y1_FrameStrobe_O[14] ;
 wire \Tile_X7Y1_FrameStrobe_O[15] ;
 wire \Tile_X7Y1_FrameStrobe_O[16] ;
 wire \Tile_X7Y1_FrameStrobe_O[17] ;
 wire \Tile_X7Y1_FrameStrobe_O[18] ;
 wire \Tile_X7Y1_FrameStrobe_O[19] ;
 wire \Tile_X7Y1_FrameStrobe_O[1] ;
 wire \Tile_X7Y1_FrameStrobe_O[2] ;
 wire \Tile_X7Y1_FrameStrobe_O[3] ;
 wire \Tile_X7Y1_FrameStrobe_O[4] ;
 wire \Tile_X7Y1_FrameStrobe_O[5] ;
 wire \Tile_X7Y1_FrameStrobe_O[6] ;
 wire \Tile_X7Y1_FrameStrobe_O[7] ;
 wire \Tile_X7Y1_FrameStrobe_O[8] ;
 wire \Tile_X7Y1_FrameStrobe_O[9] ;
 wire \Tile_X7Y1_N1BEG[0] ;
 wire \Tile_X7Y1_N1BEG[1] ;
 wire \Tile_X7Y1_N1BEG[2] ;
 wire \Tile_X7Y1_N1BEG[3] ;
 wire \Tile_X7Y1_N2BEG[0] ;
 wire \Tile_X7Y1_N2BEG[1] ;
 wire \Tile_X7Y1_N2BEG[2] ;
 wire \Tile_X7Y1_N2BEG[3] ;
 wire \Tile_X7Y1_N2BEG[4] ;
 wire \Tile_X7Y1_N2BEG[5] ;
 wire \Tile_X7Y1_N2BEG[6] ;
 wire \Tile_X7Y1_N2BEG[7] ;
 wire \Tile_X7Y1_N2BEGb[0] ;
 wire \Tile_X7Y1_N2BEGb[1] ;
 wire \Tile_X7Y1_N2BEGb[2] ;
 wire \Tile_X7Y1_N2BEGb[3] ;
 wire \Tile_X7Y1_N2BEGb[4] ;
 wire \Tile_X7Y1_N2BEGb[5] ;
 wire \Tile_X7Y1_N2BEGb[6] ;
 wire \Tile_X7Y1_N2BEGb[7] ;
 wire \Tile_X7Y1_N4BEG[0] ;
 wire \Tile_X7Y1_N4BEG[10] ;
 wire \Tile_X7Y1_N4BEG[11] ;
 wire \Tile_X7Y1_N4BEG[12] ;
 wire \Tile_X7Y1_N4BEG[13] ;
 wire \Tile_X7Y1_N4BEG[14] ;
 wire \Tile_X7Y1_N4BEG[15] ;
 wire \Tile_X7Y1_N4BEG[1] ;
 wire \Tile_X7Y1_N4BEG[2] ;
 wire \Tile_X7Y1_N4BEG[3] ;
 wire \Tile_X7Y1_N4BEG[4] ;
 wire \Tile_X7Y1_N4BEG[5] ;
 wire \Tile_X7Y1_N4BEG[6] ;
 wire \Tile_X7Y1_N4BEG[7] ;
 wire \Tile_X7Y1_N4BEG[8] ;
 wire \Tile_X7Y1_N4BEG[9] ;
 wire \Tile_X7Y1_NN4BEG[0] ;
 wire \Tile_X7Y1_NN4BEG[10] ;
 wire \Tile_X7Y1_NN4BEG[11] ;
 wire \Tile_X7Y1_NN4BEG[12] ;
 wire \Tile_X7Y1_NN4BEG[13] ;
 wire \Tile_X7Y1_NN4BEG[14] ;
 wire \Tile_X7Y1_NN4BEG[15] ;
 wire \Tile_X7Y1_NN4BEG[1] ;
 wire \Tile_X7Y1_NN4BEG[2] ;
 wire \Tile_X7Y1_NN4BEG[3] ;
 wire \Tile_X7Y1_NN4BEG[4] ;
 wire \Tile_X7Y1_NN4BEG[5] ;
 wire \Tile_X7Y1_NN4BEG[6] ;
 wire \Tile_X7Y1_NN4BEG[7] ;
 wire \Tile_X7Y1_NN4BEG[8] ;
 wire \Tile_X7Y1_NN4BEG[9] ;
 wire Tile_X7Y1_UserCLKo;
 wire \Tile_X7Y1_W1BEG[0] ;
 wire \Tile_X7Y1_W1BEG[1] ;
 wire \Tile_X7Y1_W1BEG[2] ;
 wire \Tile_X7Y1_W1BEG[3] ;
 wire \Tile_X7Y1_W2BEG[0] ;
 wire \Tile_X7Y1_W2BEG[1] ;
 wire \Tile_X7Y1_W2BEG[2] ;
 wire \Tile_X7Y1_W2BEG[3] ;
 wire \Tile_X7Y1_W2BEG[4] ;
 wire \Tile_X7Y1_W2BEG[5] ;
 wire \Tile_X7Y1_W2BEG[6] ;
 wire \Tile_X7Y1_W2BEG[7] ;
 wire \Tile_X7Y1_W2BEGb[0] ;
 wire \Tile_X7Y1_W2BEGb[1] ;
 wire \Tile_X7Y1_W2BEGb[2] ;
 wire \Tile_X7Y1_W2BEGb[3] ;
 wire \Tile_X7Y1_W2BEGb[4] ;
 wire \Tile_X7Y1_W2BEGb[5] ;
 wire \Tile_X7Y1_W2BEGb[6] ;
 wire \Tile_X7Y1_W2BEGb[7] ;
 wire \Tile_X7Y1_W6BEG[0] ;
 wire \Tile_X7Y1_W6BEG[10] ;
 wire \Tile_X7Y1_W6BEG[11] ;
 wire \Tile_X7Y1_W6BEG[1] ;
 wire \Tile_X7Y1_W6BEG[2] ;
 wire \Tile_X7Y1_W6BEG[3] ;
 wire \Tile_X7Y1_W6BEG[4] ;
 wire \Tile_X7Y1_W6BEG[5] ;
 wire \Tile_X7Y1_W6BEG[6] ;
 wire \Tile_X7Y1_W6BEG[7] ;
 wire \Tile_X7Y1_W6BEG[8] ;
 wire \Tile_X7Y1_W6BEG[9] ;
 wire \Tile_X7Y1_WW4BEG[0] ;
 wire \Tile_X7Y1_WW4BEG[10] ;
 wire \Tile_X7Y1_WW4BEG[11] ;
 wire \Tile_X7Y1_WW4BEG[12] ;
 wire \Tile_X7Y1_WW4BEG[13] ;
 wire \Tile_X7Y1_WW4BEG[14] ;
 wire \Tile_X7Y1_WW4BEG[15] ;
 wire \Tile_X7Y1_WW4BEG[1] ;
 wire \Tile_X7Y1_WW4BEG[2] ;
 wire \Tile_X7Y1_WW4BEG[3] ;
 wire \Tile_X7Y1_WW4BEG[4] ;
 wire \Tile_X7Y1_WW4BEG[5] ;
 wire \Tile_X7Y1_WW4BEG[6] ;
 wire \Tile_X7Y1_WW4BEG[7] ;
 wire \Tile_X7Y1_WW4BEG[8] ;
 wire \Tile_X7Y1_WW4BEG[9] ;
 wire \Tile_X7Y2_E1BEG[0] ;
 wire \Tile_X7Y2_E1BEG[1] ;
 wire \Tile_X7Y2_E1BEG[2] ;
 wire \Tile_X7Y2_E1BEG[3] ;
 wire \Tile_X7Y2_E2BEG[0] ;
 wire \Tile_X7Y2_E2BEG[1] ;
 wire \Tile_X7Y2_E2BEG[2] ;
 wire \Tile_X7Y2_E2BEG[3] ;
 wire \Tile_X7Y2_E2BEG[4] ;
 wire \Tile_X7Y2_E2BEG[5] ;
 wire \Tile_X7Y2_E2BEG[6] ;
 wire \Tile_X7Y2_E2BEG[7] ;
 wire \Tile_X7Y2_E2BEGb[0] ;
 wire \Tile_X7Y2_E2BEGb[1] ;
 wire \Tile_X7Y2_E2BEGb[2] ;
 wire \Tile_X7Y2_E2BEGb[3] ;
 wire \Tile_X7Y2_E2BEGb[4] ;
 wire \Tile_X7Y2_E2BEGb[5] ;
 wire \Tile_X7Y2_E2BEGb[6] ;
 wire \Tile_X7Y2_E2BEGb[7] ;
 wire \Tile_X7Y2_E6BEG[0] ;
 wire \Tile_X7Y2_E6BEG[10] ;
 wire \Tile_X7Y2_E6BEG[11] ;
 wire \Tile_X7Y2_E6BEG[1] ;
 wire \Tile_X7Y2_E6BEG[2] ;
 wire \Tile_X7Y2_E6BEG[3] ;
 wire \Tile_X7Y2_E6BEG[4] ;
 wire \Tile_X7Y2_E6BEG[5] ;
 wire \Tile_X7Y2_E6BEG[6] ;
 wire \Tile_X7Y2_E6BEG[7] ;
 wire \Tile_X7Y2_E6BEG[8] ;
 wire \Tile_X7Y2_E6BEG[9] ;
 wire \Tile_X7Y2_EE4BEG[0] ;
 wire \Tile_X7Y2_EE4BEG[10] ;
 wire \Tile_X7Y2_EE4BEG[11] ;
 wire \Tile_X7Y2_EE4BEG[12] ;
 wire \Tile_X7Y2_EE4BEG[13] ;
 wire \Tile_X7Y2_EE4BEG[14] ;
 wire \Tile_X7Y2_EE4BEG[15] ;
 wire \Tile_X7Y2_EE4BEG[1] ;
 wire \Tile_X7Y2_EE4BEG[2] ;
 wire \Tile_X7Y2_EE4BEG[3] ;
 wire \Tile_X7Y2_EE4BEG[4] ;
 wire \Tile_X7Y2_EE4BEG[5] ;
 wire \Tile_X7Y2_EE4BEG[6] ;
 wire \Tile_X7Y2_EE4BEG[7] ;
 wire \Tile_X7Y2_EE4BEG[8] ;
 wire \Tile_X7Y2_EE4BEG[9] ;
 wire \Tile_X7Y2_FrameData_O[0] ;
 wire \Tile_X7Y2_FrameData_O[10] ;
 wire \Tile_X7Y2_FrameData_O[11] ;
 wire \Tile_X7Y2_FrameData_O[12] ;
 wire \Tile_X7Y2_FrameData_O[13] ;
 wire \Tile_X7Y2_FrameData_O[14] ;
 wire \Tile_X7Y2_FrameData_O[15] ;
 wire \Tile_X7Y2_FrameData_O[16] ;
 wire \Tile_X7Y2_FrameData_O[17] ;
 wire \Tile_X7Y2_FrameData_O[18] ;
 wire \Tile_X7Y2_FrameData_O[19] ;
 wire \Tile_X7Y2_FrameData_O[1] ;
 wire \Tile_X7Y2_FrameData_O[20] ;
 wire \Tile_X7Y2_FrameData_O[21] ;
 wire \Tile_X7Y2_FrameData_O[22] ;
 wire \Tile_X7Y2_FrameData_O[23] ;
 wire \Tile_X7Y2_FrameData_O[24] ;
 wire \Tile_X7Y2_FrameData_O[25] ;
 wire \Tile_X7Y2_FrameData_O[26] ;
 wire \Tile_X7Y2_FrameData_O[27] ;
 wire \Tile_X7Y2_FrameData_O[28] ;
 wire \Tile_X7Y2_FrameData_O[29] ;
 wire \Tile_X7Y2_FrameData_O[2] ;
 wire \Tile_X7Y2_FrameData_O[30] ;
 wire \Tile_X7Y2_FrameData_O[31] ;
 wire \Tile_X7Y2_FrameData_O[3] ;
 wire \Tile_X7Y2_FrameData_O[4] ;
 wire \Tile_X7Y2_FrameData_O[5] ;
 wire \Tile_X7Y2_FrameData_O[6] ;
 wire \Tile_X7Y2_FrameData_O[7] ;
 wire \Tile_X7Y2_FrameData_O[8] ;
 wire \Tile_X7Y2_FrameData_O[9] ;
 wire \Tile_X7Y2_S1BEG[0] ;
 wire \Tile_X7Y2_S1BEG[1] ;
 wire \Tile_X7Y2_S1BEG[2] ;
 wire \Tile_X7Y2_S1BEG[3] ;
 wire \Tile_X7Y2_S2BEG[0] ;
 wire \Tile_X7Y2_S2BEG[1] ;
 wire \Tile_X7Y2_S2BEG[2] ;
 wire \Tile_X7Y2_S2BEG[3] ;
 wire \Tile_X7Y2_S2BEG[4] ;
 wire \Tile_X7Y2_S2BEG[5] ;
 wire \Tile_X7Y2_S2BEG[6] ;
 wire \Tile_X7Y2_S2BEG[7] ;
 wire \Tile_X7Y2_S2BEGb[0] ;
 wire \Tile_X7Y2_S2BEGb[1] ;
 wire \Tile_X7Y2_S2BEGb[2] ;
 wire \Tile_X7Y2_S2BEGb[3] ;
 wire \Tile_X7Y2_S2BEGb[4] ;
 wire \Tile_X7Y2_S2BEGb[5] ;
 wire \Tile_X7Y2_S2BEGb[6] ;
 wire \Tile_X7Y2_S2BEGb[7] ;
 wire \Tile_X7Y2_S4BEG[0] ;
 wire \Tile_X7Y2_S4BEG[10] ;
 wire \Tile_X7Y2_S4BEG[11] ;
 wire \Tile_X7Y2_S4BEG[12] ;
 wire \Tile_X7Y2_S4BEG[13] ;
 wire \Tile_X7Y2_S4BEG[14] ;
 wire \Tile_X7Y2_S4BEG[15] ;
 wire \Tile_X7Y2_S4BEG[1] ;
 wire \Tile_X7Y2_S4BEG[2] ;
 wire \Tile_X7Y2_S4BEG[3] ;
 wire \Tile_X7Y2_S4BEG[4] ;
 wire \Tile_X7Y2_S4BEG[5] ;
 wire \Tile_X7Y2_S4BEG[6] ;
 wire \Tile_X7Y2_S4BEG[7] ;
 wire \Tile_X7Y2_S4BEG[8] ;
 wire \Tile_X7Y2_S4BEG[9] ;
 wire \Tile_X7Y2_SS4BEG[0] ;
 wire \Tile_X7Y2_SS4BEG[10] ;
 wire \Tile_X7Y2_SS4BEG[11] ;
 wire \Tile_X7Y2_SS4BEG[12] ;
 wire \Tile_X7Y2_SS4BEG[13] ;
 wire \Tile_X7Y2_SS4BEG[14] ;
 wire \Tile_X7Y2_SS4BEG[15] ;
 wire \Tile_X7Y2_SS4BEG[1] ;
 wire \Tile_X7Y2_SS4BEG[2] ;
 wire \Tile_X7Y2_SS4BEG[3] ;
 wire \Tile_X7Y2_SS4BEG[4] ;
 wire \Tile_X7Y2_SS4BEG[5] ;
 wire \Tile_X7Y2_SS4BEG[6] ;
 wire \Tile_X7Y2_SS4BEG[7] ;
 wire \Tile_X7Y2_SS4BEG[8] ;
 wire \Tile_X7Y2_SS4BEG[9] ;
 wire \Tile_X7Y2_W1BEG[0] ;
 wire \Tile_X7Y2_W1BEG[1] ;
 wire \Tile_X7Y2_W1BEG[2] ;
 wire \Tile_X7Y2_W1BEG[3] ;
 wire \Tile_X7Y2_W2BEG[0] ;
 wire \Tile_X7Y2_W2BEG[1] ;
 wire \Tile_X7Y2_W2BEG[2] ;
 wire \Tile_X7Y2_W2BEG[3] ;
 wire \Tile_X7Y2_W2BEG[4] ;
 wire \Tile_X7Y2_W2BEG[5] ;
 wire \Tile_X7Y2_W2BEG[6] ;
 wire \Tile_X7Y2_W2BEG[7] ;
 wire \Tile_X7Y2_W2BEGb[0] ;
 wire \Tile_X7Y2_W2BEGb[1] ;
 wire \Tile_X7Y2_W2BEGb[2] ;
 wire \Tile_X7Y2_W2BEGb[3] ;
 wire \Tile_X7Y2_W2BEGb[4] ;
 wire \Tile_X7Y2_W2BEGb[5] ;
 wire \Tile_X7Y2_W2BEGb[6] ;
 wire \Tile_X7Y2_W2BEGb[7] ;
 wire \Tile_X7Y2_W6BEG[0] ;
 wire \Tile_X7Y2_W6BEG[10] ;
 wire \Tile_X7Y2_W6BEG[11] ;
 wire \Tile_X7Y2_W6BEG[1] ;
 wire \Tile_X7Y2_W6BEG[2] ;
 wire \Tile_X7Y2_W6BEG[3] ;
 wire \Tile_X7Y2_W6BEG[4] ;
 wire \Tile_X7Y2_W6BEG[5] ;
 wire \Tile_X7Y2_W6BEG[6] ;
 wire \Tile_X7Y2_W6BEG[7] ;
 wire \Tile_X7Y2_W6BEG[8] ;
 wire \Tile_X7Y2_W6BEG[9] ;
 wire \Tile_X7Y2_WW4BEG[0] ;
 wire \Tile_X7Y2_WW4BEG[10] ;
 wire \Tile_X7Y2_WW4BEG[11] ;
 wire \Tile_X7Y2_WW4BEG[12] ;
 wire \Tile_X7Y2_WW4BEG[13] ;
 wire \Tile_X7Y2_WW4BEG[14] ;
 wire \Tile_X7Y2_WW4BEG[15] ;
 wire \Tile_X7Y2_WW4BEG[1] ;
 wire \Tile_X7Y2_WW4BEG[2] ;
 wire \Tile_X7Y2_WW4BEG[3] ;
 wire \Tile_X7Y2_WW4BEG[4] ;
 wire \Tile_X7Y2_WW4BEG[5] ;
 wire \Tile_X7Y2_WW4BEG[6] ;
 wire \Tile_X7Y2_WW4BEG[7] ;
 wire \Tile_X7Y2_WW4BEG[8] ;
 wire \Tile_X7Y2_WW4BEG[9] ;
 wire \Tile_X7Y3_E1BEG[0] ;
 wire \Tile_X7Y3_E1BEG[1] ;
 wire \Tile_X7Y3_E1BEG[2] ;
 wire \Tile_X7Y3_E1BEG[3] ;
 wire \Tile_X7Y3_E2BEG[0] ;
 wire \Tile_X7Y3_E2BEG[1] ;
 wire \Tile_X7Y3_E2BEG[2] ;
 wire \Tile_X7Y3_E2BEG[3] ;
 wire \Tile_X7Y3_E2BEG[4] ;
 wire \Tile_X7Y3_E2BEG[5] ;
 wire \Tile_X7Y3_E2BEG[6] ;
 wire \Tile_X7Y3_E2BEG[7] ;
 wire \Tile_X7Y3_E2BEGb[0] ;
 wire \Tile_X7Y3_E2BEGb[1] ;
 wire \Tile_X7Y3_E2BEGb[2] ;
 wire \Tile_X7Y3_E2BEGb[3] ;
 wire \Tile_X7Y3_E2BEGb[4] ;
 wire \Tile_X7Y3_E2BEGb[5] ;
 wire \Tile_X7Y3_E2BEGb[6] ;
 wire \Tile_X7Y3_E2BEGb[7] ;
 wire \Tile_X7Y3_E6BEG[0] ;
 wire \Tile_X7Y3_E6BEG[10] ;
 wire \Tile_X7Y3_E6BEG[11] ;
 wire \Tile_X7Y3_E6BEG[1] ;
 wire \Tile_X7Y3_E6BEG[2] ;
 wire \Tile_X7Y3_E6BEG[3] ;
 wire \Tile_X7Y3_E6BEG[4] ;
 wire \Tile_X7Y3_E6BEG[5] ;
 wire \Tile_X7Y3_E6BEG[6] ;
 wire \Tile_X7Y3_E6BEG[7] ;
 wire \Tile_X7Y3_E6BEG[8] ;
 wire \Tile_X7Y3_E6BEG[9] ;
 wire \Tile_X7Y3_EE4BEG[0] ;
 wire \Tile_X7Y3_EE4BEG[10] ;
 wire \Tile_X7Y3_EE4BEG[11] ;
 wire \Tile_X7Y3_EE4BEG[12] ;
 wire \Tile_X7Y3_EE4BEG[13] ;
 wire \Tile_X7Y3_EE4BEG[14] ;
 wire \Tile_X7Y3_EE4BEG[15] ;
 wire \Tile_X7Y3_EE4BEG[1] ;
 wire \Tile_X7Y3_EE4BEG[2] ;
 wire \Tile_X7Y3_EE4BEG[3] ;
 wire \Tile_X7Y3_EE4BEG[4] ;
 wire \Tile_X7Y3_EE4BEG[5] ;
 wire \Tile_X7Y3_EE4BEG[6] ;
 wire \Tile_X7Y3_EE4BEG[7] ;
 wire \Tile_X7Y3_EE4BEG[8] ;
 wire \Tile_X7Y3_EE4BEG[9] ;
 wire \Tile_X7Y3_FrameData_O[0] ;
 wire \Tile_X7Y3_FrameData_O[10] ;
 wire \Tile_X7Y3_FrameData_O[11] ;
 wire \Tile_X7Y3_FrameData_O[12] ;
 wire \Tile_X7Y3_FrameData_O[13] ;
 wire \Tile_X7Y3_FrameData_O[14] ;
 wire \Tile_X7Y3_FrameData_O[15] ;
 wire \Tile_X7Y3_FrameData_O[16] ;
 wire \Tile_X7Y3_FrameData_O[17] ;
 wire \Tile_X7Y3_FrameData_O[18] ;
 wire \Tile_X7Y3_FrameData_O[19] ;
 wire \Tile_X7Y3_FrameData_O[1] ;
 wire \Tile_X7Y3_FrameData_O[20] ;
 wire \Tile_X7Y3_FrameData_O[21] ;
 wire \Tile_X7Y3_FrameData_O[22] ;
 wire \Tile_X7Y3_FrameData_O[23] ;
 wire \Tile_X7Y3_FrameData_O[24] ;
 wire \Tile_X7Y3_FrameData_O[25] ;
 wire \Tile_X7Y3_FrameData_O[26] ;
 wire \Tile_X7Y3_FrameData_O[27] ;
 wire \Tile_X7Y3_FrameData_O[28] ;
 wire \Tile_X7Y3_FrameData_O[29] ;
 wire \Tile_X7Y3_FrameData_O[2] ;
 wire \Tile_X7Y3_FrameData_O[30] ;
 wire \Tile_X7Y3_FrameData_O[31] ;
 wire \Tile_X7Y3_FrameData_O[3] ;
 wire \Tile_X7Y3_FrameData_O[4] ;
 wire \Tile_X7Y3_FrameData_O[5] ;
 wire \Tile_X7Y3_FrameData_O[6] ;
 wire \Tile_X7Y3_FrameData_O[7] ;
 wire \Tile_X7Y3_FrameData_O[8] ;
 wire \Tile_X7Y3_FrameData_O[9] ;
 wire \Tile_X7Y3_FrameStrobe_O[0] ;
 wire \Tile_X7Y3_FrameStrobe_O[10] ;
 wire \Tile_X7Y3_FrameStrobe_O[11] ;
 wire \Tile_X7Y3_FrameStrobe_O[12] ;
 wire \Tile_X7Y3_FrameStrobe_O[13] ;
 wire \Tile_X7Y3_FrameStrobe_O[14] ;
 wire \Tile_X7Y3_FrameStrobe_O[15] ;
 wire \Tile_X7Y3_FrameStrobe_O[16] ;
 wire \Tile_X7Y3_FrameStrobe_O[17] ;
 wire \Tile_X7Y3_FrameStrobe_O[18] ;
 wire \Tile_X7Y3_FrameStrobe_O[19] ;
 wire \Tile_X7Y3_FrameStrobe_O[1] ;
 wire \Tile_X7Y3_FrameStrobe_O[2] ;
 wire \Tile_X7Y3_FrameStrobe_O[3] ;
 wire \Tile_X7Y3_FrameStrobe_O[4] ;
 wire \Tile_X7Y3_FrameStrobe_O[5] ;
 wire \Tile_X7Y3_FrameStrobe_O[6] ;
 wire \Tile_X7Y3_FrameStrobe_O[7] ;
 wire \Tile_X7Y3_FrameStrobe_O[8] ;
 wire \Tile_X7Y3_FrameStrobe_O[9] ;
 wire \Tile_X7Y3_N1BEG[0] ;
 wire \Tile_X7Y3_N1BEG[1] ;
 wire \Tile_X7Y3_N1BEG[2] ;
 wire \Tile_X7Y3_N1BEG[3] ;
 wire \Tile_X7Y3_N2BEG[0] ;
 wire \Tile_X7Y3_N2BEG[1] ;
 wire \Tile_X7Y3_N2BEG[2] ;
 wire \Tile_X7Y3_N2BEG[3] ;
 wire \Tile_X7Y3_N2BEG[4] ;
 wire \Tile_X7Y3_N2BEG[5] ;
 wire \Tile_X7Y3_N2BEG[6] ;
 wire \Tile_X7Y3_N2BEG[7] ;
 wire \Tile_X7Y3_N2BEGb[0] ;
 wire \Tile_X7Y3_N2BEGb[1] ;
 wire \Tile_X7Y3_N2BEGb[2] ;
 wire \Tile_X7Y3_N2BEGb[3] ;
 wire \Tile_X7Y3_N2BEGb[4] ;
 wire \Tile_X7Y3_N2BEGb[5] ;
 wire \Tile_X7Y3_N2BEGb[6] ;
 wire \Tile_X7Y3_N2BEGb[7] ;
 wire \Tile_X7Y3_N4BEG[0] ;
 wire \Tile_X7Y3_N4BEG[10] ;
 wire \Tile_X7Y3_N4BEG[11] ;
 wire \Tile_X7Y3_N4BEG[12] ;
 wire \Tile_X7Y3_N4BEG[13] ;
 wire \Tile_X7Y3_N4BEG[14] ;
 wire \Tile_X7Y3_N4BEG[15] ;
 wire \Tile_X7Y3_N4BEG[1] ;
 wire \Tile_X7Y3_N4BEG[2] ;
 wire \Tile_X7Y3_N4BEG[3] ;
 wire \Tile_X7Y3_N4BEG[4] ;
 wire \Tile_X7Y3_N4BEG[5] ;
 wire \Tile_X7Y3_N4BEG[6] ;
 wire \Tile_X7Y3_N4BEG[7] ;
 wire \Tile_X7Y3_N4BEG[8] ;
 wire \Tile_X7Y3_N4BEG[9] ;
 wire \Tile_X7Y3_NN4BEG[0] ;
 wire \Tile_X7Y3_NN4BEG[10] ;
 wire \Tile_X7Y3_NN4BEG[11] ;
 wire \Tile_X7Y3_NN4BEG[12] ;
 wire \Tile_X7Y3_NN4BEG[13] ;
 wire \Tile_X7Y3_NN4BEG[14] ;
 wire \Tile_X7Y3_NN4BEG[15] ;
 wire \Tile_X7Y3_NN4BEG[1] ;
 wire \Tile_X7Y3_NN4BEG[2] ;
 wire \Tile_X7Y3_NN4BEG[3] ;
 wire \Tile_X7Y3_NN4BEG[4] ;
 wire \Tile_X7Y3_NN4BEG[5] ;
 wire \Tile_X7Y3_NN4BEG[6] ;
 wire \Tile_X7Y3_NN4BEG[7] ;
 wire \Tile_X7Y3_NN4BEG[8] ;
 wire \Tile_X7Y3_NN4BEG[9] ;
 wire Tile_X7Y3_UserCLKo;
 wire \Tile_X7Y3_W1BEG[0] ;
 wire \Tile_X7Y3_W1BEG[1] ;
 wire \Tile_X7Y3_W1BEG[2] ;
 wire \Tile_X7Y3_W1BEG[3] ;
 wire \Tile_X7Y3_W2BEG[0] ;
 wire \Tile_X7Y3_W2BEG[1] ;
 wire \Tile_X7Y3_W2BEG[2] ;
 wire \Tile_X7Y3_W2BEG[3] ;
 wire \Tile_X7Y3_W2BEG[4] ;
 wire \Tile_X7Y3_W2BEG[5] ;
 wire \Tile_X7Y3_W2BEG[6] ;
 wire \Tile_X7Y3_W2BEG[7] ;
 wire \Tile_X7Y3_W2BEGb[0] ;
 wire \Tile_X7Y3_W2BEGb[1] ;
 wire \Tile_X7Y3_W2BEGb[2] ;
 wire \Tile_X7Y3_W2BEGb[3] ;
 wire \Tile_X7Y3_W2BEGb[4] ;
 wire \Tile_X7Y3_W2BEGb[5] ;
 wire \Tile_X7Y3_W2BEGb[6] ;
 wire \Tile_X7Y3_W2BEGb[7] ;
 wire \Tile_X7Y3_W6BEG[0] ;
 wire \Tile_X7Y3_W6BEG[10] ;
 wire \Tile_X7Y3_W6BEG[11] ;
 wire \Tile_X7Y3_W6BEG[1] ;
 wire \Tile_X7Y3_W6BEG[2] ;
 wire \Tile_X7Y3_W6BEG[3] ;
 wire \Tile_X7Y3_W6BEG[4] ;
 wire \Tile_X7Y3_W6BEG[5] ;
 wire \Tile_X7Y3_W6BEG[6] ;
 wire \Tile_X7Y3_W6BEG[7] ;
 wire \Tile_X7Y3_W6BEG[8] ;
 wire \Tile_X7Y3_W6BEG[9] ;
 wire \Tile_X7Y3_WW4BEG[0] ;
 wire \Tile_X7Y3_WW4BEG[10] ;
 wire \Tile_X7Y3_WW4BEG[11] ;
 wire \Tile_X7Y3_WW4BEG[12] ;
 wire \Tile_X7Y3_WW4BEG[13] ;
 wire \Tile_X7Y3_WW4BEG[14] ;
 wire \Tile_X7Y3_WW4BEG[15] ;
 wire \Tile_X7Y3_WW4BEG[1] ;
 wire \Tile_X7Y3_WW4BEG[2] ;
 wire \Tile_X7Y3_WW4BEG[3] ;
 wire \Tile_X7Y3_WW4BEG[4] ;
 wire \Tile_X7Y3_WW4BEG[5] ;
 wire \Tile_X7Y3_WW4BEG[6] ;
 wire \Tile_X7Y3_WW4BEG[7] ;
 wire \Tile_X7Y3_WW4BEG[8] ;
 wire \Tile_X7Y3_WW4BEG[9] ;
 wire \Tile_X7Y4_E1BEG[0] ;
 wire \Tile_X7Y4_E1BEG[1] ;
 wire \Tile_X7Y4_E1BEG[2] ;
 wire \Tile_X7Y4_E1BEG[3] ;
 wire \Tile_X7Y4_E2BEG[0] ;
 wire \Tile_X7Y4_E2BEG[1] ;
 wire \Tile_X7Y4_E2BEG[2] ;
 wire \Tile_X7Y4_E2BEG[3] ;
 wire \Tile_X7Y4_E2BEG[4] ;
 wire \Tile_X7Y4_E2BEG[5] ;
 wire \Tile_X7Y4_E2BEG[6] ;
 wire \Tile_X7Y4_E2BEG[7] ;
 wire \Tile_X7Y4_E2BEGb[0] ;
 wire \Tile_X7Y4_E2BEGb[1] ;
 wire \Tile_X7Y4_E2BEGb[2] ;
 wire \Tile_X7Y4_E2BEGb[3] ;
 wire \Tile_X7Y4_E2BEGb[4] ;
 wire \Tile_X7Y4_E2BEGb[5] ;
 wire \Tile_X7Y4_E2BEGb[6] ;
 wire \Tile_X7Y4_E2BEGb[7] ;
 wire \Tile_X7Y4_E6BEG[0] ;
 wire \Tile_X7Y4_E6BEG[10] ;
 wire \Tile_X7Y4_E6BEG[11] ;
 wire \Tile_X7Y4_E6BEG[1] ;
 wire \Tile_X7Y4_E6BEG[2] ;
 wire \Tile_X7Y4_E6BEG[3] ;
 wire \Tile_X7Y4_E6BEG[4] ;
 wire \Tile_X7Y4_E6BEG[5] ;
 wire \Tile_X7Y4_E6BEG[6] ;
 wire \Tile_X7Y4_E6BEG[7] ;
 wire \Tile_X7Y4_E6BEG[8] ;
 wire \Tile_X7Y4_E6BEG[9] ;
 wire \Tile_X7Y4_EE4BEG[0] ;
 wire \Tile_X7Y4_EE4BEG[10] ;
 wire \Tile_X7Y4_EE4BEG[11] ;
 wire \Tile_X7Y4_EE4BEG[12] ;
 wire \Tile_X7Y4_EE4BEG[13] ;
 wire \Tile_X7Y4_EE4BEG[14] ;
 wire \Tile_X7Y4_EE4BEG[15] ;
 wire \Tile_X7Y4_EE4BEG[1] ;
 wire \Tile_X7Y4_EE4BEG[2] ;
 wire \Tile_X7Y4_EE4BEG[3] ;
 wire \Tile_X7Y4_EE4BEG[4] ;
 wire \Tile_X7Y4_EE4BEG[5] ;
 wire \Tile_X7Y4_EE4BEG[6] ;
 wire \Tile_X7Y4_EE4BEG[7] ;
 wire \Tile_X7Y4_EE4BEG[8] ;
 wire \Tile_X7Y4_EE4BEG[9] ;
 wire \Tile_X7Y4_FrameData_O[0] ;
 wire \Tile_X7Y4_FrameData_O[10] ;
 wire \Tile_X7Y4_FrameData_O[11] ;
 wire \Tile_X7Y4_FrameData_O[12] ;
 wire \Tile_X7Y4_FrameData_O[13] ;
 wire \Tile_X7Y4_FrameData_O[14] ;
 wire \Tile_X7Y4_FrameData_O[15] ;
 wire \Tile_X7Y4_FrameData_O[16] ;
 wire \Tile_X7Y4_FrameData_O[17] ;
 wire \Tile_X7Y4_FrameData_O[18] ;
 wire \Tile_X7Y4_FrameData_O[19] ;
 wire \Tile_X7Y4_FrameData_O[1] ;
 wire \Tile_X7Y4_FrameData_O[20] ;
 wire \Tile_X7Y4_FrameData_O[21] ;
 wire \Tile_X7Y4_FrameData_O[22] ;
 wire \Tile_X7Y4_FrameData_O[23] ;
 wire \Tile_X7Y4_FrameData_O[24] ;
 wire \Tile_X7Y4_FrameData_O[25] ;
 wire \Tile_X7Y4_FrameData_O[26] ;
 wire \Tile_X7Y4_FrameData_O[27] ;
 wire \Tile_X7Y4_FrameData_O[28] ;
 wire \Tile_X7Y4_FrameData_O[29] ;
 wire \Tile_X7Y4_FrameData_O[2] ;
 wire \Tile_X7Y4_FrameData_O[30] ;
 wire \Tile_X7Y4_FrameData_O[31] ;
 wire \Tile_X7Y4_FrameData_O[3] ;
 wire \Tile_X7Y4_FrameData_O[4] ;
 wire \Tile_X7Y4_FrameData_O[5] ;
 wire \Tile_X7Y4_FrameData_O[6] ;
 wire \Tile_X7Y4_FrameData_O[7] ;
 wire \Tile_X7Y4_FrameData_O[8] ;
 wire \Tile_X7Y4_FrameData_O[9] ;
 wire \Tile_X7Y4_S1BEG[0] ;
 wire \Tile_X7Y4_S1BEG[1] ;
 wire \Tile_X7Y4_S1BEG[2] ;
 wire \Tile_X7Y4_S1BEG[3] ;
 wire \Tile_X7Y4_S2BEG[0] ;
 wire \Tile_X7Y4_S2BEG[1] ;
 wire \Tile_X7Y4_S2BEG[2] ;
 wire \Tile_X7Y4_S2BEG[3] ;
 wire \Tile_X7Y4_S2BEG[4] ;
 wire \Tile_X7Y4_S2BEG[5] ;
 wire \Tile_X7Y4_S2BEG[6] ;
 wire \Tile_X7Y4_S2BEG[7] ;
 wire \Tile_X7Y4_S2BEGb[0] ;
 wire \Tile_X7Y4_S2BEGb[1] ;
 wire \Tile_X7Y4_S2BEGb[2] ;
 wire \Tile_X7Y4_S2BEGb[3] ;
 wire \Tile_X7Y4_S2BEGb[4] ;
 wire \Tile_X7Y4_S2BEGb[5] ;
 wire \Tile_X7Y4_S2BEGb[6] ;
 wire \Tile_X7Y4_S2BEGb[7] ;
 wire \Tile_X7Y4_S4BEG[0] ;
 wire \Tile_X7Y4_S4BEG[10] ;
 wire \Tile_X7Y4_S4BEG[11] ;
 wire \Tile_X7Y4_S4BEG[12] ;
 wire \Tile_X7Y4_S4BEG[13] ;
 wire \Tile_X7Y4_S4BEG[14] ;
 wire \Tile_X7Y4_S4BEG[15] ;
 wire \Tile_X7Y4_S4BEG[1] ;
 wire \Tile_X7Y4_S4BEG[2] ;
 wire \Tile_X7Y4_S4BEG[3] ;
 wire \Tile_X7Y4_S4BEG[4] ;
 wire \Tile_X7Y4_S4BEG[5] ;
 wire \Tile_X7Y4_S4BEG[6] ;
 wire \Tile_X7Y4_S4BEG[7] ;
 wire \Tile_X7Y4_S4BEG[8] ;
 wire \Tile_X7Y4_S4BEG[9] ;
 wire \Tile_X7Y4_SS4BEG[0] ;
 wire \Tile_X7Y4_SS4BEG[10] ;
 wire \Tile_X7Y4_SS4BEG[11] ;
 wire \Tile_X7Y4_SS4BEG[12] ;
 wire \Tile_X7Y4_SS4BEG[13] ;
 wire \Tile_X7Y4_SS4BEG[14] ;
 wire \Tile_X7Y4_SS4BEG[15] ;
 wire \Tile_X7Y4_SS4BEG[1] ;
 wire \Tile_X7Y4_SS4BEG[2] ;
 wire \Tile_X7Y4_SS4BEG[3] ;
 wire \Tile_X7Y4_SS4BEG[4] ;
 wire \Tile_X7Y4_SS4BEG[5] ;
 wire \Tile_X7Y4_SS4BEG[6] ;
 wire \Tile_X7Y4_SS4BEG[7] ;
 wire \Tile_X7Y4_SS4BEG[8] ;
 wire \Tile_X7Y4_SS4BEG[9] ;
 wire \Tile_X7Y4_W1BEG[0] ;
 wire \Tile_X7Y4_W1BEG[1] ;
 wire \Tile_X7Y4_W1BEG[2] ;
 wire \Tile_X7Y4_W1BEG[3] ;
 wire \Tile_X7Y4_W2BEG[0] ;
 wire \Tile_X7Y4_W2BEG[1] ;
 wire \Tile_X7Y4_W2BEG[2] ;
 wire \Tile_X7Y4_W2BEG[3] ;
 wire \Tile_X7Y4_W2BEG[4] ;
 wire \Tile_X7Y4_W2BEG[5] ;
 wire \Tile_X7Y4_W2BEG[6] ;
 wire \Tile_X7Y4_W2BEG[7] ;
 wire \Tile_X7Y4_W2BEGb[0] ;
 wire \Tile_X7Y4_W2BEGb[1] ;
 wire \Tile_X7Y4_W2BEGb[2] ;
 wire \Tile_X7Y4_W2BEGb[3] ;
 wire \Tile_X7Y4_W2BEGb[4] ;
 wire \Tile_X7Y4_W2BEGb[5] ;
 wire \Tile_X7Y4_W2BEGb[6] ;
 wire \Tile_X7Y4_W2BEGb[7] ;
 wire \Tile_X7Y4_W6BEG[0] ;
 wire \Tile_X7Y4_W6BEG[10] ;
 wire \Tile_X7Y4_W6BEG[11] ;
 wire \Tile_X7Y4_W6BEG[1] ;
 wire \Tile_X7Y4_W6BEG[2] ;
 wire \Tile_X7Y4_W6BEG[3] ;
 wire \Tile_X7Y4_W6BEG[4] ;
 wire \Tile_X7Y4_W6BEG[5] ;
 wire \Tile_X7Y4_W6BEG[6] ;
 wire \Tile_X7Y4_W6BEG[7] ;
 wire \Tile_X7Y4_W6BEG[8] ;
 wire \Tile_X7Y4_W6BEG[9] ;
 wire \Tile_X7Y4_WW4BEG[0] ;
 wire \Tile_X7Y4_WW4BEG[10] ;
 wire \Tile_X7Y4_WW4BEG[11] ;
 wire \Tile_X7Y4_WW4BEG[12] ;
 wire \Tile_X7Y4_WW4BEG[13] ;
 wire \Tile_X7Y4_WW4BEG[14] ;
 wire \Tile_X7Y4_WW4BEG[15] ;
 wire \Tile_X7Y4_WW4BEG[1] ;
 wire \Tile_X7Y4_WW4BEG[2] ;
 wire \Tile_X7Y4_WW4BEG[3] ;
 wire \Tile_X7Y4_WW4BEG[4] ;
 wire \Tile_X7Y4_WW4BEG[5] ;
 wire \Tile_X7Y4_WW4BEG[6] ;
 wire \Tile_X7Y4_WW4BEG[7] ;
 wire \Tile_X7Y4_WW4BEG[8] ;
 wire \Tile_X7Y4_WW4BEG[9] ;
 wire \Tile_X7Y5_E1BEG[0] ;
 wire \Tile_X7Y5_E1BEG[1] ;
 wire \Tile_X7Y5_E1BEG[2] ;
 wire \Tile_X7Y5_E1BEG[3] ;
 wire \Tile_X7Y5_E2BEG[0] ;
 wire \Tile_X7Y5_E2BEG[1] ;
 wire \Tile_X7Y5_E2BEG[2] ;
 wire \Tile_X7Y5_E2BEG[3] ;
 wire \Tile_X7Y5_E2BEG[4] ;
 wire \Tile_X7Y5_E2BEG[5] ;
 wire \Tile_X7Y5_E2BEG[6] ;
 wire \Tile_X7Y5_E2BEG[7] ;
 wire \Tile_X7Y5_E2BEGb[0] ;
 wire \Tile_X7Y5_E2BEGb[1] ;
 wire \Tile_X7Y5_E2BEGb[2] ;
 wire \Tile_X7Y5_E2BEGb[3] ;
 wire \Tile_X7Y5_E2BEGb[4] ;
 wire \Tile_X7Y5_E2BEGb[5] ;
 wire \Tile_X7Y5_E2BEGb[6] ;
 wire \Tile_X7Y5_E2BEGb[7] ;
 wire \Tile_X7Y5_E6BEG[0] ;
 wire \Tile_X7Y5_E6BEG[10] ;
 wire \Tile_X7Y5_E6BEG[11] ;
 wire \Tile_X7Y5_E6BEG[1] ;
 wire \Tile_X7Y5_E6BEG[2] ;
 wire \Tile_X7Y5_E6BEG[3] ;
 wire \Tile_X7Y5_E6BEG[4] ;
 wire \Tile_X7Y5_E6BEG[5] ;
 wire \Tile_X7Y5_E6BEG[6] ;
 wire \Tile_X7Y5_E6BEG[7] ;
 wire \Tile_X7Y5_E6BEG[8] ;
 wire \Tile_X7Y5_E6BEG[9] ;
 wire \Tile_X7Y5_EE4BEG[0] ;
 wire \Tile_X7Y5_EE4BEG[10] ;
 wire \Tile_X7Y5_EE4BEG[11] ;
 wire \Tile_X7Y5_EE4BEG[12] ;
 wire \Tile_X7Y5_EE4BEG[13] ;
 wire \Tile_X7Y5_EE4BEG[14] ;
 wire \Tile_X7Y5_EE4BEG[15] ;
 wire \Tile_X7Y5_EE4BEG[1] ;
 wire \Tile_X7Y5_EE4BEG[2] ;
 wire \Tile_X7Y5_EE4BEG[3] ;
 wire \Tile_X7Y5_EE4BEG[4] ;
 wire \Tile_X7Y5_EE4BEG[5] ;
 wire \Tile_X7Y5_EE4BEG[6] ;
 wire \Tile_X7Y5_EE4BEG[7] ;
 wire \Tile_X7Y5_EE4BEG[8] ;
 wire \Tile_X7Y5_EE4BEG[9] ;
 wire \Tile_X7Y5_FrameData_O[0] ;
 wire \Tile_X7Y5_FrameData_O[10] ;
 wire \Tile_X7Y5_FrameData_O[11] ;
 wire \Tile_X7Y5_FrameData_O[12] ;
 wire \Tile_X7Y5_FrameData_O[13] ;
 wire \Tile_X7Y5_FrameData_O[14] ;
 wire \Tile_X7Y5_FrameData_O[15] ;
 wire \Tile_X7Y5_FrameData_O[16] ;
 wire \Tile_X7Y5_FrameData_O[17] ;
 wire \Tile_X7Y5_FrameData_O[18] ;
 wire \Tile_X7Y5_FrameData_O[19] ;
 wire \Tile_X7Y5_FrameData_O[1] ;
 wire \Tile_X7Y5_FrameData_O[20] ;
 wire \Tile_X7Y5_FrameData_O[21] ;
 wire \Tile_X7Y5_FrameData_O[22] ;
 wire \Tile_X7Y5_FrameData_O[23] ;
 wire \Tile_X7Y5_FrameData_O[24] ;
 wire \Tile_X7Y5_FrameData_O[25] ;
 wire \Tile_X7Y5_FrameData_O[26] ;
 wire \Tile_X7Y5_FrameData_O[27] ;
 wire \Tile_X7Y5_FrameData_O[28] ;
 wire \Tile_X7Y5_FrameData_O[29] ;
 wire \Tile_X7Y5_FrameData_O[2] ;
 wire \Tile_X7Y5_FrameData_O[30] ;
 wire \Tile_X7Y5_FrameData_O[31] ;
 wire \Tile_X7Y5_FrameData_O[3] ;
 wire \Tile_X7Y5_FrameData_O[4] ;
 wire \Tile_X7Y5_FrameData_O[5] ;
 wire \Tile_X7Y5_FrameData_O[6] ;
 wire \Tile_X7Y5_FrameData_O[7] ;
 wire \Tile_X7Y5_FrameData_O[8] ;
 wire \Tile_X7Y5_FrameData_O[9] ;
 wire \Tile_X7Y5_FrameStrobe_O[0] ;
 wire \Tile_X7Y5_FrameStrobe_O[10] ;
 wire \Tile_X7Y5_FrameStrobe_O[11] ;
 wire \Tile_X7Y5_FrameStrobe_O[12] ;
 wire \Tile_X7Y5_FrameStrobe_O[13] ;
 wire \Tile_X7Y5_FrameStrobe_O[14] ;
 wire \Tile_X7Y5_FrameStrobe_O[15] ;
 wire \Tile_X7Y5_FrameStrobe_O[16] ;
 wire \Tile_X7Y5_FrameStrobe_O[17] ;
 wire \Tile_X7Y5_FrameStrobe_O[18] ;
 wire \Tile_X7Y5_FrameStrobe_O[19] ;
 wire \Tile_X7Y5_FrameStrobe_O[1] ;
 wire \Tile_X7Y5_FrameStrobe_O[2] ;
 wire \Tile_X7Y5_FrameStrobe_O[3] ;
 wire \Tile_X7Y5_FrameStrobe_O[4] ;
 wire \Tile_X7Y5_FrameStrobe_O[5] ;
 wire \Tile_X7Y5_FrameStrobe_O[6] ;
 wire \Tile_X7Y5_FrameStrobe_O[7] ;
 wire \Tile_X7Y5_FrameStrobe_O[8] ;
 wire \Tile_X7Y5_FrameStrobe_O[9] ;
 wire \Tile_X7Y5_N1BEG[0] ;
 wire \Tile_X7Y5_N1BEG[1] ;
 wire \Tile_X7Y5_N1BEG[2] ;
 wire \Tile_X7Y5_N1BEG[3] ;
 wire \Tile_X7Y5_N2BEG[0] ;
 wire \Tile_X7Y5_N2BEG[1] ;
 wire \Tile_X7Y5_N2BEG[2] ;
 wire \Tile_X7Y5_N2BEG[3] ;
 wire \Tile_X7Y5_N2BEG[4] ;
 wire \Tile_X7Y5_N2BEG[5] ;
 wire \Tile_X7Y5_N2BEG[6] ;
 wire \Tile_X7Y5_N2BEG[7] ;
 wire \Tile_X7Y5_N2BEGb[0] ;
 wire \Tile_X7Y5_N2BEGb[1] ;
 wire \Tile_X7Y5_N2BEGb[2] ;
 wire \Tile_X7Y5_N2BEGb[3] ;
 wire \Tile_X7Y5_N2BEGb[4] ;
 wire \Tile_X7Y5_N2BEGb[5] ;
 wire \Tile_X7Y5_N2BEGb[6] ;
 wire \Tile_X7Y5_N2BEGb[7] ;
 wire \Tile_X7Y5_N4BEG[0] ;
 wire \Tile_X7Y5_N4BEG[10] ;
 wire \Tile_X7Y5_N4BEG[11] ;
 wire \Tile_X7Y5_N4BEG[12] ;
 wire \Tile_X7Y5_N4BEG[13] ;
 wire \Tile_X7Y5_N4BEG[14] ;
 wire \Tile_X7Y5_N4BEG[15] ;
 wire \Tile_X7Y5_N4BEG[1] ;
 wire \Tile_X7Y5_N4BEG[2] ;
 wire \Tile_X7Y5_N4BEG[3] ;
 wire \Tile_X7Y5_N4BEG[4] ;
 wire \Tile_X7Y5_N4BEG[5] ;
 wire \Tile_X7Y5_N4BEG[6] ;
 wire \Tile_X7Y5_N4BEG[7] ;
 wire \Tile_X7Y5_N4BEG[8] ;
 wire \Tile_X7Y5_N4BEG[9] ;
 wire \Tile_X7Y5_NN4BEG[0] ;
 wire \Tile_X7Y5_NN4BEG[10] ;
 wire \Tile_X7Y5_NN4BEG[11] ;
 wire \Tile_X7Y5_NN4BEG[12] ;
 wire \Tile_X7Y5_NN4BEG[13] ;
 wire \Tile_X7Y5_NN4BEG[14] ;
 wire \Tile_X7Y5_NN4BEG[15] ;
 wire \Tile_X7Y5_NN4BEG[1] ;
 wire \Tile_X7Y5_NN4BEG[2] ;
 wire \Tile_X7Y5_NN4BEG[3] ;
 wire \Tile_X7Y5_NN4BEG[4] ;
 wire \Tile_X7Y5_NN4BEG[5] ;
 wire \Tile_X7Y5_NN4BEG[6] ;
 wire \Tile_X7Y5_NN4BEG[7] ;
 wire \Tile_X7Y5_NN4BEG[8] ;
 wire \Tile_X7Y5_NN4BEG[9] ;
 wire Tile_X7Y5_UserCLKo;
 wire \Tile_X7Y5_W1BEG[0] ;
 wire \Tile_X7Y5_W1BEG[1] ;
 wire \Tile_X7Y5_W1BEG[2] ;
 wire \Tile_X7Y5_W1BEG[3] ;
 wire \Tile_X7Y5_W2BEG[0] ;
 wire \Tile_X7Y5_W2BEG[1] ;
 wire \Tile_X7Y5_W2BEG[2] ;
 wire \Tile_X7Y5_W2BEG[3] ;
 wire \Tile_X7Y5_W2BEG[4] ;
 wire \Tile_X7Y5_W2BEG[5] ;
 wire \Tile_X7Y5_W2BEG[6] ;
 wire \Tile_X7Y5_W2BEG[7] ;
 wire \Tile_X7Y5_W2BEGb[0] ;
 wire \Tile_X7Y5_W2BEGb[1] ;
 wire \Tile_X7Y5_W2BEGb[2] ;
 wire \Tile_X7Y5_W2BEGb[3] ;
 wire \Tile_X7Y5_W2BEGb[4] ;
 wire \Tile_X7Y5_W2BEGb[5] ;
 wire \Tile_X7Y5_W2BEGb[6] ;
 wire \Tile_X7Y5_W2BEGb[7] ;
 wire \Tile_X7Y5_W6BEG[0] ;
 wire \Tile_X7Y5_W6BEG[10] ;
 wire \Tile_X7Y5_W6BEG[11] ;
 wire \Tile_X7Y5_W6BEG[1] ;
 wire \Tile_X7Y5_W6BEG[2] ;
 wire \Tile_X7Y5_W6BEG[3] ;
 wire \Tile_X7Y5_W6BEG[4] ;
 wire \Tile_X7Y5_W6BEG[5] ;
 wire \Tile_X7Y5_W6BEG[6] ;
 wire \Tile_X7Y5_W6BEG[7] ;
 wire \Tile_X7Y5_W6BEG[8] ;
 wire \Tile_X7Y5_W6BEG[9] ;
 wire \Tile_X7Y5_WW4BEG[0] ;
 wire \Tile_X7Y5_WW4BEG[10] ;
 wire \Tile_X7Y5_WW4BEG[11] ;
 wire \Tile_X7Y5_WW4BEG[12] ;
 wire \Tile_X7Y5_WW4BEG[13] ;
 wire \Tile_X7Y5_WW4BEG[14] ;
 wire \Tile_X7Y5_WW4BEG[15] ;
 wire \Tile_X7Y5_WW4BEG[1] ;
 wire \Tile_X7Y5_WW4BEG[2] ;
 wire \Tile_X7Y5_WW4BEG[3] ;
 wire \Tile_X7Y5_WW4BEG[4] ;
 wire \Tile_X7Y5_WW4BEG[5] ;
 wire \Tile_X7Y5_WW4BEG[6] ;
 wire \Tile_X7Y5_WW4BEG[7] ;
 wire \Tile_X7Y5_WW4BEG[8] ;
 wire \Tile_X7Y5_WW4BEG[9] ;
 wire \Tile_X7Y6_E1BEG[0] ;
 wire \Tile_X7Y6_E1BEG[1] ;
 wire \Tile_X7Y6_E1BEG[2] ;
 wire \Tile_X7Y6_E1BEG[3] ;
 wire \Tile_X7Y6_E2BEG[0] ;
 wire \Tile_X7Y6_E2BEG[1] ;
 wire \Tile_X7Y6_E2BEG[2] ;
 wire \Tile_X7Y6_E2BEG[3] ;
 wire \Tile_X7Y6_E2BEG[4] ;
 wire \Tile_X7Y6_E2BEG[5] ;
 wire \Tile_X7Y6_E2BEG[6] ;
 wire \Tile_X7Y6_E2BEG[7] ;
 wire \Tile_X7Y6_E2BEGb[0] ;
 wire \Tile_X7Y6_E2BEGb[1] ;
 wire \Tile_X7Y6_E2BEGb[2] ;
 wire \Tile_X7Y6_E2BEGb[3] ;
 wire \Tile_X7Y6_E2BEGb[4] ;
 wire \Tile_X7Y6_E2BEGb[5] ;
 wire \Tile_X7Y6_E2BEGb[6] ;
 wire \Tile_X7Y6_E2BEGb[7] ;
 wire \Tile_X7Y6_E6BEG[0] ;
 wire \Tile_X7Y6_E6BEG[10] ;
 wire \Tile_X7Y6_E6BEG[11] ;
 wire \Tile_X7Y6_E6BEG[1] ;
 wire \Tile_X7Y6_E6BEG[2] ;
 wire \Tile_X7Y6_E6BEG[3] ;
 wire \Tile_X7Y6_E6BEG[4] ;
 wire \Tile_X7Y6_E6BEG[5] ;
 wire \Tile_X7Y6_E6BEG[6] ;
 wire \Tile_X7Y6_E6BEG[7] ;
 wire \Tile_X7Y6_E6BEG[8] ;
 wire \Tile_X7Y6_E6BEG[9] ;
 wire \Tile_X7Y6_EE4BEG[0] ;
 wire \Tile_X7Y6_EE4BEG[10] ;
 wire \Tile_X7Y6_EE4BEG[11] ;
 wire \Tile_X7Y6_EE4BEG[12] ;
 wire \Tile_X7Y6_EE4BEG[13] ;
 wire \Tile_X7Y6_EE4BEG[14] ;
 wire \Tile_X7Y6_EE4BEG[15] ;
 wire \Tile_X7Y6_EE4BEG[1] ;
 wire \Tile_X7Y6_EE4BEG[2] ;
 wire \Tile_X7Y6_EE4BEG[3] ;
 wire \Tile_X7Y6_EE4BEG[4] ;
 wire \Tile_X7Y6_EE4BEG[5] ;
 wire \Tile_X7Y6_EE4BEG[6] ;
 wire \Tile_X7Y6_EE4BEG[7] ;
 wire \Tile_X7Y6_EE4BEG[8] ;
 wire \Tile_X7Y6_EE4BEG[9] ;
 wire \Tile_X7Y6_FrameData_O[0] ;
 wire \Tile_X7Y6_FrameData_O[10] ;
 wire \Tile_X7Y6_FrameData_O[11] ;
 wire \Tile_X7Y6_FrameData_O[12] ;
 wire \Tile_X7Y6_FrameData_O[13] ;
 wire \Tile_X7Y6_FrameData_O[14] ;
 wire \Tile_X7Y6_FrameData_O[15] ;
 wire \Tile_X7Y6_FrameData_O[16] ;
 wire \Tile_X7Y6_FrameData_O[17] ;
 wire \Tile_X7Y6_FrameData_O[18] ;
 wire \Tile_X7Y6_FrameData_O[19] ;
 wire \Tile_X7Y6_FrameData_O[1] ;
 wire \Tile_X7Y6_FrameData_O[20] ;
 wire \Tile_X7Y6_FrameData_O[21] ;
 wire \Tile_X7Y6_FrameData_O[22] ;
 wire \Tile_X7Y6_FrameData_O[23] ;
 wire \Tile_X7Y6_FrameData_O[24] ;
 wire \Tile_X7Y6_FrameData_O[25] ;
 wire \Tile_X7Y6_FrameData_O[26] ;
 wire \Tile_X7Y6_FrameData_O[27] ;
 wire \Tile_X7Y6_FrameData_O[28] ;
 wire \Tile_X7Y6_FrameData_O[29] ;
 wire \Tile_X7Y6_FrameData_O[2] ;
 wire \Tile_X7Y6_FrameData_O[30] ;
 wire \Tile_X7Y6_FrameData_O[31] ;
 wire \Tile_X7Y6_FrameData_O[3] ;
 wire \Tile_X7Y6_FrameData_O[4] ;
 wire \Tile_X7Y6_FrameData_O[5] ;
 wire \Tile_X7Y6_FrameData_O[6] ;
 wire \Tile_X7Y6_FrameData_O[7] ;
 wire \Tile_X7Y6_FrameData_O[8] ;
 wire \Tile_X7Y6_FrameData_O[9] ;
 wire \Tile_X7Y6_S1BEG[0] ;
 wire \Tile_X7Y6_S1BEG[1] ;
 wire \Tile_X7Y6_S1BEG[2] ;
 wire \Tile_X7Y6_S1BEG[3] ;
 wire \Tile_X7Y6_S2BEG[0] ;
 wire \Tile_X7Y6_S2BEG[1] ;
 wire \Tile_X7Y6_S2BEG[2] ;
 wire \Tile_X7Y6_S2BEG[3] ;
 wire \Tile_X7Y6_S2BEG[4] ;
 wire \Tile_X7Y6_S2BEG[5] ;
 wire \Tile_X7Y6_S2BEG[6] ;
 wire \Tile_X7Y6_S2BEG[7] ;
 wire \Tile_X7Y6_S2BEGb[0] ;
 wire \Tile_X7Y6_S2BEGb[1] ;
 wire \Tile_X7Y6_S2BEGb[2] ;
 wire \Tile_X7Y6_S2BEGb[3] ;
 wire \Tile_X7Y6_S2BEGb[4] ;
 wire \Tile_X7Y6_S2BEGb[5] ;
 wire \Tile_X7Y6_S2BEGb[6] ;
 wire \Tile_X7Y6_S2BEGb[7] ;
 wire \Tile_X7Y6_S4BEG[0] ;
 wire \Tile_X7Y6_S4BEG[10] ;
 wire \Tile_X7Y6_S4BEG[11] ;
 wire \Tile_X7Y6_S4BEG[12] ;
 wire \Tile_X7Y6_S4BEG[13] ;
 wire \Tile_X7Y6_S4BEG[14] ;
 wire \Tile_X7Y6_S4BEG[15] ;
 wire \Tile_X7Y6_S4BEG[1] ;
 wire \Tile_X7Y6_S4BEG[2] ;
 wire \Tile_X7Y6_S4BEG[3] ;
 wire \Tile_X7Y6_S4BEG[4] ;
 wire \Tile_X7Y6_S4BEG[5] ;
 wire \Tile_X7Y6_S4BEG[6] ;
 wire \Tile_X7Y6_S4BEG[7] ;
 wire \Tile_X7Y6_S4BEG[8] ;
 wire \Tile_X7Y6_S4BEG[9] ;
 wire \Tile_X7Y6_SS4BEG[0] ;
 wire \Tile_X7Y6_SS4BEG[10] ;
 wire \Tile_X7Y6_SS4BEG[11] ;
 wire \Tile_X7Y6_SS4BEG[12] ;
 wire \Tile_X7Y6_SS4BEG[13] ;
 wire \Tile_X7Y6_SS4BEG[14] ;
 wire \Tile_X7Y6_SS4BEG[15] ;
 wire \Tile_X7Y6_SS4BEG[1] ;
 wire \Tile_X7Y6_SS4BEG[2] ;
 wire \Tile_X7Y6_SS4BEG[3] ;
 wire \Tile_X7Y6_SS4BEG[4] ;
 wire \Tile_X7Y6_SS4BEG[5] ;
 wire \Tile_X7Y6_SS4BEG[6] ;
 wire \Tile_X7Y6_SS4BEG[7] ;
 wire \Tile_X7Y6_SS4BEG[8] ;
 wire \Tile_X7Y6_SS4BEG[9] ;
 wire \Tile_X7Y6_W1BEG[0] ;
 wire \Tile_X7Y6_W1BEG[1] ;
 wire \Tile_X7Y6_W1BEG[2] ;
 wire \Tile_X7Y6_W1BEG[3] ;
 wire \Tile_X7Y6_W2BEG[0] ;
 wire \Tile_X7Y6_W2BEG[1] ;
 wire \Tile_X7Y6_W2BEG[2] ;
 wire \Tile_X7Y6_W2BEG[3] ;
 wire \Tile_X7Y6_W2BEG[4] ;
 wire \Tile_X7Y6_W2BEG[5] ;
 wire \Tile_X7Y6_W2BEG[6] ;
 wire \Tile_X7Y6_W2BEG[7] ;
 wire \Tile_X7Y6_W2BEGb[0] ;
 wire \Tile_X7Y6_W2BEGb[1] ;
 wire \Tile_X7Y6_W2BEGb[2] ;
 wire \Tile_X7Y6_W2BEGb[3] ;
 wire \Tile_X7Y6_W2BEGb[4] ;
 wire \Tile_X7Y6_W2BEGb[5] ;
 wire \Tile_X7Y6_W2BEGb[6] ;
 wire \Tile_X7Y6_W2BEGb[7] ;
 wire \Tile_X7Y6_W6BEG[0] ;
 wire \Tile_X7Y6_W6BEG[10] ;
 wire \Tile_X7Y6_W6BEG[11] ;
 wire \Tile_X7Y6_W6BEG[1] ;
 wire \Tile_X7Y6_W6BEG[2] ;
 wire \Tile_X7Y6_W6BEG[3] ;
 wire \Tile_X7Y6_W6BEG[4] ;
 wire \Tile_X7Y6_W6BEG[5] ;
 wire \Tile_X7Y6_W6BEG[6] ;
 wire \Tile_X7Y6_W6BEG[7] ;
 wire \Tile_X7Y6_W6BEG[8] ;
 wire \Tile_X7Y6_W6BEG[9] ;
 wire \Tile_X7Y6_WW4BEG[0] ;
 wire \Tile_X7Y6_WW4BEG[10] ;
 wire \Tile_X7Y6_WW4BEG[11] ;
 wire \Tile_X7Y6_WW4BEG[12] ;
 wire \Tile_X7Y6_WW4BEG[13] ;
 wire \Tile_X7Y6_WW4BEG[14] ;
 wire \Tile_X7Y6_WW4BEG[15] ;
 wire \Tile_X7Y6_WW4BEG[1] ;
 wire \Tile_X7Y6_WW4BEG[2] ;
 wire \Tile_X7Y6_WW4BEG[3] ;
 wire \Tile_X7Y6_WW4BEG[4] ;
 wire \Tile_X7Y6_WW4BEG[5] ;
 wire \Tile_X7Y6_WW4BEG[6] ;
 wire \Tile_X7Y6_WW4BEG[7] ;
 wire \Tile_X7Y6_WW4BEG[8] ;
 wire \Tile_X7Y6_WW4BEG[9] ;
 wire \Tile_X7Y7_E1BEG[0] ;
 wire \Tile_X7Y7_E1BEG[1] ;
 wire \Tile_X7Y7_E1BEG[2] ;
 wire \Tile_X7Y7_E1BEG[3] ;
 wire \Tile_X7Y7_E2BEG[0] ;
 wire \Tile_X7Y7_E2BEG[1] ;
 wire \Tile_X7Y7_E2BEG[2] ;
 wire \Tile_X7Y7_E2BEG[3] ;
 wire \Tile_X7Y7_E2BEG[4] ;
 wire \Tile_X7Y7_E2BEG[5] ;
 wire \Tile_X7Y7_E2BEG[6] ;
 wire \Tile_X7Y7_E2BEG[7] ;
 wire \Tile_X7Y7_E2BEGb[0] ;
 wire \Tile_X7Y7_E2BEGb[1] ;
 wire \Tile_X7Y7_E2BEGb[2] ;
 wire \Tile_X7Y7_E2BEGb[3] ;
 wire \Tile_X7Y7_E2BEGb[4] ;
 wire \Tile_X7Y7_E2BEGb[5] ;
 wire \Tile_X7Y7_E2BEGb[6] ;
 wire \Tile_X7Y7_E2BEGb[7] ;
 wire \Tile_X7Y7_E6BEG[0] ;
 wire \Tile_X7Y7_E6BEG[10] ;
 wire \Tile_X7Y7_E6BEG[11] ;
 wire \Tile_X7Y7_E6BEG[1] ;
 wire \Tile_X7Y7_E6BEG[2] ;
 wire \Tile_X7Y7_E6BEG[3] ;
 wire \Tile_X7Y7_E6BEG[4] ;
 wire \Tile_X7Y7_E6BEG[5] ;
 wire \Tile_X7Y7_E6BEG[6] ;
 wire \Tile_X7Y7_E6BEG[7] ;
 wire \Tile_X7Y7_E6BEG[8] ;
 wire \Tile_X7Y7_E6BEG[9] ;
 wire \Tile_X7Y7_EE4BEG[0] ;
 wire \Tile_X7Y7_EE4BEG[10] ;
 wire \Tile_X7Y7_EE4BEG[11] ;
 wire \Tile_X7Y7_EE4BEG[12] ;
 wire \Tile_X7Y7_EE4BEG[13] ;
 wire \Tile_X7Y7_EE4BEG[14] ;
 wire \Tile_X7Y7_EE4BEG[15] ;
 wire \Tile_X7Y7_EE4BEG[1] ;
 wire \Tile_X7Y7_EE4BEG[2] ;
 wire \Tile_X7Y7_EE4BEG[3] ;
 wire \Tile_X7Y7_EE4BEG[4] ;
 wire \Tile_X7Y7_EE4BEG[5] ;
 wire \Tile_X7Y7_EE4BEG[6] ;
 wire \Tile_X7Y7_EE4BEG[7] ;
 wire \Tile_X7Y7_EE4BEG[8] ;
 wire \Tile_X7Y7_EE4BEG[9] ;
 wire \Tile_X7Y7_FrameData_O[0] ;
 wire \Tile_X7Y7_FrameData_O[10] ;
 wire \Tile_X7Y7_FrameData_O[11] ;
 wire \Tile_X7Y7_FrameData_O[12] ;
 wire \Tile_X7Y7_FrameData_O[13] ;
 wire \Tile_X7Y7_FrameData_O[14] ;
 wire \Tile_X7Y7_FrameData_O[15] ;
 wire \Tile_X7Y7_FrameData_O[16] ;
 wire \Tile_X7Y7_FrameData_O[17] ;
 wire \Tile_X7Y7_FrameData_O[18] ;
 wire \Tile_X7Y7_FrameData_O[19] ;
 wire \Tile_X7Y7_FrameData_O[1] ;
 wire \Tile_X7Y7_FrameData_O[20] ;
 wire \Tile_X7Y7_FrameData_O[21] ;
 wire \Tile_X7Y7_FrameData_O[22] ;
 wire \Tile_X7Y7_FrameData_O[23] ;
 wire \Tile_X7Y7_FrameData_O[24] ;
 wire \Tile_X7Y7_FrameData_O[25] ;
 wire \Tile_X7Y7_FrameData_O[26] ;
 wire \Tile_X7Y7_FrameData_O[27] ;
 wire \Tile_X7Y7_FrameData_O[28] ;
 wire \Tile_X7Y7_FrameData_O[29] ;
 wire \Tile_X7Y7_FrameData_O[2] ;
 wire \Tile_X7Y7_FrameData_O[30] ;
 wire \Tile_X7Y7_FrameData_O[31] ;
 wire \Tile_X7Y7_FrameData_O[3] ;
 wire \Tile_X7Y7_FrameData_O[4] ;
 wire \Tile_X7Y7_FrameData_O[5] ;
 wire \Tile_X7Y7_FrameData_O[6] ;
 wire \Tile_X7Y7_FrameData_O[7] ;
 wire \Tile_X7Y7_FrameData_O[8] ;
 wire \Tile_X7Y7_FrameData_O[9] ;
 wire \Tile_X7Y7_FrameStrobe_O[0] ;
 wire \Tile_X7Y7_FrameStrobe_O[10] ;
 wire \Tile_X7Y7_FrameStrobe_O[11] ;
 wire \Tile_X7Y7_FrameStrobe_O[12] ;
 wire \Tile_X7Y7_FrameStrobe_O[13] ;
 wire \Tile_X7Y7_FrameStrobe_O[14] ;
 wire \Tile_X7Y7_FrameStrobe_O[15] ;
 wire \Tile_X7Y7_FrameStrobe_O[16] ;
 wire \Tile_X7Y7_FrameStrobe_O[17] ;
 wire \Tile_X7Y7_FrameStrobe_O[18] ;
 wire \Tile_X7Y7_FrameStrobe_O[19] ;
 wire \Tile_X7Y7_FrameStrobe_O[1] ;
 wire \Tile_X7Y7_FrameStrobe_O[2] ;
 wire \Tile_X7Y7_FrameStrobe_O[3] ;
 wire \Tile_X7Y7_FrameStrobe_O[4] ;
 wire \Tile_X7Y7_FrameStrobe_O[5] ;
 wire \Tile_X7Y7_FrameStrobe_O[6] ;
 wire \Tile_X7Y7_FrameStrobe_O[7] ;
 wire \Tile_X7Y7_FrameStrobe_O[8] ;
 wire \Tile_X7Y7_FrameStrobe_O[9] ;
 wire \Tile_X7Y7_N1BEG[0] ;
 wire \Tile_X7Y7_N1BEG[1] ;
 wire \Tile_X7Y7_N1BEG[2] ;
 wire \Tile_X7Y7_N1BEG[3] ;
 wire \Tile_X7Y7_N2BEG[0] ;
 wire \Tile_X7Y7_N2BEG[1] ;
 wire \Tile_X7Y7_N2BEG[2] ;
 wire \Tile_X7Y7_N2BEG[3] ;
 wire \Tile_X7Y7_N2BEG[4] ;
 wire \Tile_X7Y7_N2BEG[5] ;
 wire \Tile_X7Y7_N2BEG[6] ;
 wire \Tile_X7Y7_N2BEG[7] ;
 wire \Tile_X7Y7_N2BEGb[0] ;
 wire \Tile_X7Y7_N2BEGb[1] ;
 wire \Tile_X7Y7_N2BEGb[2] ;
 wire \Tile_X7Y7_N2BEGb[3] ;
 wire \Tile_X7Y7_N2BEGb[4] ;
 wire \Tile_X7Y7_N2BEGb[5] ;
 wire \Tile_X7Y7_N2BEGb[6] ;
 wire \Tile_X7Y7_N2BEGb[7] ;
 wire \Tile_X7Y7_N4BEG[0] ;
 wire \Tile_X7Y7_N4BEG[10] ;
 wire \Tile_X7Y7_N4BEG[11] ;
 wire \Tile_X7Y7_N4BEG[12] ;
 wire \Tile_X7Y7_N4BEG[13] ;
 wire \Tile_X7Y7_N4BEG[14] ;
 wire \Tile_X7Y7_N4BEG[15] ;
 wire \Tile_X7Y7_N4BEG[1] ;
 wire \Tile_X7Y7_N4BEG[2] ;
 wire \Tile_X7Y7_N4BEG[3] ;
 wire \Tile_X7Y7_N4BEG[4] ;
 wire \Tile_X7Y7_N4BEG[5] ;
 wire \Tile_X7Y7_N4BEG[6] ;
 wire \Tile_X7Y7_N4BEG[7] ;
 wire \Tile_X7Y7_N4BEG[8] ;
 wire \Tile_X7Y7_N4BEG[9] ;
 wire \Tile_X7Y7_NN4BEG[0] ;
 wire \Tile_X7Y7_NN4BEG[10] ;
 wire \Tile_X7Y7_NN4BEG[11] ;
 wire \Tile_X7Y7_NN4BEG[12] ;
 wire \Tile_X7Y7_NN4BEG[13] ;
 wire \Tile_X7Y7_NN4BEG[14] ;
 wire \Tile_X7Y7_NN4BEG[15] ;
 wire \Tile_X7Y7_NN4BEG[1] ;
 wire \Tile_X7Y7_NN4BEG[2] ;
 wire \Tile_X7Y7_NN4BEG[3] ;
 wire \Tile_X7Y7_NN4BEG[4] ;
 wire \Tile_X7Y7_NN4BEG[5] ;
 wire \Tile_X7Y7_NN4BEG[6] ;
 wire \Tile_X7Y7_NN4BEG[7] ;
 wire \Tile_X7Y7_NN4BEG[8] ;
 wire \Tile_X7Y7_NN4BEG[9] ;
 wire Tile_X7Y7_UserCLKo;
 wire \Tile_X7Y7_W1BEG[0] ;
 wire \Tile_X7Y7_W1BEG[1] ;
 wire \Tile_X7Y7_W1BEG[2] ;
 wire \Tile_X7Y7_W1BEG[3] ;
 wire \Tile_X7Y7_W2BEG[0] ;
 wire \Tile_X7Y7_W2BEG[1] ;
 wire \Tile_X7Y7_W2BEG[2] ;
 wire \Tile_X7Y7_W2BEG[3] ;
 wire \Tile_X7Y7_W2BEG[4] ;
 wire \Tile_X7Y7_W2BEG[5] ;
 wire \Tile_X7Y7_W2BEG[6] ;
 wire \Tile_X7Y7_W2BEG[7] ;
 wire \Tile_X7Y7_W2BEGb[0] ;
 wire \Tile_X7Y7_W2BEGb[1] ;
 wire \Tile_X7Y7_W2BEGb[2] ;
 wire \Tile_X7Y7_W2BEGb[3] ;
 wire \Tile_X7Y7_W2BEGb[4] ;
 wire \Tile_X7Y7_W2BEGb[5] ;
 wire \Tile_X7Y7_W2BEGb[6] ;
 wire \Tile_X7Y7_W2BEGb[7] ;
 wire \Tile_X7Y7_W6BEG[0] ;
 wire \Tile_X7Y7_W6BEG[10] ;
 wire \Tile_X7Y7_W6BEG[11] ;
 wire \Tile_X7Y7_W6BEG[1] ;
 wire \Tile_X7Y7_W6BEG[2] ;
 wire \Tile_X7Y7_W6BEG[3] ;
 wire \Tile_X7Y7_W6BEG[4] ;
 wire \Tile_X7Y7_W6BEG[5] ;
 wire \Tile_X7Y7_W6BEG[6] ;
 wire \Tile_X7Y7_W6BEG[7] ;
 wire \Tile_X7Y7_W6BEG[8] ;
 wire \Tile_X7Y7_W6BEG[9] ;
 wire \Tile_X7Y7_WW4BEG[0] ;
 wire \Tile_X7Y7_WW4BEG[10] ;
 wire \Tile_X7Y7_WW4BEG[11] ;
 wire \Tile_X7Y7_WW4BEG[12] ;
 wire \Tile_X7Y7_WW4BEG[13] ;
 wire \Tile_X7Y7_WW4BEG[14] ;
 wire \Tile_X7Y7_WW4BEG[15] ;
 wire \Tile_X7Y7_WW4BEG[1] ;
 wire \Tile_X7Y7_WW4BEG[2] ;
 wire \Tile_X7Y7_WW4BEG[3] ;
 wire \Tile_X7Y7_WW4BEG[4] ;
 wire \Tile_X7Y7_WW4BEG[5] ;
 wire \Tile_X7Y7_WW4BEG[6] ;
 wire \Tile_X7Y7_WW4BEG[7] ;
 wire \Tile_X7Y7_WW4BEG[8] ;
 wire \Tile_X7Y7_WW4BEG[9] ;
 wire \Tile_X7Y8_E1BEG[0] ;
 wire \Tile_X7Y8_E1BEG[1] ;
 wire \Tile_X7Y8_E1BEG[2] ;
 wire \Tile_X7Y8_E1BEG[3] ;
 wire \Tile_X7Y8_E2BEG[0] ;
 wire \Tile_X7Y8_E2BEG[1] ;
 wire \Tile_X7Y8_E2BEG[2] ;
 wire \Tile_X7Y8_E2BEG[3] ;
 wire \Tile_X7Y8_E2BEG[4] ;
 wire \Tile_X7Y8_E2BEG[5] ;
 wire \Tile_X7Y8_E2BEG[6] ;
 wire \Tile_X7Y8_E2BEG[7] ;
 wire \Tile_X7Y8_E2BEGb[0] ;
 wire \Tile_X7Y8_E2BEGb[1] ;
 wire \Tile_X7Y8_E2BEGb[2] ;
 wire \Tile_X7Y8_E2BEGb[3] ;
 wire \Tile_X7Y8_E2BEGb[4] ;
 wire \Tile_X7Y8_E2BEGb[5] ;
 wire \Tile_X7Y8_E2BEGb[6] ;
 wire \Tile_X7Y8_E2BEGb[7] ;
 wire \Tile_X7Y8_E6BEG[0] ;
 wire \Tile_X7Y8_E6BEG[10] ;
 wire \Tile_X7Y8_E6BEG[11] ;
 wire \Tile_X7Y8_E6BEG[1] ;
 wire \Tile_X7Y8_E6BEG[2] ;
 wire \Tile_X7Y8_E6BEG[3] ;
 wire \Tile_X7Y8_E6BEG[4] ;
 wire \Tile_X7Y8_E6BEG[5] ;
 wire \Tile_X7Y8_E6BEG[6] ;
 wire \Tile_X7Y8_E6BEG[7] ;
 wire \Tile_X7Y8_E6BEG[8] ;
 wire \Tile_X7Y8_E6BEG[9] ;
 wire \Tile_X7Y8_EE4BEG[0] ;
 wire \Tile_X7Y8_EE4BEG[10] ;
 wire \Tile_X7Y8_EE4BEG[11] ;
 wire \Tile_X7Y8_EE4BEG[12] ;
 wire \Tile_X7Y8_EE4BEG[13] ;
 wire \Tile_X7Y8_EE4BEG[14] ;
 wire \Tile_X7Y8_EE4BEG[15] ;
 wire \Tile_X7Y8_EE4BEG[1] ;
 wire \Tile_X7Y8_EE4BEG[2] ;
 wire \Tile_X7Y8_EE4BEG[3] ;
 wire \Tile_X7Y8_EE4BEG[4] ;
 wire \Tile_X7Y8_EE4BEG[5] ;
 wire \Tile_X7Y8_EE4BEG[6] ;
 wire \Tile_X7Y8_EE4BEG[7] ;
 wire \Tile_X7Y8_EE4BEG[8] ;
 wire \Tile_X7Y8_EE4BEG[9] ;
 wire \Tile_X7Y8_FrameData_O[0] ;
 wire \Tile_X7Y8_FrameData_O[10] ;
 wire \Tile_X7Y8_FrameData_O[11] ;
 wire \Tile_X7Y8_FrameData_O[12] ;
 wire \Tile_X7Y8_FrameData_O[13] ;
 wire \Tile_X7Y8_FrameData_O[14] ;
 wire \Tile_X7Y8_FrameData_O[15] ;
 wire \Tile_X7Y8_FrameData_O[16] ;
 wire \Tile_X7Y8_FrameData_O[17] ;
 wire \Tile_X7Y8_FrameData_O[18] ;
 wire \Tile_X7Y8_FrameData_O[19] ;
 wire \Tile_X7Y8_FrameData_O[1] ;
 wire \Tile_X7Y8_FrameData_O[20] ;
 wire \Tile_X7Y8_FrameData_O[21] ;
 wire \Tile_X7Y8_FrameData_O[22] ;
 wire \Tile_X7Y8_FrameData_O[23] ;
 wire \Tile_X7Y8_FrameData_O[24] ;
 wire \Tile_X7Y8_FrameData_O[25] ;
 wire \Tile_X7Y8_FrameData_O[26] ;
 wire \Tile_X7Y8_FrameData_O[27] ;
 wire \Tile_X7Y8_FrameData_O[28] ;
 wire \Tile_X7Y8_FrameData_O[29] ;
 wire \Tile_X7Y8_FrameData_O[2] ;
 wire \Tile_X7Y8_FrameData_O[30] ;
 wire \Tile_X7Y8_FrameData_O[31] ;
 wire \Tile_X7Y8_FrameData_O[3] ;
 wire \Tile_X7Y8_FrameData_O[4] ;
 wire \Tile_X7Y8_FrameData_O[5] ;
 wire \Tile_X7Y8_FrameData_O[6] ;
 wire \Tile_X7Y8_FrameData_O[7] ;
 wire \Tile_X7Y8_FrameData_O[8] ;
 wire \Tile_X7Y8_FrameData_O[9] ;
 wire \Tile_X7Y8_S1BEG[0] ;
 wire \Tile_X7Y8_S1BEG[1] ;
 wire \Tile_X7Y8_S1BEG[2] ;
 wire \Tile_X7Y8_S1BEG[3] ;
 wire \Tile_X7Y8_S2BEG[0] ;
 wire \Tile_X7Y8_S2BEG[1] ;
 wire \Tile_X7Y8_S2BEG[2] ;
 wire \Tile_X7Y8_S2BEG[3] ;
 wire \Tile_X7Y8_S2BEG[4] ;
 wire \Tile_X7Y8_S2BEG[5] ;
 wire \Tile_X7Y8_S2BEG[6] ;
 wire \Tile_X7Y8_S2BEG[7] ;
 wire \Tile_X7Y8_S2BEGb[0] ;
 wire \Tile_X7Y8_S2BEGb[1] ;
 wire \Tile_X7Y8_S2BEGb[2] ;
 wire \Tile_X7Y8_S2BEGb[3] ;
 wire \Tile_X7Y8_S2BEGb[4] ;
 wire \Tile_X7Y8_S2BEGb[5] ;
 wire \Tile_X7Y8_S2BEGb[6] ;
 wire \Tile_X7Y8_S2BEGb[7] ;
 wire \Tile_X7Y8_S4BEG[0] ;
 wire \Tile_X7Y8_S4BEG[10] ;
 wire \Tile_X7Y8_S4BEG[11] ;
 wire \Tile_X7Y8_S4BEG[12] ;
 wire \Tile_X7Y8_S4BEG[13] ;
 wire \Tile_X7Y8_S4BEG[14] ;
 wire \Tile_X7Y8_S4BEG[15] ;
 wire \Tile_X7Y8_S4BEG[1] ;
 wire \Tile_X7Y8_S4BEG[2] ;
 wire \Tile_X7Y8_S4BEG[3] ;
 wire \Tile_X7Y8_S4BEG[4] ;
 wire \Tile_X7Y8_S4BEG[5] ;
 wire \Tile_X7Y8_S4BEG[6] ;
 wire \Tile_X7Y8_S4BEG[7] ;
 wire \Tile_X7Y8_S4BEG[8] ;
 wire \Tile_X7Y8_S4BEG[9] ;
 wire \Tile_X7Y8_SS4BEG[0] ;
 wire \Tile_X7Y8_SS4BEG[10] ;
 wire \Tile_X7Y8_SS4BEG[11] ;
 wire \Tile_X7Y8_SS4BEG[12] ;
 wire \Tile_X7Y8_SS4BEG[13] ;
 wire \Tile_X7Y8_SS4BEG[14] ;
 wire \Tile_X7Y8_SS4BEG[15] ;
 wire \Tile_X7Y8_SS4BEG[1] ;
 wire \Tile_X7Y8_SS4BEG[2] ;
 wire \Tile_X7Y8_SS4BEG[3] ;
 wire \Tile_X7Y8_SS4BEG[4] ;
 wire \Tile_X7Y8_SS4BEG[5] ;
 wire \Tile_X7Y8_SS4BEG[6] ;
 wire \Tile_X7Y8_SS4BEG[7] ;
 wire \Tile_X7Y8_SS4BEG[8] ;
 wire \Tile_X7Y8_SS4BEG[9] ;
 wire \Tile_X7Y8_W1BEG[0] ;
 wire \Tile_X7Y8_W1BEG[1] ;
 wire \Tile_X7Y8_W1BEG[2] ;
 wire \Tile_X7Y8_W1BEG[3] ;
 wire \Tile_X7Y8_W2BEG[0] ;
 wire \Tile_X7Y8_W2BEG[1] ;
 wire \Tile_X7Y8_W2BEG[2] ;
 wire \Tile_X7Y8_W2BEG[3] ;
 wire \Tile_X7Y8_W2BEG[4] ;
 wire \Tile_X7Y8_W2BEG[5] ;
 wire \Tile_X7Y8_W2BEG[6] ;
 wire \Tile_X7Y8_W2BEG[7] ;
 wire \Tile_X7Y8_W2BEGb[0] ;
 wire \Tile_X7Y8_W2BEGb[1] ;
 wire \Tile_X7Y8_W2BEGb[2] ;
 wire \Tile_X7Y8_W2BEGb[3] ;
 wire \Tile_X7Y8_W2BEGb[4] ;
 wire \Tile_X7Y8_W2BEGb[5] ;
 wire \Tile_X7Y8_W2BEGb[6] ;
 wire \Tile_X7Y8_W2BEGb[7] ;
 wire \Tile_X7Y8_W6BEG[0] ;
 wire \Tile_X7Y8_W6BEG[10] ;
 wire \Tile_X7Y8_W6BEG[11] ;
 wire \Tile_X7Y8_W6BEG[1] ;
 wire \Tile_X7Y8_W6BEG[2] ;
 wire \Tile_X7Y8_W6BEG[3] ;
 wire \Tile_X7Y8_W6BEG[4] ;
 wire \Tile_X7Y8_W6BEG[5] ;
 wire \Tile_X7Y8_W6BEG[6] ;
 wire \Tile_X7Y8_W6BEG[7] ;
 wire \Tile_X7Y8_W6BEG[8] ;
 wire \Tile_X7Y8_W6BEG[9] ;
 wire \Tile_X7Y8_WW4BEG[0] ;
 wire \Tile_X7Y8_WW4BEG[10] ;
 wire \Tile_X7Y8_WW4BEG[11] ;
 wire \Tile_X7Y8_WW4BEG[12] ;
 wire \Tile_X7Y8_WW4BEG[13] ;
 wire \Tile_X7Y8_WW4BEG[14] ;
 wire \Tile_X7Y8_WW4BEG[15] ;
 wire \Tile_X7Y8_WW4BEG[1] ;
 wire \Tile_X7Y8_WW4BEG[2] ;
 wire \Tile_X7Y8_WW4BEG[3] ;
 wire \Tile_X7Y8_WW4BEG[4] ;
 wire \Tile_X7Y8_WW4BEG[5] ;
 wire \Tile_X7Y8_WW4BEG[6] ;
 wire \Tile_X7Y8_WW4BEG[7] ;
 wire \Tile_X7Y8_WW4BEG[8] ;
 wire \Tile_X7Y8_WW4BEG[9] ;
 wire \Tile_X7Y9_E1BEG[0] ;
 wire \Tile_X7Y9_E1BEG[1] ;
 wire \Tile_X7Y9_E1BEG[2] ;
 wire \Tile_X7Y9_E1BEG[3] ;
 wire \Tile_X7Y9_E2BEG[0] ;
 wire \Tile_X7Y9_E2BEG[1] ;
 wire \Tile_X7Y9_E2BEG[2] ;
 wire \Tile_X7Y9_E2BEG[3] ;
 wire \Tile_X7Y9_E2BEG[4] ;
 wire \Tile_X7Y9_E2BEG[5] ;
 wire \Tile_X7Y9_E2BEG[6] ;
 wire \Tile_X7Y9_E2BEG[7] ;
 wire \Tile_X7Y9_E2BEGb[0] ;
 wire \Tile_X7Y9_E2BEGb[1] ;
 wire \Tile_X7Y9_E2BEGb[2] ;
 wire \Tile_X7Y9_E2BEGb[3] ;
 wire \Tile_X7Y9_E2BEGb[4] ;
 wire \Tile_X7Y9_E2BEGb[5] ;
 wire \Tile_X7Y9_E2BEGb[6] ;
 wire \Tile_X7Y9_E2BEGb[7] ;
 wire \Tile_X7Y9_E6BEG[0] ;
 wire \Tile_X7Y9_E6BEG[10] ;
 wire \Tile_X7Y9_E6BEG[11] ;
 wire \Tile_X7Y9_E6BEG[1] ;
 wire \Tile_X7Y9_E6BEG[2] ;
 wire \Tile_X7Y9_E6BEG[3] ;
 wire \Tile_X7Y9_E6BEG[4] ;
 wire \Tile_X7Y9_E6BEG[5] ;
 wire \Tile_X7Y9_E6BEG[6] ;
 wire \Tile_X7Y9_E6BEG[7] ;
 wire \Tile_X7Y9_E6BEG[8] ;
 wire \Tile_X7Y9_E6BEG[9] ;
 wire \Tile_X7Y9_EE4BEG[0] ;
 wire \Tile_X7Y9_EE4BEG[10] ;
 wire \Tile_X7Y9_EE4BEG[11] ;
 wire \Tile_X7Y9_EE4BEG[12] ;
 wire \Tile_X7Y9_EE4BEG[13] ;
 wire \Tile_X7Y9_EE4BEG[14] ;
 wire \Tile_X7Y9_EE4BEG[15] ;
 wire \Tile_X7Y9_EE4BEG[1] ;
 wire \Tile_X7Y9_EE4BEG[2] ;
 wire \Tile_X7Y9_EE4BEG[3] ;
 wire \Tile_X7Y9_EE4BEG[4] ;
 wire \Tile_X7Y9_EE4BEG[5] ;
 wire \Tile_X7Y9_EE4BEG[6] ;
 wire \Tile_X7Y9_EE4BEG[7] ;
 wire \Tile_X7Y9_EE4BEG[8] ;
 wire \Tile_X7Y9_EE4BEG[9] ;
 wire \Tile_X7Y9_FrameData_O[0] ;
 wire \Tile_X7Y9_FrameData_O[10] ;
 wire \Tile_X7Y9_FrameData_O[11] ;
 wire \Tile_X7Y9_FrameData_O[12] ;
 wire \Tile_X7Y9_FrameData_O[13] ;
 wire \Tile_X7Y9_FrameData_O[14] ;
 wire \Tile_X7Y9_FrameData_O[15] ;
 wire \Tile_X7Y9_FrameData_O[16] ;
 wire \Tile_X7Y9_FrameData_O[17] ;
 wire \Tile_X7Y9_FrameData_O[18] ;
 wire \Tile_X7Y9_FrameData_O[19] ;
 wire \Tile_X7Y9_FrameData_O[1] ;
 wire \Tile_X7Y9_FrameData_O[20] ;
 wire \Tile_X7Y9_FrameData_O[21] ;
 wire \Tile_X7Y9_FrameData_O[22] ;
 wire \Tile_X7Y9_FrameData_O[23] ;
 wire \Tile_X7Y9_FrameData_O[24] ;
 wire \Tile_X7Y9_FrameData_O[25] ;
 wire \Tile_X7Y9_FrameData_O[26] ;
 wire \Tile_X7Y9_FrameData_O[27] ;
 wire \Tile_X7Y9_FrameData_O[28] ;
 wire \Tile_X7Y9_FrameData_O[29] ;
 wire \Tile_X7Y9_FrameData_O[2] ;
 wire \Tile_X7Y9_FrameData_O[30] ;
 wire \Tile_X7Y9_FrameData_O[31] ;
 wire \Tile_X7Y9_FrameData_O[3] ;
 wire \Tile_X7Y9_FrameData_O[4] ;
 wire \Tile_X7Y9_FrameData_O[5] ;
 wire \Tile_X7Y9_FrameData_O[6] ;
 wire \Tile_X7Y9_FrameData_O[7] ;
 wire \Tile_X7Y9_FrameData_O[8] ;
 wire \Tile_X7Y9_FrameData_O[9] ;
 wire \Tile_X7Y9_FrameStrobe_O[0] ;
 wire \Tile_X7Y9_FrameStrobe_O[10] ;
 wire \Tile_X7Y9_FrameStrobe_O[11] ;
 wire \Tile_X7Y9_FrameStrobe_O[12] ;
 wire \Tile_X7Y9_FrameStrobe_O[13] ;
 wire \Tile_X7Y9_FrameStrobe_O[14] ;
 wire \Tile_X7Y9_FrameStrobe_O[15] ;
 wire \Tile_X7Y9_FrameStrobe_O[16] ;
 wire \Tile_X7Y9_FrameStrobe_O[17] ;
 wire \Tile_X7Y9_FrameStrobe_O[18] ;
 wire \Tile_X7Y9_FrameStrobe_O[19] ;
 wire \Tile_X7Y9_FrameStrobe_O[1] ;
 wire \Tile_X7Y9_FrameStrobe_O[2] ;
 wire \Tile_X7Y9_FrameStrobe_O[3] ;
 wire \Tile_X7Y9_FrameStrobe_O[4] ;
 wire \Tile_X7Y9_FrameStrobe_O[5] ;
 wire \Tile_X7Y9_FrameStrobe_O[6] ;
 wire \Tile_X7Y9_FrameStrobe_O[7] ;
 wire \Tile_X7Y9_FrameStrobe_O[8] ;
 wire \Tile_X7Y9_FrameStrobe_O[9] ;
 wire \Tile_X7Y9_N1BEG[0] ;
 wire \Tile_X7Y9_N1BEG[1] ;
 wire \Tile_X7Y9_N1BEG[2] ;
 wire \Tile_X7Y9_N1BEG[3] ;
 wire \Tile_X7Y9_N2BEG[0] ;
 wire \Tile_X7Y9_N2BEG[1] ;
 wire \Tile_X7Y9_N2BEG[2] ;
 wire \Tile_X7Y9_N2BEG[3] ;
 wire \Tile_X7Y9_N2BEG[4] ;
 wire \Tile_X7Y9_N2BEG[5] ;
 wire \Tile_X7Y9_N2BEG[6] ;
 wire \Tile_X7Y9_N2BEG[7] ;
 wire \Tile_X7Y9_N2BEGb[0] ;
 wire \Tile_X7Y9_N2BEGb[1] ;
 wire \Tile_X7Y9_N2BEGb[2] ;
 wire \Tile_X7Y9_N2BEGb[3] ;
 wire \Tile_X7Y9_N2BEGb[4] ;
 wire \Tile_X7Y9_N2BEGb[5] ;
 wire \Tile_X7Y9_N2BEGb[6] ;
 wire \Tile_X7Y9_N2BEGb[7] ;
 wire \Tile_X7Y9_N4BEG[0] ;
 wire \Tile_X7Y9_N4BEG[10] ;
 wire \Tile_X7Y9_N4BEG[11] ;
 wire \Tile_X7Y9_N4BEG[12] ;
 wire \Tile_X7Y9_N4BEG[13] ;
 wire \Tile_X7Y9_N4BEG[14] ;
 wire \Tile_X7Y9_N4BEG[15] ;
 wire \Tile_X7Y9_N4BEG[1] ;
 wire \Tile_X7Y9_N4BEG[2] ;
 wire \Tile_X7Y9_N4BEG[3] ;
 wire \Tile_X7Y9_N4BEG[4] ;
 wire \Tile_X7Y9_N4BEG[5] ;
 wire \Tile_X7Y9_N4BEG[6] ;
 wire \Tile_X7Y9_N4BEG[7] ;
 wire \Tile_X7Y9_N4BEG[8] ;
 wire \Tile_X7Y9_N4BEG[9] ;
 wire \Tile_X7Y9_NN4BEG[0] ;
 wire \Tile_X7Y9_NN4BEG[10] ;
 wire \Tile_X7Y9_NN4BEG[11] ;
 wire \Tile_X7Y9_NN4BEG[12] ;
 wire \Tile_X7Y9_NN4BEG[13] ;
 wire \Tile_X7Y9_NN4BEG[14] ;
 wire \Tile_X7Y9_NN4BEG[15] ;
 wire \Tile_X7Y9_NN4BEG[1] ;
 wire \Tile_X7Y9_NN4BEG[2] ;
 wire \Tile_X7Y9_NN4BEG[3] ;
 wire \Tile_X7Y9_NN4BEG[4] ;
 wire \Tile_X7Y9_NN4BEG[5] ;
 wire \Tile_X7Y9_NN4BEG[6] ;
 wire \Tile_X7Y9_NN4BEG[7] ;
 wire \Tile_X7Y9_NN4BEG[8] ;
 wire \Tile_X7Y9_NN4BEG[9] ;
 wire Tile_X7Y9_UserCLKo;
 wire \Tile_X7Y9_W1BEG[0] ;
 wire \Tile_X7Y9_W1BEG[1] ;
 wire \Tile_X7Y9_W1BEG[2] ;
 wire \Tile_X7Y9_W1BEG[3] ;
 wire \Tile_X7Y9_W2BEG[0] ;
 wire \Tile_X7Y9_W2BEG[1] ;
 wire \Tile_X7Y9_W2BEG[2] ;
 wire \Tile_X7Y9_W2BEG[3] ;
 wire \Tile_X7Y9_W2BEG[4] ;
 wire \Tile_X7Y9_W2BEG[5] ;
 wire \Tile_X7Y9_W2BEG[6] ;
 wire \Tile_X7Y9_W2BEG[7] ;
 wire \Tile_X7Y9_W2BEGb[0] ;
 wire \Tile_X7Y9_W2BEGb[1] ;
 wire \Tile_X7Y9_W2BEGb[2] ;
 wire \Tile_X7Y9_W2BEGb[3] ;
 wire \Tile_X7Y9_W2BEGb[4] ;
 wire \Tile_X7Y9_W2BEGb[5] ;
 wire \Tile_X7Y9_W2BEGb[6] ;
 wire \Tile_X7Y9_W2BEGb[7] ;
 wire \Tile_X7Y9_W6BEG[0] ;
 wire \Tile_X7Y9_W6BEG[10] ;
 wire \Tile_X7Y9_W6BEG[11] ;
 wire \Tile_X7Y9_W6BEG[1] ;
 wire \Tile_X7Y9_W6BEG[2] ;
 wire \Tile_X7Y9_W6BEG[3] ;
 wire \Tile_X7Y9_W6BEG[4] ;
 wire \Tile_X7Y9_W6BEG[5] ;
 wire \Tile_X7Y9_W6BEG[6] ;
 wire \Tile_X7Y9_W6BEG[7] ;
 wire \Tile_X7Y9_W6BEG[8] ;
 wire \Tile_X7Y9_W6BEG[9] ;
 wire \Tile_X7Y9_WW4BEG[0] ;
 wire \Tile_X7Y9_WW4BEG[10] ;
 wire \Tile_X7Y9_WW4BEG[11] ;
 wire \Tile_X7Y9_WW4BEG[12] ;
 wire \Tile_X7Y9_WW4BEG[13] ;
 wire \Tile_X7Y9_WW4BEG[14] ;
 wire \Tile_X7Y9_WW4BEG[15] ;
 wire \Tile_X7Y9_WW4BEG[1] ;
 wire \Tile_X7Y9_WW4BEG[2] ;
 wire \Tile_X7Y9_WW4BEG[3] ;
 wire \Tile_X7Y9_WW4BEG[4] ;
 wire \Tile_X7Y9_WW4BEG[5] ;
 wire \Tile_X7Y9_WW4BEG[6] ;
 wire \Tile_X7Y9_WW4BEG[7] ;
 wire \Tile_X7Y9_WW4BEG[8] ;
 wire \Tile_X7Y9_WW4BEG[9] ;
 wire \Tile_X8Y0_FrameData_O[0] ;
 wire \Tile_X8Y0_FrameData_O[10] ;
 wire \Tile_X8Y0_FrameData_O[11] ;
 wire \Tile_X8Y0_FrameData_O[12] ;
 wire \Tile_X8Y0_FrameData_O[13] ;
 wire \Tile_X8Y0_FrameData_O[14] ;
 wire \Tile_X8Y0_FrameData_O[15] ;
 wire \Tile_X8Y0_FrameData_O[16] ;
 wire \Tile_X8Y0_FrameData_O[17] ;
 wire \Tile_X8Y0_FrameData_O[18] ;
 wire \Tile_X8Y0_FrameData_O[19] ;
 wire \Tile_X8Y0_FrameData_O[1] ;
 wire \Tile_X8Y0_FrameData_O[20] ;
 wire \Tile_X8Y0_FrameData_O[21] ;
 wire \Tile_X8Y0_FrameData_O[22] ;
 wire \Tile_X8Y0_FrameData_O[23] ;
 wire \Tile_X8Y0_FrameData_O[24] ;
 wire \Tile_X8Y0_FrameData_O[25] ;
 wire \Tile_X8Y0_FrameData_O[26] ;
 wire \Tile_X8Y0_FrameData_O[27] ;
 wire \Tile_X8Y0_FrameData_O[28] ;
 wire \Tile_X8Y0_FrameData_O[29] ;
 wire \Tile_X8Y0_FrameData_O[2] ;
 wire \Tile_X8Y0_FrameData_O[30] ;
 wire \Tile_X8Y0_FrameData_O[31] ;
 wire \Tile_X8Y0_FrameData_O[3] ;
 wire \Tile_X8Y0_FrameData_O[4] ;
 wire \Tile_X8Y0_FrameData_O[5] ;
 wire \Tile_X8Y0_FrameData_O[6] ;
 wire \Tile_X8Y0_FrameData_O[7] ;
 wire \Tile_X8Y0_FrameData_O[8] ;
 wire \Tile_X8Y0_FrameData_O[9] ;
 wire \Tile_X8Y0_FrameStrobe_O[0] ;
 wire \Tile_X8Y0_FrameStrobe_O[10] ;
 wire \Tile_X8Y0_FrameStrobe_O[11] ;
 wire \Tile_X8Y0_FrameStrobe_O[12] ;
 wire \Tile_X8Y0_FrameStrobe_O[13] ;
 wire \Tile_X8Y0_FrameStrobe_O[14] ;
 wire \Tile_X8Y0_FrameStrobe_O[15] ;
 wire \Tile_X8Y0_FrameStrobe_O[16] ;
 wire \Tile_X8Y0_FrameStrobe_O[17] ;
 wire \Tile_X8Y0_FrameStrobe_O[18] ;
 wire \Tile_X8Y0_FrameStrobe_O[19] ;
 wire \Tile_X8Y0_FrameStrobe_O[1] ;
 wire \Tile_X8Y0_FrameStrobe_O[2] ;
 wire \Tile_X8Y0_FrameStrobe_O[3] ;
 wire \Tile_X8Y0_FrameStrobe_O[4] ;
 wire \Tile_X8Y0_FrameStrobe_O[5] ;
 wire \Tile_X8Y0_FrameStrobe_O[6] ;
 wire \Tile_X8Y0_FrameStrobe_O[7] ;
 wire \Tile_X8Y0_FrameStrobe_O[8] ;
 wire \Tile_X8Y0_FrameStrobe_O[9] ;
 wire \Tile_X8Y0_S1BEG[0] ;
 wire \Tile_X8Y0_S1BEG[1] ;
 wire \Tile_X8Y0_S1BEG[2] ;
 wire \Tile_X8Y0_S1BEG[3] ;
 wire \Tile_X8Y0_S2BEG[0] ;
 wire \Tile_X8Y0_S2BEG[1] ;
 wire \Tile_X8Y0_S2BEG[2] ;
 wire \Tile_X8Y0_S2BEG[3] ;
 wire \Tile_X8Y0_S2BEG[4] ;
 wire \Tile_X8Y0_S2BEG[5] ;
 wire \Tile_X8Y0_S2BEG[6] ;
 wire \Tile_X8Y0_S2BEG[7] ;
 wire \Tile_X8Y0_S2BEGb[0] ;
 wire \Tile_X8Y0_S2BEGb[1] ;
 wire \Tile_X8Y0_S2BEGb[2] ;
 wire \Tile_X8Y0_S2BEGb[3] ;
 wire \Tile_X8Y0_S2BEGb[4] ;
 wire \Tile_X8Y0_S2BEGb[5] ;
 wire \Tile_X8Y0_S2BEGb[6] ;
 wire \Tile_X8Y0_S2BEGb[7] ;
 wire \Tile_X8Y0_S4BEG[0] ;
 wire \Tile_X8Y0_S4BEG[10] ;
 wire \Tile_X8Y0_S4BEG[11] ;
 wire \Tile_X8Y0_S4BEG[12] ;
 wire \Tile_X8Y0_S4BEG[13] ;
 wire \Tile_X8Y0_S4BEG[14] ;
 wire \Tile_X8Y0_S4BEG[15] ;
 wire \Tile_X8Y0_S4BEG[1] ;
 wire \Tile_X8Y0_S4BEG[2] ;
 wire \Tile_X8Y0_S4BEG[3] ;
 wire \Tile_X8Y0_S4BEG[4] ;
 wire \Tile_X8Y0_S4BEG[5] ;
 wire \Tile_X8Y0_S4BEG[6] ;
 wire \Tile_X8Y0_S4BEG[7] ;
 wire \Tile_X8Y0_S4BEG[8] ;
 wire \Tile_X8Y0_S4BEG[9] ;
 wire \Tile_X8Y0_SS4BEG[0] ;
 wire \Tile_X8Y0_SS4BEG[10] ;
 wire \Tile_X8Y0_SS4BEG[11] ;
 wire \Tile_X8Y0_SS4BEG[12] ;
 wire \Tile_X8Y0_SS4BEG[13] ;
 wire \Tile_X8Y0_SS4BEG[14] ;
 wire \Tile_X8Y0_SS4BEG[15] ;
 wire \Tile_X8Y0_SS4BEG[1] ;
 wire \Tile_X8Y0_SS4BEG[2] ;
 wire \Tile_X8Y0_SS4BEG[3] ;
 wire \Tile_X8Y0_SS4BEG[4] ;
 wire \Tile_X8Y0_SS4BEG[5] ;
 wire \Tile_X8Y0_SS4BEG[6] ;
 wire \Tile_X8Y0_SS4BEG[7] ;
 wire \Tile_X8Y0_SS4BEG[8] ;
 wire \Tile_X8Y0_SS4BEG[9] ;
 wire Tile_X8Y0_UserCLKo;
 wire Tile_X8Y10_Co;
 wire \Tile_X8Y10_E1BEG[0] ;
 wire \Tile_X8Y10_E1BEG[1] ;
 wire \Tile_X8Y10_E1BEG[2] ;
 wire \Tile_X8Y10_E1BEG[3] ;
 wire \Tile_X8Y10_E2BEG[0] ;
 wire \Tile_X8Y10_E2BEG[1] ;
 wire \Tile_X8Y10_E2BEG[2] ;
 wire \Tile_X8Y10_E2BEG[3] ;
 wire \Tile_X8Y10_E2BEG[4] ;
 wire \Tile_X8Y10_E2BEG[5] ;
 wire \Tile_X8Y10_E2BEG[6] ;
 wire \Tile_X8Y10_E2BEG[7] ;
 wire \Tile_X8Y10_E2BEGb[0] ;
 wire \Tile_X8Y10_E2BEGb[1] ;
 wire \Tile_X8Y10_E2BEGb[2] ;
 wire \Tile_X8Y10_E2BEGb[3] ;
 wire \Tile_X8Y10_E2BEGb[4] ;
 wire \Tile_X8Y10_E2BEGb[5] ;
 wire \Tile_X8Y10_E2BEGb[6] ;
 wire \Tile_X8Y10_E2BEGb[7] ;
 wire \Tile_X8Y10_E6BEG[0] ;
 wire \Tile_X8Y10_E6BEG[10] ;
 wire \Tile_X8Y10_E6BEG[11] ;
 wire \Tile_X8Y10_E6BEG[1] ;
 wire \Tile_X8Y10_E6BEG[2] ;
 wire \Tile_X8Y10_E6BEG[3] ;
 wire \Tile_X8Y10_E6BEG[4] ;
 wire \Tile_X8Y10_E6BEG[5] ;
 wire \Tile_X8Y10_E6BEG[6] ;
 wire \Tile_X8Y10_E6BEG[7] ;
 wire \Tile_X8Y10_E6BEG[8] ;
 wire \Tile_X8Y10_E6BEG[9] ;
 wire \Tile_X8Y10_EE4BEG[0] ;
 wire \Tile_X8Y10_EE4BEG[10] ;
 wire \Tile_X8Y10_EE4BEG[11] ;
 wire \Tile_X8Y10_EE4BEG[12] ;
 wire \Tile_X8Y10_EE4BEG[13] ;
 wire \Tile_X8Y10_EE4BEG[14] ;
 wire \Tile_X8Y10_EE4BEG[15] ;
 wire \Tile_X8Y10_EE4BEG[1] ;
 wire \Tile_X8Y10_EE4BEG[2] ;
 wire \Tile_X8Y10_EE4BEG[3] ;
 wire \Tile_X8Y10_EE4BEG[4] ;
 wire \Tile_X8Y10_EE4BEG[5] ;
 wire \Tile_X8Y10_EE4BEG[6] ;
 wire \Tile_X8Y10_EE4BEG[7] ;
 wire \Tile_X8Y10_EE4BEG[8] ;
 wire \Tile_X8Y10_EE4BEG[9] ;
 wire \Tile_X8Y10_FrameData_O[0] ;
 wire \Tile_X8Y10_FrameData_O[10] ;
 wire \Tile_X8Y10_FrameData_O[11] ;
 wire \Tile_X8Y10_FrameData_O[12] ;
 wire \Tile_X8Y10_FrameData_O[13] ;
 wire \Tile_X8Y10_FrameData_O[14] ;
 wire \Tile_X8Y10_FrameData_O[15] ;
 wire \Tile_X8Y10_FrameData_O[16] ;
 wire \Tile_X8Y10_FrameData_O[17] ;
 wire \Tile_X8Y10_FrameData_O[18] ;
 wire \Tile_X8Y10_FrameData_O[19] ;
 wire \Tile_X8Y10_FrameData_O[1] ;
 wire \Tile_X8Y10_FrameData_O[20] ;
 wire \Tile_X8Y10_FrameData_O[21] ;
 wire \Tile_X8Y10_FrameData_O[22] ;
 wire \Tile_X8Y10_FrameData_O[23] ;
 wire \Tile_X8Y10_FrameData_O[24] ;
 wire \Tile_X8Y10_FrameData_O[25] ;
 wire \Tile_X8Y10_FrameData_O[26] ;
 wire \Tile_X8Y10_FrameData_O[27] ;
 wire \Tile_X8Y10_FrameData_O[28] ;
 wire \Tile_X8Y10_FrameData_O[29] ;
 wire \Tile_X8Y10_FrameData_O[2] ;
 wire \Tile_X8Y10_FrameData_O[30] ;
 wire \Tile_X8Y10_FrameData_O[31] ;
 wire \Tile_X8Y10_FrameData_O[3] ;
 wire \Tile_X8Y10_FrameData_O[4] ;
 wire \Tile_X8Y10_FrameData_O[5] ;
 wire \Tile_X8Y10_FrameData_O[6] ;
 wire \Tile_X8Y10_FrameData_O[7] ;
 wire \Tile_X8Y10_FrameData_O[8] ;
 wire \Tile_X8Y10_FrameData_O[9] ;
 wire \Tile_X8Y10_FrameStrobe_O[0] ;
 wire \Tile_X8Y10_FrameStrobe_O[10] ;
 wire \Tile_X8Y10_FrameStrobe_O[11] ;
 wire \Tile_X8Y10_FrameStrobe_O[12] ;
 wire \Tile_X8Y10_FrameStrobe_O[13] ;
 wire \Tile_X8Y10_FrameStrobe_O[14] ;
 wire \Tile_X8Y10_FrameStrobe_O[15] ;
 wire \Tile_X8Y10_FrameStrobe_O[16] ;
 wire \Tile_X8Y10_FrameStrobe_O[17] ;
 wire \Tile_X8Y10_FrameStrobe_O[18] ;
 wire \Tile_X8Y10_FrameStrobe_O[19] ;
 wire \Tile_X8Y10_FrameStrobe_O[1] ;
 wire \Tile_X8Y10_FrameStrobe_O[2] ;
 wire \Tile_X8Y10_FrameStrobe_O[3] ;
 wire \Tile_X8Y10_FrameStrobe_O[4] ;
 wire \Tile_X8Y10_FrameStrobe_O[5] ;
 wire \Tile_X8Y10_FrameStrobe_O[6] ;
 wire \Tile_X8Y10_FrameStrobe_O[7] ;
 wire \Tile_X8Y10_FrameStrobe_O[8] ;
 wire \Tile_X8Y10_FrameStrobe_O[9] ;
 wire \Tile_X8Y10_N1BEG[0] ;
 wire \Tile_X8Y10_N1BEG[1] ;
 wire \Tile_X8Y10_N1BEG[2] ;
 wire \Tile_X8Y10_N1BEG[3] ;
 wire \Tile_X8Y10_N2BEG[0] ;
 wire \Tile_X8Y10_N2BEG[1] ;
 wire \Tile_X8Y10_N2BEG[2] ;
 wire \Tile_X8Y10_N2BEG[3] ;
 wire \Tile_X8Y10_N2BEG[4] ;
 wire \Tile_X8Y10_N2BEG[5] ;
 wire \Tile_X8Y10_N2BEG[6] ;
 wire \Tile_X8Y10_N2BEG[7] ;
 wire \Tile_X8Y10_N2BEGb[0] ;
 wire \Tile_X8Y10_N2BEGb[1] ;
 wire \Tile_X8Y10_N2BEGb[2] ;
 wire \Tile_X8Y10_N2BEGb[3] ;
 wire \Tile_X8Y10_N2BEGb[4] ;
 wire \Tile_X8Y10_N2BEGb[5] ;
 wire \Tile_X8Y10_N2BEGb[6] ;
 wire \Tile_X8Y10_N2BEGb[7] ;
 wire \Tile_X8Y10_N4BEG[0] ;
 wire \Tile_X8Y10_N4BEG[10] ;
 wire \Tile_X8Y10_N4BEG[11] ;
 wire \Tile_X8Y10_N4BEG[12] ;
 wire \Tile_X8Y10_N4BEG[13] ;
 wire \Tile_X8Y10_N4BEG[14] ;
 wire \Tile_X8Y10_N4BEG[15] ;
 wire \Tile_X8Y10_N4BEG[1] ;
 wire \Tile_X8Y10_N4BEG[2] ;
 wire \Tile_X8Y10_N4BEG[3] ;
 wire \Tile_X8Y10_N4BEG[4] ;
 wire \Tile_X8Y10_N4BEG[5] ;
 wire \Tile_X8Y10_N4BEG[6] ;
 wire \Tile_X8Y10_N4BEG[7] ;
 wire \Tile_X8Y10_N4BEG[8] ;
 wire \Tile_X8Y10_N4BEG[9] ;
 wire \Tile_X8Y10_NN4BEG[0] ;
 wire \Tile_X8Y10_NN4BEG[10] ;
 wire \Tile_X8Y10_NN4BEG[11] ;
 wire \Tile_X8Y10_NN4BEG[12] ;
 wire \Tile_X8Y10_NN4BEG[13] ;
 wire \Tile_X8Y10_NN4BEG[14] ;
 wire \Tile_X8Y10_NN4BEG[15] ;
 wire \Tile_X8Y10_NN4BEG[1] ;
 wire \Tile_X8Y10_NN4BEG[2] ;
 wire \Tile_X8Y10_NN4BEG[3] ;
 wire \Tile_X8Y10_NN4BEG[4] ;
 wire \Tile_X8Y10_NN4BEG[5] ;
 wire \Tile_X8Y10_NN4BEG[6] ;
 wire \Tile_X8Y10_NN4BEG[7] ;
 wire \Tile_X8Y10_NN4BEG[8] ;
 wire \Tile_X8Y10_NN4BEG[9] ;
 wire \Tile_X8Y10_S1BEG[0] ;
 wire \Tile_X8Y10_S1BEG[1] ;
 wire \Tile_X8Y10_S1BEG[2] ;
 wire \Tile_X8Y10_S1BEG[3] ;
 wire \Tile_X8Y10_S2BEG[0] ;
 wire \Tile_X8Y10_S2BEG[1] ;
 wire \Tile_X8Y10_S2BEG[2] ;
 wire \Tile_X8Y10_S2BEG[3] ;
 wire \Tile_X8Y10_S2BEG[4] ;
 wire \Tile_X8Y10_S2BEG[5] ;
 wire \Tile_X8Y10_S2BEG[6] ;
 wire \Tile_X8Y10_S2BEG[7] ;
 wire \Tile_X8Y10_S2BEGb[0] ;
 wire \Tile_X8Y10_S2BEGb[1] ;
 wire \Tile_X8Y10_S2BEGb[2] ;
 wire \Tile_X8Y10_S2BEGb[3] ;
 wire \Tile_X8Y10_S2BEGb[4] ;
 wire \Tile_X8Y10_S2BEGb[5] ;
 wire \Tile_X8Y10_S2BEGb[6] ;
 wire \Tile_X8Y10_S2BEGb[7] ;
 wire \Tile_X8Y10_S4BEG[0] ;
 wire \Tile_X8Y10_S4BEG[10] ;
 wire \Tile_X8Y10_S4BEG[11] ;
 wire \Tile_X8Y10_S4BEG[12] ;
 wire \Tile_X8Y10_S4BEG[13] ;
 wire \Tile_X8Y10_S4BEG[14] ;
 wire \Tile_X8Y10_S4BEG[15] ;
 wire \Tile_X8Y10_S4BEG[1] ;
 wire \Tile_X8Y10_S4BEG[2] ;
 wire \Tile_X8Y10_S4BEG[3] ;
 wire \Tile_X8Y10_S4BEG[4] ;
 wire \Tile_X8Y10_S4BEG[5] ;
 wire \Tile_X8Y10_S4BEG[6] ;
 wire \Tile_X8Y10_S4BEG[7] ;
 wire \Tile_X8Y10_S4BEG[8] ;
 wire \Tile_X8Y10_S4BEG[9] ;
 wire \Tile_X8Y10_SS4BEG[0] ;
 wire \Tile_X8Y10_SS4BEG[10] ;
 wire \Tile_X8Y10_SS4BEG[11] ;
 wire \Tile_X8Y10_SS4BEG[12] ;
 wire \Tile_X8Y10_SS4BEG[13] ;
 wire \Tile_X8Y10_SS4BEG[14] ;
 wire \Tile_X8Y10_SS4BEG[15] ;
 wire \Tile_X8Y10_SS4BEG[1] ;
 wire \Tile_X8Y10_SS4BEG[2] ;
 wire \Tile_X8Y10_SS4BEG[3] ;
 wire \Tile_X8Y10_SS4BEG[4] ;
 wire \Tile_X8Y10_SS4BEG[5] ;
 wire \Tile_X8Y10_SS4BEG[6] ;
 wire \Tile_X8Y10_SS4BEG[7] ;
 wire \Tile_X8Y10_SS4BEG[8] ;
 wire \Tile_X8Y10_SS4BEG[9] ;
 wire Tile_X8Y10_UserCLKo;
 wire \Tile_X8Y10_W1BEG[0] ;
 wire \Tile_X8Y10_W1BEG[1] ;
 wire \Tile_X8Y10_W1BEG[2] ;
 wire \Tile_X8Y10_W1BEG[3] ;
 wire \Tile_X8Y10_W2BEG[0] ;
 wire \Tile_X8Y10_W2BEG[1] ;
 wire \Tile_X8Y10_W2BEG[2] ;
 wire \Tile_X8Y10_W2BEG[3] ;
 wire \Tile_X8Y10_W2BEG[4] ;
 wire \Tile_X8Y10_W2BEG[5] ;
 wire \Tile_X8Y10_W2BEG[6] ;
 wire \Tile_X8Y10_W2BEG[7] ;
 wire \Tile_X8Y10_W2BEGb[0] ;
 wire \Tile_X8Y10_W2BEGb[1] ;
 wire \Tile_X8Y10_W2BEGb[2] ;
 wire \Tile_X8Y10_W2BEGb[3] ;
 wire \Tile_X8Y10_W2BEGb[4] ;
 wire \Tile_X8Y10_W2BEGb[5] ;
 wire \Tile_X8Y10_W2BEGb[6] ;
 wire \Tile_X8Y10_W2BEGb[7] ;
 wire \Tile_X8Y10_W6BEG[0] ;
 wire \Tile_X8Y10_W6BEG[10] ;
 wire \Tile_X8Y10_W6BEG[11] ;
 wire \Tile_X8Y10_W6BEG[1] ;
 wire \Tile_X8Y10_W6BEG[2] ;
 wire \Tile_X8Y10_W6BEG[3] ;
 wire \Tile_X8Y10_W6BEG[4] ;
 wire \Tile_X8Y10_W6BEG[5] ;
 wire \Tile_X8Y10_W6BEG[6] ;
 wire \Tile_X8Y10_W6BEG[7] ;
 wire \Tile_X8Y10_W6BEG[8] ;
 wire \Tile_X8Y10_W6BEG[9] ;
 wire \Tile_X8Y10_WW4BEG[0] ;
 wire \Tile_X8Y10_WW4BEG[10] ;
 wire \Tile_X8Y10_WW4BEG[11] ;
 wire \Tile_X8Y10_WW4BEG[12] ;
 wire \Tile_X8Y10_WW4BEG[13] ;
 wire \Tile_X8Y10_WW4BEG[14] ;
 wire \Tile_X8Y10_WW4BEG[15] ;
 wire \Tile_X8Y10_WW4BEG[1] ;
 wire \Tile_X8Y10_WW4BEG[2] ;
 wire \Tile_X8Y10_WW4BEG[3] ;
 wire \Tile_X8Y10_WW4BEG[4] ;
 wire \Tile_X8Y10_WW4BEG[5] ;
 wire \Tile_X8Y10_WW4BEG[6] ;
 wire \Tile_X8Y10_WW4BEG[7] ;
 wire \Tile_X8Y10_WW4BEG[8] ;
 wire \Tile_X8Y10_WW4BEG[9] ;
 wire Tile_X8Y11_Co;
 wire \Tile_X8Y11_E1BEG[0] ;
 wire \Tile_X8Y11_E1BEG[1] ;
 wire \Tile_X8Y11_E1BEG[2] ;
 wire \Tile_X8Y11_E1BEG[3] ;
 wire \Tile_X8Y11_E2BEG[0] ;
 wire \Tile_X8Y11_E2BEG[1] ;
 wire \Tile_X8Y11_E2BEG[2] ;
 wire \Tile_X8Y11_E2BEG[3] ;
 wire \Tile_X8Y11_E2BEG[4] ;
 wire \Tile_X8Y11_E2BEG[5] ;
 wire \Tile_X8Y11_E2BEG[6] ;
 wire \Tile_X8Y11_E2BEG[7] ;
 wire \Tile_X8Y11_E2BEGb[0] ;
 wire \Tile_X8Y11_E2BEGb[1] ;
 wire \Tile_X8Y11_E2BEGb[2] ;
 wire \Tile_X8Y11_E2BEGb[3] ;
 wire \Tile_X8Y11_E2BEGb[4] ;
 wire \Tile_X8Y11_E2BEGb[5] ;
 wire \Tile_X8Y11_E2BEGb[6] ;
 wire \Tile_X8Y11_E2BEGb[7] ;
 wire \Tile_X8Y11_E6BEG[0] ;
 wire \Tile_X8Y11_E6BEG[10] ;
 wire \Tile_X8Y11_E6BEG[11] ;
 wire \Tile_X8Y11_E6BEG[1] ;
 wire \Tile_X8Y11_E6BEG[2] ;
 wire \Tile_X8Y11_E6BEG[3] ;
 wire \Tile_X8Y11_E6BEG[4] ;
 wire \Tile_X8Y11_E6BEG[5] ;
 wire \Tile_X8Y11_E6BEG[6] ;
 wire \Tile_X8Y11_E6BEG[7] ;
 wire \Tile_X8Y11_E6BEG[8] ;
 wire \Tile_X8Y11_E6BEG[9] ;
 wire \Tile_X8Y11_EE4BEG[0] ;
 wire \Tile_X8Y11_EE4BEG[10] ;
 wire \Tile_X8Y11_EE4BEG[11] ;
 wire \Tile_X8Y11_EE4BEG[12] ;
 wire \Tile_X8Y11_EE4BEG[13] ;
 wire \Tile_X8Y11_EE4BEG[14] ;
 wire \Tile_X8Y11_EE4BEG[15] ;
 wire \Tile_X8Y11_EE4BEG[1] ;
 wire \Tile_X8Y11_EE4BEG[2] ;
 wire \Tile_X8Y11_EE4BEG[3] ;
 wire \Tile_X8Y11_EE4BEG[4] ;
 wire \Tile_X8Y11_EE4BEG[5] ;
 wire \Tile_X8Y11_EE4BEG[6] ;
 wire \Tile_X8Y11_EE4BEG[7] ;
 wire \Tile_X8Y11_EE4BEG[8] ;
 wire \Tile_X8Y11_EE4BEG[9] ;
 wire \Tile_X8Y11_FrameData_O[0] ;
 wire \Tile_X8Y11_FrameData_O[10] ;
 wire \Tile_X8Y11_FrameData_O[11] ;
 wire \Tile_X8Y11_FrameData_O[12] ;
 wire \Tile_X8Y11_FrameData_O[13] ;
 wire \Tile_X8Y11_FrameData_O[14] ;
 wire \Tile_X8Y11_FrameData_O[15] ;
 wire \Tile_X8Y11_FrameData_O[16] ;
 wire \Tile_X8Y11_FrameData_O[17] ;
 wire \Tile_X8Y11_FrameData_O[18] ;
 wire \Tile_X8Y11_FrameData_O[19] ;
 wire \Tile_X8Y11_FrameData_O[1] ;
 wire \Tile_X8Y11_FrameData_O[20] ;
 wire \Tile_X8Y11_FrameData_O[21] ;
 wire \Tile_X8Y11_FrameData_O[22] ;
 wire \Tile_X8Y11_FrameData_O[23] ;
 wire \Tile_X8Y11_FrameData_O[24] ;
 wire \Tile_X8Y11_FrameData_O[25] ;
 wire \Tile_X8Y11_FrameData_O[26] ;
 wire \Tile_X8Y11_FrameData_O[27] ;
 wire \Tile_X8Y11_FrameData_O[28] ;
 wire \Tile_X8Y11_FrameData_O[29] ;
 wire \Tile_X8Y11_FrameData_O[2] ;
 wire \Tile_X8Y11_FrameData_O[30] ;
 wire \Tile_X8Y11_FrameData_O[31] ;
 wire \Tile_X8Y11_FrameData_O[3] ;
 wire \Tile_X8Y11_FrameData_O[4] ;
 wire \Tile_X8Y11_FrameData_O[5] ;
 wire \Tile_X8Y11_FrameData_O[6] ;
 wire \Tile_X8Y11_FrameData_O[7] ;
 wire \Tile_X8Y11_FrameData_O[8] ;
 wire \Tile_X8Y11_FrameData_O[9] ;
 wire \Tile_X8Y11_FrameStrobe_O[0] ;
 wire \Tile_X8Y11_FrameStrobe_O[10] ;
 wire \Tile_X8Y11_FrameStrobe_O[11] ;
 wire \Tile_X8Y11_FrameStrobe_O[12] ;
 wire \Tile_X8Y11_FrameStrobe_O[13] ;
 wire \Tile_X8Y11_FrameStrobe_O[14] ;
 wire \Tile_X8Y11_FrameStrobe_O[15] ;
 wire \Tile_X8Y11_FrameStrobe_O[16] ;
 wire \Tile_X8Y11_FrameStrobe_O[17] ;
 wire \Tile_X8Y11_FrameStrobe_O[18] ;
 wire \Tile_X8Y11_FrameStrobe_O[19] ;
 wire \Tile_X8Y11_FrameStrobe_O[1] ;
 wire \Tile_X8Y11_FrameStrobe_O[2] ;
 wire \Tile_X8Y11_FrameStrobe_O[3] ;
 wire \Tile_X8Y11_FrameStrobe_O[4] ;
 wire \Tile_X8Y11_FrameStrobe_O[5] ;
 wire \Tile_X8Y11_FrameStrobe_O[6] ;
 wire \Tile_X8Y11_FrameStrobe_O[7] ;
 wire \Tile_X8Y11_FrameStrobe_O[8] ;
 wire \Tile_X8Y11_FrameStrobe_O[9] ;
 wire \Tile_X8Y11_N1BEG[0] ;
 wire \Tile_X8Y11_N1BEG[1] ;
 wire \Tile_X8Y11_N1BEG[2] ;
 wire \Tile_X8Y11_N1BEG[3] ;
 wire \Tile_X8Y11_N2BEG[0] ;
 wire \Tile_X8Y11_N2BEG[1] ;
 wire \Tile_X8Y11_N2BEG[2] ;
 wire \Tile_X8Y11_N2BEG[3] ;
 wire \Tile_X8Y11_N2BEG[4] ;
 wire \Tile_X8Y11_N2BEG[5] ;
 wire \Tile_X8Y11_N2BEG[6] ;
 wire \Tile_X8Y11_N2BEG[7] ;
 wire \Tile_X8Y11_N2BEGb[0] ;
 wire \Tile_X8Y11_N2BEGb[1] ;
 wire \Tile_X8Y11_N2BEGb[2] ;
 wire \Tile_X8Y11_N2BEGb[3] ;
 wire \Tile_X8Y11_N2BEGb[4] ;
 wire \Tile_X8Y11_N2BEGb[5] ;
 wire \Tile_X8Y11_N2BEGb[6] ;
 wire \Tile_X8Y11_N2BEGb[7] ;
 wire \Tile_X8Y11_N4BEG[0] ;
 wire \Tile_X8Y11_N4BEG[10] ;
 wire \Tile_X8Y11_N4BEG[11] ;
 wire \Tile_X8Y11_N4BEG[12] ;
 wire \Tile_X8Y11_N4BEG[13] ;
 wire \Tile_X8Y11_N4BEG[14] ;
 wire \Tile_X8Y11_N4BEG[15] ;
 wire \Tile_X8Y11_N4BEG[1] ;
 wire \Tile_X8Y11_N4BEG[2] ;
 wire \Tile_X8Y11_N4BEG[3] ;
 wire \Tile_X8Y11_N4BEG[4] ;
 wire \Tile_X8Y11_N4BEG[5] ;
 wire \Tile_X8Y11_N4BEG[6] ;
 wire \Tile_X8Y11_N4BEG[7] ;
 wire \Tile_X8Y11_N4BEG[8] ;
 wire \Tile_X8Y11_N4BEG[9] ;
 wire \Tile_X8Y11_NN4BEG[0] ;
 wire \Tile_X8Y11_NN4BEG[10] ;
 wire \Tile_X8Y11_NN4BEG[11] ;
 wire \Tile_X8Y11_NN4BEG[12] ;
 wire \Tile_X8Y11_NN4BEG[13] ;
 wire \Tile_X8Y11_NN4BEG[14] ;
 wire \Tile_X8Y11_NN4BEG[15] ;
 wire \Tile_X8Y11_NN4BEG[1] ;
 wire \Tile_X8Y11_NN4BEG[2] ;
 wire \Tile_X8Y11_NN4BEG[3] ;
 wire \Tile_X8Y11_NN4BEG[4] ;
 wire \Tile_X8Y11_NN4BEG[5] ;
 wire \Tile_X8Y11_NN4BEG[6] ;
 wire \Tile_X8Y11_NN4BEG[7] ;
 wire \Tile_X8Y11_NN4BEG[8] ;
 wire \Tile_X8Y11_NN4BEG[9] ;
 wire \Tile_X8Y11_S1BEG[0] ;
 wire \Tile_X8Y11_S1BEG[1] ;
 wire \Tile_X8Y11_S1BEG[2] ;
 wire \Tile_X8Y11_S1BEG[3] ;
 wire \Tile_X8Y11_S2BEG[0] ;
 wire \Tile_X8Y11_S2BEG[1] ;
 wire \Tile_X8Y11_S2BEG[2] ;
 wire \Tile_X8Y11_S2BEG[3] ;
 wire \Tile_X8Y11_S2BEG[4] ;
 wire \Tile_X8Y11_S2BEG[5] ;
 wire \Tile_X8Y11_S2BEG[6] ;
 wire \Tile_X8Y11_S2BEG[7] ;
 wire \Tile_X8Y11_S2BEGb[0] ;
 wire \Tile_X8Y11_S2BEGb[1] ;
 wire \Tile_X8Y11_S2BEGb[2] ;
 wire \Tile_X8Y11_S2BEGb[3] ;
 wire \Tile_X8Y11_S2BEGb[4] ;
 wire \Tile_X8Y11_S2BEGb[5] ;
 wire \Tile_X8Y11_S2BEGb[6] ;
 wire \Tile_X8Y11_S2BEGb[7] ;
 wire \Tile_X8Y11_S4BEG[0] ;
 wire \Tile_X8Y11_S4BEG[10] ;
 wire \Tile_X8Y11_S4BEG[11] ;
 wire \Tile_X8Y11_S4BEG[12] ;
 wire \Tile_X8Y11_S4BEG[13] ;
 wire \Tile_X8Y11_S4BEG[14] ;
 wire \Tile_X8Y11_S4BEG[15] ;
 wire \Tile_X8Y11_S4BEG[1] ;
 wire \Tile_X8Y11_S4BEG[2] ;
 wire \Tile_X8Y11_S4BEG[3] ;
 wire \Tile_X8Y11_S4BEG[4] ;
 wire \Tile_X8Y11_S4BEG[5] ;
 wire \Tile_X8Y11_S4BEG[6] ;
 wire \Tile_X8Y11_S4BEG[7] ;
 wire \Tile_X8Y11_S4BEG[8] ;
 wire \Tile_X8Y11_S4BEG[9] ;
 wire \Tile_X8Y11_SS4BEG[0] ;
 wire \Tile_X8Y11_SS4BEG[10] ;
 wire \Tile_X8Y11_SS4BEG[11] ;
 wire \Tile_X8Y11_SS4BEG[12] ;
 wire \Tile_X8Y11_SS4BEG[13] ;
 wire \Tile_X8Y11_SS4BEG[14] ;
 wire \Tile_X8Y11_SS4BEG[15] ;
 wire \Tile_X8Y11_SS4BEG[1] ;
 wire \Tile_X8Y11_SS4BEG[2] ;
 wire \Tile_X8Y11_SS4BEG[3] ;
 wire \Tile_X8Y11_SS4BEG[4] ;
 wire \Tile_X8Y11_SS4BEG[5] ;
 wire \Tile_X8Y11_SS4BEG[6] ;
 wire \Tile_X8Y11_SS4BEG[7] ;
 wire \Tile_X8Y11_SS4BEG[8] ;
 wire \Tile_X8Y11_SS4BEG[9] ;
 wire Tile_X8Y11_UserCLKo;
 wire \Tile_X8Y11_W1BEG[0] ;
 wire \Tile_X8Y11_W1BEG[1] ;
 wire \Tile_X8Y11_W1BEG[2] ;
 wire \Tile_X8Y11_W1BEG[3] ;
 wire \Tile_X8Y11_W2BEG[0] ;
 wire \Tile_X8Y11_W2BEG[1] ;
 wire \Tile_X8Y11_W2BEG[2] ;
 wire \Tile_X8Y11_W2BEG[3] ;
 wire \Tile_X8Y11_W2BEG[4] ;
 wire \Tile_X8Y11_W2BEG[5] ;
 wire \Tile_X8Y11_W2BEG[6] ;
 wire \Tile_X8Y11_W2BEG[7] ;
 wire \Tile_X8Y11_W2BEGb[0] ;
 wire \Tile_X8Y11_W2BEGb[1] ;
 wire \Tile_X8Y11_W2BEGb[2] ;
 wire \Tile_X8Y11_W2BEGb[3] ;
 wire \Tile_X8Y11_W2BEGb[4] ;
 wire \Tile_X8Y11_W2BEGb[5] ;
 wire \Tile_X8Y11_W2BEGb[6] ;
 wire \Tile_X8Y11_W2BEGb[7] ;
 wire \Tile_X8Y11_W6BEG[0] ;
 wire \Tile_X8Y11_W6BEG[10] ;
 wire \Tile_X8Y11_W6BEG[11] ;
 wire \Tile_X8Y11_W6BEG[1] ;
 wire \Tile_X8Y11_W6BEG[2] ;
 wire \Tile_X8Y11_W6BEG[3] ;
 wire \Tile_X8Y11_W6BEG[4] ;
 wire \Tile_X8Y11_W6BEG[5] ;
 wire \Tile_X8Y11_W6BEG[6] ;
 wire \Tile_X8Y11_W6BEG[7] ;
 wire \Tile_X8Y11_W6BEG[8] ;
 wire \Tile_X8Y11_W6BEG[9] ;
 wire \Tile_X8Y11_WW4BEG[0] ;
 wire \Tile_X8Y11_WW4BEG[10] ;
 wire \Tile_X8Y11_WW4BEG[11] ;
 wire \Tile_X8Y11_WW4BEG[12] ;
 wire \Tile_X8Y11_WW4BEG[13] ;
 wire \Tile_X8Y11_WW4BEG[14] ;
 wire \Tile_X8Y11_WW4BEG[15] ;
 wire \Tile_X8Y11_WW4BEG[1] ;
 wire \Tile_X8Y11_WW4BEG[2] ;
 wire \Tile_X8Y11_WW4BEG[3] ;
 wire \Tile_X8Y11_WW4BEG[4] ;
 wire \Tile_X8Y11_WW4BEG[5] ;
 wire \Tile_X8Y11_WW4BEG[6] ;
 wire \Tile_X8Y11_WW4BEG[7] ;
 wire \Tile_X8Y11_WW4BEG[8] ;
 wire \Tile_X8Y11_WW4BEG[9] ;
 wire Tile_X8Y12_Co;
 wire \Tile_X8Y12_E1BEG[0] ;
 wire \Tile_X8Y12_E1BEG[1] ;
 wire \Tile_X8Y12_E1BEG[2] ;
 wire \Tile_X8Y12_E1BEG[3] ;
 wire \Tile_X8Y12_E2BEG[0] ;
 wire \Tile_X8Y12_E2BEG[1] ;
 wire \Tile_X8Y12_E2BEG[2] ;
 wire \Tile_X8Y12_E2BEG[3] ;
 wire \Tile_X8Y12_E2BEG[4] ;
 wire \Tile_X8Y12_E2BEG[5] ;
 wire \Tile_X8Y12_E2BEG[6] ;
 wire \Tile_X8Y12_E2BEG[7] ;
 wire \Tile_X8Y12_E2BEGb[0] ;
 wire \Tile_X8Y12_E2BEGb[1] ;
 wire \Tile_X8Y12_E2BEGb[2] ;
 wire \Tile_X8Y12_E2BEGb[3] ;
 wire \Tile_X8Y12_E2BEGb[4] ;
 wire \Tile_X8Y12_E2BEGb[5] ;
 wire \Tile_X8Y12_E2BEGb[6] ;
 wire \Tile_X8Y12_E2BEGb[7] ;
 wire \Tile_X8Y12_E6BEG[0] ;
 wire \Tile_X8Y12_E6BEG[10] ;
 wire \Tile_X8Y12_E6BEG[11] ;
 wire \Tile_X8Y12_E6BEG[1] ;
 wire \Tile_X8Y12_E6BEG[2] ;
 wire \Tile_X8Y12_E6BEG[3] ;
 wire \Tile_X8Y12_E6BEG[4] ;
 wire \Tile_X8Y12_E6BEG[5] ;
 wire \Tile_X8Y12_E6BEG[6] ;
 wire \Tile_X8Y12_E6BEG[7] ;
 wire \Tile_X8Y12_E6BEG[8] ;
 wire \Tile_X8Y12_E6BEG[9] ;
 wire \Tile_X8Y12_EE4BEG[0] ;
 wire \Tile_X8Y12_EE4BEG[10] ;
 wire \Tile_X8Y12_EE4BEG[11] ;
 wire \Tile_X8Y12_EE4BEG[12] ;
 wire \Tile_X8Y12_EE4BEG[13] ;
 wire \Tile_X8Y12_EE4BEG[14] ;
 wire \Tile_X8Y12_EE4BEG[15] ;
 wire \Tile_X8Y12_EE4BEG[1] ;
 wire \Tile_X8Y12_EE4BEG[2] ;
 wire \Tile_X8Y12_EE4BEG[3] ;
 wire \Tile_X8Y12_EE4BEG[4] ;
 wire \Tile_X8Y12_EE4BEG[5] ;
 wire \Tile_X8Y12_EE4BEG[6] ;
 wire \Tile_X8Y12_EE4BEG[7] ;
 wire \Tile_X8Y12_EE4BEG[8] ;
 wire \Tile_X8Y12_EE4BEG[9] ;
 wire \Tile_X8Y12_FrameData_O[0] ;
 wire \Tile_X8Y12_FrameData_O[10] ;
 wire \Tile_X8Y12_FrameData_O[11] ;
 wire \Tile_X8Y12_FrameData_O[12] ;
 wire \Tile_X8Y12_FrameData_O[13] ;
 wire \Tile_X8Y12_FrameData_O[14] ;
 wire \Tile_X8Y12_FrameData_O[15] ;
 wire \Tile_X8Y12_FrameData_O[16] ;
 wire \Tile_X8Y12_FrameData_O[17] ;
 wire \Tile_X8Y12_FrameData_O[18] ;
 wire \Tile_X8Y12_FrameData_O[19] ;
 wire \Tile_X8Y12_FrameData_O[1] ;
 wire \Tile_X8Y12_FrameData_O[20] ;
 wire \Tile_X8Y12_FrameData_O[21] ;
 wire \Tile_X8Y12_FrameData_O[22] ;
 wire \Tile_X8Y12_FrameData_O[23] ;
 wire \Tile_X8Y12_FrameData_O[24] ;
 wire \Tile_X8Y12_FrameData_O[25] ;
 wire \Tile_X8Y12_FrameData_O[26] ;
 wire \Tile_X8Y12_FrameData_O[27] ;
 wire \Tile_X8Y12_FrameData_O[28] ;
 wire \Tile_X8Y12_FrameData_O[29] ;
 wire \Tile_X8Y12_FrameData_O[2] ;
 wire \Tile_X8Y12_FrameData_O[30] ;
 wire \Tile_X8Y12_FrameData_O[31] ;
 wire \Tile_X8Y12_FrameData_O[3] ;
 wire \Tile_X8Y12_FrameData_O[4] ;
 wire \Tile_X8Y12_FrameData_O[5] ;
 wire \Tile_X8Y12_FrameData_O[6] ;
 wire \Tile_X8Y12_FrameData_O[7] ;
 wire \Tile_X8Y12_FrameData_O[8] ;
 wire \Tile_X8Y12_FrameData_O[9] ;
 wire \Tile_X8Y12_FrameStrobe_O[0] ;
 wire \Tile_X8Y12_FrameStrobe_O[10] ;
 wire \Tile_X8Y12_FrameStrobe_O[11] ;
 wire \Tile_X8Y12_FrameStrobe_O[12] ;
 wire \Tile_X8Y12_FrameStrobe_O[13] ;
 wire \Tile_X8Y12_FrameStrobe_O[14] ;
 wire \Tile_X8Y12_FrameStrobe_O[15] ;
 wire \Tile_X8Y12_FrameStrobe_O[16] ;
 wire \Tile_X8Y12_FrameStrobe_O[17] ;
 wire \Tile_X8Y12_FrameStrobe_O[18] ;
 wire \Tile_X8Y12_FrameStrobe_O[19] ;
 wire \Tile_X8Y12_FrameStrobe_O[1] ;
 wire \Tile_X8Y12_FrameStrobe_O[2] ;
 wire \Tile_X8Y12_FrameStrobe_O[3] ;
 wire \Tile_X8Y12_FrameStrobe_O[4] ;
 wire \Tile_X8Y12_FrameStrobe_O[5] ;
 wire \Tile_X8Y12_FrameStrobe_O[6] ;
 wire \Tile_X8Y12_FrameStrobe_O[7] ;
 wire \Tile_X8Y12_FrameStrobe_O[8] ;
 wire \Tile_X8Y12_FrameStrobe_O[9] ;
 wire \Tile_X8Y12_N1BEG[0] ;
 wire \Tile_X8Y12_N1BEG[1] ;
 wire \Tile_X8Y12_N1BEG[2] ;
 wire \Tile_X8Y12_N1BEG[3] ;
 wire \Tile_X8Y12_N2BEG[0] ;
 wire \Tile_X8Y12_N2BEG[1] ;
 wire \Tile_X8Y12_N2BEG[2] ;
 wire \Tile_X8Y12_N2BEG[3] ;
 wire \Tile_X8Y12_N2BEG[4] ;
 wire \Tile_X8Y12_N2BEG[5] ;
 wire \Tile_X8Y12_N2BEG[6] ;
 wire \Tile_X8Y12_N2BEG[7] ;
 wire \Tile_X8Y12_N2BEGb[0] ;
 wire \Tile_X8Y12_N2BEGb[1] ;
 wire \Tile_X8Y12_N2BEGb[2] ;
 wire \Tile_X8Y12_N2BEGb[3] ;
 wire \Tile_X8Y12_N2BEGb[4] ;
 wire \Tile_X8Y12_N2BEGb[5] ;
 wire \Tile_X8Y12_N2BEGb[6] ;
 wire \Tile_X8Y12_N2BEGb[7] ;
 wire \Tile_X8Y12_N4BEG[0] ;
 wire \Tile_X8Y12_N4BEG[10] ;
 wire \Tile_X8Y12_N4BEG[11] ;
 wire \Tile_X8Y12_N4BEG[12] ;
 wire \Tile_X8Y12_N4BEG[13] ;
 wire \Tile_X8Y12_N4BEG[14] ;
 wire \Tile_X8Y12_N4BEG[15] ;
 wire \Tile_X8Y12_N4BEG[1] ;
 wire \Tile_X8Y12_N4BEG[2] ;
 wire \Tile_X8Y12_N4BEG[3] ;
 wire \Tile_X8Y12_N4BEG[4] ;
 wire \Tile_X8Y12_N4BEG[5] ;
 wire \Tile_X8Y12_N4BEG[6] ;
 wire \Tile_X8Y12_N4BEG[7] ;
 wire \Tile_X8Y12_N4BEG[8] ;
 wire \Tile_X8Y12_N4BEG[9] ;
 wire \Tile_X8Y12_NN4BEG[0] ;
 wire \Tile_X8Y12_NN4BEG[10] ;
 wire \Tile_X8Y12_NN4BEG[11] ;
 wire \Tile_X8Y12_NN4BEG[12] ;
 wire \Tile_X8Y12_NN4BEG[13] ;
 wire \Tile_X8Y12_NN4BEG[14] ;
 wire \Tile_X8Y12_NN4BEG[15] ;
 wire \Tile_X8Y12_NN4BEG[1] ;
 wire \Tile_X8Y12_NN4BEG[2] ;
 wire \Tile_X8Y12_NN4BEG[3] ;
 wire \Tile_X8Y12_NN4BEG[4] ;
 wire \Tile_X8Y12_NN4BEG[5] ;
 wire \Tile_X8Y12_NN4BEG[6] ;
 wire \Tile_X8Y12_NN4BEG[7] ;
 wire \Tile_X8Y12_NN4BEG[8] ;
 wire \Tile_X8Y12_NN4BEG[9] ;
 wire \Tile_X8Y12_S1BEG[0] ;
 wire \Tile_X8Y12_S1BEG[1] ;
 wire \Tile_X8Y12_S1BEG[2] ;
 wire \Tile_X8Y12_S1BEG[3] ;
 wire \Tile_X8Y12_S2BEG[0] ;
 wire \Tile_X8Y12_S2BEG[1] ;
 wire \Tile_X8Y12_S2BEG[2] ;
 wire \Tile_X8Y12_S2BEG[3] ;
 wire \Tile_X8Y12_S2BEG[4] ;
 wire \Tile_X8Y12_S2BEG[5] ;
 wire \Tile_X8Y12_S2BEG[6] ;
 wire \Tile_X8Y12_S2BEG[7] ;
 wire \Tile_X8Y12_S2BEGb[0] ;
 wire \Tile_X8Y12_S2BEGb[1] ;
 wire \Tile_X8Y12_S2BEGb[2] ;
 wire \Tile_X8Y12_S2BEGb[3] ;
 wire \Tile_X8Y12_S2BEGb[4] ;
 wire \Tile_X8Y12_S2BEGb[5] ;
 wire \Tile_X8Y12_S2BEGb[6] ;
 wire \Tile_X8Y12_S2BEGb[7] ;
 wire \Tile_X8Y12_S4BEG[0] ;
 wire \Tile_X8Y12_S4BEG[10] ;
 wire \Tile_X8Y12_S4BEG[11] ;
 wire \Tile_X8Y12_S4BEG[12] ;
 wire \Tile_X8Y12_S4BEG[13] ;
 wire \Tile_X8Y12_S4BEG[14] ;
 wire \Tile_X8Y12_S4BEG[15] ;
 wire \Tile_X8Y12_S4BEG[1] ;
 wire \Tile_X8Y12_S4BEG[2] ;
 wire \Tile_X8Y12_S4BEG[3] ;
 wire \Tile_X8Y12_S4BEG[4] ;
 wire \Tile_X8Y12_S4BEG[5] ;
 wire \Tile_X8Y12_S4BEG[6] ;
 wire \Tile_X8Y12_S4BEG[7] ;
 wire \Tile_X8Y12_S4BEG[8] ;
 wire \Tile_X8Y12_S4BEG[9] ;
 wire \Tile_X8Y12_SS4BEG[0] ;
 wire \Tile_X8Y12_SS4BEG[10] ;
 wire \Tile_X8Y12_SS4BEG[11] ;
 wire \Tile_X8Y12_SS4BEG[12] ;
 wire \Tile_X8Y12_SS4BEG[13] ;
 wire \Tile_X8Y12_SS4BEG[14] ;
 wire \Tile_X8Y12_SS4BEG[15] ;
 wire \Tile_X8Y12_SS4BEG[1] ;
 wire \Tile_X8Y12_SS4BEG[2] ;
 wire \Tile_X8Y12_SS4BEG[3] ;
 wire \Tile_X8Y12_SS4BEG[4] ;
 wire \Tile_X8Y12_SS4BEG[5] ;
 wire \Tile_X8Y12_SS4BEG[6] ;
 wire \Tile_X8Y12_SS4BEG[7] ;
 wire \Tile_X8Y12_SS4BEG[8] ;
 wire \Tile_X8Y12_SS4BEG[9] ;
 wire Tile_X8Y12_UserCLKo;
 wire \Tile_X8Y12_W1BEG[0] ;
 wire \Tile_X8Y12_W1BEG[1] ;
 wire \Tile_X8Y12_W1BEG[2] ;
 wire \Tile_X8Y12_W1BEG[3] ;
 wire \Tile_X8Y12_W2BEG[0] ;
 wire \Tile_X8Y12_W2BEG[1] ;
 wire \Tile_X8Y12_W2BEG[2] ;
 wire \Tile_X8Y12_W2BEG[3] ;
 wire \Tile_X8Y12_W2BEG[4] ;
 wire \Tile_X8Y12_W2BEG[5] ;
 wire \Tile_X8Y12_W2BEG[6] ;
 wire \Tile_X8Y12_W2BEG[7] ;
 wire \Tile_X8Y12_W2BEGb[0] ;
 wire \Tile_X8Y12_W2BEGb[1] ;
 wire \Tile_X8Y12_W2BEGb[2] ;
 wire \Tile_X8Y12_W2BEGb[3] ;
 wire \Tile_X8Y12_W2BEGb[4] ;
 wire \Tile_X8Y12_W2BEGb[5] ;
 wire \Tile_X8Y12_W2BEGb[6] ;
 wire \Tile_X8Y12_W2BEGb[7] ;
 wire \Tile_X8Y12_W6BEG[0] ;
 wire \Tile_X8Y12_W6BEG[10] ;
 wire \Tile_X8Y12_W6BEG[11] ;
 wire \Tile_X8Y12_W6BEG[1] ;
 wire \Tile_X8Y12_W6BEG[2] ;
 wire \Tile_X8Y12_W6BEG[3] ;
 wire \Tile_X8Y12_W6BEG[4] ;
 wire \Tile_X8Y12_W6BEG[5] ;
 wire \Tile_X8Y12_W6BEG[6] ;
 wire \Tile_X8Y12_W6BEG[7] ;
 wire \Tile_X8Y12_W6BEG[8] ;
 wire \Tile_X8Y12_W6BEG[9] ;
 wire \Tile_X8Y12_WW4BEG[0] ;
 wire \Tile_X8Y12_WW4BEG[10] ;
 wire \Tile_X8Y12_WW4BEG[11] ;
 wire \Tile_X8Y12_WW4BEG[12] ;
 wire \Tile_X8Y12_WW4BEG[13] ;
 wire \Tile_X8Y12_WW4BEG[14] ;
 wire \Tile_X8Y12_WW4BEG[15] ;
 wire \Tile_X8Y12_WW4BEG[1] ;
 wire \Tile_X8Y12_WW4BEG[2] ;
 wire \Tile_X8Y12_WW4BEG[3] ;
 wire \Tile_X8Y12_WW4BEG[4] ;
 wire \Tile_X8Y12_WW4BEG[5] ;
 wire \Tile_X8Y12_WW4BEG[6] ;
 wire \Tile_X8Y12_WW4BEG[7] ;
 wire \Tile_X8Y12_WW4BEG[8] ;
 wire \Tile_X8Y12_WW4BEG[9] ;
 wire Tile_X8Y13_Co;
 wire \Tile_X8Y13_E1BEG[0] ;
 wire \Tile_X8Y13_E1BEG[1] ;
 wire \Tile_X8Y13_E1BEG[2] ;
 wire \Tile_X8Y13_E1BEG[3] ;
 wire \Tile_X8Y13_E2BEG[0] ;
 wire \Tile_X8Y13_E2BEG[1] ;
 wire \Tile_X8Y13_E2BEG[2] ;
 wire \Tile_X8Y13_E2BEG[3] ;
 wire \Tile_X8Y13_E2BEG[4] ;
 wire \Tile_X8Y13_E2BEG[5] ;
 wire \Tile_X8Y13_E2BEG[6] ;
 wire \Tile_X8Y13_E2BEG[7] ;
 wire \Tile_X8Y13_E2BEGb[0] ;
 wire \Tile_X8Y13_E2BEGb[1] ;
 wire \Tile_X8Y13_E2BEGb[2] ;
 wire \Tile_X8Y13_E2BEGb[3] ;
 wire \Tile_X8Y13_E2BEGb[4] ;
 wire \Tile_X8Y13_E2BEGb[5] ;
 wire \Tile_X8Y13_E2BEGb[6] ;
 wire \Tile_X8Y13_E2BEGb[7] ;
 wire \Tile_X8Y13_E6BEG[0] ;
 wire \Tile_X8Y13_E6BEG[10] ;
 wire \Tile_X8Y13_E6BEG[11] ;
 wire \Tile_X8Y13_E6BEG[1] ;
 wire \Tile_X8Y13_E6BEG[2] ;
 wire \Tile_X8Y13_E6BEG[3] ;
 wire \Tile_X8Y13_E6BEG[4] ;
 wire \Tile_X8Y13_E6BEG[5] ;
 wire \Tile_X8Y13_E6BEG[6] ;
 wire \Tile_X8Y13_E6BEG[7] ;
 wire \Tile_X8Y13_E6BEG[8] ;
 wire \Tile_X8Y13_E6BEG[9] ;
 wire \Tile_X8Y13_EE4BEG[0] ;
 wire \Tile_X8Y13_EE4BEG[10] ;
 wire \Tile_X8Y13_EE4BEG[11] ;
 wire \Tile_X8Y13_EE4BEG[12] ;
 wire \Tile_X8Y13_EE4BEG[13] ;
 wire \Tile_X8Y13_EE4BEG[14] ;
 wire \Tile_X8Y13_EE4BEG[15] ;
 wire \Tile_X8Y13_EE4BEG[1] ;
 wire \Tile_X8Y13_EE4BEG[2] ;
 wire \Tile_X8Y13_EE4BEG[3] ;
 wire \Tile_X8Y13_EE4BEG[4] ;
 wire \Tile_X8Y13_EE4BEG[5] ;
 wire \Tile_X8Y13_EE4BEG[6] ;
 wire \Tile_X8Y13_EE4BEG[7] ;
 wire \Tile_X8Y13_EE4BEG[8] ;
 wire \Tile_X8Y13_EE4BEG[9] ;
 wire \Tile_X8Y13_FrameData_O[0] ;
 wire \Tile_X8Y13_FrameData_O[10] ;
 wire \Tile_X8Y13_FrameData_O[11] ;
 wire \Tile_X8Y13_FrameData_O[12] ;
 wire \Tile_X8Y13_FrameData_O[13] ;
 wire \Tile_X8Y13_FrameData_O[14] ;
 wire \Tile_X8Y13_FrameData_O[15] ;
 wire \Tile_X8Y13_FrameData_O[16] ;
 wire \Tile_X8Y13_FrameData_O[17] ;
 wire \Tile_X8Y13_FrameData_O[18] ;
 wire \Tile_X8Y13_FrameData_O[19] ;
 wire \Tile_X8Y13_FrameData_O[1] ;
 wire \Tile_X8Y13_FrameData_O[20] ;
 wire \Tile_X8Y13_FrameData_O[21] ;
 wire \Tile_X8Y13_FrameData_O[22] ;
 wire \Tile_X8Y13_FrameData_O[23] ;
 wire \Tile_X8Y13_FrameData_O[24] ;
 wire \Tile_X8Y13_FrameData_O[25] ;
 wire \Tile_X8Y13_FrameData_O[26] ;
 wire \Tile_X8Y13_FrameData_O[27] ;
 wire \Tile_X8Y13_FrameData_O[28] ;
 wire \Tile_X8Y13_FrameData_O[29] ;
 wire \Tile_X8Y13_FrameData_O[2] ;
 wire \Tile_X8Y13_FrameData_O[30] ;
 wire \Tile_X8Y13_FrameData_O[31] ;
 wire \Tile_X8Y13_FrameData_O[3] ;
 wire \Tile_X8Y13_FrameData_O[4] ;
 wire \Tile_X8Y13_FrameData_O[5] ;
 wire \Tile_X8Y13_FrameData_O[6] ;
 wire \Tile_X8Y13_FrameData_O[7] ;
 wire \Tile_X8Y13_FrameData_O[8] ;
 wire \Tile_X8Y13_FrameData_O[9] ;
 wire \Tile_X8Y13_FrameStrobe_O[0] ;
 wire \Tile_X8Y13_FrameStrobe_O[10] ;
 wire \Tile_X8Y13_FrameStrobe_O[11] ;
 wire \Tile_X8Y13_FrameStrobe_O[12] ;
 wire \Tile_X8Y13_FrameStrobe_O[13] ;
 wire \Tile_X8Y13_FrameStrobe_O[14] ;
 wire \Tile_X8Y13_FrameStrobe_O[15] ;
 wire \Tile_X8Y13_FrameStrobe_O[16] ;
 wire \Tile_X8Y13_FrameStrobe_O[17] ;
 wire \Tile_X8Y13_FrameStrobe_O[18] ;
 wire \Tile_X8Y13_FrameStrobe_O[19] ;
 wire \Tile_X8Y13_FrameStrobe_O[1] ;
 wire \Tile_X8Y13_FrameStrobe_O[2] ;
 wire \Tile_X8Y13_FrameStrobe_O[3] ;
 wire \Tile_X8Y13_FrameStrobe_O[4] ;
 wire \Tile_X8Y13_FrameStrobe_O[5] ;
 wire \Tile_X8Y13_FrameStrobe_O[6] ;
 wire \Tile_X8Y13_FrameStrobe_O[7] ;
 wire \Tile_X8Y13_FrameStrobe_O[8] ;
 wire \Tile_X8Y13_FrameStrobe_O[9] ;
 wire \Tile_X8Y13_N1BEG[0] ;
 wire \Tile_X8Y13_N1BEG[1] ;
 wire \Tile_X8Y13_N1BEG[2] ;
 wire \Tile_X8Y13_N1BEG[3] ;
 wire \Tile_X8Y13_N2BEG[0] ;
 wire \Tile_X8Y13_N2BEG[1] ;
 wire \Tile_X8Y13_N2BEG[2] ;
 wire \Tile_X8Y13_N2BEG[3] ;
 wire \Tile_X8Y13_N2BEG[4] ;
 wire \Tile_X8Y13_N2BEG[5] ;
 wire \Tile_X8Y13_N2BEG[6] ;
 wire \Tile_X8Y13_N2BEG[7] ;
 wire \Tile_X8Y13_N2BEGb[0] ;
 wire \Tile_X8Y13_N2BEGb[1] ;
 wire \Tile_X8Y13_N2BEGb[2] ;
 wire \Tile_X8Y13_N2BEGb[3] ;
 wire \Tile_X8Y13_N2BEGb[4] ;
 wire \Tile_X8Y13_N2BEGb[5] ;
 wire \Tile_X8Y13_N2BEGb[6] ;
 wire \Tile_X8Y13_N2BEGb[7] ;
 wire \Tile_X8Y13_N4BEG[0] ;
 wire \Tile_X8Y13_N4BEG[10] ;
 wire \Tile_X8Y13_N4BEG[11] ;
 wire \Tile_X8Y13_N4BEG[12] ;
 wire \Tile_X8Y13_N4BEG[13] ;
 wire \Tile_X8Y13_N4BEG[14] ;
 wire \Tile_X8Y13_N4BEG[15] ;
 wire \Tile_X8Y13_N4BEG[1] ;
 wire \Tile_X8Y13_N4BEG[2] ;
 wire \Tile_X8Y13_N4BEG[3] ;
 wire \Tile_X8Y13_N4BEG[4] ;
 wire \Tile_X8Y13_N4BEG[5] ;
 wire \Tile_X8Y13_N4BEG[6] ;
 wire \Tile_X8Y13_N4BEG[7] ;
 wire \Tile_X8Y13_N4BEG[8] ;
 wire \Tile_X8Y13_N4BEG[9] ;
 wire \Tile_X8Y13_NN4BEG[0] ;
 wire \Tile_X8Y13_NN4BEG[10] ;
 wire \Tile_X8Y13_NN4BEG[11] ;
 wire \Tile_X8Y13_NN4BEG[12] ;
 wire \Tile_X8Y13_NN4BEG[13] ;
 wire \Tile_X8Y13_NN4BEG[14] ;
 wire \Tile_X8Y13_NN4BEG[15] ;
 wire \Tile_X8Y13_NN4BEG[1] ;
 wire \Tile_X8Y13_NN4BEG[2] ;
 wire \Tile_X8Y13_NN4BEG[3] ;
 wire \Tile_X8Y13_NN4BEG[4] ;
 wire \Tile_X8Y13_NN4BEG[5] ;
 wire \Tile_X8Y13_NN4BEG[6] ;
 wire \Tile_X8Y13_NN4BEG[7] ;
 wire \Tile_X8Y13_NN4BEG[8] ;
 wire \Tile_X8Y13_NN4BEG[9] ;
 wire \Tile_X8Y13_S1BEG[0] ;
 wire \Tile_X8Y13_S1BEG[1] ;
 wire \Tile_X8Y13_S1BEG[2] ;
 wire \Tile_X8Y13_S1BEG[3] ;
 wire \Tile_X8Y13_S2BEG[0] ;
 wire \Tile_X8Y13_S2BEG[1] ;
 wire \Tile_X8Y13_S2BEG[2] ;
 wire \Tile_X8Y13_S2BEG[3] ;
 wire \Tile_X8Y13_S2BEG[4] ;
 wire \Tile_X8Y13_S2BEG[5] ;
 wire \Tile_X8Y13_S2BEG[6] ;
 wire \Tile_X8Y13_S2BEG[7] ;
 wire \Tile_X8Y13_S2BEGb[0] ;
 wire \Tile_X8Y13_S2BEGb[1] ;
 wire \Tile_X8Y13_S2BEGb[2] ;
 wire \Tile_X8Y13_S2BEGb[3] ;
 wire \Tile_X8Y13_S2BEGb[4] ;
 wire \Tile_X8Y13_S2BEGb[5] ;
 wire \Tile_X8Y13_S2BEGb[6] ;
 wire \Tile_X8Y13_S2BEGb[7] ;
 wire \Tile_X8Y13_S4BEG[0] ;
 wire \Tile_X8Y13_S4BEG[10] ;
 wire \Tile_X8Y13_S4BEG[11] ;
 wire \Tile_X8Y13_S4BEG[12] ;
 wire \Tile_X8Y13_S4BEG[13] ;
 wire \Tile_X8Y13_S4BEG[14] ;
 wire \Tile_X8Y13_S4BEG[15] ;
 wire \Tile_X8Y13_S4BEG[1] ;
 wire \Tile_X8Y13_S4BEG[2] ;
 wire \Tile_X8Y13_S4BEG[3] ;
 wire \Tile_X8Y13_S4BEG[4] ;
 wire \Tile_X8Y13_S4BEG[5] ;
 wire \Tile_X8Y13_S4BEG[6] ;
 wire \Tile_X8Y13_S4BEG[7] ;
 wire \Tile_X8Y13_S4BEG[8] ;
 wire \Tile_X8Y13_S4BEG[9] ;
 wire \Tile_X8Y13_SS4BEG[0] ;
 wire \Tile_X8Y13_SS4BEG[10] ;
 wire \Tile_X8Y13_SS4BEG[11] ;
 wire \Tile_X8Y13_SS4BEG[12] ;
 wire \Tile_X8Y13_SS4BEG[13] ;
 wire \Tile_X8Y13_SS4BEG[14] ;
 wire \Tile_X8Y13_SS4BEG[15] ;
 wire \Tile_X8Y13_SS4BEG[1] ;
 wire \Tile_X8Y13_SS4BEG[2] ;
 wire \Tile_X8Y13_SS4BEG[3] ;
 wire \Tile_X8Y13_SS4BEG[4] ;
 wire \Tile_X8Y13_SS4BEG[5] ;
 wire \Tile_X8Y13_SS4BEG[6] ;
 wire \Tile_X8Y13_SS4BEG[7] ;
 wire \Tile_X8Y13_SS4BEG[8] ;
 wire \Tile_X8Y13_SS4BEG[9] ;
 wire Tile_X8Y13_UserCLKo;
 wire \Tile_X8Y13_W1BEG[0] ;
 wire \Tile_X8Y13_W1BEG[1] ;
 wire \Tile_X8Y13_W1BEG[2] ;
 wire \Tile_X8Y13_W1BEG[3] ;
 wire \Tile_X8Y13_W2BEG[0] ;
 wire \Tile_X8Y13_W2BEG[1] ;
 wire \Tile_X8Y13_W2BEG[2] ;
 wire \Tile_X8Y13_W2BEG[3] ;
 wire \Tile_X8Y13_W2BEG[4] ;
 wire \Tile_X8Y13_W2BEG[5] ;
 wire \Tile_X8Y13_W2BEG[6] ;
 wire \Tile_X8Y13_W2BEG[7] ;
 wire \Tile_X8Y13_W2BEGb[0] ;
 wire \Tile_X8Y13_W2BEGb[1] ;
 wire \Tile_X8Y13_W2BEGb[2] ;
 wire \Tile_X8Y13_W2BEGb[3] ;
 wire \Tile_X8Y13_W2BEGb[4] ;
 wire \Tile_X8Y13_W2BEGb[5] ;
 wire \Tile_X8Y13_W2BEGb[6] ;
 wire \Tile_X8Y13_W2BEGb[7] ;
 wire \Tile_X8Y13_W6BEG[0] ;
 wire \Tile_X8Y13_W6BEG[10] ;
 wire \Tile_X8Y13_W6BEG[11] ;
 wire \Tile_X8Y13_W6BEG[1] ;
 wire \Tile_X8Y13_W6BEG[2] ;
 wire \Tile_X8Y13_W6BEG[3] ;
 wire \Tile_X8Y13_W6BEG[4] ;
 wire \Tile_X8Y13_W6BEG[5] ;
 wire \Tile_X8Y13_W6BEG[6] ;
 wire \Tile_X8Y13_W6BEG[7] ;
 wire \Tile_X8Y13_W6BEG[8] ;
 wire \Tile_X8Y13_W6BEG[9] ;
 wire \Tile_X8Y13_WW4BEG[0] ;
 wire \Tile_X8Y13_WW4BEG[10] ;
 wire \Tile_X8Y13_WW4BEG[11] ;
 wire \Tile_X8Y13_WW4BEG[12] ;
 wire \Tile_X8Y13_WW4BEG[13] ;
 wire \Tile_X8Y13_WW4BEG[14] ;
 wire \Tile_X8Y13_WW4BEG[15] ;
 wire \Tile_X8Y13_WW4BEG[1] ;
 wire \Tile_X8Y13_WW4BEG[2] ;
 wire \Tile_X8Y13_WW4BEG[3] ;
 wire \Tile_X8Y13_WW4BEG[4] ;
 wire \Tile_X8Y13_WW4BEG[5] ;
 wire \Tile_X8Y13_WW4BEG[6] ;
 wire \Tile_X8Y13_WW4BEG[7] ;
 wire \Tile_X8Y13_WW4BEG[8] ;
 wire \Tile_X8Y13_WW4BEG[9] ;
 wire Tile_X8Y14_Co;
 wire \Tile_X8Y14_E1BEG[0] ;
 wire \Tile_X8Y14_E1BEG[1] ;
 wire \Tile_X8Y14_E1BEG[2] ;
 wire \Tile_X8Y14_E1BEG[3] ;
 wire \Tile_X8Y14_E2BEG[0] ;
 wire \Tile_X8Y14_E2BEG[1] ;
 wire \Tile_X8Y14_E2BEG[2] ;
 wire \Tile_X8Y14_E2BEG[3] ;
 wire \Tile_X8Y14_E2BEG[4] ;
 wire \Tile_X8Y14_E2BEG[5] ;
 wire \Tile_X8Y14_E2BEG[6] ;
 wire \Tile_X8Y14_E2BEG[7] ;
 wire \Tile_X8Y14_E2BEGb[0] ;
 wire \Tile_X8Y14_E2BEGb[1] ;
 wire \Tile_X8Y14_E2BEGb[2] ;
 wire \Tile_X8Y14_E2BEGb[3] ;
 wire \Tile_X8Y14_E2BEGb[4] ;
 wire \Tile_X8Y14_E2BEGb[5] ;
 wire \Tile_X8Y14_E2BEGb[6] ;
 wire \Tile_X8Y14_E2BEGb[7] ;
 wire \Tile_X8Y14_E6BEG[0] ;
 wire \Tile_X8Y14_E6BEG[10] ;
 wire \Tile_X8Y14_E6BEG[11] ;
 wire \Tile_X8Y14_E6BEG[1] ;
 wire \Tile_X8Y14_E6BEG[2] ;
 wire \Tile_X8Y14_E6BEG[3] ;
 wire \Tile_X8Y14_E6BEG[4] ;
 wire \Tile_X8Y14_E6BEG[5] ;
 wire \Tile_X8Y14_E6BEG[6] ;
 wire \Tile_X8Y14_E6BEG[7] ;
 wire \Tile_X8Y14_E6BEG[8] ;
 wire \Tile_X8Y14_E6BEG[9] ;
 wire \Tile_X8Y14_EE4BEG[0] ;
 wire \Tile_X8Y14_EE4BEG[10] ;
 wire \Tile_X8Y14_EE4BEG[11] ;
 wire \Tile_X8Y14_EE4BEG[12] ;
 wire \Tile_X8Y14_EE4BEG[13] ;
 wire \Tile_X8Y14_EE4BEG[14] ;
 wire \Tile_X8Y14_EE4BEG[15] ;
 wire \Tile_X8Y14_EE4BEG[1] ;
 wire \Tile_X8Y14_EE4BEG[2] ;
 wire \Tile_X8Y14_EE4BEG[3] ;
 wire \Tile_X8Y14_EE4BEG[4] ;
 wire \Tile_X8Y14_EE4BEG[5] ;
 wire \Tile_X8Y14_EE4BEG[6] ;
 wire \Tile_X8Y14_EE4BEG[7] ;
 wire \Tile_X8Y14_EE4BEG[8] ;
 wire \Tile_X8Y14_EE4BEG[9] ;
 wire \Tile_X8Y14_FrameData_O[0] ;
 wire \Tile_X8Y14_FrameData_O[10] ;
 wire \Tile_X8Y14_FrameData_O[11] ;
 wire \Tile_X8Y14_FrameData_O[12] ;
 wire \Tile_X8Y14_FrameData_O[13] ;
 wire \Tile_X8Y14_FrameData_O[14] ;
 wire \Tile_X8Y14_FrameData_O[15] ;
 wire \Tile_X8Y14_FrameData_O[16] ;
 wire \Tile_X8Y14_FrameData_O[17] ;
 wire \Tile_X8Y14_FrameData_O[18] ;
 wire \Tile_X8Y14_FrameData_O[19] ;
 wire \Tile_X8Y14_FrameData_O[1] ;
 wire \Tile_X8Y14_FrameData_O[20] ;
 wire \Tile_X8Y14_FrameData_O[21] ;
 wire \Tile_X8Y14_FrameData_O[22] ;
 wire \Tile_X8Y14_FrameData_O[23] ;
 wire \Tile_X8Y14_FrameData_O[24] ;
 wire \Tile_X8Y14_FrameData_O[25] ;
 wire \Tile_X8Y14_FrameData_O[26] ;
 wire \Tile_X8Y14_FrameData_O[27] ;
 wire \Tile_X8Y14_FrameData_O[28] ;
 wire \Tile_X8Y14_FrameData_O[29] ;
 wire \Tile_X8Y14_FrameData_O[2] ;
 wire \Tile_X8Y14_FrameData_O[30] ;
 wire \Tile_X8Y14_FrameData_O[31] ;
 wire \Tile_X8Y14_FrameData_O[3] ;
 wire \Tile_X8Y14_FrameData_O[4] ;
 wire \Tile_X8Y14_FrameData_O[5] ;
 wire \Tile_X8Y14_FrameData_O[6] ;
 wire \Tile_X8Y14_FrameData_O[7] ;
 wire \Tile_X8Y14_FrameData_O[8] ;
 wire \Tile_X8Y14_FrameData_O[9] ;
 wire \Tile_X8Y14_FrameStrobe_O[0] ;
 wire \Tile_X8Y14_FrameStrobe_O[10] ;
 wire \Tile_X8Y14_FrameStrobe_O[11] ;
 wire \Tile_X8Y14_FrameStrobe_O[12] ;
 wire \Tile_X8Y14_FrameStrobe_O[13] ;
 wire \Tile_X8Y14_FrameStrobe_O[14] ;
 wire \Tile_X8Y14_FrameStrobe_O[15] ;
 wire \Tile_X8Y14_FrameStrobe_O[16] ;
 wire \Tile_X8Y14_FrameStrobe_O[17] ;
 wire \Tile_X8Y14_FrameStrobe_O[18] ;
 wire \Tile_X8Y14_FrameStrobe_O[19] ;
 wire \Tile_X8Y14_FrameStrobe_O[1] ;
 wire \Tile_X8Y14_FrameStrobe_O[2] ;
 wire \Tile_X8Y14_FrameStrobe_O[3] ;
 wire \Tile_X8Y14_FrameStrobe_O[4] ;
 wire \Tile_X8Y14_FrameStrobe_O[5] ;
 wire \Tile_X8Y14_FrameStrobe_O[6] ;
 wire \Tile_X8Y14_FrameStrobe_O[7] ;
 wire \Tile_X8Y14_FrameStrobe_O[8] ;
 wire \Tile_X8Y14_FrameStrobe_O[9] ;
 wire \Tile_X8Y14_N1BEG[0] ;
 wire \Tile_X8Y14_N1BEG[1] ;
 wire \Tile_X8Y14_N1BEG[2] ;
 wire \Tile_X8Y14_N1BEG[3] ;
 wire \Tile_X8Y14_N2BEG[0] ;
 wire \Tile_X8Y14_N2BEG[1] ;
 wire \Tile_X8Y14_N2BEG[2] ;
 wire \Tile_X8Y14_N2BEG[3] ;
 wire \Tile_X8Y14_N2BEG[4] ;
 wire \Tile_X8Y14_N2BEG[5] ;
 wire \Tile_X8Y14_N2BEG[6] ;
 wire \Tile_X8Y14_N2BEG[7] ;
 wire \Tile_X8Y14_N2BEGb[0] ;
 wire \Tile_X8Y14_N2BEGb[1] ;
 wire \Tile_X8Y14_N2BEGb[2] ;
 wire \Tile_X8Y14_N2BEGb[3] ;
 wire \Tile_X8Y14_N2BEGb[4] ;
 wire \Tile_X8Y14_N2BEGb[5] ;
 wire \Tile_X8Y14_N2BEGb[6] ;
 wire \Tile_X8Y14_N2BEGb[7] ;
 wire \Tile_X8Y14_N4BEG[0] ;
 wire \Tile_X8Y14_N4BEG[10] ;
 wire \Tile_X8Y14_N4BEG[11] ;
 wire \Tile_X8Y14_N4BEG[12] ;
 wire \Tile_X8Y14_N4BEG[13] ;
 wire \Tile_X8Y14_N4BEG[14] ;
 wire \Tile_X8Y14_N4BEG[15] ;
 wire \Tile_X8Y14_N4BEG[1] ;
 wire \Tile_X8Y14_N4BEG[2] ;
 wire \Tile_X8Y14_N4BEG[3] ;
 wire \Tile_X8Y14_N4BEG[4] ;
 wire \Tile_X8Y14_N4BEG[5] ;
 wire \Tile_X8Y14_N4BEG[6] ;
 wire \Tile_X8Y14_N4BEG[7] ;
 wire \Tile_X8Y14_N4BEG[8] ;
 wire \Tile_X8Y14_N4BEG[9] ;
 wire \Tile_X8Y14_NN4BEG[0] ;
 wire \Tile_X8Y14_NN4BEG[10] ;
 wire \Tile_X8Y14_NN4BEG[11] ;
 wire \Tile_X8Y14_NN4BEG[12] ;
 wire \Tile_X8Y14_NN4BEG[13] ;
 wire \Tile_X8Y14_NN4BEG[14] ;
 wire \Tile_X8Y14_NN4BEG[15] ;
 wire \Tile_X8Y14_NN4BEG[1] ;
 wire \Tile_X8Y14_NN4BEG[2] ;
 wire \Tile_X8Y14_NN4BEG[3] ;
 wire \Tile_X8Y14_NN4BEG[4] ;
 wire \Tile_X8Y14_NN4BEG[5] ;
 wire \Tile_X8Y14_NN4BEG[6] ;
 wire \Tile_X8Y14_NN4BEG[7] ;
 wire \Tile_X8Y14_NN4BEG[8] ;
 wire \Tile_X8Y14_NN4BEG[9] ;
 wire \Tile_X8Y14_S1BEG[0] ;
 wire \Tile_X8Y14_S1BEG[1] ;
 wire \Tile_X8Y14_S1BEG[2] ;
 wire \Tile_X8Y14_S1BEG[3] ;
 wire \Tile_X8Y14_S2BEG[0] ;
 wire \Tile_X8Y14_S2BEG[1] ;
 wire \Tile_X8Y14_S2BEG[2] ;
 wire \Tile_X8Y14_S2BEG[3] ;
 wire \Tile_X8Y14_S2BEG[4] ;
 wire \Tile_X8Y14_S2BEG[5] ;
 wire \Tile_X8Y14_S2BEG[6] ;
 wire \Tile_X8Y14_S2BEG[7] ;
 wire \Tile_X8Y14_S2BEGb[0] ;
 wire \Tile_X8Y14_S2BEGb[1] ;
 wire \Tile_X8Y14_S2BEGb[2] ;
 wire \Tile_X8Y14_S2BEGb[3] ;
 wire \Tile_X8Y14_S2BEGb[4] ;
 wire \Tile_X8Y14_S2BEGb[5] ;
 wire \Tile_X8Y14_S2BEGb[6] ;
 wire \Tile_X8Y14_S2BEGb[7] ;
 wire \Tile_X8Y14_S4BEG[0] ;
 wire \Tile_X8Y14_S4BEG[10] ;
 wire \Tile_X8Y14_S4BEG[11] ;
 wire \Tile_X8Y14_S4BEG[12] ;
 wire \Tile_X8Y14_S4BEG[13] ;
 wire \Tile_X8Y14_S4BEG[14] ;
 wire \Tile_X8Y14_S4BEG[15] ;
 wire \Tile_X8Y14_S4BEG[1] ;
 wire \Tile_X8Y14_S4BEG[2] ;
 wire \Tile_X8Y14_S4BEG[3] ;
 wire \Tile_X8Y14_S4BEG[4] ;
 wire \Tile_X8Y14_S4BEG[5] ;
 wire \Tile_X8Y14_S4BEG[6] ;
 wire \Tile_X8Y14_S4BEG[7] ;
 wire \Tile_X8Y14_S4BEG[8] ;
 wire \Tile_X8Y14_S4BEG[9] ;
 wire \Tile_X8Y14_SS4BEG[0] ;
 wire \Tile_X8Y14_SS4BEG[10] ;
 wire \Tile_X8Y14_SS4BEG[11] ;
 wire \Tile_X8Y14_SS4BEG[12] ;
 wire \Tile_X8Y14_SS4BEG[13] ;
 wire \Tile_X8Y14_SS4BEG[14] ;
 wire \Tile_X8Y14_SS4BEG[15] ;
 wire \Tile_X8Y14_SS4BEG[1] ;
 wire \Tile_X8Y14_SS4BEG[2] ;
 wire \Tile_X8Y14_SS4BEG[3] ;
 wire \Tile_X8Y14_SS4BEG[4] ;
 wire \Tile_X8Y14_SS4BEG[5] ;
 wire \Tile_X8Y14_SS4BEG[6] ;
 wire \Tile_X8Y14_SS4BEG[7] ;
 wire \Tile_X8Y14_SS4BEG[8] ;
 wire \Tile_X8Y14_SS4BEG[9] ;
 wire Tile_X8Y14_UserCLKo;
 wire \Tile_X8Y14_W1BEG[0] ;
 wire \Tile_X8Y14_W1BEG[1] ;
 wire \Tile_X8Y14_W1BEG[2] ;
 wire \Tile_X8Y14_W1BEG[3] ;
 wire \Tile_X8Y14_W2BEG[0] ;
 wire \Tile_X8Y14_W2BEG[1] ;
 wire \Tile_X8Y14_W2BEG[2] ;
 wire \Tile_X8Y14_W2BEG[3] ;
 wire \Tile_X8Y14_W2BEG[4] ;
 wire \Tile_X8Y14_W2BEG[5] ;
 wire \Tile_X8Y14_W2BEG[6] ;
 wire \Tile_X8Y14_W2BEG[7] ;
 wire \Tile_X8Y14_W2BEGb[0] ;
 wire \Tile_X8Y14_W2BEGb[1] ;
 wire \Tile_X8Y14_W2BEGb[2] ;
 wire \Tile_X8Y14_W2BEGb[3] ;
 wire \Tile_X8Y14_W2BEGb[4] ;
 wire \Tile_X8Y14_W2BEGb[5] ;
 wire \Tile_X8Y14_W2BEGb[6] ;
 wire \Tile_X8Y14_W2BEGb[7] ;
 wire \Tile_X8Y14_W6BEG[0] ;
 wire \Tile_X8Y14_W6BEG[10] ;
 wire \Tile_X8Y14_W6BEG[11] ;
 wire \Tile_X8Y14_W6BEG[1] ;
 wire \Tile_X8Y14_W6BEG[2] ;
 wire \Tile_X8Y14_W6BEG[3] ;
 wire \Tile_X8Y14_W6BEG[4] ;
 wire \Tile_X8Y14_W6BEG[5] ;
 wire \Tile_X8Y14_W6BEG[6] ;
 wire \Tile_X8Y14_W6BEG[7] ;
 wire \Tile_X8Y14_W6BEG[8] ;
 wire \Tile_X8Y14_W6BEG[9] ;
 wire \Tile_X8Y14_WW4BEG[0] ;
 wire \Tile_X8Y14_WW4BEG[10] ;
 wire \Tile_X8Y14_WW4BEG[11] ;
 wire \Tile_X8Y14_WW4BEG[12] ;
 wire \Tile_X8Y14_WW4BEG[13] ;
 wire \Tile_X8Y14_WW4BEG[14] ;
 wire \Tile_X8Y14_WW4BEG[15] ;
 wire \Tile_X8Y14_WW4BEG[1] ;
 wire \Tile_X8Y14_WW4BEG[2] ;
 wire \Tile_X8Y14_WW4BEG[3] ;
 wire \Tile_X8Y14_WW4BEG[4] ;
 wire \Tile_X8Y14_WW4BEG[5] ;
 wire \Tile_X8Y14_WW4BEG[6] ;
 wire \Tile_X8Y14_WW4BEG[7] ;
 wire \Tile_X8Y14_WW4BEG[8] ;
 wire \Tile_X8Y14_WW4BEG[9] ;
 wire Tile_X8Y15_Co;
 wire \Tile_X8Y15_FrameData_O[0] ;
 wire \Tile_X8Y15_FrameData_O[10] ;
 wire \Tile_X8Y15_FrameData_O[11] ;
 wire \Tile_X8Y15_FrameData_O[12] ;
 wire \Tile_X8Y15_FrameData_O[13] ;
 wire \Tile_X8Y15_FrameData_O[14] ;
 wire \Tile_X8Y15_FrameData_O[15] ;
 wire \Tile_X8Y15_FrameData_O[16] ;
 wire \Tile_X8Y15_FrameData_O[17] ;
 wire \Tile_X8Y15_FrameData_O[18] ;
 wire \Tile_X8Y15_FrameData_O[19] ;
 wire \Tile_X8Y15_FrameData_O[1] ;
 wire \Tile_X8Y15_FrameData_O[20] ;
 wire \Tile_X8Y15_FrameData_O[21] ;
 wire \Tile_X8Y15_FrameData_O[22] ;
 wire \Tile_X8Y15_FrameData_O[23] ;
 wire \Tile_X8Y15_FrameData_O[24] ;
 wire \Tile_X8Y15_FrameData_O[25] ;
 wire \Tile_X8Y15_FrameData_O[26] ;
 wire \Tile_X8Y15_FrameData_O[27] ;
 wire \Tile_X8Y15_FrameData_O[28] ;
 wire \Tile_X8Y15_FrameData_O[29] ;
 wire \Tile_X8Y15_FrameData_O[2] ;
 wire \Tile_X8Y15_FrameData_O[30] ;
 wire \Tile_X8Y15_FrameData_O[31] ;
 wire \Tile_X8Y15_FrameData_O[3] ;
 wire \Tile_X8Y15_FrameData_O[4] ;
 wire \Tile_X8Y15_FrameData_O[5] ;
 wire \Tile_X8Y15_FrameData_O[6] ;
 wire \Tile_X8Y15_FrameData_O[7] ;
 wire \Tile_X8Y15_FrameData_O[8] ;
 wire \Tile_X8Y15_FrameData_O[9] ;
 wire \Tile_X8Y15_FrameStrobe_O[0] ;
 wire \Tile_X8Y15_FrameStrobe_O[10] ;
 wire \Tile_X8Y15_FrameStrobe_O[11] ;
 wire \Tile_X8Y15_FrameStrobe_O[12] ;
 wire \Tile_X8Y15_FrameStrobe_O[13] ;
 wire \Tile_X8Y15_FrameStrobe_O[14] ;
 wire \Tile_X8Y15_FrameStrobe_O[15] ;
 wire \Tile_X8Y15_FrameStrobe_O[16] ;
 wire \Tile_X8Y15_FrameStrobe_O[17] ;
 wire \Tile_X8Y15_FrameStrobe_O[18] ;
 wire \Tile_X8Y15_FrameStrobe_O[19] ;
 wire \Tile_X8Y15_FrameStrobe_O[1] ;
 wire \Tile_X8Y15_FrameStrobe_O[2] ;
 wire \Tile_X8Y15_FrameStrobe_O[3] ;
 wire \Tile_X8Y15_FrameStrobe_O[4] ;
 wire \Tile_X8Y15_FrameStrobe_O[5] ;
 wire \Tile_X8Y15_FrameStrobe_O[6] ;
 wire \Tile_X8Y15_FrameStrobe_O[7] ;
 wire \Tile_X8Y15_FrameStrobe_O[8] ;
 wire \Tile_X8Y15_FrameStrobe_O[9] ;
 wire \Tile_X8Y15_N1BEG[0] ;
 wire \Tile_X8Y15_N1BEG[1] ;
 wire \Tile_X8Y15_N1BEG[2] ;
 wire \Tile_X8Y15_N1BEG[3] ;
 wire \Tile_X8Y15_N2BEG[0] ;
 wire \Tile_X8Y15_N2BEG[1] ;
 wire \Tile_X8Y15_N2BEG[2] ;
 wire \Tile_X8Y15_N2BEG[3] ;
 wire \Tile_X8Y15_N2BEG[4] ;
 wire \Tile_X8Y15_N2BEG[5] ;
 wire \Tile_X8Y15_N2BEG[6] ;
 wire \Tile_X8Y15_N2BEG[7] ;
 wire \Tile_X8Y15_N2BEGb[0] ;
 wire \Tile_X8Y15_N2BEGb[1] ;
 wire \Tile_X8Y15_N2BEGb[2] ;
 wire \Tile_X8Y15_N2BEGb[3] ;
 wire \Tile_X8Y15_N2BEGb[4] ;
 wire \Tile_X8Y15_N2BEGb[5] ;
 wire \Tile_X8Y15_N2BEGb[6] ;
 wire \Tile_X8Y15_N2BEGb[7] ;
 wire \Tile_X8Y15_N4BEG[0] ;
 wire \Tile_X8Y15_N4BEG[10] ;
 wire \Tile_X8Y15_N4BEG[11] ;
 wire \Tile_X8Y15_N4BEG[12] ;
 wire \Tile_X8Y15_N4BEG[13] ;
 wire \Tile_X8Y15_N4BEG[14] ;
 wire \Tile_X8Y15_N4BEG[15] ;
 wire \Tile_X8Y15_N4BEG[1] ;
 wire \Tile_X8Y15_N4BEG[2] ;
 wire \Tile_X8Y15_N4BEG[3] ;
 wire \Tile_X8Y15_N4BEG[4] ;
 wire \Tile_X8Y15_N4BEG[5] ;
 wire \Tile_X8Y15_N4BEG[6] ;
 wire \Tile_X8Y15_N4BEG[7] ;
 wire \Tile_X8Y15_N4BEG[8] ;
 wire \Tile_X8Y15_N4BEG[9] ;
 wire \Tile_X8Y15_NN4BEG[0] ;
 wire \Tile_X8Y15_NN4BEG[10] ;
 wire \Tile_X8Y15_NN4BEG[11] ;
 wire \Tile_X8Y15_NN4BEG[12] ;
 wire \Tile_X8Y15_NN4BEG[13] ;
 wire \Tile_X8Y15_NN4BEG[14] ;
 wire \Tile_X8Y15_NN4BEG[15] ;
 wire \Tile_X8Y15_NN4BEG[1] ;
 wire \Tile_X8Y15_NN4BEG[2] ;
 wire \Tile_X8Y15_NN4BEG[3] ;
 wire \Tile_X8Y15_NN4BEG[4] ;
 wire \Tile_X8Y15_NN4BEG[5] ;
 wire \Tile_X8Y15_NN4BEG[6] ;
 wire \Tile_X8Y15_NN4BEG[7] ;
 wire \Tile_X8Y15_NN4BEG[8] ;
 wire \Tile_X8Y15_NN4BEG[9] ;
 wire Tile_X8Y15_UserCLKo;
 wire Tile_X8Y1_Co;
 wire \Tile_X8Y1_E1BEG[0] ;
 wire \Tile_X8Y1_E1BEG[1] ;
 wire \Tile_X8Y1_E1BEG[2] ;
 wire \Tile_X8Y1_E1BEG[3] ;
 wire \Tile_X8Y1_E2BEG[0] ;
 wire \Tile_X8Y1_E2BEG[1] ;
 wire \Tile_X8Y1_E2BEG[2] ;
 wire \Tile_X8Y1_E2BEG[3] ;
 wire \Tile_X8Y1_E2BEG[4] ;
 wire \Tile_X8Y1_E2BEG[5] ;
 wire \Tile_X8Y1_E2BEG[6] ;
 wire \Tile_X8Y1_E2BEG[7] ;
 wire \Tile_X8Y1_E2BEGb[0] ;
 wire \Tile_X8Y1_E2BEGb[1] ;
 wire \Tile_X8Y1_E2BEGb[2] ;
 wire \Tile_X8Y1_E2BEGb[3] ;
 wire \Tile_X8Y1_E2BEGb[4] ;
 wire \Tile_X8Y1_E2BEGb[5] ;
 wire \Tile_X8Y1_E2BEGb[6] ;
 wire \Tile_X8Y1_E2BEGb[7] ;
 wire \Tile_X8Y1_E6BEG[0] ;
 wire \Tile_X8Y1_E6BEG[10] ;
 wire \Tile_X8Y1_E6BEG[11] ;
 wire \Tile_X8Y1_E6BEG[1] ;
 wire \Tile_X8Y1_E6BEG[2] ;
 wire \Tile_X8Y1_E6BEG[3] ;
 wire \Tile_X8Y1_E6BEG[4] ;
 wire \Tile_X8Y1_E6BEG[5] ;
 wire \Tile_X8Y1_E6BEG[6] ;
 wire \Tile_X8Y1_E6BEG[7] ;
 wire \Tile_X8Y1_E6BEG[8] ;
 wire \Tile_X8Y1_E6BEG[9] ;
 wire \Tile_X8Y1_EE4BEG[0] ;
 wire \Tile_X8Y1_EE4BEG[10] ;
 wire \Tile_X8Y1_EE4BEG[11] ;
 wire \Tile_X8Y1_EE4BEG[12] ;
 wire \Tile_X8Y1_EE4BEG[13] ;
 wire \Tile_X8Y1_EE4BEG[14] ;
 wire \Tile_X8Y1_EE4BEG[15] ;
 wire \Tile_X8Y1_EE4BEG[1] ;
 wire \Tile_X8Y1_EE4BEG[2] ;
 wire \Tile_X8Y1_EE4BEG[3] ;
 wire \Tile_X8Y1_EE4BEG[4] ;
 wire \Tile_X8Y1_EE4BEG[5] ;
 wire \Tile_X8Y1_EE4BEG[6] ;
 wire \Tile_X8Y1_EE4BEG[7] ;
 wire \Tile_X8Y1_EE4BEG[8] ;
 wire \Tile_X8Y1_EE4BEG[9] ;
 wire \Tile_X8Y1_FrameData_O[0] ;
 wire \Tile_X8Y1_FrameData_O[10] ;
 wire \Tile_X8Y1_FrameData_O[11] ;
 wire \Tile_X8Y1_FrameData_O[12] ;
 wire \Tile_X8Y1_FrameData_O[13] ;
 wire \Tile_X8Y1_FrameData_O[14] ;
 wire \Tile_X8Y1_FrameData_O[15] ;
 wire \Tile_X8Y1_FrameData_O[16] ;
 wire \Tile_X8Y1_FrameData_O[17] ;
 wire \Tile_X8Y1_FrameData_O[18] ;
 wire \Tile_X8Y1_FrameData_O[19] ;
 wire \Tile_X8Y1_FrameData_O[1] ;
 wire \Tile_X8Y1_FrameData_O[20] ;
 wire \Tile_X8Y1_FrameData_O[21] ;
 wire \Tile_X8Y1_FrameData_O[22] ;
 wire \Tile_X8Y1_FrameData_O[23] ;
 wire \Tile_X8Y1_FrameData_O[24] ;
 wire \Tile_X8Y1_FrameData_O[25] ;
 wire \Tile_X8Y1_FrameData_O[26] ;
 wire \Tile_X8Y1_FrameData_O[27] ;
 wire \Tile_X8Y1_FrameData_O[28] ;
 wire \Tile_X8Y1_FrameData_O[29] ;
 wire \Tile_X8Y1_FrameData_O[2] ;
 wire \Tile_X8Y1_FrameData_O[30] ;
 wire \Tile_X8Y1_FrameData_O[31] ;
 wire \Tile_X8Y1_FrameData_O[3] ;
 wire \Tile_X8Y1_FrameData_O[4] ;
 wire \Tile_X8Y1_FrameData_O[5] ;
 wire \Tile_X8Y1_FrameData_O[6] ;
 wire \Tile_X8Y1_FrameData_O[7] ;
 wire \Tile_X8Y1_FrameData_O[8] ;
 wire \Tile_X8Y1_FrameData_O[9] ;
 wire \Tile_X8Y1_FrameStrobe_O[0] ;
 wire \Tile_X8Y1_FrameStrobe_O[10] ;
 wire \Tile_X8Y1_FrameStrobe_O[11] ;
 wire \Tile_X8Y1_FrameStrobe_O[12] ;
 wire \Tile_X8Y1_FrameStrobe_O[13] ;
 wire \Tile_X8Y1_FrameStrobe_O[14] ;
 wire \Tile_X8Y1_FrameStrobe_O[15] ;
 wire \Tile_X8Y1_FrameStrobe_O[16] ;
 wire \Tile_X8Y1_FrameStrobe_O[17] ;
 wire \Tile_X8Y1_FrameStrobe_O[18] ;
 wire \Tile_X8Y1_FrameStrobe_O[19] ;
 wire \Tile_X8Y1_FrameStrobe_O[1] ;
 wire \Tile_X8Y1_FrameStrobe_O[2] ;
 wire \Tile_X8Y1_FrameStrobe_O[3] ;
 wire \Tile_X8Y1_FrameStrobe_O[4] ;
 wire \Tile_X8Y1_FrameStrobe_O[5] ;
 wire \Tile_X8Y1_FrameStrobe_O[6] ;
 wire \Tile_X8Y1_FrameStrobe_O[7] ;
 wire \Tile_X8Y1_FrameStrobe_O[8] ;
 wire \Tile_X8Y1_FrameStrobe_O[9] ;
 wire \Tile_X8Y1_N1BEG[0] ;
 wire \Tile_X8Y1_N1BEG[1] ;
 wire \Tile_X8Y1_N1BEG[2] ;
 wire \Tile_X8Y1_N1BEG[3] ;
 wire \Tile_X8Y1_N2BEG[0] ;
 wire \Tile_X8Y1_N2BEG[1] ;
 wire \Tile_X8Y1_N2BEG[2] ;
 wire \Tile_X8Y1_N2BEG[3] ;
 wire \Tile_X8Y1_N2BEG[4] ;
 wire \Tile_X8Y1_N2BEG[5] ;
 wire \Tile_X8Y1_N2BEG[6] ;
 wire \Tile_X8Y1_N2BEG[7] ;
 wire \Tile_X8Y1_N2BEGb[0] ;
 wire \Tile_X8Y1_N2BEGb[1] ;
 wire \Tile_X8Y1_N2BEGb[2] ;
 wire \Tile_X8Y1_N2BEGb[3] ;
 wire \Tile_X8Y1_N2BEGb[4] ;
 wire \Tile_X8Y1_N2BEGb[5] ;
 wire \Tile_X8Y1_N2BEGb[6] ;
 wire \Tile_X8Y1_N2BEGb[7] ;
 wire \Tile_X8Y1_N4BEG[0] ;
 wire \Tile_X8Y1_N4BEG[10] ;
 wire \Tile_X8Y1_N4BEG[11] ;
 wire \Tile_X8Y1_N4BEG[12] ;
 wire \Tile_X8Y1_N4BEG[13] ;
 wire \Tile_X8Y1_N4BEG[14] ;
 wire \Tile_X8Y1_N4BEG[15] ;
 wire \Tile_X8Y1_N4BEG[1] ;
 wire \Tile_X8Y1_N4BEG[2] ;
 wire \Tile_X8Y1_N4BEG[3] ;
 wire \Tile_X8Y1_N4BEG[4] ;
 wire \Tile_X8Y1_N4BEG[5] ;
 wire \Tile_X8Y1_N4BEG[6] ;
 wire \Tile_X8Y1_N4BEG[7] ;
 wire \Tile_X8Y1_N4BEG[8] ;
 wire \Tile_X8Y1_N4BEG[9] ;
 wire \Tile_X8Y1_NN4BEG[0] ;
 wire \Tile_X8Y1_NN4BEG[10] ;
 wire \Tile_X8Y1_NN4BEG[11] ;
 wire \Tile_X8Y1_NN4BEG[12] ;
 wire \Tile_X8Y1_NN4BEG[13] ;
 wire \Tile_X8Y1_NN4BEG[14] ;
 wire \Tile_X8Y1_NN4BEG[15] ;
 wire \Tile_X8Y1_NN4BEG[1] ;
 wire \Tile_X8Y1_NN4BEG[2] ;
 wire \Tile_X8Y1_NN4BEG[3] ;
 wire \Tile_X8Y1_NN4BEG[4] ;
 wire \Tile_X8Y1_NN4BEG[5] ;
 wire \Tile_X8Y1_NN4BEG[6] ;
 wire \Tile_X8Y1_NN4BEG[7] ;
 wire \Tile_X8Y1_NN4BEG[8] ;
 wire \Tile_X8Y1_NN4BEG[9] ;
 wire \Tile_X8Y1_S1BEG[0] ;
 wire \Tile_X8Y1_S1BEG[1] ;
 wire \Tile_X8Y1_S1BEG[2] ;
 wire \Tile_X8Y1_S1BEG[3] ;
 wire \Tile_X8Y1_S2BEG[0] ;
 wire \Tile_X8Y1_S2BEG[1] ;
 wire \Tile_X8Y1_S2BEG[2] ;
 wire \Tile_X8Y1_S2BEG[3] ;
 wire \Tile_X8Y1_S2BEG[4] ;
 wire \Tile_X8Y1_S2BEG[5] ;
 wire \Tile_X8Y1_S2BEG[6] ;
 wire \Tile_X8Y1_S2BEG[7] ;
 wire \Tile_X8Y1_S2BEGb[0] ;
 wire \Tile_X8Y1_S2BEGb[1] ;
 wire \Tile_X8Y1_S2BEGb[2] ;
 wire \Tile_X8Y1_S2BEGb[3] ;
 wire \Tile_X8Y1_S2BEGb[4] ;
 wire \Tile_X8Y1_S2BEGb[5] ;
 wire \Tile_X8Y1_S2BEGb[6] ;
 wire \Tile_X8Y1_S2BEGb[7] ;
 wire \Tile_X8Y1_S4BEG[0] ;
 wire \Tile_X8Y1_S4BEG[10] ;
 wire \Tile_X8Y1_S4BEG[11] ;
 wire \Tile_X8Y1_S4BEG[12] ;
 wire \Tile_X8Y1_S4BEG[13] ;
 wire \Tile_X8Y1_S4BEG[14] ;
 wire \Tile_X8Y1_S4BEG[15] ;
 wire \Tile_X8Y1_S4BEG[1] ;
 wire \Tile_X8Y1_S4BEG[2] ;
 wire \Tile_X8Y1_S4BEG[3] ;
 wire \Tile_X8Y1_S4BEG[4] ;
 wire \Tile_X8Y1_S4BEG[5] ;
 wire \Tile_X8Y1_S4BEG[6] ;
 wire \Tile_X8Y1_S4BEG[7] ;
 wire \Tile_X8Y1_S4BEG[8] ;
 wire \Tile_X8Y1_S4BEG[9] ;
 wire \Tile_X8Y1_SS4BEG[0] ;
 wire \Tile_X8Y1_SS4BEG[10] ;
 wire \Tile_X8Y1_SS4BEG[11] ;
 wire \Tile_X8Y1_SS4BEG[12] ;
 wire \Tile_X8Y1_SS4BEG[13] ;
 wire \Tile_X8Y1_SS4BEG[14] ;
 wire \Tile_X8Y1_SS4BEG[15] ;
 wire \Tile_X8Y1_SS4BEG[1] ;
 wire \Tile_X8Y1_SS4BEG[2] ;
 wire \Tile_X8Y1_SS4BEG[3] ;
 wire \Tile_X8Y1_SS4BEG[4] ;
 wire \Tile_X8Y1_SS4BEG[5] ;
 wire \Tile_X8Y1_SS4BEG[6] ;
 wire \Tile_X8Y1_SS4BEG[7] ;
 wire \Tile_X8Y1_SS4BEG[8] ;
 wire \Tile_X8Y1_SS4BEG[9] ;
 wire Tile_X8Y1_UserCLKo;
 wire \Tile_X8Y1_W1BEG[0] ;
 wire \Tile_X8Y1_W1BEG[1] ;
 wire \Tile_X8Y1_W1BEG[2] ;
 wire \Tile_X8Y1_W1BEG[3] ;
 wire \Tile_X8Y1_W2BEG[0] ;
 wire \Tile_X8Y1_W2BEG[1] ;
 wire \Tile_X8Y1_W2BEG[2] ;
 wire \Tile_X8Y1_W2BEG[3] ;
 wire \Tile_X8Y1_W2BEG[4] ;
 wire \Tile_X8Y1_W2BEG[5] ;
 wire \Tile_X8Y1_W2BEG[6] ;
 wire \Tile_X8Y1_W2BEG[7] ;
 wire \Tile_X8Y1_W2BEGb[0] ;
 wire \Tile_X8Y1_W2BEGb[1] ;
 wire \Tile_X8Y1_W2BEGb[2] ;
 wire \Tile_X8Y1_W2BEGb[3] ;
 wire \Tile_X8Y1_W2BEGb[4] ;
 wire \Tile_X8Y1_W2BEGb[5] ;
 wire \Tile_X8Y1_W2BEGb[6] ;
 wire \Tile_X8Y1_W2BEGb[7] ;
 wire \Tile_X8Y1_W6BEG[0] ;
 wire \Tile_X8Y1_W6BEG[10] ;
 wire \Tile_X8Y1_W6BEG[11] ;
 wire \Tile_X8Y1_W6BEG[1] ;
 wire \Tile_X8Y1_W6BEG[2] ;
 wire \Tile_X8Y1_W6BEG[3] ;
 wire \Tile_X8Y1_W6BEG[4] ;
 wire \Tile_X8Y1_W6BEG[5] ;
 wire \Tile_X8Y1_W6BEG[6] ;
 wire \Tile_X8Y1_W6BEG[7] ;
 wire \Tile_X8Y1_W6BEG[8] ;
 wire \Tile_X8Y1_W6BEG[9] ;
 wire \Tile_X8Y1_WW4BEG[0] ;
 wire \Tile_X8Y1_WW4BEG[10] ;
 wire \Tile_X8Y1_WW4BEG[11] ;
 wire \Tile_X8Y1_WW4BEG[12] ;
 wire \Tile_X8Y1_WW4BEG[13] ;
 wire \Tile_X8Y1_WW4BEG[14] ;
 wire \Tile_X8Y1_WW4BEG[15] ;
 wire \Tile_X8Y1_WW4BEG[1] ;
 wire \Tile_X8Y1_WW4BEG[2] ;
 wire \Tile_X8Y1_WW4BEG[3] ;
 wire \Tile_X8Y1_WW4BEG[4] ;
 wire \Tile_X8Y1_WW4BEG[5] ;
 wire \Tile_X8Y1_WW4BEG[6] ;
 wire \Tile_X8Y1_WW4BEG[7] ;
 wire \Tile_X8Y1_WW4BEG[8] ;
 wire \Tile_X8Y1_WW4BEG[9] ;
 wire Tile_X8Y2_Co;
 wire \Tile_X8Y2_E1BEG[0] ;
 wire \Tile_X8Y2_E1BEG[1] ;
 wire \Tile_X8Y2_E1BEG[2] ;
 wire \Tile_X8Y2_E1BEG[3] ;
 wire \Tile_X8Y2_E2BEG[0] ;
 wire \Tile_X8Y2_E2BEG[1] ;
 wire \Tile_X8Y2_E2BEG[2] ;
 wire \Tile_X8Y2_E2BEG[3] ;
 wire \Tile_X8Y2_E2BEG[4] ;
 wire \Tile_X8Y2_E2BEG[5] ;
 wire \Tile_X8Y2_E2BEG[6] ;
 wire \Tile_X8Y2_E2BEG[7] ;
 wire \Tile_X8Y2_E2BEGb[0] ;
 wire \Tile_X8Y2_E2BEGb[1] ;
 wire \Tile_X8Y2_E2BEGb[2] ;
 wire \Tile_X8Y2_E2BEGb[3] ;
 wire \Tile_X8Y2_E2BEGb[4] ;
 wire \Tile_X8Y2_E2BEGb[5] ;
 wire \Tile_X8Y2_E2BEGb[6] ;
 wire \Tile_X8Y2_E2BEGb[7] ;
 wire \Tile_X8Y2_E6BEG[0] ;
 wire \Tile_X8Y2_E6BEG[10] ;
 wire \Tile_X8Y2_E6BEG[11] ;
 wire \Tile_X8Y2_E6BEG[1] ;
 wire \Tile_X8Y2_E6BEG[2] ;
 wire \Tile_X8Y2_E6BEG[3] ;
 wire \Tile_X8Y2_E6BEG[4] ;
 wire \Tile_X8Y2_E6BEG[5] ;
 wire \Tile_X8Y2_E6BEG[6] ;
 wire \Tile_X8Y2_E6BEG[7] ;
 wire \Tile_X8Y2_E6BEG[8] ;
 wire \Tile_X8Y2_E6BEG[9] ;
 wire \Tile_X8Y2_EE4BEG[0] ;
 wire \Tile_X8Y2_EE4BEG[10] ;
 wire \Tile_X8Y2_EE4BEG[11] ;
 wire \Tile_X8Y2_EE4BEG[12] ;
 wire \Tile_X8Y2_EE4BEG[13] ;
 wire \Tile_X8Y2_EE4BEG[14] ;
 wire \Tile_X8Y2_EE4BEG[15] ;
 wire \Tile_X8Y2_EE4BEG[1] ;
 wire \Tile_X8Y2_EE4BEG[2] ;
 wire \Tile_X8Y2_EE4BEG[3] ;
 wire \Tile_X8Y2_EE4BEG[4] ;
 wire \Tile_X8Y2_EE4BEG[5] ;
 wire \Tile_X8Y2_EE4BEG[6] ;
 wire \Tile_X8Y2_EE4BEG[7] ;
 wire \Tile_X8Y2_EE4BEG[8] ;
 wire \Tile_X8Y2_EE4BEG[9] ;
 wire \Tile_X8Y2_FrameData_O[0] ;
 wire \Tile_X8Y2_FrameData_O[10] ;
 wire \Tile_X8Y2_FrameData_O[11] ;
 wire \Tile_X8Y2_FrameData_O[12] ;
 wire \Tile_X8Y2_FrameData_O[13] ;
 wire \Tile_X8Y2_FrameData_O[14] ;
 wire \Tile_X8Y2_FrameData_O[15] ;
 wire \Tile_X8Y2_FrameData_O[16] ;
 wire \Tile_X8Y2_FrameData_O[17] ;
 wire \Tile_X8Y2_FrameData_O[18] ;
 wire \Tile_X8Y2_FrameData_O[19] ;
 wire \Tile_X8Y2_FrameData_O[1] ;
 wire \Tile_X8Y2_FrameData_O[20] ;
 wire \Tile_X8Y2_FrameData_O[21] ;
 wire \Tile_X8Y2_FrameData_O[22] ;
 wire \Tile_X8Y2_FrameData_O[23] ;
 wire \Tile_X8Y2_FrameData_O[24] ;
 wire \Tile_X8Y2_FrameData_O[25] ;
 wire \Tile_X8Y2_FrameData_O[26] ;
 wire \Tile_X8Y2_FrameData_O[27] ;
 wire \Tile_X8Y2_FrameData_O[28] ;
 wire \Tile_X8Y2_FrameData_O[29] ;
 wire \Tile_X8Y2_FrameData_O[2] ;
 wire \Tile_X8Y2_FrameData_O[30] ;
 wire \Tile_X8Y2_FrameData_O[31] ;
 wire \Tile_X8Y2_FrameData_O[3] ;
 wire \Tile_X8Y2_FrameData_O[4] ;
 wire \Tile_X8Y2_FrameData_O[5] ;
 wire \Tile_X8Y2_FrameData_O[6] ;
 wire \Tile_X8Y2_FrameData_O[7] ;
 wire \Tile_X8Y2_FrameData_O[8] ;
 wire \Tile_X8Y2_FrameData_O[9] ;
 wire \Tile_X8Y2_FrameStrobe_O[0] ;
 wire \Tile_X8Y2_FrameStrobe_O[10] ;
 wire \Tile_X8Y2_FrameStrobe_O[11] ;
 wire \Tile_X8Y2_FrameStrobe_O[12] ;
 wire \Tile_X8Y2_FrameStrobe_O[13] ;
 wire \Tile_X8Y2_FrameStrobe_O[14] ;
 wire \Tile_X8Y2_FrameStrobe_O[15] ;
 wire \Tile_X8Y2_FrameStrobe_O[16] ;
 wire \Tile_X8Y2_FrameStrobe_O[17] ;
 wire \Tile_X8Y2_FrameStrobe_O[18] ;
 wire \Tile_X8Y2_FrameStrobe_O[19] ;
 wire \Tile_X8Y2_FrameStrobe_O[1] ;
 wire \Tile_X8Y2_FrameStrobe_O[2] ;
 wire \Tile_X8Y2_FrameStrobe_O[3] ;
 wire \Tile_X8Y2_FrameStrobe_O[4] ;
 wire \Tile_X8Y2_FrameStrobe_O[5] ;
 wire \Tile_X8Y2_FrameStrobe_O[6] ;
 wire \Tile_X8Y2_FrameStrobe_O[7] ;
 wire \Tile_X8Y2_FrameStrobe_O[8] ;
 wire \Tile_X8Y2_FrameStrobe_O[9] ;
 wire \Tile_X8Y2_N1BEG[0] ;
 wire \Tile_X8Y2_N1BEG[1] ;
 wire \Tile_X8Y2_N1BEG[2] ;
 wire \Tile_X8Y2_N1BEG[3] ;
 wire \Tile_X8Y2_N2BEG[0] ;
 wire \Tile_X8Y2_N2BEG[1] ;
 wire \Tile_X8Y2_N2BEG[2] ;
 wire \Tile_X8Y2_N2BEG[3] ;
 wire \Tile_X8Y2_N2BEG[4] ;
 wire \Tile_X8Y2_N2BEG[5] ;
 wire \Tile_X8Y2_N2BEG[6] ;
 wire \Tile_X8Y2_N2BEG[7] ;
 wire \Tile_X8Y2_N2BEGb[0] ;
 wire \Tile_X8Y2_N2BEGb[1] ;
 wire \Tile_X8Y2_N2BEGb[2] ;
 wire \Tile_X8Y2_N2BEGb[3] ;
 wire \Tile_X8Y2_N2BEGb[4] ;
 wire \Tile_X8Y2_N2BEGb[5] ;
 wire \Tile_X8Y2_N2BEGb[6] ;
 wire \Tile_X8Y2_N2BEGb[7] ;
 wire \Tile_X8Y2_N4BEG[0] ;
 wire \Tile_X8Y2_N4BEG[10] ;
 wire \Tile_X8Y2_N4BEG[11] ;
 wire \Tile_X8Y2_N4BEG[12] ;
 wire \Tile_X8Y2_N4BEG[13] ;
 wire \Tile_X8Y2_N4BEG[14] ;
 wire \Tile_X8Y2_N4BEG[15] ;
 wire \Tile_X8Y2_N4BEG[1] ;
 wire \Tile_X8Y2_N4BEG[2] ;
 wire \Tile_X8Y2_N4BEG[3] ;
 wire \Tile_X8Y2_N4BEG[4] ;
 wire \Tile_X8Y2_N4BEG[5] ;
 wire \Tile_X8Y2_N4BEG[6] ;
 wire \Tile_X8Y2_N4BEG[7] ;
 wire \Tile_X8Y2_N4BEG[8] ;
 wire \Tile_X8Y2_N4BEG[9] ;
 wire \Tile_X8Y2_NN4BEG[0] ;
 wire \Tile_X8Y2_NN4BEG[10] ;
 wire \Tile_X8Y2_NN4BEG[11] ;
 wire \Tile_X8Y2_NN4BEG[12] ;
 wire \Tile_X8Y2_NN4BEG[13] ;
 wire \Tile_X8Y2_NN4BEG[14] ;
 wire \Tile_X8Y2_NN4BEG[15] ;
 wire \Tile_X8Y2_NN4BEG[1] ;
 wire \Tile_X8Y2_NN4BEG[2] ;
 wire \Tile_X8Y2_NN4BEG[3] ;
 wire \Tile_X8Y2_NN4BEG[4] ;
 wire \Tile_X8Y2_NN4BEG[5] ;
 wire \Tile_X8Y2_NN4BEG[6] ;
 wire \Tile_X8Y2_NN4BEG[7] ;
 wire \Tile_X8Y2_NN4BEG[8] ;
 wire \Tile_X8Y2_NN4BEG[9] ;
 wire \Tile_X8Y2_S1BEG[0] ;
 wire \Tile_X8Y2_S1BEG[1] ;
 wire \Tile_X8Y2_S1BEG[2] ;
 wire \Tile_X8Y2_S1BEG[3] ;
 wire \Tile_X8Y2_S2BEG[0] ;
 wire \Tile_X8Y2_S2BEG[1] ;
 wire \Tile_X8Y2_S2BEG[2] ;
 wire \Tile_X8Y2_S2BEG[3] ;
 wire \Tile_X8Y2_S2BEG[4] ;
 wire \Tile_X8Y2_S2BEG[5] ;
 wire \Tile_X8Y2_S2BEG[6] ;
 wire \Tile_X8Y2_S2BEG[7] ;
 wire \Tile_X8Y2_S2BEGb[0] ;
 wire \Tile_X8Y2_S2BEGb[1] ;
 wire \Tile_X8Y2_S2BEGb[2] ;
 wire \Tile_X8Y2_S2BEGb[3] ;
 wire \Tile_X8Y2_S2BEGb[4] ;
 wire \Tile_X8Y2_S2BEGb[5] ;
 wire \Tile_X8Y2_S2BEGb[6] ;
 wire \Tile_X8Y2_S2BEGb[7] ;
 wire \Tile_X8Y2_S4BEG[0] ;
 wire \Tile_X8Y2_S4BEG[10] ;
 wire \Tile_X8Y2_S4BEG[11] ;
 wire \Tile_X8Y2_S4BEG[12] ;
 wire \Tile_X8Y2_S4BEG[13] ;
 wire \Tile_X8Y2_S4BEG[14] ;
 wire \Tile_X8Y2_S4BEG[15] ;
 wire \Tile_X8Y2_S4BEG[1] ;
 wire \Tile_X8Y2_S4BEG[2] ;
 wire \Tile_X8Y2_S4BEG[3] ;
 wire \Tile_X8Y2_S4BEG[4] ;
 wire \Tile_X8Y2_S4BEG[5] ;
 wire \Tile_X8Y2_S4BEG[6] ;
 wire \Tile_X8Y2_S4BEG[7] ;
 wire \Tile_X8Y2_S4BEG[8] ;
 wire \Tile_X8Y2_S4BEG[9] ;
 wire \Tile_X8Y2_SS4BEG[0] ;
 wire \Tile_X8Y2_SS4BEG[10] ;
 wire \Tile_X8Y2_SS4BEG[11] ;
 wire \Tile_X8Y2_SS4BEG[12] ;
 wire \Tile_X8Y2_SS4BEG[13] ;
 wire \Tile_X8Y2_SS4BEG[14] ;
 wire \Tile_X8Y2_SS4BEG[15] ;
 wire \Tile_X8Y2_SS4BEG[1] ;
 wire \Tile_X8Y2_SS4BEG[2] ;
 wire \Tile_X8Y2_SS4BEG[3] ;
 wire \Tile_X8Y2_SS4BEG[4] ;
 wire \Tile_X8Y2_SS4BEG[5] ;
 wire \Tile_X8Y2_SS4BEG[6] ;
 wire \Tile_X8Y2_SS4BEG[7] ;
 wire \Tile_X8Y2_SS4BEG[8] ;
 wire \Tile_X8Y2_SS4BEG[9] ;
 wire Tile_X8Y2_UserCLKo;
 wire \Tile_X8Y2_W1BEG[0] ;
 wire \Tile_X8Y2_W1BEG[1] ;
 wire \Tile_X8Y2_W1BEG[2] ;
 wire \Tile_X8Y2_W1BEG[3] ;
 wire \Tile_X8Y2_W2BEG[0] ;
 wire \Tile_X8Y2_W2BEG[1] ;
 wire \Tile_X8Y2_W2BEG[2] ;
 wire \Tile_X8Y2_W2BEG[3] ;
 wire \Tile_X8Y2_W2BEG[4] ;
 wire \Tile_X8Y2_W2BEG[5] ;
 wire \Tile_X8Y2_W2BEG[6] ;
 wire \Tile_X8Y2_W2BEG[7] ;
 wire \Tile_X8Y2_W2BEGb[0] ;
 wire \Tile_X8Y2_W2BEGb[1] ;
 wire \Tile_X8Y2_W2BEGb[2] ;
 wire \Tile_X8Y2_W2BEGb[3] ;
 wire \Tile_X8Y2_W2BEGb[4] ;
 wire \Tile_X8Y2_W2BEGb[5] ;
 wire \Tile_X8Y2_W2BEGb[6] ;
 wire \Tile_X8Y2_W2BEGb[7] ;
 wire \Tile_X8Y2_W6BEG[0] ;
 wire \Tile_X8Y2_W6BEG[10] ;
 wire \Tile_X8Y2_W6BEG[11] ;
 wire \Tile_X8Y2_W6BEG[1] ;
 wire \Tile_X8Y2_W6BEG[2] ;
 wire \Tile_X8Y2_W6BEG[3] ;
 wire \Tile_X8Y2_W6BEG[4] ;
 wire \Tile_X8Y2_W6BEG[5] ;
 wire \Tile_X8Y2_W6BEG[6] ;
 wire \Tile_X8Y2_W6BEG[7] ;
 wire \Tile_X8Y2_W6BEG[8] ;
 wire \Tile_X8Y2_W6BEG[9] ;
 wire \Tile_X8Y2_WW4BEG[0] ;
 wire \Tile_X8Y2_WW4BEG[10] ;
 wire \Tile_X8Y2_WW4BEG[11] ;
 wire \Tile_X8Y2_WW4BEG[12] ;
 wire \Tile_X8Y2_WW4BEG[13] ;
 wire \Tile_X8Y2_WW4BEG[14] ;
 wire \Tile_X8Y2_WW4BEG[15] ;
 wire \Tile_X8Y2_WW4BEG[1] ;
 wire \Tile_X8Y2_WW4BEG[2] ;
 wire \Tile_X8Y2_WW4BEG[3] ;
 wire \Tile_X8Y2_WW4BEG[4] ;
 wire \Tile_X8Y2_WW4BEG[5] ;
 wire \Tile_X8Y2_WW4BEG[6] ;
 wire \Tile_X8Y2_WW4BEG[7] ;
 wire \Tile_X8Y2_WW4BEG[8] ;
 wire \Tile_X8Y2_WW4BEG[9] ;
 wire Tile_X8Y3_Co;
 wire \Tile_X8Y3_E1BEG[0] ;
 wire \Tile_X8Y3_E1BEG[1] ;
 wire \Tile_X8Y3_E1BEG[2] ;
 wire \Tile_X8Y3_E1BEG[3] ;
 wire \Tile_X8Y3_E2BEG[0] ;
 wire \Tile_X8Y3_E2BEG[1] ;
 wire \Tile_X8Y3_E2BEG[2] ;
 wire \Tile_X8Y3_E2BEG[3] ;
 wire \Tile_X8Y3_E2BEG[4] ;
 wire \Tile_X8Y3_E2BEG[5] ;
 wire \Tile_X8Y3_E2BEG[6] ;
 wire \Tile_X8Y3_E2BEG[7] ;
 wire \Tile_X8Y3_E2BEGb[0] ;
 wire \Tile_X8Y3_E2BEGb[1] ;
 wire \Tile_X8Y3_E2BEGb[2] ;
 wire \Tile_X8Y3_E2BEGb[3] ;
 wire \Tile_X8Y3_E2BEGb[4] ;
 wire \Tile_X8Y3_E2BEGb[5] ;
 wire \Tile_X8Y3_E2BEGb[6] ;
 wire \Tile_X8Y3_E2BEGb[7] ;
 wire \Tile_X8Y3_E6BEG[0] ;
 wire \Tile_X8Y3_E6BEG[10] ;
 wire \Tile_X8Y3_E6BEG[11] ;
 wire \Tile_X8Y3_E6BEG[1] ;
 wire \Tile_X8Y3_E6BEG[2] ;
 wire \Tile_X8Y3_E6BEG[3] ;
 wire \Tile_X8Y3_E6BEG[4] ;
 wire \Tile_X8Y3_E6BEG[5] ;
 wire \Tile_X8Y3_E6BEG[6] ;
 wire \Tile_X8Y3_E6BEG[7] ;
 wire \Tile_X8Y3_E6BEG[8] ;
 wire \Tile_X8Y3_E6BEG[9] ;
 wire \Tile_X8Y3_EE4BEG[0] ;
 wire \Tile_X8Y3_EE4BEG[10] ;
 wire \Tile_X8Y3_EE4BEG[11] ;
 wire \Tile_X8Y3_EE4BEG[12] ;
 wire \Tile_X8Y3_EE4BEG[13] ;
 wire \Tile_X8Y3_EE4BEG[14] ;
 wire \Tile_X8Y3_EE4BEG[15] ;
 wire \Tile_X8Y3_EE4BEG[1] ;
 wire \Tile_X8Y3_EE4BEG[2] ;
 wire \Tile_X8Y3_EE4BEG[3] ;
 wire \Tile_X8Y3_EE4BEG[4] ;
 wire \Tile_X8Y3_EE4BEG[5] ;
 wire \Tile_X8Y3_EE4BEG[6] ;
 wire \Tile_X8Y3_EE4BEG[7] ;
 wire \Tile_X8Y3_EE4BEG[8] ;
 wire \Tile_X8Y3_EE4BEG[9] ;
 wire \Tile_X8Y3_FrameData_O[0] ;
 wire \Tile_X8Y3_FrameData_O[10] ;
 wire \Tile_X8Y3_FrameData_O[11] ;
 wire \Tile_X8Y3_FrameData_O[12] ;
 wire \Tile_X8Y3_FrameData_O[13] ;
 wire \Tile_X8Y3_FrameData_O[14] ;
 wire \Tile_X8Y3_FrameData_O[15] ;
 wire \Tile_X8Y3_FrameData_O[16] ;
 wire \Tile_X8Y3_FrameData_O[17] ;
 wire \Tile_X8Y3_FrameData_O[18] ;
 wire \Tile_X8Y3_FrameData_O[19] ;
 wire \Tile_X8Y3_FrameData_O[1] ;
 wire \Tile_X8Y3_FrameData_O[20] ;
 wire \Tile_X8Y3_FrameData_O[21] ;
 wire \Tile_X8Y3_FrameData_O[22] ;
 wire \Tile_X8Y3_FrameData_O[23] ;
 wire \Tile_X8Y3_FrameData_O[24] ;
 wire \Tile_X8Y3_FrameData_O[25] ;
 wire \Tile_X8Y3_FrameData_O[26] ;
 wire \Tile_X8Y3_FrameData_O[27] ;
 wire \Tile_X8Y3_FrameData_O[28] ;
 wire \Tile_X8Y3_FrameData_O[29] ;
 wire \Tile_X8Y3_FrameData_O[2] ;
 wire \Tile_X8Y3_FrameData_O[30] ;
 wire \Tile_X8Y3_FrameData_O[31] ;
 wire \Tile_X8Y3_FrameData_O[3] ;
 wire \Tile_X8Y3_FrameData_O[4] ;
 wire \Tile_X8Y3_FrameData_O[5] ;
 wire \Tile_X8Y3_FrameData_O[6] ;
 wire \Tile_X8Y3_FrameData_O[7] ;
 wire \Tile_X8Y3_FrameData_O[8] ;
 wire \Tile_X8Y3_FrameData_O[9] ;
 wire \Tile_X8Y3_FrameStrobe_O[0] ;
 wire \Tile_X8Y3_FrameStrobe_O[10] ;
 wire \Tile_X8Y3_FrameStrobe_O[11] ;
 wire \Tile_X8Y3_FrameStrobe_O[12] ;
 wire \Tile_X8Y3_FrameStrobe_O[13] ;
 wire \Tile_X8Y3_FrameStrobe_O[14] ;
 wire \Tile_X8Y3_FrameStrobe_O[15] ;
 wire \Tile_X8Y3_FrameStrobe_O[16] ;
 wire \Tile_X8Y3_FrameStrobe_O[17] ;
 wire \Tile_X8Y3_FrameStrobe_O[18] ;
 wire \Tile_X8Y3_FrameStrobe_O[19] ;
 wire \Tile_X8Y3_FrameStrobe_O[1] ;
 wire \Tile_X8Y3_FrameStrobe_O[2] ;
 wire \Tile_X8Y3_FrameStrobe_O[3] ;
 wire \Tile_X8Y3_FrameStrobe_O[4] ;
 wire \Tile_X8Y3_FrameStrobe_O[5] ;
 wire \Tile_X8Y3_FrameStrobe_O[6] ;
 wire \Tile_X8Y3_FrameStrobe_O[7] ;
 wire \Tile_X8Y3_FrameStrobe_O[8] ;
 wire \Tile_X8Y3_FrameStrobe_O[9] ;
 wire \Tile_X8Y3_N1BEG[0] ;
 wire \Tile_X8Y3_N1BEG[1] ;
 wire \Tile_X8Y3_N1BEG[2] ;
 wire \Tile_X8Y3_N1BEG[3] ;
 wire \Tile_X8Y3_N2BEG[0] ;
 wire \Tile_X8Y3_N2BEG[1] ;
 wire \Tile_X8Y3_N2BEG[2] ;
 wire \Tile_X8Y3_N2BEG[3] ;
 wire \Tile_X8Y3_N2BEG[4] ;
 wire \Tile_X8Y3_N2BEG[5] ;
 wire \Tile_X8Y3_N2BEG[6] ;
 wire \Tile_X8Y3_N2BEG[7] ;
 wire \Tile_X8Y3_N2BEGb[0] ;
 wire \Tile_X8Y3_N2BEGb[1] ;
 wire \Tile_X8Y3_N2BEGb[2] ;
 wire \Tile_X8Y3_N2BEGb[3] ;
 wire \Tile_X8Y3_N2BEGb[4] ;
 wire \Tile_X8Y3_N2BEGb[5] ;
 wire \Tile_X8Y3_N2BEGb[6] ;
 wire \Tile_X8Y3_N2BEGb[7] ;
 wire \Tile_X8Y3_N4BEG[0] ;
 wire \Tile_X8Y3_N4BEG[10] ;
 wire \Tile_X8Y3_N4BEG[11] ;
 wire \Tile_X8Y3_N4BEG[12] ;
 wire \Tile_X8Y3_N4BEG[13] ;
 wire \Tile_X8Y3_N4BEG[14] ;
 wire \Tile_X8Y3_N4BEG[15] ;
 wire \Tile_X8Y3_N4BEG[1] ;
 wire \Tile_X8Y3_N4BEG[2] ;
 wire \Tile_X8Y3_N4BEG[3] ;
 wire \Tile_X8Y3_N4BEG[4] ;
 wire \Tile_X8Y3_N4BEG[5] ;
 wire \Tile_X8Y3_N4BEG[6] ;
 wire \Tile_X8Y3_N4BEG[7] ;
 wire \Tile_X8Y3_N4BEG[8] ;
 wire \Tile_X8Y3_N4BEG[9] ;
 wire \Tile_X8Y3_NN4BEG[0] ;
 wire \Tile_X8Y3_NN4BEG[10] ;
 wire \Tile_X8Y3_NN4BEG[11] ;
 wire \Tile_X8Y3_NN4BEG[12] ;
 wire \Tile_X8Y3_NN4BEG[13] ;
 wire \Tile_X8Y3_NN4BEG[14] ;
 wire \Tile_X8Y3_NN4BEG[15] ;
 wire \Tile_X8Y3_NN4BEG[1] ;
 wire \Tile_X8Y3_NN4BEG[2] ;
 wire \Tile_X8Y3_NN4BEG[3] ;
 wire \Tile_X8Y3_NN4BEG[4] ;
 wire \Tile_X8Y3_NN4BEG[5] ;
 wire \Tile_X8Y3_NN4BEG[6] ;
 wire \Tile_X8Y3_NN4BEG[7] ;
 wire \Tile_X8Y3_NN4BEG[8] ;
 wire \Tile_X8Y3_NN4BEG[9] ;
 wire \Tile_X8Y3_S1BEG[0] ;
 wire \Tile_X8Y3_S1BEG[1] ;
 wire \Tile_X8Y3_S1BEG[2] ;
 wire \Tile_X8Y3_S1BEG[3] ;
 wire \Tile_X8Y3_S2BEG[0] ;
 wire \Tile_X8Y3_S2BEG[1] ;
 wire \Tile_X8Y3_S2BEG[2] ;
 wire \Tile_X8Y3_S2BEG[3] ;
 wire \Tile_X8Y3_S2BEG[4] ;
 wire \Tile_X8Y3_S2BEG[5] ;
 wire \Tile_X8Y3_S2BEG[6] ;
 wire \Tile_X8Y3_S2BEG[7] ;
 wire \Tile_X8Y3_S2BEGb[0] ;
 wire \Tile_X8Y3_S2BEGb[1] ;
 wire \Tile_X8Y3_S2BEGb[2] ;
 wire \Tile_X8Y3_S2BEGb[3] ;
 wire \Tile_X8Y3_S2BEGb[4] ;
 wire \Tile_X8Y3_S2BEGb[5] ;
 wire \Tile_X8Y3_S2BEGb[6] ;
 wire \Tile_X8Y3_S2BEGb[7] ;
 wire \Tile_X8Y3_S4BEG[0] ;
 wire \Tile_X8Y3_S4BEG[10] ;
 wire \Tile_X8Y3_S4BEG[11] ;
 wire \Tile_X8Y3_S4BEG[12] ;
 wire \Tile_X8Y3_S4BEG[13] ;
 wire \Tile_X8Y3_S4BEG[14] ;
 wire \Tile_X8Y3_S4BEG[15] ;
 wire \Tile_X8Y3_S4BEG[1] ;
 wire \Tile_X8Y3_S4BEG[2] ;
 wire \Tile_X8Y3_S4BEG[3] ;
 wire \Tile_X8Y3_S4BEG[4] ;
 wire \Tile_X8Y3_S4BEG[5] ;
 wire \Tile_X8Y3_S4BEG[6] ;
 wire \Tile_X8Y3_S4BEG[7] ;
 wire \Tile_X8Y3_S4BEG[8] ;
 wire \Tile_X8Y3_S4BEG[9] ;
 wire \Tile_X8Y3_SS4BEG[0] ;
 wire \Tile_X8Y3_SS4BEG[10] ;
 wire \Tile_X8Y3_SS4BEG[11] ;
 wire \Tile_X8Y3_SS4BEG[12] ;
 wire \Tile_X8Y3_SS4BEG[13] ;
 wire \Tile_X8Y3_SS4BEG[14] ;
 wire \Tile_X8Y3_SS4BEG[15] ;
 wire \Tile_X8Y3_SS4BEG[1] ;
 wire \Tile_X8Y3_SS4BEG[2] ;
 wire \Tile_X8Y3_SS4BEG[3] ;
 wire \Tile_X8Y3_SS4BEG[4] ;
 wire \Tile_X8Y3_SS4BEG[5] ;
 wire \Tile_X8Y3_SS4BEG[6] ;
 wire \Tile_X8Y3_SS4BEG[7] ;
 wire \Tile_X8Y3_SS4BEG[8] ;
 wire \Tile_X8Y3_SS4BEG[9] ;
 wire Tile_X8Y3_UserCLKo;
 wire \Tile_X8Y3_W1BEG[0] ;
 wire \Tile_X8Y3_W1BEG[1] ;
 wire \Tile_X8Y3_W1BEG[2] ;
 wire \Tile_X8Y3_W1BEG[3] ;
 wire \Tile_X8Y3_W2BEG[0] ;
 wire \Tile_X8Y3_W2BEG[1] ;
 wire \Tile_X8Y3_W2BEG[2] ;
 wire \Tile_X8Y3_W2BEG[3] ;
 wire \Tile_X8Y3_W2BEG[4] ;
 wire \Tile_X8Y3_W2BEG[5] ;
 wire \Tile_X8Y3_W2BEG[6] ;
 wire \Tile_X8Y3_W2BEG[7] ;
 wire \Tile_X8Y3_W2BEGb[0] ;
 wire \Tile_X8Y3_W2BEGb[1] ;
 wire \Tile_X8Y3_W2BEGb[2] ;
 wire \Tile_X8Y3_W2BEGb[3] ;
 wire \Tile_X8Y3_W2BEGb[4] ;
 wire \Tile_X8Y3_W2BEGb[5] ;
 wire \Tile_X8Y3_W2BEGb[6] ;
 wire \Tile_X8Y3_W2BEGb[7] ;
 wire \Tile_X8Y3_W6BEG[0] ;
 wire \Tile_X8Y3_W6BEG[10] ;
 wire \Tile_X8Y3_W6BEG[11] ;
 wire \Tile_X8Y3_W6BEG[1] ;
 wire \Tile_X8Y3_W6BEG[2] ;
 wire \Tile_X8Y3_W6BEG[3] ;
 wire \Tile_X8Y3_W6BEG[4] ;
 wire \Tile_X8Y3_W6BEG[5] ;
 wire \Tile_X8Y3_W6BEG[6] ;
 wire \Tile_X8Y3_W6BEG[7] ;
 wire \Tile_X8Y3_W6BEG[8] ;
 wire \Tile_X8Y3_W6BEG[9] ;
 wire \Tile_X8Y3_WW4BEG[0] ;
 wire \Tile_X8Y3_WW4BEG[10] ;
 wire \Tile_X8Y3_WW4BEG[11] ;
 wire \Tile_X8Y3_WW4BEG[12] ;
 wire \Tile_X8Y3_WW4BEG[13] ;
 wire \Tile_X8Y3_WW4BEG[14] ;
 wire \Tile_X8Y3_WW4BEG[15] ;
 wire \Tile_X8Y3_WW4BEG[1] ;
 wire \Tile_X8Y3_WW4BEG[2] ;
 wire \Tile_X8Y3_WW4BEG[3] ;
 wire \Tile_X8Y3_WW4BEG[4] ;
 wire \Tile_X8Y3_WW4BEG[5] ;
 wire \Tile_X8Y3_WW4BEG[6] ;
 wire \Tile_X8Y3_WW4BEG[7] ;
 wire \Tile_X8Y3_WW4BEG[8] ;
 wire \Tile_X8Y3_WW4BEG[9] ;
 wire Tile_X8Y4_Co;
 wire \Tile_X8Y4_E1BEG[0] ;
 wire \Tile_X8Y4_E1BEG[1] ;
 wire \Tile_X8Y4_E1BEG[2] ;
 wire \Tile_X8Y4_E1BEG[3] ;
 wire \Tile_X8Y4_E2BEG[0] ;
 wire \Tile_X8Y4_E2BEG[1] ;
 wire \Tile_X8Y4_E2BEG[2] ;
 wire \Tile_X8Y4_E2BEG[3] ;
 wire \Tile_X8Y4_E2BEG[4] ;
 wire \Tile_X8Y4_E2BEG[5] ;
 wire \Tile_X8Y4_E2BEG[6] ;
 wire \Tile_X8Y4_E2BEG[7] ;
 wire \Tile_X8Y4_E2BEGb[0] ;
 wire \Tile_X8Y4_E2BEGb[1] ;
 wire \Tile_X8Y4_E2BEGb[2] ;
 wire \Tile_X8Y4_E2BEGb[3] ;
 wire \Tile_X8Y4_E2BEGb[4] ;
 wire \Tile_X8Y4_E2BEGb[5] ;
 wire \Tile_X8Y4_E2BEGb[6] ;
 wire \Tile_X8Y4_E2BEGb[7] ;
 wire \Tile_X8Y4_E6BEG[0] ;
 wire \Tile_X8Y4_E6BEG[10] ;
 wire \Tile_X8Y4_E6BEG[11] ;
 wire \Tile_X8Y4_E6BEG[1] ;
 wire \Tile_X8Y4_E6BEG[2] ;
 wire \Tile_X8Y4_E6BEG[3] ;
 wire \Tile_X8Y4_E6BEG[4] ;
 wire \Tile_X8Y4_E6BEG[5] ;
 wire \Tile_X8Y4_E6BEG[6] ;
 wire \Tile_X8Y4_E6BEG[7] ;
 wire \Tile_X8Y4_E6BEG[8] ;
 wire \Tile_X8Y4_E6BEG[9] ;
 wire \Tile_X8Y4_EE4BEG[0] ;
 wire \Tile_X8Y4_EE4BEG[10] ;
 wire \Tile_X8Y4_EE4BEG[11] ;
 wire \Tile_X8Y4_EE4BEG[12] ;
 wire \Tile_X8Y4_EE4BEG[13] ;
 wire \Tile_X8Y4_EE4BEG[14] ;
 wire \Tile_X8Y4_EE4BEG[15] ;
 wire \Tile_X8Y4_EE4BEG[1] ;
 wire \Tile_X8Y4_EE4BEG[2] ;
 wire \Tile_X8Y4_EE4BEG[3] ;
 wire \Tile_X8Y4_EE4BEG[4] ;
 wire \Tile_X8Y4_EE4BEG[5] ;
 wire \Tile_X8Y4_EE4BEG[6] ;
 wire \Tile_X8Y4_EE4BEG[7] ;
 wire \Tile_X8Y4_EE4BEG[8] ;
 wire \Tile_X8Y4_EE4BEG[9] ;
 wire \Tile_X8Y4_FrameData_O[0] ;
 wire \Tile_X8Y4_FrameData_O[10] ;
 wire \Tile_X8Y4_FrameData_O[11] ;
 wire \Tile_X8Y4_FrameData_O[12] ;
 wire \Tile_X8Y4_FrameData_O[13] ;
 wire \Tile_X8Y4_FrameData_O[14] ;
 wire \Tile_X8Y4_FrameData_O[15] ;
 wire \Tile_X8Y4_FrameData_O[16] ;
 wire \Tile_X8Y4_FrameData_O[17] ;
 wire \Tile_X8Y4_FrameData_O[18] ;
 wire \Tile_X8Y4_FrameData_O[19] ;
 wire \Tile_X8Y4_FrameData_O[1] ;
 wire \Tile_X8Y4_FrameData_O[20] ;
 wire \Tile_X8Y4_FrameData_O[21] ;
 wire \Tile_X8Y4_FrameData_O[22] ;
 wire \Tile_X8Y4_FrameData_O[23] ;
 wire \Tile_X8Y4_FrameData_O[24] ;
 wire \Tile_X8Y4_FrameData_O[25] ;
 wire \Tile_X8Y4_FrameData_O[26] ;
 wire \Tile_X8Y4_FrameData_O[27] ;
 wire \Tile_X8Y4_FrameData_O[28] ;
 wire \Tile_X8Y4_FrameData_O[29] ;
 wire \Tile_X8Y4_FrameData_O[2] ;
 wire \Tile_X8Y4_FrameData_O[30] ;
 wire \Tile_X8Y4_FrameData_O[31] ;
 wire \Tile_X8Y4_FrameData_O[3] ;
 wire \Tile_X8Y4_FrameData_O[4] ;
 wire \Tile_X8Y4_FrameData_O[5] ;
 wire \Tile_X8Y4_FrameData_O[6] ;
 wire \Tile_X8Y4_FrameData_O[7] ;
 wire \Tile_X8Y4_FrameData_O[8] ;
 wire \Tile_X8Y4_FrameData_O[9] ;
 wire \Tile_X8Y4_FrameStrobe_O[0] ;
 wire \Tile_X8Y4_FrameStrobe_O[10] ;
 wire \Tile_X8Y4_FrameStrobe_O[11] ;
 wire \Tile_X8Y4_FrameStrobe_O[12] ;
 wire \Tile_X8Y4_FrameStrobe_O[13] ;
 wire \Tile_X8Y4_FrameStrobe_O[14] ;
 wire \Tile_X8Y4_FrameStrobe_O[15] ;
 wire \Tile_X8Y4_FrameStrobe_O[16] ;
 wire \Tile_X8Y4_FrameStrobe_O[17] ;
 wire \Tile_X8Y4_FrameStrobe_O[18] ;
 wire \Tile_X8Y4_FrameStrobe_O[19] ;
 wire \Tile_X8Y4_FrameStrobe_O[1] ;
 wire \Tile_X8Y4_FrameStrobe_O[2] ;
 wire \Tile_X8Y4_FrameStrobe_O[3] ;
 wire \Tile_X8Y4_FrameStrobe_O[4] ;
 wire \Tile_X8Y4_FrameStrobe_O[5] ;
 wire \Tile_X8Y4_FrameStrobe_O[6] ;
 wire \Tile_X8Y4_FrameStrobe_O[7] ;
 wire \Tile_X8Y4_FrameStrobe_O[8] ;
 wire \Tile_X8Y4_FrameStrobe_O[9] ;
 wire \Tile_X8Y4_N1BEG[0] ;
 wire \Tile_X8Y4_N1BEG[1] ;
 wire \Tile_X8Y4_N1BEG[2] ;
 wire \Tile_X8Y4_N1BEG[3] ;
 wire \Tile_X8Y4_N2BEG[0] ;
 wire \Tile_X8Y4_N2BEG[1] ;
 wire \Tile_X8Y4_N2BEG[2] ;
 wire \Tile_X8Y4_N2BEG[3] ;
 wire \Tile_X8Y4_N2BEG[4] ;
 wire \Tile_X8Y4_N2BEG[5] ;
 wire \Tile_X8Y4_N2BEG[6] ;
 wire \Tile_X8Y4_N2BEG[7] ;
 wire \Tile_X8Y4_N2BEGb[0] ;
 wire \Tile_X8Y4_N2BEGb[1] ;
 wire \Tile_X8Y4_N2BEGb[2] ;
 wire \Tile_X8Y4_N2BEGb[3] ;
 wire \Tile_X8Y4_N2BEGb[4] ;
 wire \Tile_X8Y4_N2BEGb[5] ;
 wire \Tile_X8Y4_N2BEGb[6] ;
 wire \Tile_X8Y4_N2BEGb[7] ;
 wire \Tile_X8Y4_N4BEG[0] ;
 wire \Tile_X8Y4_N4BEG[10] ;
 wire \Tile_X8Y4_N4BEG[11] ;
 wire \Tile_X8Y4_N4BEG[12] ;
 wire \Tile_X8Y4_N4BEG[13] ;
 wire \Tile_X8Y4_N4BEG[14] ;
 wire \Tile_X8Y4_N4BEG[15] ;
 wire \Tile_X8Y4_N4BEG[1] ;
 wire \Tile_X8Y4_N4BEG[2] ;
 wire \Tile_X8Y4_N4BEG[3] ;
 wire \Tile_X8Y4_N4BEG[4] ;
 wire \Tile_X8Y4_N4BEG[5] ;
 wire \Tile_X8Y4_N4BEG[6] ;
 wire \Tile_X8Y4_N4BEG[7] ;
 wire \Tile_X8Y4_N4BEG[8] ;
 wire \Tile_X8Y4_N4BEG[9] ;
 wire \Tile_X8Y4_NN4BEG[0] ;
 wire \Tile_X8Y4_NN4BEG[10] ;
 wire \Tile_X8Y4_NN4BEG[11] ;
 wire \Tile_X8Y4_NN4BEG[12] ;
 wire \Tile_X8Y4_NN4BEG[13] ;
 wire \Tile_X8Y4_NN4BEG[14] ;
 wire \Tile_X8Y4_NN4BEG[15] ;
 wire \Tile_X8Y4_NN4BEG[1] ;
 wire \Tile_X8Y4_NN4BEG[2] ;
 wire \Tile_X8Y4_NN4BEG[3] ;
 wire \Tile_X8Y4_NN4BEG[4] ;
 wire \Tile_X8Y4_NN4BEG[5] ;
 wire \Tile_X8Y4_NN4BEG[6] ;
 wire \Tile_X8Y4_NN4BEG[7] ;
 wire \Tile_X8Y4_NN4BEG[8] ;
 wire \Tile_X8Y4_NN4BEG[9] ;
 wire \Tile_X8Y4_S1BEG[0] ;
 wire \Tile_X8Y4_S1BEG[1] ;
 wire \Tile_X8Y4_S1BEG[2] ;
 wire \Tile_X8Y4_S1BEG[3] ;
 wire \Tile_X8Y4_S2BEG[0] ;
 wire \Tile_X8Y4_S2BEG[1] ;
 wire \Tile_X8Y4_S2BEG[2] ;
 wire \Tile_X8Y4_S2BEG[3] ;
 wire \Tile_X8Y4_S2BEG[4] ;
 wire \Tile_X8Y4_S2BEG[5] ;
 wire \Tile_X8Y4_S2BEG[6] ;
 wire \Tile_X8Y4_S2BEG[7] ;
 wire \Tile_X8Y4_S2BEGb[0] ;
 wire \Tile_X8Y4_S2BEGb[1] ;
 wire \Tile_X8Y4_S2BEGb[2] ;
 wire \Tile_X8Y4_S2BEGb[3] ;
 wire \Tile_X8Y4_S2BEGb[4] ;
 wire \Tile_X8Y4_S2BEGb[5] ;
 wire \Tile_X8Y4_S2BEGb[6] ;
 wire \Tile_X8Y4_S2BEGb[7] ;
 wire \Tile_X8Y4_S4BEG[0] ;
 wire \Tile_X8Y4_S4BEG[10] ;
 wire \Tile_X8Y4_S4BEG[11] ;
 wire \Tile_X8Y4_S4BEG[12] ;
 wire \Tile_X8Y4_S4BEG[13] ;
 wire \Tile_X8Y4_S4BEG[14] ;
 wire \Tile_X8Y4_S4BEG[15] ;
 wire \Tile_X8Y4_S4BEG[1] ;
 wire \Tile_X8Y4_S4BEG[2] ;
 wire \Tile_X8Y4_S4BEG[3] ;
 wire \Tile_X8Y4_S4BEG[4] ;
 wire \Tile_X8Y4_S4BEG[5] ;
 wire \Tile_X8Y4_S4BEG[6] ;
 wire \Tile_X8Y4_S4BEG[7] ;
 wire \Tile_X8Y4_S4BEG[8] ;
 wire \Tile_X8Y4_S4BEG[9] ;
 wire \Tile_X8Y4_SS4BEG[0] ;
 wire \Tile_X8Y4_SS4BEG[10] ;
 wire \Tile_X8Y4_SS4BEG[11] ;
 wire \Tile_X8Y4_SS4BEG[12] ;
 wire \Tile_X8Y4_SS4BEG[13] ;
 wire \Tile_X8Y4_SS4BEG[14] ;
 wire \Tile_X8Y4_SS4BEG[15] ;
 wire \Tile_X8Y4_SS4BEG[1] ;
 wire \Tile_X8Y4_SS4BEG[2] ;
 wire \Tile_X8Y4_SS4BEG[3] ;
 wire \Tile_X8Y4_SS4BEG[4] ;
 wire \Tile_X8Y4_SS4BEG[5] ;
 wire \Tile_X8Y4_SS4BEG[6] ;
 wire \Tile_X8Y4_SS4BEG[7] ;
 wire \Tile_X8Y4_SS4BEG[8] ;
 wire \Tile_X8Y4_SS4BEG[9] ;
 wire Tile_X8Y4_UserCLKo;
 wire \Tile_X8Y4_W1BEG[0] ;
 wire \Tile_X8Y4_W1BEG[1] ;
 wire \Tile_X8Y4_W1BEG[2] ;
 wire \Tile_X8Y4_W1BEG[3] ;
 wire \Tile_X8Y4_W2BEG[0] ;
 wire \Tile_X8Y4_W2BEG[1] ;
 wire \Tile_X8Y4_W2BEG[2] ;
 wire \Tile_X8Y4_W2BEG[3] ;
 wire \Tile_X8Y4_W2BEG[4] ;
 wire \Tile_X8Y4_W2BEG[5] ;
 wire \Tile_X8Y4_W2BEG[6] ;
 wire \Tile_X8Y4_W2BEG[7] ;
 wire \Tile_X8Y4_W2BEGb[0] ;
 wire \Tile_X8Y4_W2BEGb[1] ;
 wire \Tile_X8Y4_W2BEGb[2] ;
 wire \Tile_X8Y4_W2BEGb[3] ;
 wire \Tile_X8Y4_W2BEGb[4] ;
 wire \Tile_X8Y4_W2BEGb[5] ;
 wire \Tile_X8Y4_W2BEGb[6] ;
 wire \Tile_X8Y4_W2BEGb[7] ;
 wire \Tile_X8Y4_W6BEG[0] ;
 wire \Tile_X8Y4_W6BEG[10] ;
 wire \Tile_X8Y4_W6BEG[11] ;
 wire \Tile_X8Y4_W6BEG[1] ;
 wire \Tile_X8Y4_W6BEG[2] ;
 wire \Tile_X8Y4_W6BEG[3] ;
 wire \Tile_X8Y4_W6BEG[4] ;
 wire \Tile_X8Y4_W6BEG[5] ;
 wire \Tile_X8Y4_W6BEG[6] ;
 wire \Tile_X8Y4_W6BEG[7] ;
 wire \Tile_X8Y4_W6BEG[8] ;
 wire \Tile_X8Y4_W6BEG[9] ;
 wire \Tile_X8Y4_WW4BEG[0] ;
 wire \Tile_X8Y4_WW4BEG[10] ;
 wire \Tile_X8Y4_WW4BEG[11] ;
 wire \Tile_X8Y4_WW4BEG[12] ;
 wire \Tile_X8Y4_WW4BEG[13] ;
 wire \Tile_X8Y4_WW4BEG[14] ;
 wire \Tile_X8Y4_WW4BEG[15] ;
 wire \Tile_X8Y4_WW4BEG[1] ;
 wire \Tile_X8Y4_WW4BEG[2] ;
 wire \Tile_X8Y4_WW4BEG[3] ;
 wire \Tile_X8Y4_WW4BEG[4] ;
 wire \Tile_X8Y4_WW4BEG[5] ;
 wire \Tile_X8Y4_WW4BEG[6] ;
 wire \Tile_X8Y4_WW4BEG[7] ;
 wire \Tile_X8Y4_WW4BEG[8] ;
 wire \Tile_X8Y4_WW4BEG[9] ;
 wire Tile_X8Y5_Co;
 wire \Tile_X8Y5_E1BEG[0] ;
 wire \Tile_X8Y5_E1BEG[1] ;
 wire \Tile_X8Y5_E1BEG[2] ;
 wire \Tile_X8Y5_E1BEG[3] ;
 wire \Tile_X8Y5_E2BEG[0] ;
 wire \Tile_X8Y5_E2BEG[1] ;
 wire \Tile_X8Y5_E2BEG[2] ;
 wire \Tile_X8Y5_E2BEG[3] ;
 wire \Tile_X8Y5_E2BEG[4] ;
 wire \Tile_X8Y5_E2BEG[5] ;
 wire \Tile_X8Y5_E2BEG[6] ;
 wire \Tile_X8Y5_E2BEG[7] ;
 wire \Tile_X8Y5_E2BEGb[0] ;
 wire \Tile_X8Y5_E2BEGb[1] ;
 wire \Tile_X8Y5_E2BEGb[2] ;
 wire \Tile_X8Y5_E2BEGb[3] ;
 wire \Tile_X8Y5_E2BEGb[4] ;
 wire \Tile_X8Y5_E2BEGb[5] ;
 wire \Tile_X8Y5_E2BEGb[6] ;
 wire \Tile_X8Y5_E2BEGb[7] ;
 wire \Tile_X8Y5_E6BEG[0] ;
 wire \Tile_X8Y5_E6BEG[10] ;
 wire \Tile_X8Y5_E6BEG[11] ;
 wire \Tile_X8Y5_E6BEG[1] ;
 wire \Tile_X8Y5_E6BEG[2] ;
 wire \Tile_X8Y5_E6BEG[3] ;
 wire \Tile_X8Y5_E6BEG[4] ;
 wire \Tile_X8Y5_E6BEG[5] ;
 wire \Tile_X8Y5_E6BEG[6] ;
 wire \Tile_X8Y5_E6BEG[7] ;
 wire \Tile_X8Y5_E6BEG[8] ;
 wire \Tile_X8Y5_E6BEG[9] ;
 wire \Tile_X8Y5_EE4BEG[0] ;
 wire \Tile_X8Y5_EE4BEG[10] ;
 wire \Tile_X8Y5_EE4BEG[11] ;
 wire \Tile_X8Y5_EE4BEG[12] ;
 wire \Tile_X8Y5_EE4BEG[13] ;
 wire \Tile_X8Y5_EE4BEG[14] ;
 wire \Tile_X8Y5_EE4BEG[15] ;
 wire \Tile_X8Y5_EE4BEG[1] ;
 wire \Tile_X8Y5_EE4BEG[2] ;
 wire \Tile_X8Y5_EE4BEG[3] ;
 wire \Tile_X8Y5_EE4BEG[4] ;
 wire \Tile_X8Y5_EE4BEG[5] ;
 wire \Tile_X8Y5_EE4BEG[6] ;
 wire \Tile_X8Y5_EE4BEG[7] ;
 wire \Tile_X8Y5_EE4BEG[8] ;
 wire \Tile_X8Y5_EE4BEG[9] ;
 wire \Tile_X8Y5_FrameData_O[0] ;
 wire \Tile_X8Y5_FrameData_O[10] ;
 wire \Tile_X8Y5_FrameData_O[11] ;
 wire \Tile_X8Y5_FrameData_O[12] ;
 wire \Tile_X8Y5_FrameData_O[13] ;
 wire \Tile_X8Y5_FrameData_O[14] ;
 wire \Tile_X8Y5_FrameData_O[15] ;
 wire \Tile_X8Y5_FrameData_O[16] ;
 wire \Tile_X8Y5_FrameData_O[17] ;
 wire \Tile_X8Y5_FrameData_O[18] ;
 wire \Tile_X8Y5_FrameData_O[19] ;
 wire \Tile_X8Y5_FrameData_O[1] ;
 wire \Tile_X8Y5_FrameData_O[20] ;
 wire \Tile_X8Y5_FrameData_O[21] ;
 wire \Tile_X8Y5_FrameData_O[22] ;
 wire \Tile_X8Y5_FrameData_O[23] ;
 wire \Tile_X8Y5_FrameData_O[24] ;
 wire \Tile_X8Y5_FrameData_O[25] ;
 wire \Tile_X8Y5_FrameData_O[26] ;
 wire \Tile_X8Y5_FrameData_O[27] ;
 wire \Tile_X8Y5_FrameData_O[28] ;
 wire \Tile_X8Y5_FrameData_O[29] ;
 wire \Tile_X8Y5_FrameData_O[2] ;
 wire \Tile_X8Y5_FrameData_O[30] ;
 wire \Tile_X8Y5_FrameData_O[31] ;
 wire \Tile_X8Y5_FrameData_O[3] ;
 wire \Tile_X8Y5_FrameData_O[4] ;
 wire \Tile_X8Y5_FrameData_O[5] ;
 wire \Tile_X8Y5_FrameData_O[6] ;
 wire \Tile_X8Y5_FrameData_O[7] ;
 wire \Tile_X8Y5_FrameData_O[8] ;
 wire \Tile_X8Y5_FrameData_O[9] ;
 wire \Tile_X8Y5_FrameStrobe_O[0] ;
 wire \Tile_X8Y5_FrameStrobe_O[10] ;
 wire \Tile_X8Y5_FrameStrobe_O[11] ;
 wire \Tile_X8Y5_FrameStrobe_O[12] ;
 wire \Tile_X8Y5_FrameStrobe_O[13] ;
 wire \Tile_X8Y5_FrameStrobe_O[14] ;
 wire \Tile_X8Y5_FrameStrobe_O[15] ;
 wire \Tile_X8Y5_FrameStrobe_O[16] ;
 wire \Tile_X8Y5_FrameStrobe_O[17] ;
 wire \Tile_X8Y5_FrameStrobe_O[18] ;
 wire \Tile_X8Y5_FrameStrobe_O[19] ;
 wire \Tile_X8Y5_FrameStrobe_O[1] ;
 wire \Tile_X8Y5_FrameStrobe_O[2] ;
 wire \Tile_X8Y5_FrameStrobe_O[3] ;
 wire \Tile_X8Y5_FrameStrobe_O[4] ;
 wire \Tile_X8Y5_FrameStrobe_O[5] ;
 wire \Tile_X8Y5_FrameStrobe_O[6] ;
 wire \Tile_X8Y5_FrameStrobe_O[7] ;
 wire \Tile_X8Y5_FrameStrobe_O[8] ;
 wire \Tile_X8Y5_FrameStrobe_O[9] ;
 wire \Tile_X8Y5_N1BEG[0] ;
 wire \Tile_X8Y5_N1BEG[1] ;
 wire \Tile_X8Y5_N1BEG[2] ;
 wire \Tile_X8Y5_N1BEG[3] ;
 wire \Tile_X8Y5_N2BEG[0] ;
 wire \Tile_X8Y5_N2BEG[1] ;
 wire \Tile_X8Y5_N2BEG[2] ;
 wire \Tile_X8Y5_N2BEG[3] ;
 wire \Tile_X8Y5_N2BEG[4] ;
 wire \Tile_X8Y5_N2BEG[5] ;
 wire \Tile_X8Y5_N2BEG[6] ;
 wire \Tile_X8Y5_N2BEG[7] ;
 wire \Tile_X8Y5_N2BEGb[0] ;
 wire \Tile_X8Y5_N2BEGb[1] ;
 wire \Tile_X8Y5_N2BEGb[2] ;
 wire \Tile_X8Y5_N2BEGb[3] ;
 wire \Tile_X8Y5_N2BEGb[4] ;
 wire \Tile_X8Y5_N2BEGb[5] ;
 wire \Tile_X8Y5_N2BEGb[6] ;
 wire \Tile_X8Y5_N2BEGb[7] ;
 wire \Tile_X8Y5_N4BEG[0] ;
 wire \Tile_X8Y5_N4BEG[10] ;
 wire \Tile_X8Y5_N4BEG[11] ;
 wire \Tile_X8Y5_N4BEG[12] ;
 wire \Tile_X8Y5_N4BEG[13] ;
 wire \Tile_X8Y5_N4BEG[14] ;
 wire \Tile_X8Y5_N4BEG[15] ;
 wire \Tile_X8Y5_N4BEG[1] ;
 wire \Tile_X8Y5_N4BEG[2] ;
 wire \Tile_X8Y5_N4BEG[3] ;
 wire \Tile_X8Y5_N4BEG[4] ;
 wire \Tile_X8Y5_N4BEG[5] ;
 wire \Tile_X8Y5_N4BEG[6] ;
 wire \Tile_X8Y5_N4BEG[7] ;
 wire \Tile_X8Y5_N4BEG[8] ;
 wire \Tile_X8Y5_N4BEG[9] ;
 wire \Tile_X8Y5_NN4BEG[0] ;
 wire \Tile_X8Y5_NN4BEG[10] ;
 wire \Tile_X8Y5_NN4BEG[11] ;
 wire \Tile_X8Y5_NN4BEG[12] ;
 wire \Tile_X8Y5_NN4BEG[13] ;
 wire \Tile_X8Y5_NN4BEG[14] ;
 wire \Tile_X8Y5_NN4BEG[15] ;
 wire \Tile_X8Y5_NN4BEG[1] ;
 wire \Tile_X8Y5_NN4BEG[2] ;
 wire \Tile_X8Y5_NN4BEG[3] ;
 wire \Tile_X8Y5_NN4BEG[4] ;
 wire \Tile_X8Y5_NN4BEG[5] ;
 wire \Tile_X8Y5_NN4BEG[6] ;
 wire \Tile_X8Y5_NN4BEG[7] ;
 wire \Tile_X8Y5_NN4BEG[8] ;
 wire \Tile_X8Y5_NN4BEG[9] ;
 wire \Tile_X8Y5_S1BEG[0] ;
 wire \Tile_X8Y5_S1BEG[1] ;
 wire \Tile_X8Y5_S1BEG[2] ;
 wire \Tile_X8Y5_S1BEG[3] ;
 wire \Tile_X8Y5_S2BEG[0] ;
 wire \Tile_X8Y5_S2BEG[1] ;
 wire \Tile_X8Y5_S2BEG[2] ;
 wire \Tile_X8Y5_S2BEG[3] ;
 wire \Tile_X8Y5_S2BEG[4] ;
 wire \Tile_X8Y5_S2BEG[5] ;
 wire \Tile_X8Y5_S2BEG[6] ;
 wire \Tile_X8Y5_S2BEG[7] ;
 wire \Tile_X8Y5_S2BEGb[0] ;
 wire \Tile_X8Y5_S2BEGb[1] ;
 wire \Tile_X8Y5_S2BEGb[2] ;
 wire \Tile_X8Y5_S2BEGb[3] ;
 wire \Tile_X8Y5_S2BEGb[4] ;
 wire \Tile_X8Y5_S2BEGb[5] ;
 wire \Tile_X8Y5_S2BEGb[6] ;
 wire \Tile_X8Y5_S2BEGb[7] ;
 wire \Tile_X8Y5_S4BEG[0] ;
 wire \Tile_X8Y5_S4BEG[10] ;
 wire \Tile_X8Y5_S4BEG[11] ;
 wire \Tile_X8Y5_S4BEG[12] ;
 wire \Tile_X8Y5_S4BEG[13] ;
 wire \Tile_X8Y5_S4BEG[14] ;
 wire \Tile_X8Y5_S4BEG[15] ;
 wire \Tile_X8Y5_S4BEG[1] ;
 wire \Tile_X8Y5_S4BEG[2] ;
 wire \Tile_X8Y5_S4BEG[3] ;
 wire \Tile_X8Y5_S4BEG[4] ;
 wire \Tile_X8Y5_S4BEG[5] ;
 wire \Tile_X8Y5_S4BEG[6] ;
 wire \Tile_X8Y5_S4BEG[7] ;
 wire \Tile_X8Y5_S4BEG[8] ;
 wire \Tile_X8Y5_S4BEG[9] ;
 wire \Tile_X8Y5_SS4BEG[0] ;
 wire \Tile_X8Y5_SS4BEG[10] ;
 wire \Tile_X8Y5_SS4BEG[11] ;
 wire \Tile_X8Y5_SS4BEG[12] ;
 wire \Tile_X8Y5_SS4BEG[13] ;
 wire \Tile_X8Y5_SS4BEG[14] ;
 wire \Tile_X8Y5_SS4BEG[15] ;
 wire \Tile_X8Y5_SS4BEG[1] ;
 wire \Tile_X8Y5_SS4BEG[2] ;
 wire \Tile_X8Y5_SS4BEG[3] ;
 wire \Tile_X8Y5_SS4BEG[4] ;
 wire \Tile_X8Y5_SS4BEG[5] ;
 wire \Tile_X8Y5_SS4BEG[6] ;
 wire \Tile_X8Y5_SS4BEG[7] ;
 wire \Tile_X8Y5_SS4BEG[8] ;
 wire \Tile_X8Y5_SS4BEG[9] ;
 wire Tile_X8Y5_UserCLKo;
 wire \Tile_X8Y5_W1BEG[0] ;
 wire \Tile_X8Y5_W1BEG[1] ;
 wire \Tile_X8Y5_W1BEG[2] ;
 wire \Tile_X8Y5_W1BEG[3] ;
 wire \Tile_X8Y5_W2BEG[0] ;
 wire \Tile_X8Y5_W2BEG[1] ;
 wire \Tile_X8Y5_W2BEG[2] ;
 wire \Tile_X8Y5_W2BEG[3] ;
 wire \Tile_X8Y5_W2BEG[4] ;
 wire \Tile_X8Y5_W2BEG[5] ;
 wire \Tile_X8Y5_W2BEG[6] ;
 wire \Tile_X8Y5_W2BEG[7] ;
 wire \Tile_X8Y5_W2BEGb[0] ;
 wire \Tile_X8Y5_W2BEGb[1] ;
 wire \Tile_X8Y5_W2BEGb[2] ;
 wire \Tile_X8Y5_W2BEGb[3] ;
 wire \Tile_X8Y5_W2BEGb[4] ;
 wire \Tile_X8Y5_W2BEGb[5] ;
 wire \Tile_X8Y5_W2BEGb[6] ;
 wire \Tile_X8Y5_W2BEGb[7] ;
 wire \Tile_X8Y5_W6BEG[0] ;
 wire \Tile_X8Y5_W6BEG[10] ;
 wire \Tile_X8Y5_W6BEG[11] ;
 wire \Tile_X8Y5_W6BEG[1] ;
 wire \Tile_X8Y5_W6BEG[2] ;
 wire \Tile_X8Y5_W6BEG[3] ;
 wire \Tile_X8Y5_W6BEG[4] ;
 wire \Tile_X8Y5_W6BEG[5] ;
 wire \Tile_X8Y5_W6BEG[6] ;
 wire \Tile_X8Y5_W6BEG[7] ;
 wire \Tile_X8Y5_W6BEG[8] ;
 wire \Tile_X8Y5_W6BEG[9] ;
 wire \Tile_X8Y5_WW4BEG[0] ;
 wire \Tile_X8Y5_WW4BEG[10] ;
 wire \Tile_X8Y5_WW4BEG[11] ;
 wire \Tile_X8Y5_WW4BEG[12] ;
 wire \Tile_X8Y5_WW4BEG[13] ;
 wire \Tile_X8Y5_WW4BEG[14] ;
 wire \Tile_X8Y5_WW4BEG[15] ;
 wire \Tile_X8Y5_WW4BEG[1] ;
 wire \Tile_X8Y5_WW4BEG[2] ;
 wire \Tile_X8Y5_WW4BEG[3] ;
 wire \Tile_X8Y5_WW4BEG[4] ;
 wire \Tile_X8Y5_WW4BEG[5] ;
 wire \Tile_X8Y5_WW4BEG[6] ;
 wire \Tile_X8Y5_WW4BEG[7] ;
 wire \Tile_X8Y5_WW4BEG[8] ;
 wire \Tile_X8Y5_WW4BEG[9] ;
 wire Tile_X8Y6_Co;
 wire \Tile_X8Y6_E1BEG[0] ;
 wire \Tile_X8Y6_E1BEG[1] ;
 wire \Tile_X8Y6_E1BEG[2] ;
 wire \Tile_X8Y6_E1BEG[3] ;
 wire \Tile_X8Y6_E2BEG[0] ;
 wire \Tile_X8Y6_E2BEG[1] ;
 wire \Tile_X8Y6_E2BEG[2] ;
 wire \Tile_X8Y6_E2BEG[3] ;
 wire \Tile_X8Y6_E2BEG[4] ;
 wire \Tile_X8Y6_E2BEG[5] ;
 wire \Tile_X8Y6_E2BEG[6] ;
 wire \Tile_X8Y6_E2BEG[7] ;
 wire \Tile_X8Y6_E2BEGb[0] ;
 wire \Tile_X8Y6_E2BEGb[1] ;
 wire \Tile_X8Y6_E2BEGb[2] ;
 wire \Tile_X8Y6_E2BEGb[3] ;
 wire \Tile_X8Y6_E2BEGb[4] ;
 wire \Tile_X8Y6_E2BEGb[5] ;
 wire \Tile_X8Y6_E2BEGb[6] ;
 wire \Tile_X8Y6_E2BEGb[7] ;
 wire \Tile_X8Y6_E6BEG[0] ;
 wire \Tile_X8Y6_E6BEG[10] ;
 wire \Tile_X8Y6_E6BEG[11] ;
 wire \Tile_X8Y6_E6BEG[1] ;
 wire \Tile_X8Y6_E6BEG[2] ;
 wire \Tile_X8Y6_E6BEG[3] ;
 wire \Tile_X8Y6_E6BEG[4] ;
 wire \Tile_X8Y6_E6BEG[5] ;
 wire \Tile_X8Y6_E6BEG[6] ;
 wire \Tile_X8Y6_E6BEG[7] ;
 wire \Tile_X8Y6_E6BEG[8] ;
 wire \Tile_X8Y6_E6BEG[9] ;
 wire \Tile_X8Y6_EE4BEG[0] ;
 wire \Tile_X8Y6_EE4BEG[10] ;
 wire \Tile_X8Y6_EE4BEG[11] ;
 wire \Tile_X8Y6_EE4BEG[12] ;
 wire \Tile_X8Y6_EE4BEG[13] ;
 wire \Tile_X8Y6_EE4BEG[14] ;
 wire \Tile_X8Y6_EE4BEG[15] ;
 wire \Tile_X8Y6_EE4BEG[1] ;
 wire \Tile_X8Y6_EE4BEG[2] ;
 wire \Tile_X8Y6_EE4BEG[3] ;
 wire \Tile_X8Y6_EE4BEG[4] ;
 wire \Tile_X8Y6_EE4BEG[5] ;
 wire \Tile_X8Y6_EE4BEG[6] ;
 wire \Tile_X8Y6_EE4BEG[7] ;
 wire \Tile_X8Y6_EE4BEG[8] ;
 wire \Tile_X8Y6_EE4BEG[9] ;
 wire \Tile_X8Y6_FrameData_O[0] ;
 wire \Tile_X8Y6_FrameData_O[10] ;
 wire \Tile_X8Y6_FrameData_O[11] ;
 wire \Tile_X8Y6_FrameData_O[12] ;
 wire \Tile_X8Y6_FrameData_O[13] ;
 wire \Tile_X8Y6_FrameData_O[14] ;
 wire \Tile_X8Y6_FrameData_O[15] ;
 wire \Tile_X8Y6_FrameData_O[16] ;
 wire \Tile_X8Y6_FrameData_O[17] ;
 wire \Tile_X8Y6_FrameData_O[18] ;
 wire \Tile_X8Y6_FrameData_O[19] ;
 wire \Tile_X8Y6_FrameData_O[1] ;
 wire \Tile_X8Y6_FrameData_O[20] ;
 wire \Tile_X8Y6_FrameData_O[21] ;
 wire \Tile_X8Y6_FrameData_O[22] ;
 wire \Tile_X8Y6_FrameData_O[23] ;
 wire \Tile_X8Y6_FrameData_O[24] ;
 wire \Tile_X8Y6_FrameData_O[25] ;
 wire \Tile_X8Y6_FrameData_O[26] ;
 wire \Tile_X8Y6_FrameData_O[27] ;
 wire \Tile_X8Y6_FrameData_O[28] ;
 wire \Tile_X8Y6_FrameData_O[29] ;
 wire \Tile_X8Y6_FrameData_O[2] ;
 wire \Tile_X8Y6_FrameData_O[30] ;
 wire \Tile_X8Y6_FrameData_O[31] ;
 wire \Tile_X8Y6_FrameData_O[3] ;
 wire \Tile_X8Y6_FrameData_O[4] ;
 wire \Tile_X8Y6_FrameData_O[5] ;
 wire \Tile_X8Y6_FrameData_O[6] ;
 wire \Tile_X8Y6_FrameData_O[7] ;
 wire \Tile_X8Y6_FrameData_O[8] ;
 wire \Tile_X8Y6_FrameData_O[9] ;
 wire \Tile_X8Y6_FrameStrobe_O[0] ;
 wire \Tile_X8Y6_FrameStrobe_O[10] ;
 wire \Tile_X8Y6_FrameStrobe_O[11] ;
 wire \Tile_X8Y6_FrameStrobe_O[12] ;
 wire \Tile_X8Y6_FrameStrobe_O[13] ;
 wire \Tile_X8Y6_FrameStrobe_O[14] ;
 wire \Tile_X8Y6_FrameStrobe_O[15] ;
 wire \Tile_X8Y6_FrameStrobe_O[16] ;
 wire \Tile_X8Y6_FrameStrobe_O[17] ;
 wire \Tile_X8Y6_FrameStrobe_O[18] ;
 wire \Tile_X8Y6_FrameStrobe_O[19] ;
 wire \Tile_X8Y6_FrameStrobe_O[1] ;
 wire \Tile_X8Y6_FrameStrobe_O[2] ;
 wire \Tile_X8Y6_FrameStrobe_O[3] ;
 wire \Tile_X8Y6_FrameStrobe_O[4] ;
 wire \Tile_X8Y6_FrameStrobe_O[5] ;
 wire \Tile_X8Y6_FrameStrobe_O[6] ;
 wire \Tile_X8Y6_FrameStrobe_O[7] ;
 wire \Tile_X8Y6_FrameStrobe_O[8] ;
 wire \Tile_X8Y6_FrameStrobe_O[9] ;
 wire \Tile_X8Y6_N1BEG[0] ;
 wire \Tile_X8Y6_N1BEG[1] ;
 wire \Tile_X8Y6_N1BEG[2] ;
 wire \Tile_X8Y6_N1BEG[3] ;
 wire \Tile_X8Y6_N2BEG[0] ;
 wire \Tile_X8Y6_N2BEG[1] ;
 wire \Tile_X8Y6_N2BEG[2] ;
 wire \Tile_X8Y6_N2BEG[3] ;
 wire \Tile_X8Y6_N2BEG[4] ;
 wire \Tile_X8Y6_N2BEG[5] ;
 wire \Tile_X8Y6_N2BEG[6] ;
 wire \Tile_X8Y6_N2BEG[7] ;
 wire \Tile_X8Y6_N2BEGb[0] ;
 wire \Tile_X8Y6_N2BEGb[1] ;
 wire \Tile_X8Y6_N2BEGb[2] ;
 wire \Tile_X8Y6_N2BEGb[3] ;
 wire \Tile_X8Y6_N2BEGb[4] ;
 wire \Tile_X8Y6_N2BEGb[5] ;
 wire \Tile_X8Y6_N2BEGb[6] ;
 wire \Tile_X8Y6_N2BEGb[7] ;
 wire \Tile_X8Y6_N4BEG[0] ;
 wire \Tile_X8Y6_N4BEG[10] ;
 wire \Tile_X8Y6_N4BEG[11] ;
 wire \Tile_X8Y6_N4BEG[12] ;
 wire \Tile_X8Y6_N4BEG[13] ;
 wire \Tile_X8Y6_N4BEG[14] ;
 wire \Tile_X8Y6_N4BEG[15] ;
 wire \Tile_X8Y6_N4BEG[1] ;
 wire \Tile_X8Y6_N4BEG[2] ;
 wire \Tile_X8Y6_N4BEG[3] ;
 wire \Tile_X8Y6_N4BEG[4] ;
 wire \Tile_X8Y6_N4BEG[5] ;
 wire \Tile_X8Y6_N4BEG[6] ;
 wire \Tile_X8Y6_N4BEG[7] ;
 wire \Tile_X8Y6_N4BEG[8] ;
 wire \Tile_X8Y6_N4BEG[9] ;
 wire \Tile_X8Y6_NN4BEG[0] ;
 wire \Tile_X8Y6_NN4BEG[10] ;
 wire \Tile_X8Y6_NN4BEG[11] ;
 wire \Tile_X8Y6_NN4BEG[12] ;
 wire \Tile_X8Y6_NN4BEG[13] ;
 wire \Tile_X8Y6_NN4BEG[14] ;
 wire \Tile_X8Y6_NN4BEG[15] ;
 wire \Tile_X8Y6_NN4BEG[1] ;
 wire \Tile_X8Y6_NN4BEG[2] ;
 wire \Tile_X8Y6_NN4BEG[3] ;
 wire \Tile_X8Y6_NN4BEG[4] ;
 wire \Tile_X8Y6_NN4BEG[5] ;
 wire \Tile_X8Y6_NN4BEG[6] ;
 wire \Tile_X8Y6_NN4BEG[7] ;
 wire \Tile_X8Y6_NN4BEG[8] ;
 wire \Tile_X8Y6_NN4BEG[9] ;
 wire \Tile_X8Y6_S1BEG[0] ;
 wire \Tile_X8Y6_S1BEG[1] ;
 wire \Tile_X8Y6_S1BEG[2] ;
 wire \Tile_X8Y6_S1BEG[3] ;
 wire \Tile_X8Y6_S2BEG[0] ;
 wire \Tile_X8Y6_S2BEG[1] ;
 wire \Tile_X8Y6_S2BEG[2] ;
 wire \Tile_X8Y6_S2BEG[3] ;
 wire \Tile_X8Y6_S2BEG[4] ;
 wire \Tile_X8Y6_S2BEG[5] ;
 wire \Tile_X8Y6_S2BEG[6] ;
 wire \Tile_X8Y6_S2BEG[7] ;
 wire \Tile_X8Y6_S2BEGb[0] ;
 wire \Tile_X8Y6_S2BEGb[1] ;
 wire \Tile_X8Y6_S2BEGb[2] ;
 wire \Tile_X8Y6_S2BEGb[3] ;
 wire \Tile_X8Y6_S2BEGb[4] ;
 wire \Tile_X8Y6_S2BEGb[5] ;
 wire \Tile_X8Y6_S2BEGb[6] ;
 wire \Tile_X8Y6_S2BEGb[7] ;
 wire \Tile_X8Y6_S4BEG[0] ;
 wire \Tile_X8Y6_S4BEG[10] ;
 wire \Tile_X8Y6_S4BEG[11] ;
 wire \Tile_X8Y6_S4BEG[12] ;
 wire \Tile_X8Y6_S4BEG[13] ;
 wire \Tile_X8Y6_S4BEG[14] ;
 wire \Tile_X8Y6_S4BEG[15] ;
 wire \Tile_X8Y6_S4BEG[1] ;
 wire \Tile_X8Y6_S4BEG[2] ;
 wire \Tile_X8Y6_S4BEG[3] ;
 wire \Tile_X8Y6_S4BEG[4] ;
 wire \Tile_X8Y6_S4BEG[5] ;
 wire \Tile_X8Y6_S4BEG[6] ;
 wire \Tile_X8Y6_S4BEG[7] ;
 wire \Tile_X8Y6_S4BEG[8] ;
 wire \Tile_X8Y6_S4BEG[9] ;
 wire \Tile_X8Y6_SS4BEG[0] ;
 wire \Tile_X8Y6_SS4BEG[10] ;
 wire \Tile_X8Y6_SS4BEG[11] ;
 wire \Tile_X8Y6_SS4BEG[12] ;
 wire \Tile_X8Y6_SS4BEG[13] ;
 wire \Tile_X8Y6_SS4BEG[14] ;
 wire \Tile_X8Y6_SS4BEG[15] ;
 wire \Tile_X8Y6_SS4BEG[1] ;
 wire \Tile_X8Y6_SS4BEG[2] ;
 wire \Tile_X8Y6_SS4BEG[3] ;
 wire \Tile_X8Y6_SS4BEG[4] ;
 wire \Tile_X8Y6_SS4BEG[5] ;
 wire \Tile_X8Y6_SS4BEG[6] ;
 wire \Tile_X8Y6_SS4BEG[7] ;
 wire \Tile_X8Y6_SS4BEG[8] ;
 wire \Tile_X8Y6_SS4BEG[9] ;
 wire Tile_X8Y6_UserCLKo;
 wire \Tile_X8Y6_W1BEG[0] ;
 wire \Tile_X8Y6_W1BEG[1] ;
 wire \Tile_X8Y6_W1BEG[2] ;
 wire \Tile_X8Y6_W1BEG[3] ;
 wire \Tile_X8Y6_W2BEG[0] ;
 wire \Tile_X8Y6_W2BEG[1] ;
 wire \Tile_X8Y6_W2BEG[2] ;
 wire \Tile_X8Y6_W2BEG[3] ;
 wire \Tile_X8Y6_W2BEG[4] ;
 wire \Tile_X8Y6_W2BEG[5] ;
 wire \Tile_X8Y6_W2BEG[6] ;
 wire \Tile_X8Y6_W2BEG[7] ;
 wire \Tile_X8Y6_W2BEGb[0] ;
 wire \Tile_X8Y6_W2BEGb[1] ;
 wire \Tile_X8Y6_W2BEGb[2] ;
 wire \Tile_X8Y6_W2BEGb[3] ;
 wire \Tile_X8Y6_W2BEGb[4] ;
 wire \Tile_X8Y6_W2BEGb[5] ;
 wire \Tile_X8Y6_W2BEGb[6] ;
 wire \Tile_X8Y6_W2BEGb[7] ;
 wire \Tile_X8Y6_W6BEG[0] ;
 wire \Tile_X8Y6_W6BEG[10] ;
 wire \Tile_X8Y6_W6BEG[11] ;
 wire \Tile_X8Y6_W6BEG[1] ;
 wire \Tile_X8Y6_W6BEG[2] ;
 wire \Tile_X8Y6_W6BEG[3] ;
 wire \Tile_X8Y6_W6BEG[4] ;
 wire \Tile_X8Y6_W6BEG[5] ;
 wire \Tile_X8Y6_W6BEG[6] ;
 wire \Tile_X8Y6_W6BEG[7] ;
 wire \Tile_X8Y6_W6BEG[8] ;
 wire \Tile_X8Y6_W6BEG[9] ;
 wire \Tile_X8Y6_WW4BEG[0] ;
 wire \Tile_X8Y6_WW4BEG[10] ;
 wire \Tile_X8Y6_WW4BEG[11] ;
 wire \Tile_X8Y6_WW4BEG[12] ;
 wire \Tile_X8Y6_WW4BEG[13] ;
 wire \Tile_X8Y6_WW4BEG[14] ;
 wire \Tile_X8Y6_WW4BEG[15] ;
 wire \Tile_X8Y6_WW4BEG[1] ;
 wire \Tile_X8Y6_WW4BEG[2] ;
 wire \Tile_X8Y6_WW4BEG[3] ;
 wire \Tile_X8Y6_WW4BEG[4] ;
 wire \Tile_X8Y6_WW4BEG[5] ;
 wire \Tile_X8Y6_WW4BEG[6] ;
 wire \Tile_X8Y6_WW4BEG[7] ;
 wire \Tile_X8Y6_WW4BEG[8] ;
 wire \Tile_X8Y6_WW4BEG[9] ;
 wire Tile_X8Y7_Co;
 wire \Tile_X8Y7_E1BEG[0] ;
 wire \Tile_X8Y7_E1BEG[1] ;
 wire \Tile_X8Y7_E1BEG[2] ;
 wire \Tile_X8Y7_E1BEG[3] ;
 wire \Tile_X8Y7_E2BEG[0] ;
 wire \Tile_X8Y7_E2BEG[1] ;
 wire \Tile_X8Y7_E2BEG[2] ;
 wire \Tile_X8Y7_E2BEG[3] ;
 wire \Tile_X8Y7_E2BEG[4] ;
 wire \Tile_X8Y7_E2BEG[5] ;
 wire \Tile_X8Y7_E2BEG[6] ;
 wire \Tile_X8Y7_E2BEG[7] ;
 wire \Tile_X8Y7_E2BEGb[0] ;
 wire \Tile_X8Y7_E2BEGb[1] ;
 wire \Tile_X8Y7_E2BEGb[2] ;
 wire \Tile_X8Y7_E2BEGb[3] ;
 wire \Tile_X8Y7_E2BEGb[4] ;
 wire \Tile_X8Y7_E2BEGb[5] ;
 wire \Tile_X8Y7_E2BEGb[6] ;
 wire \Tile_X8Y7_E2BEGb[7] ;
 wire \Tile_X8Y7_E6BEG[0] ;
 wire \Tile_X8Y7_E6BEG[10] ;
 wire \Tile_X8Y7_E6BEG[11] ;
 wire \Tile_X8Y7_E6BEG[1] ;
 wire \Tile_X8Y7_E6BEG[2] ;
 wire \Tile_X8Y7_E6BEG[3] ;
 wire \Tile_X8Y7_E6BEG[4] ;
 wire \Tile_X8Y7_E6BEG[5] ;
 wire \Tile_X8Y7_E6BEG[6] ;
 wire \Tile_X8Y7_E6BEG[7] ;
 wire \Tile_X8Y7_E6BEG[8] ;
 wire \Tile_X8Y7_E6BEG[9] ;
 wire \Tile_X8Y7_EE4BEG[0] ;
 wire \Tile_X8Y7_EE4BEG[10] ;
 wire \Tile_X8Y7_EE4BEG[11] ;
 wire \Tile_X8Y7_EE4BEG[12] ;
 wire \Tile_X8Y7_EE4BEG[13] ;
 wire \Tile_X8Y7_EE4BEG[14] ;
 wire \Tile_X8Y7_EE4BEG[15] ;
 wire \Tile_X8Y7_EE4BEG[1] ;
 wire \Tile_X8Y7_EE4BEG[2] ;
 wire \Tile_X8Y7_EE4BEG[3] ;
 wire \Tile_X8Y7_EE4BEG[4] ;
 wire \Tile_X8Y7_EE4BEG[5] ;
 wire \Tile_X8Y7_EE4BEG[6] ;
 wire \Tile_X8Y7_EE4BEG[7] ;
 wire \Tile_X8Y7_EE4BEG[8] ;
 wire \Tile_X8Y7_EE4BEG[9] ;
 wire \Tile_X8Y7_FrameData_O[0] ;
 wire \Tile_X8Y7_FrameData_O[10] ;
 wire \Tile_X8Y7_FrameData_O[11] ;
 wire \Tile_X8Y7_FrameData_O[12] ;
 wire \Tile_X8Y7_FrameData_O[13] ;
 wire \Tile_X8Y7_FrameData_O[14] ;
 wire \Tile_X8Y7_FrameData_O[15] ;
 wire \Tile_X8Y7_FrameData_O[16] ;
 wire \Tile_X8Y7_FrameData_O[17] ;
 wire \Tile_X8Y7_FrameData_O[18] ;
 wire \Tile_X8Y7_FrameData_O[19] ;
 wire \Tile_X8Y7_FrameData_O[1] ;
 wire \Tile_X8Y7_FrameData_O[20] ;
 wire \Tile_X8Y7_FrameData_O[21] ;
 wire \Tile_X8Y7_FrameData_O[22] ;
 wire \Tile_X8Y7_FrameData_O[23] ;
 wire \Tile_X8Y7_FrameData_O[24] ;
 wire \Tile_X8Y7_FrameData_O[25] ;
 wire \Tile_X8Y7_FrameData_O[26] ;
 wire \Tile_X8Y7_FrameData_O[27] ;
 wire \Tile_X8Y7_FrameData_O[28] ;
 wire \Tile_X8Y7_FrameData_O[29] ;
 wire \Tile_X8Y7_FrameData_O[2] ;
 wire \Tile_X8Y7_FrameData_O[30] ;
 wire \Tile_X8Y7_FrameData_O[31] ;
 wire \Tile_X8Y7_FrameData_O[3] ;
 wire \Tile_X8Y7_FrameData_O[4] ;
 wire \Tile_X8Y7_FrameData_O[5] ;
 wire \Tile_X8Y7_FrameData_O[6] ;
 wire \Tile_X8Y7_FrameData_O[7] ;
 wire \Tile_X8Y7_FrameData_O[8] ;
 wire \Tile_X8Y7_FrameData_O[9] ;
 wire \Tile_X8Y7_FrameStrobe_O[0] ;
 wire \Tile_X8Y7_FrameStrobe_O[10] ;
 wire \Tile_X8Y7_FrameStrobe_O[11] ;
 wire \Tile_X8Y7_FrameStrobe_O[12] ;
 wire \Tile_X8Y7_FrameStrobe_O[13] ;
 wire \Tile_X8Y7_FrameStrobe_O[14] ;
 wire \Tile_X8Y7_FrameStrobe_O[15] ;
 wire \Tile_X8Y7_FrameStrobe_O[16] ;
 wire \Tile_X8Y7_FrameStrobe_O[17] ;
 wire \Tile_X8Y7_FrameStrobe_O[18] ;
 wire \Tile_X8Y7_FrameStrobe_O[19] ;
 wire \Tile_X8Y7_FrameStrobe_O[1] ;
 wire \Tile_X8Y7_FrameStrobe_O[2] ;
 wire \Tile_X8Y7_FrameStrobe_O[3] ;
 wire \Tile_X8Y7_FrameStrobe_O[4] ;
 wire \Tile_X8Y7_FrameStrobe_O[5] ;
 wire \Tile_X8Y7_FrameStrobe_O[6] ;
 wire \Tile_X8Y7_FrameStrobe_O[7] ;
 wire \Tile_X8Y7_FrameStrobe_O[8] ;
 wire \Tile_X8Y7_FrameStrobe_O[9] ;
 wire \Tile_X8Y7_N1BEG[0] ;
 wire \Tile_X8Y7_N1BEG[1] ;
 wire \Tile_X8Y7_N1BEG[2] ;
 wire \Tile_X8Y7_N1BEG[3] ;
 wire \Tile_X8Y7_N2BEG[0] ;
 wire \Tile_X8Y7_N2BEG[1] ;
 wire \Tile_X8Y7_N2BEG[2] ;
 wire \Tile_X8Y7_N2BEG[3] ;
 wire \Tile_X8Y7_N2BEG[4] ;
 wire \Tile_X8Y7_N2BEG[5] ;
 wire \Tile_X8Y7_N2BEG[6] ;
 wire \Tile_X8Y7_N2BEG[7] ;
 wire \Tile_X8Y7_N2BEGb[0] ;
 wire \Tile_X8Y7_N2BEGb[1] ;
 wire \Tile_X8Y7_N2BEGb[2] ;
 wire \Tile_X8Y7_N2BEGb[3] ;
 wire \Tile_X8Y7_N2BEGb[4] ;
 wire \Tile_X8Y7_N2BEGb[5] ;
 wire \Tile_X8Y7_N2BEGb[6] ;
 wire \Tile_X8Y7_N2BEGb[7] ;
 wire \Tile_X8Y7_N4BEG[0] ;
 wire \Tile_X8Y7_N4BEG[10] ;
 wire \Tile_X8Y7_N4BEG[11] ;
 wire \Tile_X8Y7_N4BEG[12] ;
 wire \Tile_X8Y7_N4BEG[13] ;
 wire \Tile_X8Y7_N4BEG[14] ;
 wire \Tile_X8Y7_N4BEG[15] ;
 wire \Tile_X8Y7_N4BEG[1] ;
 wire \Tile_X8Y7_N4BEG[2] ;
 wire \Tile_X8Y7_N4BEG[3] ;
 wire \Tile_X8Y7_N4BEG[4] ;
 wire \Tile_X8Y7_N4BEG[5] ;
 wire \Tile_X8Y7_N4BEG[6] ;
 wire \Tile_X8Y7_N4BEG[7] ;
 wire \Tile_X8Y7_N4BEG[8] ;
 wire \Tile_X8Y7_N4BEG[9] ;
 wire \Tile_X8Y7_NN4BEG[0] ;
 wire \Tile_X8Y7_NN4BEG[10] ;
 wire \Tile_X8Y7_NN4BEG[11] ;
 wire \Tile_X8Y7_NN4BEG[12] ;
 wire \Tile_X8Y7_NN4BEG[13] ;
 wire \Tile_X8Y7_NN4BEG[14] ;
 wire \Tile_X8Y7_NN4BEG[15] ;
 wire \Tile_X8Y7_NN4BEG[1] ;
 wire \Tile_X8Y7_NN4BEG[2] ;
 wire \Tile_X8Y7_NN4BEG[3] ;
 wire \Tile_X8Y7_NN4BEG[4] ;
 wire \Tile_X8Y7_NN4BEG[5] ;
 wire \Tile_X8Y7_NN4BEG[6] ;
 wire \Tile_X8Y7_NN4BEG[7] ;
 wire \Tile_X8Y7_NN4BEG[8] ;
 wire \Tile_X8Y7_NN4BEG[9] ;
 wire \Tile_X8Y7_S1BEG[0] ;
 wire \Tile_X8Y7_S1BEG[1] ;
 wire \Tile_X8Y7_S1BEG[2] ;
 wire \Tile_X8Y7_S1BEG[3] ;
 wire \Tile_X8Y7_S2BEG[0] ;
 wire \Tile_X8Y7_S2BEG[1] ;
 wire \Tile_X8Y7_S2BEG[2] ;
 wire \Tile_X8Y7_S2BEG[3] ;
 wire \Tile_X8Y7_S2BEG[4] ;
 wire \Tile_X8Y7_S2BEG[5] ;
 wire \Tile_X8Y7_S2BEG[6] ;
 wire \Tile_X8Y7_S2BEG[7] ;
 wire \Tile_X8Y7_S2BEGb[0] ;
 wire \Tile_X8Y7_S2BEGb[1] ;
 wire \Tile_X8Y7_S2BEGb[2] ;
 wire \Tile_X8Y7_S2BEGb[3] ;
 wire \Tile_X8Y7_S2BEGb[4] ;
 wire \Tile_X8Y7_S2BEGb[5] ;
 wire \Tile_X8Y7_S2BEGb[6] ;
 wire \Tile_X8Y7_S2BEGb[7] ;
 wire \Tile_X8Y7_S4BEG[0] ;
 wire \Tile_X8Y7_S4BEG[10] ;
 wire \Tile_X8Y7_S4BEG[11] ;
 wire \Tile_X8Y7_S4BEG[12] ;
 wire \Tile_X8Y7_S4BEG[13] ;
 wire \Tile_X8Y7_S4BEG[14] ;
 wire \Tile_X8Y7_S4BEG[15] ;
 wire \Tile_X8Y7_S4BEG[1] ;
 wire \Tile_X8Y7_S4BEG[2] ;
 wire \Tile_X8Y7_S4BEG[3] ;
 wire \Tile_X8Y7_S4BEG[4] ;
 wire \Tile_X8Y7_S4BEG[5] ;
 wire \Tile_X8Y7_S4BEG[6] ;
 wire \Tile_X8Y7_S4BEG[7] ;
 wire \Tile_X8Y7_S4BEG[8] ;
 wire \Tile_X8Y7_S4BEG[9] ;
 wire \Tile_X8Y7_SS4BEG[0] ;
 wire \Tile_X8Y7_SS4BEG[10] ;
 wire \Tile_X8Y7_SS4BEG[11] ;
 wire \Tile_X8Y7_SS4BEG[12] ;
 wire \Tile_X8Y7_SS4BEG[13] ;
 wire \Tile_X8Y7_SS4BEG[14] ;
 wire \Tile_X8Y7_SS4BEG[15] ;
 wire \Tile_X8Y7_SS4BEG[1] ;
 wire \Tile_X8Y7_SS4BEG[2] ;
 wire \Tile_X8Y7_SS4BEG[3] ;
 wire \Tile_X8Y7_SS4BEG[4] ;
 wire \Tile_X8Y7_SS4BEG[5] ;
 wire \Tile_X8Y7_SS4BEG[6] ;
 wire \Tile_X8Y7_SS4BEG[7] ;
 wire \Tile_X8Y7_SS4BEG[8] ;
 wire \Tile_X8Y7_SS4BEG[9] ;
 wire Tile_X8Y7_UserCLKo;
 wire \Tile_X8Y7_W1BEG[0] ;
 wire \Tile_X8Y7_W1BEG[1] ;
 wire \Tile_X8Y7_W1BEG[2] ;
 wire \Tile_X8Y7_W1BEG[3] ;
 wire \Tile_X8Y7_W2BEG[0] ;
 wire \Tile_X8Y7_W2BEG[1] ;
 wire \Tile_X8Y7_W2BEG[2] ;
 wire \Tile_X8Y7_W2BEG[3] ;
 wire \Tile_X8Y7_W2BEG[4] ;
 wire \Tile_X8Y7_W2BEG[5] ;
 wire \Tile_X8Y7_W2BEG[6] ;
 wire \Tile_X8Y7_W2BEG[7] ;
 wire \Tile_X8Y7_W2BEGb[0] ;
 wire \Tile_X8Y7_W2BEGb[1] ;
 wire \Tile_X8Y7_W2BEGb[2] ;
 wire \Tile_X8Y7_W2BEGb[3] ;
 wire \Tile_X8Y7_W2BEGb[4] ;
 wire \Tile_X8Y7_W2BEGb[5] ;
 wire \Tile_X8Y7_W2BEGb[6] ;
 wire \Tile_X8Y7_W2BEGb[7] ;
 wire \Tile_X8Y7_W6BEG[0] ;
 wire \Tile_X8Y7_W6BEG[10] ;
 wire \Tile_X8Y7_W6BEG[11] ;
 wire \Tile_X8Y7_W6BEG[1] ;
 wire \Tile_X8Y7_W6BEG[2] ;
 wire \Tile_X8Y7_W6BEG[3] ;
 wire \Tile_X8Y7_W6BEG[4] ;
 wire \Tile_X8Y7_W6BEG[5] ;
 wire \Tile_X8Y7_W6BEG[6] ;
 wire \Tile_X8Y7_W6BEG[7] ;
 wire \Tile_X8Y7_W6BEG[8] ;
 wire \Tile_X8Y7_W6BEG[9] ;
 wire \Tile_X8Y7_WW4BEG[0] ;
 wire \Tile_X8Y7_WW4BEG[10] ;
 wire \Tile_X8Y7_WW4BEG[11] ;
 wire \Tile_X8Y7_WW4BEG[12] ;
 wire \Tile_X8Y7_WW4BEG[13] ;
 wire \Tile_X8Y7_WW4BEG[14] ;
 wire \Tile_X8Y7_WW4BEG[15] ;
 wire \Tile_X8Y7_WW4BEG[1] ;
 wire \Tile_X8Y7_WW4BEG[2] ;
 wire \Tile_X8Y7_WW4BEG[3] ;
 wire \Tile_X8Y7_WW4BEG[4] ;
 wire \Tile_X8Y7_WW4BEG[5] ;
 wire \Tile_X8Y7_WW4BEG[6] ;
 wire \Tile_X8Y7_WW4BEG[7] ;
 wire \Tile_X8Y7_WW4BEG[8] ;
 wire \Tile_X8Y7_WW4BEG[9] ;
 wire Tile_X8Y8_Co;
 wire \Tile_X8Y8_E1BEG[0] ;
 wire \Tile_X8Y8_E1BEG[1] ;
 wire \Tile_X8Y8_E1BEG[2] ;
 wire \Tile_X8Y8_E1BEG[3] ;
 wire \Tile_X8Y8_E2BEG[0] ;
 wire \Tile_X8Y8_E2BEG[1] ;
 wire \Tile_X8Y8_E2BEG[2] ;
 wire \Tile_X8Y8_E2BEG[3] ;
 wire \Tile_X8Y8_E2BEG[4] ;
 wire \Tile_X8Y8_E2BEG[5] ;
 wire \Tile_X8Y8_E2BEG[6] ;
 wire \Tile_X8Y8_E2BEG[7] ;
 wire \Tile_X8Y8_E2BEGb[0] ;
 wire \Tile_X8Y8_E2BEGb[1] ;
 wire \Tile_X8Y8_E2BEGb[2] ;
 wire \Tile_X8Y8_E2BEGb[3] ;
 wire \Tile_X8Y8_E2BEGb[4] ;
 wire \Tile_X8Y8_E2BEGb[5] ;
 wire \Tile_X8Y8_E2BEGb[6] ;
 wire \Tile_X8Y8_E2BEGb[7] ;
 wire \Tile_X8Y8_E6BEG[0] ;
 wire \Tile_X8Y8_E6BEG[10] ;
 wire \Tile_X8Y8_E6BEG[11] ;
 wire \Tile_X8Y8_E6BEG[1] ;
 wire \Tile_X8Y8_E6BEG[2] ;
 wire \Tile_X8Y8_E6BEG[3] ;
 wire \Tile_X8Y8_E6BEG[4] ;
 wire \Tile_X8Y8_E6BEG[5] ;
 wire \Tile_X8Y8_E6BEG[6] ;
 wire \Tile_X8Y8_E6BEG[7] ;
 wire \Tile_X8Y8_E6BEG[8] ;
 wire \Tile_X8Y8_E6BEG[9] ;
 wire \Tile_X8Y8_EE4BEG[0] ;
 wire \Tile_X8Y8_EE4BEG[10] ;
 wire \Tile_X8Y8_EE4BEG[11] ;
 wire \Tile_X8Y8_EE4BEG[12] ;
 wire \Tile_X8Y8_EE4BEG[13] ;
 wire \Tile_X8Y8_EE4BEG[14] ;
 wire \Tile_X8Y8_EE4BEG[15] ;
 wire \Tile_X8Y8_EE4BEG[1] ;
 wire \Tile_X8Y8_EE4BEG[2] ;
 wire \Tile_X8Y8_EE4BEG[3] ;
 wire \Tile_X8Y8_EE4BEG[4] ;
 wire \Tile_X8Y8_EE4BEG[5] ;
 wire \Tile_X8Y8_EE4BEG[6] ;
 wire \Tile_X8Y8_EE4BEG[7] ;
 wire \Tile_X8Y8_EE4BEG[8] ;
 wire \Tile_X8Y8_EE4BEG[9] ;
 wire \Tile_X8Y8_FrameData_O[0] ;
 wire \Tile_X8Y8_FrameData_O[10] ;
 wire \Tile_X8Y8_FrameData_O[11] ;
 wire \Tile_X8Y8_FrameData_O[12] ;
 wire \Tile_X8Y8_FrameData_O[13] ;
 wire \Tile_X8Y8_FrameData_O[14] ;
 wire \Tile_X8Y8_FrameData_O[15] ;
 wire \Tile_X8Y8_FrameData_O[16] ;
 wire \Tile_X8Y8_FrameData_O[17] ;
 wire \Tile_X8Y8_FrameData_O[18] ;
 wire \Tile_X8Y8_FrameData_O[19] ;
 wire \Tile_X8Y8_FrameData_O[1] ;
 wire \Tile_X8Y8_FrameData_O[20] ;
 wire \Tile_X8Y8_FrameData_O[21] ;
 wire \Tile_X8Y8_FrameData_O[22] ;
 wire \Tile_X8Y8_FrameData_O[23] ;
 wire \Tile_X8Y8_FrameData_O[24] ;
 wire \Tile_X8Y8_FrameData_O[25] ;
 wire \Tile_X8Y8_FrameData_O[26] ;
 wire \Tile_X8Y8_FrameData_O[27] ;
 wire \Tile_X8Y8_FrameData_O[28] ;
 wire \Tile_X8Y8_FrameData_O[29] ;
 wire \Tile_X8Y8_FrameData_O[2] ;
 wire \Tile_X8Y8_FrameData_O[30] ;
 wire \Tile_X8Y8_FrameData_O[31] ;
 wire \Tile_X8Y8_FrameData_O[3] ;
 wire \Tile_X8Y8_FrameData_O[4] ;
 wire \Tile_X8Y8_FrameData_O[5] ;
 wire \Tile_X8Y8_FrameData_O[6] ;
 wire \Tile_X8Y8_FrameData_O[7] ;
 wire \Tile_X8Y8_FrameData_O[8] ;
 wire \Tile_X8Y8_FrameData_O[9] ;
 wire \Tile_X8Y8_FrameStrobe_O[0] ;
 wire \Tile_X8Y8_FrameStrobe_O[10] ;
 wire \Tile_X8Y8_FrameStrobe_O[11] ;
 wire \Tile_X8Y8_FrameStrobe_O[12] ;
 wire \Tile_X8Y8_FrameStrobe_O[13] ;
 wire \Tile_X8Y8_FrameStrobe_O[14] ;
 wire \Tile_X8Y8_FrameStrobe_O[15] ;
 wire \Tile_X8Y8_FrameStrobe_O[16] ;
 wire \Tile_X8Y8_FrameStrobe_O[17] ;
 wire \Tile_X8Y8_FrameStrobe_O[18] ;
 wire \Tile_X8Y8_FrameStrobe_O[19] ;
 wire \Tile_X8Y8_FrameStrobe_O[1] ;
 wire \Tile_X8Y8_FrameStrobe_O[2] ;
 wire \Tile_X8Y8_FrameStrobe_O[3] ;
 wire \Tile_X8Y8_FrameStrobe_O[4] ;
 wire \Tile_X8Y8_FrameStrobe_O[5] ;
 wire \Tile_X8Y8_FrameStrobe_O[6] ;
 wire \Tile_X8Y8_FrameStrobe_O[7] ;
 wire \Tile_X8Y8_FrameStrobe_O[8] ;
 wire \Tile_X8Y8_FrameStrobe_O[9] ;
 wire \Tile_X8Y8_N1BEG[0] ;
 wire \Tile_X8Y8_N1BEG[1] ;
 wire \Tile_X8Y8_N1BEG[2] ;
 wire \Tile_X8Y8_N1BEG[3] ;
 wire \Tile_X8Y8_N2BEG[0] ;
 wire \Tile_X8Y8_N2BEG[1] ;
 wire \Tile_X8Y8_N2BEG[2] ;
 wire \Tile_X8Y8_N2BEG[3] ;
 wire \Tile_X8Y8_N2BEG[4] ;
 wire \Tile_X8Y8_N2BEG[5] ;
 wire \Tile_X8Y8_N2BEG[6] ;
 wire \Tile_X8Y8_N2BEG[7] ;
 wire \Tile_X8Y8_N2BEGb[0] ;
 wire \Tile_X8Y8_N2BEGb[1] ;
 wire \Tile_X8Y8_N2BEGb[2] ;
 wire \Tile_X8Y8_N2BEGb[3] ;
 wire \Tile_X8Y8_N2BEGb[4] ;
 wire \Tile_X8Y8_N2BEGb[5] ;
 wire \Tile_X8Y8_N2BEGb[6] ;
 wire \Tile_X8Y8_N2BEGb[7] ;
 wire \Tile_X8Y8_N4BEG[0] ;
 wire \Tile_X8Y8_N4BEG[10] ;
 wire \Tile_X8Y8_N4BEG[11] ;
 wire \Tile_X8Y8_N4BEG[12] ;
 wire \Tile_X8Y8_N4BEG[13] ;
 wire \Tile_X8Y8_N4BEG[14] ;
 wire \Tile_X8Y8_N4BEG[15] ;
 wire \Tile_X8Y8_N4BEG[1] ;
 wire \Tile_X8Y8_N4BEG[2] ;
 wire \Tile_X8Y8_N4BEG[3] ;
 wire \Tile_X8Y8_N4BEG[4] ;
 wire \Tile_X8Y8_N4BEG[5] ;
 wire \Tile_X8Y8_N4BEG[6] ;
 wire \Tile_X8Y8_N4BEG[7] ;
 wire \Tile_X8Y8_N4BEG[8] ;
 wire \Tile_X8Y8_N4BEG[9] ;
 wire \Tile_X8Y8_NN4BEG[0] ;
 wire \Tile_X8Y8_NN4BEG[10] ;
 wire \Tile_X8Y8_NN4BEG[11] ;
 wire \Tile_X8Y8_NN4BEG[12] ;
 wire \Tile_X8Y8_NN4BEG[13] ;
 wire \Tile_X8Y8_NN4BEG[14] ;
 wire \Tile_X8Y8_NN4BEG[15] ;
 wire \Tile_X8Y8_NN4BEG[1] ;
 wire \Tile_X8Y8_NN4BEG[2] ;
 wire \Tile_X8Y8_NN4BEG[3] ;
 wire \Tile_X8Y8_NN4BEG[4] ;
 wire \Tile_X8Y8_NN4BEG[5] ;
 wire \Tile_X8Y8_NN4BEG[6] ;
 wire \Tile_X8Y8_NN4BEG[7] ;
 wire \Tile_X8Y8_NN4BEG[8] ;
 wire \Tile_X8Y8_NN4BEG[9] ;
 wire \Tile_X8Y8_S1BEG[0] ;
 wire \Tile_X8Y8_S1BEG[1] ;
 wire \Tile_X8Y8_S1BEG[2] ;
 wire \Tile_X8Y8_S1BEG[3] ;
 wire \Tile_X8Y8_S2BEG[0] ;
 wire \Tile_X8Y8_S2BEG[1] ;
 wire \Tile_X8Y8_S2BEG[2] ;
 wire \Tile_X8Y8_S2BEG[3] ;
 wire \Tile_X8Y8_S2BEG[4] ;
 wire \Tile_X8Y8_S2BEG[5] ;
 wire \Tile_X8Y8_S2BEG[6] ;
 wire \Tile_X8Y8_S2BEG[7] ;
 wire \Tile_X8Y8_S2BEGb[0] ;
 wire \Tile_X8Y8_S2BEGb[1] ;
 wire \Tile_X8Y8_S2BEGb[2] ;
 wire \Tile_X8Y8_S2BEGb[3] ;
 wire \Tile_X8Y8_S2BEGb[4] ;
 wire \Tile_X8Y8_S2BEGb[5] ;
 wire \Tile_X8Y8_S2BEGb[6] ;
 wire \Tile_X8Y8_S2BEGb[7] ;
 wire \Tile_X8Y8_S4BEG[0] ;
 wire \Tile_X8Y8_S4BEG[10] ;
 wire \Tile_X8Y8_S4BEG[11] ;
 wire \Tile_X8Y8_S4BEG[12] ;
 wire \Tile_X8Y8_S4BEG[13] ;
 wire \Tile_X8Y8_S4BEG[14] ;
 wire \Tile_X8Y8_S4BEG[15] ;
 wire \Tile_X8Y8_S4BEG[1] ;
 wire \Tile_X8Y8_S4BEG[2] ;
 wire \Tile_X8Y8_S4BEG[3] ;
 wire \Tile_X8Y8_S4BEG[4] ;
 wire \Tile_X8Y8_S4BEG[5] ;
 wire \Tile_X8Y8_S4BEG[6] ;
 wire \Tile_X8Y8_S4BEG[7] ;
 wire \Tile_X8Y8_S4BEG[8] ;
 wire \Tile_X8Y8_S4BEG[9] ;
 wire \Tile_X8Y8_SS4BEG[0] ;
 wire \Tile_X8Y8_SS4BEG[10] ;
 wire \Tile_X8Y8_SS4BEG[11] ;
 wire \Tile_X8Y8_SS4BEG[12] ;
 wire \Tile_X8Y8_SS4BEG[13] ;
 wire \Tile_X8Y8_SS4BEG[14] ;
 wire \Tile_X8Y8_SS4BEG[15] ;
 wire \Tile_X8Y8_SS4BEG[1] ;
 wire \Tile_X8Y8_SS4BEG[2] ;
 wire \Tile_X8Y8_SS4BEG[3] ;
 wire \Tile_X8Y8_SS4BEG[4] ;
 wire \Tile_X8Y8_SS4BEG[5] ;
 wire \Tile_X8Y8_SS4BEG[6] ;
 wire \Tile_X8Y8_SS4BEG[7] ;
 wire \Tile_X8Y8_SS4BEG[8] ;
 wire \Tile_X8Y8_SS4BEG[9] ;
 wire Tile_X8Y8_UserCLKo;
 wire \Tile_X8Y8_W1BEG[0] ;
 wire \Tile_X8Y8_W1BEG[1] ;
 wire \Tile_X8Y8_W1BEG[2] ;
 wire \Tile_X8Y8_W1BEG[3] ;
 wire \Tile_X8Y8_W2BEG[0] ;
 wire \Tile_X8Y8_W2BEG[1] ;
 wire \Tile_X8Y8_W2BEG[2] ;
 wire \Tile_X8Y8_W2BEG[3] ;
 wire \Tile_X8Y8_W2BEG[4] ;
 wire \Tile_X8Y8_W2BEG[5] ;
 wire \Tile_X8Y8_W2BEG[6] ;
 wire \Tile_X8Y8_W2BEG[7] ;
 wire \Tile_X8Y8_W2BEGb[0] ;
 wire \Tile_X8Y8_W2BEGb[1] ;
 wire \Tile_X8Y8_W2BEGb[2] ;
 wire \Tile_X8Y8_W2BEGb[3] ;
 wire \Tile_X8Y8_W2BEGb[4] ;
 wire \Tile_X8Y8_W2BEGb[5] ;
 wire \Tile_X8Y8_W2BEGb[6] ;
 wire \Tile_X8Y8_W2BEGb[7] ;
 wire \Tile_X8Y8_W6BEG[0] ;
 wire \Tile_X8Y8_W6BEG[10] ;
 wire \Tile_X8Y8_W6BEG[11] ;
 wire \Tile_X8Y8_W6BEG[1] ;
 wire \Tile_X8Y8_W6BEG[2] ;
 wire \Tile_X8Y8_W6BEG[3] ;
 wire \Tile_X8Y8_W6BEG[4] ;
 wire \Tile_X8Y8_W6BEG[5] ;
 wire \Tile_X8Y8_W6BEG[6] ;
 wire \Tile_X8Y8_W6BEG[7] ;
 wire \Tile_X8Y8_W6BEG[8] ;
 wire \Tile_X8Y8_W6BEG[9] ;
 wire \Tile_X8Y8_WW4BEG[0] ;
 wire \Tile_X8Y8_WW4BEG[10] ;
 wire \Tile_X8Y8_WW4BEG[11] ;
 wire \Tile_X8Y8_WW4BEG[12] ;
 wire \Tile_X8Y8_WW4BEG[13] ;
 wire \Tile_X8Y8_WW4BEG[14] ;
 wire \Tile_X8Y8_WW4BEG[15] ;
 wire \Tile_X8Y8_WW4BEG[1] ;
 wire \Tile_X8Y8_WW4BEG[2] ;
 wire \Tile_X8Y8_WW4BEG[3] ;
 wire \Tile_X8Y8_WW4BEG[4] ;
 wire \Tile_X8Y8_WW4BEG[5] ;
 wire \Tile_X8Y8_WW4BEG[6] ;
 wire \Tile_X8Y8_WW4BEG[7] ;
 wire \Tile_X8Y8_WW4BEG[8] ;
 wire \Tile_X8Y8_WW4BEG[9] ;
 wire Tile_X8Y9_Co;
 wire \Tile_X8Y9_E1BEG[0] ;
 wire \Tile_X8Y9_E1BEG[1] ;
 wire \Tile_X8Y9_E1BEG[2] ;
 wire \Tile_X8Y9_E1BEG[3] ;
 wire \Tile_X8Y9_E2BEG[0] ;
 wire \Tile_X8Y9_E2BEG[1] ;
 wire \Tile_X8Y9_E2BEG[2] ;
 wire \Tile_X8Y9_E2BEG[3] ;
 wire \Tile_X8Y9_E2BEG[4] ;
 wire \Tile_X8Y9_E2BEG[5] ;
 wire \Tile_X8Y9_E2BEG[6] ;
 wire \Tile_X8Y9_E2BEG[7] ;
 wire \Tile_X8Y9_E2BEGb[0] ;
 wire \Tile_X8Y9_E2BEGb[1] ;
 wire \Tile_X8Y9_E2BEGb[2] ;
 wire \Tile_X8Y9_E2BEGb[3] ;
 wire \Tile_X8Y9_E2BEGb[4] ;
 wire \Tile_X8Y9_E2BEGb[5] ;
 wire \Tile_X8Y9_E2BEGb[6] ;
 wire \Tile_X8Y9_E2BEGb[7] ;
 wire \Tile_X8Y9_E6BEG[0] ;
 wire \Tile_X8Y9_E6BEG[10] ;
 wire \Tile_X8Y9_E6BEG[11] ;
 wire \Tile_X8Y9_E6BEG[1] ;
 wire \Tile_X8Y9_E6BEG[2] ;
 wire \Tile_X8Y9_E6BEG[3] ;
 wire \Tile_X8Y9_E6BEG[4] ;
 wire \Tile_X8Y9_E6BEG[5] ;
 wire \Tile_X8Y9_E6BEG[6] ;
 wire \Tile_X8Y9_E6BEG[7] ;
 wire \Tile_X8Y9_E6BEG[8] ;
 wire \Tile_X8Y9_E6BEG[9] ;
 wire \Tile_X8Y9_EE4BEG[0] ;
 wire \Tile_X8Y9_EE4BEG[10] ;
 wire \Tile_X8Y9_EE4BEG[11] ;
 wire \Tile_X8Y9_EE4BEG[12] ;
 wire \Tile_X8Y9_EE4BEG[13] ;
 wire \Tile_X8Y9_EE4BEG[14] ;
 wire \Tile_X8Y9_EE4BEG[15] ;
 wire \Tile_X8Y9_EE4BEG[1] ;
 wire \Tile_X8Y9_EE4BEG[2] ;
 wire \Tile_X8Y9_EE4BEG[3] ;
 wire \Tile_X8Y9_EE4BEG[4] ;
 wire \Tile_X8Y9_EE4BEG[5] ;
 wire \Tile_X8Y9_EE4BEG[6] ;
 wire \Tile_X8Y9_EE4BEG[7] ;
 wire \Tile_X8Y9_EE4BEG[8] ;
 wire \Tile_X8Y9_EE4BEG[9] ;
 wire \Tile_X8Y9_FrameData_O[0] ;
 wire \Tile_X8Y9_FrameData_O[10] ;
 wire \Tile_X8Y9_FrameData_O[11] ;
 wire \Tile_X8Y9_FrameData_O[12] ;
 wire \Tile_X8Y9_FrameData_O[13] ;
 wire \Tile_X8Y9_FrameData_O[14] ;
 wire \Tile_X8Y9_FrameData_O[15] ;
 wire \Tile_X8Y9_FrameData_O[16] ;
 wire \Tile_X8Y9_FrameData_O[17] ;
 wire \Tile_X8Y9_FrameData_O[18] ;
 wire \Tile_X8Y9_FrameData_O[19] ;
 wire \Tile_X8Y9_FrameData_O[1] ;
 wire \Tile_X8Y9_FrameData_O[20] ;
 wire \Tile_X8Y9_FrameData_O[21] ;
 wire \Tile_X8Y9_FrameData_O[22] ;
 wire \Tile_X8Y9_FrameData_O[23] ;
 wire \Tile_X8Y9_FrameData_O[24] ;
 wire \Tile_X8Y9_FrameData_O[25] ;
 wire \Tile_X8Y9_FrameData_O[26] ;
 wire \Tile_X8Y9_FrameData_O[27] ;
 wire \Tile_X8Y9_FrameData_O[28] ;
 wire \Tile_X8Y9_FrameData_O[29] ;
 wire \Tile_X8Y9_FrameData_O[2] ;
 wire \Tile_X8Y9_FrameData_O[30] ;
 wire \Tile_X8Y9_FrameData_O[31] ;
 wire \Tile_X8Y9_FrameData_O[3] ;
 wire \Tile_X8Y9_FrameData_O[4] ;
 wire \Tile_X8Y9_FrameData_O[5] ;
 wire \Tile_X8Y9_FrameData_O[6] ;
 wire \Tile_X8Y9_FrameData_O[7] ;
 wire \Tile_X8Y9_FrameData_O[8] ;
 wire \Tile_X8Y9_FrameData_O[9] ;
 wire \Tile_X8Y9_FrameStrobe_O[0] ;
 wire \Tile_X8Y9_FrameStrobe_O[10] ;
 wire \Tile_X8Y9_FrameStrobe_O[11] ;
 wire \Tile_X8Y9_FrameStrobe_O[12] ;
 wire \Tile_X8Y9_FrameStrobe_O[13] ;
 wire \Tile_X8Y9_FrameStrobe_O[14] ;
 wire \Tile_X8Y9_FrameStrobe_O[15] ;
 wire \Tile_X8Y9_FrameStrobe_O[16] ;
 wire \Tile_X8Y9_FrameStrobe_O[17] ;
 wire \Tile_X8Y9_FrameStrobe_O[18] ;
 wire \Tile_X8Y9_FrameStrobe_O[19] ;
 wire \Tile_X8Y9_FrameStrobe_O[1] ;
 wire \Tile_X8Y9_FrameStrobe_O[2] ;
 wire \Tile_X8Y9_FrameStrobe_O[3] ;
 wire \Tile_X8Y9_FrameStrobe_O[4] ;
 wire \Tile_X8Y9_FrameStrobe_O[5] ;
 wire \Tile_X8Y9_FrameStrobe_O[6] ;
 wire \Tile_X8Y9_FrameStrobe_O[7] ;
 wire \Tile_X8Y9_FrameStrobe_O[8] ;
 wire \Tile_X8Y9_FrameStrobe_O[9] ;
 wire \Tile_X8Y9_N1BEG[0] ;
 wire \Tile_X8Y9_N1BEG[1] ;
 wire \Tile_X8Y9_N1BEG[2] ;
 wire \Tile_X8Y9_N1BEG[3] ;
 wire \Tile_X8Y9_N2BEG[0] ;
 wire \Tile_X8Y9_N2BEG[1] ;
 wire \Tile_X8Y9_N2BEG[2] ;
 wire \Tile_X8Y9_N2BEG[3] ;
 wire \Tile_X8Y9_N2BEG[4] ;
 wire \Tile_X8Y9_N2BEG[5] ;
 wire \Tile_X8Y9_N2BEG[6] ;
 wire \Tile_X8Y9_N2BEG[7] ;
 wire \Tile_X8Y9_N2BEGb[0] ;
 wire \Tile_X8Y9_N2BEGb[1] ;
 wire \Tile_X8Y9_N2BEGb[2] ;
 wire \Tile_X8Y9_N2BEGb[3] ;
 wire \Tile_X8Y9_N2BEGb[4] ;
 wire \Tile_X8Y9_N2BEGb[5] ;
 wire \Tile_X8Y9_N2BEGb[6] ;
 wire \Tile_X8Y9_N2BEGb[7] ;
 wire \Tile_X8Y9_N4BEG[0] ;
 wire \Tile_X8Y9_N4BEG[10] ;
 wire \Tile_X8Y9_N4BEG[11] ;
 wire \Tile_X8Y9_N4BEG[12] ;
 wire \Tile_X8Y9_N4BEG[13] ;
 wire \Tile_X8Y9_N4BEG[14] ;
 wire \Tile_X8Y9_N4BEG[15] ;
 wire \Tile_X8Y9_N4BEG[1] ;
 wire \Tile_X8Y9_N4BEG[2] ;
 wire \Tile_X8Y9_N4BEG[3] ;
 wire \Tile_X8Y9_N4BEG[4] ;
 wire \Tile_X8Y9_N4BEG[5] ;
 wire \Tile_X8Y9_N4BEG[6] ;
 wire \Tile_X8Y9_N4BEG[7] ;
 wire \Tile_X8Y9_N4BEG[8] ;
 wire \Tile_X8Y9_N4BEG[9] ;
 wire \Tile_X8Y9_NN4BEG[0] ;
 wire \Tile_X8Y9_NN4BEG[10] ;
 wire \Tile_X8Y9_NN4BEG[11] ;
 wire \Tile_X8Y9_NN4BEG[12] ;
 wire \Tile_X8Y9_NN4BEG[13] ;
 wire \Tile_X8Y9_NN4BEG[14] ;
 wire \Tile_X8Y9_NN4BEG[15] ;
 wire \Tile_X8Y9_NN4BEG[1] ;
 wire \Tile_X8Y9_NN4BEG[2] ;
 wire \Tile_X8Y9_NN4BEG[3] ;
 wire \Tile_X8Y9_NN4BEG[4] ;
 wire \Tile_X8Y9_NN4BEG[5] ;
 wire \Tile_X8Y9_NN4BEG[6] ;
 wire \Tile_X8Y9_NN4BEG[7] ;
 wire \Tile_X8Y9_NN4BEG[8] ;
 wire \Tile_X8Y9_NN4BEG[9] ;
 wire \Tile_X8Y9_S1BEG[0] ;
 wire \Tile_X8Y9_S1BEG[1] ;
 wire \Tile_X8Y9_S1BEG[2] ;
 wire \Tile_X8Y9_S1BEG[3] ;
 wire \Tile_X8Y9_S2BEG[0] ;
 wire \Tile_X8Y9_S2BEG[1] ;
 wire \Tile_X8Y9_S2BEG[2] ;
 wire \Tile_X8Y9_S2BEG[3] ;
 wire \Tile_X8Y9_S2BEG[4] ;
 wire \Tile_X8Y9_S2BEG[5] ;
 wire \Tile_X8Y9_S2BEG[6] ;
 wire \Tile_X8Y9_S2BEG[7] ;
 wire \Tile_X8Y9_S2BEGb[0] ;
 wire \Tile_X8Y9_S2BEGb[1] ;
 wire \Tile_X8Y9_S2BEGb[2] ;
 wire \Tile_X8Y9_S2BEGb[3] ;
 wire \Tile_X8Y9_S2BEGb[4] ;
 wire \Tile_X8Y9_S2BEGb[5] ;
 wire \Tile_X8Y9_S2BEGb[6] ;
 wire \Tile_X8Y9_S2BEGb[7] ;
 wire \Tile_X8Y9_S4BEG[0] ;
 wire \Tile_X8Y9_S4BEG[10] ;
 wire \Tile_X8Y9_S4BEG[11] ;
 wire \Tile_X8Y9_S4BEG[12] ;
 wire \Tile_X8Y9_S4BEG[13] ;
 wire \Tile_X8Y9_S4BEG[14] ;
 wire \Tile_X8Y9_S4BEG[15] ;
 wire \Tile_X8Y9_S4BEG[1] ;
 wire \Tile_X8Y9_S4BEG[2] ;
 wire \Tile_X8Y9_S4BEG[3] ;
 wire \Tile_X8Y9_S4BEG[4] ;
 wire \Tile_X8Y9_S4BEG[5] ;
 wire \Tile_X8Y9_S4BEG[6] ;
 wire \Tile_X8Y9_S4BEG[7] ;
 wire \Tile_X8Y9_S4BEG[8] ;
 wire \Tile_X8Y9_S4BEG[9] ;
 wire \Tile_X8Y9_SS4BEG[0] ;
 wire \Tile_X8Y9_SS4BEG[10] ;
 wire \Tile_X8Y9_SS4BEG[11] ;
 wire \Tile_X8Y9_SS4BEG[12] ;
 wire \Tile_X8Y9_SS4BEG[13] ;
 wire \Tile_X8Y9_SS4BEG[14] ;
 wire \Tile_X8Y9_SS4BEG[15] ;
 wire \Tile_X8Y9_SS4BEG[1] ;
 wire \Tile_X8Y9_SS4BEG[2] ;
 wire \Tile_X8Y9_SS4BEG[3] ;
 wire \Tile_X8Y9_SS4BEG[4] ;
 wire \Tile_X8Y9_SS4BEG[5] ;
 wire \Tile_X8Y9_SS4BEG[6] ;
 wire \Tile_X8Y9_SS4BEG[7] ;
 wire \Tile_X8Y9_SS4BEG[8] ;
 wire \Tile_X8Y9_SS4BEG[9] ;
 wire Tile_X8Y9_UserCLKo;
 wire \Tile_X8Y9_W1BEG[0] ;
 wire \Tile_X8Y9_W1BEG[1] ;
 wire \Tile_X8Y9_W1BEG[2] ;
 wire \Tile_X8Y9_W1BEG[3] ;
 wire \Tile_X8Y9_W2BEG[0] ;
 wire \Tile_X8Y9_W2BEG[1] ;
 wire \Tile_X8Y9_W2BEG[2] ;
 wire \Tile_X8Y9_W2BEG[3] ;
 wire \Tile_X8Y9_W2BEG[4] ;
 wire \Tile_X8Y9_W2BEG[5] ;
 wire \Tile_X8Y9_W2BEG[6] ;
 wire \Tile_X8Y9_W2BEG[7] ;
 wire \Tile_X8Y9_W2BEGb[0] ;
 wire \Tile_X8Y9_W2BEGb[1] ;
 wire \Tile_X8Y9_W2BEGb[2] ;
 wire \Tile_X8Y9_W2BEGb[3] ;
 wire \Tile_X8Y9_W2BEGb[4] ;
 wire \Tile_X8Y9_W2BEGb[5] ;
 wire \Tile_X8Y9_W2BEGb[6] ;
 wire \Tile_X8Y9_W2BEGb[7] ;
 wire \Tile_X8Y9_W6BEG[0] ;
 wire \Tile_X8Y9_W6BEG[10] ;
 wire \Tile_X8Y9_W6BEG[11] ;
 wire \Tile_X8Y9_W6BEG[1] ;
 wire \Tile_X8Y9_W6BEG[2] ;
 wire \Tile_X8Y9_W6BEG[3] ;
 wire \Tile_X8Y9_W6BEG[4] ;
 wire \Tile_X8Y9_W6BEG[5] ;
 wire \Tile_X8Y9_W6BEG[6] ;
 wire \Tile_X8Y9_W6BEG[7] ;
 wire \Tile_X8Y9_W6BEG[8] ;
 wire \Tile_X8Y9_W6BEG[9] ;
 wire \Tile_X8Y9_WW4BEG[0] ;
 wire \Tile_X8Y9_WW4BEG[10] ;
 wire \Tile_X8Y9_WW4BEG[11] ;
 wire \Tile_X8Y9_WW4BEG[12] ;
 wire \Tile_X8Y9_WW4BEG[13] ;
 wire \Tile_X8Y9_WW4BEG[14] ;
 wire \Tile_X8Y9_WW4BEG[15] ;
 wire \Tile_X8Y9_WW4BEG[1] ;
 wire \Tile_X8Y9_WW4BEG[2] ;
 wire \Tile_X8Y9_WW4BEG[3] ;
 wire \Tile_X8Y9_WW4BEG[4] ;
 wire \Tile_X8Y9_WW4BEG[5] ;
 wire \Tile_X8Y9_WW4BEG[6] ;
 wire \Tile_X8Y9_WW4BEG[7] ;
 wire \Tile_X8Y9_WW4BEG[8] ;
 wire \Tile_X8Y9_WW4BEG[9] ;
 wire \Tile_X9Y0_FrameData_O[0] ;
 wire \Tile_X9Y0_FrameData_O[10] ;
 wire \Tile_X9Y0_FrameData_O[11] ;
 wire \Tile_X9Y0_FrameData_O[12] ;
 wire \Tile_X9Y0_FrameData_O[13] ;
 wire \Tile_X9Y0_FrameData_O[14] ;
 wire \Tile_X9Y0_FrameData_O[15] ;
 wire \Tile_X9Y0_FrameData_O[16] ;
 wire \Tile_X9Y0_FrameData_O[17] ;
 wire \Tile_X9Y0_FrameData_O[18] ;
 wire \Tile_X9Y0_FrameData_O[19] ;
 wire \Tile_X9Y0_FrameData_O[1] ;
 wire \Tile_X9Y0_FrameData_O[20] ;
 wire \Tile_X9Y0_FrameData_O[21] ;
 wire \Tile_X9Y0_FrameData_O[22] ;
 wire \Tile_X9Y0_FrameData_O[23] ;
 wire \Tile_X9Y0_FrameData_O[24] ;
 wire \Tile_X9Y0_FrameData_O[25] ;
 wire \Tile_X9Y0_FrameData_O[26] ;
 wire \Tile_X9Y0_FrameData_O[27] ;
 wire \Tile_X9Y0_FrameData_O[28] ;
 wire \Tile_X9Y0_FrameData_O[29] ;
 wire \Tile_X9Y0_FrameData_O[2] ;
 wire \Tile_X9Y0_FrameData_O[30] ;
 wire \Tile_X9Y0_FrameData_O[31] ;
 wire \Tile_X9Y0_FrameData_O[3] ;
 wire \Tile_X9Y0_FrameData_O[4] ;
 wire \Tile_X9Y0_FrameData_O[5] ;
 wire \Tile_X9Y0_FrameData_O[6] ;
 wire \Tile_X9Y0_FrameData_O[7] ;
 wire \Tile_X9Y0_FrameData_O[8] ;
 wire \Tile_X9Y0_FrameData_O[9] ;
 wire \Tile_X9Y0_FrameStrobe_O[0] ;
 wire \Tile_X9Y0_FrameStrobe_O[10] ;
 wire \Tile_X9Y0_FrameStrobe_O[11] ;
 wire \Tile_X9Y0_FrameStrobe_O[12] ;
 wire \Tile_X9Y0_FrameStrobe_O[13] ;
 wire \Tile_X9Y0_FrameStrobe_O[14] ;
 wire \Tile_X9Y0_FrameStrobe_O[15] ;
 wire \Tile_X9Y0_FrameStrobe_O[16] ;
 wire \Tile_X9Y0_FrameStrobe_O[17] ;
 wire \Tile_X9Y0_FrameStrobe_O[18] ;
 wire \Tile_X9Y0_FrameStrobe_O[19] ;
 wire \Tile_X9Y0_FrameStrobe_O[1] ;
 wire \Tile_X9Y0_FrameStrobe_O[2] ;
 wire \Tile_X9Y0_FrameStrobe_O[3] ;
 wire \Tile_X9Y0_FrameStrobe_O[4] ;
 wire \Tile_X9Y0_FrameStrobe_O[5] ;
 wire \Tile_X9Y0_FrameStrobe_O[6] ;
 wire \Tile_X9Y0_FrameStrobe_O[7] ;
 wire \Tile_X9Y0_FrameStrobe_O[8] ;
 wire \Tile_X9Y0_FrameStrobe_O[9] ;
 wire \Tile_X9Y0_S1BEG[0] ;
 wire \Tile_X9Y0_S1BEG[1] ;
 wire \Tile_X9Y0_S1BEG[2] ;
 wire \Tile_X9Y0_S1BEG[3] ;
 wire \Tile_X9Y0_S2BEG[0] ;
 wire \Tile_X9Y0_S2BEG[1] ;
 wire \Tile_X9Y0_S2BEG[2] ;
 wire \Tile_X9Y0_S2BEG[3] ;
 wire \Tile_X9Y0_S2BEG[4] ;
 wire \Tile_X9Y0_S2BEG[5] ;
 wire \Tile_X9Y0_S2BEG[6] ;
 wire \Tile_X9Y0_S2BEG[7] ;
 wire \Tile_X9Y0_S2BEGb[0] ;
 wire \Tile_X9Y0_S2BEGb[1] ;
 wire \Tile_X9Y0_S2BEGb[2] ;
 wire \Tile_X9Y0_S2BEGb[3] ;
 wire \Tile_X9Y0_S2BEGb[4] ;
 wire \Tile_X9Y0_S2BEGb[5] ;
 wire \Tile_X9Y0_S2BEGb[6] ;
 wire \Tile_X9Y0_S2BEGb[7] ;
 wire \Tile_X9Y0_S4BEG[0] ;
 wire \Tile_X9Y0_S4BEG[10] ;
 wire \Tile_X9Y0_S4BEG[11] ;
 wire \Tile_X9Y0_S4BEG[12] ;
 wire \Tile_X9Y0_S4BEG[13] ;
 wire \Tile_X9Y0_S4BEG[14] ;
 wire \Tile_X9Y0_S4BEG[15] ;
 wire \Tile_X9Y0_S4BEG[1] ;
 wire \Tile_X9Y0_S4BEG[2] ;
 wire \Tile_X9Y0_S4BEG[3] ;
 wire \Tile_X9Y0_S4BEG[4] ;
 wire \Tile_X9Y0_S4BEG[5] ;
 wire \Tile_X9Y0_S4BEG[6] ;
 wire \Tile_X9Y0_S4BEG[7] ;
 wire \Tile_X9Y0_S4BEG[8] ;
 wire \Tile_X9Y0_S4BEG[9] ;
 wire \Tile_X9Y0_SS4BEG[0] ;
 wire \Tile_X9Y0_SS4BEG[10] ;
 wire \Tile_X9Y0_SS4BEG[11] ;
 wire \Tile_X9Y0_SS4BEG[12] ;
 wire \Tile_X9Y0_SS4BEG[13] ;
 wire \Tile_X9Y0_SS4BEG[14] ;
 wire \Tile_X9Y0_SS4BEG[15] ;
 wire \Tile_X9Y0_SS4BEG[1] ;
 wire \Tile_X9Y0_SS4BEG[2] ;
 wire \Tile_X9Y0_SS4BEG[3] ;
 wire \Tile_X9Y0_SS4BEG[4] ;
 wire \Tile_X9Y0_SS4BEG[5] ;
 wire \Tile_X9Y0_SS4BEG[6] ;
 wire \Tile_X9Y0_SS4BEG[7] ;
 wire \Tile_X9Y0_SS4BEG[8] ;
 wire \Tile_X9Y0_SS4BEG[9] ;
 wire Tile_X9Y0_UserCLKo;
 wire Tile_X9Y10_Co;
 wire \Tile_X9Y10_E1BEG[0] ;
 wire \Tile_X9Y10_E1BEG[1] ;
 wire \Tile_X9Y10_E1BEG[2] ;
 wire \Tile_X9Y10_E1BEG[3] ;
 wire \Tile_X9Y10_E2BEG[0] ;
 wire \Tile_X9Y10_E2BEG[1] ;
 wire \Tile_X9Y10_E2BEG[2] ;
 wire \Tile_X9Y10_E2BEG[3] ;
 wire \Tile_X9Y10_E2BEG[4] ;
 wire \Tile_X9Y10_E2BEG[5] ;
 wire \Tile_X9Y10_E2BEG[6] ;
 wire \Tile_X9Y10_E2BEG[7] ;
 wire \Tile_X9Y10_E2BEGb[0] ;
 wire \Tile_X9Y10_E2BEGb[1] ;
 wire \Tile_X9Y10_E2BEGb[2] ;
 wire \Tile_X9Y10_E2BEGb[3] ;
 wire \Tile_X9Y10_E2BEGb[4] ;
 wire \Tile_X9Y10_E2BEGb[5] ;
 wire \Tile_X9Y10_E2BEGb[6] ;
 wire \Tile_X9Y10_E2BEGb[7] ;
 wire \Tile_X9Y10_E6BEG[0] ;
 wire \Tile_X9Y10_E6BEG[10] ;
 wire \Tile_X9Y10_E6BEG[11] ;
 wire \Tile_X9Y10_E6BEG[1] ;
 wire \Tile_X9Y10_E6BEG[2] ;
 wire \Tile_X9Y10_E6BEG[3] ;
 wire \Tile_X9Y10_E6BEG[4] ;
 wire \Tile_X9Y10_E6BEG[5] ;
 wire \Tile_X9Y10_E6BEG[6] ;
 wire \Tile_X9Y10_E6BEG[7] ;
 wire \Tile_X9Y10_E6BEG[8] ;
 wire \Tile_X9Y10_E6BEG[9] ;
 wire \Tile_X9Y10_EE4BEG[0] ;
 wire \Tile_X9Y10_EE4BEG[10] ;
 wire \Tile_X9Y10_EE4BEG[11] ;
 wire \Tile_X9Y10_EE4BEG[12] ;
 wire \Tile_X9Y10_EE4BEG[13] ;
 wire \Tile_X9Y10_EE4BEG[14] ;
 wire \Tile_X9Y10_EE4BEG[15] ;
 wire \Tile_X9Y10_EE4BEG[1] ;
 wire \Tile_X9Y10_EE4BEG[2] ;
 wire \Tile_X9Y10_EE4BEG[3] ;
 wire \Tile_X9Y10_EE4BEG[4] ;
 wire \Tile_X9Y10_EE4BEG[5] ;
 wire \Tile_X9Y10_EE4BEG[6] ;
 wire \Tile_X9Y10_EE4BEG[7] ;
 wire \Tile_X9Y10_EE4BEG[8] ;
 wire \Tile_X9Y10_EE4BEG[9] ;
 wire \Tile_X9Y10_FrameData_O[0] ;
 wire \Tile_X9Y10_FrameData_O[10] ;
 wire \Tile_X9Y10_FrameData_O[11] ;
 wire \Tile_X9Y10_FrameData_O[12] ;
 wire \Tile_X9Y10_FrameData_O[13] ;
 wire \Tile_X9Y10_FrameData_O[14] ;
 wire \Tile_X9Y10_FrameData_O[15] ;
 wire \Tile_X9Y10_FrameData_O[16] ;
 wire \Tile_X9Y10_FrameData_O[17] ;
 wire \Tile_X9Y10_FrameData_O[18] ;
 wire \Tile_X9Y10_FrameData_O[19] ;
 wire \Tile_X9Y10_FrameData_O[1] ;
 wire \Tile_X9Y10_FrameData_O[20] ;
 wire \Tile_X9Y10_FrameData_O[21] ;
 wire \Tile_X9Y10_FrameData_O[22] ;
 wire \Tile_X9Y10_FrameData_O[23] ;
 wire \Tile_X9Y10_FrameData_O[24] ;
 wire \Tile_X9Y10_FrameData_O[25] ;
 wire \Tile_X9Y10_FrameData_O[26] ;
 wire \Tile_X9Y10_FrameData_O[27] ;
 wire \Tile_X9Y10_FrameData_O[28] ;
 wire \Tile_X9Y10_FrameData_O[29] ;
 wire \Tile_X9Y10_FrameData_O[2] ;
 wire \Tile_X9Y10_FrameData_O[30] ;
 wire \Tile_X9Y10_FrameData_O[31] ;
 wire \Tile_X9Y10_FrameData_O[3] ;
 wire \Tile_X9Y10_FrameData_O[4] ;
 wire \Tile_X9Y10_FrameData_O[5] ;
 wire \Tile_X9Y10_FrameData_O[6] ;
 wire \Tile_X9Y10_FrameData_O[7] ;
 wire \Tile_X9Y10_FrameData_O[8] ;
 wire \Tile_X9Y10_FrameData_O[9] ;
 wire \Tile_X9Y10_FrameStrobe_O[0] ;
 wire \Tile_X9Y10_FrameStrobe_O[10] ;
 wire \Tile_X9Y10_FrameStrobe_O[11] ;
 wire \Tile_X9Y10_FrameStrobe_O[12] ;
 wire \Tile_X9Y10_FrameStrobe_O[13] ;
 wire \Tile_X9Y10_FrameStrobe_O[14] ;
 wire \Tile_X9Y10_FrameStrobe_O[15] ;
 wire \Tile_X9Y10_FrameStrobe_O[16] ;
 wire \Tile_X9Y10_FrameStrobe_O[17] ;
 wire \Tile_X9Y10_FrameStrobe_O[18] ;
 wire \Tile_X9Y10_FrameStrobe_O[19] ;
 wire \Tile_X9Y10_FrameStrobe_O[1] ;
 wire \Tile_X9Y10_FrameStrobe_O[2] ;
 wire \Tile_X9Y10_FrameStrobe_O[3] ;
 wire \Tile_X9Y10_FrameStrobe_O[4] ;
 wire \Tile_X9Y10_FrameStrobe_O[5] ;
 wire \Tile_X9Y10_FrameStrobe_O[6] ;
 wire \Tile_X9Y10_FrameStrobe_O[7] ;
 wire \Tile_X9Y10_FrameStrobe_O[8] ;
 wire \Tile_X9Y10_FrameStrobe_O[9] ;
 wire \Tile_X9Y10_N1BEG[0] ;
 wire \Tile_X9Y10_N1BEG[1] ;
 wire \Tile_X9Y10_N1BEG[2] ;
 wire \Tile_X9Y10_N1BEG[3] ;
 wire \Tile_X9Y10_N2BEG[0] ;
 wire \Tile_X9Y10_N2BEG[1] ;
 wire \Tile_X9Y10_N2BEG[2] ;
 wire \Tile_X9Y10_N2BEG[3] ;
 wire \Tile_X9Y10_N2BEG[4] ;
 wire \Tile_X9Y10_N2BEG[5] ;
 wire \Tile_X9Y10_N2BEG[6] ;
 wire \Tile_X9Y10_N2BEG[7] ;
 wire \Tile_X9Y10_N2BEGb[0] ;
 wire \Tile_X9Y10_N2BEGb[1] ;
 wire \Tile_X9Y10_N2BEGb[2] ;
 wire \Tile_X9Y10_N2BEGb[3] ;
 wire \Tile_X9Y10_N2BEGb[4] ;
 wire \Tile_X9Y10_N2BEGb[5] ;
 wire \Tile_X9Y10_N2BEGb[6] ;
 wire \Tile_X9Y10_N2BEGb[7] ;
 wire \Tile_X9Y10_N4BEG[0] ;
 wire \Tile_X9Y10_N4BEG[10] ;
 wire \Tile_X9Y10_N4BEG[11] ;
 wire \Tile_X9Y10_N4BEG[12] ;
 wire \Tile_X9Y10_N4BEG[13] ;
 wire \Tile_X9Y10_N4BEG[14] ;
 wire \Tile_X9Y10_N4BEG[15] ;
 wire \Tile_X9Y10_N4BEG[1] ;
 wire \Tile_X9Y10_N4BEG[2] ;
 wire \Tile_X9Y10_N4BEG[3] ;
 wire \Tile_X9Y10_N4BEG[4] ;
 wire \Tile_X9Y10_N4BEG[5] ;
 wire \Tile_X9Y10_N4BEG[6] ;
 wire \Tile_X9Y10_N4BEG[7] ;
 wire \Tile_X9Y10_N4BEG[8] ;
 wire \Tile_X9Y10_N4BEG[9] ;
 wire \Tile_X9Y10_NN4BEG[0] ;
 wire \Tile_X9Y10_NN4BEG[10] ;
 wire \Tile_X9Y10_NN4BEG[11] ;
 wire \Tile_X9Y10_NN4BEG[12] ;
 wire \Tile_X9Y10_NN4BEG[13] ;
 wire \Tile_X9Y10_NN4BEG[14] ;
 wire \Tile_X9Y10_NN4BEG[15] ;
 wire \Tile_X9Y10_NN4BEG[1] ;
 wire \Tile_X9Y10_NN4BEG[2] ;
 wire \Tile_X9Y10_NN4BEG[3] ;
 wire \Tile_X9Y10_NN4BEG[4] ;
 wire \Tile_X9Y10_NN4BEG[5] ;
 wire \Tile_X9Y10_NN4BEG[6] ;
 wire \Tile_X9Y10_NN4BEG[7] ;
 wire \Tile_X9Y10_NN4BEG[8] ;
 wire \Tile_X9Y10_NN4BEG[9] ;
 wire \Tile_X9Y10_S1BEG[0] ;
 wire \Tile_X9Y10_S1BEG[1] ;
 wire \Tile_X9Y10_S1BEG[2] ;
 wire \Tile_X9Y10_S1BEG[3] ;
 wire \Tile_X9Y10_S2BEG[0] ;
 wire \Tile_X9Y10_S2BEG[1] ;
 wire \Tile_X9Y10_S2BEG[2] ;
 wire \Tile_X9Y10_S2BEG[3] ;
 wire \Tile_X9Y10_S2BEG[4] ;
 wire \Tile_X9Y10_S2BEG[5] ;
 wire \Tile_X9Y10_S2BEG[6] ;
 wire \Tile_X9Y10_S2BEG[7] ;
 wire \Tile_X9Y10_S2BEGb[0] ;
 wire \Tile_X9Y10_S2BEGb[1] ;
 wire \Tile_X9Y10_S2BEGb[2] ;
 wire \Tile_X9Y10_S2BEGb[3] ;
 wire \Tile_X9Y10_S2BEGb[4] ;
 wire \Tile_X9Y10_S2BEGb[5] ;
 wire \Tile_X9Y10_S2BEGb[6] ;
 wire \Tile_X9Y10_S2BEGb[7] ;
 wire \Tile_X9Y10_S4BEG[0] ;
 wire \Tile_X9Y10_S4BEG[10] ;
 wire \Tile_X9Y10_S4BEG[11] ;
 wire \Tile_X9Y10_S4BEG[12] ;
 wire \Tile_X9Y10_S4BEG[13] ;
 wire \Tile_X9Y10_S4BEG[14] ;
 wire \Tile_X9Y10_S4BEG[15] ;
 wire \Tile_X9Y10_S4BEG[1] ;
 wire \Tile_X9Y10_S4BEG[2] ;
 wire \Tile_X9Y10_S4BEG[3] ;
 wire \Tile_X9Y10_S4BEG[4] ;
 wire \Tile_X9Y10_S4BEG[5] ;
 wire \Tile_X9Y10_S4BEG[6] ;
 wire \Tile_X9Y10_S4BEG[7] ;
 wire \Tile_X9Y10_S4BEG[8] ;
 wire \Tile_X9Y10_S4BEG[9] ;
 wire \Tile_X9Y10_SS4BEG[0] ;
 wire \Tile_X9Y10_SS4BEG[10] ;
 wire \Tile_X9Y10_SS4BEG[11] ;
 wire \Tile_X9Y10_SS4BEG[12] ;
 wire \Tile_X9Y10_SS4BEG[13] ;
 wire \Tile_X9Y10_SS4BEG[14] ;
 wire \Tile_X9Y10_SS4BEG[15] ;
 wire \Tile_X9Y10_SS4BEG[1] ;
 wire \Tile_X9Y10_SS4BEG[2] ;
 wire \Tile_X9Y10_SS4BEG[3] ;
 wire \Tile_X9Y10_SS4BEG[4] ;
 wire \Tile_X9Y10_SS4BEG[5] ;
 wire \Tile_X9Y10_SS4BEG[6] ;
 wire \Tile_X9Y10_SS4BEG[7] ;
 wire \Tile_X9Y10_SS4BEG[8] ;
 wire \Tile_X9Y10_SS4BEG[9] ;
 wire Tile_X9Y10_UserCLKo;
 wire \Tile_X9Y10_W1BEG[0] ;
 wire \Tile_X9Y10_W1BEG[1] ;
 wire \Tile_X9Y10_W1BEG[2] ;
 wire \Tile_X9Y10_W1BEG[3] ;
 wire \Tile_X9Y10_W2BEG[0] ;
 wire \Tile_X9Y10_W2BEG[1] ;
 wire \Tile_X9Y10_W2BEG[2] ;
 wire \Tile_X9Y10_W2BEG[3] ;
 wire \Tile_X9Y10_W2BEG[4] ;
 wire \Tile_X9Y10_W2BEG[5] ;
 wire \Tile_X9Y10_W2BEG[6] ;
 wire \Tile_X9Y10_W2BEG[7] ;
 wire \Tile_X9Y10_W2BEGb[0] ;
 wire \Tile_X9Y10_W2BEGb[1] ;
 wire \Tile_X9Y10_W2BEGb[2] ;
 wire \Tile_X9Y10_W2BEGb[3] ;
 wire \Tile_X9Y10_W2BEGb[4] ;
 wire \Tile_X9Y10_W2BEGb[5] ;
 wire \Tile_X9Y10_W2BEGb[6] ;
 wire \Tile_X9Y10_W2BEGb[7] ;
 wire \Tile_X9Y10_W6BEG[0] ;
 wire \Tile_X9Y10_W6BEG[10] ;
 wire \Tile_X9Y10_W6BEG[11] ;
 wire \Tile_X9Y10_W6BEG[1] ;
 wire \Tile_X9Y10_W6BEG[2] ;
 wire \Tile_X9Y10_W6BEG[3] ;
 wire \Tile_X9Y10_W6BEG[4] ;
 wire \Tile_X9Y10_W6BEG[5] ;
 wire \Tile_X9Y10_W6BEG[6] ;
 wire \Tile_X9Y10_W6BEG[7] ;
 wire \Tile_X9Y10_W6BEG[8] ;
 wire \Tile_X9Y10_W6BEG[9] ;
 wire \Tile_X9Y10_WW4BEG[0] ;
 wire \Tile_X9Y10_WW4BEG[10] ;
 wire \Tile_X9Y10_WW4BEG[11] ;
 wire \Tile_X9Y10_WW4BEG[12] ;
 wire \Tile_X9Y10_WW4BEG[13] ;
 wire \Tile_X9Y10_WW4BEG[14] ;
 wire \Tile_X9Y10_WW4BEG[15] ;
 wire \Tile_X9Y10_WW4BEG[1] ;
 wire \Tile_X9Y10_WW4BEG[2] ;
 wire \Tile_X9Y10_WW4BEG[3] ;
 wire \Tile_X9Y10_WW4BEG[4] ;
 wire \Tile_X9Y10_WW4BEG[5] ;
 wire \Tile_X9Y10_WW4BEG[6] ;
 wire \Tile_X9Y10_WW4BEG[7] ;
 wire \Tile_X9Y10_WW4BEG[8] ;
 wire \Tile_X9Y10_WW4BEG[9] ;
 wire Tile_X9Y11_Co;
 wire \Tile_X9Y11_E1BEG[0] ;
 wire \Tile_X9Y11_E1BEG[1] ;
 wire \Tile_X9Y11_E1BEG[2] ;
 wire \Tile_X9Y11_E1BEG[3] ;
 wire \Tile_X9Y11_E2BEG[0] ;
 wire \Tile_X9Y11_E2BEG[1] ;
 wire \Tile_X9Y11_E2BEG[2] ;
 wire \Tile_X9Y11_E2BEG[3] ;
 wire \Tile_X9Y11_E2BEG[4] ;
 wire \Tile_X9Y11_E2BEG[5] ;
 wire \Tile_X9Y11_E2BEG[6] ;
 wire \Tile_X9Y11_E2BEG[7] ;
 wire \Tile_X9Y11_E2BEGb[0] ;
 wire \Tile_X9Y11_E2BEGb[1] ;
 wire \Tile_X9Y11_E2BEGb[2] ;
 wire \Tile_X9Y11_E2BEGb[3] ;
 wire \Tile_X9Y11_E2BEGb[4] ;
 wire \Tile_X9Y11_E2BEGb[5] ;
 wire \Tile_X9Y11_E2BEGb[6] ;
 wire \Tile_X9Y11_E2BEGb[7] ;
 wire \Tile_X9Y11_E6BEG[0] ;
 wire \Tile_X9Y11_E6BEG[10] ;
 wire \Tile_X9Y11_E6BEG[11] ;
 wire \Tile_X9Y11_E6BEG[1] ;
 wire \Tile_X9Y11_E6BEG[2] ;
 wire \Tile_X9Y11_E6BEG[3] ;
 wire \Tile_X9Y11_E6BEG[4] ;
 wire \Tile_X9Y11_E6BEG[5] ;
 wire \Tile_X9Y11_E6BEG[6] ;
 wire \Tile_X9Y11_E6BEG[7] ;
 wire \Tile_X9Y11_E6BEG[8] ;
 wire \Tile_X9Y11_E6BEG[9] ;
 wire \Tile_X9Y11_EE4BEG[0] ;
 wire \Tile_X9Y11_EE4BEG[10] ;
 wire \Tile_X9Y11_EE4BEG[11] ;
 wire \Tile_X9Y11_EE4BEG[12] ;
 wire \Tile_X9Y11_EE4BEG[13] ;
 wire \Tile_X9Y11_EE4BEG[14] ;
 wire \Tile_X9Y11_EE4BEG[15] ;
 wire \Tile_X9Y11_EE4BEG[1] ;
 wire \Tile_X9Y11_EE4BEG[2] ;
 wire \Tile_X9Y11_EE4BEG[3] ;
 wire \Tile_X9Y11_EE4BEG[4] ;
 wire \Tile_X9Y11_EE4BEG[5] ;
 wire \Tile_X9Y11_EE4BEG[6] ;
 wire \Tile_X9Y11_EE4BEG[7] ;
 wire \Tile_X9Y11_EE4BEG[8] ;
 wire \Tile_X9Y11_EE4BEG[9] ;
 wire \Tile_X9Y11_FrameData_O[0] ;
 wire \Tile_X9Y11_FrameData_O[10] ;
 wire \Tile_X9Y11_FrameData_O[11] ;
 wire \Tile_X9Y11_FrameData_O[12] ;
 wire \Tile_X9Y11_FrameData_O[13] ;
 wire \Tile_X9Y11_FrameData_O[14] ;
 wire \Tile_X9Y11_FrameData_O[15] ;
 wire \Tile_X9Y11_FrameData_O[16] ;
 wire \Tile_X9Y11_FrameData_O[17] ;
 wire \Tile_X9Y11_FrameData_O[18] ;
 wire \Tile_X9Y11_FrameData_O[19] ;
 wire \Tile_X9Y11_FrameData_O[1] ;
 wire \Tile_X9Y11_FrameData_O[20] ;
 wire \Tile_X9Y11_FrameData_O[21] ;
 wire \Tile_X9Y11_FrameData_O[22] ;
 wire \Tile_X9Y11_FrameData_O[23] ;
 wire \Tile_X9Y11_FrameData_O[24] ;
 wire \Tile_X9Y11_FrameData_O[25] ;
 wire \Tile_X9Y11_FrameData_O[26] ;
 wire \Tile_X9Y11_FrameData_O[27] ;
 wire \Tile_X9Y11_FrameData_O[28] ;
 wire \Tile_X9Y11_FrameData_O[29] ;
 wire \Tile_X9Y11_FrameData_O[2] ;
 wire \Tile_X9Y11_FrameData_O[30] ;
 wire \Tile_X9Y11_FrameData_O[31] ;
 wire \Tile_X9Y11_FrameData_O[3] ;
 wire \Tile_X9Y11_FrameData_O[4] ;
 wire \Tile_X9Y11_FrameData_O[5] ;
 wire \Tile_X9Y11_FrameData_O[6] ;
 wire \Tile_X9Y11_FrameData_O[7] ;
 wire \Tile_X9Y11_FrameData_O[8] ;
 wire \Tile_X9Y11_FrameData_O[9] ;
 wire \Tile_X9Y11_FrameStrobe_O[0] ;
 wire \Tile_X9Y11_FrameStrobe_O[10] ;
 wire \Tile_X9Y11_FrameStrobe_O[11] ;
 wire \Tile_X9Y11_FrameStrobe_O[12] ;
 wire \Tile_X9Y11_FrameStrobe_O[13] ;
 wire \Tile_X9Y11_FrameStrobe_O[14] ;
 wire \Tile_X9Y11_FrameStrobe_O[15] ;
 wire \Tile_X9Y11_FrameStrobe_O[16] ;
 wire \Tile_X9Y11_FrameStrobe_O[17] ;
 wire \Tile_X9Y11_FrameStrobe_O[18] ;
 wire \Tile_X9Y11_FrameStrobe_O[19] ;
 wire \Tile_X9Y11_FrameStrobe_O[1] ;
 wire \Tile_X9Y11_FrameStrobe_O[2] ;
 wire \Tile_X9Y11_FrameStrobe_O[3] ;
 wire \Tile_X9Y11_FrameStrobe_O[4] ;
 wire \Tile_X9Y11_FrameStrobe_O[5] ;
 wire \Tile_X9Y11_FrameStrobe_O[6] ;
 wire \Tile_X9Y11_FrameStrobe_O[7] ;
 wire \Tile_X9Y11_FrameStrobe_O[8] ;
 wire \Tile_X9Y11_FrameStrobe_O[9] ;
 wire \Tile_X9Y11_N1BEG[0] ;
 wire \Tile_X9Y11_N1BEG[1] ;
 wire \Tile_X9Y11_N1BEG[2] ;
 wire \Tile_X9Y11_N1BEG[3] ;
 wire \Tile_X9Y11_N2BEG[0] ;
 wire \Tile_X9Y11_N2BEG[1] ;
 wire \Tile_X9Y11_N2BEG[2] ;
 wire \Tile_X9Y11_N2BEG[3] ;
 wire \Tile_X9Y11_N2BEG[4] ;
 wire \Tile_X9Y11_N2BEG[5] ;
 wire \Tile_X9Y11_N2BEG[6] ;
 wire \Tile_X9Y11_N2BEG[7] ;
 wire \Tile_X9Y11_N2BEGb[0] ;
 wire \Tile_X9Y11_N2BEGb[1] ;
 wire \Tile_X9Y11_N2BEGb[2] ;
 wire \Tile_X9Y11_N2BEGb[3] ;
 wire \Tile_X9Y11_N2BEGb[4] ;
 wire \Tile_X9Y11_N2BEGb[5] ;
 wire \Tile_X9Y11_N2BEGb[6] ;
 wire \Tile_X9Y11_N2BEGb[7] ;
 wire \Tile_X9Y11_N4BEG[0] ;
 wire \Tile_X9Y11_N4BEG[10] ;
 wire \Tile_X9Y11_N4BEG[11] ;
 wire \Tile_X9Y11_N4BEG[12] ;
 wire \Tile_X9Y11_N4BEG[13] ;
 wire \Tile_X9Y11_N4BEG[14] ;
 wire \Tile_X9Y11_N4BEG[15] ;
 wire \Tile_X9Y11_N4BEG[1] ;
 wire \Tile_X9Y11_N4BEG[2] ;
 wire \Tile_X9Y11_N4BEG[3] ;
 wire \Tile_X9Y11_N4BEG[4] ;
 wire \Tile_X9Y11_N4BEG[5] ;
 wire \Tile_X9Y11_N4BEG[6] ;
 wire \Tile_X9Y11_N4BEG[7] ;
 wire \Tile_X9Y11_N4BEG[8] ;
 wire \Tile_X9Y11_N4BEG[9] ;
 wire \Tile_X9Y11_NN4BEG[0] ;
 wire \Tile_X9Y11_NN4BEG[10] ;
 wire \Tile_X9Y11_NN4BEG[11] ;
 wire \Tile_X9Y11_NN4BEG[12] ;
 wire \Tile_X9Y11_NN4BEG[13] ;
 wire \Tile_X9Y11_NN4BEG[14] ;
 wire \Tile_X9Y11_NN4BEG[15] ;
 wire \Tile_X9Y11_NN4BEG[1] ;
 wire \Tile_X9Y11_NN4BEG[2] ;
 wire \Tile_X9Y11_NN4BEG[3] ;
 wire \Tile_X9Y11_NN4BEG[4] ;
 wire \Tile_X9Y11_NN4BEG[5] ;
 wire \Tile_X9Y11_NN4BEG[6] ;
 wire \Tile_X9Y11_NN4BEG[7] ;
 wire \Tile_X9Y11_NN4BEG[8] ;
 wire \Tile_X9Y11_NN4BEG[9] ;
 wire \Tile_X9Y11_S1BEG[0] ;
 wire \Tile_X9Y11_S1BEG[1] ;
 wire \Tile_X9Y11_S1BEG[2] ;
 wire \Tile_X9Y11_S1BEG[3] ;
 wire \Tile_X9Y11_S2BEG[0] ;
 wire \Tile_X9Y11_S2BEG[1] ;
 wire \Tile_X9Y11_S2BEG[2] ;
 wire \Tile_X9Y11_S2BEG[3] ;
 wire \Tile_X9Y11_S2BEG[4] ;
 wire \Tile_X9Y11_S2BEG[5] ;
 wire \Tile_X9Y11_S2BEG[6] ;
 wire \Tile_X9Y11_S2BEG[7] ;
 wire \Tile_X9Y11_S2BEGb[0] ;
 wire \Tile_X9Y11_S2BEGb[1] ;
 wire \Tile_X9Y11_S2BEGb[2] ;
 wire \Tile_X9Y11_S2BEGb[3] ;
 wire \Tile_X9Y11_S2BEGb[4] ;
 wire \Tile_X9Y11_S2BEGb[5] ;
 wire \Tile_X9Y11_S2BEGb[6] ;
 wire \Tile_X9Y11_S2BEGb[7] ;
 wire \Tile_X9Y11_S4BEG[0] ;
 wire \Tile_X9Y11_S4BEG[10] ;
 wire \Tile_X9Y11_S4BEG[11] ;
 wire \Tile_X9Y11_S4BEG[12] ;
 wire \Tile_X9Y11_S4BEG[13] ;
 wire \Tile_X9Y11_S4BEG[14] ;
 wire \Tile_X9Y11_S4BEG[15] ;
 wire \Tile_X9Y11_S4BEG[1] ;
 wire \Tile_X9Y11_S4BEG[2] ;
 wire \Tile_X9Y11_S4BEG[3] ;
 wire \Tile_X9Y11_S4BEG[4] ;
 wire \Tile_X9Y11_S4BEG[5] ;
 wire \Tile_X9Y11_S4BEG[6] ;
 wire \Tile_X9Y11_S4BEG[7] ;
 wire \Tile_X9Y11_S4BEG[8] ;
 wire \Tile_X9Y11_S4BEG[9] ;
 wire \Tile_X9Y11_SS4BEG[0] ;
 wire \Tile_X9Y11_SS4BEG[10] ;
 wire \Tile_X9Y11_SS4BEG[11] ;
 wire \Tile_X9Y11_SS4BEG[12] ;
 wire \Tile_X9Y11_SS4BEG[13] ;
 wire \Tile_X9Y11_SS4BEG[14] ;
 wire \Tile_X9Y11_SS4BEG[15] ;
 wire \Tile_X9Y11_SS4BEG[1] ;
 wire \Tile_X9Y11_SS4BEG[2] ;
 wire \Tile_X9Y11_SS4BEG[3] ;
 wire \Tile_X9Y11_SS4BEG[4] ;
 wire \Tile_X9Y11_SS4BEG[5] ;
 wire \Tile_X9Y11_SS4BEG[6] ;
 wire \Tile_X9Y11_SS4BEG[7] ;
 wire \Tile_X9Y11_SS4BEG[8] ;
 wire \Tile_X9Y11_SS4BEG[9] ;
 wire Tile_X9Y11_UserCLKo;
 wire \Tile_X9Y11_W1BEG[0] ;
 wire \Tile_X9Y11_W1BEG[1] ;
 wire \Tile_X9Y11_W1BEG[2] ;
 wire \Tile_X9Y11_W1BEG[3] ;
 wire \Tile_X9Y11_W2BEG[0] ;
 wire \Tile_X9Y11_W2BEG[1] ;
 wire \Tile_X9Y11_W2BEG[2] ;
 wire \Tile_X9Y11_W2BEG[3] ;
 wire \Tile_X9Y11_W2BEG[4] ;
 wire \Tile_X9Y11_W2BEG[5] ;
 wire \Tile_X9Y11_W2BEG[6] ;
 wire \Tile_X9Y11_W2BEG[7] ;
 wire \Tile_X9Y11_W2BEGb[0] ;
 wire \Tile_X9Y11_W2BEGb[1] ;
 wire \Tile_X9Y11_W2BEGb[2] ;
 wire \Tile_X9Y11_W2BEGb[3] ;
 wire \Tile_X9Y11_W2BEGb[4] ;
 wire \Tile_X9Y11_W2BEGb[5] ;
 wire \Tile_X9Y11_W2BEGb[6] ;
 wire \Tile_X9Y11_W2BEGb[7] ;
 wire \Tile_X9Y11_W6BEG[0] ;
 wire \Tile_X9Y11_W6BEG[10] ;
 wire \Tile_X9Y11_W6BEG[11] ;
 wire \Tile_X9Y11_W6BEG[1] ;
 wire \Tile_X9Y11_W6BEG[2] ;
 wire \Tile_X9Y11_W6BEG[3] ;
 wire \Tile_X9Y11_W6BEG[4] ;
 wire \Tile_X9Y11_W6BEG[5] ;
 wire \Tile_X9Y11_W6BEG[6] ;
 wire \Tile_X9Y11_W6BEG[7] ;
 wire \Tile_X9Y11_W6BEG[8] ;
 wire \Tile_X9Y11_W6BEG[9] ;
 wire \Tile_X9Y11_WW4BEG[0] ;
 wire \Tile_X9Y11_WW4BEG[10] ;
 wire \Tile_X9Y11_WW4BEG[11] ;
 wire \Tile_X9Y11_WW4BEG[12] ;
 wire \Tile_X9Y11_WW4BEG[13] ;
 wire \Tile_X9Y11_WW4BEG[14] ;
 wire \Tile_X9Y11_WW4BEG[15] ;
 wire \Tile_X9Y11_WW4BEG[1] ;
 wire \Tile_X9Y11_WW4BEG[2] ;
 wire \Tile_X9Y11_WW4BEG[3] ;
 wire \Tile_X9Y11_WW4BEG[4] ;
 wire \Tile_X9Y11_WW4BEG[5] ;
 wire \Tile_X9Y11_WW4BEG[6] ;
 wire \Tile_X9Y11_WW4BEG[7] ;
 wire \Tile_X9Y11_WW4BEG[8] ;
 wire \Tile_X9Y11_WW4BEG[9] ;
 wire Tile_X9Y12_Co;
 wire \Tile_X9Y12_E1BEG[0] ;
 wire \Tile_X9Y12_E1BEG[1] ;
 wire \Tile_X9Y12_E1BEG[2] ;
 wire \Tile_X9Y12_E1BEG[3] ;
 wire \Tile_X9Y12_E2BEG[0] ;
 wire \Tile_X9Y12_E2BEG[1] ;
 wire \Tile_X9Y12_E2BEG[2] ;
 wire \Tile_X9Y12_E2BEG[3] ;
 wire \Tile_X9Y12_E2BEG[4] ;
 wire \Tile_X9Y12_E2BEG[5] ;
 wire \Tile_X9Y12_E2BEG[6] ;
 wire \Tile_X9Y12_E2BEG[7] ;
 wire \Tile_X9Y12_E2BEGb[0] ;
 wire \Tile_X9Y12_E2BEGb[1] ;
 wire \Tile_X9Y12_E2BEGb[2] ;
 wire \Tile_X9Y12_E2BEGb[3] ;
 wire \Tile_X9Y12_E2BEGb[4] ;
 wire \Tile_X9Y12_E2BEGb[5] ;
 wire \Tile_X9Y12_E2BEGb[6] ;
 wire \Tile_X9Y12_E2BEGb[7] ;
 wire \Tile_X9Y12_E6BEG[0] ;
 wire \Tile_X9Y12_E6BEG[10] ;
 wire \Tile_X9Y12_E6BEG[11] ;
 wire \Tile_X9Y12_E6BEG[1] ;
 wire \Tile_X9Y12_E6BEG[2] ;
 wire \Tile_X9Y12_E6BEG[3] ;
 wire \Tile_X9Y12_E6BEG[4] ;
 wire \Tile_X9Y12_E6BEG[5] ;
 wire \Tile_X9Y12_E6BEG[6] ;
 wire \Tile_X9Y12_E6BEG[7] ;
 wire \Tile_X9Y12_E6BEG[8] ;
 wire \Tile_X9Y12_E6BEG[9] ;
 wire \Tile_X9Y12_EE4BEG[0] ;
 wire \Tile_X9Y12_EE4BEG[10] ;
 wire \Tile_X9Y12_EE4BEG[11] ;
 wire \Tile_X9Y12_EE4BEG[12] ;
 wire \Tile_X9Y12_EE4BEG[13] ;
 wire \Tile_X9Y12_EE4BEG[14] ;
 wire \Tile_X9Y12_EE4BEG[15] ;
 wire \Tile_X9Y12_EE4BEG[1] ;
 wire \Tile_X9Y12_EE4BEG[2] ;
 wire \Tile_X9Y12_EE4BEG[3] ;
 wire \Tile_X9Y12_EE4BEG[4] ;
 wire \Tile_X9Y12_EE4BEG[5] ;
 wire \Tile_X9Y12_EE4BEG[6] ;
 wire \Tile_X9Y12_EE4BEG[7] ;
 wire \Tile_X9Y12_EE4BEG[8] ;
 wire \Tile_X9Y12_EE4BEG[9] ;
 wire \Tile_X9Y12_FrameData_O[0] ;
 wire \Tile_X9Y12_FrameData_O[10] ;
 wire \Tile_X9Y12_FrameData_O[11] ;
 wire \Tile_X9Y12_FrameData_O[12] ;
 wire \Tile_X9Y12_FrameData_O[13] ;
 wire \Tile_X9Y12_FrameData_O[14] ;
 wire \Tile_X9Y12_FrameData_O[15] ;
 wire \Tile_X9Y12_FrameData_O[16] ;
 wire \Tile_X9Y12_FrameData_O[17] ;
 wire \Tile_X9Y12_FrameData_O[18] ;
 wire \Tile_X9Y12_FrameData_O[19] ;
 wire \Tile_X9Y12_FrameData_O[1] ;
 wire \Tile_X9Y12_FrameData_O[20] ;
 wire \Tile_X9Y12_FrameData_O[21] ;
 wire \Tile_X9Y12_FrameData_O[22] ;
 wire \Tile_X9Y12_FrameData_O[23] ;
 wire \Tile_X9Y12_FrameData_O[24] ;
 wire \Tile_X9Y12_FrameData_O[25] ;
 wire \Tile_X9Y12_FrameData_O[26] ;
 wire \Tile_X9Y12_FrameData_O[27] ;
 wire \Tile_X9Y12_FrameData_O[28] ;
 wire \Tile_X9Y12_FrameData_O[29] ;
 wire \Tile_X9Y12_FrameData_O[2] ;
 wire \Tile_X9Y12_FrameData_O[30] ;
 wire \Tile_X9Y12_FrameData_O[31] ;
 wire \Tile_X9Y12_FrameData_O[3] ;
 wire \Tile_X9Y12_FrameData_O[4] ;
 wire \Tile_X9Y12_FrameData_O[5] ;
 wire \Tile_X9Y12_FrameData_O[6] ;
 wire \Tile_X9Y12_FrameData_O[7] ;
 wire \Tile_X9Y12_FrameData_O[8] ;
 wire \Tile_X9Y12_FrameData_O[9] ;
 wire \Tile_X9Y12_FrameStrobe_O[0] ;
 wire \Tile_X9Y12_FrameStrobe_O[10] ;
 wire \Tile_X9Y12_FrameStrobe_O[11] ;
 wire \Tile_X9Y12_FrameStrobe_O[12] ;
 wire \Tile_X9Y12_FrameStrobe_O[13] ;
 wire \Tile_X9Y12_FrameStrobe_O[14] ;
 wire \Tile_X9Y12_FrameStrobe_O[15] ;
 wire \Tile_X9Y12_FrameStrobe_O[16] ;
 wire \Tile_X9Y12_FrameStrobe_O[17] ;
 wire \Tile_X9Y12_FrameStrobe_O[18] ;
 wire \Tile_X9Y12_FrameStrobe_O[19] ;
 wire \Tile_X9Y12_FrameStrobe_O[1] ;
 wire \Tile_X9Y12_FrameStrobe_O[2] ;
 wire \Tile_X9Y12_FrameStrobe_O[3] ;
 wire \Tile_X9Y12_FrameStrobe_O[4] ;
 wire \Tile_X9Y12_FrameStrobe_O[5] ;
 wire \Tile_X9Y12_FrameStrobe_O[6] ;
 wire \Tile_X9Y12_FrameStrobe_O[7] ;
 wire \Tile_X9Y12_FrameStrobe_O[8] ;
 wire \Tile_X9Y12_FrameStrobe_O[9] ;
 wire \Tile_X9Y12_N1BEG[0] ;
 wire \Tile_X9Y12_N1BEG[1] ;
 wire \Tile_X9Y12_N1BEG[2] ;
 wire \Tile_X9Y12_N1BEG[3] ;
 wire \Tile_X9Y12_N2BEG[0] ;
 wire \Tile_X9Y12_N2BEG[1] ;
 wire \Tile_X9Y12_N2BEG[2] ;
 wire \Tile_X9Y12_N2BEG[3] ;
 wire \Tile_X9Y12_N2BEG[4] ;
 wire \Tile_X9Y12_N2BEG[5] ;
 wire \Tile_X9Y12_N2BEG[6] ;
 wire \Tile_X9Y12_N2BEG[7] ;
 wire \Tile_X9Y12_N2BEGb[0] ;
 wire \Tile_X9Y12_N2BEGb[1] ;
 wire \Tile_X9Y12_N2BEGb[2] ;
 wire \Tile_X9Y12_N2BEGb[3] ;
 wire \Tile_X9Y12_N2BEGb[4] ;
 wire \Tile_X9Y12_N2BEGb[5] ;
 wire \Tile_X9Y12_N2BEGb[6] ;
 wire \Tile_X9Y12_N2BEGb[7] ;
 wire \Tile_X9Y12_N4BEG[0] ;
 wire \Tile_X9Y12_N4BEG[10] ;
 wire \Tile_X9Y12_N4BEG[11] ;
 wire \Tile_X9Y12_N4BEG[12] ;
 wire \Tile_X9Y12_N4BEG[13] ;
 wire \Tile_X9Y12_N4BEG[14] ;
 wire \Tile_X9Y12_N4BEG[15] ;
 wire \Tile_X9Y12_N4BEG[1] ;
 wire \Tile_X9Y12_N4BEG[2] ;
 wire \Tile_X9Y12_N4BEG[3] ;
 wire \Tile_X9Y12_N4BEG[4] ;
 wire \Tile_X9Y12_N4BEG[5] ;
 wire \Tile_X9Y12_N4BEG[6] ;
 wire \Tile_X9Y12_N4BEG[7] ;
 wire \Tile_X9Y12_N4BEG[8] ;
 wire \Tile_X9Y12_N4BEG[9] ;
 wire \Tile_X9Y12_NN4BEG[0] ;
 wire \Tile_X9Y12_NN4BEG[10] ;
 wire \Tile_X9Y12_NN4BEG[11] ;
 wire \Tile_X9Y12_NN4BEG[12] ;
 wire \Tile_X9Y12_NN4BEG[13] ;
 wire \Tile_X9Y12_NN4BEG[14] ;
 wire \Tile_X9Y12_NN4BEG[15] ;
 wire \Tile_X9Y12_NN4BEG[1] ;
 wire \Tile_X9Y12_NN4BEG[2] ;
 wire \Tile_X9Y12_NN4BEG[3] ;
 wire \Tile_X9Y12_NN4BEG[4] ;
 wire \Tile_X9Y12_NN4BEG[5] ;
 wire \Tile_X9Y12_NN4BEG[6] ;
 wire \Tile_X9Y12_NN4BEG[7] ;
 wire \Tile_X9Y12_NN4BEG[8] ;
 wire \Tile_X9Y12_NN4BEG[9] ;
 wire \Tile_X9Y12_S1BEG[0] ;
 wire \Tile_X9Y12_S1BEG[1] ;
 wire \Tile_X9Y12_S1BEG[2] ;
 wire \Tile_X9Y12_S1BEG[3] ;
 wire \Tile_X9Y12_S2BEG[0] ;
 wire \Tile_X9Y12_S2BEG[1] ;
 wire \Tile_X9Y12_S2BEG[2] ;
 wire \Tile_X9Y12_S2BEG[3] ;
 wire \Tile_X9Y12_S2BEG[4] ;
 wire \Tile_X9Y12_S2BEG[5] ;
 wire \Tile_X9Y12_S2BEG[6] ;
 wire \Tile_X9Y12_S2BEG[7] ;
 wire \Tile_X9Y12_S2BEGb[0] ;
 wire \Tile_X9Y12_S2BEGb[1] ;
 wire \Tile_X9Y12_S2BEGb[2] ;
 wire \Tile_X9Y12_S2BEGb[3] ;
 wire \Tile_X9Y12_S2BEGb[4] ;
 wire \Tile_X9Y12_S2BEGb[5] ;
 wire \Tile_X9Y12_S2BEGb[6] ;
 wire \Tile_X9Y12_S2BEGb[7] ;
 wire \Tile_X9Y12_S4BEG[0] ;
 wire \Tile_X9Y12_S4BEG[10] ;
 wire \Tile_X9Y12_S4BEG[11] ;
 wire \Tile_X9Y12_S4BEG[12] ;
 wire \Tile_X9Y12_S4BEG[13] ;
 wire \Tile_X9Y12_S4BEG[14] ;
 wire \Tile_X9Y12_S4BEG[15] ;
 wire \Tile_X9Y12_S4BEG[1] ;
 wire \Tile_X9Y12_S4BEG[2] ;
 wire \Tile_X9Y12_S4BEG[3] ;
 wire \Tile_X9Y12_S4BEG[4] ;
 wire \Tile_X9Y12_S4BEG[5] ;
 wire \Tile_X9Y12_S4BEG[6] ;
 wire \Tile_X9Y12_S4BEG[7] ;
 wire \Tile_X9Y12_S4BEG[8] ;
 wire \Tile_X9Y12_S4BEG[9] ;
 wire \Tile_X9Y12_SS4BEG[0] ;
 wire \Tile_X9Y12_SS4BEG[10] ;
 wire \Tile_X9Y12_SS4BEG[11] ;
 wire \Tile_X9Y12_SS4BEG[12] ;
 wire \Tile_X9Y12_SS4BEG[13] ;
 wire \Tile_X9Y12_SS4BEG[14] ;
 wire \Tile_X9Y12_SS4BEG[15] ;
 wire \Tile_X9Y12_SS4BEG[1] ;
 wire \Tile_X9Y12_SS4BEG[2] ;
 wire \Tile_X9Y12_SS4BEG[3] ;
 wire \Tile_X9Y12_SS4BEG[4] ;
 wire \Tile_X9Y12_SS4BEG[5] ;
 wire \Tile_X9Y12_SS4BEG[6] ;
 wire \Tile_X9Y12_SS4BEG[7] ;
 wire \Tile_X9Y12_SS4BEG[8] ;
 wire \Tile_X9Y12_SS4BEG[9] ;
 wire Tile_X9Y12_UserCLKo;
 wire \Tile_X9Y12_W1BEG[0] ;
 wire \Tile_X9Y12_W1BEG[1] ;
 wire \Tile_X9Y12_W1BEG[2] ;
 wire \Tile_X9Y12_W1BEG[3] ;
 wire \Tile_X9Y12_W2BEG[0] ;
 wire \Tile_X9Y12_W2BEG[1] ;
 wire \Tile_X9Y12_W2BEG[2] ;
 wire \Tile_X9Y12_W2BEG[3] ;
 wire \Tile_X9Y12_W2BEG[4] ;
 wire \Tile_X9Y12_W2BEG[5] ;
 wire \Tile_X9Y12_W2BEG[6] ;
 wire \Tile_X9Y12_W2BEG[7] ;
 wire \Tile_X9Y12_W2BEGb[0] ;
 wire \Tile_X9Y12_W2BEGb[1] ;
 wire \Tile_X9Y12_W2BEGb[2] ;
 wire \Tile_X9Y12_W2BEGb[3] ;
 wire \Tile_X9Y12_W2BEGb[4] ;
 wire \Tile_X9Y12_W2BEGb[5] ;
 wire \Tile_X9Y12_W2BEGb[6] ;
 wire \Tile_X9Y12_W2BEGb[7] ;
 wire \Tile_X9Y12_W6BEG[0] ;
 wire \Tile_X9Y12_W6BEG[10] ;
 wire \Tile_X9Y12_W6BEG[11] ;
 wire \Tile_X9Y12_W6BEG[1] ;
 wire \Tile_X9Y12_W6BEG[2] ;
 wire \Tile_X9Y12_W6BEG[3] ;
 wire \Tile_X9Y12_W6BEG[4] ;
 wire \Tile_X9Y12_W6BEG[5] ;
 wire \Tile_X9Y12_W6BEG[6] ;
 wire \Tile_X9Y12_W6BEG[7] ;
 wire \Tile_X9Y12_W6BEG[8] ;
 wire \Tile_X9Y12_W6BEG[9] ;
 wire \Tile_X9Y12_WW4BEG[0] ;
 wire \Tile_X9Y12_WW4BEG[10] ;
 wire \Tile_X9Y12_WW4BEG[11] ;
 wire \Tile_X9Y12_WW4BEG[12] ;
 wire \Tile_X9Y12_WW4BEG[13] ;
 wire \Tile_X9Y12_WW4BEG[14] ;
 wire \Tile_X9Y12_WW4BEG[15] ;
 wire \Tile_X9Y12_WW4BEG[1] ;
 wire \Tile_X9Y12_WW4BEG[2] ;
 wire \Tile_X9Y12_WW4BEG[3] ;
 wire \Tile_X9Y12_WW4BEG[4] ;
 wire \Tile_X9Y12_WW4BEG[5] ;
 wire \Tile_X9Y12_WW4BEG[6] ;
 wire \Tile_X9Y12_WW4BEG[7] ;
 wire \Tile_X9Y12_WW4BEG[8] ;
 wire \Tile_X9Y12_WW4BEG[9] ;
 wire Tile_X9Y13_Co;
 wire \Tile_X9Y13_E1BEG[0] ;
 wire \Tile_X9Y13_E1BEG[1] ;
 wire \Tile_X9Y13_E1BEG[2] ;
 wire \Tile_X9Y13_E1BEG[3] ;
 wire \Tile_X9Y13_E2BEG[0] ;
 wire \Tile_X9Y13_E2BEG[1] ;
 wire \Tile_X9Y13_E2BEG[2] ;
 wire \Tile_X9Y13_E2BEG[3] ;
 wire \Tile_X9Y13_E2BEG[4] ;
 wire \Tile_X9Y13_E2BEG[5] ;
 wire \Tile_X9Y13_E2BEG[6] ;
 wire \Tile_X9Y13_E2BEG[7] ;
 wire \Tile_X9Y13_E2BEGb[0] ;
 wire \Tile_X9Y13_E2BEGb[1] ;
 wire \Tile_X9Y13_E2BEGb[2] ;
 wire \Tile_X9Y13_E2BEGb[3] ;
 wire \Tile_X9Y13_E2BEGb[4] ;
 wire \Tile_X9Y13_E2BEGb[5] ;
 wire \Tile_X9Y13_E2BEGb[6] ;
 wire \Tile_X9Y13_E2BEGb[7] ;
 wire \Tile_X9Y13_E6BEG[0] ;
 wire \Tile_X9Y13_E6BEG[10] ;
 wire \Tile_X9Y13_E6BEG[11] ;
 wire \Tile_X9Y13_E6BEG[1] ;
 wire \Tile_X9Y13_E6BEG[2] ;
 wire \Tile_X9Y13_E6BEG[3] ;
 wire \Tile_X9Y13_E6BEG[4] ;
 wire \Tile_X9Y13_E6BEG[5] ;
 wire \Tile_X9Y13_E6BEG[6] ;
 wire \Tile_X9Y13_E6BEG[7] ;
 wire \Tile_X9Y13_E6BEG[8] ;
 wire \Tile_X9Y13_E6BEG[9] ;
 wire \Tile_X9Y13_EE4BEG[0] ;
 wire \Tile_X9Y13_EE4BEG[10] ;
 wire \Tile_X9Y13_EE4BEG[11] ;
 wire \Tile_X9Y13_EE4BEG[12] ;
 wire \Tile_X9Y13_EE4BEG[13] ;
 wire \Tile_X9Y13_EE4BEG[14] ;
 wire \Tile_X9Y13_EE4BEG[15] ;
 wire \Tile_X9Y13_EE4BEG[1] ;
 wire \Tile_X9Y13_EE4BEG[2] ;
 wire \Tile_X9Y13_EE4BEG[3] ;
 wire \Tile_X9Y13_EE4BEG[4] ;
 wire \Tile_X9Y13_EE4BEG[5] ;
 wire \Tile_X9Y13_EE4BEG[6] ;
 wire \Tile_X9Y13_EE4BEG[7] ;
 wire \Tile_X9Y13_EE4BEG[8] ;
 wire \Tile_X9Y13_EE4BEG[9] ;
 wire \Tile_X9Y13_FrameData_O[0] ;
 wire \Tile_X9Y13_FrameData_O[10] ;
 wire \Tile_X9Y13_FrameData_O[11] ;
 wire \Tile_X9Y13_FrameData_O[12] ;
 wire \Tile_X9Y13_FrameData_O[13] ;
 wire \Tile_X9Y13_FrameData_O[14] ;
 wire \Tile_X9Y13_FrameData_O[15] ;
 wire \Tile_X9Y13_FrameData_O[16] ;
 wire \Tile_X9Y13_FrameData_O[17] ;
 wire \Tile_X9Y13_FrameData_O[18] ;
 wire \Tile_X9Y13_FrameData_O[19] ;
 wire \Tile_X9Y13_FrameData_O[1] ;
 wire \Tile_X9Y13_FrameData_O[20] ;
 wire \Tile_X9Y13_FrameData_O[21] ;
 wire \Tile_X9Y13_FrameData_O[22] ;
 wire \Tile_X9Y13_FrameData_O[23] ;
 wire \Tile_X9Y13_FrameData_O[24] ;
 wire \Tile_X9Y13_FrameData_O[25] ;
 wire \Tile_X9Y13_FrameData_O[26] ;
 wire \Tile_X9Y13_FrameData_O[27] ;
 wire \Tile_X9Y13_FrameData_O[28] ;
 wire \Tile_X9Y13_FrameData_O[29] ;
 wire \Tile_X9Y13_FrameData_O[2] ;
 wire \Tile_X9Y13_FrameData_O[30] ;
 wire \Tile_X9Y13_FrameData_O[31] ;
 wire \Tile_X9Y13_FrameData_O[3] ;
 wire \Tile_X9Y13_FrameData_O[4] ;
 wire \Tile_X9Y13_FrameData_O[5] ;
 wire \Tile_X9Y13_FrameData_O[6] ;
 wire \Tile_X9Y13_FrameData_O[7] ;
 wire \Tile_X9Y13_FrameData_O[8] ;
 wire \Tile_X9Y13_FrameData_O[9] ;
 wire \Tile_X9Y13_FrameStrobe_O[0] ;
 wire \Tile_X9Y13_FrameStrobe_O[10] ;
 wire \Tile_X9Y13_FrameStrobe_O[11] ;
 wire \Tile_X9Y13_FrameStrobe_O[12] ;
 wire \Tile_X9Y13_FrameStrobe_O[13] ;
 wire \Tile_X9Y13_FrameStrobe_O[14] ;
 wire \Tile_X9Y13_FrameStrobe_O[15] ;
 wire \Tile_X9Y13_FrameStrobe_O[16] ;
 wire \Tile_X9Y13_FrameStrobe_O[17] ;
 wire \Tile_X9Y13_FrameStrobe_O[18] ;
 wire \Tile_X9Y13_FrameStrobe_O[19] ;
 wire \Tile_X9Y13_FrameStrobe_O[1] ;
 wire \Tile_X9Y13_FrameStrobe_O[2] ;
 wire \Tile_X9Y13_FrameStrobe_O[3] ;
 wire \Tile_X9Y13_FrameStrobe_O[4] ;
 wire \Tile_X9Y13_FrameStrobe_O[5] ;
 wire \Tile_X9Y13_FrameStrobe_O[6] ;
 wire \Tile_X9Y13_FrameStrobe_O[7] ;
 wire \Tile_X9Y13_FrameStrobe_O[8] ;
 wire \Tile_X9Y13_FrameStrobe_O[9] ;
 wire \Tile_X9Y13_N1BEG[0] ;
 wire \Tile_X9Y13_N1BEG[1] ;
 wire \Tile_X9Y13_N1BEG[2] ;
 wire \Tile_X9Y13_N1BEG[3] ;
 wire \Tile_X9Y13_N2BEG[0] ;
 wire \Tile_X9Y13_N2BEG[1] ;
 wire \Tile_X9Y13_N2BEG[2] ;
 wire \Tile_X9Y13_N2BEG[3] ;
 wire \Tile_X9Y13_N2BEG[4] ;
 wire \Tile_X9Y13_N2BEG[5] ;
 wire \Tile_X9Y13_N2BEG[6] ;
 wire \Tile_X9Y13_N2BEG[7] ;
 wire \Tile_X9Y13_N2BEGb[0] ;
 wire \Tile_X9Y13_N2BEGb[1] ;
 wire \Tile_X9Y13_N2BEGb[2] ;
 wire \Tile_X9Y13_N2BEGb[3] ;
 wire \Tile_X9Y13_N2BEGb[4] ;
 wire \Tile_X9Y13_N2BEGb[5] ;
 wire \Tile_X9Y13_N2BEGb[6] ;
 wire \Tile_X9Y13_N2BEGb[7] ;
 wire \Tile_X9Y13_N4BEG[0] ;
 wire \Tile_X9Y13_N4BEG[10] ;
 wire \Tile_X9Y13_N4BEG[11] ;
 wire \Tile_X9Y13_N4BEG[12] ;
 wire \Tile_X9Y13_N4BEG[13] ;
 wire \Tile_X9Y13_N4BEG[14] ;
 wire \Tile_X9Y13_N4BEG[15] ;
 wire \Tile_X9Y13_N4BEG[1] ;
 wire \Tile_X9Y13_N4BEG[2] ;
 wire \Tile_X9Y13_N4BEG[3] ;
 wire \Tile_X9Y13_N4BEG[4] ;
 wire \Tile_X9Y13_N4BEG[5] ;
 wire \Tile_X9Y13_N4BEG[6] ;
 wire \Tile_X9Y13_N4BEG[7] ;
 wire \Tile_X9Y13_N4BEG[8] ;
 wire \Tile_X9Y13_N4BEG[9] ;
 wire \Tile_X9Y13_NN4BEG[0] ;
 wire \Tile_X9Y13_NN4BEG[10] ;
 wire \Tile_X9Y13_NN4BEG[11] ;
 wire \Tile_X9Y13_NN4BEG[12] ;
 wire \Tile_X9Y13_NN4BEG[13] ;
 wire \Tile_X9Y13_NN4BEG[14] ;
 wire \Tile_X9Y13_NN4BEG[15] ;
 wire \Tile_X9Y13_NN4BEG[1] ;
 wire \Tile_X9Y13_NN4BEG[2] ;
 wire \Tile_X9Y13_NN4BEG[3] ;
 wire \Tile_X9Y13_NN4BEG[4] ;
 wire \Tile_X9Y13_NN4BEG[5] ;
 wire \Tile_X9Y13_NN4BEG[6] ;
 wire \Tile_X9Y13_NN4BEG[7] ;
 wire \Tile_X9Y13_NN4BEG[8] ;
 wire \Tile_X9Y13_NN4BEG[9] ;
 wire \Tile_X9Y13_S1BEG[0] ;
 wire \Tile_X9Y13_S1BEG[1] ;
 wire \Tile_X9Y13_S1BEG[2] ;
 wire \Tile_X9Y13_S1BEG[3] ;
 wire \Tile_X9Y13_S2BEG[0] ;
 wire \Tile_X9Y13_S2BEG[1] ;
 wire \Tile_X9Y13_S2BEG[2] ;
 wire \Tile_X9Y13_S2BEG[3] ;
 wire \Tile_X9Y13_S2BEG[4] ;
 wire \Tile_X9Y13_S2BEG[5] ;
 wire \Tile_X9Y13_S2BEG[6] ;
 wire \Tile_X9Y13_S2BEG[7] ;
 wire \Tile_X9Y13_S2BEGb[0] ;
 wire \Tile_X9Y13_S2BEGb[1] ;
 wire \Tile_X9Y13_S2BEGb[2] ;
 wire \Tile_X9Y13_S2BEGb[3] ;
 wire \Tile_X9Y13_S2BEGb[4] ;
 wire \Tile_X9Y13_S2BEGb[5] ;
 wire \Tile_X9Y13_S2BEGb[6] ;
 wire \Tile_X9Y13_S2BEGb[7] ;
 wire \Tile_X9Y13_S4BEG[0] ;
 wire \Tile_X9Y13_S4BEG[10] ;
 wire \Tile_X9Y13_S4BEG[11] ;
 wire \Tile_X9Y13_S4BEG[12] ;
 wire \Tile_X9Y13_S4BEG[13] ;
 wire \Tile_X9Y13_S4BEG[14] ;
 wire \Tile_X9Y13_S4BEG[15] ;
 wire \Tile_X9Y13_S4BEG[1] ;
 wire \Tile_X9Y13_S4BEG[2] ;
 wire \Tile_X9Y13_S4BEG[3] ;
 wire \Tile_X9Y13_S4BEG[4] ;
 wire \Tile_X9Y13_S4BEG[5] ;
 wire \Tile_X9Y13_S4BEG[6] ;
 wire \Tile_X9Y13_S4BEG[7] ;
 wire \Tile_X9Y13_S4BEG[8] ;
 wire \Tile_X9Y13_S4BEG[9] ;
 wire \Tile_X9Y13_SS4BEG[0] ;
 wire \Tile_X9Y13_SS4BEG[10] ;
 wire \Tile_X9Y13_SS4BEG[11] ;
 wire \Tile_X9Y13_SS4BEG[12] ;
 wire \Tile_X9Y13_SS4BEG[13] ;
 wire \Tile_X9Y13_SS4BEG[14] ;
 wire \Tile_X9Y13_SS4BEG[15] ;
 wire \Tile_X9Y13_SS4BEG[1] ;
 wire \Tile_X9Y13_SS4BEG[2] ;
 wire \Tile_X9Y13_SS4BEG[3] ;
 wire \Tile_X9Y13_SS4BEG[4] ;
 wire \Tile_X9Y13_SS4BEG[5] ;
 wire \Tile_X9Y13_SS4BEG[6] ;
 wire \Tile_X9Y13_SS4BEG[7] ;
 wire \Tile_X9Y13_SS4BEG[8] ;
 wire \Tile_X9Y13_SS4BEG[9] ;
 wire Tile_X9Y13_UserCLKo;
 wire \Tile_X9Y13_W1BEG[0] ;
 wire \Tile_X9Y13_W1BEG[1] ;
 wire \Tile_X9Y13_W1BEG[2] ;
 wire \Tile_X9Y13_W1BEG[3] ;
 wire \Tile_X9Y13_W2BEG[0] ;
 wire \Tile_X9Y13_W2BEG[1] ;
 wire \Tile_X9Y13_W2BEG[2] ;
 wire \Tile_X9Y13_W2BEG[3] ;
 wire \Tile_X9Y13_W2BEG[4] ;
 wire \Tile_X9Y13_W2BEG[5] ;
 wire \Tile_X9Y13_W2BEG[6] ;
 wire \Tile_X9Y13_W2BEG[7] ;
 wire \Tile_X9Y13_W2BEGb[0] ;
 wire \Tile_X9Y13_W2BEGb[1] ;
 wire \Tile_X9Y13_W2BEGb[2] ;
 wire \Tile_X9Y13_W2BEGb[3] ;
 wire \Tile_X9Y13_W2BEGb[4] ;
 wire \Tile_X9Y13_W2BEGb[5] ;
 wire \Tile_X9Y13_W2BEGb[6] ;
 wire \Tile_X9Y13_W2BEGb[7] ;
 wire \Tile_X9Y13_W6BEG[0] ;
 wire \Tile_X9Y13_W6BEG[10] ;
 wire \Tile_X9Y13_W6BEG[11] ;
 wire \Tile_X9Y13_W6BEG[1] ;
 wire \Tile_X9Y13_W6BEG[2] ;
 wire \Tile_X9Y13_W6BEG[3] ;
 wire \Tile_X9Y13_W6BEG[4] ;
 wire \Tile_X9Y13_W6BEG[5] ;
 wire \Tile_X9Y13_W6BEG[6] ;
 wire \Tile_X9Y13_W6BEG[7] ;
 wire \Tile_X9Y13_W6BEG[8] ;
 wire \Tile_X9Y13_W6BEG[9] ;
 wire \Tile_X9Y13_WW4BEG[0] ;
 wire \Tile_X9Y13_WW4BEG[10] ;
 wire \Tile_X9Y13_WW4BEG[11] ;
 wire \Tile_X9Y13_WW4BEG[12] ;
 wire \Tile_X9Y13_WW4BEG[13] ;
 wire \Tile_X9Y13_WW4BEG[14] ;
 wire \Tile_X9Y13_WW4BEG[15] ;
 wire \Tile_X9Y13_WW4BEG[1] ;
 wire \Tile_X9Y13_WW4BEG[2] ;
 wire \Tile_X9Y13_WW4BEG[3] ;
 wire \Tile_X9Y13_WW4BEG[4] ;
 wire \Tile_X9Y13_WW4BEG[5] ;
 wire \Tile_X9Y13_WW4BEG[6] ;
 wire \Tile_X9Y13_WW4BEG[7] ;
 wire \Tile_X9Y13_WW4BEG[8] ;
 wire \Tile_X9Y13_WW4BEG[9] ;
 wire Tile_X9Y14_Co;
 wire \Tile_X9Y14_E1BEG[0] ;
 wire \Tile_X9Y14_E1BEG[1] ;
 wire \Tile_X9Y14_E1BEG[2] ;
 wire \Tile_X9Y14_E1BEG[3] ;
 wire \Tile_X9Y14_E2BEG[0] ;
 wire \Tile_X9Y14_E2BEG[1] ;
 wire \Tile_X9Y14_E2BEG[2] ;
 wire \Tile_X9Y14_E2BEG[3] ;
 wire \Tile_X9Y14_E2BEG[4] ;
 wire \Tile_X9Y14_E2BEG[5] ;
 wire \Tile_X9Y14_E2BEG[6] ;
 wire \Tile_X9Y14_E2BEG[7] ;
 wire \Tile_X9Y14_E2BEGb[0] ;
 wire \Tile_X9Y14_E2BEGb[1] ;
 wire \Tile_X9Y14_E2BEGb[2] ;
 wire \Tile_X9Y14_E2BEGb[3] ;
 wire \Tile_X9Y14_E2BEGb[4] ;
 wire \Tile_X9Y14_E2BEGb[5] ;
 wire \Tile_X9Y14_E2BEGb[6] ;
 wire \Tile_X9Y14_E2BEGb[7] ;
 wire \Tile_X9Y14_E6BEG[0] ;
 wire \Tile_X9Y14_E6BEG[10] ;
 wire \Tile_X9Y14_E6BEG[11] ;
 wire \Tile_X9Y14_E6BEG[1] ;
 wire \Tile_X9Y14_E6BEG[2] ;
 wire \Tile_X9Y14_E6BEG[3] ;
 wire \Tile_X9Y14_E6BEG[4] ;
 wire \Tile_X9Y14_E6BEG[5] ;
 wire \Tile_X9Y14_E6BEG[6] ;
 wire \Tile_X9Y14_E6BEG[7] ;
 wire \Tile_X9Y14_E6BEG[8] ;
 wire \Tile_X9Y14_E6BEG[9] ;
 wire \Tile_X9Y14_EE4BEG[0] ;
 wire \Tile_X9Y14_EE4BEG[10] ;
 wire \Tile_X9Y14_EE4BEG[11] ;
 wire \Tile_X9Y14_EE4BEG[12] ;
 wire \Tile_X9Y14_EE4BEG[13] ;
 wire \Tile_X9Y14_EE4BEG[14] ;
 wire \Tile_X9Y14_EE4BEG[15] ;
 wire \Tile_X9Y14_EE4BEG[1] ;
 wire \Tile_X9Y14_EE4BEG[2] ;
 wire \Tile_X9Y14_EE4BEG[3] ;
 wire \Tile_X9Y14_EE4BEG[4] ;
 wire \Tile_X9Y14_EE4BEG[5] ;
 wire \Tile_X9Y14_EE4BEG[6] ;
 wire \Tile_X9Y14_EE4BEG[7] ;
 wire \Tile_X9Y14_EE4BEG[8] ;
 wire \Tile_X9Y14_EE4BEG[9] ;
 wire \Tile_X9Y14_FrameData_O[0] ;
 wire \Tile_X9Y14_FrameData_O[10] ;
 wire \Tile_X9Y14_FrameData_O[11] ;
 wire \Tile_X9Y14_FrameData_O[12] ;
 wire \Tile_X9Y14_FrameData_O[13] ;
 wire \Tile_X9Y14_FrameData_O[14] ;
 wire \Tile_X9Y14_FrameData_O[15] ;
 wire \Tile_X9Y14_FrameData_O[16] ;
 wire \Tile_X9Y14_FrameData_O[17] ;
 wire \Tile_X9Y14_FrameData_O[18] ;
 wire \Tile_X9Y14_FrameData_O[19] ;
 wire \Tile_X9Y14_FrameData_O[1] ;
 wire \Tile_X9Y14_FrameData_O[20] ;
 wire \Tile_X9Y14_FrameData_O[21] ;
 wire \Tile_X9Y14_FrameData_O[22] ;
 wire \Tile_X9Y14_FrameData_O[23] ;
 wire \Tile_X9Y14_FrameData_O[24] ;
 wire \Tile_X9Y14_FrameData_O[25] ;
 wire \Tile_X9Y14_FrameData_O[26] ;
 wire \Tile_X9Y14_FrameData_O[27] ;
 wire \Tile_X9Y14_FrameData_O[28] ;
 wire \Tile_X9Y14_FrameData_O[29] ;
 wire \Tile_X9Y14_FrameData_O[2] ;
 wire \Tile_X9Y14_FrameData_O[30] ;
 wire \Tile_X9Y14_FrameData_O[31] ;
 wire \Tile_X9Y14_FrameData_O[3] ;
 wire \Tile_X9Y14_FrameData_O[4] ;
 wire \Tile_X9Y14_FrameData_O[5] ;
 wire \Tile_X9Y14_FrameData_O[6] ;
 wire \Tile_X9Y14_FrameData_O[7] ;
 wire \Tile_X9Y14_FrameData_O[8] ;
 wire \Tile_X9Y14_FrameData_O[9] ;
 wire \Tile_X9Y14_FrameStrobe_O[0] ;
 wire \Tile_X9Y14_FrameStrobe_O[10] ;
 wire \Tile_X9Y14_FrameStrobe_O[11] ;
 wire \Tile_X9Y14_FrameStrobe_O[12] ;
 wire \Tile_X9Y14_FrameStrobe_O[13] ;
 wire \Tile_X9Y14_FrameStrobe_O[14] ;
 wire \Tile_X9Y14_FrameStrobe_O[15] ;
 wire \Tile_X9Y14_FrameStrobe_O[16] ;
 wire \Tile_X9Y14_FrameStrobe_O[17] ;
 wire \Tile_X9Y14_FrameStrobe_O[18] ;
 wire \Tile_X9Y14_FrameStrobe_O[19] ;
 wire \Tile_X9Y14_FrameStrobe_O[1] ;
 wire \Tile_X9Y14_FrameStrobe_O[2] ;
 wire \Tile_X9Y14_FrameStrobe_O[3] ;
 wire \Tile_X9Y14_FrameStrobe_O[4] ;
 wire \Tile_X9Y14_FrameStrobe_O[5] ;
 wire \Tile_X9Y14_FrameStrobe_O[6] ;
 wire \Tile_X9Y14_FrameStrobe_O[7] ;
 wire \Tile_X9Y14_FrameStrobe_O[8] ;
 wire \Tile_X9Y14_FrameStrobe_O[9] ;
 wire \Tile_X9Y14_N1BEG[0] ;
 wire \Tile_X9Y14_N1BEG[1] ;
 wire \Tile_X9Y14_N1BEG[2] ;
 wire \Tile_X9Y14_N1BEG[3] ;
 wire \Tile_X9Y14_N2BEG[0] ;
 wire \Tile_X9Y14_N2BEG[1] ;
 wire \Tile_X9Y14_N2BEG[2] ;
 wire \Tile_X9Y14_N2BEG[3] ;
 wire \Tile_X9Y14_N2BEG[4] ;
 wire \Tile_X9Y14_N2BEG[5] ;
 wire \Tile_X9Y14_N2BEG[6] ;
 wire \Tile_X9Y14_N2BEG[7] ;
 wire \Tile_X9Y14_N2BEGb[0] ;
 wire \Tile_X9Y14_N2BEGb[1] ;
 wire \Tile_X9Y14_N2BEGb[2] ;
 wire \Tile_X9Y14_N2BEGb[3] ;
 wire \Tile_X9Y14_N2BEGb[4] ;
 wire \Tile_X9Y14_N2BEGb[5] ;
 wire \Tile_X9Y14_N2BEGb[6] ;
 wire \Tile_X9Y14_N2BEGb[7] ;
 wire \Tile_X9Y14_N4BEG[0] ;
 wire \Tile_X9Y14_N4BEG[10] ;
 wire \Tile_X9Y14_N4BEG[11] ;
 wire \Tile_X9Y14_N4BEG[12] ;
 wire \Tile_X9Y14_N4BEG[13] ;
 wire \Tile_X9Y14_N4BEG[14] ;
 wire \Tile_X9Y14_N4BEG[15] ;
 wire \Tile_X9Y14_N4BEG[1] ;
 wire \Tile_X9Y14_N4BEG[2] ;
 wire \Tile_X9Y14_N4BEG[3] ;
 wire \Tile_X9Y14_N4BEG[4] ;
 wire \Tile_X9Y14_N4BEG[5] ;
 wire \Tile_X9Y14_N4BEG[6] ;
 wire \Tile_X9Y14_N4BEG[7] ;
 wire \Tile_X9Y14_N4BEG[8] ;
 wire \Tile_X9Y14_N4BEG[9] ;
 wire \Tile_X9Y14_NN4BEG[0] ;
 wire \Tile_X9Y14_NN4BEG[10] ;
 wire \Tile_X9Y14_NN4BEG[11] ;
 wire \Tile_X9Y14_NN4BEG[12] ;
 wire \Tile_X9Y14_NN4BEG[13] ;
 wire \Tile_X9Y14_NN4BEG[14] ;
 wire \Tile_X9Y14_NN4BEG[15] ;
 wire \Tile_X9Y14_NN4BEG[1] ;
 wire \Tile_X9Y14_NN4BEG[2] ;
 wire \Tile_X9Y14_NN4BEG[3] ;
 wire \Tile_X9Y14_NN4BEG[4] ;
 wire \Tile_X9Y14_NN4BEG[5] ;
 wire \Tile_X9Y14_NN4BEG[6] ;
 wire \Tile_X9Y14_NN4BEG[7] ;
 wire \Tile_X9Y14_NN4BEG[8] ;
 wire \Tile_X9Y14_NN4BEG[9] ;
 wire \Tile_X9Y14_S1BEG[0] ;
 wire \Tile_X9Y14_S1BEG[1] ;
 wire \Tile_X9Y14_S1BEG[2] ;
 wire \Tile_X9Y14_S1BEG[3] ;
 wire \Tile_X9Y14_S2BEG[0] ;
 wire \Tile_X9Y14_S2BEG[1] ;
 wire \Tile_X9Y14_S2BEG[2] ;
 wire \Tile_X9Y14_S2BEG[3] ;
 wire \Tile_X9Y14_S2BEG[4] ;
 wire \Tile_X9Y14_S2BEG[5] ;
 wire \Tile_X9Y14_S2BEG[6] ;
 wire \Tile_X9Y14_S2BEG[7] ;
 wire \Tile_X9Y14_S2BEGb[0] ;
 wire \Tile_X9Y14_S2BEGb[1] ;
 wire \Tile_X9Y14_S2BEGb[2] ;
 wire \Tile_X9Y14_S2BEGb[3] ;
 wire \Tile_X9Y14_S2BEGb[4] ;
 wire \Tile_X9Y14_S2BEGb[5] ;
 wire \Tile_X9Y14_S2BEGb[6] ;
 wire \Tile_X9Y14_S2BEGb[7] ;
 wire \Tile_X9Y14_S4BEG[0] ;
 wire \Tile_X9Y14_S4BEG[10] ;
 wire \Tile_X9Y14_S4BEG[11] ;
 wire \Tile_X9Y14_S4BEG[12] ;
 wire \Tile_X9Y14_S4BEG[13] ;
 wire \Tile_X9Y14_S4BEG[14] ;
 wire \Tile_X9Y14_S4BEG[15] ;
 wire \Tile_X9Y14_S4BEG[1] ;
 wire \Tile_X9Y14_S4BEG[2] ;
 wire \Tile_X9Y14_S4BEG[3] ;
 wire \Tile_X9Y14_S4BEG[4] ;
 wire \Tile_X9Y14_S4BEG[5] ;
 wire \Tile_X9Y14_S4BEG[6] ;
 wire \Tile_X9Y14_S4BEG[7] ;
 wire \Tile_X9Y14_S4BEG[8] ;
 wire \Tile_X9Y14_S4BEG[9] ;
 wire \Tile_X9Y14_SS4BEG[0] ;
 wire \Tile_X9Y14_SS4BEG[10] ;
 wire \Tile_X9Y14_SS4BEG[11] ;
 wire \Tile_X9Y14_SS4BEG[12] ;
 wire \Tile_X9Y14_SS4BEG[13] ;
 wire \Tile_X9Y14_SS4BEG[14] ;
 wire \Tile_X9Y14_SS4BEG[15] ;
 wire \Tile_X9Y14_SS4BEG[1] ;
 wire \Tile_X9Y14_SS4BEG[2] ;
 wire \Tile_X9Y14_SS4BEG[3] ;
 wire \Tile_X9Y14_SS4BEG[4] ;
 wire \Tile_X9Y14_SS4BEG[5] ;
 wire \Tile_X9Y14_SS4BEG[6] ;
 wire \Tile_X9Y14_SS4BEG[7] ;
 wire \Tile_X9Y14_SS4BEG[8] ;
 wire \Tile_X9Y14_SS4BEG[9] ;
 wire Tile_X9Y14_UserCLKo;
 wire \Tile_X9Y14_W1BEG[0] ;
 wire \Tile_X9Y14_W1BEG[1] ;
 wire \Tile_X9Y14_W1BEG[2] ;
 wire \Tile_X9Y14_W1BEG[3] ;
 wire \Tile_X9Y14_W2BEG[0] ;
 wire \Tile_X9Y14_W2BEG[1] ;
 wire \Tile_X9Y14_W2BEG[2] ;
 wire \Tile_X9Y14_W2BEG[3] ;
 wire \Tile_X9Y14_W2BEG[4] ;
 wire \Tile_X9Y14_W2BEG[5] ;
 wire \Tile_X9Y14_W2BEG[6] ;
 wire \Tile_X9Y14_W2BEG[7] ;
 wire \Tile_X9Y14_W2BEGb[0] ;
 wire \Tile_X9Y14_W2BEGb[1] ;
 wire \Tile_X9Y14_W2BEGb[2] ;
 wire \Tile_X9Y14_W2BEGb[3] ;
 wire \Tile_X9Y14_W2BEGb[4] ;
 wire \Tile_X9Y14_W2BEGb[5] ;
 wire \Tile_X9Y14_W2BEGb[6] ;
 wire \Tile_X9Y14_W2BEGb[7] ;
 wire \Tile_X9Y14_W6BEG[0] ;
 wire \Tile_X9Y14_W6BEG[10] ;
 wire \Tile_X9Y14_W6BEG[11] ;
 wire \Tile_X9Y14_W6BEG[1] ;
 wire \Tile_X9Y14_W6BEG[2] ;
 wire \Tile_X9Y14_W6BEG[3] ;
 wire \Tile_X9Y14_W6BEG[4] ;
 wire \Tile_X9Y14_W6BEG[5] ;
 wire \Tile_X9Y14_W6BEG[6] ;
 wire \Tile_X9Y14_W6BEG[7] ;
 wire \Tile_X9Y14_W6BEG[8] ;
 wire \Tile_X9Y14_W6BEG[9] ;
 wire \Tile_X9Y14_WW4BEG[0] ;
 wire \Tile_X9Y14_WW4BEG[10] ;
 wire \Tile_X9Y14_WW4BEG[11] ;
 wire \Tile_X9Y14_WW4BEG[12] ;
 wire \Tile_X9Y14_WW4BEG[13] ;
 wire \Tile_X9Y14_WW4BEG[14] ;
 wire \Tile_X9Y14_WW4BEG[15] ;
 wire \Tile_X9Y14_WW4BEG[1] ;
 wire \Tile_X9Y14_WW4BEG[2] ;
 wire \Tile_X9Y14_WW4BEG[3] ;
 wire \Tile_X9Y14_WW4BEG[4] ;
 wire \Tile_X9Y14_WW4BEG[5] ;
 wire \Tile_X9Y14_WW4BEG[6] ;
 wire \Tile_X9Y14_WW4BEG[7] ;
 wire \Tile_X9Y14_WW4BEG[8] ;
 wire \Tile_X9Y14_WW4BEG[9] ;
 wire Tile_X9Y15_Co;
 wire \Tile_X9Y15_FrameData_O[0] ;
 wire \Tile_X9Y15_FrameData_O[10] ;
 wire \Tile_X9Y15_FrameData_O[11] ;
 wire \Tile_X9Y15_FrameData_O[12] ;
 wire \Tile_X9Y15_FrameData_O[13] ;
 wire \Tile_X9Y15_FrameData_O[14] ;
 wire \Tile_X9Y15_FrameData_O[15] ;
 wire \Tile_X9Y15_FrameData_O[16] ;
 wire \Tile_X9Y15_FrameData_O[17] ;
 wire \Tile_X9Y15_FrameData_O[18] ;
 wire \Tile_X9Y15_FrameData_O[19] ;
 wire \Tile_X9Y15_FrameData_O[1] ;
 wire \Tile_X9Y15_FrameData_O[20] ;
 wire \Tile_X9Y15_FrameData_O[21] ;
 wire \Tile_X9Y15_FrameData_O[22] ;
 wire \Tile_X9Y15_FrameData_O[23] ;
 wire \Tile_X9Y15_FrameData_O[24] ;
 wire \Tile_X9Y15_FrameData_O[25] ;
 wire \Tile_X9Y15_FrameData_O[26] ;
 wire \Tile_X9Y15_FrameData_O[27] ;
 wire \Tile_X9Y15_FrameData_O[28] ;
 wire \Tile_X9Y15_FrameData_O[29] ;
 wire \Tile_X9Y15_FrameData_O[2] ;
 wire \Tile_X9Y15_FrameData_O[30] ;
 wire \Tile_X9Y15_FrameData_O[31] ;
 wire \Tile_X9Y15_FrameData_O[3] ;
 wire \Tile_X9Y15_FrameData_O[4] ;
 wire \Tile_X9Y15_FrameData_O[5] ;
 wire \Tile_X9Y15_FrameData_O[6] ;
 wire \Tile_X9Y15_FrameData_O[7] ;
 wire \Tile_X9Y15_FrameData_O[8] ;
 wire \Tile_X9Y15_FrameData_O[9] ;
 wire \Tile_X9Y15_FrameStrobe_O[0] ;
 wire \Tile_X9Y15_FrameStrobe_O[10] ;
 wire \Tile_X9Y15_FrameStrobe_O[11] ;
 wire \Tile_X9Y15_FrameStrobe_O[12] ;
 wire \Tile_X9Y15_FrameStrobe_O[13] ;
 wire \Tile_X9Y15_FrameStrobe_O[14] ;
 wire \Tile_X9Y15_FrameStrobe_O[15] ;
 wire \Tile_X9Y15_FrameStrobe_O[16] ;
 wire \Tile_X9Y15_FrameStrobe_O[17] ;
 wire \Tile_X9Y15_FrameStrobe_O[18] ;
 wire \Tile_X9Y15_FrameStrobe_O[19] ;
 wire \Tile_X9Y15_FrameStrobe_O[1] ;
 wire \Tile_X9Y15_FrameStrobe_O[2] ;
 wire \Tile_X9Y15_FrameStrobe_O[3] ;
 wire \Tile_X9Y15_FrameStrobe_O[4] ;
 wire \Tile_X9Y15_FrameStrobe_O[5] ;
 wire \Tile_X9Y15_FrameStrobe_O[6] ;
 wire \Tile_X9Y15_FrameStrobe_O[7] ;
 wire \Tile_X9Y15_FrameStrobe_O[8] ;
 wire \Tile_X9Y15_FrameStrobe_O[9] ;
 wire \Tile_X9Y15_N1BEG[0] ;
 wire \Tile_X9Y15_N1BEG[1] ;
 wire \Tile_X9Y15_N1BEG[2] ;
 wire \Tile_X9Y15_N1BEG[3] ;
 wire \Tile_X9Y15_N2BEG[0] ;
 wire \Tile_X9Y15_N2BEG[1] ;
 wire \Tile_X9Y15_N2BEG[2] ;
 wire \Tile_X9Y15_N2BEG[3] ;
 wire \Tile_X9Y15_N2BEG[4] ;
 wire \Tile_X9Y15_N2BEG[5] ;
 wire \Tile_X9Y15_N2BEG[6] ;
 wire \Tile_X9Y15_N2BEG[7] ;
 wire \Tile_X9Y15_N2BEGb[0] ;
 wire \Tile_X9Y15_N2BEGb[1] ;
 wire \Tile_X9Y15_N2BEGb[2] ;
 wire \Tile_X9Y15_N2BEGb[3] ;
 wire \Tile_X9Y15_N2BEGb[4] ;
 wire \Tile_X9Y15_N2BEGb[5] ;
 wire \Tile_X9Y15_N2BEGb[6] ;
 wire \Tile_X9Y15_N2BEGb[7] ;
 wire \Tile_X9Y15_N4BEG[0] ;
 wire \Tile_X9Y15_N4BEG[10] ;
 wire \Tile_X9Y15_N4BEG[11] ;
 wire \Tile_X9Y15_N4BEG[12] ;
 wire \Tile_X9Y15_N4BEG[13] ;
 wire \Tile_X9Y15_N4BEG[14] ;
 wire \Tile_X9Y15_N4BEG[15] ;
 wire \Tile_X9Y15_N4BEG[1] ;
 wire \Tile_X9Y15_N4BEG[2] ;
 wire \Tile_X9Y15_N4BEG[3] ;
 wire \Tile_X9Y15_N4BEG[4] ;
 wire \Tile_X9Y15_N4BEG[5] ;
 wire \Tile_X9Y15_N4BEG[6] ;
 wire \Tile_X9Y15_N4BEG[7] ;
 wire \Tile_X9Y15_N4BEG[8] ;
 wire \Tile_X9Y15_N4BEG[9] ;
 wire \Tile_X9Y15_NN4BEG[0] ;
 wire \Tile_X9Y15_NN4BEG[10] ;
 wire \Tile_X9Y15_NN4BEG[11] ;
 wire \Tile_X9Y15_NN4BEG[12] ;
 wire \Tile_X9Y15_NN4BEG[13] ;
 wire \Tile_X9Y15_NN4BEG[14] ;
 wire \Tile_X9Y15_NN4BEG[15] ;
 wire \Tile_X9Y15_NN4BEG[1] ;
 wire \Tile_X9Y15_NN4BEG[2] ;
 wire \Tile_X9Y15_NN4BEG[3] ;
 wire \Tile_X9Y15_NN4BEG[4] ;
 wire \Tile_X9Y15_NN4BEG[5] ;
 wire \Tile_X9Y15_NN4BEG[6] ;
 wire \Tile_X9Y15_NN4BEG[7] ;
 wire \Tile_X9Y15_NN4BEG[8] ;
 wire \Tile_X9Y15_NN4BEG[9] ;
 wire Tile_X9Y15_UserCLKo;
 wire Tile_X9Y1_Co;
 wire \Tile_X9Y1_E1BEG[0] ;
 wire \Tile_X9Y1_E1BEG[1] ;
 wire \Tile_X9Y1_E1BEG[2] ;
 wire \Tile_X9Y1_E1BEG[3] ;
 wire \Tile_X9Y1_E2BEG[0] ;
 wire \Tile_X9Y1_E2BEG[1] ;
 wire \Tile_X9Y1_E2BEG[2] ;
 wire \Tile_X9Y1_E2BEG[3] ;
 wire \Tile_X9Y1_E2BEG[4] ;
 wire \Tile_X9Y1_E2BEG[5] ;
 wire \Tile_X9Y1_E2BEG[6] ;
 wire \Tile_X9Y1_E2BEG[7] ;
 wire \Tile_X9Y1_E2BEGb[0] ;
 wire \Tile_X9Y1_E2BEGb[1] ;
 wire \Tile_X9Y1_E2BEGb[2] ;
 wire \Tile_X9Y1_E2BEGb[3] ;
 wire \Tile_X9Y1_E2BEGb[4] ;
 wire \Tile_X9Y1_E2BEGb[5] ;
 wire \Tile_X9Y1_E2BEGb[6] ;
 wire \Tile_X9Y1_E2BEGb[7] ;
 wire \Tile_X9Y1_E6BEG[0] ;
 wire \Tile_X9Y1_E6BEG[10] ;
 wire \Tile_X9Y1_E6BEG[11] ;
 wire \Tile_X9Y1_E6BEG[1] ;
 wire \Tile_X9Y1_E6BEG[2] ;
 wire \Tile_X9Y1_E6BEG[3] ;
 wire \Tile_X9Y1_E6BEG[4] ;
 wire \Tile_X9Y1_E6BEG[5] ;
 wire \Tile_X9Y1_E6BEG[6] ;
 wire \Tile_X9Y1_E6BEG[7] ;
 wire \Tile_X9Y1_E6BEG[8] ;
 wire \Tile_X9Y1_E6BEG[9] ;
 wire \Tile_X9Y1_EE4BEG[0] ;
 wire \Tile_X9Y1_EE4BEG[10] ;
 wire \Tile_X9Y1_EE4BEG[11] ;
 wire \Tile_X9Y1_EE4BEG[12] ;
 wire \Tile_X9Y1_EE4BEG[13] ;
 wire \Tile_X9Y1_EE4BEG[14] ;
 wire \Tile_X9Y1_EE4BEG[15] ;
 wire \Tile_X9Y1_EE4BEG[1] ;
 wire \Tile_X9Y1_EE4BEG[2] ;
 wire \Tile_X9Y1_EE4BEG[3] ;
 wire \Tile_X9Y1_EE4BEG[4] ;
 wire \Tile_X9Y1_EE4BEG[5] ;
 wire \Tile_X9Y1_EE4BEG[6] ;
 wire \Tile_X9Y1_EE4BEG[7] ;
 wire \Tile_X9Y1_EE4BEG[8] ;
 wire \Tile_X9Y1_EE4BEG[9] ;
 wire \Tile_X9Y1_FrameData_O[0] ;
 wire \Tile_X9Y1_FrameData_O[10] ;
 wire \Tile_X9Y1_FrameData_O[11] ;
 wire \Tile_X9Y1_FrameData_O[12] ;
 wire \Tile_X9Y1_FrameData_O[13] ;
 wire \Tile_X9Y1_FrameData_O[14] ;
 wire \Tile_X9Y1_FrameData_O[15] ;
 wire \Tile_X9Y1_FrameData_O[16] ;
 wire \Tile_X9Y1_FrameData_O[17] ;
 wire \Tile_X9Y1_FrameData_O[18] ;
 wire \Tile_X9Y1_FrameData_O[19] ;
 wire \Tile_X9Y1_FrameData_O[1] ;
 wire \Tile_X9Y1_FrameData_O[20] ;
 wire \Tile_X9Y1_FrameData_O[21] ;
 wire \Tile_X9Y1_FrameData_O[22] ;
 wire \Tile_X9Y1_FrameData_O[23] ;
 wire \Tile_X9Y1_FrameData_O[24] ;
 wire \Tile_X9Y1_FrameData_O[25] ;
 wire \Tile_X9Y1_FrameData_O[26] ;
 wire \Tile_X9Y1_FrameData_O[27] ;
 wire \Tile_X9Y1_FrameData_O[28] ;
 wire \Tile_X9Y1_FrameData_O[29] ;
 wire \Tile_X9Y1_FrameData_O[2] ;
 wire \Tile_X9Y1_FrameData_O[30] ;
 wire \Tile_X9Y1_FrameData_O[31] ;
 wire \Tile_X9Y1_FrameData_O[3] ;
 wire \Tile_X9Y1_FrameData_O[4] ;
 wire \Tile_X9Y1_FrameData_O[5] ;
 wire \Tile_X9Y1_FrameData_O[6] ;
 wire \Tile_X9Y1_FrameData_O[7] ;
 wire \Tile_X9Y1_FrameData_O[8] ;
 wire \Tile_X9Y1_FrameData_O[9] ;
 wire \Tile_X9Y1_FrameStrobe_O[0] ;
 wire \Tile_X9Y1_FrameStrobe_O[10] ;
 wire \Tile_X9Y1_FrameStrobe_O[11] ;
 wire \Tile_X9Y1_FrameStrobe_O[12] ;
 wire \Tile_X9Y1_FrameStrobe_O[13] ;
 wire \Tile_X9Y1_FrameStrobe_O[14] ;
 wire \Tile_X9Y1_FrameStrobe_O[15] ;
 wire \Tile_X9Y1_FrameStrobe_O[16] ;
 wire \Tile_X9Y1_FrameStrobe_O[17] ;
 wire \Tile_X9Y1_FrameStrobe_O[18] ;
 wire \Tile_X9Y1_FrameStrobe_O[19] ;
 wire \Tile_X9Y1_FrameStrobe_O[1] ;
 wire \Tile_X9Y1_FrameStrobe_O[2] ;
 wire \Tile_X9Y1_FrameStrobe_O[3] ;
 wire \Tile_X9Y1_FrameStrobe_O[4] ;
 wire \Tile_X9Y1_FrameStrobe_O[5] ;
 wire \Tile_X9Y1_FrameStrobe_O[6] ;
 wire \Tile_X9Y1_FrameStrobe_O[7] ;
 wire \Tile_X9Y1_FrameStrobe_O[8] ;
 wire \Tile_X9Y1_FrameStrobe_O[9] ;
 wire \Tile_X9Y1_N1BEG[0] ;
 wire \Tile_X9Y1_N1BEG[1] ;
 wire \Tile_X9Y1_N1BEG[2] ;
 wire \Tile_X9Y1_N1BEG[3] ;
 wire \Tile_X9Y1_N2BEG[0] ;
 wire \Tile_X9Y1_N2BEG[1] ;
 wire \Tile_X9Y1_N2BEG[2] ;
 wire \Tile_X9Y1_N2BEG[3] ;
 wire \Tile_X9Y1_N2BEG[4] ;
 wire \Tile_X9Y1_N2BEG[5] ;
 wire \Tile_X9Y1_N2BEG[6] ;
 wire \Tile_X9Y1_N2BEG[7] ;
 wire \Tile_X9Y1_N2BEGb[0] ;
 wire \Tile_X9Y1_N2BEGb[1] ;
 wire \Tile_X9Y1_N2BEGb[2] ;
 wire \Tile_X9Y1_N2BEGb[3] ;
 wire \Tile_X9Y1_N2BEGb[4] ;
 wire \Tile_X9Y1_N2BEGb[5] ;
 wire \Tile_X9Y1_N2BEGb[6] ;
 wire \Tile_X9Y1_N2BEGb[7] ;
 wire \Tile_X9Y1_N4BEG[0] ;
 wire \Tile_X9Y1_N4BEG[10] ;
 wire \Tile_X9Y1_N4BEG[11] ;
 wire \Tile_X9Y1_N4BEG[12] ;
 wire \Tile_X9Y1_N4BEG[13] ;
 wire \Tile_X9Y1_N4BEG[14] ;
 wire \Tile_X9Y1_N4BEG[15] ;
 wire \Tile_X9Y1_N4BEG[1] ;
 wire \Tile_X9Y1_N4BEG[2] ;
 wire \Tile_X9Y1_N4BEG[3] ;
 wire \Tile_X9Y1_N4BEG[4] ;
 wire \Tile_X9Y1_N4BEG[5] ;
 wire \Tile_X9Y1_N4BEG[6] ;
 wire \Tile_X9Y1_N4BEG[7] ;
 wire \Tile_X9Y1_N4BEG[8] ;
 wire \Tile_X9Y1_N4BEG[9] ;
 wire \Tile_X9Y1_NN4BEG[0] ;
 wire \Tile_X9Y1_NN4BEG[10] ;
 wire \Tile_X9Y1_NN4BEG[11] ;
 wire \Tile_X9Y1_NN4BEG[12] ;
 wire \Tile_X9Y1_NN4BEG[13] ;
 wire \Tile_X9Y1_NN4BEG[14] ;
 wire \Tile_X9Y1_NN4BEG[15] ;
 wire \Tile_X9Y1_NN4BEG[1] ;
 wire \Tile_X9Y1_NN4BEG[2] ;
 wire \Tile_X9Y1_NN4BEG[3] ;
 wire \Tile_X9Y1_NN4BEG[4] ;
 wire \Tile_X9Y1_NN4BEG[5] ;
 wire \Tile_X9Y1_NN4BEG[6] ;
 wire \Tile_X9Y1_NN4BEG[7] ;
 wire \Tile_X9Y1_NN4BEG[8] ;
 wire \Tile_X9Y1_NN4BEG[9] ;
 wire \Tile_X9Y1_S1BEG[0] ;
 wire \Tile_X9Y1_S1BEG[1] ;
 wire \Tile_X9Y1_S1BEG[2] ;
 wire \Tile_X9Y1_S1BEG[3] ;
 wire \Tile_X9Y1_S2BEG[0] ;
 wire \Tile_X9Y1_S2BEG[1] ;
 wire \Tile_X9Y1_S2BEG[2] ;
 wire \Tile_X9Y1_S2BEG[3] ;
 wire \Tile_X9Y1_S2BEG[4] ;
 wire \Tile_X9Y1_S2BEG[5] ;
 wire \Tile_X9Y1_S2BEG[6] ;
 wire \Tile_X9Y1_S2BEG[7] ;
 wire \Tile_X9Y1_S2BEGb[0] ;
 wire \Tile_X9Y1_S2BEGb[1] ;
 wire \Tile_X9Y1_S2BEGb[2] ;
 wire \Tile_X9Y1_S2BEGb[3] ;
 wire \Tile_X9Y1_S2BEGb[4] ;
 wire \Tile_X9Y1_S2BEGb[5] ;
 wire \Tile_X9Y1_S2BEGb[6] ;
 wire \Tile_X9Y1_S2BEGb[7] ;
 wire \Tile_X9Y1_S4BEG[0] ;
 wire \Tile_X9Y1_S4BEG[10] ;
 wire \Tile_X9Y1_S4BEG[11] ;
 wire \Tile_X9Y1_S4BEG[12] ;
 wire \Tile_X9Y1_S4BEG[13] ;
 wire \Tile_X9Y1_S4BEG[14] ;
 wire \Tile_X9Y1_S4BEG[15] ;
 wire \Tile_X9Y1_S4BEG[1] ;
 wire \Tile_X9Y1_S4BEG[2] ;
 wire \Tile_X9Y1_S4BEG[3] ;
 wire \Tile_X9Y1_S4BEG[4] ;
 wire \Tile_X9Y1_S4BEG[5] ;
 wire \Tile_X9Y1_S4BEG[6] ;
 wire \Tile_X9Y1_S4BEG[7] ;
 wire \Tile_X9Y1_S4BEG[8] ;
 wire \Tile_X9Y1_S4BEG[9] ;
 wire \Tile_X9Y1_SS4BEG[0] ;
 wire \Tile_X9Y1_SS4BEG[10] ;
 wire \Tile_X9Y1_SS4BEG[11] ;
 wire \Tile_X9Y1_SS4BEG[12] ;
 wire \Tile_X9Y1_SS4BEG[13] ;
 wire \Tile_X9Y1_SS4BEG[14] ;
 wire \Tile_X9Y1_SS4BEG[15] ;
 wire \Tile_X9Y1_SS4BEG[1] ;
 wire \Tile_X9Y1_SS4BEG[2] ;
 wire \Tile_X9Y1_SS4BEG[3] ;
 wire \Tile_X9Y1_SS4BEG[4] ;
 wire \Tile_X9Y1_SS4BEG[5] ;
 wire \Tile_X9Y1_SS4BEG[6] ;
 wire \Tile_X9Y1_SS4BEG[7] ;
 wire \Tile_X9Y1_SS4BEG[8] ;
 wire \Tile_X9Y1_SS4BEG[9] ;
 wire Tile_X9Y1_UserCLKo;
 wire \Tile_X9Y1_W1BEG[0] ;
 wire \Tile_X9Y1_W1BEG[1] ;
 wire \Tile_X9Y1_W1BEG[2] ;
 wire \Tile_X9Y1_W1BEG[3] ;
 wire \Tile_X9Y1_W2BEG[0] ;
 wire \Tile_X9Y1_W2BEG[1] ;
 wire \Tile_X9Y1_W2BEG[2] ;
 wire \Tile_X9Y1_W2BEG[3] ;
 wire \Tile_X9Y1_W2BEG[4] ;
 wire \Tile_X9Y1_W2BEG[5] ;
 wire \Tile_X9Y1_W2BEG[6] ;
 wire \Tile_X9Y1_W2BEG[7] ;
 wire \Tile_X9Y1_W2BEGb[0] ;
 wire \Tile_X9Y1_W2BEGb[1] ;
 wire \Tile_X9Y1_W2BEGb[2] ;
 wire \Tile_X9Y1_W2BEGb[3] ;
 wire \Tile_X9Y1_W2BEGb[4] ;
 wire \Tile_X9Y1_W2BEGb[5] ;
 wire \Tile_X9Y1_W2BEGb[6] ;
 wire \Tile_X9Y1_W2BEGb[7] ;
 wire \Tile_X9Y1_W6BEG[0] ;
 wire \Tile_X9Y1_W6BEG[10] ;
 wire \Tile_X9Y1_W6BEG[11] ;
 wire \Tile_X9Y1_W6BEG[1] ;
 wire \Tile_X9Y1_W6BEG[2] ;
 wire \Tile_X9Y1_W6BEG[3] ;
 wire \Tile_X9Y1_W6BEG[4] ;
 wire \Tile_X9Y1_W6BEG[5] ;
 wire \Tile_X9Y1_W6BEG[6] ;
 wire \Tile_X9Y1_W6BEG[7] ;
 wire \Tile_X9Y1_W6BEG[8] ;
 wire \Tile_X9Y1_W6BEG[9] ;
 wire \Tile_X9Y1_WW4BEG[0] ;
 wire \Tile_X9Y1_WW4BEG[10] ;
 wire \Tile_X9Y1_WW4BEG[11] ;
 wire \Tile_X9Y1_WW4BEG[12] ;
 wire \Tile_X9Y1_WW4BEG[13] ;
 wire \Tile_X9Y1_WW4BEG[14] ;
 wire \Tile_X9Y1_WW4BEG[15] ;
 wire \Tile_X9Y1_WW4BEG[1] ;
 wire \Tile_X9Y1_WW4BEG[2] ;
 wire \Tile_X9Y1_WW4BEG[3] ;
 wire \Tile_X9Y1_WW4BEG[4] ;
 wire \Tile_X9Y1_WW4BEG[5] ;
 wire \Tile_X9Y1_WW4BEG[6] ;
 wire \Tile_X9Y1_WW4BEG[7] ;
 wire \Tile_X9Y1_WW4BEG[8] ;
 wire \Tile_X9Y1_WW4BEG[9] ;
 wire Tile_X9Y2_Co;
 wire \Tile_X9Y2_E1BEG[0] ;
 wire \Tile_X9Y2_E1BEG[1] ;
 wire \Tile_X9Y2_E1BEG[2] ;
 wire \Tile_X9Y2_E1BEG[3] ;
 wire \Tile_X9Y2_E2BEG[0] ;
 wire \Tile_X9Y2_E2BEG[1] ;
 wire \Tile_X9Y2_E2BEG[2] ;
 wire \Tile_X9Y2_E2BEG[3] ;
 wire \Tile_X9Y2_E2BEG[4] ;
 wire \Tile_X9Y2_E2BEG[5] ;
 wire \Tile_X9Y2_E2BEG[6] ;
 wire \Tile_X9Y2_E2BEG[7] ;
 wire \Tile_X9Y2_E2BEGb[0] ;
 wire \Tile_X9Y2_E2BEGb[1] ;
 wire \Tile_X9Y2_E2BEGb[2] ;
 wire \Tile_X9Y2_E2BEGb[3] ;
 wire \Tile_X9Y2_E2BEGb[4] ;
 wire \Tile_X9Y2_E2BEGb[5] ;
 wire \Tile_X9Y2_E2BEGb[6] ;
 wire \Tile_X9Y2_E2BEGb[7] ;
 wire \Tile_X9Y2_E6BEG[0] ;
 wire \Tile_X9Y2_E6BEG[10] ;
 wire \Tile_X9Y2_E6BEG[11] ;
 wire \Tile_X9Y2_E6BEG[1] ;
 wire \Tile_X9Y2_E6BEG[2] ;
 wire \Tile_X9Y2_E6BEG[3] ;
 wire \Tile_X9Y2_E6BEG[4] ;
 wire \Tile_X9Y2_E6BEG[5] ;
 wire \Tile_X9Y2_E6BEG[6] ;
 wire \Tile_X9Y2_E6BEG[7] ;
 wire \Tile_X9Y2_E6BEG[8] ;
 wire \Tile_X9Y2_E6BEG[9] ;
 wire \Tile_X9Y2_EE4BEG[0] ;
 wire \Tile_X9Y2_EE4BEG[10] ;
 wire \Tile_X9Y2_EE4BEG[11] ;
 wire \Tile_X9Y2_EE4BEG[12] ;
 wire \Tile_X9Y2_EE4BEG[13] ;
 wire \Tile_X9Y2_EE4BEG[14] ;
 wire \Tile_X9Y2_EE4BEG[15] ;
 wire \Tile_X9Y2_EE4BEG[1] ;
 wire \Tile_X9Y2_EE4BEG[2] ;
 wire \Tile_X9Y2_EE4BEG[3] ;
 wire \Tile_X9Y2_EE4BEG[4] ;
 wire \Tile_X9Y2_EE4BEG[5] ;
 wire \Tile_X9Y2_EE4BEG[6] ;
 wire \Tile_X9Y2_EE4BEG[7] ;
 wire \Tile_X9Y2_EE4BEG[8] ;
 wire \Tile_X9Y2_EE4BEG[9] ;
 wire \Tile_X9Y2_FrameData_O[0] ;
 wire \Tile_X9Y2_FrameData_O[10] ;
 wire \Tile_X9Y2_FrameData_O[11] ;
 wire \Tile_X9Y2_FrameData_O[12] ;
 wire \Tile_X9Y2_FrameData_O[13] ;
 wire \Tile_X9Y2_FrameData_O[14] ;
 wire \Tile_X9Y2_FrameData_O[15] ;
 wire \Tile_X9Y2_FrameData_O[16] ;
 wire \Tile_X9Y2_FrameData_O[17] ;
 wire \Tile_X9Y2_FrameData_O[18] ;
 wire \Tile_X9Y2_FrameData_O[19] ;
 wire \Tile_X9Y2_FrameData_O[1] ;
 wire \Tile_X9Y2_FrameData_O[20] ;
 wire \Tile_X9Y2_FrameData_O[21] ;
 wire \Tile_X9Y2_FrameData_O[22] ;
 wire \Tile_X9Y2_FrameData_O[23] ;
 wire \Tile_X9Y2_FrameData_O[24] ;
 wire \Tile_X9Y2_FrameData_O[25] ;
 wire \Tile_X9Y2_FrameData_O[26] ;
 wire \Tile_X9Y2_FrameData_O[27] ;
 wire \Tile_X9Y2_FrameData_O[28] ;
 wire \Tile_X9Y2_FrameData_O[29] ;
 wire \Tile_X9Y2_FrameData_O[2] ;
 wire \Tile_X9Y2_FrameData_O[30] ;
 wire \Tile_X9Y2_FrameData_O[31] ;
 wire \Tile_X9Y2_FrameData_O[3] ;
 wire \Tile_X9Y2_FrameData_O[4] ;
 wire \Tile_X9Y2_FrameData_O[5] ;
 wire \Tile_X9Y2_FrameData_O[6] ;
 wire \Tile_X9Y2_FrameData_O[7] ;
 wire \Tile_X9Y2_FrameData_O[8] ;
 wire \Tile_X9Y2_FrameData_O[9] ;
 wire \Tile_X9Y2_FrameStrobe_O[0] ;
 wire \Tile_X9Y2_FrameStrobe_O[10] ;
 wire \Tile_X9Y2_FrameStrobe_O[11] ;
 wire \Tile_X9Y2_FrameStrobe_O[12] ;
 wire \Tile_X9Y2_FrameStrobe_O[13] ;
 wire \Tile_X9Y2_FrameStrobe_O[14] ;
 wire \Tile_X9Y2_FrameStrobe_O[15] ;
 wire \Tile_X9Y2_FrameStrobe_O[16] ;
 wire \Tile_X9Y2_FrameStrobe_O[17] ;
 wire \Tile_X9Y2_FrameStrobe_O[18] ;
 wire \Tile_X9Y2_FrameStrobe_O[19] ;
 wire \Tile_X9Y2_FrameStrobe_O[1] ;
 wire \Tile_X9Y2_FrameStrobe_O[2] ;
 wire \Tile_X9Y2_FrameStrobe_O[3] ;
 wire \Tile_X9Y2_FrameStrobe_O[4] ;
 wire \Tile_X9Y2_FrameStrobe_O[5] ;
 wire \Tile_X9Y2_FrameStrobe_O[6] ;
 wire \Tile_X9Y2_FrameStrobe_O[7] ;
 wire \Tile_X9Y2_FrameStrobe_O[8] ;
 wire \Tile_X9Y2_FrameStrobe_O[9] ;
 wire \Tile_X9Y2_N1BEG[0] ;
 wire \Tile_X9Y2_N1BEG[1] ;
 wire \Tile_X9Y2_N1BEG[2] ;
 wire \Tile_X9Y2_N1BEG[3] ;
 wire \Tile_X9Y2_N2BEG[0] ;
 wire \Tile_X9Y2_N2BEG[1] ;
 wire \Tile_X9Y2_N2BEG[2] ;
 wire \Tile_X9Y2_N2BEG[3] ;
 wire \Tile_X9Y2_N2BEG[4] ;
 wire \Tile_X9Y2_N2BEG[5] ;
 wire \Tile_X9Y2_N2BEG[6] ;
 wire \Tile_X9Y2_N2BEG[7] ;
 wire \Tile_X9Y2_N2BEGb[0] ;
 wire \Tile_X9Y2_N2BEGb[1] ;
 wire \Tile_X9Y2_N2BEGb[2] ;
 wire \Tile_X9Y2_N2BEGb[3] ;
 wire \Tile_X9Y2_N2BEGb[4] ;
 wire \Tile_X9Y2_N2BEGb[5] ;
 wire \Tile_X9Y2_N2BEGb[6] ;
 wire \Tile_X9Y2_N2BEGb[7] ;
 wire \Tile_X9Y2_N4BEG[0] ;
 wire \Tile_X9Y2_N4BEG[10] ;
 wire \Tile_X9Y2_N4BEG[11] ;
 wire \Tile_X9Y2_N4BEG[12] ;
 wire \Tile_X9Y2_N4BEG[13] ;
 wire \Tile_X9Y2_N4BEG[14] ;
 wire \Tile_X9Y2_N4BEG[15] ;
 wire \Tile_X9Y2_N4BEG[1] ;
 wire \Tile_X9Y2_N4BEG[2] ;
 wire \Tile_X9Y2_N4BEG[3] ;
 wire \Tile_X9Y2_N4BEG[4] ;
 wire \Tile_X9Y2_N4BEG[5] ;
 wire \Tile_X9Y2_N4BEG[6] ;
 wire \Tile_X9Y2_N4BEG[7] ;
 wire \Tile_X9Y2_N4BEG[8] ;
 wire \Tile_X9Y2_N4BEG[9] ;
 wire \Tile_X9Y2_NN4BEG[0] ;
 wire \Tile_X9Y2_NN4BEG[10] ;
 wire \Tile_X9Y2_NN4BEG[11] ;
 wire \Tile_X9Y2_NN4BEG[12] ;
 wire \Tile_X9Y2_NN4BEG[13] ;
 wire \Tile_X9Y2_NN4BEG[14] ;
 wire \Tile_X9Y2_NN4BEG[15] ;
 wire \Tile_X9Y2_NN4BEG[1] ;
 wire \Tile_X9Y2_NN4BEG[2] ;
 wire \Tile_X9Y2_NN4BEG[3] ;
 wire \Tile_X9Y2_NN4BEG[4] ;
 wire \Tile_X9Y2_NN4BEG[5] ;
 wire \Tile_X9Y2_NN4BEG[6] ;
 wire \Tile_X9Y2_NN4BEG[7] ;
 wire \Tile_X9Y2_NN4BEG[8] ;
 wire \Tile_X9Y2_NN4BEG[9] ;
 wire \Tile_X9Y2_S1BEG[0] ;
 wire \Tile_X9Y2_S1BEG[1] ;
 wire \Tile_X9Y2_S1BEG[2] ;
 wire \Tile_X9Y2_S1BEG[3] ;
 wire \Tile_X9Y2_S2BEG[0] ;
 wire \Tile_X9Y2_S2BEG[1] ;
 wire \Tile_X9Y2_S2BEG[2] ;
 wire \Tile_X9Y2_S2BEG[3] ;
 wire \Tile_X9Y2_S2BEG[4] ;
 wire \Tile_X9Y2_S2BEG[5] ;
 wire \Tile_X9Y2_S2BEG[6] ;
 wire \Tile_X9Y2_S2BEG[7] ;
 wire \Tile_X9Y2_S2BEGb[0] ;
 wire \Tile_X9Y2_S2BEGb[1] ;
 wire \Tile_X9Y2_S2BEGb[2] ;
 wire \Tile_X9Y2_S2BEGb[3] ;
 wire \Tile_X9Y2_S2BEGb[4] ;
 wire \Tile_X9Y2_S2BEGb[5] ;
 wire \Tile_X9Y2_S2BEGb[6] ;
 wire \Tile_X9Y2_S2BEGb[7] ;
 wire \Tile_X9Y2_S4BEG[0] ;
 wire \Tile_X9Y2_S4BEG[10] ;
 wire \Tile_X9Y2_S4BEG[11] ;
 wire \Tile_X9Y2_S4BEG[12] ;
 wire \Tile_X9Y2_S4BEG[13] ;
 wire \Tile_X9Y2_S4BEG[14] ;
 wire \Tile_X9Y2_S4BEG[15] ;
 wire \Tile_X9Y2_S4BEG[1] ;
 wire \Tile_X9Y2_S4BEG[2] ;
 wire \Tile_X9Y2_S4BEG[3] ;
 wire \Tile_X9Y2_S4BEG[4] ;
 wire \Tile_X9Y2_S4BEG[5] ;
 wire \Tile_X9Y2_S4BEG[6] ;
 wire \Tile_X9Y2_S4BEG[7] ;
 wire \Tile_X9Y2_S4BEG[8] ;
 wire \Tile_X9Y2_S4BEG[9] ;
 wire \Tile_X9Y2_SS4BEG[0] ;
 wire \Tile_X9Y2_SS4BEG[10] ;
 wire \Tile_X9Y2_SS4BEG[11] ;
 wire \Tile_X9Y2_SS4BEG[12] ;
 wire \Tile_X9Y2_SS4BEG[13] ;
 wire \Tile_X9Y2_SS4BEG[14] ;
 wire \Tile_X9Y2_SS4BEG[15] ;
 wire \Tile_X9Y2_SS4BEG[1] ;
 wire \Tile_X9Y2_SS4BEG[2] ;
 wire \Tile_X9Y2_SS4BEG[3] ;
 wire \Tile_X9Y2_SS4BEG[4] ;
 wire \Tile_X9Y2_SS4BEG[5] ;
 wire \Tile_X9Y2_SS4BEG[6] ;
 wire \Tile_X9Y2_SS4BEG[7] ;
 wire \Tile_X9Y2_SS4BEG[8] ;
 wire \Tile_X9Y2_SS4BEG[9] ;
 wire Tile_X9Y2_UserCLKo;
 wire \Tile_X9Y2_W1BEG[0] ;
 wire \Tile_X9Y2_W1BEG[1] ;
 wire \Tile_X9Y2_W1BEG[2] ;
 wire \Tile_X9Y2_W1BEG[3] ;
 wire \Tile_X9Y2_W2BEG[0] ;
 wire \Tile_X9Y2_W2BEG[1] ;
 wire \Tile_X9Y2_W2BEG[2] ;
 wire \Tile_X9Y2_W2BEG[3] ;
 wire \Tile_X9Y2_W2BEG[4] ;
 wire \Tile_X9Y2_W2BEG[5] ;
 wire \Tile_X9Y2_W2BEG[6] ;
 wire \Tile_X9Y2_W2BEG[7] ;
 wire \Tile_X9Y2_W2BEGb[0] ;
 wire \Tile_X9Y2_W2BEGb[1] ;
 wire \Tile_X9Y2_W2BEGb[2] ;
 wire \Tile_X9Y2_W2BEGb[3] ;
 wire \Tile_X9Y2_W2BEGb[4] ;
 wire \Tile_X9Y2_W2BEGb[5] ;
 wire \Tile_X9Y2_W2BEGb[6] ;
 wire \Tile_X9Y2_W2BEGb[7] ;
 wire \Tile_X9Y2_W6BEG[0] ;
 wire \Tile_X9Y2_W6BEG[10] ;
 wire \Tile_X9Y2_W6BEG[11] ;
 wire \Tile_X9Y2_W6BEG[1] ;
 wire \Tile_X9Y2_W6BEG[2] ;
 wire \Tile_X9Y2_W6BEG[3] ;
 wire \Tile_X9Y2_W6BEG[4] ;
 wire \Tile_X9Y2_W6BEG[5] ;
 wire \Tile_X9Y2_W6BEG[6] ;
 wire \Tile_X9Y2_W6BEG[7] ;
 wire \Tile_X9Y2_W6BEG[8] ;
 wire \Tile_X9Y2_W6BEG[9] ;
 wire \Tile_X9Y2_WW4BEG[0] ;
 wire \Tile_X9Y2_WW4BEG[10] ;
 wire \Tile_X9Y2_WW4BEG[11] ;
 wire \Tile_X9Y2_WW4BEG[12] ;
 wire \Tile_X9Y2_WW4BEG[13] ;
 wire \Tile_X9Y2_WW4BEG[14] ;
 wire \Tile_X9Y2_WW4BEG[15] ;
 wire \Tile_X9Y2_WW4BEG[1] ;
 wire \Tile_X9Y2_WW4BEG[2] ;
 wire \Tile_X9Y2_WW4BEG[3] ;
 wire \Tile_X9Y2_WW4BEG[4] ;
 wire \Tile_X9Y2_WW4BEG[5] ;
 wire \Tile_X9Y2_WW4BEG[6] ;
 wire \Tile_X9Y2_WW4BEG[7] ;
 wire \Tile_X9Y2_WW4BEG[8] ;
 wire \Tile_X9Y2_WW4BEG[9] ;
 wire Tile_X9Y3_Co;
 wire \Tile_X9Y3_E1BEG[0] ;
 wire \Tile_X9Y3_E1BEG[1] ;
 wire \Tile_X9Y3_E1BEG[2] ;
 wire \Tile_X9Y3_E1BEG[3] ;
 wire \Tile_X9Y3_E2BEG[0] ;
 wire \Tile_X9Y3_E2BEG[1] ;
 wire \Tile_X9Y3_E2BEG[2] ;
 wire \Tile_X9Y3_E2BEG[3] ;
 wire \Tile_X9Y3_E2BEG[4] ;
 wire \Tile_X9Y3_E2BEG[5] ;
 wire \Tile_X9Y3_E2BEG[6] ;
 wire \Tile_X9Y3_E2BEG[7] ;
 wire \Tile_X9Y3_E2BEGb[0] ;
 wire \Tile_X9Y3_E2BEGb[1] ;
 wire \Tile_X9Y3_E2BEGb[2] ;
 wire \Tile_X9Y3_E2BEGb[3] ;
 wire \Tile_X9Y3_E2BEGb[4] ;
 wire \Tile_X9Y3_E2BEGb[5] ;
 wire \Tile_X9Y3_E2BEGb[6] ;
 wire \Tile_X9Y3_E2BEGb[7] ;
 wire \Tile_X9Y3_E6BEG[0] ;
 wire \Tile_X9Y3_E6BEG[10] ;
 wire \Tile_X9Y3_E6BEG[11] ;
 wire \Tile_X9Y3_E6BEG[1] ;
 wire \Tile_X9Y3_E6BEG[2] ;
 wire \Tile_X9Y3_E6BEG[3] ;
 wire \Tile_X9Y3_E6BEG[4] ;
 wire \Tile_X9Y3_E6BEG[5] ;
 wire \Tile_X9Y3_E6BEG[6] ;
 wire \Tile_X9Y3_E6BEG[7] ;
 wire \Tile_X9Y3_E6BEG[8] ;
 wire \Tile_X9Y3_E6BEG[9] ;
 wire \Tile_X9Y3_EE4BEG[0] ;
 wire \Tile_X9Y3_EE4BEG[10] ;
 wire \Tile_X9Y3_EE4BEG[11] ;
 wire \Tile_X9Y3_EE4BEG[12] ;
 wire \Tile_X9Y3_EE4BEG[13] ;
 wire \Tile_X9Y3_EE4BEG[14] ;
 wire \Tile_X9Y3_EE4BEG[15] ;
 wire \Tile_X9Y3_EE4BEG[1] ;
 wire \Tile_X9Y3_EE4BEG[2] ;
 wire \Tile_X9Y3_EE4BEG[3] ;
 wire \Tile_X9Y3_EE4BEG[4] ;
 wire \Tile_X9Y3_EE4BEG[5] ;
 wire \Tile_X9Y3_EE4BEG[6] ;
 wire \Tile_X9Y3_EE4BEG[7] ;
 wire \Tile_X9Y3_EE4BEG[8] ;
 wire \Tile_X9Y3_EE4BEG[9] ;
 wire \Tile_X9Y3_FrameData_O[0] ;
 wire \Tile_X9Y3_FrameData_O[10] ;
 wire \Tile_X9Y3_FrameData_O[11] ;
 wire \Tile_X9Y3_FrameData_O[12] ;
 wire \Tile_X9Y3_FrameData_O[13] ;
 wire \Tile_X9Y3_FrameData_O[14] ;
 wire \Tile_X9Y3_FrameData_O[15] ;
 wire \Tile_X9Y3_FrameData_O[16] ;
 wire \Tile_X9Y3_FrameData_O[17] ;
 wire \Tile_X9Y3_FrameData_O[18] ;
 wire \Tile_X9Y3_FrameData_O[19] ;
 wire \Tile_X9Y3_FrameData_O[1] ;
 wire \Tile_X9Y3_FrameData_O[20] ;
 wire \Tile_X9Y3_FrameData_O[21] ;
 wire \Tile_X9Y3_FrameData_O[22] ;
 wire \Tile_X9Y3_FrameData_O[23] ;
 wire \Tile_X9Y3_FrameData_O[24] ;
 wire \Tile_X9Y3_FrameData_O[25] ;
 wire \Tile_X9Y3_FrameData_O[26] ;
 wire \Tile_X9Y3_FrameData_O[27] ;
 wire \Tile_X9Y3_FrameData_O[28] ;
 wire \Tile_X9Y3_FrameData_O[29] ;
 wire \Tile_X9Y3_FrameData_O[2] ;
 wire \Tile_X9Y3_FrameData_O[30] ;
 wire \Tile_X9Y3_FrameData_O[31] ;
 wire \Tile_X9Y3_FrameData_O[3] ;
 wire \Tile_X9Y3_FrameData_O[4] ;
 wire \Tile_X9Y3_FrameData_O[5] ;
 wire \Tile_X9Y3_FrameData_O[6] ;
 wire \Tile_X9Y3_FrameData_O[7] ;
 wire \Tile_X9Y3_FrameData_O[8] ;
 wire \Tile_X9Y3_FrameData_O[9] ;
 wire \Tile_X9Y3_FrameStrobe_O[0] ;
 wire \Tile_X9Y3_FrameStrobe_O[10] ;
 wire \Tile_X9Y3_FrameStrobe_O[11] ;
 wire \Tile_X9Y3_FrameStrobe_O[12] ;
 wire \Tile_X9Y3_FrameStrobe_O[13] ;
 wire \Tile_X9Y3_FrameStrobe_O[14] ;
 wire \Tile_X9Y3_FrameStrobe_O[15] ;
 wire \Tile_X9Y3_FrameStrobe_O[16] ;
 wire \Tile_X9Y3_FrameStrobe_O[17] ;
 wire \Tile_X9Y3_FrameStrobe_O[18] ;
 wire \Tile_X9Y3_FrameStrobe_O[19] ;
 wire \Tile_X9Y3_FrameStrobe_O[1] ;
 wire \Tile_X9Y3_FrameStrobe_O[2] ;
 wire \Tile_X9Y3_FrameStrobe_O[3] ;
 wire \Tile_X9Y3_FrameStrobe_O[4] ;
 wire \Tile_X9Y3_FrameStrobe_O[5] ;
 wire \Tile_X9Y3_FrameStrobe_O[6] ;
 wire \Tile_X9Y3_FrameStrobe_O[7] ;
 wire \Tile_X9Y3_FrameStrobe_O[8] ;
 wire \Tile_X9Y3_FrameStrobe_O[9] ;
 wire \Tile_X9Y3_N1BEG[0] ;
 wire \Tile_X9Y3_N1BEG[1] ;
 wire \Tile_X9Y3_N1BEG[2] ;
 wire \Tile_X9Y3_N1BEG[3] ;
 wire \Tile_X9Y3_N2BEG[0] ;
 wire \Tile_X9Y3_N2BEG[1] ;
 wire \Tile_X9Y3_N2BEG[2] ;
 wire \Tile_X9Y3_N2BEG[3] ;
 wire \Tile_X9Y3_N2BEG[4] ;
 wire \Tile_X9Y3_N2BEG[5] ;
 wire \Tile_X9Y3_N2BEG[6] ;
 wire \Tile_X9Y3_N2BEG[7] ;
 wire \Tile_X9Y3_N2BEGb[0] ;
 wire \Tile_X9Y3_N2BEGb[1] ;
 wire \Tile_X9Y3_N2BEGb[2] ;
 wire \Tile_X9Y3_N2BEGb[3] ;
 wire \Tile_X9Y3_N2BEGb[4] ;
 wire \Tile_X9Y3_N2BEGb[5] ;
 wire \Tile_X9Y3_N2BEGb[6] ;
 wire \Tile_X9Y3_N2BEGb[7] ;
 wire \Tile_X9Y3_N4BEG[0] ;
 wire \Tile_X9Y3_N4BEG[10] ;
 wire \Tile_X9Y3_N4BEG[11] ;
 wire \Tile_X9Y3_N4BEG[12] ;
 wire \Tile_X9Y3_N4BEG[13] ;
 wire \Tile_X9Y3_N4BEG[14] ;
 wire \Tile_X9Y3_N4BEG[15] ;
 wire \Tile_X9Y3_N4BEG[1] ;
 wire \Tile_X9Y3_N4BEG[2] ;
 wire \Tile_X9Y3_N4BEG[3] ;
 wire \Tile_X9Y3_N4BEG[4] ;
 wire \Tile_X9Y3_N4BEG[5] ;
 wire \Tile_X9Y3_N4BEG[6] ;
 wire \Tile_X9Y3_N4BEG[7] ;
 wire \Tile_X9Y3_N4BEG[8] ;
 wire \Tile_X9Y3_N4BEG[9] ;
 wire \Tile_X9Y3_NN4BEG[0] ;
 wire \Tile_X9Y3_NN4BEG[10] ;
 wire \Tile_X9Y3_NN4BEG[11] ;
 wire \Tile_X9Y3_NN4BEG[12] ;
 wire \Tile_X9Y3_NN4BEG[13] ;
 wire \Tile_X9Y3_NN4BEG[14] ;
 wire \Tile_X9Y3_NN4BEG[15] ;
 wire \Tile_X9Y3_NN4BEG[1] ;
 wire \Tile_X9Y3_NN4BEG[2] ;
 wire \Tile_X9Y3_NN4BEG[3] ;
 wire \Tile_X9Y3_NN4BEG[4] ;
 wire \Tile_X9Y3_NN4BEG[5] ;
 wire \Tile_X9Y3_NN4BEG[6] ;
 wire \Tile_X9Y3_NN4BEG[7] ;
 wire \Tile_X9Y3_NN4BEG[8] ;
 wire \Tile_X9Y3_NN4BEG[9] ;
 wire \Tile_X9Y3_S1BEG[0] ;
 wire \Tile_X9Y3_S1BEG[1] ;
 wire \Tile_X9Y3_S1BEG[2] ;
 wire \Tile_X9Y3_S1BEG[3] ;
 wire \Tile_X9Y3_S2BEG[0] ;
 wire \Tile_X9Y3_S2BEG[1] ;
 wire \Tile_X9Y3_S2BEG[2] ;
 wire \Tile_X9Y3_S2BEG[3] ;
 wire \Tile_X9Y3_S2BEG[4] ;
 wire \Tile_X9Y3_S2BEG[5] ;
 wire \Tile_X9Y3_S2BEG[6] ;
 wire \Tile_X9Y3_S2BEG[7] ;
 wire \Tile_X9Y3_S2BEGb[0] ;
 wire \Tile_X9Y3_S2BEGb[1] ;
 wire \Tile_X9Y3_S2BEGb[2] ;
 wire \Tile_X9Y3_S2BEGb[3] ;
 wire \Tile_X9Y3_S2BEGb[4] ;
 wire \Tile_X9Y3_S2BEGb[5] ;
 wire \Tile_X9Y3_S2BEGb[6] ;
 wire \Tile_X9Y3_S2BEGb[7] ;
 wire \Tile_X9Y3_S4BEG[0] ;
 wire \Tile_X9Y3_S4BEG[10] ;
 wire \Tile_X9Y3_S4BEG[11] ;
 wire \Tile_X9Y3_S4BEG[12] ;
 wire \Tile_X9Y3_S4BEG[13] ;
 wire \Tile_X9Y3_S4BEG[14] ;
 wire \Tile_X9Y3_S4BEG[15] ;
 wire \Tile_X9Y3_S4BEG[1] ;
 wire \Tile_X9Y3_S4BEG[2] ;
 wire \Tile_X9Y3_S4BEG[3] ;
 wire \Tile_X9Y3_S4BEG[4] ;
 wire \Tile_X9Y3_S4BEG[5] ;
 wire \Tile_X9Y3_S4BEG[6] ;
 wire \Tile_X9Y3_S4BEG[7] ;
 wire \Tile_X9Y3_S4BEG[8] ;
 wire \Tile_X9Y3_S4BEG[9] ;
 wire \Tile_X9Y3_SS4BEG[0] ;
 wire \Tile_X9Y3_SS4BEG[10] ;
 wire \Tile_X9Y3_SS4BEG[11] ;
 wire \Tile_X9Y3_SS4BEG[12] ;
 wire \Tile_X9Y3_SS4BEG[13] ;
 wire \Tile_X9Y3_SS4BEG[14] ;
 wire \Tile_X9Y3_SS4BEG[15] ;
 wire \Tile_X9Y3_SS4BEG[1] ;
 wire \Tile_X9Y3_SS4BEG[2] ;
 wire \Tile_X9Y3_SS4BEG[3] ;
 wire \Tile_X9Y3_SS4BEG[4] ;
 wire \Tile_X9Y3_SS4BEG[5] ;
 wire \Tile_X9Y3_SS4BEG[6] ;
 wire \Tile_X9Y3_SS4BEG[7] ;
 wire \Tile_X9Y3_SS4BEG[8] ;
 wire \Tile_X9Y3_SS4BEG[9] ;
 wire Tile_X9Y3_UserCLKo;
 wire \Tile_X9Y3_W1BEG[0] ;
 wire \Tile_X9Y3_W1BEG[1] ;
 wire \Tile_X9Y3_W1BEG[2] ;
 wire \Tile_X9Y3_W1BEG[3] ;
 wire \Tile_X9Y3_W2BEG[0] ;
 wire \Tile_X9Y3_W2BEG[1] ;
 wire \Tile_X9Y3_W2BEG[2] ;
 wire \Tile_X9Y3_W2BEG[3] ;
 wire \Tile_X9Y3_W2BEG[4] ;
 wire \Tile_X9Y3_W2BEG[5] ;
 wire \Tile_X9Y3_W2BEG[6] ;
 wire \Tile_X9Y3_W2BEG[7] ;
 wire \Tile_X9Y3_W2BEGb[0] ;
 wire \Tile_X9Y3_W2BEGb[1] ;
 wire \Tile_X9Y3_W2BEGb[2] ;
 wire \Tile_X9Y3_W2BEGb[3] ;
 wire \Tile_X9Y3_W2BEGb[4] ;
 wire \Tile_X9Y3_W2BEGb[5] ;
 wire \Tile_X9Y3_W2BEGb[6] ;
 wire \Tile_X9Y3_W2BEGb[7] ;
 wire \Tile_X9Y3_W6BEG[0] ;
 wire \Tile_X9Y3_W6BEG[10] ;
 wire \Tile_X9Y3_W6BEG[11] ;
 wire \Tile_X9Y3_W6BEG[1] ;
 wire \Tile_X9Y3_W6BEG[2] ;
 wire \Tile_X9Y3_W6BEG[3] ;
 wire \Tile_X9Y3_W6BEG[4] ;
 wire \Tile_X9Y3_W6BEG[5] ;
 wire \Tile_X9Y3_W6BEG[6] ;
 wire \Tile_X9Y3_W6BEG[7] ;
 wire \Tile_X9Y3_W6BEG[8] ;
 wire \Tile_X9Y3_W6BEG[9] ;
 wire \Tile_X9Y3_WW4BEG[0] ;
 wire \Tile_X9Y3_WW4BEG[10] ;
 wire \Tile_X9Y3_WW4BEG[11] ;
 wire \Tile_X9Y3_WW4BEG[12] ;
 wire \Tile_X9Y3_WW4BEG[13] ;
 wire \Tile_X9Y3_WW4BEG[14] ;
 wire \Tile_X9Y3_WW4BEG[15] ;
 wire \Tile_X9Y3_WW4BEG[1] ;
 wire \Tile_X9Y3_WW4BEG[2] ;
 wire \Tile_X9Y3_WW4BEG[3] ;
 wire \Tile_X9Y3_WW4BEG[4] ;
 wire \Tile_X9Y3_WW4BEG[5] ;
 wire \Tile_X9Y3_WW4BEG[6] ;
 wire \Tile_X9Y3_WW4BEG[7] ;
 wire \Tile_X9Y3_WW4BEG[8] ;
 wire \Tile_X9Y3_WW4BEG[9] ;
 wire Tile_X9Y4_Co;
 wire \Tile_X9Y4_E1BEG[0] ;
 wire \Tile_X9Y4_E1BEG[1] ;
 wire \Tile_X9Y4_E1BEG[2] ;
 wire \Tile_X9Y4_E1BEG[3] ;
 wire \Tile_X9Y4_E2BEG[0] ;
 wire \Tile_X9Y4_E2BEG[1] ;
 wire \Tile_X9Y4_E2BEG[2] ;
 wire \Tile_X9Y4_E2BEG[3] ;
 wire \Tile_X9Y4_E2BEG[4] ;
 wire \Tile_X9Y4_E2BEG[5] ;
 wire \Tile_X9Y4_E2BEG[6] ;
 wire \Tile_X9Y4_E2BEG[7] ;
 wire \Tile_X9Y4_E2BEGb[0] ;
 wire \Tile_X9Y4_E2BEGb[1] ;
 wire \Tile_X9Y4_E2BEGb[2] ;
 wire \Tile_X9Y4_E2BEGb[3] ;
 wire \Tile_X9Y4_E2BEGb[4] ;
 wire \Tile_X9Y4_E2BEGb[5] ;
 wire \Tile_X9Y4_E2BEGb[6] ;
 wire \Tile_X9Y4_E2BEGb[7] ;
 wire \Tile_X9Y4_E6BEG[0] ;
 wire \Tile_X9Y4_E6BEG[10] ;
 wire \Tile_X9Y4_E6BEG[11] ;
 wire \Tile_X9Y4_E6BEG[1] ;
 wire \Tile_X9Y4_E6BEG[2] ;
 wire \Tile_X9Y4_E6BEG[3] ;
 wire \Tile_X9Y4_E6BEG[4] ;
 wire \Tile_X9Y4_E6BEG[5] ;
 wire \Tile_X9Y4_E6BEG[6] ;
 wire \Tile_X9Y4_E6BEG[7] ;
 wire \Tile_X9Y4_E6BEG[8] ;
 wire \Tile_X9Y4_E6BEG[9] ;
 wire \Tile_X9Y4_EE4BEG[0] ;
 wire \Tile_X9Y4_EE4BEG[10] ;
 wire \Tile_X9Y4_EE4BEG[11] ;
 wire \Tile_X9Y4_EE4BEG[12] ;
 wire \Tile_X9Y4_EE4BEG[13] ;
 wire \Tile_X9Y4_EE4BEG[14] ;
 wire \Tile_X9Y4_EE4BEG[15] ;
 wire \Tile_X9Y4_EE4BEG[1] ;
 wire \Tile_X9Y4_EE4BEG[2] ;
 wire \Tile_X9Y4_EE4BEG[3] ;
 wire \Tile_X9Y4_EE4BEG[4] ;
 wire \Tile_X9Y4_EE4BEG[5] ;
 wire \Tile_X9Y4_EE4BEG[6] ;
 wire \Tile_X9Y4_EE4BEG[7] ;
 wire \Tile_X9Y4_EE4BEG[8] ;
 wire \Tile_X9Y4_EE4BEG[9] ;
 wire \Tile_X9Y4_FrameData_O[0] ;
 wire \Tile_X9Y4_FrameData_O[10] ;
 wire \Tile_X9Y4_FrameData_O[11] ;
 wire \Tile_X9Y4_FrameData_O[12] ;
 wire \Tile_X9Y4_FrameData_O[13] ;
 wire \Tile_X9Y4_FrameData_O[14] ;
 wire \Tile_X9Y4_FrameData_O[15] ;
 wire \Tile_X9Y4_FrameData_O[16] ;
 wire \Tile_X9Y4_FrameData_O[17] ;
 wire \Tile_X9Y4_FrameData_O[18] ;
 wire \Tile_X9Y4_FrameData_O[19] ;
 wire \Tile_X9Y4_FrameData_O[1] ;
 wire \Tile_X9Y4_FrameData_O[20] ;
 wire \Tile_X9Y4_FrameData_O[21] ;
 wire \Tile_X9Y4_FrameData_O[22] ;
 wire \Tile_X9Y4_FrameData_O[23] ;
 wire \Tile_X9Y4_FrameData_O[24] ;
 wire \Tile_X9Y4_FrameData_O[25] ;
 wire \Tile_X9Y4_FrameData_O[26] ;
 wire \Tile_X9Y4_FrameData_O[27] ;
 wire \Tile_X9Y4_FrameData_O[28] ;
 wire \Tile_X9Y4_FrameData_O[29] ;
 wire \Tile_X9Y4_FrameData_O[2] ;
 wire \Tile_X9Y4_FrameData_O[30] ;
 wire \Tile_X9Y4_FrameData_O[31] ;
 wire \Tile_X9Y4_FrameData_O[3] ;
 wire \Tile_X9Y4_FrameData_O[4] ;
 wire \Tile_X9Y4_FrameData_O[5] ;
 wire \Tile_X9Y4_FrameData_O[6] ;
 wire \Tile_X9Y4_FrameData_O[7] ;
 wire \Tile_X9Y4_FrameData_O[8] ;
 wire \Tile_X9Y4_FrameData_O[9] ;
 wire \Tile_X9Y4_FrameStrobe_O[0] ;
 wire \Tile_X9Y4_FrameStrobe_O[10] ;
 wire \Tile_X9Y4_FrameStrobe_O[11] ;
 wire \Tile_X9Y4_FrameStrobe_O[12] ;
 wire \Tile_X9Y4_FrameStrobe_O[13] ;
 wire \Tile_X9Y4_FrameStrobe_O[14] ;
 wire \Tile_X9Y4_FrameStrobe_O[15] ;
 wire \Tile_X9Y4_FrameStrobe_O[16] ;
 wire \Tile_X9Y4_FrameStrobe_O[17] ;
 wire \Tile_X9Y4_FrameStrobe_O[18] ;
 wire \Tile_X9Y4_FrameStrobe_O[19] ;
 wire \Tile_X9Y4_FrameStrobe_O[1] ;
 wire \Tile_X9Y4_FrameStrobe_O[2] ;
 wire \Tile_X9Y4_FrameStrobe_O[3] ;
 wire \Tile_X9Y4_FrameStrobe_O[4] ;
 wire \Tile_X9Y4_FrameStrobe_O[5] ;
 wire \Tile_X9Y4_FrameStrobe_O[6] ;
 wire \Tile_X9Y4_FrameStrobe_O[7] ;
 wire \Tile_X9Y4_FrameStrobe_O[8] ;
 wire \Tile_X9Y4_FrameStrobe_O[9] ;
 wire \Tile_X9Y4_N1BEG[0] ;
 wire \Tile_X9Y4_N1BEG[1] ;
 wire \Tile_X9Y4_N1BEG[2] ;
 wire \Tile_X9Y4_N1BEG[3] ;
 wire \Tile_X9Y4_N2BEG[0] ;
 wire \Tile_X9Y4_N2BEG[1] ;
 wire \Tile_X9Y4_N2BEG[2] ;
 wire \Tile_X9Y4_N2BEG[3] ;
 wire \Tile_X9Y4_N2BEG[4] ;
 wire \Tile_X9Y4_N2BEG[5] ;
 wire \Tile_X9Y4_N2BEG[6] ;
 wire \Tile_X9Y4_N2BEG[7] ;
 wire \Tile_X9Y4_N2BEGb[0] ;
 wire \Tile_X9Y4_N2BEGb[1] ;
 wire \Tile_X9Y4_N2BEGb[2] ;
 wire \Tile_X9Y4_N2BEGb[3] ;
 wire \Tile_X9Y4_N2BEGb[4] ;
 wire \Tile_X9Y4_N2BEGb[5] ;
 wire \Tile_X9Y4_N2BEGb[6] ;
 wire \Tile_X9Y4_N2BEGb[7] ;
 wire \Tile_X9Y4_N4BEG[0] ;
 wire \Tile_X9Y4_N4BEG[10] ;
 wire \Tile_X9Y4_N4BEG[11] ;
 wire \Tile_X9Y4_N4BEG[12] ;
 wire \Tile_X9Y4_N4BEG[13] ;
 wire \Tile_X9Y4_N4BEG[14] ;
 wire \Tile_X9Y4_N4BEG[15] ;
 wire \Tile_X9Y4_N4BEG[1] ;
 wire \Tile_X9Y4_N4BEG[2] ;
 wire \Tile_X9Y4_N4BEG[3] ;
 wire \Tile_X9Y4_N4BEG[4] ;
 wire \Tile_X9Y4_N4BEG[5] ;
 wire \Tile_X9Y4_N4BEG[6] ;
 wire \Tile_X9Y4_N4BEG[7] ;
 wire \Tile_X9Y4_N4BEG[8] ;
 wire \Tile_X9Y4_N4BEG[9] ;
 wire \Tile_X9Y4_NN4BEG[0] ;
 wire \Tile_X9Y4_NN4BEG[10] ;
 wire \Tile_X9Y4_NN4BEG[11] ;
 wire \Tile_X9Y4_NN4BEG[12] ;
 wire \Tile_X9Y4_NN4BEG[13] ;
 wire \Tile_X9Y4_NN4BEG[14] ;
 wire \Tile_X9Y4_NN4BEG[15] ;
 wire \Tile_X9Y4_NN4BEG[1] ;
 wire \Tile_X9Y4_NN4BEG[2] ;
 wire \Tile_X9Y4_NN4BEG[3] ;
 wire \Tile_X9Y4_NN4BEG[4] ;
 wire \Tile_X9Y4_NN4BEG[5] ;
 wire \Tile_X9Y4_NN4BEG[6] ;
 wire \Tile_X9Y4_NN4BEG[7] ;
 wire \Tile_X9Y4_NN4BEG[8] ;
 wire \Tile_X9Y4_NN4BEG[9] ;
 wire \Tile_X9Y4_S1BEG[0] ;
 wire \Tile_X9Y4_S1BEG[1] ;
 wire \Tile_X9Y4_S1BEG[2] ;
 wire \Tile_X9Y4_S1BEG[3] ;
 wire \Tile_X9Y4_S2BEG[0] ;
 wire \Tile_X9Y4_S2BEG[1] ;
 wire \Tile_X9Y4_S2BEG[2] ;
 wire \Tile_X9Y4_S2BEG[3] ;
 wire \Tile_X9Y4_S2BEG[4] ;
 wire \Tile_X9Y4_S2BEG[5] ;
 wire \Tile_X9Y4_S2BEG[6] ;
 wire \Tile_X9Y4_S2BEG[7] ;
 wire \Tile_X9Y4_S2BEGb[0] ;
 wire \Tile_X9Y4_S2BEGb[1] ;
 wire \Tile_X9Y4_S2BEGb[2] ;
 wire \Tile_X9Y4_S2BEGb[3] ;
 wire \Tile_X9Y4_S2BEGb[4] ;
 wire \Tile_X9Y4_S2BEGb[5] ;
 wire \Tile_X9Y4_S2BEGb[6] ;
 wire \Tile_X9Y4_S2BEGb[7] ;
 wire \Tile_X9Y4_S4BEG[0] ;
 wire \Tile_X9Y4_S4BEG[10] ;
 wire \Tile_X9Y4_S4BEG[11] ;
 wire \Tile_X9Y4_S4BEG[12] ;
 wire \Tile_X9Y4_S4BEG[13] ;
 wire \Tile_X9Y4_S4BEG[14] ;
 wire \Tile_X9Y4_S4BEG[15] ;
 wire \Tile_X9Y4_S4BEG[1] ;
 wire \Tile_X9Y4_S4BEG[2] ;
 wire \Tile_X9Y4_S4BEG[3] ;
 wire \Tile_X9Y4_S4BEG[4] ;
 wire \Tile_X9Y4_S4BEG[5] ;
 wire \Tile_X9Y4_S4BEG[6] ;
 wire \Tile_X9Y4_S4BEG[7] ;
 wire \Tile_X9Y4_S4BEG[8] ;
 wire \Tile_X9Y4_S4BEG[9] ;
 wire \Tile_X9Y4_SS4BEG[0] ;
 wire \Tile_X9Y4_SS4BEG[10] ;
 wire \Tile_X9Y4_SS4BEG[11] ;
 wire \Tile_X9Y4_SS4BEG[12] ;
 wire \Tile_X9Y4_SS4BEG[13] ;
 wire \Tile_X9Y4_SS4BEG[14] ;
 wire \Tile_X9Y4_SS4BEG[15] ;
 wire \Tile_X9Y4_SS4BEG[1] ;
 wire \Tile_X9Y4_SS4BEG[2] ;
 wire \Tile_X9Y4_SS4BEG[3] ;
 wire \Tile_X9Y4_SS4BEG[4] ;
 wire \Tile_X9Y4_SS4BEG[5] ;
 wire \Tile_X9Y4_SS4BEG[6] ;
 wire \Tile_X9Y4_SS4BEG[7] ;
 wire \Tile_X9Y4_SS4BEG[8] ;
 wire \Tile_X9Y4_SS4BEG[9] ;
 wire Tile_X9Y4_UserCLKo;
 wire \Tile_X9Y4_W1BEG[0] ;
 wire \Tile_X9Y4_W1BEG[1] ;
 wire \Tile_X9Y4_W1BEG[2] ;
 wire \Tile_X9Y4_W1BEG[3] ;
 wire \Tile_X9Y4_W2BEG[0] ;
 wire \Tile_X9Y4_W2BEG[1] ;
 wire \Tile_X9Y4_W2BEG[2] ;
 wire \Tile_X9Y4_W2BEG[3] ;
 wire \Tile_X9Y4_W2BEG[4] ;
 wire \Tile_X9Y4_W2BEG[5] ;
 wire \Tile_X9Y4_W2BEG[6] ;
 wire \Tile_X9Y4_W2BEG[7] ;
 wire \Tile_X9Y4_W2BEGb[0] ;
 wire \Tile_X9Y4_W2BEGb[1] ;
 wire \Tile_X9Y4_W2BEGb[2] ;
 wire \Tile_X9Y4_W2BEGb[3] ;
 wire \Tile_X9Y4_W2BEGb[4] ;
 wire \Tile_X9Y4_W2BEGb[5] ;
 wire \Tile_X9Y4_W2BEGb[6] ;
 wire \Tile_X9Y4_W2BEGb[7] ;
 wire \Tile_X9Y4_W6BEG[0] ;
 wire \Tile_X9Y4_W6BEG[10] ;
 wire \Tile_X9Y4_W6BEG[11] ;
 wire \Tile_X9Y4_W6BEG[1] ;
 wire \Tile_X9Y4_W6BEG[2] ;
 wire \Tile_X9Y4_W6BEG[3] ;
 wire \Tile_X9Y4_W6BEG[4] ;
 wire \Tile_X9Y4_W6BEG[5] ;
 wire \Tile_X9Y4_W6BEG[6] ;
 wire \Tile_X9Y4_W6BEG[7] ;
 wire \Tile_X9Y4_W6BEG[8] ;
 wire \Tile_X9Y4_W6BEG[9] ;
 wire \Tile_X9Y4_WW4BEG[0] ;
 wire \Tile_X9Y4_WW4BEG[10] ;
 wire \Tile_X9Y4_WW4BEG[11] ;
 wire \Tile_X9Y4_WW4BEG[12] ;
 wire \Tile_X9Y4_WW4BEG[13] ;
 wire \Tile_X9Y4_WW4BEG[14] ;
 wire \Tile_X9Y4_WW4BEG[15] ;
 wire \Tile_X9Y4_WW4BEG[1] ;
 wire \Tile_X9Y4_WW4BEG[2] ;
 wire \Tile_X9Y4_WW4BEG[3] ;
 wire \Tile_X9Y4_WW4BEG[4] ;
 wire \Tile_X9Y4_WW4BEG[5] ;
 wire \Tile_X9Y4_WW4BEG[6] ;
 wire \Tile_X9Y4_WW4BEG[7] ;
 wire \Tile_X9Y4_WW4BEG[8] ;
 wire \Tile_X9Y4_WW4BEG[9] ;
 wire Tile_X9Y5_Co;
 wire \Tile_X9Y5_E1BEG[0] ;
 wire \Tile_X9Y5_E1BEG[1] ;
 wire \Tile_X9Y5_E1BEG[2] ;
 wire \Tile_X9Y5_E1BEG[3] ;
 wire \Tile_X9Y5_E2BEG[0] ;
 wire \Tile_X9Y5_E2BEG[1] ;
 wire \Tile_X9Y5_E2BEG[2] ;
 wire \Tile_X9Y5_E2BEG[3] ;
 wire \Tile_X9Y5_E2BEG[4] ;
 wire \Tile_X9Y5_E2BEG[5] ;
 wire \Tile_X9Y5_E2BEG[6] ;
 wire \Tile_X9Y5_E2BEG[7] ;
 wire \Tile_X9Y5_E2BEGb[0] ;
 wire \Tile_X9Y5_E2BEGb[1] ;
 wire \Tile_X9Y5_E2BEGb[2] ;
 wire \Tile_X9Y5_E2BEGb[3] ;
 wire \Tile_X9Y5_E2BEGb[4] ;
 wire \Tile_X9Y5_E2BEGb[5] ;
 wire \Tile_X9Y5_E2BEGb[6] ;
 wire \Tile_X9Y5_E2BEGb[7] ;
 wire \Tile_X9Y5_E6BEG[0] ;
 wire \Tile_X9Y5_E6BEG[10] ;
 wire \Tile_X9Y5_E6BEG[11] ;
 wire \Tile_X9Y5_E6BEG[1] ;
 wire \Tile_X9Y5_E6BEG[2] ;
 wire \Tile_X9Y5_E6BEG[3] ;
 wire \Tile_X9Y5_E6BEG[4] ;
 wire \Tile_X9Y5_E6BEG[5] ;
 wire \Tile_X9Y5_E6BEG[6] ;
 wire \Tile_X9Y5_E6BEG[7] ;
 wire \Tile_X9Y5_E6BEG[8] ;
 wire \Tile_X9Y5_E6BEG[9] ;
 wire \Tile_X9Y5_EE4BEG[0] ;
 wire \Tile_X9Y5_EE4BEG[10] ;
 wire \Tile_X9Y5_EE4BEG[11] ;
 wire \Tile_X9Y5_EE4BEG[12] ;
 wire \Tile_X9Y5_EE4BEG[13] ;
 wire \Tile_X9Y5_EE4BEG[14] ;
 wire \Tile_X9Y5_EE4BEG[15] ;
 wire \Tile_X9Y5_EE4BEG[1] ;
 wire \Tile_X9Y5_EE4BEG[2] ;
 wire \Tile_X9Y5_EE4BEG[3] ;
 wire \Tile_X9Y5_EE4BEG[4] ;
 wire \Tile_X9Y5_EE4BEG[5] ;
 wire \Tile_X9Y5_EE4BEG[6] ;
 wire \Tile_X9Y5_EE4BEG[7] ;
 wire \Tile_X9Y5_EE4BEG[8] ;
 wire \Tile_X9Y5_EE4BEG[9] ;
 wire \Tile_X9Y5_FrameData_O[0] ;
 wire \Tile_X9Y5_FrameData_O[10] ;
 wire \Tile_X9Y5_FrameData_O[11] ;
 wire \Tile_X9Y5_FrameData_O[12] ;
 wire \Tile_X9Y5_FrameData_O[13] ;
 wire \Tile_X9Y5_FrameData_O[14] ;
 wire \Tile_X9Y5_FrameData_O[15] ;
 wire \Tile_X9Y5_FrameData_O[16] ;
 wire \Tile_X9Y5_FrameData_O[17] ;
 wire \Tile_X9Y5_FrameData_O[18] ;
 wire \Tile_X9Y5_FrameData_O[19] ;
 wire \Tile_X9Y5_FrameData_O[1] ;
 wire \Tile_X9Y5_FrameData_O[20] ;
 wire \Tile_X9Y5_FrameData_O[21] ;
 wire \Tile_X9Y5_FrameData_O[22] ;
 wire \Tile_X9Y5_FrameData_O[23] ;
 wire \Tile_X9Y5_FrameData_O[24] ;
 wire \Tile_X9Y5_FrameData_O[25] ;
 wire \Tile_X9Y5_FrameData_O[26] ;
 wire \Tile_X9Y5_FrameData_O[27] ;
 wire \Tile_X9Y5_FrameData_O[28] ;
 wire \Tile_X9Y5_FrameData_O[29] ;
 wire \Tile_X9Y5_FrameData_O[2] ;
 wire \Tile_X9Y5_FrameData_O[30] ;
 wire \Tile_X9Y5_FrameData_O[31] ;
 wire \Tile_X9Y5_FrameData_O[3] ;
 wire \Tile_X9Y5_FrameData_O[4] ;
 wire \Tile_X9Y5_FrameData_O[5] ;
 wire \Tile_X9Y5_FrameData_O[6] ;
 wire \Tile_X9Y5_FrameData_O[7] ;
 wire \Tile_X9Y5_FrameData_O[8] ;
 wire \Tile_X9Y5_FrameData_O[9] ;
 wire \Tile_X9Y5_FrameStrobe_O[0] ;
 wire \Tile_X9Y5_FrameStrobe_O[10] ;
 wire \Tile_X9Y5_FrameStrobe_O[11] ;
 wire \Tile_X9Y5_FrameStrobe_O[12] ;
 wire \Tile_X9Y5_FrameStrobe_O[13] ;
 wire \Tile_X9Y5_FrameStrobe_O[14] ;
 wire \Tile_X9Y5_FrameStrobe_O[15] ;
 wire \Tile_X9Y5_FrameStrobe_O[16] ;
 wire \Tile_X9Y5_FrameStrobe_O[17] ;
 wire \Tile_X9Y5_FrameStrobe_O[18] ;
 wire \Tile_X9Y5_FrameStrobe_O[19] ;
 wire \Tile_X9Y5_FrameStrobe_O[1] ;
 wire \Tile_X9Y5_FrameStrobe_O[2] ;
 wire \Tile_X9Y5_FrameStrobe_O[3] ;
 wire \Tile_X9Y5_FrameStrobe_O[4] ;
 wire \Tile_X9Y5_FrameStrobe_O[5] ;
 wire \Tile_X9Y5_FrameStrobe_O[6] ;
 wire \Tile_X9Y5_FrameStrobe_O[7] ;
 wire \Tile_X9Y5_FrameStrobe_O[8] ;
 wire \Tile_X9Y5_FrameStrobe_O[9] ;
 wire \Tile_X9Y5_N1BEG[0] ;
 wire \Tile_X9Y5_N1BEG[1] ;
 wire \Tile_X9Y5_N1BEG[2] ;
 wire \Tile_X9Y5_N1BEG[3] ;
 wire \Tile_X9Y5_N2BEG[0] ;
 wire \Tile_X9Y5_N2BEG[1] ;
 wire \Tile_X9Y5_N2BEG[2] ;
 wire \Tile_X9Y5_N2BEG[3] ;
 wire \Tile_X9Y5_N2BEG[4] ;
 wire \Tile_X9Y5_N2BEG[5] ;
 wire \Tile_X9Y5_N2BEG[6] ;
 wire \Tile_X9Y5_N2BEG[7] ;
 wire \Tile_X9Y5_N2BEGb[0] ;
 wire \Tile_X9Y5_N2BEGb[1] ;
 wire \Tile_X9Y5_N2BEGb[2] ;
 wire \Tile_X9Y5_N2BEGb[3] ;
 wire \Tile_X9Y5_N2BEGb[4] ;
 wire \Tile_X9Y5_N2BEGb[5] ;
 wire \Tile_X9Y5_N2BEGb[6] ;
 wire \Tile_X9Y5_N2BEGb[7] ;
 wire \Tile_X9Y5_N4BEG[0] ;
 wire \Tile_X9Y5_N4BEG[10] ;
 wire \Tile_X9Y5_N4BEG[11] ;
 wire \Tile_X9Y5_N4BEG[12] ;
 wire \Tile_X9Y5_N4BEG[13] ;
 wire \Tile_X9Y5_N4BEG[14] ;
 wire \Tile_X9Y5_N4BEG[15] ;
 wire \Tile_X9Y5_N4BEG[1] ;
 wire \Tile_X9Y5_N4BEG[2] ;
 wire \Tile_X9Y5_N4BEG[3] ;
 wire \Tile_X9Y5_N4BEG[4] ;
 wire \Tile_X9Y5_N4BEG[5] ;
 wire \Tile_X9Y5_N4BEG[6] ;
 wire \Tile_X9Y5_N4BEG[7] ;
 wire \Tile_X9Y5_N4BEG[8] ;
 wire \Tile_X9Y5_N4BEG[9] ;
 wire \Tile_X9Y5_NN4BEG[0] ;
 wire \Tile_X9Y5_NN4BEG[10] ;
 wire \Tile_X9Y5_NN4BEG[11] ;
 wire \Tile_X9Y5_NN4BEG[12] ;
 wire \Tile_X9Y5_NN4BEG[13] ;
 wire \Tile_X9Y5_NN4BEG[14] ;
 wire \Tile_X9Y5_NN4BEG[15] ;
 wire \Tile_X9Y5_NN4BEG[1] ;
 wire \Tile_X9Y5_NN4BEG[2] ;
 wire \Tile_X9Y5_NN4BEG[3] ;
 wire \Tile_X9Y5_NN4BEG[4] ;
 wire \Tile_X9Y5_NN4BEG[5] ;
 wire \Tile_X9Y5_NN4BEG[6] ;
 wire \Tile_X9Y5_NN4BEG[7] ;
 wire \Tile_X9Y5_NN4BEG[8] ;
 wire \Tile_X9Y5_NN4BEG[9] ;
 wire \Tile_X9Y5_S1BEG[0] ;
 wire \Tile_X9Y5_S1BEG[1] ;
 wire \Tile_X9Y5_S1BEG[2] ;
 wire \Tile_X9Y5_S1BEG[3] ;
 wire \Tile_X9Y5_S2BEG[0] ;
 wire \Tile_X9Y5_S2BEG[1] ;
 wire \Tile_X9Y5_S2BEG[2] ;
 wire \Tile_X9Y5_S2BEG[3] ;
 wire \Tile_X9Y5_S2BEG[4] ;
 wire \Tile_X9Y5_S2BEG[5] ;
 wire \Tile_X9Y5_S2BEG[6] ;
 wire \Tile_X9Y5_S2BEG[7] ;
 wire \Tile_X9Y5_S2BEGb[0] ;
 wire \Tile_X9Y5_S2BEGb[1] ;
 wire \Tile_X9Y5_S2BEGb[2] ;
 wire \Tile_X9Y5_S2BEGb[3] ;
 wire \Tile_X9Y5_S2BEGb[4] ;
 wire \Tile_X9Y5_S2BEGb[5] ;
 wire \Tile_X9Y5_S2BEGb[6] ;
 wire \Tile_X9Y5_S2BEGb[7] ;
 wire \Tile_X9Y5_S4BEG[0] ;
 wire \Tile_X9Y5_S4BEG[10] ;
 wire \Tile_X9Y5_S4BEG[11] ;
 wire \Tile_X9Y5_S4BEG[12] ;
 wire \Tile_X9Y5_S4BEG[13] ;
 wire \Tile_X9Y5_S4BEG[14] ;
 wire \Tile_X9Y5_S4BEG[15] ;
 wire \Tile_X9Y5_S4BEG[1] ;
 wire \Tile_X9Y5_S4BEG[2] ;
 wire \Tile_X9Y5_S4BEG[3] ;
 wire \Tile_X9Y5_S4BEG[4] ;
 wire \Tile_X9Y5_S4BEG[5] ;
 wire \Tile_X9Y5_S4BEG[6] ;
 wire \Tile_X9Y5_S4BEG[7] ;
 wire \Tile_X9Y5_S4BEG[8] ;
 wire \Tile_X9Y5_S4BEG[9] ;
 wire \Tile_X9Y5_SS4BEG[0] ;
 wire \Tile_X9Y5_SS4BEG[10] ;
 wire \Tile_X9Y5_SS4BEG[11] ;
 wire \Tile_X9Y5_SS4BEG[12] ;
 wire \Tile_X9Y5_SS4BEG[13] ;
 wire \Tile_X9Y5_SS4BEG[14] ;
 wire \Tile_X9Y5_SS4BEG[15] ;
 wire \Tile_X9Y5_SS4BEG[1] ;
 wire \Tile_X9Y5_SS4BEG[2] ;
 wire \Tile_X9Y5_SS4BEG[3] ;
 wire \Tile_X9Y5_SS4BEG[4] ;
 wire \Tile_X9Y5_SS4BEG[5] ;
 wire \Tile_X9Y5_SS4BEG[6] ;
 wire \Tile_X9Y5_SS4BEG[7] ;
 wire \Tile_X9Y5_SS4BEG[8] ;
 wire \Tile_X9Y5_SS4BEG[9] ;
 wire Tile_X9Y5_UserCLKo;
 wire \Tile_X9Y5_W1BEG[0] ;
 wire \Tile_X9Y5_W1BEG[1] ;
 wire \Tile_X9Y5_W1BEG[2] ;
 wire \Tile_X9Y5_W1BEG[3] ;
 wire \Tile_X9Y5_W2BEG[0] ;
 wire \Tile_X9Y5_W2BEG[1] ;
 wire \Tile_X9Y5_W2BEG[2] ;
 wire \Tile_X9Y5_W2BEG[3] ;
 wire \Tile_X9Y5_W2BEG[4] ;
 wire \Tile_X9Y5_W2BEG[5] ;
 wire \Tile_X9Y5_W2BEG[6] ;
 wire \Tile_X9Y5_W2BEG[7] ;
 wire \Tile_X9Y5_W2BEGb[0] ;
 wire \Tile_X9Y5_W2BEGb[1] ;
 wire \Tile_X9Y5_W2BEGb[2] ;
 wire \Tile_X9Y5_W2BEGb[3] ;
 wire \Tile_X9Y5_W2BEGb[4] ;
 wire \Tile_X9Y5_W2BEGb[5] ;
 wire \Tile_X9Y5_W2BEGb[6] ;
 wire \Tile_X9Y5_W2BEGb[7] ;
 wire \Tile_X9Y5_W6BEG[0] ;
 wire \Tile_X9Y5_W6BEG[10] ;
 wire \Tile_X9Y5_W6BEG[11] ;
 wire \Tile_X9Y5_W6BEG[1] ;
 wire \Tile_X9Y5_W6BEG[2] ;
 wire \Tile_X9Y5_W6BEG[3] ;
 wire \Tile_X9Y5_W6BEG[4] ;
 wire \Tile_X9Y5_W6BEG[5] ;
 wire \Tile_X9Y5_W6BEG[6] ;
 wire \Tile_X9Y5_W6BEG[7] ;
 wire \Tile_X9Y5_W6BEG[8] ;
 wire \Tile_X9Y5_W6BEG[9] ;
 wire \Tile_X9Y5_WW4BEG[0] ;
 wire \Tile_X9Y5_WW4BEG[10] ;
 wire \Tile_X9Y5_WW4BEG[11] ;
 wire \Tile_X9Y5_WW4BEG[12] ;
 wire \Tile_X9Y5_WW4BEG[13] ;
 wire \Tile_X9Y5_WW4BEG[14] ;
 wire \Tile_X9Y5_WW4BEG[15] ;
 wire \Tile_X9Y5_WW4BEG[1] ;
 wire \Tile_X9Y5_WW4BEG[2] ;
 wire \Tile_X9Y5_WW4BEG[3] ;
 wire \Tile_X9Y5_WW4BEG[4] ;
 wire \Tile_X9Y5_WW4BEG[5] ;
 wire \Tile_X9Y5_WW4BEG[6] ;
 wire \Tile_X9Y5_WW4BEG[7] ;
 wire \Tile_X9Y5_WW4BEG[8] ;
 wire \Tile_X9Y5_WW4BEG[9] ;
 wire Tile_X9Y6_Co;
 wire \Tile_X9Y6_E1BEG[0] ;
 wire \Tile_X9Y6_E1BEG[1] ;
 wire \Tile_X9Y6_E1BEG[2] ;
 wire \Tile_X9Y6_E1BEG[3] ;
 wire \Tile_X9Y6_E2BEG[0] ;
 wire \Tile_X9Y6_E2BEG[1] ;
 wire \Tile_X9Y6_E2BEG[2] ;
 wire \Tile_X9Y6_E2BEG[3] ;
 wire \Tile_X9Y6_E2BEG[4] ;
 wire \Tile_X9Y6_E2BEG[5] ;
 wire \Tile_X9Y6_E2BEG[6] ;
 wire \Tile_X9Y6_E2BEG[7] ;
 wire \Tile_X9Y6_E2BEGb[0] ;
 wire \Tile_X9Y6_E2BEGb[1] ;
 wire \Tile_X9Y6_E2BEGb[2] ;
 wire \Tile_X9Y6_E2BEGb[3] ;
 wire \Tile_X9Y6_E2BEGb[4] ;
 wire \Tile_X9Y6_E2BEGb[5] ;
 wire \Tile_X9Y6_E2BEGb[6] ;
 wire \Tile_X9Y6_E2BEGb[7] ;
 wire \Tile_X9Y6_E6BEG[0] ;
 wire \Tile_X9Y6_E6BEG[10] ;
 wire \Tile_X9Y6_E6BEG[11] ;
 wire \Tile_X9Y6_E6BEG[1] ;
 wire \Tile_X9Y6_E6BEG[2] ;
 wire \Tile_X9Y6_E6BEG[3] ;
 wire \Tile_X9Y6_E6BEG[4] ;
 wire \Tile_X9Y6_E6BEG[5] ;
 wire \Tile_X9Y6_E6BEG[6] ;
 wire \Tile_X9Y6_E6BEG[7] ;
 wire \Tile_X9Y6_E6BEG[8] ;
 wire \Tile_X9Y6_E6BEG[9] ;
 wire \Tile_X9Y6_EE4BEG[0] ;
 wire \Tile_X9Y6_EE4BEG[10] ;
 wire \Tile_X9Y6_EE4BEG[11] ;
 wire \Tile_X9Y6_EE4BEG[12] ;
 wire \Tile_X9Y6_EE4BEG[13] ;
 wire \Tile_X9Y6_EE4BEG[14] ;
 wire \Tile_X9Y6_EE4BEG[15] ;
 wire \Tile_X9Y6_EE4BEG[1] ;
 wire \Tile_X9Y6_EE4BEG[2] ;
 wire \Tile_X9Y6_EE4BEG[3] ;
 wire \Tile_X9Y6_EE4BEG[4] ;
 wire \Tile_X9Y6_EE4BEG[5] ;
 wire \Tile_X9Y6_EE4BEG[6] ;
 wire \Tile_X9Y6_EE4BEG[7] ;
 wire \Tile_X9Y6_EE4BEG[8] ;
 wire \Tile_X9Y6_EE4BEG[9] ;
 wire \Tile_X9Y6_FrameData_O[0] ;
 wire \Tile_X9Y6_FrameData_O[10] ;
 wire \Tile_X9Y6_FrameData_O[11] ;
 wire \Tile_X9Y6_FrameData_O[12] ;
 wire \Tile_X9Y6_FrameData_O[13] ;
 wire \Tile_X9Y6_FrameData_O[14] ;
 wire \Tile_X9Y6_FrameData_O[15] ;
 wire \Tile_X9Y6_FrameData_O[16] ;
 wire \Tile_X9Y6_FrameData_O[17] ;
 wire \Tile_X9Y6_FrameData_O[18] ;
 wire \Tile_X9Y6_FrameData_O[19] ;
 wire \Tile_X9Y6_FrameData_O[1] ;
 wire \Tile_X9Y6_FrameData_O[20] ;
 wire \Tile_X9Y6_FrameData_O[21] ;
 wire \Tile_X9Y6_FrameData_O[22] ;
 wire \Tile_X9Y6_FrameData_O[23] ;
 wire \Tile_X9Y6_FrameData_O[24] ;
 wire \Tile_X9Y6_FrameData_O[25] ;
 wire \Tile_X9Y6_FrameData_O[26] ;
 wire \Tile_X9Y6_FrameData_O[27] ;
 wire \Tile_X9Y6_FrameData_O[28] ;
 wire \Tile_X9Y6_FrameData_O[29] ;
 wire \Tile_X9Y6_FrameData_O[2] ;
 wire \Tile_X9Y6_FrameData_O[30] ;
 wire \Tile_X9Y6_FrameData_O[31] ;
 wire \Tile_X9Y6_FrameData_O[3] ;
 wire \Tile_X9Y6_FrameData_O[4] ;
 wire \Tile_X9Y6_FrameData_O[5] ;
 wire \Tile_X9Y6_FrameData_O[6] ;
 wire \Tile_X9Y6_FrameData_O[7] ;
 wire \Tile_X9Y6_FrameData_O[8] ;
 wire \Tile_X9Y6_FrameData_O[9] ;
 wire \Tile_X9Y6_FrameStrobe_O[0] ;
 wire \Tile_X9Y6_FrameStrobe_O[10] ;
 wire \Tile_X9Y6_FrameStrobe_O[11] ;
 wire \Tile_X9Y6_FrameStrobe_O[12] ;
 wire \Tile_X9Y6_FrameStrobe_O[13] ;
 wire \Tile_X9Y6_FrameStrobe_O[14] ;
 wire \Tile_X9Y6_FrameStrobe_O[15] ;
 wire \Tile_X9Y6_FrameStrobe_O[16] ;
 wire \Tile_X9Y6_FrameStrobe_O[17] ;
 wire \Tile_X9Y6_FrameStrobe_O[18] ;
 wire \Tile_X9Y6_FrameStrobe_O[19] ;
 wire \Tile_X9Y6_FrameStrobe_O[1] ;
 wire \Tile_X9Y6_FrameStrobe_O[2] ;
 wire \Tile_X9Y6_FrameStrobe_O[3] ;
 wire \Tile_X9Y6_FrameStrobe_O[4] ;
 wire \Tile_X9Y6_FrameStrobe_O[5] ;
 wire \Tile_X9Y6_FrameStrobe_O[6] ;
 wire \Tile_X9Y6_FrameStrobe_O[7] ;
 wire \Tile_X9Y6_FrameStrobe_O[8] ;
 wire \Tile_X9Y6_FrameStrobe_O[9] ;
 wire \Tile_X9Y6_N1BEG[0] ;
 wire \Tile_X9Y6_N1BEG[1] ;
 wire \Tile_X9Y6_N1BEG[2] ;
 wire \Tile_X9Y6_N1BEG[3] ;
 wire \Tile_X9Y6_N2BEG[0] ;
 wire \Tile_X9Y6_N2BEG[1] ;
 wire \Tile_X9Y6_N2BEG[2] ;
 wire \Tile_X9Y6_N2BEG[3] ;
 wire \Tile_X9Y6_N2BEG[4] ;
 wire \Tile_X9Y6_N2BEG[5] ;
 wire \Tile_X9Y6_N2BEG[6] ;
 wire \Tile_X9Y6_N2BEG[7] ;
 wire \Tile_X9Y6_N2BEGb[0] ;
 wire \Tile_X9Y6_N2BEGb[1] ;
 wire \Tile_X9Y6_N2BEGb[2] ;
 wire \Tile_X9Y6_N2BEGb[3] ;
 wire \Tile_X9Y6_N2BEGb[4] ;
 wire \Tile_X9Y6_N2BEGb[5] ;
 wire \Tile_X9Y6_N2BEGb[6] ;
 wire \Tile_X9Y6_N2BEGb[7] ;
 wire \Tile_X9Y6_N4BEG[0] ;
 wire \Tile_X9Y6_N4BEG[10] ;
 wire \Tile_X9Y6_N4BEG[11] ;
 wire \Tile_X9Y6_N4BEG[12] ;
 wire \Tile_X9Y6_N4BEG[13] ;
 wire \Tile_X9Y6_N4BEG[14] ;
 wire \Tile_X9Y6_N4BEG[15] ;
 wire \Tile_X9Y6_N4BEG[1] ;
 wire \Tile_X9Y6_N4BEG[2] ;
 wire \Tile_X9Y6_N4BEG[3] ;
 wire \Tile_X9Y6_N4BEG[4] ;
 wire \Tile_X9Y6_N4BEG[5] ;
 wire \Tile_X9Y6_N4BEG[6] ;
 wire \Tile_X9Y6_N4BEG[7] ;
 wire \Tile_X9Y6_N4BEG[8] ;
 wire \Tile_X9Y6_N4BEG[9] ;
 wire \Tile_X9Y6_NN4BEG[0] ;
 wire \Tile_X9Y6_NN4BEG[10] ;
 wire \Tile_X9Y6_NN4BEG[11] ;
 wire \Tile_X9Y6_NN4BEG[12] ;
 wire \Tile_X9Y6_NN4BEG[13] ;
 wire \Tile_X9Y6_NN4BEG[14] ;
 wire \Tile_X9Y6_NN4BEG[15] ;
 wire \Tile_X9Y6_NN4BEG[1] ;
 wire \Tile_X9Y6_NN4BEG[2] ;
 wire \Tile_X9Y6_NN4BEG[3] ;
 wire \Tile_X9Y6_NN4BEG[4] ;
 wire \Tile_X9Y6_NN4BEG[5] ;
 wire \Tile_X9Y6_NN4BEG[6] ;
 wire \Tile_X9Y6_NN4BEG[7] ;
 wire \Tile_X9Y6_NN4BEG[8] ;
 wire \Tile_X9Y6_NN4BEG[9] ;
 wire \Tile_X9Y6_S1BEG[0] ;
 wire \Tile_X9Y6_S1BEG[1] ;
 wire \Tile_X9Y6_S1BEG[2] ;
 wire \Tile_X9Y6_S1BEG[3] ;
 wire \Tile_X9Y6_S2BEG[0] ;
 wire \Tile_X9Y6_S2BEG[1] ;
 wire \Tile_X9Y6_S2BEG[2] ;
 wire \Tile_X9Y6_S2BEG[3] ;
 wire \Tile_X9Y6_S2BEG[4] ;
 wire \Tile_X9Y6_S2BEG[5] ;
 wire \Tile_X9Y6_S2BEG[6] ;
 wire \Tile_X9Y6_S2BEG[7] ;
 wire \Tile_X9Y6_S2BEGb[0] ;
 wire \Tile_X9Y6_S2BEGb[1] ;
 wire \Tile_X9Y6_S2BEGb[2] ;
 wire \Tile_X9Y6_S2BEGb[3] ;
 wire \Tile_X9Y6_S2BEGb[4] ;
 wire \Tile_X9Y6_S2BEGb[5] ;
 wire \Tile_X9Y6_S2BEGb[6] ;
 wire \Tile_X9Y6_S2BEGb[7] ;
 wire \Tile_X9Y6_S4BEG[0] ;
 wire \Tile_X9Y6_S4BEG[10] ;
 wire \Tile_X9Y6_S4BEG[11] ;
 wire \Tile_X9Y6_S4BEG[12] ;
 wire \Tile_X9Y6_S4BEG[13] ;
 wire \Tile_X9Y6_S4BEG[14] ;
 wire \Tile_X9Y6_S4BEG[15] ;
 wire \Tile_X9Y6_S4BEG[1] ;
 wire \Tile_X9Y6_S4BEG[2] ;
 wire \Tile_X9Y6_S4BEG[3] ;
 wire \Tile_X9Y6_S4BEG[4] ;
 wire \Tile_X9Y6_S4BEG[5] ;
 wire \Tile_X9Y6_S4BEG[6] ;
 wire \Tile_X9Y6_S4BEG[7] ;
 wire \Tile_X9Y6_S4BEG[8] ;
 wire \Tile_X9Y6_S4BEG[9] ;
 wire \Tile_X9Y6_SS4BEG[0] ;
 wire \Tile_X9Y6_SS4BEG[10] ;
 wire \Tile_X9Y6_SS4BEG[11] ;
 wire \Tile_X9Y6_SS4BEG[12] ;
 wire \Tile_X9Y6_SS4BEG[13] ;
 wire \Tile_X9Y6_SS4BEG[14] ;
 wire \Tile_X9Y6_SS4BEG[15] ;
 wire \Tile_X9Y6_SS4BEG[1] ;
 wire \Tile_X9Y6_SS4BEG[2] ;
 wire \Tile_X9Y6_SS4BEG[3] ;
 wire \Tile_X9Y6_SS4BEG[4] ;
 wire \Tile_X9Y6_SS4BEG[5] ;
 wire \Tile_X9Y6_SS4BEG[6] ;
 wire \Tile_X9Y6_SS4BEG[7] ;
 wire \Tile_X9Y6_SS4BEG[8] ;
 wire \Tile_X9Y6_SS4BEG[9] ;
 wire Tile_X9Y6_UserCLKo;
 wire \Tile_X9Y6_W1BEG[0] ;
 wire \Tile_X9Y6_W1BEG[1] ;
 wire \Tile_X9Y6_W1BEG[2] ;
 wire \Tile_X9Y6_W1BEG[3] ;
 wire \Tile_X9Y6_W2BEG[0] ;
 wire \Tile_X9Y6_W2BEG[1] ;
 wire \Tile_X9Y6_W2BEG[2] ;
 wire \Tile_X9Y6_W2BEG[3] ;
 wire \Tile_X9Y6_W2BEG[4] ;
 wire \Tile_X9Y6_W2BEG[5] ;
 wire \Tile_X9Y6_W2BEG[6] ;
 wire \Tile_X9Y6_W2BEG[7] ;
 wire \Tile_X9Y6_W2BEGb[0] ;
 wire \Tile_X9Y6_W2BEGb[1] ;
 wire \Tile_X9Y6_W2BEGb[2] ;
 wire \Tile_X9Y6_W2BEGb[3] ;
 wire \Tile_X9Y6_W2BEGb[4] ;
 wire \Tile_X9Y6_W2BEGb[5] ;
 wire \Tile_X9Y6_W2BEGb[6] ;
 wire \Tile_X9Y6_W2BEGb[7] ;
 wire \Tile_X9Y6_W6BEG[0] ;
 wire \Tile_X9Y6_W6BEG[10] ;
 wire \Tile_X9Y6_W6BEG[11] ;
 wire \Tile_X9Y6_W6BEG[1] ;
 wire \Tile_X9Y6_W6BEG[2] ;
 wire \Tile_X9Y6_W6BEG[3] ;
 wire \Tile_X9Y6_W6BEG[4] ;
 wire \Tile_X9Y6_W6BEG[5] ;
 wire \Tile_X9Y6_W6BEG[6] ;
 wire \Tile_X9Y6_W6BEG[7] ;
 wire \Tile_X9Y6_W6BEG[8] ;
 wire \Tile_X9Y6_W6BEG[9] ;
 wire \Tile_X9Y6_WW4BEG[0] ;
 wire \Tile_X9Y6_WW4BEG[10] ;
 wire \Tile_X9Y6_WW4BEG[11] ;
 wire \Tile_X9Y6_WW4BEG[12] ;
 wire \Tile_X9Y6_WW4BEG[13] ;
 wire \Tile_X9Y6_WW4BEG[14] ;
 wire \Tile_X9Y6_WW4BEG[15] ;
 wire \Tile_X9Y6_WW4BEG[1] ;
 wire \Tile_X9Y6_WW4BEG[2] ;
 wire \Tile_X9Y6_WW4BEG[3] ;
 wire \Tile_X9Y6_WW4BEG[4] ;
 wire \Tile_X9Y6_WW4BEG[5] ;
 wire \Tile_X9Y6_WW4BEG[6] ;
 wire \Tile_X9Y6_WW4BEG[7] ;
 wire \Tile_X9Y6_WW4BEG[8] ;
 wire \Tile_X9Y6_WW4BEG[9] ;
 wire Tile_X9Y7_Co;
 wire \Tile_X9Y7_E1BEG[0] ;
 wire \Tile_X9Y7_E1BEG[1] ;
 wire \Tile_X9Y7_E1BEG[2] ;
 wire \Tile_X9Y7_E1BEG[3] ;
 wire \Tile_X9Y7_E2BEG[0] ;
 wire \Tile_X9Y7_E2BEG[1] ;
 wire \Tile_X9Y7_E2BEG[2] ;
 wire \Tile_X9Y7_E2BEG[3] ;
 wire \Tile_X9Y7_E2BEG[4] ;
 wire \Tile_X9Y7_E2BEG[5] ;
 wire \Tile_X9Y7_E2BEG[6] ;
 wire \Tile_X9Y7_E2BEG[7] ;
 wire \Tile_X9Y7_E2BEGb[0] ;
 wire \Tile_X9Y7_E2BEGb[1] ;
 wire \Tile_X9Y7_E2BEGb[2] ;
 wire \Tile_X9Y7_E2BEGb[3] ;
 wire \Tile_X9Y7_E2BEGb[4] ;
 wire \Tile_X9Y7_E2BEGb[5] ;
 wire \Tile_X9Y7_E2BEGb[6] ;
 wire \Tile_X9Y7_E2BEGb[7] ;
 wire \Tile_X9Y7_E6BEG[0] ;
 wire \Tile_X9Y7_E6BEG[10] ;
 wire \Tile_X9Y7_E6BEG[11] ;
 wire \Tile_X9Y7_E6BEG[1] ;
 wire \Tile_X9Y7_E6BEG[2] ;
 wire \Tile_X9Y7_E6BEG[3] ;
 wire \Tile_X9Y7_E6BEG[4] ;
 wire \Tile_X9Y7_E6BEG[5] ;
 wire \Tile_X9Y7_E6BEG[6] ;
 wire \Tile_X9Y7_E6BEG[7] ;
 wire \Tile_X9Y7_E6BEG[8] ;
 wire \Tile_X9Y7_E6BEG[9] ;
 wire \Tile_X9Y7_EE4BEG[0] ;
 wire \Tile_X9Y7_EE4BEG[10] ;
 wire \Tile_X9Y7_EE4BEG[11] ;
 wire \Tile_X9Y7_EE4BEG[12] ;
 wire \Tile_X9Y7_EE4BEG[13] ;
 wire \Tile_X9Y7_EE4BEG[14] ;
 wire \Tile_X9Y7_EE4BEG[15] ;
 wire \Tile_X9Y7_EE4BEG[1] ;
 wire \Tile_X9Y7_EE4BEG[2] ;
 wire \Tile_X9Y7_EE4BEG[3] ;
 wire \Tile_X9Y7_EE4BEG[4] ;
 wire \Tile_X9Y7_EE4BEG[5] ;
 wire \Tile_X9Y7_EE4BEG[6] ;
 wire \Tile_X9Y7_EE4BEG[7] ;
 wire \Tile_X9Y7_EE4BEG[8] ;
 wire \Tile_X9Y7_EE4BEG[9] ;
 wire \Tile_X9Y7_FrameData_O[0] ;
 wire \Tile_X9Y7_FrameData_O[10] ;
 wire \Tile_X9Y7_FrameData_O[11] ;
 wire \Tile_X9Y7_FrameData_O[12] ;
 wire \Tile_X9Y7_FrameData_O[13] ;
 wire \Tile_X9Y7_FrameData_O[14] ;
 wire \Tile_X9Y7_FrameData_O[15] ;
 wire \Tile_X9Y7_FrameData_O[16] ;
 wire \Tile_X9Y7_FrameData_O[17] ;
 wire \Tile_X9Y7_FrameData_O[18] ;
 wire \Tile_X9Y7_FrameData_O[19] ;
 wire \Tile_X9Y7_FrameData_O[1] ;
 wire \Tile_X9Y7_FrameData_O[20] ;
 wire \Tile_X9Y7_FrameData_O[21] ;
 wire \Tile_X9Y7_FrameData_O[22] ;
 wire \Tile_X9Y7_FrameData_O[23] ;
 wire \Tile_X9Y7_FrameData_O[24] ;
 wire \Tile_X9Y7_FrameData_O[25] ;
 wire \Tile_X9Y7_FrameData_O[26] ;
 wire \Tile_X9Y7_FrameData_O[27] ;
 wire \Tile_X9Y7_FrameData_O[28] ;
 wire \Tile_X9Y7_FrameData_O[29] ;
 wire \Tile_X9Y7_FrameData_O[2] ;
 wire \Tile_X9Y7_FrameData_O[30] ;
 wire \Tile_X9Y7_FrameData_O[31] ;
 wire \Tile_X9Y7_FrameData_O[3] ;
 wire \Tile_X9Y7_FrameData_O[4] ;
 wire \Tile_X9Y7_FrameData_O[5] ;
 wire \Tile_X9Y7_FrameData_O[6] ;
 wire \Tile_X9Y7_FrameData_O[7] ;
 wire \Tile_X9Y7_FrameData_O[8] ;
 wire \Tile_X9Y7_FrameData_O[9] ;
 wire \Tile_X9Y7_FrameStrobe_O[0] ;
 wire \Tile_X9Y7_FrameStrobe_O[10] ;
 wire \Tile_X9Y7_FrameStrobe_O[11] ;
 wire \Tile_X9Y7_FrameStrobe_O[12] ;
 wire \Tile_X9Y7_FrameStrobe_O[13] ;
 wire \Tile_X9Y7_FrameStrobe_O[14] ;
 wire \Tile_X9Y7_FrameStrobe_O[15] ;
 wire \Tile_X9Y7_FrameStrobe_O[16] ;
 wire \Tile_X9Y7_FrameStrobe_O[17] ;
 wire \Tile_X9Y7_FrameStrobe_O[18] ;
 wire \Tile_X9Y7_FrameStrobe_O[19] ;
 wire \Tile_X9Y7_FrameStrobe_O[1] ;
 wire \Tile_X9Y7_FrameStrobe_O[2] ;
 wire \Tile_X9Y7_FrameStrobe_O[3] ;
 wire \Tile_X9Y7_FrameStrobe_O[4] ;
 wire \Tile_X9Y7_FrameStrobe_O[5] ;
 wire \Tile_X9Y7_FrameStrobe_O[6] ;
 wire \Tile_X9Y7_FrameStrobe_O[7] ;
 wire \Tile_X9Y7_FrameStrobe_O[8] ;
 wire \Tile_X9Y7_FrameStrobe_O[9] ;
 wire \Tile_X9Y7_N1BEG[0] ;
 wire \Tile_X9Y7_N1BEG[1] ;
 wire \Tile_X9Y7_N1BEG[2] ;
 wire \Tile_X9Y7_N1BEG[3] ;
 wire \Tile_X9Y7_N2BEG[0] ;
 wire \Tile_X9Y7_N2BEG[1] ;
 wire \Tile_X9Y7_N2BEG[2] ;
 wire \Tile_X9Y7_N2BEG[3] ;
 wire \Tile_X9Y7_N2BEG[4] ;
 wire \Tile_X9Y7_N2BEG[5] ;
 wire \Tile_X9Y7_N2BEG[6] ;
 wire \Tile_X9Y7_N2BEG[7] ;
 wire \Tile_X9Y7_N2BEGb[0] ;
 wire \Tile_X9Y7_N2BEGb[1] ;
 wire \Tile_X9Y7_N2BEGb[2] ;
 wire \Tile_X9Y7_N2BEGb[3] ;
 wire \Tile_X9Y7_N2BEGb[4] ;
 wire \Tile_X9Y7_N2BEGb[5] ;
 wire \Tile_X9Y7_N2BEGb[6] ;
 wire \Tile_X9Y7_N2BEGb[7] ;
 wire \Tile_X9Y7_N4BEG[0] ;
 wire \Tile_X9Y7_N4BEG[10] ;
 wire \Tile_X9Y7_N4BEG[11] ;
 wire \Tile_X9Y7_N4BEG[12] ;
 wire \Tile_X9Y7_N4BEG[13] ;
 wire \Tile_X9Y7_N4BEG[14] ;
 wire \Tile_X9Y7_N4BEG[15] ;
 wire \Tile_X9Y7_N4BEG[1] ;
 wire \Tile_X9Y7_N4BEG[2] ;
 wire \Tile_X9Y7_N4BEG[3] ;
 wire \Tile_X9Y7_N4BEG[4] ;
 wire \Tile_X9Y7_N4BEG[5] ;
 wire \Tile_X9Y7_N4BEG[6] ;
 wire \Tile_X9Y7_N4BEG[7] ;
 wire \Tile_X9Y7_N4BEG[8] ;
 wire \Tile_X9Y7_N4BEG[9] ;
 wire \Tile_X9Y7_NN4BEG[0] ;
 wire \Tile_X9Y7_NN4BEG[10] ;
 wire \Tile_X9Y7_NN4BEG[11] ;
 wire \Tile_X9Y7_NN4BEG[12] ;
 wire \Tile_X9Y7_NN4BEG[13] ;
 wire \Tile_X9Y7_NN4BEG[14] ;
 wire \Tile_X9Y7_NN4BEG[15] ;
 wire \Tile_X9Y7_NN4BEG[1] ;
 wire \Tile_X9Y7_NN4BEG[2] ;
 wire \Tile_X9Y7_NN4BEG[3] ;
 wire \Tile_X9Y7_NN4BEG[4] ;
 wire \Tile_X9Y7_NN4BEG[5] ;
 wire \Tile_X9Y7_NN4BEG[6] ;
 wire \Tile_X9Y7_NN4BEG[7] ;
 wire \Tile_X9Y7_NN4BEG[8] ;
 wire \Tile_X9Y7_NN4BEG[9] ;
 wire \Tile_X9Y7_S1BEG[0] ;
 wire \Tile_X9Y7_S1BEG[1] ;
 wire \Tile_X9Y7_S1BEG[2] ;
 wire \Tile_X9Y7_S1BEG[3] ;
 wire \Tile_X9Y7_S2BEG[0] ;
 wire \Tile_X9Y7_S2BEG[1] ;
 wire \Tile_X9Y7_S2BEG[2] ;
 wire \Tile_X9Y7_S2BEG[3] ;
 wire \Tile_X9Y7_S2BEG[4] ;
 wire \Tile_X9Y7_S2BEG[5] ;
 wire \Tile_X9Y7_S2BEG[6] ;
 wire \Tile_X9Y7_S2BEG[7] ;
 wire \Tile_X9Y7_S2BEGb[0] ;
 wire \Tile_X9Y7_S2BEGb[1] ;
 wire \Tile_X9Y7_S2BEGb[2] ;
 wire \Tile_X9Y7_S2BEGb[3] ;
 wire \Tile_X9Y7_S2BEGb[4] ;
 wire \Tile_X9Y7_S2BEGb[5] ;
 wire \Tile_X9Y7_S2BEGb[6] ;
 wire \Tile_X9Y7_S2BEGb[7] ;
 wire \Tile_X9Y7_S4BEG[0] ;
 wire \Tile_X9Y7_S4BEG[10] ;
 wire \Tile_X9Y7_S4BEG[11] ;
 wire \Tile_X9Y7_S4BEG[12] ;
 wire \Tile_X9Y7_S4BEG[13] ;
 wire \Tile_X9Y7_S4BEG[14] ;
 wire \Tile_X9Y7_S4BEG[15] ;
 wire \Tile_X9Y7_S4BEG[1] ;
 wire \Tile_X9Y7_S4BEG[2] ;
 wire \Tile_X9Y7_S4BEG[3] ;
 wire \Tile_X9Y7_S4BEG[4] ;
 wire \Tile_X9Y7_S4BEG[5] ;
 wire \Tile_X9Y7_S4BEG[6] ;
 wire \Tile_X9Y7_S4BEG[7] ;
 wire \Tile_X9Y7_S4BEG[8] ;
 wire \Tile_X9Y7_S4BEG[9] ;
 wire \Tile_X9Y7_SS4BEG[0] ;
 wire \Tile_X9Y7_SS4BEG[10] ;
 wire \Tile_X9Y7_SS4BEG[11] ;
 wire \Tile_X9Y7_SS4BEG[12] ;
 wire \Tile_X9Y7_SS4BEG[13] ;
 wire \Tile_X9Y7_SS4BEG[14] ;
 wire \Tile_X9Y7_SS4BEG[15] ;
 wire \Tile_X9Y7_SS4BEG[1] ;
 wire \Tile_X9Y7_SS4BEG[2] ;
 wire \Tile_X9Y7_SS4BEG[3] ;
 wire \Tile_X9Y7_SS4BEG[4] ;
 wire \Tile_X9Y7_SS4BEG[5] ;
 wire \Tile_X9Y7_SS4BEG[6] ;
 wire \Tile_X9Y7_SS4BEG[7] ;
 wire \Tile_X9Y7_SS4BEG[8] ;
 wire \Tile_X9Y7_SS4BEG[9] ;
 wire Tile_X9Y7_UserCLKo;
 wire \Tile_X9Y7_W1BEG[0] ;
 wire \Tile_X9Y7_W1BEG[1] ;
 wire \Tile_X9Y7_W1BEG[2] ;
 wire \Tile_X9Y7_W1BEG[3] ;
 wire \Tile_X9Y7_W2BEG[0] ;
 wire \Tile_X9Y7_W2BEG[1] ;
 wire \Tile_X9Y7_W2BEG[2] ;
 wire \Tile_X9Y7_W2BEG[3] ;
 wire \Tile_X9Y7_W2BEG[4] ;
 wire \Tile_X9Y7_W2BEG[5] ;
 wire \Tile_X9Y7_W2BEG[6] ;
 wire \Tile_X9Y7_W2BEG[7] ;
 wire \Tile_X9Y7_W2BEGb[0] ;
 wire \Tile_X9Y7_W2BEGb[1] ;
 wire \Tile_X9Y7_W2BEGb[2] ;
 wire \Tile_X9Y7_W2BEGb[3] ;
 wire \Tile_X9Y7_W2BEGb[4] ;
 wire \Tile_X9Y7_W2BEGb[5] ;
 wire \Tile_X9Y7_W2BEGb[6] ;
 wire \Tile_X9Y7_W2BEGb[7] ;
 wire \Tile_X9Y7_W6BEG[0] ;
 wire \Tile_X9Y7_W6BEG[10] ;
 wire \Tile_X9Y7_W6BEG[11] ;
 wire \Tile_X9Y7_W6BEG[1] ;
 wire \Tile_X9Y7_W6BEG[2] ;
 wire \Tile_X9Y7_W6BEG[3] ;
 wire \Tile_X9Y7_W6BEG[4] ;
 wire \Tile_X9Y7_W6BEG[5] ;
 wire \Tile_X9Y7_W6BEG[6] ;
 wire \Tile_X9Y7_W6BEG[7] ;
 wire \Tile_X9Y7_W6BEG[8] ;
 wire \Tile_X9Y7_W6BEG[9] ;
 wire \Tile_X9Y7_WW4BEG[0] ;
 wire \Tile_X9Y7_WW4BEG[10] ;
 wire \Tile_X9Y7_WW4BEG[11] ;
 wire \Tile_X9Y7_WW4BEG[12] ;
 wire \Tile_X9Y7_WW4BEG[13] ;
 wire \Tile_X9Y7_WW4BEG[14] ;
 wire \Tile_X9Y7_WW4BEG[15] ;
 wire \Tile_X9Y7_WW4BEG[1] ;
 wire \Tile_X9Y7_WW4BEG[2] ;
 wire \Tile_X9Y7_WW4BEG[3] ;
 wire \Tile_X9Y7_WW4BEG[4] ;
 wire \Tile_X9Y7_WW4BEG[5] ;
 wire \Tile_X9Y7_WW4BEG[6] ;
 wire \Tile_X9Y7_WW4BEG[7] ;
 wire \Tile_X9Y7_WW4BEG[8] ;
 wire \Tile_X9Y7_WW4BEG[9] ;
 wire Tile_X9Y8_Co;
 wire \Tile_X9Y8_E1BEG[0] ;
 wire \Tile_X9Y8_E1BEG[1] ;
 wire \Tile_X9Y8_E1BEG[2] ;
 wire \Tile_X9Y8_E1BEG[3] ;
 wire \Tile_X9Y8_E2BEG[0] ;
 wire \Tile_X9Y8_E2BEG[1] ;
 wire \Tile_X9Y8_E2BEG[2] ;
 wire \Tile_X9Y8_E2BEG[3] ;
 wire \Tile_X9Y8_E2BEG[4] ;
 wire \Tile_X9Y8_E2BEG[5] ;
 wire \Tile_X9Y8_E2BEG[6] ;
 wire \Tile_X9Y8_E2BEG[7] ;
 wire \Tile_X9Y8_E2BEGb[0] ;
 wire \Tile_X9Y8_E2BEGb[1] ;
 wire \Tile_X9Y8_E2BEGb[2] ;
 wire \Tile_X9Y8_E2BEGb[3] ;
 wire \Tile_X9Y8_E2BEGb[4] ;
 wire \Tile_X9Y8_E2BEGb[5] ;
 wire \Tile_X9Y8_E2BEGb[6] ;
 wire \Tile_X9Y8_E2BEGb[7] ;
 wire \Tile_X9Y8_E6BEG[0] ;
 wire \Tile_X9Y8_E6BEG[10] ;
 wire \Tile_X9Y8_E6BEG[11] ;
 wire \Tile_X9Y8_E6BEG[1] ;
 wire \Tile_X9Y8_E6BEG[2] ;
 wire \Tile_X9Y8_E6BEG[3] ;
 wire \Tile_X9Y8_E6BEG[4] ;
 wire \Tile_X9Y8_E6BEG[5] ;
 wire \Tile_X9Y8_E6BEG[6] ;
 wire \Tile_X9Y8_E6BEG[7] ;
 wire \Tile_X9Y8_E6BEG[8] ;
 wire \Tile_X9Y8_E6BEG[9] ;
 wire \Tile_X9Y8_EE4BEG[0] ;
 wire \Tile_X9Y8_EE4BEG[10] ;
 wire \Tile_X9Y8_EE4BEG[11] ;
 wire \Tile_X9Y8_EE4BEG[12] ;
 wire \Tile_X9Y8_EE4BEG[13] ;
 wire \Tile_X9Y8_EE4BEG[14] ;
 wire \Tile_X9Y8_EE4BEG[15] ;
 wire \Tile_X9Y8_EE4BEG[1] ;
 wire \Tile_X9Y8_EE4BEG[2] ;
 wire \Tile_X9Y8_EE4BEG[3] ;
 wire \Tile_X9Y8_EE4BEG[4] ;
 wire \Tile_X9Y8_EE4BEG[5] ;
 wire \Tile_X9Y8_EE4BEG[6] ;
 wire \Tile_X9Y8_EE4BEG[7] ;
 wire \Tile_X9Y8_EE4BEG[8] ;
 wire \Tile_X9Y8_EE4BEG[9] ;
 wire \Tile_X9Y8_FrameData_O[0] ;
 wire \Tile_X9Y8_FrameData_O[10] ;
 wire \Tile_X9Y8_FrameData_O[11] ;
 wire \Tile_X9Y8_FrameData_O[12] ;
 wire \Tile_X9Y8_FrameData_O[13] ;
 wire \Tile_X9Y8_FrameData_O[14] ;
 wire \Tile_X9Y8_FrameData_O[15] ;
 wire \Tile_X9Y8_FrameData_O[16] ;
 wire \Tile_X9Y8_FrameData_O[17] ;
 wire \Tile_X9Y8_FrameData_O[18] ;
 wire \Tile_X9Y8_FrameData_O[19] ;
 wire \Tile_X9Y8_FrameData_O[1] ;
 wire \Tile_X9Y8_FrameData_O[20] ;
 wire \Tile_X9Y8_FrameData_O[21] ;
 wire \Tile_X9Y8_FrameData_O[22] ;
 wire \Tile_X9Y8_FrameData_O[23] ;
 wire \Tile_X9Y8_FrameData_O[24] ;
 wire \Tile_X9Y8_FrameData_O[25] ;
 wire \Tile_X9Y8_FrameData_O[26] ;
 wire \Tile_X9Y8_FrameData_O[27] ;
 wire \Tile_X9Y8_FrameData_O[28] ;
 wire \Tile_X9Y8_FrameData_O[29] ;
 wire \Tile_X9Y8_FrameData_O[2] ;
 wire \Tile_X9Y8_FrameData_O[30] ;
 wire \Tile_X9Y8_FrameData_O[31] ;
 wire \Tile_X9Y8_FrameData_O[3] ;
 wire \Tile_X9Y8_FrameData_O[4] ;
 wire \Tile_X9Y8_FrameData_O[5] ;
 wire \Tile_X9Y8_FrameData_O[6] ;
 wire \Tile_X9Y8_FrameData_O[7] ;
 wire \Tile_X9Y8_FrameData_O[8] ;
 wire \Tile_X9Y8_FrameData_O[9] ;
 wire \Tile_X9Y8_FrameStrobe_O[0] ;
 wire \Tile_X9Y8_FrameStrobe_O[10] ;
 wire \Tile_X9Y8_FrameStrobe_O[11] ;
 wire \Tile_X9Y8_FrameStrobe_O[12] ;
 wire \Tile_X9Y8_FrameStrobe_O[13] ;
 wire \Tile_X9Y8_FrameStrobe_O[14] ;
 wire \Tile_X9Y8_FrameStrobe_O[15] ;
 wire \Tile_X9Y8_FrameStrobe_O[16] ;
 wire \Tile_X9Y8_FrameStrobe_O[17] ;
 wire \Tile_X9Y8_FrameStrobe_O[18] ;
 wire \Tile_X9Y8_FrameStrobe_O[19] ;
 wire \Tile_X9Y8_FrameStrobe_O[1] ;
 wire \Tile_X9Y8_FrameStrobe_O[2] ;
 wire \Tile_X9Y8_FrameStrobe_O[3] ;
 wire \Tile_X9Y8_FrameStrobe_O[4] ;
 wire \Tile_X9Y8_FrameStrobe_O[5] ;
 wire \Tile_X9Y8_FrameStrobe_O[6] ;
 wire \Tile_X9Y8_FrameStrobe_O[7] ;
 wire \Tile_X9Y8_FrameStrobe_O[8] ;
 wire \Tile_X9Y8_FrameStrobe_O[9] ;
 wire \Tile_X9Y8_N1BEG[0] ;
 wire \Tile_X9Y8_N1BEG[1] ;
 wire \Tile_X9Y8_N1BEG[2] ;
 wire \Tile_X9Y8_N1BEG[3] ;
 wire \Tile_X9Y8_N2BEG[0] ;
 wire \Tile_X9Y8_N2BEG[1] ;
 wire \Tile_X9Y8_N2BEG[2] ;
 wire \Tile_X9Y8_N2BEG[3] ;
 wire \Tile_X9Y8_N2BEG[4] ;
 wire \Tile_X9Y8_N2BEG[5] ;
 wire \Tile_X9Y8_N2BEG[6] ;
 wire \Tile_X9Y8_N2BEG[7] ;
 wire \Tile_X9Y8_N2BEGb[0] ;
 wire \Tile_X9Y8_N2BEGb[1] ;
 wire \Tile_X9Y8_N2BEGb[2] ;
 wire \Tile_X9Y8_N2BEGb[3] ;
 wire \Tile_X9Y8_N2BEGb[4] ;
 wire \Tile_X9Y8_N2BEGb[5] ;
 wire \Tile_X9Y8_N2BEGb[6] ;
 wire \Tile_X9Y8_N2BEGb[7] ;
 wire \Tile_X9Y8_N4BEG[0] ;
 wire \Tile_X9Y8_N4BEG[10] ;
 wire \Tile_X9Y8_N4BEG[11] ;
 wire \Tile_X9Y8_N4BEG[12] ;
 wire \Tile_X9Y8_N4BEG[13] ;
 wire \Tile_X9Y8_N4BEG[14] ;
 wire \Tile_X9Y8_N4BEG[15] ;
 wire \Tile_X9Y8_N4BEG[1] ;
 wire \Tile_X9Y8_N4BEG[2] ;
 wire \Tile_X9Y8_N4BEG[3] ;
 wire \Tile_X9Y8_N4BEG[4] ;
 wire \Tile_X9Y8_N4BEG[5] ;
 wire \Tile_X9Y8_N4BEG[6] ;
 wire \Tile_X9Y8_N4BEG[7] ;
 wire \Tile_X9Y8_N4BEG[8] ;
 wire \Tile_X9Y8_N4BEG[9] ;
 wire \Tile_X9Y8_NN4BEG[0] ;
 wire \Tile_X9Y8_NN4BEG[10] ;
 wire \Tile_X9Y8_NN4BEG[11] ;
 wire \Tile_X9Y8_NN4BEG[12] ;
 wire \Tile_X9Y8_NN4BEG[13] ;
 wire \Tile_X9Y8_NN4BEG[14] ;
 wire \Tile_X9Y8_NN4BEG[15] ;
 wire \Tile_X9Y8_NN4BEG[1] ;
 wire \Tile_X9Y8_NN4BEG[2] ;
 wire \Tile_X9Y8_NN4BEG[3] ;
 wire \Tile_X9Y8_NN4BEG[4] ;
 wire \Tile_X9Y8_NN4BEG[5] ;
 wire \Tile_X9Y8_NN4BEG[6] ;
 wire \Tile_X9Y8_NN4BEG[7] ;
 wire \Tile_X9Y8_NN4BEG[8] ;
 wire \Tile_X9Y8_NN4BEG[9] ;
 wire \Tile_X9Y8_S1BEG[0] ;
 wire \Tile_X9Y8_S1BEG[1] ;
 wire \Tile_X9Y8_S1BEG[2] ;
 wire \Tile_X9Y8_S1BEG[3] ;
 wire \Tile_X9Y8_S2BEG[0] ;
 wire \Tile_X9Y8_S2BEG[1] ;
 wire \Tile_X9Y8_S2BEG[2] ;
 wire \Tile_X9Y8_S2BEG[3] ;
 wire \Tile_X9Y8_S2BEG[4] ;
 wire \Tile_X9Y8_S2BEG[5] ;
 wire \Tile_X9Y8_S2BEG[6] ;
 wire \Tile_X9Y8_S2BEG[7] ;
 wire \Tile_X9Y8_S2BEGb[0] ;
 wire \Tile_X9Y8_S2BEGb[1] ;
 wire \Tile_X9Y8_S2BEGb[2] ;
 wire \Tile_X9Y8_S2BEGb[3] ;
 wire \Tile_X9Y8_S2BEGb[4] ;
 wire \Tile_X9Y8_S2BEGb[5] ;
 wire \Tile_X9Y8_S2BEGb[6] ;
 wire \Tile_X9Y8_S2BEGb[7] ;
 wire \Tile_X9Y8_S4BEG[0] ;
 wire \Tile_X9Y8_S4BEG[10] ;
 wire \Tile_X9Y8_S4BEG[11] ;
 wire \Tile_X9Y8_S4BEG[12] ;
 wire \Tile_X9Y8_S4BEG[13] ;
 wire \Tile_X9Y8_S4BEG[14] ;
 wire \Tile_X9Y8_S4BEG[15] ;
 wire \Tile_X9Y8_S4BEG[1] ;
 wire \Tile_X9Y8_S4BEG[2] ;
 wire \Tile_X9Y8_S4BEG[3] ;
 wire \Tile_X9Y8_S4BEG[4] ;
 wire \Tile_X9Y8_S4BEG[5] ;
 wire \Tile_X9Y8_S4BEG[6] ;
 wire \Tile_X9Y8_S4BEG[7] ;
 wire \Tile_X9Y8_S4BEG[8] ;
 wire \Tile_X9Y8_S4BEG[9] ;
 wire \Tile_X9Y8_SS4BEG[0] ;
 wire \Tile_X9Y8_SS4BEG[10] ;
 wire \Tile_X9Y8_SS4BEG[11] ;
 wire \Tile_X9Y8_SS4BEG[12] ;
 wire \Tile_X9Y8_SS4BEG[13] ;
 wire \Tile_X9Y8_SS4BEG[14] ;
 wire \Tile_X9Y8_SS4BEG[15] ;
 wire \Tile_X9Y8_SS4BEG[1] ;
 wire \Tile_X9Y8_SS4BEG[2] ;
 wire \Tile_X9Y8_SS4BEG[3] ;
 wire \Tile_X9Y8_SS4BEG[4] ;
 wire \Tile_X9Y8_SS4BEG[5] ;
 wire \Tile_X9Y8_SS4BEG[6] ;
 wire \Tile_X9Y8_SS4BEG[7] ;
 wire \Tile_X9Y8_SS4BEG[8] ;
 wire \Tile_X9Y8_SS4BEG[9] ;
 wire Tile_X9Y8_UserCLKo;
 wire \Tile_X9Y8_W1BEG[0] ;
 wire \Tile_X9Y8_W1BEG[1] ;
 wire \Tile_X9Y8_W1BEG[2] ;
 wire \Tile_X9Y8_W1BEG[3] ;
 wire \Tile_X9Y8_W2BEG[0] ;
 wire \Tile_X9Y8_W2BEG[1] ;
 wire \Tile_X9Y8_W2BEG[2] ;
 wire \Tile_X9Y8_W2BEG[3] ;
 wire \Tile_X9Y8_W2BEG[4] ;
 wire \Tile_X9Y8_W2BEG[5] ;
 wire \Tile_X9Y8_W2BEG[6] ;
 wire \Tile_X9Y8_W2BEG[7] ;
 wire \Tile_X9Y8_W2BEGb[0] ;
 wire \Tile_X9Y8_W2BEGb[1] ;
 wire \Tile_X9Y8_W2BEGb[2] ;
 wire \Tile_X9Y8_W2BEGb[3] ;
 wire \Tile_X9Y8_W2BEGb[4] ;
 wire \Tile_X9Y8_W2BEGb[5] ;
 wire \Tile_X9Y8_W2BEGb[6] ;
 wire \Tile_X9Y8_W2BEGb[7] ;
 wire \Tile_X9Y8_W6BEG[0] ;
 wire \Tile_X9Y8_W6BEG[10] ;
 wire \Tile_X9Y8_W6BEG[11] ;
 wire \Tile_X9Y8_W6BEG[1] ;
 wire \Tile_X9Y8_W6BEG[2] ;
 wire \Tile_X9Y8_W6BEG[3] ;
 wire \Tile_X9Y8_W6BEG[4] ;
 wire \Tile_X9Y8_W6BEG[5] ;
 wire \Tile_X9Y8_W6BEG[6] ;
 wire \Tile_X9Y8_W6BEG[7] ;
 wire \Tile_X9Y8_W6BEG[8] ;
 wire \Tile_X9Y8_W6BEG[9] ;
 wire \Tile_X9Y8_WW4BEG[0] ;
 wire \Tile_X9Y8_WW4BEG[10] ;
 wire \Tile_X9Y8_WW4BEG[11] ;
 wire \Tile_X9Y8_WW4BEG[12] ;
 wire \Tile_X9Y8_WW4BEG[13] ;
 wire \Tile_X9Y8_WW4BEG[14] ;
 wire \Tile_X9Y8_WW4BEG[15] ;
 wire \Tile_X9Y8_WW4BEG[1] ;
 wire \Tile_X9Y8_WW4BEG[2] ;
 wire \Tile_X9Y8_WW4BEG[3] ;
 wire \Tile_X9Y8_WW4BEG[4] ;
 wire \Tile_X9Y8_WW4BEG[5] ;
 wire \Tile_X9Y8_WW4BEG[6] ;
 wire \Tile_X9Y8_WW4BEG[7] ;
 wire \Tile_X9Y8_WW4BEG[8] ;
 wire \Tile_X9Y8_WW4BEG[9] ;
 wire Tile_X9Y9_Co;
 wire \Tile_X9Y9_E1BEG[0] ;
 wire \Tile_X9Y9_E1BEG[1] ;
 wire \Tile_X9Y9_E1BEG[2] ;
 wire \Tile_X9Y9_E1BEG[3] ;
 wire \Tile_X9Y9_E2BEG[0] ;
 wire \Tile_X9Y9_E2BEG[1] ;
 wire \Tile_X9Y9_E2BEG[2] ;
 wire \Tile_X9Y9_E2BEG[3] ;
 wire \Tile_X9Y9_E2BEG[4] ;
 wire \Tile_X9Y9_E2BEG[5] ;
 wire \Tile_X9Y9_E2BEG[6] ;
 wire \Tile_X9Y9_E2BEG[7] ;
 wire \Tile_X9Y9_E2BEGb[0] ;
 wire \Tile_X9Y9_E2BEGb[1] ;
 wire \Tile_X9Y9_E2BEGb[2] ;
 wire \Tile_X9Y9_E2BEGb[3] ;
 wire \Tile_X9Y9_E2BEGb[4] ;
 wire \Tile_X9Y9_E2BEGb[5] ;
 wire \Tile_X9Y9_E2BEGb[6] ;
 wire \Tile_X9Y9_E2BEGb[7] ;
 wire \Tile_X9Y9_E6BEG[0] ;
 wire \Tile_X9Y9_E6BEG[10] ;
 wire \Tile_X9Y9_E6BEG[11] ;
 wire \Tile_X9Y9_E6BEG[1] ;
 wire \Tile_X9Y9_E6BEG[2] ;
 wire \Tile_X9Y9_E6BEG[3] ;
 wire \Tile_X9Y9_E6BEG[4] ;
 wire \Tile_X9Y9_E6BEG[5] ;
 wire \Tile_X9Y9_E6BEG[6] ;
 wire \Tile_X9Y9_E6BEG[7] ;
 wire \Tile_X9Y9_E6BEG[8] ;
 wire \Tile_X9Y9_E6BEG[9] ;
 wire \Tile_X9Y9_EE4BEG[0] ;
 wire \Tile_X9Y9_EE4BEG[10] ;
 wire \Tile_X9Y9_EE4BEG[11] ;
 wire \Tile_X9Y9_EE4BEG[12] ;
 wire \Tile_X9Y9_EE4BEG[13] ;
 wire \Tile_X9Y9_EE4BEG[14] ;
 wire \Tile_X9Y9_EE4BEG[15] ;
 wire \Tile_X9Y9_EE4BEG[1] ;
 wire \Tile_X9Y9_EE4BEG[2] ;
 wire \Tile_X9Y9_EE4BEG[3] ;
 wire \Tile_X9Y9_EE4BEG[4] ;
 wire \Tile_X9Y9_EE4BEG[5] ;
 wire \Tile_X9Y9_EE4BEG[6] ;
 wire \Tile_X9Y9_EE4BEG[7] ;
 wire \Tile_X9Y9_EE4BEG[8] ;
 wire \Tile_X9Y9_EE4BEG[9] ;
 wire \Tile_X9Y9_FrameData_O[0] ;
 wire \Tile_X9Y9_FrameData_O[10] ;
 wire \Tile_X9Y9_FrameData_O[11] ;
 wire \Tile_X9Y9_FrameData_O[12] ;
 wire \Tile_X9Y9_FrameData_O[13] ;
 wire \Tile_X9Y9_FrameData_O[14] ;
 wire \Tile_X9Y9_FrameData_O[15] ;
 wire \Tile_X9Y9_FrameData_O[16] ;
 wire \Tile_X9Y9_FrameData_O[17] ;
 wire \Tile_X9Y9_FrameData_O[18] ;
 wire \Tile_X9Y9_FrameData_O[19] ;
 wire \Tile_X9Y9_FrameData_O[1] ;
 wire \Tile_X9Y9_FrameData_O[20] ;
 wire \Tile_X9Y9_FrameData_O[21] ;
 wire \Tile_X9Y9_FrameData_O[22] ;
 wire \Tile_X9Y9_FrameData_O[23] ;
 wire \Tile_X9Y9_FrameData_O[24] ;
 wire \Tile_X9Y9_FrameData_O[25] ;
 wire \Tile_X9Y9_FrameData_O[26] ;
 wire \Tile_X9Y9_FrameData_O[27] ;
 wire \Tile_X9Y9_FrameData_O[28] ;
 wire \Tile_X9Y9_FrameData_O[29] ;
 wire \Tile_X9Y9_FrameData_O[2] ;
 wire \Tile_X9Y9_FrameData_O[30] ;
 wire \Tile_X9Y9_FrameData_O[31] ;
 wire \Tile_X9Y9_FrameData_O[3] ;
 wire \Tile_X9Y9_FrameData_O[4] ;
 wire \Tile_X9Y9_FrameData_O[5] ;
 wire \Tile_X9Y9_FrameData_O[6] ;
 wire \Tile_X9Y9_FrameData_O[7] ;
 wire \Tile_X9Y9_FrameData_O[8] ;
 wire \Tile_X9Y9_FrameData_O[9] ;
 wire \Tile_X9Y9_FrameStrobe_O[0] ;
 wire \Tile_X9Y9_FrameStrobe_O[10] ;
 wire \Tile_X9Y9_FrameStrobe_O[11] ;
 wire \Tile_X9Y9_FrameStrobe_O[12] ;
 wire \Tile_X9Y9_FrameStrobe_O[13] ;
 wire \Tile_X9Y9_FrameStrobe_O[14] ;
 wire \Tile_X9Y9_FrameStrobe_O[15] ;
 wire \Tile_X9Y9_FrameStrobe_O[16] ;
 wire \Tile_X9Y9_FrameStrobe_O[17] ;
 wire \Tile_X9Y9_FrameStrobe_O[18] ;
 wire \Tile_X9Y9_FrameStrobe_O[19] ;
 wire \Tile_X9Y9_FrameStrobe_O[1] ;
 wire \Tile_X9Y9_FrameStrobe_O[2] ;
 wire \Tile_X9Y9_FrameStrobe_O[3] ;
 wire \Tile_X9Y9_FrameStrobe_O[4] ;
 wire \Tile_X9Y9_FrameStrobe_O[5] ;
 wire \Tile_X9Y9_FrameStrobe_O[6] ;
 wire \Tile_X9Y9_FrameStrobe_O[7] ;
 wire \Tile_X9Y9_FrameStrobe_O[8] ;
 wire \Tile_X9Y9_FrameStrobe_O[9] ;
 wire \Tile_X9Y9_N1BEG[0] ;
 wire \Tile_X9Y9_N1BEG[1] ;
 wire \Tile_X9Y9_N1BEG[2] ;
 wire \Tile_X9Y9_N1BEG[3] ;
 wire \Tile_X9Y9_N2BEG[0] ;
 wire \Tile_X9Y9_N2BEG[1] ;
 wire \Tile_X9Y9_N2BEG[2] ;
 wire \Tile_X9Y9_N2BEG[3] ;
 wire \Tile_X9Y9_N2BEG[4] ;
 wire \Tile_X9Y9_N2BEG[5] ;
 wire \Tile_X9Y9_N2BEG[6] ;
 wire \Tile_X9Y9_N2BEG[7] ;
 wire \Tile_X9Y9_N2BEGb[0] ;
 wire \Tile_X9Y9_N2BEGb[1] ;
 wire \Tile_X9Y9_N2BEGb[2] ;
 wire \Tile_X9Y9_N2BEGb[3] ;
 wire \Tile_X9Y9_N2BEGb[4] ;
 wire \Tile_X9Y9_N2BEGb[5] ;
 wire \Tile_X9Y9_N2BEGb[6] ;
 wire \Tile_X9Y9_N2BEGb[7] ;
 wire \Tile_X9Y9_N4BEG[0] ;
 wire \Tile_X9Y9_N4BEG[10] ;
 wire \Tile_X9Y9_N4BEG[11] ;
 wire \Tile_X9Y9_N4BEG[12] ;
 wire \Tile_X9Y9_N4BEG[13] ;
 wire \Tile_X9Y9_N4BEG[14] ;
 wire \Tile_X9Y9_N4BEG[15] ;
 wire \Tile_X9Y9_N4BEG[1] ;
 wire \Tile_X9Y9_N4BEG[2] ;
 wire \Tile_X9Y9_N4BEG[3] ;
 wire \Tile_X9Y9_N4BEG[4] ;
 wire \Tile_X9Y9_N4BEG[5] ;
 wire \Tile_X9Y9_N4BEG[6] ;
 wire \Tile_X9Y9_N4BEG[7] ;
 wire \Tile_X9Y9_N4BEG[8] ;
 wire \Tile_X9Y9_N4BEG[9] ;
 wire \Tile_X9Y9_NN4BEG[0] ;
 wire \Tile_X9Y9_NN4BEG[10] ;
 wire \Tile_X9Y9_NN4BEG[11] ;
 wire \Tile_X9Y9_NN4BEG[12] ;
 wire \Tile_X9Y9_NN4BEG[13] ;
 wire \Tile_X9Y9_NN4BEG[14] ;
 wire \Tile_X9Y9_NN4BEG[15] ;
 wire \Tile_X9Y9_NN4BEG[1] ;
 wire \Tile_X9Y9_NN4BEG[2] ;
 wire \Tile_X9Y9_NN4BEG[3] ;
 wire \Tile_X9Y9_NN4BEG[4] ;
 wire \Tile_X9Y9_NN4BEG[5] ;
 wire \Tile_X9Y9_NN4BEG[6] ;
 wire \Tile_X9Y9_NN4BEG[7] ;
 wire \Tile_X9Y9_NN4BEG[8] ;
 wire \Tile_X9Y9_NN4BEG[9] ;
 wire \Tile_X9Y9_S1BEG[0] ;
 wire \Tile_X9Y9_S1BEG[1] ;
 wire \Tile_X9Y9_S1BEG[2] ;
 wire \Tile_X9Y9_S1BEG[3] ;
 wire \Tile_X9Y9_S2BEG[0] ;
 wire \Tile_X9Y9_S2BEG[1] ;
 wire \Tile_X9Y9_S2BEG[2] ;
 wire \Tile_X9Y9_S2BEG[3] ;
 wire \Tile_X9Y9_S2BEG[4] ;
 wire \Tile_X9Y9_S2BEG[5] ;
 wire \Tile_X9Y9_S2BEG[6] ;
 wire \Tile_X9Y9_S2BEG[7] ;
 wire \Tile_X9Y9_S2BEGb[0] ;
 wire \Tile_X9Y9_S2BEGb[1] ;
 wire \Tile_X9Y9_S2BEGb[2] ;
 wire \Tile_X9Y9_S2BEGb[3] ;
 wire \Tile_X9Y9_S2BEGb[4] ;
 wire \Tile_X9Y9_S2BEGb[5] ;
 wire \Tile_X9Y9_S2BEGb[6] ;
 wire \Tile_X9Y9_S2BEGb[7] ;
 wire \Tile_X9Y9_S4BEG[0] ;
 wire \Tile_X9Y9_S4BEG[10] ;
 wire \Tile_X9Y9_S4BEG[11] ;
 wire \Tile_X9Y9_S4BEG[12] ;
 wire \Tile_X9Y9_S4BEG[13] ;
 wire \Tile_X9Y9_S4BEG[14] ;
 wire \Tile_X9Y9_S4BEG[15] ;
 wire \Tile_X9Y9_S4BEG[1] ;
 wire \Tile_X9Y9_S4BEG[2] ;
 wire \Tile_X9Y9_S4BEG[3] ;
 wire \Tile_X9Y9_S4BEG[4] ;
 wire \Tile_X9Y9_S4BEG[5] ;
 wire \Tile_X9Y9_S4BEG[6] ;
 wire \Tile_X9Y9_S4BEG[7] ;
 wire \Tile_X9Y9_S4BEG[8] ;
 wire \Tile_X9Y9_S4BEG[9] ;
 wire \Tile_X9Y9_SS4BEG[0] ;
 wire \Tile_X9Y9_SS4BEG[10] ;
 wire \Tile_X9Y9_SS4BEG[11] ;
 wire \Tile_X9Y9_SS4BEG[12] ;
 wire \Tile_X9Y9_SS4BEG[13] ;
 wire \Tile_X9Y9_SS4BEG[14] ;
 wire \Tile_X9Y9_SS4BEG[15] ;
 wire \Tile_X9Y9_SS4BEG[1] ;
 wire \Tile_X9Y9_SS4BEG[2] ;
 wire \Tile_X9Y9_SS4BEG[3] ;
 wire \Tile_X9Y9_SS4BEG[4] ;
 wire \Tile_X9Y9_SS4BEG[5] ;
 wire \Tile_X9Y9_SS4BEG[6] ;
 wire \Tile_X9Y9_SS4BEG[7] ;
 wire \Tile_X9Y9_SS4BEG[8] ;
 wire \Tile_X9Y9_SS4BEG[9] ;
 wire Tile_X9Y9_UserCLKo;
 wire \Tile_X9Y9_W1BEG[0] ;
 wire \Tile_X9Y9_W1BEG[1] ;
 wire \Tile_X9Y9_W1BEG[2] ;
 wire \Tile_X9Y9_W1BEG[3] ;
 wire \Tile_X9Y9_W2BEG[0] ;
 wire \Tile_X9Y9_W2BEG[1] ;
 wire \Tile_X9Y9_W2BEG[2] ;
 wire \Tile_X9Y9_W2BEG[3] ;
 wire \Tile_X9Y9_W2BEG[4] ;
 wire \Tile_X9Y9_W2BEG[5] ;
 wire \Tile_X9Y9_W2BEG[6] ;
 wire \Tile_X9Y9_W2BEG[7] ;
 wire \Tile_X9Y9_W2BEGb[0] ;
 wire \Tile_X9Y9_W2BEGb[1] ;
 wire \Tile_X9Y9_W2BEGb[2] ;
 wire \Tile_X9Y9_W2BEGb[3] ;
 wire \Tile_X9Y9_W2BEGb[4] ;
 wire \Tile_X9Y9_W2BEGb[5] ;
 wire \Tile_X9Y9_W2BEGb[6] ;
 wire \Tile_X9Y9_W2BEGb[7] ;
 wire \Tile_X9Y9_W6BEG[0] ;
 wire \Tile_X9Y9_W6BEG[10] ;
 wire \Tile_X9Y9_W6BEG[11] ;
 wire \Tile_X9Y9_W6BEG[1] ;
 wire \Tile_X9Y9_W6BEG[2] ;
 wire \Tile_X9Y9_W6BEG[3] ;
 wire \Tile_X9Y9_W6BEG[4] ;
 wire \Tile_X9Y9_W6BEG[5] ;
 wire \Tile_X9Y9_W6BEG[6] ;
 wire \Tile_X9Y9_W6BEG[7] ;
 wire \Tile_X9Y9_W6BEG[8] ;
 wire \Tile_X9Y9_W6BEG[9] ;
 wire \Tile_X9Y9_WW4BEG[0] ;
 wire \Tile_X9Y9_WW4BEG[10] ;
 wire \Tile_X9Y9_WW4BEG[11] ;
 wire \Tile_X9Y9_WW4BEG[12] ;
 wire \Tile_X9Y9_WW4BEG[13] ;
 wire \Tile_X9Y9_WW4BEG[14] ;
 wire \Tile_X9Y9_WW4BEG[15] ;
 wire \Tile_X9Y9_WW4BEG[1] ;
 wire \Tile_X9Y9_WW4BEG[2] ;
 wire \Tile_X9Y9_WW4BEG[3] ;
 wire \Tile_X9Y9_WW4BEG[4] ;
 wire \Tile_X9Y9_WW4BEG[5] ;
 wire \Tile_X9Y9_WW4BEG[6] ;
 wire \Tile_X9Y9_WW4BEG[7] ;
 wire \Tile_X9Y9_WW4BEG[8] ;
 wire \Tile_X9Y9_WW4BEG[9] ;

 W_IO Tile_X0Y10_W_IO (.A_I_top(Tile_X0Y10_A_I_top),
    .A_O_top(Tile_X0Y10_A_O_top),
    .A_T_top(Tile_X0Y10_A_T_top),
    .A_config_C_bit0(Tile_X0Y10_A_config_C_bit0),
    .A_config_C_bit1(Tile_X0Y10_A_config_C_bit1),
    .A_config_C_bit2(Tile_X0Y10_A_config_C_bit2),
    .A_config_C_bit3(Tile_X0Y10_A_config_C_bit3),
    .B_I_top(Tile_X0Y10_B_I_top),
    .B_O_top(Tile_X0Y10_B_O_top),
    .B_T_top(Tile_X0Y10_B_T_top),
    .B_config_C_bit0(Tile_X0Y10_B_config_C_bit0),
    .B_config_C_bit1(Tile_X0Y10_B_config_C_bit1),
    .B_config_C_bit2(Tile_X0Y10_B_config_C_bit2),
    .B_config_C_bit3(Tile_X0Y10_B_config_C_bit3),
    .UserCLK(Tile_X0Y11_UserCLKo),
    .UserCLKo(Tile_X0Y10_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X0Y10_E1BEG[3] ,
    \Tile_X0Y10_E1BEG[2] ,
    \Tile_X0Y10_E1BEG[1] ,
    \Tile_X0Y10_E1BEG[0] }),
    .E2BEG({\Tile_X0Y10_E2BEG[7] ,
    \Tile_X0Y10_E2BEG[6] ,
    \Tile_X0Y10_E2BEG[5] ,
    \Tile_X0Y10_E2BEG[4] ,
    \Tile_X0Y10_E2BEG[3] ,
    \Tile_X0Y10_E2BEG[2] ,
    \Tile_X0Y10_E2BEG[1] ,
    \Tile_X0Y10_E2BEG[0] }),
    .E2BEGb({\Tile_X0Y10_E2BEGb[7] ,
    \Tile_X0Y10_E2BEGb[6] ,
    \Tile_X0Y10_E2BEGb[5] ,
    \Tile_X0Y10_E2BEGb[4] ,
    \Tile_X0Y10_E2BEGb[3] ,
    \Tile_X0Y10_E2BEGb[2] ,
    \Tile_X0Y10_E2BEGb[1] ,
    \Tile_X0Y10_E2BEGb[0] }),
    .E6BEG({\Tile_X0Y10_E6BEG[11] ,
    \Tile_X0Y10_E6BEG[10] ,
    \Tile_X0Y10_E6BEG[9] ,
    \Tile_X0Y10_E6BEG[8] ,
    \Tile_X0Y10_E6BEG[7] ,
    \Tile_X0Y10_E6BEG[6] ,
    \Tile_X0Y10_E6BEG[5] ,
    \Tile_X0Y10_E6BEG[4] ,
    \Tile_X0Y10_E6BEG[3] ,
    \Tile_X0Y10_E6BEG[2] ,
    \Tile_X0Y10_E6BEG[1] ,
    \Tile_X0Y10_E6BEG[0] }),
    .EE4BEG({\Tile_X0Y10_EE4BEG[15] ,
    \Tile_X0Y10_EE4BEG[14] ,
    \Tile_X0Y10_EE4BEG[13] ,
    \Tile_X0Y10_EE4BEG[12] ,
    \Tile_X0Y10_EE4BEG[11] ,
    \Tile_X0Y10_EE4BEG[10] ,
    \Tile_X0Y10_EE4BEG[9] ,
    \Tile_X0Y10_EE4BEG[8] ,
    \Tile_X0Y10_EE4BEG[7] ,
    \Tile_X0Y10_EE4BEG[6] ,
    \Tile_X0Y10_EE4BEG[5] ,
    \Tile_X0Y10_EE4BEG[4] ,
    \Tile_X0Y10_EE4BEG[3] ,
    \Tile_X0Y10_EE4BEG[2] ,
    \Tile_X0Y10_EE4BEG[1] ,
    \Tile_X0Y10_EE4BEG[0] }),
    .FrameData({FrameData[351],
    FrameData[350],
    FrameData[349],
    FrameData[348],
    FrameData[347],
    FrameData[346],
    FrameData[345],
    FrameData[344],
    FrameData[343],
    FrameData[342],
    FrameData[341],
    FrameData[340],
    FrameData[339],
    FrameData[338],
    FrameData[337],
    FrameData[336],
    FrameData[335],
    FrameData[334],
    FrameData[333],
    FrameData[332],
    FrameData[331],
    FrameData[330],
    FrameData[329],
    FrameData[328],
    FrameData[327],
    FrameData[326],
    FrameData[325],
    FrameData[324],
    FrameData[323],
    FrameData[322],
    FrameData[321],
    FrameData[320]}),
    .FrameData_O({\Tile_X0Y10_FrameData_O[31] ,
    \Tile_X0Y10_FrameData_O[30] ,
    \Tile_X0Y10_FrameData_O[29] ,
    \Tile_X0Y10_FrameData_O[28] ,
    \Tile_X0Y10_FrameData_O[27] ,
    \Tile_X0Y10_FrameData_O[26] ,
    \Tile_X0Y10_FrameData_O[25] ,
    \Tile_X0Y10_FrameData_O[24] ,
    \Tile_X0Y10_FrameData_O[23] ,
    \Tile_X0Y10_FrameData_O[22] ,
    \Tile_X0Y10_FrameData_O[21] ,
    \Tile_X0Y10_FrameData_O[20] ,
    \Tile_X0Y10_FrameData_O[19] ,
    \Tile_X0Y10_FrameData_O[18] ,
    \Tile_X0Y10_FrameData_O[17] ,
    \Tile_X0Y10_FrameData_O[16] ,
    \Tile_X0Y10_FrameData_O[15] ,
    \Tile_X0Y10_FrameData_O[14] ,
    \Tile_X0Y10_FrameData_O[13] ,
    \Tile_X0Y10_FrameData_O[12] ,
    \Tile_X0Y10_FrameData_O[11] ,
    \Tile_X0Y10_FrameData_O[10] ,
    \Tile_X0Y10_FrameData_O[9] ,
    \Tile_X0Y10_FrameData_O[8] ,
    \Tile_X0Y10_FrameData_O[7] ,
    \Tile_X0Y10_FrameData_O[6] ,
    \Tile_X0Y10_FrameData_O[5] ,
    \Tile_X0Y10_FrameData_O[4] ,
    \Tile_X0Y10_FrameData_O[3] ,
    \Tile_X0Y10_FrameData_O[2] ,
    \Tile_X0Y10_FrameData_O[1] ,
    \Tile_X0Y10_FrameData_O[0] }),
    .FrameStrobe({\Tile_X0Y11_FrameStrobe_O[19] ,
    \Tile_X0Y11_FrameStrobe_O[18] ,
    \Tile_X0Y11_FrameStrobe_O[17] ,
    \Tile_X0Y11_FrameStrobe_O[16] ,
    \Tile_X0Y11_FrameStrobe_O[15] ,
    \Tile_X0Y11_FrameStrobe_O[14] ,
    \Tile_X0Y11_FrameStrobe_O[13] ,
    \Tile_X0Y11_FrameStrobe_O[12] ,
    \Tile_X0Y11_FrameStrobe_O[11] ,
    \Tile_X0Y11_FrameStrobe_O[10] ,
    \Tile_X0Y11_FrameStrobe_O[9] ,
    \Tile_X0Y11_FrameStrobe_O[8] ,
    \Tile_X0Y11_FrameStrobe_O[7] ,
    \Tile_X0Y11_FrameStrobe_O[6] ,
    \Tile_X0Y11_FrameStrobe_O[5] ,
    \Tile_X0Y11_FrameStrobe_O[4] ,
    \Tile_X0Y11_FrameStrobe_O[3] ,
    \Tile_X0Y11_FrameStrobe_O[2] ,
    \Tile_X0Y11_FrameStrobe_O[1] ,
    \Tile_X0Y11_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X0Y10_FrameStrobe_O[19] ,
    \Tile_X0Y10_FrameStrobe_O[18] ,
    \Tile_X0Y10_FrameStrobe_O[17] ,
    \Tile_X0Y10_FrameStrobe_O[16] ,
    \Tile_X0Y10_FrameStrobe_O[15] ,
    \Tile_X0Y10_FrameStrobe_O[14] ,
    \Tile_X0Y10_FrameStrobe_O[13] ,
    \Tile_X0Y10_FrameStrobe_O[12] ,
    \Tile_X0Y10_FrameStrobe_O[11] ,
    \Tile_X0Y10_FrameStrobe_O[10] ,
    \Tile_X0Y10_FrameStrobe_O[9] ,
    \Tile_X0Y10_FrameStrobe_O[8] ,
    \Tile_X0Y10_FrameStrobe_O[7] ,
    \Tile_X0Y10_FrameStrobe_O[6] ,
    \Tile_X0Y10_FrameStrobe_O[5] ,
    \Tile_X0Y10_FrameStrobe_O[4] ,
    \Tile_X0Y10_FrameStrobe_O[3] ,
    \Tile_X0Y10_FrameStrobe_O[2] ,
    \Tile_X0Y10_FrameStrobe_O[1] ,
    \Tile_X0Y10_FrameStrobe_O[0] }),
    .W1END({\Tile_X1Y10_W1BEG[3] ,
    \Tile_X1Y10_W1BEG[2] ,
    \Tile_X1Y10_W1BEG[1] ,
    \Tile_X1Y10_W1BEG[0] }),
    .W2END({\Tile_X1Y10_W2BEGb[7] ,
    \Tile_X1Y10_W2BEGb[6] ,
    \Tile_X1Y10_W2BEGb[5] ,
    \Tile_X1Y10_W2BEGb[4] ,
    \Tile_X1Y10_W2BEGb[3] ,
    \Tile_X1Y10_W2BEGb[2] ,
    \Tile_X1Y10_W2BEGb[1] ,
    \Tile_X1Y10_W2BEGb[0] }),
    .W2MID({\Tile_X1Y10_W2BEG[7] ,
    \Tile_X1Y10_W2BEG[6] ,
    \Tile_X1Y10_W2BEG[5] ,
    \Tile_X1Y10_W2BEG[4] ,
    \Tile_X1Y10_W2BEG[3] ,
    \Tile_X1Y10_W2BEG[2] ,
    \Tile_X1Y10_W2BEG[1] ,
    \Tile_X1Y10_W2BEG[0] }),
    .W6END({\Tile_X1Y10_W6BEG[11] ,
    \Tile_X1Y10_W6BEG[10] ,
    \Tile_X1Y10_W6BEG[9] ,
    \Tile_X1Y10_W6BEG[8] ,
    \Tile_X1Y10_W6BEG[7] ,
    \Tile_X1Y10_W6BEG[6] ,
    \Tile_X1Y10_W6BEG[5] ,
    \Tile_X1Y10_W6BEG[4] ,
    \Tile_X1Y10_W6BEG[3] ,
    \Tile_X1Y10_W6BEG[2] ,
    \Tile_X1Y10_W6BEG[1] ,
    \Tile_X1Y10_W6BEG[0] }),
    .WW4END({\Tile_X1Y10_WW4BEG[15] ,
    \Tile_X1Y10_WW4BEG[14] ,
    \Tile_X1Y10_WW4BEG[13] ,
    \Tile_X1Y10_WW4BEG[12] ,
    \Tile_X1Y10_WW4BEG[11] ,
    \Tile_X1Y10_WW4BEG[10] ,
    \Tile_X1Y10_WW4BEG[9] ,
    \Tile_X1Y10_WW4BEG[8] ,
    \Tile_X1Y10_WW4BEG[7] ,
    \Tile_X1Y10_WW4BEG[6] ,
    \Tile_X1Y10_WW4BEG[5] ,
    \Tile_X1Y10_WW4BEG[4] ,
    \Tile_X1Y10_WW4BEG[3] ,
    \Tile_X1Y10_WW4BEG[2] ,
    \Tile_X1Y10_WW4BEG[1] ,
    \Tile_X1Y10_WW4BEG[0] }));
 W_IO Tile_X0Y11_W_IO (.A_I_top(Tile_X0Y11_A_I_top),
    .A_O_top(Tile_X0Y11_A_O_top),
    .A_T_top(Tile_X0Y11_A_T_top),
    .A_config_C_bit0(Tile_X0Y11_A_config_C_bit0),
    .A_config_C_bit1(Tile_X0Y11_A_config_C_bit1),
    .A_config_C_bit2(Tile_X0Y11_A_config_C_bit2),
    .A_config_C_bit3(Tile_X0Y11_A_config_C_bit3),
    .B_I_top(Tile_X0Y11_B_I_top),
    .B_O_top(Tile_X0Y11_B_O_top),
    .B_T_top(Tile_X0Y11_B_T_top),
    .B_config_C_bit0(Tile_X0Y11_B_config_C_bit0),
    .B_config_C_bit1(Tile_X0Y11_B_config_C_bit1),
    .B_config_C_bit2(Tile_X0Y11_B_config_C_bit2),
    .B_config_C_bit3(Tile_X0Y11_B_config_C_bit3),
    .UserCLK(Tile_X0Y12_UserCLKo),
    .UserCLKo(Tile_X0Y11_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X0Y11_E1BEG[3] ,
    \Tile_X0Y11_E1BEG[2] ,
    \Tile_X0Y11_E1BEG[1] ,
    \Tile_X0Y11_E1BEG[0] }),
    .E2BEG({\Tile_X0Y11_E2BEG[7] ,
    \Tile_X0Y11_E2BEG[6] ,
    \Tile_X0Y11_E2BEG[5] ,
    \Tile_X0Y11_E2BEG[4] ,
    \Tile_X0Y11_E2BEG[3] ,
    \Tile_X0Y11_E2BEG[2] ,
    \Tile_X0Y11_E2BEG[1] ,
    \Tile_X0Y11_E2BEG[0] }),
    .E2BEGb({\Tile_X0Y11_E2BEGb[7] ,
    \Tile_X0Y11_E2BEGb[6] ,
    \Tile_X0Y11_E2BEGb[5] ,
    \Tile_X0Y11_E2BEGb[4] ,
    \Tile_X0Y11_E2BEGb[3] ,
    \Tile_X0Y11_E2BEGb[2] ,
    \Tile_X0Y11_E2BEGb[1] ,
    \Tile_X0Y11_E2BEGb[0] }),
    .E6BEG({\Tile_X0Y11_E6BEG[11] ,
    \Tile_X0Y11_E6BEG[10] ,
    \Tile_X0Y11_E6BEG[9] ,
    \Tile_X0Y11_E6BEG[8] ,
    \Tile_X0Y11_E6BEG[7] ,
    \Tile_X0Y11_E6BEG[6] ,
    \Tile_X0Y11_E6BEG[5] ,
    \Tile_X0Y11_E6BEG[4] ,
    \Tile_X0Y11_E6BEG[3] ,
    \Tile_X0Y11_E6BEG[2] ,
    \Tile_X0Y11_E6BEG[1] ,
    \Tile_X0Y11_E6BEG[0] }),
    .EE4BEG({\Tile_X0Y11_EE4BEG[15] ,
    \Tile_X0Y11_EE4BEG[14] ,
    \Tile_X0Y11_EE4BEG[13] ,
    \Tile_X0Y11_EE4BEG[12] ,
    \Tile_X0Y11_EE4BEG[11] ,
    \Tile_X0Y11_EE4BEG[10] ,
    \Tile_X0Y11_EE4BEG[9] ,
    \Tile_X0Y11_EE4BEG[8] ,
    \Tile_X0Y11_EE4BEG[7] ,
    \Tile_X0Y11_EE4BEG[6] ,
    \Tile_X0Y11_EE4BEG[5] ,
    \Tile_X0Y11_EE4BEG[4] ,
    \Tile_X0Y11_EE4BEG[3] ,
    \Tile_X0Y11_EE4BEG[2] ,
    \Tile_X0Y11_EE4BEG[1] ,
    \Tile_X0Y11_EE4BEG[0] }),
    .FrameData({FrameData[383],
    FrameData[382],
    FrameData[381],
    FrameData[380],
    FrameData[379],
    FrameData[378],
    FrameData[377],
    FrameData[376],
    FrameData[375],
    FrameData[374],
    FrameData[373],
    FrameData[372],
    FrameData[371],
    FrameData[370],
    FrameData[369],
    FrameData[368],
    FrameData[367],
    FrameData[366],
    FrameData[365],
    FrameData[364],
    FrameData[363],
    FrameData[362],
    FrameData[361],
    FrameData[360],
    FrameData[359],
    FrameData[358],
    FrameData[357],
    FrameData[356],
    FrameData[355],
    FrameData[354],
    FrameData[353],
    FrameData[352]}),
    .FrameData_O({\Tile_X0Y11_FrameData_O[31] ,
    \Tile_X0Y11_FrameData_O[30] ,
    \Tile_X0Y11_FrameData_O[29] ,
    \Tile_X0Y11_FrameData_O[28] ,
    \Tile_X0Y11_FrameData_O[27] ,
    \Tile_X0Y11_FrameData_O[26] ,
    \Tile_X0Y11_FrameData_O[25] ,
    \Tile_X0Y11_FrameData_O[24] ,
    \Tile_X0Y11_FrameData_O[23] ,
    \Tile_X0Y11_FrameData_O[22] ,
    \Tile_X0Y11_FrameData_O[21] ,
    \Tile_X0Y11_FrameData_O[20] ,
    \Tile_X0Y11_FrameData_O[19] ,
    \Tile_X0Y11_FrameData_O[18] ,
    \Tile_X0Y11_FrameData_O[17] ,
    \Tile_X0Y11_FrameData_O[16] ,
    \Tile_X0Y11_FrameData_O[15] ,
    \Tile_X0Y11_FrameData_O[14] ,
    \Tile_X0Y11_FrameData_O[13] ,
    \Tile_X0Y11_FrameData_O[12] ,
    \Tile_X0Y11_FrameData_O[11] ,
    \Tile_X0Y11_FrameData_O[10] ,
    \Tile_X0Y11_FrameData_O[9] ,
    \Tile_X0Y11_FrameData_O[8] ,
    \Tile_X0Y11_FrameData_O[7] ,
    \Tile_X0Y11_FrameData_O[6] ,
    \Tile_X0Y11_FrameData_O[5] ,
    \Tile_X0Y11_FrameData_O[4] ,
    \Tile_X0Y11_FrameData_O[3] ,
    \Tile_X0Y11_FrameData_O[2] ,
    \Tile_X0Y11_FrameData_O[1] ,
    \Tile_X0Y11_FrameData_O[0] }),
    .FrameStrobe({\Tile_X0Y12_FrameStrobe_O[19] ,
    \Tile_X0Y12_FrameStrobe_O[18] ,
    \Tile_X0Y12_FrameStrobe_O[17] ,
    \Tile_X0Y12_FrameStrobe_O[16] ,
    \Tile_X0Y12_FrameStrobe_O[15] ,
    \Tile_X0Y12_FrameStrobe_O[14] ,
    \Tile_X0Y12_FrameStrobe_O[13] ,
    \Tile_X0Y12_FrameStrobe_O[12] ,
    \Tile_X0Y12_FrameStrobe_O[11] ,
    \Tile_X0Y12_FrameStrobe_O[10] ,
    \Tile_X0Y12_FrameStrobe_O[9] ,
    \Tile_X0Y12_FrameStrobe_O[8] ,
    \Tile_X0Y12_FrameStrobe_O[7] ,
    \Tile_X0Y12_FrameStrobe_O[6] ,
    \Tile_X0Y12_FrameStrobe_O[5] ,
    \Tile_X0Y12_FrameStrobe_O[4] ,
    \Tile_X0Y12_FrameStrobe_O[3] ,
    \Tile_X0Y12_FrameStrobe_O[2] ,
    \Tile_X0Y12_FrameStrobe_O[1] ,
    \Tile_X0Y12_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X0Y11_FrameStrobe_O[19] ,
    \Tile_X0Y11_FrameStrobe_O[18] ,
    \Tile_X0Y11_FrameStrobe_O[17] ,
    \Tile_X0Y11_FrameStrobe_O[16] ,
    \Tile_X0Y11_FrameStrobe_O[15] ,
    \Tile_X0Y11_FrameStrobe_O[14] ,
    \Tile_X0Y11_FrameStrobe_O[13] ,
    \Tile_X0Y11_FrameStrobe_O[12] ,
    \Tile_X0Y11_FrameStrobe_O[11] ,
    \Tile_X0Y11_FrameStrobe_O[10] ,
    \Tile_X0Y11_FrameStrobe_O[9] ,
    \Tile_X0Y11_FrameStrobe_O[8] ,
    \Tile_X0Y11_FrameStrobe_O[7] ,
    \Tile_X0Y11_FrameStrobe_O[6] ,
    \Tile_X0Y11_FrameStrobe_O[5] ,
    \Tile_X0Y11_FrameStrobe_O[4] ,
    \Tile_X0Y11_FrameStrobe_O[3] ,
    \Tile_X0Y11_FrameStrobe_O[2] ,
    \Tile_X0Y11_FrameStrobe_O[1] ,
    \Tile_X0Y11_FrameStrobe_O[0] }),
    .W1END({\Tile_X1Y11_W1BEG[3] ,
    \Tile_X1Y11_W1BEG[2] ,
    \Tile_X1Y11_W1BEG[1] ,
    \Tile_X1Y11_W1BEG[0] }),
    .W2END({\Tile_X1Y11_W2BEGb[7] ,
    \Tile_X1Y11_W2BEGb[6] ,
    \Tile_X1Y11_W2BEGb[5] ,
    \Tile_X1Y11_W2BEGb[4] ,
    \Tile_X1Y11_W2BEGb[3] ,
    \Tile_X1Y11_W2BEGb[2] ,
    \Tile_X1Y11_W2BEGb[1] ,
    \Tile_X1Y11_W2BEGb[0] }),
    .W2MID({\Tile_X1Y11_W2BEG[7] ,
    \Tile_X1Y11_W2BEG[6] ,
    \Tile_X1Y11_W2BEG[5] ,
    \Tile_X1Y11_W2BEG[4] ,
    \Tile_X1Y11_W2BEG[3] ,
    \Tile_X1Y11_W2BEG[2] ,
    \Tile_X1Y11_W2BEG[1] ,
    \Tile_X1Y11_W2BEG[0] }),
    .W6END({\Tile_X1Y11_W6BEG[11] ,
    \Tile_X1Y11_W6BEG[10] ,
    \Tile_X1Y11_W6BEG[9] ,
    \Tile_X1Y11_W6BEG[8] ,
    \Tile_X1Y11_W6BEG[7] ,
    \Tile_X1Y11_W6BEG[6] ,
    \Tile_X1Y11_W6BEG[5] ,
    \Tile_X1Y11_W6BEG[4] ,
    \Tile_X1Y11_W6BEG[3] ,
    \Tile_X1Y11_W6BEG[2] ,
    \Tile_X1Y11_W6BEG[1] ,
    \Tile_X1Y11_W6BEG[0] }),
    .WW4END({\Tile_X1Y11_WW4BEG[15] ,
    \Tile_X1Y11_WW4BEG[14] ,
    \Tile_X1Y11_WW4BEG[13] ,
    \Tile_X1Y11_WW4BEG[12] ,
    \Tile_X1Y11_WW4BEG[11] ,
    \Tile_X1Y11_WW4BEG[10] ,
    \Tile_X1Y11_WW4BEG[9] ,
    \Tile_X1Y11_WW4BEG[8] ,
    \Tile_X1Y11_WW4BEG[7] ,
    \Tile_X1Y11_WW4BEG[6] ,
    \Tile_X1Y11_WW4BEG[5] ,
    \Tile_X1Y11_WW4BEG[4] ,
    \Tile_X1Y11_WW4BEG[3] ,
    \Tile_X1Y11_WW4BEG[2] ,
    \Tile_X1Y11_WW4BEG[1] ,
    \Tile_X1Y11_WW4BEG[0] }));
 W_IO Tile_X0Y12_W_IO (.A_I_top(Tile_X0Y12_A_I_top),
    .A_O_top(Tile_X0Y12_A_O_top),
    .A_T_top(Tile_X0Y12_A_T_top),
    .A_config_C_bit0(Tile_X0Y12_A_config_C_bit0),
    .A_config_C_bit1(Tile_X0Y12_A_config_C_bit1),
    .A_config_C_bit2(Tile_X0Y12_A_config_C_bit2),
    .A_config_C_bit3(Tile_X0Y12_A_config_C_bit3),
    .B_I_top(Tile_X0Y12_B_I_top),
    .B_O_top(Tile_X0Y12_B_O_top),
    .B_T_top(Tile_X0Y12_B_T_top),
    .B_config_C_bit0(Tile_X0Y12_B_config_C_bit0),
    .B_config_C_bit1(Tile_X0Y12_B_config_C_bit1),
    .B_config_C_bit2(Tile_X0Y12_B_config_C_bit2),
    .B_config_C_bit3(Tile_X0Y12_B_config_C_bit3),
    .UserCLK(Tile_X0Y13_UserCLKo),
    .UserCLKo(Tile_X0Y12_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X0Y12_E1BEG[3] ,
    \Tile_X0Y12_E1BEG[2] ,
    \Tile_X0Y12_E1BEG[1] ,
    \Tile_X0Y12_E1BEG[0] }),
    .E2BEG({\Tile_X0Y12_E2BEG[7] ,
    \Tile_X0Y12_E2BEG[6] ,
    \Tile_X0Y12_E2BEG[5] ,
    \Tile_X0Y12_E2BEG[4] ,
    \Tile_X0Y12_E2BEG[3] ,
    \Tile_X0Y12_E2BEG[2] ,
    \Tile_X0Y12_E2BEG[1] ,
    \Tile_X0Y12_E2BEG[0] }),
    .E2BEGb({\Tile_X0Y12_E2BEGb[7] ,
    \Tile_X0Y12_E2BEGb[6] ,
    \Tile_X0Y12_E2BEGb[5] ,
    \Tile_X0Y12_E2BEGb[4] ,
    \Tile_X0Y12_E2BEGb[3] ,
    \Tile_X0Y12_E2BEGb[2] ,
    \Tile_X0Y12_E2BEGb[1] ,
    \Tile_X0Y12_E2BEGb[0] }),
    .E6BEG({\Tile_X0Y12_E6BEG[11] ,
    \Tile_X0Y12_E6BEG[10] ,
    \Tile_X0Y12_E6BEG[9] ,
    \Tile_X0Y12_E6BEG[8] ,
    \Tile_X0Y12_E6BEG[7] ,
    \Tile_X0Y12_E6BEG[6] ,
    \Tile_X0Y12_E6BEG[5] ,
    \Tile_X0Y12_E6BEG[4] ,
    \Tile_X0Y12_E6BEG[3] ,
    \Tile_X0Y12_E6BEG[2] ,
    \Tile_X0Y12_E6BEG[1] ,
    \Tile_X0Y12_E6BEG[0] }),
    .EE4BEG({\Tile_X0Y12_EE4BEG[15] ,
    \Tile_X0Y12_EE4BEG[14] ,
    \Tile_X0Y12_EE4BEG[13] ,
    \Tile_X0Y12_EE4BEG[12] ,
    \Tile_X0Y12_EE4BEG[11] ,
    \Tile_X0Y12_EE4BEG[10] ,
    \Tile_X0Y12_EE4BEG[9] ,
    \Tile_X0Y12_EE4BEG[8] ,
    \Tile_X0Y12_EE4BEG[7] ,
    \Tile_X0Y12_EE4BEG[6] ,
    \Tile_X0Y12_EE4BEG[5] ,
    \Tile_X0Y12_EE4BEG[4] ,
    \Tile_X0Y12_EE4BEG[3] ,
    \Tile_X0Y12_EE4BEG[2] ,
    \Tile_X0Y12_EE4BEG[1] ,
    \Tile_X0Y12_EE4BEG[0] }),
    .FrameData({FrameData[415],
    FrameData[414],
    FrameData[413],
    FrameData[412],
    FrameData[411],
    FrameData[410],
    FrameData[409],
    FrameData[408],
    FrameData[407],
    FrameData[406],
    FrameData[405],
    FrameData[404],
    FrameData[403],
    FrameData[402],
    FrameData[401],
    FrameData[400],
    FrameData[399],
    FrameData[398],
    FrameData[397],
    FrameData[396],
    FrameData[395],
    FrameData[394],
    FrameData[393],
    FrameData[392],
    FrameData[391],
    FrameData[390],
    FrameData[389],
    FrameData[388],
    FrameData[387],
    FrameData[386],
    FrameData[385],
    FrameData[384]}),
    .FrameData_O({\Tile_X0Y12_FrameData_O[31] ,
    \Tile_X0Y12_FrameData_O[30] ,
    \Tile_X0Y12_FrameData_O[29] ,
    \Tile_X0Y12_FrameData_O[28] ,
    \Tile_X0Y12_FrameData_O[27] ,
    \Tile_X0Y12_FrameData_O[26] ,
    \Tile_X0Y12_FrameData_O[25] ,
    \Tile_X0Y12_FrameData_O[24] ,
    \Tile_X0Y12_FrameData_O[23] ,
    \Tile_X0Y12_FrameData_O[22] ,
    \Tile_X0Y12_FrameData_O[21] ,
    \Tile_X0Y12_FrameData_O[20] ,
    \Tile_X0Y12_FrameData_O[19] ,
    \Tile_X0Y12_FrameData_O[18] ,
    \Tile_X0Y12_FrameData_O[17] ,
    \Tile_X0Y12_FrameData_O[16] ,
    \Tile_X0Y12_FrameData_O[15] ,
    \Tile_X0Y12_FrameData_O[14] ,
    \Tile_X0Y12_FrameData_O[13] ,
    \Tile_X0Y12_FrameData_O[12] ,
    \Tile_X0Y12_FrameData_O[11] ,
    \Tile_X0Y12_FrameData_O[10] ,
    \Tile_X0Y12_FrameData_O[9] ,
    \Tile_X0Y12_FrameData_O[8] ,
    \Tile_X0Y12_FrameData_O[7] ,
    \Tile_X0Y12_FrameData_O[6] ,
    \Tile_X0Y12_FrameData_O[5] ,
    \Tile_X0Y12_FrameData_O[4] ,
    \Tile_X0Y12_FrameData_O[3] ,
    \Tile_X0Y12_FrameData_O[2] ,
    \Tile_X0Y12_FrameData_O[1] ,
    \Tile_X0Y12_FrameData_O[0] }),
    .FrameStrobe({\Tile_X0Y13_FrameStrobe_O[19] ,
    \Tile_X0Y13_FrameStrobe_O[18] ,
    \Tile_X0Y13_FrameStrobe_O[17] ,
    \Tile_X0Y13_FrameStrobe_O[16] ,
    \Tile_X0Y13_FrameStrobe_O[15] ,
    \Tile_X0Y13_FrameStrobe_O[14] ,
    \Tile_X0Y13_FrameStrobe_O[13] ,
    \Tile_X0Y13_FrameStrobe_O[12] ,
    \Tile_X0Y13_FrameStrobe_O[11] ,
    \Tile_X0Y13_FrameStrobe_O[10] ,
    \Tile_X0Y13_FrameStrobe_O[9] ,
    \Tile_X0Y13_FrameStrobe_O[8] ,
    \Tile_X0Y13_FrameStrobe_O[7] ,
    \Tile_X0Y13_FrameStrobe_O[6] ,
    \Tile_X0Y13_FrameStrobe_O[5] ,
    \Tile_X0Y13_FrameStrobe_O[4] ,
    \Tile_X0Y13_FrameStrobe_O[3] ,
    \Tile_X0Y13_FrameStrobe_O[2] ,
    \Tile_X0Y13_FrameStrobe_O[1] ,
    \Tile_X0Y13_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X0Y12_FrameStrobe_O[19] ,
    \Tile_X0Y12_FrameStrobe_O[18] ,
    \Tile_X0Y12_FrameStrobe_O[17] ,
    \Tile_X0Y12_FrameStrobe_O[16] ,
    \Tile_X0Y12_FrameStrobe_O[15] ,
    \Tile_X0Y12_FrameStrobe_O[14] ,
    \Tile_X0Y12_FrameStrobe_O[13] ,
    \Tile_X0Y12_FrameStrobe_O[12] ,
    \Tile_X0Y12_FrameStrobe_O[11] ,
    \Tile_X0Y12_FrameStrobe_O[10] ,
    \Tile_X0Y12_FrameStrobe_O[9] ,
    \Tile_X0Y12_FrameStrobe_O[8] ,
    \Tile_X0Y12_FrameStrobe_O[7] ,
    \Tile_X0Y12_FrameStrobe_O[6] ,
    \Tile_X0Y12_FrameStrobe_O[5] ,
    \Tile_X0Y12_FrameStrobe_O[4] ,
    \Tile_X0Y12_FrameStrobe_O[3] ,
    \Tile_X0Y12_FrameStrobe_O[2] ,
    \Tile_X0Y12_FrameStrobe_O[1] ,
    \Tile_X0Y12_FrameStrobe_O[0] }),
    .W1END({\Tile_X1Y12_W1BEG[3] ,
    \Tile_X1Y12_W1BEG[2] ,
    \Tile_X1Y12_W1BEG[1] ,
    \Tile_X1Y12_W1BEG[0] }),
    .W2END({\Tile_X1Y12_W2BEGb[7] ,
    \Tile_X1Y12_W2BEGb[6] ,
    \Tile_X1Y12_W2BEGb[5] ,
    \Tile_X1Y12_W2BEGb[4] ,
    \Tile_X1Y12_W2BEGb[3] ,
    \Tile_X1Y12_W2BEGb[2] ,
    \Tile_X1Y12_W2BEGb[1] ,
    \Tile_X1Y12_W2BEGb[0] }),
    .W2MID({\Tile_X1Y12_W2BEG[7] ,
    \Tile_X1Y12_W2BEG[6] ,
    \Tile_X1Y12_W2BEG[5] ,
    \Tile_X1Y12_W2BEG[4] ,
    \Tile_X1Y12_W2BEG[3] ,
    \Tile_X1Y12_W2BEG[2] ,
    \Tile_X1Y12_W2BEG[1] ,
    \Tile_X1Y12_W2BEG[0] }),
    .W6END({\Tile_X1Y12_W6BEG[11] ,
    \Tile_X1Y12_W6BEG[10] ,
    \Tile_X1Y12_W6BEG[9] ,
    \Tile_X1Y12_W6BEG[8] ,
    \Tile_X1Y12_W6BEG[7] ,
    \Tile_X1Y12_W6BEG[6] ,
    \Tile_X1Y12_W6BEG[5] ,
    \Tile_X1Y12_W6BEG[4] ,
    \Tile_X1Y12_W6BEG[3] ,
    \Tile_X1Y12_W6BEG[2] ,
    \Tile_X1Y12_W6BEG[1] ,
    \Tile_X1Y12_W6BEG[0] }),
    .WW4END({\Tile_X1Y12_WW4BEG[15] ,
    \Tile_X1Y12_WW4BEG[14] ,
    \Tile_X1Y12_WW4BEG[13] ,
    \Tile_X1Y12_WW4BEG[12] ,
    \Tile_X1Y12_WW4BEG[11] ,
    \Tile_X1Y12_WW4BEG[10] ,
    \Tile_X1Y12_WW4BEG[9] ,
    \Tile_X1Y12_WW4BEG[8] ,
    \Tile_X1Y12_WW4BEG[7] ,
    \Tile_X1Y12_WW4BEG[6] ,
    \Tile_X1Y12_WW4BEG[5] ,
    \Tile_X1Y12_WW4BEG[4] ,
    \Tile_X1Y12_WW4BEG[3] ,
    \Tile_X1Y12_WW4BEG[2] ,
    \Tile_X1Y12_WW4BEG[1] ,
    \Tile_X1Y12_WW4BEG[0] }));
 W_IO Tile_X0Y13_W_IO (.A_I_top(Tile_X0Y13_A_I_top),
    .A_O_top(Tile_X0Y13_A_O_top),
    .A_T_top(Tile_X0Y13_A_T_top),
    .A_config_C_bit0(Tile_X0Y13_A_config_C_bit0),
    .A_config_C_bit1(Tile_X0Y13_A_config_C_bit1),
    .A_config_C_bit2(Tile_X0Y13_A_config_C_bit2),
    .A_config_C_bit3(Tile_X0Y13_A_config_C_bit3),
    .B_I_top(Tile_X0Y13_B_I_top),
    .B_O_top(Tile_X0Y13_B_O_top),
    .B_T_top(Tile_X0Y13_B_T_top),
    .B_config_C_bit0(Tile_X0Y13_B_config_C_bit0),
    .B_config_C_bit1(Tile_X0Y13_B_config_C_bit1),
    .B_config_C_bit2(Tile_X0Y13_B_config_C_bit2),
    .B_config_C_bit3(Tile_X0Y13_B_config_C_bit3),
    .UserCLK(Tile_X0Y14_UserCLKo),
    .UserCLKo(Tile_X0Y13_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X0Y13_E1BEG[3] ,
    \Tile_X0Y13_E1BEG[2] ,
    \Tile_X0Y13_E1BEG[1] ,
    \Tile_X0Y13_E1BEG[0] }),
    .E2BEG({\Tile_X0Y13_E2BEG[7] ,
    \Tile_X0Y13_E2BEG[6] ,
    \Tile_X0Y13_E2BEG[5] ,
    \Tile_X0Y13_E2BEG[4] ,
    \Tile_X0Y13_E2BEG[3] ,
    \Tile_X0Y13_E2BEG[2] ,
    \Tile_X0Y13_E2BEG[1] ,
    \Tile_X0Y13_E2BEG[0] }),
    .E2BEGb({\Tile_X0Y13_E2BEGb[7] ,
    \Tile_X0Y13_E2BEGb[6] ,
    \Tile_X0Y13_E2BEGb[5] ,
    \Tile_X0Y13_E2BEGb[4] ,
    \Tile_X0Y13_E2BEGb[3] ,
    \Tile_X0Y13_E2BEGb[2] ,
    \Tile_X0Y13_E2BEGb[1] ,
    \Tile_X0Y13_E2BEGb[0] }),
    .E6BEG({\Tile_X0Y13_E6BEG[11] ,
    \Tile_X0Y13_E6BEG[10] ,
    \Tile_X0Y13_E6BEG[9] ,
    \Tile_X0Y13_E6BEG[8] ,
    \Tile_X0Y13_E6BEG[7] ,
    \Tile_X0Y13_E6BEG[6] ,
    \Tile_X0Y13_E6BEG[5] ,
    \Tile_X0Y13_E6BEG[4] ,
    \Tile_X0Y13_E6BEG[3] ,
    \Tile_X0Y13_E6BEG[2] ,
    \Tile_X0Y13_E6BEG[1] ,
    \Tile_X0Y13_E6BEG[0] }),
    .EE4BEG({\Tile_X0Y13_EE4BEG[15] ,
    \Tile_X0Y13_EE4BEG[14] ,
    \Tile_X0Y13_EE4BEG[13] ,
    \Tile_X0Y13_EE4BEG[12] ,
    \Tile_X0Y13_EE4BEG[11] ,
    \Tile_X0Y13_EE4BEG[10] ,
    \Tile_X0Y13_EE4BEG[9] ,
    \Tile_X0Y13_EE4BEG[8] ,
    \Tile_X0Y13_EE4BEG[7] ,
    \Tile_X0Y13_EE4BEG[6] ,
    \Tile_X0Y13_EE4BEG[5] ,
    \Tile_X0Y13_EE4BEG[4] ,
    \Tile_X0Y13_EE4BEG[3] ,
    \Tile_X0Y13_EE4BEG[2] ,
    \Tile_X0Y13_EE4BEG[1] ,
    \Tile_X0Y13_EE4BEG[0] }),
    .FrameData({FrameData[447],
    FrameData[446],
    FrameData[445],
    FrameData[444],
    FrameData[443],
    FrameData[442],
    FrameData[441],
    FrameData[440],
    FrameData[439],
    FrameData[438],
    FrameData[437],
    FrameData[436],
    FrameData[435],
    FrameData[434],
    FrameData[433],
    FrameData[432],
    FrameData[431],
    FrameData[430],
    FrameData[429],
    FrameData[428],
    FrameData[427],
    FrameData[426],
    FrameData[425],
    FrameData[424],
    FrameData[423],
    FrameData[422],
    FrameData[421],
    FrameData[420],
    FrameData[419],
    FrameData[418],
    FrameData[417],
    FrameData[416]}),
    .FrameData_O({\Tile_X0Y13_FrameData_O[31] ,
    \Tile_X0Y13_FrameData_O[30] ,
    \Tile_X0Y13_FrameData_O[29] ,
    \Tile_X0Y13_FrameData_O[28] ,
    \Tile_X0Y13_FrameData_O[27] ,
    \Tile_X0Y13_FrameData_O[26] ,
    \Tile_X0Y13_FrameData_O[25] ,
    \Tile_X0Y13_FrameData_O[24] ,
    \Tile_X0Y13_FrameData_O[23] ,
    \Tile_X0Y13_FrameData_O[22] ,
    \Tile_X0Y13_FrameData_O[21] ,
    \Tile_X0Y13_FrameData_O[20] ,
    \Tile_X0Y13_FrameData_O[19] ,
    \Tile_X0Y13_FrameData_O[18] ,
    \Tile_X0Y13_FrameData_O[17] ,
    \Tile_X0Y13_FrameData_O[16] ,
    \Tile_X0Y13_FrameData_O[15] ,
    \Tile_X0Y13_FrameData_O[14] ,
    \Tile_X0Y13_FrameData_O[13] ,
    \Tile_X0Y13_FrameData_O[12] ,
    \Tile_X0Y13_FrameData_O[11] ,
    \Tile_X0Y13_FrameData_O[10] ,
    \Tile_X0Y13_FrameData_O[9] ,
    \Tile_X0Y13_FrameData_O[8] ,
    \Tile_X0Y13_FrameData_O[7] ,
    \Tile_X0Y13_FrameData_O[6] ,
    \Tile_X0Y13_FrameData_O[5] ,
    \Tile_X0Y13_FrameData_O[4] ,
    \Tile_X0Y13_FrameData_O[3] ,
    \Tile_X0Y13_FrameData_O[2] ,
    \Tile_X0Y13_FrameData_O[1] ,
    \Tile_X0Y13_FrameData_O[0] }),
    .FrameStrobe({\Tile_X0Y14_FrameStrobe_O[19] ,
    \Tile_X0Y14_FrameStrobe_O[18] ,
    \Tile_X0Y14_FrameStrobe_O[17] ,
    \Tile_X0Y14_FrameStrobe_O[16] ,
    \Tile_X0Y14_FrameStrobe_O[15] ,
    \Tile_X0Y14_FrameStrobe_O[14] ,
    \Tile_X0Y14_FrameStrobe_O[13] ,
    \Tile_X0Y14_FrameStrobe_O[12] ,
    \Tile_X0Y14_FrameStrobe_O[11] ,
    \Tile_X0Y14_FrameStrobe_O[10] ,
    \Tile_X0Y14_FrameStrobe_O[9] ,
    \Tile_X0Y14_FrameStrobe_O[8] ,
    \Tile_X0Y14_FrameStrobe_O[7] ,
    \Tile_X0Y14_FrameStrobe_O[6] ,
    \Tile_X0Y14_FrameStrobe_O[5] ,
    \Tile_X0Y14_FrameStrobe_O[4] ,
    \Tile_X0Y14_FrameStrobe_O[3] ,
    \Tile_X0Y14_FrameStrobe_O[2] ,
    \Tile_X0Y14_FrameStrobe_O[1] ,
    \Tile_X0Y14_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X0Y13_FrameStrobe_O[19] ,
    \Tile_X0Y13_FrameStrobe_O[18] ,
    \Tile_X0Y13_FrameStrobe_O[17] ,
    \Tile_X0Y13_FrameStrobe_O[16] ,
    \Tile_X0Y13_FrameStrobe_O[15] ,
    \Tile_X0Y13_FrameStrobe_O[14] ,
    \Tile_X0Y13_FrameStrobe_O[13] ,
    \Tile_X0Y13_FrameStrobe_O[12] ,
    \Tile_X0Y13_FrameStrobe_O[11] ,
    \Tile_X0Y13_FrameStrobe_O[10] ,
    \Tile_X0Y13_FrameStrobe_O[9] ,
    \Tile_X0Y13_FrameStrobe_O[8] ,
    \Tile_X0Y13_FrameStrobe_O[7] ,
    \Tile_X0Y13_FrameStrobe_O[6] ,
    \Tile_X0Y13_FrameStrobe_O[5] ,
    \Tile_X0Y13_FrameStrobe_O[4] ,
    \Tile_X0Y13_FrameStrobe_O[3] ,
    \Tile_X0Y13_FrameStrobe_O[2] ,
    \Tile_X0Y13_FrameStrobe_O[1] ,
    \Tile_X0Y13_FrameStrobe_O[0] }),
    .W1END({\Tile_X1Y13_W1BEG[3] ,
    \Tile_X1Y13_W1BEG[2] ,
    \Tile_X1Y13_W1BEG[1] ,
    \Tile_X1Y13_W1BEG[0] }),
    .W2END({\Tile_X1Y13_W2BEGb[7] ,
    \Tile_X1Y13_W2BEGb[6] ,
    \Tile_X1Y13_W2BEGb[5] ,
    \Tile_X1Y13_W2BEGb[4] ,
    \Tile_X1Y13_W2BEGb[3] ,
    \Tile_X1Y13_W2BEGb[2] ,
    \Tile_X1Y13_W2BEGb[1] ,
    \Tile_X1Y13_W2BEGb[0] }),
    .W2MID({\Tile_X1Y13_W2BEG[7] ,
    \Tile_X1Y13_W2BEG[6] ,
    \Tile_X1Y13_W2BEG[5] ,
    \Tile_X1Y13_W2BEG[4] ,
    \Tile_X1Y13_W2BEG[3] ,
    \Tile_X1Y13_W2BEG[2] ,
    \Tile_X1Y13_W2BEG[1] ,
    \Tile_X1Y13_W2BEG[0] }),
    .W6END({\Tile_X1Y13_W6BEG[11] ,
    \Tile_X1Y13_W6BEG[10] ,
    \Tile_X1Y13_W6BEG[9] ,
    \Tile_X1Y13_W6BEG[8] ,
    \Tile_X1Y13_W6BEG[7] ,
    \Tile_X1Y13_W6BEG[6] ,
    \Tile_X1Y13_W6BEG[5] ,
    \Tile_X1Y13_W6BEG[4] ,
    \Tile_X1Y13_W6BEG[3] ,
    \Tile_X1Y13_W6BEG[2] ,
    \Tile_X1Y13_W6BEG[1] ,
    \Tile_X1Y13_W6BEG[0] }),
    .WW4END({\Tile_X1Y13_WW4BEG[15] ,
    \Tile_X1Y13_WW4BEG[14] ,
    \Tile_X1Y13_WW4BEG[13] ,
    \Tile_X1Y13_WW4BEG[12] ,
    \Tile_X1Y13_WW4BEG[11] ,
    \Tile_X1Y13_WW4BEG[10] ,
    \Tile_X1Y13_WW4BEG[9] ,
    \Tile_X1Y13_WW4BEG[8] ,
    \Tile_X1Y13_WW4BEG[7] ,
    \Tile_X1Y13_WW4BEG[6] ,
    \Tile_X1Y13_WW4BEG[5] ,
    \Tile_X1Y13_WW4BEG[4] ,
    \Tile_X1Y13_WW4BEG[3] ,
    \Tile_X1Y13_WW4BEG[2] ,
    \Tile_X1Y13_WW4BEG[1] ,
    \Tile_X1Y13_WW4BEG[0] }));
 W_IO Tile_X0Y14_W_IO (.A_I_top(Tile_X0Y14_A_I_top),
    .A_O_top(Tile_X0Y14_A_O_top),
    .A_T_top(Tile_X0Y14_A_T_top),
    .A_config_C_bit0(Tile_X0Y14_A_config_C_bit0),
    .A_config_C_bit1(Tile_X0Y14_A_config_C_bit1),
    .A_config_C_bit2(Tile_X0Y14_A_config_C_bit2),
    .A_config_C_bit3(Tile_X0Y14_A_config_C_bit3),
    .B_I_top(Tile_X0Y14_B_I_top),
    .B_O_top(Tile_X0Y14_B_O_top),
    .B_T_top(Tile_X0Y14_B_T_top),
    .B_config_C_bit0(Tile_X0Y14_B_config_C_bit0),
    .B_config_C_bit1(Tile_X0Y14_B_config_C_bit1),
    .B_config_C_bit2(Tile_X0Y14_B_config_C_bit2),
    .B_config_C_bit3(Tile_X0Y14_B_config_C_bit3),
    .UserCLK(UserCLK),
    .UserCLKo(Tile_X0Y14_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X0Y14_E1BEG[3] ,
    \Tile_X0Y14_E1BEG[2] ,
    \Tile_X0Y14_E1BEG[1] ,
    \Tile_X0Y14_E1BEG[0] }),
    .E2BEG({\Tile_X0Y14_E2BEG[7] ,
    \Tile_X0Y14_E2BEG[6] ,
    \Tile_X0Y14_E2BEG[5] ,
    \Tile_X0Y14_E2BEG[4] ,
    \Tile_X0Y14_E2BEG[3] ,
    \Tile_X0Y14_E2BEG[2] ,
    \Tile_X0Y14_E2BEG[1] ,
    \Tile_X0Y14_E2BEG[0] }),
    .E2BEGb({\Tile_X0Y14_E2BEGb[7] ,
    \Tile_X0Y14_E2BEGb[6] ,
    \Tile_X0Y14_E2BEGb[5] ,
    \Tile_X0Y14_E2BEGb[4] ,
    \Tile_X0Y14_E2BEGb[3] ,
    \Tile_X0Y14_E2BEGb[2] ,
    \Tile_X0Y14_E2BEGb[1] ,
    \Tile_X0Y14_E2BEGb[0] }),
    .E6BEG({\Tile_X0Y14_E6BEG[11] ,
    \Tile_X0Y14_E6BEG[10] ,
    \Tile_X0Y14_E6BEG[9] ,
    \Tile_X0Y14_E6BEG[8] ,
    \Tile_X0Y14_E6BEG[7] ,
    \Tile_X0Y14_E6BEG[6] ,
    \Tile_X0Y14_E6BEG[5] ,
    \Tile_X0Y14_E6BEG[4] ,
    \Tile_X0Y14_E6BEG[3] ,
    \Tile_X0Y14_E6BEG[2] ,
    \Tile_X0Y14_E6BEG[1] ,
    \Tile_X0Y14_E6BEG[0] }),
    .EE4BEG({\Tile_X0Y14_EE4BEG[15] ,
    \Tile_X0Y14_EE4BEG[14] ,
    \Tile_X0Y14_EE4BEG[13] ,
    \Tile_X0Y14_EE4BEG[12] ,
    \Tile_X0Y14_EE4BEG[11] ,
    \Tile_X0Y14_EE4BEG[10] ,
    \Tile_X0Y14_EE4BEG[9] ,
    \Tile_X0Y14_EE4BEG[8] ,
    \Tile_X0Y14_EE4BEG[7] ,
    \Tile_X0Y14_EE4BEG[6] ,
    \Tile_X0Y14_EE4BEG[5] ,
    \Tile_X0Y14_EE4BEG[4] ,
    \Tile_X0Y14_EE4BEG[3] ,
    \Tile_X0Y14_EE4BEG[2] ,
    \Tile_X0Y14_EE4BEG[1] ,
    \Tile_X0Y14_EE4BEG[0] }),
    .FrameData({FrameData[479],
    FrameData[478],
    FrameData[477],
    FrameData[476],
    FrameData[475],
    FrameData[474],
    FrameData[473],
    FrameData[472],
    FrameData[471],
    FrameData[470],
    FrameData[469],
    FrameData[468],
    FrameData[467],
    FrameData[466],
    FrameData[465],
    FrameData[464],
    FrameData[463],
    FrameData[462],
    FrameData[461],
    FrameData[460],
    FrameData[459],
    FrameData[458],
    FrameData[457],
    FrameData[456],
    FrameData[455],
    FrameData[454],
    FrameData[453],
    FrameData[452],
    FrameData[451],
    FrameData[450],
    FrameData[449],
    FrameData[448]}),
    .FrameData_O({\Tile_X0Y14_FrameData_O[31] ,
    \Tile_X0Y14_FrameData_O[30] ,
    \Tile_X0Y14_FrameData_O[29] ,
    \Tile_X0Y14_FrameData_O[28] ,
    \Tile_X0Y14_FrameData_O[27] ,
    \Tile_X0Y14_FrameData_O[26] ,
    \Tile_X0Y14_FrameData_O[25] ,
    \Tile_X0Y14_FrameData_O[24] ,
    \Tile_X0Y14_FrameData_O[23] ,
    \Tile_X0Y14_FrameData_O[22] ,
    \Tile_X0Y14_FrameData_O[21] ,
    \Tile_X0Y14_FrameData_O[20] ,
    \Tile_X0Y14_FrameData_O[19] ,
    \Tile_X0Y14_FrameData_O[18] ,
    \Tile_X0Y14_FrameData_O[17] ,
    \Tile_X0Y14_FrameData_O[16] ,
    \Tile_X0Y14_FrameData_O[15] ,
    \Tile_X0Y14_FrameData_O[14] ,
    \Tile_X0Y14_FrameData_O[13] ,
    \Tile_X0Y14_FrameData_O[12] ,
    \Tile_X0Y14_FrameData_O[11] ,
    \Tile_X0Y14_FrameData_O[10] ,
    \Tile_X0Y14_FrameData_O[9] ,
    \Tile_X0Y14_FrameData_O[8] ,
    \Tile_X0Y14_FrameData_O[7] ,
    \Tile_X0Y14_FrameData_O[6] ,
    \Tile_X0Y14_FrameData_O[5] ,
    \Tile_X0Y14_FrameData_O[4] ,
    \Tile_X0Y14_FrameData_O[3] ,
    \Tile_X0Y14_FrameData_O[2] ,
    \Tile_X0Y14_FrameData_O[1] ,
    \Tile_X0Y14_FrameData_O[0] }),
    .FrameStrobe({FrameStrobe[19],
    FrameStrobe[18],
    FrameStrobe[17],
    FrameStrobe[16],
    FrameStrobe[15],
    FrameStrobe[14],
    FrameStrobe[13],
    FrameStrobe[12],
    FrameStrobe[11],
    FrameStrobe[10],
    FrameStrobe[9],
    FrameStrobe[8],
    FrameStrobe[7],
    FrameStrobe[6],
    FrameStrobe[5],
    FrameStrobe[4],
    FrameStrobe[3],
    FrameStrobe[2],
    FrameStrobe[1],
    FrameStrobe[0]}),
    .FrameStrobe_O({\Tile_X0Y14_FrameStrobe_O[19] ,
    \Tile_X0Y14_FrameStrobe_O[18] ,
    \Tile_X0Y14_FrameStrobe_O[17] ,
    \Tile_X0Y14_FrameStrobe_O[16] ,
    \Tile_X0Y14_FrameStrobe_O[15] ,
    \Tile_X0Y14_FrameStrobe_O[14] ,
    \Tile_X0Y14_FrameStrobe_O[13] ,
    \Tile_X0Y14_FrameStrobe_O[12] ,
    \Tile_X0Y14_FrameStrobe_O[11] ,
    \Tile_X0Y14_FrameStrobe_O[10] ,
    \Tile_X0Y14_FrameStrobe_O[9] ,
    \Tile_X0Y14_FrameStrobe_O[8] ,
    \Tile_X0Y14_FrameStrobe_O[7] ,
    \Tile_X0Y14_FrameStrobe_O[6] ,
    \Tile_X0Y14_FrameStrobe_O[5] ,
    \Tile_X0Y14_FrameStrobe_O[4] ,
    \Tile_X0Y14_FrameStrobe_O[3] ,
    \Tile_X0Y14_FrameStrobe_O[2] ,
    \Tile_X0Y14_FrameStrobe_O[1] ,
    \Tile_X0Y14_FrameStrobe_O[0] }),
    .W1END({\Tile_X1Y14_W1BEG[3] ,
    \Tile_X1Y14_W1BEG[2] ,
    \Tile_X1Y14_W1BEG[1] ,
    \Tile_X1Y14_W1BEG[0] }),
    .W2END({\Tile_X1Y14_W2BEGb[7] ,
    \Tile_X1Y14_W2BEGb[6] ,
    \Tile_X1Y14_W2BEGb[5] ,
    \Tile_X1Y14_W2BEGb[4] ,
    \Tile_X1Y14_W2BEGb[3] ,
    \Tile_X1Y14_W2BEGb[2] ,
    \Tile_X1Y14_W2BEGb[1] ,
    \Tile_X1Y14_W2BEGb[0] }),
    .W2MID({\Tile_X1Y14_W2BEG[7] ,
    \Tile_X1Y14_W2BEG[6] ,
    \Tile_X1Y14_W2BEG[5] ,
    \Tile_X1Y14_W2BEG[4] ,
    \Tile_X1Y14_W2BEG[3] ,
    \Tile_X1Y14_W2BEG[2] ,
    \Tile_X1Y14_W2BEG[1] ,
    \Tile_X1Y14_W2BEG[0] }),
    .W6END({\Tile_X1Y14_W6BEG[11] ,
    \Tile_X1Y14_W6BEG[10] ,
    \Tile_X1Y14_W6BEG[9] ,
    \Tile_X1Y14_W6BEG[8] ,
    \Tile_X1Y14_W6BEG[7] ,
    \Tile_X1Y14_W6BEG[6] ,
    \Tile_X1Y14_W6BEG[5] ,
    \Tile_X1Y14_W6BEG[4] ,
    \Tile_X1Y14_W6BEG[3] ,
    \Tile_X1Y14_W6BEG[2] ,
    \Tile_X1Y14_W6BEG[1] ,
    \Tile_X1Y14_W6BEG[0] }),
    .WW4END({\Tile_X1Y14_WW4BEG[15] ,
    \Tile_X1Y14_WW4BEG[14] ,
    \Tile_X1Y14_WW4BEG[13] ,
    \Tile_X1Y14_WW4BEG[12] ,
    \Tile_X1Y14_WW4BEG[11] ,
    \Tile_X1Y14_WW4BEG[10] ,
    \Tile_X1Y14_WW4BEG[9] ,
    \Tile_X1Y14_WW4BEG[8] ,
    \Tile_X1Y14_WW4BEG[7] ,
    \Tile_X1Y14_WW4BEG[6] ,
    \Tile_X1Y14_WW4BEG[5] ,
    \Tile_X1Y14_WW4BEG[4] ,
    \Tile_X1Y14_WW4BEG[3] ,
    \Tile_X1Y14_WW4BEG[2] ,
    \Tile_X1Y14_WW4BEG[1] ,
    \Tile_X1Y14_WW4BEG[0] }));
 W_IO Tile_X0Y1_W_IO (.A_I_top(Tile_X0Y1_A_I_top),
    .A_O_top(Tile_X0Y1_A_O_top),
    .A_T_top(Tile_X0Y1_A_T_top),
    .A_config_C_bit0(Tile_X0Y1_A_config_C_bit0),
    .A_config_C_bit1(Tile_X0Y1_A_config_C_bit1),
    .A_config_C_bit2(Tile_X0Y1_A_config_C_bit2),
    .A_config_C_bit3(Tile_X0Y1_A_config_C_bit3),
    .B_I_top(Tile_X0Y1_B_I_top),
    .B_O_top(Tile_X0Y1_B_O_top),
    .B_T_top(Tile_X0Y1_B_T_top),
    .B_config_C_bit0(Tile_X0Y1_B_config_C_bit0),
    .B_config_C_bit1(Tile_X0Y1_B_config_C_bit1),
    .B_config_C_bit2(Tile_X0Y1_B_config_C_bit2),
    .B_config_C_bit3(Tile_X0Y1_B_config_C_bit3),
    .UserCLK(Tile_X0Y2_UserCLKo),
    .UserCLKo(Tile_X0Y1_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X0Y1_E1BEG[3] ,
    \Tile_X0Y1_E1BEG[2] ,
    \Tile_X0Y1_E1BEG[1] ,
    \Tile_X0Y1_E1BEG[0] }),
    .E2BEG({\Tile_X0Y1_E2BEG[7] ,
    \Tile_X0Y1_E2BEG[6] ,
    \Tile_X0Y1_E2BEG[5] ,
    \Tile_X0Y1_E2BEG[4] ,
    \Tile_X0Y1_E2BEG[3] ,
    \Tile_X0Y1_E2BEG[2] ,
    \Tile_X0Y1_E2BEG[1] ,
    \Tile_X0Y1_E2BEG[0] }),
    .E2BEGb({\Tile_X0Y1_E2BEGb[7] ,
    \Tile_X0Y1_E2BEGb[6] ,
    \Tile_X0Y1_E2BEGb[5] ,
    \Tile_X0Y1_E2BEGb[4] ,
    \Tile_X0Y1_E2BEGb[3] ,
    \Tile_X0Y1_E2BEGb[2] ,
    \Tile_X0Y1_E2BEGb[1] ,
    \Tile_X0Y1_E2BEGb[0] }),
    .E6BEG({\Tile_X0Y1_E6BEG[11] ,
    \Tile_X0Y1_E6BEG[10] ,
    \Tile_X0Y1_E6BEG[9] ,
    \Tile_X0Y1_E6BEG[8] ,
    \Tile_X0Y1_E6BEG[7] ,
    \Tile_X0Y1_E6BEG[6] ,
    \Tile_X0Y1_E6BEG[5] ,
    \Tile_X0Y1_E6BEG[4] ,
    \Tile_X0Y1_E6BEG[3] ,
    \Tile_X0Y1_E6BEG[2] ,
    \Tile_X0Y1_E6BEG[1] ,
    \Tile_X0Y1_E6BEG[0] }),
    .EE4BEG({\Tile_X0Y1_EE4BEG[15] ,
    \Tile_X0Y1_EE4BEG[14] ,
    \Tile_X0Y1_EE4BEG[13] ,
    \Tile_X0Y1_EE4BEG[12] ,
    \Tile_X0Y1_EE4BEG[11] ,
    \Tile_X0Y1_EE4BEG[10] ,
    \Tile_X0Y1_EE4BEG[9] ,
    \Tile_X0Y1_EE4BEG[8] ,
    \Tile_X0Y1_EE4BEG[7] ,
    \Tile_X0Y1_EE4BEG[6] ,
    \Tile_X0Y1_EE4BEG[5] ,
    \Tile_X0Y1_EE4BEG[4] ,
    \Tile_X0Y1_EE4BEG[3] ,
    \Tile_X0Y1_EE4BEG[2] ,
    \Tile_X0Y1_EE4BEG[1] ,
    \Tile_X0Y1_EE4BEG[0] }),
    .FrameData({FrameData[63],
    FrameData[62],
    FrameData[61],
    FrameData[60],
    FrameData[59],
    FrameData[58],
    FrameData[57],
    FrameData[56],
    FrameData[55],
    FrameData[54],
    FrameData[53],
    FrameData[52],
    FrameData[51],
    FrameData[50],
    FrameData[49],
    FrameData[48],
    FrameData[47],
    FrameData[46],
    FrameData[45],
    FrameData[44],
    FrameData[43],
    FrameData[42],
    FrameData[41],
    FrameData[40],
    FrameData[39],
    FrameData[38],
    FrameData[37],
    FrameData[36],
    FrameData[35],
    FrameData[34],
    FrameData[33],
    FrameData[32]}),
    .FrameData_O({\Tile_X0Y1_FrameData_O[31] ,
    \Tile_X0Y1_FrameData_O[30] ,
    \Tile_X0Y1_FrameData_O[29] ,
    \Tile_X0Y1_FrameData_O[28] ,
    \Tile_X0Y1_FrameData_O[27] ,
    \Tile_X0Y1_FrameData_O[26] ,
    \Tile_X0Y1_FrameData_O[25] ,
    \Tile_X0Y1_FrameData_O[24] ,
    \Tile_X0Y1_FrameData_O[23] ,
    \Tile_X0Y1_FrameData_O[22] ,
    \Tile_X0Y1_FrameData_O[21] ,
    \Tile_X0Y1_FrameData_O[20] ,
    \Tile_X0Y1_FrameData_O[19] ,
    \Tile_X0Y1_FrameData_O[18] ,
    \Tile_X0Y1_FrameData_O[17] ,
    \Tile_X0Y1_FrameData_O[16] ,
    \Tile_X0Y1_FrameData_O[15] ,
    \Tile_X0Y1_FrameData_O[14] ,
    \Tile_X0Y1_FrameData_O[13] ,
    \Tile_X0Y1_FrameData_O[12] ,
    \Tile_X0Y1_FrameData_O[11] ,
    \Tile_X0Y1_FrameData_O[10] ,
    \Tile_X0Y1_FrameData_O[9] ,
    \Tile_X0Y1_FrameData_O[8] ,
    \Tile_X0Y1_FrameData_O[7] ,
    \Tile_X0Y1_FrameData_O[6] ,
    \Tile_X0Y1_FrameData_O[5] ,
    \Tile_X0Y1_FrameData_O[4] ,
    \Tile_X0Y1_FrameData_O[3] ,
    \Tile_X0Y1_FrameData_O[2] ,
    \Tile_X0Y1_FrameData_O[1] ,
    \Tile_X0Y1_FrameData_O[0] }),
    .FrameStrobe({\Tile_X0Y2_FrameStrobe_O[19] ,
    \Tile_X0Y2_FrameStrobe_O[18] ,
    \Tile_X0Y2_FrameStrobe_O[17] ,
    \Tile_X0Y2_FrameStrobe_O[16] ,
    \Tile_X0Y2_FrameStrobe_O[15] ,
    \Tile_X0Y2_FrameStrobe_O[14] ,
    \Tile_X0Y2_FrameStrobe_O[13] ,
    \Tile_X0Y2_FrameStrobe_O[12] ,
    \Tile_X0Y2_FrameStrobe_O[11] ,
    \Tile_X0Y2_FrameStrobe_O[10] ,
    \Tile_X0Y2_FrameStrobe_O[9] ,
    \Tile_X0Y2_FrameStrobe_O[8] ,
    \Tile_X0Y2_FrameStrobe_O[7] ,
    \Tile_X0Y2_FrameStrobe_O[6] ,
    \Tile_X0Y2_FrameStrobe_O[5] ,
    \Tile_X0Y2_FrameStrobe_O[4] ,
    \Tile_X0Y2_FrameStrobe_O[3] ,
    \Tile_X0Y2_FrameStrobe_O[2] ,
    \Tile_X0Y2_FrameStrobe_O[1] ,
    \Tile_X0Y2_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X0Y1_FrameStrobe_O[19] ,
    \Tile_X0Y1_FrameStrobe_O[18] ,
    \Tile_X0Y1_FrameStrobe_O[17] ,
    \Tile_X0Y1_FrameStrobe_O[16] ,
    \Tile_X0Y1_FrameStrobe_O[15] ,
    \Tile_X0Y1_FrameStrobe_O[14] ,
    \Tile_X0Y1_FrameStrobe_O[13] ,
    \Tile_X0Y1_FrameStrobe_O[12] ,
    \Tile_X0Y1_FrameStrobe_O[11] ,
    \Tile_X0Y1_FrameStrobe_O[10] ,
    \Tile_X0Y1_FrameStrobe_O[9] ,
    \Tile_X0Y1_FrameStrobe_O[8] ,
    \Tile_X0Y1_FrameStrobe_O[7] ,
    \Tile_X0Y1_FrameStrobe_O[6] ,
    \Tile_X0Y1_FrameStrobe_O[5] ,
    \Tile_X0Y1_FrameStrobe_O[4] ,
    \Tile_X0Y1_FrameStrobe_O[3] ,
    \Tile_X0Y1_FrameStrobe_O[2] ,
    \Tile_X0Y1_FrameStrobe_O[1] ,
    \Tile_X0Y1_FrameStrobe_O[0] }),
    .W1END({\Tile_X1Y1_W1BEG[3] ,
    \Tile_X1Y1_W1BEG[2] ,
    \Tile_X1Y1_W1BEG[1] ,
    \Tile_X1Y1_W1BEG[0] }),
    .W2END({\Tile_X1Y1_W2BEGb[7] ,
    \Tile_X1Y1_W2BEGb[6] ,
    \Tile_X1Y1_W2BEGb[5] ,
    \Tile_X1Y1_W2BEGb[4] ,
    \Tile_X1Y1_W2BEGb[3] ,
    \Tile_X1Y1_W2BEGb[2] ,
    \Tile_X1Y1_W2BEGb[1] ,
    \Tile_X1Y1_W2BEGb[0] }),
    .W2MID({\Tile_X1Y1_W2BEG[7] ,
    \Tile_X1Y1_W2BEG[6] ,
    \Tile_X1Y1_W2BEG[5] ,
    \Tile_X1Y1_W2BEG[4] ,
    \Tile_X1Y1_W2BEG[3] ,
    \Tile_X1Y1_W2BEG[2] ,
    \Tile_X1Y1_W2BEG[1] ,
    \Tile_X1Y1_W2BEG[0] }),
    .W6END({\Tile_X1Y1_W6BEG[11] ,
    \Tile_X1Y1_W6BEG[10] ,
    \Tile_X1Y1_W6BEG[9] ,
    \Tile_X1Y1_W6BEG[8] ,
    \Tile_X1Y1_W6BEG[7] ,
    \Tile_X1Y1_W6BEG[6] ,
    \Tile_X1Y1_W6BEG[5] ,
    \Tile_X1Y1_W6BEG[4] ,
    \Tile_X1Y1_W6BEG[3] ,
    \Tile_X1Y1_W6BEG[2] ,
    \Tile_X1Y1_W6BEG[1] ,
    \Tile_X1Y1_W6BEG[0] }),
    .WW4END({\Tile_X1Y1_WW4BEG[15] ,
    \Tile_X1Y1_WW4BEG[14] ,
    \Tile_X1Y1_WW4BEG[13] ,
    \Tile_X1Y1_WW4BEG[12] ,
    \Tile_X1Y1_WW4BEG[11] ,
    \Tile_X1Y1_WW4BEG[10] ,
    \Tile_X1Y1_WW4BEG[9] ,
    \Tile_X1Y1_WW4BEG[8] ,
    \Tile_X1Y1_WW4BEG[7] ,
    \Tile_X1Y1_WW4BEG[6] ,
    \Tile_X1Y1_WW4BEG[5] ,
    \Tile_X1Y1_WW4BEG[4] ,
    \Tile_X1Y1_WW4BEG[3] ,
    \Tile_X1Y1_WW4BEG[2] ,
    \Tile_X1Y1_WW4BEG[1] ,
    \Tile_X1Y1_WW4BEG[0] }));
 W_IO Tile_X0Y2_W_IO (.A_I_top(Tile_X0Y2_A_I_top),
    .A_O_top(Tile_X0Y2_A_O_top),
    .A_T_top(Tile_X0Y2_A_T_top),
    .A_config_C_bit0(Tile_X0Y2_A_config_C_bit0),
    .A_config_C_bit1(Tile_X0Y2_A_config_C_bit1),
    .A_config_C_bit2(Tile_X0Y2_A_config_C_bit2),
    .A_config_C_bit3(Tile_X0Y2_A_config_C_bit3),
    .B_I_top(Tile_X0Y2_B_I_top),
    .B_O_top(Tile_X0Y2_B_O_top),
    .B_T_top(Tile_X0Y2_B_T_top),
    .B_config_C_bit0(Tile_X0Y2_B_config_C_bit0),
    .B_config_C_bit1(Tile_X0Y2_B_config_C_bit1),
    .B_config_C_bit2(Tile_X0Y2_B_config_C_bit2),
    .B_config_C_bit3(Tile_X0Y2_B_config_C_bit3),
    .UserCLK(Tile_X0Y3_UserCLKo),
    .UserCLKo(Tile_X0Y2_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X0Y2_E1BEG[3] ,
    \Tile_X0Y2_E1BEG[2] ,
    \Tile_X0Y2_E1BEG[1] ,
    \Tile_X0Y2_E1BEG[0] }),
    .E2BEG({\Tile_X0Y2_E2BEG[7] ,
    \Tile_X0Y2_E2BEG[6] ,
    \Tile_X0Y2_E2BEG[5] ,
    \Tile_X0Y2_E2BEG[4] ,
    \Tile_X0Y2_E2BEG[3] ,
    \Tile_X0Y2_E2BEG[2] ,
    \Tile_X0Y2_E2BEG[1] ,
    \Tile_X0Y2_E2BEG[0] }),
    .E2BEGb({\Tile_X0Y2_E2BEGb[7] ,
    \Tile_X0Y2_E2BEGb[6] ,
    \Tile_X0Y2_E2BEGb[5] ,
    \Tile_X0Y2_E2BEGb[4] ,
    \Tile_X0Y2_E2BEGb[3] ,
    \Tile_X0Y2_E2BEGb[2] ,
    \Tile_X0Y2_E2BEGb[1] ,
    \Tile_X0Y2_E2BEGb[0] }),
    .E6BEG({\Tile_X0Y2_E6BEG[11] ,
    \Tile_X0Y2_E6BEG[10] ,
    \Tile_X0Y2_E6BEG[9] ,
    \Tile_X0Y2_E6BEG[8] ,
    \Tile_X0Y2_E6BEG[7] ,
    \Tile_X0Y2_E6BEG[6] ,
    \Tile_X0Y2_E6BEG[5] ,
    \Tile_X0Y2_E6BEG[4] ,
    \Tile_X0Y2_E6BEG[3] ,
    \Tile_X0Y2_E6BEG[2] ,
    \Tile_X0Y2_E6BEG[1] ,
    \Tile_X0Y2_E6BEG[0] }),
    .EE4BEG({\Tile_X0Y2_EE4BEG[15] ,
    \Tile_X0Y2_EE4BEG[14] ,
    \Tile_X0Y2_EE4BEG[13] ,
    \Tile_X0Y2_EE4BEG[12] ,
    \Tile_X0Y2_EE4BEG[11] ,
    \Tile_X0Y2_EE4BEG[10] ,
    \Tile_X0Y2_EE4BEG[9] ,
    \Tile_X0Y2_EE4BEG[8] ,
    \Tile_X0Y2_EE4BEG[7] ,
    \Tile_X0Y2_EE4BEG[6] ,
    \Tile_X0Y2_EE4BEG[5] ,
    \Tile_X0Y2_EE4BEG[4] ,
    \Tile_X0Y2_EE4BEG[3] ,
    \Tile_X0Y2_EE4BEG[2] ,
    \Tile_X0Y2_EE4BEG[1] ,
    \Tile_X0Y2_EE4BEG[0] }),
    .FrameData({FrameData[95],
    FrameData[94],
    FrameData[93],
    FrameData[92],
    FrameData[91],
    FrameData[90],
    FrameData[89],
    FrameData[88],
    FrameData[87],
    FrameData[86],
    FrameData[85],
    FrameData[84],
    FrameData[83],
    FrameData[82],
    FrameData[81],
    FrameData[80],
    FrameData[79],
    FrameData[78],
    FrameData[77],
    FrameData[76],
    FrameData[75],
    FrameData[74],
    FrameData[73],
    FrameData[72],
    FrameData[71],
    FrameData[70],
    FrameData[69],
    FrameData[68],
    FrameData[67],
    FrameData[66],
    FrameData[65],
    FrameData[64]}),
    .FrameData_O({\Tile_X0Y2_FrameData_O[31] ,
    \Tile_X0Y2_FrameData_O[30] ,
    \Tile_X0Y2_FrameData_O[29] ,
    \Tile_X0Y2_FrameData_O[28] ,
    \Tile_X0Y2_FrameData_O[27] ,
    \Tile_X0Y2_FrameData_O[26] ,
    \Tile_X0Y2_FrameData_O[25] ,
    \Tile_X0Y2_FrameData_O[24] ,
    \Tile_X0Y2_FrameData_O[23] ,
    \Tile_X0Y2_FrameData_O[22] ,
    \Tile_X0Y2_FrameData_O[21] ,
    \Tile_X0Y2_FrameData_O[20] ,
    \Tile_X0Y2_FrameData_O[19] ,
    \Tile_X0Y2_FrameData_O[18] ,
    \Tile_X0Y2_FrameData_O[17] ,
    \Tile_X0Y2_FrameData_O[16] ,
    \Tile_X0Y2_FrameData_O[15] ,
    \Tile_X0Y2_FrameData_O[14] ,
    \Tile_X0Y2_FrameData_O[13] ,
    \Tile_X0Y2_FrameData_O[12] ,
    \Tile_X0Y2_FrameData_O[11] ,
    \Tile_X0Y2_FrameData_O[10] ,
    \Tile_X0Y2_FrameData_O[9] ,
    \Tile_X0Y2_FrameData_O[8] ,
    \Tile_X0Y2_FrameData_O[7] ,
    \Tile_X0Y2_FrameData_O[6] ,
    \Tile_X0Y2_FrameData_O[5] ,
    \Tile_X0Y2_FrameData_O[4] ,
    \Tile_X0Y2_FrameData_O[3] ,
    \Tile_X0Y2_FrameData_O[2] ,
    \Tile_X0Y2_FrameData_O[1] ,
    \Tile_X0Y2_FrameData_O[0] }),
    .FrameStrobe({\Tile_X0Y3_FrameStrobe_O[19] ,
    \Tile_X0Y3_FrameStrobe_O[18] ,
    \Tile_X0Y3_FrameStrobe_O[17] ,
    \Tile_X0Y3_FrameStrobe_O[16] ,
    \Tile_X0Y3_FrameStrobe_O[15] ,
    \Tile_X0Y3_FrameStrobe_O[14] ,
    \Tile_X0Y3_FrameStrobe_O[13] ,
    \Tile_X0Y3_FrameStrobe_O[12] ,
    \Tile_X0Y3_FrameStrobe_O[11] ,
    \Tile_X0Y3_FrameStrobe_O[10] ,
    \Tile_X0Y3_FrameStrobe_O[9] ,
    \Tile_X0Y3_FrameStrobe_O[8] ,
    \Tile_X0Y3_FrameStrobe_O[7] ,
    \Tile_X0Y3_FrameStrobe_O[6] ,
    \Tile_X0Y3_FrameStrobe_O[5] ,
    \Tile_X0Y3_FrameStrobe_O[4] ,
    \Tile_X0Y3_FrameStrobe_O[3] ,
    \Tile_X0Y3_FrameStrobe_O[2] ,
    \Tile_X0Y3_FrameStrobe_O[1] ,
    \Tile_X0Y3_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X0Y2_FrameStrobe_O[19] ,
    \Tile_X0Y2_FrameStrobe_O[18] ,
    \Tile_X0Y2_FrameStrobe_O[17] ,
    \Tile_X0Y2_FrameStrobe_O[16] ,
    \Tile_X0Y2_FrameStrobe_O[15] ,
    \Tile_X0Y2_FrameStrobe_O[14] ,
    \Tile_X0Y2_FrameStrobe_O[13] ,
    \Tile_X0Y2_FrameStrobe_O[12] ,
    \Tile_X0Y2_FrameStrobe_O[11] ,
    \Tile_X0Y2_FrameStrobe_O[10] ,
    \Tile_X0Y2_FrameStrobe_O[9] ,
    \Tile_X0Y2_FrameStrobe_O[8] ,
    \Tile_X0Y2_FrameStrobe_O[7] ,
    \Tile_X0Y2_FrameStrobe_O[6] ,
    \Tile_X0Y2_FrameStrobe_O[5] ,
    \Tile_X0Y2_FrameStrobe_O[4] ,
    \Tile_X0Y2_FrameStrobe_O[3] ,
    \Tile_X0Y2_FrameStrobe_O[2] ,
    \Tile_X0Y2_FrameStrobe_O[1] ,
    \Tile_X0Y2_FrameStrobe_O[0] }),
    .W1END({\Tile_X1Y2_W1BEG[3] ,
    \Tile_X1Y2_W1BEG[2] ,
    \Tile_X1Y2_W1BEG[1] ,
    \Tile_X1Y2_W1BEG[0] }),
    .W2END({\Tile_X1Y2_W2BEGb[7] ,
    \Tile_X1Y2_W2BEGb[6] ,
    \Tile_X1Y2_W2BEGb[5] ,
    \Tile_X1Y2_W2BEGb[4] ,
    \Tile_X1Y2_W2BEGb[3] ,
    \Tile_X1Y2_W2BEGb[2] ,
    \Tile_X1Y2_W2BEGb[1] ,
    \Tile_X1Y2_W2BEGb[0] }),
    .W2MID({\Tile_X1Y2_W2BEG[7] ,
    \Tile_X1Y2_W2BEG[6] ,
    \Tile_X1Y2_W2BEG[5] ,
    \Tile_X1Y2_W2BEG[4] ,
    \Tile_X1Y2_W2BEG[3] ,
    \Tile_X1Y2_W2BEG[2] ,
    \Tile_X1Y2_W2BEG[1] ,
    \Tile_X1Y2_W2BEG[0] }),
    .W6END({\Tile_X1Y2_W6BEG[11] ,
    \Tile_X1Y2_W6BEG[10] ,
    \Tile_X1Y2_W6BEG[9] ,
    \Tile_X1Y2_W6BEG[8] ,
    \Tile_X1Y2_W6BEG[7] ,
    \Tile_X1Y2_W6BEG[6] ,
    \Tile_X1Y2_W6BEG[5] ,
    \Tile_X1Y2_W6BEG[4] ,
    \Tile_X1Y2_W6BEG[3] ,
    \Tile_X1Y2_W6BEG[2] ,
    \Tile_X1Y2_W6BEG[1] ,
    \Tile_X1Y2_W6BEG[0] }),
    .WW4END({\Tile_X1Y2_WW4BEG[15] ,
    \Tile_X1Y2_WW4BEG[14] ,
    \Tile_X1Y2_WW4BEG[13] ,
    \Tile_X1Y2_WW4BEG[12] ,
    \Tile_X1Y2_WW4BEG[11] ,
    \Tile_X1Y2_WW4BEG[10] ,
    \Tile_X1Y2_WW4BEG[9] ,
    \Tile_X1Y2_WW4BEG[8] ,
    \Tile_X1Y2_WW4BEG[7] ,
    \Tile_X1Y2_WW4BEG[6] ,
    \Tile_X1Y2_WW4BEG[5] ,
    \Tile_X1Y2_WW4BEG[4] ,
    \Tile_X1Y2_WW4BEG[3] ,
    \Tile_X1Y2_WW4BEG[2] ,
    \Tile_X1Y2_WW4BEG[1] ,
    \Tile_X1Y2_WW4BEG[0] }));
 W_IO Tile_X0Y3_W_IO (.A_I_top(Tile_X0Y3_A_I_top),
    .A_O_top(Tile_X0Y3_A_O_top),
    .A_T_top(Tile_X0Y3_A_T_top),
    .A_config_C_bit0(Tile_X0Y3_A_config_C_bit0),
    .A_config_C_bit1(Tile_X0Y3_A_config_C_bit1),
    .A_config_C_bit2(Tile_X0Y3_A_config_C_bit2),
    .A_config_C_bit3(Tile_X0Y3_A_config_C_bit3),
    .B_I_top(Tile_X0Y3_B_I_top),
    .B_O_top(Tile_X0Y3_B_O_top),
    .B_T_top(Tile_X0Y3_B_T_top),
    .B_config_C_bit0(Tile_X0Y3_B_config_C_bit0),
    .B_config_C_bit1(Tile_X0Y3_B_config_C_bit1),
    .B_config_C_bit2(Tile_X0Y3_B_config_C_bit2),
    .B_config_C_bit3(Tile_X0Y3_B_config_C_bit3),
    .UserCLK(Tile_X0Y4_UserCLKo),
    .UserCLKo(Tile_X0Y3_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X0Y3_E1BEG[3] ,
    \Tile_X0Y3_E1BEG[2] ,
    \Tile_X0Y3_E1BEG[1] ,
    \Tile_X0Y3_E1BEG[0] }),
    .E2BEG({\Tile_X0Y3_E2BEG[7] ,
    \Tile_X0Y3_E2BEG[6] ,
    \Tile_X0Y3_E2BEG[5] ,
    \Tile_X0Y3_E2BEG[4] ,
    \Tile_X0Y3_E2BEG[3] ,
    \Tile_X0Y3_E2BEG[2] ,
    \Tile_X0Y3_E2BEG[1] ,
    \Tile_X0Y3_E2BEG[0] }),
    .E2BEGb({\Tile_X0Y3_E2BEGb[7] ,
    \Tile_X0Y3_E2BEGb[6] ,
    \Tile_X0Y3_E2BEGb[5] ,
    \Tile_X0Y3_E2BEGb[4] ,
    \Tile_X0Y3_E2BEGb[3] ,
    \Tile_X0Y3_E2BEGb[2] ,
    \Tile_X0Y3_E2BEGb[1] ,
    \Tile_X0Y3_E2BEGb[0] }),
    .E6BEG({\Tile_X0Y3_E6BEG[11] ,
    \Tile_X0Y3_E6BEG[10] ,
    \Tile_X0Y3_E6BEG[9] ,
    \Tile_X0Y3_E6BEG[8] ,
    \Tile_X0Y3_E6BEG[7] ,
    \Tile_X0Y3_E6BEG[6] ,
    \Tile_X0Y3_E6BEG[5] ,
    \Tile_X0Y3_E6BEG[4] ,
    \Tile_X0Y3_E6BEG[3] ,
    \Tile_X0Y3_E6BEG[2] ,
    \Tile_X0Y3_E6BEG[1] ,
    \Tile_X0Y3_E6BEG[0] }),
    .EE4BEG({\Tile_X0Y3_EE4BEG[15] ,
    \Tile_X0Y3_EE4BEG[14] ,
    \Tile_X0Y3_EE4BEG[13] ,
    \Tile_X0Y3_EE4BEG[12] ,
    \Tile_X0Y3_EE4BEG[11] ,
    \Tile_X0Y3_EE4BEG[10] ,
    \Tile_X0Y3_EE4BEG[9] ,
    \Tile_X0Y3_EE4BEG[8] ,
    \Tile_X0Y3_EE4BEG[7] ,
    \Tile_X0Y3_EE4BEG[6] ,
    \Tile_X0Y3_EE4BEG[5] ,
    \Tile_X0Y3_EE4BEG[4] ,
    \Tile_X0Y3_EE4BEG[3] ,
    \Tile_X0Y3_EE4BEG[2] ,
    \Tile_X0Y3_EE4BEG[1] ,
    \Tile_X0Y3_EE4BEG[0] }),
    .FrameData({FrameData[127],
    FrameData[126],
    FrameData[125],
    FrameData[124],
    FrameData[123],
    FrameData[122],
    FrameData[121],
    FrameData[120],
    FrameData[119],
    FrameData[118],
    FrameData[117],
    FrameData[116],
    FrameData[115],
    FrameData[114],
    FrameData[113],
    FrameData[112],
    FrameData[111],
    FrameData[110],
    FrameData[109],
    FrameData[108],
    FrameData[107],
    FrameData[106],
    FrameData[105],
    FrameData[104],
    FrameData[103],
    FrameData[102],
    FrameData[101],
    FrameData[100],
    FrameData[99],
    FrameData[98],
    FrameData[97],
    FrameData[96]}),
    .FrameData_O({\Tile_X0Y3_FrameData_O[31] ,
    \Tile_X0Y3_FrameData_O[30] ,
    \Tile_X0Y3_FrameData_O[29] ,
    \Tile_X0Y3_FrameData_O[28] ,
    \Tile_X0Y3_FrameData_O[27] ,
    \Tile_X0Y3_FrameData_O[26] ,
    \Tile_X0Y3_FrameData_O[25] ,
    \Tile_X0Y3_FrameData_O[24] ,
    \Tile_X0Y3_FrameData_O[23] ,
    \Tile_X0Y3_FrameData_O[22] ,
    \Tile_X0Y3_FrameData_O[21] ,
    \Tile_X0Y3_FrameData_O[20] ,
    \Tile_X0Y3_FrameData_O[19] ,
    \Tile_X0Y3_FrameData_O[18] ,
    \Tile_X0Y3_FrameData_O[17] ,
    \Tile_X0Y3_FrameData_O[16] ,
    \Tile_X0Y3_FrameData_O[15] ,
    \Tile_X0Y3_FrameData_O[14] ,
    \Tile_X0Y3_FrameData_O[13] ,
    \Tile_X0Y3_FrameData_O[12] ,
    \Tile_X0Y3_FrameData_O[11] ,
    \Tile_X0Y3_FrameData_O[10] ,
    \Tile_X0Y3_FrameData_O[9] ,
    \Tile_X0Y3_FrameData_O[8] ,
    \Tile_X0Y3_FrameData_O[7] ,
    \Tile_X0Y3_FrameData_O[6] ,
    \Tile_X0Y3_FrameData_O[5] ,
    \Tile_X0Y3_FrameData_O[4] ,
    \Tile_X0Y3_FrameData_O[3] ,
    \Tile_X0Y3_FrameData_O[2] ,
    \Tile_X0Y3_FrameData_O[1] ,
    \Tile_X0Y3_FrameData_O[0] }),
    .FrameStrobe({\Tile_X0Y4_FrameStrobe_O[19] ,
    \Tile_X0Y4_FrameStrobe_O[18] ,
    \Tile_X0Y4_FrameStrobe_O[17] ,
    \Tile_X0Y4_FrameStrobe_O[16] ,
    \Tile_X0Y4_FrameStrobe_O[15] ,
    \Tile_X0Y4_FrameStrobe_O[14] ,
    \Tile_X0Y4_FrameStrobe_O[13] ,
    \Tile_X0Y4_FrameStrobe_O[12] ,
    \Tile_X0Y4_FrameStrobe_O[11] ,
    \Tile_X0Y4_FrameStrobe_O[10] ,
    \Tile_X0Y4_FrameStrobe_O[9] ,
    \Tile_X0Y4_FrameStrobe_O[8] ,
    \Tile_X0Y4_FrameStrobe_O[7] ,
    \Tile_X0Y4_FrameStrobe_O[6] ,
    \Tile_X0Y4_FrameStrobe_O[5] ,
    \Tile_X0Y4_FrameStrobe_O[4] ,
    \Tile_X0Y4_FrameStrobe_O[3] ,
    \Tile_X0Y4_FrameStrobe_O[2] ,
    \Tile_X0Y4_FrameStrobe_O[1] ,
    \Tile_X0Y4_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X0Y3_FrameStrobe_O[19] ,
    \Tile_X0Y3_FrameStrobe_O[18] ,
    \Tile_X0Y3_FrameStrobe_O[17] ,
    \Tile_X0Y3_FrameStrobe_O[16] ,
    \Tile_X0Y3_FrameStrobe_O[15] ,
    \Tile_X0Y3_FrameStrobe_O[14] ,
    \Tile_X0Y3_FrameStrobe_O[13] ,
    \Tile_X0Y3_FrameStrobe_O[12] ,
    \Tile_X0Y3_FrameStrobe_O[11] ,
    \Tile_X0Y3_FrameStrobe_O[10] ,
    \Tile_X0Y3_FrameStrobe_O[9] ,
    \Tile_X0Y3_FrameStrobe_O[8] ,
    \Tile_X0Y3_FrameStrobe_O[7] ,
    \Tile_X0Y3_FrameStrobe_O[6] ,
    \Tile_X0Y3_FrameStrobe_O[5] ,
    \Tile_X0Y3_FrameStrobe_O[4] ,
    \Tile_X0Y3_FrameStrobe_O[3] ,
    \Tile_X0Y3_FrameStrobe_O[2] ,
    \Tile_X0Y3_FrameStrobe_O[1] ,
    \Tile_X0Y3_FrameStrobe_O[0] }),
    .W1END({\Tile_X1Y3_W1BEG[3] ,
    \Tile_X1Y3_W1BEG[2] ,
    \Tile_X1Y3_W1BEG[1] ,
    \Tile_X1Y3_W1BEG[0] }),
    .W2END({\Tile_X1Y3_W2BEGb[7] ,
    \Tile_X1Y3_W2BEGb[6] ,
    \Tile_X1Y3_W2BEGb[5] ,
    \Tile_X1Y3_W2BEGb[4] ,
    \Tile_X1Y3_W2BEGb[3] ,
    \Tile_X1Y3_W2BEGb[2] ,
    \Tile_X1Y3_W2BEGb[1] ,
    \Tile_X1Y3_W2BEGb[0] }),
    .W2MID({\Tile_X1Y3_W2BEG[7] ,
    \Tile_X1Y3_W2BEG[6] ,
    \Tile_X1Y3_W2BEG[5] ,
    \Tile_X1Y3_W2BEG[4] ,
    \Tile_X1Y3_W2BEG[3] ,
    \Tile_X1Y3_W2BEG[2] ,
    \Tile_X1Y3_W2BEG[1] ,
    \Tile_X1Y3_W2BEG[0] }),
    .W6END({\Tile_X1Y3_W6BEG[11] ,
    \Tile_X1Y3_W6BEG[10] ,
    \Tile_X1Y3_W6BEG[9] ,
    \Tile_X1Y3_W6BEG[8] ,
    \Tile_X1Y3_W6BEG[7] ,
    \Tile_X1Y3_W6BEG[6] ,
    \Tile_X1Y3_W6BEG[5] ,
    \Tile_X1Y3_W6BEG[4] ,
    \Tile_X1Y3_W6BEG[3] ,
    \Tile_X1Y3_W6BEG[2] ,
    \Tile_X1Y3_W6BEG[1] ,
    \Tile_X1Y3_W6BEG[0] }),
    .WW4END({\Tile_X1Y3_WW4BEG[15] ,
    \Tile_X1Y3_WW4BEG[14] ,
    \Tile_X1Y3_WW4BEG[13] ,
    \Tile_X1Y3_WW4BEG[12] ,
    \Tile_X1Y3_WW4BEG[11] ,
    \Tile_X1Y3_WW4BEG[10] ,
    \Tile_X1Y3_WW4BEG[9] ,
    \Tile_X1Y3_WW4BEG[8] ,
    \Tile_X1Y3_WW4BEG[7] ,
    \Tile_X1Y3_WW4BEG[6] ,
    \Tile_X1Y3_WW4BEG[5] ,
    \Tile_X1Y3_WW4BEG[4] ,
    \Tile_X1Y3_WW4BEG[3] ,
    \Tile_X1Y3_WW4BEG[2] ,
    \Tile_X1Y3_WW4BEG[1] ,
    \Tile_X1Y3_WW4BEG[0] }));
 W_IO Tile_X0Y4_W_IO (.A_I_top(Tile_X0Y4_A_I_top),
    .A_O_top(Tile_X0Y4_A_O_top),
    .A_T_top(Tile_X0Y4_A_T_top),
    .A_config_C_bit0(Tile_X0Y4_A_config_C_bit0),
    .A_config_C_bit1(Tile_X0Y4_A_config_C_bit1),
    .A_config_C_bit2(Tile_X0Y4_A_config_C_bit2),
    .A_config_C_bit3(Tile_X0Y4_A_config_C_bit3),
    .B_I_top(Tile_X0Y4_B_I_top),
    .B_O_top(Tile_X0Y4_B_O_top),
    .B_T_top(Tile_X0Y4_B_T_top),
    .B_config_C_bit0(Tile_X0Y4_B_config_C_bit0),
    .B_config_C_bit1(Tile_X0Y4_B_config_C_bit1),
    .B_config_C_bit2(Tile_X0Y4_B_config_C_bit2),
    .B_config_C_bit3(Tile_X0Y4_B_config_C_bit3),
    .UserCLK(Tile_X0Y5_UserCLKo),
    .UserCLKo(Tile_X0Y4_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X0Y4_E1BEG[3] ,
    \Tile_X0Y4_E1BEG[2] ,
    \Tile_X0Y4_E1BEG[1] ,
    \Tile_X0Y4_E1BEG[0] }),
    .E2BEG({\Tile_X0Y4_E2BEG[7] ,
    \Tile_X0Y4_E2BEG[6] ,
    \Tile_X0Y4_E2BEG[5] ,
    \Tile_X0Y4_E2BEG[4] ,
    \Tile_X0Y4_E2BEG[3] ,
    \Tile_X0Y4_E2BEG[2] ,
    \Tile_X0Y4_E2BEG[1] ,
    \Tile_X0Y4_E2BEG[0] }),
    .E2BEGb({\Tile_X0Y4_E2BEGb[7] ,
    \Tile_X0Y4_E2BEGb[6] ,
    \Tile_X0Y4_E2BEGb[5] ,
    \Tile_X0Y4_E2BEGb[4] ,
    \Tile_X0Y4_E2BEGb[3] ,
    \Tile_X0Y4_E2BEGb[2] ,
    \Tile_X0Y4_E2BEGb[1] ,
    \Tile_X0Y4_E2BEGb[0] }),
    .E6BEG({\Tile_X0Y4_E6BEG[11] ,
    \Tile_X0Y4_E6BEG[10] ,
    \Tile_X0Y4_E6BEG[9] ,
    \Tile_X0Y4_E6BEG[8] ,
    \Tile_X0Y4_E6BEG[7] ,
    \Tile_X0Y4_E6BEG[6] ,
    \Tile_X0Y4_E6BEG[5] ,
    \Tile_X0Y4_E6BEG[4] ,
    \Tile_X0Y4_E6BEG[3] ,
    \Tile_X0Y4_E6BEG[2] ,
    \Tile_X0Y4_E6BEG[1] ,
    \Tile_X0Y4_E6BEG[0] }),
    .EE4BEG({\Tile_X0Y4_EE4BEG[15] ,
    \Tile_X0Y4_EE4BEG[14] ,
    \Tile_X0Y4_EE4BEG[13] ,
    \Tile_X0Y4_EE4BEG[12] ,
    \Tile_X0Y4_EE4BEG[11] ,
    \Tile_X0Y4_EE4BEG[10] ,
    \Tile_X0Y4_EE4BEG[9] ,
    \Tile_X0Y4_EE4BEG[8] ,
    \Tile_X0Y4_EE4BEG[7] ,
    \Tile_X0Y4_EE4BEG[6] ,
    \Tile_X0Y4_EE4BEG[5] ,
    \Tile_X0Y4_EE4BEG[4] ,
    \Tile_X0Y4_EE4BEG[3] ,
    \Tile_X0Y4_EE4BEG[2] ,
    \Tile_X0Y4_EE4BEG[1] ,
    \Tile_X0Y4_EE4BEG[0] }),
    .FrameData({FrameData[159],
    FrameData[158],
    FrameData[157],
    FrameData[156],
    FrameData[155],
    FrameData[154],
    FrameData[153],
    FrameData[152],
    FrameData[151],
    FrameData[150],
    FrameData[149],
    FrameData[148],
    FrameData[147],
    FrameData[146],
    FrameData[145],
    FrameData[144],
    FrameData[143],
    FrameData[142],
    FrameData[141],
    FrameData[140],
    FrameData[139],
    FrameData[138],
    FrameData[137],
    FrameData[136],
    FrameData[135],
    FrameData[134],
    FrameData[133],
    FrameData[132],
    FrameData[131],
    FrameData[130],
    FrameData[129],
    FrameData[128]}),
    .FrameData_O({\Tile_X0Y4_FrameData_O[31] ,
    \Tile_X0Y4_FrameData_O[30] ,
    \Tile_X0Y4_FrameData_O[29] ,
    \Tile_X0Y4_FrameData_O[28] ,
    \Tile_X0Y4_FrameData_O[27] ,
    \Tile_X0Y4_FrameData_O[26] ,
    \Tile_X0Y4_FrameData_O[25] ,
    \Tile_X0Y4_FrameData_O[24] ,
    \Tile_X0Y4_FrameData_O[23] ,
    \Tile_X0Y4_FrameData_O[22] ,
    \Tile_X0Y4_FrameData_O[21] ,
    \Tile_X0Y4_FrameData_O[20] ,
    \Tile_X0Y4_FrameData_O[19] ,
    \Tile_X0Y4_FrameData_O[18] ,
    \Tile_X0Y4_FrameData_O[17] ,
    \Tile_X0Y4_FrameData_O[16] ,
    \Tile_X0Y4_FrameData_O[15] ,
    \Tile_X0Y4_FrameData_O[14] ,
    \Tile_X0Y4_FrameData_O[13] ,
    \Tile_X0Y4_FrameData_O[12] ,
    \Tile_X0Y4_FrameData_O[11] ,
    \Tile_X0Y4_FrameData_O[10] ,
    \Tile_X0Y4_FrameData_O[9] ,
    \Tile_X0Y4_FrameData_O[8] ,
    \Tile_X0Y4_FrameData_O[7] ,
    \Tile_X0Y4_FrameData_O[6] ,
    \Tile_X0Y4_FrameData_O[5] ,
    \Tile_X0Y4_FrameData_O[4] ,
    \Tile_X0Y4_FrameData_O[3] ,
    \Tile_X0Y4_FrameData_O[2] ,
    \Tile_X0Y4_FrameData_O[1] ,
    \Tile_X0Y4_FrameData_O[0] }),
    .FrameStrobe({\Tile_X0Y5_FrameStrobe_O[19] ,
    \Tile_X0Y5_FrameStrobe_O[18] ,
    \Tile_X0Y5_FrameStrobe_O[17] ,
    \Tile_X0Y5_FrameStrobe_O[16] ,
    \Tile_X0Y5_FrameStrobe_O[15] ,
    \Tile_X0Y5_FrameStrobe_O[14] ,
    \Tile_X0Y5_FrameStrobe_O[13] ,
    \Tile_X0Y5_FrameStrobe_O[12] ,
    \Tile_X0Y5_FrameStrobe_O[11] ,
    \Tile_X0Y5_FrameStrobe_O[10] ,
    \Tile_X0Y5_FrameStrobe_O[9] ,
    \Tile_X0Y5_FrameStrobe_O[8] ,
    \Tile_X0Y5_FrameStrobe_O[7] ,
    \Tile_X0Y5_FrameStrobe_O[6] ,
    \Tile_X0Y5_FrameStrobe_O[5] ,
    \Tile_X0Y5_FrameStrobe_O[4] ,
    \Tile_X0Y5_FrameStrobe_O[3] ,
    \Tile_X0Y5_FrameStrobe_O[2] ,
    \Tile_X0Y5_FrameStrobe_O[1] ,
    \Tile_X0Y5_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X0Y4_FrameStrobe_O[19] ,
    \Tile_X0Y4_FrameStrobe_O[18] ,
    \Tile_X0Y4_FrameStrobe_O[17] ,
    \Tile_X0Y4_FrameStrobe_O[16] ,
    \Tile_X0Y4_FrameStrobe_O[15] ,
    \Tile_X0Y4_FrameStrobe_O[14] ,
    \Tile_X0Y4_FrameStrobe_O[13] ,
    \Tile_X0Y4_FrameStrobe_O[12] ,
    \Tile_X0Y4_FrameStrobe_O[11] ,
    \Tile_X0Y4_FrameStrobe_O[10] ,
    \Tile_X0Y4_FrameStrobe_O[9] ,
    \Tile_X0Y4_FrameStrobe_O[8] ,
    \Tile_X0Y4_FrameStrobe_O[7] ,
    \Tile_X0Y4_FrameStrobe_O[6] ,
    \Tile_X0Y4_FrameStrobe_O[5] ,
    \Tile_X0Y4_FrameStrobe_O[4] ,
    \Tile_X0Y4_FrameStrobe_O[3] ,
    \Tile_X0Y4_FrameStrobe_O[2] ,
    \Tile_X0Y4_FrameStrobe_O[1] ,
    \Tile_X0Y4_FrameStrobe_O[0] }),
    .W1END({\Tile_X1Y4_W1BEG[3] ,
    \Tile_X1Y4_W1BEG[2] ,
    \Tile_X1Y4_W1BEG[1] ,
    \Tile_X1Y4_W1BEG[0] }),
    .W2END({\Tile_X1Y4_W2BEGb[7] ,
    \Tile_X1Y4_W2BEGb[6] ,
    \Tile_X1Y4_W2BEGb[5] ,
    \Tile_X1Y4_W2BEGb[4] ,
    \Tile_X1Y4_W2BEGb[3] ,
    \Tile_X1Y4_W2BEGb[2] ,
    \Tile_X1Y4_W2BEGb[1] ,
    \Tile_X1Y4_W2BEGb[0] }),
    .W2MID({\Tile_X1Y4_W2BEG[7] ,
    \Tile_X1Y4_W2BEG[6] ,
    \Tile_X1Y4_W2BEG[5] ,
    \Tile_X1Y4_W2BEG[4] ,
    \Tile_X1Y4_W2BEG[3] ,
    \Tile_X1Y4_W2BEG[2] ,
    \Tile_X1Y4_W2BEG[1] ,
    \Tile_X1Y4_W2BEG[0] }),
    .W6END({\Tile_X1Y4_W6BEG[11] ,
    \Tile_X1Y4_W6BEG[10] ,
    \Tile_X1Y4_W6BEG[9] ,
    \Tile_X1Y4_W6BEG[8] ,
    \Tile_X1Y4_W6BEG[7] ,
    \Tile_X1Y4_W6BEG[6] ,
    \Tile_X1Y4_W6BEG[5] ,
    \Tile_X1Y4_W6BEG[4] ,
    \Tile_X1Y4_W6BEG[3] ,
    \Tile_X1Y4_W6BEG[2] ,
    \Tile_X1Y4_W6BEG[1] ,
    \Tile_X1Y4_W6BEG[0] }),
    .WW4END({\Tile_X1Y4_WW4BEG[15] ,
    \Tile_X1Y4_WW4BEG[14] ,
    \Tile_X1Y4_WW4BEG[13] ,
    \Tile_X1Y4_WW4BEG[12] ,
    \Tile_X1Y4_WW4BEG[11] ,
    \Tile_X1Y4_WW4BEG[10] ,
    \Tile_X1Y4_WW4BEG[9] ,
    \Tile_X1Y4_WW4BEG[8] ,
    \Tile_X1Y4_WW4BEG[7] ,
    \Tile_X1Y4_WW4BEG[6] ,
    \Tile_X1Y4_WW4BEG[5] ,
    \Tile_X1Y4_WW4BEG[4] ,
    \Tile_X1Y4_WW4BEG[3] ,
    \Tile_X1Y4_WW4BEG[2] ,
    \Tile_X1Y4_WW4BEG[1] ,
    \Tile_X1Y4_WW4BEG[0] }));
 W_IO Tile_X0Y5_W_IO (.A_I_top(Tile_X0Y5_A_I_top),
    .A_O_top(Tile_X0Y5_A_O_top),
    .A_T_top(Tile_X0Y5_A_T_top),
    .A_config_C_bit0(Tile_X0Y5_A_config_C_bit0),
    .A_config_C_bit1(Tile_X0Y5_A_config_C_bit1),
    .A_config_C_bit2(Tile_X0Y5_A_config_C_bit2),
    .A_config_C_bit3(Tile_X0Y5_A_config_C_bit3),
    .B_I_top(Tile_X0Y5_B_I_top),
    .B_O_top(Tile_X0Y5_B_O_top),
    .B_T_top(Tile_X0Y5_B_T_top),
    .B_config_C_bit0(Tile_X0Y5_B_config_C_bit0),
    .B_config_C_bit1(Tile_X0Y5_B_config_C_bit1),
    .B_config_C_bit2(Tile_X0Y5_B_config_C_bit2),
    .B_config_C_bit3(Tile_X0Y5_B_config_C_bit3),
    .UserCLK(Tile_X0Y6_UserCLKo),
    .UserCLKo(Tile_X0Y5_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X0Y5_E1BEG[3] ,
    \Tile_X0Y5_E1BEG[2] ,
    \Tile_X0Y5_E1BEG[1] ,
    \Tile_X0Y5_E1BEG[0] }),
    .E2BEG({\Tile_X0Y5_E2BEG[7] ,
    \Tile_X0Y5_E2BEG[6] ,
    \Tile_X0Y5_E2BEG[5] ,
    \Tile_X0Y5_E2BEG[4] ,
    \Tile_X0Y5_E2BEG[3] ,
    \Tile_X0Y5_E2BEG[2] ,
    \Tile_X0Y5_E2BEG[1] ,
    \Tile_X0Y5_E2BEG[0] }),
    .E2BEGb({\Tile_X0Y5_E2BEGb[7] ,
    \Tile_X0Y5_E2BEGb[6] ,
    \Tile_X0Y5_E2BEGb[5] ,
    \Tile_X0Y5_E2BEGb[4] ,
    \Tile_X0Y5_E2BEGb[3] ,
    \Tile_X0Y5_E2BEGb[2] ,
    \Tile_X0Y5_E2BEGb[1] ,
    \Tile_X0Y5_E2BEGb[0] }),
    .E6BEG({\Tile_X0Y5_E6BEG[11] ,
    \Tile_X0Y5_E6BEG[10] ,
    \Tile_X0Y5_E6BEG[9] ,
    \Tile_X0Y5_E6BEG[8] ,
    \Tile_X0Y5_E6BEG[7] ,
    \Tile_X0Y5_E6BEG[6] ,
    \Tile_X0Y5_E6BEG[5] ,
    \Tile_X0Y5_E6BEG[4] ,
    \Tile_X0Y5_E6BEG[3] ,
    \Tile_X0Y5_E6BEG[2] ,
    \Tile_X0Y5_E6BEG[1] ,
    \Tile_X0Y5_E6BEG[0] }),
    .EE4BEG({\Tile_X0Y5_EE4BEG[15] ,
    \Tile_X0Y5_EE4BEG[14] ,
    \Tile_X0Y5_EE4BEG[13] ,
    \Tile_X0Y5_EE4BEG[12] ,
    \Tile_X0Y5_EE4BEG[11] ,
    \Tile_X0Y5_EE4BEG[10] ,
    \Tile_X0Y5_EE4BEG[9] ,
    \Tile_X0Y5_EE4BEG[8] ,
    \Tile_X0Y5_EE4BEG[7] ,
    \Tile_X0Y5_EE4BEG[6] ,
    \Tile_X0Y5_EE4BEG[5] ,
    \Tile_X0Y5_EE4BEG[4] ,
    \Tile_X0Y5_EE4BEG[3] ,
    \Tile_X0Y5_EE4BEG[2] ,
    \Tile_X0Y5_EE4BEG[1] ,
    \Tile_X0Y5_EE4BEG[0] }),
    .FrameData({FrameData[191],
    FrameData[190],
    FrameData[189],
    FrameData[188],
    FrameData[187],
    FrameData[186],
    FrameData[185],
    FrameData[184],
    FrameData[183],
    FrameData[182],
    FrameData[181],
    FrameData[180],
    FrameData[179],
    FrameData[178],
    FrameData[177],
    FrameData[176],
    FrameData[175],
    FrameData[174],
    FrameData[173],
    FrameData[172],
    FrameData[171],
    FrameData[170],
    FrameData[169],
    FrameData[168],
    FrameData[167],
    FrameData[166],
    FrameData[165],
    FrameData[164],
    FrameData[163],
    FrameData[162],
    FrameData[161],
    FrameData[160]}),
    .FrameData_O({\Tile_X0Y5_FrameData_O[31] ,
    \Tile_X0Y5_FrameData_O[30] ,
    \Tile_X0Y5_FrameData_O[29] ,
    \Tile_X0Y5_FrameData_O[28] ,
    \Tile_X0Y5_FrameData_O[27] ,
    \Tile_X0Y5_FrameData_O[26] ,
    \Tile_X0Y5_FrameData_O[25] ,
    \Tile_X0Y5_FrameData_O[24] ,
    \Tile_X0Y5_FrameData_O[23] ,
    \Tile_X0Y5_FrameData_O[22] ,
    \Tile_X0Y5_FrameData_O[21] ,
    \Tile_X0Y5_FrameData_O[20] ,
    \Tile_X0Y5_FrameData_O[19] ,
    \Tile_X0Y5_FrameData_O[18] ,
    \Tile_X0Y5_FrameData_O[17] ,
    \Tile_X0Y5_FrameData_O[16] ,
    \Tile_X0Y5_FrameData_O[15] ,
    \Tile_X0Y5_FrameData_O[14] ,
    \Tile_X0Y5_FrameData_O[13] ,
    \Tile_X0Y5_FrameData_O[12] ,
    \Tile_X0Y5_FrameData_O[11] ,
    \Tile_X0Y5_FrameData_O[10] ,
    \Tile_X0Y5_FrameData_O[9] ,
    \Tile_X0Y5_FrameData_O[8] ,
    \Tile_X0Y5_FrameData_O[7] ,
    \Tile_X0Y5_FrameData_O[6] ,
    \Tile_X0Y5_FrameData_O[5] ,
    \Tile_X0Y5_FrameData_O[4] ,
    \Tile_X0Y5_FrameData_O[3] ,
    \Tile_X0Y5_FrameData_O[2] ,
    \Tile_X0Y5_FrameData_O[1] ,
    \Tile_X0Y5_FrameData_O[0] }),
    .FrameStrobe({\Tile_X0Y6_FrameStrobe_O[19] ,
    \Tile_X0Y6_FrameStrobe_O[18] ,
    \Tile_X0Y6_FrameStrobe_O[17] ,
    \Tile_X0Y6_FrameStrobe_O[16] ,
    \Tile_X0Y6_FrameStrobe_O[15] ,
    \Tile_X0Y6_FrameStrobe_O[14] ,
    \Tile_X0Y6_FrameStrobe_O[13] ,
    \Tile_X0Y6_FrameStrobe_O[12] ,
    \Tile_X0Y6_FrameStrobe_O[11] ,
    \Tile_X0Y6_FrameStrobe_O[10] ,
    \Tile_X0Y6_FrameStrobe_O[9] ,
    \Tile_X0Y6_FrameStrobe_O[8] ,
    \Tile_X0Y6_FrameStrobe_O[7] ,
    \Tile_X0Y6_FrameStrobe_O[6] ,
    \Tile_X0Y6_FrameStrobe_O[5] ,
    \Tile_X0Y6_FrameStrobe_O[4] ,
    \Tile_X0Y6_FrameStrobe_O[3] ,
    \Tile_X0Y6_FrameStrobe_O[2] ,
    \Tile_X0Y6_FrameStrobe_O[1] ,
    \Tile_X0Y6_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X0Y5_FrameStrobe_O[19] ,
    \Tile_X0Y5_FrameStrobe_O[18] ,
    \Tile_X0Y5_FrameStrobe_O[17] ,
    \Tile_X0Y5_FrameStrobe_O[16] ,
    \Tile_X0Y5_FrameStrobe_O[15] ,
    \Tile_X0Y5_FrameStrobe_O[14] ,
    \Tile_X0Y5_FrameStrobe_O[13] ,
    \Tile_X0Y5_FrameStrobe_O[12] ,
    \Tile_X0Y5_FrameStrobe_O[11] ,
    \Tile_X0Y5_FrameStrobe_O[10] ,
    \Tile_X0Y5_FrameStrobe_O[9] ,
    \Tile_X0Y5_FrameStrobe_O[8] ,
    \Tile_X0Y5_FrameStrobe_O[7] ,
    \Tile_X0Y5_FrameStrobe_O[6] ,
    \Tile_X0Y5_FrameStrobe_O[5] ,
    \Tile_X0Y5_FrameStrobe_O[4] ,
    \Tile_X0Y5_FrameStrobe_O[3] ,
    \Tile_X0Y5_FrameStrobe_O[2] ,
    \Tile_X0Y5_FrameStrobe_O[1] ,
    \Tile_X0Y5_FrameStrobe_O[0] }),
    .W1END({\Tile_X1Y5_W1BEG[3] ,
    \Tile_X1Y5_W1BEG[2] ,
    \Tile_X1Y5_W1BEG[1] ,
    \Tile_X1Y5_W1BEG[0] }),
    .W2END({\Tile_X1Y5_W2BEGb[7] ,
    \Tile_X1Y5_W2BEGb[6] ,
    \Tile_X1Y5_W2BEGb[5] ,
    \Tile_X1Y5_W2BEGb[4] ,
    \Tile_X1Y5_W2BEGb[3] ,
    \Tile_X1Y5_W2BEGb[2] ,
    \Tile_X1Y5_W2BEGb[1] ,
    \Tile_X1Y5_W2BEGb[0] }),
    .W2MID({\Tile_X1Y5_W2BEG[7] ,
    \Tile_X1Y5_W2BEG[6] ,
    \Tile_X1Y5_W2BEG[5] ,
    \Tile_X1Y5_W2BEG[4] ,
    \Tile_X1Y5_W2BEG[3] ,
    \Tile_X1Y5_W2BEG[2] ,
    \Tile_X1Y5_W2BEG[1] ,
    \Tile_X1Y5_W2BEG[0] }),
    .W6END({\Tile_X1Y5_W6BEG[11] ,
    \Tile_X1Y5_W6BEG[10] ,
    \Tile_X1Y5_W6BEG[9] ,
    \Tile_X1Y5_W6BEG[8] ,
    \Tile_X1Y5_W6BEG[7] ,
    \Tile_X1Y5_W6BEG[6] ,
    \Tile_X1Y5_W6BEG[5] ,
    \Tile_X1Y5_W6BEG[4] ,
    \Tile_X1Y5_W6BEG[3] ,
    \Tile_X1Y5_W6BEG[2] ,
    \Tile_X1Y5_W6BEG[1] ,
    \Tile_X1Y5_W6BEG[0] }),
    .WW4END({\Tile_X1Y5_WW4BEG[15] ,
    \Tile_X1Y5_WW4BEG[14] ,
    \Tile_X1Y5_WW4BEG[13] ,
    \Tile_X1Y5_WW4BEG[12] ,
    \Tile_X1Y5_WW4BEG[11] ,
    \Tile_X1Y5_WW4BEG[10] ,
    \Tile_X1Y5_WW4BEG[9] ,
    \Tile_X1Y5_WW4BEG[8] ,
    \Tile_X1Y5_WW4BEG[7] ,
    \Tile_X1Y5_WW4BEG[6] ,
    \Tile_X1Y5_WW4BEG[5] ,
    \Tile_X1Y5_WW4BEG[4] ,
    \Tile_X1Y5_WW4BEG[3] ,
    \Tile_X1Y5_WW4BEG[2] ,
    \Tile_X1Y5_WW4BEG[1] ,
    \Tile_X1Y5_WW4BEG[0] }));
 W_IO Tile_X0Y6_W_IO (.A_I_top(Tile_X0Y6_A_I_top),
    .A_O_top(Tile_X0Y6_A_O_top),
    .A_T_top(Tile_X0Y6_A_T_top),
    .A_config_C_bit0(Tile_X0Y6_A_config_C_bit0),
    .A_config_C_bit1(Tile_X0Y6_A_config_C_bit1),
    .A_config_C_bit2(Tile_X0Y6_A_config_C_bit2),
    .A_config_C_bit3(Tile_X0Y6_A_config_C_bit3),
    .B_I_top(Tile_X0Y6_B_I_top),
    .B_O_top(Tile_X0Y6_B_O_top),
    .B_T_top(Tile_X0Y6_B_T_top),
    .B_config_C_bit0(Tile_X0Y6_B_config_C_bit0),
    .B_config_C_bit1(Tile_X0Y6_B_config_C_bit1),
    .B_config_C_bit2(Tile_X0Y6_B_config_C_bit2),
    .B_config_C_bit3(Tile_X0Y6_B_config_C_bit3),
    .UserCLK(Tile_X0Y7_UserCLKo),
    .UserCLKo(Tile_X0Y6_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X0Y6_E1BEG[3] ,
    \Tile_X0Y6_E1BEG[2] ,
    \Tile_X0Y6_E1BEG[1] ,
    \Tile_X0Y6_E1BEG[0] }),
    .E2BEG({\Tile_X0Y6_E2BEG[7] ,
    \Tile_X0Y6_E2BEG[6] ,
    \Tile_X0Y6_E2BEG[5] ,
    \Tile_X0Y6_E2BEG[4] ,
    \Tile_X0Y6_E2BEG[3] ,
    \Tile_X0Y6_E2BEG[2] ,
    \Tile_X0Y6_E2BEG[1] ,
    \Tile_X0Y6_E2BEG[0] }),
    .E2BEGb({\Tile_X0Y6_E2BEGb[7] ,
    \Tile_X0Y6_E2BEGb[6] ,
    \Tile_X0Y6_E2BEGb[5] ,
    \Tile_X0Y6_E2BEGb[4] ,
    \Tile_X0Y6_E2BEGb[3] ,
    \Tile_X0Y6_E2BEGb[2] ,
    \Tile_X0Y6_E2BEGb[1] ,
    \Tile_X0Y6_E2BEGb[0] }),
    .E6BEG({\Tile_X0Y6_E6BEG[11] ,
    \Tile_X0Y6_E6BEG[10] ,
    \Tile_X0Y6_E6BEG[9] ,
    \Tile_X0Y6_E6BEG[8] ,
    \Tile_X0Y6_E6BEG[7] ,
    \Tile_X0Y6_E6BEG[6] ,
    \Tile_X0Y6_E6BEG[5] ,
    \Tile_X0Y6_E6BEG[4] ,
    \Tile_X0Y6_E6BEG[3] ,
    \Tile_X0Y6_E6BEG[2] ,
    \Tile_X0Y6_E6BEG[1] ,
    \Tile_X0Y6_E6BEG[0] }),
    .EE4BEG({\Tile_X0Y6_EE4BEG[15] ,
    \Tile_X0Y6_EE4BEG[14] ,
    \Tile_X0Y6_EE4BEG[13] ,
    \Tile_X0Y6_EE4BEG[12] ,
    \Tile_X0Y6_EE4BEG[11] ,
    \Tile_X0Y6_EE4BEG[10] ,
    \Tile_X0Y6_EE4BEG[9] ,
    \Tile_X0Y6_EE4BEG[8] ,
    \Tile_X0Y6_EE4BEG[7] ,
    \Tile_X0Y6_EE4BEG[6] ,
    \Tile_X0Y6_EE4BEG[5] ,
    \Tile_X0Y6_EE4BEG[4] ,
    \Tile_X0Y6_EE4BEG[3] ,
    \Tile_X0Y6_EE4BEG[2] ,
    \Tile_X0Y6_EE4BEG[1] ,
    \Tile_X0Y6_EE4BEG[0] }),
    .FrameData({FrameData[223],
    FrameData[222],
    FrameData[221],
    FrameData[220],
    FrameData[219],
    FrameData[218],
    FrameData[217],
    FrameData[216],
    FrameData[215],
    FrameData[214],
    FrameData[213],
    FrameData[212],
    FrameData[211],
    FrameData[210],
    FrameData[209],
    FrameData[208],
    FrameData[207],
    FrameData[206],
    FrameData[205],
    FrameData[204],
    FrameData[203],
    FrameData[202],
    FrameData[201],
    FrameData[200],
    FrameData[199],
    FrameData[198],
    FrameData[197],
    FrameData[196],
    FrameData[195],
    FrameData[194],
    FrameData[193],
    FrameData[192]}),
    .FrameData_O({\Tile_X0Y6_FrameData_O[31] ,
    \Tile_X0Y6_FrameData_O[30] ,
    \Tile_X0Y6_FrameData_O[29] ,
    \Tile_X0Y6_FrameData_O[28] ,
    \Tile_X0Y6_FrameData_O[27] ,
    \Tile_X0Y6_FrameData_O[26] ,
    \Tile_X0Y6_FrameData_O[25] ,
    \Tile_X0Y6_FrameData_O[24] ,
    \Tile_X0Y6_FrameData_O[23] ,
    \Tile_X0Y6_FrameData_O[22] ,
    \Tile_X0Y6_FrameData_O[21] ,
    \Tile_X0Y6_FrameData_O[20] ,
    \Tile_X0Y6_FrameData_O[19] ,
    \Tile_X0Y6_FrameData_O[18] ,
    \Tile_X0Y6_FrameData_O[17] ,
    \Tile_X0Y6_FrameData_O[16] ,
    \Tile_X0Y6_FrameData_O[15] ,
    \Tile_X0Y6_FrameData_O[14] ,
    \Tile_X0Y6_FrameData_O[13] ,
    \Tile_X0Y6_FrameData_O[12] ,
    \Tile_X0Y6_FrameData_O[11] ,
    \Tile_X0Y6_FrameData_O[10] ,
    \Tile_X0Y6_FrameData_O[9] ,
    \Tile_X0Y6_FrameData_O[8] ,
    \Tile_X0Y6_FrameData_O[7] ,
    \Tile_X0Y6_FrameData_O[6] ,
    \Tile_X0Y6_FrameData_O[5] ,
    \Tile_X0Y6_FrameData_O[4] ,
    \Tile_X0Y6_FrameData_O[3] ,
    \Tile_X0Y6_FrameData_O[2] ,
    \Tile_X0Y6_FrameData_O[1] ,
    \Tile_X0Y6_FrameData_O[0] }),
    .FrameStrobe({\Tile_X0Y7_FrameStrobe_O[19] ,
    \Tile_X0Y7_FrameStrobe_O[18] ,
    \Tile_X0Y7_FrameStrobe_O[17] ,
    \Tile_X0Y7_FrameStrobe_O[16] ,
    \Tile_X0Y7_FrameStrobe_O[15] ,
    \Tile_X0Y7_FrameStrobe_O[14] ,
    \Tile_X0Y7_FrameStrobe_O[13] ,
    \Tile_X0Y7_FrameStrobe_O[12] ,
    \Tile_X0Y7_FrameStrobe_O[11] ,
    \Tile_X0Y7_FrameStrobe_O[10] ,
    \Tile_X0Y7_FrameStrobe_O[9] ,
    \Tile_X0Y7_FrameStrobe_O[8] ,
    \Tile_X0Y7_FrameStrobe_O[7] ,
    \Tile_X0Y7_FrameStrobe_O[6] ,
    \Tile_X0Y7_FrameStrobe_O[5] ,
    \Tile_X0Y7_FrameStrobe_O[4] ,
    \Tile_X0Y7_FrameStrobe_O[3] ,
    \Tile_X0Y7_FrameStrobe_O[2] ,
    \Tile_X0Y7_FrameStrobe_O[1] ,
    \Tile_X0Y7_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X0Y6_FrameStrobe_O[19] ,
    \Tile_X0Y6_FrameStrobe_O[18] ,
    \Tile_X0Y6_FrameStrobe_O[17] ,
    \Tile_X0Y6_FrameStrobe_O[16] ,
    \Tile_X0Y6_FrameStrobe_O[15] ,
    \Tile_X0Y6_FrameStrobe_O[14] ,
    \Tile_X0Y6_FrameStrobe_O[13] ,
    \Tile_X0Y6_FrameStrobe_O[12] ,
    \Tile_X0Y6_FrameStrobe_O[11] ,
    \Tile_X0Y6_FrameStrobe_O[10] ,
    \Tile_X0Y6_FrameStrobe_O[9] ,
    \Tile_X0Y6_FrameStrobe_O[8] ,
    \Tile_X0Y6_FrameStrobe_O[7] ,
    \Tile_X0Y6_FrameStrobe_O[6] ,
    \Tile_X0Y6_FrameStrobe_O[5] ,
    \Tile_X0Y6_FrameStrobe_O[4] ,
    \Tile_X0Y6_FrameStrobe_O[3] ,
    \Tile_X0Y6_FrameStrobe_O[2] ,
    \Tile_X0Y6_FrameStrobe_O[1] ,
    \Tile_X0Y6_FrameStrobe_O[0] }),
    .W1END({\Tile_X1Y6_W1BEG[3] ,
    \Tile_X1Y6_W1BEG[2] ,
    \Tile_X1Y6_W1BEG[1] ,
    \Tile_X1Y6_W1BEG[0] }),
    .W2END({\Tile_X1Y6_W2BEGb[7] ,
    \Tile_X1Y6_W2BEGb[6] ,
    \Tile_X1Y6_W2BEGb[5] ,
    \Tile_X1Y6_W2BEGb[4] ,
    \Tile_X1Y6_W2BEGb[3] ,
    \Tile_X1Y6_W2BEGb[2] ,
    \Tile_X1Y6_W2BEGb[1] ,
    \Tile_X1Y6_W2BEGb[0] }),
    .W2MID({\Tile_X1Y6_W2BEG[7] ,
    \Tile_X1Y6_W2BEG[6] ,
    \Tile_X1Y6_W2BEG[5] ,
    \Tile_X1Y6_W2BEG[4] ,
    \Tile_X1Y6_W2BEG[3] ,
    \Tile_X1Y6_W2BEG[2] ,
    \Tile_X1Y6_W2BEG[1] ,
    \Tile_X1Y6_W2BEG[0] }),
    .W6END({\Tile_X1Y6_W6BEG[11] ,
    \Tile_X1Y6_W6BEG[10] ,
    \Tile_X1Y6_W6BEG[9] ,
    \Tile_X1Y6_W6BEG[8] ,
    \Tile_X1Y6_W6BEG[7] ,
    \Tile_X1Y6_W6BEG[6] ,
    \Tile_X1Y6_W6BEG[5] ,
    \Tile_X1Y6_W6BEG[4] ,
    \Tile_X1Y6_W6BEG[3] ,
    \Tile_X1Y6_W6BEG[2] ,
    \Tile_X1Y6_W6BEG[1] ,
    \Tile_X1Y6_W6BEG[0] }),
    .WW4END({\Tile_X1Y6_WW4BEG[15] ,
    \Tile_X1Y6_WW4BEG[14] ,
    \Tile_X1Y6_WW4BEG[13] ,
    \Tile_X1Y6_WW4BEG[12] ,
    \Tile_X1Y6_WW4BEG[11] ,
    \Tile_X1Y6_WW4BEG[10] ,
    \Tile_X1Y6_WW4BEG[9] ,
    \Tile_X1Y6_WW4BEG[8] ,
    \Tile_X1Y6_WW4BEG[7] ,
    \Tile_X1Y6_WW4BEG[6] ,
    \Tile_X1Y6_WW4BEG[5] ,
    \Tile_X1Y6_WW4BEG[4] ,
    \Tile_X1Y6_WW4BEG[3] ,
    \Tile_X1Y6_WW4BEG[2] ,
    \Tile_X1Y6_WW4BEG[1] ,
    \Tile_X1Y6_WW4BEG[0] }));
 W_IO Tile_X0Y7_W_IO (.A_I_top(Tile_X0Y7_A_I_top),
    .A_O_top(Tile_X0Y7_A_O_top),
    .A_T_top(Tile_X0Y7_A_T_top),
    .A_config_C_bit0(Tile_X0Y7_A_config_C_bit0),
    .A_config_C_bit1(Tile_X0Y7_A_config_C_bit1),
    .A_config_C_bit2(Tile_X0Y7_A_config_C_bit2),
    .A_config_C_bit3(Tile_X0Y7_A_config_C_bit3),
    .B_I_top(Tile_X0Y7_B_I_top),
    .B_O_top(Tile_X0Y7_B_O_top),
    .B_T_top(Tile_X0Y7_B_T_top),
    .B_config_C_bit0(Tile_X0Y7_B_config_C_bit0),
    .B_config_C_bit1(Tile_X0Y7_B_config_C_bit1),
    .B_config_C_bit2(Tile_X0Y7_B_config_C_bit2),
    .B_config_C_bit3(Tile_X0Y7_B_config_C_bit3),
    .UserCLK(Tile_X0Y8_UserCLKo),
    .UserCLKo(Tile_X0Y7_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X0Y7_E1BEG[3] ,
    \Tile_X0Y7_E1BEG[2] ,
    \Tile_X0Y7_E1BEG[1] ,
    \Tile_X0Y7_E1BEG[0] }),
    .E2BEG({\Tile_X0Y7_E2BEG[7] ,
    \Tile_X0Y7_E2BEG[6] ,
    \Tile_X0Y7_E2BEG[5] ,
    \Tile_X0Y7_E2BEG[4] ,
    \Tile_X0Y7_E2BEG[3] ,
    \Tile_X0Y7_E2BEG[2] ,
    \Tile_X0Y7_E2BEG[1] ,
    \Tile_X0Y7_E2BEG[0] }),
    .E2BEGb({\Tile_X0Y7_E2BEGb[7] ,
    \Tile_X0Y7_E2BEGb[6] ,
    \Tile_X0Y7_E2BEGb[5] ,
    \Tile_X0Y7_E2BEGb[4] ,
    \Tile_X0Y7_E2BEGb[3] ,
    \Tile_X0Y7_E2BEGb[2] ,
    \Tile_X0Y7_E2BEGb[1] ,
    \Tile_X0Y7_E2BEGb[0] }),
    .E6BEG({\Tile_X0Y7_E6BEG[11] ,
    \Tile_X0Y7_E6BEG[10] ,
    \Tile_X0Y7_E6BEG[9] ,
    \Tile_X0Y7_E6BEG[8] ,
    \Tile_X0Y7_E6BEG[7] ,
    \Tile_X0Y7_E6BEG[6] ,
    \Tile_X0Y7_E6BEG[5] ,
    \Tile_X0Y7_E6BEG[4] ,
    \Tile_X0Y7_E6BEG[3] ,
    \Tile_X0Y7_E6BEG[2] ,
    \Tile_X0Y7_E6BEG[1] ,
    \Tile_X0Y7_E6BEG[0] }),
    .EE4BEG({\Tile_X0Y7_EE4BEG[15] ,
    \Tile_X0Y7_EE4BEG[14] ,
    \Tile_X0Y7_EE4BEG[13] ,
    \Tile_X0Y7_EE4BEG[12] ,
    \Tile_X0Y7_EE4BEG[11] ,
    \Tile_X0Y7_EE4BEG[10] ,
    \Tile_X0Y7_EE4BEG[9] ,
    \Tile_X0Y7_EE4BEG[8] ,
    \Tile_X0Y7_EE4BEG[7] ,
    \Tile_X0Y7_EE4BEG[6] ,
    \Tile_X0Y7_EE4BEG[5] ,
    \Tile_X0Y7_EE4BEG[4] ,
    \Tile_X0Y7_EE4BEG[3] ,
    \Tile_X0Y7_EE4BEG[2] ,
    \Tile_X0Y7_EE4BEG[1] ,
    \Tile_X0Y7_EE4BEG[0] }),
    .FrameData({FrameData[255],
    FrameData[254],
    FrameData[253],
    FrameData[252],
    FrameData[251],
    FrameData[250],
    FrameData[249],
    FrameData[248],
    FrameData[247],
    FrameData[246],
    FrameData[245],
    FrameData[244],
    FrameData[243],
    FrameData[242],
    FrameData[241],
    FrameData[240],
    FrameData[239],
    FrameData[238],
    FrameData[237],
    FrameData[236],
    FrameData[235],
    FrameData[234],
    FrameData[233],
    FrameData[232],
    FrameData[231],
    FrameData[230],
    FrameData[229],
    FrameData[228],
    FrameData[227],
    FrameData[226],
    FrameData[225],
    FrameData[224]}),
    .FrameData_O({\Tile_X0Y7_FrameData_O[31] ,
    \Tile_X0Y7_FrameData_O[30] ,
    \Tile_X0Y7_FrameData_O[29] ,
    \Tile_X0Y7_FrameData_O[28] ,
    \Tile_X0Y7_FrameData_O[27] ,
    \Tile_X0Y7_FrameData_O[26] ,
    \Tile_X0Y7_FrameData_O[25] ,
    \Tile_X0Y7_FrameData_O[24] ,
    \Tile_X0Y7_FrameData_O[23] ,
    \Tile_X0Y7_FrameData_O[22] ,
    \Tile_X0Y7_FrameData_O[21] ,
    \Tile_X0Y7_FrameData_O[20] ,
    \Tile_X0Y7_FrameData_O[19] ,
    \Tile_X0Y7_FrameData_O[18] ,
    \Tile_X0Y7_FrameData_O[17] ,
    \Tile_X0Y7_FrameData_O[16] ,
    \Tile_X0Y7_FrameData_O[15] ,
    \Tile_X0Y7_FrameData_O[14] ,
    \Tile_X0Y7_FrameData_O[13] ,
    \Tile_X0Y7_FrameData_O[12] ,
    \Tile_X0Y7_FrameData_O[11] ,
    \Tile_X0Y7_FrameData_O[10] ,
    \Tile_X0Y7_FrameData_O[9] ,
    \Tile_X0Y7_FrameData_O[8] ,
    \Tile_X0Y7_FrameData_O[7] ,
    \Tile_X0Y7_FrameData_O[6] ,
    \Tile_X0Y7_FrameData_O[5] ,
    \Tile_X0Y7_FrameData_O[4] ,
    \Tile_X0Y7_FrameData_O[3] ,
    \Tile_X0Y7_FrameData_O[2] ,
    \Tile_X0Y7_FrameData_O[1] ,
    \Tile_X0Y7_FrameData_O[0] }),
    .FrameStrobe({\Tile_X0Y8_FrameStrobe_O[19] ,
    \Tile_X0Y8_FrameStrobe_O[18] ,
    \Tile_X0Y8_FrameStrobe_O[17] ,
    \Tile_X0Y8_FrameStrobe_O[16] ,
    \Tile_X0Y8_FrameStrobe_O[15] ,
    \Tile_X0Y8_FrameStrobe_O[14] ,
    \Tile_X0Y8_FrameStrobe_O[13] ,
    \Tile_X0Y8_FrameStrobe_O[12] ,
    \Tile_X0Y8_FrameStrobe_O[11] ,
    \Tile_X0Y8_FrameStrobe_O[10] ,
    \Tile_X0Y8_FrameStrobe_O[9] ,
    \Tile_X0Y8_FrameStrobe_O[8] ,
    \Tile_X0Y8_FrameStrobe_O[7] ,
    \Tile_X0Y8_FrameStrobe_O[6] ,
    \Tile_X0Y8_FrameStrobe_O[5] ,
    \Tile_X0Y8_FrameStrobe_O[4] ,
    \Tile_X0Y8_FrameStrobe_O[3] ,
    \Tile_X0Y8_FrameStrobe_O[2] ,
    \Tile_X0Y8_FrameStrobe_O[1] ,
    \Tile_X0Y8_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X0Y7_FrameStrobe_O[19] ,
    \Tile_X0Y7_FrameStrobe_O[18] ,
    \Tile_X0Y7_FrameStrobe_O[17] ,
    \Tile_X0Y7_FrameStrobe_O[16] ,
    \Tile_X0Y7_FrameStrobe_O[15] ,
    \Tile_X0Y7_FrameStrobe_O[14] ,
    \Tile_X0Y7_FrameStrobe_O[13] ,
    \Tile_X0Y7_FrameStrobe_O[12] ,
    \Tile_X0Y7_FrameStrobe_O[11] ,
    \Tile_X0Y7_FrameStrobe_O[10] ,
    \Tile_X0Y7_FrameStrobe_O[9] ,
    \Tile_X0Y7_FrameStrobe_O[8] ,
    \Tile_X0Y7_FrameStrobe_O[7] ,
    \Tile_X0Y7_FrameStrobe_O[6] ,
    \Tile_X0Y7_FrameStrobe_O[5] ,
    \Tile_X0Y7_FrameStrobe_O[4] ,
    \Tile_X0Y7_FrameStrobe_O[3] ,
    \Tile_X0Y7_FrameStrobe_O[2] ,
    \Tile_X0Y7_FrameStrobe_O[1] ,
    \Tile_X0Y7_FrameStrobe_O[0] }),
    .W1END({\Tile_X1Y7_W1BEG[3] ,
    \Tile_X1Y7_W1BEG[2] ,
    \Tile_X1Y7_W1BEG[1] ,
    \Tile_X1Y7_W1BEG[0] }),
    .W2END({\Tile_X1Y7_W2BEGb[7] ,
    \Tile_X1Y7_W2BEGb[6] ,
    \Tile_X1Y7_W2BEGb[5] ,
    \Tile_X1Y7_W2BEGb[4] ,
    \Tile_X1Y7_W2BEGb[3] ,
    \Tile_X1Y7_W2BEGb[2] ,
    \Tile_X1Y7_W2BEGb[1] ,
    \Tile_X1Y7_W2BEGb[0] }),
    .W2MID({\Tile_X1Y7_W2BEG[7] ,
    \Tile_X1Y7_W2BEG[6] ,
    \Tile_X1Y7_W2BEG[5] ,
    \Tile_X1Y7_W2BEG[4] ,
    \Tile_X1Y7_W2BEG[3] ,
    \Tile_X1Y7_W2BEG[2] ,
    \Tile_X1Y7_W2BEG[1] ,
    \Tile_X1Y7_W2BEG[0] }),
    .W6END({\Tile_X1Y7_W6BEG[11] ,
    \Tile_X1Y7_W6BEG[10] ,
    \Tile_X1Y7_W6BEG[9] ,
    \Tile_X1Y7_W6BEG[8] ,
    \Tile_X1Y7_W6BEG[7] ,
    \Tile_X1Y7_W6BEG[6] ,
    \Tile_X1Y7_W6BEG[5] ,
    \Tile_X1Y7_W6BEG[4] ,
    \Tile_X1Y7_W6BEG[3] ,
    \Tile_X1Y7_W6BEG[2] ,
    \Tile_X1Y7_W6BEG[1] ,
    \Tile_X1Y7_W6BEG[0] }),
    .WW4END({\Tile_X1Y7_WW4BEG[15] ,
    \Tile_X1Y7_WW4BEG[14] ,
    \Tile_X1Y7_WW4BEG[13] ,
    \Tile_X1Y7_WW4BEG[12] ,
    \Tile_X1Y7_WW4BEG[11] ,
    \Tile_X1Y7_WW4BEG[10] ,
    \Tile_X1Y7_WW4BEG[9] ,
    \Tile_X1Y7_WW4BEG[8] ,
    \Tile_X1Y7_WW4BEG[7] ,
    \Tile_X1Y7_WW4BEG[6] ,
    \Tile_X1Y7_WW4BEG[5] ,
    \Tile_X1Y7_WW4BEG[4] ,
    \Tile_X1Y7_WW4BEG[3] ,
    \Tile_X1Y7_WW4BEG[2] ,
    \Tile_X1Y7_WW4BEG[1] ,
    \Tile_X1Y7_WW4BEG[0] }));
 W_IO Tile_X0Y8_W_IO (.A_I_top(Tile_X0Y8_A_I_top),
    .A_O_top(Tile_X0Y8_A_O_top),
    .A_T_top(Tile_X0Y8_A_T_top),
    .A_config_C_bit0(Tile_X0Y8_A_config_C_bit0),
    .A_config_C_bit1(Tile_X0Y8_A_config_C_bit1),
    .A_config_C_bit2(Tile_X0Y8_A_config_C_bit2),
    .A_config_C_bit3(Tile_X0Y8_A_config_C_bit3),
    .B_I_top(Tile_X0Y8_B_I_top),
    .B_O_top(Tile_X0Y8_B_O_top),
    .B_T_top(Tile_X0Y8_B_T_top),
    .B_config_C_bit0(Tile_X0Y8_B_config_C_bit0),
    .B_config_C_bit1(Tile_X0Y8_B_config_C_bit1),
    .B_config_C_bit2(Tile_X0Y8_B_config_C_bit2),
    .B_config_C_bit3(Tile_X0Y8_B_config_C_bit3),
    .UserCLK(Tile_X0Y9_UserCLKo),
    .UserCLKo(Tile_X0Y8_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X0Y8_E1BEG[3] ,
    \Tile_X0Y8_E1BEG[2] ,
    \Tile_X0Y8_E1BEG[1] ,
    \Tile_X0Y8_E1BEG[0] }),
    .E2BEG({\Tile_X0Y8_E2BEG[7] ,
    \Tile_X0Y8_E2BEG[6] ,
    \Tile_X0Y8_E2BEG[5] ,
    \Tile_X0Y8_E2BEG[4] ,
    \Tile_X0Y8_E2BEG[3] ,
    \Tile_X0Y8_E2BEG[2] ,
    \Tile_X0Y8_E2BEG[1] ,
    \Tile_X0Y8_E2BEG[0] }),
    .E2BEGb({\Tile_X0Y8_E2BEGb[7] ,
    \Tile_X0Y8_E2BEGb[6] ,
    \Tile_X0Y8_E2BEGb[5] ,
    \Tile_X0Y8_E2BEGb[4] ,
    \Tile_X0Y8_E2BEGb[3] ,
    \Tile_X0Y8_E2BEGb[2] ,
    \Tile_X0Y8_E2BEGb[1] ,
    \Tile_X0Y8_E2BEGb[0] }),
    .E6BEG({\Tile_X0Y8_E6BEG[11] ,
    \Tile_X0Y8_E6BEG[10] ,
    \Tile_X0Y8_E6BEG[9] ,
    \Tile_X0Y8_E6BEG[8] ,
    \Tile_X0Y8_E6BEG[7] ,
    \Tile_X0Y8_E6BEG[6] ,
    \Tile_X0Y8_E6BEG[5] ,
    \Tile_X0Y8_E6BEG[4] ,
    \Tile_X0Y8_E6BEG[3] ,
    \Tile_X0Y8_E6BEG[2] ,
    \Tile_X0Y8_E6BEG[1] ,
    \Tile_X0Y8_E6BEG[0] }),
    .EE4BEG({\Tile_X0Y8_EE4BEG[15] ,
    \Tile_X0Y8_EE4BEG[14] ,
    \Tile_X0Y8_EE4BEG[13] ,
    \Tile_X0Y8_EE4BEG[12] ,
    \Tile_X0Y8_EE4BEG[11] ,
    \Tile_X0Y8_EE4BEG[10] ,
    \Tile_X0Y8_EE4BEG[9] ,
    \Tile_X0Y8_EE4BEG[8] ,
    \Tile_X0Y8_EE4BEG[7] ,
    \Tile_X0Y8_EE4BEG[6] ,
    \Tile_X0Y8_EE4BEG[5] ,
    \Tile_X0Y8_EE4BEG[4] ,
    \Tile_X0Y8_EE4BEG[3] ,
    \Tile_X0Y8_EE4BEG[2] ,
    \Tile_X0Y8_EE4BEG[1] ,
    \Tile_X0Y8_EE4BEG[0] }),
    .FrameData({FrameData[287],
    FrameData[286],
    FrameData[285],
    FrameData[284],
    FrameData[283],
    FrameData[282],
    FrameData[281],
    FrameData[280],
    FrameData[279],
    FrameData[278],
    FrameData[277],
    FrameData[276],
    FrameData[275],
    FrameData[274],
    FrameData[273],
    FrameData[272],
    FrameData[271],
    FrameData[270],
    FrameData[269],
    FrameData[268],
    FrameData[267],
    FrameData[266],
    FrameData[265],
    FrameData[264],
    FrameData[263],
    FrameData[262],
    FrameData[261],
    FrameData[260],
    FrameData[259],
    FrameData[258],
    FrameData[257],
    FrameData[256]}),
    .FrameData_O({\Tile_X0Y8_FrameData_O[31] ,
    \Tile_X0Y8_FrameData_O[30] ,
    \Tile_X0Y8_FrameData_O[29] ,
    \Tile_X0Y8_FrameData_O[28] ,
    \Tile_X0Y8_FrameData_O[27] ,
    \Tile_X0Y8_FrameData_O[26] ,
    \Tile_X0Y8_FrameData_O[25] ,
    \Tile_X0Y8_FrameData_O[24] ,
    \Tile_X0Y8_FrameData_O[23] ,
    \Tile_X0Y8_FrameData_O[22] ,
    \Tile_X0Y8_FrameData_O[21] ,
    \Tile_X0Y8_FrameData_O[20] ,
    \Tile_X0Y8_FrameData_O[19] ,
    \Tile_X0Y8_FrameData_O[18] ,
    \Tile_X0Y8_FrameData_O[17] ,
    \Tile_X0Y8_FrameData_O[16] ,
    \Tile_X0Y8_FrameData_O[15] ,
    \Tile_X0Y8_FrameData_O[14] ,
    \Tile_X0Y8_FrameData_O[13] ,
    \Tile_X0Y8_FrameData_O[12] ,
    \Tile_X0Y8_FrameData_O[11] ,
    \Tile_X0Y8_FrameData_O[10] ,
    \Tile_X0Y8_FrameData_O[9] ,
    \Tile_X0Y8_FrameData_O[8] ,
    \Tile_X0Y8_FrameData_O[7] ,
    \Tile_X0Y8_FrameData_O[6] ,
    \Tile_X0Y8_FrameData_O[5] ,
    \Tile_X0Y8_FrameData_O[4] ,
    \Tile_X0Y8_FrameData_O[3] ,
    \Tile_X0Y8_FrameData_O[2] ,
    \Tile_X0Y8_FrameData_O[1] ,
    \Tile_X0Y8_FrameData_O[0] }),
    .FrameStrobe({\Tile_X0Y9_FrameStrobe_O[19] ,
    \Tile_X0Y9_FrameStrobe_O[18] ,
    \Tile_X0Y9_FrameStrobe_O[17] ,
    \Tile_X0Y9_FrameStrobe_O[16] ,
    \Tile_X0Y9_FrameStrobe_O[15] ,
    \Tile_X0Y9_FrameStrobe_O[14] ,
    \Tile_X0Y9_FrameStrobe_O[13] ,
    \Tile_X0Y9_FrameStrobe_O[12] ,
    \Tile_X0Y9_FrameStrobe_O[11] ,
    \Tile_X0Y9_FrameStrobe_O[10] ,
    \Tile_X0Y9_FrameStrobe_O[9] ,
    \Tile_X0Y9_FrameStrobe_O[8] ,
    \Tile_X0Y9_FrameStrobe_O[7] ,
    \Tile_X0Y9_FrameStrobe_O[6] ,
    \Tile_X0Y9_FrameStrobe_O[5] ,
    \Tile_X0Y9_FrameStrobe_O[4] ,
    \Tile_X0Y9_FrameStrobe_O[3] ,
    \Tile_X0Y9_FrameStrobe_O[2] ,
    \Tile_X0Y9_FrameStrobe_O[1] ,
    \Tile_X0Y9_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X0Y8_FrameStrobe_O[19] ,
    \Tile_X0Y8_FrameStrobe_O[18] ,
    \Tile_X0Y8_FrameStrobe_O[17] ,
    \Tile_X0Y8_FrameStrobe_O[16] ,
    \Tile_X0Y8_FrameStrobe_O[15] ,
    \Tile_X0Y8_FrameStrobe_O[14] ,
    \Tile_X0Y8_FrameStrobe_O[13] ,
    \Tile_X0Y8_FrameStrobe_O[12] ,
    \Tile_X0Y8_FrameStrobe_O[11] ,
    \Tile_X0Y8_FrameStrobe_O[10] ,
    \Tile_X0Y8_FrameStrobe_O[9] ,
    \Tile_X0Y8_FrameStrobe_O[8] ,
    \Tile_X0Y8_FrameStrobe_O[7] ,
    \Tile_X0Y8_FrameStrobe_O[6] ,
    \Tile_X0Y8_FrameStrobe_O[5] ,
    \Tile_X0Y8_FrameStrobe_O[4] ,
    \Tile_X0Y8_FrameStrobe_O[3] ,
    \Tile_X0Y8_FrameStrobe_O[2] ,
    \Tile_X0Y8_FrameStrobe_O[1] ,
    \Tile_X0Y8_FrameStrobe_O[0] }),
    .W1END({\Tile_X1Y8_W1BEG[3] ,
    \Tile_X1Y8_W1BEG[2] ,
    \Tile_X1Y8_W1BEG[1] ,
    \Tile_X1Y8_W1BEG[0] }),
    .W2END({\Tile_X1Y8_W2BEGb[7] ,
    \Tile_X1Y8_W2BEGb[6] ,
    \Tile_X1Y8_W2BEGb[5] ,
    \Tile_X1Y8_W2BEGb[4] ,
    \Tile_X1Y8_W2BEGb[3] ,
    \Tile_X1Y8_W2BEGb[2] ,
    \Tile_X1Y8_W2BEGb[1] ,
    \Tile_X1Y8_W2BEGb[0] }),
    .W2MID({\Tile_X1Y8_W2BEG[7] ,
    \Tile_X1Y8_W2BEG[6] ,
    \Tile_X1Y8_W2BEG[5] ,
    \Tile_X1Y8_W2BEG[4] ,
    \Tile_X1Y8_W2BEG[3] ,
    \Tile_X1Y8_W2BEG[2] ,
    \Tile_X1Y8_W2BEG[1] ,
    \Tile_X1Y8_W2BEG[0] }),
    .W6END({\Tile_X1Y8_W6BEG[11] ,
    \Tile_X1Y8_W6BEG[10] ,
    \Tile_X1Y8_W6BEG[9] ,
    \Tile_X1Y8_W6BEG[8] ,
    \Tile_X1Y8_W6BEG[7] ,
    \Tile_X1Y8_W6BEG[6] ,
    \Tile_X1Y8_W6BEG[5] ,
    \Tile_X1Y8_W6BEG[4] ,
    \Tile_X1Y8_W6BEG[3] ,
    \Tile_X1Y8_W6BEG[2] ,
    \Tile_X1Y8_W6BEG[1] ,
    \Tile_X1Y8_W6BEG[0] }),
    .WW4END({\Tile_X1Y8_WW4BEG[15] ,
    \Tile_X1Y8_WW4BEG[14] ,
    \Tile_X1Y8_WW4BEG[13] ,
    \Tile_X1Y8_WW4BEG[12] ,
    \Tile_X1Y8_WW4BEG[11] ,
    \Tile_X1Y8_WW4BEG[10] ,
    \Tile_X1Y8_WW4BEG[9] ,
    \Tile_X1Y8_WW4BEG[8] ,
    \Tile_X1Y8_WW4BEG[7] ,
    \Tile_X1Y8_WW4BEG[6] ,
    \Tile_X1Y8_WW4BEG[5] ,
    \Tile_X1Y8_WW4BEG[4] ,
    \Tile_X1Y8_WW4BEG[3] ,
    \Tile_X1Y8_WW4BEG[2] ,
    \Tile_X1Y8_WW4BEG[1] ,
    \Tile_X1Y8_WW4BEG[0] }));
 W_IO Tile_X0Y9_W_IO (.A_I_top(Tile_X0Y9_A_I_top),
    .A_O_top(Tile_X0Y9_A_O_top),
    .A_T_top(Tile_X0Y9_A_T_top),
    .A_config_C_bit0(Tile_X0Y9_A_config_C_bit0),
    .A_config_C_bit1(Tile_X0Y9_A_config_C_bit1),
    .A_config_C_bit2(Tile_X0Y9_A_config_C_bit2),
    .A_config_C_bit3(Tile_X0Y9_A_config_C_bit3),
    .B_I_top(Tile_X0Y9_B_I_top),
    .B_O_top(Tile_X0Y9_B_O_top),
    .B_T_top(Tile_X0Y9_B_T_top),
    .B_config_C_bit0(Tile_X0Y9_B_config_C_bit0),
    .B_config_C_bit1(Tile_X0Y9_B_config_C_bit1),
    .B_config_C_bit2(Tile_X0Y9_B_config_C_bit2),
    .B_config_C_bit3(Tile_X0Y9_B_config_C_bit3),
    .UserCLK(Tile_X0Y10_UserCLKo),
    .UserCLKo(Tile_X0Y9_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X0Y9_E1BEG[3] ,
    \Tile_X0Y9_E1BEG[2] ,
    \Tile_X0Y9_E1BEG[1] ,
    \Tile_X0Y9_E1BEG[0] }),
    .E2BEG({\Tile_X0Y9_E2BEG[7] ,
    \Tile_X0Y9_E2BEG[6] ,
    \Tile_X0Y9_E2BEG[5] ,
    \Tile_X0Y9_E2BEG[4] ,
    \Tile_X0Y9_E2BEG[3] ,
    \Tile_X0Y9_E2BEG[2] ,
    \Tile_X0Y9_E2BEG[1] ,
    \Tile_X0Y9_E2BEG[0] }),
    .E2BEGb({\Tile_X0Y9_E2BEGb[7] ,
    \Tile_X0Y9_E2BEGb[6] ,
    \Tile_X0Y9_E2BEGb[5] ,
    \Tile_X0Y9_E2BEGb[4] ,
    \Tile_X0Y9_E2BEGb[3] ,
    \Tile_X0Y9_E2BEGb[2] ,
    \Tile_X0Y9_E2BEGb[1] ,
    \Tile_X0Y9_E2BEGb[0] }),
    .E6BEG({\Tile_X0Y9_E6BEG[11] ,
    \Tile_X0Y9_E6BEG[10] ,
    \Tile_X0Y9_E6BEG[9] ,
    \Tile_X0Y9_E6BEG[8] ,
    \Tile_X0Y9_E6BEG[7] ,
    \Tile_X0Y9_E6BEG[6] ,
    \Tile_X0Y9_E6BEG[5] ,
    \Tile_X0Y9_E6BEG[4] ,
    \Tile_X0Y9_E6BEG[3] ,
    \Tile_X0Y9_E6BEG[2] ,
    \Tile_X0Y9_E6BEG[1] ,
    \Tile_X0Y9_E6BEG[0] }),
    .EE4BEG({\Tile_X0Y9_EE4BEG[15] ,
    \Tile_X0Y9_EE4BEG[14] ,
    \Tile_X0Y9_EE4BEG[13] ,
    \Tile_X0Y9_EE4BEG[12] ,
    \Tile_X0Y9_EE4BEG[11] ,
    \Tile_X0Y9_EE4BEG[10] ,
    \Tile_X0Y9_EE4BEG[9] ,
    \Tile_X0Y9_EE4BEG[8] ,
    \Tile_X0Y9_EE4BEG[7] ,
    \Tile_X0Y9_EE4BEG[6] ,
    \Tile_X0Y9_EE4BEG[5] ,
    \Tile_X0Y9_EE4BEG[4] ,
    \Tile_X0Y9_EE4BEG[3] ,
    \Tile_X0Y9_EE4BEG[2] ,
    \Tile_X0Y9_EE4BEG[1] ,
    \Tile_X0Y9_EE4BEG[0] }),
    .FrameData({FrameData[319],
    FrameData[318],
    FrameData[317],
    FrameData[316],
    FrameData[315],
    FrameData[314],
    FrameData[313],
    FrameData[312],
    FrameData[311],
    FrameData[310],
    FrameData[309],
    FrameData[308],
    FrameData[307],
    FrameData[306],
    FrameData[305],
    FrameData[304],
    FrameData[303],
    FrameData[302],
    FrameData[301],
    FrameData[300],
    FrameData[299],
    FrameData[298],
    FrameData[297],
    FrameData[296],
    FrameData[295],
    FrameData[294],
    FrameData[293],
    FrameData[292],
    FrameData[291],
    FrameData[290],
    FrameData[289],
    FrameData[288]}),
    .FrameData_O({\Tile_X0Y9_FrameData_O[31] ,
    \Tile_X0Y9_FrameData_O[30] ,
    \Tile_X0Y9_FrameData_O[29] ,
    \Tile_X0Y9_FrameData_O[28] ,
    \Tile_X0Y9_FrameData_O[27] ,
    \Tile_X0Y9_FrameData_O[26] ,
    \Tile_X0Y9_FrameData_O[25] ,
    \Tile_X0Y9_FrameData_O[24] ,
    \Tile_X0Y9_FrameData_O[23] ,
    \Tile_X0Y9_FrameData_O[22] ,
    \Tile_X0Y9_FrameData_O[21] ,
    \Tile_X0Y9_FrameData_O[20] ,
    \Tile_X0Y9_FrameData_O[19] ,
    \Tile_X0Y9_FrameData_O[18] ,
    \Tile_X0Y9_FrameData_O[17] ,
    \Tile_X0Y9_FrameData_O[16] ,
    \Tile_X0Y9_FrameData_O[15] ,
    \Tile_X0Y9_FrameData_O[14] ,
    \Tile_X0Y9_FrameData_O[13] ,
    \Tile_X0Y9_FrameData_O[12] ,
    \Tile_X0Y9_FrameData_O[11] ,
    \Tile_X0Y9_FrameData_O[10] ,
    \Tile_X0Y9_FrameData_O[9] ,
    \Tile_X0Y9_FrameData_O[8] ,
    \Tile_X0Y9_FrameData_O[7] ,
    \Tile_X0Y9_FrameData_O[6] ,
    \Tile_X0Y9_FrameData_O[5] ,
    \Tile_X0Y9_FrameData_O[4] ,
    \Tile_X0Y9_FrameData_O[3] ,
    \Tile_X0Y9_FrameData_O[2] ,
    \Tile_X0Y9_FrameData_O[1] ,
    \Tile_X0Y9_FrameData_O[0] }),
    .FrameStrobe({\Tile_X0Y10_FrameStrobe_O[19] ,
    \Tile_X0Y10_FrameStrobe_O[18] ,
    \Tile_X0Y10_FrameStrobe_O[17] ,
    \Tile_X0Y10_FrameStrobe_O[16] ,
    \Tile_X0Y10_FrameStrobe_O[15] ,
    \Tile_X0Y10_FrameStrobe_O[14] ,
    \Tile_X0Y10_FrameStrobe_O[13] ,
    \Tile_X0Y10_FrameStrobe_O[12] ,
    \Tile_X0Y10_FrameStrobe_O[11] ,
    \Tile_X0Y10_FrameStrobe_O[10] ,
    \Tile_X0Y10_FrameStrobe_O[9] ,
    \Tile_X0Y10_FrameStrobe_O[8] ,
    \Tile_X0Y10_FrameStrobe_O[7] ,
    \Tile_X0Y10_FrameStrobe_O[6] ,
    \Tile_X0Y10_FrameStrobe_O[5] ,
    \Tile_X0Y10_FrameStrobe_O[4] ,
    \Tile_X0Y10_FrameStrobe_O[3] ,
    \Tile_X0Y10_FrameStrobe_O[2] ,
    \Tile_X0Y10_FrameStrobe_O[1] ,
    \Tile_X0Y10_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X0Y9_FrameStrobe_O[19] ,
    \Tile_X0Y9_FrameStrobe_O[18] ,
    \Tile_X0Y9_FrameStrobe_O[17] ,
    \Tile_X0Y9_FrameStrobe_O[16] ,
    \Tile_X0Y9_FrameStrobe_O[15] ,
    \Tile_X0Y9_FrameStrobe_O[14] ,
    \Tile_X0Y9_FrameStrobe_O[13] ,
    \Tile_X0Y9_FrameStrobe_O[12] ,
    \Tile_X0Y9_FrameStrobe_O[11] ,
    \Tile_X0Y9_FrameStrobe_O[10] ,
    \Tile_X0Y9_FrameStrobe_O[9] ,
    \Tile_X0Y9_FrameStrobe_O[8] ,
    \Tile_X0Y9_FrameStrobe_O[7] ,
    \Tile_X0Y9_FrameStrobe_O[6] ,
    \Tile_X0Y9_FrameStrobe_O[5] ,
    \Tile_X0Y9_FrameStrobe_O[4] ,
    \Tile_X0Y9_FrameStrobe_O[3] ,
    \Tile_X0Y9_FrameStrobe_O[2] ,
    \Tile_X0Y9_FrameStrobe_O[1] ,
    \Tile_X0Y9_FrameStrobe_O[0] }),
    .W1END({\Tile_X1Y9_W1BEG[3] ,
    \Tile_X1Y9_W1BEG[2] ,
    \Tile_X1Y9_W1BEG[1] ,
    \Tile_X1Y9_W1BEG[0] }),
    .W2END({\Tile_X1Y9_W2BEGb[7] ,
    \Tile_X1Y9_W2BEGb[6] ,
    \Tile_X1Y9_W2BEGb[5] ,
    \Tile_X1Y9_W2BEGb[4] ,
    \Tile_X1Y9_W2BEGb[3] ,
    \Tile_X1Y9_W2BEGb[2] ,
    \Tile_X1Y9_W2BEGb[1] ,
    \Tile_X1Y9_W2BEGb[0] }),
    .W2MID({\Tile_X1Y9_W2BEG[7] ,
    \Tile_X1Y9_W2BEG[6] ,
    \Tile_X1Y9_W2BEG[5] ,
    \Tile_X1Y9_W2BEG[4] ,
    \Tile_X1Y9_W2BEG[3] ,
    \Tile_X1Y9_W2BEG[2] ,
    \Tile_X1Y9_W2BEG[1] ,
    \Tile_X1Y9_W2BEG[0] }),
    .W6END({\Tile_X1Y9_W6BEG[11] ,
    \Tile_X1Y9_W6BEG[10] ,
    \Tile_X1Y9_W6BEG[9] ,
    \Tile_X1Y9_W6BEG[8] ,
    \Tile_X1Y9_W6BEG[7] ,
    \Tile_X1Y9_W6BEG[6] ,
    \Tile_X1Y9_W6BEG[5] ,
    \Tile_X1Y9_W6BEG[4] ,
    \Tile_X1Y9_W6BEG[3] ,
    \Tile_X1Y9_W6BEG[2] ,
    \Tile_X1Y9_W6BEG[1] ,
    \Tile_X1Y9_W6BEG[0] }),
    .WW4END({\Tile_X1Y9_WW4BEG[15] ,
    \Tile_X1Y9_WW4BEG[14] ,
    \Tile_X1Y9_WW4BEG[13] ,
    \Tile_X1Y9_WW4BEG[12] ,
    \Tile_X1Y9_WW4BEG[11] ,
    \Tile_X1Y9_WW4BEG[10] ,
    \Tile_X1Y9_WW4BEG[9] ,
    \Tile_X1Y9_WW4BEG[8] ,
    \Tile_X1Y9_WW4BEG[7] ,
    \Tile_X1Y9_WW4BEG[6] ,
    \Tile_X1Y9_WW4BEG[5] ,
    \Tile_X1Y9_WW4BEG[4] ,
    \Tile_X1Y9_WW4BEG[3] ,
    \Tile_X1Y9_WW4BEG[2] ,
    \Tile_X1Y9_WW4BEG[1] ,
    \Tile_X1Y9_WW4BEG[0] }));
 N_term_IHP_SRAM Tile_X10Y0_N_term_IHP_SRAM (.UserCLK(Tile_X10Y1_UserCLKo),
    .UserCLKo(Tile_X10Y0_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .FrameData({\Tile_X9Y0_FrameData_O[31] ,
    \Tile_X9Y0_FrameData_O[30] ,
    \Tile_X9Y0_FrameData_O[29] ,
    \Tile_X9Y0_FrameData_O[28] ,
    \Tile_X9Y0_FrameData_O[27] ,
    \Tile_X9Y0_FrameData_O[26] ,
    \Tile_X9Y0_FrameData_O[25] ,
    \Tile_X9Y0_FrameData_O[24] ,
    \Tile_X9Y0_FrameData_O[23] ,
    \Tile_X9Y0_FrameData_O[22] ,
    \Tile_X9Y0_FrameData_O[21] ,
    \Tile_X9Y0_FrameData_O[20] ,
    \Tile_X9Y0_FrameData_O[19] ,
    \Tile_X9Y0_FrameData_O[18] ,
    \Tile_X9Y0_FrameData_O[17] ,
    \Tile_X9Y0_FrameData_O[16] ,
    \Tile_X9Y0_FrameData_O[15] ,
    \Tile_X9Y0_FrameData_O[14] ,
    \Tile_X9Y0_FrameData_O[13] ,
    \Tile_X9Y0_FrameData_O[12] ,
    \Tile_X9Y0_FrameData_O[11] ,
    \Tile_X9Y0_FrameData_O[10] ,
    \Tile_X9Y0_FrameData_O[9] ,
    \Tile_X9Y0_FrameData_O[8] ,
    \Tile_X9Y0_FrameData_O[7] ,
    \Tile_X9Y0_FrameData_O[6] ,
    \Tile_X9Y0_FrameData_O[5] ,
    \Tile_X9Y0_FrameData_O[4] ,
    \Tile_X9Y0_FrameData_O[3] ,
    \Tile_X9Y0_FrameData_O[2] ,
    \Tile_X9Y0_FrameData_O[1] ,
    \Tile_X9Y0_FrameData_O[0] }),
    .FrameData_O({\Tile_X10Y0_FrameData_O[31] ,
    \Tile_X10Y0_FrameData_O[30] ,
    \Tile_X10Y0_FrameData_O[29] ,
    \Tile_X10Y0_FrameData_O[28] ,
    \Tile_X10Y0_FrameData_O[27] ,
    \Tile_X10Y0_FrameData_O[26] ,
    \Tile_X10Y0_FrameData_O[25] ,
    \Tile_X10Y0_FrameData_O[24] ,
    \Tile_X10Y0_FrameData_O[23] ,
    \Tile_X10Y0_FrameData_O[22] ,
    \Tile_X10Y0_FrameData_O[21] ,
    \Tile_X10Y0_FrameData_O[20] ,
    \Tile_X10Y0_FrameData_O[19] ,
    \Tile_X10Y0_FrameData_O[18] ,
    \Tile_X10Y0_FrameData_O[17] ,
    \Tile_X10Y0_FrameData_O[16] ,
    \Tile_X10Y0_FrameData_O[15] ,
    \Tile_X10Y0_FrameData_O[14] ,
    \Tile_X10Y0_FrameData_O[13] ,
    \Tile_X10Y0_FrameData_O[12] ,
    \Tile_X10Y0_FrameData_O[11] ,
    \Tile_X10Y0_FrameData_O[10] ,
    \Tile_X10Y0_FrameData_O[9] ,
    \Tile_X10Y0_FrameData_O[8] ,
    \Tile_X10Y0_FrameData_O[7] ,
    \Tile_X10Y0_FrameData_O[6] ,
    \Tile_X10Y0_FrameData_O[5] ,
    \Tile_X10Y0_FrameData_O[4] ,
    \Tile_X10Y0_FrameData_O[3] ,
    \Tile_X10Y0_FrameData_O[2] ,
    \Tile_X10Y0_FrameData_O[1] ,
    \Tile_X10Y0_FrameData_O[0] }),
    .FrameStrobe({\Tile_X10Y1_FrameStrobe_O[19] ,
    \Tile_X10Y1_FrameStrobe_O[18] ,
    \Tile_X10Y1_FrameStrobe_O[17] ,
    \Tile_X10Y1_FrameStrobe_O[16] ,
    \Tile_X10Y1_FrameStrobe_O[15] ,
    \Tile_X10Y1_FrameStrobe_O[14] ,
    \Tile_X10Y1_FrameStrobe_O[13] ,
    \Tile_X10Y1_FrameStrobe_O[12] ,
    \Tile_X10Y1_FrameStrobe_O[11] ,
    \Tile_X10Y1_FrameStrobe_O[10] ,
    \Tile_X10Y1_FrameStrobe_O[9] ,
    \Tile_X10Y1_FrameStrobe_O[8] ,
    \Tile_X10Y1_FrameStrobe_O[7] ,
    \Tile_X10Y1_FrameStrobe_O[6] ,
    \Tile_X10Y1_FrameStrobe_O[5] ,
    \Tile_X10Y1_FrameStrobe_O[4] ,
    \Tile_X10Y1_FrameStrobe_O[3] ,
    \Tile_X10Y1_FrameStrobe_O[2] ,
    \Tile_X10Y1_FrameStrobe_O[1] ,
    \Tile_X10Y1_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X10Y0_FrameStrobe_O[19] ,
    \Tile_X10Y0_FrameStrobe_O[18] ,
    \Tile_X10Y0_FrameStrobe_O[17] ,
    \Tile_X10Y0_FrameStrobe_O[16] ,
    \Tile_X10Y0_FrameStrobe_O[15] ,
    \Tile_X10Y0_FrameStrobe_O[14] ,
    \Tile_X10Y0_FrameStrobe_O[13] ,
    \Tile_X10Y0_FrameStrobe_O[12] ,
    \Tile_X10Y0_FrameStrobe_O[11] ,
    \Tile_X10Y0_FrameStrobe_O[10] ,
    \Tile_X10Y0_FrameStrobe_O[9] ,
    \Tile_X10Y0_FrameStrobe_O[8] ,
    \Tile_X10Y0_FrameStrobe_O[7] ,
    \Tile_X10Y0_FrameStrobe_O[6] ,
    \Tile_X10Y0_FrameStrobe_O[5] ,
    \Tile_X10Y0_FrameStrobe_O[4] ,
    \Tile_X10Y0_FrameStrobe_O[3] ,
    \Tile_X10Y0_FrameStrobe_O[2] ,
    \Tile_X10Y0_FrameStrobe_O[1] ,
    \Tile_X10Y0_FrameStrobe_O[0] }),
    .N1END({\Tile_X10Y1_N1BEG[3] ,
    \Tile_X10Y1_N1BEG[2] ,
    \Tile_X10Y1_N1BEG[1] ,
    \Tile_X10Y1_N1BEG[0] }),
    .N2END({\Tile_X10Y1_N2BEGb[7] ,
    \Tile_X10Y1_N2BEGb[6] ,
    \Tile_X10Y1_N2BEGb[5] ,
    \Tile_X10Y1_N2BEGb[4] ,
    \Tile_X10Y1_N2BEGb[3] ,
    \Tile_X10Y1_N2BEGb[2] ,
    \Tile_X10Y1_N2BEGb[1] ,
    \Tile_X10Y1_N2BEGb[0] }),
    .N2MID({\Tile_X10Y1_N2BEG[7] ,
    \Tile_X10Y1_N2BEG[6] ,
    \Tile_X10Y1_N2BEG[5] ,
    \Tile_X10Y1_N2BEG[4] ,
    \Tile_X10Y1_N2BEG[3] ,
    \Tile_X10Y1_N2BEG[2] ,
    \Tile_X10Y1_N2BEG[1] ,
    \Tile_X10Y1_N2BEG[0] }),
    .N4END({\Tile_X10Y1_N4BEG[15] ,
    \Tile_X10Y1_N4BEG[14] ,
    \Tile_X10Y1_N4BEG[13] ,
    \Tile_X10Y1_N4BEG[12] ,
    \Tile_X10Y1_N4BEG[11] ,
    \Tile_X10Y1_N4BEG[10] ,
    \Tile_X10Y1_N4BEG[9] ,
    \Tile_X10Y1_N4BEG[8] ,
    \Tile_X10Y1_N4BEG[7] ,
    \Tile_X10Y1_N4BEG[6] ,
    \Tile_X10Y1_N4BEG[5] ,
    \Tile_X10Y1_N4BEG[4] ,
    \Tile_X10Y1_N4BEG[3] ,
    \Tile_X10Y1_N4BEG[2] ,
    \Tile_X10Y1_N4BEG[1] ,
    \Tile_X10Y1_N4BEG[0] }),
    .S1BEG({\Tile_X10Y0_S1BEG[3] ,
    \Tile_X10Y0_S1BEG[2] ,
    \Tile_X10Y0_S1BEG[1] ,
    \Tile_X10Y0_S1BEG[0] }),
    .S2BEG({\Tile_X10Y0_S2BEG[7] ,
    \Tile_X10Y0_S2BEG[6] ,
    \Tile_X10Y0_S2BEG[5] ,
    \Tile_X10Y0_S2BEG[4] ,
    \Tile_X10Y0_S2BEG[3] ,
    \Tile_X10Y0_S2BEG[2] ,
    \Tile_X10Y0_S2BEG[1] ,
    \Tile_X10Y0_S2BEG[0] }),
    .S2BEGb({\Tile_X10Y0_S2BEGb[7] ,
    \Tile_X10Y0_S2BEGb[6] ,
    \Tile_X10Y0_S2BEGb[5] ,
    \Tile_X10Y0_S2BEGb[4] ,
    \Tile_X10Y0_S2BEGb[3] ,
    \Tile_X10Y0_S2BEGb[2] ,
    \Tile_X10Y0_S2BEGb[1] ,
    \Tile_X10Y0_S2BEGb[0] }),
    .S4BEG({\Tile_X10Y0_S4BEG[15] ,
    \Tile_X10Y0_S4BEG[14] ,
    \Tile_X10Y0_S4BEG[13] ,
    \Tile_X10Y0_S4BEG[12] ,
    \Tile_X10Y0_S4BEG[11] ,
    \Tile_X10Y0_S4BEG[10] ,
    \Tile_X10Y0_S4BEG[9] ,
    \Tile_X10Y0_S4BEG[8] ,
    \Tile_X10Y0_S4BEG[7] ,
    \Tile_X10Y0_S4BEG[6] ,
    \Tile_X10Y0_S4BEG[5] ,
    \Tile_X10Y0_S4BEG[4] ,
    \Tile_X10Y0_S4BEG[3] ,
    \Tile_X10Y0_S4BEG[2] ,
    \Tile_X10Y0_S4BEG[1] ,
    \Tile_X10Y0_S4BEG[0] }));
 IHP_SRAM Tile_X10Y11_IHP_SRAM (.ADDR_SRAM0(Tile_X10Y12_ADDR_SRAM0),
    .ADDR_SRAM1(Tile_X10Y12_ADDR_SRAM1),
    .ADDR_SRAM2(Tile_X10Y12_ADDR_SRAM2),
    .ADDR_SRAM3(Tile_X10Y12_ADDR_SRAM3),
    .ADDR_SRAM4(Tile_X10Y12_ADDR_SRAM4),
    .ADDR_SRAM5(Tile_X10Y12_ADDR_SRAM5),
    .ADDR_SRAM6(Tile_X10Y12_ADDR_SRAM6),
    .ADDR_SRAM7(Tile_X10Y12_ADDR_SRAM7),
    .ADDR_SRAM8(Tile_X10Y12_ADDR_SRAM8),
    .ADDR_SRAM9(Tile_X10Y12_ADDR_SRAM9),
    .BM_SRAM0(Tile_X10Y12_BM_SRAM0),
    .BM_SRAM1(Tile_X10Y12_BM_SRAM1),
    .BM_SRAM10(Tile_X10Y12_BM_SRAM10),
    .BM_SRAM11(Tile_X10Y12_BM_SRAM11),
    .BM_SRAM12(Tile_X10Y12_BM_SRAM12),
    .BM_SRAM13(Tile_X10Y12_BM_SRAM13),
    .BM_SRAM14(Tile_X10Y12_BM_SRAM14),
    .BM_SRAM15(Tile_X10Y12_BM_SRAM15),
    .BM_SRAM16(Tile_X10Y12_BM_SRAM16),
    .BM_SRAM17(Tile_X10Y12_BM_SRAM17),
    .BM_SRAM18(Tile_X10Y12_BM_SRAM18),
    .BM_SRAM19(Tile_X10Y12_BM_SRAM19),
    .BM_SRAM2(Tile_X10Y12_BM_SRAM2),
    .BM_SRAM20(Tile_X10Y12_BM_SRAM20),
    .BM_SRAM21(Tile_X10Y12_BM_SRAM21),
    .BM_SRAM22(Tile_X10Y12_BM_SRAM22),
    .BM_SRAM23(Tile_X10Y12_BM_SRAM23),
    .BM_SRAM24(Tile_X10Y12_BM_SRAM24),
    .BM_SRAM25(Tile_X10Y12_BM_SRAM25),
    .BM_SRAM26(Tile_X10Y12_BM_SRAM26),
    .BM_SRAM27(Tile_X10Y12_BM_SRAM27),
    .BM_SRAM28(Tile_X10Y12_BM_SRAM28),
    .BM_SRAM29(Tile_X10Y12_BM_SRAM29),
    .BM_SRAM3(Tile_X10Y12_BM_SRAM3),
    .BM_SRAM30(Tile_X10Y12_BM_SRAM30),
    .BM_SRAM31(Tile_X10Y12_BM_SRAM31),
    .BM_SRAM4(Tile_X10Y12_BM_SRAM4),
    .BM_SRAM5(Tile_X10Y12_BM_SRAM5),
    .BM_SRAM6(Tile_X10Y12_BM_SRAM6),
    .BM_SRAM7(Tile_X10Y12_BM_SRAM7),
    .BM_SRAM8(Tile_X10Y12_BM_SRAM8),
    .BM_SRAM9(Tile_X10Y12_BM_SRAM9),
    .CLK_SRAM(Tile_X10Y12_CLK_SRAM),
    .CONFIGURED_top(Tile_X10Y12_CONFIGURED_top),
    .DIN_SRAM0(Tile_X10Y12_DIN_SRAM0),
    .DIN_SRAM1(Tile_X10Y12_DIN_SRAM1),
    .DIN_SRAM10(Tile_X10Y12_DIN_SRAM10),
    .DIN_SRAM11(Tile_X10Y12_DIN_SRAM11),
    .DIN_SRAM12(Tile_X10Y12_DIN_SRAM12),
    .DIN_SRAM13(Tile_X10Y12_DIN_SRAM13),
    .DIN_SRAM14(Tile_X10Y12_DIN_SRAM14),
    .DIN_SRAM15(Tile_X10Y12_DIN_SRAM15),
    .DIN_SRAM16(Tile_X10Y12_DIN_SRAM16),
    .DIN_SRAM17(Tile_X10Y12_DIN_SRAM17),
    .DIN_SRAM18(Tile_X10Y12_DIN_SRAM18),
    .DIN_SRAM19(Tile_X10Y12_DIN_SRAM19),
    .DIN_SRAM2(Tile_X10Y12_DIN_SRAM2),
    .DIN_SRAM20(Tile_X10Y12_DIN_SRAM20),
    .DIN_SRAM21(Tile_X10Y12_DIN_SRAM21),
    .DIN_SRAM22(Tile_X10Y12_DIN_SRAM22),
    .DIN_SRAM23(Tile_X10Y12_DIN_SRAM23),
    .DIN_SRAM24(Tile_X10Y12_DIN_SRAM24),
    .DIN_SRAM25(Tile_X10Y12_DIN_SRAM25),
    .DIN_SRAM26(Tile_X10Y12_DIN_SRAM26),
    .DIN_SRAM27(Tile_X10Y12_DIN_SRAM27),
    .DIN_SRAM28(Tile_X10Y12_DIN_SRAM28),
    .DIN_SRAM29(Tile_X10Y12_DIN_SRAM29),
    .DIN_SRAM3(Tile_X10Y12_DIN_SRAM3),
    .DIN_SRAM30(Tile_X10Y12_DIN_SRAM30),
    .DIN_SRAM31(Tile_X10Y12_DIN_SRAM31),
    .DIN_SRAM4(Tile_X10Y12_DIN_SRAM4),
    .DIN_SRAM5(Tile_X10Y12_DIN_SRAM5),
    .DIN_SRAM6(Tile_X10Y12_DIN_SRAM6),
    .DIN_SRAM7(Tile_X10Y12_DIN_SRAM7),
    .DIN_SRAM8(Tile_X10Y12_DIN_SRAM8),
    .DIN_SRAM9(Tile_X10Y12_DIN_SRAM9),
    .DOUT_SRAM0(Tile_X10Y12_DOUT_SRAM0),
    .DOUT_SRAM1(Tile_X10Y12_DOUT_SRAM1),
    .DOUT_SRAM10(Tile_X10Y12_DOUT_SRAM10),
    .DOUT_SRAM11(Tile_X10Y12_DOUT_SRAM11),
    .DOUT_SRAM12(Tile_X10Y12_DOUT_SRAM12),
    .DOUT_SRAM13(Tile_X10Y12_DOUT_SRAM13),
    .DOUT_SRAM14(Tile_X10Y12_DOUT_SRAM14),
    .DOUT_SRAM15(Tile_X10Y12_DOUT_SRAM15),
    .DOUT_SRAM16(Tile_X10Y12_DOUT_SRAM16),
    .DOUT_SRAM17(Tile_X10Y12_DOUT_SRAM17),
    .DOUT_SRAM18(Tile_X10Y12_DOUT_SRAM18),
    .DOUT_SRAM19(Tile_X10Y12_DOUT_SRAM19),
    .DOUT_SRAM2(Tile_X10Y12_DOUT_SRAM2),
    .DOUT_SRAM20(Tile_X10Y12_DOUT_SRAM20),
    .DOUT_SRAM21(Tile_X10Y12_DOUT_SRAM21),
    .DOUT_SRAM22(Tile_X10Y12_DOUT_SRAM22),
    .DOUT_SRAM23(Tile_X10Y12_DOUT_SRAM23),
    .DOUT_SRAM24(Tile_X10Y12_DOUT_SRAM24),
    .DOUT_SRAM25(Tile_X10Y12_DOUT_SRAM25),
    .DOUT_SRAM26(Tile_X10Y12_DOUT_SRAM26),
    .DOUT_SRAM27(Tile_X10Y12_DOUT_SRAM27),
    .DOUT_SRAM28(Tile_X10Y12_DOUT_SRAM28),
    .DOUT_SRAM29(Tile_X10Y12_DOUT_SRAM29),
    .DOUT_SRAM3(Tile_X10Y12_DOUT_SRAM3),
    .DOUT_SRAM30(Tile_X10Y12_DOUT_SRAM30),
    .DOUT_SRAM31(Tile_X10Y12_DOUT_SRAM31),
    .DOUT_SRAM4(Tile_X10Y12_DOUT_SRAM4),
    .DOUT_SRAM5(Tile_X10Y12_DOUT_SRAM5),
    .DOUT_SRAM6(Tile_X10Y12_DOUT_SRAM6),
    .DOUT_SRAM7(Tile_X10Y12_DOUT_SRAM7),
    .DOUT_SRAM8(Tile_X10Y12_DOUT_SRAM8),
    .DOUT_SRAM9(Tile_X10Y12_DOUT_SRAM9),
    .MEN_SRAM(Tile_X10Y12_MEN_SRAM),
    .REN_SRAM(Tile_X10Y12_REN_SRAM),
    .TIE_HIGH_SRAM(Tile_X10Y12_TIE_HIGH_SRAM),
    .TIE_LOW_SRAM(Tile_X10Y12_TIE_LOW_SRAM),
    .Tile_X0Y0_UserCLKo(Tile_X10Y11_UserCLKo),
    .Tile_X0Y1_UserCLK(Tile_X10Y13_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .WEN_SRAM(Tile_X10Y12_WEN_SRAM),
    .Tile_X0Y0_E1END({\Tile_X9Y11_E1BEG[3] ,
    \Tile_X9Y11_E1BEG[2] ,
    \Tile_X9Y11_E1BEG[1] ,
    \Tile_X9Y11_E1BEG[0] }),
    .Tile_X0Y0_E2END({\Tile_X9Y11_E2BEGb[7] ,
    \Tile_X9Y11_E2BEGb[6] ,
    \Tile_X9Y11_E2BEGb[5] ,
    \Tile_X9Y11_E2BEGb[4] ,
    \Tile_X9Y11_E2BEGb[3] ,
    \Tile_X9Y11_E2BEGb[2] ,
    \Tile_X9Y11_E2BEGb[1] ,
    \Tile_X9Y11_E2BEGb[0] }),
    .Tile_X0Y0_E2MID({\Tile_X9Y11_E2BEG[7] ,
    \Tile_X9Y11_E2BEG[6] ,
    \Tile_X9Y11_E2BEG[5] ,
    \Tile_X9Y11_E2BEG[4] ,
    \Tile_X9Y11_E2BEG[3] ,
    \Tile_X9Y11_E2BEG[2] ,
    \Tile_X9Y11_E2BEG[1] ,
    \Tile_X9Y11_E2BEG[0] }),
    .Tile_X0Y0_E6END({\Tile_X9Y11_E6BEG[11] ,
    \Tile_X9Y11_E6BEG[10] ,
    \Tile_X9Y11_E6BEG[9] ,
    \Tile_X9Y11_E6BEG[8] ,
    \Tile_X9Y11_E6BEG[7] ,
    \Tile_X9Y11_E6BEG[6] ,
    \Tile_X9Y11_E6BEG[5] ,
    \Tile_X9Y11_E6BEG[4] ,
    \Tile_X9Y11_E6BEG[3] ,
    \Tile_X9Y11_E6BEG[2] ,
    \Tile_X9Y11_E6BEG[1] ,
    \Tile_X9Y11_E6BEG[0] }),
    .Tile_X0Y0_EE4END({\Tile_X9Y11_EE4BEG[15] ,
    \Tile_X9Y11_EE4BEG[14] ,
    \Tile_X9Y11_EE4BEG[13] ,
    \Tile_X9Y11_EE4BEG[12] ,
    \Tile_X9Y11_EE4BEG[11] ,
    \Tile_X9Y11_EE4BEG[10] ,
    \Tile_X9Y11_EE4BEG[9] ,
    \Tile_X9Y11_EE4BEG[8] ,
    \Tile_X9Y11_EE4BEG[7] ,
    \Tile_X9Y11_EE4BEG[6] ,
    \Tile_X9Y11_EE4BEG[5] ,
    \Tile_X9Y11_EE4BEG[4] ,
    \Tile_X9Y11_EE4BEG[3] ,
    \Tile_X9Y11_EE4BEG[2] ,
    \Tile_X9Y11_EE4BEG[1] ,
    \Tile_X9Y11_EE4BEG[0] }),
    .Tile_X0Y0_FrameData({\Tile_X9Y11_FrameData_O[31] ,
    \Tile_X9Y11_FrameData_O[30] ,
    \Tile_X9Y11_FrameData_O[29] ,
    \Tile_X9Y11_FrameData_O[28] ,
    \Tile_X9Y11_FrameData_O[27] ,
    \Tile_X9Y11_FrameData_O[26] ,
    \Tile_X9Y11_FrameData_O[25] ,
    \Tile_X9Y11_FrameData_O[24] ,
    \Tile_X9Y11_FrameData_O[23] ,
    \Tile_X9Y11_FrameData_O[22] ,
    \Tile_X9Y11_FrameData_O[21] ,
    \Tile_X9Y11_FrameData_O[20] ,
    \Tile_X9Y11_FrameData_O[19] ,
    \Tile_X9Y11_FrameData_O[18] ,
    \Tile_X9Y11_FrameData_O[17] ,
    \Tile_X9Y11_FrameData_O[16] ,
    \Tile_X9Y11_FrameData_O[15] ,
    \Tile_X9Y11_FrameData_O[14] ,
    \Tile_X9Y11_FrameData_O[13] ,
    \Tile_X9Y11_FrameData_O[12] ,
    \Tile_X9Y11_FrameData_O[11] ,
    \Tile_X9Y11_FrameData_O[10] ,
    \Tile_X9Y11_FrameData_O[9] ,
    \Tile_X9Y11_FrameData_O[8] ,
    \Tile_X9Y11_FrameData_O[7] ,
    \Tile_X9Y11_FrameData_O[6] ,
    \Tile_X9Y11_FrameData_O[5] ,
    \Tile_X9Y11_FrameData_O[4] ,
    \Tile_X9Y11_FrameData_O[3] ,
    \Tile_X9Y11_FrameData_O[2] ,
    \Tile_X9Y11_FrameData_O[1] ,
    \Tile_X9Y11_FrameData_O[0] }),
    .Tile_X0Y0_FrameData_O({\Tile_X10Y11_FrameData_O[31] ,
    \Tile_X10Y11_FrameData_O[30] ,
    \Tile_X10Y11_FrameData_O[29] ,
    \Tile_X10Y11_FrameData_O[28] ,
    \Tile_X10Y11_FrameData_O[27] ,
    \Tile_X10Y11_FrameData_O[26] ,
    \Tile_X10Y11_FrameData_O[25] ,
    \Tile_X10Y11_FrameData_O[24] ,
    \Tile_X10Y11_FrameData_O[23] ,
    \Tile_X10Y11_FrameData_O[22] ,
    \Tile_X10Y11_FrameData_O[21] ,
    \Tile_X10Y11_FrameData_O[20] ,
    \Tile_X10Y11_FrameData_O[19] ,
    \Tile_X10Y11_FrameData_O[18] ,
    \Tile_X10Y11_FrameData_O[17] ,
    \Tile_X10Y11_FrameData_O[16] ,
    \Tile_X10Y11_FrameData_O[15] ,
    \Tile_X10Y11_FrameData_O[14] ,
    \Tile_X10Y11_FrameData_O[13] ,
    \Tile_X10Y11_FrameData_O[12] ,
    \Tile_X10Y11_FrameData_O[11] ,
    \Tile_X10Y11_FrameData_O[10] ,
    \Tile_X10Y11_FrameData_O[9] ,
    \Tile_X10Y11_FrameData_O[8] ,
    \Tile_X10Y11_FrameData_O[7] ,
    \Tile_X10Y11_FrameData_O[6] ,
    \Tile_X10Y11_FrameData_O[5] ,
    \Tile_X10Y11_FrameData_O[4] ,
    \Tile_X10Y11_FrameData_O[3] ,
    \Tile_X10Y11_FrameData_O[2] ,
    \Tile_X10Y11_FrameData_O[1] ,
    \Tile_X10Y11_FrameData_O[0] }),
    .Tile_X0Y0_FrameStrobe_O({\Tile_X10Y11_FrameStrobe_O[19] ,
    \Tile_X10Y11_FrameStrobe_O[18] ,
    \Tile_X10Y11_FrameStrobe_O[17] ,
    \Tile_X10Y11_FrameStrobe_O[16] ,
    \Tile_X10Y11_FrameStrobe_O[15] ,
    \Tile_X10Y11_FrameStrobe_O[14] ,
    \Tile_X10Y11_FrameStrobe_O[13] ,
    \Tile_X10Y11_FrameStrobe_O[12] ,
    \Tile_X10Y11_FrameStrobe_O[11] ,
    \Tile_X10Y11_FrameStrobe_O[10] ,
    \Tile_X10Y11_FrameStrobe_O[9] ,
    \Tile_X10Y11_FrameStrobe_O[8] ,
    \Tile_X10Y11_FrameStrobe_O[7] ,
    \Tile_X10Y11_FrameStrobe_O[6] ,
    \Tile_X10Y11_FrameStrobe_O[5] ,
    \Tile_X10Y11_FrameStrobe_O[4] ,
    \Tile_X10Y11_FrameStrobe_O[3] ,
    \Tile_X10Y11_FrameStrobe_O[2] ,
    \Tile_X10Y11_FrameStrobe_O[1] ,
    \Tile_X10Y11_FrameStrobe_O[0] }),
    .Tile_X0Y0_N1BEG({\Tile_X10Y11_N1BEG[3] ,
    \Tile_X10Y11_N1BEG[2] ,
    \Tile_X10Y11_N1BEG[1] ,
    \Tile_X10Y11_N1BEG[0] }),
    .Tile_X0Y0_N2BEG({\Tile_X10Y11_N2BEG[7] ,
    \Tile_X10Y11_N2BEG[6] ,
    \Tile_X10Y11_N2BEG[5] ,
    \Tile_X10Y11_N2BEG[4] ,
    \Tile_X10Y11_N2BEG[3] ,
    \Tile_X10Y11_N2BEG[2] ,
    \Tile_X10Y11_N2BEG[1] ,
    \Tile_X10Y11_N2BEG[0] }),
    .Tile_X0Y0_N2BEGb({\Tile_X10Y11_N2BEGb[7] ,
    \Tile_X10Y11_N2BEGb[6] ,
    \Tile_X10Y11_N2BEGb[5] ,
    \Tile_X10Y11_N2BEGb[4] ,
    \Tile_X10Y11_N2BEGb[3] ,
    \Tile_X10Y11_N2BEGb[2] ,
    \Tile_X10Y11_N2BEGb[1] ,
    \Tile_X10Y11_N2BEGb[0] }),
    .Tile_X0Y0_N4BEG({\Tile_X10Y11_N4BEG[15] ,
    \Tile_X10Y11_N4BEG[14] ,
    \Tile_X10Y11_N4BEG[13] ,
    \Tile_X10Y11_N4BEG[12] ,
    \Tile_X10Y11_N4BEG[11] ,
    \Tile_X10Y11_N4BEG[10] ,
    \Tile_X10Y11_N4BEG[9] ,
    \Tile_X10Y11_N4BEG[8] ,
    \Tile_X10Y11_N4BEG[7] ,
    \Tile_X10Y11_N4BEG[6] ,
    \Tile_X10Y11_N4BEG[5] ,
    \Tile_X10Y11_N4BEG[4] ,
    \Tile_X10Y11_N4BEG[3] ,
    \Tile_X10Y11_N4BEG[2] ,
    \Tile_X10Y11_N4BEG[1] ,
    \Tile_X10Y11_N4BEG[0] }),
    .Tile_X0Y0_S1END({\Tile_X10Y10_S1BEG[3] ,
    \Tile_X10Y10_S1BEG[2] ,
    \Tile_X10Y10_S1BEG[1] ,
    \Tile_X10Y10_S1BEG[0] }),
    .Tile_X0Y0_S2END({\Tile_X10Y10_S2BEGb[7] ,
    \Tile_X10Y10_S2BEGb[6] ,
    \Tile_X10Y10_S2BEGb[5] ,
    \Tile_X10Y10_S2BEGb[4] ,
    \Tile_X10Y10_S2BEGb[3] ,
    \Tile_X10Y10_S2BEGb[2] ,
    \Tile_X10Y10_S2BEGb[1] ,
    \Tile_X10Y10_S2BEGb[0] }),
    .Tile_X0Y0_S2MID({\Tile_X10Y10_S2BEG[7] ,
    \Tile_X10Y10_S2BEG[6] ,
    \Tile_X10Y10_S2BEG[5] ,
    \Tile_X10Y10_S2BEG[4] ,
    \Tile_X10Y10_S2BEG[3] ,
    \Tile_X10Y10_S2BEG[2] ,
    \Tile_X10Y10_S2BEG[1] ,
    \Tile_X10Y10_S2BEG[0] }),
    .Tile_X0Y0_S4END({\Tile_X10Y10_S4BEG[15] ,
    \Tile_X10Y10_S4BEG[14] ,
    \Tile_X10Y10_S4BEG[13] ,
    \Tile_X10Y10_S4BEG[12] ,
    \Tile_X10Y10_S4BEG[11] ,
    \Tile_X10Y10_S4BEG[10] ,
    \Tile_X10Y10_S4BEG[9] ,
    \Tile_X10Y10_S4BEG[8] ,
    \Tile_X10Y10_S4BEG[7] ,
    \Tile_X10Y10_S4BEG[6] ,
    \Tile_X10Y10_S4BEG[5] ,
    \Tile_X10Y10_S4BEG[4] ,
    \Tile_X10Y10_S4BEG[3] ,
    \Tile_X10Y10_S4BEG[2] ,
    \Tile_X10Y10_S4BEG[1] ,
    \Tile_X10Y10_S4BEG[0] }),
    .Tile_X0Y0_W1BEG({\Tile_X10Y11_W1BEG[3] ,
    \Tile_X10Y11_W1BEG[2] ,
    \Tile_X10Y11_W1BEG[1] ,
    \Tile_X10Y11_W1BEG[0] }),
    .Tile_X0Y0_W2BEG({\Tile_X10Y11_W2BEG[7] ,
    \Tile_X10Y11_W2BEG[6] ,
    \Tile_X10Y11_W2BEG[5] ,
    \Tile_X10Y11_W2BEG[4] ,
    \Tile_X10Y11_W2BEG[3] ,
    \Tile_X10Y11_W2BEG[2] ,
    \Tile_X10Y11_W2BEG[1] ,
    \Tile_X10Y11_W2BEG[0] }),
    .Tile_X0Y0_W2BEGb({\Tile_X10Y11_W2BEGb[7] ,
    \Tile_X10Y11_W2BEGb[6] ,
    \Tile_X10Y11_W2BEGb[5] ,
    \Tile_X10Y11_W2BEGb[4] ,
    \Tile_X10Y11_W2BEGb[3] ,
    \Tile_X10Y11_W2BEGb[2] ,
    \Tile_X10Y11_W2BEGb[1] ,
    \Tile_X10Y11_W2BEGb[0] }),
    .Tile_X0Y0_W6BEG({\Tile_X10Y11_W6BEG[11] ,
    \Tile_X10Y11_W6BEG[10] ,
    \Tile_X10Y11_W6BEG[9] ,
    \Tile_X10Y11_W6BEG[8] ,
    \Tile_X10Y11_W6BEG[7] ,
    \Tile_X10Y11_W6BEG[6] ,
    \Tile_X10Y11_W6BEG[5] ,
    \Tile_X10Y11_W6BEG[4] ,
    \Tile_X10Y11_W6BEG[3] ,
    \Tile_X10Y11_W6BEG[2] ,
    \Tile_X10Y11_W6BEG[1] ,
    \Tile_X10Y11_W6BEG[0] }),
    .Tile_X0Y0_WW4BEG({\Tile_X10Y11_WW4BEG[15] ,
    \Tile_X10Y11_WW4BEG[14] ,
    \Tile_X10Y11_WW4BEG[13] ,
    \Tile_X10Y11_WW4BEG[12] ,
    \Tile_X10Y11_WW4BEG[11] ,
    \Tile_X10Y11_WW4BEG[10] ,
    \Tile_X10Y11_WW4BEG[9] ,
    \Tile_X10Y11_WW4BEG[8] ,
    \Tile_X10Y11_WW4BEG[7] ,
    \Tile_X10Y11_WW4BEG[6] ,
    \Tile_X10Y11_WW4BEG[5] ,
    \Tile_X10Y11_WW4BEG[4] ,
    \Tile_X10Y11_WW4BEG[3] ,
    \Tile_X10Y11_WW4BEG[2] ,
    \Tile_X10Y11_WW4BEG[1] ,
    \Tile_X10Y11_WW4BEG[0] }),
    .Tile_X0Y1_E1END({\Tile_X9Y12_E1BEG[3] ,
    \Tile_X9Y12_E1BEG[2] ,
    \Tile_X9Y12_E1BEG[1] ,
    \Tile_X9Y12_E1BEG[0] }),
    .Tile_X0Y1_E2END({\Tile_X9Y12_E2BEGb[7] ,
    \Tile_X9Y12_E2BEGb[6] ,
    \Tile_X9Y12_E2BEGb[5] ,
    \Tile_X9Y12_E2BEGb[4] ,
    \Tile_X9Y12_E2BEGb[3] ,
    \Tile_X9Y12_E2BEGb[2] ,
    \Tile_X9Y12_E2BEGb[1] ,
    \Tile_X9Y12_E2BEGb[0] }),
    .Tile_X0Y1_E2MID({\Tile_X9Y12_E2BEG[7] ,
    \Tile_X9Y12_E2BEG[6] ,
    \Tile_X9Y12_E2BEG[5] ,
    \Tile_X9Y12_E2BEG[4] ,
    \Tile_X9Y12_E2BEG[3] ,
    \Tile_X9Y12_E2BEG[2] ,
    \Tile_X9Y12_E2BEG[1] ,
    \Tile_X9Y12_E2BEG[0] }),
    .Tile_X0Y1_E6END({\Tile_X9Y12_E6BEG[11] ,
    \Tile_X9Y12_E6BEG[10] ,
    \Tile_X9Y12_E6BEG[9] ,
    \Tile_X9Y12_E6BEG[8] ,
    \Tile_X9Y12_E6BEG[7] ,
    \Tile_X9Y12_E6BEG[6] ,
    \Tile_X9Y12_E6BEG[5] ,
    \Tile_X9Y12_E6BEG[4] ,
    \Tile_X9Y12_E6BEG[3] ,
    \Tile_X9Y12_E6BEG[2] ,
    \Tile_X9Y12_E6BEG[1] ,
    \Tile_X9Y12_E6BEG[0] }),
    .Tile_X0Y1_EE4END({\Tile_X9Y12_EE4BEG[15] ,
    \Tile_X9Y12_EE4BEG[14] ,
    \Tile_X9Y12_EE4BEG[13] ,
    \Tile_X9Y12_EE4BEG[12] ,
    \Tile_X9Y12_EE4BEG[11] ,
    \Tile_X9Y12_EE4BEG[10] ,
    \Tile_X9Y12_EE4BEG[9] ,
    \Tile_X9Y12_EE4BEG[8] ,
    \Tile_X9Y12_EE4BEG[7] ,
    \Tile_X9Y12_EE4BEG[6] ,
    \Tile_X9Y12_EE4BEG[5] ,
    \Tile_X9Y12_EE4BEG[4] ,
    \Tile_X9Y12_EE4BEG[3] ,
    \Tile_X9Y12_EE4BEG[2] ,
    \Tile_X9Y12_EE4BEG[1] ,
    \Tile_X9Y12_EE4BEG[0] }),
    .Tile_X0Y1_FrameData({\Tile_X9Y12_FrameData_O[31] ,
    \Tile_X9Y12_FrameData_O[30] ,
    \Tile_X9Y12_FrameData_O[29] ,
    \Tile_X9Y12_FrameData_O[28] ,
    \Tile_X9Y12_FrameData_O[27] ,
    \Tile_X9Y12_FrameData_O[26] ,
    \Tile_X9Y12_FrameData_O[25] ,
    \Tile_X9Y12_FrameData_O[24] ,
    \Tile_X9Y12_FrameData_O[23] ,
    \Tile_X9Y12_FrameData_O[22] ,
    \Tile_X9Y12_FrameData_O[21] ,
    \Tile_X9Y12_FrameData_O[20] ,
    \Tile_X9Y12_FrameData_O[19] ,
    \Tile_X9Y12_FrameData_O[18] ,
    \Tile_X9Y12_FrameData_O[17] ,
    \Tile_X9Y12_FrameData_O[16] ,
    \Tile_X9Y12_FrameData_O[15] ,
    \Tile_X9Y12_FrameData_O[14] ,
    \Tile_X9Y12_FrameData_O[13] ,
    \Tile_X9Y12_FrameData_O[12] ,
    \Tile_X9Y12_FrameData_O[11] ,
    \Tile_X9Y12_FrameData_O[10] ,
    \Tile_X9Y12_FrameData_O[9] ,
    \Tile_X9Y12_FrameData_O[8] ,
    \Tile_X9Y12_FrameData_O[7] ,
    \Tile_X9Y12_FrameData_O[6] ,
    \Tile_X9Y12_FrameData_O[5] ,
    \Tile_X9Y12_FrameData_O[4] ,
    \Tile_X9Y12_FrameData_O[3] ,
    \Tile_X9Y12_FrameData_O[2] ,
    \Tile_X9Y12_FrameData_O[1] ,
    \Tile_X9Y12_FrameData_O[0] }),
    .Tile_X0Y1_FrameData_O({\Tile_X10Y12_FrameData_O[31] ,
    \Tile_X10Y12_FrameData_O[30] ,
    \Tile_X10Y12_FrameData_O[29] ,
    \Tile_X10Y12_FrameData_O[28] ,
    \Tile_X10Y12_FrameData_O[27] ,
    \Tile_X10Y12_FrameData_O[26] ,
    \Tile_X10Y12_FrameData_O[25] ,
    \Tile_X10Y12_FrameData_O[24] ,
    \Tile_X10Y12_FrameData_O[23] ,
    \Tile_X10Y12_FrameData_O[22] ,
    \Tile_X10Y12_FrameData_O[21] ,
    \Tile_X10Y12_FrameData_O[20] ,
    \Tile_X10Y12_FrameData_O[19] ,
    \Tile_X10Y12_FrameData_O[18] ,
    \Tile_X10Y12_FrameData_O[17] ,
    \Tile_X10Y12_FrameData_O[16] ,
    \Tile_X10Y12_FrameData_O[15] ,
    \Tile_X10Y12_FrameData_O[14] ,
    \Tile_X10Y12_FrameData_O[13] ,
    \Tile_X10Y12_FrameData_O[12] ,
    \Tile_X10Y12_FrameData_O[11] ,
    \Tile_X10Y12_FrameData_O[10] ,
    \Tile_X10Y12_FrameData_O[9] ,
    \Tile_X10Y12_FrameData_O[8] ,
    \Tile_X10Y12_FrameData_O[7] ,
    \Tile_X10Y12_FrameData_O[6] ,
    \Tile_X10Y12_FrameData_O[5] ,
    \Tile_X10Y12_FrameData_O[4] ,
    \Tile_X10Y12_FrameData_O[3] ,
    \Tile_X10Y12_FrameData_O[2] ,
    \Tile_X10Y12_FrameData_O[1] ,
    \Tile_X10Y12_FrameData_O[0] }),
    .Tile_X0Y1_FrameStrobe({\Tile_X10Y13_FrameStrobe_O[19] ,
    \Tile_X10Y13_FrameStrobe_O[18] ,
    \Tile_X10Y13_FrameStrobe_O[17] ,
    \Tile_X10Y13_FrameStrobe_O[16] ,
    \Tile_X10Y13_FrameStrobe_O[15] ,
    \Tile_X10Y13_FrameStrobe_O[14] ,
    \Tile_X10Y13_FrameStrobe_O[13] ,
    \Tile_X10Y13_FrameStrobe_O[12] ,
    \Tile_X10Y13_FrameStrobe_O[11] ,
    \Tile_X10Y13_FrameStrobe_O[10] ,
    \Tile_X10Y13_FrameStrobe_O[9] ,
    \Tile_X10Y13_FrameStrobe_O[8] ,
    \Tile_X10Y13_FrameStrobe_O[7] ,
    \Tile_X10Y13_FrameStrobe_O[6] ,
    \Tile_X10Y13_FrameStrobe_O[5] ,
    \Tile_X10Y13_FrameStrobe_O[4] ,
    \Tile_X10Y13_FrameStrobe_O[3] ,
    \Tile_X10Y13_FrameStrobe_O[2] ,
    \Tile_X10Y13_FrameStrobe_O[1] ,
    \Tile_X10Y13_FrameStrobe_O[0] }),
    .Tile_X0Y1_N1END({\Tile_X10Y13_N1BEG[3] ,
    \Tile_X10Y13_N1BEG[2] ,
    \Tile_X10Y13_N1BEG[1] ,
    \Tile_X10Y13_N1BEG[0] }),
    .Tile_X0Y1_N2END({\Tile_X10Y13_N2BEGb[7] ,
    \Tile_X10Y13_N2BEGb[6] ,
    \Tile_X10Y13_N2BEGb[5] ,
    \Tile_X10Y13_N2BEGb[4] ,
    \Tile_X10Y13_N2BEGb[3] ,
    \Tile_X10Y13_N2BEGb[2] ,
    \Tile_X10Y13_N2BEGb[1] ,
    \Tile_X10Y13_N2BEGb[0] }),
    .Tile_X0Y1_N2MID({\Tile_X10Y13_N2BEG[7] ,
    \Tile_X10Y13_N2BEG[6] ,
    \Tile_X10Y13_N2BEG[5] ,
    \Tile_X10Y13_N2BEG[4] ,
    \Tile_X10Y13_N2BEG[3] ,
    \Tile_X10Y13_N2BEG[2] ,
    \Tile_X10Y13_N2BEG[1] ,
    \Tile_X10Y13_N2BEG[0] }),
    .Tile_X0Y1_N4END({\Tile_X10Y13_N4BEG[15] ,
    \Tile_X10Y13_N4BEG[14] ,
    \Tile_X10Y13_N4BEG[13] ,
    \Tile_X10Y13_N4BEG[12] ,
    \Tile_X10Y13_N4BEG[11] ,
    \Tile_X10Y13_N4BEG[10] ,
    \Tile_X10Y13_N4BEG[9] ,
    \Tile_X10Y13_N4BEG[8] ,
    \Tile_X10Y13_N4BEG[7] ,
    \Tile_X10Y13_N4BEG[6] ,
    \Tile_X10Y13_N4BEG[5] ,
    \Tile_X10Y13_N4BEG[4] ,
    \Tile_X10Y13_N4BEG[3] ,
    \Tile_X10Y13_N4BEG[2] ,
    \Tile_X10Y13_N4BEG[1] ,
    \Tile_X10Y13_N4BEG[0] }),
    .Tile_X0Y1_S1BEG({\Tile_X10Y12_S1BEG[3] ,
    \Tile_X10Y12_S1BEG[2] ,
    \Tile_X10Y12_S1BEG[1] ,
    \Tile_X10Y12_S1BEG[0] }),
    .Tile_X0Y1_S2BEG({\Tile_X10Y12_S2BEG[7] ,
    \Tile_X10Y12_S2BEG[6] ,
    \Tile_X10Y12_S2BEG[5] ,
    \Tile_X10Y12_S2BEG[4] ,
    \Tile_X10Y12_S2BEG[3] ,
    \Tile_X10Y12_S2BEG[2] ,
    \Tile_X10Y12_S2BEG[1] ,
    \Tile_X10Y12_S2BEG[0] }),
    .Tile_X0Y1_S2BEGb({\Tile_X10Y12_S2BEGb[7] ,
    \Tile_X10Y12_S2BEGb[6] ,
    \Tile_X10Y12_S2BEGb[5] ,
    \Tile_X10Y12_S2BEGb[4] ,
    \Tile_X10Y12_S2BEGb[3] ,
    \Tile_X10Y12_S2BEGb[2] ,
    \Tile_X10Y12_S2BEGb[1] ,
    \Tile_X10Y12_S2BEGb[0] }),
    .Tile_X0Y1_S4BEG({\Tile_X10Y12_S4BEG[15] ,
    \Tile_X10Y12_S4BEG[14] ,
    \Tile_X10Y12_S4BEG[13] ,
    \Tile_X10Y12_S4BEG[12] ,
    \Tile_X10Y12_S4BEG[11] ,
    \Tile_X10Y12_S4BEG[10] ,
    \Tile_X10Y12_S4BEG[9] ,
    \Tile_X10Y12_S4BEG[8] ,
    \Tile_X10Y12_S4BEG[7] ,
    \Tile_X10Y12_S4BEG[6] ,
    \Tile_X10Y12_S4BEG[5] ,
    \Tile_X10Y12_S4BEG[4] ,
    \Tile_X10Y12_S4BEG[3] ,
    \Tile_X10Y12_S4BEG[2] ,
    \Tile_X10Y12_S4BEG[1] ,
    \Tile_X10Y12_S4BEG[0] }),
    .Tile_X0Y1_W1BEG({\Tile_X10Y12_W1BEG[3] ,
    \Tile_X10Y12_W1BEG[2] ,
    \Tile_X10Y12_W1BEG[1] ,
    \Tile_X10Y12_W1BEG[0] }),
    .Tile_X0Y1_W2BEG({\Tile_X10Y12_W2BEG[7] ,
    \Tile_X10Y12_W2BEG[6] ,
    \Tile_X10Y12_W2BEG[5] ,
    \Tile_X10Y12_W2BEG[4] ,
    \Tile_X10Y12_W2BEG[3] ,
    \Tile_X10Y12_W2BEG[2] ,
    \Tile_X10Y12_W2BEG[1] ,
    \Tile_X10Y12_W2BEG[0] }),
    .Tile_X0Y1_W2BEGb({\Tile_X10Y12_W2BEGb[7] ,
    \Tile_X10Y12_W2BEGb[6] ,
    \Tile_X10Y12_W2BEGb[5] ,
    \Tile_X10Y12_W2BEGb[4] ,
    \Tile_X10Y12_W2BEGb[3] ,
    \Tile_X10Y12_W2BEGb[2] ,
    \Tile_X10Y12_W2BEGb[1] ,
    \Tile_X10Y12_W2BEGb[0] }),
    .Tile_X0Y1_W6BEG({\Tile_X10Y12_W6BEG[11] ,
    \Tile_X10Y12_W6BEG[10] ,
    \Tile_X10Y12_W6BEG[9] ,
    \Tile_X10Y12_W6BEG[8] ,
    \Tile_X10Y12_W6BEG[7] ,
    \Tile_X10Y12_W6BEG[6] ,
    \Tile_X10Y12_W6BEG[5] ,
    \Tile_X10Y12_W6BEG[4] ,
    \Tile_X10Y12_W6BEG[3] ,
    \Tile_X10Y12_W6BEG[2] ,
    \Tile_X10Y12_W6BEG[1] ,
    \Tile_X10Y12_W6BEG[0] }),
    .Tile_X0Y1_WW4BEG({\Tile_X10Y12_WW4BEG[15] ,
    \Tile_X10Y12_WW4BEG[14] ,
    \Tile_X10Y12_WW4BEG[13] ,
    \Tile_X10Y12_WW4BEG[12] ,
    \Tile_X10Y12_WW4BEG[11] ,
    \Tile_X10Y12_WW4BEG[10] ,
    \Tile_X10Y12_WW4BEG[9] ,
    \Tile_X10Y12_WW4BEG[8] ,
    \Tile_X10Y12_WW4BEG[7] ,
    \Tile_X10Y12_WW4BEG[6] ,
    \Tile_X10Y12_WW4BEG[5] ,
    \Tile_X10Y12_WW4BEG[4] ,
    \Tile_X10Y12_WW4BEG[3] ,
    \Tile_X10Y12_WW4BEG[2] ,
    \Tile_X10Y12_WW4BEG[1] ,
    \Tile_X10Y12_WW4BEG[0] }));
 IHP_SRAM Tile_X10Y13_IHP_SRAM (.ADDR_SRAM0(Tile_X10Y14_ADDR_SRAM0),
    .ADDR_SRAM1(Tile_X10Y14_ADDR_SRAM1),
    .ADDR_SRAM2(Tile_X10Y14_ADDR_SRAM2),
    .ADDR_SRAM3(Tile_X10Y14_ADDR_SRAM3),
    .ADDR_SRAM4(Tile_X10Y14_ADDR_SRAM4),
    .ADDR_SRAM5(Tile_X10Y14_ADDR_SRAM5),
    .ADDR_SRAM6(Tile_X10Y14_ADDR_SRAM6),
    .ADDR_SRAM7(Tile_X10Y14_ADDR_SRAM7),
    .ADDR_SRAM8(Tile_X10Y14_ADDR_SRAM8),
    .ADDR_SRAM9(Tile_X10Y14_ADDR_SRAM9),
    .BM_SRAM0(Tile_X10Y14_BM_SRAM0),
    .BM_SRAM1(Tile_X10Y14_BM_SRAM1),
    .BM_SRAM10(Tile_X10Y14_BM_SRAM10),
    .BM_SRAM11(Tile_X10Y14_BM_SRAM11),
    .BM_SRAM12(Tile_X10Y14_BM_SRAM12),
    .BM_SRAM13(Tile_X10Y14_BM_SRAM13),
    .BM_SRAM14(Tile_X10Y14_BM_SRAM14),
    .BM_SRAM15(Tile_X10Y14_BM_SRAM15),
    .BM_SRAM16(Tile_X10Y14_BM_SRAM16),
    .BM_SRAM17(Tile_X10Y14_BM_SRAM17),
    .BM_SRAM18(Tile_X10Y14_BM_SRAM18),
    .BM_SRAM19(Tile_X10Y14_BM_SRAM19),
    .BM_SRAM2(Tile_X10Y14_BM_SRAM2),
    .BM_SRAM20(Tile_X10Y14_BM_SRAM20),
    .BM_SRAM21(Tile_X10Y14_BM_SRAM21),
    .BM_SRAM22(Tile_X10Y14_BM_SRAM22),
    .BM_SRAM23(Tile_X10Y14_BM_SRAM23),
    .BM_SRAM24(Tile_X10Y14_BM_SRAM24),
    .BM_SRAM25(Tile_X10Y14_BM_SRAM25),
    .BM_SRAM26(Tile_X10Y14_BM_SRAM26),
    .BM_SRAM27(Tile_X10Y14_BM_SRAM27),
    .BM_SRAM28(Tile_X10Y14_BM_SRAM28),
    .BM_SRAM29(Tile_X10Y14_BM_SRAM29),
    .BM_SRAM3(Tile_X10Y14_BM_SRAM3),
    .BM_SRAM30(Tile_X10Y14_BM_SRAM30),
    .BM_SRAM31(Tile_X10Y14_BM_SRAM31),
    .BM_SRAM4(Tile_X10Y14_BM_SRAM4),
    .BM_SRAM5(Tile_X10Y14_BM_SRAM5),
    .BM_SRAM6(Tile_X10Y14_BM_SRAM6),
    .BM_SRAM7(Tile_X10Y14_BM_SRAM7),
    .BM_SRAM8(Tile_X10Y14_BM_SRAM8),
    .BM_SRAM9(Tile_X10Y14_BM_SRAM9),
    .CLK_SRAM(Tile_X10Y14_CLK_SRAM),
    .CONFIGURED_top(Tile_X10Y14_CONFIGURED_top),
    .DIN_SRAM0(Tile_X10Y14_DIN_SRAM0),
    .DIN_SRAM1(Tile_X10Y14_DIN_SRAM1),
    .DIN_SRAM10(Tile_X10Y14_DIN_SRAM10),
    .DIN_SRAM11(Tile_X10Y14_DIN_SRAM11),
    .DIN_SRAM12(Tile_X10Y14_DIN_SRAM12),
    .DIN_SRAM13(Tile_X10Y14_DIN_SRAM13),
    .DIN_SRAM14(Tile_X10Y14_DIN_SRAM14),
    .DIN_SRAM15(Tile_X10Y14_DIN_SRAM15),
    .DIN_SRAM16(Tile_X10Y14_DIN_SRAM16),
    .DIN_SRAM17(Tile_X10Y14_DIN_SRAM17),
    .DIN_SRAM18(Tile_X10Y14_DIN_SRAM18),
    .DIN_SRAM19(Tile_X10Y14_DIN_SRAM19),
    .DIN_SRAM2(Tile_X10Y14_DIN_SRAM2),
    .DIN_SRAM20(Tile_X10Y14_DIN_SRAM20),
    .DIN_SRAM21(Tile_X10Y14_DIN_SRAM21),
    .DIN_SRAM22(Tile_X10Y14_DIN_SRAM22),
    .DIN_SRAM23(Tile_X10Y14_DIN_SRAM23),
    .DIN_SRAM24(Tile_X10Y14_DIN_SRAM24),
    .DIN_SRAM25(Tile_X10Y14_DIN_SRAM25),
    .DIN_SRAM26(Tile_X10Y14_DIN_SRAM26),
    .DIN_SRAM27(Tile_X10Y14_DIN_SRAM27),
    .DIN_SRAM28(Tile_X10Y14_DIN_SRAM28),
    .DIN_SRAM29(Tile_X10Y14_DIN_SRAM29),
    .DIN_SRAM3(Tile_X10Y14_DIN_SRAM3),
    .DIN_SRAM30(Tile_X10Y14_DIN_SRAM30),
    .DIN_SRAM31(Tile_X10Y14_DIN_SRAM31),
    .DIN_SRAM4(Tile_X10Y14_DIN_SRAM4),
    .DIN_SRAM5(Tile_X10Y14_DIN_SRAM5),
    .DIN_SRAM6(Tile_X10Y14_DIN_SRAM6),
    .DIN_SRAM7(Tile_X10Y14_DIN_SRAM7),
    .DIN_SRAM8(Tile_X10Y14_DIN_SRAM8),
    .DIN_SRAM9(Tile_X10Y14_DIN_SRAM9),
    .DOUT_SRAM0(Tile_X10Y14_DOUT_SRAM0),
    .DOUT_SRAM1(Tile_X10Y14_DOUT_SRAM1),
    .DOUT_SRAM10(Tile_X10Y14_DOUT_SRAM10),
    .DOUT_SRAM11(Tile_X10Y14_DOUT_SRAM11),
    .DOUT_SRAM12(Tile_X10Y14_DOUT_SRAM12),
    .DOUT_SRAM13(Tile_X10Y14_DOUT_SRAM13),
    .DOUT_SRAM14(Tile_X10Y14_DOUT_SRAM14),
    .DOUT_SRAM15(Tile_X10Y14_DOUT_SRAM15),
    .DOUT_SRAM16(Tile_X10Y14_DOUT_SRAM16),
    .DOUT_SRAM17(Tile_X10Y14_DOUT_SRAM17),
    .DOUT_SRAM18(Tile_X10Y14_DOUT_SRAM18),
    .DOUT_SRAM19(Tile_X10Y14_DOUT_SRAM19),
    .DOUT_SRAM2(Tile_X10Y14_DOUT_SRAM2),
    .DOUT_SRAM20(Tile_X10Y14_DOUT_SRAM20),
    .DOUT_SRAM21(Tile_X10Y14_DOUT_SRAM21),
    .DOUT_SRAM22(Tile_X10Y14_DOUT_SRAM22),
    .DOUT_SRAM23(Tile_X10Y14_DOUT_SRAM23),
    .DOUT_SRAM24(Tile_X10Y14_DOUT_SRAM24),
    .DOUT_SRAM25(Tile_X10Y14_DOUT_SRAM25),
    .DOUT_SRAM26(Tile_X10Y14_DOUT_SRAM26),
    .DOUT_SRAM27(Tile_X10Y14_DOUT_SRAM27),
    .DOUT_SRAM28(Tile_X10Y14_DOUT_SRAM28),
    .DOUT_SRAM29(Tile_X10Y14_DOUT_SRAM29),
    .DOUT_SRAM3(Tile_X10Y14_DOUT_SRAM3),
    .DOUT_SRAM30(Tile_X10Y14_DOUT_SRAM30),
    .DOUT_SRAM31(Tile_X10Y14_DOUT_SRAM31),
    .DOUT_SRAM4(Tile_X10Y14_DOUT_SRAM4),
    .DOUT_SRAM5(Tile_X10Y14_DOUT_SRAM5),
    .DOUT_SRAM6(Tile_X10Y14_DOUT_SRAM6),
    .DOUT_SRAM7(Tile_X10Y14_DOUT_SRAM7),
    .DOUT_SRAM8(Tile_X10Y14_DOUT_SRAM8),
    .DOUT_SRAM9(Tile_X10Y14_DOUT_SRAM9),
    .MEN_SRAM(Tile_X10Y14_MEN_SRAM),
    .REN_SRAM(Tile_X10Y14_REN_SRAM),
    .TIE_HIGH_SRAM(Tile_X10Y14_TIE_HIGH_SRAM),
    .TIE_LOW_SRAM(Tile_X10Y14_TIE_LOW_SRAM),
    .Tile_X0Y0_UserCLKo(Tile_X10Y13_UserCLKo),
    .Tile_X0Y1_UserCLK(Tile_X10Y15_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .WEN_SRAM(Tile_X10Y14_WEN_SRAM),
    .Tile_X0Y0_E1END({\Tile_X9Y13_E1BEG[3] ,
    \Tile_X9Y13_E1BEG[2] ,
    \Tile_X9Y13_E1BEG[1] ,
    \Tile_X9Y13_E1BEG[0] }),
    .Tile_X0Y0_E2END({\Tile_X9Y13_E2BEGb[7] ,
    \Tile_X9Y13_E2BEGb[6] ,
    \Tile_X9Y13_E2BEGb[5] ,
    \Tile_X9Y13_E2BEGb[4] ,
    \Tile_X9Y13_E2BEGb[3] ,
    \Tile_X9Y13_E2BEGb[2] ,
    \Tile_X9Y13_E2BEGb[1] ,
    \Tile_X9Y13_E2BEGb[0] }),
    .Tile_X0Y0_E2MID({\Tile_X9Y13_E2BEG[7] ,
    \Tile_X9Y13_E2BEG[6] ,
    \Tile_X9Y13_E2BEG[5] ,
    \Tile_X9Y13_E2BEG[4] ,
    \Tile_X9Y13_E2BEG[3] ,
    \Tile_X9Y13_E2BEG[2] ,
    \Tile_X9Y13_E2BEG[1] ,
    \Tile_X9Y13_E2BEG[0] }),
    .Tile_X0Y0_E6END({\Tile_X9Y13_E6BEG[11] ,
    \Tile_X9Y13_E6BEG[10] ,
    \Tile_X9Y13_E6BEG[9] ,
    \Tile_X9Y13_E6BEG[8] ,
    \Tile_X9Y13_E6BEG[7] ,
    \Tile_X9Y13_E6BEG[6] ,
    \Tile_X9Y13_E6BEG[5] ,
    \Tile_X9Y13_E6BEG[4] ,
    \Tile_X9Y13_E6BEG[3] ,
    \Tile_X9Y13_E6BEG[2] ,
    \Tile_X9Y13_E6BEG[1] ,
    \Tile_X9Y13_E6BEG[0] }),
    .Tile_X0Y0_EE4END({\Tile_X9Y13_EE4BEG[15] ,
    \Tile_X9Y13_EE4BEG[14] ,
    \Tile_X9Y13_EE4BEG[13] ,
    \Tile_X9Y13_EE4BEG[12] ,
    \Tile_X9Y13_EE4BEG[11] ,
    \Tile_X9Y13_EE4BEG[10] ,
    \Tile_X9Y13_EE4BEG[9] ,
    \Tile_X9Y13_EE4BEG[8] ,
    \Tile_X9Y13_EE4BEG[7] ,
    \Tile_X9Y13_EE4BEG[6] ,
    \Tile_X9Y13_EE4BEG[5] ,
    \Tile_X9Y13_EE4BEG[4] ,
    \Tile_X9Y13_EE4BEG[3] ,
    \Tile_X9Y13_EE4BEG[2] ,
    \Tile_X9Y13_EE4BEG[1] ,
    \Tile_X9Y13_EE4BEG[0] }),
    .Tile_X0Y0_FrameData({\Tile_X9Y13_FrameData_O[31] ,
    \Tile_X9Y13_FrameData_O[30] ,
    \Tile_X9Y13_FrameData_O[29] ,
    \Tile_X9Y13_FrameData_O[28] ,
    \Tile_X9Y13_FrameData_O[27] ,
    \Tile_X9Y13_FrameData_O[26] ,
    \Tile_X9Y13_FrameData_O[25] ,
    \Tile_X9Y13_FrameData_O[24] ,
    \Tile_X9Y13_FrameData_O[23] ,
    \Tile_X9Y13_FrameData_O[22] ,
    \Tile_X9Y13_FrameData_O[21] ,
    \Tile_X9Y13_FrameData_O[20] ,
    \Tile_X9Y13_FrameData_O[19] ,
    \Tile_X9Y13_FrameData_O[18] ,
    \Tile_X9Y13_FrameData_O[17] ,
    \Tile_X9Y13_FrameData_O[16] ,
    \Tile_X9Y13_FrameData_O[15] ,
    \Tile_X9Y13_FrameData_O[14] ,
    \Tile_X9Y13_FrameData_O[13] ,
    \Tile_X9Y13_FrameData_O[12] ,
    \Tile_X9Y13_FrameData_O[11] ,
    \Tile_X9Y13_FrameData_O[10] ,
    \Tile_X9Y13_FrameData_O[9] ,
    \Tile_X9Y13_FrameData_O[8] ,
    \Tile_X9Y13_FrameData_O[7] ,
    \Tile_X9Y13_FrameData_O[6] ,
    \Tile_X9Y13_FrameData_O[5] ,
    \Tile_X9Y13_FrameData_O[4] ,
    \Tile_X9Y13_FrameData_O[3] ,
    \Tile_X9Y13_FrameData_O[2] ,
    \Tile_X9Y13_FrameData_O[1] ,
    \Tile_X9Y13_FrameData_O[0] }),
    .Tile_X0Y0_FrameData_O({\Tile_X10Y13_FrameData_O[31] ,
    \Tile_X10Y13_FrameData_O[30] ,
    \Tile_X10Y13_FrameData_O[29] ,
    \Tile_X10Y13_FrameData_O[28] ,
    \Tile_X10Y13_FrameData_O[27] ,
    \Tile_X10Y13_FrameData_O[26] ,
    \Tile_X10Y13_FrameData_O[25] ,
    \Tile_X10Y13_FrameData_O[24] ,
    \Tile_X10Y13_FrameData_O[23] ,
    \Tile_X10Y13_FrameData_O[22] ,
    \Tile_X10Y13_FrameData_O[21] ,
    \Tile_X10Y13_FrameData_O[20] ,
    \Tile_X10Y13_FrameData_O[19] ,
    \Tile_X10Y13_FrameData_O[18] ,
    \Tile_X10Y13_FrameData_O[17] ,
    \Tile_X10Y13_FrameData_O[16] ,
    \Tile_X10Y13_FrameData_O[15] ,
    \Tile_X10Y13_FrameData_O[14] ,
    \Tile_X10Y13_FrameData_O[13] ,
    \Tile_X10Y13_FrameData_O[12] ,
    \Tile_X10Y13_FrameData_O[11] ,
    \Tile_X10Y13_FrameData_O[10] ,
    \Tile_X10Y13_FrameData_O[9] ,
    \Tile_X10Y13_FrameData_O[8] ,
    \Tile_X10Y13_FrameData_O[7] ,
    \Tile_X10Y13_FrameData_O[6] ,
    \Tile_X10Y13_FrameData_O[5] ,
    \Tile_X10Y13_FrameData_O[4] ,
    \Tile_X10Y13_FrameData_O[3] ,
    \Tile_X10Y13_FrameData_O[2] ,
    \Tile_X10Y13_FrameData_O[1] ,
    \Tile_X10Y13_FrameData_O[0] }),
    .Tile_X0Y0_FrameStrobe_O({\Tile_X10Y13_FrameStrobe_O[19] ,
    \Tile_X10Y13_FrameStrobe_O[18] ,
    \Tile_X10Y13_FrameStrobe_O[17] ,
    \Tile_X10Y13_FrameStrobe_O[16] ,
    \Tile_X10Y13_FrameStrobe_O[15] ,
    \Tile_X10Y13_FrameStrobe_O[14] ,
    \Tile_X10Y13_FrameStrobe_O[13] ,
    \Tile_X10Y13_FrameStrobe_O[12] ,
    \Tile_X10Y13_FrameStrobe_O[11] ,
    \Tile_X10Y13_FrameStrobe_O[10] ,
    \Tile_X10Y13_FrameStrobe_O[9] ,
    \Tile_X10Y13_FrameStrobe_O[8] ,
    \Tile_X10Y13_FrameStrobe_O[7] ,
    \Tile_X10Y13_FrameStrobe_O[6] ,
    \Tile_X10Y13_FrameStrobe_O[5] ,
    \Tile_X10Y13_FrameStrobe_O[4] ,
    \Tile_X10Y13_FrameStrobe_O[3] ,
    \Tile_X10Y13_FrameStrobe_O[2] ,
    \Tile_X10Y13_FrameStrobe_O[1] ,
    \Tile_X10Y13_FrameStrobe_O[0] }),
    .Tile_X0Y0_N1BEG({\Tile_X10Y13_N1BEG[3] ,
    \Tile_X10Y13_N1BEG[2] ,
    \Tile_X10Y13_N1BEG[1] ,
    \Tile_X10Y13_N1BEG[0] }),
    .Tile_X0Y0_N2BEG({\Tile_X10Y13_N2BEG[7] ,
    \Tile_X10Y13_N2BEG[6] ,
    \Tile_X10Y13_N2BEG[5] ,
    \Tile_X10Y13_N2BEG[4] ,
    \Tile_X10Y13_N2BEG[3] ,
    \Tile_X10Y13_N2BEG[2] ,
    \Tile_X10Y13_N2BEG[1] ,
    \Tile_X10Y13_N2BEG[0] }),
    .Tile_X0Y0_N2BEGb({\Tile_X10Y13_N2BEGb[7] ,
    \Tile_X10Y13_N2BEGb[6] ,
    \Tile_X10Y13_N2BEGb[5] ,
    \Tile_X10Y13_N2BEGb[4] ,
    \Tile_X10Y13_N2BEGb[3] ,
    \Tile_X10Y13_N2BEGb[2] ,
    \Tile_X10Y13_N2BEGb[1] ,
    \Tile_X10Y13_N2BEGb[0] }),
    .Tile_X0Y0_N4BEG({\Tile_X10Y13_N4BEG[15] ,
    \Tile_X10Y13_N4BEG[14] ,
    \Tile_X10Y13_N4BEG[13] ,
    \Tile_X10Y13_N4BEG[12] ,
    \Tile_X10Y13_N4BEG[11] ,
    \Tile_X10Y13_N4BEG[10] ,
    \Tile_X10Y13_N4BEG[9] ,
    \Tile_X10Y13_N4BEG[8] ,
    \Tile_X10Y13_N4BEG[7] ,
    \Tile_X10Y13_N4BEG[6] ,
    \Tile_X10Y13_N4BEG[5] ,
    \Tile_X10Y13_N4BEG[4] ,
    \Tile_X10Y13_N4BEG[3] ,
    \Tile_X10Y13_N4BEG[2] ,
    \Tile_X10Y13_N4BEG[1] ,
    \Tile_X10Y13_N4BEG[0] }),
    .Tile_X0Y0_S1END({\Tile_X10Y12_S1BEG[3] ,
    \Tile_X10Y12_S1BEG[2] ,
    \Tile_X10Y12_S1BEG[1] ,
    \Tile_X10Y12_S1BEG[0] }),
    .Tile_X0Y0_S2END({\Tile_X10Y12_S2BEGb[7] ,
    \Tile_X10Y12_S2BEGb[6] ,
    \Tile_X10Y12_S2BEGb[5] ,
    \Tile_X10Y12_S2BEGb[4] ,
    \Tile_X10Y12_S2BEGb[3] ,
    \Tile_X10Y12_S2BEGb[2] ,
    \Tile_X10Y12_S2BEGb[1] ,
    \Tile_X10Y12_S2BEGb[0] }),
    .Tile_X0Y0_S2MID({\Tile_X10Y12_S2BEG[7] ,
    \Tile_X10Y12_S2BEG[6] ,
    \Tile_X10Y12_S2BEG[5] ,
    \Tile_X10Y12_S2BEG[4] ,
    \Tile_X10Y12_S2BEG[3] ,
    \Tile_X10Y12_S2BEG[2] ,
    \Tile_X10Y12_S2BEG[1] ,
    \Tile_X10Y12_S2BEG[0] }),
    .Tile_X0Y0_S4END({\Tile_X10Y12_S4BEG[15] ,
    \Tile_X10Y12_S4BEG[14] ,
    \Tile_X10Y12_S4BEG[13] ,
    \Tile_X10Y12_S4BEG[12] ,
    \Tile_X10Y12_S4BEG[11] ,
    \Tile_X10Y12_S4BEG[10] ,
    \Tile_X10Y12_S4BEG[9] ,
    \Tile_X10Y12_S4BEG[8] ,
    \Tile_X10Y12_S4BEG[7] ,
    \Tile_X10Y12_S4BEG[6] ,
    \Tile_X10Y12_S4BEG[5] ,
    \Tile_X10Y12_S4BEG[4] ,
    \Tile_X10Y12_S4BEG[3] ,
    \Tile_X10Y12_S4BEG[2] ,
    \Tile_X10Y12_S4BEG[1] ,
    \Tile_X10Y12_S4BEG[0] }),
    .Tile_X0Y0_W1BEG({\Tile_X10Y13_W1BEG[3] ,
    \Tile_X10Y13_W1BEG[2] ,
    \Tile_X10Y13_W1BEG[1] ,
    \Tile_X10Y13_W1BEG[0] }),
    .Tile_X0Y0_W2BEG({\Tile_X10Y13_W2BEG[7] ,
    \Tile_X10Y13_W2BEG[6] ,
    \Tile_X10Y13_W2BEG[5] ,
    \Tile_X10Y13_W2BEG[4] ,
    \Tile_X10Y13_W2BEG[3] ,
    \Tile_X10Y13_W2BEG[2] ,
    \Tile_X10Y13_W2BEG[1] ,
    \Tile_X10Y13_W2BEG[0] }),
    .Tile_X0Y0_W2BEGb({\Tile_X10Y13_W2BEGb[7] ,
    \Tile_X10Y13_W2BEGb[6] ,
    \Tile_X10Y13_W2BEGb[5] ,
    \Tile_X10Y13_W2BEGb[4] ,
    \Tile_X10Y13_W2BEGb[3] ,
    \Tile_X10Y13_W2BEGb[2] ,
    \Tile_X10Y13_W2BEGb[1] ,
    \Tile_X10Y13_W2BEGb[0] }),
    .Tile_X0Y0_W6BEG({\Tile_X10Y13_W6BEG[11] ,
    \Tile_X10Y13_W6BEG[10] ,
    \Tile_X10Y13_W6BEG[9] ,
    \Tile_X10Y13_W6BEG[8] ,
    \Tile_X10Y13_W6BEG[7] ,
    \Tile_X10Y13_W6BEG[6] ,
    \Tile_X10Y13_W6BEG[5] ,
    \Tile_X10Y13_W6BEG[4] ,
    \Tile_X10Y13_W6BEG[3] ,
    \Tile_X10Y13_W6BEG[2] ,
    \Tile_X10Y13_W6BEG[1] ,
    \Tile_X10Y13_W6BEG[0] }),
    .Tile_X0Y0_WW4BEG({\Tile_X10Y13_WW4BEG[15] ,
    \Tile_X10Y13_WW4BEG[14] ,
    \Tile_X10Y13_WW4BEG[13] ,
    \Tile_X10Y13_WW4BEG[12] ,
    \Tile_X10Y13_WW4BEG[11] ,
    \Tile_X10Y13_WW4BEG[10] ,
    \Tile_X10Y13_WW4BEG[9] ,
    \Tile_X10Y13_WW4BEG[8] ,
    \Tile_X10Y13_WW4BEG[7] ,
    \Tile_X10Y13_WW4BEG[6] ,
    \Tile_X10Y13_WW4BEG[5] ,
    \Tile_X10Y13_WW4BEG[4] ,
    \Tile_X10Y13_WW4BEG[3] ,
    \Tile_X10Y13_WW4BEG[2] ,
    \Tile_X10Y13_WW4BEG[1] ,
    \Tile_X10Y13_WW4BEG[0] }),
    .Tile_X0Y1_E1END({\Tile_X9Y14_E1BEG[3] ,
    \Tile_X9Y14_E1BEG[2] ,
    \Tile_X9Y14_E1BEG[1] ,
    \Tile_X9Y14_E1BEG[0] }),
    .Tile_X0Y1_E2END({\Tile_X9Y14_E2BEGb[7] ,
    \Tile_X9Y14_E2BEGb[6] ,
    \Tile_X9Y14_E2BEGb[5] ,
    \Tile_X9Y14_E2BEGb[4] ,
    \Tile_X9Y14_E2BEGb[3] ,
    \Tile_X9Y14_E2BEGb[2] ,
    \Tile_X9Y14_E2BEGb[1] ,
    \Tile_X9Y14_E2BEGb[0] }),
    .Tile_X0Y1_E2MID({\Tile_X9Y14_E2BEG[7] ,
    \Tile_X9Y14_E2BEG[6] ,
    \Tile_X9Y14_E2BEG[5] ,
    \Tile_X9Y14_E2BEG[4] ,
    \Tile_X9Y14_E2BEG[3] ,
    \Tile_X9Y14_E2BEG[2] ,
    \Tile_X9Y14_E2BEG[1] ,
    \Tile_X9Y14_E2BEG[0] }),
    .Tile_X0Y1_E6END({\Tile_X9Y14_E6BEG[11] ,
    \Tile_X9Y14_E6BEG[10] ,
    \Tile_X9Y14_E6BEG[9] ,
    \Tile_X9Y14_E6BEG[8] ,
    \Tile_X9Y14_E6BEG[7] ,
    \Tile_X9Y14_E6BEG[6] ,
    \Tile_X9Y14_E6BEG[5] ,
    \Tile_X9Y14_E6BEG[4] ,
    \Tile_X9Y14_E6BEG[3] ,
    \Tile_X9Y14_E6BEG[2] ,
    \Tile_X9Y14_E6BEG[1] ,
    \Tile_X9Y14_E6BEG[0] }),
    .Tile_X0Y1_EE4END({\Tile_X9Y14_EE4BEG[15] ,
    \Tile_X9Y14_EE4BEG[14] ,
    \Tile_X9Y14_EE4BEG[13] ,
    \Tile_X9Y14_EE4BEG[12] ,
    \Tile_X9Y14_EE4BEG[11] ,
    \Tile_X9Y14_EE4BEG[10] ,
    \Tile_X9Y14_EE4BEG[9] ,
    \Tile_X9Y14_EE4BEG[8] ,
    \Tile_X9Y14_EE4BEG[7] ,
    \Tile_X9Y14_EE4BEG[6] ,
    \Tile_X9Y14_EE4BEG[5] ,
    \Tile_X9Y14_EE4BEG[4] ,
    \Tile_X9Y14_EE4BEG[3] ,
    \Tile_X9Y14_EE4BEG[2] ,
    \Tile_X9Y14_EE4BEG[1] ,
    \Tile_X9Y14_EE4BEG[0] }),
    .Tile_X0Y1_FrameData({\Tile_X9Y14_FrameData_O[31] ,
    \Tile_X9Y14_FrameData_O[30] ,
    \Tile_X9Y14_FrameData_O[29] ,
    \Tile_X9Y14_FrameData_O[28] ,
    \Tile_X9Y14_FrameData_O[27] ,
    \Tile_X9Y14_FrameData_O[26] ,
    \Tile_X9Y14_FrameData_O[25] ,
    \Tile_X9Y14_FrameData_O[24] ,
    \Tile_X9Y14_FrameData_O[23] ,
    \Tile_X9Y14_FrameData_O[22] ,
    \Tile_X9Y14_FrameData_O[21] ,
    \Tile_X9Y14_FrameData_O[20] ,
    \Tile_X9Y14_FrameData_O[19] ,
    \Tile_X9Y14_FrameData_O[18] ,
    \Tile_X9Y14_FrameData_O[17] ,
    \Tile_X9Y14_FrameData_O[16] ,
    \Tile_X9Y14_FrameData_O[15] ,
    \Tile_X9Y14_FrameData_O[14] ,
    \Tile_X9Y14_FrameData_O[13] ,
    \Tile_X9Y14_FrameData_O[12] ,
    \Tile_X9Y14_FrameData_O[11] ,
    \Tile_X9Y14_FrameData_O[10] ,
    \Tile_X9Y14_FrameData_O[9] ,
    \Tile_X9Y14_FrameData_O[8] ,
    \Tile_X9Y14_FrameData_O[7] ,
    \Tile_X9Y14_FrameData_O[6] ,
    \Tile_X9Y14_FrameData_O[5] ,
    \Tile_X9Y14_FrameData_O[4] ,
    \Tile_X9Y14_FrameData_O[3] ,
    \Tile_X9Y14_FrameData_O[2] ,
    \Tile_X9Y14_FrameData_O[1] ,
    \Tile_X9Y14_FrameData_O[0] }),
    .Tile_X0Y1_FrameData_O({\Tile_X10Y14_FrameData_O[31] ,
    \Tile_X10Y14_FrameData_O[30] ,
    \Tile_X10Y14_FrameData_O[29] ,
    \Tile_X10Y14_FrameData_O[28] ,
    \Tile_X10Y14_FrameData_O[27] ,
    \Tile_X10Y14_FrameData_O[26] ,
    \Tile_X10Y14_FrameData_O[25] ,
    \Tile_X10Y14_FrameData_O[24] ,
    \Tile_X10Y14_FrameData_O[23] ,
    \Tile_X10Y14_FrameData_O[22] ,
    \Tile_X10Y14_FrameData_O[21] ,
    \Tile_X10Y14_FrameData_O[20] ,
    \Tile_X10Y14_FrameData_O[19] ,
    \Tile_X10Y14_FrameData_O[18] ,
    \Tile_X10Y14_FrameData_O[17] ,
    \Tile_X10Y14_FrameData_O[16] ,
    \Tile_X10Y14_FrameData_O[15] ,
    \Tile_X10Y14_FrameData_O[14] ,
    \Tile_X10Y14_FrameData_O[13] ,
    \Tile_X10Y14_FrameData_O[12] ,
    \Tile_X10Y14_FrameData_O[11] ,
    \Tile_X10Y14_FrameData_O[10] ,
    \Tile_X10Y14_FrameData_O[9] ,
    \Tile_X10Y14_FrameData_O[8] ,
    \Tile_X10Y14_FrameData_O[7] ,
    \Tile_X10Y14_FrameData_O[6] ,
    \Tile_X10Y14_FrameData_O[5] ,
    \Tile_X10Y14_FrameData_O[4] ,
    \Tile_X10Y14_FrameData_O[3] ,
    \Tile_X10Y14_FrameData_O[2] ,
    \Tile_X10Y14_FrameData_O[1] ,
    \Tile_X10Y14_FrameData_O[0] }),
    .Tile_X0Y1_FrameStrobe({\Tile_X10Y15_FrameStrobe_O[19] ,
    \Tile_X10Y15_FrameStrobe_O[18] ,
    \Tile_X10Y15_FrameStrobe_O[17] ,
    \Tile_X10Y15_FrameStrobe_O[16] ,
    \Tile_X10Y15_FrameStrobe_O[15] ,
    \Tile_X10Y15_FrameStrobe_O[14] ,
    \Tile_X10Y15_FrameStrobe_O[13] ,
    \Tile_X10Y15_FrameStrobe_O[12] ,
    \Tile_X10Y15_FrameStrobe_O[11] ,
    \Tile_X10Y15_FrameStrobe_O[10] ,
    \Tile_X10Y15_FrameStrobe_O[9] ,
    \Tile_X10Y15_FrameStrobe_O[8] ,
    \Tile_X10Y15_FrameStrobe_O[7] ,
    \Tile_X10Y15_FrameStrobe_O[6] ,
    \Tile_X10Y15_FrameStrobe_O[5] ,
    \Tile_X10Y15_FrameStrobe_O[4] ,
    \Tile_X10Y15_FrameStrobe_O[3] ,
    \Tile_X10Y15_FrameStrobe_O[2] ,
    \Tile_X10Y15_FrameStrobe_O[1] ,
    \Tile_X10Y15_FrameStrobe_O[0] }),
    .Tile_X0Y1_N1END({\Tile_X10Y15_N1BEG[3] ,
    \Tile_X10Y15_N1BEG[2] ,
    \Tile_X10Y15_N1BEG[1] ,
    \Tile_X10Y15_N1BEG[0] }),
    .Tile_X0Y1_N2END({\Tile_X10Y15_N2BEGb[7] ,
    \Tile_X10Y15_N2BEGb[6] ,
    \Tile_X10Y15_N2BEGb[5] ,
    \Tile_X10Y15_N2BEGb[4] ,
    \Tile_X10Y15_N2BEGb[3] ,
    \Tile_X10Y15_N2BEGb[2] ,
    \Tile_X10Y15_N2BEGb[1] ,
    \Tile_X10Y15_N2BEGb[0] }),
    .Tile_X0Y1_N2MID({\Tile_X10Y15_N2BEG[7] ,
    \Tile_X10Y15_N2BEG[6] ,
    \Tile_X10Y15_N2BEG[5] ,
    \Tile_X10Y15_N2BEG[4] ,
    \Tile_X10Y15_N2BEG[3] ,
    \Tile_X10Y15_N2BEG[2] ,
    \Tile_X10Y15_N2BEG[1] ,
    \Tile_X10Y15_N2BEG[0] }),
    .Tile_X0Y1_N4END({\Tile_X10Y15_N4BEG[15] ,
    \Tile_X10Y15_N4BEG[14] ,
    \Tile_X10Y15_N4BEG[13] ,
    \Tile_X10Y15_N4BEG[12] ,
    \Tile_X10Y15_N4BEG[11] ,
    \Tile_X10Y15_N4BEG[10] ,
    \Tile_X10Y15_N4BEG[9] ,
    \Tile_X10Y15_N4BEG[8] ,
    \Tile_X10Y15_N4BEG[7] ,
    \Tile_X10Y15_N4BEG[6] ,
    \Tile_X10Y15_N4BEG[5] ,
    \Tile_X10Y15_N4BEG[4] ,
    \Tile_X10Y15_N4BEG[3] ,
    \Tile_X10Y15_N4BEG[2] ,
    \Tile_X10Y15_N4BEG[1] ,
    \Tile_X10Y15_N4BEG[0] }),
    .Tile_X0Y1_S1BEG({\Tile_X10Y14_S1BEG[3] ,
    \Tile_X10Y14_S1BEG[2] ,
    \Tile_X10Y14_S1BEG[1] ,
    \Tile_X10Y14_S1BEG[0] }),
    .Tile_X0Y1_S2BEG({\Tile_X10Y14_S2BEG[7] ,
    \Tile_X10Y14_S2BEG[6] ,
    \Tile_X10Y14_S2BEG[5] ,
    \Tile_X10Y14_S2BEG[4] ,
    \Tile_X10Y14_S2BEG[3] ,
    \Tile_X10Y14_S2BEG[2] ,
    \Tile_X10Y14_S2BEG[1] ,
    \Tile_X10Y14_S2BEG[0] }),
    .Tile_X0Y1_S2BEGb({\Tile_X10Y14_S2BEGb[7] ,
    \Tile_X10Y14_S2BEGb[6] ,
    \Tile_X10Y14_S2BEGb[5] ,
    \Tile_X10Y14_S2BEGb[4] ,
    \Tile_X10Y14_S2BEGb[3] ,
    \Tile_X10Y14_S2BEGb[2] ,
    \Tile_X10Y14_S2BEGb[1] ,
    \Tile_X10Y14_S2BEGb[0] }),
    .Tile_X0Y1_S4BEG({\Tile_X10Y14_S4BEG[15] ,
    \Tile_X10Y14_S4BEG[14] ,
    \Tile_X10Y14_S4BEG[13] ,
    \Tile_X10Y14_S4BEG[12] ,
    \Tile_X10Y14_S4BEG[11] ,
    \Tile_X10Y14_S4BEG[10] ,
    \Tile_X10Y14_S4BEG[9] ,
    \Tile_X10Y14_S4BEG[8] ,
    \Tile_X10Y14_S4BEG[7] ,
    \Tile_X10Y14_S4BEG[6] ,
    \Tile_X10Y14_S4BEG[5] ,
    \Tile_X10Y14_S4BEG[4] ,
    \Tile_X10Y14_S4BEG[3] ,
    \Tile_X10Y14_S4BEG[2] ,
    \Tile_X10Y14_S4BEG[1] ,
    \Tile_X10Y14_S4BEG[0] }),
    .Tile_X0Y1_W1BEG({\Tile_X10Y14_W1BEG[3] ,
    \Tile_X10Y14_W1BEG[2] ,
    \Tile_X10Y14_W1BEG[1] ,
    \Tile_X10Y14_W1BEG[0] }),
    .Tile_X0Y1_W2BEG({\Tile_X10Y14_W2BEG[7] ,
    \Tile_X10Y14_W2BEG[6] ,
    \Tile_X10Y14_W2BEG[5] ,
    \Tile_X10Y14_W2BEG[4] ,
    \Tile_X10Y14_W2BEG[3] ,
    \Tile_X10Y14_W2BEG[2] ,
    \Tile_X10Y14_W2BEG[1] ,
    \Tile_X10Y14_W2BEG[0] }),
    .Tile_X0Y1_W2BEGb({\Tile_X10Y14_W2BEGb[7] ,
    \Tile_X10Y14_W2BEGb[6] ,
    \Tile_X10Y14_W2BEGb[5] ,
    \Tile_X10Y14_W2BEGb[4] ,
    \Tile_X10Y14_W2BEGb[3] ,
    \Tile_X10Y14_W2BEGb[2] ,
    \Tile_X10Y14_W2BEGb[1] ,
    \Tile_X10Y14_W2BEGb[0] }),
    .Tile_X0Y1_W6BEG({\Tile_X10Y14_W6BEG[11] ,
    \Tile_X10Y14_W6BEG[10] ,
    \Tile_X10Y14_W6BEG[9] ,
    \Tile_X10Y14_W6BEG[8] ,
    \Tile_X10Y14_W6BEG[7] ,
    \Tile_X10Y14_W6BEG[6] ,
    \Tile_X10Y14_W6BEG[5] ,
    \Tile_X10Y14_W6BEG[4] ,
    \Tile_X10Y14_W6BEG[3] ,
    \Tile_X10Y14_W6BEG[2] ,
    \Tile_X10Y14_W6BEG[1] ,
    \Tile_X10Y14_W6BEG[0] }),
    .Tile_X0Y1_WW4BEG({\Tile_X10Y14_WW4BEG[15] ,
    \Tile_X10Y14_WW4BEG[14] ,
    \Tile_X10Y14_WW4BEG[13] ,
    \Tile_X10Y14_WW4BEG[12] ,
    \Tile_X10Y14_WW4BEG[11] ,
    \Tile_X10Y14_WW4BEG[10] ,
    \Tile_X10Y14_WW4BEG[9] ,
    \Tile_X10Y14_WW4BEG[8] ,
    \Tile_X10Y14_WW4BEG[7] ,
    \Tile_X10Y14_WW4BEG[6] ,
    \Tile_X10Y14_WW4BEG[5] ,
    \Tile_X10Y14_WW4BEG[4] ,
    \Tile_X10Y14_WW4BEG[3] ,
    \Tile_X10Y14_WW4BEG[2] ,
    \Tile_X10Y14_WW4BEG[1] ,
    \Tile_X10Y14_WW4BEG[0] }));
 S_term_IHP_SRAM Tile_X10Y15_S_term_IHP_SRAM (.UserCLK(UserCLK),
    .UserCLKo(Tile_X10Y15_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .FrameData({\Tile_X9Y15_FrameData_O[31] ,
    \Tile_X9Y15_FrameData_O[30] ,
    \Tile_X9Y15_FrameData_O[29] ,
    \Tile_X9Y15_FrameData_O[28] ,
    \Tile_X9Y15_FrameData_O[27] ,
    \Tile_X9Y15_FrameData_O[26] ,
    \Tile_X9Y15_FrameData_O[25] ,
    \Tile_X9Y15_FrameData_O[24] ,
    \Tile_X9Y15_FrameData_O[23] ,
    \Tile_X9Y15_FrameData_O[22] ,
    \Tile_X9Y15_FrameData_O[21] ,
    \Tile_X9Y15_FrameData_O[20] ,
    \Tile_X9Y15_FrameData_O[19] ,
    \Tile_X9Y15_FrameData_O[18] ,
    \Tile_X9Y15_FrameData_O[17] ,
    \Tile_X9Y15_FrameData_O[16] ,
    \Tile_X9Y15_FrameData_O[15] ,
    \Tile_X9Y15_FrameData_O[14] ,
    \Tile_X9Y15_FrameData_O[13] ,
    \Tile_X9Y15_FrameData_O[12] ,
    \Tile_X9Y15_FrameData_O[11] ,
    \Tile_X9Y15_FrameData_O[10] ,
    \Tile_X9Y15_FrameData_O[9] ,
    \Tile_X9Y15_FrameData_O[8] ,
    \Tile_X9Y15_FrameData_O[7] ,
    \Tile_X9Y15_FrameData_O[6] ,
    \Tile_X9Y15_FrameData_O[5] ,
    \Tile_X9Y15_FrameData_O[4] ,
    \Tile_X9Y15_FrameData_O[3] ,
    \Tile_X9Y15_FrameData_O[2] ,
    \Tile_X9Y15_FrameData_O[1] ,
    \Tile_X9Y15_FrameData_O[0] }),
    .FrameData_O({\Tile_X10Y15_FrameData_O[31] ,
    \Tile_X10Y15_FrameData_O[30] ,
    \Tile_X10Y15_FrameData_O[29] ,
    \Tile_X10Y15_FrameData_O[28] ,
    \Tile_X10Y15_FrameData_O[27] ,
    \Tile_X10Y15_FrameData_O[26] ,
    \Tile_X10Y15_FrameData_O[25] ,
    \Tile_X10Y15_FrameData_O[24] ,
    \Tile_X10Y15_FrameData_O[23] ,
    \Tile_X10Y15_FrameData_O[22] ,
    \Tile_X10Y15_FrameData_O[21] ,
    \Tile_X10Y15_FrameData_O[20] ,
    \Tile_X10Y15_FrameData_O[19] ,
    \Tile_X10Y15_FrameData_O[18] ,
    \Tile_X10Y15_FrameData_O[17] ,
    \Tile_X10Y15_FrameData_O[16] ,
    \Tile_X10Y15_FrameData_O[15] ,
    \Tile_X10Y15_FrameData_O[14] ,
    \Tile_X10Y15_FrameData_O[13] ,
    \Tile_X10Y15_FrameData_O[12] ,
    \Tile_X10Y15_FrameData_O[11] ,
    \Tile_X10Y15_FrameData_O[10] ,
    \Tile_X10Y15_FrameData_O[9] ,
    \Tile_X10Y15_FrameData_O[8] ,
    \Tile_X10Y15_FrameData_O[7] ,
    \Tile_X10Y15_FrameData_O[6] ,
    \Tile_X10Y15_FrameData_O[5] ,
    \Tile_X10Y15_FrameData_O[4] ,
    \Tile_X10Y15_FrameData_O[3] ,
    \Tile_X10Y15_FrameData_O[2] ,
    \Tile_X10Y15_FrameData_O[1] ,
    \Tile_X10Y15_FrameData_O[0] }),
    .FrameStrobe({FrameStrobe[219],
    FrameStrobe[218],
    FrameStrobe[217],
    FrameStrobe[216],
    FrameStrobe[215],
    FrameStrobe[214],
    FrameStrobe[213],
    FrameStrobe[212],
    FrameStrobe[211],
    FrameStrobe[210],
    FrameStrobe[209],
    FrameStrobe[208],
    FrameStrobe[207],
    FrameStrobe[206],
    FrameStrobe[205],
    FrameStrobe[204],
    FrameStrobe[203],
    FrameStrobe[202],
    FrameStrobe[201],
    FrameStrobe[200]}),
    .FrameStrobe_O({\Tile_X10Y15_FrameStrobe_O[19] ,
    \Tile_X10Y15_FrameStrobe_O[18] ,
    \Tile_X10Y15_FrameStrobe_O[17] ,
    \Tile_X10Y15_FrameStrobe_O[16] ,
    \Tile_X10Y15_FrameStrobe_O[15] ,
    \Tile_X10Y15_FrameStrobe_O[14] ,
    \Tile_X10Y15_FrameStrobe_O[13] ,
    \Tile_X10Y15_FrameStrobe_O[12] ,
    \Tile_X10Y15_FrameStrobe_O[11] ,
    \Tile_X10Y15_FrameStrobe_O[10] ,
    \Tile_X10Y15_FrameStrobe_O[9] ,
    \Tile_X10Y15_FrameStrobe_O[8] ,
    \Tile_X10Y15_FrameStrobe_O[7] ,
    \Tile_X10Y15_FrameStrobe_O[6] ,
    \Tile_X10Y15_FrameStrobe_O[5] ,
    \Tile_X10Y15_FrameStrobe_O[4] ,
    \Tile_X10Y15_FrameStrobe_O[3] ,
    \Tile_X10Y15_FrameStrobe_O[2] ,
    \Tile_X10Y15_FrameStrobe_O[1] ,
    \Tile_X10Y15_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X10Y15_N1BEG[3] ,
    \Tile_X10Y15_N1BEG[2] ,
    \Tile_X10Y15_N1BEG[1] ,
    \Tile_X10Y15_N1BEG[0] }),
    .N2BEG({\Tile_X10Y15_N2BEG[7] ,
    \Tile_X10Y15_N2BEG[6] ,
    \Tile_X10Y15_N2BEG[5] ,
    \Tile_X10Y15_N2BEG[4] ,
    \Tile_X10Y15_N2BEG[3] ,
    \Tile_X10Y15_N2BEG[2] ,
    \Tile_X10Y15_N2BEG[1] ,
    \Tile_X10Y15_N2BEG[0] }),
    .N2BEGb({\Tile_X10Y15_N2BEGb[7] ,
    \Tile_X10Y15_N2BEGb[6] ,
    \Tile_X10Y15_N2BEGb[5] ,
    \Tile_X10Y15_N2BEGb[4] ,
    \Tile_X10Y15_N2BEGb[3] ,
    \Tile_X10Y15_N2BEGb[2] ,
    \Tile_X10Y15_N2BEGb[1] ,
    \Tile_X10Y15_N2BEGb[0] }),
    .N4BEG({\Tile_X10Y15_N4BEG[15] ,
    \Tile_X10Y15_N4BEG[14] ,
    \Tile_X10Y15_N4BEG[13] ,
    \Tile_X10Y15_N4BEG[12] ,
    \Tile_X10Y15_N4BEG[11] ,
    \Tile_X10Y15_N4BEG[10] ,
    \Tile_X10Y15_N4BEG[9] ,
    \Tile_X10Y15_N4BEG[8] ,
    \Tile_X10Y15_N4BEG[7] ,
    \Tile_X10Y15_N4BEG[6] ,
    \Tile_X10Y15_N4BEG[5] ,
    \Tile_X10Y15_N4BEG[4] ,
    \Tile_X10Y15_N4BEG[3] ,
    \Tile_X10Y15_N4BEG[2] ,
    \Tile_X10Y15_N4BEG[1] ,
    \Tile_X10Y15_N4BEG[0] }),
    .S1END({\Tile_X10Y14_S1BEG[3] ,
    \Tile_X10Y14_S1BEG[2] ,
    \Tile_X10Y14_S1BEG[1] ,
    \Tile_X10Y14_S1BEG[0] }),
    .S2END({\Tile_X10Y14_S2BEGb[7] ,
    \Tile_X10Y14_S2BEGb[6] ,
    \Tile_X10Y14_S2BEGb[5] ,
    \Tile_X10Y14_S2BEGb[4] ,
    \Tile_X10Y14_S2BEGb[3] ,
    \Tile_X10Y14_S2BEGb[2] ,
    \Tile_X10Y14_S2BEGb[1] ,
    \Tile_X10Y14_S2BEGb[0] }),
    .S2MID({\Tile_X10Y14_S2BEG[7] ,
    \Tile_X10Y14_S2BEG[6] ,
    \Tile_X10Y14_S2BEG[5] ,
    \Tile_X10Y14_S2BEG[4] ,
    \Tile_X10Y14_S2BEG[3] ,
    \Tile_X10Y14_S2BEG[2] ,
    \Tile_X10Y14_S2BEG[1] ,
    \Tile_X10Y14_S2BEG[0] }),
    .S4END({\Tile_X10Y14_S4BEG[15] ,
    \Tile_X10Y14_S4BEG[14] ,
    \Tile_X10Y14_S4BEG[13] ,
    \Tile_X10Y14_S4BEG[12] ,
    \Tile_X10Y14_S4BEG[11] ,
    \Tile_X10Y14_S4BEG[10] ,
    \Tile_X10Y14_S4BEG[9] ,
    \Tile_X10Y14_S4BEG[8] ,
    \Tile_X10Y14_S4BEG[7] ,
    \Tile_X10Y14_S4BEG[6] ,
    \Tile_X10Y14_S4BEG[5] ,
    \Tile_X10Y14_S4BEG[4] ,
    \Tile_X10Y14_S4BEG[3] ,
    \Tile_X10Y14_S4BEG[2] ,
    \Tile_X10Y14_S4BEG[1] ,
    \Tile_X10Y14_S4BEG[0] }));
 IHP_SRAM Tile_X10Y1_IHP_SRAM (.ADDR_SRAM0(Tile_X10Y2_ADDR_SRAM0),
    .ADDR_SRAM1(Tile_X10Y2_ADDR_SRAM1),
    .ADDR_SRAM2(Tile_X10Y2_ADDR_SRAM2),
    .ADDR_SRAM3(Tile_X10Y2_ADDR_SRAM3),
    .ADDR_SRAM4(Tile_X10Y2_ADDR_SRAM4),
    .ADDR_SRAM5(Tile_X10Y2_ADDR_SRAM5),
    .ADDR_SRAM6(Tile_X10Y2_ADDR_SRAM6),
    .ADDR_SRAM7(Tile_X10Y2_ADDR_SRAM7),
    .ADDR_SRAM8(Tile_X10Y2_ADDR_SRAM8),
    .ADDR_SRAM9(Tile_X10Y2_ADDR_SRAM9),
    .BM_SRAM0(Tile_X10Y2_BM_SRAM0),
    .BM_SRAM1(Tile_X10Y2_BM_SRAM1),
    .BM_SRAM10(Tile_X10Y2_BM_SRAM10),
    .BM_SRAM11(Tile_X10Y2_BM_SRAM11),
    .BM_SRAM12(Tile_X10Y2_BM_SRAM12),
    .BM_SRAM13(Tile_X10Y2_BM_SRAM13),
    .BM_SRAM14(Tile_X10Y2_BM_SRAM14),
    .BM_SRAM15(Tile_X10Y2_BM_SRAM15),
    .BM_SRAM16(Tile_X10Y2_BM_SRAM16),
    .BM_SRAM17(Tile_X10Y2_BM_SRAM17),
    .BM_SRAM18(Tile_X10Y2_BM_SRAM18),
    .BM_SRAM19(Tile_X10Y2_BM_SRAM19),
    .BM_SRAM2(Tile_X10Y2_BM_SRAM2),
    .BM_SRAM20(Tile_X10Y2_BM_SRAM20),
    .BM_SRAM21(Tile_X10Y2_BM_SRAM21),
    .BM_SRAM22(Tile_X10Y2_BM_SRAM22),
    .BM_SRAM23(Tile_X10Y2_BM_SRAM23),
    .BM_SRAM24(Tile_X10Y2_BM_SRAM24),
    .BM_SRAM25(Tile_X10Y2_BM_SRAM25),
    .BM_SRAM26(Tile_X10Y2_BM_SRAM26),
    .BM_SRAM27(Tile_X10Y2_BM_SRAM27),
    .BM_SRAM28(Tile_X10Y2_BM_SRAM28),
    .BM_SRAM29(Tile_X10Y2_BM_SRAM29),
    .BM_SRAM3(Tile_X10Y2_BM_SRAM3),
    .BM_SRAM30(Tile_X10Y2_BM_SRAM30),
    .BM_SRAM31(Tile_X10Y2_BM_SRAM31),
    .BM_SRAM4(Tile_X10Y2_BM_SRAM4),
    .BM_SRAM5(Tile_X10Y2_BM_SRAM5),
    .BM_SRAM6(Tile_X10Y2_BM_SRAM6),
    .BM_SRAM7(Tile_X10Y2_BM_SRAM7),
    .BM_SRAM8(Tile_X10Y2_BM_SRAM8),
    .BM_SRAM9(Tile_X10Y2_BM_SRAM9),
    .CLK_SRAM(Tile_X10Y2_CLK_SRAM),
    .CONFIGURED_top(Tile_X10Y2_CONFIGURED_top),
    .DIN_SRAM0(Tile_X10Y2_DIN_SRAM0),
    .DIN_SRAM1(Tile_X10Y2_DIN_SRAM1),
    .DIN_SRAM10(Tile_X10Y2_DIN_SRAM10),
    .DIN_SRAM11(Tile_X10Y2_DIN_SRAM11),
    .DIN_SRAM12(Tile_X10Y2_DIN_SRAM12),
    .DIN_SRAM13(Tile_X10Y2_DIN_SRAM13),
    .DIN_SRAM14(Tile_X10Y2_DIN_SRAM14),
    .DIN_SRAM15(Tile_X10Y2_DIN_SRAM15),
    .DIN_SRAM16(Tile_X10Y2_DIN_SRAM16),
    .DIN_SRAM17(Tile_X10Y2_DIN_SRAM17),
    .DIN_SRAM18(Tile_X10Y2_DIN_SRAM18),
    .DIN_SRAM19(Tile_X10Y2_DIN_SRAM19),
    .DIN_SRAM2(Tile_X10Y2_DIN_SRAM2),
    .DIN_SRAM20(Tile_X10Y2_DIN_SRAM20),
    .DIN_SRAM21(Tile_X10Y2_DIN_SRAM21),
    .DIN_SRAM22(Tile_X10Y2_DIN_SRAM22),
    .DIN_SRAM23(Tile_X10Y2_DIN_SRAM23),
    .DIN_SRAM24(Tile_X10Y2_DIN_SRAM24),
    .DIN_SRAM25(Tile_X10Y2_DIN_SRAM25),
    .DIN_SRAM26(Tile_X10Y2_DIN_SRAM26),
    .DIN_SRAM27(Tile_X10Y2_DIN_SRAM27),
    .DIN_SRAM28(Tile_X10Y2_DIN_SRAM28),
    .DIN_SRAM29(Tile_X10Y2_DIN_SRAM29),
    .DIN_SRAM3(Tile_X10Y2_DIN_SRAM3),
    .DIN_SRAM30(Tile_X10Y2_DIN_SRAM30),
    .DIN_SRAM31(Tile_X10Y2_DIN_SRAM31),
    .DIN_SRAM4(Tile_X10Y2_DIN_SRAM4),
    .DIN_SRAM5(Tile_X10Y2_DIN_SRAM5),
    .DIN_SRAM6(Tile_X10Y2_DIN_SRAM6),
    .DIN_SRAM7(Tile_X10Y2_DIN_SRAM7),
    .DIN_SRAM8(Tile_X10Y2_DIN_SRAM8),
    .DIN_SRAM9(Tile_X10Y2_DIN_SRAM9),
    .DOUT_SRAM0(Tile_X10Y2_DOUT_SRAM0),
    .DOUT_SRAM1(Tile_X10Y2_DOUT_SRAM1),
    .DOUT_SRAM10(Tile_X10Y2_DOUT_SRAM10),
    .DOUT_SRAM11(Tile_X10Y2_DOUT_SRAM11),
    .DOUT_SRAM12(Tile_X10Y2_DOUT_SRAM12),
    .DOUT_SRAM13(Tile_X10Y2_DOUT_SRAM13),
    .DOUT_SRAM14(Tile_X10Y2_DOUT_SRAM14),
    .DOUT_SRAM15(Tile_X10Y2_DOUT_SRAM15),
    .DOUT_SRAM16(Tile_X10Y2_DOUT_SRAM16),
    .DOUT_SRAM17(Tile_X10Y2_DOUT_SRAM17),
    .DOUT_SRAM18(Tile_X10Y2_DOUT_SRAM18),
    .DOUT_SRAM19(Tile_X10Y2_DOUT_SRAM19),
    .DOUT_SRAM2(Tile_X10Y2_DOUT_SRAM2),
    .DOUT_SRAM20(Tile_X10Y2_DOUT_SRAM20),
    .DOUT_SRAM21(Tile_X10Y2_DOUT_SRAM21),
    .DOUT_SRAM22(Tile_X10Y2_DOUT_SRAM22),
    .DOUT_SRAM23(Tile_X10Y2_DOUT_SRAM23),
    .DOUT_SRAM24(Tile_X10Y2_DOUT_SRAM24),
    .DOUT_SRAM25(Tile_X10Y2_DOUT_SRAM25),
    .DOUT_SRAM26(Tile_X10Y2_DOUT_SRAM26),
    .DOUT_SRAM27(Tile_X10Y2_DOUT_SRAM27),
    .DOUT_SRAM28(Tile_X10Y2_DOUT_SRAM28),
    .DOUT_SRAM29(Tile_X10Y2_DOUT_SRAM29),
    .DOUT_SRAM3(Tile_X10Y2_DOUT_SRAM3),
    .DOUT_SRAM30(Tile_X10Y2_DOUT_SRAM30),
    .DOUT_SRAM31(Tile_X10Y2_DOUT_SRAM31),
    .DOUT_SRAM4(Tile_X10Y2_DOUT_SRAM4),
    .DOUT_SRAM5(Tile_X10Y2_DOUT_SRAM5),
    .DOUT_SRAM6(Tile_X10Y2_DOUT_SRAM6),
    .DOUT_SRAM7(Tile_X10Y2_DOUT_SRAM7),
    .DOUT_SRAM8(Tile_X10Y2_DOUT_SRAM8),
    .DOUT_SRAM9(Tile_X10Y2_DOUT_SRAM9),
    .MEN_SRAM(Tile_X10Y2_MEN_SRAM),
    .REN_SRAM(Tile_X10Y2_REN_SRAM),
    .TIE_HIGH_SRAM(Tile_X10Y2_TIE_HIGH_SRAM),
    .TIE_LOW_SRAM(Tile_X10Y2_TIE_LOW_SRAM),
    .Tile_X0Y0_UserCLKo(Tile_X10Y1_UserCLKo),
    .Tile_X0Y1_UserCLK(Tile_X10Y3_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .WEN_SRAM(Tile_X10Y2_WEN_SRAM),
    .Tile_X0Y0_E1END({\Tile_X9Y1_E1BEG[3] ,
    \Tile_X9Y1_E1BEG[2] ,
    \Tile_X9Y1_E1BEG[1] ,
    \Tile_X9Y1_E1BEG[0] }),
    .Tile_X0Y0_E2END({\Tile_X9Y1_E2BEGb[7] ,
    \Tile_X9Y1_E2BEGb[6] ,
    \Tile_X9Y1_E2BEGb[5] ,
    \Tile_X9Y1_E2BEGb[4] ,
    \Tile_X9Y1_E2BEGb[3] ,
    \Tile_X9Y1_E2BEGb[2] ,
    \Tile_X9Y1_E2BEGb[1] ,
    \Tile_X9Y1_E2BEGb[0] }),
    .Tile_X0Y0_E2MID({\Tile_X9Y1_E2BEG[7] ,
    \Tile_X9Y1_E2BEG[6] ,
    \Tile_X9Y1_E2BEG[5] ,
    \Tile_X9Y1_E2BEG[4] ,
    \Tile_X9Y1_E2BEG[3] ,
    \Tile_X9Y1_E2BEG[2] ,
    \Tile_X9Y1_E2BEG[1] ,
    \Tile_X9Y1_E2BEG[0] }),
    .Tile_X0Y0_E6END({\Tile_X9Y1_E6BEG[11] ,
    \Tile_X9Y1_E6BEG[10] ,
    \Tile_X9Y1_E6BEG[9] ,
    \Tile_X9Y1_E6BEG[8] ,
    \Tile_X9Y1_E6BEG[7] ,
    \Tile_X9Y1_E6BEG[6] ,
    \Tile_X9Y1_E6BEG[5] ,
    \Tile_X9Y1_E6BEG[4] ,
    \Tile_X9Y1_E6BEG[3] ,
    \Tile_X9Y1_E6BEG[2] ,
    \Tile_X9Y1_E6BEG[1] ,
    \Tile_X9Y1_E6BEG[0] }),
    .Tile_X0Y0_EE4END({\Tile_X9Y1_EE4BEG[15] ,
    \Tile_X9Y1_EE4BEG[14] ,
    \Tile_X9Y1_EE4BEG[13] ,
    \Tile_X9Y1_EE4BEG[12] ,
    \Tile_X9Y1_EE4BEG[11] ,
    \Tile_X9Y1_EE4BEG[10] ,
    \Tile_X9Y1_EE4BEG[9] ,
    \Tile_X9Y1_EE4BEG[8] ,
    \Tile_X9Y1_EE4BEG[7] ,
    \Tile_X9Y1_EE4BEG[6] ,
    \Tile_X9Y1_EE4BEG[5] ,
    \Tile_X9Y1_EE4BEG[4] ,
    \Tile_X9Y1_EE4BEG[3] ,
    \Tile_X9Y1_EE4BEG[2] ,
    \Tile_X9Y1_EE4BEG[1] ,
    \Tile_X9Y1_EE4BEG[0] }),
    .Tile_X0Y0_FrameData({\Tile_X9Y1_FrameData_O[31] ,
    \Tile_X9Y1_FrameData_O[30] ,
    \Tile_X9Y1_FrameData_O[29] ,
    \Tile_X9Y1_FrameData_O[28] ,
    \Tile_X9Y1_FrameData_O[27] ,
    \Tile_X9Y1_FrameData_O[26] ,
    \Tile_X9Y1_FrameData_O[25] ,
    \Tile_X9Y1_FrameData_O[24] ,
    \Tile_X9Y1_FrameData_O[23] ,
    \Tile_X9Y1_FrameData_O[22] ,
    \Tile_X9Y1_FrameData_O[21] ,
    \Tile_X9Y1_FrameData_O[20] ,
    \Tile_X9Y1_FrameData_O[19] ,
    \Tile_X9Y1_FrameData_O[18] ,
    \Tile_X9Y1_FrameData_O[17] ,
    \Tile_X9Y1_FrameData_O[16] ,
    \Tile_X9Y1_FrameData_O[15] ,
    \Tile_X9Y1_FrameData_O[14] ,
    \Tile_X9Y1_FrameData_O[13] ,
    \Tile_X9Y1_FrameData_O[12] ,
    \Tile_X9Y1_FrameData_O[11] ,
    \Tile_X9Y1_FrameData_O[10] ,
    \Tile_X9Y1_FrameData_O[9] ,
    \Tile_X9Y1_FrameData_O[8] ,
    \Tile_X9Y1_FrameData_O[7] ,
    \Tile_X9Y1_FrameData_O[6] ,
    \Tile_X9Y1_FrameData_O[5] ,
    \Tile_X9Y1_FrameData_O[4] ,
    \Tile_X9Y1_FrameData_O[3] ,
    \Tile_X9Y1_FrameData_O[2] ,
    \Tile_X9Y1_FrameData_O[1] ,
    \Tile_X9Y1_FrameData_O[0] }),
    .Tile_X0Y0_FrameData_O({\Tile_X10Y1_FrameData_O[31] ,
    \Tile_X10Y1_FrameData_O[30] ,
    \Tile_X10Y1_FrameData_O[29] ,
    \Tile_X10Y1_FrameData_O[28] ,
    \Tile_X10Y1_FrameData_O[27] ,
    \Tile_X10Y1_FrameData_O[26] ,
    \Tile_X10Y1_FrameData_O[25] ,
    \Tile_X10Y1_FrameData_O[24] ,
    \Tile_X10Y1_FrameData_O[23] ,
    \Tile_X10Y1_FrameData_O[22] ,
    \Tile_X10Y1_FrameData_O[21] ,
    \Tile_X10Y1_FrameData_O[20] ,
    \Tile_X10Y1_FrameData_O[19] ,
    \Tile_X10Y1_FrameData_O[18] ,
    \Tile_X10Y1_FrameData_O[17] ,
    \Tile_X10Y1_FrameData_O[16] ,
    \Tile_X10Y1_FrameData_O[15] ,
    \Tile_X10Y1_FrameData_O[14] ,
    \Tile_X10Y1_FrameData_O[13] ,
    \Tile_X10Y1_FrameData_O[12] ,
    \Tile_X10Y1_FrameData_O[11] ,
    \Tile_X10Y1_FrameData_O[10] ,
    \Tile_X10Y1_FrameData_O[9] ,
    \Tile_X10Y1_FrameData_O[8] ,
    \Tile_X10Y1_FrameData_O[7] ,
    \Tile_X10Y1_FrameData_O[6] ,
    \Tile_X10Y1_FrameData_O[5] ,
    \Tile_X10Y1_FrameData_O[4] ,
    \Tile_X10Y1_FrameData_O[3] ,
    \Tile_X10Y1_FrameData_O[2] ,
    \Tile_X10Y1_FrameData_O[1] ,
    \Tile_X10Y1_FrameData_O[0] }),
    .Tile_X0Y0_FrameStrobe_O({\Tile_X10Y1_FrameStrobe_O[19] ,
    \Tile_X10Y1_FrameStrobe_O[18] ,
    \Tile_X10Y1_FrameStrobe_O[17] ,
    \Tile_X10Y1_FrameStrobe_O[16] ,
    \Tile_X10Y1_FrameStrobe_O[15] ,
    \Tile_X10Y1_FrameStrobe_O[14] ,
    \Tile_X10Y1_FrameStrobe_O[13] ,
    \Tile_X10Y1_FrameStrobe_O[12] ,
    \Tile_X10Y1_FrameStrobe_O[11] ,
    \Tile_X10Y1_FrameStrobe_O[10] ,
    \Tile_X10Y1_FrameStrobe_O[9] ,
    \Tile_X10Y1_FrameStrobe_O[8] ,
    \Tile_X10Y1_FrameStrobe_O[7] ,
    \Tile_X10Y1_FrameStrobe_O[6] ,
    \Tile_X10Y1_FrameStrobe_O[5] ,
    \Tile_X10Y1_FrameStrobe_O[4] ,
    \Tile_X10Y1_FrameStrobe_O[3] ,
    \Tile_X10Y1_FrameStrobe_O[2] ,
    \Tile_X10Y1_FrameStrobe_O[1] ,
    \Tile_X10Y1_FrameStrobe_O[0] }),
    .Tile_X0Y0_N1BEG({\Tile_X10Y1_N1BEG[3] ,
    \Tile_X10Y1_N1BEG[2] ,
    \Tile_X10Y1_N1BEG[1] ,
    \Tile_X10Y1_N1BEG[0] }),
    .Tile_X0Y0_N2BEG({\Tile_X10Y1_N2BEG[7] ,
    \Tile_X10Y1_N2BEG[6] ,
    \Tile_X10Y1_N2BEG[5] ,
    \Tile_X10Y1_N2BEG[4] ,
    \Tile_X10Y1_N2BEG[3] ,
    \Tile_X10Y1_N2BEG[2] ,
    \Tile_X10Y1_N2BEG[1] ,
    \Tile_X10Y1_N2BEG[0] }),
    .Tile_X0Y0_N2BEGb({\Tile_X10Y1_N2BEGb[7] ,
    \Tile_X10Y1_N2BEGb[6] ,
    \Tile_X10Y1_N2BEGb[5] ,
    \Tile_X10Y1_N2BEGb[4] ,
    \Tile_X10Y1_N2BEGb[3] ,
    \Tile_X10Y1_N2BEGb[2] ,
    \Tile_X10Y1_N2BEGb[1] ,
    \Tile_X10Y1_N2BEGb[0] }),
    .Tile_X0Y0_N4BEG({\Tile_X10Y1_N4BEG[15] ,
    \Tile_X10Y1_N4BEG[14] ,
    \Tile_X10Y1_N4BEG[13] ,
    \Tile_X10Y1_N4BEG[12] ,
    \Tile_X10Y1_N4BEG[11] ,
    \Tile_X10Y1_N4BEG[10] ,
    \Tile_X10Y1_N4BEG[9] ,
    \Tile_X10Y1_N4BEG[8] ,
    \Tile_X10Y1_N4BEG[7] ,
    \Tile_X10Y1_N4BEG[6] ,
    \Tile_X10Y1_N4BEG[5] ,
    \Tile_X10Y1_N4BEG[4] ,
    \Tile_X10Y1_N4BEG[3] ,
    \Tile_X10Y1_N4BEG[2] ,
    \Tile_X10Y1_N4BEG[1] ,
    \Tile_X10Y1_N4BEG[0] }),
    .Tile_X0Y0_S1END({\Tile_X10Y0_S1BEG[3] ,
    \Tile_X10Y0_S1BEG[2] ,
    \Tile_X10Y0_S1BEG[1] ,
    \Tile_X10Y0_S1BEG[0] }),
    .Tile_X0Y0_S2END({\Tile_X10Y0_S2BEGb[7] ,
    \Tile_X10Y0_S2BEGb[6] ,
    \Tile_X10Y0_S2BEGb[5] ,
    \Tile_X10Y0_S2BEGb[4] ,
    \Tile_X10Y0_S2BEGb[3] ,
    \Tile_X10Y0_S2BEGb[2] ,
    \Tile_X10Y0_S2BEGb[1] ,
    \Tile_X10Y0_S2BEGb[0] }),
    .Tile_X0Y0_S2MID({\Tile_X10Y0_S2BEG[7] ,
    \Tile_X10Y0_S2BEG[6] ,
    \Tile_X10Y0_S2BEG[5] ,
    \Tile_X10Y0_S2BEG[4] ,
    \Tile_X10Y0_S2BEG[3] ,
    \Tile_X10Y0_S2BEG[2] ,
    \Tile_X10Y0_S2BEG[1] ,
    \Tile_X10Y0_S2BEG[0] }),
    .Tile_X0Y0_S4END({\Tile_X10Y0_S4BEG[15] ,
    \Tile_X10Y0_S4BEG[14] ,
    \Tile_X10Y0_S4BEG[13] ,
    \Tile_X10Y0_S4BEG[12] ,
    \Tile_X10Y0_S4BEG[11] ,
    \Tile_X10Y0_S4BEG[10] ,
    \Tile_X10Y0_S4BEG[9] ,
    \Tile_X10Y0_S4BEG[8] ,
    \Tile_X10Y0_S4BEG[7] ,
    \Tile_X10Y0_S4BEG[6] ,
    \Tile_X10Y0_S4BEG[5] ,
    \Tile_X10Y0_S4BEG[4] ,
    \Tile_X10Y0_S4BEG[3] ,
    \Tile_X10Y0_S4BEG[2] ,
    \Tile_X10Y0_S4BEG[1] ,
    \Tile_X10Y0_S4BEG[0] }),
    .Tile_X0Y0_W1BEG({\Tile_X10Y1_W1BEG[3] ,
    \Tile_X10Y1_W1BEG[2] ,
    \Tile_X10Y1_W1BEG[1] ,
    \Tile_X10Y1_W1BEG[0] }),
    .Tile_X0Y0_W2BEG({\Tile_X10Y1_W2BEG[7] ,
    \Tile_X10Y1_W2BEG[6] ,
    \Tile_X10Y1_W2BEG[5] ,
    \Tile_X10Y1_W2BEG[4] ,
    \Tile_X10Y1_W2BEG[3] ,
    \Tile_X10Y1_W2BEG[2] ,
    \Tile_X10Y1_W2BEG[1] ,
    \Tile_X10Y1_W2BEG[0] }),
    .Tile_X0Y0_W2BEGb({\Tile_X10Y1_W2BEGb[7] ,
    \Tile_X10Y1_W2BEGb[6] ,
    \Tile_X10Y1_W2BEGb[5] ,
    \Tile_X10Y1_W2BEGb[4] ,
    \Tile_X10Y1_W2BEGb[3] ,
    \Tile_X10Y1_W2BEGb[2] ,
    \Tile_X10Y1_W2BEGb[1] ,
    \Tile_X10Y1_W2BEGb[0] }),
    .Tile_X0Y0_W6BEG({\Tile_X10Y1_W6BEG[11] ,
    \Tile_X10Y1_W6BEG[10] ,
    \Tile_X10Y1_W6BEG[9] ,
    \Tile_X10Y1_W6BEG[8] ,
    \Tile_X10Y1_W6BEG[7] ,
    \Tile_X10Y1_W6BEG[6] ,
    \Tile_X10Y1_W6BEG[5] ,
    \Tile_X10Y1_W6BEG[4] ,
    \Tile_X10Y1_W6BEG[3] ,
    \Tile_X10Y1_W6BEG[2] ,
    \Tile_X10Y1_W6BEG[1] ,
    \Tile_X10Y1_W6BEG[0] }),
    .Tile_X0Y0_WW4BEG({\Tile_X10Y1_WW4BEG[15] ,
    \Tile_X10Y1_WW4BEG[14] ,
    \Tile_X10Y1_WW4BEG[13] ,
    \Tile_X10Y1_WW4BEG[12] ,
    \Tile_X10Y1_WW4BEG[11] ,
    \Tile_X10Y1_WW4BEG[10] ,
    \Tile_X10Y1_WW4BEG[9] ,
    \Tile_X10Y1_WW4BEG[8] ,
    \Tile_X10Y1_WW4BEG[7] ,
    \Tile_X10Y1_WW4BEG[6] ,
    \Tile_X10Y1_WW4BEG[5] ,
    \Tile_X10Y1_WW4BEG[4] ,
    \Tile_X10Y1_WW4BEG[3] ,
    \Tile_X10Y1_WW4BEG[2] ,
    \Tile_X10Y1_WW4BEG[1] ,
    \Tile_X10Y1_WW4BEG[0] }),
    .Tile_X0Y1_E1END({\Tile_X9Y2_E1BEG[3] ,
    \Tile_X9Y2_E1BEG[2] ,
    \Tile_X9Y2_E1BEG[1] ,
    \Tile_X9Y2_E1BEG[0] }),
    .Tile_X0Y1_E2END({\Tile_X9Y2_E2BEGb[7] ,
    \Tile_X9Y2_E2BEGb[6] ,
    \Tile_X9Y2_E2BEGb[5] ,
    \Tile_X9Y2_E2BEGb[4] ,
    \Tile_X9Y2_E2BEGb[3] ,
    \Tile_X9Y2_E2BEGb[2] ,
    \Tile_X9Y2_E2BEGb[1] ,
    \Tile_X9Y2_E2BEGb[0] }),
    .Tile_X0Y1_E2MID({\Tile_X9Y2_E2BEG[7] ,
    \Tile_X9Y2_E2BEG[6] ,
    \Tile_X9Y2_E2BEG[5] ,
    \Tile_X9Y2_E2BEG[4] ,
    \Tile_X9Y2_E2BEG[3] ,
    \Tile_X9Y2_E2BEG[2] ,
    \Tile_X9Y2_E2BEG[1] ,
    \Tile_X9Y2_E2BEG[0] }),
    .Tile_X0Y1_E6END({\Tile_X9Y2_E6BEG[11] ,
    \Tile_X9Y2_E6BEG[10] ,
    \Tile_X9Y2_E6BEG[9] ,
    \Tile_X9Y2_E6BEG[8] ,
    \Tile_X9Y2_E6BEG[7] ,
    \Tile_X9Y2_E6BEG[6] ,
    \Tile_X9Y2_E6BEG[5] ,
    \Tile_X9Y2_E6BEG[4] ,
    \Tile_X9Y2_E6BEG[3] ,
    \Tile_X9Y2_E6BEG[2] ,
    \Tile_X9Y2_E6BEG[1] ,
    \Tile_X9Y2_E6BEG[0] }),
    .Tile_X0Y1_EE4END({\Tile_X9Y2_EE4BEG[15] ,
    \Tile_X9Y2_EE4BEG[14] ,
    \Tile_X9Y2_EE4BEG[13] ,
    \Tile_X9Y2_EE4BEG[12] ,
    \Tile_X9Y2_EE4BEG[11] ,
    \Tile_X9Y2_EE4BEG[10] ,
    \Tile_X9Y2_EE4BEG[9] ,
    \Tile_X9Y2_EE4BEG[8] ,
    \Tile_X9Y2_EE4BEG[7] ,
    \Tile_X9Y2_EE4BEG[6] ,
    \Tile_X9Y2_EE4BEG[5] ,
    \Tile_X9Y2_EE4BEG[4] ,
    \Tile_X9Y2_EE4BEG[3] ,
    \Tile_X9Y2_EE4BEG[2] ,
    \Tile_X9Y2_EE4BEG[1] ,
    \Tile_X9Y2_EE4BEG[0] }),
    .Tile_X0Y1_FrameData({\Tile_X9Y2_FrameData_O[31] ,
    \Tile_X9Y2_FrameData_O[30] ,
    \Tile_X9Y2_FrameData_O[29] ,
    \Tile_X9Y2_FrameData_O[28] ,
    \Tile_X9Y2_FrameData_O[27] ,
    \Tile_X9Y2_FrameData_O[26] ,
    \Tile_X9Y2_FrameData_O[25] ,
    \Tile_X9Y2_FrameData_O[24] ,
    \Tile_X9Y2_FrameData_O[23] ,
    \Tile_X9Y2_FrameData_O[22] ,
    \Tile_X9Y2_FrameData_O[21] ,
    \Tile_X9Y2_FrameData_O[20] ,
    \Tile_X9Y2_FrameData_O[19] ,
    \Tile_X9Y2_FrameData_O[18] ,
    \Tile_X9Y2_FrameData_O[17] ,
    \Tile_X9Y2_FrameData_O[16] ,
    \Tile_X9Y2_FrameData_O[15] ,
    \Tile_X9Y2_FrameData_O[14] ,
    \Tile_X9Y2_FrameData_O[13] ,
    \Tile_X9Y2_FrameData_O[12] ,
    \Tile_X9Y2_FrameData_O[11] ,
    \Tile_X9Y2_FrameData_O[10] ,
    \Tile_X9Y2_FrameData_O[9] ,
    \Tile_X9Y2_FrameData_O[8] ,
    \Tile_X9Y2_FrameData_O[7] ,
    \Tile_X9Y2_FrameData_O[6] ,
    \Tile_X9Y2_FrameData_O[5] ,
    \Tile_X9Y2_FrameData_O[4] ,
    \Tile_X9Y2_FrameData_O[3] ,
    \Tile_X9Y2_FrameData_O[2] ,
    \Tile_X9Y2_FrameData_O[1] ,
    \Tile_X9Y2_FrameData_O[0] }),
    .Tile_X0Y1_FrameData_O({\Tile_X10Y2_FrameData_O[31] ,
    \Tile_X10Y2_FrameData_O[30] ,
    \Tile_X10Y2_FrameData_O[29] ,
    \Tile_X10Y2_FrameData_O[28] ,
    \Tile_X10Y2_FrameData_O[27] ,
    \Tile_X10Y2_FrameData_O[26] ,
    \Tile_X10Y2_FrameData_O[25] ,
    \Tile_X10Y2_FrameData_O[24] ,
    \Tile_X10Y2_FrameData_O[23] ,
    \Tile_X10Y2_FrameData_O[22] ,
    \Tile_X10Y2_FrameData_O[21] ,
    \Tile_X10Y2_FrameData_O[20] ,
    \Tile_X10Y2_FrameData_O[19] ,
    \Tile_X10Y2_FrameData_O[18] ,
    \Tile_X10Y2_FrameData_O[17] ,
    \Tile_X10Y2_FrameData_O[16] ,
    \Tile_X10Y2_FrameData_O[15] ,
    \Tile_X10Y2_FrameData_O[14] ,
    \Tile_X10Y2_FrameData_O[13] ,
    \Tile_X10Y2_FrameData_O[12] ,
    \Tile_X10Y2_FrameData_O[11] ,
    \Tile_X10Y2_FrameData_O[10] ,
    \Tile_X10Y2_FrameData_O[9] ,
    \Tile_X10Y2_FrameData_O[8] ,
    \Tile_X10Y2_FrameData_O[7] ,
    \Tile_X10Y2_FrameData_O[6] ,
    \Tile_X10Y2_FrameData_O[5] ,
    \Tile_X10Y2_FrameData_O[4] ,
    \Tile_X10Y2_FrameData_O[3] ,
    \Tile_X10Y2_FrameData_O[2] ,
    \Tile_X10Y2_FrameData_O[1] ,
    \Tile_X10Y2_FrameData_O[0] }),
    .Tile_X0Y1_FrameStrobe({\Tile_X10Y3_FrameStrobe_O[19] ,
    \Tile_X10Y3_FrameStrobe_O[18] ,
    \Tile_X10Y3_FrameStrobe_O[17] ,
    \Tile_X10Y3_FrameStrobe_O[16] ,
    \Tile_X10Y3_FrameStrobe_O[15] ,
    \Tile_X10Y3_FrameStrobe_O[14] ,
    \Tile_X10Y3_FrameStrobe_O[13] ,
    \Tile_X10Y3_FrameStrobe_O[12] ,
    \Tile_X10Y3_FrameStrobe_O[11] ,
    \Tile_X10Y3_FrameStrobe_O[10] ,
    \Tile_X10Y3_FrameStrobe_O[9] ,
    \Tile_X10Y3_FrameStrobe_O[8] ,
    \Tile_X10Y3_FrameStrobe_O[7] ,
    \Tile_X10Y3_FrameStrobe_O[6] ,
    \Tile_X10Y3_FrameStrobe_O[5] ,
    \Tile_X10Y3_FrameStrobe_O[4] ,
    \Tile_X10Y3_FrameStrobe_O[3] ,
    \Tile_X10Y3_FrameStrobe_O[2] ,
    \Tile_X10Y3_FrameStrobe_O[1] ,
    \Tile_X10Y3_FrameStrobe_O[0] }),
    .Tile_X0Y1_N1END({\Tile_X10Y3_N1BEG[3] ,
    \Tile_X10Y3_N1BEG[2] ,
    \Tile_X10Y3_N1BEG[1] ,
    \Tile_X10Y3_N1BEG[0] }),
    .Tile_X0Y1_N2END({\Tile_X10Y3_N2BEGb[7] ,
    \Tile_X10Y3_N2BEGb[6] ,
    \Tile_X10Y3_N2BEGb[5] ,
    \Tile_X10Y3_N2BEGb[4] ,
    \Tile_X10Y3_N2BEGb[3] ,
    \Tile_X10Y3_N2BEGb[2] ,
    \Tile_X10Y3_N2BEGb[1] ,
    \Tile_X10Y3_N2BEGb[0] }),
    .Tile_X0Y1_N2MID({\Tile_X10Y3_N2BEG[7] ,
    \Tile_X10Y3_N2BEG[6] ,
    \Tile_X10Y3_N2BEG[5] ,
    \Tile_X10Y3_N2BEG[4] ,
    \Tile_X10Y3_N2BEG[3] ,
    \Tile_X10Y3_N2BEG[2] ,
    \Tile_X10Y3_N2BEG[1] ,
    \Tile_X10Y3_N2BEG[0] }),
    .Tile_X0Y1_N4END({\Tile_X10Y3_N4BEG[15] ,
    \Tile_X10Y3_N4BEG[14] ,
    \Tile_X10Y3_N4BEG[13] ,
    \Tile_X10Y3_N4BEG[12] ,
    \Tile_X10Y3_N4BEG[11] ,
    \Tile_X10Y3_N4BEG[10] ,
    \Tile_X10Y3_N4BEG[9] ,
    \Tile_X10Y3_N4BEG[8] ,
    \Tile_X10Y3_N4BEG[7] ,
    \Tile_X10Y3_N4BEG[6] ,
    \Tile_X10Y3_N4BEG[5] ,
    \Tile_X10Y3_N4BEG[4] ,
    \Tile_X10Y3_N4BEG[3] ,
    \Tile_X10Y3_N4BEG[2] ,
    \Tile_X10Y3_N4BEG[1] ,
    \Tile_X10Y3_N4BEG[0] }),
    .Tile_X0Y1_S1BEG({\Tile_X10Y2_S1BEG[3] ,
    \Tile_X10Y2_S1BEG[2] ,
    \Tile_X10Y2_S1BEG[1] ,
    \Tile_X10Y2_S1BEG[0] }),
    .Tile_X0Y1_S2BEG({\Tile_X10Y2_S2BEG[7] ,
    \Tile_X10Y2_S2BEG[6] ,
    \Tile_X10Y2_S2BEG[5] ,
    \Tile_X10Y2_S2BEG[4] ,
    \Tile_X10Y2_S2BEG[3] ,
    \Tile_X10Y2_S2BEG[2] ,
    \Tile_X10Y2_S2BEG[1] ,
    \Tile_X10Y2_S2BEG[0] }),
    .Tile_X0Y1_S2BEGb({\Tile_X10Y2_S2BEGb[7] ,
    \Tile_X10Y2_S2BEGb[6] ,
    \Tile_X10Y2_S2BEGb[5] ,
    \Tile_X10Y2_S2BEGb[4] ,
    \Tile_X10Y2_S2BEGb[3] ,
    \Tile_X10Y2_S2BEGb[2] ,
    \Tile_X10Y2_S2BEGb[1] ,
    \Tile_X10Y2_S2BEGb[0] }),
    .Tile_X0Y1_S4BEG({\Tile_X10Y2_S4BEG[15] ,
    \Tile_X10Y2_S4BEG[14] ,
    \Tile_X10Y2_S4BEG[13] ,
    \Tile_X10Y2_S4BEG[12] ,
    \Tile_X10Y2_S4BEG[11] ,
    \Tile_X10Y2_S4BEG[10] ,
    \Tile_X10Y2_S4BEG[9] ,
    \Tile_X10Y2_S4BEG[8] ,
    \Tile_X10Y2_S4BEG[7] ,
    \Tile_X10Y2_S4BEG[6] ,
    \Tile_X10Y2_S4BEG[5] ,
    \Tile_X10Y2_S4BEG[4] ,
    \Tile_X10Y2_S4BEG[3] ,
    \Tile_X10Y2_S4BEG[2] ,
    \Tile_X10Y2_S4BEG[1] ,
    \Tile_X10Y2_S4BEG[0] }),
    .Tile_X0Y1_W1BEG({\Tile_X10Y2_W1BEG[3] ,
    \Tile_X10Y2_W1BEG[2] ,
    \Tile_X10Y2_W1BEG[1] ,
    \Tile_X10Y2_W1BEG[0] }),
    .Tile_X0Y1_W2BEG({\Tile_X10Y2_W2BEG[7] ,
    \Tile_X10Y2_W2BEG[6] ,
    \Tile_X10Y2_W2BEG[5] ,
    \Tile_X10Y2_W2BEG[4] ,
    \Tile_X10Y2_W2BEG[3] ,
    \Tile_X10Y2_W2BEG[2] ,
    \Tile_X10Y2_W2BEG[1] ,
    \Tile_X10Y2_W2BEG[0] }),
    .Tile_X0Y1_W2BEGb({\Tile_X10Y2_W2BEGb[7] ,
    \Tile_X10Y2_W2BEGb[6] ,
    \Tile_X10Y2_W2BEGb[5] ,
    \Tile_X10Y2_W2BEGb[4] ,
    \Tile_X10Y2_W2BEGb[3] ,
    \Tile_X10Y2_W2BEGb[2] ,
    \Tile_X10Y2_W2BEGb[1] ,
    \Tile_X10Y2_W2BEGb[0] }),
    .Tile_X0Y1_W6BEG({\Tile_X10Y2_W6BEG[11] ,
    \Tile_X10Y2_W6BEG[10] ,
    \Tile_X10Y2_W6BEG[9] ,
    \Tile_X10Y2_W6BEG[8] ,
    \Tile_X10Y2_W6BEG[7] ,
    \Tile_X10Y2_W6BEG[6] ,
    \Tile_X10Y2_W6BEG[5] ,
    \Tile_X10Y2_W6BEG[4] ,
    \Tile_X10Y2_W6BEG[3] ,
    \Tile_X10Y2_W6BEG[2] ,
    \Tile_X10Y2_W6BEG[1] ,
    \Tile_X10Y2_W6BEG[0] }),
    .Tile_X0Y1_WW4BEG({\Tile_X10Y2_WW4BEG[15] ,
    \Tile_X10Y2_WW4BEG[14] ,
    \Tile_X10Y2_WW4BEG[13] ,
    \Tile_X10Y2_WW4BEG[12] ,
    \Tile_X10Y2_WW4BEG[11] ,
    \Tile_X10Y2_WW4BEG[10] ,
    \Tile_X10Y2_WW4BEG[9] ,
    \Tile_X10Y2_WW4BEG[8] ,
    \Tile_X10Y2_WW4BEG[7] ,
    \Tile_X10Y2_WW4BEG[6] ,
    \Tile_X10Y2_WW4BEG[5] ,
    \Tile_X10Y2_WW4BEG[4] ,
    \Tile_X10Y2_WW4BEG[3] ,
    \Tile_X10Y2_WW4BEG[2] ,
    \Tile_X10Y2_WW4BEG[1] ,
    \Tile_X10Y2_WW4BEG[0] }));
 IHP_SRAM Tile_X10Y3_IHP_SRAM (.ADDR_SRAM0(Tile_X10Y4_ADDR_SRAM0),
    .ADDR_SRAM1(Tile_X10Y4_ADDR_SRAM1),
    .ADDR_SRAM2(Tile_X10Y4_ADDR_SRAM2),
    .ADDR_SRAM3(Tile_X10Y4_ADDR_SRAM3),
    .ADDR_SRAM4(Tile_X10Y4_ADDR_SRAM4),
    .ADDR_SRAM5(Tile_X10Y4_ADDR_SRAM5),
    .ADDR_SRAM6(Tile_X10Y4_ADDR_SRAM6),
    .ADDR_SRAM7(Tile_X10Y4_ADDR_SRAM7),
    .ADDR_SRAM8(Tile_X10Y4_ADDR_SRAM8),
    .ADDR_SRAM9(Tile_X10Y4_ADDR_SRAM9),
    .BM_SRAM0(Tile_X10Y4_BM_SRAM0),
    .BM_SRAM1(Tile_X10Y4_BM_SRAM1),
    .BM_SRAM10(Tile_X10Y4_BM_SRAM10),
    .BM_SRAM11(Tile_X10Y4_BM_SRAM11),
    .BM_SRAM12(Tile_X10Y4_BM_SRAM12),
    .BM_SRAM13(Tile_X10Y4_BM_SRAM13),
    .BM_SRAM14(Tile_X10Y4_BM_SRAM14),
    .BM_SRAM15(Tile_X10Y4_BM_SRAM15),
    .BM_SRAM16(Tile_X10Y4_BM_SRAM16),
    .BM_SRAM17(Tile_X10Y4_BM_SRAM17),
    .BM_SRAM18(Tile_X10Y4_BM_SRAM18),
    .BM_SRAM19(Tile_X10Y4_BM_SRAM19),
    .BM_SRAM2(Tile_X10Y4_BM_SRAM2),
    .BM_SRAM20(Tile_X10Y4_BM_SRAM20),
    .BM_SRAM21(Tile_X10Y4_BM_SRAM21),
    .BM_SRAM22(Tile_X10Y4_BM_SRAM22),
    .BM_SRAM23(Tile_X10Y4_BM_SRAM23),
    .BM_SRAM24(Tile_X10Y4_BM_SRAM24),
    .BM_SRAM25(Tile_X10Y4_BM_SRAM25),
    .BM_SRAM26(Tile_X10Y4_BM_SRAM26),
    .BM_SRAM27(Tile_X10Y4_BM_SRAM27),
    .BM_SRAM28(Tile_X10Y4_BM_SRAM28),
    .BM_SRAM29(Tile_X10Y4_BM_SRAM29),
    .BM_SRAM3(Tile_X10Y4_BM_SRAM3),
    .BM_SRAM30(Tile_X10Y4_BM_SRAM30),
    .BM_SRAM31(Tile_X10Y4_BM_SRAM31),
    .BM_SRAM4(Tile_X10Y4_BM_SRAM4),
    .BM_SRAM5(Tile_X10Y4_BM_SRAM5),
    .BM_SRAM6(Tile_X10Y4_BM_SRAM6),
    .BM_SRAM7(Tile_X10Y4_BM_SRAM7),
    .BM_SRAM8(Tile_X10Y4_BM_SRAM8),
    .BM_SRAM9(Tile_X10Y4_BM_SRAM9),
    .CLK_SRAM(Tile_X10Y4_CLK_SRAM),
    .CONFIGURED_top(Tile_X10Y4_CONFIGURED_top),
    .DIN_SRAM0(Tile_X10Y4_DIN_SRAM0),
    .DIN_SRAM1(Tile_X10Y4_DIN_SRAM1),
    .DIN_SRAM10(Tile_X10Y4_DIN_SRAM10),
    .DIN_SRAM11(Tile_X10Y4_DIN_SRAM11),
    .DIN_SRAM12(Tile_X10Y4_DIN_SRAM12),
    .DIN_SRAM13(Tile_X10Y4_DIN_SRAM13),
    .DIN_SRAM14(Tile_X10Y4_DIN_SRAM14),
    .DIN_SRAM15(Tile_X10Y4_DIN_SRAM15),
    .DIN_SRAM16(Tile_X10Y4_DIN_SRAM16),
    .DIN_SRAM17(Tile_X10Y4_DIN_SRAM17),
    .DIN_SRAM18(Tile_X10Y4_DIN_SRAM18),
    .DIN_SRAM19(Tile_X10Y4_DIN_SRAM19),
    .DIN_SRAM2(Tile_X10Y4_DIN_SRAM2),
    .DIN_SRAM20(Tile_X10Y4_DIN_SRAM20),
    .DIN_SRAM21(Tile_X10Y4_DIN_SRAM21),
    .DIN_SRAM22(Tile_X10Y4_DIN_SRAM22),
    .DIN_SRAM23(Tile_X10Y4_DIN_SRAM23),
    .DIN_SRAM24(Tile_X10Y4_DIN_SRAM24),
    .DIN_SRAM25(Tile_X10Y4_DIN_SRAM25),
    .DIN_SRAM26(Tile_X10Y4_DIN_SRAM26),
    .DIN_SRAM27(Tile_X10Y4_DIN_SRAM27),
    .DIN_SRAM28(Tile_X10Y4_DIN_SRAM28),
    .DIN_SRAM29(Tile_X10Y4_DIN_SRAM29),
    .DIN_SRAM3(Tile_X10Y4_DIN_SRAM3),
    .DIN_SRAM30(Tile_X10Y4_DIN_SRAM30),
    .DIN_SRAM31(Tile_X10Y4_DIN_SRAM31),
    .DIN_SRAM4(Tile_X10Y4_DIN_SRAM4),
    .DIN_SRAM5(Tile_X10Y4_DIN_SRAM5),
    .DIN_SRAM6(Tile_X10Y4_DIN_SRAM6),
    .DIN_SRAM7(Tile_X10Y4_DIN_SRAM7),
    .DIN_SRAM8(Tile_X10Y4_DIN_SRAM8),
    .DIN_SRAM9(Tile_X10Y4_DIN_SRAM9),
    .DOUT_SRAM0(Tile_X10Y4_DOUT_SRAM0),
    .DOUT_SRAM1(Tile_X10Y4_DOUT_SRAM1),
    .DOUT_SRAM10(Tile_X10Y4_DOUT_SRAM10),
    .DOUT_SRAM11(Tile_X10Y4_DOUT_SRAM11),
    .DOUT_SRAM12(Tile_X10Y4_DOUT_SRAM12),
    .DOUT_SRAM13(Tile_X10Y4_DOUT_SRAM13),
    .DOUT_SRAM14(Tile_X10Y4_DOUT_SRAM14),
    .DOUT_SRAM15(Tile_X10Y4_DOUT_SRAM15),
    .DOUT_SRAM16(Tile_X10Y4_DOUT_SRAM16),
    .DOUT_SRAM17(Tile_X10Y4_DOUT_SRAM17),
    .DOUT_SRAM18(Tile_X10Y4_DOUT_SRAM18),
    .DOUT_SRAM19(Tile_X10Y4_DOUT_SRAM19),
    .DOUT_SRAM2(Tile_X10Y4_DOUT_SRAM2),
    .DOUT_SRAM20(Tile_X10Y4_DOUT_SRAM20),
    .DOUT_SRAM21(Tile_X10Y4_DOUT_SRAM21),
    .DOUT_SRAM22(Tile_X10Y4_DOUT_SRAM22),
    .DOUT_SRAM23(Tile_X10Y4_DOUT_SRAM23),
    .DOUT_SRAM24(Tile_X10Y4_DOUT_SRAM24),
    .DOUT_SRAM25(Tile_X10Y4_DOUT_SRAM25),
    .DOUT_SRAM26(Tile_X10Y4_DOUT_SRAM26),
    .DOUT_SRAM27(Tile_X10Y4_DOUT_SRAM27),
    .DOUT_SRAM28(Tile_X10Y4_DOUT_SRAM28),
    .DOUT_SRAM29(Tile_X10Y4_DOUT_SRAM29),
    .DOUT_SRAM3(Tile_X10Y4_DOUT_SRAM3),
    .DOUT_SRAM30(Tile_X10Y4_DOUT_SRAM30),
    .DOUT_SRAM31(Tile_X10Y4_DOUT_SRAM31),
    .DOUT_SRAM4(Tile_X10Y4_DOUT_SRAM4),
    .DOUT_SRAM5(Tile_X10Y4_DOUT_SRAM5),
    .DOUT_SRAM6(Tile_X10Y4_DOUT_SRAM6),
    .DOUT_SRAM7(Tile_X10Y4_DOUT_SRAM7),
    .DOUT_SRAM8(Tile_X10Y4_DOUT_SRAM8),
    .DOUT_SRAM9(Tile_X10Y4_DOUT_SRAM9),
    .MEN_SRAM(Tile_X10Y4_MEN_SRAM),
    .REN_SRAM(Tile_X10Y4_REN_SRAM),
    .TIE_HIGH_SRAM(Tile_X10Y4_TIE_HIGH_SRAM),
    .TIE_LOW_SRAM(Tile_X10Y4_TIE_LOW_SRAM),
    .Tile_X0Y0_UserCLKo(Tile_X10Y3_UserCLKo),
    .Tile_X0Y1_UserCLK(Tile_X10Y5_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .WEN_SRAM(Tile_X10Y4_WEN_SRAM),
    .Tile_X0Y0_E1END({\Tile_X9Y3_E1BEG[3] ,
    \Tile_X9Y3_E1BEG[2] ,
    \Tile_X9Y3_E1BEG[1] ,
    \Tile_X9Y3_E1BEG[0] }),
    .Tile_X0Y0_E2END({\Tile_X9Y3_E2BEGb[7] ,
    \Tile_X9Y3_E2BEGb[6] ,
    \Tile_X9Y3_E2BEGb[5] ,
    \Tile_X9Y3_E2BEGb[4] ,
    \Tile_X9Y3_E2BEGb[3] ,
    \Tile_X9Y3_E2BEGb[2] ,
    \Tile_X9Y3_E2BEGb[1] ,
    \Tile_X9Y3_E2BEGb[0] }),
    .Tile_X0Y0_E2MID({\Tile_X9Y3_E2BEG[7] ,
    \Tile_X9Y3_E2BEG[6] ,
    \Tile_X9Y3_E2BEG[5] ,
    \Tile_X9Y3_E2BEG[4] ,
    \Tile_X9Y3_E2BEG[3] ,
    \Tile_X9Y3_E2BEG[2] ,
    \Tile_X9Y3_E2BEG[1] ,
    \Tile_X9Y3_E2BEG[0] }),
    .Tile_X0Y0_E6END({\Tile_X9Y3_E6BEG[11] ,
    \Tile_X9Y3_E6BEG[10] ,
    \Tile_X9Y3_E6BEG[9] ,
    \Tile_X9Y3_E6BEG[8] ,
    \Tile_X9Y3_E6BEG[7] ,
    \Tile_X9Y3_E6BEG[6] ,
    \Tile_X9Y3_E6BEG[5] ,
    \Tile_X9Y3_E6BEG[4] ,
    \Tile_X9Y3_E6BEG[3] ,
    \Tile_X9Y3_E6BEG[2] ,
    \Tile_X9Y3_E6BEG[1] ,
    \Tile_X9Y3_E6BEG[0] }),
    .Tile_X0Y0_EE4END({\Tile_X9Y3_EE4BEG[15] ,
    \Tile_X9Y3_EE4BEG[14] ,
    \Tile_X9Y3_EE4BEG[13] ,
    \Tile_X9Y3_EE4BEG[12] ,
    \Tile_X9Y3_EE4BEG[11] ,
    \Tile_X9Y3_EE4BEG[10] ,
    \Tile_X9Y3_EE4BEG[9] ,
    \Tile_X9Y3_EE4BEG[8] ,
    \Tile_X9Y3_EE4BEG[7] ,
    \Tile_X9Y3_EE4BEG[6] ,
    \Tile_X9Y3_EE4BEG[5] ,
    \Tile_X9Y3_EE4BEG[4] ,
    \Tile_X9Y3_EE4BEG[3] ,
    \Tile_X9Y3_EE4BEG[2] ,
    \Tile_X9Y3_EE4BEG[1] ,
    \Tile_X9Y3_EE4BEG[0] }),
    .Tile_X0Y0_FrameData({\Tile_X9Y3_FrameData_O[31] ,
    \Tile_X9Y3_FrameData_O[30] ,
    \Tile_X9Y3_FrameData_O[29] ,
    \Tile_X9Y3_FrameData_O[28] ,
    \Tile_X9Y3_FrameData_O[27] ,
    \Tile_X9Y3_FrameData_O[26] ,
    \Tile_X9Y3_FrameData_O[25] ,
    \Tile_X9Y3_FrameData_O[24] ,
    \Tile_X9Y3_FrameData_O[23] ,
    \Tile_X9Y3_FrameData_O[22] ,
    \Tile_X9Y3_FrameData_O[21] ,
    \Tile_X9Y3_FrameData_O[20] ,
    \Tile_X9Y3_FrameData_O[19] ,
    \Tile_X9Y3_FrameData_O[18] ,
    \Tile_X9Y3_FrameData_O[17] ,
    \Tile_X9Y3_FrameData_O[16] ,
    \Tile_X9Y3_FrameData_O[15] ,
    \Tile_X9Y3_FrameData_O[14] ,
    \Tile_X9Y3_FrameData_O[13] ,
    \Tile_X9Y3_FrameData_O[12] ,
    \Tile_X9Y3_FrameData_O[11] ,
    \Tile_X9Y3_FrameData_O[10] ,
    \Tile_X9Y3_FrameData_O[9] ,
    \Tile_X9Y3_FrameData_O[8] ,
    \Tile_X9Y3_FrameData_O[7] ,
    \Tile_X9Y3_FrameData_O[6] ,
    \Tile_X9Y3_FrameData_O[5] ,
    \Tile_X9Y3_FrameData_O[4] ,
    \Tile_X9Y3_FrameData_O[3] ,
    \Tile_X9Y3_FrameData_O[2] ,
    \Tile_X9Y3_FrameData_O[1] ,
    \Tile_X9Y3_FrameData_O[0] }),
    .Tile_X0Y0_FrameData_O({\Tile_X10Y3_FrameData_O[31] ,
    \Tile_X10Y3_FrameData_O[30] ,
    \Tile_X10Y3_FrameData_O[29] ,
    \Tile_X10Y3_FrameData_O[28] ,
    \Tile_X10Y3_FrameData_O[27] ,
    \Tile_X10Y3_FrameData_O[26] ,
    \Tile_X10Y3_FrameData_O[25] ,
    \Tile_X10Y3_FrameData_O[24] ,
    \Tile_X10Y3_FrameData_O[23] ,
    \Tile_X10Y3_FrameData_O[22] ,
    \Tile_X10Y3_FrameData_O[21] ,
    \Tile_X10Y3_FrameData_O[20] ,
    \Tile_X10Y3_FrameData_O[19] ,
    \Tile_X10Y3_FrameData_O[18] ,
    \Tile_X10Y3_FrameData_O[17] ,
    \Tile_X10Y3_FrameData_O[16] ,
    \Tile_X10Y3_FrameData_O[15] ,
    \Tile_X10Y3_FrameData_O[14] ,
    \Tile_X10Y3_FrameData_O[13] ,
    \Tile_X10Y3_FrameData_O[12] ,
    \Tile_X10Y3_FrameData_O[11] ,
    \Tile_X10Y3_FrameData_O[10] ,
    \Tile_X10Y3_FrameData_O[9] ,
    \Tile_X10Y3_FrameData_O[8] ,
    \Tile_X10Y3_FrameData_O[7] ,
    \Tile_X10Y3_FrameData_O[6] ,
    \Tile_X10Y3_FrameData_O[5] ,
    \Tile_X10Y3_FrameData_O[4] ,
    \Tile_X10Y3_FrameData_O[3] ,
    \Tile_X10Y3_FrameData_O[2] ,
    \Tile_X10Y3_FrameData_O[1] ,
    \Tile_X10Y3_FrameData_O[0] }),
    .Tile_X0Y0_FrameStrobe_O({\Tile_X10Y3_FrameStrobe_O[19] ,
    \Tile_X10Y3_FrameStrobe_O[18] ,
    \Tile_X10Y3_FrameStrobe_O[17] ,
    \Tile_X10Y3_FrameStrobe_O[16] ,
    \Tile_X10Y3_FrameStrobe_O[15] ,
    \Tile_X10Y3_FrameStrobe_O[14] ,
    \Tile_X10Y3_FrameStrobe_O[13] ,
    \Tile_X10Y3_FrameStrobe_O[12] ,
    \Tile_X10Y3_FrameStrobe_O[11] ,
    \Tile_X10Y3_FrameStrobe_O[10] ,
    \Tile_X10Y3_FrameStrobe_O[9] ,
    \Tile_X10Y3_FrameStrobe_O[8] ,
    \Tile_X10Y3_FrameStrobe_O[7] ,
    \Tile_X10Y3_FrameStrobe_O[6] ,
    \Tile_X10Y3_FrameStrobe_O[5] ,
    \Tile_X10Y3_FrameStrobe_O[4] ,
    \Tile_X10Y3_FrameStrobe_O[3] ,
    \Tile_X10Y3_FrameStrobe_O[2] ,
    \Tile_X10Y3_FrameStrobe_O[1] ,
    \Tile_X10Y3_FrameStrobe_O[0] }),
    .Tile_X0Y0_N1BEG({\Tile_X10Y3_N1BEG[3] ,
    \Tile_X10Y3_N1BEG[2] ,
    \Tile_X10Y3_N1BEG[1] ,
    \Tile_X10Y3_N1BEG[0] }),
    .Tile_X0Y0_N2BEG({\Tile_X10Y3_N2BEG[7] ,
    \Tile_X10Y3_N2BEG[6] ,
    \Tile_X10Y3_N2BEG[5] ,
    \Tile_X10Y3_N2BEG[4] ,
    \Tile_X10Y3_N2BEG[3] ,
    \Tile_X10Y3_N2BEG[2] ,
    \Tile_X10Y3_N2BEG[1] ,
    \Tile_X10Y3_N2BEG[0] }),
    .Tile_X0Y0_N2BEGb({\Tile_X10Y3_N2BEGb[7] ,
    \Tile_X10Y3_N2BEGb[6] ,
    \Tile_X10Y3_N2BEGb[5] ,
    \Tile_X10Y3_N2BEGb[4] ,
    \Tile_X10Y3_N2BEGb[3] ,
    \Tile_X10Y3_N2BEGb[2] ,
    \Tile_X10Y3_N2BEGb[1] ,
    \Tile_X10Y3_N2BEGb[0] }),
    .Tile_X0Y0_N4BEG({\Tile_X10Y3_N4BEG[15] ,
    \Tile_X10Y3_N4BEG[14] ,
    \Tile_X10Y3_N4BEG[13] ,
    \Tile_X10Y3_N4BEG[12] ,
    \Tile_X10Y3_N4BEG[11] ,
    \Tile_X10Y3_N4BEG[10] ,
    \Tile_X10Y3_N4BEG[9] ,
    \Tile_X10Y3_N4BEG[8] ,
    \Tile_X10Y3_N4BEG[7] ,
    \Tile_X10Y3_N4BEG[6] ,
    \Tile_X10Y3_N4BEG[5] ,
    \Tile_X10Y3_N4BEG[4] ,
    \Tile_X10Y3_N4BEG[3] ,
    \Tile_X10Y3_N4BEG[2] ,
    \Tile_X10Y3_N4BEG[1] ,
    \Tile_X10Y3_N4BEG[0] }),
    .Tile_X0Y0_S1END({\Tile_X10Y2_S1BEG[3] ,
    \Tile_X10Y2_S1BEG[2] ,
    \Tile_X10Y2_S1BEG[1] ,
    \Tile_X10Y2_S1BEG[0] }),
    .Tile_X0Y0_S2END({\Tile_X10Y2_S2BEGb[7] ,
    \Tile_X10Y2_S2BEGb[6] ,
    \Tile_X10Y2_S2BEGb[5] ,
    \Tile_X10Y2_S2BEGb[4] ,
    \Tile_X10Y2_S2BEGb[3] ,
    \Tile_X10Y2_S2BEGb[2] ,
    \Tile_X10Y2_S2BEGb[1] ,
    \Tile_X10Y2_S2BEGb[0] }),
    .Tile_X0Y0_S2MID({\Tile_X10Y2_S2BEG[7] ,
    \Tile_X10Y2_S2BEG[6] ,
    \Tile_X10Y2_S2BEG[5] ,
    \Tile_X10Y2_S2BEG[4] ,
    \Tile_X10Y2_S2BEG[3] ,
    \Tile_X10Y2_S2BEG[2] ,
    \Tile_X10Y2_S2BEG[1] ,
    \Tile_X10Y2_S2BEG[0] }),
    .Tile_X0Y0_S4END({\Tile_X10Y2_S4BEG[15] ,
    \Tile_X10Y2_S4BEG[14] ,
    \Tile_X10Y2_S4BEG[13] ,
    \Tile_X10Y2_S4BEG[12] ,
    \Tile_X10Y2_S4BEG[11] ,
    \Tile_X10Y2_S4BEG[10] ,
    \Tile_X10Y2_S4BEG[9] ,
    \Tile_X10Y2_S4BEG[8] ,
    \Tile_X10Y2_S4BEG[7] ,
    \Tile_X10Y2_S4BEG[6] ,
    \Tile_X10Y2_S4BEG[5] ,
    \Tile_X10Y2_S4BEG[4] ,
    \Tile_X10Y2_S4BEG[3] ,
    \Tile_X10Y2_S4BEG[2] ,
    \Tile_X10Y2_S4BEG[1] ,
    \Tile_X10Y2_S4BEG[0] }),
    .Tile_X0Y0_W1BEG({\Tile_X10Y3_W1BEG[3] ,
    \Tile_X10Y3_W1BEG[2] ,
    \Tile_X10Y3_W1BEG[1] ,
    \Tile_X10Y3_W1BEG[0] }),
    .Tile_X0Y0_W2BEG({\Tile_X10Y3_W2BEG[7] ,
    \Tile_X10Y3_W2BEG[6] ,
    \Tile_X10Y3_W2BEG[5] ,
    \Tile_X10Y3_W2BEG[4] ,
    \Tile_X10Y3_W2BEG[3] ,
    \Tile_X10Y3_W2BEG[2] ,
    \Tile_X10Y3_W2BEG[1] ,
    \Tile_X10Y3_W2BEG[0] }),
    .Tile_X0Y0_W2BEGb({\Tile_X10Y3_W2BEGb[7] ,
    \Tile_X10Y3_W2BEGb[6] ,
    \Tile_X10Y3_W2BEGb[5] ,
    \Tile_X10Y3_W2BEGb[4] ,
    \Tile_X10Y3_W2BEGb[3] ,
    \Tile_X10Y3_W2BEGb[2] ,
    \Tile_X10Y3_W2BEGb[1] ,
    \Tile_X10Y3_W2BEGb[0] }),
    .Tile_X0Y0_W6BEG({\Tile_X10Y3_W6BEG[11] ,
    \Tile_X10Y3_W6BEG[10] ,
    \Tile_X10Y3_W6BEG[9] ,
    \Tile_X10Y3_W6BEG[8] ,
    \Tile_X10Y3_W6BEG[7] ,
    \Tile_X10Y3_W6BEG[6] ,
    \Tile_X10Y3_W6BEG[5] ,
    \Tile_X10Y3_W6BEG[4] ,
    \Tile_X10Y3_W6BEG[3] ,
    \Tile_X10Y3_W6BEG[2] ,
    \Tile_X10Y3_W6BEG[1] ,
    \Tile_X10Y3_W6BEG[0] }),
    .Tile_X0Y0_WW4BEG({\Tile_X10Y3_WW4BEG[15] ,
    \Tile_X10Y3_WW4BEG[14] ,
    \Tile_X10Y3_WW4BEG[13] ,
    \Tile_X10Y3_WW4BEG[12] ,
    \Tile_X10Y3_WW4BEG[11] ,
    \Tile_X10Y3_WW4BEG[10] ,
    \Tile_X10Y3_WW4BEG[9] ,
    \Tile_X10Y3_WW4BEG[8] ,
    \Tile_X10Y3_WW4BEG[7] ,
    \Tile_X10Y3_WW4BEG[6] ,
    \Tile_X10Y3_WW4BEG[5] ,
    \Tile_X10Y3_WW4BEG[4] ,
    \Tile_X10Y3_WW4BEG[3] ,
    \Tile_X10Y3_WW4BEG[2] ,
    \Tile_X10Y3_WW4BEG[1] ,
    \Tile_X10Y3_WW4BEG[0] }),
    .Tile_X0Y1_E1END({\Tile_X9Y4_E1BEG[3] ,
    \Tile_X9Y4_E1BEG[2] ,
    \Tile_X9Y4_E1BEG[1] ,
    \Tile_X9Y4_E1BEG[0] }),
    .Tile_X0Y1_E2END({\Tile_X9Y4_E2BEGb[7] ,
    \Tile_X9Y4_E2BEGb[6] ,
    \Tile_X9Y4_E2BEGb[5] ,
    \Tile_X9Y4_E2BEGb[4] ,
    \Tile_X9Y4_E2BEGb[3] ,
    \Tile_X9Y4_E2BEGb[2] ,
    \Tile_X9Y4_E2BEGb[1] ,
    \Tile_X9Y4_E2BEGb[0] }),
    .Tile_X0Y1_E2MID({\Tile_X9Y4_E2BEG[7] ,
    \Tile_X9Y4_E2BEG[6] ,
    \Tile_X9Y4_E2BEG[5] ,
    \Tile_X9Y4_E2BEG[4] ,
    \Tile_X9Y4_E2BEG[3] ,
    \Tile_X9Y4_E2BEG[2] ,
    \Tile_X9Y4_E2BEG[1] ,
    \Tile_X9Y4_E2BEG[0] }),
    .Tile_X0Y1_E6END({\Tile_X9Y4_E6BEG[11] ,
    \Tile_X9Y4_E6BEG[10] ,
    \Tile_X9Y4_E6BEG[9] ,
    \Tile_X9Y4_E6BEG[8] ,
    \Tile_X9Y4_E6BEG[7] ,
    \Tile_X9Y4_E6BEG[6] ,
    \Tile_X9Y4_E6BEG[5] ,
    \Tile_X9Y4_E6BEG[4] ,
    \Tile_X9Y4_E6BEG[3] ,
    \Tile_X9Y4_E6BEG[2] ,
    \Tile_X9Y4_E6BEG[1] ,
    \Tile_X9Y4_E6BEG[0] }),
    .Tile_X0Y1_EE4END({\Tile_X9Y4_EE4BEG[15] ,
    \Tile_X9Y4_EE4BEG[14] ,
    \Tile_X9Y4_EE4BEG[13] ,
    \Tile_X9Y4_EE4BEG[12] ,
    \Tile_X9Y4_EE4BEG[11] ,
    \Tile_X9Y4_EE4BEG[10] ,
    \Tile_X9Y4_EE4BEG[9] ,
    \Tile_X9Y4_EE4BEG[8] ,
    \Tile_X9Y4_EE4BEG[7] ,
    \Tile_X9Y4_EE4BEG[6] ,
    \Tile_X9Y4_EE4BEG[5] ,
    \Tile_X9Y4_EE4BEG[4] ,
    \Tile_X9Y4_EE4BEG[3] ,
    \Tile_X9Y4_EE4BEG[2] ,
    \Tile_X9Y4_EE4BEG[1] ,
    \Tile_X9Y4_EE4BEG[0] }),
    .Tile_X0Y1_FrameData({\Tile_X9Y4_FrameData_O[31] ,
    \Tile_X9Y4_FrameData_O[30] ,
    \Tile_X9Y4_FrameData_O[29] ,
    \Tile_X9Y4_FrameData_O[28] ,
    \Tile_X9Y4_FrameData_O[27] ,
    \Tile_X9Y4_FrameData_O[26] ,
    \Tile_X9Y4_FrameData_O[25] ,
    \Tile_X9Y4_FrameData_O[24] ,
    \Tile_X9Y4_FrameData_O[23] ,
    \Tile_X9Y4_FrameData_O[22] ,
    \Tile_X9Y4_FrameData_O[21] ,
    \Tile_X9Y4_FrameData_O[20] ,
    \Tile_X9Y4_FrameData_O[19] ,
    \Tile_X9Y4_FrameData_O[18] ,
    \Tile_X9Y4_FrameData_O[17] ,
    \Tile_X9Y4_FrameData_O[16] ,
    \Tile_X9Y4_FrameData_O[15] ,
    \Tile_X9Y4_FrameData_O[14] ,
    \Tile_X9Y4_FrameData_O[13] ,
    \Tile_X9Y4_FrameData_O[12] ,
    \Tile_X9Y4_FrameData_O[11] ,
    \Tile_X9Y4_FrameData_O[10] ,
    \Tile_X9Y4_FrameData_O[9] ,
    \Tile_X9Y4_FrameData_O[8] ,
    \Tile_X9Y4_FrameData_O[7] ,
    \Tile_X9Y4_FrameData_O[6] ,
    \Tile_X9Y4_FrameData_O[5] ,
    \Tile_X9Y4_FrameData_O[4] ,
    \Tile_X9Y4_FrameData_O[3] ,
    \Tile_X9Y4_FrameData_O[2] ,
    \Tile_X9Y4_FrameData_O[1] ,
    \Tile_X9Y4_FrameData_O[0] }),
    .Tile_X0Y1_FrameData_O({\Tile_X10Y4_FrameData_O[31] ,
    \Tile_X10Y4_FrameData_O[30] ,
    \Tile_X10Y4_FrameData_O[29] ,
    \Tile_X10Y4_FrameData_O[28] ,
    \Tile_X10Y4_FrameData_O[27] ,
    \Tile_X10Y4_FrameData_O[26] ,
    \Tile_X10Y4_FrameData_O[25] ,
    \Tile_X10Y4_FrameData_O[24] ,
    \Tile_X10Y4_FrameData_O[23] ,
    \Tile_X10Y4_FrameData_O[22] ,
    \Tile_X10Y4_FrameData_O[21] ,
    \Tile_X10Y4_FrameData_O[20] ,
    \Tile_X10Y4_FrameData_O[19] ,
    \Tile_X10Y4_FrameData_O[18] ,
    \Tile_X10Y4_FrameData_O[17] ,
    \Tile_X10Y4_FrameData_O[16] ,
    \Tile_X10Y4_FrameData_O[15] ,
    \Tile_X10Y4_FrameData_O[14] ,
    \Tile_X10Y4_FrameData_O[13] ,
    \Tile_X10Y4_FrameData_O[12] ,
    \Tile_X10Y4_FrameData_O[11] ,
    \Tile_X10Y4_FrameData_O[10] ,
    \Tile_X10Y4_FrameData_O[9] ,
    \Tile_X10Y4_FrameData_O[8] ,
    \Tile_X10Y4_FrameData_O[7] ,
    \Tile_X10Y4_FrameData_O[6] ,
    \Tile_X10Y4_FrameData_O[5] ,
    \Tile_X10Y4_FrameData_O[4] ,
    \Tile_X10Y4_FrameData_O[3] ,
    \Tile_X10Y4_FrameData_O[2] ,
    \Tile_X10Y4_FrameData_O[1] ,
    \Tile_X10Y4_FrameData_O[0] }),
    .Tile_X0Y1_FrameStrobe({\Tile_X10Y5_FrameStrobe_O[19] ,
    \Tile_X10Y5_FrameStrobe_O[18] ,
    \Tile_X10Y5_FrameStrobe_O[17] ,
    \Tile_X10Y5_FrameStrobe_O[16] ,
    \Tile_X10Y5_FrameStrobe_O[15] ,
    \Tile_X10Y5_FrameStrobe_O[14] ,
    \Tile_X10Y5_FrameStrobe_O[13] ,
    \Tile_X10Y5_FrameStrobe_O[12] ,
    \Tile_X10Y5_FrameStrobe_O[11] ,
    \Tile_X10Y5_FrameStrobe_O[10] ,
    \Tile_X10Y5_FrameStrobe_O[9] ,
    \Tile_X10Y5_FrameStrobe_O[8] ,
    \Tile_X10Y5_FrameStrobe_O[7] ,
    \Tile_X10Y5_FrameStrobe_O[6] ,
    \Tile_X10Y5_FrameStrobe_O[5] ,
    \Tile_X10Y5_FrameStrobe_O[4] ,
    \Tile_X10Y5_FrameStrobe_O[3] ,
    \Tile_X10Y5_FrameStrobe_O[2] ,
    \Tile_X10Y5_FrameStrobe_O[1] ,
    \Tile_X10Y5_FrameStrobe_O[0] }),
    .Tile_X0Y1_N1END({\Tile_X10Y5_N1BEG[3] ,
    \Tile_X10Y5_N1BEG[2] ,
    \Tile_X10Y5_N1BEG[1] ,
    \Tile_X10Y5_N1BEG[0] }),
    .Tile_X0Y1_N2END({\Tile_X10Y5_N2BEGb[7] ,
    \Tile_X10Y5_N2BEGb[6] ,
    \Tile_X10Y5_N2BEGb[5] ,
    \Tile_X10Y5_N2BEGb[4] ,
    \Tile_X10Y5_N2BEGb[3] ,
    \Tile_X10Y5_N2BEGb[2] ,
    \Tile_X10Y5_N2BEGb[1] ,
    \Tile_X10Y5_N2BEGb[0] }),
    .Tile_X0Y1_N2MID({\Tile_X10Y5_N2BEG[7] ,
    \Tile_X10Y5_N2BEG[6] ,
    \Tile_X10Y5_N2BEG[5] ,
    \Tile_X10Y5_N2BEG[4] ,
    \Tile_X10Y5_N2BEG[3] ,
    \Tile_X10Y5_N2BEG[2] ,
    \Tile_X10Y5_N2BEG[1] ,
    \Tile_X10Y5_N2BEG[0] }),
    .Tile_X0Y1_N4END({\Tile_X10Y5_N4BEG[15] ,
    \Tile_X10Y5_N4BEG[14] ,
    \Tile_X10Y5_N4BEG[13] ,
    \Tile_X10Y5_N4BEG[12] ,
    \Tile_X10Y5_N4BEG[11] ,
    \Tile_X10Y5_N4BEG[10] ,
    \Tile_X10Y5_N4BEG[9] ,
    \Tile_X10Y5_N4BEG[8] ,
    \Tile_X10Y5_N4BEG[7] ,
    \Tile_X10Y5_N4BEG[6] ,
    \Tile_X10Y5_N4BEG[5] ,
    \Tile_X10Y5_N4BEG[4] ,
    \Tile_X10Y5_N4BEG[3] ,
    \Tile_X10Y5_N4BEG[2] ,
    \Tile_X10Y5_N4BEG[1] ,
    \Tile_X10Y5_N4BEG[0] }),
    .Tile_X0Y1_S1BEG({\Tile_X10Y4_S1BEG[3] ,
    \Tile_X10Y4_S1BEG[2] ,
    \Tile_X10Y4_S1BEG[1] ,
    \Tile_X10Y4_S1BEG[0] }),
    .Tile_X0Y1_S2BEG({\Tile_X10Y4_S2BEG[7] ,
    \Tile_X10Y4_S2BEG[6] ,
    \Tile_X10Y4_S2BEG[5] ,
    \Tile_X10Y4_S2BEG[4] ,
    \Tile_X10Y4_S2BEG[3] ,
    \Tile_X10Y4_S2BEG[2] ,
    \Tile_X10Y4_S2BEG[1] ,
    \Tile_X10Y4_S2BEG[0] }),
    .Tile_X0Y1_S2BEGb({\Tile_X10Y4_S2BEGb[7] ,
    \Tile_X10Y4_S2BEGb[6] ,
    \Tile_X10Y4_S2BEGb[5] ,
    \Tile_X10Y4_S2BEGb[4] ,
    \Tile_X10Y4_S2BEGb[3] ,
    \Tile_X10Y4_S2BEGb[2] ,
    \Tile_X10Y4_S2BEGb[1] ,
    \Tile_X10Y4_S2BEGb[0] }),
    .Tile_X0Y1_S4BEG({\Tile_X10Y4_S4BEG[15] ,
    \Tile_X10Y4_S4BEG[14] ,
    \Tile_X10Y4_S4BEG[13] ,
    \Tile_X10Y4_S4BEG[12] ,
    \Tile_X10Y4_S4BEG[11] ,
    \Tile_X10Y4_S4BEG[10] ,
    \Tile_X10Y4_S4BEG[9] ,
    \Tile_X10Y4_S4BEG[8] ,
    \Tile_X10Y4_S4BEG[7] ,
    \Tile_X10Y4_S4BEG[6] ,
    \Tile_X10Y4_S4BEG[5] ,
    \Tile_X10Y4_S4BEG[4] ,
    \Tile_X10Y4_S4BEG[3] ,
    \Tile_X10Y4_S4BEG[2] ,
    \Tile_X10Y4_S4BEG[1] ,
    \Tile_X10Y4_S4BEG[0] }),
    .Tile_X0Y1_W1BEG({\Tile_X10Y4_W1BEG[3] ,
    \Tile_X10Y4_W1BEG[2] ,
    \Tile_X10Y4_W1BEG[1] ,
    \Tile_X10Y4_W1BEG[0] }),
    .Tile_X0Y1_W2BEG({\Tile_X10Y4_W2BEG[7] ,
    \Tile_X10Y4_W2BEG[6] ,
    \Tile_X10Y4_W2BEG[5] ,
    \Tile_X10Y4_W2BEG[4] ,
    \Tile_X10Y4_W2BEG[3] ,
    \Tile_X10Y4_W2BEG[2] ,
    \Tile_X10Y4_W2BEG[1] ,
    \Tile_X10Y4_W2BEG[0] }),
    .Tile_X0Y1_W2BEGb({\Tile_X10Y4_W2BEGb[7] ,
    \Tile_X10Y4_W2BEGb[6] ,
    \Tile_X10Y4_W2BEGb[5] ,
    \Tile_X10Y4_W2BEGb[4] ,
    \Tile_X10Y4_W2BEGb[3] ,
    \Tile_X10Y4_W2BEGb[2] ,
    \Tile_X10Y4_W2BEGb[1] ,
    \Tile_X10Y4_W2BEGb[0] }),
    .Tile_X0Y1_W6BEG({\Tile_X10Y4_W6BEG[11] ,
    \Tile_X10Y4_W6BEG[10] ,
    \Tile_X10Y4_W6BEG[9] ,
    \Tile_X10Y4_W6BEG[8] ,
    \Tile_X10Y4_W6BEG[7] ,
    \Tile_X10Y4_W6BEG[6] ,
    \Tile_X10Y4_W6BEG[5] ,
    \Tile_X10Y4_W6BEG[4] ,
    \Tile_X10Y4_W6BEG[3] ,
    \Tile_X10Y4_W6BEG[2] ,
    \Tile_X10Y4_W6BEG[1] ,
    \Tile_X10Y4_W6BEG[0] }),
    .Tile_X0Y1_WW4BEG({\Tile_X10Y4_WW4BEG[15] ,
    \Tile_X10Y4_WW4BEG[14] ,
    \Tile_X10Y4_WW4BEG[13] ,
    \Tile_X10Y4_WW4BEG[12] ,
    \Tile_X10Y4_WW4BEG[11] ,
    \Tile_X10Y4_WW4BEG[10] ,
    \Tile_X10Y4_WW4BEG[9] ,
    \Tile_X10Y4_WW4BEG[8] ,
    \Tile_X10Y4_WW4BEG[7] ,
    \Tile_X10Y4_WW4BEG[6] ,
    \Tile_X10Y4_WW4BEG[5] ,
    \Tile_X10Y4_WW4BEG[4] ,
    \Tile_X10Y4_WW4BEG[3] ,
    \Tile_X10Y4_WW4BEG[2] ,
    \Tile_X10Y4_WW4BEG[1] ,
    \Tile_X10Y4_WW4BEG[0] }));
 IHP_SRAM Tile_X10Y5_IHP_SRAM (.ADDR_SRAM0(Tile_X10Y6_ADDR_SRAM0),
    .ADDR_SRAM1(Tile_X10Y6_ADDR_SRAM1),
    .ADDR_SRAM2(Tile_X10Y6_ADDR_SRAM2),
    .ADDR_SRAM3(Tile_X10Y6_ADDR_SRAM3),
    .ADDR_SRAM4(Tile_X10Y6_ADDR_SRAM4),
    .ADDR_SRAM5(Tile_X10Y6_ADDR_SRAM5),
    .ADDR_SRAM6(Tile_X10Y6_ADDR_SRAM6),
    .ADDR_SRAM7(Tile_X10Y6_ADDR_SRAM7),
    .ADDR_SRAM8(Tile_X10Y6_ADDR_SRAM8),
    .ADDR_SRAM9(Tile_X10Y6_ADDR_SRAM9),
    .BM_SRAM0(Tile_X10Y6_BM_SRAM0),
    .BM_SRAM1(Tile_X10Y6_BM_SRAM1),
    .BM_SRAM10(Tile_X10Y6_BM_SRAM10),
    .BM_SRAM11(Tile_X10Y6_BM_SRAM11),
    .BM_SRAM12(Tile_X10Y6_BM_SRAM12),
    .BM_SRAM13(Tile_X10Y6_BM_SRAM13),
    .BM_SRAM14(Tile_X10Y6_BM_SRAM14),
    .BM_SRAM15(Tile_X10Y6_BM_SRAM15),
    .BM_SRAM16(Tile_X10Y6_BM_SRAM16),
    .BM_SRAM17(Tile_X10Y6_BM_SRAM17),
    .BM_SRAM18(Tile_X10Y6_BM_SRAM18),
    .BM_SRAM19(Tile_X10Y6_BM_SRAM19),
    .BM_SRAM2(Tile_X10Y6_BM_SRAM2),
    .BM_SRAM20(Tile_X10Y6_BM_SRAM20),
    .BM_SRAM21(Tile_X10Y6_BM_SRAM21),
    .BM_SRAM22(Tile_X10Y6_BM_SRAM22),
    .BM_SRAM23(Tile_X10Y6_BM_SRAM23),
    .BM_SRAM24(Tile_X10Y6_BM_SRAM24),
    .BM_SRAM25(Tile_X10Y6_BM_SRAM25),
    .BM_SRAM26(Tile_X10Y6_BM_SRAM26),
    .BM_SRAM27(Tile_X10Y6_BM_SRAM27),
    .BM_SRAM28(Tile_X10Y6_BM_SRAM28),
    .BM_SRAM29(Tile_X10Y6_BM_SRAM29),
    .BM_SRAM3(Tile_X10Y6_BM_SRAM3),
    .BM_SRAM30(Tile_X10Y6_BM_SRAM30),
    .BM_SRAM31(Tile_X10Y6_BM_SRAM31),
    .BM_SRAM4(Tile_X10Y6_BM_SRAM4),
    .BM_SRAM5(Tile_X10Y6_BM_SRAM5),
    .BM_SRAM6(Tile_X10Y6_BM_SRAM6),
    .BM_SRAM7(Tile_X10Y6_BM_SRAM7),
    .BM_SRAM8(Tile_X10Y6_BM_SRAM8),
    .BM_SRAM9(Tile_X10Y6_BM_SRAM9),
    .CLK_SRAM(Tile_X10Y6_CLK_SRAM),
    .CONFIGURED_top(Tile_X10Y6_CONFIGURED_top),
    .DIN_SRAM0(Tile_X10Y6_DIN_SRAM0),
    .DIN_SRAM1(Tile_X10Y6_DIN_SRAM1),
    .DIN_SRAM10(Tile_X10Y6_DIN_SRAM10),
    .DIN_SRAM11(Tile_X10Y6_DIN_SRAM11),
    .DIN_SRAM12(Tile_X10Y6_DIN_SRAM12),
    .DIN_SRAM13(Tile_X10Y6_DIN_SRAM13),
    .DIN_SRAM14(Tile_X10Y6_DIN_SRAM14),
    .DIN_SRAM15(Tile_X10Y6_DIN_SRAM15),
    .DIN_SRAM16(Tile_X10Y6_DIN_SRAM16),
    .DIN_SRAM17(Tile_X10Y6_DIN_SRAM17),
    .DIN_SRAM18(Tile_X10Y6_DIN_SRAM18),
    .DIN_SRAM19(Tile_X10Y6_DIN_SRAM19),
    .DIN_SRAM2(Tile_X10Y6_DIN_SRAM2),
    .DIN_SRAM20(Tile_X10Y6_DIN_SRAM20),
    .DIN_SRAM21(Tile_X10Y6_DIN_SRAM21),
    .DIN_SRAM22(Tile_X10Y6_DIN_SRAM22),
    .DIN_SRAM23(Tile_X10Y6_DIN_SRAM23),
    .DIN_SRAM24(Tile_X10Y6_DIN_SRAM24),
    .DIN_SRAM25(Tile_X10Y6_DIN_SRAM25),
    .DIN_SRAM26(Tile_X10Y6_DIN_SRAM26),
    .DIN_SRAM27(Tile_X10Y6_DIN_SRAM27),
    .DIN_SRAM28(Tile_X10Y6_DIN_SRAM28),
    .DIN_SRAM29(Tile_X10Y6_DIN_SRAM29),
    .DIN_SRAM3(Tile_X10Y6_DIN_SRAM3),
    .DIN_SRAM30(Tile_X10Y6_DIN_SRAM30),
    .DIN_SRAM31(Tile_X10Y6_DIN_SRAM31),
    .DIN_SRAM4(Tile_X10Y6_DIN_SRAM4),
    .DIN_SRAM5(Tile_X10Y6_DIN_SRAM5),
    .DIN_SRAM6(Tile_X10Y6_DIN_SRAM6),
    .DIN_SRAM7(Tile_X10Y6_DIN_SRAM7),
    .DIN_SRAM8(Tile_X10Y6_DIN_SRAM8),
    .DIN_SRAM9(Tile_X10Y6_DIN_SRAM9),
    .DOUT_SRAM0(Tile_X10Y6_DOUT_SRAM0),
    .DOUT_SRAM1(Tile_X10Y6_DOUT_SRAM1),
    .DOUT_SRAM10(Tile_X10Y6_DOUT_SRAM10),
    .DOUT_SRAM11(Tile_X10Y6_DOUT_SRAM11),
    .DOUT_SRAM12(Tile_X10Y6_DOUT_SRAM12),
    .DOUT_SRAM13(Tile_X10Y6_DOUT_SRAM13),
    .DOUT_SRAM14(Tile_X10Y6_DOUT_SRAM14),
    .DOUT_SRAM15(Tile_X10Y6_DOUT_SRAM15),
    .DOUT_SRAM16(Tile_X10Y6_DOUT_SRAM16),
    .DOUT_SRAM17(Tile_X10Y6_DOUT_SRAM17),
    .DOUT_SRAM18(Tile_X10Y6_DOUT_SRAM18),
    .DOUT_SRAM19(Tile_X10Y6_DOUT_SRAM19),
    .DOUT_SRAM2(Tile_X10Y6_DOUT_SRAM2),
    .DOUT_SRAM20(Tile_X10Y6_DOUT_SRAM20),
    .DOUT_SRAM21(Tile_X10Y6_DOUT_SRAM21),
    .DOUT_SRAM22(Tile_X10Y6_DOUT_SRAM22),
    .DOUT_SRAM23(Tile_X10Y6_DOUT_SRAM23),
    .DOUT_SRAM24(Tile_X10Y6_DOUT_SRAM24),
    .DOUT_SRAM25(Tile_X10Y6_DOUT_SRAM25),
    .DOUT_SRAM26(Tile_X10Y6_DOUT_SRAM26),
    .DOUT_SRAM27(Tile_X10Y6_DOUT_SRAM27),
    .DOUT_SRAM28(Tile_X10Y6_DOUT_SRAM28),
    .DOUT_SRAM29(Tile_X10Y6_DOUT_SRAM29),
    .DOUT_SRAM3(Tile_X10Y6_DOUT_SRAM3),
    .DOUT_SRAM30(Tile_X10Y6_DOUT_SRAM30),
    .DOUT_SRAM31(Tile_X10Y6_DOUT_SRAM31),
    .DOUT_SRAM4(Tile_X10Y6_DOUT_SRAM4),
    .DOUT_SRAM5(Tile_X10Y6_DOUT_SRAM5),
    .DOUT_SRAM6(Tile_X10Y6_DOUT_SRAM6),
    .DOUT_SRAM7(Tile_X10Y6_DOUT_SRAM7),
    .DOUT_SRAM8(Tile_X10Y6_DOUT_SRAM8),
    .DOUT_SRAM9(Tile_X10Y6_DOUT_SRAM9),
    .MEN_SRAM(Tile_X10Y6_MEN_SRAM),
    .REN_SRAM(Tile_X10Y6_REN_SRAM),
    .TIE_HIGH_SRAM(Tile_X10Y6_TIE_HIGH_SRAM),
    .TIE_LOW_SRAM(Tile_X10Y6_TIE_LOW_SRAM),
    .Tile_X0Y0_UserCLKo(Tile_X10Y5_UserCLKo),
    .Tile_X0Y1_UserCLK(Tile_X10Y7_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .WEN_SRAM(Tile_X10Y6_WEN_SRAM),
    .Tile_X0Y0_E1END({\Tile_X9Y5_E1BEG[3] ,
    \Tile_X9Y5_E1BEG[2] ,
    \Tile_X9Y5_E1BEG[1] ,
    \Tile_X9Y5_E1BEG[0] }),
    .Tile_X0Y0_E2END({\Tile_X9Y5_E2BEGb[7] ,
    \Tile_X9Y5_E2BEGb[6] ,
    \Tile_X9Y5_E2BEGb[5] ,
    \Tile_X9Y5_E2BEGb[4] ,
    \Tile_X9Y5_E2BEGb[3] ,
    \Tile_X9Y5_E2BEGb[2] ,
    \Tile_X9Y5_E2BEGb[1] ,
    \Tile_X9Y5_E2BEGb[0] }),
    .Tile_X0Y0_E2MID({\Tile_X9Y5_E2BEG[7] ,
    \Tile_X9Y5_E2BEG[6] ,
    \Tile_X9Y5_E2BEG[5] ,
    \Tile_X9Y5_E2BEG[4] ,
    \Tile_X9Y5_E2BEG[3] ,
    \Tile_X9Y5_E2BEG[2] ,
    \Tile_X9Y5_E2BEG[1] ,
    \Tile_X9Y5_E2BEG[0] }),
    .Tile_X0Y0_E6END({\Tile_X9Y5_E6BEG[11] ,
    \Tile_X9Y5_E6BEG[10] ,
    \Tile_X9Y5_E6BEG[9] ,
    \Tile_X9Y5_E6BEG[8] ,
    \Tile_X9Y5_E6BEG[7] ,
    \Tile_X9Y5_E6BEG[6] ,
    \Tile_X9Y5_E6BEG[5] ,
    \Tile_X9Y5_E6BEG[4] ,
    \Tile_X9Y5_E6BEG[3] ,
    \Tile_X9Y5_E6BEG[2] ,
    \Tile_X9Y5_E6BEG[1] ,
    \Tile_X9Y5_E6BEG[0] }),
    .Tile_X0Y0_EE4END({\Tile_X9Y5_EE4BEG[15] ,
    \Tile_X9Y5_EE4BEG[14] ,
    \Tile_X9Y5_EE4BEG[13] ,
    \Tile_X9Y5_EE4BEG[12] ,
    \Tile_X9Y5_EE4BEG[11] ,
    \Tile_X9Y5_EE4BEG[10] ,
    \Tile_X9Y5_EE4BEG[9] ,
    \Tile_X9Y5_EE4BEG[8] ,
    \Tile_X9Y5_EE4BEG[7] ,
    \Tile_X9Y5_EE4BEG[6] ,
    \Tile_X9Y5_EE4BEG[5] ,
    \Tile_X9Y5_EE4BEG[4] ,
    \Tile_X9Y5_EE4BEG[3] ,
    \Tile_X9Y5_EE4BEG[2] ,
    \Tile_X9Y5_EE4BEG[1] ,
    \Tile_X9Y5_EE4BEG[0] }),
    .Tile_X0Y0_FrameData({\Tile_X9Y5_FrameData_O[31] ,
    \Tile_X9Y5_FrameData_O[30] ,
    \Tile_X9Y5_FrameData_O[29] ,
    \Tile_X9Y5_FrameData_O[28] ,
    \Tile_X9Y5_FrameData_O[27] ,
    \Tile_X9Y5_FrameData_O[26] ,
    \Tile_X9Y5_FrameData_O[25] ,
    \Tile_X9Y5_FrameData_O[24] ,
    \Tile_X9Y5_FrameData_O[23] ,
    \Tile_X9Y5_FrameData_O[22] ,
    \Tile_X9Y5_FrameData_O[21] ,
    \Tile_X9Y5_FrameData_O[20] ,
    \Tile_X9Y5_FrameData_O[19] ,
    \Tile_X9Y5_FrameData_O[18] ,
    \Tile_X9Y5_FrameData_O[17] ,
    \Tile_X9Y5_FrameData_O[16] ,
    \Tile_X9Y5_FrameData_O[15] ,
    \Tile_X9Y5_FrameData_O[14] ,
    \Tile_X9Y5_FrameData_O[13] ,
    \Tile_X9Y5_FrameData_O[12] ,
    \Tile_X9Y5_FrameData_O[11] ,
    \Tile_X9Y5_FrameData_O[10] ,
    \Tile_X9Y5_FrameData_O[9] ,
    \Tile_X9Y5_FrameData_O[8] ,
    \Tile_X9Y5_FrameData_O[7] ,
    \Tile_X9Y5_FrameData_O[6] ,
    \Tile_X9Y5_FrameData_O[5] ,
    \Tile_X9Y5_FrameData_O[4] ,
    \Tile_X9Y5_FrameData_O[3] ,
    \Tile_X9Y5_FrameData_O[2] ,
    \Tile_X9Y5_FrameData_O[1] ,
    \Tile_X9Y5_FrameData_O[0] }),
    .Tile_X0Y0_FrameData_O({\Tile_X10Y5_FrameData_O[31] ,
    \Tile_X10Y5_FrameData_O[30] ,
    \Tile_X10Y5_FrameData_O[29] ,
    \Tile_X10Y5_FrameData_O[28] ,
    \Tile_X10Y5_FrameData_O[27] ,
    \Tile_X10Y5_FrameData_O[26] ,
    \Tile_X10Y5_FrameData_O[25] ,
    \Tile_X10Y5_FrameData_O[24] ,
    \Tile_X10Y5_FrameData_O[23] ,
    \Tile_X10Y5_FrameData_O[22] ,
    \Tile_X10Y5_FrameData_O[21] ,
    \Tile_X10Y5_FrameData_O[20] ,
    \Tile_X10Y5_FrameData_O[19] ,
    \Tile_X10Y5_FrameData_O[18] ,
    \Tile_X10Y5_FrameData_O[17] ,
    \Tile_X10Y5_FrameData_O[16] ,
    \Tile_X10Y5_FrameData_O[15] ,
    \Tile_X10Y5_FrameData_O[14] ,
    \Tile_X10Y5_FrameData_O[13] ,
    \Tile_X10Y5_FrameData_O[12] ,
    \Tile_X10Y5_FrameData_O[11] ,
    \Tile_X10Y5_FrameData_O[10] ,
    \Tile_X10Y5_FrameData_O[9] ,
    \Tile_X10Y5_FrameData_O[8] ,
    \Tile_X10Y5_FrameData_O[7] ,
    \Tile_X10Y5_FrameData_O[6] ,
    \Tile_X10Y5_FrameData_O[5] ,
    \Tile_X10Y5_FrameData_O[4] ,
    \Tile_X10Y5_FrameData_O[3] ,
    \Tile_X10Y5_FrameData_O[2] ,
    \Tile_X10Y5_FrameData_O[1] ,
    \Tile_X10Y5_FrameData_O[0] }),
    .Tile_X0Y0_FrameStrobe_O({\Tile_X10Y5_FrameStrobe_O[19] ,
    \Tile_X10Y5_FrameStrobe_O[18] ,
    \Tile_X10Y5_FrameStrobe_O[17] ,
    \Tile_X10Y5_FrameStrobe_O[16] ,
    \Tile_X10Y5_FrameStrobe_O[15] ,
    \Tile_X10Y5_FrameStrobe_O[14] ,
    \Tile_X10Y5_FrameStrobe_O[13] ,
    \Tile_X10Y5_FrameStrobe_O[12] ,
    \Tile_X10Y5_FrameStrobe_O[11] ,
    \Tile_X10Y5_FrameStrobe_O[10] ,
    \Tile_X10Y5_FrameStrobe_O[9] ,
    \Tile_X10Y5_FrameStrobe_O[8] ,
    \Tile_X10Y5_FrameStrobe_O[7] ,
    \Tile_X10Y5_FrameStrobe_O[6] ,
    \Tile_X10Y5_FrameStrobe_O[5] ,
    \Tile_X10Y5_FrameStrobe_O[4] ,
    \Tile_X10Y5_FrameStrobe_O[3] ,
    \Tile_X10Y5_FrameStrobe_O[2] ,
    \Tile_X10Y5_FrameStrobe_O[1] ,
    \Tile_X10Y5_FrameStrobe_O[0] }),
    .Tile_X0Y0_N1BEG({\Tile_X10Y5_N1BEG[3] ,
    \Tile_X10Y5_N1BEG[2] ,
    \Tile_X10Y5_N1BEG[1] ,
    \Tile_X10Y5_N1BEG[0] }),
    .Tile_X0Y0_N2BEG({\Tile_X10Y5_N2BEG[7] ,
    \Tile_X10Y5_N2BEG[6] ,
    \Tile_X10Y5_N2BEG[5] ,
    \Tile_X10Y5_N2BEG[4] ,
    \Tile_X10Y5_N2BEG[3] ,
    \Tile_X10Y5_N2BEG[2] ,
    \Tile_X10Y5_N2BEG[1] ,
    \Tile_X10Y5_N2BEG[0] }),
    .Tile_X0Y0_N2BEGb({\Tile_X10Y5_N2BEGb[7] ,
    \Tile_X10Y5_N2BEGb[6] ,
    \Tile_X10Y5_N2BEGb[5] ,
    \Tile_X10Y5_N2BEGb[4] ,
    \Tile_X10Y5_N2BEGb[3] ,
    \Tile_X10Y5_N2BEGb[2] ,
    \Tile_X10Y5_N2BEGb[1] ,
    \Tile_X10Y5_N2BEGb[0] }),
    .Tile_X0Y0_N4BEG({\Tile_X10Y5_N4BEG[15] ,
    \Tile_X10Y5_N4BEG[14] ,
    \Tile_X10Y5_N4BEG[13] ,
    \Tile_X10Y5_N4BEG[12] ,
    \Tile_X10Y5_N4BEG[11] ,
    \Tile_X10Y5_N4BEG[10] ,
    \Tile_X10Y5_N4BEG[9] ,
    \Tile_X10Y5_N4BEG[8] ,
    \Tile_X10Y5_N4BEG[7] ,
    \Tile_X10Y5_N4BEG[6] ,
    \Tile_X10Y5_N4BEG[5] ,
    \Tile_X10Y5_N4BEG[4] ,
    \Tile_X10Y5_N4BEG[3] ,
    \Tile_X10Y5_N4BEG[2] ,
    \Tile_X10Y5_N4BEG[1] ,
    \Tile_X10Y5_N4BEG[0] }),
    .Tile_X0Y0_S1END({\Tile_X10Y4_S1BEG[3] ,
    \Tile_X10Y4_S1BEG[2] ,
    \Tile_X10Y4_S1BEG[1] ,
    \Tile_X10Y4_S1BEG[0] }),
    .Tile_X0Y0_S2END({\Tile_X10Y4_S2BEGb[7] ,
    \Tile_X10Y4_S2BEGb[6] ,
    \Tile_X10Y4_S2BEGb[5] ,
    \Tile_X10Y4_S2BEGb[4] ,
    \Tile_X10Y4_S2BEGb[3] ,
    \Tile_X10Y4_S2BEGb[2] ,
    \Tile_X10Y4_S2BEGb[1] ,
    \Tile_X10Y4_S2BEGb[0] }),
    .Tile_X0Y0_S2MID({\Tile_X10Y4_S2BEG[7] ,
    \Tile_X10Y4_S2BEG[6] ,
    \Tile_X10Y4_S2BEG[5] ,
    \Tile_X10Y4_S2BEG[4] ,
    \Tile_X10Y4_S2BEG[3] ,
    \Tile_X10Y4_S2BEG[2] ,
    \Tile_X10Y4_S2BEG[1] ,
    \Tile_X10Y4_S2BEG[0] }),
    .Tile_X0Y0_S4END({\Tile_X10Y4_S4BEG[15] ,
    \Tile_X10Y4_S4BEG[14] ,
    \Tile_X10Y4_S4BEG[13] ,
    \Tile_X10Y4_S4BEG[12] ,
    \Tile_X10Y4_S4BEG[11] ,
    \Tile_X10Y4_S4BEG[10] ,
    \Tile_X10Y4_S4BEG[9] ,
    \Tile_X10Y4_S4BEG[8] ,
    \Tile_X10Y4_S4BEG[7] ,
    \Tile_X10Y4_S4BEG[6] ,
    \Tile_X10Y4_S4BEG[5] ,
    \Tile_X10Y4_S4BEG[4] ,
    \Tile_X10Y4_S4BEG[3] ,
    \Tile_X10Y4_S4BEG[2] ,
    \Tile_X10Y4_S4BEG[1] ,
    \Tile_X10Y4_S4BEG[0] }),
    .Tile_X0Y0_W1BEG({\Tile_X10Y5_W1BEG[3] ,
    \Tile_X10Y5_W1BEG[2] ,
    \Tile_X10Y5_W1BEG[1] ,
    \Tile_X10Y5_W1BEG[0] }),
    .Tile_X0Y0_W2BEG({\Tile_X10Y5_W2BEG[7] ,
    \Tile_X10Y5_W2BEG[6] ,
    \Tile_X10Y5_W2BEG[5] ,
    \Tile_X10Y5_W2BEG[4] ,
    \Tile_X10Y5_W2BEG[3] ,
    \Tile_X10Y5_W2BEG[2] ,
    \Tile_X10Y5_W2BEG[1] ,
    \Tile_X10Y5_W2BEG[0] }),
    .Tile_X0Y0_W2BEGb({\Tile_X10Y5_W2BEGb[7] ,
    \Tile_X10Y5_W2BEGb[6] ,
    \Tile_X10Y5_W2BEGb[5] ,
    \Tile_X10Y5_W2BEGb[4] ,
    \Tile_X10Y5_W2BEGb[3] ,
    \Tile_X10Y5_W2BEGb[2] ,
    \Tile_X10Y5_W2BEGb[1] ,
    \Tile_X10Y5_W2BEGb[0] }),
    .Tile_X0Y0_W6BEG({\Tile_X10Y5_W6BEG[11] ,
    \Tile_X10Y5_W6BEG[10] ,
    \Tile_X10Y5_W6BEG[9] ,
    \Tile_X10Y5_W6BEG[8] ,
    \Tile_X10Y5_W6BEG[7] ,
    \Tile_X10Y5_W6BEG[6] ,
    \Tile_X10Y5_W6BEG[5] ,
    \Tile_X10Y5_W6BEG[4] ,
    \Tile_X10Y5_W6BEG[3] ,
    \Tile_X10Y5_W6BEG[2] ,
    \Tile_X10Y5_W6BEG[1] ,
    \Tile_X10Y5_W6BEG[0] }),
    .Tile_X0Y0_WW4BEG({\Tile_X10Y5_WW4BEG[15] ,
    \Tile_X10Y5_WW4BEG[14] ,
    \Tile_X10Y5_WW4BEG[13] ,
    \Tile_X10Y5_WW4BEG[12] ,
    \Tile_X10Y5_WW4BEG[11] ,
    \Tile_X10Y5_WW4BEG[10] ,
    \Tile_X10Y5_WW4BEG[9] ,
    \Tile_X10Y5_WW4BEG[8] ,
    \Tile_X10Y5_WW4BEG[7] ,
    \Tile_X10Y5_WW4BEG[6] ,
    \Tile_X10Y5_WW4BEG[5] ,
    \Tile_X10Y5_WW4BEG[4] ,
    \Tile_X10Y5_WW4BEG[3] ,
    \Tile_X10Y5_WW4BEG[2] ,
    \Tile_X10Y5_WW4BEG[1] ,
    \Tile_X10Y5_WW4BEG[0] }),
    .Tile_X0Y1_E1END({\Tile_X9Y6_E1BEG[3] ,
    \Tile_X9Y6_E1BEG[2] ,
    \Tile_X9Y6_E1BEG[1] ,
    \Tile_X9Y6_E1BEG[0] }),
    .Tile_X0Y1_E2END({\Tile_X9Y6_E2BEGb[7] ,
    \Tile_X9Y6_E2BEGb[6] ,
    \Tile_X9Y6_E2BEGb[5] ,
    \Tile_X9Y6_E2BEGb[4] ,
    \Tile_X9Y6_E2BEGb[3] ,
    \Tile_X9Y6_E2BEGb[2] ,
    \Tile_X9Y6_E2BEGb[1] ,
    \Tile_X9Y6_E2BEGb[0] }),
    .Tile_X0Y1_E2MID({\Tile_X9Y6_E2BEG[7] ,
    \Tile_X9Y6_E2BEG[6] ,
    \Tile_X9Y6_E2BEG[5] ,
    \Tile_X9Y6_E2BEG[4] ,
    \Tile_X9Y6_E2BEG[3] ,
    \Tile_X9Y6_E2BEG[2] ,
    \Tile_X9Y6_E2BEG[1] ,
    \Tile_X9Y6_E2BEG[0] }),
    .Tile_X0Y1_E6END({\Tile_X9Y6_E6BEG[11] ,
    \Tile_X9Y6_E6BEG[10] ,
    \Tile_X9Y6_E6BEG[9] ,
    \Tile_X9Y6_E6BEG[8] ,
    \Tile_X9Y6_E6BEG[7] ,
    \Tile_X9Y6_E6BEG[6] ,
    \Tile_X9Y6_E6BEG[5] ,
    \Tile_X9Y6_E6BEG[4] ,
    \Tile_X9Y6_E6BEG[3] ,
    \Tile_X9Y6_E6BEG[2] ,
    \Tile_X9Y6_E6BEG[1] ,
    \Tile_X9Y6_E6BEG[0] }),
    .Tile_X0Y1_EE4END({\Tile_X9Y6_EE4BEG[15] ,
    \Tile_X9Y6_EE4BEG[14] ,
    \Tile_X9Y6_EE4BEG[13] ,
    \Tile_X9Y6_EE4BEG[12] ,
    \Tile_X9Y6_EE4BEG[11] ,
    \Tile_X9Y6_EE4BEG[10] ,
    \Tile_X9Y6_EE4BEG[9] ,
    \Tile_X9Y6_EE4BEG[8] ,
    \Tile_X9Y6_EE4BEG[7] ,
    \Tile_X9Y6_EE4BEG[6] ,
    \Tile_X9Y6_EE4BEG[5] ,
    \Tile_X9Y6_EE4BEG[4] ,
    \Tile_X9Y6_EE4BEG[3] ,
    \Tile_X9Y6_EE4BEG[2] ,
    \Tile_X9Y6_EE4BEG[1] ,
    \Tile_X9Y6_EE4BEG[0] }),
    .Tile_X0Y1_FrameData({\Tile_X9Y6_FrameData_O[31] ,
    \Tile_X9Y6_FrameData_O[30] ,
    \Tile_X9Y6_FrameData_O[29] ,
    \Tile_X9Y6_FrameData_O[28] ,
    \Tile_X9Y6_FrameData_O[27] ,
    \Tile_X9Y6_FrameData_O[26] ,
    \Tile_X9Y6_FrameData_O[25] ,
    \Tile_X9Y6_FrameData_O[24] ,
    \Tile_X9Y6_FrameData_O[23] ,
    \Tile_X9Y6_FrameData_O[22] ,
    \Tile_X9Y6_FrameData_O[21] ,
    \Tile_X9Y6_FrameData_O[20] ,
    \Tile_X9Y6_FrameData_O[19] ,
    \Tile_X9Y6_FrameData_O[18] ,
    \Tile_X9Y6_FrameData_O[17] ,
    \Tile_X9Y6_FrameData_O[16] ,
    \Tile_X9Y6_FrameData_O[15] ,
    \Tile_X9Y6_FrameData_O[14] ,
    \Tile_X9Y6_FrameData_O[13] ,
    \Tile_X9Y6_FrameData_O[12] ,
    \Tile_X9Y6_FrameData_O[11] ,
    \Tile_X9Y6_FrameData_O[10] ,
    \Tile_X9Y6_FrameData_O[9] ,
    \Tile_X9Y6_FrameData_O[8] ,
    \Tile_X9Y6_FrameData_O[7] ,
    \Tile_X9Y6_FrameData_O[6] ,
    \Tile_X9Y6_FrameData_O[5] ,
    \Tile_X9Y6_FrameData_O[4] ,
    \Tile_X9Y6_FrameData_O[3] ,
    \Tile_X9Y6_FrameData_O[2] ,
    \Tile_X9Y6_FrameData_O[1] ,
    \Tile_X9Y6_FrameData_O[0] }),
    .Tile_X0Y1_FrameData_O({\Tile_X10Y6_FrameData_O[31] ,
    \Tile_X10Y6_FrameData_O[30] ,
    \Tile_X10Y6_FrameData_O[29] ,
    \Tile_X10Y6_FrameData_O[28] ,
    \Tile_X10Y6_FrameData_O[27] ,
    \Tile_X10Y6_FrameData_O[26] ,
    \Tile_X10Y6_FrameData_O[25] ,
    \Tile_X10Y6_FrameData_O[24] ,
    \Tile_X10Y6_FrameData_O[23] ,
    \Tile_X10Y6_FrameData_O[22] ,
    \Tile_X10Y6_FrameData_O[21] ,
    \Tile_X10Y6_FrameData_O[20] ,
    \Tile_X10Y6_FrameData_O[19] ,
    \Tile_X10Y6_FrameData_O[18] ,
    \Tile_X10Y6_FrameData_O[17] ,
    \Tile_X10Y6_FrameData_O[16] ,
    \Tile_X10Y6_FrameData_O[15] ,
    \Tile_X10Y6_FrameData_O[14] ,
    \Tile_X10Y6_FrameData_O[13] ,
    \Tile_X10Y6_FrameData_O[12] ,
    \Tile_X10Y6_FrameData_O[11] ,
    \Tile_X10Y6_FrameData_O[10] ,
    \Tile_X10Y6_FrameData_O[9] ,
    \Tile_X10Y6_FrameData_O[8] ,
    \Tile_X10Y6_FrameData_O[7] ,
    \Tile_X10Y6_FrameData_O[6] ,
    \Tile_X10Y6_FrameData_O[5] ,
    \Tile_X10Y6_FrameData_O[4] ,
    \Tile_X10Y6_FrameData_O[3] ,
    \Tile_X10Y6_FrameData_O[2] ,
    \Tile_X10Y6_FrameData_O[1] ,
    \Tile_X10Y6_FrameData_O[0] }),
    .Tile_X0Y1_FrameStrobe({\Tile_X10Y7_FrameStrobe_O[19] ,
    \Tile_X10Y7_FrameStrobe_O[18] ,
    \Tile_X10Y7_FrameStrobe_O[17] ,
    \Tile_X10Y7_FrameStrobe_O[16] ,
    \Tile_X10Y7_FrameStrobe_O[15] ,
    \Tile_X10Y7_FrameStrobe_O[14] ,
    \Tile_X10Y7_FrameStrobe_O[13] ,
    \Tile_X10Y7_FrameStrobe_O[12] ,
    \Tile_X10Y7_FrameStrobe_O[11] ,
    \Tile_X10Y7_FrameStrobe_O[10] ,
    \Tile_X10Y7_FrameStrobe_O[9] ,
    \Tile_X10Y7_FrameStrobe_O[8] ,
    \Tile_X10Y7_FrameStrobe_O[7] ,
    \Tile_X10Y7_FrameStrobe_O[6] ,
    \Tile_X10Y7_FrameStrobe_O[5] ,
    \Tile_X10Y7_FrameStrobe_O[4] ,
    \Tile_X10Y7_FrameStrobe_O[3] ,
    \Tile_X10Y7_FrameStrobe_O[2] ,
    \Tile_X10Y7_FrameStrobe_O[1] ,
    \Tile_X10Y7_FrameStrobe_O[0] }),
    .Tile_X0Y1_N1END({\Tile_X10Y7_N1BEG[3] ,
    \Tile_X10Y7_N1BEG[2] ,
    \Tile_X10Y7_N1BEG[1] ,
    \Tile_X10Y7_N1BEG[0] }),
    .Tile_X0Y1_N2END({\Tile_X10Y7_N2BEGb[7] ,
    \Tile_X10Y7_N2BEGb[6] ,
    \Tile_X10Y7_N2BEGb[5] ,
    \Tile_X10Y7_N2BEGb[4] ,
    \Tile_X10Y7_N2BEGb[3] ,
    \Tile_X10Y7_N2BEGb[2] ,
    \Tile_X10Y7_N2BEGb[1] ,
    \Tile_X10Y7_N2BEGb[0] }),
    .Tile_X0Y1_N2MID({\Tile_X10Y7_N2BEG[7] ,
    \Tile_X10Y7_N2BEG[6] ,
    \Tile_X10Y7_N2BEG[5] ,
    \Tile_X10Y7_N2BEG[4] ,
    \Tile_X10Y7_N2BEG[3] ,
    \Tile_X10Y7_N2BEG[2] ,
    \Tile_X10Y7_N2BEG[1] ,
    \Tile_X10Y7_N2BEG[0] }),
    .Tile_X0Y1_N4END({\Tile_X10Y7_N4BEG[15] ,
    \Tile_X10Y7_N4BEG[14] ,
    \Tile_X10Y7_N4BEG[13] ,
    \Tile_X10Y7_N4BEG[12] ,
    \Tile_X10Y7_N4BEG[11] ,
    \Tile_X10Y7_N4BEG[10] ,
    \Tile_X10Y7_N4BEG[9] ,
    \Tile_X10Y7_N4BEG[8] ,
    \Tile_X10Y7_N4BEG[7] ,
    \Tile_X10Y7_N4BEG[6] ,
    \Tile_X10Y7_N4BEG[5] ,
    \Tile_X10Y7_N4BEG[4] ,
    \Tile_X10Y7_N4BEG[3] ,
    \Tile_X10Y7_N4BEG[2] ,
    \Tile_X10Y7_N4BEG[1] ,
    \Tile_X10Y7_N4BEG[0] }),
    .Tile_X0Y1_S1BEG({\Tile_X10Y6_S1BEG[3] ,
    \Tile_X10Y6_S1BEG[2] ,
    \Tile_X10Y6_S1BEG[1] ,
    \Tile_X10Y6_S1BEG[0] }),
    .Tile_X0Y1_S2BEG({\Tile_X10Y6_S2BEG[7] ,
    \Tile_X10Y6_S2BEG[6] ,
    \Tile_X10Y6_S2BEG[5] ,
    \Tile_X10Y6_S2BEG[4] ,
    \Tile_X10Y6_S2BEG[3] ,
    \Tile_X10Y6_S2BEG[2] ,
    \Tile_X10Y6_S2BEG[1] ,
    \Tile_X10Y6_S2BEG[0] }),
    .Tile_X0Y1_S2BEGb({\Tile_X10Y6_S2BEGb[7] ,
    \Tile_X10Y6_S2BEGb[6] ,
    \Tile_X10Y6_S2BEGb[5] ,
    \Tile_X10Y6_S2BEGb[4] ,
    \Tile_X10Y6_S2BEGb[3] ,
    \Tile_X10Y6_S2BEGb[2] ,
    \Tile_X10Y6_S2BEGb[1] ,
    \Tile_X10Y6_S2BEGb[0] }),
    .Tile_X0Y1_S4BEG({\Tile_X10Y6_S4BEG[15] ,
    \Tile_X10Y6_S4BEG[14] ,
    \Tile_X10Y6_S4BEG[13] ,
    \Tile_X10Y6_S4BEG[12] ,
    \Tile_X10Y6_S4BEG[11] ,
    \Tile_X10Y6_S4BEG[10] ,
    \Tile_X10Y6_S4BEG[9] ,
    \Tile_X10Y6_S4BEG[8] ,
    \Tile_X10Y6_S4BEG[7] ,
    \Tile_X10Y6_S4BEG[6] ,
    \Tile_X10Y6_S4BEG[5] ,
    \Tile_X10Y6_S4BEG[4] ,
    \Tile_X10Y6_S4BEG[3] ,
    \Tile_X10Y6_S4BEG[2] ,
    \Tile_X10Y6_S4BEG[1] ,
    \Tile_X10Y6_S4BEG[0] }),
    .Tile_X0Y1_W1BEG({\Tile_X10Y6_W1BEG[3] ,
    \Tile_X10Y6_W1BEG[2] ,
    \Tile_X10Y6_W1BEG[1] ,
    \Tile_X10Y6_W1BEG[0] }),
    .Tile_X0Y1_W2BEG({\Tile_X10Y6_W2BEG[7] ,
    \Tile_X10Y6_W2BEG[6] ,
    \Tile_X10Y6_W2BEG[5] ,
    \Tile_X10Y6_W2BEG[4] ,
    \Tile_X10Y6_W2BEG[3] ,
    \Tile_X10Y6_W2BEG[2] ,
    \Tile_X10Y6_W2BEG[1] ,
    \Tile_X10Y6_W2BEG[0] }),
    .Tile_X0Y1_W2BEGb({\Tile_X10Y6_W2BEGb[7] ,
    \Tile_X10Y6_W2BEGb[6] ,
    \Tile_X10Y6_W2BEGb[5] ,
    \Tile_X10Y6_W2BEGb[4] ,
    \Tile_X10Y6_W2BEGb[3] ,
    \Tile_X10Y6_W2BEGb[2] ,
    \Tile_X10Y6_W2BEGb[1] ,
    \Tile_X10Y6_W2BEGb[0] }),
    .Tile_X0Y1_W6BEG({\Tile_X10Y6_W6BEG[11] ,
    \Tile_X10Y6_W6BEG[10] ,
    \Tile_X10Y6_W6BEG[9] ,
    \Tile_X10Y6_W6BEG[8] ,
    \Tile_X10Y6_W6BEG[7] ,
    \Tile_X10Y6_W6BEG[6] ,
    \Tile_X10Y6_W6BEG[5] ,
    \Tile_X10Y6_W6BEG[4] ,
    \Tile_X10Y6_W6BEG[3] ,
    \Tile_X10Y6_W6BEG[2] ,
    \Tile_X10Y6_W6BEG[1] ,
    \Tile_X10Y6_W6BEG[0] }),
    .Tile_X0Y1_WW4BEG({\Tile_X10Y6_WW4BEG[15] ,
    \Tile_X10Y6_WW4BEG[14] ,
    \Tile_X10Y6_WW4BEG[13] ,
    \Tile_X10Y6_WW4BEG[12] ,
    \Tile_X10Y6_WW4BEG[11] ,
    \Tile_X10Y6_WW4BEG[10] ,
    \Tile_X10Y6_WW4BEG[9] ,
    \Tile_X10Y6_WW4BEG[8] ,
    \Tile_X10Y6_WW4BEG[7] ,
    \Tile_X10Y6_WW4BEG[6] ,
    \Tile_X10Y6_WW4BEG[5] ,
    \Tile_X10Y6_WW4BEG[4] ,
    \Tile_X10Y6_WW4BEG[3] ,
    \Tile_X10Y6_WW4BEG[2] ,
    \Tile_X10Y6_WW4BEG[1] ,
    \Tile_X10Y6_WW4BEG[0] }));
 IHP_SRAM Tile_X10Y7_IHP_SRAM (.ADDR_SRAM0(Tile_X10Y8_ADDR_SRAM0),
    .ADDR_SRAM1(Tile_X10Y8_ADDR_SRAM1),
    .ADDR_SRAM2(Tile_X10Y8_ADDR_SRAM2),
    .ADDR_SRAM3(Tile_X10Y8_ADDR_SRAM3),
    .ADDR_SRAM4(Tile_X10Y8_ADDR_SRAM4),
    .ADDR_SRAM5(Tile_X10Y8_ADDR_SRAM5),
    .ADDR_SRAM6(Tile_X10Y8_ADDR_SRAM6),
    .ADDR_SRAM7(Tile_X10Y8_ADDR_SRAM7),
    .ADDR_SRAM8(Tile_X10Y8_ADDR_SRAM8),
    .ADDR_SRAM9(Tile_X10Y8_ADDR_SRAM9),
    .BM_SRAM0(Tile_X10Y8_BM_SRAM0),
    .BM_SRAM1(Tile_X10Y8_BM_SRAM1),
    .BM_SRAM10(Tile_X10Y8_BM_SRAM10),
    .BM_SRAM11(Tile_X10Y8_BM_SRAM11),
    .BM_SRAM12(Tile_X10Y8_BM_SRAM12),
    .BM_SRAM13(Tile_X10Y8_BM_SRAM13),
    .BM_SRAM14(Tile_X10Y8_BM_SRAM14),
    .BM_SRAM15(Tile_X10Y8_BM_SRAM15),
    .BM_SRAM16(Tile_X10Y8_BM_SRAM16),
    .BM_SRAM17(Tile_X10Y8_BM_SRAM17),
    .BM_SRAM18(Tile_X10Y8_BM_SRAM18),
    .BM_SRAM19(Tile_X10Y8_BM_SRAM19),
    .BM_SRAM2(Tile_X10Y8_BM_SRAM2),
    .BM_SRAM20(Tile_X10Y8_BM_SRAM20),
    .BM_SRAM21(Tile_X10Y8_BM_SRAM21),
    .BM_SRAM22(Tile_X10Y8_BM_SRAM22),
    .BM_SRAM23(Tile_X10Y8_BM_SRAM23),
    .BM_SRAM24(Tile_X10Y8_BM_SRAM24),
    .BM_SRAM25(Tile_X10Y8_BM_SRAM25),
    .BM_SRAM26(Tile_X10Y8_BM_SRAM26),
    .BM_SRAM27(Tile_X10Y8_BM_SRAM27),
    .BM_SRAM28(Tile_X10Y8_BM_SRAM28),
    .BM_SRAM29(Tile_X10Y8_BM_SRAM29),
    .BM_SRAM3(Tile_X10Y8_BM_SRAM3),
    .BM_SRAM30(Tile_X10Y8_BM_SRAM30),
    .BM_SRAM31(Tile_X10Y8_BM_SRAM31),
    .BM_SRAM4(Tile_X10Y8_BM_SRAM4),
    .BM_SRAM5(Tile_X10Y8_BM_SRAM5),
    .BM_SRAM6(Tile_X10Y8_BM_SRAM6),
    .BM_SRAM7(Tile_X10Y8_BM_SRAM7),
    .BM_SRAM8(Tile_X10Y8_BM_SRAM8),
    .BM_SRAM9(Tile_X10Y8_BM_SRAM9),
    .CLK_SRAM(Tile_X10Y8_CLK_SRAM),
    .CONFIGURED_top(Tile_X10Y8_CONFIGURED_top),
    .DIN_SRAM0(Tile_X10Y8_DIN_SRAM0),
    .DIN_SRAM1(Tile_X10Y8_DIN_SRAM1),
    .DIN_SRAM10(Tile_X10Y8_DIN_SRAM10),
    .DIN_SRAM11(Tile_X10Y8_DIN_SRAM11),
    .DIN_SRAM12(Tile_X10Y8_DIN_SRAM12),
    .DIN_SRAM13(Tile_X10Y8_DIN_SRAM13),
    .DIN_SRAM14(Tile_X10Y8_DIN_SRAM14),
    .DIN_SRAM15(Tile_X10Y8_DIN_SRAM15),
    .DIN_SRAM16(Tile_X10Y8_DIN_SRAM16),
    .DIN_SRAM17(Tile_X10Y8_DIN_SRAM17),
    .DIN_SRAM18(Tile_X10Y8_DIN_SRAM18),
    .DIN_SRAM19(Tile_X10Y8_DIN_SRAM19),
    .DIN_SRAM2(Tile_X10Y8_DIN_SRAM2),
    .DIN_SRAM20(Tile_X10Y8_DIN_SRAM20),
    .DIN_SRAM21(Tile_X10Y8_DIN_SRAM21),
    .DIN_SRAM22(Tile_X10Y8_DIN_SRAM22),
    .DIN_SRAM23(Tile_X10Y8_DIN_SRAM23),
    .DIN_SRAM24(Tile_X10Y8_DIN_SRAM24),
    .DIN_SRAM25(Tile_X10Y8_DIN_SRAM25),
    .DIN_SRAM26(Tile_X10Y8_DIN_SRAM26),
    .DIN_SRAM27(Tile_X10Y8_DIN_SRAM27),
    .DIN_SRAM28(Tile_X10Y8_DIN_SRAM28),
    .DIN_SRAM29(Tile_X10Y8_DIN_SRAM29),
    .DIN_SRAM3(Tile_X10Y8_DIN_SRAM3),
    .DIN_SRAM30(Tile_X10Y8_DIN_SRAM30),
    .DIN_SRAM31(Tile_X10Y8_DIN_SRAM31),
    .DIN_SRAM4(Tile_X10Y8_DIN_SRAM4),
    .DIN_SRAM5(Tile_X10Y8_DIN_SRAM5),
    .DIN_SRAM6(Tile_X10Y8_DIN_SRAM6),
    .DIN_SRAM7(Tile_X10Y8_DIN_SRAM7),
    .DIN_SRAM8(Tile_X10Y8_DIN_SRAM8),
    .DIN_SRAM9(Tile_X10Y8_DIN_SRAM9),
    .DOUT_SRAM0(Tile_X10Y8_DOUT_SRAM0),
    .DOUT_SRAM1(Tile_X10Y8_DOUT_SRAM1),
    .DOUT_SRAM10(Tile_X10Y8_DOUT_SRAM10),
    .DOUT_SRAM11(Tile_X10Y8_DOUT_SRAM11),
    .DOUT_SRAM12(Tile_X10Y8_DOUT_SRAM12),
    .DOUT_SRAM13(Tile_X10Y8_DOUT_SRAM13),
    .DOUT_SRAM14(Tile_X10Y8_DOUT_SRAM14),
    .DOUT_SRAM15(Tile_X10Y8_DOUT_SRAM15),
    .DOUT_SRAM16(Tile_X10Y8_DOUT_SRAM16),
    .DOUT_SRAM17(Tile_X10Y8_DOUT_SRAM17),
    .DOUT_SRAM18(Tile_X10Y8_DOUT_SRAM18),
    .DOUT_SRAM19(Tile_X10Y8_DOUT_SRAM19),
    .DOUT_SRAM2(Tile_X10Y8_DOUT_SRAM2),
    .DOUT_SRAM20(Tile_X10Y8_DOUT_SRAM20),
    .DOUT_SRAM21(Tile_X10Y8_DOUT_SRAM21),
    .DOUT_SRAM22(Tile_X10Y8_DOUT_SRAM22),
    .DOUT_SRAM23(Tile_X10Y8_DOUT_SRAM23),
    .DOUT_SRAM24(Tile_X10Y8_DOUT_SRAM24),
    .DOUT_SRAM25(Tile_X10Y8_DOUT_SRAM25),
    .DOUT_SRAM26(Tile_X10Y8_DOUT_SRAM26),
    .DOUT_SRAM27(Tile_X10Y8_DOUT_SRAM27),
    .DOUT_SRAM28(Tile_X10Y8_DOUT_SRAM28),
    .DOUT_SRAM29(Tile_X10Y8_DOUT_SRAM29),
    .DOUT_SRAM3(Tile_X10Y8_DOUT_SRAM3),
    .DOUT_SRAM30(Tile_X10Y8_DOUT_SRAM30),
    .DOUT_SRAM31(Tile_X10Y8_DOUT_SRAM31),
    .DOUT_SRAM4(Tile_X10Y8_DOUT_SRAM4),
    .DOUT_SRAM5(Tile_X10Y8_DOUT_SRAM5),
    .DOUT_SRAM6(Tile_X10Y8_DOUT_SRAM6),
    .DOUT_SRAM7(Tile_X10Y8_DOUT_SRAM7),
    .DOUT_SRAM8(Tile_X10Y8_DOUT_SRAM8),
    .DOUT_SRAM9(Tile_X10Y8_DOUT_SRAM9),
    .MEN_SRAM(Tile_X10Y8_MEN_SRAM),
    .REN_SRAM(Tile_X10Y8_REN_SRAM),
    .TIE_HIGH_SRAM(Tile_X10Y8_TIE_HIGH_SRAM),
    .TIE_LOW_SRAM(Tile_X10Y8_TIE_LOW_SRAM),
    .Tile_X0Y0_UserCLKo(Tile_X10Y7_UserCLKo),
    .Tile_X0Y1_UserCLK(Tile_X10Y9_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .WEN_SRAM(Tile_X10Y8_WEN_SRAM),
    .Tile_X0Y0_E1END({\Tile_X9Y7_E1BEG[3] ,
    \Tile_X9Y7_E1BEG[2] ,
    \Tile_X9Y7_E1BEG[1] ,
    \Tile_X9Y7_E1BEG[0] }),
    .Tile_X0Y0_E2END({\Tile_X9Y7_E2BEGb[7] ,
    \Tile_X9Y7_E2BEGb[6] ,
    \Tile_X9Y7_E2BEGb[5] ,
    \Tile_X9Y7_E2BEGb[4] ,
    \Tile_X9Y7_E2BEGb[3] ,
    \Tile_X9Y7_E2BEGb[2] ,
    \Tile_X9Y7_E2BEGb[1] ,
    \Tile_X9Y7_E2BEGb[0] }),
    .Tile_X0Y0_E2MID({\Tile_X9Y7_E2BEG[7] ,
    \Tile_X9Y7_E2BEG[6] ,
    \Tile_X9Y7_E2BEG[5] ,
    \Tile_X9Y7_E2BEG[4] ,
    \Tile_X9Y7_E2BEG[3] ,
    \Tile_X9Y7_E2BEG[2] ,
    \Tile_X9Y7_E2BEG[1] ,
    \Tile_X9Y7_E2BEG[0] }),
    .Tile_X0Y0_E6END({\Tile_X9Y7_E6BEG[11] ,
    \Tile_X9Y7_E6BEG[10] ,
    \Tile_X9Y7_E6BEG[9] ,
    \Tile_X9Y7_E6BEG[8] ,
    \Tile_X9Y7_E6BEG[7] ,
    \Tile_X9Y7_E6BEG[6] ,
    \Tile_X9Y7_E6BEG[5] ,
    \Tile_X9Y7_E6BEG[4] ,
    \Tile_X9Y7_E6BEG[3] ,
    \Tile_X9Y7_E6BEG[2] ,
    \Tile_X9Y7_E6BEG[1] ,
    \Tile_X9Y7_E6BEG[0] }),
    .Tile_X0Y0_EE4END({\Tile_X9Y7_EE4BEG[15] ,
    \Tile_X9Y7_EE4BEG[14] ,
    \Tile_X9Y7_EE4BEG[13] ,
    \Tile_X9Y7_EE4BEG[12] ,
    \Tile_X9Y7_EE4BEG[11] ,
    \Tile_X9Y7_EE4BEG[10] ,
    \Tile_X9Y7_EE4BEG[9] ,
    \Tile_X9Y7_EE4BEG[8] ,
    \Tile_X9Y7_EE4BEG[7] ,
    \Tile_X9Y7_EE4BEG[6] ,
    \Tile_X9Y7_EE4BEG[5] ,
    \Tile_X9Y7_EE4BEG[4] ,
    \Tile_X9Y7_EE4BEG[3] ,
    \Tile_X9Y7_EE4BEG[2] ,
    \Tile_X9Y7_EE4BEG[1] ,
    \Tile_X9Y7_EE4BEG[0] }),
    .Tile_X0Y0_FrameData({\Tile_X9Y7_FrameData_O[31] ,
    \Tile_X9Y7_FrameData_O[30] ,
    \Tile_X9Y7_FrameData_O[29] ,
    \Tile_X9Y7_FrameData_O[28] ,
    \Tile_X9Y7_FrameData_O[27] ,
    \Tile_X9Y7_FrameData_O[26] ,
    \Tile_X9Y7_FrameData_O[25] ,
    \Tile_X9Y7_FrameData_O[24] ,
    \Tile_X9Y7_FrameData_O[23] ,
    \Tile_X9Y7_FrameData_O[22] ,
    \Tile_X9Y7_FrameData_O[21] ,
    \Tile_X9Y7_FrameData_O[20] ,
    \Tile_X9Y7_FrameData_O[19] ,
    \Tile_X9Y7_FrameData_O[18] ,
    \Tile_X9Y7_FrameData_O[17] ,
    \Tile_X9Y7_FrameData_O[16] ,
    \Tile_X9Y7_FrameData_O[15] ,
    \Tile_X9Y7_FrameData_O[14] ,
    \Tile_X9Y7_FrameData_O[13] ,
    \Tile_X9Y7_FrameData_O[12] ,
    \Tile_X9Y7_FrameData_O[11] ,
    \Tile_X9Y7_FrameData_O[10] ,
    \Tile_X9Y7_FrameData_O[9] ,
    \Tile_X9Y7_FrameData_O[8] ,
    \Tile_X9Y7_FrameData_O[7] ,
    \Tile_X9Y7_FrameData_O[6] ,
    \Tile_X9Y7_FrameData_O[5] ,
    \Tile_X9Y7_FrameData_O[4] ,
    \Tile_X9Y7_FrameData_O[3] ,
    \Tile_X9Y7_FrameData_O[2] ,
    \Tile_X9Y7_FrameData_O[1] ,
    \Tile_X9Y7_FrameData_O[0] }),
    .Tile_X0Y0_FrameData_O({\Tile_X10Y7_FrameData_O[31] ,
    \Tile_X10Y7_FrameData_O[30] ,
    \Tile_X10Y7_FrameData_O[29] ,
    \Tile_X10Y7_FrameData_O[28] ,
    \Tile_X10Y7_FrameData_O[27] ,
    \Tile_X10Y7_FrameData_O[26] ,
    \Tile_X10Y7_FrameData_O[25] ,
    \Tile_X10Y7_FrameData_O[24] ,
    \Tile_X10Y7_FrameData_O[23] ,
    \Tile_X10Y7_FrameData_O[22] ,
    \Tile_X10Y7_FrameData_O[21] ,
    \Tile_X10Y7_FrameData_O[20] ,
    \Tile_X10Y7_FrameData_O[19] ,
    \Tile_X10Y7_FrameData_O[18] ,
    \Tile_X10Y7_FrameData_O[17] ,
    \Tile_X10Y7_FrameData_O[16] ,
    \Tile_X10Y7_FrameData_O[15] ,
    \Tile_X10Y7_FrameData_O[14] ,
    \Tile_X10Y7_FrameData_O[13] ,
    \Tile_X10Y7_FrameData_O[12] ,
    \Tile_X10Y7_FrameData_O[11] ,
    \Tile_X10Y7_FrameData_O[10] ,
    \Tile_X10Y7_FrameData_O[9] ,
    \Tile_X10Y7_FrameData_O[8] ,
    \Tile_X10Y7_FrameData_O[7] ,
    \Tile_X10Y7_FrameData_O[6] ,
    \Tile_X10Y7_FrameData_O[5] ,
    \Tile_X10Y7_FrameData_O[4] ,
    \Tile_X10Y7_FrameData_O[3] ,
    \Tile_X10Y7_FrameData_O[2] ,
    \Tile_X10Y7_FrameData_O[1] ,
    \Tile_X10Y7_FrameData_O[0] }),
    .Tile_X0Y0_FrameStrobe_O({\Tile_X10Y7_FrameStrobe_O[19] ,
    \Tile_X10Y7_FrameStrobe_O[18] ,
    \Tile_X10Y7_FrameStrobe_O[17] ,
    \Tile_X10Y7_FrameStrobe_O[16] ,
    \Tile_X10Y7_FrameStrobe_O[15] ,
    \Tile_X10Y7_FrameStrobe_O[14] ,
    \Tile_X10Y7_FrameStrobe_O[13] ,
    \Tile_X10Y7_FrameStrobe_O[12] ,
    \Tile_X10Y7_FrameStrobe_O[11] ,
    \Tile_X10Y7_FrameStrobe_O[10] ,
    \Tile_X10Y7_FrameStrobe_O[9] ,
    \Tile_X10Y7_FrameStrobe_O[8] ,
    \Tile_X10Y7_FrameStrobe_O[7] ,
    \Tile_X10Y7_FrameStrobe_O[6] ,
    \Tile_X10Y7_FrameStrobe_O[5] ,
    \Tile_X10Y7_FrameStrobe_O[4] ,
    \Tile_X10Y7_FrameStrobe_O[3] ,
    \Tile_X10Y7_FrameStrobe_O[2] ,
    \Tile_X10Y7_FrameStrobe_O[1] ,
    \Tile_X10Y7_FrameStrobe_O[0] }),
    .Tile_X0Y0_N1BEG({\Tile_X10Y7_N1BEG[3] ,
    \Tile_X10Y7_N1BEG[2] ,
    \Tile_X10Y7_N1BEG[1] ,
    \Tile_X10Y7_N1BEG[0] }),
    .Tile_X0Y0_N2BEG({\Tile_X10Y7_N2BEG[7] ,
    \Tile_X10Y7_N2BEG[6] ,
    \Tile_X10Y7_N2BEG[5] ,
    \Tile_X10Y7_N2BEG[4] ,
    \Tile_X10Y7_N2BEG[3] ,
    \Tile_X10Y7_N2BEG[2] ,
    \Tile_X10Y7_N2BEG[1] ,
    \Tile_X10Y7_N2BEG[0] }),
    .Tile_X0Y0_N2BEGb({\Tile_X10Y7_N2BEGb[7] ,
    \Tile_X10Y7_N2BEGb[6] ,
    \Tile_X10Y7_N2BEGb[5] ,
    \Tile_X10Y7_N2BEGb[4] ,
    \Tile_X10Y7_N2BEGb[3] ,
    \Tile_X10Y7_N2BEGb[2] ,
    \Tile_X10Y7_N2BEGb[1] ,
    \Tile_X10Y7_N2BEGb[0] }),
    .Tile_X0Y0_N4BEG({\Tile_X10Y7_N4BEG[15] ,
    \Tile_X10Y7_N4BEG[14] ,
    \Tile_X10Y7_N4BEG[13] ,
    \Tile_X10Y7_N4BEG[12] ,
    \Tile_X10Y7_N4BEG[11] ,
    \Tile_X10Y7_N4BEG[10] ,
    \Tile_X10Y7_N4BEG[9] ,
    \Tile_X10Y7_N4BEG[8] ,
    \Tile_X10Y7_N4BEG[7] ,
    \Tile_X10Y7_N4BEG[6] ,
    \Tile_X10Y7_N4BEG[5] ,
    \Tile_X10Y7_N4BEG[4] ,
    \Tile_X10Y7_N4BEG[3] ,
    \Tile_X10Y7_N4BEG[2] ,
    \Tile_X10Y7_N4BEG[1] ,
    \Tile_X10Y7_N4BEG[0] }),
    .Tile_X0Y0_S1END({\Tile_X10Y6_S1BEG[3] ,
    \Tile_X10Y6_S1BEG[2] ,
    \Tile_X10Y6_S1BEG[1] ,
    \Tile_X10Y6_S1BEG[0] }),
    .Tile_X0Y0_S2END({\Tile_X10Y6_S2BEGb[7] ,
    \Tile_X10Y6_S2BEGb[6] ,
    \Tile_X10Y6_S2BEGb[5] ,
    \Tile_X10Y6_S2BEGb[4] ,
    \Tile_X10Y6_S2BEGb[3] ,
    \Tile_X10Y6_S2BEGb[2] ,
    \Tile_X10Y6_S2BEGb[1] ,
    \Tile_X10Y6_S2BEGb[0] }),
    .Tile_X0Y0_S2MID({\Tile_X10Y6_S2BEG[7] ,
    \Tile_X10Y6_S2BEG[6] ,
    \Tile_X10Y6_S2BEG[5] ,
    \Tile_X10Y6_S2BEG[4] ,
    \Tile_X10Y6_S2BEG[3] ,
    \Tile_X10Y6_S2BEG[2] ,
    \Tile_X10Y6_S2BEG[1] ,
    \Tile_X10Y6_S2BEG[0] }),
    .Tile_X0Y0_S4END({\Tile_X10Y6_S4BEG[15] ,
    \Tile_X10Y6_S4BEG[14] ,
    \Tile_X10Y6_S4BEG[13] ,
    \Tile_X10Y6_S4BEG[12] ,
    \Tile_X10Y6_S4BEG[11] ,
    \Tile_X10Y6_S4BEG[10] ,
    \Tile_X10Y6_S4BEG[9] ,
    \Tile_X10Y6_S4BEG[8] ,
    \Tile_X10Y6_S4BEG[7] ,
    \Tile_X10Y6_S4BEG[6] ,
    \Tile_X10Y6_S4BEG[5] ,
    \Tile_X10Y6_S4BEG[4] ,
    \Tile_X10Y6_S4BEG[3] ,
    \Tile_X10Y6_S4BEG[2] ,
    \Tile_X10Y6_S4BEG[1] ,
    \Tile_X10Y6_S4BEG[0] }),
    .Tile_X0Y0_W1BEG({\Tile_X10Y7_W1BEG[3] ,
    \Tile_X10Y7_W1BEG[2] ,
    \Tile_X10Y7_W1BEG[1] ,
    \Tile_X10Y7_W1BEG[0] }),
    .Tile_X0Y0_W2BEG({\Tile_X10Y7_W2BEG[7] ,
    \Tile_X10Y7_W2BEG[6] ,
    \Tile_X10Y7_W2BEG[5] ,
    \Tile_X10Y7_W2BEG[4] ,
    \Tile_X10Y7_W2BEG[3] ,
    \Tile_X10Y7_W2BEG[2] ,
    \Tile_X10Y7_W2BEG[1] ,
    \Tile_X10Y7_W2BEG[0] }),
    .Tile_X0Y0_W2BEGb({\Tile_X10Y7_W2BEGb[7] ,
    \Tile_X10Y7_W2BEGb[6] ,
    \Tile_X10Y7_W2BEGb[5] ,
    \Tile_X10Y7_W2BEGb[4] ,
    \Tile_X10Y7_W2BEGb[3] ,
    \Tile_X10Y7_W2BEGb[2] ,
    \Tile_X10Y7_W2BEGb[1] ,
    \Tile_X10Y7_W2BEGb[0] }),
    .Tile_X0Y0_W6BEG({\Tile_X10Y7_W6BEG[11] ,
    \Tile_X10Y7_W6BEG[10] ,
    \Tile_X10Y7_W6BEG[9] ,
    \Tile_X10Y7_W6BEG[8] ,
    \Tile_X10Y7_W6BEG[7] ,
    \Tile_X10Y7_W6BEG[6] ,
    \Tile_X10Y7_W6BEG[5] ,
    \Tile_X10Y7_W6BEG[4] ,
    \Tile_X10Y7_W6BEG[3] ,
    \Tile_X10Y7_W6BEG[2] ,
    \Tile_X10Y7_W6BEG[1] ,
    \Tile_X10Y7_W6BEG[0] }),
    .Tile_X0Y0_WW4BEG({\Tile_X10Y7_WW4BEG[15] ,
    \Tile_X10Y7_WW4BEG[14] ,
    \Tile_X10Y7_WW4BEG[13] ,
    \Tile_X10Y7_WW4BEG[12] ,
    \Tile_X10Y7_WW4BEG[11] ,
    \Tile_X10Y7_WW4BEG[10] ,
    \Tile_X10Y7_WW4BEG[9] ,
    \Tile_X10Y7_WW4BEG[8] ,
    \Tile_X10Y7_WW4BEG[7] ,
    \Tile_X10Y7_WW4BEG[6] ,
    \Tile_X10Y7_WW4BEG[5] ,
    \Tile_X10Y7_WW4BEG[4] ,
    \Tile_X10Y7_WW4BEG[3] ,
    \Tile_X10Y7_WW4BEG[2] ,
    \Tile_X10Y7_WW4BEG[1] ,
    \Tile_X10Y7_WW4BEG[0] }),
    .Tile_X0Y1_E1END({\Tile_X9Y8_E1BEG[3] ,
    \Tile_X9Y8_E1BEG[2] ,
    \Tile_X9Y8_E1BEG[1] ,
    \Tile_X9Y8_E1BEG[0] }),
    .Tile_X0Y1_E2END({\Tile_X9Y8_E2BEGb[7] ,
    \Tile_X9Y8_E2BEGb[6] ,
    \Tile_X9Y8_E2BEGb[5] ,
    \Tile_X9Y8_E2BEGb[4] ,
    \Tile_X9Y8_E2BEGb[3] ,
    \Tile_X9Y8_E2BEGb[2] ,
    \Tile_X9Y8_E2BEGb[1] ,
    \Tile_X9Y8_E2BEGb[0] }),
    .Tile_X0Y1_E2MID({\Tile_X9Y8_E2BEG[7] ,
    \Tile_X9Y8_E2BEG[6] ,
    \Tile_X9Y8_E2BEG[5] ,
    \Tile_X9Y8_E2BEG[4] ,
    \Tile_X9Y8_E2BEG[3] ,
    \Tile_X9Y8_E2BEG[2] ,
    \Tile_X9Y8_E2BEG[1] ,
    \Tile_X9Y8_E2BEG[0] }),
    .Tile_X0Y1_E6END({\Tile_X9Y8_E6BEG[11] ,
    \Tile_X9Y8_E6BEG[10] ,
    \Tile_X9Y8_E6BEG[9] ,
    \Tile_X9Y8_E6BEG[8] ,
    \Tile_X9Y8_E6BEG[7] ,
    \Tile_X9Y8_E6BEG[6] ,
    \Tile_X9Y8_E6BEG[5] ,
    \Tile_X9Y8_E6BEG[4] ,
    \Tile_X9Y8_E6BEG[3] ,
    \Tile_X9Y8_E6BEG[2] ,
    \Tile_X9Y8_E6BEG[1] ,
    \Tile_X9Y8_E6BEG[0] }),
    .Tile_X0Y1_EE4END({\Tile_X9Y8_EE4BEG[15] ,
    \Tile_X9Y8_EE4BEG[14] ,
    \Tile_X9Y8_EE4BEG[13] ,
    \Tile_X9Y8_EE4BEG[12] ,
    \Tile_X9Y8_EE4BEG[11] ,
    \Tile_X9Y8_EE4BEG[10] ,
    \Tile_X9Y8_EE4BEG[9] ,
    \Tile_X9Y8_EE4BEG[8] ,
    \Tile_X9Y8_EE4BEG[7] ,
    \Tile_X9Y8_EE4BEG[6] ,
    \Tile_X9Y8_EE4BEG[5] ,
    \Tile_X9Y8_EE4BEG[4] ,
    \Tile_X9Y8_EE4BEG[3] ,
    \Tile_X9Y8_EE4BEG[2] ,
    \Tile_X9Y8_EE4BEG[1] ,
    \Tile_X9Y8_EE4BEG[0] }),
    .Tile_X0Y1_FrameData({\Tile_X9Y8_FrameData_O[31] ,
    \Tile_X9Y8_FrameData_O[30] ,
    \Tile_X9Y8_FrameData_O[29] ,
    \Tile_X9Y8_FrameData_O[28] ,
    \Tile_X9Y8_FrameData_O[27] ,
    \Tile_X9Y8_FrameData_O[26] ,
    \Tile_X9Y8_FrameData_O[25] ,
    \Tile_X9Y8_FrameData_O[24] ,
    \Tile_X9Y8_FrameData_O[23] ,
    \Tile_X9Y8_FrameData_O[22] ,
    \Tile_X9Y8_FrameData_O[21] ,
    \Tile_X9Y8_FrameData_O[20] ,
    \Tile_X9Y8_FrameData_O[19] ,
    \Tile_X9Y8_FrameData_O[18] ,
    \Tile_X9Y8_FrameData_O[17] ,
    \Tile_X9Y8_FrameData_O[16] ,
    \Tile_X9Y8_FrameData_O[15] ,
    \Tile_X9Y8_FrameData_O[14] ,
    \Tile_X9Y8_FrameData_O[13] ,
    \Tile_X9Y8_FrameData_O[12] ,
    \Tile_X9Y8_FrameData_O[11] ,
    \Tile_X9Y8_FrameData_O[10] ,
    \Tile_X9Y8_FrameData_O[9] ,
    \Tile_X9Y8_FrameData_O[8] ,
    \Tile_X9Y8_FrameData_O[7] ,
    \Tile_X9Y8_FrameData_O[6] ,
    \Tile_X9Y8_FrameData_O[5] ,
    \Tile_X9Y8_FrameData_O[4] ,
    \Tile_X9Y8_FrameData_O[3] ,
    \Tile_X9Y8_FrameData_O[2] ,
    \Tile_X9Y8_FrameData_O[1] ,
    \Tile_X9Y8_FrameData_O[0] }),
    .Tile_X0Y1_FrameData_O({\Tile_X10Y8_FrameData_O[31] ,
    \Tile_X10Y8_FrameData_O[30] ,
    \Tile_X10Y8_FrameData_O[29] ,
    \Tile_X10Y8_FrameData_O[28] ,
    \Tile_X10Y8_FrameData_O[27] ,
    \Tile_X10Y8_FrameData_O[26] ,
    \Tile_X10Y8_FrameData_O[25] ,
    \Tile_X10Y8_FrameData_O[24] ,
    \Tile_X10Y8_FrameData_O[23] ,
    \Tile_X10Y8_FrameData_O[22] ,
    \Tile_X10Y8_FrameData_O[21] ,
    \Tile_X10Y8_FrameData_O[20] ,
    \Tile_X10Y8_FrameData_O[19] ,
    \Tile_X10Y8_FrameData_O[18] ,
    \Tile_X10Y8_FrameData_O[17] ,
    \Tile_X10Y8_FrameData_O[16] ,
    \Tile_X10Y8_FrameData_O[15] ,
    \Tile_X10Y8_FrameData_O[14] ,
    \Tile_X10Y8_FrameData_O[13] ,
    \Tile_X10Y8_FrameData_O[12] ,
    \Tile_X10Y8_FrameData_O[11] ,
    \Tile_X10Y8_FrameData_O[10] ,
    \Tile_X10Y8_FrameData_O[9] ,
    \Tile_X10Y8_FrameData_O[8] ,
    \Tile_X10Y8_FrameData_O[7] ,
    \Tile_X10Y8_FrameData_O[6] ,
    \Tile_X10Y8_FrameData_O[5] ,
    \Tile_X10Y8_FrameData_O[4] ,
    \Tile_X10Y8_FrameData_O[3] ,
    \Tile_X10Y8_FrameData_O[2] ,
    \Tile_X10Y8_FrameData_O[1] ,
    \Tile_X10Y8_FrameData_O[0] }),
    .Tile_X0Y1_FrameStrobe({\Tile_X10Y9_FrameStrobe_O[19] ,
    \Tile_X10Y9_FrameStrobe_O[18] ,
    \Tile_X10Y9_FrameStrobe_O[17] ,
    \Tile_X10Y9_FrameStrobe_O[16] ,
    \Tile_X10Y9_FrameStrobe_O[15] ,
    \Tile_X10Y9_FrameStrobe_O[14] ,
    \Tile_X10Y9_FrameStrobe_O[13] ,
    \Tile_X10Y9_FrameStrobe_O[12] ,
    \Tile_X10Y9_FrameStrobe_O[11] ,
    \Tile_X10Y9_FrameStrobe_O[10] ,
    \Tile_X10Y9_FrameStrobe_O[9] ,
    \Tile_X10Y9_FrameStrobe_O[8] ,
    \Tile_X10Y9_FrameStrobe_O[7] ,
    \Tile_X10Y9_FrameStrobe_O[6] ,
    \Tile_X10Y9_FrameStrobe_O[5] ,
    \Tile_X10Y9_FrameStrobe_O[4] ,
    \Tile_X10Y9_FrameStrobe_O[3] ,
    \Tile_X10Y9_FrameStrobe_O[2] ,
    \Tile_X10Y9_FrameStrobe_O[1] ,
    \Tile_X10Y9_FrameStrobe_O[0] }),
    .Tile_X0Y1_N1END({\Tile_X10Y9_N1BEG[3] ,
    \Tile_X10Y9_N1BEG[2] ,
    \Tile_X10Y9_N1BEG[1] ,
    \Tile_X10Y9_N1BEG[0] }),
    .Tile_X0Y1_N2END({\Tile_X10Y9_N2BEGb[7] ,
    \Tile_X10Y9_N2BEGb[6] ,
    \Tile_X10Y9_N2BEGb[5] ,
    \Tile_X10Y9_N2BEGb[4] ,
    \Tile_X10Y9_N2BEGb[3] ,
    \Tile_X10Y9_N2BEGb[2] ,
    \Tile_X10Y9_N2BEGb[1] ,
    \Tile_X10Y9_N2BEGb[0] }),
    .Tile_X0Y1_N2MID({\Tile_X10Y9_N2BEG[7] ,
    \Tile_X10Y9_N2BEG[6] ,
    \Tile_X10Y9_N2BEG[5] ,
    \Tile_X10Y9_N2BEG[4] ,
    \Tile_X10Y9_N2BEG[3] ,
    \Tile_X10Y9_N2BEG[2] ,
    \Tile_X10Y9_N2BEG[1] ,
    \Tile_X10Y9_N2BEG[0] }),
    .Tile_X0Y1_N4END({\Tile_X10Y9_N4BEG[15] ,
    \Tile_X10Y9_N4BEG[14] ,
    \Tile_X10Y9_N4BEG[13] ,
    \Tile_X10Y9_N4BEG[12] ,
    \Tile_X10Y9_N4BEG[11] ,
    \Tile_X10Y9_N4BEG[10] ,
    \Tile_X10Y9_N4BEG[9] ,
    \Tile_X10Y9_N4BEG[8] ,
    \Tile_X10Y9_N4BEG[7] ,
    \Tile_X10Y9_N4BEG[6] ,
    \Tile_X10Y9_N4BEG[5] ,
    \Tile_X10Y9_N4BEG[4] ,
    \Tile_X10Y9_N4BEG[3] ,
    \Tile_X10Y9_N4BEG[2] ,
    \Tile_X10Y9_N4BEG[1] ,
    \Tile_X10Y9_N4BEG[0] }),
    .Tile_X0Y1_S1BEG({\Tile_X10Y8_S1BEG[3] ,
    \Tile_X10Y8_S1BEG[2] ,
    \Tile_X10Y8_S1BEG[1] ,
    \Tile_X10Y8_S1BEG[0] }),
    .Tile_X0Y1_S2BEG({\Tile_X10Y8_S2BEG[7] ,
    \Tile_X10Y8_S2BEG[6] ,
    \Tile_X10Y8_S2BEG[5] ,
    \Tile_X10Y8_S2BEG[4] ,
    \Tile_X10Y8_S2BEG[3] ,
    \Tile_X10Y8_S2BEG[2] ,
    \Tile_X10Y8_S2BEG[1] ,
    \Tile_X10Y8_S2BEG[0] }),
    .Tile_X0Y1_S2BEGb({\Tile_X10Y8_S2BEGb[7] ,
    \Tile_X10Y8_S2BEGb[6] ,
    \Tile_X10Y8_S2BEGb[5] ,
    \Tile_X10Y8_S2BEGb[4] ,
    \Tile_X10Y8_S2BEGb[3] ,
    \Tile_X10Y8_S2BEGb[2] ,
    \Tile_X10Y8_S2BEGb[1] ,
    \Tile_X10Y8_S2BEGb[0] }),
    .Tile_X0Y1_S4BEG({\Tile_X10Y8_S4BEG[15] ,
    \Tile_X10Y8_S4BEG[14] ,
    \Tile_X10Y8_S4BEG[13] ,
    \Tile_X10Y8_S4BEG[12] ,
    \Tile_X10Y8_S4BEG[11] ,
    \Tile_X10Y8_S4BEG[10] ,
    \Tile_X10Y8_S4BEG[9] ,
    \Tile_X10Y8_S4BEG[8] ,
    \Tile_X10Y8_S4BEG[7] ,
    \Tile_X10Y8_S4BEG[6] ,
    \Tile_X10Y8_S4BEG[5] ,
    \Tile_X10Y8_S4BEG[4] ,
    \Tile_X10Y8_S4BEG[3] ,
    \Tile_X10Y8_S4BEG[2] ,
    \Tile_X10Y8_S4BEG[1] ,
    \Tile_X10Y8_S4BEG[0] }),
    .Tile_X0Y1_W1BEG({\Tile_X10Y8_W1BEG[3] ,
    \Tile_X10Y8_W1BEG[2] ,
    \Tile_X10Y8_W1BEG[1] ,
    \Tile_X10Y8_W1BEG[0] }),
    .Tile_X0Y1_W2BEG({\Tile_X10Y8_W2BEG[7] ,
    \Tile_X10Y8_W2BEG[6] ,
    \Tile_X10Y8_W2BEG[5] ,
    \Tile_X10Y8_W2BEG[4] ,
    \Tile_X10Y8_W2BEG[3] ,
    \Tile_X10Y8_W2BEG[2] ,
    \Tile_X10Y8_W2BEG[1] ,
    \Tile_X10Y8_W2BEG[0] }),
    .Tile_X0Y1_W2BEGb({\Tile_X10Y8_W2BEGb[7] ,
    \Tile_X10Y8_W2BEGb[6] ,
    \Tile_X10Y8_W2BEGb[5] ,
    \Tile_X10Y8_W2BEGb[4] ,
    \Tile_X10Y8_W2BEGb[3] ,
    \Tile_X10Y8_W2BEGb[2] ,
    \Tile_X10Y8_W2BEGb[1] ,
    \Tile_X10Y8_W2BEGb[0] }),
    .Tile_X0Y1_W6BEG({\Tile_X10Y8_W6BEG[11] ,
    \Tile_X10Y8_W6BEG[10] ,
    \Tile_X10Y8_W6BEG[9] ,
    \Tile_X10Y8_W6BEG[8] ,
    \Tile_X10Y8_W6BEG[7] ,
    \Tile_X10Y8_W6BEG[6] ,
    \Tile_X10Y8_W6BEG[5] ,
    \Tile_X10Y8_W6BEG[4] ,
    \Tile_X10Y8_W6BEG[3] ,
    \Tile_X10Y8_W6BEG[2] ,
    \Tile_X10Y8_W6BEG[1] ,
    \Tile_X10Y8_W6BEG[0] }),
    .Tile_X0Y1_WW4BEG({\Tile_X10Y8_WW4BEG[15] ,
    \Tile_X10Y8_WW4BEG[14] ,
    \Tile_X10Y8_WW4BEG[13] ,
    \Tile_X10Y8_WW4BEG[12] ,
    \Tile_X10Y8_WW4BEG[11] ,
    \Tile_X10Y8_WW4BEG[10] ,
    \Tile_X10Y8_WW4BEG[9] ,
    \Tile_X10Y8_WW4BEG[8] ,
    \Tile_X10Y8_WW4BEG[7] ,
    \Tile_X10Y8_WW4BEG[6] ,
    \Tile_X10Y8_WW4BEG[5] ,
    \Tile_X10Y8_WW4BEG[4] ,
    \Tile_X10Y8_WW4BEG[3] ,
    \Tile_X10Y8_WW4BEG[2] ,
    \Tile_X10Y8_WW4BEG[1] ,
    \Tile_X10Y8_WW4BEG[0] }));
 IHP_SRAM Tile_X10Y9_IHP_SRAM (.ADDR_SRAM0(Tile_X10Y10_ADDR_SRAM0),
    .ADDR_SRAM1(Tile_X10Y10_ADDR_SRAM1),
    .ADDR_SRAM2(Tile_X10Y10_ADDR_SRAM2),
    .ADDR_SRAM3(Tile_X10Y10_ADDR_SRAM3),
    .ADDR_SRAM4(Tile_X10Y10_ADDR_SRAM4),
    .ADDR_SRAM5(Tile_X10Y10_ADDR_SRAM5),
    .ADDR_SRAM6(Tile_X10Y10_ADDR_SRAM6),
    .ADDR_SRAM7(Tile_X10Y10_ADDR_SRAM7),
    .ADDR_SRAM8(Tile_X10Y10_ADDR_SRAM8),
    .ADDR_SRAM9(Tile_X10Y10_ADDR_SRAM9),
    .BM_SRAM0(Tile_X10Y10_BM_SRAM0),
    .BM_SRAM1(Tile_X10Y10_BM_SRAM1),
    .BM_SRAM10(Tile_X10Y10_BM_SRAM10),
    .BM_SRAM11(Tile_X10Y10_BM_SRAM11),
    .BM_SRAM12(Tile_X10Y10_BM_SRAM12),
    .BM_SRAM13(Tile_X10Y10_BM_SRAM13),
    .BM_SRAM14(Tile_X10Y10_BM_SRAM14),
    .BM_SRAM15(Tile_X10Y10_BM_SRAM15),
    .BM_SRAM16(Tile_X10Y10_BM_SRAM16),
    .BM_SRAM17(Tile_X10Y10_BM_SRAM17),
    .BM_SRAM18(Tile_X10Y10_BM_SRAM18),
    .BM_SRAM19(Tile_X10Y10_BM_SRAM19),
    .BM_SRAM2(Tile_X10Y10_BM_SRAM2),
    .BM_SRAM20(Tile_X10Y10_BM_SRAM20),
    .BM_SRAM21(Tile_X10Y10_BM_SRAM21),
    .BM_SRAM22(Tile_X10Y10_BM_SRAM22),
    .BM_SRAM23(Tile_X10Y10_BM_SRAM23),
    .BM_SRAM24(Tile_X10Y10_BM_SRAM24),
    .BM_SRAM25(Tile_X10Y10_BM_SRAM25),
    .BM_SRAM26(Tile_X10Y10_BM_SRAM26),
    .BM_SRAM27(Tile_X10Y10_BM_SRAM27),
    .BM_SRAM28(Tile_X10Y10_BM_SRAM28),
    .BM_SRAM29(Tile_X10Y10_BM_SRAM29),
    .BM_SRAM3(Tile_X10Y10_BM_SRAM3),
    .BM_SRAM30(Tile_X10Y10_BM_SRAM30),
    .BM_SRAM31(Tile_X10Y10_BM_SRAM31),
    .BM_SRAM4(Tile_X10Y10_BM_SRAM4),
    .BM_SRAM5(Tile_X10Y10_BM_SRAM5),
    .BM_SRAM6(Tile_X10Y10_BM_SRAM6),
    .BM_SRAM7(Tile_X10Y10_BM_SRAM7),
    .BM_SRAM8(Tile_X10Y10_BM_SRAM8),
    .BM_SRAM9(Tile_X10Y10_BM_SRAM9),
    .CLK_SRAM(Tile_X10Y10_CLK_SRAM),
    .CONFIGURED_top(Tile_X10Y10_CONFIGURED_top),
    .DIN_SRAM0(Tile_X10Y10_DIN_SRAM0),
    .DIN_SRAM1(Tile_X10Y10_DIN_SRAM1),
    .DIN_SRAM10(Tile_X10Y10_DIN_SRAM10),
    .DIN_SRAM11(Tile_X10Y10_DIN_SRAM11),
    .DIN_SRAM12(Tile_X10Y10_DIN_SRAM12),
    .DIN_SRAM13(Tile_X10Y10_DIN_SRAM13),
    .DIN_SRAM14(Tile_X10Y10_DIN_SRAM14),
    .DIN_SRAM15(Tile_X10Y10_DIN_SRAM15),
    .DIN_SRAM16(Tile_X10Y10_DIN_SRAM16),
    .DIN_SRAM17(Tile_X10Y10_DIN_SRAM17),
    .DIN_SRAM18(Tile_X10Y10_DIN_SRAM18),
    .DIN_SRAM19(Tile_X10Y10_DIN_SRAM19),
    .DIN_SRAM2(Tile_X10Y10_DIN_SRAM2),
    .DIN_SRAM20(Tile_X10Y10_DIN_SRAM20),
    .DIN_SRAM21(Tile_X10Y10_DIN_SRAM21),
    .DIN_SRAM22(Tile_X10Y10_DIN_SRAM22),
    .DIN_SRAM23(Tile_X10Y10_DIN_SRAM23),
    .DIN_SRAM24(Tile_X10Y10_DIN_SRAM24),
    .DIN_SRAM25(Tile_X10Y10_DIN_SRAM25),
    .DIN_SRAM26(Tile_X10Y10_DIN_SRAM26),
    .DIN_SRAM27(Tile_X10Y10_DIN_SRAM27),
    .DIN_SRAM28(Tile_X10Y10_DIN_SRAM28),
    .DIN_SRAM29(Tile_X10Y10_DIN_SRAM29),
    .DIN_SRAM3(Tile_X10Y10_DIN_SRAM3),
    .DIN_SRAM30(Tile_X10Y10_DIN_SRAM30),
    .DIN_SRAM31(Tile_X10Y10_DIN_SRAM31),
    .DIN_SRAM4(Tile_X10Y10_DIN_SRAM4),
    .DIN_SRAM5(Tile_X10Y10_DIN_SRAM5),
    .DIN_SRAM6(Tile_X10Y10_DIN_SRAM6),
    .DIN_SRAM7(Tile_X10Y10_DIN_SRAM7),
    .DIN_SRAM8(Tile_X10Y10_DIN_SRAM8),
    .DIN_SRAM9(Tile_X10Y10_DIN_SRAM9),
    .DOUT_SRAM0(Tile_X10Y10_DOUT_SRAM0),
    .DOUT_SRAM1(Tile_X10Y10_DOUT_SRAM1),
    .DOUT_SRAM10(Tile_X10Y10_DOUT_SRAM10),
    .DOUT_SRAM11(Tile_X10Y10_DOUT_SRAM11),
    .DOUT_SRAM12(Tile_X10Y10_DOUT_SRAM12),
    .DOUT_SRAM13(Tile_X10Y10_DOUT_SRAM13),
    .DOUT_SRAM14(Tile_X10Y10_DOUT_SRAM14),
    .DOUT_SRAM15(Tile_X10Y10_DOUT_SRAM15),
    .DOUT_SRAM16(Tile_X10Y10_DOUT_SRAM16),
    .DOUT_SRAM17(Tile_X10Y10_DOUT_SRAM17),
    .DOUT_SRAM18(Tile_X10Y10_DOUT_SRAM18),
    .DOUT_SRAM19(Tile_X10Y10_DOUT_SRAM19),
    .DOUT_SRAM2(Tile_X10Y10_DOUT_SRAM2),
    .DOUT_SRAM20(Tile_X10Y10_DOUT_SRAM20),
    .DOUT_SRAM21(Tile_X10Y10_DOUT_SRAM21),
    .DOUT_SRAM22(Tile_X10Y10_DOUT_SRAM22),
    .DOUT_SRAM23(Tile_X10Y10_DOUT_SRAM23),
    .DOUT_SRAM24(Tile_X10Y10_DOUT_SRAM24),
    .DOUT_SRAM25(Tile_X10Y10_DOUT_SRAM25),
    .DOUT_SRAM26(Tile_X10Y10_DOUT_SRAM26),
    .DOUT_SRAM27(Tile_X10Y10_DOUT_SRAM27),
    .DOUT_SRAM28(Tile_X10Y10_DOUT_SRAM28),
    .DOUT_SRAM29(Tile_X10Y10_DOUT_SRAM29),
    .DOUT_SRAM3(Tile_X10Y10_DOUT_SRAM3),
    .DOUT_SRAM30(Tile_X10Y10_DOUT_SRAM30),
    .DOUT_SRAM31(Tile_X10Y10_DOUT_SRAM31),
    .DOUT_SRAM4(Tile_X10Y10_DOUT_SRAM4),
    .DOUT_SRAM5(Tile_X10Y10_DOUT_SRAM5),
    .DOUT_SRAM6(Tile_X10Y10_DOUT_SRAM6),
    .DOUT_SRAM7(Tile_X10Y10_DOUT_SRAM7),
    .DOUT_SRAM8(Tile_X10Y10_DOUT_SRAM8),
    .DOUT_SRAM9(Tile_X10Y10_DOUT_SRAM9),
    .MEN_SRAM(Tile_X10Y10_MEN_SRAM),
    .REN_SRAM(Tile_X10Y10_REN_SRAM),
    .TIE_HIGH_SRAM(Tile_X10Y10_TIE_HIGH_SRAM),
    .TIE_LOW_SRAM(Tile_X10Y10_TIE_LOW_SRAM),
    .Tile_X0Y0_UserCLKo(Tile_X10Y9_UserCLKo),
    .Tile_X0Y1_UserCLK(Tile_X10Y11_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .WEN_SRAM(Tile_X10Y10_WEN_SRAM),
    .Tile_X0Y0_E1END({\Tile_X9Y9_E1BEG[3] ,
    \Tile_X9Y9_E1BEG[2] ,
    \Tile_X9Y9_E1BEG[1] ,
    \Tile_X9Y9_E1BEG[0] }),
    .Tile_X0Y0_E2END({\Tile_X9Y9_E2BEGb[7] ,
    \Tile_X9Y9_E2BEGb[6] ,
    \Tile_X9Y9_E2BEGb[5] ,
    \Tile_X9Y9_E2BEGb[4] ,
    \Tile_X9Y9_E2BEGb[3] ,
    \Tile_X9Y9_E2BEGb[2] ,
    \Tile_X9Y9_E2BEGb[1] ,
    \Tile_X9Y9_E2BEGb[0] }),
    .Tile_X0Y0_E2MID({\Tile_X9Y9_E2BEG[7] ,
    \Tile_X9Y9_E2BEG[6] ,
    \Tile_X9Y9_E2BEG[5] ,
    \Tile_X9Y9_E2BEG[4] ,
    \Tile_X9Y9_E2BEG[3] ,
    \Tile_X9Y9_E2BEG[2] ,
    \Tile_X9Y9_E2BEG[1] ,
    \Tile_X9Y9_E2BEG[0] }),
    .Tile_X0Y0_E6END({\Tile_X9Y9_E6BEG[11] ,
    \Tile_X9Y9_E6BEG[10] ,
    \Tile_X9Y9_E6BEG[9] ,
    \Tile_X9Y9_E6BEG[8] ,
    \Tile_X9Y9_E6BEG[7] ,
    \Tile_X9Y9_E6BEG[6] ,
    \Tile_X9Y9_E6BEG[5] ,
    \Tile_X9Y9_E6BEG[4] ,
    \Tile_X9Y9_E6BEG[3] ,
    \Tile_X9Y9_E6BEG[2] ,
    \Tile_X9Y9_E6BEG[1] ,
    \Tile_X9Y9_E6BEG[0] }),
    .Tile_X0Y0_EE4END({\Tile_X9Y9_EE4BEG[15] ,
    \Tile_X9Y9_EE4BEG[14] ,
    \Tile_X9Y9_EE4BEG[13] ,
    \Tile_X9Y9_EE4BEG[12] ,
    \Tile_X9Y9_EE4BEG[11] ,
    \Tile_X9Y9_EE4BEG[10] ,
    \Tile_X9Y9_EE4BEG[9] ,
    \Tile_X9Y9_EE4BEG[8] ,
    \Tile_X9Y9_EE4BEG[7] ,
    \Tile_X9Y9_EE4BEG[6] ,
    \Tile_X9Y9_EE4BEG[5] ,
    \Tile_X9Y9_EE4BEG[4] ,
    \Tile_X9Y9_EE4BEG[3] ,
    \Tile_X9Y9_EE4BEG[2] ,
    \Tile_X9Y9_EE4BEG[1] ,
    \Tile_X9Y9_EE4BEG[0] }),
    .Tile_X0Y0_FrameData({\Tile_X9Y9_FrameData_O[31] ,
    \Tile_X9Y9_FrameData_O[30] ,
    \Tile_X9Y9_FrameData_O[29] ,
    \Tile_X9Y9_FrameData_O[28] ,
    \Tile_X9Y9_FrameData_O[27] ,
    \Tile_X9Y9_FrameData_O[26] ,
    \Tile_X9Y9_FrameData_O[25] ,
    \Tile_X9Y9_FrameData_O[24] ,
    \Tile_X9Y9_FrameData_O[23] ,
    \Tile_X9Y9_FrameData_O[22] ,
    \Tile_X9Y9_FrameData_O[21] ,
    \Tile_X9Y9_FrameData_O[20] ,
    \Tile_X9Y9_FrameData_O[19] ,
    \Tile_X9Y9_FrameData_O[18] ,
    \Tile_X9Y9_FrameData_O[17] ,
    \Tile_X9Y9_FrameData_O[16] ,
    \Tile_X9Y9_FrameData_O[15] ,
    \Tile_X9Y9_FrameData_O[14] ,
    \Tile_X9Y9_FrameData_O[13] ,
    \Tile_X9Y9_FrameData_O[12] ,
    \Tile_X9Y9_FrameData_O[11] ,
    \Tile_X9Y9_FrameData_O[10] ,
    \Tile_X9Y9_FrameData_O[9] ,
    \Tile_X9Y9_FrameData_O[8] ,
    \Tile_X9Y9_FrameData_O[7] ,
    \Tile_X9Y9_FrameData_O[6] ,
    \Tile_X9Y9_FrameData_O[5] ,
    \Tile_X9Y9_FrameData_O[4] ,
    \Tile_X9Y9_FrameData_O[3] ,
    \Tile_X9Y9_FrameData_O[2] ,
    \Tile_X9Y9_FrameData_O[1] ,
    \Tile_X9Y9_FrameData_O[0] }),
    .Tile_X0Y0_FrameData_O({\Tile_X10Y9_FrameData_O[31] ,
    \Tile_X10Y9_FrameData_O[30] ,
    \Tile_X10Y9_FrameData_O[29] ,
    \Tile_X10Y9_FrameData_O[28] ,
    \Tile_X10Y9_FrameData_O[27] ,
    \Tile_X10Y9_FrameData_O[26] ,
    \Tile_X10Y9_FrameData_O[25] ,
    \Tile_X10Y9_FrameData_O[24] ,
    \Tile_X10Y9_FrameData_O[23] ,
    \Tile_X10Y9_FrameData_O[22] ,
    \Tile_X10Y9_FrameData_O[21] ,
    \Tile_X10Y9_FrameData_O[20] ,
    \Tile_X10Y9_FrameData_O[19] ,
    \Tile_X10Y9_FrameData_O[18] ,
    \Tile_X10Y9_FrameData_O[17] ,
    \Tile_X10Y9_FrameData_O[16] ,
    \Tile_X10Y9_FrameData_O[15] ,
    \Tile_X10Y9_FrameData_O[14] ,
    \Tile_X10Y9_FrameData_O[13] ,
    \Tile_X10Y9_FrameData_O[12] ,
    \Tile_X10Y9_FrameData_O[11] ,
    \Tile_X10Y9_FrameData_O[10] ,
    \Tile_X10Y9_FrameData_O[9] ,
    \Tile_X10Y9_FrameData_O[8] ,
    \Tile_X10Y9_FrameData_O[7] ,
    \Tile_X10Y9_FrameData_O[6] ,
    \Tile_X10Y9_FrameData_O[5] ,
    \Tile_X10Y9_FrameData_O[4] ,
    \Tile_X10Y9_FrameData_O[3] ,
    \Tile_X10Y9_FrameData_O[2] ,
    \Tile_X10Y9_FrameData_O[1] ,
    \Tile_X10Y9_FrameData_O[0] }),
    .Tile_X0Y0_FrameStrobe_O({\Tile_X10Y9_FrameStrobe_O[19] ,
    \Tile_X10Y9_FrameStrobe_O[18] ,
    \Tile_X10Y9_FrameStrobe_O[17] ,
    \Tile_X10Y9_FrameStrobe_O[16] ,
    \Tile_X10Y9_FrameStrobe_O[15] ,
    \Tile_X10Y9_FrameStrobe_O[14] ,
    \Tile_X10Y9_FrameStrobe_O[13] ,
    \Tile_X10Y9_FrameStrobe_O[12] ,
    \Tile_X10Y9_FrameStrobe_O[11] ,
    \Tile_X10Y9_FrameStrobe_O[10] ,
    \Tile_X10Y9_FrameStrobe_O[9] ,
    \Tile_X10Y9_FrameStrobe_O[8] ,
    \Tile_X10Y9_FrameStrobe_O[7] ,
    \Tile_X10Y9_FrameStrobe_O[6] ,
    \Tile_X10Y9_FrameStrobe_O[5] ,
    \Tile_X10Y9_FrameStrobe_O[4] ,
    \Tile_X10Y9_FrameStrobe_O[3] ,
    \Tile_X10Y9_FrameStrobe_O[2] ,
    \Tile_X10Y9_FrameStrobe_O[1] ,
    \Tile_X10Y9_FrameStrobe_O[0] }),
    .Tile_X0Y0_N1BEG({\Tile_X10Y9_N1BEG[3] ,
    \Tile_X10Y9_N1BEG[2] ,
    \Tile_X10Y9_N1BEG[1] ,
    \Tile_X10Y9_N1BEG[0] }),
    .Tile_X0Y0_N2BEG({\Tile_X10Y9_N2BEG[7] ,
    \Tile_X10Y9_N2BEG[6] ,
    \Tile_X10Y9_N2BEG[5] ,
    \Tile_X10Y9_N2BEG[4] ,
    \Tile_X10Y9_N2BEG[3] ,
    \Tile_X10Y9_N2BEG[2] ,
    \Tile_X10Y9_N2BEG[1] ,
    \Tile_X10Y9_N2BEG[0] }),
    .Tile_X0Y0_N2BEGb({\Tile_X10Y9_N2BEGb[7] ,
    \Tile_X10Y9_N2BEGb[6] ,
    \Tile_X10Y9_N2BEGb[5] ,
    \Tile_X10Y9_N2BEGb[4] ,
    \Tile_X10Y9_N2BEGb[3] ,
    \Tile_X10Y9_N2BEGb[2] ,
    \Tile_X10Y9_N2BEGb[1] ,
    \Tile_X10Y9_N2BEGb[0] }),
    .Tile_X0Y0_N4BEG({\Tile_X10Y9_N4BEG[15] ,
    \Tile_X10Y9_N4BEG[14] ,
    \Tile_X10Y9_N4BEG[13] ,
    \Tile_X10Y9_N4BEG[12] ,
    \Tile_X10Y9_N4BEG[11] ,
    \Tile_X10Y9_N4BEG[10] ,
    \Tile_X10Y9_N4BEG[9] ,
    \Tile_X10Y9_N4BEG[8] ,
    \Tile_X10Y9_N4BEG[7] ,
    \Tile_X10Y9_N4BEG[6] ,
    \Tile_X10Y9_N4BEG[5] ,
    \Tile_X10Y9_N4BEG[4] ,
    \Tile_X10Y9_N4BEG[3] ,
    \Tile_X10Y9_N4BEG[2] ,
    \Tile_X10Y9_N4BEG[1] ,
    \Tile_X10Y9_N4BEG[0] }),
    .Tile_X0Y0_S1END({\Tile_X10Y8_S1BEG[3] ,
    \Tile_X10Y8_S1BEG[2] ,
    \Tile_X10Y8_S1BEG[1] ,
    \Tile_X10Y8_S1BEG[0] }),
    .Tile_X0Y0_S2END({\Tile_X10Y8_S2BEGb[7] ,
    \Tile_X10Y8_S2BEGb[6] ,
    \Tile_X10Y8_S2BEGb[5] ,
    \Tile_X10Y8_S2BEGb[4] ,
    \Tile_X10Y8_S2BEGb[3] ,
    \Tile_X10Y8_S2BEGb[2] ,
    \Tile_X10Y8_S2BEGb[1] ,
    \Tile_X10Y8_S2BEGb[0] }),
    .Tile_X0Y0_S2MID({\Tile_X10Y8_S2BEG[7] ,
    \Tile_X10Y8_S2BEG[6] ,
    \Tile_X10Y8_S2BEG[5] ,
    \Tile_X10Y8_S2BEG[4] ,
    \Tile_X10Y8_S2BEG[3] ,
    \Tile_X10Y8_S2BEG[2] ,
    \Tile_X10Y8_S2BEG[1] ,
    \Tile_X10Y8_S2BEG[0] }),
    .Tile_X0Y0_S4END({\Tile_X10Y8_S4BEG[15] ,
    \Tile_X10Y8_S4BEG[14] ,
    \Tile_X10Y8_S4BEG[13] ,
    \Tile_X10Y8_S4BEG[12] ,
    \Tile_X10Y8_S4BEG[11] ,
    \Tile_X10Y8_S4BEG[10] ,
    \Tile_X10Y8_S4BEG[9] ,
    \Tile_X10Y8_S4BEG[8] ,
    \Tile_X10Y8_S4BEG[7] ,
    \Tile_X10Y8_S4BEG[6] ,
    \Tile_X10Y8_S4BEG[5] ,
    \Tile_X10Y8_S4BEG[4] ,
    \Tile_X10Y8_S4BEG[3] ,
    \Tile_X10Y8_S4BEG[2] ,
    \Tile_X10Y8_S4BEG[1] ,
    \Tile_X10Y8_S4BEG[0] }),
    .Tile_X0Y0_W1BEG({\Tile_X10Y9_W1BEG[3] ,
    \Tile_X10Y9_W1BEG[2] ,
    \Tile_X10Y9_W1BEG[1] ,
    \Tile_X10Y9_W1BEG[0] }),
    .Tile_X0Y0_W2BEG({\Tile_X10Y9_W2BEG[7] ,
    \Tile_X10Y9_W2BEG[6] ,
    \Tile_X10Y9_W2BEG[5] ,
    \Tile_X10Y9_W2BEG[4] ,
    \Tile_X10Y9_W2BEG[3] ,
    \Tile_X10Y9_W2BEG[2] ,
    \Tile_X10Y9_W2BEG[1] ,
    \Tile_X10Y9_W2BEG[0] }),
    .Tile_X0Y0_W2BEGb({\Tile_X10Y9_W2BEGb[7] ,
    \Tile_X10Y9_W2BEGb[6] ,
    \Tile_X10Y9_W2BEGb[5] ,
    \Tile_X10Y9_W2BEGb[4] ,
    \Tile_X10Y9_W2BEGb[3] ,
    \Tile_X10Y9_W2BEGb[2] ,
    \Tile_X10Y9_W2BEGb[1] ,
    \Tile_X10Y9_W2BEGb[0] }),
    .Tile_X0Y0_W6BEG({\Tile_X10Y9_W6BEG[11] ,
    \Tile_X10Y9_W6BEG[10] ,
    \Tile_X10Y9_W6BEG[9] ,
    \Tile_X10Y9_W6BEG[8] ,
    \Tile_X10Y9_W6BEG[7] ,
    \Tile_X10Y9_W6BEG[6] ,
    \Tile_X10Y9_W6BEG[5] ,
    \Tile_X10Y9_W6BEG[4] ,
    \Tile_X10Y9_W6BEG[3] ,
    \Tile_X10Y9_W6BEG[2] ,
    \Tile_X10Y9_W6BEG[1] ,
    \Tile_X10Y9_W6BEG[0] }),
    .Tile_X0Y0_WW4BEG({\Tile_X10Y9_WW4BEG[15] ,
    \Tile_X10Y9_WW4BEG[14] ,
    \Tile_X10Y9_WW4BEG[13] ,
    \Tile_X10Y9_WW4BEG[12] ,
    \Tile_X10Y9_WW4BEG[11] ,
    \Tile_X10Y9_WW4BEG[10] ,
    \Tile_X10Y9_WW4BEG[9] ,
    \Tile_X10Y9_WW4BEG[8] ,
    \Tile_X10Y9_WW4BEG[7] ,
    \Tile_X10Y9_WW4BEG[6] ,
    \Tile_X10Y9_WW4BEG[5] ,
    \Tile_X10Y9_WW4BEG[4] ,
    \Tile_X10Y9_WW4BEG[3] ,
    \Tile_X10Y9_WW4BEG[2] ,
    \Tile_X10Y9_WW4BEG[1] ,
    \Tile_X10Y9_WW4BEG[0] }),
    .Tile_X0Y1_E1END({\Tile_X9Y10_E1BEG[3] ,
    \Tile_X9Y10_E1BEG[2] ,
    \Tile_X9Y10_E1BEG[1] ,
    \Tile_X9Y10_E1BEG[0] }),
    .Tile_X0Y1_E2END({\Tile_X9Y10_E2BEGb[7] ,
    \Tile_X9Y10_E2BEGb[6] ,
    \Tile_X9Y10_E2BEGb[5] ,
    \Tile_X9Y10_E2BEGb[4] ,
    \Tile_X9Y10_E2BEGb[3] ,
    \Tile_X9Y10_E2BEGb[2] ,
    \Tile_X9Y10_E2BEGb[1] ,
    \Tile_X9Y10_E2BEGb[0] }),
    .Tile_X0Y1_E2MID({\Tile_X9Y10_E2BEG[7] ,
    \Tile_X9Y10_E2BEG[6] ,
    \Tile_X9Y10_E2BEG[5] ,
    \Tile_X9Y10_E2BEG[4] ,
    \Tile_X9Y10_E2BEG[3] ,
    \Tile_X9Y10_E2BEG[2] ,
    \Tile_X9Y10_E2BEG[1] ,
    \Tile_X9Y10_E2BEG[0] }),
    .Tile_X0Y1_E6END({\Tile_X9Y10_E6BEG[11] ,
    \Tile_X9Y10_E6BEG[10] ,
    \Tile_X9Y10_E6BEG[9] ,
    \Tile_X9Y10_E6BEG[8] ,
    \Tile_X9Y10_E6BEG[7] ,
    \Tile_X9Y10_E6BEG[6] ,
    \Tile_X9Y10_E6BEG[5] ,
    \Tile_X9Y10_E6BEG[4] ,
    \Tile_X9Y10_E6BEG[3] ,
    \Tile_X9Y10_E6BEG[2] ,
    \Tile_X9Y10_E6BEG[1] ,
    \Tile_X9Y10_E6BEG[0] }),
    .Tile_X0Y1_EE4END({\Tile_X9Y10_EE4BEG[15] ,
    \Tile_X9Y10_EE4BEG[14] ,
    \Tile_X9Y10_EE4BEG[13] ,
    \Tile_X9Y10_EE4BEG[12] ,
    \Tile_X9Y10_EE4BEG[11] ,
    \Tile_X9Y10_EE4BEG[10] ,
    \Tile_X9Y10_EE4BEG[9] ,
    \Tile_X9Y10_EE4BEG[8] ,
    \Tile_X9Y10_EE4BEG[7] ,
    \Tile_X9Y10_EE4BEG[6] ,
    \Tile_X9Y10_EE4BEG[5] ,
    \Tile_X9Y10_EE4BEG[4] ,
    \Tile_X9Y10_EE4BEG[3] ,
    \Tile_X9Y10_EE4BEG[2] ,
    \Tile_X9Y10_EE4BEG[1] ,
    \Tile_X9Y10_EE4BEG[0] }),
    .Tile_X0Y1_FrameData({\Tile_X9Y10_FrameData_O[31] ,
    \Tile_X9Y10_FrameData_O[30] ,
    \Tile_X9Y10_FrameData_O[29] ,
    \Tile_X9Y10_FrameData_O[28] ,
    \Tile_X9Y10_FrameData_O[27] ,
    \Tile_X9Y10_FrameData_O[26] ,
    \Tile_X9Y10_FrameData_O[25] ,
    \Tile_X9Y10_FrameData_O[24] ,
    \Tile_X9Y10_FrameData_O[23] ,
    \Tile_X9Y10_FrameData_O[22] ,
    \Tile_X9Y10_FrameData_O[21] ,
    \Tile_X9Y10_FrameData_O[20] ,
    \Tile_X9Y10_FrameData_O[19] ,
    \Tile_X9Y10_FrameData_O[18] ,
    \Tile_X9Y10_FrameData_O[17] ,
    \Tile_X9Y10_FrameData_O[16] ,
    \Tile_X9Y10_FrameData_O[15] ,
    \Tile_X9Y10_FrameData_O[14] ,
    \Tile_X9Y10_FrameData_O[13] ,
    \Tile_X9Y10_FrameData_O[12] ,
    \Tile_X9Y10_FrameData_O[11] ,
    \Tile_X9Y10_FrameData_O[10] ,
    \Tile_X9Y10_FrameData_O[9] ,
    \Tile_X9Y10_FrameData_O[8] ,
    \Tile_X9Y10_FrameData_O[7] ,
    \Tile_X9Y10_FrameData_O[6] ,
    \Tile_X9Y10_FrameData_O[5] ,
    \Tile_X9Y10_FrameData_O[4] ,
    \Tile_X9Y10_FrameData_O[3] ,
    \Tile_X9Y10_FrameData_O[2] ,
    \Tile_X9Y10_FrameData_O[1] ,
    \Tile_X9Y10_FrameData_O[0] }),
    .Tile_X0Y1_FrameData_O({\Tile_X10Y10_FrameData_O[31] ,
    \Tile_X10Y10_FrameData_O[30] ,
    \Tile_X10Y10_FrameData_O[29] ,
    \Tile_X10Y10_FrameData_O[28] ,
    \Tile_X10Y10_FrameData_O[27] ,
    \Tile_X10Y10_FrameData_O[26] ,
    \Tile_X10Y10_FrameData_O[25] ,
    \Tile_X10Y10_FrameData_O[24] ,
    \Tile_X10Y10_FrameData_O[23] ,
    \Tile_X10Y10_FrameData_O[22] ,
    \Tile_X10Y10_FrameData_O[21] ,
    \Tile_X10Y10_FrameData_O[20] ,
    \Tile_X10Y10_FrameData_O[19] ,
    \Tile_X10Y10_FrameData_O[18] ,
    \Tile_X10Y10_FrameData_O[17] ,
    \Tile_X10Y10_FrameData_O[16] ,
    \Tile_X10Y10_FrameData_O[15] ,
    \Tile_X10Y10_FrameData_O[14] ,
    \Tile_X10Y10_FrameData_O[13] ,
    \Tile_X10Y10_FrameData_O[12] ,
    \Tile_X10Y10_FrameData_O[11] ,
    \Tile_X10Y10_FrameData_O[10] ,
    \Tile_X10Y10_FrameData_O[9] ,
    \Tile_X10Y10_FrameData_O[8] ,
    \Tile_X10Y10_FrameData_O[7] ,
    \Tile_X10Y10_FrameData_O[6] ,
    \Tile_X10Y10_FrameData_O[5] ,
    \Tile_X10Y10_FrameData_O[4] ,
    \Tile_X10Y10_FrameData_O[3] ,
    \Tile_X10Y10_FrameData_O[2] ,
    \Tile_X10Y10_FrameData_O[1] ,
    \Tile_X10Y10_FrameData_O[0] }),
    .Tile_X0Y1_FrameStrobe({\Tile_X10Y11_FrameStrobe_O[19] ,
    \Tile_X10Y11_FrameStrobe_O[18] ,
    \Tile_X10Y11_FrameStrobe_O[17] ,
    \Tile_X10Y11_FrameStrobe_O[16] ,
    \Tile_X10Y11_FrameStrobe_O[15] ,
    \Tile_X10Y11_FrameStrobe_O[14] ,
    \Tile_X10Y11_FrameStrobe_O[13] ,
    \Tile_X10Y11_FrameStrobe_O[12] ,
    \Tile_X10Y11_FrameStrobe_O[11] ,
    \Tile_X10Y11_FrameStrobe_O[10] ,
    \Tile_X10Y11_FrameStrobe_O[9] ,
    \Tile_X10Y11_FrameStrobe_O[8] ,
    \Tile_X10Y11_FrameStrobe_O[7] ,
    \Tile_X10Y11_FrameStrobe_O[6] ,
    \Tile_X10Y11_FrameStrobe_O[5] ,
    \Tile_X10Y11_FrameStrobe_O[4] ,
    \Tile_X10Y11_FrameStrobe_O[3] ,
    \Tile_X10Y11_FrameStrobe_O[2] ,
    \Tile_X10Y11_FrameStrobe_O[1] ,
    \Tile_X10Y11_FrameStrobe_O[0] }),
    .Tile_X0Y1_N1END({\Tile_X10Y11_N1BEG[3] ,
    \Tile_X10Y11_N1BEG[2] ,
    \Tile_X10Y11_N1BEG[1] ,
    \Tile_X10Y11_N1BEG[0] }),
    .Tile_X0Y1_N2END({\Tile_X10Y11_N2BEGb[7] ,
    \Tile_X10Y11_N2BEGb[6] ,
    \Tile_X10Y11_N2BEGb[5] ,
    \Tile_X10Y11_N2BEGb[4] ,
    \Tile_X10Y11_N2BEGb[3] ,
    \Tile_X10Y11_N2BEGb[2] ,
    \Tile_X10Y11_N2BEGb[1] ,
    \Tile_X10Y11_N2BEGb[0] }),
    .Tile_X0Y1_N2MID({\Tile_X10Y11_N2BEG[7] ,
    \Tile_X10Y11_N2BEG[6] ,
    \Tile_X10Y11_N2BEG[5] ,
    \Tile_X10Y11_N2BEG[4] ,
    \Tile_X10Y11_N2BEG[3] ,
    \Tile_X10Y11_N2BEG[2] ,
    \Tile_X10Y11_N2BEG[1] ,
    \Tile_X10Y11_N2BEG[0] }),
    .Tile_X0Y1_N4END({\Tile_X10Y11_N4BEG[15] ,
    \Tile_X10Y11_N4BEG[14] ,
    \Tile_X10Y11_N4BEG[13] ,
    \Tile_X10Y11_N4BEG[12] ,
    \Tile_X10Y11_N4BEG[11] ,
    \Tile_X10Y11_N4BEG[10] ,
    \Tile_X10Y11_N4BEG[9] ,
    \Tile_X10Y11_N4BEG[8] ,
    \Tile_X10Y11_N4BEG[7] ,
    \Tile_X10Y11_N4BEG[6] ,
    \Tile_X10Y11_N4BEG[5] ,
    \Tile_X10Y11_N4BEG[4] ,
    \Tile_X10Y11_N4BEG[3] ,
    \Tile_X10Y11_N4BEG[2] ,
    \Tile_X10Y11_N4BEG[1] ,
    \Tile_X10Y11_N4BEG[0] }),
    .Tile_X0Y1_S1BEG({\Tile_X10Y10_S1BEG[3] ,
    \Tile_X10Y10_S1BEG[2] ,
    \Tile_X10Y10_S1BEG[1] ,
    \Tile_X10Y10_S1BEG[0] }),
    .Tile_X0Y1_S2BEG({\Tile_X10Y10_S2BEG[7] ,
    \Tile_X10Y10_S2BEG[6] ,
    \Tile_X10Y10_S2BEG[5] ,
    \Tile_X10Y10_S2BEG[4] ,
    \Tile_X10Y10_S2BEG[3] ,
    \Tile_X10Y10_S2BEG[2] ,
    \Tile_X10Y10_S2BEG[1] ,
    \Tile_X10Y10_S2BEG[0] }),
    .Tile_X0Y1_S2BEGb({\Tile_X10Y10_S2BEGb[7] ,
    \Tile_X10Y10_S2BEGb[6] ,
    \Tile_X10Y10_S2BEGb[5] ,
    \Tile_X10Y10_S2BEGb[4] ,
    \Tile_X10Y10_S2BEGb[3] ,
    \Tile_X10Y10_S2BEGb[2] ,
    \Tile_X10Y10_S2BEGb[1] ,
    \Tile_X10Y10_S2BEGb[0] }),
    .Tile_X0Y1_S4BEG({\Tile_X10Y10_S4BEG[15] ,
    \Tile_X10Y10_S4BEG[14] ,
    \Tile_X10Y10_S4BEG[13] ,
    \Tile_X10Y10_S4BEG[12] ,
    \Tile_X10Y10_S4BEG[11] ,
    \Tile_X10Y10_S4BEG[10] ,
    \Tile_X10Y10_S4BEG[9] ,
    \Tile_X10Y10_S4BEG[8] ,
    \Tile_X10Y10_S4BEG[7] ,
    \Tile_X10Y10_S4BEG[6] ,
    \Tile_X10Y10_S4BEG[5] ,
    \Tile_X10Y10_S4BEG[4] ,
    \Tile_X10Y10_S4BEG[3] ,
    \Tile_X10Y10_S4BEG[2] ,
    \Tile_X10Y10_S4BEG[1] ,
    \Tile_X10Y10_S4BEG[0] }),
    .Tile_X0Y1_W1BEG({\Tile_X10Y10_W1BEG[3] ,
    \Tile_X10Y10_W1BEG[2] ,
    \Tile_X10Y10_W1BEG[1] ,
    \Tile_X10Y10_W1BEG[0] }),
    .Tile_X0Y1_W2BEG({\Tile_X10Y10_W2BEG[7] ,
    \Tile_X10Y10_W2BEG[6] ,
    \Tile_X10Y10_W2BEG[5] ,
    \Tile_X10Y10_W2BEG[4] ,
    \Tile_X10Y10_W2BEG[3] ,
    \Tile_X10Y10_W2BEG[2] ,
    \Tile_X10Y10_W2BEG[1] ,
    \Tile_X10Y10_W2BEG[0] }),
    .Tile_X0Y1_W2BEGb({\Tile_X10Y10_W2BEGb[7] ,
    \Tile_X10Y10_W2BEGb[6] ,
    \Tile_X10Y10_W2BEGb[5] ,
    \Tile_X10Y10_W2BEGb[4] ,
    \Tile_X10Y10_W2BEGb[3] ,
    \Tile_X10Y10_W2BEGb[2] ,
    \Tile_X10Y10_W2BEGb[1] ,
    \Tile_X10Y10_W2BEGb[0] }),
    .Tile_X0Y1_W6BEG({\Tile_X10Y10_W6BEG[11] ,
    \Tile_X10Y10_W6BEG[10] ,
    \Tile_X10Y10_W6BEG[9] ,
    \Tile_X10Y10_W6BEG[8] ,
    \Tile_X10Y10_W6BEG[7] ,
    \Tile_X10Y10_W6BEG[6] ,
    \Tile_X10Y10_W6BEG[5] ,
    \Tile_X10Y10_W6BEG[4] ,
    \Tile_X10Y10_W6BEG[3] ,
    \Tile_X10Y10_W6BEG[2] ,
    \Tile_X10Y10_W6BEG[1] ,
    \Tile_X10Y10_W6BEG[0] }),
    .Tile_X0Y1_WW4BEG({\Tile_X10Y10_WW4BEG[15] ,
    \Tile_X10Y10_WW4BEG[14] ,
    \Tile_X10Y10_WW4BEG[13] ,
    \Tile_X10Y10_WW4BEG[12] ,
    \Tile_X10Y10_WW4BEG[11] ,
    \Tile_X10Y10_WW4BEG[10] ,
    \Tile_X10Y10_WW4BEG[9] ,
    \Tile_X10Y10_WW4BEG[8] ,
    \Tile_X10Y10_WW4BEG[7] ,
    \Tile_X10Y10_WW4BEG[6] ,
    \Tile_X10Y10_WW4BEG[5] ,
    \Tile_X10Y10_WW4BEG[4] ,
    \Tile_X10Y10_WW4BEG[3] ,
    \Tile_X10Y10_WW4BEG[2] ,
    \Tile_X10Y10_WW4BEG[1] ,
    \Tile_X10Y10_WW4BEG[0] }));
 N_IO Tile_X1Y0_N_IO (.A_I_top(Tile_X1Y0_A_I_top),
    .A_O_top(Tile_X1Y0_A_O_top),
    .A_T_top(Tile_X1Y0_A_T_top),
    .A_config_C_bit0(Tile_X1Y0_A_config_C_bit0),
    .A_config_C_bit1(Tile_X1Y0_A_config_C_bit1),
    .A_config_C_bit2(Tile_X1Y0_A_config_C_bit2),
    .A_config_C_bit3(Tile_X1Y0_A_config_C_bit3),
    .B_I_top(Tile_X1Y0_B_I_top),
    .B_O_top(Tile_X1Y0_B_O_top),
    .B_T_top(Tile_X1Y0_B_T_top),
    .B_config_C_bit0(Tile_X1Y0_B_config_C_bit0),
    .B_config_C_bit1(Tile_X1Y0_B_config_C_bit1),
    .B_config_C_bit2(Tile_X1Y0_B_config_C_bit2),
    .B_config_C_bit3(Tile_X1Y0_B_config_C_bit3),
    .Ci(Tile_X1Y1_Co),
    .UserCLK(Tile_X1Y1_UserCLKo),
    .UserCLKo(Tile_X1Y0_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .FrameData({FrameData[31],
    FrameData[30],
    FrameData[29],
    FrameData[28],
    FrameData[27],
    FrameData[26],
    FrameData[25],
    FrameData[24],
    FrameData[23],
    FrameData[22],
    FrameData[21],
    FrameData[20],
    FrameData[19],
    FrameData[18],
    FrameData[17],
    FrameData[16],
    FrameData[15],
    FrameData[14],
    FrameData[13],
    FrameData[12],
    FrameData[11],
    FrameData[10],
    FrameData[9],
    FrameData[8],
    FrameData[7],
    FrameData[6],
    FrameData[5],
    FrameData[4],
    FrameData[3],
    FrameData[2],
    FrameData[1],
    FrameData[0]}),
    .FrameData_O({\Tile_X1Y0_FrameData_O[31] ,
    \Tile_X1Y0_FrameData_O[30] ,
    \Tile_X1Y0_FrameData_O[29] ,
    \Tile_X1Y0_FrameData_O[28] ,
    \Tile_X1Y0_FrameData_O[27] ,
    \Tile_X1Y0_FrameData_O[26] ,
    \Tile_X1Y0_FrameData_O[25] ,
    \Tile_X1Y0_FrameData_O[24] ,
    \Tile_X1Y0_FrameData_O[23] ,
    \Tile_X1Y0_FrameData_O[22] ,
    \Tile_X1Y0_FrameData_O[21] ,
    \Tile_X1Y0_FrameData_O[20] ,
    \Tile_X1Y0_FrameData_O[19] ,
    \Tile_X1Y0_FrameData_O[18] ,
    \Tile_X1Y0_FrameData_O[17] ,
    \Tile_X1Y0_FrameData_O[16] ,
    \Tile_X1Y0_FrameData_O[15] ,
    \Tile_X1Y0_FrameData_O[14] ,
    \Tile_X1Y0_FrameData_O[13] ,
    \Tile_X1Y0_FrameData_O[12] ,
    \Tile_X1Y0_FrameData_O[11] ,
    \Tile_X1Y0_FrameData_O[10] ,
    \Tile_X1Y0_FrameData_O[9] ,
    \Tile_X1Y0_FrameData_O[8] ,
    \Tile_X1Y0_FrameData_O[7] ,
    \Tile_X1Y0_FrameData_O[6] ,
    \Tile_X1Y0_FrameData_O[5] ,
    \Tile_X1Y0_FrameData_O[4] ,
    \Tile_X1Y0_FrameData_O[3] ,
    \Tile_X1Y0_FrameData_O[2] ,
    \Tile_X1Y0_FrameData_O[1] ,
    \Tile_X1Y0_FrameData_O[0] }),
    .FrameStrobe({\Tile_X1Y1_FrameStrobe_O[19] ,
    \Tile_X1Y1_FrameStrobe_O[18] ,
    \Tile_X1Y1_FrameStrobe_O[17] ,
    \Tile_X1Y1_FrameStrobe_O[16] ,
    \Tile_X1Y1_FrameStrobe_O[15] ,
    \Tile_X1Y1_FrameStrobe_O[14] ,
    \Tile_X1Y1_FrameStrobe_O[13] ,
    \Tile_X1Y1_FrameStrobe_O[12] ,
    \Tile_X1Y1_FrameStrobe_O[11] ,
    \Tile_X1Y1_FrameStrobe_O[10] ,
    \Tile_X1Y1_FrameStrobe_O[9] ,
    \Tile_X1Y1_FrameStrobe_O[8] ,
    \Tile_X1Y1_FrameStrobe_O[7] ,
    \Tile_X1Y1_FrameStrobe_O[6] ,
    \Tile_X1Y1_FrameStrobe_O[5] ,
    \Tile_X1Y1_FrameStrobe_O[4] ,
    \Tile_X1Y1_FrameStrobe_O[3] ,
    \Tile_X1Y1_FrameStrobe_O[2] ,
    \Tile_X1Y1_FrameStrobe_O[1] ,
    \Tile_X1Y1_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X1Y0_FrameStrobe_O[19] ,
    \Tile_X1Y0_FrameStrobe_O[18] ,
    \Tile_X1Y0_FrameStrobe_O[17] ,
    \Tile_X1Y0_FrameStrobe_O[16] ,
    \Tile_X1Y0_FrameStrobe_O[15] ,
    \Tile_X1Y0_FrameStrobe_O[14] ,
    \Tile_X1Y0_FrameStrobe_O[13] ,
    \Tile_X1Y0_FrameStrobe_O[12] ,
    \Tile_X1Y0_FrameStrobe_O[11] ,
    \Tile_X1Y0_FrameStrobe_O[10] ,
    \Tile_X1Y0_FrameStrobe_O[9] ,
    \Tile_X1Y0_FrameStrobe_O[8] ,
    \Tile_X1Y0_FrameStrobe_O[7] ,
    \Tile_X1Y0_FrameStrobe_O[6] ,
    \Tile_X1Y0_FrameStrobe_O[5] ,
    \Tile_X1Y0_FrameStrobe_O[4] ,
    \Tile_X1Y0_FrameStrobe_O[3] ,
    \Tile_X1Y0_FrameStrobe_O[2] ,
    \Tile_X1Y0_FrameStrobe_O[1] ,
    \Tile_X1Y0_FrameStrobe_O[0] }),
    .N1END({\Tile_X1Y1_N1BEG[3] ,
    \Tile_X1Y1_N1BEG[2] ,
    \Tile_X1Y1_N1BEG[1] ,
    \Tile_X1Y1_N1BEG[0] }),
    .N2END({\Tile_X1Y1_N2BEGb[7] ,
    \Tile_X1Y1_N2BEGb[6] ,
    \Tile_X1Y1_N2BEGb[5] ,
    \Tile_X1Y1_N2BEGb[4] ,
    \Tile_X1Y1_N2BEGb[3] ,
    \Tile_X1Y1_N2BEGb[2] ,
    \Tile_X1Y1_N2BEGb[1] ,
    \Tile_X1Y1_N2BEGb[0] }),
    .N2MID({\Tile_X1Y1_N2BEG[7] ,
    \Tile_X1Y1_N2BEG[6] ,
    \Tile_X1Y1_N2BEG[5] ,
    \Tile_X1Y1_N2BEG[4] ,
    \Tile_X1Y1_N2BEG[3] ,
    \Tile_X1Y1_N2BEG[2] ,
    \Tile_X1Y1_N2BEG[1] ,
    \Tile_X1Y1_N2BEG[0] }),
    .N4END({\Tile_X1Y1_N4BEG[15] ,
    \Tile_X1Y1_N4BEG[14] ,
    \Tile_X1Y1_N4BEG[13] ,
    \Tile_X1Y1_N4BEG[12] ,
    \Tile_X1Y1_N4BEG[11] ,
    \Tile_X1Y1_N4BEG[10] ,
    \Tile_X1Y1_N4BEG[9] ,
    \Tile_X1Y1_N4BEG[8] ,
    \Tile_X1Y1_N4BEG[7] ,
    \Tile_X1Y1_N4BEG[6] ,
    \Tile_X1Y1_N4BEG[5] ,
    \Tile_X1Y1_N4BEG[4] ,
    \Tile_X1Y1_N4BEG[3] ,
    \Tile_X1Y1_N4BEG[2] ,
    \Tile_X1Y1_N4BEG[1] ,
    \Tile_X1Y1_N4BEG[0] }),
    .NN4END({\Tile_X1Y1_NN4BEG[15] ,
    \Tile_X1Y1_NN4BEG[14] ,
    \Tile_X1Y1_NN4BEG[13] ,
    \Tile_X1Y1_NN4BEG[12] ,
    \Tile_X1Y1_NN4BEG[11] ,
    \Tile_X1Y1_NN4BEG[10] ,
    \Tile_X1Y1_NN4BEG[9] ,
    \Tile_X1Y1_NN4BEG[8] ,
    \Tile_X1Y1_NN4BEG[7] ,
    \Tile_X1Y1_NN4BEG[6] ,
    \Tile_X1Y1_NN4BEG[5] ,
    \Tile_X1Y1_NN4BEG[4] ,
    \Tile_X1Y1_NN4BEG[3] ,
    \Tile_X1Y1_NN4BEG[2] ,
    \Tile_X1Y1_NN4BEG[1] ,
    \Tile_X1Y1_NN4BEG[0] }),
    .S1BEG({\Tile_X1Y0_S1BEG[3] ,
    \Tile_X1Y0_S1BEG[2] ,
    \Tile_X1Y0_S1BEG[1] ,
    \Tile_X1Y0_S1BEG[0] }),
    .S2BEG({\Tile_X1Y0_S2BEG[7] ,
    \Tile_X1Y0_S2BEG[6] ,
    \Tile_X1Y0_S2BEG[5] ,
    \Tile_X1Y0_S2BEG[4] ,
    \Tile_X1Y0_S2BEG[3] ,
    \Tile_X1Y0_S2BEG[2] ,
    \Tile_X1Y0_S2BEG[1] ,
    \Tile_X1Y0_S2BEG[0] }),
    .S2BEGb({\Tile_X1Y0_S2BEGb[7] ,
    \Tile_X1Y0_S2BEGb[6] ,
    \Tile_X1Y0_S2BEGb[5] ,
    \Tile_X1Y0_S2BEGb[4] ,
    \Tile_X1Y0_S2BEGb[3] ,
    \Tile_X1Y0_S2BEGb[2] ,
    \Tile_X1Y0_S2BEGb[1] ,
    \Tile_X1Y0_S2BEGb[0] }),
    .S4BEG({\Tile_X1Y0_S4BEG[15] ,
    \Tile_X1Y0_S4BEG[14] ,
    \Tile_X1Y0_S4BEG[13] ,
    \Tile_X1Y0_S4BEG[12] ,
    \Tile_X1Y0_S4BEG[11] ,
    \Tile_X1Y0_S4BEG[10] ,
    \Tile_X1Y0_S4BEG[9] ,
    \Tile_X1Y0_S4BEG[8] ,
    \Tile_X1Y0_S4BEG[7] ,
    \Tile_X1Y0_S4BEG[6] ,
    \Tile_X1Y0_S4BEG[5] ,
    \Tile_X1Y0_S4BEG[4] ,
    \Tile_X1Y0_S4BEG[3] ,
    \Tile_X1Y0_S4BEG[2] ,
    \Tile_X1Y0_S4BEG[1] ,
    \Tile_X1Y0_S4BEG[0] }),
    .SS4BEG({\Tile_X1Y0_SS4BEG[15] ,
    \Tile_X1Y0_SS4BEG[14] ,
    \Tile_X1Y0_SS4BEG[13] ,
    \Tile_X1Y0_SS4BEG[12] ,
    \Tile_X1Y0_SS4BEG[11] ,
    \Tile_X1Y0_SS4BEG[10] ,
    \Tile_X1Y0_SS4BEG[9] ,
    \Tile_X1Y0_SS4BEG[8] ,
    \Tile_X1Y0_SS4BEG[7] ,
    \Tile_X1Y0_SS4BEG[6] ,
    \Tile_X1Y0_SS4BEG[5] ,
    \Tile_X1Y0_SS4BEG[4] ,
    \Tile_X1Y0_SS4BEG[3] ,
    \Tile_X1Y0_SS4BEG[2] ,
    \Tile_X1Y0_SS4BEG[1] ,
    \Tile_X1Y0_SS4BEG[0] }));
 LUT4AB Tile_X1Y10_LUT4AB (.Ci(Tile_X1Y11_Co),
    .Co(Tile_X1Y10_Co),
    .UserCLK(Tile_X1Y11_UserCLKo),
    .UserCLKo(Tile_X1Y10_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X1Y10_E1BEG[3] ,
    \Tile_X1Y10_E1BEG[2] ,
    \Tile_X1Y10_E1BEG[1] ,
    \Tile_X1Y10_E1BEG[0] }),
    .E1END({\Tile_X0Y10_E1BEG[3] ,
    \Tile_X0Y10_E1BEG[2] ,
    \Tile_X0Y10_E1BEG[1] ,
    \Tile_X0Y10_E1BEG[0] }),
    .E2BEG({\Tile_X1Y10_E2BEG[7] ,
    \Tile_X1Y10_E2BEG[6] ,
    \Tile_X1Y10_E2BEG[5] ,
    \Tile_X1Y10_E2BEG[4] ,
    \Tile_X1Y10_E2BEG[3] ,
    \Tile_X1Y10_E2BEG[2] ,
    \Tile_X1Y10_E2BEG[1] ,
    \Tile_X1Y10_E2BEG[0] }),
    .E2BEGb({\Tile_X1Y10_E2BEGb[7] ,
    \Tile_X1Y10_E2BEGb[6] ,
    \Tile_X1Y10_E2BEGb[5] ,
    \Tile_X1Y10_E2BEGb[4] ,
    \Tile_X1Y10_E2BEGb[3] ,
    \Tile_X1Y10_E2BEGb[2] ,
    \Tile_X1Y10_E2BEGb[1] ,
    \Tile_X1Y10_E2BEGb[0] }),
    .E2END({\Tile_X0Y10_E2BEGb[7] ,
    \Tile_X0Y10_E2BEGb[6] ,
    \Tile_X0Y10_E2BEGb[5] ,
    \Tile_X0Y10_E2BEGb[4] ,
    \Tile_X0Y10_E2BEGb[3] ,
    \Tile_X0Y10_E2BEGb[2] ,
    \Tile_X0Y10_E2BEGb[1] ,
    \Tile_X0Y10_E2BEGb[0] }),
    .E2MID({\Tile_X0Y10_E2BEG[7] ,
    \Tile_X0Y10_E2BEG[6] ,
    \Tile_X0Y10_E2BEG[5] ,
    \Tile_X0Y10_E2BEG[4] ,
    \Tile_X0Y10_E2BEG[3] ,
    \Tile_X0Y10_E2BEG[2] ,
    \Tile_X0Y10_E2BEG[1] ,
    \Tile_X0Y10_E2BEG[0] }),
    .E6BEG({\Tile_X1Y10_E6BEG[11] ,
    \Tile_X1Y10_E6BEG[10] ,
    \Tile_X1Y10_E6BEG[9] ,
    \Tile_X1Y10_E6BEG[8] ,
    \Tile_X1Y10_E6BEG[7] ,
    \Tile_X1Y10_E6BEG[6] ,
    \Tile_X1Y10_E6BEG[5] ,
    \Tile_X1Y10_E6BEG[4] ,
    \Tile_X1Y10_E6BEG[3] ,
    \Tile_X1Y10_E6BEG[2] ,
    \Tile_X1Y10_E6BEG[1] ,
    \Tile_X1Y10_E6BEG[0] }),
    .E6END({\Tile_X0Y10_E6BEG[11] ,
    \Tile_X0Y10_E6BEG[10] ,
    \Tile_X0Y10_E6BEG[9] ,
    \Tile_X0Y10_E6BEG[8] ,
    \Tile_X0Y10_E6BEG[7] ,
    \Tile_X0Y10_E6BEG[6] ,
    \Tile_X0Y10_E6BEG[5] ,
    \Tile_X0Y10_E6BEG[4] ,
    \Tile_X0Y10_E6BEG[3] ,
    \Tile_X0Y10_E6BEG[2] ,
    \Tile_X0Y10_E6BEG[1] ,
    \Tile_X0Y10_E6BEG[0] }),
    .EE4BEG({\Tile_X1Y10_EE4BEG[15] ,
    \Tile_X1Y10_EE4BEG[14] ,
    \Tile_X1Y10_EE4BEG[13] ,
    \Tile_X1Y10_EE4BEG[12] ,
    \Tile_X1Y10_EE4BEG[11] ,
    \Tile_X1Y10_EE4BEG[10] ,
    \Tile_X1Y10_EE4BEG[9] ,
    \Tile_X1Y10_EE4BEG[8] ,
    \Tile_X1Y10_EE4BEG[7] ,
    \Tile_X1Y10_EE4BEG[6] ,
    \Tile_X1Y10_EE4BEG[5] ,
    \Tile_X1Y10_EE4BEG[4] ,
    \Tile_X1Y10_EE4BEG[3] ,
    \Tile_X1Y10_EE4BEG[2] ,
    \Tile_X1Y10_EE4BEG[1] ,
    \Tile_X1Y10_EE4BEG[0] }),
    .EE4END({\Tile_X0Y10_EE4BEG[15] ,
    \Tile_X0Y10_EE4BEG[14] ,
    \Tile_X0Y10_EE4BEG[13] ,
    \Tile_X0Y10_EE4BEG[12] ,
    \Tile_X0Y10_EE4BEG[11] ,
    \Tile_X0Y10_EE4BEG[10] ,
    \Tile_X0Y10_EE4BEG[9] ,
    \Tile_X0Y10_EE4BEG[8] ,
    \Tile_X0Y10_EE4BEG[7] ,
    \Tile_X0Y10_EE4BEG[6] ,
    \Tile_X0Y10_EE4BEG[5] ,
    \Tile_X0Y10_EE4BEG[4] ,
    \Tile_X0Y10_EE4BEG[3] ,
    \Tile_X0Y10_EE4BEG[2] ,
    \Tile_X0Y10_EE4BEG[1] ,
    \Tile_X0Y10_EE4BEG[0] }),
    .FrameData({\Tile_X0Y10_FrameData_O[31] ,
    \Tile_X0Y10_FrameData_O[30] ,
    \Tile_X0Y10_FrameData_O[29] ,
    \Tile_X0Y10_FrameData_O[28] ,
    \Tile_X0Y10_FrameData_O[27] ,
    \Tile_X0Y10_FrameData_O[26] ,
    \Tile_X0Y10_FrameData_O[25] ,
    \Tile_X0Y10_FrameData_O[24] ,
    \Tile_X0Y10_FrameData_O[23] ,
    \Tile_X0Y10_FrameData_O[22] ,
    \Tile_X0Y10_FrameData_O[21] ,
    \Tile_X0Y10_FrameData_O[20] ,
    \Tile_X0Y10_FrameData_O[19] ,
    \Tile_X0Y10_FrameData_O[18] ,
    \Tile_X0Y10_FrameData_O[17] ,
    \Tile_X0Y10_FrameData_O[16] ,
    \Tile_X0Y10_FrameData_O[15] ,
    \Tile_X0Y10_FrameData_O[14] ,
    \Tile_X0Y10_FrameData_O[13] ,
    \Tile_X0Y10_FrameData_O[12] ,
    \Tile_X0Y10_FrameData_O[11] ,
    \Tile_X0Y10_FrameData_O[10] ,
    \Tile_X0Y10_FrameData_O[9] ,
    \Tile_X0Y10_FrameData_O[8] ,
    \Tile_X0Y10_FrameData_O[7] ,
    \Tile_X0Y10_FrameData_O[6] ,
    \Tile_X0Y10_FrameData_O[5] ,
    \Tile_X0Y10_FrameData_O[4] ,
    \Tile_X0Y10_FrameData_O[3] ,
    \Tile_X0Y10_FrameData_O[2] ,
    \Tile_X0Y10_FrameData_O[1] ,
    \Tile_X0Y10_FrameData_O[0] }),
    .FrameData_O({\Tile_X1Y10_FrameData_O[31] ,
    \Tile_X1Y10_FrameData_O[30] ,
    \Tile_X1Y10_FrameData_O[29] ,
    \Tile_X1Y10_FrameData_O[28] ,
    \Tile_X1Y10_FrameData_O[27] ,
    \Tile_X1Y10_FrameData_O[26] ,
    \Tile_X1Y10_FrameData_O[25] ,
    \Tile_X1Y10_FrameData_O[24] ,
    \Tile_X1Y10_FrameData_O[23] ,
    \Tile_X1Y10_FrameData_O[22] ,
    \Tile_X1Y10_FrameData_O[21] ,
    \Tile_X1Y10_FrameData_O[20] ,
    \Tile_X1Y10_FrameData_O[19] ,
    \Tile_X1Y10_FrameData_O[18] ,
    \Tile_X1Y10_FrameData_O[17] ,
    \Tile_X1Y10_FrameData_O[16] ,
    \Tile_X1Y10_FrameData_O[15] ,
    \Tile_X1Y10_FrameData_O[14] ,
    \Tile_X1Y10_FrameData_O[13] ,
    \Tile_X1Y10_FrameData_O[12] ,
    \Tile_X1Y10_FrameData_O[11] ,
    \Tile_X1Y10_FrameData_O[10] ,
    \Tile_X1Y10_FrameData_O[9] ,
    \Tile_X1Y10_FrameData_O[8] ,
    \Tile_X1Y10_FrameData_O[7] ,
    \Tile_X1Y10_FrameData_O[6] ,
    \Tile_X1Y10_FrameData_O[5] ,
    \Tile_X1Y10_FrameData_O[4] ,
    \Tile_X1Y10_FrameData_O[3] ,
    \Tile_X1Y10_FrameData_O[2] ,
    \Tile_X1Y10_FrameData_O[1] ,
    \Tile_X1Y10_FrameData_O[0] }),
    .FrameStrobe({\Tile_X1Y11_FrameStrobe_O[19] ,
    \Tile_X1Y11_FrameStrobe_O[18] ,
    \Tile_X1Y11_FrameStrobe_O[17] ,
    \Tile_X1Y11_FrameStrobe_O[16] ,
    \Tile_X1Y11_FrameStrobe_O[15] ,
    \Tile_X1Y11_FrameStrobe_O[14] ,
    \Tile_X1Y11_FrameStrobe_O[13] ,
    \Tile_X1Y11_FrameStrobe_O[12] ,
    \Tile_X1Y11_FrameStrobe_O[11] ,
    \Tile_X1Y11_FrameStrobe_O[10] ,
    \Tile_X1Y11_FrameStrobe_O[9] ,
    \Tile_X1Y11_FrameStrobe_O[8] ,
    \Tile_X1Y11_FrameStrobe_O[7] ,
    \Tile_X1Y11_FrameStrobe_O[6] ,
    \Tile_X1Y11_FrameStrobe_O[5] ,
    \Tile_X1Y11_FrameStrobe_O[4] ,
    \Tile_X1Y11_FrameStrobe_O[3] ,
    \Tile_X1Y11_FrameStrobe_O[2] ,
    \Tile_X1Y11_FrameStrobe_O[1] ,
    \Tile_X1Y11_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X1Y10_FrameStrobe_O[19] ,
    \Tile_X1Y10_FrameStrobe_O[18] ,
    \Tile_X1Y10_FrameStrobe_O[17] ,
    \Tile_X1Y10_FrameStrobe_O[16] ,
    \Tile_X1Y10_FrameStrobe_O[15] ,
    \Tile_X1Y10_FrameStrobe_O[14] ,
    \Tile_X1Y10_FrameStrobe_O[13] ,
    \Tile_X1Y10_FrameStrobe_O[12] ,
    \Tile_X1Y10_FrameStrobe_O[11] ,
    \Tile_X1Y10_FrameStrobe_O[10] ,
    \Tile_X1Y10_FrameStrobe_O[9] ,
    \Tile_X1Y10_FrameStrobe_O[8] ,
    \Tile_X1Y10_FrameStrobe_O[7] ,
    \Tile_X1Y10_FrameStrobe_O[6] ,
    \Tile_X1Y10_FrameStrobe_O[5] ,
    \Tile_X1Y10_FrameStrobe_O[4] ,
    \Tile_X1Y10_FrameStrobe_O[3] ,
    \Tile_X1Y10_FrameStrobe_O[2] ,
    \Tile_X1Y10_FrameStrobe_O[1] ,
    \Tile_X1Y10_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X1Y10_N1BEG[3] ,
    \Tile_X1Y10_N1BEG[2] ,
    \Tile_X1Y10_N1BEG[1] ,
    \Tile_X1Y10_N1BEG[0] }),
    .N1END({\Tile_X1Y11_N1BEG[3] ,
    \Tile_X1Y11_N1BEG[2] ,
    \Tile_X1Y11_N1BEG[1] ,
    \Tile_X1Y11_N1BEG[0] }),
    .N2BEG({\Tile_X1Y10_N2BEG[7] ,
    \Tile_X1Y10_N2BEG[6] ,
    \Tile_X1Y10_N2BEG[5] ,
    \Tile_X1Y10_N2BEG[4] ,
    \Tile_X1Y10_N2BEG[3] ,
    \Tile_X1Y10_N2BEG[2] ,
    \Tile_X1Y10_N2BEG[1] ,
    \Tile_X1Y10_N2BEG[0] }),
    .N2BEGb({\Tile_X1Y10_N2BEGb[7] ,
    \Tile_X1Y10_N2BEGb[6] ,
    \Tile_X1Y10_N2BEGb[5] ,
    \Tile_X1Y10_N2BEGb[4] ,
    \Tile_X1Y10_N2BEGb[3] ,
    \Tile_X1Y10_N2BEGb[2] ,
    \Tile_X1Y10_N2BEGb[1] ,
    \Tile_X1Y10_N2BEGb[0] }),
    .N2END({\Tile_X1Y11_N2BEGb[7] ,
    \Tile_X1Y11_N2BEGb[6] ,
    \Tile_X1Y11_N2BEGb[5] ,
    \Tile_X1Y11_N2BEGb[4] ,
    \Tile_X1Y11_N2BEGb[3] ,
    \Tile_X1Y11_N2BEGb[2] ,
    \Tile_X1Y11_N2BEGb[1] ,
    \Tile_X1Y11_N2BEGb[0] }),
    .N2MID({\Tile_X1Y11_N2BEG[7] ,
    \Tile_X1Y11_N2BEG[6] ,
    \Tile_X1Y11_N2BEG[5] ,
    \Tile_X1Y11_N2BEG[4] ,
    \Tile_X1Y11_N2BEG[3] ,
    \Tile_X1Y11_N2BEG[2] ,
    \Tile_X1Y11_N2BEG[1] ,
    \Tile_X1Y11_N2BEG[0] }),
    .N4BEG({\Tile_X1Y10_N4BEG[15] ,
    \Tile_X1Y10_N4BEG[14] ,
    \Tile_X1Y10_N4BEG[13] ,
    \Tile_X1Y10_N4BEG[12] ,
    \Tile_X1Y10_N4BEG[11] ,
    \Tile_X1Y10_N4BEG[10] ,
    \Tile_X1Y10_N4BEG[9] ,
    \Tile_X1Y10_N4BEG[8] ,
    \Tile_X1Y10_N4BEG[7] ,
    \Tile_X1Y10_N4BEG[6] ,
    \Tile_X1Y10_N4BEG[5] ,
    \Tile_X1Y10_N4BEG[4] ,
    \Tile_X1Y10_N4BEG[3] ,
    \Tile_X1Y10_N4BEG[2] ,
    \Tile_X1Y10_N4BEG[1] ,
    \Tile_X1Y10_N4BEG[0] }),
    .N4END({\Tile_X1Y11_N4BEG[15] ,
    \Tile_X1Y11_N4BEG[14] ,
    \Tile_X1Y11_N4BEG[13] ,
    \Tile_X1Y11_N4BEG[12] ,
    \Tile_X1Y11_N4BEG[11] ,
    \Tile_X1Y11_N4BEG[10] ,
    \Tile_X1Y11_N4BEG[9] ,
    \Tile_X1Y11_N4BEG[8] ,
    \Tile_X1Y11_N4BEG[7] ,
    \Tile_X1Y11_N4BEG[6] ,
    \Tile_X1Y11_N4BEG[5] ,
    \Tile_X1Y11_N4BEG[4] ,
    \Tile_X1Y11_N4BEG[3] ,
    \Tile_X1Y11_N4BEG[2] ,
    \Tile_X1Y11_N4BEG[1] ,
    \Tile_X1Y11_N4BEG[0] }),
    .NN4BEG({\Tile_X1Y10_NN4BEG[15] ,
    \Tile_X1Y10_NN4BEG[14] ,
    \Tile_X1Y10_NN4BEG[13] ,
    \Tile_X1Y10_NN4BEG[12] ,
    \Tile_X1Y10_NN4BEG[11] ,
    \Tile_X1Y10_NN4BEG[10] ,
    \Tile_X1Y10_NN4BEG[9] ,
    \Tile_X1Y10_NN4BEG[8] ,
    \Tile_X1Y10_NN4BEG[7] ,
    \Tile_X1Y10_NN4BEG[6] ,
    \Tile_X1Y10_NN4BEG[5] ,
    \Tile_X1Y10_NN4BEG[4] ,
    \Tile_X1Y10_NN4BEG[3] ,
    \Tile_X1Y10_NN4BEG[2] ,
    \Tile_X1Y10_NN4BEG[1] ,
    \Tile_X1Y10_NN4BEG[0] }),
    .NN4END({\Tile_X1Y11_NN4BEG[15] ,
    \Tile_X1Y11_NN4BEG[14] ,
    \Tile_X1Y11_NN4BEG[13] ,
    \Tile_X1Y11_NN4BEG[12] ,
    \Tile_X1Y11_NN4BEG[11] ,
    \Tile_X1Y11_NN4BEG[10] ,
    \Tile_X1Y11_NN4BEG[9] ,
    \Tile_X1Y11_NN4BEG[8] ,
    \Tile_X1Y11_NN4BEG[7] ,
    \Tile_X1Y11_NN4BEG[6] ,
    \Tile_X1Y11_NN4BEG[5] ,
    \Tile_X1Y11_NN4BEG[4] ,
    \Tile_X1Y11_NN4BEG[3] ,
    \Tile_X1Y11_NN4BEG[2] ,
    \Tile_X1Y11_NN4BEG[1] ,
    \Tile_X1Y11_NN4BEG[0] }),
    .S1BEG({\Tile_X1Y10_S1BEG[3] ,
    \Tile_X1Y10_S1BEG[2] ,
    \Tile_X1Y10_S1BEG[1] ,
    \Tile_X1Y10_S1BEG[0] }),
    .S1END({\Tile_X1Y9_S1BEG[3] ,
    \Tile_X1Y9_S1BEG[2] ,
    \Tile_X1Y9_S1BEG[1] ,
    \Tile_X1Y9_S1BEG[0] }),
    .S2BEG({\Tile_X1Y10_S2BEG[7] ,
    \Tile_X1Y10_S2BEG[6] ,
    \Tile_X1Y10_S2BEG[5] ,
    \Tile_X1Y10_S2BEG[4] ,
    \Tile_X1Y10_S2BEG[3] ,
    \Tile_X1Y10_S2BEG[2] ,
    \Tile_X1Y10_S2BEG[1] ,
    \Tile_X1Y10_S2BEG[0] }),
    .S2BEGb({\Tile_X1Y10_S2BEGb[7] ,
    \Tile_X1Y10_S2BEGb[6] ,
    \Tile_X1Y10_S2BEGb[5] ,
    \Tile_X1Y10_S2BEGb[4] ,
    \Tile_X1Y10_S2BEGb[3] ,
    \Tile_X1Y10_S2BEGb[2] ,
    \Tile_X1Y10_S2BEGb[1] ,
    \Tile_X1Y10_S2BEGb[0] }),
    .S2END({\Tile_X1Y9_S2BEGb[7] ,
    \Tile_X1Y9_S2BEGb[6] ,
    \Tile_X1Y9_S2BEGb[5] ,
    \Tile_X1Y9_S2BEGb[4] ,
    \Tile_X1Y9_S2BEGb[3] ,
    \Tile_X1Y9_S2BEGb[2] ,
    \Tile_X1Y9_S2BEGb[1] ,
    \Tile_X1Y9_S2BEGb[0] }),
    .S2MID({\Tile_X1Y9_S2BEG[7] ,
    \Tile_X1Y9_S2BEG[6] ,
    \Tile_X1Y9_S2BEG[5] ,
    \Tile_X1Y9_S2BEG[4] ,
    \Tile_X1Y9_S2BEG[3] ,
    \Tile_X1Y9_S2BEG[2] ,
    \Tile_X1Y9_S2BEG[1] ,
    \Tile_X1Y9_S2BEG[0] }),
    .S4BEG({\Tile_X1Y10_S4BEG[15] ,
    \Tile_X1Y10_S4BEG[14] ,
    \Tile_X1Y10_S4BEG[13] ,
    \Tile_X1Y10_S4BEG[12] ,
    \Tile_X1Y10_S4BEG[11] ,
    \Tile_X1Y10_S4BEG[10] ,
    \Tile_X1Y10_S4BEG[9] ,
    \Tile_X1Y10_S4BEG[8] ,
    \Tile_X1Y10_S4BEG[7] ,
    \Tile_X1Y10_S4BEG[6] ,
    \Tile_X1Y10_S4BEG[5] ,
    \Tile_X1Y10_S4BEG[4] ,
    \Tile_X1Y10_S4BEG[3] ,
    \Tile_X1Y10_S4BEG[2] ,
    \Tile_X1Y10_S4BEG[1] ,
    \Tile_X1Y10_S4BEG[0] }),
    .S4END({\Tile_X1Y9_S4BEG[15] ,
    \Tile_X1Y9_S4BEG[14] ,
    \Tile_X1Y9_S4BEG[13] ,
    \Tile_X1Y9_S4BEG[12] ,
    \Tile_X1Y9_S4BEG[11] ,
    \Tile_X1Y9_S4BEG[10] ,
    \Tile_X1Y9_S4BEG[9] ,
    \Tile_X1Y9_S4BEG[8] ,
    \Tile_X1Y9_S4BEG[7] ,
    \Tile_X1Y9_S4BEG[6] ,
    \Tile_X1Y9_S4BEG[5] ,
    \Tile_X1Y9_S4BEG[4] ,
    \Tile_X1Y9_S4BEG[3] ,
    \Tile_X1Y9_S4BEG[2] ,
    \Tile_X1Y9_S4BEG[1] ,
    \Tile_X1Y9_S4BEG[0] }),
    .SS4BEG({\Tile_X1Y10_SS4BEG[15] ,
    \Tile_X1Y10_SS4BEG[14] ,
    \Tile_X1Y10_SS4BEG[13] ,
    \Tile_X1Y10_SS4BEG[12] ,
    \Tile_X1Y10_SS4BEG[11] ,
    \Tile_X1Y10_SS4BEG[10] ,
    \Tile_X1Y10_SS4BEG[9] ,
    \Tile_X1Y10_SS4BEG[8] ,
    \Tile_X1Y10_SS4BEG[7] ,
    \Tile_X1Y10_SS4BEG[6] ,
    \Tile_X1Y10_SS4BEG[5] ,
    \Tile_X1Y10_SS4BEG[4] ,
    \Tile_X1Y10_SS4BEG[3] ,
    \Tile_X1Y10_SS4BEG[2] ,
    \Tile_X1Y10_SS4BEG[1] ,
    \Tile_X1Y10_SS4BEG[0] }),
    .SS4END({\Tile_X1Y9_SS4BEG[15] ,
    \Tile_X1Y9_SS4BEG[14] ,
    \Tile_X1Y9_SS4BEG[13] ,
    \Tile_X1Y9_SS4BEG[12] ,
    \Tile_X1Y9_SS4BEG[11] ,
    \Tile_X1Y9_SS4BEG[10] ,
    \Tile_X1Y9_SS4BEG[9] ,
    \Tile_X1Y9_SS4BEG[8] ,
    \Tile_X1Y9_SS4BEG[7] ,
    \Tile_X1Y9_SS4BEG[6] ,
    \Tile_X1Y9_SS4BEG[5] ,
    \Tile_X1Y9_SS4BEG[4] ,
    \Tile_X1Y9_SS4BEG[3] ,
    \Tile_X1Y9_SS4BEG[2] ,
    \Tile_X1Y9_SS4BEG[1] ,
    \Tile_X1Y9_SS4BEG[0] }),
    .W1BEG({\Tile_X1Y10_W1BEG[3] ,
    \Tile_X1Y10_W1BEG[2] ,
    \Tile_X1Y10_W1BEG[1] ,
    \Tile_X1Y10_W1BEG[0] }),
    .W1END({\Tile_X2Y10_W1BEG[3] ,
    \Tile_X2Y10_W1BEG[2] ,
    \Tile_X2Y10_W1BEG[1] ,
    \Tile_X2Y10_W1BEG[0] }),
    .W2BEG({\Tile_X1Y10_W2BEG[7] ,
    \Tile_X1Y10_W2BEG[6] ,
    \Tile_X1Y10_W2BEG[5] ,
    \Tile_X1Y10_W2BEG[4] ,
    \Tile_X1Y10_W2BEG[3] ,
    \Tile_X1Y10_W2BEG[2] ,
    \Tile_X1Y10_W2BEG[1] ,
    \Tile_X1Y10_W2BEG[0] }),
    .W2BEGb({\Tile_X1Y10_W2BEGb[7] ,
    \Tile_X1Y10_W2BEGb[6] ,
    \Tile_X1Y10_W2BEGb[5] ,
    \Tile_X1Y10_W2BEGb[4] ,
    \Tile_X1Y10_W2BEGb[3] ,
    \Tile_X1Y10_W2BEGb[2] ,
    \Tile_X1Y10_W2BEGb[1] ,
    \Tile_X1Y10_W2BEGb[0] }),
    .W2END({\Tile_X2Y10_W2BEGb[7] ,
    \Tile_X2Y10_W2BEGb[6] ,
    \Tile_X2Y10_W2BEGb[5] ,
    \Tile_X2Y10_W2BEGb[4] ,
    \Tile_X2Y10_W2BEGb[3] ,
    \Tile_X2Y10_W2BEGb[2] ,
    \Tile_X2Y10_W2BEGb[1] ,
    \Tile_X2Y10_W2BEGb[0] }),
    .W2MID({\Tile_X2Y10_W2BEG[7] ,
    \Tile_X2Y10_W2BEG[6] ,
    \Tile_X2Y10_W2BEG[5] ,
    \Tile_X2Y10_W2BEG[4] ,
    \Tile_X2Y10_W2BEG[3] ,
    \Tile_X2Y10_W2BEG[2] ,
    \Tile_X2Y10_W2BEG[1] ,
    \Tile_X2Y10_W2BEG[0] }),
    .W6BEG({\Tile_X1Y10_W6BEG[11] ,
    \Tile_X1Y10_W6BEG[10] ,
    \Tile_X1Y10_W6BEG[9] ,
    \Tile_X1Y10_W6BEG[8] ,
    \Tile_X1Y10_W6BEG[7] ,
    \Tile_X1Y10_W6BEG[6] ,
    \Tile_X1Y10_W6BEG[5] ,
    \Tile_X1Y10_W6BEG[4] ,
    \Tile_X1Y10_W6BEG[3] ,
    \Tile_X1Y10_W6BEG[2] ,
    \Tile_X1Y10_W6BEG[1] ,
    \Tile_X1Y10_W6BEG[0] }),
    .W6END({\Tile_X2Y10_W6BEG[11] ,
    \Tile_X2Y10_W6BEG[10] ,
    \Tile_X2Y10_W6BEG[9] ,
    \Tile_X2Y10_W6BEG[8] ,
    \Tile_X2Y10_W6BEG[7] ,
    \Tile_X2Y10_W6BEG[6] ,
    \Tile_X2Y10_W6BEG[5] ,
    \Tile_X2Y10_W6BEG[4] ,
    \Tile_X2Y10_W6BEG[3] ,
    \Tile_X2Y10_W6BEG[2] ,
    \Tile_X2Y10_W6BEG[1] ,
    \Tile_X2Y10_W6BEG[0] }),
    .WW4BEG({\Tile_X1Y10_WW4BEG[15] ,
    \Tile_X1Y10_WW4BEG[14] ,
    \Tile_X1Y10_WW4BEG[13] ,
    \Tile_X1Y10_WW4BEG[12] ,
    \Tile_X1Y10_WW4BEG[11] ,
    \Tile_X1Y10_WW4BEG[10] ,
    \Tile_X1Y10_WW4BEG[9] ,
    \Tile_X1Y10_WW4BEG[8] ,
    \Tile_X1Y10_WW4BEG[7] ,
    \Tile_X1Y10_WW4BEG[6] ,
    \Tile_X1Y10_WW4BEG[5] ,
    \Tile_X1Y10_WW4BEG[4] ,
    \Tile_X1Y10_WW4BEG[3] ,
    \Tile_X1Y10_WW4BEG[2] ,
    \Tile_X1Y10_WW4BEG[1] ,
    \Tile_X1Y10_WW4BEG[0] }),
    .WW4END({\Tile_X2Y10_WW4BEG[15] ,
    \Tile_X2Y10_WW4BEG[14] ,
    \Tile_X2Y10_WW4BEG[13] ,
    \Tile_X2Y10_WW4BEG[12] ,
    \Tile_X2Y10_WW4BEG[11] ,
    \Tile_X2Y10_WW4BEG[10] ,
    \Tile_X2Y10_WW4BEG[9] ,
    \Tile_X2Y10_WW4BEG[8] ,
    \Tile_X2Y10_WW4BEG[7] ,
    \Tile_X2Y10_WW4BEG[6] ,
    \Tile_X2Y10_WW4BEG[5] ,
    \Tile_X2Y10_WW4BEG[4] ,
    \Tile_X2Y10_WW4BEG[3] ,
    \Tile_X2Y10_WW4BEG[2] ,
    \Tile_X2Y10_WW4BEG[1] ,
    \Tile_X2Y10_WW4BEG[0] }));
 LUT4AB Tile_X1Y11_LUT4AB (.Ci(Tile_X1Y12_Co),
    .Co(Tile_X1Y11_Co),
    .UserCLK(Tile_X1Y12_UserCLKo),
    .UserCLKo(Tile_X1Y11_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X1Y11_E1BEG[3] ,
    \Tile_X1Y11_E1BEG[2] ,
    \Tile_X1Y11_E1BEG[1] ,
    \Tile_X1Y11_E1BEG[0] }),
    .E1END({\Tile_X0Y11_E1BEG[3] ,
    \Tile_X0Y11_E1BEG[2] ,
    \Tile_X0Y11_E1BEG[1] ,
    \Tile_X0Y11_E1BEG[0] }),
    .E2BEG({\Tile_X1Y11_E2BEG[7] ,
    \Tile_X1Y11_E2BEG[6] ,
    \Tile_X1Y11_E2BEG[5] ,
    \Tile_X1Y11_E2BEG[4] ,
    \Tile_X1Y11_E2BEG[3] ,
    \Tile_X1Y11_E2BEG[2] ,
    \Tile_X1Y11_E2BEG[1] ,
    \Tile_X1Y11_E2BEG[0] }),
    .E2BEGb({\Tile_X1Y11_E2BEGb[7] ,
    \Tile_X1Y11_E2BEGb[6] ,
    \Tile_X1Y11_E2BEGb[5] ,
    \Tile_X1Y11_E2BEGb[4] ,
    \Tile_X1Y11_E2BEGb[3] ,
    \Tile_X1Y11_E2BEGb[2] ,
    \Tile_X1Y11_E2BEGb[1] ,
    \Tile_X1Y11_E2BEGb[0] }),
    .E2END({\Tile_X0Y11_E2BEGb[7] ,
    \Tile_X0Y11_E2BEGb[6] ,
    \Tile_X0Y11_E2BEGb[5] ,
    \Tile_X0Y11_E2BEGb[4] ,
    \Tile_X0Y11_E2BEGb[3] ,
    \Tile_X0Y11_E2BEGb[2] ,
    \Tile_X0Y11_E2BEGb[1] ,
    \Tile_X0Y11_E2BEGb[0] }),
    .E2MID({\Tile_X0Y11_E2BEG[7] ,
    \Tile_X0Y11_E2BEG[6] ,
    \Tile_X0Y11_E2BEG[5] ,
    \Tile_X0Y11_E2BEG[4] ,
    \Tile_X0Y11_E2BEG[3] ,
    \Tile_X0Y11_E2BEG[2] ,
    \Tile_X0Y11_E2BEG[1] ,
    \Tile_X0Y11_E2BEG[0] }),
    .E6BEG({\Tile_X1Y11_E6BEG[11] ,
    \Tile_X1Y11_E6BEG[10] ,
    \Tile_X1Y11_E6BEG[9] ,
    \Tile_X1Y11_E6BEG[8] ,
    \Tile_X1Y11_E6BEG[7] ,
    \Tile_X1Y11_E6BEG[6] ,
    \Tile_X1Y11_E6BEG[5] ,
    \Tile_X1Y11_E6BEG[4] ,
    \Tile_X1Y11_E6BEG[3] ,
    \Tile_X1Y11_E6BEG[2] ,
    \Tile_X1Y11_E6BEG[1] ,
    \Tile_X1Y11_E6BEG[0] }),
    .E6END({\Tile_X0Y11_E6BEG[11] ,
    \Tile_X0Y11_E6BEG[10] ,
    \Tile_X0Y11_E6BEG[9] ,
    \Tile_X0Y11_E6BEG[8] ,
    \Tile_X0Y11_E6BEG[7] ,
    \Tile_X0Y11_E6BEG[6] ,
    \Tile_X0Y11_E6BEG[5] ,
    \Tile_X0Y11_E6BEG[4] ,
    \Tile_X0Y11_E6BEG[3] ,
    \Tile_X0Y11_E6BEG[2] ,
    \Tile_X0Y11_E6BEG[1] ,
    \Tile_X0Y11_E6BEG[0] }),
    .EE4BEG({\Tile_X1Y11_EE4BEG[15] ,
    \Tile_X1Y11_EE4BEG[14] ,
    \Tile_X1Y11_EE4BEG[13] ,
    \Tile_X1Y11_EE4BEG[12] ,
    \Tile_X1Y11_EE4BEG[11] ,
    \Tile_X1Y11_EE4BEG[10] ,
    \Tile_X1Y11_EE4BEG[9] ,
    \Tile_X1Y11_EE4BEG[8] ,
    \Tile_X1Y11_EE4BEG[7] ,
    \Tile_X1Y11_EE4BEG[6] ,
    \Tile_X1Y11_EE4BEG[5] ,
    \Tile_X1Y11_EE4BEG[4] ,
    \Tile_X1Y11_EE4BEG[3] ,
    \Tile_X1Y11_EE4BEG[2] ,
    \Tile_X1Y11_EE4BEG[1] ,
    \Tile_X1Y11_EE4BEG[0] }),
    .EE4END({\Tile_X0Y11_EE4BEG[15] ,
    \Tile_X0Y11_EE4BEG[14] ,
    \Tile_X0Y11_EE4BEG[13] ,
    \Tile_X0Y11_EE4BEG[12] ,
    \Tile_X0Y11_EE4BEG[11] ,
    \Tile_X0Y11_EE4BEG[10] ,
    \Tile_X0Y11_EE4BEG[9] ,
    \Tile_X0Y11_EE4BEG[8] ,
    \Tile_X0Y11_EE4BEG[7] ,
    \Tile_X0Y11_EE4BEG[6] ,
    \Tile_X0Y11_EE4BEG[5] ,
    \Tile_X0Y11_EE4BEG[4] ,
    \Tile_X0Y11_EE4BEG[3] ,
    \Tile_X0Y11_EE4BEG[2] ,
    \Tile_X0Y11_EE4BEG[1] ,
    \Tile_X0Y11_EE4BEG[0] }),
    .FrameData({\Tile_X0Y11_FrameData_O[31] ,
    \Tile_X0Y11_FrameData_O[30] ,
    \Tile_X0Y11_FrameData_O[29] ,
    \Tile_X0Y11_FrameData_O[28] ,
    \Tile_X0Y11_FrameData_O[27] ,
    \Tile_X0Y11_FrameData_O[26] ,
    \Tile_X0Y11_FrameData_O[25] ,
    \Tile_X0Y11_FrameData_O[24] ,
    \Tile_X0Y11_FrameData_O[23] ,
    \Tile_X0Y11_FrameData_O[22] ,
    \Tile_X0Y11_FrameData_O[21] ,
    \Tile_X0Y11_FrameData_O[20] ,
    \Tile_X0Y11_FrameData_O[19] ,
    \Tile_X0Y11_FrameData_O[18] ,
    \Tile_X0Y11_FrameData_O[17] ,
    \Tile_X0Y11_FrameData_O[16] ,
    \Tile_X0Y11_FrameData_O[15] ,
    \Tile_X0Y11_FrameData_O[14] ,
    \Tile_X0Y11_FrameData_O[13] ,
    \Tile_X0Y11_FrameData_O[12] ,
    \Tile_X0Y11_FrameData_O[11] ,
    \Tile_X0Y11_FrameData_O[10] ,
    \Tile_X0Y11_FrameData_O[9] ,
    \Tile_X0Y11_FrameData_O[8] ,
    \Tile_X0Y11_FrameData_O[7] ,
    \Tile_X0Y11_FrameData_O[6] ,
    \Tile_X0Y11_FrameData_O[5] ,
    \Tile_X0Y11_FrameData_O[4] ,
    \Tile_X0Y11_FrameData_O[3] ,
    \Tile_X0Y11_FrameData_O[2] ,
    \Tile_X0Y11_FrameData_O[1] ,
    \Tile_X0Y11_FrameData_O[0] }),
    .FrameData_O({\Tile_X1Y11_FrameData_O[31] ,
    \Tile_X1Y11_FrameData_O[30] ,
    \Tile_X1Y11_FrameData_O[29] ,
    \Tile_X1Y11_FrameData_O[28] ,
    \Tile_X1Y11_FrameData_O[27] ,
    \Tile_X1Y11_FrameData_O[26] ,
    \Tile_X1Y11_FrameData_O[25] ,
    \Tile_X1Y11_FrameData_O[24] ,
    \Tile_X1Y11_FrameData_O[23] ,
    \Tile_X1Y11_FrameData_O[22] ,
    \Tile_X1Y11_FrameData_O[21] ,
    \Tile_X1Y11_FrameData_O[20] ,
    \Tile_X1Y11_FrameData_O[19] ,
    \Tile_X1Y11_FrameData_O[18] ,
    \Tile_X1Y11_FrameData_O[17] ,
    \Tile_X1Y11_FrameData_O[16] ,
    \Tile_X1Y11_FrameData_O[15] ,
    \Tile_X1Y11_FrameData_O[14] ,
    \Tile_X1Y11_FrameData_O[13] ,
    \Tile_X1Y11_FrameData_O[12] ,
    \Tile_X1Y11_FrameData_O[11] ,
    \Tile_X1Y11_FrameData_O[10] ,
    \Tile_X1Y11_FrameData_O[9] ,
    \Tile_X1Y11_FrameData_O[8] ,
    \Tile_X1Y11_FrameData_O[7] ,
    \Tile_X1Y11_FrameData_O[6] ,
    \Tile_X1Y11_FrameData_O[5] ,
    \Tile_X1Y11_FrameData_O[4] ,
    \Tile_X1Y11_FrameData_O[3] ,
    \Tile_X1Y11_FrameData_O[2] ,
    \Tile_X1Y11_FrameData_O[1] ,
    \Tile_X1Y11_FrameData_O[0] }),
    .FrameStrobe({\Tile_X1Y12_FrameStrobe_O[19] ,
    \Tile_X1Y12_FrameStrobe_O[18] ,
    \Tile_X1Y12_FrameStrobe_O[17] ,
    \Tile_X1Y12_FrameStrobe_O[16] ,
    \Tile_X1Y12_FrameStrobe_O[15] ,
    \Tile_X1Y12_FrameStrobe_O[14] ,
    \Tile_X1Y12_FrameStrobe_O[13] ,
    \Tile_X1Y12_FrameStrobe_O[12] ,
    \Tile_X1Y12_FrameStrobe_O[11] ,
    \Tile_X1Y12_FrameStrobe_O[10] ,
    \Tile_X1Y12_FrameStrobe_O[9] ,
    \Tile_X1Y12_FrameStrobe_O[8] ,
    \Tile_X1Y12_FrameStrobe_O[7] ,
    \Tile_X1Y12_FrameStrobe_O[6] ,
    \Tile_X1Y12_FrameStrobe_O[5] ,
    \Tile_X1Y12_FrameStrobe_O[4] ,
    \Tile_X1Y12_FrameStrobe_O[3] ,
    \Tile_X1Y12_FrameStrobe_O[2] ,
    \Tile_X1Y12_FrameStrobe_O[1] ,
    \Tile_X1Y12_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X1Y11_FrameStrobe_O[19] ,
    \Tile_X1Y11_FrameStrobe_O[18] ,
    \Tile_X1Y11_FrameStrobe_O[17] ,
    \Tile_X1Y11_FrameStrobe_O[16] ,
    \Tile_X1Y11_FrameStrobe_O[15] ,
    \Tile_X1Y11_FrameStrobe_O[14] ,
    \Tile_X1Y11_FrameStrobe_O[13] ,
    \Tile_X1Y11_FrameStrobe_O[12] ,
    \Tile_X1Y11_FrameStrobe_O[11] ,
    \Tile_X1Y11_FrameStrobe_O[10] ,
    \Tile_X1Y11_FrameStrobe_O[9] ,
    \Tile_X1Y11_FrameStrobe_O[8] ,
    \Tile_X1Y11_FrameStrobe_O[7] ,
    \Tile_X1Y11_FrameStrobe_O[6] ,
    \Tile_X1Y11_FrameStrobe_O[5] ,
    \Tile_X1Y11_FrameStrobe_O[4] ,
    \Tile_X1Y11_FrameStrobe_O[3] ,
    \Tile_X1Y11_FrameStrobe_O[2] ,
    \Tile_X1Y11_FrameStrobe_O[1] ,
    \Tile_X1Y11_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X1Y11_N1BEG[3] ,
    \Tile_X1Y11_N1BEG[2] ,
    \Tile_X1Y11_N1BEG[1] ,
    \Tile_X1Y11_N1BEG[0] }),
    .N1END({\Tile_X1Y12_N1BEG[3] ,
    \Tile_X1Y12_N1BEG[2] ,
    \Tile_X1Y12_N1BEG[1] ,
    \Tile_X1Y12_N1BEG[0] }),
    .N2BEG({\Tile_X1Y11_N2BEG[7] ,
    \Tile_X1Y11_N2BEG[6] ,
    \Tile_X1Y11_N2BEG[5] ,
    \Tile_X1Y11_N2BEG[4] ,
    \Tile_X1Y11_N2BEG[3] ,
    \Tile_X1Y11_N2BEG[2] ,
    \Tile_X1Y11_N2BEG[1] ,
    \Tile_X1Y11_N2BEG[0] }),
    .N2BEGb({\Tile_X1Y11_N2BEGb[7] ,
    \Tile_X1Y11_N2BEGb[6] ,
    \Tile_X1Y11_N2BEGb[5] ,
    \Tile_X1Y11_N2BEGb[4] ,
    \Tile_X1Y11_N2BEGb[3] ,
    \Tile_X1Y11_N2BEGb[2] ,
    \Tile_X1Y11_N2BEGb[1] ,
    \Tile_X1Y11_N2BEGb[0] }),
    .N2END({\Tile_X1Y12_N2BEGb[7] ,
    \Tile_X1Y12_N2BEGb[6] ,
    \Tile_X1Y12_N2BEGb[5] ,
    \Tile_X1Y12_N2BEGb[4] ,
    \Tile_X1Y12_N2BEGb[3] ,
    \Tile_X1Y12_N2BEGb[2] ,
    \Tile_X1Y12_N2BEGb[1] ,
    \Tile_X1Y12_N2BEGb[0] }),
    .N2MID({\Tile_X1Y12_N2BEG[7] ,
    \Tile_X1Y12_N2BEG[6] ,
    \Tile_X1Y12_N2BEG[5] ,
    \Tile_X1Y12_N2BEG[4] ,
    \Tile_X1Y12_N2BEG[3] ,
    \Tile_X1Y12_N2BEG[2] ,
    \Tile_X1Y12_N2BEG[1] ,
    \Tile_X1Y12_N2BEG[0] }),
    .N4BEG({\Tile_X1Y11_N4BEG[15] ,
    \Tile_X1Y11_N4BEG[14] ,
    \Tile_X1Y11_N4BEG[13] ,
    \Tile_X1Y11_N4BEG[12] ,
    \Tile_X1Y11_N4BEG[11] ,
    \Tile_X1Y11_N4BEG[10] ,
    \Tile_X1Y11_N4BEG[9] ,
    \Tile_X1Y11_N4BEG[8] ,
    \Tile_X1Y11_N4BEG[7] ,
    \Tile_X1Y11_N4BEG[6] ,
    \Tile_X1Y11_N4BEG[5] ,
    \Tile_X1Y11_N4BEG[4] ,
    \Tile_X1Y11_N4BEG[3] ,
    \Tile_X1Y11_N4BEG[2] ,
    \Tile_X1Y11_N4BEG[1] ,
    \Tile_X1Y11_N4BEG[0] }),
    .N4END({\Tile_X1Y12_N4BEG[15] ,
    \Tile_X1Y12_N4BEG[14] ,
    \Tile_X1Y12_N4BEG[13] ,
    \Tile_X1Y12_N4BEG[12] ,
    \Tile_X1Y12_N4BEG[11] ,
    \Tile_X1Y12_N4BEG[10] ,
    \Tile_X1Y12_N4BEG[9] ,
    \Tile_X1Y12_N4BEG[8] ,
    \Tile_X1Y12_N4BEG[7] ,
    \Tile_X1Y12_N4BEG[6] ,
    \Tile_X1Y12_N4BEG[5] ,
    \Tile_X1Y12_N4BEG[4] ,
    \Tile_X1Y12_N4BEG[3] ,
    \Tile_X1Y12_N4BEG[2] ,
    \Tile_X1Y12_N4BEG[1] ,
    \Tile_X1Y12_N4BEG[0] }),
    .NN4BEG({\Tile_X1Y11_NN4BEG[15] ,
    \Tile_X1Y11_NN4BEG[14] ,
    \Tile_X1Y11_NN4BEG[13] ,
    \Tile_X1Y11_NN4BEG[12] ,
    \Tile_X1Y11_NN4BEG[11] ,
    \Tile_X1Y11_NN4BEG[10] ,
    \Tile_X1Y11_NN4BEG[9] ,
    \Tile_X1Y11_NN4BEG[8] ,
    \Tile_X1Y11_NN4BEG[7] ,
    \Tile_X1Y11_NN4BEG[6] ,
    \Tile_X1Y11_NN4BEG[5] ,
    \Tile_X1Y11_NN4BEG[4] ,
    \Tile_X1Y11_NN4BEG[3] ,
    \Tile_X1Y11_NN4BEG[2] ,
    \Tile_X1Y11_NN4BEG[1] ,
    \Tile_X1Y11_NN4BEG[0] }),
    .NN4END({\Tile_X1Y12_NN4BEG[15] ,
    \Tile_X1Y12_NN4BEG[14] ,
    \Tile_X1Y12_NN4BEG[13] ,
    \Tile_X1Y12_NN4BEG[12] ,
    \Tile_X1Y12_NN4BEG[11] ,
    \Tile_X1Y12_NN4BEG[10] ,
    \Tile_X1Y12_NN4BEG[9] ,
    \Tile_X1Y12_NN4BEG[8] ,
    \Tile_X1Y12_NN4BEG[7] ,
    \Tile_X1Y12_NN4BEG[6] ,
    \Tile_X1Y12_NN4BEG[5] ,
    \Tile_X1Y12_NN4BEG[4] ,
    \Tile_X1Y12_NN4BEG[3] ,
    \Tile_X1Y12_NN4BEG[2] ,
    \Tile_X1Y12_NN4BEG[1] ,
    \Tile_X1Y12_NN4BEG[0] }),
    .S1BEG({\Tile_X1Y11_S1BEG[3] ,
    \Tile_X1Y11_S1BEG[2] ,
    \Tile_X1Y11_S1BEG[1] ,
    \Tile_X1Y11_S1BEG[0] }),
    .S1END({\Tile_X1Y10_S1BEG[3] ,
    \Tile_X1Y10_S1BEG[2] ,
    \Tile_X1Y10_S1BEG[1] ,
    \Tile_X1Y10_S1BEG[0] }),
    .S2BEG({\Tile_X1Y11_S2BEG[7] ,
    \Tile_X1Y11_S2BEG[6] ,
    \Tile_X1Y11_S2BEG[5] ,
    \Tile_X1Y11_S2BEG[4] ,
    \Tile_X1Y11_S2BEG[3] ,
    \Tile_X1Y11_S2BEG[2] ,
    \Tile_X1Y11_S2BEG[1] ,
    \Tile_X1Y11_S2BEG[0] }),
    .S2BEGb({\Tile_X1Y11_S2BEGb[7] ,
    \Tile_X1Y11_S2BEGb[6] ,
    \Tile_X1Y11_S2BEGb[5] ,
    \Tile_X1Y11_S2BEGb[4] ,
    \Tile_X1Y11_S2BEGb[3] ,
    \Tile_X1Y11_S2BEGb[2] ,
    \Tile_X1Y11_S2BEGb[1] ,
    \Tile_X1Y11_S2BEGb[0] }),
    .S2END({\Tile_X1Y10_S2BEGb[7] ,
    \Tile_X1Y10_S2BEGb[6] ,
    \Tile_X1Y10_S2BEGb[5] ,
    \Tile_X1Y10_S2BEGb[4] ,
    \Tile_X1Y10_S2BEGb[3] ,
    \Tile_X1Y10_S2BEGb[2] ,
    \Tile_X1Y10_S2BEGb[1] ,
    \Tile_X1Y10_S2BEGb[0] }),
    .S2MID({\Tile_X1Y10_S2BEG[7] ,
    \Tile_X1Y10_S2BEG[6] ,
    \Tile_X1Y10_S2BEG[5] ,
    \Tile_X1Y10_S2BEG[4] ,
    \Tile_X1Y10_S2BEG[3] ,
    \Tile_X1Y10_S2BEG[2] ,
    \Tile_X1Y10_S2BEG[1] ,
    \Tile_X1Y10_S2BEG[0] }),
    .S4BEG({\Tile_X1Y11_S4BEG[15] ,
    \Tile_X1Y11_S4BEG[14] ,
    \Tile_X1Y11_S4BEG[13] ,
    \Tile_X1Y11_S4BEG[12] ,
    \Tile_X1Y11_S4BEG[11] ,
    \Tile_X1Y11_S4BEG[10] ,
    \Tile_X1Y11_S4BEG[9] ,
    \Tile_X1Y11_S4BEG[8] ,
    \Tile_X1Y11_S4BEG[7] ,
    \Tile_X1Y11_S4BEG[6] ,
    \Tile_X1Y11_S4BEG[5] ,
    \Tile_X1Y11_S4BEG[4] ,
    \Tile_X1Y11_S4BEG[3] ,
    \Tile_X1Y11_S4BEG[2] ,
    \Tile_X1Y11_S4BEG[1] ,
    \Tile_X1Y11_S4BEG[0] }),
    .S4END({\Tile_X1Y10_S4BEG[15] ,
    \Tile_X1Y10_S4BEG[14] ,
    \Tile_X1Y10_S4BEG[13] ,
    \Tile_X1Y10_S4BEG[12] ,
    \Tile_X1Y10_S4BEG[11] ,
    \Tile_X1Y10_S4BEG[10] ,
    \Tile_X1Y10_S4BEG[9] ,
    \Tile_X1Y10_S4BEG[8] ,
    \Tile_X1Y10_S4BEG[7] ,
    \Tile_X1Y10_S4BEG[6] ,
    \Tile_X1Y10_S4BEG[5] ,
    \Tile_X1Y10_S4BEG[4] ,
    \Tile_X1Y10_S4BEG[3] ,
    \Tile_X1Y10_S4BEG[2] ,
    \Tile_X1Y10_S4BEG[1] ,
    \Tile_X1Y10_S4BEG[0] }),
    .SS4BEG({\Tile_X1Y11_SS4BEG[15] ,
    \Tile_X1Y11_SS4BEG[14] ,
    \Tile_X1Y11_SS4BEG[13] ,
    \Tile_X1Y11_SS4BEG[12] ,
    \Tile_X1Y11_SS4BEG[11] ,
    \Tile_X1Y11_SS4BEG[10] ,
    \Tile_X1Y11_SS4BEG[9] ,
    \Tile_X1Y11_SS4BEG[8] ,
    \Tile_X1Y11_SS4BEG[7] ,
    \Tile_X1Y11_SS4BEG[6] ,
    \Tile_X1Y11_SS4BEG[5] ,
    \Tile_X1Y11_SS4BEG[4] ,
    \Tile_X1Y11_SS4BEG[3] ,
    \Tile_X1Y11_SS4BEG[2] ,
    \Tile_X1Y11_SS4BEG[1] ,
    \Tile_X1Y11_SS4BEG[0] }),
    .SS4END({\Tile_X1Y10_SS4BEG[15] ,
    \Tile_X1Y10_SS4BEG[14] ,
    \Tile_X1Y10_SS4BEG[13] ,
    \Tile_X1Y10_SS4BEG[12] ,
    \Tile_X1Y10_SS4BEG[11] ,
    \Tile_X1Y10_SS4BEG[10] ,
    \Tile_X1Y10_SS4BEG[9] ,
    \Tile_X1Y10_SS4BEG[8] ,
    \Tile_X1Y10_SS4BEG[7] ,
    \Tile_X1Y10_SS4BEG[6] ,
    \Tile_X1Y10_SS4BEG[5] ,
    \Tile_X1Y10_SS4BEG[4] ,
    \Tile_X1Y10_SS4BEG[3] ,
    \Tile_X1Y10_SS4BEG[2] ,
    \Tile_X1Y10_SS4BEG[1] ,
    \Tile_X1Y10_SS4BEG[0] }),
    .W1BEG({\Tile_X1Y11_W1BEG[3] ,
    \Tile_X1Y11_W1BEG[2] ,
    \Tile_X1Y11_W1BEG[1] ,
    \Tile_X1Y11_W1BEG[0] }),
    .W1END({\Tile_X2Y11_W1BEG[3] ,
    \Tile_X2Y11_W1BEG[2] ,
    \Tile_X2Y11_W1BEG[1] ,
    \Tile_X2Y11_W1BEG[0] }),
    .W2BEG({\Tile_X1Y11_W2BEG[7] ,
    \Tile_X1Y11_W2BEG[6] ,
    \Tile_X1Y11_W2BEG[5] ,
    \Tile_X1Y11_W2BEG[4] ,
    \Tile_X1Y11_W2BEG[3] ,
    \Tile_X1Y11_W2BEG[2] ,
    \Tile_X1Y11_W2BEG[1] ,
    \Tile_X1Y11_W2BEG[0] }),
    .W2BEGb({\Tile_X1Y11_W2BEGb[7] ,
    \Tile_X1Y11_W2BEGb[6] ,
    \Tile_X1Y11_W2BEGb[5] ,
    \Tile_X1Y11_W2BEGb[4] ,
    \Tile_X1Y11_W2BEGb[3] ,
    \Tile_X1Y11_W2BEGb[2] ,
    \Tile_X1Y11_W2BEGb[1] ,
    \Tile_X1Y11_W2BEGb[0] }),
    .W2END({\Tile_X2Y11_W2BEGb[7] ,
    \Tile_X2Y11_W2BEGb[6] ,
    \Tile_X2Y11_W2BEGb[5] ,
    \Tile_X2Y11_W2BEGb[4] ,
    \Tile_X2Y11_W2BEGb[3] ,
    \Tile_X2Y11_W2BEGb[2] ,
    \Tile_X2Y11_W2BEGb[1] ,
    \Tile_X2Y11_W2BEGb[0] }),
    .W2MID({\Tile_X2Y11_W2BEG[7] ,
    \Tile_X2Y11_W2BEG[6] ,
    \Tile_X2Y11_W2BEG[5] ,
    \Tile_X2Y11_W2BEG[4] ,
    \Tile_X2Y11_W2BEG[3] ,
    \Tile_X2Y11_W2BEG[2] ,
    \Tile_X2Y11_W2BEG[1] ,
    \Tile_X2Y11_W2BEG[0] }),
    .W6BEG({\Tile_X1Y11_W6BEG[11] ,
    \Tile_X1Y11_W6BEG[10] ,
    \Tile_X1Y11_W6BEG[9] ,
    \Tile_X1Y11_W6BEG[8] ,
    \Tile_X1Y11_W6BEG[7] ,
    \Tile_X1Y11_W6BEG[6] ,
    \Tile_X1Y11_W6BEG[5] ,
    \Tile_X1Y11_W6BEG[4] ,
    \Tile_X1Y11_W6BEG[3] ,
    \Tile_X1Y11_W6BEG[2] ,
    \Tile_X1Y11_W6BEG[1] ,
    \Tile_X1Y11_W6BEG[0] }),
    .W6END({\Tile_X2Y11_W6BEG[11] ,
    \Tile_X2Y11_W6BEG[10] ,
    \Tile_X2Y11_W6BEG[9] ,
    \Tile_X2Y11_W6BEG[8] ,
    \Tile_X2Y11_W6BEG[7] ,
    \Tile_X2Y11_W6BEG[6] ,
    \Tile_X2Y11_W6BEG[5] ,
    \Tile_X2Y11_W6BEG[4] ,
    \Tile_X2Y11_W6BEG[3] ,
    \Tile_X2Y11_W6BEG[2] ,
    \Tile_X2Y11_W6BEG[1] ,
    \Tile_X2Y11_W6BEG[0] }),
    .WW4BEG({\Tile_X1Y11_WW4BEG[15] ,
    \Tile_X1Y11_WW4BEG[14] ,
    \Tile_X1Y11_WW4BEG[13] ,
    \Tile_X1Y11_WW4BEG[12] ,
    \Tile_X1Y11_WW4BEG[11] ,
    \Tile_X1Y11_WW4BEG[10] ,
    \Tile_X1Y11_WW4BEG[9] ,
    \Tile_X1Y11_WW4BEG[8] ,
    \Tile_X1Y11_WW4BEG[7] ,
    \Tile_X1Y11_WW4BEG[6] ,
    \Tile_X1Y11_WW4BEG[5] ,
    \Tile_X1Y11_WW4BEG[4] ,
    \Tile_X1Y11_WW4BEG[3] ,
    \Tile_X1Y11_WW4BEG[2] ,
    \Tile_X1Y11_WW4BEG[1] ,
    \Tile_X1Y11_WW4BEG[0] }),
    .WW4END({\Tile_X2Y11_WW4BEG[15] ,
    \Tile_X2Y11_WW4BEG[14] ,
    \Tile_X2Y11_WW4BEG[13] ,
    \Tile_X2Y11_WW4BEG[12] ,
    \Tile_X2Y11_WW4BEG[11] ,
    \Tile_X2Y11_WW4BEG[10] ,
    \Tile_X2Y11_WW4BEG[9] ,
    \Tile_X2Y11_WW4BEG[8] ,
    \Tile_X2Y11_WW4BEG[7] ,
    \Tile_X2Y11_WW4BEG[6] ,
    \Tile_X2Y11_WW4BEG[5] ,
    \Tile_X2Y11_WW4BEG[4] ,
    \Tile_X2Y11_WW4BEG[3] ,
    \Tile_X2Y11_WW4BEG[2] ,
    \Tile_X2Y11_WW4BEG[1] ,
    \Tile_X2Y11_WW4BEG[0] }));
 LUT4AB Tile_X1Y12_LUT4AB (.Ci(Tile_X1Y13_Co),
    .Co(Tile_X1Y12_Co),
    .UserCLK(Tile_X1Y13_UserCLKo),
    .UserCLKo(Tile_X1Y12_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X1Y12_E1BEG[3] ,
    \Tile_X1Y12_E1BEG[2] ,
    \Tile_X1Y12_E1BEG[1] ,
    \Tile_X1Y12_E1BEG[0] }),
    .E1END({\Tile_X0Y12_E1BEG[3] ,
    \Tile_X0Y12_E1BEG[2] ,
    \Tile_X0Y12_E1BEG[1] ,
    \Tile_X0Y12_E1BEG[0] }),
    .E2BEG({\Tile_X1Y12_E2BEG[7] ,
    \Tile_X1Y12_E2BEG[6] ,
    \Tile_X1Y12_E2BEG[5] ,
    \Tile_X1Y12_E2BEG[4] ,
    \Tile_X1Y12_E2BEG[3] ,
    \Tile_X1Y12_E2BEG[2] ,
    \Tile_X1Y12_E2BEG[1] ,
    \Tile_X1Y12_E2BEG[0] }),
    .E2BEGb({\Tile_X1Y12_E2BEGb[7] ,
    \Tile_X1Y12_E2BEGb[6] ,
    \Tile_X1Y12_E2BEGb[5] ,
    \Tile_X1Y12_E2BEGb[4] ,
    \Tile_X1Y12_E2BEGb[3] ,
    \Tile_X1Y12_E2BEGb[2] ,
    \Tile_X1Y12_E2BEGb[1] ,
    \Tile_X1Y12_E2BEGb[0] }),
    .E2END({\Tile_X0Y12_E2BEGb[7] ,
    \Tile_X0Y12_E2BEGb[6] ,
    \Tile_X0Y12_E2BEGb[5] ,
    \Tile_X0Y12_E2BEGb[4] ,
    \Tile_X0Y12_E2BEGb[3] ,
    \Tile_X0Y12_E2BEGb[2] ,
    \Tile_X0Y12_E2BEGb[1] ,
    \Tile_X0Y12_E2BEGb[0] }),
    .E2MID({\Tile_X0Y12_E2BEG[7] ,
    \Tile_X0Y12_E2BEG[6] ,
    \Tile_X0Y12_E2BEG[5] ,
    \Tile_X0Y12_E2BEG[4] ,
    \Tile_X0Y12_E2BEG[3] ,
    \Tile_X0Y12_E2BEG[2] ,
    \Tile_X0Y12_E2BEG[1] ,
    \Tile_X0Y12_E2BEG[0] }),
    .E6BEG({\Tile_X1Y12_E6BEG[11] ,
    \Tile_X1Y12_E6BEG[10] ,
    \Tile_X1Y12_E6BEG[9] ,
    \Tile_X1Y12_E6BEG[8] ,
    \Tile_X1Y12_E6BEG[7] ,
    \Tile_X1Y12_E6BEG[6] ,
    \Tile_X1Y12_E6BEG[5] ,
    \Tile_X1Y12_E6BEG[4] ,
    \Tile_X1Y12_E6BEG[3] ,
    \Tile_X1Y12_E6BEG[2] ,
    \Tile_X1Y12_E6BEG[1] ,
    \Tile_X1Y12_E6BEG[0] }),
    .E6END({\Tile_X0Y12_E6BEG[11] ,
    \Tile_X0Y12_E6BEG[10] ,
    \Tile_X0Y12_E6BEG[9] ,
    \Tile_X0Y12_E6BEG[8] ,
    \Tile_X0Y12_E6BEG[7] ,
    \Tile_X0Y12_E6BEG[6] ,
    \Tile_X0Y12_E6BEG[5] ,
    \Tile_X0Y12_E6BEG[4] ,
    \Tile_X0Y12_E6BEG[3] ,
    \Tile_X0Y12_E6BEG[2] ,
    \Tile_X0Y12_E6BEG[1] ,
    \Tile_X0Y12_E6BEG[0] }),
    .EE4BEG({\Tile_X1Y12_EE4BEG[15] ,
    \Tile_X1Y12_EE4BEG[14] ,
    \Tile_X1Y12_EE4BEG[13] ,
    \Tile_X1Y12_EE4BEG[12] ,
    \Tile_X1Y12_EE4BEG[11] ,
    \Tile_X1Y12_EE4BEG[10] ,
    \Tile_X1Y12_EE4BEG[9] ,
    \Tile_X1Y12_EE4BEG[8] ,
    \Tile_X1Y12_EE4BEG[7] ,
    \Tile_X1Y12_EE4BEG[6] ,
    \Tile_X1Y12_EE4BEG[5] ,
    \Tile_X1Y12_EE4BEG[4] ,
    \Tile_X1Y12_EE4BEG[3] ,
    \Tile_X1Y12_EE4BEG[2] ,
    \Tile_X1Y12_EE4BEG[1] ,
    \Tile_X1Y12_EE4BEG[0] }),
    .EE4END({\Tile_X0Y12_EE4BEG[15] ,
    \Tile_X0Y12_EE4BEG[14] ,
    \Tile_X0Y12_EE4BEG[13] ,
    \Tile_X0Y12_EE4BEG[12] ,
    \Tile_X0Y12_EE4BEG[11] ,
    \Tile_X0Y12_EE4BEG[10] ,
    \Tile_X0Y12_EE4BEG[9] ,
    \Tile_X0Y12_EE4BEG[8] ,
    \Tile_X0Y12_EE4BEG[7] ,
    \Tile_X0Y12_EE4BEG[6] ,
    \Tile_X0Y12_EE4BEG[5] ,
    \Tile_X0Y12_EE4BEG[4] ,
    \Tile_X0Y12_EE4BEG[3] ,
    \Tile_X0Y12_EE4BEG[2] ,
    \Tile_X0Y12_EE4BEG[1] ,
    \Tile_X0Y12_EE4BEG[0] }),
    .FrameData({\Tile_X0Y12_FrameData_O[31] ,
    \Tile_X0Y12_FrameData_O[30] ,
    \Tile_X0Y12_FrameData_O[29] ,
    \Tile_X0Y12_FrameData_O[28] ,
    \Tile_X0Y12_FrameData_O[27] ,
    \Tile_X0Y12_FrameData_O[26] ,
    \Tile_X0Y12_FrameData_O[25] ,
    \Tile_X0Y12_FrameData_O[24] ,
    \Tile_X0Y12_FrameData_O[23] ,
    \Tile_X0Y12_FrameData_O[22] ,
    \Tile_X0Y12_FrameData_O[21] ,
    \Tile_X0Y12_FrameData_O[20] ,
    \Tile_X0Y12_FrameData_O[19] ,
    \Tile_X0Y12_FrameData_O[18] ,
    \Tile_X0Y12_FrameData_O[17] ,
    \Tile_X0Y12_FrameData_O[16] ,
    \Tile_X0Y12_FrameData_O[15] ,
    \Tile_X0Y12_FrameData_O[14] ,
    \Tile_X0Y12_FrameData_O[13] ,
    \Tile_X0Y12_FrameData_O[12] ,
    \Tile_X0Y12_FrameData_O[11] ,
    \Tile_X0Y12_FrameData_O[10] ,
    \Tile_X0Y12_FrameData_O[9] ,
    \Tile_X0Y12_FrameData_O[8] ,
    \Tile_X0Y12_FrameData_O[7] ,
    \Tile_X0Y12_FrameData_O[6] ,
    \Tile_X0Y12_FrameData_O[5] ,
    \Tile_X0Y12_FrameData_O[4] ,
    \Tile_X0Y12_FrameData_O[3] ,
    \Tile_X0Y12_FrameData_O[2] ,
    \Tile_X0Y12_FrameData_O[1] ,
    \Tile_X0Y12_FrameData_O[0] }),
    .FrameData_O({\Tile_X1Y12_FrameData_O[31] ,
    \Tile_X1Y12_FrameData_O[30] ,
    \Tile_X1Y12_FrameData_O[29] ,
    \Tile_X1Y12_FrameData_O[28] ,
    \Tile_X1Y12_FrameData_O[27] ,
    \Tile_X1Y12_FrameData_O[26] ,
    \Tile_X1Y12_FrameData_O[25] ,
    \Tile_X1Y12_FrameData_O[24] ,
    \Tile_X1Y12_FrameData_O[23] ,
    \Tile_X1Y12_FrameData_O[22] ,
    \Tile_X1Y12_FrameData_O[21] ,
    \Tile_X1Y12_FrameData_O[20] ,
    \Tile_X1Y12_FrameData_O[19] ,
    \Tile_X1Y12_FrameData_O[18] ,
    \Tile_X1Y12_FrameData_O[17] ,
    \Tile_X1Y12_FrameData_O[16] ,
    \Tile_X1Y12_FrameData_O[15] ,
    \Tile_X1Y12_FrameData_O[14] ,
    \Tile_X1Y12_FrameData_O[13] ,
    \Tile_X1Y12_FrameData_O[12] ,
    \Tile_X1Y12_FrameData_O[11] ,
    \Tile_X1Y12_FrameData_O[10] ,
    \Tile_X1Y12_FrameData_O[9] ,
    \Tile_X1Y12_FrameData_O[8] ,
    \Tile_X1Y12_FrameData_O[7] ,
    \Tile_X1Y12_FrameData_O[6] ,
    \Tile_X1Y12_FrameData_O[5] ,
    \Tile_X1Y12_FrameData_O[4] ,
    \Tile_X1Y12_FrameData_O[3] ,
    \Tile_X1Y12_FrameData_O[2] ,
    \Tile_X1Y12_FrameData_O[1] ,
    \Tile_X1Y12_FrameData_O[0] }),
    .FrameStrobe({\Tile_X1Y13_FrameStrobe_O[19] ,
    \Tile_X1Y13_FrameStrobe_O[18] ,
    \Tile_X1Y13_FrameStrobe_O[17] ,
    \Tile_X1Y13_FrameStrobe_O[16] ,
    \Tile_X1Y13_FrameStrobe_O[15] ,
    \Tile_X1Y13_FrameStrobe_O[14] ,
    \Tile_X1Y13_FrameStrobe_O[13] ,
    \Tile_X1Y13_FrameStrobe_O[12] ,
    \Tile_X1Y13_FrameStrobe_O[11] ,
    \Tile_X1Y13_FrameStrobe_O[10] ,
    \Tile_X1Y13_FrameStrobe_O[9] ,
    \Tile_X1Y13_FrameStrobe_O[8] ,
    \Tile_X1Y13_FrameStrobe_O[7] ,
    \Tile_X1Y13_FrameStrobe_O[6] ,
    \Tile_X1Y13_FrameStrobe_O[5] ,
    \Tile_X1Y13_FrameStrobe_O[4] ,
    \Tile_X1Y13_FrameStrobe_O[3] ,
    \Tile_X1Y13_FrameStrobe_O[2] ,
    \Tile_X1Y13_FrameStrobe_O[1] ,
    \Tile_X1Y13_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X1Y12_FrameStrobe_O[19] ,
    \Tile_X1Y12_FrameStrobe_O[18] ,
    \Tile_X1Y12_FrameStrobe_O[17] ,
    \Tile_X1Y12_FrameStrobe_O[16] ,
    \Tile_X1Y12_FrameStrobe_O[15] ,
    \Tile_X1Y12_FrameStrobe_O[14] ,
    \Tile_X1Y12_FrameStrobe_O[13] ,
    \Tile_X1Y12_FrameStrobe_O[12] ,
    \Tile_X1Y12_FrameStrobe_O[11] ,
    \Tile_X1Y12_FrameStrobe_O[10] ,
    \Tile_X1Y12_FrameStrobe_O[9] ,
    \Tile_X1Y12_FrameStrobe_O[8] ,
    \Tile_X1Y12_FrameStrobe_O[7] ,
    \Tile_X1Y12_FrameStrobe_O[6] ,
    \Tile_X1Y12_FrameStrobe_O[5] ,
    \Tile_X1Y12_FrameStrobe_O[4] ,
    \Tile_X1Y12_FrameStrobe_O[3] ,
    \Tile_X1Y12_FrameStrobe_O[2] ,
    \Tile_X1Y12_FrameStrobe_O[1] ,
    \Tile_X1Y12_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X1Y12_N1BEG[3] ,
    \Tile_X1Y12_N1BEG[2] ,
    \Tile_X1Y12_N1BEG[1] ,
    \Tile_X1Y12_N1BEG[0] }),
    .N1END({\Tile_X1Y13_N1BEG[3] ,
    \Tile_X1Y13_N1BEG[2] ,
    \Tile_X1Y13_N1BEG[1] ,
    \Tile_X1Y13_N1BEG[0] }),
    .N2BEG({\Tile_X1Y12_N2BEG[7] ,
    \Tile_X1Y12_N2BEG[6] ,
    \Tile_X1Y12_N2BEG[5] ,
    \Tile_X1Y12_N2BEG[4] ,
    \Tile_X1Y12_N2BEG[3] ,
    \Tile_X1Y12_N2BEG[2] ,
    \Tile_X1Y12_N2BEG[1] ,
    \Tile_X1Y12_N2BEG[0] }),
    .N2BEGb({\Tile_X1Y12_N2BEGb[7] ,
    \Tile_X1Y12_N2BEGb[6] ,
    \Tile_X1Y12_N2BEGb[5] ,
    \Tile_X1Y12_N2BEGb[4] ,
    \Tile_X1Y12_N2BEGb[3] ,
    \Tile_X1Y12_N2BEGb[2] ,
    \Tile_X1Y12_N2BEGb[1] ,
    \Tile_X1Y12_N2BEGb[0] }),
    .N2END({\Tile_X1Y13_N2BEGb[7] ,
    \Tile_X1Y13_N2BEGb[6] ,
    \Tile_X1Y13_N2BEGb[5] ,
    \Tile_X1Y13_N2BEGb[4] ,
    \Tile_X1Y13_N2BEGb[3] ,
    \Tile_X1Y13_N2BEGb[2] ,
    \Tile_X1Y13_N2BEGb[1] ,
    \Tile_X1Y13_N2BEGb[0] }),
    .N2MID({\Tile_X1Y13_N2BEG[7] ,
    \Tile_X1Y13_N2BEG[6] ,
    \Tile_X1Y13_N2BEG[5] ,
    \Tile_X1Y13_N2BEG[4] ,
    \Tile_X1Y13_N2BEG[3] ,
    \Tile_X1Y13_N2BEG[2] ,
    \Tile_X1Y13_N2BEG[1] ,
    \Tile_X1Y13_N2BEG[0] }),
    .N4BEG({\Tile_X1Y12_N4BEG[15] ,
    \Tile_X1Y12_N4BEG[14] ,
    \Tile_X1Y12_N4BEG[13] ,
    \Tile_X1Y12_N4BEG[12] ,
    \Tile_X1Y12_N4BEG[11] ,
    \Tile_X1Y12_N4BEG[10] ,
    \Tile_X1Y12_N4BEG[9] ,
    \Tile_X1Y12_N4BEG[8] ,
    \Tile_X1Y12_N4BEG[7] ,
    \Tile_X1Y12_N4BEG[6] ,
    \Tile_X1Y12_N4BEG[5] ,
    \Tile_X1Y12_N4BEG[4] ,
    \Tile_X1Y12_N4BEG[3] ,
    \Tile_X1Y12_N4BEG[2] ,
    \Tile_X1Y12_N4BEG[1] ,
    \Tile_X1Y12_N4BEG[0] }),
    .N4END({\Tile_X1Y13_N4BEG[15] ,
    \Tile_X1Y13_N4BEG[14] ,
    \Tile_X1Y13_N4BEG[13] ,
    \Tile_X1Y13_N4BEG[12] ,
    \Tile_X1Y13_N4BEG[11] ,
    \Tile_X1Y13_N4BEG[10] ,
    \Tile_X1Y13_N4BEG[9] ,
    \Tile_X1Y13_N4BEG[8] ,
    \Tile_X1Y13_N4BEG[7] ,
    \Tile_X1Y13_N4BEG[6] ,
    \Tile_X1Y13_N4BEG[5] ,
    \Tile_X1Y13_N4BEG[4] ,
    \Tile_X1Y13_N4BEG[3] ,
    \Tile_X1Y13_N4BEG[2] ,
    \Tile_X1Y13_N4BEG[1] ,
    \Tile_X1Y13_N4BEG[0] }),
    .NN4BEG({\Tile_X1Y12_NN4BEG[15] ,
    \Tile_X1Y12_NN4BEG[14] ,
    \Tile_X1Y12_NN4BEG[13] ,
    \Tile_X1Y12_NN4BEG[12] ,
    \Tile_X1Y12_NN4BEG[11] ,
    \Tile_X1Y12_NN4BEG[10] ,
    \Tile_X1Y12_NN4BEG[9] ,
    \Tile_X1Y12_NN4BEG[8] ,
    \Tile_X1Y12_NN4BEG[7] ,
    \Tile_X1Y12_NN4BEG[6] ,
    \Tile_X1Y12_NN4BEG[5] ,
    \Tile_X1Y12_NN4BEG[4] ,
    \Tile_X1Y12_NN4BEG[3] ,
    \Tile_X1Y12_NN4BEG[2] ,
    \Tile_X1Y12_NN4BEG[1] ,
    \Tile_X1Y12_NN4BEG[0] }),
    .NN4END({\Tile_X1Y13_NN4BEG[15] ,
    \Tile_X1Y13_NN4BEG[14] ,
    \Tile_X1Y13_NN4BEG[13] ,
    \Tile_X1Y13_NN4BEG[12] ,
    \Tile_X1Y13_NN4BEG[11] ,
    \Tile_X1Y13_NN4BEG[10] ,
    \Tile_X1Y13_NN4BEG[9] ,
    \Tile_X1Y13_NN4BEG[8] ,
    \Tile_X1Y13_NN4BEG[7] ,
    \Tile_X1Y13_NN4BEG[6] ,
    \Tile_X1Y13_NN4BEG[5] ,
    \Tile_X1Y13_NN4BEG[4] ,
    \Tile_X1Y13_NN4BEG[3] ,
    \Tile_X1Y13_NN4BEG[2] ,
    \Tile_X1Y13_NN4BEG[1] ,
    \Tile_X1Y13_NN4BEG[0] }),
    .S1BEG({\Tile_X1Y12_S1BEG[3] ,
    \Tile_X1Y12_S1BEG[2] ,
    \Tile_X1Y12_S1BEG[1] ,
    \Tile_X1Y12_S1BEG[0] }),
    .S1END({\Tile_X1Y11_S1BEG[3] ,
    \Tile_X1Y11_S1BEG[2] ,
    \Tile_X1Y11_S1BEG[1] ,
    \Tile_X1Y11_S1BEG[0] }),
    .S2BEG({\Tile_X1Y12_S2BEG[7] ,
    \Tile_X1Y12_S2BEG[6] ,
    \Tile_X1Y12_S2BEG[5] ,
    \Tile_X1Y12_S2BEG[4] ,
    \Tile_X1Y12_S2BEG[3] ,
    \Tile_X1Y12_S2BEG[2] ,
    \Tile_X1Y12_S2BEG[1] ,
    \Tile_X1Y12_S2BEG[0] }),
    .S2BEGb({\Tile_X1Y12_S2BEGb[7] ,
    \Tile_X1Y12_S2BEGb[6] ,
    \Tile_X1Y12_S2BEGb[5] ,
    \Tile_X1Y12_S2BEGb[4] ,
    \Tile_X1Y12_S2BEGb[3] ,
    \Tile_X1Y12_S2BEGb[2] ,
    \Tile_X1Y12_S2BEGb[1] ,
    \Tile_X1Y12_S2BEGb[0] }),
    .S2END({\Tile_X1Y11_S2BEGb[7] ,
    \Tile_X1Y11_S2BEGb[6] ,
    \Tile_X1Y11_S2BEGb[5] ,
    \Tile_X1Y11_S2BEGb[4] ,
    \Tile_X1Y11_S2BEGb[3] ,
    \Tile_X1Y11_S2BEGb[2] ,
    \Tile_X1Y11_S2BEGb[1] ,
    \Tile_X1Y11_S2BEGb[0] }),
    .S2MID({\Tile_X1Y11_S2BEG[7] ,
    \Tile_X1Y11_S2BEG[6] ,
    \Tile_X1Y11_S2BEG[5] ,
    \Tile_X1Y11_S2BEG[4] ,
    \Tile_X1Y11_S2BEG[3] ,
    \Tile_X1Y11_S2BEG[2] ,
    \Tile_X1Y11_S2BEG[1] ,
    \Tile_X1Y11_S2BEG[0] }),
    .S4BEG({\Tile_X1Y12_S4BEG[15] ,
    \Tile_X1Y12_S4BEG[14] ,
    \Tile_X1Y12_S4BEG[13] ,
    \Tile_X1Y12_S4BEG[12] ,
    \Tile_X1Y12_S4BEG[11] ,
    \Tile_X1Y12_S4BEG[10] ,
    \Tile_X1Y12_S4BEG[9] ,
    \Tile_X1Y12_S4BEG[8] ,
    \Tile_X1Y12_S4BEG[7] ,
    \Tile_X1Y12_S4BEG[6] ,
    \Tile_X1Y12_S4BEG[5] ,
    \Tile_X1Y12_S4BEG[4] ,
    \Tile_X1Y12_S4BEG[3] ,
    \Tile_X1Y12_S4BEG[2] ,
    \Tile_X1Y12_S4BEG[1] ,
    \Tile_X1Y12_S4BEG[0] }),
    .S4END({\Tile_X1Y11_S4BEG[15] ,
    \Tile_X1Y11_S4BEG[14] ,
    \Tile_X1Y11_S4BEG[13] ,
    \Tile_X1Y11_S4BEG[12] ,
    \Tile_X1Y11_S4BEG[11] ,
    \Tile_X1Y11_S4BEG[10] ,
    \Tile_X1Y11_S4BEG[9] ,
    \Tile_X1Y11_S4BEG[8] ,
    \Tile_X1Y11_S4BEG[7] ,
    \Tile_X1Y11_S4BEG[6] ,
    \Tile_X1Y11_S4BEG[5] ,
    \Tile_X1Y11_S4BEG[4] ,
    \Tile_X1Y11_S4BEG[3] ,
    \Tile_X1Y11_S4BEG[2] ,
    \Tile_X1Y11_S4BEG[1] ,
    \Tile_X1Y11_S4BEG[0] }),
    .SS4BEG({\Tile_X1Y12_SS4BEG[15] ,
    \Tile_X1Y12_SS4BEG[14] ,
    \Tile_X1Y12_SS4BEG[13] ,
    \Tile_X1Y12_SS4BEG[12] ,
    \Tile_X1Y12_SS4BEG[11] ,
    \Tile_X1Y12_SS4BEG[10] ,
    \Tile_X1Y12_SS4BEG[9] ,
    \Tile_X1Y12_SS4BEG[8] ,
    \Tile_X1Y12_SS4BEG[7] ,
    \Tile_X1Y12_SS4BEG[6] ,
    \Tile_X1Y12_SS4BEG[5] ,
    \Tile_X1Y12_SS4BEG[4] ,
    \Tile_X1Y12_SS4BEG[3] ,
    \Tile_X1Y12_SS4BEG[2] ,
    \Tile_X1Y12_SS4BEG[1] ,
    \Tile_X1Y12_SS4BEG[0] }),
    .SS4END({\Tile_X1Y11_SS4BEG[15] ,
    \Tile_X1Y11_SS4BEG[14] ,
    \Tile_X1Y11_SS4BEG[13] ,
    \Tile_X1Y11_SS4BEG[12] ,
    \Tile_X1Y11_SS4BEG[11] ,
    \Tile_X1Y11_SS4BEG[10] ,
    \Tile_X1Y11_SS4BEG[9] ,
    \Tile_X1Y11_SS4BEG[8] ,
    \Tile_X1Y11_SS4BEG[7] ,
    \Tile_X1Y11_SS4BEG[6] ,
    \Tile_X1Y11_SS4BEG[5] ,
    \Tile_X1Y11_SS4BEG[4] ,
    \Tile_X1Y11_SS4BEG[3] ,
    \Tile_X1Y11_SS4BEG[2] ,
    \Tile_X1Y11_SS4BEG[1] ,
    \Tile_X1Y11_SS4BEG[0] }),
    .W1BEG({\Tile_X1Y12_W1BEG[3] ,
    \Tile_X1Y12_W1BEG[2] ,
    \Tile_X1Y12_W1BEG[1] ,
    \Tile_X1Y12_W1BEG[0] }),
    .W1END({\Tile_X2Y12_W1BEG[3] ,
    \Tile_X2Y12_W1BEG[2] ,
    \Tile_X2Y12_W1BEG[1] ,
    \Tile_X2Y12_W1BEG[0] }),
    .W2BEG({\Tile_X1Y12_W2BEG[7] ,
    \Tile_X1Y12_W2BEG[6] ,
    \Tile_X1Y12_W2BEG[5] ,
    \Tile_X1Y12_W2BEG[4] ,
    \Tile_X1Y12_W2BEG[3] ,
    \Tile_X1Y12_W2BEG[2] ,
    \Tile_X1Y12_W2BEG[1] ,
    \Tile_X1Y12_W2BEG[0] }),
    .W2BEGb({\Tile_X1Y12_W2BEGb[7] ,
    \Tile_X1Y12_W2BEGb[6] ,
    \Tile_X1Y12_W2BEGb[5] ,
    \Tile_X1Y12_W2BEGb[4] ,
    \Tile_X1Y12_W2BEGb[3] ,
    \Tile_X1Y12_W2BEGb[2] ,
    \Tile_X1Y12_W2BEGb[1] ,
    \Tile_X1Y12_W2BEGb[0] }),
    .W2END({\Tile_X2Y12_W2BEGb[7] ,
    \Tile_X2Y12_W2BEGb[6] ,
    \Tile_X2Y12_W2BEGb[5] ,
    \Tile_X2Y12_W2BEGb[4] ,
    \Tile_X2Y12_W2BEGb[3] ,
    \Tile_X2Y12_W2BEGb[2] ,
    \Tile_X2Y12_W2BEGb[1] ,
    \Tile_X2Y12_W2BEGb[0] }),
    .W2MID({\Tile_X2Y12_W2BEG[7] ,
    \Tile_X2Y12_W2BEG[6] ,
    \Tile_X2Y12_W2BEG[5] ,
    \Tile_X2Y12_W2BEG[4] ,
    \Tile_X2Y12_W2BEG[3] ,
    \Tile_X2Y12_W2BEG[2] ,
    \Tile_X2Y12_W2BEG[1] ,
    \Tile_X2Y12_W2BEG[0] }),
    .W6BEG({\Tile_X1Y12_W6BEG[11] ,
    \Tile_X1Y12_W6BEG[10] ,
    \Tile_X1Y12_W6BEG[9] ,
    \Tile_X1Y12_W6BEG[8] ,
    \Tile_X1Y12_W6BEG[7] ,
    \Tile_X1Y12_W6BEG[6] ,
    \Tile_X1Y12_W6BEG[5] ,
    \Tile_X1Y12_W6BEG[4] ,
    \Tile_X1Y12_W6BEG[3] ,
    \Tile_X1Y12_W6BEG[2] ,
    \Tile_X1Y12_W6BEG[1] ,
    \Tile_X1Y12_W6BEG[0] }),
    .W6END({\Tile_X2Y12_W6BEG[11] ,
    \Tile_X2Y12_W6BEG[10] ,
    \Tile_X2Y12_W6BEG[9] ,
    \Tile_X2Y12_W6BEG[8] ,
    \Tile_X2Y12_W6BEG[7] ,
    \Tile_X2Y12_W6BEG[6] ,
    \Tile_X2Y12_W6BEG[5] ,
    \Tile_X2Y12_W6BEG[4] ,
    \Tile_X2Y12_W6BEG[3] ,
    \Tile_X2Y12_W6BEG[2] ,
    \Tile_X2Y12_W6BEG[1] ,
    \Tile_X2Y12_W6BEG[0] }),
    .WW4BEG({\Tile_X1Y12_WW4BEG[15] ,
    \Tile_X1Y12_WW4BEG[14] ,
    \Tile_X1Y12_WW4BEG[13] ,
    \Tile_X1Y12_WW4BEG[12] ,
    \Tile_X1Y12_WW4BEG[11] ,
    \Tile_X1Y12_WW4BEG[10] ,
    \Tile_X1Y12_WW4BEG[9] ,
    \Tile_X1Y12_WW4BEG[8] ,
    \Tile_X1Y12_WW4BEG[7] ,
    \Tile_X1Y12_WW4BEG[6] ,
    \Tile_X1Y12_WW4BEG[5] ,
    \Tile_X1Y12_WW4BEG[4] ,
    \Tile_X1Y12_WW4BEG[3] ,
    \Tile_X1Y12_WW4BEG[2] ,
    \Tile_X1Y12_WW4BEG[1] ,
    \Tile_X1Y12_WW4BEG[0] }),
    .WW4END({\Tile_X2Y12_WW4BEG[15] ,
    \Tile_X2Y12_WW4BEG[14] ,
    \Tile_X2Y12_WW4BEG[13] ,
    \Tile_X2Y12_WW4BEG[12] ,
    \Tile_X2Y12_WW4BEG[11] ,
    \Tile_X2Y12_WW4BEG[10] ,
    \Tile_X2Y12_WW4BEG[9] ,
    \Tile_X2Y12_WW4BEG[8] ,
    \Tile_X2Y12_WW4BEG[7] ,
    \Tile_X2Y12_WW4BEG[6] ,
    \Tile_X2Y12_WW4BEG[5] ,
    \Tile_X2Y12_WW4BEG[4] ,
    \Tile_X2Y12_WW4BEG[3] ,
    \Tile_X2Y12_WW4BEG[2] ,
    \Tile_X2Y12_WW4BEG[1] ,
    \Tile_X2Y12_WW4BEG[0] }));
 LUT4AB Tile_X1Y13_LUT4AB (.Ci(Tile_X1Y14_Co),
    .Co(Tile_X1Y13_Co),
    .UserCLK(Tile_X1Y14_UserCLKo),
    .UserCLKo(Tile_X1Y13_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X1Y13_E1BEG[3] ,
    \Tile_X1Y13_E1BEG[2] ,
    \Tile_X1Y13_E1BEG[1] ,
    \Tile_X1Y13_E1BEG[0] }),
    .E1END({\Tile_X0Y13_E1BEG[3] ,
    \Tile_X0Y13_E1BEG[2] ,
    \Tile_X0Y13_E1BEG[1] ,
    \Tile_X0Y13_E1BEG[0] }),
    .E2BEG({\Tile_X1Y13_E2BEG[7] ,
    \Tile_X1Y13_E2BEG[6] ,
    \Tile_X1Y13_E2BEG[5] ,
    \Tile_X1Y13_E2BEG[4] ,
    \Tile_X1Y13_E2BEG[3] ,
    \Tile_X1Y13_E2BEG[2] ,
    \Tile_X1Y13_E2BEG[1] ,
    \Tile_X1Y13_E2BEG[0] }),
    .E2BEGb({\Tile_X1Y13_E2BEGb[7] ,
    \Tile_X1Y13_E2BEGb[6] ,
    \Tile_X1Y13_E2BEGb[5] ,
    \Tile_X1Y13_E2BEGb[4] ,
    \Tile_X1Y13_E2BEGb[3] ,
    \Tile_X1Y13_E2BEGb[2] ,
    \Tile_X1Y13_E2BEGb[1] ,
    \Tile_X1Y13_E2BEGb[0] }),
    .E2END({\Tile_X0Y13_E2BEGb[7] ,
    \Tile_X0Y13_E2BEGb[6] ,
    \Tile_X0Y13_E2BEGb[5] ,
    \Tile_X0Y13_E2BEGb[4] ,
    \Tile_X0Y13_E2BEGb[3] ,
    \Tile_X0Y13_E2BEGb[2] ,
    \Tile_X0Y13_E2BEGb[1] ,
    \Tile_X0Y13_E2BEGb[0] }),
    .E2MID({\Tile_X0Y13_E2BEG[7] ,
    \Tile_X0Y13_E2BEG[6] ,
    \Tile_X0Y13_E2BEG[5] ,
    \Tile_X0Y13_E2BEG[4] ,
    \Tile_X0Y13_E2BEG[3] ,
    \Tile_X0Y13_E2BEG[2] ,
    \Tile_X0Y13_E2BEG[1] ,
    \Tile_X0Y13_E2BEG[0] }),
    .E6BEG({\Tile_X1Y13_E6BEG[11] ,
    \Tile_X1Y13_E6BEG[10] ,
    \Tile_X1Y13_E6BEG[9] ,
    \Tile_X1Y13_E6BEG[8] ,
    \Tile_X1Y13_E6BEG[7] ,
    \Tile_X1Y13_E6BEG[6] ,
    \Tile_X1Y13_E6BEG[5] ,
    \Tile_X1Y13_E6BEG[4] ,
    \Tile_X1Y13_E6BEG[3] ,
    \Tile_X1Y13_E6BEG[2] ,
    \Tile_X1Y13_E6BEG[1] ,
    \Tile_X1Y13_E6BEG[0] }),
    .E6END({\Tile_X0Y13_E6BEG[11] ,
    \Tile_X0Y13_E6BEG[10] ,
    \Tile_X0Y13_E6BEG[9] ,
    \Tile_X0Y13_E6BEG[8] ,
    \Tile_X0Y13_E6BEG[7] ,
    \Tile_X0Y13_E6BEG[6] ,
    \Tile_X0Y13_E6BEG[5] ,
    \Tile_X0Y13_E6BEG[4] ,
    \Tile_X0Y13_E6BEG[3] ,
    \Tile_X0Y13_E6BEG[2] ,
    \Tile_X0Y13_E6BEG[1] ,
    \Tile_X0Y13_E6BEG[0] }),
    .EE4BEG({\Tile_X1Y13_EE4BEG[15] ,
    \Tile_X1Y13_EE4BEG[14] ,
    \Tile_X1Y13_EE4BEG[13] ,
    \Tile_X1Y13_EE4BEG[12] ,
    \Tile_X1Y13_EE4BEG[11] ,
    \Tile_X1Y13_EE4BEG[10] ,
    \Tile_X1Y13_EE4BEG[9] ,
    \Tile_X1Y13_EE4BEG[8] ,
    \Tile_X1Y13_EE4BEG[7] ,
    \Tile_X1Y13_EE4BEG[6] ,
    \Tile_X1Y13_EE4BEG[5] ,
    \Tile_X1Y13_EE4BEG[4] ,
    \Tile_X1Y13_EE4BEG[3] ,
    \Tile_X1Y13_EE4BEG[2] ,
    \Tile_X1Y13_EE4BEG[1] ,
    \Tile_X1Y13_EE4BEG[0] }),
    .EE4END({\Tile_X0Y13_EE4BEG[15] ,
    \Tile_X0Y13_EE4BEG[14] ,
    \Tile_X0Y13_EE4BEG[13] ,
    \Tile_X0Y13_EE4BEG[12] ,
    \Tile_X0Y13_EE4BEG[11] ,
    \Tile_X0Y13_EE4BEG[10] ,
    \Tile_X0Y13_EE4BEG[9] ,
    \Tile_X0Y13_EE4BEG[8] ,
    \Tile_X0Y13_EE4BEG[7] ,
    \Tile_X0Y13_EE4BEG[6] ,
    \Tile_X0Y13_EE4BEG[5] ,
    \Tile_X0Y13_EE4BEG[4] ,
    \Tile_X0Y13_EE4BEG[3] ,
    \Tile_X0Y13_EE4BEG[2] ,
    \Tile_X0Y13_EE4BEG[1] ,
    \Tile_X0Y13_EE4BEG[0] }),
    .FrameData({\Tile_X0Y13_FrameData_O[31] ,
    \Tile_X0Y13_FrameData_O[30] ,
    \Tile_X0Y13_FrameData_O[29] ,
    \Tile_X0Y13_FrameData_O[28] ,
    \Tile_X0Y13_FrameData_O[27] ,
    \Tile_X0Y13_FrameData_O[26] ,
    \Tile_X0Y13_FrameData_O[25] ,
    \Tile_X0Y13_FrameData_O[24] ,
    \Tile_X0Y13_FrameData_O[23] ,
    \Tile_X0Y13_FrameData_O[22] ,
    \Tile_X0Y13_FrameData_O[21] ,
    \Tile_X0Y13_FrameData_O[20] ,
    \Tile_X0Y13_FrameData_O[19] ,
    \Tile_X0Y13_FrameData_O[18] ,
    \Tile_X0Y13_FrameData_O[17] ,
    \Tile_X0Y13_FrameData_O[16] ,
    \Tile_X0Y13_FrameData_O[15] ,
    \Tile_X0Y13_FrameData_O[14] ,
    \Tile_X0Y13_FrameData_O[13] ,
    \Tile_X0Y13_FrameData_O[12] ,
    \Tile_X0Y13_FrameData_O[11] ,
    \Tile_X0Y13_FrameData_O[10] ,
    \Tile_X0Y13_FrameData_O[9] ,
    \Tile_X0Y13_FrameData_O[8] ,
    \Tile_X0Y13_FrameData_O[7] ,
    \Tile_X0Y13_FrameData_O[6] ,
    \Tile_X0Y13_FrameData_O[5] ,
    \Tile_X0Y13_FrameData_O[4] ,
    \Tile_X0Y13_FrameData_O[3] ,
    \Tile_X0Y13_FrameData_O[2] ,
    \Tile_X0Y13_FrameData_O[1] ,
    \Tile_X0Y13_FrameData_O[0] }),
    .FrameData_O({\Tile_X1Y13_FrameData_O[31] ,
    \Tile_X1Y13_FrameData_O[30] ,
    \Tile_X1Y13_FrameData_O[29] ,
    \Tile_X1Y13_FrameData_O[28] ,
    \Tile_X1Y13_FrameData_O[27] ,
    \Tile_X1Y13_FrameData_O[26] ,
    \Tile_X1Y13_FrameData_O[25] ,
    \Tile_X1Y13_FrameData_O[24] ,
    \Tile_X1Y13_FrameData_O[23] ,
    \Tile_X1Y13_FrameData_O[22] ,
    \Tile_X1Y13_FrameData_O[21] ,
    \Tile_X1Y13_FrameData_O[20] ,
    \Tile_X1Y13_FrameData_O[19] ,
    \Tile_X1Y13_FrameData_O[18] ,
    \Tile_X1Y13_FrameData_O[17] ,
    \Tile_X1Y13_FrameData_O[16] ,
    \Tile_X1Y13_FrameData_O[15] ,
    \Tile_X1Y13_FrameData_O[14] ,
    \Tile_X1Y13_FrameData_O[13] ,
    \Tile_X1Y13_FrameData_O[12] ,
    \Tile_X1Y13_FrameData_O[11] ,
    \Tile_X1Y13_FrameData_O[10] ,
    \Tile_X1Y13_FrameData_O[9] ,
    \Tile_X1Y13_FrameData_O[8] ,
    \Tile_X1Y13_FrameData_O[7] ,
    \Tile_X1Y13_FrameData_O[6] ,
    \Tile_X1Y13_FrameData_O[5] ,
    \Tile_X1Y13_FrameData_O[4] ,
    \Tile_X1Y13_FrameData_O[3] ,
    \Tile_X1Y13_FrameData_O[2] ,
    \Tile_X1Y13_FrameData_O[1] ,
    \Tile_X1Y13_FrameData_O[0] }),
    .FrameStrobe({\Tile_X1Y14_FrameStrobe_O[19] ,
    \Tile_X1Y14_FrameStrobe_O[18] ,
    \Tile_X1Y14_FrameStrobe_O[17] ,
    \Tile_X1Y14_FrameStrobe_O[16] ,
    \Tile_X1Y14_FrameStrobe_O[15] ,
    \Tile_X1Y14_FrameStrobe_O[14] ,
    \Tile_X1Y14_FrameStrobe_O[13] ,
    \Tile_X1Y14_FrameStrobe_O[12] ,
    \Tile_X1Y14_FrameStrobe_O[11] ,
    \Tile_X1Y14_FrameStrobe_O[10] ,
    \Tile_X1Y14_FrameStrobe_O[9] ,
    \Tile_X1Y14_FrameStrobe_O[8] ,
    \Tile_X1Y14_FrameStrobe_O[7] ,
    \Tile_X1Y14_FrameStrobe_O[6] ,
    \Tile_X1Y14_FrameStrobe_O[5] ,
    \Tile_X1Y14_FrameStrobe_O[4] ,
    \Tile_X1Y14_FrameStrobe_O[3] ,
    \Tile_X1Y14_FrameStrobe_O[2] ,
    \Tile_X1Y14_FrameStrobe_O[1] ,
    \Tile_X1Y14_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X1Y13_FrameStrobe_O[19] ,
    \Tile_X1Y13_FrameStrobe_O[18] ,
    \Tile_X1Y13_FrameStrobe_O[17] ,
    \Tile_X1Y13_FrameStrobe_O[16] ,
    \Tile_X1Y13_FrameStrobe_O[15] ,
    \Tile_X1Y13_FrameStrobe_O[14] ,
    \Tile_X1Y13_FrameStrobe_O[13] ,
    \Tile_X1Y13_FrameStrobe_O[12] ,
    \Tile_X1Y13_FrameStrobe_O[11] ,
    \Tile_X1Y13_FrameStrobe_O[10] ,
    \Tile_X1Y13_FrameStrobe_O[9] ,
    \Tile_X1Y13_FrameStrobe_O[8] ,
    \Tile_X1Y13_FrameStrobe_O[7] ,
    \Tile_X1Y13_FrameStrobe_O[6] ,
    \Tile_X1Y13_FrameStrobe_O[5] ,
    \Tile_X1Y13_FrameStrobe_O[4] ,
    \Tile_X1Y13_FrameStrobe_O[3] ,
    \Tile_X1Y13_FrameStrobe_O[2] ,
    \Tile_X1Y13_FrameStrobe_O[1] ,
    \Tile_X1Y13_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X1Y13_N1BEG[3] ,
    \Tile_X1Y13_N1BEG[2] ,
    \Tile_X1Y13_N1BEG[1] ,
    \Tile_X1Y13_N1BEG[0] }),
    .N1END({\Tile_X1Y14_N1BEG[3] ,
    \Tile_X1Y14_N1BEG[2] ,
    \Tile_X1Y14_N1BEG[1] ,
    \Tile_X1Y14_N1BEG[0] }),
    .N2BEG({\Tile_X1Y13_N2BEG[7] ,
    \Tile_X1Y13_N2BEG[6] ,
    \Tile_X1Y13_N2BEG[5] ,
    \Tile_X1Y13_N2BEG[4] ,
    \Tile_X1Y13_N2BEG[3] ,
    \Tile_X1Y13_N2BEG[2] ,
    \Tile_X1Y13_N2BEG[1] ,
    \Tile_X1Y13_N2BEG[0] }),
    .N2BEGb({\Tile_X1Y13_N2BEGb[7] ,
    \Tile_X1Y13_N2BEGb[6] ,
    \Tile_X1Y13_N2BEGb[5] ,
    \Tile_X1Y13_N2BEGb[4] ,
    \Tile_X1Y13_N2BEGb[3] ,
    \Tile_X1Y13_N2BEGb[2] ,
    \Tile_X1Y13_N2BEGb[1] ,
    \Tile_X1Y13_N2BEGb[0] }),
    .N2END({\Tile_X1Y14_N2BEGb[7] ,
    \Tile_X1Y14_N2BEGb[6] ,
    \Tile_X1Y14_N2BEGb[5] ,
    \Tile_X1Y14_N2BEGb[4] ,
    \Tile_X1Y14_N2BEGb[3] ,
    \Tile_X1Y14_N2BEGb[2] ,
    \Tile_X1Y14_N2BEGb[1] ,
    \Tile_X1Y14_N2BEGb[0] }),
    .N2MID({\Tile_X1Y14_N2BEG[7] ,
    \Tile_X1Y14_N2BEG[6] ,
    \Tile_X1Y14_N2BEG[5] ,
    \Tile_X1Y14_N2BEG[4] ,
    \Tile_X1Y14_N2BEG[3] ,
    \Tile_X1Y14_N2BEG[2] ,
    \Tile_X1Y14_N2BEG[1] ,
    \Tile_X1Y14_N2BEG[0] }),
    .N4BEG({\Tile_X1Y13_N4BEG[15] ,
    \Tile_X1Y13_N4BEG[14] ,
    \Tile_X1Y13_N4BEG[13] ,
    \Tile_X1Y13_N4BEG[12] ,
    \Tile_X1Y13_N4BEG[11] ,
    \Tile_X1Y13_N4BEG[10] ,
    \Tile_X1Y13_N4BEG[9] ,
    \Tile_X1Y13_N4BEG[8] ,
    \Tile_X1Y13_N4BEG[7] ,
    \Tile_X1Y13_N4BEG[6] ,
    \Tile_X1Y13_N4BEG[5] ,
    \Tile_X1Y13_N4BEG[4] ,
    \Tile_X1Y13_N4BEG[3] ,
    \Tile_X1Y13_N4BEG[2] ,
    \Tile_X1Y13_N4BEG[1] ,
    \Tile_X1Y13_N4BEG[0] }),
    .N4END({\Tile_X1Y14_N4BEG[15] ,
    \Tile_X1Y14_N4BEG[14] ,
    \Tile_X1Y14_N4BEG[13] ,
    \Tile_X1Y14_N4BEG[12] ,
    \Tile_X1Y14_N4BEG[11] ,
    \Tile_X1Y14_N4BEG[10] ,
    \Tile_X1Y14_N4BEG[9] ,
    \Tile_X1Y14_N4BEG[8] ,
    \Tile_X1Y14_N4BEG[7] ,
    \Tile_X1Y14_N4BEG[6] ,
    \Tile_X1Y14_N4BEG[5] ,
    \Tile_X1Y14_N4BEG[4] ,
    \Tile_X1Y14_N4BEG[3] ,
    \Tile_X1Y14_N4BEG[2] ,
    \Tile_X1Y14_N4BEG[1] ,
    \Tile_X1Y14_N4BEG[0] }),
    .NN4BEG({\Tile_X1Y13_NN4BEG[15] ,
    \Tile_X1Y13_NN4BEG[14] ,
    \Tile_X1Y13_NN4BEG[13] ,
    \Tile_X1Y13_NN4BEG[12] ,
    \Tile_X1Y13_NN4BEG[11] ,
    \Tile_X1Y13_NN4BEG[10] ,
    \Tile_X1Y13_NN4BEG[9] ,
    \Tile_X1Y13_NN4BEG[8] ,
    \Tile_X1Y13_NN4BEG[7] ,
    \Tile_X1Y13_NN4BEG[6] ,
    \Tile_X1Y13_NN4BEG[5] ,
    \Tile_X1Y13_NN4BEG[4] ,
    \Tile_X1Y13_NN4BEG[3] ,
    \Tile_X1Y13_NN4BEG[2] ,
    \Tile_X1Y13_NN4BEG[1] ,
    \Tile_X1Y13_NN4BEG[0] }),
    .NN4END({\Tile_X1Y14_NN4BEG[15] ,
    \Tile_X1Y14_NN4BEG[14] ,
    \Tile_X1Y14_NN4BEG[13] ,
    \Tile_X1Y14_NN4BEG[12] ,
    \Tile_X1Y14_NN4BEG[11] ,
    \Tile_X1Y14_NN4BEG[10] ,
    \Tile_X1Y14_NN4BEG[9] ,
    \Tile_X1Y14_NN4BEG[8] ,
    \Tile_X1Y14_NN4BEG[7] ,
    \Tile_X1Y14_NN4BEG[6] ,
    \Tile_X1Y14_NN4BEG[5] ,
    \Tile_X1Y14_NN4BEG[4] ,
    \Tile_X1Y14_NN4BEG[3] ,
    \Tile_X1Y14_NN4BEG[2] ,
    \Tile_X1Y14_NN4BEG[1] ,
    \Tile_X1Y14_NN4BEG[0] }),
    .S1BEG({\Tile_X1Y13_S1BEG[3] ,
    \Tile_X1Y13_S1BEG[2] ,
    \Tile_X1Y13_S1BEG[1] ,
    \Tile_X1Y13_S1BEG[0] }),
    .S1END({\Tile_X1Y12_S1BEG[3] ,
    \Tile_X1Y12_S1BEG[2] ,
    \Tile_X1Y12_S1BEG[1] ,
    \Tile_X1Y12_S1BEG[0] }),
    .S2BEG({\Tile_X1Y13_S2BEG[7] ,
    \Tile_X1Y13_S2BEG[6] ,
    \Tile_X1Y13_S2BEG[5] ,
    \Tile_X1Y13_S2BEG[4] ,
    \Tile_X1Y13_S2BEG[3] ,
    \Tile_X1Y13_S2BEG[2] ,
    \Tile_X1Y13_S2BEG[1] ,
    \Tile_X1Y13_S2BEG[0] }),
    .S2BEGb({\Tile_X1Y13_S2BEGb[7] ,
    \Tile_X1Y13_S2BEGb[6] ,
    \Tile_X1Y13_S2BEGb[5] ,
    \Tile_X1Y13_S2BEGb[4] ,
    \Tile_X1Y13_S2BEGb[3] ,
    \Tile_X1Y13_S2BEGb[2] ,
    \Tile_X1Y13_S2BEGb[1] ,
    \Tile_X1Y13_S2BEGb[0] }),
    .S2END({\Tile_X1Y12_S2BEGb[7] ,
    \Tile_X1Y12_S2BEGb[6] ,
    \Tile_X1Y12_S2BEGb[5] ,
    \Tile_X1Y12_S2BEGb[4] ,
    \Tile_X1Y12_S2BEGb[3] ,
    \Tile_X1Y12_S2BEGb[2] ,
    \Tile_X1Y12_S2BEGb[1] ,
    \Tile_X1Y12_S2BEGb[0] }),
    .S2MID({\Tile_X1Y12_S2BEG[7] ,
    \Tile_X1Y12_S2BEG[6] ,
    \Tile_X1Y12_S2BEG[5] ,
    \Tile_X1Y12_S2BEG[4] ,
    \Tile_X1Y12_S2BEG[3] ,
    \Tile_X1Y12_S2BEG[2] ,
    \Tile_X1Y12_S2BEG[1] ,
    \Tile_X1Y12_S2BEG[0] }),
    .S4BEG({\Tile_X1Y13_S4BEG[15] ,
    \Tile_X1Y13_S4BEG[14] ,
    \Tile_X1Y13_S4BEG[13] ,
    \Tile_X1Y13_S4BEG[12] ,
    \Tile_X1Y13_S4BEG[11] ,
    \Tile_X1Y13_S4BEG[10] ,
    \Tile_X1Y13_S4BEG[9] ,
    \Tile_X1Y13_S4BEG[8] ,
    \Tile_X1Y13_S4BEG[7] ,
    \Tile_X1Y13_S4BEG[6] ,
    \Tile_X1Y13_S4BEG[5] ,
    \Tile_X1Y13_S4BEG[4] ,
    \Tile_X1Y13_S4BEG[3] ,
    \Tile_X1Y13_S4BEG[2] ,
    \Tile_X1Y13_S4BEG[1] ,
    \Tile_X1Y13_S4BEG[0] }),
    .S4END({\Tile_X1Y12_S4BEG[15] ,
    \Tile_X1Y12_S4BEG[14] ,
    \Tile_X1Y12_S4BEG[13] ,
    \Tile_X1Y12_S4BEG[12] ,
    \Tile_X1Y12_S4BEG[11] ,
    \Tile_X1Y12_S4BEG[10] ,
    \Tile_X1Y12_S4BEG[9] ,
    \Tile_X1Y12_S4BEG[8] ,
    \Tile_X1Y12_S4BEG[7] ,
    \Tile_X1Y12_S4BEG[6] ,
    \Tile_X1Y12_S4BEG[5] ,
    \Tile_X1Y12_S4BEG[4] ,
    \Tile_X1Y12_S4BEG[3] ,
    \Tile_X1Y12_S4BEG[2] ,
    \Tile_X1Y12_S4BEG[1] ,
    \Tile_X1Y12_S4BEG[0] }),
    .SS4BEG({\Tile_X1Y13_SS4BEG[15] ,
    \Tile_X1Y13_SS4BEG[14] ,
    \Tile_X1Y13_SS4BEG[13] ,
    \Tile_X1Y13_SS4BEG[12] ,
    \Tile_X1Y13_SS4BEG[11] ,
    \Tile_X1Y13_SS4BEG[10] ,
    \Tile_X1Y13_SS4BEG[9] ,
    \Tile_X1Y13_SS4BEG[8] ,
    \Tile_X1Y13_SS4BEG[7] ,
    \Tile_X1Y13_SS4BEG[6] ,
    \Tile_X1Y13_SS4BEG[5] ,
    \Tile_X1Y13_SS4BEG[4] ,
    \Tile_X1Y13_SS4BEG[3] ,
    \Tile_X1Y13_SS4BEG[2] ,
    \Tile_X1Y13_SS4BEG[1] ,
    \Tile_X1Y13_SS4BEG[0] }),
    .SS4END({\Tile_X1Y12_SS4BEG[15] ,
    \Tile_X1Y12_SS4BEG[14] ,
    \Tile_X1Y12_SS4BEG[13] ,
    \Tile_X1Y12_SS4BEG[12] ,
    \Tile_X1Y12_SS4BEG[11] ,
    \Tile_X1Y12_SS4BEG[10] ,
    \Tile_X1Y12_SS4BEG[9] ,
    \Tile_X1Y12_SS4BEG[8] ,
    \Tile_X1Y12_SS4BEG[7] ,
    \Tile_X1Y12_SS4BEG[6] ,
    \Tile_X1Y12_SS4BEG[5] ,
    \Tile_X1Y12_SS4BEG[4] ,
    \Tile_X1Y12_SS4BEG[3] ,
    \Tile_X1Y12_SS4BEG[2] ,
    \Tile_X1Y12_SS4BEG[1] ,
    \Tile_X1Y12_SS4BEG[0] }),
    .W1BEG({\Tile_X1Y13_W1BEG[3] ,
    \Tile_X1Y13_W1BEG[2] ,
    \Tile_X1Y13_W1BEG[1] ,
    \Tile_X1Y13_W1BEG[0] }),
    .W1END({\Tile_X2Y13_W1BEG[3] ,
    \Tile_X2Y13_W1BEG[2] ,
    \Tile_X2Y13_W1BEG[1] ,
    \Tile_X2Y13_W1BEG[0] }),
    .W2BEG({\Tile_X1Y13_W2BEG[7] ,
    \Tile_X1Y13_W2BEG[6] ,
    \Tile_X1Y13_W2BEG[5] ,
    \Tile_X1Y13_W2BEG[4] ,
    \Tile_X1Y13_W2BEG[3] ,
    \Tile_X1Y13_W2BEG[2] ,
    \Tile_X1Y13_W2BEG[1] ,
    \Tile_X1Y13_W2BEG[0] }),
    .W2BEGb({\Tile_X1Y13_W2BEGb[7] ,
    \Tile_X1Y13_W2BEGb[6] ,
    \Tile_X1Y13_W2BEGb[5] ,
    \Tile_X1Y13_W2BEGb[4] ,
    \Tile_X1Y13_W2BEGb[3] ,
    \Tile_X1Y13_W2BEGb[2] ,
    \Tile_X1Y13_W2BEGb[1] ,
    \Tile_X1Y13_W2BEGb[0] }),
    .W2END({\Tile_X2Y13_W2BEGb[7] ,
    \Tile_X2Y13_W2BEGb[6] ,
    \Tile_X2Y13_W2BEGb[5] ,
    \Tile_X2Y13_W2BEGb[4] ,
    \Tile_X2Y13_W2BEGb[3] ,
    \Tile_X2Y13_W2BEGb[2] ,
    \Tile_X2Y13_W2BEGb[1] ,
    \Tile_X2Y13_W2BEGb[0] }),
    .W2MID({\Tile_X2Y13_W2BEG[7] ,
    \Tile_X2Y13_W2BEG[6] ,
    \Tile_X2Y13_W2BEG[5] ,
    \Tile_X2Y13_W2BEG[4] ,
    \Tile_X2Y13_W2BEG[3] ,
    \Tile_X2Y13_W2BEG[2] ,
    \Tile_X2Y13_W2BEG[1] ,
    \Tile_X2Y13_W2BEG[0] }),
    .W6BEG({\Tile_X1Y13_W6BEG[11] ,
    \Tile_X1Y13_W6BEG[10] ,
    \Tile_X1Y13_W6BEG[9] ,
    \Tile_X1Y13_W6BEG[8] ,
    \Tile_X1Y13_W6BEG[7] ,
    \Tile_X1Y13_W6BEG[6] ,
    \Tile_X1Y13_W6BEG[5] ,
    \Tile_X1Y13_W6BEG[4] ,
    \Tile_X1Y13_W6BEG[3] ,
    \Tile_X1Y13_W6BEG[2] ,
    \Tile_X1Y13_W6BEG[1] ,
    \Tile_X1Y13_W6BEG[0] }),
    .W6END({\Tile_X2Y13_W6BEG[11] ,
    \Tile_X2Y13_W6BEG[10] ,
    \Tile_X2Y13_W6BEG[9] ,
    \Tile_X2Y13_W6BEG[8] ,
    \Tile_X2Y13_W6BEG[7] ,
    \Tile_X2Y13_W6BEG[6] ,
    \Tile_X2Y13_W6BEG[5] ,
    \Tile_X2Y13_W6BEG[4] ,
    \Tile_X2Y13_W6BEG[3] ,
    \Tile_X2Y13_W6BEG[2] ,
    \Tile_X2Y13_W6BEG[1] ,
    \Tile_X2Y13_W6BEG[0] }),
    .WW4BEG({\Tile_X1Y13_WW4BEG[15] ,
    \Tile_X1Y13_WW4BEG[14] ,
    \Tile_X1Y13_WW4BEG[13] ,
    \Tile_X1Y13_WW4BEG[12] ,
    \Tile_X1Y13_WW4BEG[11] ,
    \Tile_X1Y13_WW4BEG[10] ,
    \Tile_X1Y13_WW4BEG[9] ,
    \Tile_X1Y13_WW4BEG[8] ,
    \Tile_X1Y13_WW4BEG[7] ,
    \Tile_X1Y13_WW4BEG[6] ,
    \Tile_X1Y13_WW4BEG[5] ,
    \Tile_X1Y13_WW4BEG[4] ,
    \Tile_X1Y13_WW4BEG[3] ,
    \Tile_X1Y13_WW4BEG[2] ,
    \Tile_X1Y13_WW4BEG[1] ,
    \Tile_X1Y13_WW4BEG[0] }),
    .WW4END({\Tile_X2Y13_WW4BEG[15] ,
    \Tile_X2Y13_WW4BEG[14] ,
    \Tile_X2Y13_WW4BEG[13] ,
    \Tile_X2Y13_WW4BEG[12] ,
    \Tile_X2Y13_WW4BEG[11] ,
    \Tile_X2Y13_WW4BEG[10] ,
    \Tile_X2Y13_WW4BEG[9] ,
    \Tile_X2Y13_WW4BEG[8] ,
    \Tile_X2Y13_WW4BEG[7] ,
    \Tile_X2Y13_WW4BEG[6] ,
    \Tile_X2Y13_WW4BEG[5] ,
    \Tile_X2Y13_WW4BEG[4] ,
    \Tile_X2Y13_WW4BEG[3] ,
    \Tile_X2Y13_WW4BEG[2] ,
    \Tile_X2Y13_WW4BEG[1] ,
    \Tile_X2Y13_WW4BEG[0] }));
 LUT4AB Tile_X1Y14_LUT4AB (.Ci(Tile_X1Y15_Co),
    .Co(Tile_X1Y14_Co),
    .UserCLK(Tile_X1Y15_UserCLKo),
    .UserCLKo(Tile_X1Y14_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X1Y14_E1BEG[3] ,
    \Tile_X1Y14_E1BEG[2] ,
    \Tile_X1Y14_E1BEG[1] ,
    \Tile_X1Y14_E1BEG[0] }),
    .E1END({\Tile_X0Y14_E1BEG[3] ,
    \Tile_X0Y14_E1BEG[2] ,
    \Tile_X0Y14_E1BEG[1] ,
    \Tile_X0Y14_E1BEG[0] }),
    .E2BEG({\Tile_X1Y14_E2BEG[7] ,
    \Tile_X1Y14_E2BEG[6] ,
    \Tile_X1Y14_E2BEG[5] ,
    \Tile_X1Y14_E2BEG[4] ,
    \Tile_X1Y14_E2BEG[3] ,
    \Tile_X1Y14_E2BEG[2] ,
    \Tile_X1Y14_E2BEG[1] ,
    \Tile_X1Y14_E2BEG[0] }),
    .E2BEGb({\Tile_X1Y14_E2BEGb[7] ,
    \Tile_X1Y14_E2BEGb[6] ,
    \Tile_X1Y14_E2BEGb[5] ,
    \Tile_X1Y14_E2BEGb[4] ,
    \Tile_X1Y14_E2BEGb[3] ,
    \Tile_X1Y14_E2BEGb[2] ,
    \Tile_X1Y14_E2BEGb[1] ,
    \Tile_X1Y14_E2BEGb[0] }),
    .E2END({\Tile_X0Y14_E2BEGb[7] ,
    \Tile_X0Y14_E2BEGb[6] ,
    \Tile_X0Y14_E2BEGb[5] ,
    \Tile_X0Y14_E2BEGb[4] ,
    \Tile_X0Y14_E2BEGb[3] ,
    \Tile_X0Y14_E2BEGb[2] ,
    \Tile_X0Y14_E2BEGb[1] ,
    \Tile_X0Y14_E2BEGb[0] }),
    .E2MID({\Tile_X0Y14_E2BEG[7] ,
    \Tile_X0Y14_E2BEG[6] ,
    \Tile_X0Y14_E2BEG[5] ,
    \Tile_X0Y14_E2BEG[4] ,
    \Tile_X0Y14_E2BEG[3] ,
    \Tile_X0Y14_E2BEG[2] ,
    \Tile_X0Y14_E2BEG[1] ,
    \Tile_X0Y14_E2BEG[0] }),
    .E6BEG({\Tile_X1Y14_E6BEG[11] ,
    \Tile_X1Y14_E6BEG[10] ,
    \Tile_X1Y14_E6BEG[9] ,
    \Tile_X1Y14_E6BEG[8] ,
    \Tile_X1Y14_E6BEG[7] ,
    \Tile_X1Y14_E6BEG[6] ,
    \Tile_X1Y14_E6BEG[5] ,
    \Tile_X1Y14_E6BEG[4] ,
    \Tile_X1Y14_E6BEG[3] ,
    \Tile_X1Y14_E6BEG[2] ,
    \Tile_X1Y14_E6BEG[1] ,
    \Tile_X1Y14_E6BEG[0] }),
    .E6END({\Tile_X0Y14_E6BEG[11] ,
    \Tile_X0Y14_E6BEG[10] ,
    \Tile_X0Y14_E6BEG[9] ,
    \Tile_X0Y14_E6BEG[8] ,
    \Tile_X0Y14_E6BEG[7] ,
    \Tile_X0Y14_E6BEG[6] ,
    \Tile_X0Y14_E6BEG[5] ,
    \Tile_X0Y14_E6BEG[4] ,
    \Tile_X0Y14_E6BEG[3] ,
    \Tile_X0Y14_E6BEG[2] ,
    \Tile_X0Y14_E6BEG[1] ,
    \Tile_X0Y14_E6BEG[0] }),
    .EE4BEG({\Tile_X1Y14_EE4BEG[15] ,
    \Tile_X1Y14_EE4BEG[14] ,
    \Tile_X1Y14_EE4BEG[13] ,
    \Tile_X1Y14_EE4BEG[12] ,
    \Tile_X1Y14_EE4BEG[11] ,
    \Tile_X1Y14_EE4BEG[10] ,
    \Tile_X1Y14_EE4BEG[9] ,
    \Tile_X1Y14_EE4BEG[8] ,
    \Tile_X1Y14_EE4BEG[7] ,
    \Tile_X1Y14_EE4BEG[6] ,
    \Tile_X1Y14_EE4BEG[5] ,
    \Tile_X1Y14_EE4BEG[4] ,
    \Tile_X1Y14_EE4BEG[3] ,
    \Tile_X1Y14_EE4BEG[2] ,
    \Tile_X1Y14_EE4BEG[1] ,
    \Tile_X1Y14_EE4BEG[0] }),
    .EE4END({\Tile_X0Y14_EE4BEG[15] ,
    \Tile_X0Y14_EE4BEG[14] ,
    \Tile_X0Y14_EE4BEG[13] ,
    \Tile_X0Y14_EE4BEG[12] ,
    \Tile_X0Y14_EE4BEG[11] ,
    \Tile_X0Y14_EE4BEG[10] ,
    \Tile_X0Y14_EE4BEG[9] ,
    \Tile_X0Y14_EE4BEG[8] ,
    \Tile_X0Y14_EE4BEG[7] ,
    \Tile_X0Y14_EE4BEG[6] ,
    \Tile_X0Y14_EE4BEG[5] ,
    \Tile_X0Y14_EE4BEG[4] ,
    \Tile_X0Y14_EE4BEG[3] ,
    \Tile_X0Y14_EE4BEG[2] ,
    \Tile_X0Y14_EE4BEG[1] ,
    \Tile_X0Y14_EE4BEG[0] }),
    .FrameData({\Tile_X0Y14_FrameData_O[31] ,
    \Tile_X0Y14_FrameData_O[30] ,
    \Tile_X0Y14_FrameData_O[29] ,
    \Tile_X0Y14_FrameData_O[28] ,
    \Tile_X0Y14_FrameData_O[27] ,
    \Tile_X0Y14_FrameData_O[26] ,
    \Tile_X0Y14_FrameData_O[25] ,
    \Tile_X0Y14_FrameData_O[24] ,
    \Tile_X0Y14_FrameData_O[23] ,
    \Tile_X0Y14_FrameData_O[22] ,
    \Tile_X0Y14_FrameData_O[21] ,
    \Tile_X0Y14_FrameData_O[20] ,
    \Tile_X0Y14_FrameData_O[19] ,
    \Tile_X0Y14_FrameData_O[18] ,
    \Tile_X0Y14_FrameData_O[17] ,
    \Tile_X0Y14_FrameData_O[16] ,
    \Tile_X0Y14_FrameData_O[15] ,
    \Tile_X0Y14_FrameData_O[14] ,
    \Tile_X0Y14_FrameData_O[13] ,
    \Tile_X0Y14_FrameData_O[12] ,
    \Tile_X0Y14_FrameData_O[11] ,
    \Tile_X0Y14_FrameData_O[10] ,
    \Tile_X0Y14_FrameData_O[9] ,
    \Tile_X0Y14_FrameData_O[8] ,
    \Tile_X0Y14_FrameData_O[7] ,
    \Tile_X0Y14_FrameData_O[6] ,
    \Tile_X0Y14_FrameData_O[5] ,
    \Tile_X0Y14_FrameData_O[4] ,
    \Tile_X0Y14_FrameData_O[3] ,
    \Tile_X0Y14_FrameData_O[2] ,
    \Tile_X0Y14_FrameData_O[1] ,
    \Tile_X0Y14_FrameData_O[0] }),
    .FrameData_O({\Tile_X1Y14_FrameData_O[31] ,
    \Tile_X1Y14_FrameData_O[30] ,
    \Tile_X1Y14_FrameData_O[29] ,
    \Tile_X1Y14_FrameData_O[28] ,
    \Tile_X1Y14_FrameData_O[27] ,
    \Tile_X1Y14_FrameData_O[26] ,
    \Tile_X1Y14_FrameData_O[25] ,
    \Tile_X1Y14_FrameData_O[24] ,
    \Tile_X1Y14_FrameData_O[23] ,
    \Tile_X1Y14_FrameData_O[22] ,
    \Tile_X1Y14_FrameData_O[21] ,
    \Tile_X1Y14_FrameData_O[20] ,
    \Tile_X1Y14_FrameData_O[19] ,
    \Tile_X1Y14_FrameData_O[18] ,
    \Tile_X1Y14_FrameData_O[17] ,
    \Tile_X1Y14_FrameData_O[16] ,
    \Tile_X1Y14_FrameData_O[15] ,
    \Tile_X1Y14_FrameData_O[14] ,
    \Tile_X1Y14_FrameData_O[13] ,
    \Tile_X1Y14_FrameData_O[12] ,
    \Tile_X1Y14_FrameData_O[11] ,
    \Tile_X1Y14_FrameData_O[10] ,
    \Tile_X1Y14_FrameData_O[9] ,
    \Tile_X1Y14_FrameData_O[8] ,
    \Tile_X1Y14_FrameData_O[7] ,
    \Tile_X1Y14_FrameData_O[6] ,
    \Tile_X1Y14_FrameData_O[5] ,
    \Tile_X1Y14_FrameData_O[4] ,
    \Tile_X1Y14_FrameData_O[3] ,
    \Tile_X1Y14_FrameData_O[2] ,
    \Tile_X1Y14_FrameData_O[1] ,
    \Tile_X1Y14_FrameData_O[0] }),
    .FrameStrobe({\Tile_X1Y15_FrameStrobe_O[19] ,
    \Tile_X1Y15_FrameStrobe_O[18] ,
    \Tile_X1Y15_FrameStrobe_O[17] ,
    \Tile_X1Y15_FrameStrobe_O[16] ,
    \Tile_X1Y15_FrameStrobe_O[15] ,
    \Tile_X1Y15_FrameStrobe_O[14] ,
    \Tile_X1Y15_FrameStrobe_O[13] ,
    \Tile_X1Y15_FrameStrobe_O[12] ,
    \Tile_X1Y15_FrameStrobe_O[11] ,
    \Tile_X1Y15_FrameStrobe_O[10] ,
    \Tile_X1Y15_FrameStrobe_O[9] ,
    \Tile_X1Y15_FrameStrobe_O[8] ,
    \Tile_X1Y15_FrameStrobe_O[7] ,
    \Tile_X1Y15_FrameStrobe_O[6] ,
    \Tile_X1Y15_FrameStrobe_O[5] ,
    \Tile_X1Y15_FrameStrobe_O[4] ,
    \Tile_X1Y15_FrameStrobe_O[3] ,
    \Tile_X1Y15_FrameStrobe_O[2] ,
    \Tile_X1Y15_FrameStrobe_O[1] ,
    \Tile_X1Y15_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X1Y14_FrameStrobe_O[19] ,
    \Tile_X1Y14_FrameStrobe_O[18] ,
    \Tile_X1Y14_FrameStrobe_O[17] ,
    \Tile_X1Y14_FrameStrobe_O[16] ,
    \Tile_X1Y14_FrameStrobe_O[15] ,
    \Tile_X1Y14_FrameStrobe_O[14] ,
    \Tile_X1Y14_FrameStrobe_O[13] ,
    \Tile_X1Y14_FrameStrobe_O[12] ,
    \Tile_X1Y14_FrameStrobe_O[11] ,
    \Tile_X1Y14_FrameStrobe_O[10] ,
    \Tile_X1Y14_FrameStrobe_O[9] ,
    \Tile_X1Y14_FrameStrobe_O[8] ,
    \Tile_X1Y14_FrameStrobe_O[7] ,
    \Tile_X1Y14_FrameStrobe_O[6] ,
    \Tile_X1Y14_FrameStrobe_O[5] ,
    \Tile_X1Y14_FrameStrobe_O[4] ,
    \Tile_X1Y14_FrameStrobe_O[3] ,
    \Tile_X1Y14_FrameStrobe_O[2] ,
    \Tile_X1Y14_FrameStrobe_O[1] ,
    \Tile_X1Y14_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X1Y14_N1BEG[3] ,
    \Tile_X1Y14_N1BEG[2] ,
    \Tile_X1Y14_N1BEG[1] ,
    \Tile_X1Y14_N1BEG[0] }),
    .N1END({\Tile_X1Y15_N1BEG[3] ,
    \Tile_X1Y15_N1BEG[2] ,
    \Tile_X1Y15_N1BEG[1] ,
    \Tile_X1Y15_N1BEG[0] }),
    .N2BEG({\Tile_X1Y14_N2BEG[7] ,
    \Tile_X1Y14_N2BEG[6] ,
    \Tile_X1Y14_N2BEG[5] ,
    \Tile_X1Y14_N2BEG[4] ,
    \Tile_X1Y14_N2BEG[3] ,
    \Tile_X1Y14_N2BEG[2] ,
    \Tile_X1Y14_N2BEG[1] ,
    \Tile_X1Y14_N2BEG[0] }),
    .N2BEGb({\Tile_X1Y14_N2BEGb[7] ,
    \Tile_X1Y14_N2BEGb[6] ,
    \Tile_X1Y14_N2BEGb[5] ,
    \Tile_X1Y14_N2BEGb[4] ,
    \Tile_X1Y14_N2BEGb[3] ,
    \Tile_X1Y14_N2BEGb[2] ,
    \Tile_X1Y14_N2BEGb[1] ,
    \Tile_X1Y14_N2BEGb[0] }),
    .N2END({\Tile_X1Y15_N2BEGb[7] ,
    \Tile_X1Y15_N2BEGb[6] ,
    \Tile_X1Y15_N2BEGb[5] ,
    \Tile_X1Y15_N2BEGb[4] ,
    \Tile_X1Y15_N2BEGb[3] ,
    \Tile_X1Y15_N2BEGb[2] ,
    \Tile_X1Y15_N2BEGb[1] ,
    \Tile_X1Y15_N2BEGb[0] }),
    .N2MID({\Tile_X1Y15_N2BEG[7] ,
    \Tile_X1Y15_N2BEG[6] ,
    \Tile_X1Y15_N2BEG[5] ,
    \Tile_X1Y15_N2BEG[4] ,
    \Tile_X1Y15_N2BEG[3] ,
    \Tile_X1Y15_N2BEG[2] ,
    \Tile_X1Y15_N2BEG[1] ,
    \Tile_X1Y15_N2BEG[0] }),
    .N4BEG({\Tile_X1Y14_N4BEG[15] ,
    \Tile_X1Y14_N4BEG[14] ,
    \Tile_X1Y14_N4BEG[13] ,
    \Tile_X1Y14_N4BEG[12] ,
    \Tile_X1Y14_N4BEG[11] ,
    \Tile_X1Y14_N4BEG[10] ,
    \Tile_X1Y14_N4BEG[9] ,
    \Tile_X1Y14_N4BEG[8] ,
    \Tile_X1Y14_N4BEG[7] ,
    \Tile_X1Y14_N4BEG[6] ,
    \Tile_X1Y14_N4BEG[5] ,
    \Tile_X1Y14_N4BEG[4] ,
    \Tile_X1Y14_N4BEG[3] ,
    \Tile_X1Y14_N4BEG[2] ,
    \Tile_X1Y14_N4BEG[1] ,
    \Tile_X1Y14_N4BEG[0] }),
    .N4END({\Tile_X1Y15_N4BEG[15] ,
    \Tile_X1Y15_N4BEG[14] ,
    \Tile_X1Y15_N4BEG[13] ,
    \Tile_X1Y15_N4BEG[12] ,
    \Tile_X1Y15_N4BEG[11] ,
    \Tile_X1Y15_N4BEG[10] ,
    \Tile_X1Y15_N4BEG[9] ,
    \Tile_X1Y15_N4BEG[8] ,
    \Tile_X1Y15_N4BEG[7] ,
    \Tile_X1Y15_N4BEG[6] ,
    \Tile_X1Y15_N4BEG[5] ,
    \Tile_X1Y15_N4BEG[4] ,
    \Tile_X1Y15_N4BEG[3] ,
    \Tile_X1Y15_N4BEG[2] ,
    \Tile_X1Y15_N4BEG[1] ,
    \Tile_X1Y15_N4BEG[0] }),
    .NN4BEG({\Tile_X1Y14_NN4BEG[15] ,
    \Tile_X1Y14_NN4BEG[14] ,
    \Tile_X1Y14_NN4BEG[13] ,
    \Tile_X1Y14_NN4BEG[12] ,
    \Tile_X1Y14_NN4BEG[11] ,
    \Tile_X1Y14_NN4BEG[10] ,
    \Tile_X1Y14_NN4BEG[9] ,
    \Tile_X1Y14_NN4BEG[8] ,
    \Tile_X1Y14_NN4BEG[7] ,
    \Tile_X1Y14_NN4BEG[6] ,
    \Tile_X1Y14_NN4BEG[5] ,
    \Tile_X1Y14_NN4BEG[4] ,
    \Tile_X1Y14_NN4BEG[3] ,
    \Tile_X1Y14_NN4BEG[2] ,
    \Tile_X1Y14_NN4BEG[1] ,
    \Tile_X1Y14_NN4BEG[0] }),
    .NN4END({\Tile_X1Y15_NN4BEG[15] ,
    \Tile_X1Y15_NN4BEG[14] ,
    \Tile_X1Y15_NN4BEG[13] ,
    \Tile_X1Y15_NN4BEG[12] ,
    \Tile_X1Y15_NN4BEG[11] ,
    \Tile_X1Y15_NN4BEG[10] ,
    \Tile_X1Y15_NN4BEG[9] ,
    \Tile_X1Y15_NN4BEG[8] ,
    \Tile_X1Y15_NN4BEG[7] ,
    \Tile_X1Y15_NN4BEG[6] ,
    \Tile_X1Y15_NN4BEG[5] ,
    \Tile_X1Y15_NN4BEG[4] ,
    \Tile_X1Y15_NN4BEG[3] ,
    \Tile_X1Y15_NN4BEG[2] ,
    \Tile_X1Y15_NN4BEG[1] ,
    \Tile_X1Y15_NN4BEG[0] }),
    .S1BEG({\Tile_X1Y14_S1BEG[3] ,
    \Tile_X1Y14_S1BEG[2] ,
    \Tile_X1Y14_S1BEG[1] ,
    \Tile_X1Y14_S1BEG[0] }),
    .S1END({\Tile_X1Y13_S1BEG[3] ,
    \Tile_X1Y13_S1BEG[2] ,
    \Tile_X1Y13_S1BEG[1] ,
    \Tile_X1Y13_S1BEG[0] }),
    .S2BEG({\Tile_X1Y14_S2BEG[7] ,
    \Tile_X1Y14_S2BEG[6] ,
    \Tile_X1Y14_S2BEG[5] ,
    \Tile_X1Y14_S2BEG[4] ,
    \Tile_X1Y14_S2BEG[3] ,
    \Tile_X1Y14_S2BEG[2] ,
    \Tile_X1Y14_S2BEG[1] ,
    \Tile_X1Y14_S2BEG[0] }),
    .S2BEGb({\Tile_X1Y14_S2BEGb[7] ,
    \Tile_X1Y14_S2BEGb[6] ,
    \Tile_X1Y14_S2BEGb[5] ,
    \Tile_X1Y14_S2BEGb[4] ,
    \Tile_X1Y14_S2BEGb[3] ,
    \Tile_X1Y14_S2BEGb[2] ,
    \Tile_X1Y14_S2BEGb[1] ,
    \Tile_X1Y14_S2BEGb[0] }),
    .S2END({\Tile_X1Y13_S2BEGb[7] ,
    \Tile_X1Y13_S2BEGb[6] ,
    \Tile_X1Y13_S2BEGb[5] ,
    \Tile_X1Y13_S2BEGb[4] ,
    \Tile_X1Y13_S2BEGb[3] ,
    \Tile_X1Y13_S2BEGb[2] ,
    \Tile_X1Y13_S2BEGb[1] ,
    \Tile_X1Y13_S2BEGb[0] }),
    .S2MID({\Tile_X1Y13_S2BEG[7] ,
    \Tile_X1Y13_S2BEG[6] ,
    \Tile_X1Y13_S2BEG[5] ,
    \Tile_X1Y13_S2BEG[4] ,
    \Tile_X1Y13_S2BEG[3] ,
    \Tile_X1Y13_S2BEG[2] ,
    \Tile_X1Y13_S2BEG[1] ,
    \Tile_X1Y13_S2BEG[0] }),
    .S4BEG({\Tile_X1Y14_S4BEG[15] ,
    \Tile_X1Y14_S4BEG[14] ,
    \Tile_X1Y14_S4BEG[13] ,
    \Tile_X1Y14_S4BEG[12] ,
    \Tile_X1Y14_S4BEG[11] ,
    \Tile_X1Y14_S4BEG[10] ,
    \Tile_X1Y14_S4BEG[9] ,
    \Tile_X1Y14_S4BEG[8] ,
    \Tile_X1Y14_S4BEG[7] ,
    \Tile_X1Y14_S4BEG[6] ,
    \Tile_X1Y14_S4BEG[5] ,
    \Tile_X1Y14_S4BEG[4] ,
    \Tile_X1Y14_S4BEG[3] ,
    \Tile_X1Y14_S4BEG[2] ,
    \Tile_X1Y14_S4BEG[1] ,
    \Tile_X1Y14_S4BEG[0] }),
    .S4END({\Tile_X1Y13_S4BEG[15] ,
    \Tile_X1Y13_S4BEG[14] ,
    \Tile_X1Y13_S4BEG[13] ,
    \Tile_X1Y13_S4BEG[12] ,
    \Tile_X1Y13_S4BEG[11] ,
    \Tile_X1Y13_S4BEG[10] ,
    \Tile_X1Y13_S4BEG[9] ,
    \Tile_X1Y13_S4BEG[8] ,
    \Tile_X1Y13_S4BEG[7] ,
    \Tile_X1Y13_S4BEG[6] ,
    \Tile_X1Y13_S4BEG[5] ,
    \Tile_X1Y13_S4BEG[4] ,
    \Tile_X1Y13_S4BEG[3] ,
    \Tile_X1Y13_S4BEG[2] ,
    \Tile_X1Y13_S4BEG[1] ,
    \Tile_X1Y13_S4BEG[0] }),
    .SS4BEG({\Tile_X1Y14_SS4BEG[15] ,
    \Tile_X1Y14_SS4BEG[14] ,
    \Tile_X1Y14_SS4BEG[13] ,
    \Tile_X1Y14_SS4BEG[12] ,
    \Tile_X1Y14_SS4BEG[11] ,
    \Tile_X1Y14_SS4BEG[10] ,
    \Tile_X1Y14_SS4BEG[9] ,
    \Tile_X1Y14_SS4BEG[8] ,
    \Tile_X1Y14_SS4BEG[7] ,
    \Tile_X1Y14_SS4BEG[6] ,
    \Tile_X1Y14_SS4BEG[5] ,
    \Tile_X1Y14_SS4BEG[4] ,
    \Tile_X1Y14_SS4BEG[3] ,
    \Tile_X1Y14_SS4BEG[2] ,
    \Tile_X1Y14_SS4BEG[1] ,
    \Tile_X1Y14_SS4BEG[0] }),
    .SS4END({\Tile_X1Y13_SS4BEG[15] ,
    \Tile_X1Y13_SS4BEG[14] ,
    \Tile_X1Y13_SS4BEG[13] ,
    \Tile_X1Y13_SS4BEG[12] ,
    \Tile_X1Y13_SS4BEG[11] ,
    \Tile_X1Y13_SS4BEG[10] ,
    \Tile_X1Y13_SS4BEG[9] ,
    \Tile_X1Y13_SS4BEG[8] ,
    \Tile_X1Y13_SS4BEG[7] ,
    \Tile_X1Y13_SS4BEG[6] ,
    \Tile_X1Y13_SS4BEG[5] ,
    \Tile_X1Y13_SS4BEG[4] ,
    \Tile_X1Y13_SS4BEG[3] ,
    \Tile_X1Y13_SS4BEG[2] ,
    \Tile_X1Y13_SS4BEG[1] ,
    \Tile_X1Y13_SS4BEG[0] }),
    .W1BEG({\Tile_X1Y14_W1BEG[3] ,
    \Tile_X1Y14_W1BEG[2] ,
    \Tile_X1Y14_W1BEG[1] ,
    \Tile_X1Y14_W1BEG[0] }),
    .W1END({\Tile_X2Y14_W1BEG[3] ,
    \Tile_X2Y14_W1BEG[2] ,
    \Tile_X2Y14_W1BEG[1] ,
    \Tile_X2Y14_W1BEG[0] }),
    .W2BEG({\Tile_X1Y14_W2BEG[7] ,
    \Tile_X1Y14_W2BEG[6] ,
    \Tile_X1Y14_W2BEG[5] ,
    \Tile_X1Y14_W2BEG[4] ,
    \Tile_X1Y14_W2BEG[3] ,
    \Tile_X1Y14_W2BEG[2] ,
    \Tile_X1Y14_W2BEG[1] ,
    \Tile_X1Y14_W2BEG[0] }),
    .W2BEGb({\Tile_X1Y14_W2BEGb[7] ,
    \Tile_X1Y14_W2BEGb[6] ,
    \Tile_X1Y14_W2BEGb[5] ,
    \Tile_X1Y14_W2BEGb[4] ,
    \Tile_X1Y14_W2BEGb[3] ,
    \Tile_X1Y14_W2BEGb[2] ,
    \Tile_X1Y14_W2BEGb[1] ,
    \Tile_X1Y14_W2BEGb[0] }),
    .W2END({\Tile_X2Y14_W2BEGb[7] ,
    \Tile_X2Y14_W2BEGb[6] ,
    \Tile_X2Y14_W2BEGb[5] ,
    \Tile_X2Y14_W2BEGb[4] ,
    \Tile_X2Y14_W2BEGb[3] ,
    \Tile_X2Y14_W2BEGb[2] ,
    \Tile_X2Y14_W2BEGb[1] ,
    \Tile_X2Y14_W2BEGb[0] }),
    .W2MID({\Tile_X2Y14_W2BEG[7] ,
    \Tile_X2Y14_W2BEG[6] ,
    \Tile_X2Y14_W2BEG[5] ,
    \Tile_X2Y14_W2BEG[4] ,
    \Tile_X2Y14_W2BEG[3] ,
    \Tile_X2Y14_W2BEG[2] ,
    \Tile_X2Y14_W2BEG[1] ,
    \Tile_X2Y14_W2BEG[0] }),
    .W6BEG({\Tile_X1Y14_W6BEG[11] ,
    \Tile_X1Y14_W6BEG[10] ,
    \Tile_X1Y14_W6BEG[9] ,
    \Tile_X1Y14_W6BEG[8] ,
    \Tile_X1Y14_W6BEG[7] ,
    \Tile_X1Y14_W6BEG[6] ,
    \Tile_X1Y14_W6BEG[5] ,
    \Tile_X1Y14_W6BEG[4] ,
    \Tile_X1Y14_W6BEG[3] ,
    \Tile_X1Y14_W6BEG[2] ,
    \Tile_X1Y14_W6BEG[1] ,
    \Tile_X1Y14_W6BEG[0] }),
    .W6END({\Tile_X2Y14_W6BEG[11] ,
    \Tile_X2Y14_W6BEG[10] ,
    \Tile_X2Y14_W6BEG[9] ,
    \Tile_X2Y14_W6BEG[8] ,
    \Tile_X2Y14_W6BEG[7] ,
    \Tile_X2Y14_W6BEG[6] ,
    \Tile_X2Y14_W6BEG[5] ,
    \Tile_X2Y14_W6BEG[4] ,
    \Tile_X2Y14_W6BEG[3] ,
    \Tile_X2Y14_W6BEG[2] ,
    \Tile_X2Y14_W6BEG[1] ,
    \Tile_X2Y14_W6BEG[0] }),
    .WW4BEG({\Tile_X1Y14_WW4BEG[15] ,
    \Tile_X1Y14_WW4BEG[14] ,
    \Tile_X1Y14_WW4BEG[13] ,
    \Tile_X1Y14_WW4BEG[12] ,
    \Tile_X1Y14_WW4BEG[11] ,
    \Tile_X1Y14_WW4BEG[10] ,
    \Tile_X1Y14_WW4BEG[9] ,
    \Tile_X1Y14_WW4BEG[8] ,
    \Tile_X1Y14_WW4BEG[7] ,
    \Tile_X1Y14_WW4BEG[6] ,
    \Tile_X1Y14_WW4BEG[5] ,
    \Tile_X1Y14_WW4BEG[4] ,
    \Tile_X1Y14_WW4BEG[3] ,
    \Tile_X1Y14_WW4BEG[2] ,
    \Tile_X1Y14_WW4BEG[1] ,
    \Tile_X1Y14_WW4BEG[0] }),
    .WW4END({\Tile_X2Y14_WW4BEG[15] ,
    \Tile_X2Y14_WW4BEG[14] ,
    \Tile_X2Y14_WW4BEG[13] ,
    \Tile_X2Y14_WW4BEG[12] ,
    \Tile_X2Y14_WW4BEG[11] ,
    \Tile_X2Y14_WW4BEG[10] ,
    \Tile_X2Y14_WW4BEG[9] ,
    \Tile_X2Y14_WW4BEG[8] ,
    \Tile_X2Y14_WW4BEG[7] ,
    \Tile_X2Y14_WW4BEG[6] ,
    \Tile_X2Y14_WW4BEG[5] ,
    \Tile_X2Y14_WW4BEG[4] ,
    \Tile_X2Y14_WW4BEG[3] ,
    \Tile_X2Y14_WW4BEG[2] ,
    \Tile_X2Y14_WW4BEG[1] ,
    \Tile_X2Y14_WW4BEG[0] }));
 S_term_single Tile_X1Y15_S_term_single (.Co(Tile_X1Y15_Co),
    .UserCLK(UserCLK),
    .UserCLKo(Tile_X1Y15_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .FrameData({FrameData[511],
    FrameData[510],
    FrameData[509],
    FrameData[508],
    FrameData[507],
    FrameData[506],
    FrameData[505],
    FrameData[504],
    FrameData[503],
    FrameData[502],
    FrameData[501],
    FrameData[500],
    FrameData[499],
    FrameData[498],
    FrameData[497],
    FrameData[496],
    FrameData[495],
    FrameData[494],
    FrameData[493],
    FrameData[492],
    FrameData[491],
    FrameData[490],
    FrameData[489],
    FrameData[488],
    FrameData[487],
    FrameData[486],
    FrameData[485],
    FrameData[484],
    FrameData[483],
    FrameData[482],
    FrameData[481],
    FrameData[480]}),
    .FrameData_O({\Tile_X1Y15_FrameData_O[31] ,
    \Tile_X1Y15_FrameData_O[30] ,
    \Tile_X1Y15_FrameData_O[29] ,
    \Tile_X1Y15_FrameData_O[28] ,
    \Tile_X1Y15_FrameData_O[27] ,
    \Tile_X1Y15_FrameData_O[26] ,
    \Tile_X1Y15_FrameData_O[25] ,
    \Tile_X1Y15_FrameData_O[24] ,
    \Tile_X1Y15_FrameData_O[23] ,
    \Tile_X1Y15_FrameData_O[22] ,
    \Tile_X1Y15_FrameData_O[21] ,
    \Tile_X1Y15_FrameData_O[20] ,
    \Tile_X1Y15_FrameData_O[19] ,
    \Tile_X1Y15_FrameData_O[18] ,
    \Tile_X1Y15_FrameData_O[17] ,
    \Tile_X1Y15_FrameData_O[16] ,
    \Tile_X1Y15_FrameData_O[15] ,
    \Tile_X1Y15_FrameData_O[14] ,
    \Tile_X1Y15_FrameData_O[13] ,
    \Tile_X1Y15_FrameData_O[12] ,
    \Tile_X1Y15_FrameData_O[11] ,
    \Tile_X1Y15_FrameData_O[10] ,
    \Tile_X1Y15_FrameData_O[9] ,
    \Tile_X1Y15_FrameData_O[8] ,
    \Tile_X1Y15_FrameData_O[7] ,
    \Tile_X1Y15_FrameData_O[6] ,
    \Tile_X1Y15_FrameData_O[5] ,
    \Tile_X1Y15_FrameData_O[4] ,
    \Tile_X1Y15_FrameData_O[3] ,
    \Tile_X1Y15_FrameData_O[2] ,
    \Tile_X1Y15_FrameData_O[1] ,
    \Tile_X1Y15_FrameData_O[0] }),
    .FrameStrobe({FrameStrobe[39],
    FrameStrobe[38],
    FrameStrobe[37],
    FrameStrobe[36],
    FrameStrobe[35],
    FrameStrobe[34],
    FrameStrobe[33],
    FrameStrobe[32],
    FrameStrobe[31],
    FrameStrobe[30],
    FrameStrobe[29],
    FrameStrobe[28],
    FrameStrobe[27],
    FrameStrobe[26],
    FrameStrobe[25],
    FrameStrobe[24],
    FrameStrobe[23],
    FrameStrobe[22],
    FrameStrobe[21],
    FrameStrobe[20]}),
    .FrameStrobe_O({\Tile_X1Y15_FrameStrobe_O[19] ,
    \Tile_X1Y15_FrameStrobe_O[18] ,
    \Tile_X1Y15_FrameStrobe_O[17] ,
    \Tile_X1Y15_FrameStrobe_O[16] ,
    \Tile_X1Y15_FrameStrobe_O[15] ,
    \Tile_X1Y15_FrameStrobe_O[14] ,
    \Tile_X1Y15_FrameStrobe_O[13] ,
    \Tile_X1Y15_FrameStrobe_O[12] ,
    \Tile_X1Y15_FrameStrobe_O[11] ,
    \Tile_X1Y15_FrameStrobe_O[10] ,
    \Tile_X1Y15_FrameStrobe_O[9] ,
    \Tile_X1Y15_FrameStrobe_O[8] ,
    \Tile_X1Y15_FrameStrobe_O[7] ,
    \Tile_X1Y15_FrameStrobe_O[6] ,
    \Tile_X1Y15_FrameStrobe_O[5] ,
    \Tile_X1Y15_FrameStrobe_O[4] ,
    \Tile_X1Y15_FrameStrobe_O[3] ,
    \Tile_X1Y15_FrameStrobe_O[2] ,
    \Tile_X1Y15_FrameStrobe_O[1] ,
    \Tile_X1Y15_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X1Y15_N1BEG[3] ,
    \Tile_X1Y15_N1BEG[2] ,
    \Tile_X1Y15_N1BEG[1] ,
    \Tile_X1Y15_N1BEG[0] }),
    .N2BEG({\Tile_X1Y15_N2BEG[7] ,
    \Tile_X1Y15_N2BEG[6] ,
    \Tile_X1Y15_N2BEG[5] ,
    \Tile_X1Y15_N2BEG[4] ,
    \Tile_X1Y15_N2BEG[3] ,
    \Tile_X1Y15_N2BEG[2] ,
    \Tile_X1Y15_N2BEG[1] ,
    \Tile_X1Y15_N2BEG[0] }),
    .N2BEGb({\Tile_X1Y15_N2BEGb[7] ,
    \Tile_X1Y15_N2BEGb[6] ,
    \Tile_X1Y15_N2BEGb[5] ,
    \Tile_X1Y15_N2BEGb[4] ,
    \Tile_X1Y15_N2BEGb[3] ,
    \Tile_X1Y15_N2BEGb[2] ,
    \Tile_X1Y15_N2BEGb[1] ,
    \Tile_X1Y15_N2BEGb[0] }),
    .N4BEG({\Tile_X1Y15_N4BEG[15] ,
    \Tile_X1Y15_N4BEG[14] ,
    \Tile_X1Y15_N4BEG[13] ,
    \Tile_X1Y15_N4BEG[12] ,
    \Tile_X1Y15_N4BEG[11] ,
    \Tile_X1Y15_N4BEG[10] ,
    \Tile_X1Y15_N4BEG[9] ,
    \Tile_X1Y15_N4BEG[8] ,
    \Tile_X1Y15_N4BEG[7] ,
    \Tile_X1Y15_N4BEG[6] ,
    \Tile_X1Y15_N4BEG[5] ,
    \Tile_X1Y15_N4BEG[4] ,
    \Tile_X1Y15_N4BEG[3] ,
    \Tile_X1Y15_N4BEG[2] ,
    \Tile_X1Y15_N4BEG[1] ,
    \Tile_X1Y15_N4BEG[0] }),
    .NN4BEG({\Tile_X1Y15_NN4BEG[15] ,
    \Tile_X1Y15_NN4BEG[14] ,
    \Tile_X1Y15_NN4BEG[13] ,
    \Tile_X1Y15_NN4BEG[12] ,
    \Tile_X1Y15_NN4BEG[11] ,
    \Tile_X1Y15_NN4BEG[10] ,
    \Tile_X1Y15_NN4BEG[9] ,
    \Tile_X1Y15_NN4BEG[8] ,
    \Tile_X1Y15_NN4BEG[7] ,
    \Tile_X1Y15_NN4BEG[6] ,
    \Tile_X1Y15_NN4BEG[5] ,
    \Tile_X1Y15_NN4BEG[4] ,
    \Tile_X1Y15_NN4BEG[3] ,
    \Tile_X1Y15_NN4BEG[2] ,
    \Tile_X1Y15_NN4BEG[1] ,
    \Tile_X1Y15_NN4BEG[0] }),
    .S1END({\Tile_X1Y14_S1BEG[3] ,
    \Tile_X1Y14_S1BEG[2] ,
    \Tile_X1Y14_S1BEG[1] ,
    \Tile_X1Y14_S1BEG[0] }),
    .S2END({\Tile_X1Y14_S2BEGb[7] ,
    \Tile_X1Y14_S2BEGb[6] ,
    \Tile_X1Y14_S2BEGb[5] ,
    \Tile_X1Y14_S2BEGb[4] ,
    \Tile_X1Y14_S2BEGb[3] ,
    \Tile_X1Y14_S2BEGb[2] ,
    \Tile_X1Y14_S2BEGb[1] ,
    \Tile_X1Y14_S2BEGb[0] }),
    .S2MID({\Tile_X1Y14_S2BEG[7] ,
    \Tile_X1Y14_S2BEG[6] ,
    \Tile_X1Y14_S2BEG[5] ,
    \Tile_X1Y14_S2BEG[4] ,
    \Tile_X1Y14_S2BEG[3] ,
    \Tile_X1Y14_S2BEG[2] ,
    \Tile_X1Y14_S2BEG[1] ,
    \Tile_X1Y14_S2BEG[0] }),
    .S4END({\Tile_X1Y14_S4BEG[15] ,
    \Tile_X1Y14_S4BEG[14] ,
    \Tile_X1Y14_S4BEG[13] ,
    \Tile_X1Y14_S4BEG[12] ,
    \Tile_X1Y14_S4BEG[11] ,
    \Tile_X1Y14_S4BEG[10] ,
    \Tile_X1Y14_S4BEG[9] ,
    \Tile_X1Y14_S4BEG[8] ,
    \Tile_X1Y14_S4BEG[7] ,
    \Tile_X1Y14_S4BEG[6] ,
    \Tile_X1Y14_S4BEG[5] ,
    \Tile_X1Y14_S4BEG[4] ,
    \Tile_X1Y14_S4BEG[3] ,
    \Tile_X1Y14_S4BEG[2] ,
    \Tile_X1Y14_S4BEG[1] ,
    \Tile_X1Y14_S4BEG[0] }),
    .SS4END({\Tile_X1Y14_SS4BEG[15] ,
    \Tile_X1Y14_SS4BEG[14] ,
    \Tile_X1Y14_SS4BEG[13] ,
    \Tile_X1Y14_SS4BEG[12] ,
    \Tile_X1Y14_SS4BEG[11] ,
    \Tile_X1Y14_SS4BEG[10] ,
    \Tile_X1Y14_SS4BEG[9] ,
    \Tile_X1Y14_SS4BEG[8] ,
    \Tile_X1Y14_SS4BEG[7] ,
    \Tile_X1Y14_SS4BEG[6] ,
    \Tile_X1Y14_SS4BEG[5] ,
    \Tile_X1Y14_SS4BEG[4] ,
    \Tile_X1Y14_SS4BEG[3] ,
    \Tile_X1Y14_SS4BEG[2] ,
    \Tile_X1Y14_SS4BEG[1] ,
    \Tile_X1Y14_SS4BEG[0] }));
 LUT4AB Tile_X1Y1_LUT4AB (.Ci(Tile_X1Y2_Co),
    .Co(Tile_X1Y1_Co),
    .UserCLK(Tile_X1Y2_UserCLKo),
    .UserCLKo(Tile_X1Y1_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X1Y1_E1BEG[3] ,
    \Tile_X1Y1_E1BEG[2] ,
    \Tile_X1Y1_E1BEG[1] ,
    \Tile_X1Y1_E1BEG[0] }),
    .E1END({\Tile_X0Y1_E1BEG[3] ,
    \Tile_X0Y1_E1BEG[2] ,
    \Tile_X0Y1_E1BEG[1] ,
    \Tile_X0Y1_E1BEG[0] }),
    .E2BEG({\Tile_X1Y1_E2BEG[7] ,
    \Tile_X1Y1_E2BEG[6] ,
    \Tile_X1Y1_E2BEG[5] ,
    \Tile_X1Y1_E2BEG[4] ,
    \Tile_X1Y1_E2BEG[3] ,
    \Tile_X1Y1_E2BEG[2] ,
    \Tile_X1Y1_E2BEG[1] ,
    \Tile_X1Y1_E2BEG[0] }),
    .E2BEGb({\Tile_X1Y1_E2BEGb[7] ,
    \Tile_X1Y1_E2BEGb[6] ,
    \Tile_X1Y1_E2BEGb[5] ,
    \Tile_X1Y1_E2BEGb[4] ,
    \Tile_X1Y1_E2BEGb[3] ,
    \Tile_X1Y1_E2BEGb[2] ,
    \Tile_X1Y1_E2BEGb[1] ,
    \Tile_X1Y1_E2BEGb[0] }),
    .E2END({\Tile_X0Y1_E2BEGb[7] ,
    \Tile_X0Y1_E2BEGb[6] ,
    \Tile_X0Y1_E2BEGb[5] ,
    \Tile_X0Y1_E2BEGb[4] ,
    \Tile_X0Y1_E2BEGb[3] ,
    \Tile_X0Y1_E2BEGb[2] ,
    \Tile_X0Y1_E2BEGb[1] ,
    \Tile_X0Y1_E2BEGb[0] }),
    .E2MID({\Tile_X0Y1_E2BEG[7] ,
    \Tile_X0Y1_E2BEG[6] ,
    \Tile_X0Y1_E2BEG[5] ,
    \Tile_X0Y1_E2BEG[4] ,
    \Tile_X0Y1_E2BEG[3] ,
    \Tile_X0Y1_E2BEG[2] ,
    \Tile_X0Y1_E2BEG[1] ,
    \Tile_X0Y1_E2BEG[0] }),
    .E6BEG({\Tile_X1Y1_E6BEG[11] ,
    \Tile_X1Y1_E6BEG[10] ,
    \Tile_X1Y1_E6BEG[9] ,
    \Tile_X1Y1_E6BEG[8] ,
    \Tile_X1Y1_E6BEG[7] ,
    \Tile_X1Y1_E6BEG[6] ,
    \Tile_X1Y1_E6BEG[5] ,
    \Tile_X1Y1_E6BEG[4] ,
    \Tile_X1Y1_E6BEG[3] ,
    \Tile_X1Y1_E6BEG[2] ,
    \Tile_X1Y1_E6BEG[1] ,
    \Tile_X1Y1_E6BEG[0] }),
    .E6END({\Tile_X0Y1_E6BEG[11] ,
    \Tile_X0Y1_E6BEG[10] ,
    \Tile_X0Y1_E6BEG[9] ,
    \Tile_X0Y1_E6BEG[8] ,
    \Tile_X0Y1_E6BEG[7] ,
    \Tile_X0Y1_E6BEG[6] ,
    \Tile_X0Y1_E6BEG[5] ,
    \Tile_X0Y1_E6BEG[4] ,
    \Tile_X0Y1_E6BEG[3] ,
    \Tile_X0Y1_E6BEG[2] ,
    \Tile_X0Y1_E6BEG[1] ,
    \Tile_X0Y1_E6BEG[0] }),
    .EE4BEG({\Tile_X1Y1_EE4BEG[15] ,
    \Tile_X1Y1_EE4BEG[14] ,
    \Tile_X1Y1_EE4BEG[13] ,
    \Tile_X1Y1_EE4BEG[12] ,
    \Tile_X1Y1_EE4BEG[11] ,
    \Tile_X1Y1_EE4BEG[10] ,
    \Tile_X1Y1_EE4BEG[9] ,
    \Tile_X1Y1_EE4BEG[8] ,
    \Tile_X1Y1_EE4BEG[7] ,
    \Tile_X1Y1_EE4BEG[6] ,
    \Tile_X1Y1_EE4BEG[5] ,
    \Tile_X1Y1_EE4BEG[4] ,
    \Tile_X1Y1_EE4BEG[3] ,
    \Tile_X1Y1_EE4BEG[2] ,
    \Tile_X1Y1_EE4BEG[1] ,
    \Tile_X1Y1_EE4BEG[0] }),
    .EE4END({\Tile_X0Y1_EE4BEG[15] ,
    \Tile_X0Y1_EE4BEG[14] ,
    \Tile_X0Y1_EE4BEG[13] ,
    \Tile_X0Y1_EE4BEG[12] ,
    \Tile_X0Y1_EE4BEG[11] ,
    \Tile_X0Y1_EE4BEG[10] ,
    \Tile_X0Y1_EE4BEG[9] ,
    \Tile_X0Y1_EE4BEG[8] ,
    \Tile_X0Y1_EE4BEG[7] ,
    \Tile_X0Y1_EE4BEG[6] ,
    \Tile_X0Y1_EE4BEG[5] ,
    \Tile_X0Y1_EE4BEG[4] ,
    \Tile_X0Y1_EE4BEG[3] ,
    \Tile_X0Y1_EE4BEG[2] ,
    \Tile_X0Y1_EE4BEG[1] ,
    \Tile_X0Y1_EE4BEG[0] }),
    .FrameData({\Tile_X0Y1_FrameData_O[31] ,
    \Tile_X0Y1_FrameData_O[30] ,
    \Tile_X0Y1_FrameData_O[29] ,
    \Tile_X0Y1_FrameData_O[28] ,
    \Tile_X0Y1_FrameData_O[27] ,
    \Tile_X0Y1_FrameData_O[26] ,
    \Tile_X0Y1_FrameData_O[25] ,
    \Tile_X0Y1_FrameData_O[24] ,
    \Tile_X0Y1_FrameData_O[23] ,
    \Tile_X0Y1_FrameData_O[22] ,
    \Tile_X0Y1_FrameData_O[21] ,
    \Tile_X0Y1_FrameData_O[20] ,
    \Tile_X0Y1_FrameData_O[19] ,
    \Tile_X0Y1_FrameData_O[18] ,
    \Tile_X0Y1_FrameData_O[17] ,
    \Tile_X0Y1_FrameData_O[16] ,
    \Tile_X0Y1_FrameData_O[15] ,
    \Tile_X0Y1_FrameData_O[14] ,
    \Tile_X0Y1_FrameData_O[13] ,
    \Tile_X0Y1_FrameData_O[12] ,
    \Tile_X0Y1_FrameData_O[11] ,
    \Tile_X0Y1_FrameData_O[10] ,
    \Tile_X0Y1_FrameData_O[9] ,
    \Tile_X0Y1_FrameData_O[8] ,
    \Tile_X0Y1_FrameData_O[7] ,
    \Tile_X0Y1_FrameData_O[6] ,
    \Tile_X0Y1_FrameData_O[5] ,
    \Tile_X0Y1_FrameData_O[4] ,
    \Tile_X0Y1_FrameData_O[3] ,
    \Tile_X0Y1_FrameData_O[2] ,
    \Tile_X0Y1_FrameData_O[1] ,
    \Tile_X0Y1_FrameData_O[0] }),
    .FrameData_O({\Tile_X1Y1_FrameData_O[31] ,
    \Tile_X1Y1_FrameData_O[30] ,
    \Tile_X1Y1_FrameData_O[29] ,
    \Tile_X1Y1_FrameData_O[28] ,
    \Tile_X1Y1_FrameData_O[27] ,
    \Tile_X1Y1_FrameData_O[26] ,
    \Tile_X1Y1_FrameData_O[25] ,
    \Tile_X1Y1_FrameData_O[24] ,
    \Tile_X1Y1_FrameData_O[23] ,
    \Tile_X1Y1_FrameData_O[22] ,
    \Tile_X1Y1_FrameData_O[21] ,
    \Tile_X1Y1_FrameData_O[20] ,
    \Tile_X1Y1_FrameData_O[19] ,
    \Tile_X1Y1_FrameData_O[18] ,
    \Tile_X1Y1_FrameData_O[17] ,
    \Tile_X1Y1_FrameData_O[16] ,
    \Tile_X1Y1_FrameData_O[15] ,
    \Tile_X1Y1_FrameData_O[14] ,
    \Tile_X1Y1_FrameData_O[13] ,
    \Tile_X1Y1_FrameData_O[12] ,
    \Tile_X1Y1_FrameData_O[11] ,
    \Tile_X1Y1_FrameData_O[10] ,
    \Tile_X1Y1_FrameData_O[9] ,
    \Tile_X1Y1_FrameData_O[8] ,
    \Tile_X1Y1_FrameData_O[7] ,
    \Tile_X1Y1_FrameData_O[6] ,
    \Tile_X1Y1_FrameData_O[5] ,
    \Tile_X1Y1_FrameData_O[4] ,
    \Tile_X1Y1_FrameData_O[3] ,
    \Tile_X1Y1_FrameData_O[2] ,
    \Tile_X1Y1_FrameData_O[1] ,
    \Tile_X1Y1_FrameData_O[0] }),
    .FrameStrobe({\Tile_X1Y2_FrameStrobe_O[19] ,
    \Tile_X1Y2_FrameStrobe_O[18] ,
    \Tile_X1Y2_FrameStrobe_O[17] ,
    \Tile_X1Y2_FrameStrobe_O[16] ,
    \Tile_X1Y2_FrameStrobe_O[15] ,
    \Tile_X1Y2_FrameStrobe_O[14] ,
    \Tile_X1Y2_FrameStrobe_O[13] ,
    \Tile_X1Y2_FrameStrobe_O[12] ,
    \Tile_X1Y2_FrameStrobe_O[11] ,
    \Tile_X1Y2_FrameStrobe_O[10] ,
    \Tile_X1Y2_FrameStrobe_O[9] ,
    \Tile_X1Y2_FrameStrobe_O[8] ,
    \Tile_X1Y2_FrameStrobe_O[7] ,
    \Tile_X1Y2_FrameStrobe_O[6] ,
    \Tile_X1Y2_FrameStrobe_O[5] ,
    \Tile_X1Y2_FrameStrobe_O[4] ,
    \Tile_X1Y2_FrameStrobe_O[3] ,
    \Tile_X1Y2_FrameStrobe_O[2] ,
    \Tile_X1Y2_FrameStrobe_O[1] ,
    \Tile_X1Y2_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X1Y1_FrameStrobe_O[19] ,
    \Tile_X1Y1_FrameStrobe_O[18] ,
    \Tile_X1Y1_FrameStrobe_O[17] ,
    \Tile_X1Y1_FrameStrobe_O[16] ,
    \Tile_X1Y1_FrameStrobe_O[15] ,
    \Tile_X1Y1_FrameStrobe_O[14] ,
    \Tile_X1Y1_FrameStrobe_O[13] ,
    \Tile_X1Y1_FrameStrobe_O[12] ,
    \Tile_X1Y1_FrameStrobe_O[11] ,
    \Tile_X1Y1_FrameStrobe_O[10] ,
    \Tile_X1Y1_FrameStrobe_O[9] ,
    \Tile_X1Y1_FrameStrobe_O[8] ,
    \Tile_X1Y1_FrameStrobe_O[7] ,
    \Tile_X1Y1_FrameStrobe_O[6] ,
    \Tile_X1Y1_FrameStrobe_O[5] ,
    \Tile_X1Y1_FrameStrobe_O[4] ,
    \Tile_X1Y1_FrameStrobe_O[3] ,
    \Tile_X1Y1_FrameStrobe_O[2] ,
    \Tile_X1Y1_FrameStrobe_O[1] ,
    \Tile_X1Y1_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X1Y1_N1BEG[3] ,
    \Tile_X1Y1_N1BEG[2] ,
    \Tile_X1Y1_N1BEG[1] ,
    \Tile_X1Y1_N1BEG[0] }),
    .N1END({\Tile_X1Y2_N1BEG[3] ,
    \Tile_X1Y2_N1BEG[2] ,
    \Tile_X1Y2_N1BEG[1] ,
    \Tile_X1Y2_N1BEG[0] }),
    .N2BEG({\Tile_X1Y1_N2BEG[7] ,
    \Tile_X1Y1_N2BEG[6] ,
    \Tile_X1Y1_N2BEG[5] ,
    \Tile_X1Y1_N2BEG[4] ,
    \Tile_X1Y1_N2BEG[3] ,
    \Tile_X1Y1_N2BEG[2] ,
    \Tile_X1Y1_N2BEG[1] ,
    \Tile_X1Y1_N2BEG[0] }),
    .N2BEGb({\Tile_X1Y1_N2BEGb[7] ,
    \Tile_X1Y1_N2BEGb[6] ,
    \Tile_X1Y1_N2BEGb[5] ,
    \Tile_X1Y1_N2BEGb[4] ,
    \Tile_X1Y1_N2BEGb[3] ,
    \Tile_X1Y1_N2BEGb[2] ,
    \Tile_X1Y1_N2BEGb[1] ,
    \Tile_X1Y1_N2BEGb[0] }),
    .N2END({\Tile_X1Y2_N2BEGb[7] ,
    \Tile_X1Y2_N2BEGb[6] ,
    \Tile_X1Y2_N2BEGb[5] ,
    \Tile_X1Y2_N2BEGb[4] ,
    \Tile_X1Y2_N2BEGb[3] ,
    \Tile_X1Y2_N2BEGb[2] ,
    \Tile_X1Y2_N2BEGb[1] ,
    \Tile_X1Y2_N2BEGb[0] }),
    .N2MID({\Tile_X1Y2_N2BEG[7] ,
    \Tile_X1Y2_N2BEG[6] ,
    \Tile_X1Y2_N2BEG[5] ,
    \Tile_X1Y2_N2BEG[4] ,
    \Tile_X1Y2_N2BEG[3] ,
    \Tile_X1Y2_N2BEG[2] ,
    \Tile_X1Y2_N2BEG[1] ,
    \Tile_X1Y2_N2BEG[0] }),
    .N4BEG({\Tile_X1Y1_N4BEG[15] ,
    \Tile_X1Y1_N4BEG[14] ,
    \Tile_X1Y1_N4BEG[13] ,
    \Tile_X1Y1_N4BEG[12] ,
    \Tile_X1Y1_N4BEG[11] ,
    \Tile_X1Y1_N4BEG[10] ,
    \Tile_X1Y1_N4BEG[9] ,
    \Tile_X1Y1_N4BEG[8] ,
    \Tile_X1Y1_N4BEG[7] ,
    \Tile_X1Y1_N4BEG[6] ,
    \Tile_X1Y1_N4BEG[5] ,
    \Tile_X1Y1_N4BEG[4] ,
    \Tile_X1Y1_N4BEG[3] ,
    \Tile_X1Y1_N4BEG[2] ,
    \Tile_X1Y1_N4BEG[1] ,
    \Tile_X1Y1_N4BEG[0] }),
    .N4END({\Tile_X1Y2_N4BEG[15] ,
    \Tile_X1Y2_N4BEG[14] ,
    \Tile_X1Y2_N4BEG[13] ,
    \Tile_X1Y2_N4BEG[12] ,
    \Tile_X1Y2_N4BEG[11] ,
    \Tile_X1Y2_N4BEG[10] ,
    \Tile_X1Y2_N4BEG[9] ,
    \Tile_X1Y2_N4BEG[8] ,
    \Tile_X1Y2_N4BEG[7] ,
    \Tile_X1Y2_N4BEG[6] ,
    \Tile_X1Y2_N4BEG[5] ,
    \Tile_X1Y2_N4BEG[4] ,
    \Tile_X1Y2_N4BEG[3] ,
    \Tile_X1Y2_N4BEG[2] ,
    \Tile_X1Y2_N4BEG[1] ,
    \Tile_X1Y2_N4BEG[0] }),
    .NN4BEG({\Tile_X1Y1_NN4BEG[15] ,
    \Tile_X1Y1_NN4BEG[14] ,
    \Tile_X1Y1_NN4BEG[13] ,
    \Tile_X1Y1_NN4BEG[12] ,
    \Tile_X1Y1_NN4BEG[11] ,
    \Tile_X1Y1_NN4BEG[10] ,
    \Tile_X1Y1_NN4BEG[9] ,
    \Tile_X1Y1_NN4BEG[8] ,
    \Tile_X1Y1_NN4BEG[7] ,
    \Tile_X1Y1_NN4BEG[6] ,
    \Tile_X1Y1_NN4BEG[5] ,
    \Tile_X1Y1_NN4BEG[4] ,
    \Tile_X1Y1_NN4BEG[3] ,
    \Tile_X1Y1_NN4BEG[2] ,
    \Tile_X1Y1_NN4BEG[1] ,
    \Tile_X1Y1_NN4BEG[0] }),
    .NN4END({\Tile_X1Y2_NN4BEG[15] ,
    \Tile_X1Y2_NN4BEG[14] ,
    \Tile_X1Y2_NN4BEG[13] ,
    \Tile_X1Y2_NN4BEG[12] ,
    \Tile_X1Y2_NN4BEG[11] ,
    \Tile_X1Y2_NN4BEG[10] ,
    \Tile_X1Y2_NN4BEG[9] ,
    \Tile_X1Y2_NN4BEG[8] ,
    \Tile_X1Y2_NN4BEG[7] ,
    \Tile_X1Y2_NN4BEG[6] ,
    \Tile_X1Y2_NN4BEG[5] ,
    \Tile_X1Y2_NN4BEG[4] ,
    \Tile_X1Y2_NN4BEG[3] ,
    \Tile_X1Y2_NN4BEG[2] ,
    \Tile_X1Y2_NN4BEG[1] ,
    \Tile_X1Y2_NN4BEG[0] }),
    .S1BEG({\Tile_X1Y1_S1BEG[3] ,
    \Tile_X1Y1_S1BEG[2] ,
    \Tile_X1Y1_S1BEG[1] ,
    \Tile_X1Y1_S1BEG[0] }),
    .S1END({\Tile_X1Y0_S1BEG[3] ,
    \Tile_X1Y0_S1BEG[2] ,
    \Tile_X1Y0_S1BEG[1] ,
    \Tile_X1Y0_S1BEG[0] }),
    .S2BEG({\Tile_X1Y1_S2BEG[7] ,
    \Tile_X1Y1_S2BEG[6] ,
    \Tile_X1Y1_S2BEG[5] ,
    \Tile_X1Y1_S2BEG[4] ,
    \Tile_X1Y1_S2BEG[3] ,
    \Tile_X1Y1_S2BEG[2] ,
    \Tile_X1Y1_S2BEG[1] ,
    \Tile_X1Y1_S2BEG[0] }),
    .S2BEGb({\Tile_X1Y1_S2BEGb[7] ,
    \Tile_X1Y1_S2BEGb[6] ,
    \Tile_X1Y1_S2BEGb[5] ,
    \Tile_X1Y1_S2BEGb[4] ,
    \Tile_X1Y1_S2BEGb[3] ,
    \Tile_X1Y1_S2BEGb[2] ,
    \Tile_X1Y1_S2BEGb[1] ,
    \Tile_X1Y1_S2BEGb[0] }),
    .S2END({\Tile_X1Y0_S2BEGb[7] ,
    \Tile_X1Y0_S2BEGb[6] ,
    \Tile_X1Y0_S2BEGb[5] ,
    \Tile_X1Y0_S2BEGb[4] ,
    \Tile_X1Y0_S2BEGb[3] ,
    \Tile_X1Y0_S2BEGb[2] ,
    \Tile_X1Y0_S2BEGb[1] ,
    \Tile_X1Y0_S2BEGb[0] }),
    .S2MID({\Tile_X1Y0_S2BEG[7] ,
    \Tile_X1Y0_S2BEG[6] ,
    \Tile_X1Y0_S2BEG[5] ,
    \Tile_X1Y0_S2BEG[4] ,
    \Tile_X1Y0_S2BEG[3] ,
    \Tile_X1Y0_S2BEG[2] ,
    \Tile_X1Y0_S2BEG[1] ,
    \Tile_X1Y0_S2BEG[0] }),
    .S4BEG({\Tile_X1Y1_S4BEG[15] ,
    \Tile_X1Y1_S4BEG[14] ,
    \Tile_X1Y1_S4BEG[13] ,
    \Tile_X1Y1_S4BEG[12] ,
    \Tile_X1Y1_S4BEG[11] ,
    \Tile_X1Y1_S4BEG[10] ,
    \Tile_X1Y1_S4BEG[9] ,
    \Tile_X1Y1_S4BEG[8] ,
    \Tile_X1Y1_S4BEG[7] ,
    \Tile_X1Y1_S4BEG[6] ,
    \Tile_X1Y1_S4BEG[5] ,
    \Tile_X1Y1_S4BEG[4] ,
    \Tile_X1Y1_S4BEG[3] ,
    \Tile_X1Y1_S4BEG[2] ,
    \Tile_X1Y1_S4BEG[1] ,
    \Tile_X1Y1_S4BEG[0] }),
    .S4END({\Tile_X1Y0_S4BEG[15] ,
    \Tile_X1Y0_S4BEG[14] ,
    \Tile_X1Y0_S4BEG[13] ,
    \Tile_X1Y0_S4BEG[12] ,
    \Tile_X1Y0_S4BEG[11] ,
    \Tile_X1Y0_S4BEG[10] ,
    \Tile_X1Y0_S4BEG[9] ,
    \Tile_X1Y0_S4BEG[8] ,
    \Tile_X1Y0_S4BEG[7] ,
    \Tile_X1Y0_S4BEG[6] ,
    \Tile_X1Y0_S4BEG[5] ,
    \Tile_X1Y0_S4BEG[4] ,
    \Tile_X1Y0_S4BEG[3] ,
    \Tile_X1Y0_S4BEG[2] ,
    \Tile_X1Y0_S4BEG[1] ,
    \Tile_X1Y0_S4BEG[0] }),
    .SS4BEG({\Tile_X1Y1_SS4BEG[15] ,
    \Tile_X1Y1_SS4BEG[14] ,
    \Tile_X1Y1_SS4BEG[13] ,
    \Tile_X1Y1_SS4BEG[12] ,
    \Tile_X1Y1_SS4BEG[11] ,
    \Tile_X1Y1_SS4BEG[10] ,
    \Tile_X1Y1_SS4BEG[9] ,
    \Tile_X1Y1_SS4BEG[8] ,
    \Tile_X1Y1_SS4BEG[7] ,
    \Tile_X1Y1_SS4BEG[6] ,
    \Tile_X1Y1_SS4BEG[5] ,
    \Tile_X1Y1_SS4BEG[4] ,
    \Tile_X1Y1_SS4BEG[3] ,
    \Tile_X1Y1_SS4BEG[2] ,
    \Tile_X1Y1_SS4BEG[1] ,
    \Tile_X1Y1_SS4BEG[0] }),
    .SS4END({\Tile_X1Y0_SS4BEG[15] ,
    \Tile_X1Y0_SS4BEG[14] ,
    \Tile_X1Y0_SS4BEG[13] ,
    \Tile_X1Y0_SS4BEG[12] ,
    \Tile_X1Y0_SS4BEG[11] ,
    \Tile_X1Y0_SS4BEG[10] ,
    \Tile_X1Y0_SS4BEG[9] ,
    \Tile_X1Y0_SS4BEG[8] ,
    \Tile_X1Y0_SS4BEG[7] ,
    \Tile_X1Y0_SS4BEG[6] ,
    \Tile_X1Y0_SS4BEG[5] ,
    \Tile_X1Y0_SS4BEG[4] ,
    \Tile_X1Y0_SS4BEG[3] ,
    \Tile_X1Y0_SS4BEG[2] ,
    \Tile_X1Y0_SS4BEG[1] ,
    \Tile_X1Y0_SS4BEG[0] }),
    .W1BEG({\Tile_X1Y1_W1BEG[3] ,
    \Tile_X1Y1_W1BEG[2] ,
    \Tile_X1Y1_W1BEG[1] ,
    \Tile_X1Y1_W1BEG[0] }),
    .W1END({\Tile_X2Y1_W1BEG[3] ,
    \Tile_X2Y1_W1BEG[2] ,
    \Tile_X2Y1_W1BEG[1] ,
    \Tile_X2Y1_W1BEG[0] }),
    .W2BEG({\Tile_X1Y1_W2BEG[7] ,
    \Tile_X1Y1_W2BEG[6] ,
    \Tile_X1Y1_W2BEG[5] ,
    \Tile_X1Y1_W2BEG[4] ,
    \Tile_X1Y1_W2BEG[3] ,
    \Tile_X1Y1_W2BEG[2] ,
    \Tile_X1Y1_W2BEG[1] ,
    \Tile_X1Y1_W2BEG[0] }),
    .W2BEGb({\Tile_X1Y1_W2BEGb[7] ,
    \Tile_X1Y1_W2BEGb[6] ,
    \Tile_X1Y1_W2BEGb[5] ,
    \Tile_X1Y1_W2BEGb[4] ,
    \Tile_X1Y1_W2BEGb[3] ,
    \Tile_X1Y1_W2BEGb[2] ,
    \Tile_X1Y1_W2BEGb[1] ,
    \Tile_X1Y1_W2BEGb[0] }),
    .W2END({\Tile_X2Y1_W2BEGb[7] ,
    \Tile_X2Y1_W2BEGb[6] ,
    \Tile_X2Y1_W2BEGb[5] ,
    \Tile_X2Y1_W2BEGb[4] ,
    \Tile_X2Y1_W2BEGb[3] ,
    \Tile_X2Y1_W2BEGb[2] ,
    \Tile_X2Y1_W2BEGb[1] ,
    \Tile_X2Y1_W2BEGb[0] }),
    .W2MID({\Tile_X2Y1_W2BEG[7] ,
    \Tile_X2Y1_W2BEG[6] ,
    \Tile_X2Y1_W2BEG[5] ,
    \Tile_X2Y1_W2BEG[4] ,
    \Tile_X2Y1_W2BEG[3] ,
    \Tile_X2Y1_W2BEG[2] ,
    \Tile_X2Y1_W2BEG[1] ,
    \Tile_X2Y1_W2BEG[0] }),
    .W6BEG({\Tile_X1Y1_W6BEG[11] ,
    \Tile_X1Y1_W6BEG[10] ,
    \Tile_X1Y1_W6BEG[9] ,
    \Tile_X1Y1_W6BEG[8] ,
    \Tile_X1Y1_W6BEG[7] ,
    \Tile_X1Y1_W6BEG[6] ,
    \Tile_X1Y1_W6BEG[5] ,
    \Tile_X1Y1_W6BEG[4] ,
    \Tile_X1Y1_W6BEG[3] ,
    \Tile_X1Y1_W6BEG[2] ,
    \Tile_X1Y1_W6BEG[1] ,
    \Tile_X1Y1_W6BEG[0] }),
    .W6END({\Tile_X2Y1_W6BEG[11] ,
    \Tile_X2Y1_W6BEG[10] ,
    \Tile_X2Y1_W6BEG[9] ,
    \Tile_X2Y1_W6BEG[8] ,
    \Tile_X2Y1_W6BEG[7] ,
    \Tile_X2Y1_W6BEG[6] ,
    \Tile_X2Y1_W6BEG[5] ,
    \Tile_X2Y1_W6BEG[4] ,
    \Tile_X2Y1_W6BEG[3] ,
    \Tile_X2Y1_W6BEG[2] ,
    \Tile_X2Y1_W6BEG[1] ,
    \Tile_X2Y1_W6BEG[0] }),
    .WW4BEG({\Tile_X1Y1_WW4BEG[15] ,
    \Tile_X1Y1_WW4BEG[14] ,
    \Tile_X1Y1_WW4BEG[13] ,
    \Tile_X1Y1_WW4BEG[12] ,
    \Tile_X1Y1_WW4BEG[11] ,
    \Tile_X1Y1_WW4BEG[10] ,
    \Tile_X1Y1_WW4BEG[9] ,
    \Tile_X1Y1_WW4BEG[8] ,
    \Tile_X1Y1_WW4BEG[7] ,
    \Tile_X1Y1_WW4BEG[6] ,
    \Tile_X1Y1_WW4BEG[5] ,
    \Tile_X1Y1_WW4BEG[4] ,
    \Tile_X1Y1_WW4BEG[3] ,
    \Tile_X1Y1_WW4BEG[2] ,
    \Tile_X1Y1_WW4BEG[1] ,
    \Tile_X1Y1_WW4BEG[0] }),
    .WW4END({\Tile_X2Y1_WW4BEG[15] ,
    \Tile_X2Y1_WW4BEG[14] ,
    \Tile_X2Y1_WW4BEG[13] ,
    \Tile_X2Y1_WW4BEG[12] ,
    \Tile_X2Y1_WW4BEG[11] ,
    \Tile_X2Y1_WW4BEG[10] ,
    \Tile_X2Y1_WW4BEG[9] ,
    \Tile_X2Y1_WW4BEG[8] ,
    \Tile_X2Y1_WW4BEG[7] ,
    \Tile_X2Y1_WW4BEG[6] ,
    \Tile_X2Y1_WW4BEG[5] ,
    \Tile_X2Y1_WW4BEG[4] ,
    \Tile_X2Y1_WW4BEG[3] ,
    \Tile_X2Y1_WW4BEG[2] ,
    \Tile_X2Y1_WW4BEG[1] ,
    \Tile_X2Y1_WW4BEG[0] }));
 LUT4AB Tile_X1Y2_LUT4AB (.Ci(Tile_X1Y3_Co),
    .Co(Tile_X1Y2_Co),
    .UserCLK(Tile_X1Y3_UserCLKo),
    .UserCLKo(Tile_X1Y2_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X1Y2_E1BEG[3] ,
    \Tile_X1Y2_E1BEG[2] ,
    \Tile_X1Y2_E1BEG[1] ,
    \Tile_X1Y2_E1BEG[0] }),
    .E1END({\Tile_X0Y2_E1BEG[3] ,
    \Tile_X0Y2_E1BEG[2] ,
    \Tile_X0Y2_E1BEG[1] ,
    \Tile_X0Y2_E1BEG[0] }),
    .E2BEG({\Tile_X1Y2_E2BEG[7] ,
    \Tile_X1Y2_E2BEG[6] ,
    \Tile_X1Y2_E2BEG[5] ,
    \Tile_X1Y2_E2BEG[4] ,
    \Tile_X1Y2_E2BEG[3] ,
    \Tile_X1Y2_E2BEG[2] ,
    \Tile_X1Y2_E2BEG[1] ,
    \Tile_X1Y2_E2BEG[0] }),
    .E2BEGb({\Tile_X1Y2_E2BEGb[7] ,
    \Tile_X1Y2_E2BEGb[6] ,
    \Tile_X1Y2_E2BEGb[5] ,
    \Tile_X1Y2_E2BEGb[4] ,
    \Tile_X1Y2_E2BEGb[3] ,
    \Tile_X1Y2_E2BEGb[2] ,
    \Tile_X1Y2_E2BEGb[1] ,
    \Tile_X1Y2_E2BEGb[0] }),
    .E2END({\Tile_X0Y2_E2BEGb[7] ,
    \Tile_X0Y2_E2BEGb[6] ,
    \Tile_X0Y2_E2BEGb[5] ,
    \Tile_X0Y2_E2BEGb[4] ,
    \Tile_X0Y2_E2BEGb[3] ,
    \Tile_X0Y2_E2BEGb[2] ,
    \Tile_X0Y2_E2BEGb[1] ,
    \Tile_X0Y2_E2BEGb[0] }),
    .E2MID({\Tile_X0Y2_E2BEG[7] ,
    \Tile_X0Y2_E2BEG[6] ,
    \Tile_X0Y2_E2BEG[5] ,
    \Tile_X0Y2_E2BEG[4] ,
    \Tile_X0Y2_E2BEG[3] ,
    \Tile_X0Y2_E2BEG[2] ,
    \Tile_X0Y2_E2BEG[1] ,
    \Tile_X0Y2_E2BEG[0] }),
    .E6BEG({\Tile_X1Y2_E6BEG[11] ,
    \Tile_X1Y2_E6BEG[10] ,
    \Tile_X1Y2_E6BEG[9] ,
    \Tile_X1Y2_E6BEG[8] ,
    \Tile_X1Y2_E6BEG[7] ,
    \Tile_X1Y2_E6BEG[6] ,
    \Tile_X1Y2_E6BEG[5] ,
    \Tile_X1Y2_E6BEG[4] ,
    \Tile_X1Y2_E6BEG[3] ,
    \Tile_X1Y2_E6BEG[2] ,
    \Tile_X1Y2_E6BEG[1] ,
    \Tile_X1Y2_E6BEG[0] }),
    .E6END({\Tile_X0Y2_E6BEG[11] ,
    \Tile_X0Y2_E6BEG[10] ,
    \Tile_X0Y2_E6BEG[9] ,
    \Tile_X0Y2_E6BEG[8] ,
    \Tile_X0Y2_E6BEG[7] ,
    \Tile_X0Y2_E6BEG[6] ,
    \Tile_X0Y2_E6BEG[5] ,
    \Tile_X0Y2_E6BEG[4] ,
    \Tile_X0Y2_E6BEG[3] ,
    \Tile_X0Y2_E6BEG[2] ,
    \Tile_X0Y2_E6BEG[1] ,
    \Tile_X0Y2_E6BEG[0] }),
    .EE4BEG({\Tile_X1Y2_EE4BEG[15] ,
    \Tile_X1Y2_EE4BEG[14] ,
    \Tile_X1Y2_EE4BEG[13] ,
    \Tile_X1Y2_EE4BEG[12] ,
    \Tile_X1Y2_EE4BEG[11] ,
    \Tile_X1Y2_EE4BEG[10] ,
    \Tile_X1Y2_EE4BEG[9] ,
    \Tile_X1Y2_EE4BEG[8] ,
    \Tile_X1Y2_EE4BEG[7] ,
    \Tile_X1Y2_EE4BEG[6] ,
    \Tile_X1Y2_EE4BEG[5] ,
    \Tile_X1Y2_EE4BEG[4] ,
    \Tile_X1Y2_EE4BEG[3] ,
    \Tile_X1Y2_EE4BEG[2] ,
    \Tile_X1Y2_EE4BEG[1] ,
    \Tile_X1Y2_EE4BEG[0] }),
    .EE4END({\Tile_X0Y2_EE4BEG[15] ,
    \Tile_X0Y2_EE4BEG[14] ,
    \Tile_X0Y2_EE4BEG[13] ,
    \Tile_X0Y2_EE4BEG[12] ,
    \Tile_X0Y2_EE4BEG[11] ,
    \Tile_X0Y2_EE4BEG[10] ,
    \Tile_X0Y2_EE4BEG[9] ,
    \Tile_X0Y2_EE4BEG[8] ,
    \Tile_X0Y2_EE4BEG[7] ,
    \Tile_X0Y2_EE4BEG[6] ,
    \Tile_X0Y2_EE4BEG[5] ,
    \Tile_X0Y2_EE4BEG[4] ,
    \Tile_X0Y2_EE4BEG[3] ,
    \Tile_X0Y2_EE4BEG[2] ,
    \Tile_X0Y2_EE4BEG[1] ,
    \Tile_X0Y2_EE4BEG[0] }),
    .FrameData({\Tile_X0Y2_FrameData_O[31] ,
    \Tile_X0Y2_FrameData_O[30] ,
    \Tile_X0Y2_FrameData_O[29] ,
    \Tile_X0Y2_FrameData_O[28] ,
    \Tile_X0Y2_FrameData_O[27] ,
    \Tile_X0Y2_FrameData_O[26] ,
    \Tile_X0Y2_FrameData_O[25] ,
    \Tile_X0Y2_FrameData_O[24] ,
    \Tile_X0Y2_FrameData_O[23] ,
    \Tile_X0Y2_FrameData_O[22] ,
    \Tile_X0Y2_FrameData_O[21] ,
    \Tile_X0Y2_FrameData_O[20] ,
    \Tile_X0Y2_FrameData_O[19] ,
    \Tile_X0Y2_FrameData_O[18] ,
    \Tile_X0Y2_FrameData_O[17] ,
    \Tile_X0Y2_FrameData_O[16] ,
    \Tile_X0Y2_FrameData_O[15] ,
    \Tile_X0Y2_FrameData_O[14] ,
    \Tile_X0Y2_FrameData_O[13] ,
    \Tile_X0Y2_FrameData_O[12] ,
    \Tile_X0Y2_FrameData_O[11] ,
    \Tile_X0Y2_FrameData_O[10] ,
    \Tile_X0Y2_FrameData_O[9] ,
    \Tile_X0Y2_FrameData_O[8] ,
    \Tile_X0Y2_FrameData_O[7] ,
    \Tile_X0Y2_FrameData_O[6] ,
    \Tile_X0Y2_FrameData_O[5] ,
    \Tile_X0Y2_FrameData_O[4] ,
    \Tile_X0Y2_FrameData_O[3] ,
    \Tile_X0Y2_FrameData_O[2] ,
    \Tile_X0Y2_FrameData_O[1] ,
    \Tile_X0Y2_FrameData_O[0] }),
    .FrameData_O({\Tile_X1Y2_FrameData_O[31] ,
    \Tile_X1Y2_FrameData_O[30] ,
    \Tile_X1Y2_FrameData_O[29] ,
    \Tile_X1Y2_FrameData_O[28] ,
    \Tile_X1Y2_FrameData_O[27] ,
    \Tile_X1Y2_FrameData_O[26] ,
    \Tile_X1Y2_FrameData_O[25] ,
    \Tile_X1Y2_FrameData_O[24] ,
    \Tile_X1Y2_FrameData_O[23] ,
    \Tile_X1Y2_FrameData_O[22] ,
    \Tile_X1Y2_FrameData_O[21] ,
    \Tile_X1Y2_FrameData_O[20] ,
    \Tile_X1Y2_FrameData_O[19] ,
    \Tile_X1Y2_FrameData_O[18] ,
    \Tile_X1Y2_FrameData_O[17] ,
    \Tile_X1Y2_FrameData_O[16] ,
    \Tile_X1Y2_FrameData_O[15] ,
    \Tile_X1Y2_FrameData_O[14] ,
    \Tile_X1Y2_FrameData_O[13] ,
    \Tile_X1Y2_FrameData_O[12] ,
    \Tile_X1Y2_FrameData_O[11] ,
    \Tile_X1Y2_FrameData_O[10] ,
    \Tile_X1Y2_FrameData_O[9] ,
    \Tile_X1Y2_FrameData_O[8] ,
    \Tile_X1Y2_FrameData_O[7] ,
    \Tile_X1Y2_FrameData_O[6] ,
    \Tile_X1Y2_FrameData_O[5] ,
    \Tile_X1Y2_FrameData_O[4] ,
    \Tile_X1Y2_FrameData_O[3] ,
    \Tile_X1Y2_FrameData_O[2] ,
    \Tile_X1Y2_FrameData_O[1] ,
    \Tile_X1Y2_FrameData_O[0] }),
    .FrameStrobe({\Tile_X1Y3_FrameStrobe_O[19] ,
    \Tile_X1Y3_FrameStrobe_O[18] ,
    \Tile_X1Y3_FrameStrobe_O[17] ,
    \Tile_X1Y3_FrameStrobe_O[16] ,
    \Tile_X1Y3_FrameStrobe_O[15] ,
    \Tile_X1Y3_FrameStrobe_O[14] ,
    \Tile_X1Y3_FrameStrobe_O[13] ,
    \Tile_X1Y3_FrameStrobe_O[12] ,
    \Tile_X1Y3_FrameStrobe_O[11] ,
    \Tile_X1Y3_FrameStrobe_O[10] ,
    \Tile_X1Y3_FrameStrobe_O[9] ,
    \Tile_X1Y3_FrameStrobe_O[8] ,
    \Tile_X1Y3_FrameStrobe_O[7] ,
    \Tile_X1Y3_FrameStrobe_O[6] ,
    \Tile_X1Y3_FrameStrobe_O[5] ,
    \Tile_X1Y3_FrameStrobe_O[4] ,
    \Tile_X1Y3_FrameStrobe_O[3] ,
    \Tile_X1Y3_FrameStrobe_O[2] ,
    \Tile_X1Y3_FrameStrobe_O[1] ,
    \Tile_X1Y3_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X1Y2_FrameStrobe_O[19] ,
    \Tile_X1Y2_FrameStrobe_O[18] ,
    \Tile_X1Y2_FrameStrobe_O[17] ,
    \Tile_X1Y2_FrameStrobe_O[16] ,
    \Tile_X1Y2_FrameStrobe_O[15] ,
    \Tile_X1Y2_FrameStrobe_O[14] ,
    \Tile_X1Y2_FrameStrobe_O[13] ,
    \Tile_X1Y2_FrameStrobe_O[12] ,
    \Tile_X1Y2_FrameStrobe_O[11] ,
    \Tile_X1Y2_FrameStrobe_O[10] ,
    \Tile_X1Y2_FrameStrobe_O[9] ,
    \Tile_X1Y2_FrameStrobe_O[8] ,
    \Tile_X1Y2_FrameStrobe_O[7] ,
    \Tile_X1Y2_FrameStrobe_O[6] ,
    \Tile_X1Y2_FrameStrobe_O[5] ,
    \Tile_X1Y2_FrameStrobe_O[4] ,
    \Tile_X1Y2_FrameStrobe_O[3] ,
    \Tile_X1Y2_FrameStrobe_O[2] ,
    \Tile_X1Y2_FrameStrobe_O[1] ,
    \Tile_X1Y2_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X1Y2_N1BEG[3] ,
    \Tile_X1Y2_N1BEG[2] ,
    \Tile_X1Y2_N1BEG[1] ,
    \Tile_X1Y2_N1BEG[0] }),
    .N1END({\Tile_X1Y3_N1BEG[3] ,
    \Tile_X1Y3_N1BEG[2] ,
    \Tile_X1Y3_N1BEG[1] ,
    \Tile_X1Y3_N1BEG[0] }),
    .N2BEG({\Tile_X1Y2_N2BEG[7] ,
    \Tile_X1Y2_N2BEG[6] ,
    \Tile_X1Y2_N2BEG[5] ,
    \Tile_X1Y2_N2BEG[4] ,
    \Tile_X1Y2_N2BEG[3] ,
    \Tile_X1Y2_N2BEG[2] ,
    \Tile_X1Y2_N2BEG[1] ,
    \Tile_X1Y2_N2BEG[0] }),
    .N2BEGb({\Tile_X1Y2_N2BEGb[7] ,
    \Tile_X1Y2_N2BEGb[6] ,
    \Tile_X1Y2_N2BEGb[5] ,
    \Tile_X1Y2_N2BEGb[4] ,
    \Tile_X1Y2_N2BEGb[3] ,
    \Tile_X1Y2_N2BEGb[2] ,
    \Tile_X1Y2_N2BEGb[1] ,
    \Tile_X1Y2_N2BEGb[0] }),
    .N2END({\Tile_X1Y3_N2BEGb[7] ,
    \Tile_X1Y3_N2BEGb[6] ,
    \Tile_X1Y3_N2BEGb[5] ,
    \Tile_X1Y3_N2BEGb[4] ,
    \Tile_X1Y3_N2BEGb[3] ,
    \Tile_X1Y3_N2BEGb[2] ,
    \Tile_X1Y3_N2BEGb[1] ,
    \Tile_X1Y3_N2BEGb[0] }),
    .N2MID({\Tile_X1Y3_N2BEG[7] ,
    \Tile_X1Y3_N2BEG[6] ,
    \Tile_X1Y3_N2BEG[5] ,
    \Tile_X1Y3_N2BEG[4] ,
    \Tile_X1Y3_N2BEG[3] ,
    \Tile_X1Y3_N2BEG[2] ,
    \Tile_X1Y3_N2BEG[1] ,
    \Tile_X1Y3_N2BEG[0] }),
    .N4BEG({\Tile_X1Y2_N4BEG[15] ,
    \Tile_X1Y2_N4BEG[14] ,
    \Tile_X1Y2_N4BEG[13] ,
    \Tile_X1Y2_N4BEG[12] ,
    \Tile_X1Y2_N4BEG[11] ,
    \Tile_X1Y2_N4BEG[10] ,
    \Tile_X1Y2_N4BEG[9] ,
    \Tile_X1Y2_N4BEG[8] ,
    \Tile_X1Y2_N4BEG[7] ,
    \Tile_X1Y2_N4BEG[6] ,
    \Tile_X1Y2_N4BEG[5] ,
    \Tile_X1Y2_N4BEG[4] ,
    \Tile_X1Y2_N4BEG[3] ,
    \Tile_X1Y2_N4BEG[2] ,
    \Tile_X1Y2_N4BEG[1] ,
    \Tile_X1Y2_N4BEG[0] }),
    .N4END({\Tile_X1Y3_N4BEG[15] ,
    \Tile_X1Y3_N4BEG[14] ,
    \Tile_X1Y3_N4BEG[13] ,
    \Tile_X1Y3_N4BEG[12] ,
    \Tile_X1Y3_N4BEG[11] ,
    \Tile_X1Y3_N4BEG[10] ,
    \Tile_X1Y3_N4BEG[9] ,
    \Tile_X1Y3_N4BEG[8] ,
    \Tile_X1Y3_N4BEG[7] ,
    \Tile_X1Y3_N4BEG[6] ,
    \Tile_X1Y3_N4BEG[5] ,
    \Tile_X1Y3_N4BEG[4] ,
    \Tile_X1Y3_N4BEG[3] ,
    \Tile_X1Y3_N4BEG[2] ,
    \Tile_X1Y3_N4BEG[1] ,
    \Tile_X1Y3_N4BEG[0] }),
    .NN4BEG({\Tile_X1Y2_NN4BEG[15] ,
    \Tile_X1Y2_NN4BEG[14] ,
    \Tile_X1Y2_NN4BEG[13] ,
    \Tile_X1Y2_NN4BEG[12] ,
    \Tile_X1Y2_NN4BEG[11] ,
    \Tile_X1Y2_NN4BEG[10] ,
    \Tile_X1Y2_NN4BEG[9] ,
    \Tile_X1Y2_NN4BEG[8] ,
    \Tile_X1Y2_NN4BEG[7] ,
    \Tile_X1Y2_NN4BEG[6] ,
    \Tile_X1Y2_NN4BEG[5] ,
    \Tile_X1Y2_NN4BEG[4] ,
    \Tile_X1Y2_NN4BEG[3] ,
    \Tile_X1Y2_NN4BEG[2] ,
    \Tile_X1Y2_NN4BEG[1] ,
    \Tile_X1Y2_NN4BEG[0] }),
    .NN4END({\Tile_X1Y3_NN4BEG[15] ,
    \Tile_X1Y3_NN4BEG[14] ,
    \Tile_X1Y3_NN4BEG[13] ,
    \Tile_X1Y3_NN4BEG[12] ,
    \Tile_X1Y3_NN4BEG[11] ,
    \Tile_X1Y3_NN4BEG[10] ,
    \Tile_X1Y3_NN4BEG[9] ,
    \Tile_X1Y3_NN4BEG[8] ,
    \Tile_X1Y3_NN4BEG[7] ,
    \Tile_X1Y3_NN4BEG[6] ,
    \Tile_X1Y3_NN4BEG[5] ,
    \Tile_X1Y3_NN4BEG[4] ,
    \Tile_X1Y3_NN4BEG[3] ,
    \Tile_X1Y3_NN4BEG[2] ,
    \Tile_X1Y3_NN4BEG[1] ,
    \Tile_X1Y3_NN4BEG[0] }),
    .S1BEG({\Tile_X1Y2_S1BEG[3] ,
    \Tile_X1Y2_S1BEG[2] ,
    \Tile_X1Y2_S1BEG[1] ,
    \Tile_X1Y2_S1BEG[0] }),
    .S1END({\Tile_X1Y1_S1BEG[3] ,
    \Tile_X1Y1_S1BEG[2] ,
    \Tile_X1Y1_S1BEG[1] ,
    \Tile_X1Y1_S1BEG[0] }),
    .S2BEG({\Tile_X1Y2_S2BEG[7] ,
    \Tile_X1Y2_S2BEG[6] ,
    \Tile_X1Y2_S2BEG[5] ,
    \Tile_X1Y2_S2BEG[4] ,
    \Tile_X1Y2_S2BEG[3] ,
    \Tile_X1Y2_S2BEG[2] ,
    \Tile_X1Y2_S2BEG[1] ,
    \Tile_X1Y2_S2BEG[0] }),
    .S2BEGb({\Tile_X1Y2_S2BEGb[7] ,
    \Tile_X1Y2_S2BEGb[6] ,
    \Tile_X1Y2_S2BEGb[5] ,
    \Tile_X1Y2_S2BEGb[4] ,
    \Tile_X1Y2_S2BEGb[3] ,
    \Tile_X1Y2_S2BEGb[2] ,
    \Tile_X1Y2_S2BEGb[1] ,
    \Tile_X1Y2_S2BEGb[0] }),
    .S2END({\Tile_X1Y1_S2BEGb[7] ,
    \Tile_X1Y1_S2BEGb[6] ,
    \Tile_X1Y1_S2BEGb[5] ,
    \Tile_X1Y1_S2BEGb[4] ,
    \Tile_X1Y1_S2BEGb[3] ,
    \Tile_X1Y1_S2BEGb[2] ,
    \Tile_X1Y1_S2BEGb[1] ,
    \Tile_X1Y1_S2BEGb[0] }),
    .S2MID({\Tile_X1Y1_S2BEG[7] ,
    \Tile_X1Y1_S2BEG[6] ,
    \Tile_X1Y1_S2BEG[5] ,
    \Tile_X1Y1_S2BEG[4] ,
    \Tile_X1Y1_S2BEG[3] ,
    \Tile_X1Y1_S2BEG[2] ,
    \Tile_X1Y1_S2BEG[1] ,
    \Tile_X1Y1_S2BEG[0] }),
    .S4BEG({\Tile_X1Y2_S4BEG[15] ,
    \Tile_X1Y2_S4BEG[14] ,
    \Tile_X1Y2_S4BEG[13] ,
    \Tile_X1Y2_S4BEG[12] ,
    \Tile_X1Y2_S4BEG[11] ,
    \Tile_X1Y2_S4BEG[10] ,
    \Tile_X1Y2_S4BEG[9] ,
    \Tile_X1Y2_S4BEG[8] ,
    \Tile_X1Y2_S4BEG[7] ,
    \Tile_X1Y2_S4BEG[6] ,
    \Tile_X1Y2_S4BEG[5] ,
    \Tile_X1Y2_S4BEG[4] ,
    \Tile_X1Y2_S4BEG[3] ,
    \Tile_X1Y2_S4BEG[2] ,
    \Tile_X1Y2_S4BEG[1] ,
    \Tile_X1Y2_S4BEG[0] }),
    .S4END({\Tile_X1Y1_S4BEG[15] ,
    \Tile_X1Y1_S4BEG[14] ,
    \Tile_X1Y1_S4BEG[13] ,
    \Tile_X1Y1_S4BEG[12] ,
    \Tile_X1Y1_S4BEG[11] ,
    \Tile_X1Y1_S4BEG[10] ,
    \Tile_X1Y1_S4BEG[9] ,
    \Tile_X1Y1_S4BEG[8] ,
    \Tile_X1Y1_S4BEG[7] ,
    \Tile_X1Y1_S4BEG[6] ,
    \Tile_X1Y1_S4BEG[5] ,
    \Tile_X1Y1_S4BEG[4] ,
    \Tile_X1Y1_S4BEG[3] ,
    \Tile_X1Y1_S4BEG[2] ,
    \Tile_X1Y1_S4BEG[1] ,
    \Tile_X1Y1_S4BEG[0] }),
    .SS4BEG({\Tile_X1Y2_SS4BEG[15] ,
    \Tile_X1Y2_SS4BEG[14] ,
    \Tile_X1Y2_SS4BEG[13] ,
    \Tile_X1Y2_SS4BEG[12] ,
    \Tile_X1Y2_SS4BEG[11] ,
    \Tile_X1Y2_SS4BEG[10] ,
    \Tile_X1Y2_SS4BEG[9] ,
    \Tile_X1Y2_SS4BEG[8] ,
    \Tile_X1Y2_SS4BEG[7] ,
    \Tile_X1Y2_SS4BEG[6] ,
    \Tile_X1Y2_SS4BEG[5] ,
    \Tile_X1Y2_SS4BEG[4] ,
    \Tile_X1Y2_SS4BEG[3] ,
    \Tile_X1Y2_SS4BEG[2] ,
    \Tile_X1Y2_SS4BEG[1] ,
    \Tile_X1Y2_SS4BEG[0] }),
    .SS4END({\Tile_X1Y1_SS4BEG[15] ,
    \Tile_X1Y1_SS4BEG[14] ,
    \Tile_X1Y1_SS4BEG[13] ,
    \Tile_X1Y1_SS4BEG[12] ,
    \Tile_X1Y1_SS4BEG[11] ,
    \Tile_X1Y1_SS4BEG[10] ,
    \Tile_X1Y1_SS4BEG[9] ,
    \Tile_X1Y1_SS4BEG[8] ,
    \Tile_X1Y1_SS4BEG[7] ,
    \Tile_X1Y1_SS4BEG[6] ,
    \Tile_X1Y1_SS4BEG[5] ,
    \Tile_X1Y1_SS4BEG[4] ,
    \Tile_X1Y1_SS4BEG[3] ,
    \Tile_X1Y1_SS4BEG[2] ,
    \Tile_X1Y1_SS4BEG[1] ,
    \Tile_X1Y1_SS4BEG[0] }),
    .W1BEG({\Tile_X1Y2_W1BEG[3] ,
    \Tile_X1Y2_W1BEG[2] ,
    \Tile_X1Y2_W1BEG[1] ,
    \Tile_X1Y2_W1BEG[0] }),
    .W1END({\Tile_X2Y2_W1BEG[3] ,
    \Tile_X2Y2_W1BEG[2] ,
    \Tile_X2Y2_W1BEG[1] ,
    \Tile_X2Y2_W1BEG[0] }),
    .W2BEG({\Tile_X1Y2_W2BEG[7] ,
    \Tile_X1Y2_W2BEG[6] ,
    \Tile_X1Y2_W2BEG[5] ,
    \Tile_X1Y2_W2BEG[4] ,
    \Tile_X1Y2_W2BEG[3] ,
    \Tile_X1Y2_W2BEG[2] ,
    \Tile_X1Y2_W2BEG[1] ,
    \Tile_X1Y2_W2BEG[0] }),
    .W2BEGb({\Tile_X1Y2_W2BEGb[7] ,
    \Tile_X1Y2_W2BEGb[6] ,
    \Tile_X1Y2_W2BEGb[5] ,
    \Tile_X1Y2_W2BEGb[4] ,
    \Tile_X1Y2_W2BEGb[3] ,
    \Tile_X1Y2_W2BEGb[2] ,
    \Tile_X1Y2_W2BEGb[1] ,
    \Tile_X1Y2_W2BEGb[0] }),
    .W2END({\Tile_X2Y2_W2BEGb[7] ,
    \Tile_X2Y2_W2BEGb[6] ,
    \Tile_X2Y2_W2BEGb[5] ,
    \Tile_X2Y2_W2BEGb[4] ,
    \Tile_X2Y2_W2BEGb[3] ,
    \Tile_X2Y2_W2BEGb[2] ,
    \Tile_X2Y2_W2BEGb[1] ,
    \Tile_X2Y2_W2BEGb[0] }),
    .W2MID({\Tile_X2Y2_W2BEG[7] ,
    \Tile_X2Y2_W2BEG[6] ,
    \Tile_X2Y2_W2BEG[5] ,
    \Tile_X2Y2_W2BEG[4] ,
    \Tile_X2Y2_W2BEG[3] ,
    \Tile_X2Y2_W2BEG[2] ,
    \Tile_X2Y2_W2BEG[1] ,
    \Tile_X2Y2_W2BEG[0] }),
    .W6BEG({\Tile_X1Y2_W6BEG[11] ,
    \Tile_X1Y2_W6BEG[10] ,
    \Tile_X1Y2_W6BEG[9] ,
    \Tile_X1Y2_W6BEG[8] ,
    \Tile_X1Y2_W6BEG[7] ,
    \Tile_X1Y2_W6BEG[6] ,
    \Tile_X1Y2_W6BEG[5] ,
    \Tile_X1Y2_W6BEG[4] ,
    \Tile_X1Y2_W6BEG[3] ,
    \Tile_X1Y2_W6BEG[2] ,
    \Tile_X1Y2_W6BEG[1] ,
    \Tile_X1Y2_W6BEG[0] }),
    .W6END({\Tile_X2Y2_W6BEG[11] ,
    \Tile_X2Y2_W6BEG[10] ,
    \Tile_X2Y2_W6BEG[9] ,
    \Tile_X2Y2_W6BEG[8] ,
    \Tile_X2Y2_W6BEG[7] ,
    \Tile_X2Y2_W6BEG[6] ,
    \Tile_X2Y2_W6BEG[5] ,
    \Tile_X2Y2_W6BEG[4] ,
    \Tile_X2Y2_W6BEG[3] ,
    \Tile_X2Y2_W6BEG[2] ,
    \Tile_X2Y2_W6BEG[1] ,
    \Tile_X2Y2_W6BEG[0] }),
    .WW4BEG({\Tile_X1Y2_WW4BEG[15] ,
    \Tile_X1Y2_WW4BEG[14] ,
    \Tile_X1Y2_WW4BEG[13] ,
    \Tile_X1Y2_WW4BEG[12] ,
    \Tile_X1Y2_WW4BEG[11] ,
    \Tile_X1Y2_WW4BEG[10] ,
    \Tile_X1Y2_WW4BEG[9] ,
    \Tile_X1Y2_WW4BEG[8] ,
    \Tile_X1Y2_WW4BEG[7] ,
    \Tile_X1Y2_WW4BEG[6] ,
    \Tile_X1Y2_WW4BEG[5] ,
    \Tile_X1Y2_WW4BEG[4] ,
    \Tile_X1Y2_WW4BEG[3] ,
    \Tile_X1Y2_WW4BEG[2] ,
    \Tile_X1Y2_WW4BEG[1] ,
    \Tile_X1Y2_WW4BEG[0] }),
    .WW4END({\Tile_X2Y2_WW4BEG[15] ,
    \Tile_X2Y2_WW4BEG[14] ,
    \Tile_X2Y2_WW4BEG[13] ,
    \Tile_X2Y2_WW4BEG[12] ,
    \Tile_X2Y2_WW4BEG[11] ,
    \Tile_X2Y2_WW4BEG[10] ,
    \Tile_X2Y2_WW4BEG[9] ,
    \Tile_X2Y2_WW4BEG[8] ,
    \Tile_X2Y2_WW4BEG[7] ,
    \Tile_X2Y2_WW4BEG[6] ,
    \Tile_X2Y2_WW4BEG[5] ,
    \Tile_X2Y2_WW4BEG[4] ,
    \Tile_X2Y2_WW4BEG[3] ,
    \Tile_X2Y2_WW4BEG[2] ,
    \Tile_X2Y2_WW4BEG[1] ,
    \Tile_X2Y2_WW4BEG[0] }));
 LUT4AB Tile_X1Y3_LUT4AB (.Ci(Tile_X1Y4_Co),
    .Co(Tile_X1Y3_Co),
    .UserCLK(Tile_X1Y4_UserCLKo),
    .UserCLKo(Tile_X1Y3_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X1Y3_E1BEG[3] ,
    \Tile_X1Y3_E1BEG[2] ,
    \Tile_X1Y3_E1BEG[1] ,
    \Tile_X1Y3_E1BEG[0] }),
    .E1END({\Tile_X0Y3_E1BEG[3] ,
    \Tile_X0Y3_E1BEG[2] ,
    \Tile_X0Y3_E1BEG[1] ,
    \Tile_X0Y3_E1BEG[0] }),
    .E2BEG({\Tile_X1Y3_E2BEG[7] ,
    \Tile_X1Y3_E2BEG[6] ,
    \Tile_X1Y3_E2BEG[5] ,
    \Tile_X1Y3_E2BEG[4] ,
    \Tile_X1Y3_E2BEG[3] ,
    \Tile_X1Y3_E2BEG[2] ,
    \Tile_X1Y3_E2BEG[1] ,
    \Tile_X1Y3_E2BEG[0] }),
    .E2BEGb({\Tile_X1Y3_E2BEGb[7] ,
    \Tile_X1Y3_E2BEGb[6] ,
    \Tile_X1Y3_E2BEGb[5] ,
    \Tile_X1Y3_E2BEGb[4] ,
    \Tile_X1Y3_E2BEGb[3] ,
    \Tile_X1Y3_E2BEGb[2] ,
    \Tile_X1Y3_E2BEGb[1] ,
    \Tile_X1Y3_E2BEGb[0] }),
    .E2END({\Tile_X0Y3_E2BEGb[7] ,
    \Tile_X0Y3_E2BEGb[6] ,
    \Tile_X0Y3_E2BEGb[5] ,
    \Tile_X0Y3_E2BEGb[4] ,
    \Tile_X0Y3_E2BEGb[3] ,
    \Tile_X0Y3_E2BEGb[2] ,
    \Tile_X0Y3_E2BEGb[1] ,
    \Tile_X0Y3_E2BEGb[0] }),
    .E2MID({\Tile_X0Y3_E2BEG[7] ,
    \Tile_X0Y3_E2BEG[6] ,
    \Tile_X0Y3_E2BEG[5] ,
    \Tile_X0Y3_E2BEG[4] ,
    \Tile_X0Y3_E2BEG[3] ,
    \Tile_X0Y3_E2BEG[2] ,
    \Tile_X0Y3_E2BEG[1] ,
    \Tile_X0Y3_E2BEG[0] }),
    .E6BEG({\Tile_X1Y3_E6BEG[11] ,
    \Tile_X1Y3_E6BEG[10] ,
    \Tile_X1Y3_E6BEG[9] ,
    \Tile_X1Y3_E6BEG[8] ,
    \Tile_X1Y3_E6BEG[7] ,
    \Tile_X1Y3_E6BEG[6] ,
    \Tile_X1Y3_E6BEG[5] ,
    \Tile_X1Y3_E6BEG[4] ,
    \Tile_X1Y3_E6BEG[3] ,
    \Tile_X1Y3_E6BEG[2] ,
    \Tile_X1Y3_E6BEG[1] ,
    \Tile_X1Y3_E6BEG[0] }),
    .E6END({\Tile_X0Y3_E6BEG[11] ,
    \Tile_X0Y3_E6BEG[10] ,
    \Tile_X0Y3_E6BEG[9] ,
    \Tile_X0Y3_E6BEG[8] ,
    \Tile_X0Y3_E6BEG[7] ,
    \Tile_X0Y3_E6BEG[6] ,
    \Tile_X0Y3_E6BEG[5] ,
    \Tile_X0Y3_E6BEG[4] ,
    \Tile_X0Y3_E6BEG[3] ,
    \Tile_X0Y3_E6BEG[2] ,
    \Tile_X0Y3_E6BEG[1] ,
    \Tile_X0Y3_E6BEG[0] }),
    .EE4BEG({\Tile_X1Y3_EE4BEG[15] ,
    \Tile_X1Y3_EE4BEG[14] ,
    \Tile_X1Y3_EE4BEG[13] ,
    \Tile_X1Y3_EE4BEG[12] ,
    \Tile_X1Y3_EE4BEG[11] ,
    \Tile_X1Y3_EE4BEG[10] ,
    \Tile_X1Y3_EE4BEG[9] ,
    \Tile_X1Y3_EE4BEG[8] ,
    \Tile_X1Y3_EE4BEG[7] ,
    \Tile_X1Y3_EE4BEG[6] ,
    \Tile_X1Y3_EE4BEG[5] ,
    \Tile_X1Y3_EE4BEG[4] ,
    \Tile_X1Y3_EE4BEG[3] ,
    \Tile_X1Y3_EE4BEG[2] ,
    \Tile_X1Y3_EE4BEG[1] ,
    \Tile_X1Y3_EE4BEG[0] }),
    .EE4END({\Tile_X0Y3_EE4BEG[15] ,
    \Tile_X0Y3_EE4BEG[14] ,
    \Tile_X0Y3_EE4BEG[13] ,
    \Tile_X0Y3_EE4BEG[12] ,
    \Tile_X0Y3_EE4BEG[11] ,
    \Tile_X0Y3_EE4BEG[10] ,
    \Tile_X0Y3_EE4BEG[9] ,
    \Tile_X0Y3_EE4BEG[8] ,
    \Tile_X0Y3_EE4BEG[7] ,
    \Tile_X0Y3_EE4BEG[6] ,
    \Tile_X0Y3_EE4BEG[5] ,
    \Tile_X0Y3_EE4BEG[4] ,
    \Tile_X0Y3_EE4BEG[3] ,
    \Tile_X0Y3_EE4BEG[2] ,
    \Tile_X0Y3_EE4BEG[1] ,
    \Tile_X0Y3_EE4BEG[0] }),
    .FrameData({\Tile_X0Y3_FrameData_O[31] ,
    \Tile_X0Y3_FrameData_O[30] ,
    \Tile_X0Y3_FrameData_O[29] ,
    \Tile_X0Y3_FrameData_O[28] ,
    \Tile_X0Y3_FrameData_O[27] ,
    \Tile_X0Y3_FrameData_O[26] ,
    \Tile_X0Y3_FrameData_O[25] ,
    \Tile_X0Y3_FrameData_O[24] ,
    \Tile_X0Y3_FrameData_O[23] ,
    \Tile_X0Y3_FrameData_O[22] ,
    \Tile_X0Y3_FrameData_O[21] ,
    \Tile_X0Y3_FrameData_O[20] ,
    \Tile_X0Y3_FrameData_O[19] ,
    \Tile_X0Y3_FrameData_O[18] ,
    \Tile_X0Y3_FrameData_O[17] ,
    \Tile_X0Y3_FrameData_O[16] ,
    \Tile_X0Y3_FrameData_O[15] ,
    \Tile_X0Y3_FrameData_O[14] ,
    \Tile_X0Y3_FrameData_O[13] ,
    \Tile_X0Y3_FrameData_O[12] ,
    \Tile_X0Y3_FrameData_O[11] ,
    \Tile_X0Y3_FrameData_O[10] ,
    \Tile_X0Y3_FrameData_O[9] ,
    \Tile_X0Y3_FrameData_O[8] ,
    \Tile_X0Y3_FrameData_O[7] ,
    \Tile_X0Y3_FrameData_O[6] ,
    \Tile_X0Y3_FrameData_O[5] ,
    \Tile_X0Y3_FrameData_O[4] ,
    \Tile_X0Y3_FrameData_O[3] ,
    \Tile_X0Y3_FrameData_O[2] ,
    \Tile_X0Y3_FrameData_O[1] ,
    \Tile_X0Y3_FrameData_O[0] }),
    .FrameData_O({\Tile_X1Y3_FrameData_O[31] ,
    \Tile_X1Y3_FrameData_O[30] ,
    \Tile_X1Y3_FrameData_O[29] ,
    \Tile_X1Y3_FrameData_O[28] ,
    \Tile_X1Y3_FrameData_O[27] ,
    \Tile_X1Y3_FrameData_O[26] ,
    \Tile_X1Y3_FrameData_O[25] ,
    \Tile_X1Y3_FrameData_O[24] ,
    \Tile_X1Y3_FrameData_O[23] ,
    \Tile_X1Y3_FrameData_O[22] ,
    \Tile_X1Y3_FrameData_O[21] ,
    \Tile_X1Y3_FrameData_O[20] ,
    \Tile_X1Y3_FrameData_O[19] ,
    \Tile_X1Y3_FrameData_O[18] ,
    \Tile_X1Y3_FrameData_O[17] ,
    \Tile_X1Y3_FrameData_O[16] ,
    \Tile_X1Y3_FrameData_O[15] ,
    \Tile_X1Y3_FrameData_O[14] ,
    \Tile_X1Y3_FrameData_O[13] ,
    \Tile_X1Y3_FrameData_O[12] ,
    \Tile_X1Y3_FrameData_O[11] ,
    \Tile_X1Y3_FrameData_O[10] ,
    \Tile_X1Y3_FrameData_O[9] ,
    \Tile_X1Y3_FrameData_O[8] ,
    \Tile_X1Y3_FrameData_O[7] ,
    \Tile_X1Y3_FrameData_O[6] ,
    \Tile_X1Y3_FrameData_O[5] ,
    \Tile_X1Y3_FrameData_O[4] ,
    \Tile_X1Y3_FrameData_O[3] ,
    \Tile_X1Y3_FrameData_O[2] ,
    \Tile_X1Y3_FrameData_O[1] ,
    \Tile_X1Y3_FrameData_O[0] }),
    .FrameStrobe({\Tile_X1Y4_FrameStrobe_O[19] ,
    \Tile_X1Y4_FrameStrobe_O[18] ,
    \Tile_X1Y4_FrameStrobe_O[17] ,
    \Tile_X1Y4_FrameStrobe_O[16] ,
    \Tile_X1Y4_FrameStrobe_O[15] ,
    \Tile_X1Y4_FrameStrobe_O[14] ,
    \Tile_X1Y4_FrameStrobe_O[13] ,
    \Tile_X1Y4_FrameStrobe_O[12] ,
    \Tile_X1Y4_FrameStrobe_O[11] ,
    \Tile_X1Y4_FrameStrobe_O[10] ,
    \Tile_X1Y4_FrameStrobe_O[9] ,
    \Tile_X1Y4_FrameStrobe_O[8] ,
    \Tile_X1Y4_FrameStrobe_O[7] ,
    \Tile_X1Y4_FrameStrobe_O[6] ,
    \Tile_X1Y4_FrameStrobe_O[5] ,
    \Tile_X1Y4_FrameStrobe_O[4] ,
    \Tile_X1Y4_FrameStrobe_O[3] ,
    \Tile_X1Y4_FrameStrobe_O[2] ,
    \Tile_X1Y4_FrameStrobe_O[1] ,
    \Tile_X1Y4_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X1Y3_FrameStrobe_O[19] ,
    \Tile_X1Y3_FrameStrobe_O[18] ,
    \Tile_X1Y3_FrameStrobe_O[17] ,
    \Tile_X1Y3_FrameStrobe_O[16] ,
    \Tile_X1Y3_FrameStrobe_O[15] ,
    \Tile_X1Y3_FrameStrobe_O[14] ,
    \Tile_X1Y3_FrameStrobe_O[13] ,
    \Tile_X1Y3_FrameStrobe_O[12] ,
    \Tile_X1Y3_FrameStrobe_O[11] ,
    \Tile_X1Y3_FrameStrobe_O[10] ,
    \Tile_X1Y3_FrameStrobe_O[9] ,
    \Tile_X1Y3_FrameStrobe_O[8] ,
    \Tile_X1Y3_FrameStrobe_O[7] ,
    \Tile_X1Y3_FrameStrobe_O[6] ,
    \Tile_X1Y3_FrameStrobe_O[5] ,
    \Tile_X1Y3_FrameStrobe_O[4] ,
    \Tile_X1Y3_FrameStrobe_O[3] ,
    \Tile_X1Y3_FrameStrobe_O[2] ,
    \Tile_X1Y3_FrameStrobe_O[1] ,
    \Tile_X1Y3_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X1Y3_N1BEG[3] ,
    \Tile_X1Y3_N1BEG[2] ,
    \Tile_X1Y3_N1BEG[1] ,
    \Tile_X1Y3_N1BEG[0] }),
    .N1END({\Tile_X1Y4_N1BEG[3] ,
    \Tile_X1Y4_N1BEG[2] ,
    \Tile_X1Y4_N1BEG[1] ,
    \Tile_X1Y4_N1BEG[0] }),
    .N2BEG({\Tile_X1Y3_N2BEG[7] ,
    \Tile_X1Y3_N2BEG[6] ,
    \Tile_X1Y3_N2BEG[5] ,
    \Tile_X1Y3_N2BEG[4] ,
    \Tile_X1Y3_N2BEG[3] ,
    \Tile_X1Y3_N2BEG[2] ,
    \Tile_X1Y3_N2BEG[1] ,
    \Tile_X1Y3_N2BEG[0] }),
    .N2BEGb({\Tile_X1Y3_N2BEGb[7] ,
    \Tile_X1Y3_N2BEGb[6] ,
    \Tile_X1Y3_N2BEGb[5] ,
    \Tile_X1Y3_N2BEGb[4] ,
    \Tile_X1Y3_N2BEGb[3] ,
    \Tile_X1Y3_N2BEGb[2] ,
    \Tile_X1Y3_N2BEGb[1] ,
    \Tile_X1Y3_N2BEGb[0] }),
    .N2END({\Tile_X1Y4_N2BEGb[7] ,
    \Tile_X1Y4_N2BEGb[6] ,
    \Tile_X1Y4_N2BEGb[5] ,
    \Tile_X1Y4_N2BEGb[4] ,
    \Tile_X1Y4_N2BEGb[3] ,
    \Tile_X1Y4_N2BEGb[2] ,
    \Tile_X1Y4_N2BEGb[1] ,
    \Tile_X1Y4_N2BEGb[0] }),
    .N2MID({\Tile_X1Y4_N2BEG[7] ,
    \Tile_X1Y4_N2BEG[6] ,
    \Tile_X1Y4_N2BEG[5] ,
    \Tile_X1Y4_N2BEG[4] ,
    \Tile_X1Y4_N2BEG[3] ,
    \Tile_X1Y4_N2BEG[2] ,
    \Tile_X1Y4_N2BEG[1] ,
    \Tile_X1Y4_N2BEG[0] }),
    .N4BEG({\Tile_X1Y3_N4BEG[15] ,
    \Tile_X1Y3_N4BEG[14] ,
    \Tile_X1Y3_N4BEG[13] ,
    \Tile_X1Y3_N4BEG[12] ,
    \Tile_X1Y3_N4BEG[11] ,
    \Tile_X1Y3_N4BEG[10] ,
    \Tile_X1Y3_N4BEG[9] ,
    \Tile_X1Y3_N4BEG[8] ,
    \Tile_X1Y3_N4BEG[7] ,
    \Tile_X1Y3_N4BEG[6] ,
    \Tile_X1Y3_N4BEG[5] ,
    \Tile_X1Y3_N4BEG[4] ,
    \Tile_X1Y3_N4BEG[3] ,
    \Tile_X1Y3_N4BEG[2] ,
    \Tile_X1Y3_N4BEG[1] ,
    \Tile_X1Y3_N4BEG[0] }),
    .N4END({\Tile_X1Y4_N4BEG[15] ,
    \Tile_X1Y4_N4BEG[14] ,
    \Tile_X1Y4_N4BEG[13] ,
    \Tile_X1Y4_N4BEG[12] ,
    \Tile_X1Y4_N4BEG[11] ,
    \Tile_X1Y4_N4BEG[10] ,
    \Tile_X1Y4_N4BEG[9] ,
    \Tile_X1Y4_N4BEG[8] ,
    \Tile_X1Y4_N4BEG[7] ,
    \Tile_X1Y4_N4BEG[6] ,
    \Tile_X1Y4_N4BEG[5] ,
    \Tile_X1Y4_N4BEG[4] ,
    \Tile_X1Y4_N4BEG[3] ,
    \Tile_X1Y4_N4BEG[2] ,
    \Tile_X1Y4_N4BEG[1] ,
    \Tile_X1Y4_N4BEG[0] }),
    .NN4BEG({\Tile_X1Y3_NN4BEG[15] ,
    \Tile_X1Y3_NN4BEG[14] ,
    \Tile_X1Y3_NN4BEG[13] ,
    \Tile_X1Y3_NN4BEG[12] ,
    \Tile_X1Y3_NN4BEG[11] ,
    \Tile_X1Y3_NN4BEG[10] ,
    \Tile_X1Y3_NN4BEG[9] ,
    \Tile_X1Y3_NN4BEG[8] ,
    \Tile_X1Y3_NN4BEG[7] ,
    \Tile_X1Y3_NN4BEG[6] ,
    \Tile_X1Y3_NN4BEG[5] ,
    \Tile_X1Y3_NN4BEG[4] ,
    \Tile_X1Y3_NN4BEG[3] ,
    \Tile_X1Y3_NN4BEG[2] ,
    \Tile_X1Y3_NN4BEG[1] ,
    \Tile_X1Y3_NN4BEG[0] }),
    .NN4END({\Tile_X1Y4_NN4BEG[15] ,
    \Tile_X1Y4_NN4BEG[14] ,
    \Tile_X1Y4_NN4BEG[13] ,
    \Tile_X1Y4_NN4BEG[12] ,
    \Tile_X1Y4_NN4BEG[11] ,
    \Tile_X1Y4_NN4BEG[10] ,
    \Tile_X1Y4_NN4BEG[9] ,
    \Tile_X1Y4_NN4BEG[8] ,
    \Tile_X1Y4_NN4BEG[7] ,
    \Tile_X1Y4_NN4BEG[6] ,
    \Tile_X1Y4_NN4BEG[5] ,
    \Tile_X1Y4_NN4BEG[4] ,
    \Tile_X1Y4_NN4BEG[3] ,
    \Tile_X1Y4_NN4BEG[2] ,
    \Tile_X1Y4_NN4BEG[1] ,
    \Tile_X1Y4_NN4BEG[0] }),
    .S1BEG({\Tile_X1Y3_S1BEG[3] ,
    \Tile_X1Y3_S1BEG[2] ,
    \Tile_X1Y3_S1BEG[1] ,
    \Tile_X1Y3_S1BEG[0] }),
    .S1END({\Tile_X1Y2_S1BEG[3] ,
    \Tile_X1Y2_S1BEG[2] ,
    \Tile_X1Y2_S1BEG[1] ,
    \Tile_X1Y2_S1BEG[0] }),
    .S2BEG({\Tile_X1Y3_S2BEG[7] ,
    \Tile_X1Y3_S2BEG[6] ,
    \Tile_X1Y3_S2BEG[5] ,
    \Tile_X1Y3_S2BEG[4] ,
    \Tile_X1Y3_S2BEG[3] ,
    \Tile_X1Y3_S2BEG[2] ,
    \Tile_X1Y3_S2BEG[1] ,
    \Tile_X1Y3_S2BEG[0] }),
    .S2BEGb({\Tile_X1Y3_S2BEGb[7] ,
    \Tile_X1Y3_S2BEGb[6] ,
    \Tile_X1Y3_S2BEGb[5] ,
    \Tile_X1Y3_S2BEGb[4] ,
    \Tile_X1Y3_S2BEGb[3] ,
    \Tile_X1Y3_S2BEGb[2] ,
    \Tile_X1Y3_S2BEGb[1] ,
    \Tile_X1Y3_S2BEGb[0] }),
    .S2END({\Tile_X1Y2_S2BEGb[7] ,
    \Tile_X1Y2_S2BEGb[6] ,
    \Tile_X1Y2_S2BEGb[5] ,
    \Tile_X1Y2_S2BEGb[4] ,
    \Tile_X1Y2_S2BEGb[3] ,
    \Tile_X1Y2_S2BEGb[2] ,
    \Tile_X1Y2_S2BEGb[1] ,
    \Tile_X1Y2_S2BEGb[0] }),
    .S2MID({\Tile_X1Y2_S2BEG[7] ,
    \Tile_X1Y2_S2BEG[6] ,
    \Tile_X1Y2_S2BEG[5] ,
    \Tile_X1Y2_S2BEG[4] ,
    \Tile_X1Y2_S2BEG[3] ,
    \Tile_X1Y2_S2BEG[2] ,
    \Tile_X1Y2_S2BEG[1] ,
    \Tile_X1Y2_S2BEG[0] }),
    .S4BEG({\Tile_X1Y3_S4BEG[15] ,
    \Tile_X1Y3_S4BEG[14] ,
    \Tile_X1Y3_S4BEG[13] ,
    \Tile_X1Y3_S4BEG[12] ,
    \Tile_X1Y3_S4BEG[11] ,
    \Tile_X1Y3_S4BEG[10] ,
    \Tile_X1Y3_S4BEG[9] ,
    \Tile_X1Y3_S4BEG[8] ,
    \Tile_X1Y3_S4BEG[7] ,
    \Tile_X1Y3_S4BEG[6] ,
    \Tile_X1Y3_S4BEG[5] ,
    \Tile_X1Y3_S4BEG[4] ,
    \Tile_X1Y3_S4BEG[3] ,
    \Tile_X1Y3_S4BEG[2] ,
    \Tile_X1Y3_S4BEG[1] ,
    \Tile_X1Y3_S4BEG[0] }),
    .S4END({\Tile_X1Y2_S4BEG[15] ,
    \Tile_X1Y2_S4BEG[14] ,
    \Tile_X1Y2_S4BEG[13] ,
    \Tile_X1Y2_S4BEG[12] ,
    \Tile_X1Y2_S4BEG[11] ,
    \Tile_X1Y2_S4BEG[10] ,
    \Tile_X1Y2_S4BEG[9] ,
    \Tile_X1Y2_S4BEG[8] ,
    \Tile_X1Y2_S4BEG[7] ,
    \Tile_X1Y2_S4BEG[6] ,
    \Tile_X1Y2_S4BEG[5] ,
    \Tile_X1Y2_S4BEG[4] ,
    \Tile_X1Y2_S4BEG[3] ,
    \Tile_X1Y2_S4BEG[2] ,
    \Tile_X1Y2_S4BEG[1] ,
    \Tile_X1Y2_S4BEG[0] }),
    .SS4BEG({\Tile_X1Y3_SS4BEG[15] ,
    \Tile_X1Y3_SS4BEG[14] ,
    \Tile_X1Y3_SS4BEG[13] ,
    \Tile_X1Y3_SS4BEG[12] ,
    \Tile_X1Y3_SS4BEG[11] ,
    \Tile_X1Y3_SS4BEG[10] ,
    \Tile_X1Y3_SS4BEG[9] ,
    \Tile_X1Y3_SS4BEG[8] ,
    \Tile_X1Y3_SS4BEG[7] ,
    \Tile_X1Y3_SS4BEG[6] ,
    \Tile_X1Y3_SS4BEG[5] ,
    \Tile_X1Y3_SS4BEG[4] ,
    \Tile_X1Y3_SS4BEG[3] ,
    \Tile_X1Y3_SS4BEG[2] ,
    \Tile_X1Y3_SS4BEG[1] ,
    \Tile_X1Y3_SS4BEG[0] }),
    .SS4END({\Tile_X1Y2_SS4BEG[15] ,
    \Tile_X1Y2_SS4BEG[14] ,
    \Tile_X1Y2_SS4BEG[13] ,
    \Tile_X1Y2_SS4BEG[12] ,
    \Tile_X1Y2_SS4BEG[11] ,
    \Tile_X1Y2_SS4BEG[10] ,
    \Tile_X1Y2_SS4BEG[9] ,
    \Tile_X1Y2_SS4BEG[8] ,
    \Tile_X1Y2_SS4BEG[7] ,
    \Tile_X1Y2_SS4BEG[6] ,
    \Tile_X1Y2_SS4BEG[5] ,
    \Tile_X1Y2_SS4BEG[4] ,
    \Tile_X1Y2_SS4BEG[3] ,
    \Tile_X1Y2_SS4BEG[2] ,
    \Tile_X1Y2_SS4BEG[1] ,
    \Tile_X1Y2_SS4BEG[0] }),
    .W1BEG({\Tile_X1Y3_W1BEG[3] ,
    \Tile_X1Y3_W1BEG[2] ,
    \Tile_X1Y3_W1BEG[1] ,
    \Tile_X1Y3_W1BEG[0] }),
    .W1END({\Tile_X2Y3_W1BEG[3] ,
    \Tile_X2Y3_W1BEG[2] ,
    \Tile_X2Y3_W1BEG[1] ,
    \Tile_X2Y3_W1BEG[0] }),
    .W2BEG({\Tile_X1Y3_W2BEG[7] ,
    \Tile_X1Y3_W2BEG[6] ,
    \Tile_X1Y3_W2BEG[5] ,
    \Tile_X1Y3_W2BEG[4] ,
    \Tile_X1Y3_W2BEG[3] ,
    \Tile_X1Y3_W2BEG[2] ,
    \Tile_X1Y3_W2BEG[1] ,
    \Tile_X1Y3_W2BEG[0] }),
    .W2BEGb({\Tile_X1Y3_W2BEGb[7] ,
    \Tile_X1Y3_W2BEGb[6] ,
    \Tile_X1Y3_W2BEGb[5] ,
    \Tile_X1Y3_W2BEGb[4] ,
    \Tile_X1Y3_W2BEGb[3] ,
    \Tile_X1Y3_W2BEGb[2] ,
    \Tile_X1Y3_W2BEGb[1] ,
    \Tile_X1Y3_W2BEGb[0] }),
    .W2END({\Tile_X2Y3_W2BEGb[7] ,
    \Tile_X2Y3_W2BEGb[6] ,
    \Tile_X2Y3_W2BEGb[5] ,
    \Tile_X2Y3_W2BEGb[4] ,
    \Tile_X2Y3_W2BEGb[3] ,
    \Tile_X2Y3_W2BEGb[2] ,
    \Tile_X2Y3_W2BEGb[1] ,
    \Tile_X2Y3_W2BEGb[0] }),
    .W2MID({\Tile_X2Y3_W2BEG[7] ,
    \Tile_X2Y3_W2BEG[6] ,
    \Tile_X2Y3_W2BEG[5] ,
    \Tile_X2Y3_W2BEG[4] ,
    \Tile_X2Y3_W2BEG[3] ,
    \Tile_X2Y3_W2BEG[2] ,
    \Tile_X2Y3_W2BEG[1] ,
    \Tile_X2Y3_W2BEG[0] }),
    .W6BEG({\Tile_X1Y3_W6BEG[11] ,
    \Tile_X1Y3_W6BEG[10] ,
    \Tile_X1Y3_W6BEG[9] ,
    \Tile_X1Y3_W6BEG[8] ,
    \Tile_X1Y3_W6BEG[7] ,
    \Tile_X1Y3_W6BEG[6] ,
    \Tile_X1Y3_W6BEG[5] ,
    \Tile_X1Y3_W6BEG[4] ,
    \Tile_X1Y3_W6BEG[3] ,
    \Tile_X1Y3_W6BEG[2] ,
    \Tile_X1Y3_W6BEG[1] ,
    \Tile_X1Y3_W6BEG[0] }),
    .W6END({\Tile_X2Y3_W6BEG[11] ,
    \Tile_X2Y3_W6BEG[10] ,
    \Tile_X2Y3_W6BEG[9] ,
    \Tile_X2Y3_W6BEG[8] ,
    \Tile_X2Y3_W6BEG[7] ,
    \Tile_X2Y3_W6BEG[6] ,
    \Tile_X2Y3_W6BEG[5] ,
    \Tile_X2Y3_W6BEG[4] ,
    \Tile_X2Y3_W6BEG[3] ,
    \Tile_X2Y3_W6BEG[2] ,
    \Tile_X2Y3_W6BEG[1] ,
    \Tile_X2Y3_W6BEG[0] }),
    .WW4BEG({\Tile_X1Y3_WW4BEG[15] ,
    \Tile_X1Y3_WW4BEG[14] ,
    \Tile_X1Y3_WW4BEG[13] ,
    \Tile_X1Y3_WW4BEG[12] ,
    \Tile_X1Y3_WW4BEG[11] ,
    \Tile_X1Y3_WW4BEG[10] ,
    \Tile_X1Y3_WW4BEG[9] ,
    \Tile_X1Y3_WW4BEG[8] ,
    \Tile_X1Y3_WW4BEG[7] ,
    \Tile_X1Y3_WW4BEG[6] ,
    \Tile_X1Y3_WW4BEG[5] ,
    \Tile_X1Y3_WW4BEG[4] ,
    \Tile_X1Y3_WW4BEG[3] ,
    \Tile_X1Y3_WW4BEG[2] ,
    \Tile_X1Y3_WW4BEG[1] ,
    \Tile_X1Y3_WW4BEG[0] }),
    .WW4END({\Tile_X2Y3_WW4BEG[15] ,
    \Tile_X2Y3_WW4BEG[14] ,
    \Tile_X2Y3_WW4BEG[13] ,
    \Tile_X2Y3_WW4BEG[12] ,
    \Tile_X2Y3_WW4BEG[11] ,
    \Tile_X2Y3_WW4BEG[10] ,
    \Tile_X2Y3_WW4BEG[9] ,
    \Tile_X2Y3_WW4BEG[8] ,
    \Tile_X2Y3_WW4BEG[7] ,
    \Tile_X2Y3_WW4BEG[6] ,
    \Tile_X2Y3_WW4BEG[5] ,
    \Tile_X2Y3_WW4BEG[4] ,
    \Tile_X2Y3_WW4BEG[3] ,
    \Tile_X2Y3_WW4BEG[2] ,
    \Tile_X2Y3_WW4BEG[1] ,
    \Tile_X2Y3_WW4BEG[0] }));
 LUT4AB Tile_X1Y4_LUT4AB (.Ci(Tile_X1Y5_Co),
    .Co(Tile_X1Y4_Co),
    .UserCLK(Tile_X1Y5_UserCLKo),
    .UserCLKo(Tile_X1Y4_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X1Y4_E1BEG[3] ,
    \Tile_X1Y4_E1BEG[2] ,
    \Tile_X1Y4_E1BEG[1] ,
    \Tile_X1Y4_E1BEG[0] }),
    .E1END({\Tile_X0Y4_E1BEG[3] ,
    \Tile_X0Y4_E1BEG[2] ,
    \Tile_X0Y4_E1BEG[1] ,
    \Tile_X0Y4_E1BEG[0] }),
    .E2BEG({\Tile_X1Y4_E2BEG[7] ,
    \Tile_X1Y4_E2BEG[6] ,
    \Tile_X1Y4_E2BEG[5] ,
    \Tile_X1Y4_E2BEG[4] ,
    \Tile_X1Y4_E2BEG[3] ,
    \Tile_X1Y4_E2BEG[2] ,
    \Tile_X1Y4_E2BEG[1] ,
    \Tile_X1Y4_E2BEG[0] }),
    .E2BEGb({\Tile_X1Y4_E2BEGb[7] ,
    \Tile_X1Y4_E2BEGb[6] ,
    \Tile_X1Y4_E2BEGb[5] ,
    \Tile_X1Y4_E2BEGb[4] ,
    \Tile_X1Y4_E2BEGb[3] ,
    \Tile_X1Y4_E2BEGb[2] ,
    \Tile_X1Y4_E2BEGb[1] ,
    \Tile_X1Y4_E2BEGb[0] }),
    .E2END({\Tile_X0Y4_E2BEGb[7] ,
    \Tile_X0Y4_E2BEGb[6] ,
    \Tile_X0Y4_E2BEGb[5] ,
    \Tile_X0Y4_E2BEGb[4] ,
    \Tile_X0Y4_E2BEGb[3] ,
    \Tile_X0Y4_E2BEGb[2] ,
    \Tile_X0Y4_E2BEGb[1] ,
    \Tile_X0Y4_E2BEGb[0] }),
    .E2MID({\Tile_X0Y4_E2BEG[7] ,
    \Tile_X0Y4_E2BEG[6] ,
    \Tile_X0Y4_E2BEG[5] ,
    \Tile_X0Y4_E2BEG[4] ,
    \Tile_X0Y4_E2BEG[3] ,
    \Tile_X0Y4_E2BEG[2] ,
    \Tile_X0Y4_E2BEG[1] ,
    \Tile_X0Y4_E2BEG[0] }),
    .E6BEG({\Tile_X1Y4_E6BEG[11] ,
    \Tile_X1Y4_E6BEG[10] ,
    \Tile_X1Y4_E6BEG[9] ,
    \Tile_X1Y4_E6BEG[8] ,
    \Tile_X1Y4_E6BEG[7] ,
    \Tile_X1Y4_E6BEG[6] ,
    \Tile_X1Y4_E6BEG[5] ,
    \Tile_X1Y4_E6BEG[4] ,
    \Tile_X1Y4_E6BEG[3] ,
    \Tile_X1Y4_E6BEG[2] ,
    \Tile_X1Y4_E6BEG[1] ,
    \Tile_X1Y4_E6BEG[0] }),
    .E6END({\Tile_X0Y4_E6BEG[11] ,
    \Tile_X0Y4_E6BEG[10] ,
    \Tile_X0Y4_E6BEG[9] ,
    \Tile_X0Y4_E6BEG[8] ,
    \Tile_X0Y4_E6BEG[7] ,
    \Tile_X0Y4_E6BEG[6] ,
    \Tile_X0Y4_E6BEG[5] ,
    \Tile_X0Y4_E6BEG[4] ,
    \Tile_X0Y4_E6BEG[3] ,
    \Tile_X0Y4_E6BEG[2] ,
    \Tile_X0Y4_E6BEG[1] ,
    \Tile_X0Y4_E6BEG[0] }),
    .EE4BEG({\Tile_X1Y4_EE4BEG[15] ,
    \Tile_X1Y4_EE4BEG[14] ,
    \Tile_X1Y4_EE4BEG[13] ,
    \Tile_X1Y4_EE4BEG[12] ,
    \Tile_X1Y4_EE4BEG[11] ,
    \Tile_X1Y4_EE4BEG[10] ,
    \Tile_X1Y4_EE4BEG[9] ,
    \Tile_X1Y4_EE4BEG[8] ,
    \Tile_X1Y4_EE4BEG[7] ,
    \Tile_X1Y4_EE4BEG[6] ,
    \Tile_X1Y4_EE4BEG[5] ,
    \Tile_X1Y4_EE4BEG[4] ,
    \Tile_X1Y4_EE4BEG[3] ,
    \Tile_X1Y4_EE4BEG[2] ,
    \Tile_X1Y4_EE4BEG[1] ,
    \Tile_X1Y4_EE4BEG[0] }),
    .EE4END({\Tile_X0Y4_EE4BEG[15] ,
    \Tile_X0Y4_EE4BEG[14] ,
    \Tile_X0Y4_EE4BEG[13] ,
    \Tile_X0Y4_EE4BEG[12] ,
    \Tile_X0Y4_EE4BEG[11] ,
    \Tile_X0Y4_EE4BEG[10] ,
    \Tile_X0Y4_EE4BEG[9] ,
    \Tile_X0Y4_EE4BEG[8] ,
    \Tile_X0Y4_EE4BEG[7] ,
    \Tile_X0Y4_EE4BEG[6] ,
    \Tile_X0Y4_EE4BEG[5] ,
    \Tile_X0Y4_EE4BEG[4] ,
    \Tile_X0Y4_EE4BEG[3] ,
    \Tile_X0Y4_EE4BEG[2] ,
    \Tile_X0Y4_EE4BEG[1] ,
    \Tile_X0Y4_EE4BEG[0] }),
    .FrameData({\Tile_X0Y4_FrameData_O[31] ,
    \Tile_X0Y4_FrameData_O[30] ,
    \Tile_X0Y4_FrameData_O[29] ,
    \Tile_X0Y4_FrameData_O[28] ,
    \Tile_X0Y4_FrameData_O[27] ,
    \Tile_X0Y4_FrameData_O[26] ,
    \Tile_X0Y4_FrameData_O[25] ,
    \Tile_X0Y4_FrameData_O[24] ,
    \Tile_X0Y4_FrameData_O[23] ,
    \Tile_X0Y4_FrameData_O[22] ,
    \Tile_X0Y4_FrameData_O[21] ,
    \Tile_X0Y4_FrameData_O[20] ,
    \Tile_X0Y4_FrameData_O[19] ,
    \Tile_X0Y4_FrameData_O[18] ,
    \Tile_X0Y4_FrameData_O[17] ,
    \Tile_X0Y4_FrameData_O[16] ,
    \Tile_X0Y4_FrameData_O[15] ,
    \Tile_X0Y4_FrameData_O[14] ,
    \Tile_X0Y4_FrameData_O[13] ,
    \Tile_X0Y4_FrameData_O[12] ,
    \Tile_X0Y4_FrameData_O[11] ,
    \Tile_X0Y4_FrameData_O[10] ,
    \Tile_X0Y4_FrameData_O[9] ,
    \Tile_X0Y4_FrameData_O[8] ,
    \Tile_X0Y4_FrameData_O[7] ,
    \Tile_X0Y4_FrameData_O[6] ,
    \Tile_X0Y4_FrameData_O[5] ,
    \Tile_X0Y4_FrameData_O[4] ,
    \Tile_X0Y4_FrameData_O[3] ,
    \Tile_X0Y4_FrameData_O[2] ,
    \Tile_X0Y4_FrameData_O[1] ,
    \Tile_X0Y4_FrameData_O[0] }),
    .FrameData_O({\Tile_X1Y4_FrameData_O[31] ,
    \Tile_X1Y4_FrameData_O[30] ,
    \Tile_X1Y4_FrameData_O[29] ,
    \Tile_X1Y4_FrameData_O[28] ,
    \Tile_X1Y4_FrameData_O[27] ,
    \Tile_X1Y4_FrameData_O[26] ,
    \Tile_X1Y4_FrameData_O[25] ,
    \Tile_X1Y4_FrameData_O[24] ,
    \Tile_X1Y4_FrameData_O[23] ,
    \Tile_X1Y4_FrameData_O[22] ,
    \Tile_X1Y4_FrameData_O[21] ,
    \Tile_X1Y4_FrameData_O[20] ,
    \Tile_X1Y4_FrameData_O[19] ,
    \Tile_X1Y4_FrameData_O[18] ,
    \Tile_X1Y4_FrameData_O[17] ,
    \Tile_X1Y4_FrameData_O[16] ,
    \Tile_X1Y4_FrameData_O[15] ,
    \Tile_X1Y4_FrameData_O[14] ,
    \Tile_X1Y4_FrameData_O[13] ,
    \Tile_X1Y4_FrameData_O[12] ,
    \Tile_X1Y4_FrameData_O[11] ,
    \Tile_X1Y4_FrameData_O[10] ,
    \Tile_X1Y4_FrameData_O[9] ,
    \Tile_X1Y4_FrameData_O[8] ,
    \Tile_X1Y4_FrameData_O[7] ,
    \Tile_X1Y4_FrameData_O[6] ,
    \Tile_X1Y4_FrameData_O[5] ,
    \Tile_X1Y4_FrameData_O[4] ,
    \Tile_X1Y4_FrameData_O[3] ,
    \Tile_X1Y4_FrameData_O[2] ,
    \Tile_X1Y4_FrameData_O[1] ,
    \Tile_X1Y4_FrameData_O[0] }),
    .FrameStrobe({\Tile_X1Y5_FrameStrobe_O[19] ,
    \Tile_X1Y5_FrameStrobe_O[18] ,
    \Tile_X1Y5_FrameStrobe_O[17] ,
    \Tile_X1Y5_FrameStrobe_O[16] ,
    \Tile_X1Y5_FrameStrobe_O[15] ,
    \Tile_X1Y5_FrameStrobe_O[14] ,
    \Tile_X1Y5_FrameStrobe_O[13] ,
    \Tile_X1Y5_FrameStrobe_O[12] ,
    \Tile_X1Y5_FrameStrobe_O[11] ,
    \Tile_X1Y5_FrameStrobe_O[10] ,
    \Tile_X1Y5_FrameStrobe_O[9] ,
    \Tile_X1Y5_FrameStrobe_O[8] ,
    \Tile_X1Y5_FrameStrobe_O[7] ,
    \Tile_X1Y5_FrameStrobe_O[6] ,
    \Tile_X1Y5_FrameStrobe_O[5] ,
    \Tile_X1Y5_FrameStrobe_O[4] ,
    \Tile_X1Y5_FrameStrobe_O[3] ,
    \Tile_X1Y5_FrameStrobe_O[2] ,
    \Tile_X1Y5_FrameStrobe_O[1] ,
    \Tile_X1Y5_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X1Y4_FrameStrobe_O[19] ,
    \Tile_X1Y4_FrameStrobe_O[18] ,
    \Tile_X1Y4_FrameStrobe_O[17] ,
    \Tile_X1Y4_FrameStrobe_O[16] ,
    \Tile_X1Y4_FrameStrobe_O[15] ,
    \Tile_X1Y4_FrameStrobe_O[14] ,
    \Tile_X1Y4_FrameStrobe_O[13] ,
    \Tile_X1Y4_FrameStrobe_O[12] ,
    \Tile_X1Y4_FrameStrobe_O[11] ,
    \Tile_X1Y4_FrameStrobe_O[10] ,
    \Tile_X1Y4_FrameStrobe_O[9] ,
    \Tile_X1Y4_FrameStrobe_O[8] ,
    \Tile_X1Y4_FrameStrobe_O[7] ,
    \Tile_X1Y4_FrameStrobe_O[6] ,
    \Tile_X1Y4_FrameStrobe_O[5] ,
    \Tile_X1Y4_FrameStrobe_O[4] ,
    \Tile_X1Y4_FrameStrobe_O[3] ,
    \Tile_X1Y4_FrameStrobe_O[2] ,
    \Tile_X1Y4_FrameStrobe_O[1] ,
    \Tile_X1Y4_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X1Y4_N1BEG[3] ,
    \Tile_X1Y4_N1BEG[2] ,
    \Tile_X1Y4_N1BEG[1] ,
    \Tile_X1Y4_N1BEG[0] }),
    .N1END({\Tile_X1Y5_N1BEG[3] ,
    \Tile_X1Y5_N1BEG[2] ,
    \Tile_X1Y5_N1BEG[1] ,
    \Tile_X1Y5_N1BEG[0] }),
    .N2BEG({\Tile_X1Y4_N2BEG[7] ,
    \Tile_X1Y4_N2BEG[6] ,
    \Tile_X1Y4_N2BEG[5] ,
    \Tile_X1Y4_N2BEG[4] ,
    \Tile_X1Y4_N2BEG[3] ,
    \Tile_X1Y4_N2BEG[2] ,
    \Tile_X1Y4_N2BEG[1] ,
    \Tile_X1Y4_N2BEG[0] }),
    .N2BEGb({\Tile_X1Y4_N2BEGb[7] ,
    \Tile_X1Y4_N2BEGb[6] ,
    \Tile_X1Y4_N2BEGb[5] ,
    \Tile_X1Y4_N2BEGb[4] ,
    \Tile_X1Y4_N2BEGb[3] ,
    \Tile_X1Y4_N2BEGb[2] ,
    \Tile_X1Y4_N2BEGb[1] ,
    \Tile_X1Y4_N2BEGb[0] }),
    .N2END({\Tile_X1Y5_N2BEGb[7] ,
    \Tile_X1Y5_N2BEGb[6] ,
    \Tile_X1Y5_N2BEGb[5] ,
    \Tile_X1Y5_N2BEGb[4] ,
    \Tile_X1Y5_N2BEGb[3] ,
    \Tile_X1Y5_N2BEGb[2] ,
    \Tile_X1Y5_N2BEGb[1] ,
    \Tile_X1Y5_N2BEGb[0] }),
    .N2MID({\Tile_X1Y5_N2BEG[7] ,
    \Tile_X1Y5_N2BEG[6] ,
    \Tile_X1Y5_N2BEG[5] ,
    \Tile_X1Y5_N2BEG[4] ,
    \Tile_X1Y5_N2BEG[3] ,
    \Tile_X1Y5_N2BEG[2] ,
    \Tile_X1Y5_N2BEG[1] ,
    \Tile_X1Y5_N2BEG[0] }),
    .N4BEG({\Tile_X1Y4_N4BEG[15] ,
    \Tile_X1Y4_N4BEG[14] ,
    \Tile_X1Y4_N4BEG[13] ,
    \Tile_X1Y4_N4BEG[12] ,
    \Tile_X1Y4_N4BEG[11] ,
    \Tile_X1Y4_N4BEG[10] ,
    \Tile_X1Y4_N4BEG[9] ,
    \Tile_X1Y4_N4BEG[8] ,
    \Tile_X1Y4_N4BEG[7] ,
    \Tile_X1Y4_N4BEG[6] ,
    \Tile_X1Y4_N4BEG[5] ,
    \Tile_X1Y4_N4BEG[4] ,
    \Tile_X1Y4_N4BEG[3] ,
    \Tile_X1Y4_N4BEG[2] ,
    \Tile_X1Y4_N4BEG[1] ,
    \Tile_X1Y4_N4BEG[0] }),
    .N4END({\Tile_X1Y5_N4BEG[15] ,
    \Tile_X1Y5_N4BEG[14] ,
    \Tile_X1Y5_N4BEG[13] ,
    \Tile_X1Y5_N4BEG[12] ,
    \Tile_X1Y5_N4BEG[11] ,
    \Tile_X1Y5_N4BEG[10] ,
    \Tile_X1Y5_N4BEG[9] ,
    \Tile_X1Y5_N4BEG[8] ,
    \Tile_X1Y5_N4BEG[7] ,
    \Tile_X1Y5_N4BEG[6] ,
    \Tile_X1Y5_N4BEG[5] ,
    \Tile_X1Y5_N4BEG[4] ,
    \Tile_X1Y5_N4BEG[3] ,
    \Tile_X1Y5_N4BEG[2] ,
    \Tile_X1Y5_N4BEG[1] ,
    \Tile_X1Y5_N4BEG[0] }),
    .NN4BEG({\Tile_X1Y4_NN4BEG[15] ,
    \Tile_X1Y4_NN4BEG[14] ,
    \Tile_X1Y4_NN4BEG[13] ,
    \Tile_X1Y4_NN4BEG[12] ,
    \Tile_X1Y4_NN4BEG[11] ,
    \Tile_X1Y4_NN4BEG[10] ,
    \Tile_X1Y4_NN4BEG[9] ,
    \Tile_X1Y4_NN4BEG[8] ,
    \Tile_X1Y4_NN4BEG[7] ,
    \Tile_X1Y4_NN4BEG[6] ,
    \Tile_X1Y4_NN4BEG[5] ,
    \Tile_X1Y4_NN4BEG[4] ,
    \Tile_X1Y4_NN4BEG[3] ,
    \Tile_X1Y4_NN4BEG[2] ,
    \Tile_X1Y4_NN4BEG[1] ,
    \Tile_X1Y4_NN4BEG[0] }),
    .NN4END({\Tile_X1Y5_NN4BEG[15] ,
    \Tile_X1Y5_NN4BEG[14] ,
    \Tile_X1Y5_NN4BEG[13] ,
    \Tile_X1Y5_NN4BEG[12] ,
    \Tile_X1Y5_NN4BEG[11] ,
    \Tile_X1Y5_NN4BEG[10] ,
    \Tile_X1Y5_NN4BEG[9] ,
    \Tile_X1Y5_NN4BEG[8] ,
    \Tile_X1Y5_NN4BEG[7] ,
    \Tile_X1Y5_NN4BEG[6] ,
    \Tile_X1Y5_NN4BEG[5] ,
    \Tile_X1Y5_NN4BEG[4] ,
    \Tile_X1Y5_NN4BEG[3] ,
    \Tile_X1Y5_NN4BEG[2] ,
    \Tile_X1Y5_NN4BEG[1] ,
    \Tile_X1Y5_NN4BEG[0] }),
    .S1BEG({\Tile_X1Y4_S1BEG[3] ,
    \Tile_X1Y4_S1BEG[2] ,
    \Tile_X1Y4_S1BEG[1] ,
    \Tile_X1Y4_S1BEG[0] }),
    .S1END({\Tile_X1Y3_S1BEG[3] ,
    \Tile_X1Y3_S1BEG[2] ,
    \Tile_X1Y3_S1BEG[1] ,
    \Tile_X1Y3_S1BEG[0] }),
    .S2BEG({\Tile_X1Y4_S2BEG[7] ,
    \Tile_X1Y4_S2BEG[6] ,
    \Tile_X1Y4_S2BEG[5] ,
    \Tile_X1Y4_S2BEG[4] ,
    \Tile_X1Y4_S2BEG[3] ,
    \Tile_X1Y4_S2BEG[2] ,
    \Tile_X1Y4_S2BEG[1] ,
    \Tile_X1Y4_S2BEG[0] }),
    .S2BEGb({\Tile_X1Y4_S2BEGb[7] ,
    \Tile_X1Y4_S2BEGb[6] ,
    \Tile_X1Y4_S2BEGb[5] ,
    \Tile_X1Y4_S2BEGb[4] ,
    \Tile_X1Y4_S2BEGb[3] ,
    \Tile_X1Y4_S2BEGb[2] ,
    \Tile_X1Y4_S2BEGb[1] ,
    \Tile_X1Y4_S2BEGb[0] }),
    .S2END({\Tile_X1Y3_S2BEGb[7] ,
    \Tile_X1Y3_S2BEGb[6] ,
    \Tile_X1Y3_S2BEGb[5] ,
    \Tile_X1Y3_S2BEGb[4] ,
    \Tile_X1Y3_S2BEGb[3] ,
    \Tile_X1Y3_S2BEGb[2] ,
    \Tile_X1Y3_S2BEGb[1] ,
    \Tile_X1Y3_S2BEGb[0] }),
    .S2MID({\Tile_X1Y3_S2BEG[7] ,
    \Tile_X1Y3_S2BEG[6] ,
    \Tile_X1Y3_S2BEG[5] ,
    \Tile_X1Y3_S2BEG[4] ,
    \Tile_X1Y3_S2BEG[3] ,
    \Tile_X1Y3_S2BEG[2] ,
    \Tile_X1Y3_S2BEG[1] ,
    \Tile_X1Y3_S2BEG[0] }),
    .S4BEG({\Tile_X1Y4_S4BEG[15] ,
    \Tile_X1Y4_S4BEG[14] ,
    \Tile_X1Y4_S4BEG[13] ,
    \Tile_X1Y4_S4BEG[12] ,
    \Tile_X1Y4_S4BEG[11] ,
    \Tile_X1Y4_S4BEG[10] ,
    \Tile_X1Y4_S4BEG[9] ,
    \Tile_X1Y4_S4BEG[8] ,
    \Tile_X1Y4_S4BEG[7] ,
    \Tile_X1Y4_S4BEG[6] ,
    \Tile_X1Y4_S4BEG[5] ,
    \Tile_X1Y4_S4BEG[4] ,
    \Tile_X1Y4_S4BEG[3] ,
    \Tile_X1Y4_S4BEG[2] ,
    \Tile_X1Y4_S4BEG[1] ,
    \Tile_X1Y4_S4BEG[0] }),
    .S4END({\Tile_X1Y3_S4BEG[15] ,
    \Tile_X1Y3_S4BEG[14] ,
    \Tile_X1Y3_S4BEG[13] ,
    \Tile_X1Y3_S4BEG[12] ,
    \Tile_X1Y3_S4BEG[11] ,
    \Tile_X1Y3_S4BEG[10] ,
    \Tile_X1Y3_S4BEG[9] ,
    \Tile_X1Y3_S4BEG[8] ,
    \Tile_X1Y3_S4BEG[7] ,
    \Tile_X1Y3_S4BEG[6] ,
    \Tile_X1Y3_S4BEG[5] ,
    \Tile_X1Y3_S4BEG[4] ,
    \Tile_X1Y3_S4BEG[3] ,
    \Tile_X1Y3_S4BEG[2] ,
    \Tile_X1Y3_S4BEG[1] ,
    \Tile_X1Y3_S4BEG[0] }),
    .SS4BEG({\Tile_X1Y4_SS4BEG[15] ,
    \Tile_X1Y4_SS4BEG[14] ,
    \Tile_X1Y4_SS4BEG[13] ,
    \Tile_X1Y4_SS4BEG[12] ,
    \Tile_X1Y4_SS4BEG[11] ,
    \Tile_X1Y4_SS4BEG[10] ,
    \Tile_X1Y4_SS4BEG[9] ,
    \Tile_X1Y4_SS4BEG[8] ,
    \Tile_X1Y4_SS4BEG[7] ,
    \Tile_X1Y4_SS4BEG[6] ,
    \Tile_X1Y4_SS4BEG[5] ,
    \Tile_X1Y4_SS4BEG[4] ,
    \Tile_X1Y4_SS4BEG[3] ,
    \Tile_X1Y4_SS4BEG[2] ,
    \Tile_X1Y4_SS4BEG[1] ,
    \Tile_X1Y4_SS4BEG[0] }),
    .SS4END({\Tile_X1Y3_SS4BEG[15] ,
    \Tile_X1Y3_SS4BEG[14] ,
    \Tile_X1Y3_SS4BEG[13] ,
    \Tile_X1Y3_SS4BEG[12] ,
    \Tile_X1Y3_SS4BEG[11] ,
    \Tile_X1Y3_SS4BEG[10] ,
    \Tile_X1Y3_SS4BEG[9] ,
    \Tile_X1Y3_SS4BEG[8] ,
    \Tile_X1Y3_SS4BEG[7] ,
    \Tile_X1Y3_SS4BEG[6] ,
    \Tile_X1Y3_SS4BEG[5] ,
    \Tile_X1Y3_SS4BEG[4] ,
    \Tile_X1Y3_SS4BEG[3] ,
    \Tile_X1Y3_SS4BEG[2] ,
    \Tile_X1Y3_SS4BEG[1] ,
    \Tile_X1Y3_SS4BEG[0] }),
    .W1BEG({\Tile_X1Y4_W1BEG[3] ,
    \Tile_X1Y4_W1BEG[2] ,
    \Tile_X1Y4_W1BEG[1] ,
    \Tile_X1Y4_W1BEG[0] }),
    .W1END({\Tile_X2Y4_W1BEG[3] ,
    \Tile_X2Y4_W1BEG[2] ,
    \Tile_X2Y4_W1BEG[1] ,
    \Tile_X2Y4_W1BEG[0] }),
    .W2BEG({\Tile_X1Y4_W2BEG[7] ,
    \Tile_X1Y4_W2BEG[6] ,
    \Tile_X1Y4_W2BEG[5] ,
    \Tile_X1Y4_W2BEG[4] ,
    \Tile_X1Y4_W2BEG[3] ,
    \Tile_X1Y4_W2BEG[2] ,
    \Tile_X1Y4_W2BEG[1] ,
    \Tile_X1Y4_W2BEG[0] }),
    .W2BEGb({\Tile_X1Y4_W2BEGb[7] ,
    \Tile_X1Y4_W2BEGb[6] ,
    \Tile_X1Y4_W2BEGb[5] ,
    \Tile_X1Y4_W2BEGb[4] ,
    \Tile_X1Y4_W2BEGb[3] ,
    \Tile_X1Y4_W2BEGb[2] ,
    \Tile_X1Y4_W2BEGb[1] ,
    \Tile_X1Y4_W2BEGb[0] }),
    .W2END({\Tile_X2Y4_W2BEGb[7] ,
    \Tile_X2Y4_W2BEGb[6] ,
    \Tile_X2Y4_W2BEGb[5] ,
    \Tile_X2Y4_W2BEGb[4] ,
    \Tile_X2Y4_W2BEGb[3] ,
    \Tile_X2Y4_W2BEGb[2] ,
    \Tile_X2Y4_W2BEGb[1] ,
    \Tile_X2Y4_W2BEGb[0] }),
    .W2MID({\Tile_X2Y4_W2BEG[7] ,
    \Tile_X2Y4_W2BEG[6] ,
    \Tile_X2Y4_W2BEG[5] ,
    \Tile_X2Y4_W2BEG[4] ,
    \Tile_X2Y4_W2BEG[3] ,
    \Tile_X2Y4_W2BEG[2] ,
    \Tile_X2Y4_W2BEG[1] ,
    \Tile_X2Y4_W2BEG[0] }),
    .W6BEG({\Tile_X1Y4_W6BEG[11] ,
    \Tile_X1Y4_W6BEG[10] ,
    \Tile_X1Y4_W6BEG[9] ,
    \Tile_X1Y4_W6BEG[8] ,
    \Tile_X1Y4_W6BEG[7] ,
    \Tile_X1Y4_W6BEG[6] ,
    \Tile_X1Y4_W6BEG[5] ,
    \Tile_X1Y4_W6BEG[4] ,
    \Tile_X1Y4_W6BEG[3] ,
    \Tile_X1Y4_W6BEG[2] ,
    \Tile_X1Y4_W6BEG[1] ,
    \Tile_X1Y4_W6BEG[0] }),
    .W6END({\Tile_X2Y4_W6BEG[11] ,
    \Tile_X2Y4_W6BEG[10] ,
    \Tile_X2Y4_W6BEG[9] ,
    \Tile_X2Y4_W6BEG[8] ,
    \Tile_X2Y4_W6BEG[7] ,
    \Tile_X2Y4_W6BEG[6] ,
    \Tile_X2Y4_W6BEG[5] ,
    \Tile_X2Y4_W6BEG[4] ,
    \Tile_X2Y4_W6BEG[3] ,
    \Tile_X2Y4_W6BEG[2] ,
    \Tile_X2Y4_W6BEG[1] ,
    \Tile_X2Y4_W6BEG[0] }),
    .WW4BEG({\Tile_X1Y4_WW4BEG[15] ,
    \Tile_X1Y4_WW4BEG[14] ,
    \Tile_X1Y4_WW4BEG[13] ,
    \Tile_X1Y4_WW4BEG[12] ,
    \Tile_X1Y4_WW4BEG[11] ,
    \Tile_X1Y4_WW4BEG[10] ,
    \Tile_X1Y4_WW4BEG[9] ,
    \Tile_X1Y4_WW4BEG[8] ,
    \Tile_X1Y4_WW4BEG[7] ,
    \Tile_X1Y4_WW4BEG[6] ,
    \Tile_X1Y4_WW4BEG[5] ,
    \Tile_X1Y4_WW4BEG[4] ,
    \Tile_X1Y4_WW4BEG[3] ,
    \Tile_X1Y4_WW4BEG[2] ,
    \Tile_X1Y4_WW4BEG[1] ,
    \Tile_X1Y4_WW4BEG[0] }),
    .WW4END({\Tile_X2Y4_WW4BEG[15] ,
    \Tile_X2Y4_WW4BEG[14] ,
    \Tile_X2Y4_WW4BEG[13] ,
    \Tile_X2Y4_WW4BEG[12] ,
    \Tile_X2Y4_WW4BEG[11] ,
    \Tile_X2Y4_WW4BEG[10] ,
    \Tile_X2Y4_WW4BEG[9] ,
    \Tile_X2Y4_WW4BEG[8] ,
    \Tile_X2Y4_WW4BEG[7] ,
    \Tile_X2Y4_WW4BEG[6] ,
    \Tile_X2Y4_WW4BEG[5] ,
    \Tile_X2Y4_WW4BEG[4] ,
    \Tile_X2Y4_WW4BEG[3] ,
    \Tile_X2Y4_WW4BEG[2] ,
    \Tile_X2Y4_WW4BEG[1] ,
    \Tile_X2Y4_WW4BEG[0] }));
 LUT4AB Tile_X1Y5_LUT4AB (.Ci(Tile_X1Y6_Co),
    .Co(Tile_X1Y5_Co),
    .UserCLK(Tile_X1Y6_UserCLKo),
    .UserCLKo(Tile_X1Y5_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X1Y5_E1BEG[3] ,
    \Tile_X1Y5_E1BEG[2] ,
    \Tile_X1Y5_E1BEG[1] ,
    \Tile_X1Y5_E1BEG[0] }),
    .E1END({\Tile_X0Y5_E1BEG[3] ,
    \Tile_X0Y5_E1BEG[2] ,
    \Tile_X0Y5_E1BEG[1] ,
    \Tile_X0Y5_E1BEG[0] }),
    .E2BEG({\Tile_X1Y5_E2BEG[7] ,
    \Tile_X1Y5_E2BEG[6] ,
    \Tile_X1Y5_E2BEG[5] ,
    \Tile_X1Y5_E2BEG[4] ,
    \Tile_X1Y5_E2BEG[3] ,
    \Tile_X1Y5_E2BEG[2] ,
    \Tile_X1Y5_E2BEG[1] ,
    \Tile_X1Y5_E2BEG[0] }),
    .E2BEGb({\Tile_X1Y5_E2BEGb[7] ,
    \Tile_X1Y5_E2BEGb[6] ,
    \Tile_X1Y5_E2BEGb[5] ,
    \Tile_X1Y5_E2BEGb[4] ,
    \Tile_X1Y5_E2BEGb[3] ,
    \Tile_X1Y5_E2BEGb[2] ,
    \Tile_X1Y5_E2BEGb[1] ,
    \Tile_X1Y5_E2BEGb[0] }),
    .E2END({\Tile_X0Y5_E2BEGb[7] ,
    \Tile_X0Y5_E2BEGb[6] ,
    \Tile_X0Y5_E2BEGb[5] ,
    \Tile_X0Y5_E2BEGb[4] ,
    \Tile_X0Y5_E2BEGb[3] ,
    \Tile_X0Y5_E2BEGb[2] ,
    \Tile_X0Y5_E2BEGb[1] ,
    \Tile_X0Y5_E2BEGb[0] }),
    .E2MID({\Tile_X0Y5_E2BEG[7] ,
    \Tile_X0Y5_E2BEG[6] ,
    \Tile_X0Y5_E2BEG[5] ,
    \Tile_X0Y5_E2BEG[4] ,
    \Tile_X0Y5_E2BEG[3] ,
    \Tile_X0Y5_E2BEG[2] ,
    \Tile_X0Y5_E2BEG[1] ,
    \Tile_X0Y5_E2BEG[0] }),
    .E6BEG({\Tile_X1Y5_E6BEG[11] ,
    \Tile_X1Y5_E6BEG[10] ,
    \Tile_X1Y5_E6BEG[9] ,
    \Tile_X1Y5_E6BEG[8] ,
    \Tile_X1Y5_E6BEG[7] ,
    \Tile_X1Y5_E6BEG[6] ,
    \Tile_X1Y5_E6BEG[5] ,
    \Tile_X1Y5_E6BEG[4] ,
    \Tile_X1Y5_E6BEG[3] ,
    \Tile_X1Y5_E6BEG[2] ,
    \Tile_X1Y5_E6BEG[1] ,
    \Tile_X1Y5_E6BEG[0] }),
    .E6END({\Tile_X0Y5_E6BEG[11] ,
    \Tile_X0Y5_E6BEG[10] ,
    \Tile_X0Y5_E6BEG[9] ,
    \Tile_X0Y5_E6BEG[8] ,
    \Tile_X0Y5_E6BEG[7] ,
    \Tile_X0Y5_E6BEG[6] ,
    \Tile_X0Y5_E6BEG[5] ,
    \Tile_X0Y5_E6BEG[4] ,
    \Tile_X0Y5_E6BEG[3] ,
    \Tile_X0Y5_E6BEG[2] ,
    \Tile_X0Y5_E6BEG[1] ,
    \Tile_X0Y5_E6BEG[0] }),
    .EE4BEG({\Tile_X1Y5_EE4BEG[15] ,
    \Tile_X1Y5_EE4BEG[14] ,
    \Tile_X1Y5_EE4BEG[13] ,
    \Tile_X1Y5_EE4BEG[12] ,
    \Tile_X1Y5_EE4BEG[11] ,
    \Tile_X1Y5_EE4BEG[10] ,
    \Tile_X1Y5_EE4BEG[9] ,
    \Tile_X1Y5_EE4BEG[8] ,
    \Tile_X1Y5_EE4BEG[7] ,
    \Tile_X1Y5_EE4BEG[6] ,
    \Tile_X1Y5_EE4BEG[5] ,
    \Tile_X1Y5_EE4BEG[4] ,
    \Tile_X1Y5_EE4BEG[3] ,
    \Tile_X1Y5_EE4BEG[2] ,
    \Tile_X1Y5_EE4BEG[1] ,
    \Tile_X1Y5_EE4BEG[0] }),
    .EE4END({\Tile_X0Y5_EE4BEG[15] ,
    \Tile_X0Y5_EE4BEG[14] ,
    \Tile_X0Y5_EE4BEG[13] ,
    \Tile_X0Y5_EE4BEG[12] ,
    \Tile_X0Y5_EE4BEG[11] ,
    \Tile_X0Y5_EE4BEG[10] ,
    \Tile_X0Y5_EE4BEG[9] ,
    \Tile_X0Y5_EE4BEG[8] ,
    \Tile_X0Y5_EE4BEG[7] ,
    \Tile_X0Y5_EE4BEG[6] ,
    \Tile_X0Y5_EE4BEG[5] ,
    \Tile_X0Y5_EE4BEG[4] ,
    \Tile_X0Y5_EE4BEG[3] ,
    \Tile_X0Y5_EE4BEG[2] ,
    \Tile_X0Y5_EE4BEG[1] ,
    \Tile_X0Y5_EE4BEG[0] }),
    .FrameData({\Tile_X0Y5_FrameData_O[31] ,
    \Tile_X0Y5_FrameData_O[30] ,
    \Tile_X0Y5_FrameData_O[29] ,
    \Tile_X0Y5_FrameData_O[28] ,
    \Tile_X0Y5_FrameData_O[27] ,
    \Tile_X0Y5_FrameData_O[26] ,
    \Tile_X0Y5_FrameData_O[25] ,
    \Tile_X0Y5_FrameData_O[24] ,
    \Tile_X0Y5_FrameData_O[23] ,
    \Tile_X0Y5_FrameData_O[22] ,
    \Tile_X0Y5_FrameData_O[21] ,
    \Tile_X0Y5_FrameData_O[20] ,
    \Tile_X0Y5_FrameData_O[19] ,
    \Tile_X0Y5_FrameData_O[18] ,
    \Tile_X0Y5_FrameData_O[17] ,
    \Tile_X0Y5_FrameData_O[16] ,
    \Tile_X0Y5_FrameData_O[15] ,
    \Tile_X0Y5_FrameData_O[14] ,
    \Tile_X0Y5_FrameData_O[13] ,
    \Tile_X0Y5_FrameData_O[12] ,
    \Tile_X0Y5_FrameData_O[11] ,
    \Tile_X0Y5_FrameData_O[10] ,
    \Tile_X0Y5_FrameData_O[9] ,
    \Tile_X0Y5_FrameData_O[8] ,
    \Tile_X0Y5_FrameData_O[7] ,
    \Tile_X0Y5_FrameData_O[6] ,
    \Tile_X0Y5_FrameData_O[5] ,
    \Tile_X0Y5_FrameData_O[4] ,
    \Tile_X0Y5_FrameData_O[3] ,
    \Tile_X0Y5_FrameData_O[2] ,
    \Tile_X0Y5_FrameData_O[1] ,
    \Tile_X0Y5_FrameData_O[0] }),
    .FrameData_O({\Tile_X1Y5_FrameData_O[31] ,
    \Tile_X1Y5_FrameData_O[30] ,
    \Tile_X1Y5_FrameData_O[29] ,
    \Tile_X1Y5_FrameData_O[28] ,
    \Tile_X1Y5_FrameData_O[27] ,
    \Tile_X1Y5_FrameData_O[26] ,
    \Tile_X1Y5_FrameData_O[25] ,
    \Tile_X1Y5_FrameData_O[24] ,
    \Tile_X1Y5_FrameData_O[23] ,
    \Tile_X1Y5_FrameData_O[22] ,
    \Tile_X1Y5_FrameData_O[21] ,
    \Tile_X1Y5_FrameData_O[20] ,
    \Tile_X1Y5_FrameData_O[19] ,
    \Tile_X1Y5_FrameData_O[18] ,
    \Tile_X1Y5_FrameData_O[17] ,
    \Tile_X1Y5_FrameData_O[16] ,
    \Tile_X1Y5_FrameData_O[15] ,
    \Tile_X1Y5_FrameData_O[14] ,
    \Tile_X1Y5_FrameData_O[13] ,
    \Tile_X1Y5_FrameData_O[12] ,
    \Tile_X1Y5_FrameData_O[11] ,
    \Tile_X1Y5_FrameData_O[10] ,
    \Tile_X1Y5_FrameData_O[9] ,
    \Tile_X1Y5_FrameData_O[8] ,
    \Tile_X1Y5_FrameData_O[7] ,
    \Tile_X1Y5_FrameData_O[6] ,
    \Tile_X1Y5_FrameData_O[5] ,
    \Tile_X1Y5_FrameData_O[4] ,
    \Tile_X1Y5_FrameData_O[3] ,
    \Tile_X1Y5_FrameData_O[2] ,
    \Tile_X1Y5_FrameData_O[1] ,
    \Tile_X1Y5_FrameData_O[0] }),
    .FrameStrobe({\Tile_X1Y6_FrameStrobe_O[19] ,
    \Tile_X1Y6_FrameStrobe_O[18] ,
    \Tile_X1Y6_FrameStrobe_O[17] ,
    \Tile_X1Y6_FrameStrobe_O[16] ,
    \Tile_X1Y6_FrameStrobe_O[15] ,
    \Tile_X1Y6_FrameStrobe_O[14] ,
    \Tile_X1Y6_FrameStrobe_O[13] ,
    \Tile_X1Y6_FrameStrobe_O[12] ,
    \Tile_X1Y6_FrameStrobe_O[11] ,
    \Tile_X1Y6_FrameStrobe_O[10] ,
    \Tile_X1Y6_FrameStrobe_O[9] ,
    \Tile_X1Y6_FrameStrobe_O[8] ,
    \Tile_X1Y6_FrameStrobe_O[7] ,
    \Tile_X1Y6_FrameStrobe_O[6] ,
    \Tile_X1Y6_FrameStrobe_O[5] ,
    \Tile_X1Y6_FrameStrobe_O[4] ,
    \Tile_X1Y6_FrameStrobe_O[3] ,
    \Tile_X1Y6_FrameStrobe_O[2] ,
    \Tile_X1Y6_FrameStrobe_O[1] ,
    \Tile_X1Y6_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X1Y5_FrameStrobe_O[19] ,
    \Tile_X1Y5_FrameStrobe_O[18] ,
    \Tile_X1Y5_FrameStrobe_O[17] ,
    \Tile_X1Y5_FrameStrobe_O[16] ,
    \Tile_X1Y5_FrameStrobe_O[15] ,
    \Tile_X1Y5_FrameStrobe_O[14] ,
    \Tile_X1Y5_FrameStrobe_O[13] ,
    \Tile_X1Y5_FrameStrobe_O[12] ,
    \Tile_X1Y5_FrameStrobe_O[11] ,
    \Tile_X1Y5_FrameStrobe_O[10] ,
    \Tile_X1Y5_FrameStrobe_O[9] ,
    \Tile_X1Y5_FrameStrobe_O[8] ,
    \Tile_X1Y5_FrameStrobe_O[7] ,
    \Tile_X1Y5_FrameStrobe_O[6] ,
    \Tile_X1Y5_FrameStrobe_O[5] ,
    \Tile_X1Y5_FrameStrobe_O[4] ,
    \Tile_X1Y5_FrameStrobe_O[3] ,
    \Tile_X1Y5_FrameStrobe_O[2] ,
    \Tile_X1Y5_FrameStrobe_O[1] ,
    \Tile_X1Y5_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X1Y5_N1BEG[3] ,
    \Tile_X1Y5_N1BEG[2] ,
    \Tile_X1Y5_N1BEG[1] ,
    \Tile_X1Y5_N1BEG[0] }),
    .N1END({\Tile_X1Y6_N1BEG[3] ,
    \Tile_X1Y6_N1BEG[2] ,
    \Tile_X1Y6_N1BEG[1] ,
    \Tile_X1Y6_N1BEG[0] }),
    .N2BEG({\Tile_X1Y5_N2BEG[7] ,
    \Tile_X1Y5_N2BEG[6] ,
    \Tile_X1Y5_N2BEG[5] ,
    \Tile_X1Y5_N2BEG[4] ,
    \Tile_X1Y5_N2BEG[3] ,
    \Tile_X1Y5_N2BEG[2] ,
    \Tile_X1Y5_N2BEG[1] ,
    \Tile_X1Y5_N2BEG[0] }),
    .N2BEGb({\Tile_X1Y5_N2BEGb[7] ,
    \Tile_X1Y5_N2BEGb[6] ,
    \Tile_X1Y5_N2BEGb[5] ,
    \Tile_X1Y5_N2BEGb[4] ,
    \Tile_X1Y5_N2BEGb[3] ,
    \Tile_X1Y5_N2BEGb[2] ,
    \Tile_X1Y5_N2BEGb[1] ,
    \Tile_X1Y5_N2BEGb[0] }),
    .N2END({\Tile_X1Y6_N2BEGb[7] ,
    \Tile_X1Y6_N2BEGb[6] ,
    \Tile_X1Y6_N2BEGb[5] ,
    \Tile_X1Y6_N2BEGb[4] ,
    \Tile_X1Y6_N2BEGb[3] ,
    \Tile_X1Y6_N2BEGb[2] ,
    \Tile_X1Y6_N2BEGb[1] ,
    \Tile_X1Y6_N2BEGb[0] }),
    .N2MID({\Tile_X1Y6_N2BEG[7] ,
    \Tile_X1Y6_N2BEG[6] ,
    \Tile_X1Y6_N2BEG[5] ,
    \Tile_X1Y6_N2BEG[4] ,
    \Tile_X1Y6_N2BEG[3] ,
    \Tile_X1Y6_N2BEG[2] ,
    \Tile_X1Y6_N2BEG[1] ,
    \Tile_X1Y6_N2BEG[0] }),
    .N4BEG({\Tile_X1Y5_N4BEG[15] ,
    \Tile_X1Y5_N4BEG[14] ,
    \Tile_X1Y5_N4BEG[13] ,
    \Tile_X1Y5_N4BEG[12] ,
    \Tile_X1Y5_N4BEG[11] ,
    \Tile_X1Y5_N4BEG[10] ,
    \Tile_X1Y5_N4BEG[9] ,
    \Tile_X1Y5_N4BEG[8] ,
    \Tile_X1Y5_N4BEG[7] ,
    \Tile_X1Y5_N4BEG[6] ,
    \Tile_X1Y5_N4BEG[5] ,
    \Tile_X1Y5_N4BEG[4] ,
    \Tile_X1Y5_N4BEG[3] ,
    \Tile_X1Y5_N4BEG[2] ,
    \Tile_X1Y5_N4BEG[1] ,
    \Tile_X1Y5_N4BEG[0] }),
    .N4END({\Tile_X1Y6_N4BEG[15] ,
    \Tile_X1Y6_N4BEG[14] ,
    \Tile_X1Y6_N4BEG[13] ,
    \Tile_X1Y6_N4BEG[12] ,
    \Tile_X1Y6_N4BEG[11] ,
    \Tile_X1Y6_N4BEG[10] ,
    \Tile_X1Y6_N4BEG[9] ,
    \Tile_X1Y6_N4BEG[8] ,
    \Tile_X1Y6_N4BEG[7] ,
    \Tile_X1Y6_N4BEG[6] ,
    \Tile_X1Y6_N4BEG[5] ,
    \Tile_X1Y6_N4BEG[4] ,
    \Tile_X1Y6_N4BEG[3] ,
    \Tile_X1Y6_N4BEG[2] ,
    \Tile_X1Y6_N4BEG[1] ,
    \Tile_X1Y6_N4BEG[0] }),
    .NN4BEG({\Tile_X1Y5_NN4BEG[15] ,
    \Tile_X1Y5_NN4BEG[14] ,
    \Tile_X1Y5_NN4BEG[13] ,
    \Tile_X1Y5_NN4BEG[12] ,
    \Tile_X1Y5_NN4BEG[11] ,
    \Tile_X1Y5_NN4BEG[10] ,
    \Tile_X1Y5_NN4BEG[9] ,
    \Tile_X1Y5_NN4BEG[8] ,
    \Tile_X1Y5_NN4BEG[7] ,
    \Tile_X1Y5_NN4BEG[6] ,
    \Tile_X1Y5_NN4BEG[5] ,
    \Tile_X1Y5_NN4BEG[4] ,
    \Tile_X1Y5_NN4BEG[3] ,
    \Tile_X1Y5_NN4BEG[2] ,
    \Tile_X1Y5_NN4BEG[1] ,
    \Tile_X1Y5_NN4BEG[0] }),
    .NN4END({\Tile_X1Y6_NN4BEG[15] ,
    \Tile_X1Y6_NN4BEG[14] ,
    \Tile_X1Y6_NN4BEG[13] ,
    \Tile_X1Y6_NN4BEG[12] ,
    \Tile_X1Y6_NN4BEG[11] ,
    \Tile_X1Y6_NN4BEG[10] ,
    \Tile_X1Y6_NN4BEG[9] ,
    \Tile_X1Y6_NN4BEG[8] ,
    \Tile_X1Y6_NN4BEG[7] ,
    \Tile_X1Y6_NN4BEG[6] ,
    \Tile_X1Y6_NN4BEG[5] ,
    \Tile_X1Y6_NN4BEG[4] ,
    \Tile_X1Y6_NN4BEG[3] ,
    \Tile_X1Y6_NN4BEG[2] ,
    \Tile_X1Y6_NN4BEG[1] ,
    \Tile_X1Y6_NN4BEG[0] }),
    .S1BEG({\Tile_X1Y5_S1BEG[3] ,
    \Tile_X1Y5_S1BEG[2] ,
    \Tile_X1Y5_S1BEG[1] ,
    \Tile_X1Y5_S1BEG[0] }),
    .S1END({\Tile_X1Y4_S1BEG[3] ,
    \Tile_X1Y4_S1BEG[2] ,
    \Tile_X1Y4_S1BEG[1] ,
    \Tile_X1Y4_S1BEG[0] }),
    .S2BEG({\Tile_X1Y5_S2BEG[7] ,
    \Tile_X1Y5_S2BEG[6] ,
    \Tile_X1Y5_S2BEG[5] ,
    \Tile_X1Y5_S2BEG[4] ,
    \Tile_X1Y5_S2BEG[3] ,
    \Tile_X1Y5_S2BEG[2] ,
    \Tile_X1Y5_S2BEG[1] ,
    \Tile_X1Y5_S2BEG[0] }),
    .S2BEGb({\Tile_X1Y5_S2BEGb[7] ,
    \Tile_X1Y5_S2BEGb[6] ,
    \Tile_X1Y5_S2BEGb[5] ,
    \Tile_X1Y5_S2BEGb[4] ,
    \Tile_X1Y5_S2BEGb[3] ,
    \Tile_X1Y5_S2BEGb[2] ,
    \Tile_X1Y5_S2BEGb[1] ,
    \Tile_X1Y5_S2BEGb[0] }),
    .S2END({\Tile_X1Y4_S2BEGb[7] ,
    \Tile_X1Y4_S2BEGb[6] ,
    \Tile_X1Y4_S2BEGb[5] ,
    \Tile_X1Y4_S2BEGb[4] ,
    \Tile_X1Y4_S2BEGb[3] ,
    \Tile_X1Y4_S2BEGb[2] ,
    \Tile_X1Y4_S2BEGb[1] ,
    \Tile_X1Y4_S2BEGb[0] }),
    .S2MID({\Tile_X1Y4_S2BEG[7] ,
    \Tile_X1Y4_S2BEG[6] ,
    \Tile_X1Y4_S2BEG[5] ,
    \Tile_X1Y4_S2BEG[4] ,
    \Tile_X1Y4_S2BEG[3] ,
    \Tile_X1Y4_S2BEG[2] ,
    \Tile_X1Y4_S2BEG[1] ,
    \Tile_X1Y4_S2BEG[0] }),
    .S4BEG({\Tile_X1Y5_S4BEG[15] ,
    \Tile_X1Y5_S4BEG[14] ,
    \Tile_X1Y5_S4BEG[13] ,
    \Tile_X1Y5_S4BEG[12] ,
    \Tile_X1Y5_S4BEG[11] ,
    \Tile_X1Y5_S4BEG[10] ,
    \Tile_X1Y5_S4BEG[9] ,
    \Tile_X1Y5_S4BEG[8] ,
    \Tile_X1Y5_S4BEG[7] ,
    \Tile_X1Y5_S4BEG[6] ,
    \Tile_X1Y5_S4BEG[5] ,
    \Tile_X1Y5_S4BEG[4] ,
    \Tile_X1Y5_S4BEG[3] ,
    \Tile_X1Y5_S4BEG[2] ,
    \Tile_X1Y5_S4BEG[1] ,
    \Tile_X1Y5_S4BEG[0] }),
    .S4END({\Tile_X1Y4_S4BEG[15] ,
    \Tile_X1Y4_S4BEG[14] ,
    \Tile_X1Y4_S4BEG[13] ,
    \Tile_X1Y4_S4BEG[12] ,
    \Tile_X1Y4_S4BEG[11] ,
    \Tile_X1Y4_S4BEG[10] ,
    \Tile_X1Y4_S4BEG[9] ,
    \Tile_X1Y4_S4BEG[8] ,
    \Tile_X1Y4_S4BEG[7] ,
    \Tile_X1Y4_S4BEG[6] ,
    \Tile_X1Y4_S4BEG[5] ,
    \Tile_X1Y4_S4BEG[4] ,
    \Tile_X1Y4_S4BEG[3] ,
    \Tile_X1Y4_S4BEG[2] ,
    \Tile_X1Y4_S4BEG[1] ,
    \Tile_X1Y4_S4BEG[0] }),
    .SS4BEG({\Tile_X1Y5_SS4BEG[15] ,
    \Tile_X1Y5_SS4BEG[14] ,
    \Tile_X1Y5_SS4BEG[13] ,
    \Tile_X1Y5_SS4BEG[12] ,
    \Tile_X1Y5_SS4BEG[11] ,
    \Tile_X1Y5_SS4BEG[10] ,
    \Tile_X1Y5_SS4BEG[9] ,
    \Tile_X1Y5_SS4BEG[8] ,
    \Tile_X1Y5_SS4BEG[7] ,
    \Tile_X1Y5_SS4BEG[6] ,
    \Tile_X1Y5_SS4BEG[5] ,
    \Tile_X1Y5_SS4BEG[4] ,
    \Tile_X1Y5_SS4BEG[3] ,
    \Tile_X1Y5_SS4BEG[2] ,
    \Tile_X1Y5_SS4BEG[1] ,
    \Tile_X1Y5_SS4BEG[0] }),
    .SS4END({\Tile_X1Y4_SS4BEG[15] ,
    \Tile_X1Y4_SS4BEG[14] ,
    \Tile_X1Y4_SS4BEG[13] ,
    \Tile_X1Y4_SS4BEG[12] ,
    \Tile_X1Y4_SS4BEG[11] ,
    \Tile_X1Y4_SS4BEG[10] ,
    \Tile_X1Y4_SS4BEG[9] ,
    \Tile_X1Y4_SS4BEG[8] ,
    \Tile_X1Y4_SS4BEG[7] ,
    \Tile_X1Y4_SS4BEG[6] ,
    \Tile_X1Y4_SS4BEG[5] ,
    \Tile_X1Y4_SS4BEG[4] ,
    \Tile_X1Y4_SS4BEG[3] ,
    \Tile_X1Y4_SS4BEG[2] ,
    \Tile_X1Y4_SS4BEG[1] ,
    \Tile_X1Y4_SS4BEG[0] }),
    .W1BEG({\Tile_X1Y5_W1BEG[3] ,
    \Tile_X1Y5_W1BEG[2] ,
    \Tile_X1Y5_W1BEG[1] ,
    \Tile_X1Y5_W1BEG[0] }),
    .W1END({\Tile_X2Y5_W1BEG[3] ,
    \Tile_X2Y5_W1BEG[2] ,
    \Tile_X2Y5_W1BEG[1] ,
    \Tile_X2Y5_W1BEG[0] }),
    .W2BEG({\Tile_X1Y5_W2BEG[7] ,
    \Tile_X1Y5_W2BEG[6] ,
    \Tile_X1Y5_W2BEG[5] ,
    \Tile_X1Y5_W2BEG[4] ,
    \Tile_X1Y5_W2BEG[3] ,
    \Tile_X1Y5_W2BEG[2] ,
    \Tile_X1Y5_W2BEG[1] ,
    \Tile_X1Y5_W2BEG[0] }),
    .W2BEGb({\Tile_X1Y5_W2BEGb[7] ,
    \Tile_X1Y5_W2BEGb[6] ,
    \Tile_X1Y5_W2BEGb[5] ,
    \Tile_X1Y5_W2BEGb[4] ,
    \Tile_X1Y5_W2BEGb[3] ,
    \Tile_X1Y5_W2BEGb[2] ,
    \Tile_X1Y5_W2BEGb[1] ,
    \Tile_X1Y5_W2BEGb[0] }),
    .W2END({\Tile_X2Y5_W2BEGb[7] ,
    \Tile_X2Y5_W2BEGb[6] ,
    \Tile_X2Y5_W2BEGb[5] ,
    \Tile_X2Y5_W2BEGb[4] ,
    \Tile_X2Y5_W2BEGb[3] ,
    \Tile_X2Y5_W2BEGb[2] ,
    \Tile_X2Y5_W2BEGb[1] ,
    \Tile_X2Y5_W2BEGb[0] }),
    .W2MID({\Tile_X2Y5_W2BEG[7] ,
    \Tile_X2Y5_W2BEG[6] ,
    \Tile_X2Y5_W2BEG[5] ,
    \Tile_X2Y5_W2BEG[4] ,
    \Tile_X2Y5_W2BEG[3] ,
    \Tile_X2Y5_W2BEG[2] ,
    \Tile_X2Y5_W2BEG[1] ,
    \Tile_X2Y5_W2BEG[0] }),
    .W6BEG({\Tile_X1Y5_W6BEG[11] ,
    \Tile_X1Y5_W6BEG[10] ,
    \Tile_X1Y5_W6BEG[9] ,
    \Tile_X1Y5_W6BEG[8] ,
    \Tile_X1Y5_W6BEG[7] ,
    \Tile_X1Y5_W6BEG[6] ,
    \Tile_X1Y5_W6BEG[5] ,
    \Tile_X1Y5_W6BEG[4] ,
    \Tile_X1Y5_W6BEG[3] ,
    \Tile_X1Y5_W6BEG[2] ,
    \Tile_X1Y5_W6BEG[1] ,
    \Tile_X1Y5_W6BEG[0] }),
    .W6END({\Tile_X2Y5_W6BEG[11] ,
    \Tile_X2Y5_W6BEG[10] ,
    \Tile_X2Y5_W6BEG[9] ,
    \Tile_X2Y5_W6BEG[8] ,
    \Tile_X2Y5_W6BEG[7] ,
    \Tile_X2Y5_W6BEG[6] ,
    \Tile_X2Y5_W6BEG[5] ,
    \Tile_X2Y5_W6BEG[4] ,
    \Tile_X2Y5_W6BEG[3] ,
    \Tile_X2Y5_W6BEG[2] ,
    \Tile_X2Y5_W6BEG[1] ,
    \Tile_X2Y5_W6BEG[0] }),
    .WW4BEG({\Tile_X1Y5_WW4BEG[15] ,
    \Tile_X1Y5_WW4BEG[14] ,
    \Tile_X1Y5_WW4BEG[13] ,
    \Tile_X1Y5_WW4BEG[12] ,
    \Tile_X1Y5_WW4BEG[11] ,
    \Tile_X1Y5_WW4BEG[10] ,
    \Tile_X1Y5_WW4BEG[9] ,
    \Tile_X1Y5_WW4BEG[8] ,
    \Tile_X1Y5_WW4BEG[7] ,
    \Tile_X1Y5_WW4BEG[6] ,
    \Tile_X1Y5_WW4BEG[5] ,
    \Tile_X1Y5_WW4BEG[4] ,
    \Tile_X1Y5_WW4BEG[3] ,
    \Tile_X1Y5_WW4BEG[2] ,
    \Tile_X1Y5_WW4BEG[1] ,
    \Tile_X1Y5_WW4BEG[0] }),
    .WW4END({\Tile_X2Y5_WW4BEG[15] ,
    \Tile_X2Y5_WW4BEG[14] ,
    \Tile_X2Y5_WW4BEG[13] ,
    \Tile_X2Y5_WW4BEG[12] ,
    \Tile_X2Y5_WW4BEG[11] ,
    \Tile_X2Y5_WW4BEG[10] ,
    \Tile_X2Y5_WW4BEG[9] ,
    \Tile_X2Y5_WW4BEG[8] ,
    \Tile_X2Y5_WW4BEG[7] ,
    \Tile_X2Y5_WW4BEG[6] ,
    \Tile_X2Y5_WW4BEG[5] ,
    \Tile_X2Y5_WW4BEG[4] ,
    \Tile_X2Y5_WW4BEG[3] ,
    \Tile_X2Y5_WW4BEG[2] ,
    \Tile_X2Y5_WW4BEG[1] ,
    \Tile_X2Y5_WW4BEG[0] }));
 LUT4AB Tile_X1Y6_LUT4AB (.Ci(Tile_X1Y7_Co),
    .Co(Tile_X1Y6_Co),
    .UserCLK(Tile_X1Y7_UserCLKo),
    .UserCLKo(Tile_X1Y6_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X1Y6_E1BEG[3] ,
    \Tile_X1Y6_E1BEG[2] ,
    \Tile_X1Y6_E1BEG[1] ,
    \Tile_X1Y6_E1BEG[0] }),
    .E1END({\Tile_X0Y6_E1BEG[3] ,
    \Tile_X0Y6_E1BEG[2] ,
    \Tile_X0Y6_E1BEG[1] ,
    \Tile_X0Y6_E1BEG[0] }),
    .E2BEG({\Tile_X1Y6_E2BEG[7] ,
    \Tile_X1Y6_E2BEG[6] ,
    \Tile_X1Y6_E2BEG[5] ,
    \Tile_X1Y6_E2BEG[4] ,
    \Tile_X1Y6_E2BEG[3] ,
    \Tile_X1Y6_E2BEG[2] ,
    \Tile_X1Y6_E2BEG[1] ,
    \Tile_X1Y6_E2BEG[0] }),
    .E2BEGb({\Tile_X1Y6_E2BEGb[7] ,
    \Tile_X1Y6_E2BEGb[6] ,
    \Tile_X1Y6_E2BEGb[5] ,
    \Tile_X1Y6_E2BEGb[4] ,
    \Tile_X1Y6_E2BEGb[3] ,
    \Tile_X1Y6_E2BEGb[2] ,
    \Tile_X1Y6_E2BEGb[1] ,
    \Tile_X1Y6_E2BEGb[0] }),
    .E2END({\Tile_X0Y6_E2BEGb[7] ,
    \Tile_X0Y6_E2BEGb[6] ,
    \Tile_X0Y6_E2BEGb[5] ,
    \Tile_X0Y6_E2BEGb[4] ,
    \Tile_X0Y6_E2BEGb[3] ,
    \Tile_X0Y6_E2BEGb[2] ,
    \Tile_X0Y6_E2BEGb[1] ,
    \Tile_X0Y6_E2BEGb[0] }),
    .E2MID({\Tile_X0Y6_E2BEG[7] ,
    \Tile_X0Y6_E2BEG[6] ,
    \Tile_X0Y6_E2BEG[5] ,
    \Tile_X0Y6_E2BEG[4] ,
    \Tile_X0Y6_E2BEG[3] ,
    \Tile_X0Y6_E2BEG[2] ,
    \Tile_X0Y6_E2BEG[1] ,
    \Tile_X0Y6_E2BEG[0] }),
    .E6BEG({\Tile_X1Y6_E6BEG[11] ,
    \Tile_X1Y6_E6BEG[10] ,
    \Tile_X1Y6_E6BEG[9] ,
    \Tile_X1Y6_E6BEG[8] ,
    \Tile_X1Y6_E6BEG[7] ,
    \Tile_X1Y6_E6BEG[6] ,
    \Tile_X1Y6_E6BEG[5] ,
    \Tile_X1Y6_E6BEG[4] ,
    \Tile_X1Y6_E6BEG[3] ,
    \Tile_X1Y6_E6BEG[2] ,
    \Tile_X1Y6_E6BEG[1] ,
    \Tile_X1Y6_E6BEG[0] }),
    .E6END({\Tile_X0Y6_E6BEG[11] ,
    \Tile_X0Y6_E6BEG[10] ,
    \Tile_X0Y6_E6BEG[9] ,
    \Tile_X0Y6_E6BEG[8] ,
    \Tile_X0Y6_E6BEG[7] ,
    \Tile_X0Y6_E6BEG[6] ,
    \Tile_X0Y6_E6BEG[5] ,
    \Tile_X0Y6_E6BEG[4] ,
    \Tile_X0Y6_E6BEG[3] ,
    \Tile_X0Y6_E6BEG[2] ,
    \Tile_X0Y6_E6BEG[1] ,
    \Tile_X0Y6_E6BEG[0] }),
    .EE4BEG({\Tile_X1Y6_EE4BEG[15] ,
    \Tile_X1Y6_EE4BEG[14] ,
    \Tile_X1Y6_EE4BEG[13] ,
    \Tile_X1Y6_EE4BEG[12] ,
    \Tile_X1Y6_EE4BEG[11] ,
    \Tile_X1Y6_EE4BEG[10] ,
    \Tile_X1Y6_EE4BEG[9] ,
    \Tile_X1Y6_EE4BEG[8] ,
    \Tile_X1Y6_EE4BEG[7] ,
    \Tile_X1Y6_EE4BEG[6] ,
    \Tile_X1Y6_EE4BEG[5] ,
    \Tile_X1Y6_EE4BEG[4] ,
    \Tile_X1Y6_EE4BEG[3] ,
    \Tile_X1Y6_EE4BEG[2] ,
    \Tile_X1Y6_EE4BEG[1] ,
    \Tile_X1Y6_EE4BEG[0] }),
    .EE4END({\Tile_X0Y6_EE4BEG[15] ,
    \Tile_X0Y6_EE4BEG[14] ,
    \Tile_X0Y6_EE4BEG[13] ,
    \Tile_X0Y6_EE4BEG[12] ,
    \Tile_X0Y6_EE4BEG[11] ,
    \Tile_X0Y6_EE4BEG[10] ,
    \Tile_X0Y6_EE4BEG[9] ,
    \Tile_X0Y6_EE4BEG[8] ,
    \Tile_X0Y6_EE4BEG[7] ,
    \Tile_X0Y6_EE4BEG[6] ,
    \Tile_X0Y6_EE4BEG[5] ,
    \Tile_X0Y6_EE4BEG[4] ,
    \Tile_X0Y6_EE4BEG[3] ,
    \Tile_X0Y6_EE4BEG[2] ,
    \Tile_X0Y6_EE4BEG[1] ,
    \Tile_X0Y6_EE4BEG[0] }),
    .FrameData({\Tile_X0Y6_FrameData_O[31] ,
    \Tile_X0Y6_FrameData_O[30] ,
    \Tile_X0Y6_FrameData_O[29] ,
    \Tile_X0Y6_FrameData_O[28] ,
    \Tile_X0Y6_FrameData_O[27] ,
    \Tile_X0Y6_FrameData_O[26] ,
    \Tile_X0Y6_FrameData_O[25] ,
    \Tile_X0Y6_FrameData_O[24] ,
    \Tile_X0Y6_FrameData_O[23] ,
    \Tile_X0Y6_FrameData_O[22] ,
    \Tile_X0Y6_FrameData_O[21] ,
    \Tile_X0Y6_FrameData_O[20] ,
    \Tile_X0Y6_FrameData_O[19] ,
    \Tile_X0Y6_FrameData_O[18] ,
    \Tile_X0Y6_FrameData_O[17] ,
    \Tile_X0Y6_FrameData_O[16] ,
    \Tile_X0Y6_FrameData_O[15] ,
    \Tile_X0Y6_FrameData_O[14] ,
    \Tile_X0Y6_FrameData_O[13] ,
    \Tile_X0Y6_FrameData_O[12] ,
    \Tile_X0Y6_FrameData_O[11] ,
    \Tile_X0Y6_FrameData_O[10] ,
    \Tile_X0Y6_FrameData_O[9] ,
    \Tile_X0Y6_FrameData_O[8] ,
    \Tile_X0Y6_FrameData_O[7] ,
    \Tile_X0Y6_FrameData_O[6] ,
    \Tile_X0Y6_FrameData_O[5] ,
    \Tile_X0Y6_FrameData_O[4] ,
    \Tile_X0Y6_FrameData_O[3] ,
    \Tile_X0Y6_FrameData_O[2] ,
    \Tile_X0Y6_FrameData_O[1] ,
    \Tile_X0Y6_FrameData_O[0] }),
    .FrameData_O({\Tile_X1Y6_FrameData_O[31] ,
    \Tile_X1Y6_FrameData_O[30] ,
    \Tile_X1Y6_FrameData_O[29] ,
    \Tile_X1Y6_FrameData_O[28] ,
    \Tile_X1Y6_FrameData_O[27] ,
    \Tile_X1Y6_FrameData_O[26] ,
    \Tile_X1Y6_FrameData_O[25] ,
    \Tile_X1Y6_FrameData_O[24] ,
    \Tile_X1Y6_FrameData_O[23] ,
    \Tile_X1Y6_FrameData_O[22] ,
    \Tile_X1Y6_FrameData_O[21] ,
    \Tile_X1Y6_FrameData_O[20] ,
    \Tile_X1Y6_FrameData_O[19] ,
    \Tile_X1Y6_FrameData_O[18] ,
    \Tile_X1Y6_FrameData_O[17] ,
    \Tile_X1Y6_FrameData_O[16] ,
    \Tile_X1Y6_FrameData_O[15] ,
    \Tile_X1Y6_FrameData_O[14] ,
    \Tile_X1Y6_FrameData_O[13] ,
    \Tile_X1Y6_FrameData_O[12] ,
    \Tile_X1Y6_FrameData_O[11] ,
    \Tile_X1Y6_FrameData_O[10] ,
    \Tile_X1Y6_FrameData_O[9] ,
    \Tile_X1Y6_FrameData_O[8] ,
    \Tile_X1Y6_FrameData_O[7] ,
    \Tile_X1Y6_FrameData_O[6] ,
    \Tile_X1Y6_FrameData_O[5] ,
    \Tile_X1Y6_FrameData_O[4] ,
    \Tile_X1Y6_FrameData_O[3] ,
    \Tile_X1Y6_FrameData_O[2] ,
    \Tile_X1Y6_FrameData_O[1] ,
    \Tile_X1Y6_FrameData_O[0] }),
    .FrameStrobe({\Tile_X1Y7_FrameStrobe_O[19] ,
    \Tile_X1Y7_FrameStrobe_O[18] ,
    \Tile_X1Y7_FrameStrobe_O[17] ,
    \Tile_X1Y7_FrameStrobe_O[16] ,
    \Tile_X1Y7_FrameStrobe_O[15] ,
    \Tile_X1Y7_FrameStrobe_O[14] ,
    \Tile_X1Y7_FrameStrobe_O[13] ,
    \Tile_X1Y7_FrameStrobe_O[12] ,
    \Tile_X1Y7_FrameStrobe_O[11] ,
    \Tile_X1Y7_FrameStrobe_O[10] ,
    \Tile_X1Y7_FrameStrobe_O[9] ,
    \Tile_X1Y7_FrameStrobe_O[8] ,
    \Tile_X1Y7_FrameStrobe_O[7] ,
    \Tile_X1Y7_FrameStrobe_O[6] ,
    \Tile_X1Y7_FrameStrobe_O[5] ,
    \Tile_X1Y7_FrameStrobe_O[4] ,
    \Tile_X1Y7_FrameStrobe_O[3] ,
    \Tile_X1Y7_FrameStrobe_O[2] ,
    \Tile_X1Y7_FrameStrobe_O[1] ,
    \Tile_X1Y7_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X1Y6_FrameStrobe_O[19] ,
    \Tile_X1Y6_FrameStrobe_O[18] ,
    \Tile_X1Y6_FrameStrobe_O[17] ,
    \Tile_X1Y6_FrameStrobe_O[16] ,
    \Tile_X1Y6_FrameStrobe_O[15] ,
    \Tile_X1Y6_FrameStrobe_O[14] ,
    \Tile_X1Y6_FrameStrobe_O[13] ,
    \Tile_X1Y6_FrameStrobe_O[12] ,
    \Tile_X1Y6_FrameStrobe_O[11] ,
    \Tile_X1Y6_FrameStrobe_O[10] ,
    \Tile_X1Y6_FrameStrobe_O[9] ,
    \Tile_X1Y6_FrameStrobe_O[8] ,
    \Tile_X1Y6_FrameStrobe_O[7] ,
    \Tile_X1Y6_FrameStrobe_O[6] ,
    \Tile_X1Y6_FrameStrobe_O[5] ,
    \Tile_X1Y6_FrameStrobe_O[4] ,
    \Tile_X1Y6_FrameStrobe_O[3] ,
    \Tile_X1Y6_FrameStrobe_O[2] ,
    \Tile_X1Y6_FrameStrobe_O[1] ,
    \Tile_X1Y6_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X1Y6_N1BEG[3] ,
    \Tile_X1Y6_N1BEG[2] ,
    \Tile_X1Y6_N1BEG[1] ,
    \Tile_X1Y6_N1BEG[0] }),
    .N1END({\Tile_X1Y7_N1BEG[3] ,
    \Tile_X1Y7_N1BEG[2] ,
    \Tile_X1Y7_N1BEG[1] ,
    \Tile_X1Y7_N1BEG[0] }),
    .N2BEG({\Tile_X1Y6_N2BEG[7] ,
    \Tile_X1Y6_N2BEG[6] ,
    \Tile_X1Y6_N2BEG[5] ,
    \Tile_X1Y6_N2BEG[4] ,
    \Tile_X1Y6_N2BEG[3] ,
    \Tile_X1Y6_N2BEG[2] ,
    \Tile_X1Y6_N2BEG[1] ,
    \Tile_X1Y6_N2BEG[0] }),
    .N2BEGb({\Tile_X1Y6_N2BEGb[7] ,
    \Tile_X1Y6_N2BEGb[6] ,
    \Tile_X1Y6_N2BEGb[5] ,
    \Tile_X1Y6_N2BEGb[4] ,
    \Tile_X1Y6_N2BEGb[3] ,
    \Tile_X1Y6_N2BEGb[2] ,
    \Tile_X1Y6_N2BEGb[1] ,
    \Tile_X1Y6_N2BEGb[0] }),
    .N2END({\Tile_X1Y7_N2BEGb[7] ,
    \Tile_X1Y7_N2BEGb[6] ,
    \Tile_X1Y7_N2BEGb[5] ,
    \Tile_X1Y7_N2BEGb[4] ,
    \Tile_X1Y7_N2BEGb[3] ,
    \Tile_X1Y7_N2BEGb[2] ,
    \Tile_X1Y7_N2BEGb[1] ,
    \Tile_X1Y7_N2BEGb[0] }),
    .N2MID({\Tile_X1Y7_N2BEG[7] ,
    \Tile_X1Y7_N2BEG[6] ,
    \Tile_X1Y7_N2BEG[5] ,
    \Tile_X1Y7_N2BEG[4] ,
    \Tile_X1Y7_N2BEG[3] ,
    \Tile_X1Y7_N2BEG[2] ,
    \Tile_X1Y7_N2BEG[1] ,
    \Tile_X1Y7_N2BEG[0] }),
    .N4BEG({\Tile_X1Y6_N4BEG[15] ,
    \Tile_X1Y6_N4BEG[14] ,
    \Tile_X1Y6_N4BEG[13] ,
    \Tile_X1Y6_N4BEG[12] ,
    \Tile_X1Y6_N4BEG[11] ,
    \Tile_X1Y6_N4BEG[10] ,
    \Tile_X1Y6_N4BEG[9] ,
    \Tile_X1Y6_N4BEG[8] ,
    \Tile_X1Y6_N4BEG[7] ,
    \Tile_X1Y6_N4BEG[6] ,
    \Tile_X1Y6_N4BEG[5] ,
    \Tile_X1Y6_N4BEG[4] ,
    \Tile_X1Y6_N4BEG[3] ,
    \Tile_X1Y6_N4BEG[2] ,
    \Tile_X1Y6_N4BEG[1] ,
    \Tile_X1Y6_N4BEG[0] }),
    .N4END({\Tile_X1Y7_N4BEG[15] ,
    \Tile_X1Y7_N4BEG[14] ,
    \Tile_X1Y7_N4BEG[13] ,
    \Tile_X1Y7_N4BEG[12] ,
    \Tile_X1Y7_N4BEG[11] ,
    \Tile_X1Y7_N4BEG[10] ,
    \Tile_X1Y7_N4BEG[9] ,
    \Tile_X1Y7_N4BEG[8] ,
    \Tile_X1Y7_N4BEG[7] ,
    \Tile_X1Y7_N4BEG[6] ,
    \Tile_X1Y7_N4BEG[5] ,
    \Tile_X1Y7_N4BEG[4] ,
    \Tile_X1Y7_N4BEG[3] ,
    \Tile_X1Y7_N4BEG[2] ,
    \Tile_X1Y7_N4BEG[1] ,
    \Tile_X1Y7_N4BEG[0] }),
    .NN4BEG({\Tile_X1Y6_NN4BEG[15] ,
    \Tile_X1Y6_NN4BEG[14] ,
    \Tile_X1Y6_NN4BEG[13] ,
    \Tile_X1Y6_NN4BEG[12] ,
    \Tile_X1Y6_NN4BEG[11] ,
    \Tile_X1Y6_NN4BEG[10] ,
    \Tile_X1Y6_NN4BEG[9] ,
    \Tile_X1Y6_NN4BEG[8] ,
    \Tile_X1Y6_NN4BEG[7] ,
    \Tile_X1Y6_NN4BEG[6] ,
    \Tile_X1Y6_NN4BEG[5] ,
    \Tile_X1Y6_NN4BEG[4] ,
    \Tile_X1Y6_NN4BEG[3] ,
    \Tile_X1Y6_NN4BEG[2] ,
    \Tile_X1Y6_NN4BEG[1] ,
    \Tile_X1Y6_NN4BEG[0] }),
    .NN4END({\Tile_X1Y7_NN4BEG[15] ,
    \Tile_X1Y7_NN4BEG[14] ,
    \Tile_X1Y7_NN4BEG[13] ,
    \Tile_X1Y7_NN4BEG[12] ,
    \Tile_X1Y7_NN4BEG[11] ,
    \Tile_X1Y7_NN4BEG[10] ,
    \Tile_X1Y7_NN4BEG[9] ,
    \Tile_X1Y7_NN4BEG[8] ,
    \Tile_X1Y7_NN4BEG[7] ,
    \Tile_X1Y7_NN4BEG[6] ,
    \Tile_X1Y7_NN4BEG[5] ,
    \Tile_X1Y7_NN4BEG[4] ,
    \Tile_X1Y7_NN4BEG[3] ,
    \Tile_X1Y7_NN4BEG[2] ,
    \Tile_X1Y7_NN4BEG[1] ,
    \Tile_X1Y7_NN4BEG[0] }),
    .S1BEG({\Tile_X1Y6_S1BEG[3] ,
    \Tile_X1Y6_S1BEG[2] ,
    \Tile_X1Y6_S1BEG[1] ,
    \Tile_X1Y6_S1BEG[0] }),
    .S1END({\Tile_X1Y5_S1BEG[3] ,
    \Tile_X1Y5_S1BEG[2] ,
    \Tile_X1Y5_S1BEG[1] ,
    \Tile_X1Y5_S1BEG[0] }),
    .S2BEG({\Tile_X1Y6_S2BEG[7] ,
    \Tile_X1Y6_S2BEG[6] ,
    \Tile_X1Y6_S2BEG[5] ,
    \Tile_X1Y6_S2BEG[4] ,
    \Tile_X1Y6_S2BEG[3] ,
    \Tile_X1Y6_S2BEG[2] ,
    \Tile_X1Y6_S2BEG[1] ,
    \Tile_X1Y6_S2BEG[0] }),
    .S2BEGb({\Tile_X1Y6_S2BEGb[7] ,
    \Tile_X1Y6_S2BEGb[6] ,
    \Tile_X1Y6_S2BEGb[5] ,
    \Tile_X1Y6_S2BEGb[4] ,
    \Tile_X1Y6_S2BEGb[3] ,
    \Tile_X1Y6_S2BEGb[2] ,
    \Tile_X1Y6_S2BEGb[1] ,
    \Tile_X1Y6_S2BEGb[0] }),
    .S2END({\Tile_X1Y5_S2BEGb[7] ,
    \Tile_X1Y5_S2BEGb[6] ,
    \Tile_X1Y5_S2BEGb[5] ,
    \Tile_X1Y5_S2BEGb[4] ,
    \Tile_X1Y5_S2BEGb[3] ,
    \Tile_X1Y5_S2BEGb[2] ,
    \Tile_X1Y5_S2BEGb[1] ,
    \Tile_X1Y5_S2BEGb[0] }),
    .S2MID({\Tile_X1Y5_S2BEG[7] ,
    \Tile_X1Y5_S2BEG[6] ,
    \Tile_X1Y5_S2BEG[5] ,
    \Tile_X1Y5_S2BEG[4] ,
    \Tile_X1Y5_S2BEG[3] ,
    \Tile_X1Y5_S2BEG[2] ,
    \Tile_X1Y5_S2BEG[1] ,
    \Tile_X1Y5_S2BEG[0] }),
    .S4BEG({\Tile_X1Y6_S4BEG[15] ,
    \Tile_X1Y6_S4BEG[14] ,
    \Tile_X1Y6_S4BEG[13] ,
    \Tile_X1Y6_S4BEG[12] ,
    \Tile_X1Y6_S4BEG[11] ,
    \Tile_X1Y6_S4BEG[10] ,
    \Tile_X1Y6_S4BEG[9] ,
    \Tile_X1Y6_S4BEG[8] ,
    \Tile_X1Y6_S4BEG[7] ,
    \Tile_X1Y6_S4BEG[6] ,
    \Tile_X1Y6_S4BEG[5] ,
    \Tile_X1Y6_S4BEG[4] ,
    \Tile_X1Y6_S4BEG[3] ,
    \Tile_X1Y6_S4BEG[2] ,
    \Tile_X1Y6_S4BEG[1] ,
    \Tile_X1Y6_S4BEG[0] }),
    .S4END({\Tile_X1Y5_S4BEG[15] ,
    \Tile_X1Y5_S4BEG[14] ,
    \Tile_X1Y5_S4BEG[13] ,
    \Tile_X1Y5_S4BEG[12] ,
    \Tile_X1Y5_S4BEG[11] ,
    \Tile_X1Y5_S4BEG[10] ,
    \Tile_X1Y5_S4BEG[9] ,
    \Tile_X1Y5_S4BEG[8] ,
    \Tile_X1Y5_S4BEG[7] ,
    \Tile_X1Y5_S4BEG[6] ,
    \Tile_X1Y5_S4BEG[5] ,
    \Tile_X1Y5_S4BEG[4] ,
    \Tile_X1Y5_S4BEG[3] ,
    \Tile_X1Y5_S4BEG[2] ,
    \Tile_X1Y5_S4BEG[1] ,
    \Tile_X1Y5_S4BEG[0] }),
    .SS4BEG({\Tile_X1Y6_SS4BEG[15] ,
    \Tile_X1Y6_SS4BEG[14] ,
    \Tile_X1Y6_SS4BEG[13] ,
    \Tile_X1Y6_SS4BEG[12] ,
    \Tile_X1Y6_SS4BEG[11] ,
    \Tile_X1Y6_SS4BEG[10] ,
    \Tile_X1Y6_SS4BEG[9] ,
    \Tile_X1Y6_SS4BEG[8] ,
    \Tile_X1Y6_SS4BEG[7] ,
    \Tile_X1Y6_SS4BEG[6] ,
    \Tile_X1Y6_SS4BEG[5] ,
    \Tile_X1Y6_SS4BEG[4] ,
    \Tile_X1Y6_SS4BEG[3] ,
    \Tile_X1Y6_SS4BEG[2] ,
    \Tile_X1Y6_SS4BEG[1] ,
    \Tile_X1Y6_SS4BEG[0] }),
    .SS4END({\Tile_X1Y5_SS4BEG[15] ,
    \Tile_X1Y5_SS4BEG[14] ,
    \Tile_X1Y5_SS4BEG[13] ,
    \Tile_X1Y5_SS4BEG[12] ,
    \Tile_X1Y5_SS4BEG[11] ,
    \Tile_X1Y5_SS4BEG[10] ,
    \Tile_X1Y5_SS4BEG[9] ,
    \Tile_X1Y5_SS4BEG[8] ,
    \Tile_X1Y5_SS4BEG[7] ,
    \Tile_X1Y5_SS4BEG[6] ,
    \Tile_X1Y5_SS4BEG[5] ,
    \Tile_X1Y5_SS4BEG[4] ,
    \Tile_X1Y5_SS4BEG[3] ,
    \Tile_X1Y5_SS4BEG[2] ,
    \Tile_X1Y5_SS4BEG[1] ,
    \Tile_X1Y5_SS4BEG[0] }),
    .W1BEG({\Tile_X1Y6_W1BEG[3] ,
    \Tile_X1Y6_W1BEG[2] ,
    \Tile_X1Y6_W1BEG[1] ,
    \Tile_X1Y6_W1BEG[0] }),
    .W1END({\Tile_X2Y6_W1BEG[3] ,
    \Tile_X2Y6_W1BEG[2] ,
    \Tile_X2Y6_W1BEG[1] ,
    \Tile_X2Y6_W1BEG[0] }),
    .W2BEG({\Tile_X1Y6_W2BEG[7] ,
    \Tile_X1Y6_W2BEG[6] ,
    \Tile_X1Y6_W2BEG[5] ,
    \Tile_X1Y6_W2BEG[4] ,
    \Tile_X1Y6_W2BEG[3] ,
    \Tile_X1Y6_W2BEG[2] ,
    \Tile_X1Y6_W2BEG[1] ,
    \Tile_X1Y6_W2BEG[0] }),
    .W2BEGb({\Tile_X1Y6_W2BEGb[7] ,
    \Tile_X1Y6_W2BEGb[6] ,
    \Tile_X1Y6_W2BEGb[5] ,
    \Tile_X1Y6_W2BEGb[4] ,
    \Tile_X1Y6_W2BEGb[3] ,
    \Tile_X1Y6_W2BEGb[2] ,
    \Tile_X1Y6_W2BEGb[1] ,
    \Tile_X1Y6_W2BEGb[0] }),
    .W2END({\Tile_X2Y6_W2BEGb[7] ,
    \Tile_X2Y6_W2BEGb[6] ,
    \Tile_X2Y6_W2BEGb[5] ,
    \Tile_X2Y6_W2BEGb[4] ,
    \Tile_X2Y6_W2BEGb[3] ,
    \Tile_X2Y6_W2BEGb[2] ,
    \Tile_X2Y6_W2BEGb[1] ,
    \Tile_X2Y6_W2BEGb[0] }),
    .W2MID({\Tile_X2Y6_W2BEG[7] ,
    \Tile_X2Y6_W2BEG[6] ,
    \Tile_X2Y6_W2BEG[5] ,
    \Tile_X2Y6_W2BEG[4] ,
    \Tile_X2Y6_W2BEG[3] ,
    \Tile_X2Y6_W2BEG[2] ,
    \Tile_X2Y6_W2BEG[1] ,
    \Tile_X2Y6_W2BEG[0] }),
    .W6BEG({\Tile_X1Y6_W6BEG[11] ,
    \Tile_X1Y6_W6BEG[10] ,
    \Tile_X1Y6_W6BEG[9] ,
    \Tile_X1Y6_W6BEG[8] ,
    \Tile_X1Y6_W6BEG[7] ,
    \Tile_X1Y6_W6BEG[6] ,
    \Tile_X1Y6_W6BEG[5] ,
    \Tile_X1Y6_W6BEG[4] ,
    \Tile_X1Y6_W6BEG[3] ,
    \Tile_X1Y6_W6BEG[2] ,
    \Tile_X1Y6_W6BEG[1] ,
    \Tile_X1Y6_W6BEG[0] }),
    .W6END({\Tile_X2Y6_W6BEG[11] ,
    \Tile_X2Y6_W6BEG[10] ,
    \Tile_X2Y6_W6BEG[9] ,
    \Tile_X2Y6_W6BEG[8] ,
    \Tile_X2Y6_W6BEG[7] ,
    \Tile_X2Y6_W6BEG[6] ,
    \Tile_X2Y6_W6BEG[5] ,
    \Tile_X2Y6_W6BEG[4] ,
    \Tile_X2Y6_W6BEG[3] ,
    \Tile_X2Y6_W6BEG[2] ,
    \Tile_X2Y6_W6BEG[1] ,
    \Tile_X2Y6_W6BEG[0] }),
    .WW4BEG({\Tile_X1Y6_WW4BEG[15] ,
    \Tile_X1Y6_WW4BEG[14] ,
    \Tile_X1Y6_WW4BEG[13] ,
    \Tile_X1Y6_WW4BEG[12] ,
    \Tile_X1Y6_WW4BEG[11] ,
    \Tile_X1Y6_WW4BEG[10] ,
    \Tile_X1Y6_WW4BEG[9] ,
    \Tile_X1Y6_WW4BEG[8] ,
    \Tile_X1Y6_WW4BEG[7] ,
    \Tile_X1Y6_WW4BEG[6] ,
    \Tile_X1Y6_WW4BEG[5] ,
    \Tile_X1Y6_WW4BEG[4] ,
    \Tile_X1Y6_WW4BEG[3] ,
    \Tile_X1Y6_WW4BEG[2] ,
    \Tile_X1Y6_WW4BEG[1] ,
    \Tile_X1Y6_WW4BEG[0] }),
    .WW4END({\Tile_X2Y6_WW4BEG[15] ,
    \Tile_X2Y6_WW4BEG[14] ,
    \Tile_X2Y6_WW4BEG[13] ,
    \Tile_X2Y6_WW4BEG[12] ,
    \Tile_X2Y6_WW4BEG[11] ,
    \Tile_X2Y6_WW4BEG[10] ,
    \Tile_X2Y6_WW4BEG[9] ,
    \Tile_X2Y6_WW4BEG[8] ,
    \Tile_X2Y6_WW4BEG[7] ,
    \Tile_X2Y6_WW4BEG[6] ,
    \Tile_X2Y6_WW4BEG[5] ,
    \Tile_X2Y6_WW4BEG[4] ,
    \Tile_X2Y6_WW4BEG[3] ,
    \Tile_X2Y6_WW4BEG[2] ,
    \Tile_X2Y6_WW4BEG[1] ,
    \Tile_X2Y6_WW4BEG[0] }));
 LUT4AB Tile_X1Y7_LUT4AB (.Ci(Tile_X1Y8_Co),
    .Co(Tile_X1Y7_Co),
    .UserCLK(Tile_X1Y8_UserCLKo),
    .UserCLKo(Tile_X1Y7_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X1Y7_E1BEG[3] ,
    \Tile_X1Y7_E1BEG[2] ,
    \Tile_X1Y7_E1BEG[1] ,
    \Tile_X1Y7_E1BEG[0] }),
    .E1END({\Tile_X0Y7_E1BEG[3] ,
    \Tile_X0Y7_E1BEG[2] ,
    \Tile_X0Y7_E1BEG[1] ,
    \Tile_X0Y7_E1BEG[0] }),
    .E2BEG({\Tile_X1Y7_E2BEG[7] ,
    \Tile_X1Y7_E2BEG[6] ,
    \Tile_X1Y7_E2BEG[5] ,
    \Tile_X1Y7_E2BEG[4] ,
    \Tile_X1Y7_E2BEG[3] ,
    \Tile_X1Y7_E2BEG[2] ,
    \Tile_X1Y7_E2BEG[1] ,
    \Tile_X1Y7_E2BEG[0] }),
    .E2BEGb({\Tile_X1Y7_E2BEGb[7] ,
    \Tile_X1Y7_E2BEGb[6] ,
    \Tile_X1Y7_E2BEGb[5] ,
    \Tile_X1Y7_E2BEGb[4] ,
    \Tile_X1Y7_E2BEGb[3] ,
    \Tile_X1Y7_E2BEGb[2] ,
    \Tile_X1Y7_E2BEGb[1] ,
    \Tile_X1Y7_E2BEGb[0] }),
    .E2END({\Tile_X0Y7_E2BEGb[7] ,
    \Tile_X0Y7_E2BEGb[6] ,
    \Tile_X0Y7_E2BEGb[5] ,
    \Tile_X0Y7_E2BEGb[4] ,
    \Tile_X0Y7_E2BEGb[3] ,
    \Tile_X0Y7_E2BEGb[2] ,
    \Tile_X0Y7_E2BEGb[1] ,
    \Tile_X0Y7_E2BEGb[0] }),
    .E2MID({\Tile_X0Y7_E2BEG[7] ,
    \Tile_X0Y7_E2BEG[6] ,
    \Tile_X0Y7_E2BEG[5] ,
    \Tile_X0Y7_E2BEG[4] ,
    \Tile_X0Y7_E2BEG[3] ,
    \Tile_X0Y7_E2BEG[2] ,
    \Tile_X0Y7_E2BEG[1] ,
    \Tile_X0Y7_E2BEG[0] }),
    .E6BEG({\Tile_X1Y7_E6BEG[11] ,
    \Tile_X1Y7_E6BEG[10] ,
    \Tile_X1Y7_E6BEG[9] ,
    \Tile_X1Y7_E6BEG[8] ,
    \Tile_X1Y7_E6BEG[7] ,
    \Tile_X1Y7_E6BEG[6] ,
    \Tile_X1Y7_E6BEG[5] ,
    \Tile_X1Y7_E6BEG[4] ,
    \Tile_X1Y7_E6BEG[3] ,
    \Tile_X1Y7_E6BEG[2] ,
    \Tile_X1Y7_E6BEG[1] ,
    \Tile_X1Y7_E6BEG[0] }),
    .E6END({\Tile_X0Y7_E6BEG[11] ,
    \Tile_X0Y7_E6BEG[10] ,
    \Tile_X0Y7_E6BEG[9] ,
    \Tile_X0Y7_E6BEG[8] ,
    \Tile_X0Y7_E6BEG[7] ,
    \Tile_X0Y7_E6BEG[6] ,
    \Tile_X0Y7_E6BEG[5] ,
    \Tile_X0Y7_E6BEG[4] ,
    \Tile_X0Y7_E6BEG[3] ,
    \Tile_X0Y7_E6BEG[2] ,
    \Tile_X0Y7_E6BEG[1] ,
    \Tile_X0Y7_E6BEG[0] }),
    .EE4BEG({\Tile_X1Y7_EE4BEG[15] ,
    \Tile_X1Y7_EE4BEG[14] ,
    \Tile_X1Y7_EE4BEG[13] ,
    \Tile_X1Y7_EE4BEG[12] ,
    \Tile_X1Y7_EE4BEG[11] ,
    \Tile_X1Y7_EE4BEG[10] ,
    \Tile_X1Y7_EE4BEG[9] ,
    \Tile_X1Y7_EE4BEG[8] ,
    \Tile_X1Y7_EE4BEG[7] ,
    \Tile_X1Y7_EE4BEG[6] ,
    \Tile_X1Y7_EE4BEG[5] ,
    \Tile_X1Y7_EE4BEG[4] ,
    \Tile_X1Y7_EE4BEG[3] ,
    \Tile_X1Y7_EE4BEG[2] ,
    \Tile_X1Y7_EE4BEG[1] ,
    \Tile_X1Y7_EE4BEG[0] }),
    .EE4END({\Tile_X0Y7_EE4BEG[15] ,
    \Tile_X0Y7_EE4BEG[14] ,
    \Tile_X0Y7_EE4BEG[13] ,
    \Tile_X0Y7_EE4BEG[12] ,
    \Tile_X0Y7_EE4BEG[11] ,
    \Tile_X0Y7_EE4BEG[10] ,
    \Tile_X0Y7_EE4BEG[9] ,
    \Tile_X0Y7_EE4BEG[8] ,
    \Tile_X0Y7_EE4BEG[7] ,
    \Tile_X0Y7_EE4BEG[6] ,
    \Tile_X0Y7_EE4BEG[5] ,
    \Tile_X0Y7_EE4BEG[4] ,
    \Tile_X0Y7_EE4BEG[3] ,
    \Tile_X0Y7_EE4BEG[2] ,
    \Tile_X0Y7_EE4BEG[1] ,
    \Tile_X0Y7_EE4BEG[0] }),
    .FrameData({\Tile_X0Y7_FrameData_O[31] ,
    \Tile_X0Y7_FrameData_O[30] ,
    \Tile_X0Y7_FrameData_O[29] ,
    \Tile_X0Y7_FrameData_O[28] ,
    \Tile_X0Y7_FrameData_O[27] ,
    \Tile_X0Y7_FrameData_O[26] ,
    \Tile_X0Y7_FrameData_O[25] ,
    \Tile_X0Y7_FrameData_O[24] ,
    \Tile_X0Y7_FrameData_O[23] ,
    \Tile_X0Y7_FrameData_O[22] ,
    \Tile_X0Y7_FrameData_O[21] ,
    \Tile_X0Y7_FrameData_O[20] ,
    \Tile_X0Y7_FrameData_O[19] ,
    \Tile_X0Y7_FrameData_O[18] ,
    \Tile_X0Y7_FrameData_O[17] ,
    \Tile_X0Y7_FrameData_O[16] ,
    \Tile_X0Y7_FrameData_O[15] ,
    \Tile_X0Y7_FrameData_O[14] ,
    \Tile_X0Y7_FrameData_O[13] ,
    \Tile_X0Y7_FrameData_O[12] ,
    \Tile_X0Y7_FrameData_O[11] ,
    \Tile_X0Y7_FrameData_O[10] ,
    \Tile_X0Y7_FrameData_O[9] ,
    \Tile_X0Y7_FrameData_O[8] ,
    \Tile_X0Y7_FrameData_O[7] ,
    \Tile_X0Y7_FrameData_O[6] ,
    \Tile_X0Y7_FrameData_O[5] ,
    \Tile_X0Y7_FrameData_O[4] ,
    \Tile_X0Y7_FrameData_O[3] ,
    \Tile_X0Y7_FrameData_O[2] ,
    \Tile_X0Y7_FrameData_O[1] ,
    \Tile_X0Y7_FrameData_O[0] }),
    .FrameData_O({\Tile_X1Y7_FrameData_O[31] ,
    \Tile_X1Y7_FrameData_O[30] ,
    \Tile_X1Y7_FrameData_O[29] ,
    \Tile_X1Y7_FrameData_O[28] ,
    \Tile_X1Y7_FrameData_O[27] ,
    \Tile_X1Y7_FrameData_O[26] ,
    \Tile_X1Y7_FrameData_O[25] ,
    \Tile_X1Y7_FrameData_O[24] ,
    \Tile_X1Y7_FrameData_O[23] ,
    \Tile_X1Y7_FrameData_O[22] ,
    \Tile_X1Y7_FrameData_O[21] ,
    \Tile_X1Y7_FrameData_O[20] ,
    \Tile_X1Y7_FrameData_O[19] ,
    \Tile_X1Y7_FrameData_O[18] ,
    \Tile_X1Y7_FrameData_O[17] ,
    \Tile_X1Y7_FrameData_O[16] ,
    \Tile_X1Y7_FrameData_O[15] ,
    \Tile_X1Y7_FrameData_O[14] ,
    \Tile_X1Y7_FrameData_O[13] ,
    \Tile_X1Y7_FrameData_O[12] ,
    \Tile_X1Y7_FrameData_O[11] ,
    \Tile_X1Y7_FrameData_O[10] ,
    \Tile_X1Y7_FrameData_O[9] ,
    \Tile_X1Y7_FrameData_O[8] ,
    \Tile_X1Y7_FrameData_O[7] ,
    \Tile_X1Y7_FrameData_O[6] ,
    \Tile_X1Y7_FrameData_O[5] ,
    \Tile_X1Y7_FrameData_O[4] ,
    \Tile_X1Y7_FrameData_O[3] ,
    \Tile_X1Y7_FrameData_O[2] ,
    \Tile_X1Y7_FrameData_O[1] ,
    \Tile_X1Y7_FrameData_O[0] }),
    .FrameStrobe({\Tile_X1Y8_FrameStrobe_O[19] ,
    \Tile_X1Y8_FrameStrobe_O[18] ,
    \Tile_X1Y8_FrameStrobe_O[17] ,
    \Tile_X1Y8_FrameStrobe_O[16] ,
    \Tile_X1Y8_FrameStrobe_O[15] ,
    \Tile_X1Y8_FrameStrobe_O[14] ,
    \Tile_X1Y8_FrameStrobe_O[13] ,
    \Tile_X1Y8_FrameStrobe_O[12] ,
    \Tile_X1Y8_FrameStrobe_O[11] ,
    \Tile_X1Y8_FrameStrobe_O[10] ,
    \Tile_X1Y8_FrameStrobe_O[9] ,
    \Tile_X1Y8_FrameStrobe_O[8] ,
    \Tile_X1Y8_FrameStrobe_O[7] ,
    \Tile_X1Y8_FrameStrobe_O[6] ,
    \Tile_X1Y8_FrameStrobe_O[5] ,
    \Tile_X1Y8_FrameStrobe_O[4] ,
    \Tile_X1Y8_FrameStrobe_O[3] ,
    \Tile_X1Y8_FrameStrobe_O[2] ,
    \Tile_X1Y8_FrameStrobe_O[1] ,
    \Tile_X1Y8_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X1Y7_FrameStrobe_O[19] ,
    \Tile_X1Y7_FrameStrobe_O[18] ,
    \Tile_X1Y7_FrameStrobe_O[17] ,
    \Tile_X1Y7_FrameStrobe_O[16] ,
    \Tile_X1Y7_FrameStrobe_O[15] ,
    \Tile_X1Y7_FrameStrobe_O[14] ,
    \Tile_X1Y7_FrameStrobe_O[13] ,
    \Tile_X1Y7_FrameStrobe_O[12] ,
    \Tile_X1Y7_FrameStrobe_O[11] ,
    \Tile_X1Y7_FrameStrobe_O[10] ,
    \Tile_X1Y7_FrameStrobe_O[9] ,
    \Tile_X1Y7_FrameStrobe_O[8] ,
    \Tile_X1Y7_FrameStrobe_O[7] ,
    \Tile_X1Y7_FrameStrobe_O[6] ,
    \Tile_X1Y7_FrameStrobe_O[5] ,
    \Tile_X1Y7_FrameStrobe_O[4] ,
    \Tile_X1Y7_FrameStrobe_O[3] ,
    \Tile_X1Y7_FrameStrobe_O[2] ,
    \Tile_X1Y7_FrameStrobe_O[1] ,
    \Tile_X1Y7_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X1Y7_N1BEG[3] ,
    \Tile_X1Y7_N1BEG[2] ,
    \Tile_X1Y7_N1BEG[1] ,
    \Tile_X1Y7_N1BEG[0] }),
    .N1END({\Tile_X1Y8_N1BEG[3] ,
    \Tile_X1Y8_N1BEG[2] ,
    \Tile_X1Y8_N1BEG[1] ,
    \Tile_X1Y8_N1BEG[0] }),
    .N2BEG({\Tile_X1Y7_N2BEG[7] ,
    \Tile_X1Y7_N2BEG[6] ,
    \Tile_X1Y7_N2BEG[5] ,
    \Tile_X1Y7_N2BEG[4] ,
    \Tile_X1Y7_N2BEG[3] ,
    \Tile_X1Y7_N2BEG[2] ,
    \Tile_X1Y7_N2BEG[1] ,
    \Tile_X1Y7_N2BEG[0] }),
    .N2BEGb({\Tile_X1Y7_N2BEGb[7] ,
    \Tile_X1Y7_N2BEGb[6] ,
    \Tile_X1Y7_N2BEGb[5] ,
    \Tile_X1Y7_N2BEGb[4] ,
    \Tile_X1Y7_N2BEGb[3] ,
    \Tile_X1Y7_N2BEGb[2] ,
    \Tile_X1Y7_N2BEGb[1] ,
    \Tile_X1Y7_N2BEGb[0] }),
    .N2END({\Tile_X1Y8_N2BEGb[7] ,
    \Tile_X1Y8_N2BEGb[6] ,
    \Tile_X1Y8_N2BEGb[5] ,
    \Tile_X1Y8_N2BEGb[4] ,
    \Tile_X1Y8_N2BEGb[3] ,
    \Tile_X1Y8_N2BEGb[2] ,
    \Tile_X1Y8_N2BEGb[1] ,
    \Tile_X1Y8_N2BEGb[0] }),
    .N2MID({\Tile_X1Y8_N2BEG[7] ,
    \Tile_X1Y8_N2BEG[6] ,
    \Tile_X1Y8_N2BEG[5] ,
    \Tile_X1Y8_N2BEG[4] ,
    \Tile_X1Y8_N2BEG[3] ,
    \Tile_X1Y8_N2BEG[2] ,
    \Tile_X1Y8_N2BEG[1] ,
    \Tile_X1Y8_N2BEG[0] }),
    .N4BEG({\Tile_X1Y7_N4BEG[15] ,
    \Tile_X1Y7_N4BEG[14] ,
    \Tile_X1Y7_N4BEG[13] ,
    \Tile_X1Y7_N4BEG[12] ,
    \Tile_X1Y7_N4BEG[11] ,
    \Tile_X1Y7_N4BEG[10] ,
    \Tile_X1Y7_N4BEG[9] ,
    \Tile_X1Y7_N4BEG[8] ,
    \Tile_X1Y7_N4BEG[7] ,
    \Tile_X1Y7_N4BEG[6] ,
    \Tile_X1Y7_N4BEG[5] ,
    \Tile_X1Y7_N4BEG[4] ,
    \Tile_X1Y7_N4BEG[3] ,
    \Tile_X1Y7_N4BEG[2] ,
    \Tile_X1Y7_N4BEG[1] ,
    \Tile_X1Y7_N4BEG[0] }),
    .N4END({\Tile_X1Y8_N4BEG[15] ,
    \Tile_X1Y8_N4BEG[14] ,
    \Tile_X1Y8_N4BEG[13] ,
    \Tile_X1Y8_N4BEG[12] ,
    \Tile_X1Y8_N4BEG[11] ,
    \Tile_X1Y8_N4BEG[10] ,
    \Tile_X1Y8_N4BEG[9] ,
    \Tile_X1Y8_N4BEG[8] ,
    \Tile_X1Y8_N4BEG[7] ,
    \Tile_X1Y8_N4BEG[6] ,
    \Tile_X1Y8_N4BEG[5] ,
    \Tile_X1Y8_N4BEG[4] ,
    \Tile_X1Y8_N4BEG[3] ,
    \Tile_X1Y8_N4BEG[2] ,
    \Tile_X1Y8_N4BEG[1] ,
    \Tile_X1Y8_N4BEG[0] }),
    .NN4BEG({\Tile_X1Y7_NN4BEG[15] ,
    \Tile_X1Y7_NN4BEG[14] ,
    \Tile_X1Y7_NN4BEG[13] ,
    \Tile_X1Y7_NN4BEG[12] ,
    \Tile_X1Y7_NN4BEG[11] ,
    \Tile_X1Y7_NN4BEG[10] ,
    \Tile_X1Y7_NN4BEG[9] ,
    \Tile_X1Y7_NN4BEG[8] ,
    \Tile_X1Y7_NN4BEG[7] ,
    \Tile_X1Y7_NN4BEG[6] ,
    \Tile_X1Y7_NN4BEG[5] ,
    \Tile_X1Y7_NN4BEG[4] ,
    \Tile_X1Y7_NN4BEG[3] ,
    \Tile_X1Y7_NN4BEG[2] ,
    \Tile_X1Y7_NN4BEG[1] ,
    \Tile_X1Y7_NN4BEG[0] }),
    .NN4END({\Tile_X1Y8_NN4BEG[15] ,
    \Tile_X1Y8_NN4BEG[14] ,
    \Tile_X1Y8_NN4BEG[13] ,
    \Tile_X1Y8_NN4BEG[12] ,
    \Tile_X1Y8_NN4BEG[11] ,
    \Tile_X1Y8_NN4BEG[10] ,
    \Tile_X1Y8_NN4BEG[9] ,
    \Tile_X1Y8_NN4BEG[8] ,
    \Tile_X1Y8_NN4BEG[7] ,
    \Tile_X1Y8_NN4BEG[6] ,
    \Tile_X1Y8_NN4BEG[5] ,
    \Tile_X1Y8_NN4BEG[4] ,
    \Tile_X1Y8_NN4BEG[3] ,
    \Tile_X1Y8_NN4BEG[2] ,
    \Tile_X1Y8_NN4BEG[1] ,
    \Tile_X1Y8_NN4BEG[0] }),
    .S1BEG({\Tile_X1Y7_S1BEG[3] ,
    \Tile_X1Y7_S1BEG[2] ,
    \Tile_X1Y7_S1BEG[1] ,
    \Tile_X1Y7_S1BEG[0] }),
    .S1END({\Tile_X1Y6_S1BEG[3] ,
    \Tile_X1Y6_S1BEG[2] ,
    \Tile_X1Y6_S1BEG[1] ,
    \Tile_X1Y6_S1BEG[0] }),
    .S2BEG({\Tile_X1Y7_S2BEG[7] ,
    \Tile_X1Y7_S2BEG[6] ,
    \Tile_X1Y7_S2BEG[5] ,
    \Tile_X1Y7_S2BEG[4] ,
    \Tile_X1Y7_S2BEG[3] ,
    \Tile_X1Y7_S2BEG[2] ,
    \Tile_X1Y7_S2BEG[1] ,
    \Tile_X1Y7_S2BEG[0] }),
    .S2BEGb({\Tile_X1Y7_S2BEGb[7] ,
    \Tile_X1Y7_S2BEGb[6] ,
    \Tile_X1Y7_S2BEGb[5] ,
    \Tile_X1Y7_S2BEGb[4] ,
    \Tile_X1Y7_S2BEGb[3] ,
    \Tile_X1Y7_S2BEGb[2] ,
    \Tile_X1Y7_S2BEGb[1] ,
    \Tile_X1Y7_S2BEGb[0] }),
    .S2END({\Tile_X1Y6_S2BEGb[7] ,
    \Tile_X1Y6_S2BEGb[6] ,
    \Tile_X1Y6_S2BEGb[5] ,
    \Tile_X1Y6_S2BEGb[4] ,
    \Tile_X1Y6_S2BEGb[3] ,
    \Tile_X1Y6_S2BEGb[2] ,
    \Tile_X1Y6_S2BEGb[1] ,
    \Tile_X1Y6_S2BEGb[0] }),
    .S2MID({\Tile_X1Y6_S2BEG[7] ,
    \Tile_X1Y6_S2BEG[6] ,
    \Tile_X1Y6_S2BEG[5] ,
    \Tile_X1Y6_S2BEG[4] ,
    \Tile_X1Y6_S2BEG[3] ,
    \Tile_X1Y6_S2BEG[2] ,
    \Tile_X1Y6_S2BEG[1] ,
    \Tile_X1Y6_S2BEG[0] }),
    .S4BEG({\Tile_X1Y7_S4BEG[15] ,
    \Tile_X1Y7_S4BEG[14] ,
    \Tile_X1Y7_S4BEG[13] ,
    \Tile_X1Y7_S4BEG[12] ,
    \Tile_X1Y7_S4BEG[11] ,
    \Tile_X1Y7_S4BEG[10] ,
    \Tile_X1Y7_S4BEG[9] ,
    \Tile_X1Y7_S4BEG[8] ,
    \Tile_X1Y7_S4BEG[7] ,
    \Tile_X1Y7_S4BEG[6] ,
    \Tile_X1Y7_S4BEG[5] ,
    \Tile_X1Y7_S4BEG[4] ,
    \Tile_X1Y7_S4BEG[3] ,
    \Tile_X1Y7_S4BEG[2] ,
    \Tile_X1Y7_S4BEG[1] ,
    \Tile_X1Y7_S4BEG[0] }),
    .S4END({\Tile_X1Y6_S4BEG[15] ,
    \Tile_X1Y6_S4BEG[14] ,
    \Tile_X1Y6_S4BEG[13] ,
    \Tile_X1Y6_S4BEG[12] ,
    \Tile_X1Y6_S4BEG[11] ,
    \Tile_X1Y6_S4BEG[10] ,
    \Tile_X1Y6_S4BEG[9] ,
    \Tile_X1Y6_S4BEG[8] ,
    \Tile_X1Y6_S4BEG[7] ,
    \Tile_X1Y6_S4BEG[6] ,
    \Tile_X1Y6_S4BEG[5] ,
    \Tile_X1Y6_S4BEG[4] ,
    \Tile_X1Y6_S4BEG[3] ,
    \Tile_X1Y6_S4BEG[2] ,
    \Tile_X1Y6_S4BEG[1] ,
    \Tile_X1Y6_S4BEG[0] }),
    .SS4BEG({\Tile_X1Y7_SS4BEG[15] ,
    \Tile_X1Y7_SS4BEG[14] ,
    \Tile_X1Y7_SS4BEG[13] ,
    \Tile_X1Y7_SS4BEG[12] ,
    \Tile_X1Y7_SS4BEG[11] ,
    \Tile_X1Y7_SS4BEG[10] ,
    \Tile_X1Y7_SS4BEG[9] ,
    \Tile_X1Y7_SS4BEG[8] ,
    \Tile_X1Y7_SS4BEG[7] ,
    \Tile_X1Y7_SS4BEG[6] ,
    \Tile_X1Y7_SS4BEG[5] ,
    \Tile_X1Y7_SS4BEG[4] ,
    \Tile_X1Y7_SS4BEG[3] ,
    \Tile_X1Y7_SS4BEG[2] ,
    \Tile_X1Y7_SS4BEG[1] ,
    \Tile_X1Y7_SS4BEG[0] }),
    .SS4END({\Tile_X1Y6_SS4BEG[15] ,
    \Tile_X1Y6_SS4BEG[14] ,
    \Tile_X1Y6_SS4BEG[13] ,
    \Tile_X1Y6_SS4BEG[12] ,
    \Tile_X1Y6_SS4BEG[11] ,
    \Tile_X1Y6_SS4BEG[10] ,
    \Tile_X1Y6_SS4BEG[9] ,
    \Tile_X1Y6_SS4BEG[8] ,
    \Tile_X1Y6_SS4BEG[7] ,
    \Tile_X1Y6_SS4BEG[6] ,
    \Tile_X1Y6_SS4BEG[5] ,
    \Tile_X1Y6_SS4BEG[4] ,
    \Tile_X1Y6_SS4BEG[3] ,
    \Tile_X1Y6_SS4BEG[2] ,
    \Tile_X1Y6_SS4BEG[1] ,
    \Tile_X1Y6_SS4BEG[0] }),
    .W1BEG({\Tile_X1Y7_W1BEG[3] ,
    \Tile_X1Y7_W1BEG[2] ,
    \Tile_X1Y7_W1BEG[1] ,
    \Tile_X1Y7_W1BEG[0] }),
    .W1END({\Tile_X2Y7_W1BEG[3] ,
    \Tile_X2Y7_W1BEG[2] ,
    \Tile_X2Y7_W1BEG[1] ,
    \Tile_X2Y7_W1BEG[0] }),
    .W2BEG({\Tile_X1Y7_W2BEG[7] ,
    \Tile_X1Y7_W2BEG[6] ,
    \Tile_X1Y7_W2BEG[5] ,
    \Tile_X1Y7_W2BEG[4] ,
    \Tile_X1Y7_W2BEG[3] ,
    \Tile_X1Y7_W2BEG[2] ,
    \Tile_X1Y7_W2BEG[1] ,
    \Tile_X1Y7_W2BEG[0] }),
    .W2BEGb({\Tile_X1Y7_W2BEGb[7] ,
    \Tile_X1Y7_W2BEGb[6] ,
    \Tile_X1Y7_W2BEGb[5] ,
    \Tile_X1Y7_W2BEGb[4] ,
    \Tile_X1Y7_W2BEGb[3] ,
    \Tile_X1Y7_W2BEGb[2] ,
    \Tile_X1Y7_W2BEGb[1] ,
    \Tile_X1Y7_W2BEGb[0] }),
    .W2END({\Tile_X2Y7_W2BEGb[7] ,
    \Tile_X2Y7_W2BEGb[6] ,
    \Tile_X2Y7_W2BEGb[5] ,
    \Tile_X2Y7_W2BEGb[4] ,
    \Tile_X2Y7_W2BEGb[3] ,
    \Tile_X2Y7_W2BEGb[2] ,
    \Tile_X2Y7_W2BEGb[1] ,
    \Tile_X2Y7_W2BEGb[0] }),
    .W2MID({\Tile_X2Y7_W2BEG[7] ,
    \Tile_X2Y7_W2BEG[6] ,
    \Tile_X2Y7_W2BEG[5] ,
    \Tile_X2Y7_W2BEG[4] ,
    \Tile_X2Y7_W2BEG[3] ,
    \Tile_X2Y7_W2BEG[2] ,
    \Tile_X2Y7_W2BEG[1] ,
    \Tile_X2Y7_W2BEG[0] }),
    .W6BEG({\Tile_X1Y7_W6BEG[11] ,
    \Tile_X1Y7_W6BEG[10] ,
    \Tile_X1Y7_W6BEG[9] ,
    \Tile_X1Y7_W6BEG[8] ,
    \Tile_X1Y7_W6BEG[7] ,
    \Tile_X1Y7_W6BEG[6] ,
    \Tile_X1Y7_W6BEG[5] ,
    \Tile_X1Y7_W6BEG[4] ,
    \Tile_X1Y7_W6BEG[3] ,
    \Tile_X1Y7_W6BEG[2] ,
    \Tile_X1Y7_W6BEG[1] ,
    \Tile_X1Y7_W6BEG[0] }),
    .W6END({\Tile_X2Y7_W6BEG[11] ,
    \Tile_X2Y7_W6BEG[10] ,
    \Tile_X2Y7_W6BEG[9] ,
    \Tile_X2Y7_W6BEG[8] ,
    \Tile_X2Y7_W6BEG[7] ,
    \Tile_X2Y7_W6BEG[6] ,
    \Tile_X2Y7_W6BEG[5] ,
    \Tile_X2Y7_W6BEG[4] ,
    \Tile_X2Y7_W6BEG[3] ,
    \Tile_X2Y7_W6BEG[2] ,
    \Tile_X2Y7_W6BEG[1] ,
    \Tile_X2Y7_W6BEG[0] }),
    .WW4BEG({\Tile_X1Y7_WW4BEG[15] ,
    \Tile_X1Y7_WW4BEG[14] ,
    \Tile_X1Y7_WW4BEG[13] ,
    \Tile_X1Y7_WW4BEG[12] ,
    \Tile_X1Y7_WW4BEG[11] ,
    \Tile_X1Y7_WW4BEG[10] ,
    \Tile_X1Y7_WW4BEG[9] ,
    \Tile_X1Y7_WW4BEG[8] ,
    \Tile_X1Y7_WW4BEG[7] ,
    \Tile_X1Y7_WW4BEG[6] ,
    \Tile_X1Y7_WW4BEG[5] ,
    \Tile_X1Y7_WW4BEG[4] ,
    \Tile_X1Y7_WW4BEG[3] ,
    \Tile_X1Y7_WW4BEG[2] ,
    \Tile_X1Y7_WW4BEG[1] ,
    \Tile_X1Y7_WW4BEG[0] }),
    .WW4END({\Tile_X2Y7_WW4BEG[15] ,
    \Tile_X2Y7_WW4BEG[14] ,
    \Tile_X2Y7_WW4BEG[13] ,
    \Tile_X2Y7_WW4BEG[12] ,
    \Tile_X2Y7_WW4BEG[11] ,
    \Tile_X2Y7_WW4BEG[10] ,
    \Tile_X2Y7_WW4BEG[9] ,
    \Tile_X2Y7_WW4BEG[8] ,
    \Tile_X2Y7_WW4BEG[7] ,
    \Tile_X2Y7_WW4BEG[6] ,
    \Tile_X2Y7_WW4BEG[5] ,
    \Tile_X2Y7_WW4BEG[4] ,
    \Tile_X2Y7_WW4BEG[3] ,
    \Tile_X2Y7_WW4BEG[2] ,
    \Tile_X2Y7_WW4BEG[1] ,
    \Tile_X2Y7_WW4BEG[0] }));
 LUT4AB Tile_X1Y8_LUT4AB (.Ci(Tile_X1Y9_Co),
    .Co(Tile_X1Y8_Co),
    .UserCLK(Tile_X1Y9_UserCLKo),
    .UserCLKo(Tile_X1Y8_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X1Y8_E1BEG[3] ,
    \Tile_X1Y8_E1BEG[2] ,
    \Tile_X1Y8_E1BEG[1] ,
    \Tile_X1Y8_E1BEG[0] }),
    .E1END({\Tile_X0Y8_E1BEG[3] ,
    \Tile_X0Y8_E1BEG[2] ,
    \Tile_X0Y8_E1BEG[1] ,
    \Tile_X0Y8_E1BEG[0] }),
    .E2BEG({\Tile_X1Y8_E2BEG[7] ,
    \Tile_X1Y8_E2BEG[6] ,
    \Tile_X1Y8_E2BEG[5] ,
    \Tile_X1Y8_E2BEG[4] ,
    \Tile_X1Y8_E2BEG[3] ,
    \Tile_X1Y8_E2BEG[2] ,
    \Tile_X1Y8_E2BEG[1] ,
    \Tile_X1Y8_E2BEG[0] }),
    .E2BEGb({\Tile_X1Y8_E2BEGb[7] ,
    \Tile_X1Y8_E2BEGb[6] ,
    \Tile_X1Y8_E2BEGb[5] ,
    \Tile_X1Y8_E2BEGb[4] ,
    \Tile_X1Y8_E2BEGb[3] ,
    \Tile_X1Y8_E2BEGb[2] ,
    \Tile_X1Y8_E2BEGb[1] ,
    \Tile_X1Y8_E2BEGb[0] }),
    .E2END({\Tile_X0Y8_E2BEGb[7] ,
    \Tile_X0Y8_E2BEGb[6] ,
    \Tile_X0Y8_E2BEGb[5] ,
    \Tile_X0Y8_E2BEGb[4] ,
    \Tile_X0Y8_E2BEGb[3] ,
    \Tile_X0Y8_E2BEGb[2] ,
    \Tile_X0Y8_E2BEGb[1] ,
    \Tile_X0Y8_E2BEGb[0] }),
    .E2MID({\Tile_X0Y8_E2BEG[7] ,
    \Tile_X0Y8_E2BEG[6] ,
    \Tile_X0Y8_E2BEG[5] ,
    \Tile_X0Y8_E2BEG[4] ,
    \Tile_X0Y8_E2BEG[3] ,
    \Tile_X0Y8_E2BEG[2] ,
    \Tile_X0Y8_E2BEG[1] ,
    \Tile_X0Y8_E2BEG[0] }),
    .E6BEG({\Tile_X1Y8_E6BEG[11] ,
    \Tile_X1Y8_E6BEG[10] ,
    \Tile_X1Y8_E6BEG[9] ,
    \Tile_X1Y8_E6BEG[8] ,
    \Tile_X1Y8_E6BEG[7] ,
    \Tile_X1Y8_E6BEG[6] ,
    \Tile_X1Y8_E6BEG[5] ,
    \Tile_X1Y8_E6BEG[4] ,
    \Tile_X1Y8_E6BEG[3] ,
    \Tile_X1Y8_E6BEG[2] ,
    \Tile_X1Y8_E6BEG[1] ,
    \Tile_X1Y8_E6BEG[0] }),
    .E6END({\Tile_X0Y8_E6BEG[11] ,
    \Tile_X0Y8_E6BEG[10] ,
    \Tile_X0Y8_E6BEG[9] ,
    \Tile_X0Y8_E6BEG[8] ,
    \Tile_X0Y8_E6BEG[7] ,
    \Tile_X0Y8_E6BEG[6] ,
    \Tile_X0Y8_E6BEG[5] ,
    \Tile_X0Y8_E6BEG[4] ,
    \Tile_X0Y8_E6BEG[3] ,
    \Tile_X0Y8_E6BEG[2] ,
    \Tile_X0Y8_E6BEG[1] ,
    \Tile_X0Y8_E6BEG[0] }),
    .EE4BEG({\Tile_X1Y8_EE4BEG[15] ,
    \Tile_X1Y8_EE4BEG[14] ,
    \Tile_X1Y8_EE4BEG[13] ,
    \Tile_X1Y8_EE4BEG[12] ,
    \Tile_X1Y8_EE4BEG[11] ,
    \Tile_X1Y8_EE4BEG[10] ,
    \Tile_X1Y8_EE4BEG[9] ,
    \Tile_X1Y8_EE4BEG[8] ,
    \Tile_X1Y8_EE4BEG[7] ,
    \Tile_X1Y8_EE4BEG[6] ,
    \Tile_X1Y8_EE4BEG[5] ,
    \Tile_X1Y8_EE4BEG[4] ,
    \Tile_X1Y8_EE4BEG[3] ,
    \Tile_X1Y8_EE4BEG[2] ,
    \Tile_X1Y8_EE4BEG[1] ,
    \Tile_X1Y8_EE4BEG[0] }),
    .EE4END({\Tile_X0Y8_EE4BEG[15] ,
    \Tile_X0Y8_EE4BEG[14] ,
    \Tile_X0Y8_EE4BEG[13] ,
    \Tile_X0Y8_EE4BEG[12] ,
    \Tile_X0Y8_EE4BEG[11] ,
    \Tile_X0Y8_EE4BEG[10] ,
    \Tile_X0Y8_EE4BEG[9] ,
    \Tile_X0Y8_EE4BEG[8] ,
    \Tile_X0Y8_EE4BEG[7] ,
    \Tile_X0Y8_EE4BEG[6] ,
    \Tile_X0Y8_EE4BEG[5] ,
    \Tile_X0Y8_EE4BEG[4] ,
    \Tile_X0Y8_EE4BEG[3] ,
    \Tile_X0Y8_EE4BEG[2] ,
    \Tile_X0Y8_EE4BEG[1] ,
    \Tile_X0Y8_EE4BEG[0] }),
    .FrameData({\Tile_X0Y8_FrameData_O[31] ,
    \Tile_X0Y8_FrameData_O[30] ,
    \Tile_X0Y8_FrameData_O[29] ,
    \Tile_X0Y8_FrameData_O[28] ,
    \Tile_X0Y8_FrameData_O[27] ,
    \Tile_X0Y8_FrameData_O[26] ,
    \Tile_X0Y8_FrameData_O[25] ,
    \Tile_X0Y8_FrameData_O[24] ,
    \Tile_X0Y8_FrameData_O[23] ,
    \Tile_X0Y8_FrameData_O[22] ,
    \Tile_X0Y8_FrameData_O[21] ,
    \Tile_X0Y8_FrameData_O[20] ,
    \Tile_X0Y8_FrameData_O[19] ,
    \Tile_X0Y8_FrameData_O[18] ,
    \Tile_X0Y8_FrameData_O[17] ,
    \Tile_X0Y8_FrameData_O[16] ,
    \Tile_X0Y8_FrameData_O[15] ,
    \Tile_X0Y8_FrameData_O[14] ,
    \Tile_X0Y8_FrameData_O[13] ,
    \Tile_X0Y8_FrameData_O[12] ,
    \Tile_X0Y8_FrameData_O[11] ,
    \Tile_X0Y8_FrameData_O[10] ,
    \Tile_X0Y8_FrameData_O[9] ,
    \Tile_X0Y8_FrameData_O[8] ,
    \Tile_X0Y8_FrameData_O[7] ,
    \Tile_X0Y8_FrameData_O[6] ,
    \Tile_X0Y8_FrameData_O[5] ,
    \Tile_X0Y8_FrameData_O[4] ,
    \Tile_X0Y8_FrameData_O[3] ,
    \Tile_X0Y8_FrameData_O[2] ,
    \Tile_X0Y8_FrameData_O[1] ,
    \Tile_X0Y8_FrameData_O[0] }),
    .FrameData_O({\Tile_X1Y8_FrameData_O[31] ,
    \Tile_X1Y8_FrameData_O[30] ,
    \Tile_X1Y8_FrameData_O[29] ,
    \Tile_X1Y8_FrameData_O[28] ,
    \Tile_X1Y8_FrameData_O[27] ,
    \Tile_X1Y8_FrameData_O[26] ,
    \Tile_X1Y8_FrameData_O[25] ,
    \Tile_X1Y8_FrameData_O[24] ,
    \Tile_X1Y8_FrameData_O[23] ,
    \Tile_X1Y8_FrameData_O[22] ,
    \Tile_X1Y8_FrameData_O[21] ,
    \Tile_X1Y8_FrameData_O[20] ,
    \Tile_X1Y8_FrameData_O[19] ,
    \Tile_X1Y8_FrameData_O[18] ,
    \Tile_X1Y8_FrameData_O[17] ,
    \Tile_X1Y8_FrameData_O[16] ,
    \Tile_X1Y8_FrameData_O[15] ,
    \Tile_X1Y8_FrameData_O[14] ,
    \Tile_X1Y8_FrameData_O[13] ,
    \Tile_X1Y8_FrameData_O[12] ,
    \Tile_X1Y8_FrameData_O[11] ,
    \Tile_X1Y8_FrameData_O[10] ,
    \Tile_X1Y8_FrameData_O[9] ,
    \Tile_X1Y8_FrameData_O[8] ,
    \Tile_X1Y8_FrameData_O[7] ,
    \Tile_X1Y8_FrameData_O[6] ,
    \Tile_X1Y8_FrameData_O[5] ,
    \Tile_X1Y8_FrameData_O[4] ,
    \Tile_X1Y8_FrameData_O[3] ,
    \Tile_X1Y8_FrameData_O[2] ,
    \Tile_X1Y8_FrameData_O[1] ,
    \Tile_X1Y8_FrameData_O[0] }),
    .FrameStrobe({\Tile_X1Y9_FrameStrobe_O[19] ,
    \Tile_X1Y9_FrameStrobe_O[18] ,
    \Tile_X1Y9_FrameStrobe_O[17] ,
    \Tile_X1Y9_FrameStrobe_O[16] ,
    \Tile_X1Y9_FrameStrobe_O[15] ,
    \Tile_X1Y9_FrameStrobe_O[14] ,
    \Tile_X1Y9_FrameStrobe_O[13] ,
    \Tile_X1Y9_FrameStrobe_O[12] ,
    \Tile_X1Y9_FrameStrobe_O[11] ,
    \Tile_X1Y9_FrameStrobe_O[10] ,
    \Tile_X1Y9_FrameStrobe_O[9] ,
    \Tile_X1Y9_FrameStrobe_O[8] ,
    \Tile_X1Y9_FrameStrobe_O[7] ,
    \Tile_X1Y9_FrameStrobe_O[6] ,
    \Tile_X1Y9_FrameStrobe_O[5] ,
    \Tile_X1Y9_FrameStrobe_O[4] ,
    \Tile_X1Y9_FrameStrobe_O[3] ,
    \Tile_X1Y9_FrameStrobe_O[2] ,
    \Tile_X1Y9_FrameStrobe_O[1] ,
    \Tile_X1Y9_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X1Y8_FrameStrobe_O[19] ,
    \Tile_X1Y8_FrameStrobe_O[18] ,
    \Tile_X1Y8_FrameStrobe_O[17] ,
    \Tile_X1Y8_FrameStrobe_O[16] ,
    \Tile_X1Y8_FrameStrobe_O[15] ,
    \Tile_X1Y8_FrameStrobe_O[14] ,
    \Tile_X1Y8_FrameStrobe_O[13] ,
    \Tile_X1Y8_FrameStrobe_O[12] ,
    \Tile_X1Y8_FrameStrobe_O[11] ,
    \Tile_X1Y8_FrameStrobe_O[10] ,
    \Tile_X1Y8_FrameStrobe_O[9] ,
    \Tile_X1Y8_FrameStrobe_O[8] ,
    \Tile_X1Y8_FrameStrobe_O[7] ,
    \Tile_X1Y8_FrameStrobe_O[6] ,
    \Tile_X1Y8_FrameStrobe_O[5] ,
    \Tile_X1Y8_FrameStrobe_O[4] ,
    \Tile_X1Y8_FrameStrobe_O[3] ,
    \Tile_X1Y8_FrameStrobe_O[2] ,
    \Tile_X1Y8_FrameStrobe_O[1] ,
    \Tile_X1Y8_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X1Y8_N1BEG[3] ,
    \Tile_X1Y8_N1BEG[2] ,
    \Tile_X1Y8_N1BEG[1] ,
    \Tile_X1Y8_N1BEG[0] }),
    .N1END({\Tile_X1Y9_N1BEG[3] ,
    \Tile_X1Y9_N1BEG[2] ,
    \Tile_X1Y9_N1BEG[1] ,
    \Tile_X1Y9_N1BEG[0] }),
    .N2BEG({\Tile_X1Y8_N2BEG[7] ,
    \Tile_X1Y8_N2BEG[6] ,
    \Tile_X1Y8_N2BEG[5] ,
    \Tile_X1Y8_N2BEG[4] ,
    \Tile_X1Y8_N2BEG[3] ,
    \Tile_X1Y8_N2BEG[2] ,
    \Tile_X1Y8_N2BEG[1] ,
    \Tile_X1Y8_N2BEG[0] }),
    .N2BEGb({\Tile_X1Y8_N2BEGb[7] ,
    \Tile_X1Y8_N2BEGb[6] ,
    \Tile_X1Y8_N2BEGb[5] ,
    \Tile_X1Y8_N2BEGb[4] ,
    \Tile_X1Y8_N2BEGb[3] ,
    \Tile_X1Y8_N2BEGb[2] ,
    \Tile_X1Y8_N2BEGb[1] ,
    \Tile_X1Y8_N2BEGb[0] }),
    .N2END({\Tile_X1Y9_N2BEGb[7] ,
    \Tile_X1Y9_N2BEGb[6] ,
    \Tile_X1Y9_N2BEGb[5] ,
    \Tile_X1Y9_N2BEGb[4] ,
    \Tile_X1Y9_N2BEGb[3] ,
    \Tile_X1Y9_N2BEGb[2] ,
    \Tile_X1Y9_N2BEGb[1] ,
    \Tile_X1Y9_N2BEGb[0] }),
    .N2MID({\Tile_X1Y9_N2BEG[7] ,
    \Tile_X1Y9_N2BEG[6] ,
    \Tile_X1Y9_N2BEG[5] ,
    \Tile_X1Y9_N2BEG[4] ,
    \Tile_X1Y9_N2BEG[3] ,
    \Tile_X1Y9_N2BEG[2] ,
    \Tile_X1Y9_N2BEG[1] ,
    \Tile_X1Y9_N2BEG[0] }),
    .N4BEG({\Tile_X1Y8_N4BEG[15] ,
    \Tile_X1Y8_N4BEG[14] ,
    \Tile_X1Y8_N4BEG[13] ,
    \Tile_X1Y8_N4BEG[12] ,
    \Tile_X1Y8_N4BEG[11] ,
    \Tile_X1Y8_N4BEG[10] ,
    \Tile_X1Y8_N4BEG[9] ,
    \Tile_X1Y8_N4BEG[8] ,
    \Tile_X1Y8_N4BEG[7] ,
    \Tile_X1Y8_N4BEG[6] ,
    \Tile_X1Y8_N4BEG[5] ,
    \Tile_X1Y8_N4BEG[4] ,
    \Tile_X1Y8_N4BEG[3] ,
    \Tile_X1Y8_N4BEG[2] ,
    \Tile_X1Y8_N4BEG[1] ,
    \Tile_X1Y8_N4BEG[0] }),
    .N4END({\Tile_X1Y9_N4BEG[15] ,
    \Tile_X1Y9_N4BEG[14] ,
    \Tile_X1Y9_N4BEG[13] ,
    \Tile_X1Y9_N4BEG[12] ,
    \Tile_X1Y9_N4BEG[11] ,
    \Tile_X1Y9_N4BEG[10] ,
    \Tile_X1Y9_N4BEG[9] ,
    \Tile_X1Y9_N4BEG[8] ,
    \Tile_X1Y9_N4BEG[7] ,
    \Tile_X1Y9_N4BEG[6] ,
    \Tile_X1Y9_N4BEG[5] ,
    \Tile_X1Y9_N4BEG[4] ,
    \Tile_X1Y9_N4BEG[3] ,
    \Tile_X1Y9_N4BEG[2] ,
    \Tile_X1Y9_N4BEG[1] ,
    \Tile_X1Y9_N4BEG[0] }),
    .NN4BEG({\Tile_X1Y8_NN4BEG[15] ,
    \Tile_X1Y8_NN4BEG[14] ,
    \Tile_X1Y8_NN4BEG[13] ,
    \Tile_X1Y8_NN4BEG[12] ,
    \Tile_X1Y8_NN4BEG[11] ,
    \Tile_X1Y8_NN4BEG[10] ,
    \Tile_X1Y8_NN4BEG[9] ,
    \Tile_X1Y8_NN4BEG[8] ,
    \Tile_X1Y8_NN4BEG[7] ,
    \Tile_X1Y8_NN4BEG[6] ,
    \Tile_X1Y8_NN4BEG[5] ,
    \Tile_X1Y8_NN4BEG[4] ,
    \Tile_X1Y8_NN4BEG[3] ,
    \Tile_X1Y8_NN4BEG[2] ,
    \Tile_X1Y8_NN4BEG[1] ,
    \Tile_X1Y8_NN4BEG[0] }),
    .NN4END({\Tile_X1Y9_NN4BEG[15] ,
    \Tile_X1Y9_NN4BEG[14] ,
    \Tile_X1Y9_NN4BEG[13] ,
    \Tile_X1Y9_NN4BEG[12] ,
    \Tile_X1Y9_NN4BEG[11] ,
    \Tile_X1Y9_NN4BEG[10] ,
    \Tile_X1Y9_NN4BEG[9] ,
    \Tile_X1Y9_NN4BEG[8] ,
    \Tile_X1Y9_NN4BEG[7] ,
    \Tile_X1Y9_NN4BEG[6] ,
    \Tile_X1Y9_NN4BEG[5] ,
    \Tile_X1Y9_NN4BEG[4] ,
    \Tile_X1Y9_NN4BEG[3] ,
    \Tile_X1Y9_NN4BEG[2] ,
    \Tile_X1Y9_NN4BEG[1] ,
    \Tile_X1Y9_NN4BEG[0] }),
    .S1BEG({\Tile_X1Y8_S1BEG[3] ,
    \Tile_X1Y8_S1BEG[2] ,
    \Tile_X1Y8_S1BEG[1] ,
    \Tile_X1Y8_S1BEG[0] }),
    .S1END({\Tile_X1Y7_S1BEG[3] ,
    \Tile_X1Y7_S1BEG[2] ,
    \Tile_X1Y7_S1BEG[1] ,
    \Tile_X1Y7_S1BEG[0] }),
    .S2BEG({\Tile_X1Y8_S2BEG[7] ,
    \Tile_X1Y8_S2BEG[6] ,
    \Tile_X1Y8_S2BEG[5] ,
    \Tile_X1Y8_S2BEG[4] ,
    \Tile_X1Y8_S2BEG[3] ,
    \Tile_X1Y8_S2BEG[2] ,
    \Tile_X1Y8_S2BEG[1] ,
    \Tile_X1Y8_S2BEG[0] }),
    .S2BEGb({\Tile_X1Y8_S2BEGb[7] ,
    \Tile_X1Y8_S2BEGb[6] ,
    \Tile_X1Y8_S2BEGb[5] ,
    \Tile_X1Y8_S2BEGb[4] ,
    \Tile_X1Y8_S2BEGb[3] ,
    \Tile_X1Y8_S2BEGb[2] ,
    \Tile_X1Y8_S2BEGb[1] ,
    \Tile_X1Y8_S2BEGb[0] }),
    .S2END({\Tile_X1Y7_S2BEGb[7] ,
    \Tile_X1Y7_S2BEGb[6] ,
    \Tile_X1Y7_S2BEGb[5] ,
    \Tile_X1Y7_S2BEGb[4] ,
    \Tile_X1Y7_S2BEGb[3] ,
    \Tile_X1Y7_S2BEGb[2] ,
    \Tile_X1Y7_S2BEGb[1] ,
    \Tile_X1Y7_S2BEGb[0] }),
    .S2MID({\Tile_X1Y7_S2BEG[7] ,
    \Tile_X1Y7_S2BEG[6] ,
    \Tile_X1Y7_S2BEG[5] ,
    \Tile_X1Y7_S2BEG[4] ,
    \Tile_X1Y7_S2BEG[3] ,
    \Tile_X1Y7_S2BEG[2] ,
    \Tile_X1Y7_S2BEG[1] ,
    \Tile_X1Y7_S2BEG[0] }),
    .S4BEG({\Tile_X1Y8_S4BEG[15] ,
    \Tile_X1Y8_S4BEG[14] ,
    \Tile_X1Y8_S4BEG[13] ,
    \Tile_X1Y8_S4BEG[12] ,
    \Tile_X1Y8_S4BEG[11] ,
    \Tile_X1Y8_S4BEG[10] ,
    \Tile_X1Y8_S4BEG[9] ,
    \Tile_X1Y8_S4BEG[8] ,
    \Tile_X1Y8_S4BEG[7] ,
    \Tile_X1Y8_S4BEG[6] ,
    \Tile_X1Y8_S4BEG[5] ,
    \Tile_X1Y8_S4BEG[4] ,
    \Tile_X1Y8_S4BEG[3] ,
    \Tile_X1Y8_S4BEG[2] ,
    \Tile_X1Y8_S4BEG[1] ,
    \Tile_X1Y8_S4BEG[0] }),
    .S4END({\Tile_X1Y7_S4BEG[15] ,
    \Tile_X1Y7_S4BEG[14] ,
    \Tile_X1Y7_S4BEG[13] ,
    \Tile_X1Y7_S4BEG[12] ,
    \Tile_X1Y7_S4BEG[11] ,
    \Tile_X1Y7_S4BEG[10] ,
    \Tile_X1Y7_S4BEG[9] ,
    \Tile_X1Y7_S4BEG[8] ,
    \Tile_X1Y7_S4BEG[7] ,
    \Tile_X1Y7_S4BEG[6] ,
    \Tile_X1Y7_S4BEG[5] ,
    \Tile_X1Y7_S4BEG[4] ,
    \Tile_X1Y7_S4BEG[3] ,
    \Tile_X1Y7_S4BEG[2] ,
    \Tile_X1Y7_S4BEG[1] ,
    \Tile_X1Y7_S4BEG[0] }),
    .SS4BEG({\Tile_X1Y8_SS4BEG[15] ,
    \Tile_X1Y8_SS4BEG[14] ,
    \Tile_X1Y8_SS4BEG[13] ,
    \Tile_X1Y8_SS4BEG[12] ,
    \Tile_X1Y8_SS4BEG[11] ,
    \Tile_X1Y8_SS4BEG[10] ,
    \Tile_X1Y8_SS4BEG[9] ,
    \Tile_X1Y8_SS4BEG[8] ,
    \Tile_X1Y8_SS4BEG[7] ,
    \Tile_X1Y8_SS4BEG[6] ,
    \Tile_X1Y8_SS4BEG[5] ,
    \Tile_X1Y8_SS4BEG[4] ,
    \Tile_X1Y8_SS4BEG[3] ,
    \Tile_X1Y8_SS4BEG[2] ,
    \Tile_X1Y8_SS4BEG[1] ,
    \Tile_X1Y8_SS4BEG[0] }),
    .SS4END({\Tile_X1Y7_SS4BEG[15] ,
    \Tile_X1Y7_SS4BEG[14] ,
    \Tile_X1Y7_SS4BEG[13] ,
    \Tile_X1Y7_SS4BEG[12] ,
    \Tile_X1Y7_SS4BEG[11] ,
    \Tile_X1Y7_SS4BEG[10] ,
    \Tile_X1Y7_SS4BEG[9] ,
    \Tile_X1Y7_SS4BEG[8] ,
    \Tile_X1Y7_SS4BEG[7] ,
    \Tile_X1Y7_SS4BEG[6] ,
    \Tile_X1Y7_SS4BEG[5] ,
    \Tile_X1Y7_SS4BEG[4] ,
    \Tile_X1Y7_SS4BEG[3] ,
    \Tile_X1Y7_SS4BEG[2] ,
    \Tile_X1Y7_SS4BEG[1] ,
    \Tile_X1Y7_SS4BEG[0] }),
    .W1BEG({\Tile_X1Y8_W1BEG[3] ,
    \Tile_X1Y8_W1BEG[2] ,
    \Tile_X1Y8_W1BEG[1] ,
    \Tile_X1Y8_W1BEG[0] }),
    .W1END({\Tile_X2Y8_W1BEG[3] ,
    \Tile_X2Y8_W1BEG[2] ,
    \Tile_X2Y8_W1BEG[1] ,
    \Tile_X2Y8_W1BEG[0] }),
    .W2BEG({\Tile_X1Y8_W2BEG[7] ,
    \Tile_X1Y8_W2BEG[6] ,
    \Tile_X1Y8_W2BEG[5] ,
    \Tile_X1Y8_W2BEG[4] ,
    \Tile_X1Y8_W2BEG[3] ,
    \Tile_X1Y8_W2BEG[2] ,
    \Tile_X1Y8_W2BEG[1] ,
    \Tile_X1Y8_W2BEG[0] }),
    .W2BEGb({\Tile_X1Y8_W2BEGb[7] ,
    \Tile_X1Y8_W2BEGb[6] ,
    \Tile_X1Y8_W2BEGb[5] ,
    \Tile_X1Y8_W2BEGb[4] ,
    \Tile_X1Y8_W2BEGb[3] ,
    \Tile_X1Y8_W2BEGb[2] ,
    \Tile_X1Y8_W2BEGb[1] ,
    \Tile_X1Y8_W2BEGb[0] }),
    .W2END({\Tile_X2Y8_W2BEGb[7] ,
    \Tile_X2Y8_W2BEGb[6] ,
    \Tile_X2Y8_W2BEGb[5] ,
    \Tile_X2Y8_W2BEGb[4] ,
    \Tile_X2Y8_W2BEGb[3] ,
    \Tile_X2Y8_W2BEGb[2] ,
    \Tile_X2Y8_W2BEGb[1] ,
    \Tile_X2Y8_W2BEGb[0] }),
    .W2MID({\Tile_X2Y8_W2BEG[7] ,
    \Tile_X2Y8_W2BEG[6] ,
    \Tile_X2Y8_W2BEG[5] ,
    \Tile_X2Y8_W2BEG[4] ,
    \Tile_X2Y8_W2BEG[3] ,
    \Tile_X2Y8_W2BEG[2] ,
    \Tile_X2Y8_W2BEG[1] ,
    \Tile_X2Y8_W2BEG[0] }),
    .W6BEG({\Tile_X1Y8_W6BEG[11] ,
    \Tile_X1Y8_W6BEG[10] ,
    \Tile_X1Y8_W6BEG[9] ,
    \Tile_X1Y8_W6BEG[8] ,
    \Tile_X1Y8_W6BEG[7] ,
    \Tile_X1Y8_W6BEG[6] ,
    \Tile_X1Y8_W6BEG[5] ,
    \Tile_X1Y8_W6BEG[4] ,
    \Tile_X1Y8_W6BEG[3] ,
    \Tile_X1Y8_W6BEG[2] ,
    \Tile_X1Y8_W6BEG[1] ,
    \Tile_X1Y8_W6BEG[0] }),
    .W6END({\Tile_X2Y8_W6BEG[11] ,
    \Tile_X2Y8_W6BEG[10] ,
    \Tile_X2Y8_W6BEG[9] ,
    \Tile_X2Y8_W6BEG[8] ,
    \Tile_X2Y8_W6BEG[7] ,
    \Tile_X2Y8_W6BEG[6] ,
    \Tile_X2Y8_W6BEG[5] ,
    \Tile_X2Y8_W6BEG[4] ,
    \Tile_X2Y8_W6BEG[3] ,
    \Tile_X2Y8_W6BEG[2] ,
    \Tile_X2Y8_W6BEG[1] ,
    \Tile_X2Y8_W6BEG[0] }),
    .WW4BEG({\Tile_X1Y8_WW4BEG[15] ,
    \Tile_X1Y8_WW4BEG[14] ,
    \Tile_X1Y8_WW4BEG[13] ,
    \Tile_X1Y8_WW4BEG[12] ,
    \Tile_X1Y8_WW4BEG[11] ,
    \Tile_X1Y8_WW4BEG[10] ,
    \Tile_X1Y8_WW4BEG[9] ,
    \Tile_X1Y8_WW4BEG[8] ,
    \Tile_X1Y8_WW4BEG[7] ,
    \Tile_X1Y8_WW4BEG[6] ,
    \Tile_X1Y8_WW4BEG[5] ,
    \Tile_X1Y8_WW4BEG[4] ,
    \Tile_X1Y8_WW4BEG[3] ,
    \Tile_X1Y8_WW4BEG[2] ,
    \Tile_X1Y8_WW4BEG[1] ,
    \Tile_X1Y8_WW4BEG[0] }),
    .WW4END({\Tile_X2Y8_WW4BEG[15] ,
    \Tile_X2Y8_WW4BEG[14] ,
    \Tile_X2Y8_WW4BEG[13] ,
    \Tile_X2Y8_WW4BEG[12] ,
    \Tile_X2Y8_WW4BEG[11] ,
    \Tile_X2Y8_WW4BEG[10] ,
    \Tile_X2Y8_WW4BEG[9] ,
    \Tile_X2Y8_WW4BEG[8] ,
    \Tile_X2Y8_WW4BEG[7] ,
    \Tile_X2Y8_WW4BEG[6] ,
    \Tile_X2Y8_WW4BEG[5] ,
    \Tile_X2Y8_WW4BEG[4] ,
    \Tile_X2Y8_WW4BEG[3] ,
    \Tile_X2Y8_WW4BEG[2] ,
    \Tile_X2Y8_WW4BEG[1] ,
    \Tile_X2Y8_WW4BEG[0] }));
 LUT4AB Tile_X1Y9_LUT4AB (.Ci(Tile_X1Y10_Co),
    .Co(Tile_X1Y9_Co),
    .UserCLK(Tile_X1Y10_UserCLKo),
    .UserCLKo(Tile_X1Y9_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X1Y9_E1BEG[3] ,
    \Tile_X1Y9_E1BEG[2] ,
    \Tile_X1Y9_E1BEG[1] ,
    \Tile_X1Y9_E1BEG[0] }),
    .E1END({\Tile_X0Y9_E1BEG[3] ,
    \Tile_X0Y9_E1BEG[2] ,
    \Tile_X0Y9_E1BEG[1] ,
    \Tile_X0Y9_E1BEG[0] }),
    .E2BEG({\Tile_X1Y9_E2BEG[7] ,
    \Tile_X1Y9_E2BEG[6] ,
    \Tile_X1Y9_E2BEG[5] ,
    \Tile_X1Y9_E2BEG[4] ,
    \Tile_X1Y9_E2BEG[3] ,
    \Tile_X1Y9_E2BEG[2] ,
    \Tile_X1Y9_E2BEG[1] ,
    \Tile_X1Y9_E2BEG[0] }),
    .E2BEGb({\Tile_X1Y9_E2BEGb[7] ,
    \Tile_X1Y9_E2BEGb[6] ,
    \Tile_X1Y9_E2BEGb[5] ,
    \Tile_X1Y9_E2BEGb[4] ,
    \Tile_X1Y9_E2BEGb[3] ,
    \Tile_X1Y9_E2BEGb[2] ,
    \Tile_X1Y9_E2BEGb[1] ,
    \Tile_X1Y9_E2BEGb[0] }),
    .E2END({\Tile_X0Y9_E2BEGb[7] ,
    \Tile_X0Y9_E2BEGb[6] ,
    \Tile_X0Y9_E2BEGb[5] ,
    \Tile_X0Y9_E2BEGb[4] ,
    \Tile_X0Y9_E2BEGb[3] ,
    \Tile_X0Y9_E2BEGb[2] ,
    \Tile_X0Y9_E2BEGb[1] ,
    \Tile_X0Y9_E2BEGb[0] }),
    .E2MID({\Tile_X0Y9_E2BEG[7] ,
    \Tile_X0Y9_E2BEG[6] ,
    \Tile_X0Y9_E2BEG[5] ,
    \Tile_X0Y9_E2BEG[4] ,
    \Tile_X0Y9_E2BEG[3] ,
    \Tile_X0Y9_E2BEG[2] ,
    \Tile_X0Y9_E2BEG[1] ,
    \Tile_X0Y9_E2BEG[0] }),
    .E6BEG({\Tile_X1Y9_E6BEG[11] ,
    \Tile_X1Y9_E6BEG[10] ,
    \Tile_X1Y9_E6BEG[9] ,
    \Tile_X1Y9_E6BEG[8] ,
    \Tile_X1Y9_E6BEG[7] ,
    \Tile_X1Y9_E6BEG[6] ,
    \Tile_X1Y9_E6BEG[5] ,
    \Tile_X1Y9_E6BEG[4] ,
    \Tile_X1Y9_E6BEG[3] ,
    \Tile_X1Y9_E6BEG[2] ,
    \Tile_X1Y9_E6BEG[1] ,
    \Tile_X1Y9_E6BEG[0] }),
    .E6END({\Tile_X0Y9_E6BEG[11] ,
    \Tile_X0Y9_E6BEG[10] ,
    \Tile_X0Y9_E6BEG[9] ,
    \Tile_X0Y9_E6BEG[8] ,
    \Tile_X0Y9_E6BEG[7] ,
    \Tile_X0Y9_E6BEG[6] ,
    \Tile_X0Y9_E6BEG[5] ,
    \Tile_X0Y9_E6BEG[4] ,
    \Tile_X0Y9_E6BEG[3] ,
    \Tile_X0Y9_E6BEG[2] ,
    \Tile_X0Y9_E6BEG[1] ,
    \Tile_X0Y9_E6BEG[0] }),
    .EE4BEG({\Tile_X1Y9_EE4BEG[15] ,
    \Tile_X1Y9_EE4BEG[14] ,
    \Tile_X1Y9_EE4BEG[13] ,
    \Tile_X1Y9_EE4BEG[12] ,
    \Tile_X1Y9_EE4BEG[11] ,
    \Tile_X1Y9_EE4BEG[10] ,
    \Tile_X1Y9_EE4BEG[9] ,
    \Tile_X1Y9_EE4BEG[8] ,
    \Tile_X1Y9_EE4BEG[7] ,
    \Tile_X1Y9_EE4BEG[6] ,
    \Tile_X1Y9_EE4BEG[5] ,
    \Tile_X1Y9_EE4BEG[4] ,
    \Tile_X1Y9_EE4BEG[3] ,
    \Tile_X1Y9_EE4BEG[2] ,
    \Tile_X1Y9_EE4BEG[1] ,
    \Tile_X1Y9_EE4BEG[0] }),
    .EE4END({\Tile_X0Y9_EE4BEG[15] ,
    \Tile_X0Y9_EE4BEG[14] ,
    \Tile_X0Y9_EE4BEG[13] ,
    \Tile_X0Y9_EE4BEG[12] ,
    \Tile_X0Y9_EE4BEG[11] ,
    \Tile_X0Y9_EE4BEG[10] ,
    \Tile_X0Y9_EE4BEG[9] ,
    \Tile_X0Y9_EE4BEG[8] ,
    \Tile_X0Y9_EE4BEG[7] ,
    \Tile_X0Y9_EE4BEG[6] ,
    \Tile_X0Y9_EE4BEG[5] ,
    \Tile_X0Y9_EE4BEG[4] ,
    \Tile_X0Y9_EE4BEG[3] ,
    \Tile_X0Y9_EE4BEG[2] ,
    \Tile_X0Y9_EE4BEG[1] ,
    \Tile_X0Y9_EE4BEG[0] }),
    .FrameData({\Tile_X0Y9_FrameData_O[31] ,
    \Tile_X0Y9_FrameData_O[30] ,
    \Tile_X0Y9_FrameData_O[29] ,
    \Tile_X0Y9_FrameData_O[28] ,
    \Tile_X0Y9_FrameData_O[27] ,
    \Tile_X0Y9_FrameData_O[26] ,
    \Tile_X0Y9_FrameData_O[25] ,
    \Tile_X0Y9_FrameData_O[24] ,
    \Tile_X0Y9_FrameData_O[23] ,
    \Tile_X0Y9_FrameData_O[22] ,
    \Tile_X0Y9_FrameData_O[21] ,
    \Tile_X0Y9_FrameData_O[20] ,
    \Tile_X0Y9_FrameData_O[19] ,
    \Tile_X0Y9_FrameData_O[18] ,
    \Tile_X0Y9_FrameData_O[17] ,
    \Tile_X0Y9_FrameData_O[16] ,
    \Tile_X0Y9_FrameData_O[15] ,
    \Tile_X0Y9_FrameData_O[14] ,
    \Tile_X0Y9_FrameData_O[13] ,
    \Tile_X0Y9_FrameData_O[12] ,
    \Tile_X0Y9_FrameData_O[11] ,
    \Tile_X0Y9_FrameData_O[10] ,
    \Tile_X0Y9_FrameData_O[9] ,
    \Tile_X0Y9_FrameData_O[8] ,
    \Tile_X0Y9_FrameData_O[7] ,
    \Tile_X0Y9_FrameData_O[6] ,
    \Tile_X0Y9_FrameData_O[5] ,
    \Tile_X0Y9_FrameData_O[4] ,
    \Tile_X0Y9_FrameData_O[3] ,
    \Tile_X0Y9_FrameData_O[2] ,
    \Tile_X0Y9_FrameData_O[1] ,
    \Tile_X0Y9_FrameData_O[0] }),
    .FrameData_O({\Tile_X1Y9_FrameData_O[31] ,
    \Tile_X1Y9_FrameData_O[30] ,
    \Tile_X1Y9_FrameData_O[29] ,
    \Tile_X1Y9_FrameData_O[28] ,
    \Tile_X1Y9_FrameData_O[27] ,
    \Tile_X1Y9_FrameData_O[26] ,
    \Tile_X1Y9_FrameData_O[25] ,
    \Tile_X1Y9_FrameData_O[24] ,
    \Tile_X1Y9_FrameData_O[23] ,
    \Tile_X1Y9_FrameData_O[22] ,
    \Tile_X1Y9_FrameData_O[21] ,
    \Tile_X1Y9_FrameData_O[20] ,
    \Tile_X1Y9_FrameData_O[19] ,
    \Tile_X1Y9_FrameData_O[18] ,
    \Tile_X1Y9_FrameData_O[17] ,
    \Tile_X1Y9_FrameData_O[16] ,
    \Tile_X1Y9_FrameData_O[15] ,
    \Tile_X1Y9_FrameData_O[14] ,
    \Tile_X1Y9_FrameData_O[13] ,
    \Tile_X1Y9_FrameData_O[12] ,
    \Tile_X1Y9_FrameData_O[11] ,
    \Tile_X1Y9_FrameData_O[10] ,
    \Tile_X1Y9_FrameData_O[9] ,
    \Tile_X1Y9_FrameData_O[8] ,
    \Tile_X1Y9_FrameData_O[7] ,
    \Tile_X1Y9_FrameData_O[6] ,
    \Tile_X1Y9_FrameData_O[5] ,
    \Tile_X1Y9_FrameData_O[4] ,
    \Tile_X1Y9_FrameData_O[3] ,
    \Tile_X1Y9_FrameData_O[2] ,
    \Tile_X1Y9_FrameData_O[1] ,
    \Tile_X1Y9_FrameData_O[0] }),
    .FrameStrobe({\Tile_X1Y10_FrameStrobe_O[19] ,
    \Tile_X1Y10_FrameStrobe_O[18] ,
    \Tile_X1Y10_FrameStrobe_O[17] ,
    \Tile_X1Y10_FrameStrobe_O[16] ,
    \Tile_X1Y10_FrameStrobe_O[15] ,
    \Tile_X1Y10_FrameStrobe_O[14] ,
    \Tile_X1Y10_FrameStrobe_O[13] ,
    \Tile_X1Y10_FrameStrobe_O[12] ,
    \Tile_X1Y10_FrameStrobe_O[11] ,
    \Tile_X1Y10_FrameStrobe_O[10] ,
    \Tile_X1Y10_FrameStrobe_O[9] ,
    \Tile_X1Y10_FrameStrobe_O[8] ,
    \Tile_X1Y10_FrameStrobe_O[7] ,
    \Tile_X1Y10_FrameStrobe_O[6] ,
    \Tile_X1Y10_FrameStrobe_O[5] ,
    \Tile_X1Y10_FrameStrobe_O[4] ,
    \Tile_X1Y10_FrameStrobe_O[3] ,
    \Tile_X1Y10_FrameStrobe_O[2] ,
    \Tile_X1Y10_FrameStrobe_O[1] ,
    \Tile_X1Y10_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X1Y9_FrameStrobe_O[19] ,
    \Tile_X1Y9_FrameStrobe_O[18] ,
    \Tile_X1Y9_FrameStrobe_O[17] ,
    \Tile_X1Y9_FrameStrobe_O[16] ,
    \Tile_X1Y9_FrameStrobe_O[15] ,
    \Tile_X1Y9_FrameStrobe_O[14] ,
    \Tile_X1Y9_FrameStrobe_O[13] ,
    \Tile_X1Y9_FrameStrobe_O[12] ,
    \Tile_X1Y9_FrameStrobe_O[11] ,
    \Tile_X1Y9_FrameStrobe_O[10] ,
    \Tile_X1Y9_FrameStrobe_O[9] ,
    \Tile_X1Y9_FrameStrobe_O[8] ,
    \Tile_X1Y9_FrameStrobe_O[7] ,
    \Tile_X1Y9_FrameStrobe_O[6] ,
    \Tile_X1Y9_FrameStrobe_O[5] ,
    \Tile_X1Y9_FrameStrobe_O[4] ,
    \Tile_X1Y9_FrameStrobe_O[3] ,
    \Tile_X1Y9_FrameStrobe_O[2] ,
    \Tile_X1Y9_FrameStrobe_O[1] ,
    \Tile_X1Y9_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X1Y9_N1BEG[3] ,
    \Tile_X1Y9_N1BEG[2] ,
    \Tile_X1Y9_N1BEG[1] ,
    \Tile_X1Y9_N1BEG[0] }),
    .N1END({\Tile_X1Y10_N1BEG[3] ,
    \Tile_X1Y10_N1BEG[2] ,
    \Tile_X1Y10_N1BEG[1] ,
    \Tile_X1Y10_N1BEG[0] }),
    .N2BEG({\Tile_X1Y9_N2BEG[7] ,
    \Tile_X1Y9_N2BEG[6] ,
    \Tile_X1Y9_N2BEG[5] ,
    \Tile_X1Y9_N2BEG[4] ,
    \Tile_X1Y9_N2BEG[3] ,
    \Tile_X1Y9_N2BEG[2] ,
    \Tile_X1Y9_N2BEG[1] ,
    \Tile_X1Y9_N2BEG[0] }),
    .N2BEGb({\Tile_X1Y9_N2BEGb[7] ,
    \Tile_X1Y9_N2BEGb[6] ,
    \Tile_X1Y9_N2BEGb[5] ,
    \Tile_X1Y9_N2BEGb[4] ,
    \Tile_X1Y9_N2BEGb[3] ,
    \Tile_X1Y9_N2BEGb[2] ,
    \Tile_X1Y9_N2BEGb[1] ,
    \Tile_X1Y9_N2BEGb[0] }),
    .N2END({\Tile_X1Y10_N2BEGb[7] ,
    \Tile_X1Y10_N2BEGb[6] ,
    \Tile_X1Y10_N2BEGb[5] ,
    \Tile_X1Y10_N2BEGb[4] ,
    \Tile_X1Y10_N2BEGb[3] ,
    \Tile_X1Y10_N2BEGb[2] ,
    \Tile_X1Y10_N2BEGb[1] ,
    \Tile_X1Y10_N2BEGb[0] }),
    .N2MID({\Tile_X1Y10_N2BEG[7] ,
    \Tile_X1Y10_N2BEG[6] ,
    \Tile_X1Y10_N2BEG[5] ,
    \Tile_X1Y10_N2BEG[4] ,
    \Tile_X1Y10_N2BEG[3] ,
    \Tile_X1Y10_N2BEG[2] ,
    \Tile_X1Y10_N2BEG[1] ,
    \Tile_X1Y10_N2BEG[0] }),
    .N4BEG({\Tile_X1Y9_N4BEG[15] ,
    \Tile_X1Y9_N4BEG[14] ,
    \Tile_X1Y9_N4BEG[13] ,
    \Tile_X1Y9_N4BEG[12] ,
    \Tile_X1Y9_N4BEG[11] ,
    \Tile_X1Y9_N4BEG[10] ,
    \Tile_X1Y9_N4BEG[9] ,
    \Tile_X1Y9_N4BEG[8] ,
    \Tile_X1Y9_N4BEG[7] ,
    \Tile_X1Y9_N4BEG[6] ,
    \Tile_X1Y9_N4BEG[5] ,
    \Tile_X1Y9_N4BEG[4] ,
    \Tile_X1Y9_N4BEG[3] ,
    \Tile_X1Y9_N4BEG[2] ,
    \Tile_X1Y9_N4BEG[1] ,
    \Tile_X1Y9_N4BEG[0] }),
    .N4END({\Tile_X1Y10_N4BEG[15] ,
    \Tile_X1Y10_N4BEG[14] ,
    \Tile_X1Y10_N4BEG[13] ,
    \Tile_X1Y10_N4BEG[12] ,
    \Tile_X1Y10_N4BEG[11] ,
    \Tile_X1Y10_N4BEG[10] ,
    \Tile_X1Y10_N4BEG[9] ,
    \Tile_X1Y10_N4BEG[8] ,
    \Tile_X1Y10_N4BEG[7] ,
    \Tile_X1Y10_N4BEG[6] ,
    \Tile_X1Y10_N4BEG[5] ,
    \Tile_X1Y10_N4BEG[4] ,
    \Tile_X1Y10_N4BEG[3] ,
    \Tile_X1Y10_N4BEG[2] ,
    \Tile_X1Y10_N4BEG[1] ,
    \Tile_X1Y10_N4BEG[0] }),
    .NN4BEG({\Tile_X1Y9_NN4BEG[15] ,
    \Tile_X1Y9_NN4BEG[14] ,
    \Tile_X1Y9_NN4BEG[13] ,
    \Tile_X1Y9_NN4BEG[12] ,
    \Tile_X1Y9_NN4BEG[11] ,
    \Tile_X1Y9_NN4BEG[10] ,
    \Tile_X1Y9_NN4BEG[9] ,
    \Tile_X1Y9_NN4BEG[8] ,
    \Tile_X1Y9_NN4BEG[7] ,
    \Tile_X1Y9_NN4BEG[6] ,
    \Tile_X1Y9_NN4BEG[5] ,
    \Tile_X1Y9_NN4BEG[4] ,
    \Tile_X1Y9_NN4BEG[3] ,
    \Tile_X1Y9_NN4BEG[2] ,
    \Tile_X1Y9_NN4BEG[1] ,
    \Tile_X1Y9_NN4BEG[0] }),
    .NN4END({\Tile_X1Y10_NN4BEG[15] ,
    \Tile_X1Y10_NN4BEG[14] ,
    \Tile_X1Y10_NN4BEG[13] ,
    \Tile_X1Y10_NN4BEG[12] ,
    \Tile_X1Y10_NN4BEG[11] ,
    \Tile_X1Y10_NN4BEG[10] ,
    \Tile_X1Y10_NN4BEG[9] ,
    \Tile_X1Y10_NN4BEG[8] ,
    \Tile_X1Y10_NN4BEG[7] ,
    \Tile_X1Y10_NN4BEG[6] ,
    \Tile_X1Y10_NN4BEG[5] ,
    \Tile_X1Y10_NN4BEG[4] ,
    \Tile_X1Y10_NN4BEG[3] ,
    \Tile_X1Y10_NN4BEG[2] ,
    \Tile_X1Y10_NN4BEG[1] ,
    \Tile_X1Y10_NN4BEG[0] }),
    .S1BEG({\Tile_X1Y9_S1BEG[3] ,
    \Tile_X1Y9_S1BEG[2] ,
    \Tile_X1Y9_S1BEG[1] ,
    \Tile_X1Y9_S1BEG[0] }),
    .S1END({\Tile_X1Y8_S1BEG[3] ,
    \Tile_X1Y8_S1BEG[2] ,
    \Tile_X1Y8_S1BEG[1] ,
    \Tile_X1Y8_S1BEG[0] }),
    .S2BEG({\Tile_X1Y9_S2BEG[7] ,
    \Tile_X1Y9_S2BEG[6] ,
    \Tile_X1Y9_S2BEG[5] ,
    \Tile_X1Y9_S2BEG[4] ,
    \Tile_X1Y9_S2BEG[3] ,
    \Tile_X1Y9_S2BEG[2] ,
    \Tile_X1Y9_S2BEG[1] ,
    \Tile_X1Y9_S2BEG[0] }),
    .S2BEGb({\Tile_X1Y9_S2BEGb[7] ,
    \Tile_X1Y9_S2BEGb[6] ,
    \Tile_X1Y9_S2BEGb[5] ,
    \Tile_X1Y9_S2BEGb[4] ,
    \Tile_X1Y9_S2BEGb[3] ,
    \Tile_X1Y9_S2BEGb[2] ,
    \Tile_X1Y9_S2BEGb[1] ,
    \Tile_X1Y9_S2BEGb[0] }),
    .S2END({\Tile_X1Y8_S2BEGb[7] ,
    \Tile_X1Y8_S2BEGb[6] ,
    \Tile_X1Y8_S2BEGb[5] ,
    \Tile_X1Y8_S2BEGb[4] ,
    \Tile_X1Y8_S2BEGb[3] ,
    \Tile_X1Y8_S2BEGb[2] ,
    \Tile_X1Y8_S2BEGb[1] ,
    \Tile_X1Y8_S2BEGb[0] }),
    .S2MID({\Tile_X1Y8_S2BEG[7] ,
    \Tile_X1Y8_S2BEG[6] ,
    \Tile_X1Y8_S2BEG[5] ,
    \Tile_X1Y8_S2BEG[4] ,
    \Tile_X1Y8_S2BEG[3] ,
    \Tile_X1Y8_S2BEG[2] ,
    \Tile_X1Y8_S2BEG[1] ,
    \Tile_X1Y8_S2BEG[0] }),
    .S4BEG({\Tile_X1Y9_S4BEG[15] ,
    \Tile_X1Y9_S4BEG[14] ,
    \Tile_X1Y9_S4BEG[13] ,
    \Tile_X1Y9_S4BEG[12] ,
    \Tile_X1Y9_S4BEG[11] ,
    \Tile_X1Y9_S4BEG[10] ,
    \Tile_X1Y9_S4BEG[9] ,
    \Tile_X1Y9_S4BEG[8] ,
    \Tile_X1Y9_S4BEG[7] ,
    \Tile_X1Y9_S4BEG[6] ,
    \Tile_X1Y9_S4BEG[5] ,
    \Tile_X1Y9_S4BEG[4] ,
    \Tile_X1Y9_S4BEG[3] ,
    \Tile_X1Y9_S4BEG[2] ,
    \Tile_X1Y9_S4BEG[1] ,
    \Tile_X1Y9_S4BEG[0] }),
    .S4END({\Tile_X1Y8_S4BEG[15] ,
    \Tile_X1Y8_S4BEG[14] ,
    \Tile_X1Y8_S4BEG[13] ,
    \Tile_X1Y8_S4BEG[12] ,
    \Tile_X1Y8_S4BEG[11] ,
    \Tile_X1Y8_S4BEG[10] ,
    \Tile_X1Y8_S4BEG[9] ,
    \Tile_X1Y8_S4BEG[8] ,
    \Tile_X1Y8_S4BEG[7] ,
    \Tile_X1Y8_S4BEG[6] ,
    \Tile_X1Y8_S4BEG[5] ,
    \Tile_X1Y8_S4BEG[4] ,
    \Tile_X1Y8_S4BEG[3] ,
    \Tile_X1Y8_S4BEG[2] ,
    \Tile_X1Y8_S4BEG[1] ,
    \Tile_X1Y8_S4BEG[0] }),
    .SS4BEG({\Tile_X1Y9_SS4BEG[15] ,
    \Tile_X1Y9_SS4BEG[14] ,
    \Tile_X1Y9_SS4BEG[13] ,
    \Tile_X1Y9_SS4BEG[12] ,
    \Tile_X1Y9_SS4BEG[11] ,
    \Tile_X1Y9_SS4BEG[10] ,
    \Tile_X1Y9_SS4BEG[9] ,
    \Tile_X1Y9_SS4BEG[8] ,
    \Tile_X1Y9_SS4BEG[7] ,
    \Tile_X1Y9_SS4BEG[6] ,
    \Tile_X1Y9_SS4BEG[5] ,
    \Tile_X1Y9_SS4BEG[4] ,
    \Tile_X1Y9_SS4BEG[3] ,
    \Tile_X1Y9_SS4BEG[2] ,
    \Tile_X1Y9_SS4BEG[1] ,
    \Tile_X1Y9_SS4BEG[0] }),
    .SS4END({\Tile_X1Y8_SS4BEG[15] ,
    \Tile_X1Y8_SS4BEG[14] ,
    \Tile_X1Y8_SS4BEG[13] ,
    \Tile_X1Y8_SS4BEG[12] ,
    \Tile_X1Y8_SS4BEG[11] ,
    \Tile_X1Y8_SS4BEG[10] ,
    \Tile_X1Y8_SS4BEG[9] ,
    \Tile_X1Y8_SS4BEG[8] ,
    \Tile_X1Y8_SS4BEG[7] ,
    \Tile_X1Y8_SS4BEG[6] ,
    \Tile_X1Y8_SS4BEG[5] ,
    \Tile_X1Y8_SS4BEG[4] ,
    \Tile_X1Y8_SS4BEG[3] ,
    \Tile_X1Y8_SS4BEG[2] ,
    \Tile_X1Y8_SS4BEG[1] ,
    \Tile_X1Y8_SS4BEG[0] }),
    .W1BEG({\Tile_X1Y9_W1BEG[3] ,
    \Tile_X1Y9_W1BEG[2] ,
    \Tile_X1Y9_W1BEG[1] ,
    \Tile_X1Y9_W1BEG[0] }),
    .W1END({\Tile_X2Y9_W1BEG[3] ,
    \Tile_X2Y9_W1BEG[2] ,
    \Tile_X2Y9_W1BEG[1] ,
    \Tile_X2Y9_W1BEG[0] }),
    .W2BEG({\Tile_X1Y9_W2BEG[7] ,
    \Tile_X1Y9_W2BEG[6] ,
    \Tile_X1Y9_W2BEG[5] ,
    \Tile_X1Y9_W2BEG[4] ,
    \Tile_X1Y9_W2BEG[3] ,
    \Tile_X1Y9_W2BEG[2] ,
    \Tile_X1Y9_W2BEG[1] ,
    \Tile_X1Y9_W2BEG[0] }),
    .W2BEGb({\Tile_X1Y9_W2BEGb[7] ,
    \Tile_X1Y9_W2BEGb[6] ,
    \Tile_X1Y9_W2BEGb[5] ,
    \Tile_X1Y9_W2BEGb[4] ,
    \Tile_X1Y9_W2BEGb[3] ,
    \Tile_X1Y9_W2BEGb[2] ,
    \Tile_X1Y9_W2BEGb[1] ,
    \Tile_X1Y9_W2BEGb[0] }),
    .W2END({\Tile_X2Y9_W2BEGb[7] ,
    \Tile_X2Y9_W2BEGb[6] ,
    \Tile_X2Y9_W2BEGb[5] ,
    \Tile_X2Y9_W2BEGb[4] ,
    \Tile_X2Y9_W2BEGb[3] ,
    \Tile_X2Y9_W2BEGb[2] ,
    \Tile_X2Y9_W2BEGb[1] ,
    \Tile_X2Y9_W2BEGb[0] }),
    .W2MID({\Tile_X2Y9_W2BEG[7] ,
    \Tile_X2Y9_W2BEG[6] ,
    \Tile_X2Y9_W2BEG[5] ,
    \Tile_X2Y9_W2BEG[4] ,
    \Tile_X2Y9_W2BEG[3] ,
    \Tile_X2Y9_W2BEG[2] ,
    \Tile_X2Y9_W2BEG[1] ,
    \Tile_X2Y9_W2BEG[0] }),
    .W6BEG({\Tile_X1Y9_W6BEG[11] ,
    \Tile_X1Y9_W6BEG[10] ,
    \Tile_X1Y9_W6BEG[9] ,
    \Tile_X1Y9_W6BEG[8] ,
    \Tile_X1Y9_W6BEG[7] ,
    \Tile_X1Y9_W6BEG[6] ,
    \Tile_X1Y9_W6BEG[5] ,
    \Tile_X1Y9_W6BEG[4] ,
    \Tile_X1Y9_W6BEG[3] ,
    \Tile_X1Y9_W6BEG[2] ,
    \Tile_X1Y9_W6BEG[1] ,
    \Tile_X1Y9_W6BEG[0] }),
    .W6END({\Tile_X2Y9_W6BEG[11] ,
    \Tile_X2Y9_W6BEG[10] ,
    \Tile_X2Y9_W6BEG[9] ,
    \Tile_X2Y9_W6BEG[8] ,
    \Tile_X2Y9_W6BEG[7] ,
    \Tile_X2Y9_W6BEG[6] ,
    \Tile_X2Y9_W6BEG[5] ,
    \Tile_X2Y9_W6BEG[4] ,
    \Tile_X2Y9_W6BEG[3] ,
    \Tile_X2Y9_W6BEG[2] ,
    \Tile_X2Y9_W6BEG[1] ,
    \Tile_X2Y9_W6BEG[0] }),
    .WW4BEG({\Tile_X1Y9_WW4BEG[15] ,
    \Tile_X1Y9_WW4BEG[14] ,
    \Tile_X1Y9_WW4BEG[13] ,
    \Tile_X1Y9_WW4BEG[12] ,
    \Tile_X1Y9_WW4BEG[11] ,
    \Tile_X1Y9_WW4BEG[10] ,
    \Tile_X1Y9_WW4BEG[9] ,
    \Tile_X1Y9_WW4BEG[8] ,
    \Tile_X1Y9_WW4BEG[7] ,
    \Tile_X1Y9_WW4BEG[6] ,
    \Tile_X1Y9_WW4BEG[5] ,
    \Tile_X1Y9_WW4BEG[4] ,
    \Tile_X1Y9_WW4BEG[3] ,
    \Tile_X1Y9_WW4BEG[2] ,
    \Tile_X1Y9_WW4BEG[1] ,
    \Tile_X1Y9_WW4BEG[0] }),
    .WW4END({\Tile_X2Y9_WW4BEG[15] ,
    \Tile_X2Y9_WW4BEG[14] ,
    \Tile_X2Y9_WW4BEG[13] ,
    \Tile_X2Y9_WW4BEG[12] ,
    \Tile_X2Y9_WW4BEG[11] ,
    \Tile_X2Y9_WW4BEG[10] ,
    \Tile_X2Y9_WW4BEG[9] ,
    \Tile_X2Y9_WW4BEG[8] ,
    \Tile_X2Y9_WW4BEG[7] ,
    \Tile_X2Y9_WW4BEG[6] ,
    \Tile_X2Y9_WW4BEG[5] ,
    \Tile_X2Y9_WW4BEG[4] ,
    \Tile_X2Y9_WW4BEG[3] ,
    \Tile_X2Y9_WW4BEG[2] ,
    \Tile_X2Y9_WW4BEG[1] ,
    \Tile_X2Y9_WW4BEG[0] }));
 N_IO Tile_X2Y0_N_IO (.A_I_top(Tile_X2Y0_A_I_top),
    .A_O_top(Tile_X2Y0_A_O_top),
    .A_T_top(Tile_X2Y0_A_T_top),
    .A_config_C_bit0(Tile_X2Y0_A_config_C_bit0),
    .A_config_C_bit1(Tile_X2Y0_A_config_C_bit1),
    .A_config_C_bit2(Tile_X2Y0_A_config_C_bit2),
    .A_config_C_bit3(Tile_X2Y0_A_config_C_bit3),
    .B_I_top(Tile_X2Y0_B_I_top),
    .B_O_top(Tile_X2Y0_B_O_top),
    .B_T_top(Tile_X2Y0_B_T_top),
    .B_config_C_bit0(Tile_X2Y0_B_config_C_bit0),
    .B_config_C_bit1(Tile_X2Y0_B_config_C_bit1),
    .B_config_C_bit2(Tile_X2Y0_B_config_C_bit2),
    .B_config_C_bit3(Tile_X2Y0_B_config_C_bit3),
    .Ci(Tile_X2Y1_Co),
    .UserCLK(Tile_X2Y1_UserCLKo),
    .UserCLKo(Tile_X2Y0_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .FrameData({\Tile_X1Y0_FrameData_O[31] ,
    \Tile_X1Y0_FrameData_O[30] ,
    \Tile_X1Y0_FrameData_O[29] ,
    \Tile_X1Y0_FrameData_O[28] ,
    \Tile_X1Y0_FrameData_O[27] ,
    \Tile_X1Y0_FrameData_O[26] ,
    \Tile_X1Y0_FrameData_O[25] ,
    \Tile_X1Y0_FrameData_O[24] ,
    \Tile_X1Y0_FrameData_O[23] ,
    \Tile_X1Y0_FrameData_O[22] ,
    \Tile_X1Y0_FrameData_O[21] ,
    \Tile_X1Y0_FrameData_O[20] ,
    \Tile_X1Y0_FrameData_O[19] ,
    \Tile_X1Y0_FrameData_O[18] ,
    \Tile_X1Y0_FrameData_O[17] ,
    \Tile_X1Y0_FrameData_O[16] ,
    \Tile_X1Y0_FrameData_O[15] ,
    \Tile_X1Y0_FrameData_O[14] ,
    \Tile_X1Y0_FrameData_O[13] ,
    \Tile_X1Y0_FrameData_O[12] ,
    \Tile_X1Y0_FrameData_O[11] ,
    \Tile_X1Y0_FrameData_O[10] ,
    \Tile_X1Y0_FrameData_O[9] ,
    \Tile_X1Y0_FrameData_O[8] ,
    \Tile_X1Y0_FrameData_O[7] ,
    \Tile_X1Y0_FrameData_O[6] ,
    \Tile_X1Y0_FrameData_O[5] ,
    \Tile_X1Y0_FrameData_O[4] ,
    \Tile_X1Y0_FrameData_O[3] ,
    \Tile_X1Y0_FrameData_O[2] ,
    \Tile_X1Y0_FrameData_O[1] ,
    \Tile_X1Y0_FrameData_O[0] }),
    .FrameData_O({\Tile_X2Y0_FrameData_O[31] ,
    \Tile_X2Y0_FrameData_O[30] ,
    \Tile_X2Y0_FrameData_O[29] ,
    \Tile_X2Y0_FrameData_O[28] ,
    \Tile_X2Y0_FrameData_O[27] ,
    \Tile_X2Y0_FrameData_O[26] ,
    \Tile_X2Y0_FrameData_O[25] ,
    \Tile_X2Y0_FrameData_O[24] ,
    \Tile_X2Y0_FrameData_O[23] ,
    \Tile_X2Y0_FrameData_O[22] ,
    \Tile_X2Y0_FrameData_O[21] ,
    \Tile_X2Y0_FrameData_O[20] ,
    \Tile_X2Y0_FrameData_O[19] ,
    \Tile_X2Y0_FrameData_O[18] ,
    \Tile_X2Y0_FrameData_O[17] ,
    \Tile_X2Y0_FrameData_O[16] ,
    \Tile_X2Y0_FrameData_O[15] ,
    \Tile_X2Y0_FrameData_O[14] ,
    \Tile_X2Y0_FrameData_O[13] ,
    \Tile_X2Y0_FrameData_O[12] ,
    \Tile_X2Y0_FrameData_O[11] ,
    \Tile_X2Y0_FrameData_O[10] ,
    \Tile_X2Y0_FrameData_O[9] ,
    \Tile_X2Y0_FrameData_O[8] ,
    \Tile_X2Y0_FrameData_O[7] ,
    \Tile_X2Y0_FrameData_O[6] ,
    \Tile_X2Y0_FrameData_O[5] ,
    \Tile_X2Y0_FrameData_O[4] ,
    \Tile_X2Y0_FrameData_O[3] ,
    \Tile_X2Y0_FrameData_O[2] ,
    \Tile_X2Y0_FrameData_O[1] ,
    \Tile_X2Y0_FrameData_O[0] }),
    .FrameStrobe({\Tile_X2Y1_FrameStrobe_O[19] ,
    \Tile_X2Y1_FrameStrobe_O[18] ,
    \Tile_X2Y1_FrameStrobe_O[17] ,
    \Tile_X2Y1_FrameStrobe_O[16] ,
    \Tile_X2Y1_FrameStrobe_O[15] ,
    \Tile_X2Y1_FrameStrobe_O[14] ,
    \Tile_X2Y1_FrameStrobe_O[13] ,
    \Tile_X2Y1_FrameStrobe_O[12] ,
    \Tile_X2Y1_FrameStrobe_O[11] ,
    \Tile_X2Y1_FrameStrobe_O[10] ,
    \Tile_X2Y1_FrameStrobe_O[9] ,
    \Tile_X2Y1_FrameStrobe_O[8] ,
    \Tile_X2Y1_FrameStrobe_O[7] ,
    \Tile_X2Y1_FrameStrobe_O[6] ,
    \Tile_X2Y1_FrameStrobe_O[5] ,
    \Tile_X2Y1_FrameStrobe_O[4] ,
    \Tile_X2Y1_FrameStrobe_O[3] ,
    \Tile_X2Y1_FrameStrobe_O[2] ,
    \Tile_X2Y1_FrameStrobe_O[1] ,
    \Tile_X2Y1_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X2Y0_FrameStrobe_O[19] ,
    \Tile_X2Y0_FrameStrobe_O[18] ,
    \Tile_X2Y0_FrameStrobe_O[17] ,
    \Tile_X2Y0_FrameStrobe_O[16] ,
    \Tile_X2Y0_FrameStrobe_O[15] ,
    \Tile_X2Y0_FrameStrobe_O[14] ,
    \Tile_X2Y0_FrameStrobe_O[13] ,
    \Tile_X2Y0_FrameStrobe_O[12] ,
    \Tile_X2Y0_FrameStrobe_O[11] ,
    \Tile_X2Y0_FrameStrobe_O[10] ,
    \Tile_X2Y0_FrameStrobe_O[9] ,
    \Tile_X2Y0_FrameStrobe_O[8] ,
    \Tile_X2Y0_FrameStrobe_O[7] ,
    \Tile_X2Y0_FrameStrobe_O[6] ,
    \Tile_X2Y0_FrameStrobe_O[5] ,
    \Tile_X2Y0_FrameStrobe_O[4] ,
    \Tile_X2Y0_FrameStrobe_O[3] ,
    \Tile_X2Y0_FrameStrobe_O[2] ,
    \Tile_X2Y0_FrameStrobe_O[1] ,
    \Tile_X2Y0_FrameStrobe_O[0] }),
    .N1END({\Tile_X2Y1_N1BEG[3] ,
    \Tile_X2Y1_N1BEG[2] ,
    \Tile_X2Y1_N1BEG[1] ,
    \Tile_X2Y1_N1BEG[0] }),
    .N2END({\Tile_X2Y1_N2BEGb[7] ,
    \Tile_X2Y1_N2BEGb[6] ,
    \Tile_X2Y1_N2BEGb[5] ,
    \Tile_X2Y1_N2BEGb[4] ,
    \Tile_X2Y1_N2BEGb[3] ,
    \Tile_X2Y1_N2BEGb[2] ,
    \Tile_X2Y1_N2BEGb[1] ,
    \Tile_X2Y1_N2BEGb[0] }),
    .N2MID({\Tile_X2Y1_N2BEG[7] ,
    \Tile_X2Y1_N2BEG[6] ,
    \Tile_X2Y1_N2BEG[5] ,
    \Tile_X2Y1_N2BEG[4] ,
    \Tile_X2Y1_N2BEG[3] ,
    \Tile_X2Y1_N2BEG[2] ,
    \Tile_X2Y1_N2BEG[1] ,
    \Tile_X2Y1_N2BEG[0] }),
    .N4END({\Tile_X2Y1_N4BEG[15] ,
    \Tile_X2Y1_N4BEG[14] ,
    \Tile_X2Y1_N4BEG[13] ,
    \Tile_X2Y1_N4BEG[12] ,
    \Tile_X2Y1_N4BEG[11] ,
    \Tile_X2Y1_N4BEG[10] ,
    \Tile_X2Y1_N4BEG[9] ,
    \Tile_X2Y1_N4BEG[8] ,
    \Tile_X2Y1_N4BEG[7] ,
    \Tile_X2Y1_N4BEG[6] ,
    \Tile_X2Y1_N4BEG[5] ,
    \Tile_X2Y1_N4BEG[4] ,
    \Tile_X2Y1_N4BEG[3] ,
    \Tile_X2Y1_N4BEG[2] ,
    \Tile_X2Y1_N4BEG[1] ,
    \Tile_X2Y1_N4BEG[0] }),
    .NN4END({\Tile_X2Y1_NN4BEG[15] ,
    \Tile_X2Y1_NN4BEG[14] ,
    \Tile_X2Y1_NN4BEG[13] ,
    \Tile_X2Y1_NN4BEG[12] ,
    \Tile_X2Y1_NN4BEG[11] ,
    \Tile_X2Y1_NN4BEG[10] ,
    \Tile_X2Y1_NN4BEG[9] ,
    \Tile_X2Y1_NN4BEG[8] ,
    \Tile_X2Y1_NN4BEG[7] ,
    \Tile_X2Y1_NN4BEG[6] ,
    \Tile_X2Y1_NN4BEG[5] ,
    \Tile_X2Y1_NN4BEG[4] ,
    \Tile_X2Y1_NN4BEG[3] ,
    \Tile_X2Y1_NN4BEG[2] ,
    \Tile_X2Y1_NN4BEG[1] ,
    \Tile_X2Y1_NN4BEG[0] }),
    .S1BEG({\Tile_X2Y0_S1BEG[3] ,
    \Tile_X2Y0_S1BEG[2] ,
    \Tile_X2Y0_S1BEG[1] ,
    \Tile_X2Y0_S1BEG[0] }),
    .S2BEG({\Tile_X2Y0_S2BEG[7] ,
    \Tile_X2Y0_S2BEG[6] ,
    \Tile_X2Y0_S2BEG[5] ,
    \Tile_X2Y0_S2BEG[4] ,
    \Tile_X2Y0_S2BEG[3] ,
    \Tile_X2Y0_S2BEG[2] ,
    \Tile_X2Y0_S2BEG[1] ,
    \Tile_X2Y0_S2BEG[0] }),
    .S2BEGb({\Tile_X2Y0_S2BEGb[7] ,
    \Tile_X2Y0_S2BEGb[6] ,
    \Tile_X2Y0_S2BEGb[5] ,
    \Tile_X2Y0_S2BEGb[4] ,
    \Tile_X2Y0_S2BEGb[3] ,
    \Tile_X2Y0_S2BEGb[2] ,
    \Tile_X2Y0_S2BEGb[1] ,
    \Tile_X2Y0_S2BEGb[0] }),
    .S4BEG({\Tile_X2Y0_S4BEG[15] ,
    \Tile_X2Y0_S4BEG[14] ,
    \Tile_X2Y0_S4BEG[13] ,
    \Tile_X2Y0_S4BEG[12] ,
    \Tile_X2Y0_S4BEG[11] ,
    \Tile_X2Y0_S4BEG[10] ,
    \Tile_X2Y0_S4BEG[9] ,
    \Tile_X2Y0_S4BEG[8] ,
    \Tile_X2Y0_S4BEG[7] ,
    \Tile_X2Y0_S4BEG[6] ,
    \Tile_X2Y0_S4BEG[5] ,
    \Tile_X2Y0_S4BEG[4] ,
    \Tile_X2Y0_S4BEG[3] ,
    \Tile_X2Y0_S4BEG[2] ,
    \Tile_X2Y0_S4BEG[1] ,
    \Tile_X2Y0_S4BEG[0] }),
    .SS4BEG({\Tile_X2Y0_SS4BEG[15] ,
    \Tile_X2Y0_SS4BEG[14] ,
    \Tile_X2Y0_SS4BEG[13] ,
    \Tile_X2Y0_SS4BEG[12] ,
    \Tile_X2Y0_SS4BEG[11] ,
    \Tile_X2Y0_SS4BEG[10] ,
    \Tile_X2Y0_SS4BEG[9] ,
    \Tile_X2Y0_SS4BEG[8] ,
    \Tile_X2Y0_SS4BEG[7] ,
    \Tile_X2Y0_SS4BEG[6] ,
    \Tile_X2Y0_SS4BEG[5] ,
    \Tile_X2Y0_SS4BEG[4] ,
    \Tile_X2Y0_SS4BEG[3] ,
    \Tile_X2Y0_SS4BEG[2] ,
    \Tile_X2Y0_SS4BEG[1] ,
    \Tile_X2Y0_SS4BEG[0] }));
 LUT4AB Tile_X2Y10_LUT4AB (.Ci(Tile_X2Y11_Co),
    .Co(Tile_X2Y10_Co),
    .UserCLK(Tile_X2Y11_UserCLKo),
    .UserCLKo(Tile_X2Y10_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X2Y10_E1BEG[3] ,
    \Tile_X2Y10_E1BEG[2] ,
    \Tile_X2Y10_E1BEG[1] ,
    \Tile_X2Y10_E1BEG[0] }),
    .E1END({\Tile_X1Y10_E1BEG[3] ,
    \Tile_X1Y10_E1BEG[2] ,
    \Tile_X1Y10_E1BEG[1] ,
    \Tile_X1Y10_E1BEG[0] }),
    .E2BEG({\Tile_X2Y10_E2BEG[7] ,
    \Tile_X2Y10_E2BEG[6] ,
    \Tile_X2Y10_E2BEG[5] ,
    \Tile_X2Y10_E2BEG[4] ,
    \Tile_X2Y10_E2BEG[3] ,
    \Tile_X2Y10_E2BEG[2] ,
    \Tile_X2Y10_E2BEG[1] ,
    \Tile_X2Y10_E2BEG[0] }),
    .E2BEGb({\Tile_X2Y10_E2BEGb[7] ,
    \Tile_X2Y10_E2BEGb[6] ,
    \Tile_X2Y10_E2BEGb[5] ,
    \Tile_X2Y10_E2BEGb[4] ,
    \Tile_X2Y10_E2BEGb[3] ,
    \Tile_X2Y10_E2BEGb[2] ,
    \Tile_X2Y10_E2BEGb[1] ,
    \Tile_X2Y10_E2BEGb[0] }),
    .E2END({\Tile_X1Y10_E2BEGb[7] ,
    \Tile_X1Y10_E2BEGb[6] ,
    \Tile_X1Y10_E2BEGb[5] ,
    \Tile_X1Y10_E2BEGb[4] ,
    \Tile_X1Y10_E2BEGb[3] ,
    \Tile_X1Y10_E2BEGb[2] ,
    \Tile_X1Y10_E2BEGb[1] ,
    \Tile_X1Y10_E2BEGb[0] }),
    .E2MID({\Tile_X1Y10_E2BEG[7] ,
    \Tile_X1Y10_E2BEG[6] ,
    \Tile_X1Y10_E2BEG[5] ,
    \Tile_X1Y10_E2BEG[4] ,
    \Tile_X1Y10_E2BEG[3] ,
    \Tile_X1Y10_E2BEG[2] ,
    \Tile_X1Y10_E2BEG[1] ,
    \Tile_X1Y10_E2BEG[0] }),
    .E6BEG({\Tile_X2Y10_E6BEG[11] ,
    \Tile_X2Y10_E6BEG[10] ,
    \Tile_X2Y10_E6BEG[9] ,
    \Tile_X2Y10_E6BEG[8] ,
    \Tile_X2Y10_E6BEG[7] ,
    \Tile_X2Y10_E6BEG[6] ,
    \Tile_X2Y10_E6BEG[5] ,
    \Tile_X2Y10_E6BEG[4] ,
    \Tile_X2Y10_E6BEG[3] ,
    \Tile_X2Y10_E6BEG[2] ,
    \Tile_X2Y10_E6BEG[1] ,
    \Tile_X2Y10_E6BEG[0] }),
    .E6END({\Tile_X1Y10_E6BEG[11] ,
    \Tile_X1Y10_E6BEG[10] ,
    \Tile_X1Y10_E6BEG[9] ,
    \Tile_X1Y10_E6BEG[8] ,
    \Tile_X1Y10_E6BEG[7] ,
    \Tile_X1Y10_E6BEG[6] ,
    \Tile_X1Y10_E6BEG[5] ,
    \Tile_X1Y10_E6BEG[4] ,
    \Tile_X1Y10_E6BEG[3] ,
    \Tile_X1Y10_E6BEG[2] ,
    \Tile_X1Y10_E6BEG[1] ,
    \Tile_X1Y10_E6BEG[0] }),
    .EE4BEG({\Tile_X2Y10_EE4BEG[15] ,
    \Tile_X2Y10_EE4BEG[14] ,
    \Tile_X2Y10_EE4BEG[13] ,
    \Tile_X2Y10_EE4BEG[12] ,
    \Tile_X2Y10_EE4BEG[11] ,
    \Tile_X2Y10_EE4BEG[10] ,
    \Tile_X2Y10_EE4BEG[9] ,
    \Tile_X2Y10_EE4BEG[8] ,
    \Tile_X2Y10_EE4BEG[7] ,
    \Tile_X2Y10_EE4BEG[6] ,
    \Tile_X2Y10_EE4BEG[5] ,
    \Tile_X2Y10_EE4BEG[4] ,
    \Tile_X2Y10_EE4BEG[3] ,
    \Tile_X2Y10_EE4BEG[2] ,
    \Tile_X2Y10_EE4BEG[1] ,
    \Tile_X2Y10_EE4BEG[0] }),
    .EE4END({\Tile_X1Y10_EE4BEG[15] ,
    \Tile_X1Y10_EE4BEG[14] ,
    \Tile_X1Y10_EE4BEG[13] ,
    \Tile_X1Y10_EE4BEG[12] ,
    \Tile_X1Y10_EE4BEG[11] ,
    \Tile_X1Y10_EE4BEG[10] ,
    \Tile_X1Y10_EE4BEG[9] ,
    \Tile_X1Y10_EE4BEG[8] ,
    \Tile_X1Y10_EE4BEG[7] ,
    \Tile_X1Y10_EE4BEG[6] ,
    \Tile_X1Y10_EE4BEG[5] ,
    \Tile_X1Y10_EE4BEG[4] ,
    \Tile_X1Y10_EE4BEG[3] ,
    \Tile_X1Y10_EE4BEG[2] ,
    \Tile_X1Y10_EE4BEG[1] ,
    \Tile_X1Y10_EE4BEG[0] }),
    .FrameData({\Tile_X1Y10_FrameData_O[31] ,
    \Tile_X1Y10_FrameData_O[30] ,
    \Tile_X1Y10_FrameData_O[29] ,
    \Tile_X1Y10_FrameData_O[28] ,
    \Tile_X1Y10_FrameData_O[27] ,
    \Tile_X1Y10_FrameData_O[26] ,
    \Tile_X1Y10_FrameData_O[25] ,
    \Tile_X1Y10_FrameData_O[24] ,
    \Tile_X1Y10_FrameData_O[23] ,
    \Tile_X1Y10_FrameData_O[22] ,
    \Tile_X1Y10_FrameData_O[21] ,
    \Tile_X1Y10_FrameData_O[20] ,
    \Tile_X1Y10_FrameData_O[19] ,
    \Tile_X1Y10_FrameData_O[18] ,
    \Tile_X1Y10_FrameData_O[17] ,
    \Tile_X1Y10_FrameData_O[16] ,
    \Tile_X1Y10_FrameData_O[15] ,
    \Tile_X1Y10_FrameData_O[14] ,
    \Tile_X1Y10_FrameData_O[13] ,
    \Tile_X1Y10_FrameData_O[12] ,
    \Tile_X1Y10_FrameData_O[11] ,
    \Tile_X1Y10_FrameData_O[10] ,
    \Tile_X1Y10_FrameData_O[9] ,
    \Tile_X1Y10_FrameData_O[8] ,
    \Tile_X1Y10_FrameData_O[7] ,
    \Tile_X1Y10_FrameData_O[6] ,
    \Tile_X1Y10_FrameData_O[5] ,
    \Tile_X1Y10_FrameData_O[4] ,
    \Tile_X1Y10_FrameData_O[3] ,
    \Tile_X1Y10_FrameData_O[2] ,
    \Tile_X1Y10_FrameData_O[1] ,
    \Tile_X1Y10_FrameData_O[0] }),
    .FrameData_O({\Tile_X2Y10_FrameData_O[31] ,
    \Tile_X2Y10_FrameData_O[30] ,
    \Tile_X2Y10_FrameData_O[29] ,
    \Tile_X2Y10_FrameData_O[28] ,
    \Tile_X2Y10_FrameData_O[27] ,
    \Tile_X2Y10_FrameData_O[26] ,
    \Tile_X2Y10_FrameData_O[25] ,
    \Tile_X2Y10_FrameData_O[24] ,
    \Tile_X2Y10_FrameData_O[23] ,
    \Tile_X2Y10_FrameData_O[22] ,
    \Tile_X2Y10_FrameData_O[21] ,
    \Tile_X2Y10_FrameData_O[20] ,
    \Tile_X2Y10_FrameData_O[19] ,
    \Tile_X2Y10_FrameData_O[18] ,
    \Tile_X2Y10_FrameData_O[17] ,
    \Tile_X2Y10_FrameData_O[16] ,
    \Tile_X2Y10_FrameData_O[15] ,
    \Tile_X2Y10_FrameData_O[14] ,
    \Tile_X2Y10_FrameData_O[13] ,
    \Tile_X2Y10_FrameData_O[12] ,
    \Tile_X2Y10_FrameData_O[11] ,
    \Tile_X2Y10_FrameData_O[10] ,
    \Tile_X2Y10_FrameData_O[9] ,
    \Tile_X2Y10_FrameData_O[8] ,
    \Tile_X2Y10_FrameData_O[7] ,
    \Tile_X2Y10_FrameData_O[6] ,
    \Tile_X2Y10_FrameData_O[5] ,
    \Tile_X2Y10_FrameData_O[4] ,
    \Tile_X2Y10_FrameData_O[3] ,
    \Tile_X2Y10_FrameData_O[2] ,
    \Tile_X2Y10_FrameData_O[1] ,
    \Tile_X2Y10_FrameData_O[0] }),
    .FrameStrobe({\Tile_X2Y11_FrameStrobe_O[19] ,
    \Tile_X2Y11_FrameStrobe_O[18] ,
    \Tile_X2Y11_FrameStrobe_O[17] ,
    \Tile_X2Y11_FrameStrobe_O[16] ,
    \Tile_X2Y11_FrameStrobe_O[15] ,
    \Tile_X2Y11_FrameStrobe_O[14] ,
    \Tile_X2Y11_FrameStrobe_O[13] ,
    \Tile_X2Y11_FrameStrobe_O[12] ,
    \Tile_X2Y11_FrameStrobe_O[11] ,
    \Tile_X2Y11_FrameStrobe_O[10] ,
    \Tile_X2Y11_FrameStrobe_O[9] ,
    \Tile_X2Y11_FrameStrobe_O[8] ,
    \Tile_X2Y11_FrameStrobe_O[7] ,
    \Tile_X2Y11_FrameStrobe_O[6] ,
    \Tile_X2Y11_FrameStrobe_O[5] ,
    \Tile_X2Y11_FrameStrobe_O[4] ,
    \Tile_X2Y11_FrameStrobe_O[3] ,
    \Tile_X2Y11_FrameStrobe_O[2] ,
    \Tile_X2Y11_FrameStrobe_O[1] ,
    \Tile_X2Y11_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X2Y10_FrameStrobe_O[19] ,
    \Tile_X2Y10_FrameStrobe_O[18] ,
    \Tile_X2Y10_FrameStrobe_O[17] ,
    \Tile_X2Y10_FrameStrobe_O[16] ,
    \Tile_X2Y10_FrameStrobe_O[15] ,
    \Tile_X2Y10_FrameStrobe_O[14] ,
    \Tile_X2Y10_FrameStrobe_O[13] ,
    \Tile_X2Y10_FrameStrobe_O[12] ,
    \Tile_X2Y10_FrameStrobe_O[11] ,
    \Tile_X2Y10_FrameStrobe_O[10] ,
    \Tile_X2Y10_FrameStrobe_O[9] ,
    \Tile_X2Y10_FrameStrobe_O[8] ,
    \Tile_X2Y10_FrameStrobe_O[7] ,
    \Tile_X2Y10_FrameStrobe_O[6] ,
    \Tile_X2Y10_FrameStrobe_O[5] ,
    \Tile_X2Y10_FrameStrobe_O[4] ,
    \Tile_X2Y10_FrameStrobe_O[3] ,
    \Tile_X2Y10_FrameStrobe_O[2] ,
    \Tile_X2Y10_FrameStrobe_O[1] ,
    \Tile_X2Y10_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X2Y10_N1BEG[3] ,
    \Tile_X2Y10_N1BEG[2] ,
    \Tile_X2Y10_N1BEG[1] ,
    \Tile_X2Y10_N1BEG[0] }),
    .N1END({\Tile_X2Y11_N1BEG[3] ,
    \Tile_X2Y11_N1BEG[2] ,
    \Tile_X2Y11_N1BEG[1] ,
    \Tile_X2Y11_N1BEG[0] }),
    .N2BEG({\Tile_X2Y10_N2BEG[7] ,
    \Tile_X2Y10_N2BEG[6] ,
    \Tile_X2Y10_N2BEG[5] ,
    \Tile_X2Y10_N2BEG[4] ,
    \Tile_X2Y10_N2BEG[3] ,
    \Tile_X2Y10_N2BEG[2] ,
    \Tile_X2Y10_N2BEG[1] ,
    \Tile_X2Y10_N2BEG[0] }),
    .N2BEGb({\Tile_X2Y10_N2BEGb[7] ,
    \Tile_X2Y10_N2BEGb[6] ,
    \Tile_X2Y10_N2BEGb[5] ,
    \Tile_X2Y10_N2BEGb[4] ,
    \Tile_X2Y10_N2BEGb[3] ,
    \Tile_X2Y10_N2BEGb[2] ,
    \Tile_X2Y10_N2BEGb[1] ,
    \Tile_X2Y10_N2BEGb[0] }),
    .N2END({\Tile_X2Y11_N2BEGb[7] ,
    \Tile_X2Y11_N2BEGb[6] ,
    \Tile_X2Y11_N2BEGb[5] ,
    \Tile_X2Y11_N2BEGb[4] ,
    \Tile_X2Y11_N2BEGb[3] ,
    \Tile_X2Y11_N2BEGb[2] ,
    \Tile_X2Y11_N2BEGb[1] ,
    \Tile_X2Y11_N2BEGb[0] }),
    .N2MID({\Tile_X2Y11_N2BEG[7] ,
    \Tile_X2Y11_N2BEG[6] ,
    \Tile_X2Y11_N2BEG[5] ,
    \Tile_X2Y11_N2BEG[4] ,
    \Tile_X2Y11_N2BEG[3] ,
    \Tile_X2Y11_N2BEG[2] ,
    \Tile_X2Y11_N2BEG[1] ,
    \Tile_X2Y11_N2BEG[0] }),
    .N4BEG({\Tile_X2Y10_N4BEG[15] ,
    \Tile_X2Y10_N4BEG[14] ,
    \Tile_X2Y10_N4BEG[13] ,
    \Tile_X2Y10_N4BEG[12] ,
    \Tile_X2Y10_N4BEG[11] ,
    \Tile_X2Y10_N4BEG[10] ,
    \Tile_X2Y10_N4BEG[9] ,
    \Tile_X2Y10_N4BEG[8] ,
    \Tile_X2Y10_N4BEG[7] ,
    \Tile_X2Y10_N4BEG[6] ,
    \Tile_X2Y10_N4BEG[5] ,
    \Tile_X2Y10_N4BEG[4] ,
    \Tile_X2Y10_N4BEG[3] ,
    \Tile_X2Y10_N4BEG[2] ,
    \Tile_X2Y10_N4BEG[1] ,
    \Tile_X2Y10_N4BEG[0] }),
    .N4END({\Tile_X2Y11_N4BEG[15] ,
    \Tile_X2Y11_N4BEG[14] ,
    \Tile_X2Y11_N4BEG[13] ,
    \Tile_X2Y11_N4BEG[12] ,
    \Tile_X2Y11_N4BEG[11] ,
    \Tile_X2Y11_N4BEG[10] ,
    \Tile_X2Y11_N4BEG[9] ,
    \Tile_X2Y11_N4BEG[8] ,
    \Tile_X2Y11_N4BEG[7] ,
    \Tile_X2Y11_N4BEG[6] ,
    \Tile_X2Y11_N4BEG[5] ,
    \Tile_X2Y11_N4BEG[4] ,
    \Tile_X2Y11_N4BEG[3] ,
    \Tile_X2Y11_N4BEG[2] ,
    \Tile_X2Y11_N4BEG[1] ,
    \Tile_X2Y11_N4BEG[0] }),
    .NN4BEG({\Tile_X2Y10_NN4BEG[15] ,
    \Tile_X2Y10_NN4BEG[14] ,
    \Tile_X2Y10_NN4BEG[13] ,
    \Tile_X2Y10_NN4BEG[12] ,
    \Tile_X2Y10_NN4BEG[11] ,
    \Tile_X2Y10_NN4BEG[10] ,
    \Tile_X2Y10_NN4BEG[9] ,
    \Tile_X2Y10_NN4BEG[8] ,
    \Tile_X2Y10_NN4BEG[7] ,
    \Tile_X2Y10_NN4BEG[6] ,
    \Tile_X2Y10_NN4BEG[5] ,
    \Tile_X2Y10_NN4BEG[4] ,
    \Tile_X2Y10_NN4BEG[3] ,
    \Tile_X2Y10_NN4BEG[2] ,
    \Tile_X2Y10_NN4BEG[1] ,
    \Tile_X2Y10_NN4BEG[0] }),
    .NN4END({\Tile_X2Y11_NN4BEG[15] ,
    \Tile_X2Y11_NN4BEG[14] ,
    \Tile_X2Y11_NN4BEG[13] ,
    \Tile_X2Y11_NN4BEG[12] ,
    \Tile_X2Y11_NN4BEG[11] ,
    \Tile_X2Y11_NN4BEG[10] ,
    \Tile_X2Y11_NN4BEG[9] ,
    \Tile_X2Y11_NN4BEG[8] ,
    \Tile_X2Y11_NN4BEG[7] ,
    \Tile_X2Y11_NN4BEG[6] ,
    \Tile_X2Y11_NN4BEG[5] ,
    \Tile_X2Y11_NN4BEG[4] ,
    \Tile_X2Y11_NN4BEG[3] ,
    \Tile_X2Y11_NN4BEG[2] ,
    \Tile_X2Y11_NN4BEG[1] ,
    \Tile_X2Y11_NN4BEG[0] }),
    .S1BEG({\Tile_X2Y10_S1BEG[3] ,
    \Tile_X2Y10_S1BEG[2] ,
    \Tile_X2Y10_S1BEG[1] ,
    \Tile_X2Y10_S1BEG[0] }),
    .S1END({\Tile_X2Y9_S1BEG[3] ,
    \Tile_X2Y9_S1BEG[2] ,
    \Tile_X2Y9_S1BEG[1] ,
    \Tile_X2Y9_S1BEG[0] }),
    .S2BEG({\Tile_X2Y10_S2BEG[7] ,
    \Tile_X2Y10_S2BEG[6] ,
    \Tile_X2Y10_S2BEG[5] ,
    \Tile_X2Y10_S2BEG[4] ,
    \Tile_X2Y10_S2BEG[3] ,
    \Tile_X2Y10_S2BEG[2] ,
    \Tile_X2Y10_S2BEG[1] ,
    \Tile_X2Y10_S2BEG[0] }),
    .S2BEGb({\Tile_X2Y10_S2BEGb[7] ,
    \Tile_X2Y10_S2BEGb[6] ,
    \Tile_X2Y10_S2BEGb[5] ,
    \Tile_X2Y10_S2BEGb[4] ,
    \Tile_X2Y10_S2BEGb[3] ,
    \Tile_X2Y10_S2BEGb[2] ,
    \Tile_X2Y10_S2BEGb[1] ,
    \Tile_X2Y10_S2BEGb[0] }),
    .S2END({\Tile_X2Y9_S2BEGb[7] ,
    \Tile_X2Y9_S2BEGb[6] ,
    \Tile_X2Y9_S2BEGb[5] ,
    \Tile_X2Y9_S2BEGb[4] ,
    \Tile_X2Y9_S2BEGb[3] ,
    \Tile_X2Y9_S2BEGb[2] ,
    \Tile_X2Y9_S2BEGb[1] ,
    \Tile_X2Y9_S2BEGb[0] }),
    .S2MID({\Tile_X2Y9_S2BEG[7] ,
    \Tile_X2Y9_S2BEG[6] ,
    \Tile_X2Y9_S2BEG[5] ,
    \Tile_X2Y9_S2BEG[4] ,
    \Tile_X2Y9_S2BEG[3] ,
    \Tile_X2Y9_S2BEG[2] ,
    \Tile_X2Y9_S2BEG[1] ,
    \Tile_X2Y9_S2BEG[0] }),
    .S4BEG({\Tile_X2Y10_S4BEG[15] ,
    \Tile_X2Y10_S4BEG[14] ,
    \Tile_X2Y10_S4BEG[13] ,
    \Tile_X2Y10_S4BEG[12] ,
    \Tile_X2Y10_S4BEG[11] ,
    \Tile_X2Y10_S4BEG[10] ,
    \Tile_X2Y10_S4BEG[9] ,
    \Tile_X2Y10_S4BEG[8] ,
    \Tile_X2Y10_S4BEG[7] ,
    \Tile_X2Y10_S4BEG[6] ,
    \Tile_X2Y10_S4BEG[5] ,
    \Tile_X2Y10_S4BEG[4] ,
    \Tile_X2Y10_S4BEG[3] ,
    \Tile_X2Y10_S4BEG[2] ,
    \Tile_X2Y10_S4BEG[1] ,
    \Tile_X2Y10_S4BEG[0] }),
    .S4END({\Tile_X2Y9_S4BEG[15] ,
    \Tile_X2Y9_S4BEG[14] ,
    \Tile_X2Y9_S4BEG[13] ,
    \Tile_X2Y9_S4BEG[12] ,
    \Tile_X2Y9_S4BEG[11] ,
    \Tile_X2Y9_S4BEG[10] ,
    \Tile_X2Y9_S4BEG[9] ,
    \Tile_X2Y9_S4BEG[8] ,
    \Tile_X2Y9_S4BEG[7] ,
    \Tile_X2Y9_S4BEG[6] ,
    \Tile_X2Y9_S4BEG[5] ,
    \Tile_X2Y9_S4BEG[4] ,
    \Tile_X2Y9_S4BEG[3] ,
    \Tile_X2Y9_S4BEG[2] ,
    \Tile_X2Y9_S4BEG[1] ,
    \Tile_X2Y9_S4BEG[0] }),
    .SS4BEG({\Tile_X2Y10_SS4BEG[15] ,
    \Tile_X2Y10_SS4BEG[14] ,
    \Tile_X2Y10_SS4BEG[13] ,
    \Tile_X2Y10_SS4BEG[12] ,
    \Tile_X2Y10_SS4BEG[11] ,
    \Tile_X2Y10_SS4BEG[10] ,
    \Tile_X2Y10_SS4BEG[9] ,
    \Tile_X2Y10_SS4BEG[8] ,
    \Tile_X2Y10_SS4BEG[7] ,
    \Tile_X2Y10_SS4BEG[6] ,
    \Tile_X2Y10_SS4BEG[5] ,
    \Tile_X2Y10_SS4BEG[4] ,
    \Tile_X2Y10_SS4BEG[3] ,
    \Tile_X2Y10_SS4BEG[2] ,
    \Tile_X2Y10_SS4BEG[1] ,
    \Tile_X2Y10_SS4BEG[0] }),
    .SS4END({\Tile_X2Y9_SS4BEG[15] ,
    \Tile_X2Y9_SS4BEG[14] ,
    \Tile_X2Y9_SS4BEG[13] ,
    \Tile_X2Y9_SS4BEG[12] ,
    \Tile_X2Y9_SS4BEG[11] ,
    \Tile_X2Y9_SS4BEG[10] ,
    \Tile_X2Y9_SS4BEG[9] ,
    \Tile_X2Y9_SS4BEG[8] ,
    \Tile_X2Y9_SS4BEG[7] ,
    \Tile_X2Y9_SS4BEG[6] ,
    \Tile_X2Y9_SS4BEG[5] ,
    \Tile_X2Y9_SS4BEG[4] ,
    \Tile_X2Y9_SS4BEG[3] ,
    \Tile_X2Y9_SS4BEG[2] ,
    \Tile_X2Y9_SS4BEG[1] ,
    \Tile_X2Y9_SS4BEG[0] }),
    .W1BEG({\Tile_X2Y10_W1BEG[3] ,
    \Tile_X2Y10_W1BEG[2] ,
    \Tile_X2Y10_W1BEG[1] ,
    \Tile_X2Y10_W1BEG[0] }),
    .W1END({\Tile_X3Y10_W1BEG[3] ,
    \Tile_X3Y10_W1BEG[2] ,
    \Tile_X3Y10_W1BEG[1] ,
    \Tile_X3Y10_W1BEG[0] }),
    .W2BEG({\Tile_X2Y10_W2BEG[7] ,
    \Tile_X2Y10_W2BEG[6] ,
    \Tile_X2Y10_W2BEG[5] ,
    \Tile_X2Y10_W2BEG[4] ,
    \Tile_X2Y10_W2BEG[3] ,
    \Tile_X2Y10_W2BEG[2] ,
    \Tile_X2Y10_W2BEG[1] ,
    \Tile_X2Y10_W2BEG[0] }),
    .W2BEGb({\Tile_X2Y10_W2BEGb[7] ,
    \Tile_X2Y10_W2BEGb[6] ,
    \Tile_X2Y10_W2BEGb[5] ,
    \Tile_X2Y10_W2BEGb[4] ,
    \Tile_X2Y10_W2BEGb[3] ,
    \Tile_X2Y10_W2BEGb[2] ,
    \Tile_X2Y10_W2BEGb[1] ,
    \Tile_X2Y10_W2BEGb[0] }),
    .W2END({\Tile_X3Y10_W2BEGb[7] ,
    \Tile_X3Y10_W2BEGb[6] ,
    \Tile_X3Y10_W2BEGb[5] ,
    \Tile_X3Y10_W2BEGb[4] ,
    \Tile_X3Y10_W2BEGb[3] ,
    \Tile_X3Y10_W2BEGb[2] ,
    \Tile_X3Y10_W2BEGb[1] ,
    \Tile_X3Y10_W2BEGb[0] }),
    .W2MID({\Tile_X3Y10_W2BEG[7] ,
    \Tile_X3Y10_W2BEG[6] ,
    \Tile_X3Y10_W2BEG[5] ,
    \Tile_X3Y10_W2BEG[4] ,
    \Tile_X3Y10_W2BEG[3] ,
    \Tile_X3Y10_W2BEG[2] ,
    \Tile_X3Y10_W2BEG[1] ,
    \Tile_X3Y10_W2BEG[0] }),
    .W6BEG({\Tile_X2Y10_W6BEG[11] ,
    \Tile_X2Y10_W6BEG[10] ,
    \Tile_X2Y10_W6BEG[9] ,
    \Tile_X2Y10_W6BEG[8] ,
    \Tile_X2Y10_W6BEG[7] ,
    \Tile_X2Y10_W6BEG[6] ,
    \Tile_X2Y10_W6BEG[5] ,
    \Tile_X2Y10_W6BEG[4] ,
    \Tile_X2Y10_W6BEG[3] ,
    \Tile_X2Y10_W6BEG[2] ,
    \Tile_X2Y10_W6BEG[1] ,
    \Tile_X2Y10_W6BEG[0] }),
    .W6END({\Tile_X3Y10_W6BEG[11] ,
    \Tile_X3Y10_W6BEG[10] ,
    \Tile_X3Y10_W6BEG[9] ,
    \Tile_X3Y10_W6BEG[8] ,
    \Tile_X3Y10_W6BEG[7] ,
    \Tile_X3Y10_W6BEG[6] ,
    \Tile_X3Y10_W6BEG[5] ,
    \Tile_X3Y10_W6BEG[4] ,
    \Tile_X3Y10_W6BEG[3] ,
    \Tile_X3Y10_W6BEG[2] ,
    \Tile_X3Y10_W6BEG[1] ,
    \Tile_X3Y10_W6BEG[0] }),
    .WW4BEG({\Tile_X2Y10_WW4BEG[15] ,
    \Tile_X2Y10_WW4BEG[14] ,
    \Tile_X2Y10_WW4BEG[13] ,
    \Tile_X2Y10_WW4BEG[12] ,
    \Tile_X2Y10_WW4BEG[11] ,
    \Tile_X2Y10_WW4BEG[10] ,
    \Tile_X2Y10_WW4BEG[9] ,
    \Tile_X2Y10_WW4BEG[8] ,
    \Tile_X2Y10_WW4BEG[7] ,
    \Tile_X2Y10_WW4BEG[6] ,
    \Tile_X2Y10_WW4BEG[5] ,
    \Tile_X2Y10_WW4BEG[4] ,
    \Tile_X2Y10_WW4BEG[3] ,
    \Tile_X2Y10_WW4BEG[2] ,
    \Tile_X2Y10_WW4BEG[1] ,
    \Tile_X2Y10_WW4BEG[0] }),
    .WW4END({\Tile_X3Y10_WW4BEG[15] ,
    \Tile_X3Y10_WW4BEG[14] ,
    \Tile_X3Y10_WW4BEG[13] ,
    \Tile_X3Y10_WW4BEG[12] ,
    \Tile_X3Y10_WW4BEG[11] ,
    \Tile_X3Y10_WW4BEG[10] ,
    \Tile_X3Y10_WW4BEG[9] ,
    \Tile_X3Y10_WW4BEG[8] ,
    \Tile_X3Y10_WW4BEG[7] ,
    \Tile_X3Y10_WW4BEG[6] ,
    \Tile_X3Y10_WW4BEG[5] ,
    \Tile_X3Y10_WW4BEG[4] ,
    \Tile_X3Y10_WW4BEG[3] ,
    \Tile_X3Y10_WW4BEG[2] ,
    \Tile_X3Y10_WW4BEG[1] ,
    \Tile_X3Y10_WW4BEG[0] }));
 LUT4AB Tile_X2Y11_LUT4AB (.Ci(Tile_X2Y12_Co),
    .Co(Tile_X2Y11_Co),
    .UserCLK(Tile_X2Y12_UserCLKo),
    .UserCLKo(Tile_X2Y11_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X2Y11_E1BEG[3] ,
    \Tile_X2Y11_E1BEG[2] ,
    \Tile_X2Y11_E1BEG[1] ,
    \Tile_X2Y11_E1BEG[0] }),
    .E1END({\Tile_X1Y11_E1BEG[3] ,
    \Tile_X1Y11_E1BEG[2] ,
    \Tile_X1Y11_E1BEG[1] ,
    \Tile_X1Y11_E1BEG[0] }),
    .E2BEG({\Tile_X2Y11_E2BEG[7] ,
    \Tile_X2Y11_E2BEG[6] ,
    \Tile_X2Y11_E2BEG[5] ,
    \Tile_X2Y11_E2BEG[4] ,
    \Tile_X2Y11_E2BEG[3] ,
    \Tile_X2Y11_E2BEG[2] ,
    \Tile_X2Y11_E2BEG[1] ,
    \Tile_X2Y11_E2BEG[0] }),
    .E2BEGb({\Tile_X2Y11_E2BEGb[7] ,
    \Tile_X2Y11_E2BEGb[6] ,
    \Tile_X2Y11_E2BEGb[5] ,
    \Tile_X2Y11_E2BEGb[4] ,
    \Tile_X2Y11_E2BEGb[3] ,
    \Tile_X2Y11_E2BEGb[2] ,
    \Tile_X2Y11_E2BEGb[1] ,
    \Tile_X2Y11_E2BEGb[0] }),
    .E2END({\Tile_X1Y11_E2BEGb[7] ,
    \Tile_X1Y11_E2BEGb[6] ,
    \Tile_X1Y11_E2BEGb[5] ,
    \Tile_X1Y11_E2BEGb[4] ,
    \Tile_X1Y11_E2BEGb[3] ,
    \Tile_X1Y11_E2BEGb[2] ,
    \Tile_X1Y11_E2BEGb[1] ,
    \Tile_X1Y11_E2BEGb[0] }),
    .E2MID({\Tile_X1Y11_E2BEG[7] ,
    \Tile_X1Y11_E2BEG[6] ,
    \Tile_X1Y11_E2BEG[5] ,
    \Tile_X1Y11_E2BEG[4] ,
    \Tile_X1Y11_E2BEG[3] ,
    \Tile_X1Y11_E2BEG[2] ,
    \Tile_X1Y11_E2BEG[1] ,
    \Tile_X1Y11_E2BEG[0] }),
    .E6BEG({\Tile_X2Y11_E6BEG[11] ,
    \Tile_X2Y11_E6BEG[10] ,
    \Tile_X2Y11_E6BEG[9] ,
    \Tile_X2Y11_E6BEG[8] ,
    \Tile_X2Y11_E6BEG[7] ,
    \Tile_X2Y11_E6BEG[6] ,
    \Tile_X2Y11_E6BEG[5] ,
    \Tile_X2Y11_E6BEG[4] ,
    \Tile_X2Y11_E6BEG[3] ,
    \Tile_X2Y11_E6BEG[2] ,
    \Tile_X2Y11_E6BEG[1] ,
    \Tile_X2Y11_E6BEG[0] }),
    .E6END({\Tile_X1Y11_E6BEG[11] ,
    \Tile_X1Y11_E6BEG[10] ,
    \Tile_X1Y11_E6BEG[9] ,
    \Tile_X1Y11_E6BEG[8] ,
    \Tile_X1Y11_E6BEG[7] ,
    \Tile_X1Y11_E6BEG[6] ,
    \Tile_X1Y11_E6BEG[5] ,
    \Tile_X1Y11_E6BEG[4] ,
    \Tile_X1Y11_E6BEG[3] ,
    \Tile_X1Y11_E6BEG[2] ,
    \Tile_X1Y11_E6BEG[1] ,
    \Tile_X1Y11_E6BEG[0] }),
    .EE4BEG({\Tile_X2Y11_EE4BEG[15] ,
    \Tile_X2Y11_EE4BEG[14] ,
    \Tile_X2Y11_EE4BEG[13] ,
    \Tile_X2Y11_EE4BEG[12] ,
    \Tile_X2Y11_EE4BEG[11] ,
    \Tile_X2Y11_EE4BEG[10] ,
    \Tile_X2Y11_EE4BEG[9] ,
    \Tile_X2Y11_EE4BEG[8] ,
    \Tile_X2Y11_EE4BEG[7] ,
    \Tile_X2Y11_EE4BEG[6] ,
    \Tile_X2Y11_EE4BEG[5] ,
    \Tile_X2Y11_EE4BEG[4] ,
    \Tile_X2Y11_EE4BEG[3] ,
    \Tile_X2Y11_EE4BEG[2] ,
    \Tile_X2Y11_EE4BEG[1] ,
    \Tile_X2Y11_EE4BEG[0] }),
    .EE4END({\Tile_X1Y11_EE4BEG[15] ,
    \Tile_X1Y11_EE4BEG[14] ,
    \Tile_X1Y11_EE4BEG[13] ,
    \Tile_X1Y11_EE4BEG[12] ,
    \Tile_X1Y11_EE4BEG[11] ,
    \Tile_X1Y11_EE4BEG[10] ,
    \Tile_X1Y11_EE4BEG[9] ,
    \Tile_X1Y11_EE4BEG[8] ,
    \Tile_X1Y11_EE4BEG[7] ,
    \Tile_X1Y11_EE4BEG[6] ,
    \Tile_X1Y11_EE4BEG[5] ,
    \Tile_X1Y11_EE4BEG[4] ,
    \Tile_X1Y11_EE4BEG[3] ,
    \Tile_X1Y11_EE4BEG[2] ,
    \Tile_X1Y11_EE4BEG[1] ,
    \Tile_X1Y11_EE4BEG[0] }),
    .FrameData({\Tile_X1Y11_FrameData_O[31] ,
    \Tile_X1Y11_FrameData_O[30] ,
    \Tile_X1Y11_FrameData_O[29] ,
    \Tile_X1Y11_FrameData_O[28] ,
    \Tile_X1Y11_FrameData_O[27] ,
    \Tile_X1Y11_FrameData_O[26] ,
    \Tile_X1Y11_FrameData_O[25] ,
    \Tile_X1Y11_FrameData_O[24] ,
    \Tile_X1Y11_FrameData_O[23] ,
    \Tile_X1Y11_FrameData_O[22] ,
    \Tile_X1Y11_FrameData_O[21] ,
    \Tile_X1Y11_FrameData_O[20] ,
    \Tile_X1Y11_FrameData_O[19] ,
    \Tile_X1Y11_FrameData_O[18] ,
    \Tile_X1Y11_FrameData_O[17] ,
    \Tile_X1Y11_FrameData_O[16] ,
    \Tile_X1Y11_FrameData_O[15] ,
    \Tile_X1Y11_FrameData_O[14] ,
    \Tile_X1Y11_FrameData_O[13] ,
    \Tile_X1Y11_FrameData_O[12] ,
    \Tile_X1Y11_FrameData_O[11] ,
    \Tile_X1Y11_FrameData_O[10] ,
    \Tile_X1Y11_FrameData_O[9] ,
    \Tile_X1Y11_FrameData_O[8] ,
    \Tile_X1Y11_FrameData_O[7] ,
    \Tile_X1Y11_FrameData_O[6] ,
    \Tile_X1Y11_FrameData_O[5] ,
    \Tile_X1Y11_FrameData_O[4] ,
    \Tile_X1Y11_FrameData_O[3] ,
    \Tile_X1Y11_FrameData_O[2] ,
    \Tile_X1Y11_FrameData_O[1] ,
    \Tile_X1Y11_FrameData_O[0] }),
    .FrameData_O({\Tile_X2Y11_FrameData_O[31] ,
    \Tile_X2Y11_FrameData_O[30] ,
    \Tile_X2Y11_FrameData_O[29] ,
    \Tile_X2Y11_FrameData_O[28] ,
    \Tile_X2Y11_FrameData_O[27] ,
    \Tile_X2Y11_FrameData_O[26] ,
    \Tile_X2Y11_FrameData_O[25] ,
    \Tile_X2Y11_FrameData_O[24] ,
    \Tile_X2Y11_FrameData_O[23] ,
    \Tile_X2Y11_FrameData_O[22] ,
    \Tile_X2Y11_FrameData_O[21] ,
    \Tile_X2Y11_FrameData_O[20] ,
    \Tile_X2Y11_FrameData_O[19] ,
    \Tile_X2Y11_FrameData_O[18] ,
    \Tile_X2Y11_FrameData_O[17] ,
    \Tile_X2Y11_FrameData_O[16] ,
    \Tile_X2Y11_FrameData_O[15] ,
    \Tile_X2Y11_FrameData_O[14] ,
    \Tile_X2Y11_FrameData_O[13] ,
    \Tile_X2Y11_FrameData_O[12] ,
    \Tile_X2Y11_FrameData_O[11] ,
    \Tile_X2Y11_FrameData_O[10] ,
    \Tile_X2Y11_FrameData_O[9] ,
    \Tile_X2Y11_FrameData_O[8] ,
    \Tile_X2Y11_FrameData_O[7] ,
    \Tile_X2Y11_FrameData_O[6] ,
    \Tile_X2Y11_FrameData_O[5] ,
    \Tile_X2Y11_FrameData_O[4] ,
    \Tile_X2Y11_FrameData_O[3] ,
    \Tile_X2Y11_FrameData_O[2] ,
    \Tile_X2Y11_FrameData_O[1] ,
    \Tile_X2Y11_FrameData_O[0] }),
    .FrameStrobe({\Tile_X2Y12_FrameStrobe_O[19] ,
    \Tile_X2Y12_FrameStrobe_O[18] ,
    \Tile_X2Y12_FrameStrobe_O[17] ,
    \Tile_X2Y12_FrameStrobe_O[16] ,
    \Tile_X2Y12_FrameStrobe_O[15] ,
    \Tile_X2Y12_FrameStrobe_O[14] ,
    \Tile_X2Y12_FrameStrobe_O[13] ,
    \Tile_X2Y12_FrameStrobe_O[12] ,
    \Tile_X2Y12_FrameStrobe_O[11] ,
    \Tile_X2Y12_FrameStrobe_O[10] ,
    \Tile_X2Y12_FrameStrobe_O[9] ,
    \Tile_X2Y12_FrameStrobe_O[8] ,
    \Tile_X2Y12_FrameStrobe_O[7] ,
    \Tile_X2Y12_FrameStrobe_O[6] ,
    \Tile_X2Y12_FrameStrobe_O[5] ,
    \Tile_X2Y12_FrameStrobe_O[4] ,
    \Tile_X2Y12_FrameStrobe_O[3] ,
    \Tile_X2Y12_FrameStrobe_O[2] ,
    \Tile_X2Y12_FrameStrobe_O[1] ,
    \Tile_X2Y12_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X2Y11_FrameStrobe_O[19] ,
    \Tile_X2Y11_FrameStrobe_O[18] ,
    \Tile_X2Y11_FrameStrobe_O[17] ,
    \Tile_X2Y11_FrameStrobe_O[16] ,
    \Tile_X2Y11_FrameStrobe_O[15] ,
    \Tile_X2Y11_FrameStrobe_O[14] ,
    \Tile_X2Y11_FrameStrobe_O[13] ,
    \Tile_X2Y11_FrameStrobe_O[12] ,
    \Tile_X2Y11_FrameStrobe_O[11] ,
    \Tile_X2Y11_FrameStrobe_O[10] ,
    \Tile_X2Y11_FrameStrobe_O[9] ,
    \Tile_X2Y11_FrameStrobe_O[8] ,
    \Tile_X2Y11_FrameStrobe_O[7] ,
    \Tile_X2Y11_FrameStrobe_O[6] ,
    \Tile_X2Y11_FrameStrobe_O[5] ,
    \Tile_X2Y11_FrameStrobe_O[4] ,
    \Tile_X2Y11_FrameStrobe_O[3] ,
    \Tile_X2Y11_FrameStrobe_O[2] ,
    \Tile_X2Y11_FrameStrobe_O[1] ,
    \Tile_X2Y11_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X2Y11_N1BEG[3] ,
    \Tile_X2Y11_N1BEG[2] ,
    \Tile_X2Y11_N1BEG[1] ,
    \Tile_X2Y11_N1BEG[0] }),
    .N1END({\Tile_X2Y12_N1BEG[3] ,
    \Tile_X2Y12_N1BEG[2] ,
    \Tile_X2Y12_N1BEG[1] ,
    \Tile_X2Y12_N1BEG[0] }),
    .N2BEG({\Tile_X2Y11_N2BEG[7] ,
    \Tile_X2Y11_N2BEG[6] ,
    \Tile_X2Y11_N2BEG[5] ,
    \Tile_X2Y11_N2BEG[4] ,
    \Tile_X2Y11_N2BEG[3] ,
    \Tile_X2Y11_N2BEG[2] ,
    \Tile_X2Y11_N2BEG[1] ,
    \Tile_X2Y11_N2BEG[0] }),
    .N2BEGb({\Tile_X2Y11_N2BEGb[7] ,
    \Tile_X2Y11_N2BEGb[6] ,
    \Tile_X2Y11_N2BEGb[5] ,
    \Tile_X2Y11_N2BEGb[4] ,
    \Tile_X2Y11_N2BEGb[3] ,
    \Tile_X2Y11_N2BEGb[2] ,
    \Tile_X2Y11_N2BEGb[1] ,
    \Tile_X2Y11_N2BEGb[0] }),
    .N2END({\Tile_X2Y12_N2BEGb[7] ,
    \Tile_X2Y12_N2BEGb[6] ,
    \Tile_X2Y12_N2BEGb[5] ,
    \Tile_X2Y12_N2BEGb[4] ,
    \Tile_X2Y12_N2BEGb[3] ,
    \Tile_X2Y12_N2BEGb[2] ,
    \Tile_X2Y12_N2BEGb[1] ,
    \Tile_X2Y12_N2BEGb[0] }),
    .N2MID({\Tile_X2Y12_N2BEG[7] ,
    \Tile_X2Y12_N2BEG[6] ,
    \Tile_X2Y12_N2BEG[5] ,
    \Tile_X2Y12_N2BEG[4] ,
    \Tile_X2Y12_N2BEG[3] ,
    \Tile_X2Y12_N2BEG[2] ,
    \Tile_X2Y12_N2BEG[1] ,
    \Tile_X2Y12_N2BEG[0] }),
    .N4BEG({\Tile_X2Y11_N4BEG[15] ,
    \Tile_X2Y11_N4BEG[14] ,
    \Tile_X2Y11_N4BEG[13] ,
    \Tile_X2Y11_N4BEG[12] ,
    \Tile_X2Y11_N4BEG[11] ,
    \Tile_X2Y11_N4BEG[10] ,
    \Tile_X2Y11_N4BEG[9] ,
    \Tile_X2Y11_N4BEG[8] ,
    \Tile_X2Y11_N4BEG[7] ,
    \Tile_X2Y11_N4BEG[6] ,
    \Tile_X2Y11_N4BEG[5] ,
    \Tile_X2Y11_N4BEG[4] ,
    \Tile_X2Y11_N4BEG[3] ,
    \Tile_X2Y11_N4BEG[2] ,
    \Tile_X2Y11_N4BEG[1] ,
    \Tile_X2Y11_N4BEG[0] }),
    .N4END({\Tile_X2Y12_N4BEG[15] ,
    \Tile_X2Y12_N4BEG[14] ,
    \Tile_X2Y12_N4BEG[13] ,
    \Tile_X2Y12_N4BEG[12] ,
    \Tile_X2Y12_N4BEG[11] ,
    \Tile_X2Y12_N4BEG[10] ,
    \Tile_X2Y12_N4BEG[9] ,
    \Tile_X2Y12_N4BEG[8] ,
    \Tile_X2Y12_N4BEG[7] ,
    \Tile_X2Y12_N4BEG[6] ,
    \Tile_X2Y12_N4BEG[5] ,
    \Tile_X2Y12_N4BEG[4] ,
    \Tile_X2Y12_N4BEG[3] ,
    \Tile_X2Y12_N4BEG[2] ,
    \Tile_X2Y12_N4BEG[1] ,
    \Tile_X2Y12_N4BEG[0] }),
    .NN4BEG({\Tile_X2Y11_NN4BEG[15] ,
    \Tile_X2Y11_NN4BEG[14] ,
    \Tile_X2Y11_NN4BEG[13] ,
    \Tile_X2Y11_NN4BEG[12] ,
    \Tile_X2Y11_NN4BEG[11] ,
    \Tile_X2Y11_NN4BEG[10] ,
    \Tile_X2Y11_NN4BEG[9] ,
    \Tile_X2Y11_NN4BEG[8] ,
    \Tile_X2Y11_NN4BEG[7] ,
    \Tile_X2Y11_NN4BEG[6] ,
    \Tile_X2Y11_NN4BEG[5] ,
    \Tile_X2Y11_NN4BEG[4] ,
    \Tile_X2Y11_NN4BEG[3] ,
    \Tile_X2Y11_NN4BEG[2] ,
    \Tile_X2Y11_NN4BEG[1] ,
    \Tile_X2Y11_NN4BEG[0] }),
    .NN4END({\Tile_X2Y12_NN4BEG[15] ,
    \Tile_X2Y12_NN4BEG[14] ,
    \Tile_X2Y12_NN4BEG[13] ,
    \Tile_X2Y12_NN4BEG[12] ,
    \Tile_X2Y12_NN4BEG[11] ,
    \Tile_X2Y12_NN4BEG[10] ,
    \Tile_X2Y12_NN4BEG[9] ,
    \Tile_X2Y12_NN4BEG[8] ,
    \Tile_X2Y12_NN4BEG[7] ,
    \Tile_X2Y12_NN4BEG[6] ,
    \Tile_X2Y12_NN4BEG[5] ,
    \Tile_X2Y12_NN4BEG[4] ,
    \Tile_X2Y12_NN4BEG[3] ,
    \Tile_X2Y12_NN4BEG[2] ,
    \Tile_X2Y12_NN4BEG[1] ,
    \Tile_X2Y12_NN4BEG[0] }),
    .S1BEG({\Tile_X2Y11_S1BEG[3] ,
    \Tile_X2Y11_S1BEG[2] ,
    \Tile_X2Y11_S1BEG[1] ,
    \Tile_X2Y11_S1BEG[0] }),
    .S1END({\Tile_X2Y10_S1BEG[3] ,
    \Tile_X2Y10_S1BEG[2] ,
    \Tile_X2Y10_S1BEG[1] ,
    \Tile_X2Y10_S1BEG[0] }),
    .S2BEG({\Tile_X2Y11_S2BEG[7] ,
    \Tile_X2Y11_S2BEG[6] ,
    \Tile_X2Y11_S2BEG[5] ,
    \Tile_X2Y11_S2BEG[4] ,
    \Tile_X2Y11_S2BEG[3] ,
    \Tile_X2Y11_S2BEG[2] ,
    \Tile_X2Y11_S2BEG[1] ,
    \Tile_X2Y11_S2BEG[0] }),
    .S2BEGb({\Tile_X2Y11_S2BEGb[7] ,
    \Tile_X2Y11_S2BEGb[6] ,
    \Tile_X2Y11_S2BEGb[5] ,
    \Tile_X2Y11_S2BEGb[4] ,
    \Tile_X2Y11_S2BEGb[3] ,
    \Tile_X2Y11_S2BEGb[2] ,
    \Tile_X2Y11_S2BEGb[1] ,
    \Tile_X2Y11_S2BEGb[0] }),
    .S2END({\Tile_X2Y10_S2BEGb[7] ,
    \Tile_X2Y10_S2BEGb[6] ,
    \Tile_X2Y10_S2BEGb[5] ,
    \Tile_X2Y10_S2BEGb[4] ,
    \Tile_X2Y10_S2BEGb[3] ,
    \Tile_X2Y10_S2BEGb[2] ,
    \Tile_X2Y10_S2BEGb[1] ,
    \Tile_X2Y10_S2BEGb[0] }),
    .S2MID({\Tile_X2Y10_S2BEG[7] ,
    \Tile_X2Y10_S2BEG[6] ,
    \Tile_X2Y10_S2BEG[5] ,
    \Tile_X2Y10_S2BEG[4] ,
    \Tile_X2Y10_S2BEG[3] ,
    \Tile_X2Y10_S2BEG[2] ,
    \Tile_X2Y10_S2BEG[1] ,
    \Tile_X2Y10_S2BEG[0] }),
    .S4BEG({\Tile_X2Y11_S4BEG[15] ,
    \Tile_X2Y11_S4BEG[14] ,
    \Tile_X2Y11_S4BEG[13] ,
    \Tile_X2Y11_S4BEG[12] ,
    \Tile_X2Y11_S4BEG[11] ,
    \Tile_X2Y11_S4BEG[10] ,
    \Tile_X2Y11_S4BEG[9] ,
    \Tile_X2Y11_S4BEG[8] ,
    \Tile_X2Y11_S4BEG[7] ,
    \Tile_X2Y11_S4BEG[6] ,
    \Tile_X2Y11_S4BEG[5] ,
    \Tile_X2Y11_S4BEG[4] ,
    \Tile_X2Y11_S4BEG[3] ,
    \Tile_X2Y11_S4BEG[2] ,
    \Tile_X2Y11_S4BEG[1] ,
    \Tile_X2Y11_S4BEG[0] }),
    .S4END({\Tile_X2Y10_S4BEG[15] ,
    \Tile_X2Y10_S4BEG[14] ,
    \Tile_X2Y10_S4BEG[13] ,
    \Tile_X2Y10_S4BEG[12] ,
    \Tile_X2Y10_S4BEG[11] ,
    \Tile_X2Y10_S4BEG[10] ,
    \Tile_X2Y10_S4BEG[9] ,
    \Tile_X2Y10_S4BEG[8] ,
    \Tile_X2Y10_S4BEG[7] ,
    \Tile_X2Y10_S4BEG[6] ,
    \Tile_X2Y10_S4BEG[5] ,
    \Tile_X2Y10_S4BEG[4] ,
    \Tile_X2Y10_S4BEG[3] ,
    \Tile_X2Y10_S4BEG[2] ,
    \Tile_X2Y10_S4BEG[1] ,
    \Tile_X2Y10_S4BEG[0] }),
    .SS4BEG({\Tile_X2Y11_SS4BEG[15] ,
    \Tile_X2Y11_SS4BEG[14] ,
    \Tile_X2Y11_SS4BEG[13] ,
    \Tile_X2Y11_SS4BEG[12] ,
    \Tile_X2Y11_SS4BEG[11] ,
    \Tile_X2Y11_SS4BEG[10] ,
    \Tile_X2Y11_SS4BEG[9] ,
    \Tile_X2Y11_SS4BEG[8] ,
    \Tile_X2Y11_SS4BEG[7] ,
    \Tile_X2Y11_SS4BEG[6] ,
    \Tile_X2Y11_SS4BEG[5] ,
    \Tile_X2Y11_SS4BEG[4] ,
    \Tile_X2Y11_SS4BEG[3] ,
    \Tile_X2Y11_SS4BEG[2] ,
    \Tile_X2Y11_SS4BEG[1] ,
    \Tile_X2Y11_SS4BEG[0] }),
    .SS4END({\Tile_X2Y10_SS4BEG[15] ,
    \Tile_X2Y10_SS4BEG[14] ,
    \Tile_X2Y10_SS4BEG[13] ,
    \Tile_X2Y10_SS4BEG[12] ,
    \Tile_X2Y10_SS4BEG[11] ,
    \Tile_X2Y10_SS4BEG[10] ,
    \Tile_X2Y10_SS4BEG[9] ,
    \Tile_X2Y10_SS4BEG[8] ,
    \Tile_X2Y10_SS4BEG[7] ,
    \Tile_X2Y10_SS4BEG[6] ,
    \Tile_X2Y10_SS4BEG[5] ,
    \Tile_X2Y10_SS4BEG[4] ,
    \Tile_X2Y10_SS4BEG[3] ,
    \Tile_X2Y10_SS4BEG[2] ,
    \Tile_X2Y10_SS4BEG[1] ,
    \Tile_X2Y10_SS4BEG[0] }),
    .W1BEG({\Tile_X2Y11_W1BEG[3] ,
    \Tile_X2Y11_W1BEG[2] ,
    \Tile_X2Y11_W1BEG[1] ,
    \Tile_X2Y11_W1BEG[0] }),
    .W1END({\Tile_X3Y11_W1BEG[3] ,
    \Tile_X3Y11_W1BEG[2] ,
    \Tile_X3Y11_W1BEG[1] ,
    \Tile_X3Y11_W1BEG[0] }),
    .W2BEG({\Tile_X2Y11_W2BEG[7] ,
    \Tile_X2Y11_W2BEG[6] ,
    \Tile_X2Y11_W2BEG[5] ,
    \Tile_X2Y11_W2BEG[4] ,
    \Tile_X2Y11_W2BEG[3] ,
    \Tile_X2Y11_W2BEG[2] ,
    \Tile_X2Y11_W2BEG[1] ,
    \Tile_X2Y11_W2BEG[0] }),
    .W2BEGb({\Tile_X2Y11_W2BEGb[7] ,
    \Tile_X2Y11_W2BEGb[6] ,
    \Tile_X2Y11_W2BEGb[5] ,
    \Tile_X2Y11_W2BEGb[4] ,
    \Tile_X2Y11_W2BEGb[3] ,
    \Tile_X2Y11_W2BEGb[2] ,
    \Tile_X2Y11_W2BEGb[1] ,
    \Tile_X2Y11_W2BEGb[0] }),
    .W2END({\Tile_X3Y11_W2BEGb[7] ,
    \Tile_X3Y11_W2BEGb[6] ,
    \Tile_X3Y11_W2BEGb[5] ,
    \Tile_X3Y11_W2BEGb[4] ,
    \Tile_X3Y11_W2BEGb[3] ,
    \Tile_X3Y11_W2BEGb[2] ,
    \Tile_X3Y11_W2BEGb[1] ,
    \Tile_X3Y11_W2BEGb[0] }),
    .W2MID({\Tile_X3Y11_W2BEG[7] ,
    \Tile_X3Y11_W2BEG[6] ,
    \Tile_X3Y11_W2BEG[5] ,
    \Tile_X3Y11_W2BEG[4] ,
    \Tile_X3Y11_W2BEG[3] ,
    \Tile_X3Y11_W2BEG[2] ,
    \Tile_X3Y11_W2BEG[1] ,
    \Tile_X3Y11_W2BEG[0] }),
    .W6BEG({\Tile_X2Y11_W6BEG[11] ,
    \Tile_X2Y11_W6BEG[10] ,
    \Tile_X2Y11_W6BEG[9] ,
    \Tile_X2Y11_W6BEG[8] ,
    \Tile_X2Y11_W6BEG[7] ,
    \Tile_X2Y11_W6BEG[6] ,
    \Tile_X2Y11_W6BEG[5] ,
    \Tile_X2Y11_W6BEG[4] ,
    \Tile_X2Y11_W6BEG[3] ,
    \Tile_X2Y11_W6BEG[2] ,
    \Tile_X2Y11_W6BEG[1] ,
    \Tile_X2Y11_W6BEG[0] }),
    .W6END({\Tile_X3Y11_W6BEG[11] ,
    \Tile_X3Y11_W6BEG[10] ,
    \Tile_X3Y11_W6BEG[9] ,
    \Tile_X3Y11_W6BEG[8] ,
    \Tile_X3Y11_W6BEG[7] ,
    \Tile_X3Y11_W6BEG[6] ,
    \Tile_X3Y11_W6BEG[5] ,
    \Tile_X3Y11_W6BEG[4] ,
    \Tile_X3Y11_W6BEG[3] ,
    \Tile_X3Y11_W6BEG[2] ,
    \Tile_X3Y11_W6BEG[1] ,
    \Tile_X3Y11_W6BEG[0] }),
    .WW4BEG({\Tile_X2Y11_WW4BEG[15] ,
    \Tile_X2Y11_WW4BEG[14] ,
    \Tile_X2Y11_WW4BEG[13] ,
    \Tile_X2Y11_WW4BEG[12] ,
    \Tile_X2Y11_WW4BEG[11] ,
    \Tile_X2Y11_WW4BEG[10] ,
    \Tile_X2Y11_WW4BEG[9] ,
    \Tile_X2Y11_WW4BEG[8] ,
    \Tile_X2Y11_WW4BEG[7] ,
    \Tile_X2Y11_WW4BEG[6] ,
    \Tile_X2Y11_WW4BEG[5] ,
    \Tile_X2Y11_WW4BEG[4] ,
    \Tile_X2Y11_WW4BEG[3] ,
    \Tile_X2Y11_WW4BEG[2] ,
    \Tile_X2Y11_WW4BEG[1] ,
    \Tile_X2Y11_WW4BEG[0] }),
    .WW4END({\Tile_X3Y11_WW4BEG[15] ,
    \Tile_X3Y11_WW4BEG[14] ,
    \Tile_X3Y11_WW4BEG[13] ,
    \Tile_X3Y11_WW4BEG[12] ,
    \Tile_X3Y11_WW4BEG[11] ,
    \Tile_X3Y11_WW4BEG[10] ,
    \Tile_X3Y11_WW4BEG[9] ,
    \Tile_X3Y11_WW4BEG[8] ,
    \Tile_X3Y11_WW4BEG[7] ,
    \Tile_X3Y11_WW4BEG[6] ,
    \Tile_X3Y11_WW4BEG[5] ,
    \Tile_X3Y11_WW4BEG[4] ,
    \Tile_X3Y11_WW4BEG[3] ,
    \Tile_X3Y11_WW4BEG[2] ,
    \Tile_X3Y11_WW4BEG[1] ,
    \Tile_X3Y11_WW4BEG[0] }));
 LUT4AB Tile_X2Y12_LUT4AB (.Ci(Tile_X2Y13_Co),
    .Co(Tile_X2Y12_Co),
    .UserCLK(Tile_X2Y13_UserCLKo),
    .UserCLKo(Tile_X2Y12_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X2Y12_E1BEG[3] ,
    \Tile_X2Y12_E1BEG[2] ,
    \Tile_X2Y12_E1BEG[1] ,
    \Tile_X2Y12_E1BEG[0] }),
    .E1END({\Tile_X1Y12_E1BEG[3] ,
    \Tile_X1Y12_E1BEG[2] ,
    \Tile_X1Y12_E1BEG[1] ,
    \Tile_X1Y12_E1BEG[0] }),
    .E2BEG({\Tile_X2Y12_E2BEG[7] ,
    \Tile_X2Y12_E2BEG[6] ,
    \Tile_X2Y12_E2BEG[5] ,
    \Tile_X2Y12_E2BEG[4] ,
    \Tile_X2Y12_E2BEG[3] ,
    \Tile_X2Y12_E2BEG[2] ,
    \Tile_X2Y12_E2BEG[1] ,
    \Tile_X2Y12_E2BEG[0] }),
    .E2BEGb({\Tile_X2Y12_E2BEGb[7] ,
    \Tile_X2Y12_E2BEGb[6] ,
    \Tile_X2Y12_E2BEGb[5] ,
    \Tile_X2Y12_E2BEGb[4] ,
    \Tile_X2Y12_E2BEGb[3] ,
    \Tile_X2Y12_E2BEGb[2] ,
    \Tile_X2Y12_E2BEGb[1] ,
    \Tile_X2Y12_E2BEGb[0] }),
    .E2END({\Tile_X1Y12_E2BEGb[7] ,
    \Tile_X1Y12_E2BEGb[6] ,
    \Tile_X1Y12_E2BEGb[5] ,
    \Tile_X1Y12_E2BEGb[4] ,
    \Tile_X1Y12_E2BEGb[3] ,
    \Tile_X1Y12_E2BEGb[2] ,
    \Tile_X1Y12_E2BEGb[1] ,
    \Tile_X1Y12_E2BEGb[0] }),
    .E2MID({\Tile_X1Y12_E2BEG[7] ,
    \Tile_X1Y12_E2BEG[6] ,
    \Tile_X1Y12_E2BEG[5] ,
    \Tile_X1Y12_E2BEG[4] ,
    \Tile_X1Y12_E2BEG[3] ,
    \Tile_X1Y12_E2BEG[2] ,
    \Tile_X1Y12_E2BEG[1] ,
    \Tile_X1Y12_E2BEG[0] }),
    .E6BEG({\Tile_X2Y12_E6BEG[11] ,
    \Tile_X2Y12_E6BEG[10] ,
    \Tile_X2Y12_E6BEG[9] ,
    \Tile_X2Y12_E6BEG[8] ,
    \Tile_X2Y12_E6BEG[7] ,
    \Tile_X2Y12_E6BEG[6] ,
    \Tile_X2Y12_E6BEG[5] ,
    \Tile_X2Y12_E6BEG[4] ,
    \Tile_X2Y12_E6BEG[3] ,
    \Tile_X2Y12_E6BEG[2] ,
    \Tile_X2Y12_E6BEG[1] ,
    \Tile_X2Y12_E6BEG[0] }),
    .E6END({\Tile_X1Y12_E6BEG[11] ,
    \Tile_X1Y12_E6BEG[10] ,
    \Tile_X1Y12_E6BEG[9] ,
    \Tile_X1Y12_E6BEG[8] ,
    \Tile_X1Y12_E6BEG[7] ,
    \Tile_X1Y12_E6BEG[6] ,
    \Tile_X1Y12_E6BEG[5] ,
    \Tile_X1Y12_E6BEG[4] ,
    \Tile_X1Y12_E6BEG[3] ,
    \Tile_X1Y12_E6BEG[2] ,
    \Tile_X1Y12_E6BEG[1] ,
    \Tile_X1Y12_E6BEG[0] }),
    .EE4BEG({\Tile_X2Y12_EE4BEG[15] ,
    \Tile_X2Y12_EE4BEG[14] ,
    \Tile_X2Y12_EE4BEG[13] ,
    \Tile_X2Y12_EE4BEG[12] ,
    \Tile_X2Y12_EE4BEG[11] ,
    \Tile_X2Y12_EE4BEG[10] ,
    \Tile_X2Y12_EE4BEG[9] ,
    \Tile_X2Y12_EE4BEG[8] ,
    \Tile_X2Y12_EE4BEG[7] ,
    \Tile_X2Y12_EE4BEG[6] ,
    \Tile_X2Y12_EE4BEG[5] ,
    \Tile_X2Y12_EE4BEG[4] ,
    \Tile_X2Y12_EE4BEG[3] ,
    \Tile_X2Y12_EE4BEG[2] ,
    \Tile_X2Y12_EE4BEG[1] ,
    \Tile_X2Y12_EE4BEG[0] }),
    .EE4END({\Tile_X1Y12_EE4BEG[15] ,
    \Tile_X1Y12_EE4BEG[14] ,
    \Tile_X1Y12_EE4BEG[13] ,
    \Tile_X1Y12_EE4BEG[12] ,
    \Tile_X1Y12_EE4BEG[11] ,
    \Tile_X1Y12_EE4BEG[10] ,
    \Tile_X1Y12_EE4BEG[9] ,
    \Tile_X1Y12_EE4BEG[8] ,
    \Tile_X1Y12_EE4BEG[7] ,
    \Tile_X1Y12_EE4BEG[6] ,
    \Tile_X1Y12_EE4BEG[5] ,
    \Tile_X1Y12_EE4BEG[4] ,
    \Tile_X1Y12_EE4BEG[3] ,
    \Tile_X1Y12_EE4BEG[2] ,
    \Tile_X1Y12_EE4BEG[1] ,
    \Tile_X1Y12_EE4BEG[0] }),
    .FrameData({\Tile_X1Y12_FrameData_O[31] ,
    \Tile_X1Y12_FrameData_O[30] ,
    \Tile_X1Y12_FrameData_O[29] ,
    \Tile_X1Y12_FrameData_O[28] ,
    \Tile_X1Y12_FrameData_O[27] ,
    \Tile_X1Y12_FrameData_O[26] ,
    \Tile_X1Y12_FrameData_O[25] ,
    \Tile_X1Y12_FrameData_O[24] ,
    \Tile_X1Y12_FrameData_O[23] ,
    \Tile_X1Y12_FrameData_O[22] ,
    \Tile_X1Y12_FrameData_O[21] ,
    \Tile_X1Y12_FrameData_O[20] ,
    \Tile_X1Y12_FrameData_O[19] ,
    \Tile_X1Y12_FrameData_O[18] ,
    \Tile_X1Y12_FrameData_O[17] ,
    \Tile_X1Y12_FrameData_O[16] ,
    \Tile_X1Y12_FrameData_O[15] ,
    \Tile_X1Y12_FrameData_O[14] ,
    \Tile_X1Y12_FrameData_O[13] ,
    \Tile_X1Y12_FrameData_O[12] ,
    \Tile_X1Y12_FrameData_O[11] ,
    \Tile_X1Y12_FrameData_O[10] ,
    \Tile_X1Y12_FrameData_O[9] ,
    \Tile_X1Y12_FrameData_O[8] ,
    \Tile_X1Y12_FrameData_O[7] ,
    \Tile_X1Y12_FrameData_O[6] ,
    \Tile_X1Y12_FrameData_O[5] ,
    \Tile_X1Y12_FrameData_O[4] ,
    \Tile_X1Y12_FrameData_O[3] ,
    \Tile_X1Y12_FrameData_O[2] ,
    \Tile_X1Y12_FrameData_O[1] ,
    \Tile_X1Y12_FrameData_O[0] }),
    .FrameData_O({\Tile_X2Y12_FrameData_O[31] ,
    \Tile_X2Y12_FrameData_O[30] ,
    \Tile_X2Y12_FrameData_O[29] ,
    \Tile_X2Y12_FrameData_O[28] ,
    \Tile_X2Y12_FrameData_O[27] ,
    \Tile_X2Y12_FrameData_O[26] ,
    \Tile_X2Y12_FrameData_O[25] ,
    \Tile_X2Y12_FrameData_O[24] ,
    \Tile_X2Y12_FrameData_O[23] ,
    \Tile_X2Y12_FrameData_O[22] ,
    \Tile_X2Y12_FrameData_O[21] ,
    \Tile_X2Y12_FrameData_O[20] ,
    \Tile_X2Y12_FrameData_O[19] ,
    \Tile_X2Y12_FrameData_O[18] ,
    \Tile_X2Y12_FrameData_O[17] ,
    \Tile_X2Y12_FrameData_O[16] ,
    \Tile_X2Y12_FrameData_O[15] ,
    \Tile_X2Y12_FrameData_O[14] ,
    \Tile_X2Y12_FrameData_O[13] ,
    \Tile_X2Y12_FrameData_O[12] ,
    \Tile_X2Y12_FrameData_O[11] ,
    \Tile_X2Y12_FrameData_O[10] ,
    \Tile_X2Y12_FrameData_O[9] ,
    \Tile_X2Y12_FrameData_O[8] ,
    \Tile_X2Y12_FrameData_O[7] ,
    \Tile_X2Y12_FrameData_O[6] ,
    \Tile_X2Y12_FrameData_O[5] ,
    \Tile_X2Y12_FrameData_O[4] ,
    \Tile_X2Y12_FrameData_O[3] ,
    \Tile_X2Y12_FrameData_O[2] ,
    \Tile_X2Y12_FrameData_O[1] ,
    \Tile_X2Y12_FrameData_O[0] }),
    .FrameStrobe({\Tile_X2Y13_FrameStrobe_O[19] ,
    \Tile_X2Y13_FrameStrobe_O[18] ,
    \Tile_X2Y13_FrameStrobe_O[17] ,
    \Tile_X2Y13_FrameStrobe_O[16] ,
    \Tile_X2Y13_FrameStrobe_O[15] ,
    \Tile_X2Y13_FrameStrobe_O[14] ,
    \Tile_X2Y13_FrameStrobe_O[13] ,
    \Tile_X2Y13_FrameStrobe_O[12] ,
    \Tile_X2Y13_FrameStrobe_O[11] ,
    \Tile_X2Y13_FrameStrobe_O[10] ,
    \Tile_X2Y13_FrameStrobe_O[9] ,
    \Tile_X2Y13_FrameStrobe_O[8] ,
    \Tile_X2Y13_FrameStrobe_O[7] ,
    \Tile_X2Y13_FrameStrobe_O[6] ,
    \Tile_X2Y13_FrameStrobe_O[5] ,
    \Tile_X2Y13_FrameStrobe_O[4] ,
    \Tile_X2Y13_FrameStrobe_O[3] ,
    \Tile_X2Y13_FrameStrobe_O[2] ,
    \Tile_X2Y13_FrameStrobe_O[1] ,
    \Tile_X2Y13_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X2Y12_FrameStrobe_O[19] ,
    \Tile_X2Y12_FrameStrobe_O[18] ,
    \Tile_X2Y12_FrameStrobe_O[17] ,
    \Tile_X2Y12_FrameStrobe_O[16] ,
    \Tile_X2Y12_FrameStrobe_O[15] ,
    \Tile_X2Y12_FrameStrobe_O[14] ,
    \Tile_X2Y12_FrameStrobe_O[13] ,
    \Tile_X2Y12_FrameStrobe_O[12] ,
    \Tile_X2Y12_FrameStrobe_O[11] ,
    \Tile_X2Y12_FrameStrobe_O[10] ,
    \Tile_X2Y12_FrameStrobe_O[9] ,
    \Tile_X2Y12_FrameStrobe_O[8] ,
    \Tile_X2Y12_FrameStrobe_O[7] ,
    \Tile_X2Y12_FrameStrobe_O[6] ,
    \Tile_X2Y12_FrameStrobe_O[5] ,
    \Tile_X2Y12_FrameStrobe_O[4] ,
    \Tile_X2Y12_FrameStrobe_O[3] ,
    \Tile_X2Y12_FrameStrobe_O[2] ,
    \Tile_X2Y12_FrameStrobe_O[1] ,
    \Tile_X2Y12_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X2Y12_N1BEG[3] ,
    \Tile_X2Y12_N1BEG[2] ,
    \Tile_X2Y12_N1BEG[1] ,
    \Tile_X2Y12_N1BEG[0] }),
    .N1END({\Tile_X2Y13_N1BEG[3] ,
    \Tile_X2Y13_N1BEG[2] ,
    \Tile_X2Y13_N1BEG[1] ,
    \Tile_X2Y13_N1BEG[0] }),
    .N2BEG({\Tile_X2Y12_N2BEG[7] ,
    \Tile_X2Y12_N2BEG[6] ,
    \Tile_X2Y12_N2BEG[5] ,
    \Tile_X2Y12_N2BEG[4] ,
    \Tile_X2Y12_N2BEG[3] ,
    \Tile_X2Y12_N2BEG[2] ,
    \Tile_X2Y12_N2BEG[1] ,
    \Tile_X2Y12_N2BEG[0] }),
    .N2BEGb({\Tile_X2Y12_N2BEGb[7] ,
    \Tile_X2Y12_N2BEGb[6] ,
    \Tile_X2Y12_N2BEGb[5] ,
    \Tile_X2Y12_N2BEGb[4] ,
    \Tile_X2Y12_N2BEGb[3] ,
    \Tile_X2Y12_N2BEGb[2] ,
    \Tile_X2Y12_N2BEGb[1] ,
    \Tile_X2Y12_N2BEGb[0] }),
    .N2END({\Tile_X2Y13_N2BEGb[7] ,
    \Tile_X2Y13_N2BEGb[6] ,
    \Tile_X2Y13_N2BEGb[5] ,
    \Tile_X2Y13_N2BEGb[4] ,
    \Tile_X2Y13_N2BEGb[3] ,
    \Tile_X2Y13_N2BEGb[2] ,
    \Tile_X2Y13_N2BEGb[1] ,
    \Tile_X2Y13_N2BEGb[0] }),
    .N2MID({\Tile_X2Y13_N2BEG[7] ,
    \Tile_X2Y13_N2BEG[6] ,
    \Tile_X2Y13_N2BEG[5] ,
    \Tile_X2Y13_N2BEG[4] ,
    \Tile_X2Y13_N2BEG[3] ,
    \Tile_X2Y13_N2BEG[2] ,
    \Tile_X2Y13_N2BEG[1] ,
    \Tile_X2Y13_N2BEG[0] }),
    .N4BEG({\Tile_X2Y12_N4BEG[15] ,
    \Tile_X2Y12_N4BEG[14] ,
    \Tile_X2Y12_N4BEG[13] ,
    \Tile_X2Y12_N4BEG[12] ,
    \Tile_X2Y12_N4BEG[11] ,
    \Tile_X2Y12_N4BEG[10] ,
    \Tile_X2Y12_N4BEG[9] ,
    \Tile_X2Y12_N4BEG[8] ,
    \Tile_X2Y12_N4BEG[7] ,
    \Tile_X2Y12_N4BEG[6] ,
    \Tile_X2Y12_N4BEG[5] ,
    \Tile_X2Y12_N4BEG[4] ,
    \Tile_X2Y12_N4BEG[3] ,
    \Tile_X2Y12_N4BEG[2] ,
    \Tile_X2Y12_N4BEG[1] ,
    \Tile_X2Y12_N4BEG[0] }),
    .N4END({\Tile_X2Y13_N4BEG[15] ,
    \Tile_X2Y13_N4BEG[14] ,
    \Tile_X2Y13_N4BEG[13] ,
    \Tile_X2Y13_N4BEG[12] ,
    \Tile_X2Y13_N4BEG[11] ,
    \Tile_X2Y13_N4BEG[10] ,
    \Tile_X2Y13_N4BEG[9] ,
    \Tile_X2Y13_N4BEG[8] ,
    \Tile_X2Y13_N4BEG[7] ,
    \Tile_X2Y13_N4BEG[6] ,
    \Tile_X2Y13_N4BEG[5] ,
    \Tile_X2Y13_N4BEG[4] ,
    \Tile_X2Y13_N4BEG[3] ,
    \Tile_X2Y13_N4BEG[2] ,
    \Tile_X2Y13_N4BEG[1] ,
    \Tile_X2Y13_N4BEG[0] }),
    .NN4BEG({\Tile_X2Y12_NN4BEG[15] ,
    \Tile_X2Y12_NN4BEG[14] ,
    \Tile_X2Y12_NN4BEG[13] ,
    \Tile_X2Y12_NN4BEG[12] ,
    \Tile_X2Y12_NN4BEG[11] ,
    \Tile_X2Y12_NN4BEG[10] ,
    \Tile_X2Y12_NN4BEG[9] ,
    \Tile_X2Y12_NN4BEG[8] ,
    \Tile_X2Y12_NN4BEG[7] ,
    \Tile_X2Y12_NN4BEG[6] ,
    \Tile_X2Y12_NN4BEG[5] ,
    \Tile_X2Y12_NN4BEG[4] ,
    \Tile_X2Y12_NN4BEG[3] ,
    \Tile_X2Y12_NN4BEG[2] ,
    \Tile_X2Y12_NN4BEG[1] ,
    \Tile_X2Y12_NN4BEG[0] }),
    .NN4END({\Tile_X2Y13_NN4BEG[15] ,
    \Tile_X2Y13_NN4BEG[14] ,
    \Tile_X2Y13_NN4BEG[13] ,
    \Tile_X2Y13_NN4BEG[12] ,
    \Tile_X2Y13_NN4BEG[11] ,
    \Tile_X2Y13_NN4BEG[10] ,
    \Tile_X2Y13_NN4BEG[9] ,
    \Tile_X2Y13_NN4BEG[8] ,
    \Tile_X2Y13_NN4BEG[7] ,
    \Tile_X2Y13_NN4BEG[6] ,
    \Tile_X2Y13_NN4BEG[5] ,
    \Tile_X2Y13_NN4BEG[4] ,
    \Tile_X2Y13_NN4BEG[3] ,
    \Tile_X2Y13_NN4BEG[2] ,
    \Tile_X2Y13_NN4BEG[1] ,
    \Tile_X2Y13_NN4BEG[0] }),
    .S1BEG({\Tile_X2Y12_S1BEG[3] ,
    \Tile_X2Y12_S1BEG[2] ,
    \Tile_X2Y12_S1BEG[1] ,
    \Tile_X2Y12_S1BEG[0] }),
    .S1END({\Tile_X2Y11_S1BEG[3] ,
    \Tile_X2Y11_S1BEG[2] ,
    \Tile_X2Y11_S1BEG[1] ,
    \Tile_X2Y11_S1BEG[0] }),
    .S2BEG({\Tile_X2Y12_S2BEG[7] ,
    \Tile_X2Y12_S2BEG[6] ,
    \Tile_X2Y12_S2BEG[5] ,
    \Tile_X2Y12_S2BEG[4] ,
    \Tile_X2Y12_S2BEG[3] ,
    \Tile_X2Y12_S2BEG[2] ,
    \Tile_X2Y12_S2BEG[1] ,
    \Tile_X2Y12_S2BEG[0] }),
    .S2BEGb({\Tile_X2Y12_S2BEGb[7] ,
    \Tile_X2Y12_S2BEGb[6] ,
    \Tile_X2Y12_S2BEGb[5] ,
    \Tile_X2Y12_S2BEGb[4] ,
    \Tile_X2Y12_S2BEGb[3] ,
    \Tile_X2Y12_S2BEGb[2] ,
    \Tile_X2Y12_S2BEGb[1] ,
    \Tile_X2Y12_S2BEGb[0] }),
    .S2END({\Tile_X2Y11_S2BEGb[7] ,
    \Tile_X2Y11_S2BEGb[6] ,
    \Tile_X2Y11_S2BEGb[5] ,
    \Tile_X2Y11_S2BEGb[4] ,
    \Tile_X2Y11_S2BEGb[3] ,
    \Tile_X2Y11_S2BEGb[2] ,
    \Tile_X2Y11_S2BEGb[1] ,
    \Tile_X2Y11_S2BEGb[0] }),
    .S2MID({\Tile_X2Y11_S2BEG[7] ,
    \Tile_X2Y11_S2BEG[6] ,
    \Tile_X2Y11_S2BEG[5] ,
    \Tile_X2Y11_S2BEG[4] ,
    \Tile_X2Y11_S2BEG[3] ,
    \Tile_X2Y11_S2BEG[2] ,
    \Tile_X2Y11_S2BEG[1] ,
    \Tile_X2Y11_S2BEG[0] }),
    .S4BEG({\Tile_X2Y12_S4BEG[15] ,
    \Tile_X2Y12_S4BEG[14] ,
    \Tile_X2Y12_S4BEG[13] ,
    \Tile_X2Y12_S4BEG[12] ,
    \Tile_X2Y12_S4BEG[11] ,
    \Tile_X2Y12_S4BEG[10] ,
    \Tile_X2Y12_S4BEG[9] ,
    \Tile_X2Y12_S4BEG[8] ,
    \Tile_X2Y12_S4BEG[7] ,
    \Tile_X2Y12_S4BEG[6] ,
    \Tile_X2Y12_S4BEG[5] ,
    \Tile_X2Y12_S4BEG[4] ,
    \Tile_X2Y12_S4BEG[3] ,
    \Tile_X2Y12_S4BEG[2] ,
    \Tile_X2Y12_S4BEG[1] ,
    \Tile_X2Y12_S4BEG[0] }),
    .S4END({\Tile_X2Y11_S4BEG[15] ,
    \Tile_X2Y11_S4BEG[14] ,
    \Tile_X2Y11_S4BEG[13] ,
    \Tile_X2Y11_S4BEG[12] ,
    \Tile_X2Y11_S4BEG[11] ,
    \Tile_X2Y11_S4BEG[10] ,
    \Tile_X2Y11_S4BEG[9] ,
    \Tile_X2Y11_S4BEG[8] ,
    \Tile_X2Y11_S4BEG[7] ,
    \Tile_X2Y11_S4BEG[6] ,
    \Tile_X2Y11_S4BEG[5] ,
    \Tile_X2Y11_S4BEG[4] ,
    \Tile_X2Y11_S4BEG[3] ,
    \Tile_X2Y11_S4BEG[2] ,
    \Tile_X2Y11_S4BEG[1] ,
    \Tile_X2Y11_S4BEG[0] }),
    .SS4BEG({\Tile_X2Y12_SS4BEG[15] ,
    \Tile_X2Y12_SS4BEG[14] ,
    \Tile_X2Y12_SS4BEG[13] ,
    \Tile_X2Y12_SS4BEG[12] ,
    \Tile_X2Y12_SS4BEG[11] ,
    \Tile_X2Y12_SS4BEG[10] ,
    \Tile_X2Y12_SS4BEG[9] ,
    \Tile_X2Y12_SS4BEG[8] ,
    \Tile_X2Y12_SS4BEG[7] ,
    \Tile_X2Y12_SS4BEG[6] ,
    \Tile_X2Y12_SS4BEG[5] ,
    \Tile_X2Y12_SS4BEG[4] ,
    \Tile_X2Y12_SS4BEG[3] ,
    \Tile_X2Y12_SS4BEG[2] ,
    \Tile_X2Y12_SS4BEG[1] ,
    \Tile_X2Y12_SS4BEG[0] }),
    .SS4END({\Tile_X2Y11_SS4BEG[15] ,
    \Tile_X2Y11_SS4BEG[14] ,
    \Tile_X2Y11_SS4BEG[13] ,
    \Tile_X2Y11_SS4BEG[12] ,
    \Tile_X2Y11_SS4BEG[11] ,
    \Tile_X2Y11_SS4BEG[10] ,
    \Tile_X2Y11_SS4BEG[9] ,
    \Tile_X2Y11_SS4BEG[8] ,
    \Tile_X2Y11_SS4BEG[7] ,
    \Tile_X2Y11_SS4BEG[6] ,
    \Tile_X2Y11_SS4BEG[5] ,
    \Tile_X2Y11_SS4BEG[4] ,
    \Tile_X2Y11_SS4BEG[3] ,
    \Tile_X2Y11_SS4BEG[2] ,
    \Tile_X2Y11_SS4BEG[1] ,
    \Tile_X2Y11_SS4BEG[0] }),
    .W1BEG({\Tile_X2Y12_W1BEG[3] ,
    \Tile_X2Y12_W1BEG[2] ,
    \Tile_X2Y12_W1BEG[1] ,
    \Tile_X2Y12_W1BEG[0] }),
    .W1END({\Tile_X3Y12_W1BEG[3] ,
    \Tile_X3Y12_W1BEG[2] ,
    \Tile_X3Y12_W1BEG[1] ,
    \Tile_X3Y12_W1BEG[0] }),
    .W2BEG({\Tile_X2Y12_W2BEG[7] ,
    \Tile_X2Y12_W2BEG[6] ,
    \Tile_X2Y12_W2BEG[5] ,
    \Tile_X2Y12_W2BEG[4] ,
    \Tile_X2Y12_W2BEG[3] ,
    \Tile_X2Y12_W2BEG[2] ,
    \Tile_X2Y12_W2BEG[1] ,
    \Tile_X2Y12_W2BEG[0] }),
    .W2BEGb({\Tile_X2Y12_W2BEGb[7] ,
    \Tile_X2Y12_W2BEGb[6] ,
    \Tile_X2Y12_W2BEGb[5] ,
    \Tile_X2Y12_W2BEGb[4] ,
    \Tile_X2Y12_W2BEGb[3] ,
    \Tile_X2Y12_W2BEGb[2] ,
    \Tile_X2Y12_W2BEGb[1] ,
    \Tile_X2Y12_W2BEGb[0] }),
    .W2END({\Tile_X3Y12_W2BEGb[7] ,
    \Tile_X3Y12_W2BEGb[6] ,
    \Tile_X3Y12_W2BEGb[5] ,
    \Tile_X3Y12_W2BEGb[4] ,
    \Tile_X3Y12_W2BEGb[3] ,
    \Tile_X3Y12_W2BEGb[2] ,
    \Tile_X3Y12_W2BEGb[1] ,
    \Tile_X3Y12_W2BEGb[0] }),
    .W2MID({\Tile_X3Y12_W2BEG[7] ,
    \Tile_X3Y12_W2BEG[6] ,
    \Tile_X3Y12_W2BEG[5] ,
    \Tile_X3Y12_W2BEG[4] ,
    \Tile_X3Y12_W2BEG[3] ,
    \Tile_X3Y12_W2BEG[2] ,
    \Tile_X3Y12_W2BEG[1] ,
    \Tile_X3Y12_W2BEG[0] }),
    .W6BEG({\Tile_X2Y12_W6BEG[11] ,
    \Tile_X2Y12_W6BEG[10] ,
    \Tile_X2Y12_W6BEG[9] ,
    \Tile_X2Y12_W6BEG[8] ,
    \Tile_X2Y12_W6BEG[7] ,
    \Tile_X2Y12_W6BEG[6] ,
    \Tile_X2Y12_W6BEG[5] ,
    \Tile_X2Y12_W6BEG[4] ,
    \Tile_X2Y12_W6BEG[3] ,
    \Tile_X2Y12_W6BEG[2] ,
    \Tile_X2Y12_W6BEG[1] ,
    \Tile_X2Y12_W6BEG[0] }),
    .W6END({\Tile_X3Y12_W6BEG[11] ,
    \Tile_X3Y12_W6BEG[10] ,
    \Tile_X3Y12_W6BEG[9] ,
    \Tile_X3Y12_W6BEG[8] ,
    \Tile_X3Y12_W6BEG[7] ,
    \Tile_X3Y12_W6BEG[6] ,
    \Tile_X3Y12_W6BEG[5] ,
    \Tile_X3Y12_W6BEG[4] ,
    \Tile_X3Y12_W6BEG[3] ,
    \Tile_X3Y12_W6BEG[2] ,
    \Tile_X3Y12_W6BEG[1] ,
    \Tile_X3Y12_W6BEG[0] }),
    .WW4BEG({\Tile_X2Y12_WW4BEG[15] ,
    \Tile_X2Y12_WW4BEG[14] ,
    \Tile_X2Y12_WW4BEG[13] ,
    \Tile_X2Y12_WW4BEG[12] ,
    \Tile_X2Y12_WW4BEG[11] ,
    \Tile_X2Y12_WW4BEG[10] ,
    \Tile_X2Y12_WW4BEG[9] ,
    \Tile_X2Y12_WW4BEG[8] ,
    \Tile_X2Y12_WW4BEG[7] ,
    \Tile_X2Y12_WW4BEG[6] ,
    \Tile_X2Y12_WW4BEG[5] ,
    \Tile_X2Y12_WW4BEG[4] ,
    \Tile_X2Y12_WW4BEG[3] ,
    \Tile_X2Y12_WW4BEG[2] ,
    \Tile_X2Y12_WW4BEG[1] ,
    \Tile_X2Y12_WW4BEG[0] }),
    .WW4END({\Tile_X3Y12_WW4BEG[15] ,
    \Tile_X3Y12_WW4BEG[14] ,
    \Tile_X3Y12_WW4BEG[13] ,
    \Tile_X3Y12_WW4BEG[12] ,
    \Tile_X3Y12_WW4BEG[11] ,
    \Tile_X3Y12_WW4BEG[10] ,
    \Tile_X3Y12_WW4BEG[9] ,
    \Tile_X3Y12_WW4BEG[8] ,
    \Tile_X3Y12_WW4BEG[7] ,
    \Tile_X3Y12_WW4BEG[6] ,
    \Tile_X3Y12_WW4BEG[5] ,
    \Tile_X3Y12_WW4BEG[4] ,
    \Tile_X3Y12_WW4BEG[3] ,
    \Tile_X3Y12_WW4BEG[2] ,
    \Tile_X3Y12_WW4BEG[1] ,
    \Tile_X3Y12_WW4BEG[0] }));
 LUT4AB Tile_X2Y13_LUT4AB (.Ci(Tile_X2Y14_Co),
    .Co(Tile_X2Y13_Co),
    .UserCLK(Tile_X2Y14_UserCLKo),
    .UserCLKo(Tile_X2Y13_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X2Y13_E1BEG[3] ,
    \Tile_X2Y13_E1BEG[2] ,
    \Tile_X2Y13_E1BEG[1] ,
    \Tile_X2Y13_E1BEG[0] }),
    .E1END({\Tile_X1Y13_E1BEG[3] ,
    \Tile_X1Y13_E1BEG[2] ,
    \Tile_X1Y13_E1BEG[1] ,
    \Tile_X1Y13_E1BEG[0] }),
    .E2BEG({\Tile_X2Y13_E2BEG[7] ,
    \Tile_X2Y13_E2BEG[6] ,
    \Tile_X2Y13_E2BEG[5] ,
    \Tile_X2Y13_E2BEG[4] ,
    \Tile_X2Y13_E2BEG[3] ,
    \Tile_X2Y13_E2BEG[2] ,
    \Tile_X2Y13_E2BEG[1] ,
    \Tile_X2Y13_E2BEG[0] }),
    .E2BEGb({\Tile_X2Y13_E2BEGb[7] ,
    \Tile_X2Y13_E2BEGb[6] ,
    \Tile_X2Y13_E2BEGb[5] ,
    \Tile_X2Y13_E2BEGb[4] ,
    \Tile_X2Y13_E2BEGb[3] ,
    \Tile_X2Y13_E2BEGb[2] ,
    \Tile_X2Y13_E2BEGb[1] ,
    \Tile_X2Y13_E2BEGb[0] }),
    .E2END({\Tile_X1Y13_E2BEGb[7] ,
    \Tile_X1Y13_E2BEGb[6] ,
    \Tile_X1Y13_E2BEGb[5] ,
    \Tile_X1Y13_E2BEGb[4] ,
    \Tile_X1Y13_E2BEGb[3] ,
    \Tile_X1Y13_E2BEGb[2] ,
    \Tile_X1Y13_E2BEGb[1] ,
    \Tile_X1Y13_E2BEGb[0] }),
    .E2MID({\Tile_X1Y13_E2BEG[7] ,
    \Tile_X1Y13_E2BEG[6] ,
    \Tile_X1Y13_E2BEG[5] ,
    \Tile_X1Y13_E2BEG[4] ,
    \Tile_X1Y13_E2BEG[3] ,
    \Tile_X1Y13_E2BEG[2] ,
    \Tile_X1Y13_E2BEG[1] ,
    \Tile_X1Y13_E2BEG[0] }),
    .E6BEG({\Tile_X2Y13_E6BEG[11] ,
    \Tile_X2Y13_E6BEG[10] ,
    \Tile_X2Y13_E6BEG[9] ,
    \Tile_X2Y13_E6BEG[8] ,
    \Tile_X2Y13_E6BEG[7] ,
    \Tile_X2Y13_E6BEG[6] ,
    \Tile_X2Y13_E6BEG[5] ,
    \Tile_X2Y13_E6BEG[4] ,
    \Tile_X2Y13_E6BEG[3] ,
    \Tile_X2Y13_E6BEG[2] ,
    \Tile_X2Y13_E6BEG[1] ,
    \Tile_X2Y13_E6BEG[0] }),
    .E6END({\Tile_X1Y13_E6BEG[11] ,
    \Tile_X1Y13_E6BEG[10] ,
    \Tile_X1Y13_E6BEG[9] ,
    \Tile_X1Y13_E6BEG[8] ,
    \Tile_X1Y13_E6BEG[7] ,
    \Tile_X1Y13_E6BEG[6] ,
    \Tile_X1Y13_E6BEG[5] ,
    \Tile_X1Y13_E6BEG[4] ,
    \Tile_X1Y13_E6BEG[3] ,
    \Tile_X1Y13_E6BEG[2] ,
    \Tile_X1Y13_E6BEG[1] ,
    \Tile_X1Y13_E6BEG[0] }),
    .EE4BEG({\Tile_X2Y13_EE4BEG[15] ,
    \Tile_X2Y13_EE4BEG[14] ,
    \Tile_X2Y13_EE4BEG[13] ,
    \Tile_X2Y13_EE4BEG[12] ,
    \Tile_X2Y13_EE4BEG[11] ,
    \Tile_X2Y13_EE4BEG[10] ,
    \Tile_X2Y13_EE4BEG[9] ,
    \Tile_X2Y13_EE4BEG[8] ,
    \Tile_X2Y13_EE4BEG[7] ,
    \Tile_X2Y13_EE4BEG[6] ,
    \Tile_X2Y13_EE4BEG[5] ,
    \Tile_X2Y13_EE4BEG[4] ,
    \Tile_X2Y13_EE4BEG[3] ,
    \Tile_X2Y13_EE4BEG[2] ,
    \Tile_X2Y13_EE4BEG[1] ,
    \Tile_X2Y13_EE4BEG[0] }),
    .EE4END({\Tile_X1Y13_EE4BEG[15] ,
    \Tile_X1Y13_EE4BEG[14] ,
    \Tile_X1Y13_EE4BEG[13] ,
    \Tile_X1Y13_EE4BEG[12] ,
    \Tile_X1Y13_EE4BEG[11] ,
    \Tile_X1Y13_EE4BEG[10] ,
    \Tile_X1Y13_EE4BEG[9] ,
    \Tile_X1Y13_EE4BEG[8] ,
    \Tile_X1Y13_EE4BEG[7] ,
    \Tile_X1Y13_EE4BEG[6] ,
    \Tile_X1Y13_EE4BEG[5] ,
    \Tile_X1Y13_EE4BEG[4] ,
    \Tile_X1Y13_EE4BEG[3] ,
    \Tile_X1Y13_EE4BEG[2] ,
    \Tile_X1Y13_EE4BEG[1] ,
    \Tile_X1Y13_EE4BEG[0] }),
    .FrameData({\Tile_X1Y13_FrameData_O[31] ,
    \Tile_X1Y13_FrameData_O[30] ,
    \Tile_X1Y13_FrameData_O[29] ,
    \Tile_X1Y13_FrameData_O[28] ,
    \Tile_X1Y13_FrameData_O[27] ,
    \Tile_X1Y13_FrameData_O[26] ,
    \Tile_X1Y13_FrameData_O[25] ,
    \Tile_X1Y13_FrameData_O[24] ,
    \Tile_X1Y13_FrameData_O[23] ,
    \Tile_X1Y13_FrameData_O[22] ,
    \Tile_X1Y13_FrameData_O[21] ,
    \Tile_X1Y13_FrameData_O[20] ,
    \Tile_X1Y13_FrameData_O[19] ,
    \Tile_X1Y13_FrameData_O[18] ,
    \Tile_X1Y13_FrameData_O[17] ,
    \Tile_X1Y13_FrameData_O[16] ,
    \Tile_X1Y13_FrameData_O[15] ,
    \Tile_X1Y13_FrameData_O[14] ,
    \Tile_X1Y13_FrameData_O[13] ,
    \Tile_X1Y13_FrameData_O[12] ,
    \Tile_X1Y13_FrameData_O[11] ,
    \Tile_X1Y13_FrameData_O[10] ,
    \Tile_X1Y13_FrameData_O[9] ,
    \Tile_X1Y13_FrameData_O[8] ,
    \Tile_X1Y13_FrameData_O[7] ,
    \Tile_X1Y13_FrameData_O[6] ,
    \Tile_X1Y13_FrameData_O[5] ,
    \Tile_X1Y13_FrameData_O[4] ,
    \Tile_X1Y13_FrameData_O[3] ,
    \Tile_X1Y13_FrameData_O[2] ,
    \Tile_X1Y13_FrameData_O[1] ,
    \Tile_X1Y13_FrameData_O[0] }),
    .FrameData_O({\Tile_X2Y13_FrameData_O[31] ,
    \Tile_X2Y13_FrameData_O[30] ,
    \Tile_X2Y13_FrameData_O[29] ,
    \Tile_X2Y13_FrameData_O[28] ,
    \Tile_X2Y13_FrameData_O[27] ,
    \Tile_X2Y13_FrameData_O[26] ,
    \Tile_X2Y13_FrameData_O[25] ,
    \Tile_X2Y13_FrameData_O[24] ,
    \Tile_X2Y13_FrameData_O[23] ,
    \Tile_X2Y13_FrameData_O[22] ,
    \Tile_X2Y13_FrameData_O[21] ,
    \Tile_X2Y13_FrameData_O[20] ,
    \Tile_X2Y13_FrameData_O[19] ,
    \Tile_X2Y13_FrameData_O[18] ,
    \Tile_X2Y13_FrameData_O[17] ,
    \Tile_X2Y13_FrameData_O[16] ,
    \Tile_X2Y13_FrameData_O[15] ,
    \Tile_X2Y13_FrameData_O[14] ,
    \Tile_X2Y13_FrameData_O[13] ,
    \Tile_X2Y13_FrameData_O[12] ,
    \Tile_X2Y13_FrameData_O[11] ,
    \Tile_X2Y13_FrameData_O[10] ,
    \Tile_X2Y13_FrameData_O[9] ,
    \Tile_X2Y13_FrameData_O[8] ,
    \Tile_X2Y13_FrameData_O[7] ,
    \Tile_X2Y13_FrameData_O[6] ,
    \Tile_X2Y13_FrameData_O[5] ,
    \Tile_X2Y13_FrameData_O[4] ,
    \Tile_X2Y13_FrameData_O[3] ,
    \Tile_X2Y13_FrameData_O[2] ,
    \Tile_X2Y13_FrameData_O[1] ,
    \Tile_X2Y13_FrameData_O[0] }),
    .FrameStrobe({\Tile_X2Y14_FrameStrobe_O[19] ,
    \Tile_X2Y14_FrameStrobe_O[18] ,
    \Tile_X2Y14_FrameStrobe_O[17] ,
    \Tile_X2Y14_FrameStrobe_O[16] ,
    \Tile_X2Y14_FrameStrobe_O[15] ,
    \Tile_X2Y14_FrameStrobe_O[14] ,
    \Tile_X2Y14_FrameStrobe_O[13] ,
    \Tile_X2Y14_FrameStrobe_O[12] ,
    \Tile_X2Y14_FrameStrobe_O[11] ,
    \Tile_X2Y14_FrameStrobe_O[10] ,
    \Tile_X2Y14_FrameStrobe_O[9] ,
    \Tile_X2Y14_FrameStrobe_O[8] ,
    \Tile_X2Y14_FrameStrobe_O[7] ,
    \Tile_X2Y14_FrameStrobe_O[6] ,
    \Tile_X2Y14_FrameStrobe_O[5] ,
    \Tile_X2Y14_FrameStrobe_O[4] ,
    \Tile_X2Y14_FrameStrobe_O[3] ,
    \Tile_X2Y14_FrameStrobe_O[2] ,
    \Tile_X2Y14_FrameStrobe_O[1] ,
    \Tile_X2Y14_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X2Y13_FrameStrobe_O[19] ,
    \Tile_X2Y13_FrameStrobe_O[18] ,
    \Tile_X2Y13_FrameStrobe_O[17] ,
    \Tile_X2Y13_FrameStrobe_O[16] ,
    \Tile_X2Y13_FrameStrobe_O[15] ,
    \Tile_X2Y13_FrameStrobe_O[14] ,
    \Tile_X2Y13_FrameStrobe_O[13] ,
    \Tile_X2Y13_FrameStrobe_O[12] ,
    \Tile_X2Y13_FrameStrobe_O[11] ,
    \Tile_X2Y13_FrameStrobe_O[10] ,
    \Tile_X2Y13_FrameStrobe_O[9] ,
    \Tile_X2Y13_FrameStrobe_O[8] ,
    \Tile_X2Y13_FrameStrobe_O[7] ,
    \Tile_X2Y13_FrameStrobe_O[6] ,
    \Tile_X2Y13_FrameStrobe_O[5] ,
    \Tile_X2Y13_FrameStrobe_O[4] ,
    \Tile_X2Y13_FrameStrobe_O[3] ,
    \Tile_X2Y13_FrameStrobe_O[2] ,
    \Tile_X2Y13_FrameStrobe_O[1] ,
    \Tile_X2Y13_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X2Y13_N1BEG[3] ,
    \Tile_X2Y13_N1BEG[2] ,
    \Tile_X2Y13_N1BEG[1] ,
    \Tile_X2Y13_N1BEG[0] }),
    .N1END({\Tile_X2Y14_N1BEG[3] ,
    \Tile_X2Y14_N1BEG[2] ,
    \Tile_X2Y14_N1BEG[1] ,
    \Tile_X2Y14_N1BEG[0] }),
    .N2BEG({\Tile_X2Y13_N2BEG[7] ,
    \Tile_X2Y13_N2BEG[6] ,
    \Tile_X2Y13_N2BEG[5] ,
    \Tile_X2Y13_N2BEG[4] ,
    \Tile_X2Y13_N2BEG[3] ,
    \Tile_X2Y13_N2BEG[2] ,
    \Tile_X2Y13_N2BEG[1] ,
    \Tile_X2Y13_N2BEG[0] }),
    .N2BEGb({\Tile_X2Y13_N2BEGb[7] ,
    \Tile_X2Y13_N2BEGb[6] ,
    \Tile_X2Y13_N2BEGb[5] ,
    \Tile_X2Y13_N2BEGb[4] ,
    \Tile_X2Y13_N2BEGb[3] ,
    \Tile_X2Y13_N2BEGb[2] ,
    \Tile_X2Y13_N2BEGb[1] ,
    \Tile_X2Y13_N2BEGb[0] }),
    .N2END({\Tile_X2Y14_N2BEGb[7] ,
    \Tile_X2Y14_N2BEGb[6] ,
    \Tile_X2Y14_N2BEGb[5] ,
    \Tile_X2Y14_N2BEGb[4] ,
    \Tile_X2Y14_N2BEGb[3] ,
    \Tile_X2Y14_N2BEGb[2] ,
    \Tile_X2Y14_N2BEGb[1] ,
    \Tile_X2Y14_N2BEGb[0] }),
    .N2MID({\Tile_X2Y14_N2BEG[7] ,
    \Tile_X2Y14_N2BEG[6] ,
    \Tile_X2Y14_N2BEG[5] ,
    \Tile_X2Y14_N2BEG[4] ,
    \Tile_X2Y14_N2BEG[3] ,
    \Tile_X2Y14_N2BEG[2] ,
    \Tile_X2Y14_N2BEG[1] ,
    \Tile_X2Y14_N2BEG[0] }),
    .N4BEG({\Tile_X2Y13_N4BEG[15] ,
    \Tile_X2Y13_N4BEG[14] ,
    \Tile_X2Y13_N4BEG[13] ,
    \Tile_X2Y13_N4BEG[12] ,
    \Tile_X2Y13_N4BEG[11] ,
    \Tile_X2Y13_N4BEG[10] ,
    \Tile_X2Y13_N4BEG[9] ,
    \Tile_X2Y13_N4BEG[8] ,
    \Tile_X2Y13_N4BEG[7] ,
    \Tile_X2Y13_N4BEG[6] ,
    \Tile_X2Y13_N4BEG[5] ,
    \Tile_X2Y13_N4BEG[4] ,
    \Tile_X2Y13_N4BEG[3] ,
    \Tile_X2Y13_N4BEG[2] ,
    \Tile_X2Y13_N4BEG[1] ,
    \Tile_X2Y13_N4BEG[0] }),
    .N4END({\Tile_X2Y14_N4BEG[15] ,
    \Tile_X2Y14_N4BEG[14] ,
    \Tile_X2Y14_N4BEG[13] ,
    \Tile_X2Y14_N4BEG[12] ,
    \Tile_X2Y14_N4BEG[11] ,
    \Tile_X2Y14_N4BEG[10] ,
    \Tile_X2Y14_N4BEG[9] ,
    \Tile_X2Y14_N4BEG[8] ,
    \Tile_X2Y14_N4BEG[7] ,
    \Tile_X2Y14_N4BEG[6] ,
    \Tile_X2Y14_N4BEG[5] ,
    \Tile_X2Y14_N4BEG[4] ,
    \Tile_X2Y14_N4BEG[3] ,
    \Tile_X2Y14_N4BEG[2] ,
    \Tile_X2Y14_N4BEG[1] ,
    \Tile_X2Y14_N4BEG[0] }),
    .NN4BEG({\Tile_X2Y13_NN4BEG[15] ,
    \Tile_X2Y13_NN4BEG[14] ,
    \Tile_X2Y13_NN4BEG[13] ,
    \Tile_X2Y13_NN4BEG[12] ,
    \Tile_X2Y13_NN4BEG[11] ,
    \Tile_X2Y13_NN4BEG[10] ,
    \Tile_X2Y13_NN4BEG[9] ,
    \Tile_X2Y13_NN4BEG[8] ,
    \Tile_X2Y13_NN4BEG[7] ,
    \Tile_X2Y13_NN4BEG[6] ,
    \Tile_X2Y13_NN4BEG[5] ,
    \Tile_X2Y13_NN4BEG[4] ,
    \Tile_X2Y13_NN4BEG[3] ,
    \Tile_X2Y13_NN4BEG[2] ,
    \Tile_X2Y13_NN4BEG[1] ,
    \Tile_X2Y13_NN4BEG[0] }),
    .NN4END({\Tile_X2Y14_NN4BEG[15] ,
    \Tile_X2Y14_NN4BEG[14] ,
    \Tile_X2Y14_NN4BEG[13] ,
    \Tile_X2Y14_NN4BEG[12] ,
    \Tile_X2Y14_NN4BEG[11] ,
    \Tile_X2Y14_NN4BEG[10] ,
    \Tile_X2Y14_NN4BEG[9] ,
    \Tile_X2Y14_NN4BEG[8] ,
    \Tile_X2Y14_NN4BEG[7] ,
    \Tile_X2Y14_NN4BEG[6] ,
    \Tile_X2Y14_NN4BEG[5] ,
    \Tile_X2Y14_NN4BEG[4] ,
    \Tile_X2Y14_NN4BEG[3] ,
    \Tile_X2Y14_NN4BEG[2] ,
    \Tile_X2Y14_NN4BEG[1] ,
    \Tile_X2Y14_NN4BEG[0] }),
    .S1BEG({\Tile_X2Y13_S1BEG[3] ,
    \Tile_X2Y13_S1BEG[2] ,
    \Tile_X2Y13_S1BEG[1] ,
    \Tile_X2Y13_S1BEG[0] }),
    .S1END({\Tile_X2Y12_S1BEG[3] ,
    \Tile_X2Y12_S1BEG[2] ,
    \Tile_X2Y12_S1BEG[1] ,
    \Tile_X2Y12_S1BEG[0] }),
    .S2BEG({\Tile_X2Y13_S2BEG[7] ,
    \Tile_X2Y13_S2BEG[6] ,
    \Tile_X2Y13_S2BEG[5] ,
    \Tile_X2Y13_S2BEG[4] ,
    \Tile_X2Y13_S2BEG[3] ,
    \Tile_X2Y13_S2BEG[2] ,
    \Tile_X2Y13_S2BEG[1] ,
    \Tile_X2Y13_S2BEG[0] }),
    .S2BEGb({\Tile_X2Y13_S2BEGb[7] ,
    \Tile_X2Y13_S2BEGb[6] ,
    \Tile_X2Y13_S2BEGb[5] ,
    \Tile_X2Y13_S2BEGb[4] ,
    \Tile_X2Y13_S2BEGb[3] ,
    \Tile_X2Y13_S2BEGb[2] ,
    \Tile_X2Y13_S2BEGb[1] ,
    \Tile_X2Y13_S2BEGb[0] }),
    .S2END({\Tile_X2Y12_S2BEGb[7] ,
    \Tile_X2Y12_S2BEGb[6] ,
    \Tile_X2Y12_S2BEGb[5] ,
    \Tile_X2Y12_S2BEGb[4] ,
    \Tile_X2Y12_S2BEGb[3] ,
    \Tile_X2Y12_S2BEGb[2] ,
    \Tile_X2Y12_S2BEGb[1] ,
    \Tile_X2Y12_S2BEGb[0] }),
    .S2MID({\Tile_X2Y12_S2BEG[7] ,
    \Tile_X2Y12_S2BEG[6] ,
    \Tile_X2Y12_S2BEG[5] ,
    \Tile_X2Y12_S2BEG[4] ,
    \Tile_X2Y12_S2BEG[3] ,
    \Tile_X2Y12_S2BEG[2] ,
    \Tile_X2Y12_S2BEG[1] ,
    \Tile_X2Y12_S2BEG[0] }),
    .S4BEG({\Tile_X2Y13_S4BEG[15] ,
    \Tile_X2Y13_S4BEG[14] ,
    \Tile_X2Y13_S4BEG[13] ,
    \Tile_X2Y13_S4BEG[12] ,
    \Tile_X2Y13_S4BEG[11] ,
    \Tile_X2Y13_S4BEG[10] ,
    \Tile_X2Y13_S4BEG[9] ,
    \Tile_X2Y13_S4BEG[8] ,
    \Tile_X2Y13_S4BEG[7] ,
    \Tile_X2Y13_S4BEG[6] ,
    \Tile_X2Y13_S4BEG[5] ,
    \Tile_X2Y13_S4BEG[4] ,
    \Tile_X2Y13_S4BEG[3] ,
    \Tile_X2Y13_S4BEG[2] ,
    \Tile_X2Y13_S4BEG[1] ,
    \Tile_X2Y13_S4BEG[0] }),
    .S4END({\Tile_X2Y12_S4BEG[15] ,
    \Tile_X2Y12_S4BEG[14] ,
    \Tile_X2Y12_S4BEG[13] ,
    \Tile_X2Y12_S4BEG[12] ,
    \Tile_X2Y12_S4BEG[11] ,
    \Tile_X2Y12_S4BEG[10] ,
    \Tile_X2Y12_S4BEG[9] ,
    \Tile_X2Y12_S4BEG[8] ,
    \Tile_X2Y12_S4BEG[7] ,
    \Tile_X2Y12_S4BEG[6] ,
    \Tile_X2Y12_S4BEG[5] ,
    \Tile_X2Y12_S4BEG[4] ,
    \Tile_X2Y12_S4BEG[3] ,
    \Tile_X2Y12_S4BEG[2] ,
    \Tile_X2Y12_S4BEG[1] ,
    \Tile_X2Y12_S4BEG[0] }),
    .SS4BEG({\Tile_X2Y13_SS4BEG[15] ,
    \Tile_X2Y13_SS4BEG[14] ,
    \Tile_X2Y13_SS4BEG[13] ,
    \Tile_X2Y13_SS4BEG[12] ,
    \Tile_X2Y13_SS4BEG[11] ,
    \Tile_X2Y13_SS4BEG[10] ,
    \Tile_X2Y13_SS4BEG[9] ,
    \Tile_X2Y13_SS4BEG[8] ,
    \Tile_X2Y13_SS4BEG[7] ,
    \Tile_X2Y13_SS4BEG[6] ,
    \Tile_X2Y13_SS4BEG[5] ,
    \Tile_X2Y13_SS4BEG[4] ,
    \Tile_X2Y13_SS4BEG[3] ,
    \Tile_X2Y13_SS4BEG[2] ,
    \Tile_X2Y13_SS4BEG[1] ,
    \Tile_X2Y13_SS4BEG[0] }),
    .SS4END({\Tile_X2Y12_SS4BEG[15] ,
    \Tile_X2Y12_SS4BEG[14] ,
    \Tile_X2Y12_SS4BEG[13] ,
    \Tile_X2Y12_SS4BEG[12] ,
    \Tile_X2Y12_SS4BEG[11] ,
    \Tile_X2Y12_SS4BEG[10] ,
    \Tile_X2Y12_SS4BEG[9] ,
    \Tile_X2Y12_SS4BEG[8] ,
    \Tile_X2Y12_SS4BEG[7] ,
    \Tile_X2Y12_SS4BEG[6] ,
    \Tile_X2Y12_SS4BEG[5] ,
    \Tile_X2Y12_SS4BEG[4] ,
    \Tile_X2Y12_SS4BEG[3] ,
    \Tile_X2Y12_SS4BEG[2] ,
    \Tile_X2Y12_SS4BEG[1] ,
    \Tile_X2Y12_SS4BEG[0] }),
    .W1BEG({\Tile_X2Y13_W1BEG[3] ,
    \Tile_X2Y13_W1BEG[2] ,
    \Tile_X2Y13_W1BEG[1] ,
    \Tile_X2Y13_W1BEG[0] }),
    .W1END({\Tile_X3Y13_W1BEG[3] ,
    \Tile_X3Y13_W1BEG[2] ,
    \Tile_X3Y13_W1BEG[1] ,
    \Tile_X3Y13_W1BEG[0] }),
    .W2BEG({\Tile_X2Y13_W2BEG[7] ,
    \Tile_X2Y13_W2BEG[6] ,
    \Tile_X2Y13_W2BEG[5] ,
    \Tile_X2Y13_W2BEG[4] ,
    \Tile_X2Y13_W2BEG[3] ,
    \Tile_X2Y13_W2BEG[2] ,
    \Tile_X2Y13_W2BEG[1] ,
    \Tile_X2Y13_W2BEG[0] }),
    .W2BEGb({\Tile_X2Y13_W2BEGb[7] ,
    \Tile_X2Y13_W2BEGb[6] ,
    \Tile_X2Y13_W2BEGb[5] ,
    \Tile_X2Y13_W2BEGb[4] ,
    \Tile_X2Y13_W2BEGb[3] ,
    \Tile_X2Y13_W2BEGb[2] ,
    \Tile_X2Y13_W2BEGb[1] ,
    \Tile_X2Y13_W2BEGb[0] }),
    .W2END({\Tile_X3Y13_W2BEGb[7] ,
    \Tile_X3Y13_W2BEGb[6] ,
    \Tile_X3Y13_W2BEGb[5] ,
    \Tile_X3Y13_W2BEGb[4] ,
    \Tile_X3Y13_W2BEGb[3] ,
    \Tile_X3Y13_W2BEGb[2] ,
    \Tile_X3Y13_W2BEGb[1] ,
    \Tile_X3Y13_W2BEGb[0] }),
    .W2MID({\Tile_X3Y13_W2BEG[7] ,
    \Tile_X3Y13_W2BEG[6] ,
    \Tile_X3Y13_W2BEG[5] ,
    \Tile_X3Y13_W2BEG[4] ,
    \Tile_X3Y13_W2BEG[3] ,
    \Tile_X3Y13_W2BEG[2] ,
    \Tile_X3Y13_W2BEG[1] ,
    \Tile_X3Y13_W2BEG[0] }),
    .W6BEG({\Tile_X2Y13_W6BEG[11] ,
    \Tile_X2Y13_W6BEG[10] ,
    \Tile_X2Y13_W6BEG[9] ,
    \Tile_X2Y13_W6BEG[8] ,
    \Tile_X2Y13_W6BEG[7] ,
    \Tile_X2Y13_W6BEG[6] ,
    \Tile_X2Y13_W6BEG[5] ,
    \Tile_X2Y13_W6BEG[4] ,
    \Tile_X2Y13_W6BEG[3] ,
    \Tile_X2Y13_W6BEG[2] ,
    \Tile_X2Y13_W6BEG[1] ,
    \Tile_X2Y13_W6BEG[0] }),
    .W6END({\Tile_X3Y13_W6BEG[11] ,
    \Tile_X3Y13_W6BEG[10] ,
    \Tile_X3Y13_W6BEG[9] ,
    \Tile_X3Y13_W6BEG[8] ,
    \Tile_X3Y13_W6BEG[7] ,
    \Tile_X3Y13_W6BEG[6] ,
    \Tile_X3Y13_W6BEG[5] ,
    \Tile_X3Y13_W6BEG[4] ,
    \Tile_X3Y13_W6BEG[3] ,
    \Tile_X3Y13_W6BEG[2] ,
    \Tile_X3Y13_W6BEG[1] ,
    \Tile_X3Y13_W6BEG[0] }),
    .WW4BEG({\Tile_X2Y13_WW4BEG[15] ,
    \Tile_X2Y13_WW4BEG[14] ,
    \Tile_X2Y13_WW4BEG[13] ,
    \Tile_X2Y13_WW4BEG[12] ,
    \Tile_X2Y13_WW4BEG[11] ,
    \Tile_X2Y13_WW4BEG[10] ,
    \Tile_X2Y13_WW4BEG[9] ,
    \Tile_X2Y13_WW4BEG[8] ,
    \Tile_X2Y13_WW4BEG[7] ,
    \Tile_X2Y13_WW4BEG[6] ,
    \Tile_X2Y13_WW4BEG[5] ,
    \Tile_X2Y13_WW4BEG[4] ,
    \Tile_X2Y13_WW4BEG[3] ,
    \Tile_X2Y13_WW4BEG[2] ,
    \Tile_X2Y13_WW4BEG[1] ,
    \Tile_X2Y13_WW4BEG[0] }),
    .WW4END({\Tile_X3Y13_WW4BEG[15] ,
    \Tile_X3Y13_WW4BEG[14] ,
    \Tile_X3Y13_WW4BEG[13] ,
    \Tile_X3Y13_WW4BEG[12] ,
    \Tile_X3Y13_WW4BEG[11] ,
    \Tile_X3Y13_WW4BEG[10] ,
    \Tile_X3Y13_WW4BEG[9] ,
    \Tile_X3Y13_WW4BEG[8] ,
    \Tile_X3Y13_WW4BEG[7] ,
    \Tile_X3Y13_WW4BEG[6] ,
    \Tile_X3Y13_WW4BEG[5] ,
    \Tile_X3Y13_WW4BEG[4] ,
    \Tile_X3Y13_WW4BEG[3] ,
    \Tile_X3Y13_WW4BEG[2] ,
    \Tile_X3Y13_WW4BEG[1] ,
    \Tile_X3Y13_WW4BEG[0] }));
 LUT4AB Tile_X2Y14_LUT4AB (.Ci(Tile_X2Y15_Co),
    .Co(Tile_X2Y14_Co),
    .UserCLK(Tile_X2Y15_UserCLKo),
    .UserCLKo(Tile_X2Y14_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X2Y14_E1BEG[3] ,
    \Tile_X2Y14_E1BEG[2] ,
    \Tile_X2Y14_E1BEG[1] ,
    \Tile_X2Y14_E1BEG[0] }),
    .E1END({\Tile_X1Y14_E1BEG[3] ,
    \Tile_X1Y14_E1BEG[2] ,
    \Tile_X1Y14_E1BEG[1] ,
    \Tile_X1Y14_E1BEG[0] }),
    .E2BEG({\Tile_X2Y14_E2BEG[7] ,
    \Tile_X2Y14_E2BEG[6] ,
    \Tile_X2Y14_E2BEG[5] ,
    \Tile_X2Y14_E2BEG[4] ,
    \Tile_X2Y14_E2BEG[3] ,
    \Tile_X2Y14_E2BEG[2] ,
    \Tile_X2Y14_E2BEG[1] ,
    \Tile_X2Y14_E2BEG[0] }),
    .E2BEGb({\Tile_X2Y14_E2BEGb[7] ,
    \Tile_X2Y14_E2BEGb[6] ,
    \Tile_X2Y14_E2BEGb[5] ,
    \Tile_X2Y14_E2BEGb[4] ,
    \Tile_X2Y14_E2BEGb[3] ,
    \Tile_X2Y14_E2BEGb[2] ,
    \Tile_X2Y14_E2BEGb[1] ,
    \Tile_X2Y14_E2BEGb[0] }),
    .E2END({\Tile_X1Y14_E2BEGb[7] ,
    \Tile_X1Y14_E2BEGb[6] ,
    \Tile_X1Y14_E2BEGb[5] ,
    \Tile_X1Y14_E2BEGb[4] ,
    \Tile_X1Y14_E2BEGb[3] ,
    \Tile_X1Y14_E2BEGb[2] ,
    \Tile_X1Y14_E2BEGb[1] ,
    \Tile_X1Y14_E2BEGb[0] }),
    .E2MID({\Tile_X1Y14_E2BEG[7] ,
    \Tile_X1Y14_E2BEG[6] ,
    \Tile_X1Y14_E2BEG[5] ,
    \Tile_X1Y14_E2BEG[4] ,
    \Tile_X1Y14_E2BEG[3] ,
    \Tile_X1Y14_E2BEG[2] ,
    \Tile_X1Y14_E2BEG[1] ,
    \Tile_X1Y14_E2BEG[0] }),
    .E6BEG({\Tile_X2Y14_E6BEG[11] ,
    \Tile_X2Y14_E6BEG[10] ,
    \Tile_X2Y14_E6BEG[9] ,
    \Tile_X2Y14_E6BEG[8] ,
    \Tile_X2Y14_E6BEG[7] ,
    \Tile_X2Y14_E6BEG[6] ,
    \Tile_X2Y14_E6BEG[5] ,
    \Tile_X2Y14_E6BEG[4] ,
    \Tile_X2Y14_E6BEG[3] ,
    \Tile_X2Y14_E6BEG[2] ,
    \Tile_X2Y14_E6BEG[1] ,
    \Tile_X2Y14_E6BEG[0] }),
    .E6END({\Tile_X1Y14_E6BEG[11] ,
    \Tile_X1Y14_E6BEG[10] ,
    \Tile_X1Y14_E6BEG[9] ,
    \Tile_X1Y14_E6BEG[8] ,
    \Tile_X1Y14_E6BEG[7] ,
    \Tile_X1Y14_E6BEG[6] ,
    \Tile_X1Y14_E6BEG[5] ,
    \Tile_X1Y14_E6BEG[4] ,
    \Tile_X1Y14_E6BEG[3] ,
    \Tile_X1Y14_E6BEG[2] ,
    \Tile_X1Y14_E6BEG[1] ,
    \Tile_X1Y14_E6BEG[0] }),
    .EE4BEG({\Tile_X2Y14_EE4BEG[15] ,
    \Tile_X2Y14_EE4BEG[14] ,
    \Tile_X2Y14_EE4BEG[13] ,
    \Tile_X2Y14_EE4BEG[12] ,
    \Tile_X2Y14_EE4BEG[11] ,
    \Tile_X2Y14_EE4BEG[10] ,
    \Tile_X2Y14_EE4BEG[9] ,
    \Tile_X2Y14_EE4BEG[8] ,
    \Tile_X2Y14_EE4BEG[7] ,
    \Tile_X2Y14_EE4BEG[6] ,
    \Tile_X2Y14_EE4BEG[5] ,
    \Tile_X2Y14_EE4BEG[4] ,
    \Tile_X2Y14_EE4BEG[3] ,
    \Tile_X2Y14_EE4BEG[2] ,
    \Tile_X2Y14_EE4BEG[1] ,
    \Tile_X2Y14_EE4BEG[0] }),
    .EE4END({\Tile_X1Y14_EE4BEG[15] ,
    \Tile_X1Y14_EE4BEG[14] ,
    \Tile_X1Y14_EE4BEG[13] ,
    \Tile_X1Y14_EE4BEG[12] ,
    \Tile_X1Y14_EE4BEG[11] ,
    \Tile_X1Y14_EE4BEG[10] ,
    \Tile_X1Y14_EE4BEG[9] ,
    \Tile_X1Y14_EE4BEG[8] ,
    \Tile_X1Y14_EE4BEG[7] ,
    \Tile_X1Y14_EE4BEG[6] ,
    \Tile_X1Y14_EE4BEG[5] ,
    \Tile_X1Y14_EE4BEG[4] ,
    \Tile_X1Y14_EE4BEG[3] ,
    \Tile_X1Y14_EE4BEG[2] ,
    \Tile_X1Y14_EE4BEG[1] ,
    \Tile_X1Y14_EE4BEG[0] }),
    .FrameData({\Tile_X1Y14_FrameData_O[31] ,
    \Tile_X1Y14_FrameData_O[30] ,
    \Tile_X1Y14_FrameData_O[29] ,
    \Tile_X1Y14_FrameData_O[28] ,
    \Tile_X1Y14_FrameData_O[27] ,
    \Tile_X1Y14_FrameData_O[26] ,
    \Tile_X1Y14_FrameData_O[25] ,
    \Tile_X1Y14_FrameData_O[24] ,
    \Tile_X1Y14_FrameData_O[23] ,
    \Tile_X1Y14_FrameData_O[22] ,
    \Tile_X1Y14_FrameData_O[21] ,
    \Tile_X1Y14_FrameData_O[20] ,
    \Tile_X1Y14_FrameData_O[19] ,
    \Tile_X1Y14_FrameData_O[18] ,
    \Tile_X1Y14_FrameData_O[17] ,
    \Tile_X1Y14_FrameData_O[16] ,
    \Tile_X1Y14_FrameData_O[15] ,
    \Tile_X1Y14_FrameData_O[14] ,
    \Tile_X1Y14_FrameData_O[13] ,
    \Tile_X1Y14_FrameData_O[12] ,
    \Tile_X1Y14_FrameData_O[11] ,
    \Tile_X1Y14_FrameData_O[10] ,
    \Tile_X1Y14_FrameData_O[9] ,
    \Tile_X1Y14_FrameData_O[8] ,
    \Tile_X1Y14_FrameData_O[7] ,
    \Tile_X1Y14_FrameData_O[6] ,
    \Tile_X1Y14_FrameData_O[5] ,
    \Tile_X1Y14_FrameData_O[4] ,
    \Tile_X1Y14_FrameData_O[3] ,
    \Tile_X1Y14_FrameData_O[2] ,
    \Tile_X1Y14_FrameData_O[1] ,
    \Tile_X1Y14_FrameData_O[0] }),
    .FrameData_O({\Tile_X2Y14_FrameData_O[31] ,
    \Tile_X2Y14_FrameData_O[30] ,
    \Tile_X2Y14_FrameData_O[29] ,
    \Tile_X2Y14_FrameData_O[28] ,
    \Tile_X2Y14_FrameData_O[27] ,
    \Tile_X2Y14_FrameData_O[26] ,
    \Tile_X2Y14_FrameData_O[25] ,
    \Tile_X2Y14_FrameData_O[24] ,
    \Tile_X2Y14_FrameData_O[23] ,
    \Tile_X2Y14_FrameData_O[22] ,
    \Tile_X2Y14_FrameData_O[21] ,
    \Tile_X2Y14_FrameData_O[20] ,
    \Tile_X2Y14_FrameData_O[19] ,
    \Tile_X2Y14_FrameData_O[18] ,
    \Tile_X2Y14_FrameData_O[17] ,
    \Tile_X2Y14_FrameData_O[16] ,
    \Tile_X2Y14_FrameData_O[15] ,
    \Tile_X2Y14_FrameData_O[14] ,
    \Tile_X2Y14_FrameData_O[13] ,
    \Tile_X2Y14_FrameData_O[12] ,
    \Tile_X2Y14_FrameData_O[11] ,
    \Tile_X2Y14_FrameData_O[10] ,
    \Tile_X2Y14_FrameData_O[9] ,
    \Tile_X2Y14_FrameData_O[8] ,
    \Tile_X2Y14_FrameData_O[7] ,
    \Tile_X2Y14_FrameData_O[6] ,
    \Tile_X2Y14_FrameData_O[5] ,
    \Tile_X2Y14_FrameData_O[4] ,
    \Tile_X2Y14_FrameData_O[3] ,
    \Tile_X2Y14_FrameData_O[2] ,
    \Tile_X2Y14_FrameData_O[1] ,
    \Tile_X2Y14_FrameData_O[0] }),
    .FrameStrobe({\Tile_X2Y15_FrameStrobe_O[19] ,
    \Tile_X2Y15_FrameStrobe_O[18] ,
    \Tile_X2Y15_FrameStrobe_O[17] ,
    \Tile_X2Y15_FrameStrobe_O[16] ,
    \Tile_X2Y15_FrameStrobe_O[15] ,
    \Tile_X2Y15_FrameStrobe_O[14] ,
    \Tile_X2Y15_FrameStrobe_O[13] ,
    \Tile_X2Y15_FrameStrobe_O[12] ,
    \Tile_X2Y15_FrameStrobe_O[11] ,
    \Tile_X2Y15_FrameStrobe_O[10] ,
    \Tile_X2Y15_FrameStrobe_O[9] ,
    \Tile_X2Y15_FrameStrobe_O[8] ,
    \Tile_X2Y15_FrameStrobe_O[7] ,
    \Tile_X2Y15_FrameStrobe_O[6] ,
    \Tile_X2Y15_FrameStrobe_O[5] ,
    \Tile_X2Y15_FrameStrobe_O[4] ,
    \Tile_X2Y15_FrameStrobe_O[3] ,
    \Tile_X2Y15_FrameStrobe_O[2] ,
    \Tile_X2Y15_FrameStrobe_O[1] ,
    \Tile_X2Y15_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X2Y14_FrameStrobe_O[19] ,
    \Tile_X2Y14_FrameStrobe_O[18] ,
    \Tile_X2Y14_FrameStrobe_O[17] ,
    \Tile_X2Y14_FrameStrobe_O[16] ,
    \Tile_X2Y14_FrameStrobe_O[15] ,
    \Tile_X2Y14_FrameStrobe_O[14] ,
    \Tile_X2Y14_FrameStrobe_O[13] ,
    \Tile_X2Y14_FrameStrobe_O[12] ,
    \Tile_X2Y14_FrameStrobe_O[11] ,
    \Tile_X2Y14_FrameStrobe_O[10] ,
    \Tile_X2Y14_FrameStrobe_O[9] ,
    \Tile_X2Y14_FrameStrobe_O[8] ,
    \Tile_X2Y14_FrameStrobe_O[7] ,
    \Tile_X2Y14_FrameStrobe_O[6] ,
    \Tile_X2Y14_FrameStrobe_O[5] ,
    \Tile_X2Y14_FrameStrobe_O[4] ,
    \Tile_X2Y14_FrameStrobe_O[3] ,
    \Tile_X2Y14_FrameStrobe_O[2] ,
    \Tile_X2Y14_FrameStrobe_O[1] ,
    \Tile_X2Y14_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X2Y14_N1BEG[3] ,
    \Tile_X2Y14_N1BEG[2] ,
    \Tile_X2Y14_N1BEG[1] ,
    \Tile_X2Y14_N1BEG[0] }),
    .N1END({\Tile_X2Y15_N1BEG[3] ,
    \Tile_X2Y15_N1BEG[2] ,
    \Tile_X2Y15_N1BEG[1] ,
    \Tile_X2Y15_N1BEG[0] }),
    .N2BEG({\Tile_X2Y14_N2BEG[7] ,
    \Tile_X2Y14_N2BEG[6] ,
    \Tile_X2Y14_N2BEG[5] ,
    \Tile_X2Y14_N2BEG[4] ,
    \Tile_X2Y14_N2BEG[3] ,
    \Tile_X2Y14_N2BEG[2] ,
    \Tile_X2Y14_N2BEG[1] ,
    \Tile_X2Y14_N2BEG[0] }),
    .N2BEGb({\Tile_X2Y14_N2BEGb[7] ,
    \Tile_X2Y14_N2BEGb[6] ,
    \Tile_X2Y14_N2BEGb[5] ,
    \Tile_X2Y14_N2BEGb[4] ,
    \Tile_X2Y14_N2BEGb[3] ,
    \Tile_X2Y14_N2BEGb[2] ,
    \Tile_X2Y14_N2BEGb[1] ,
    \Tile_X2Y14_N2BEGb[0] }),
    .N2END({\Tile_X2Y15_N2BEGb[7] ,
    \Tile_X2Y15_N2BEGb[6] ,
    \Tile_X2Y15_N2BEGb[5] ,
    \Tile_X2Y15_N2BEGb[4] ,
    \Tile_X2Y15_N2BEGb[3] ,
    \Tile_X2Y15_N2BEGb[2] ,
    \Tile_X2Y15_N2BEGb[1] ,
    \Tile_X2Y15_N2BEGb[0] }),
    .N2MID({\Tile_X2Y15_N2BEG[7] ,
    \Tile_X2Y15_N2BEG[6] ,
    \Tile_X2Y15_N2BEG[5] ,
    \Tile_X2Y15_N2BEG[4] ,
    \Tile_X2Y15_N2BEG[3] ,
    \Tile_X2Y15_N2BEG[2] ,
    \Tile_X2Y15_N2BEG[1] ,
    \Tile_X2Y15_N2BEG[0] }),
    .N4BEG({\Tile_X2Y14_N4BEG[15] ,
    \Tile_X2Y14_N4BEG[14] ,
    \Tile_X2Y14_N4BEG[13] ,
    \Tile_X2Y14_N4BEG[12] ,
    \Tile_X2Y14_N4BEG[11] ,
    \Tile_X2Y14_N4BEG[10] ,
    \Tile_X2Y14_N4BEG[9] ,
    \Tile_X2Y14_N4BEG[8] ,
    \Tile_X2Y14_N4BEG[7] ,
    \Tile_X2Y14_N4BEG[6] ,
    \Tile_X2Y14_N4BEG[5] ,
    \Tile_X2Y14_N4BEG[4] ,
    \Tile_X2Y14_N4BEG[3] ,
    \Tile_X2Y14_N4BEG[2] ,
    \Tile_X2Y14_N4BEG[1] ,
    \Tile_X2Y14_N4BEG[0] }),
    .N4END({\Tile_X2Y15_N4BEG[15] ,
    \Tile_X2Y15_N4BEG[14] ,
    \Tile_X2Y15_N4BEG[13] ,
    \Tile_X2Y15_N4BEG[12] ,
    \Tile_X2Y15_N4BEG[11] ,
    \Tile_X2Y15_N4BEG[10] ,
    \Tile_X2Y15_N4BEG[9] ,
    \Tile_X2Y15_N4BEG[8] ,
    \Tile_X2Y15_N4BEG[7] ,
    \Tile_X2Y15_N4BEG[6] ,
    \Tile_X2Y15_N4BEG[5] ,
    \Tile_X2Y15_N4BEG[4] ,
    \Tile_X2Y15_N4BEG[3] ,
    \Tile_X2Y15_N4BEG[2] ,
    \Tile_X2Y15_N4BEG[1] ,
    \Tile_X2Y15_N4BEG[0] }),
    .NN4BEG({\Tile_X2Y14_NN4BEG[15] ,
    \Tile_X2Y14_NN4BEG[14] ,
    \Tile_X2Y14_NN4BEG[13] ,
    \Tile_X2Y14_NN4BEG[12] ,
    \Tile_X2Y14_NN4BEG[11] ,
    \Tile_X2Y14_NN4BEG[10] ,
    \Tile_X2Y14_NN4BEG[9] ,
    \Tile_X2Y14_NN4BEG[8] ,
    \Tile_X2Y14_NN4BEG[7] ,
    \Tile_X2Y14_NN4BEG[6] ,
    \Tile_X2Y14_NN4BEG[5] ,
    \Tile_X2Y14_NN4BEG[4] ,
    \Tile_X2Y14_NN4BEG[3] ,
    \Tile_X2Y14_NN4BEG[2] ,
    \Tile_X2Y14_NN4BEG[1] ,
    \Tile_X2Y14_NN4BEG[0] }),
    .NN4END({\Tile_X2Y15_NN4BEG[15] ,
    \Tile_X2Y15_NN4BEG[14] ,
    \Tile_X2Y15_NN4BEG[13] ,
    \Tile_X2Y15_NN4BEG[12] ,
    \Tile_X2Y15_NN4BEG[11] ,
    \Tile_X2Y15_NN4BEG[10] ,
    \Tile_X2Y15_NN4BEG[9] ,
    \Tile_X2Y15_NN4BEG[8] ,
    \Tile_X2Y15_NN4BEG[7] ,
    \Tile_X2Y15_NN4BEG[6] ,
    \Tile_X2Y15_NN4BEG[5] ,
    \Tile_X2Y15_NN4BEG[4] ,
    \Tile_X2Y15_NN4BEG[3] ,
    \Tile_X2Y15_NN4BEG[2] ,
    \Tile_X2Y15_NN4BEG[1] ,
    \Tile_X2Y15_NN4BEG[0] }),
    .S1BEG({\Tile_X2Y14_S1BEG[3] ,
    \Tile_X2Y14_S1BEG[2] ,
    \Tile_X2Y14_S1BEG[1] ,
    \Tile_X2Y14_S1BEG[0] }),
    .S1END({\Tile_X2Y13_S1BEG[3] ,
    \Tile_X2Y13_S1BEG[2] ,
    \Tile_X2Y13_S1BEG[1] ,
    \Tile_X2Y13_S1BEG[0] }),
    .S2BEG({\Tile_X2Y14_S2BEG[7] ,
    \Tile_X2Y14_S2BEG[6] ,
    \Tile_X2Y14_S2BEG[5] ,
    \Tile_X2Y14_S2BEG[4] ,
    \Tile_X2Y14_S2BEG[3] ,
    \Tile_X2Y14_S2BEG[2] ,
    \Tile_X2Y14_S2BEG[1] ,
    \Tile_X2Y14_S2BEG[0] }),
    .S2BEGb({\Tile_X2Y14_S2BEGb[7] ,
    \Tile_X2Y14_S2BEGb[6] ,
    \Tile_X2Y14_S2BEGb[5] ,
    \Tile_X2Y14_S2BEGb[4] ,
    \Tile_X2Y14_S2BEGb[3] ,
    \Tile_X2Y14_S2BEGb[2] ,
    \Tile_X2Y14_S2BEGb[1] ,
    \Tile_X2Y14_S2BEGb[0] }),
    .S2END({\Tile_X2Y13_S2BEGb[7] ,
    \Tile_X2Y13_S2BEGb[6] ,
    \Tile_X2Y13_S2BEGb[5] ,
    \Tile_X2Y13_S2BEGb[4] ,
    \Tile_X2Y13_S2BEGb[3] ,
    \Tile_X2Y13_S2BEGb[2] ,
    \Tile_X2Y13_S2BEGb[1] ,
    \Tile_X2Y13_S2BEGb[0] }),
    .S2MID({\Tile_X2Y13_S2BEG[7] ,
    \Tile_X2Y13_S2BEG[6] ,
    \Tile_X2Y13_S2BEG[5] ,
    \Tile_X2Y13_S2BEG[4] ,
    \Tile_X2Y13_S2BEG[3] ,
    \Tile_X2Y13_S2BEG[2] ,
    \Tile_X2Y13_S2BEG[1] ,
    \Tile_X2Y13_S2BEG[0] }),
    .S4BEG({\Tile_X2Y14_S4BEG[15] ,
    \Tile_X2Y14_S4BEG[14] ,
    \Tile_X2Y14_S4BEG[13] ,
    \Tile_X2Y14_S4BEG[12] ,
    \Tile_X2Y14_S4BEG[11] ,
    \Tile_X2Y14_S4BEG[10] ,
    \Tile_X2Y14_S4BEG[9] ,
    \Tile_X2Y14_S4BEG[8] ,
    \Tile_X2Y14_S4BEG[7] ,
    \Tile_X2Y14_S4BEG[6] ,
    \Tile_X2Y14_S4BEG[5] ,
    \Tile_X2Y14_S4BEG[4] ,
    \Tile_X2Y14_S4BEG[3] ,
    \Tile_X2Y14_S4BEG[2] ,
    \Tile_X2Y14_S4BEG[1] ,
    \Tile_X2Y14_S4BEG[0] }),
    .S4END({\Tile_X2Y13_S4BEG[15] ,
    \Tile_X2Y13_S4BEG[14] ,
    \Tile_X2Y13_S4BEG[13] ,
    \Tile_X2Y13_S4BEG[12] ,
    \Tile_X2Y13_S4BEG[11] ,
    \Tile_X2Y13_S4BEG[10] ,
    \Tile_X2Y13_S4BEG[9] ,
    \Tile_X2Y13_S4BEG[8] ,
    \Tile_X2Y13_S4BEG[7] ,
    \Tile_X2Y13_S4BEG[6] ,
    \Tile_X2Y13_S4BEG[5] ,
    \Tile_X2Y13_S4BEG[4] ,
    \Tile_X2Y13_S4BEG[3] ,
    \Tile_X2Y13_S4BEG[2] ,
    \Tile_X2Y13_S4BEG[1] ,
    \Tile_X2Y13_S4BEG[0] }),
    .SS4BEG({\Tile_X2Y14_SS4BEG[15] ,
    \Tile_X2Y14_SS4BEG[14] ,
    \Tile_X2Y14_SS4BEG[13] ,
    \Tile_X2Y14_SS4BEG[12] ,
    \Tile_X2Y14_SS4BEG[11] ,
    \Tile_X2Y14_SS4BEG[10] ,
    \Tile_X2Y14_SS4BEG[9] ,
    \Tile_X2Y14_SS4BEG[8] ,
    \Tile_X2Y14_SS4BEG[7] ,
    \Tile_X2Y14_SS4BEG[6] ,
    \Tile_X2Y14_SS4BEG[5] ,
    \Tile_X2Y14_SS4BEG[4] ,
    \Tile_X2Y14_SS4BEG[3] ,
    \Tile_X2Y14_SS4BEG[2] ,
    \Tile_X2Y14_SS4BEG[1] ,
    \Tile_X2Y14_SS4BEG[0] }),
    .SS4END({\Tile_X2Y13_SS4BEG[15] ,
    \Tile_X2Y13_SS4BEG[14] ,
    \Tile_X2Y13_SS4BEG[13] ,
    \Tile_X2Y13_SS4BEG[12] ,
    \Tile_X2Y13_SS4BEG[11] ,
    \Tile_X2Y13_SS4BEG[10] ,
    \Tile_X2Y13_SS4BEG[9] ,
    \Tile_X2Y13_SS4BEG[8] ,
    \Tile_X2Y13_SS4BEG[7] ,
    \Tile_X2Y13_SS4BEG[6] ,
    \Tile_X2Y13_SS4BEG[5] ,
    \Tile_X2Y13_SS4BEG[4] ,
    \Tile_X2Y13_SS4BEG[3] ,
    \Tile_X2Y13_SS4BEG[2] ,
    \Tile_X2Y13_SS4BEG[1] ,
    \Tile_X2Y13_SS4BEG[0] }),
    .W1BEG({\Tile_X2Y14_W1BEG[3] ,
    \Tile_X2Y14_W1BEG[2] ,
    \Tile_X2Y14_W1BEG[1] ,
    \Tile_X2Y14_W1BEG[0] }),
    .W1END({\Tile_X3Y14_W1BEG[3] ,
    \Tile_X3Y14_W1BEG[2] ,
    \Tile_X3Y14_W1BEG[1] ,
    \Tile_X3Y14_W1BEG[0] }),
    .W2BEG({\Tile_X2Y14_W2BEG[7] ,
    \Tile_X2Y14_W2BEG[6] ,
    \Tile_X2Y14_W2BEG[5] ,
    \Tile_X2Y14_W2BEG[4] ,
    \Tile_X2Y14_W2BEG[3] ,
    \Tile_X2Y14_W2BEG[2] ,
    \Tile_X2Y14_W2BEG[1] ,
    \Tile_X2Y14_W2BEG[0] }),
    .W2BEGb({\Tile_X2Y14_W2BEGb[7] ,
    \Tile_X2Y14_W2BEGb[6] ,
    \Tile_X2Y14_W2BEGb[5] ,
    \Tile_X2Y14_W2BEGb[4] ,
    \Tile_X2Y14_W2BEGb[3] ,
    \Tile_X2Y14_W2BEGb[2] ,
    \Tile_X2Y14_W2BEGb[1] ,
    \Tile_X2Y14_W2BEGb[0] }),
    .W2END({\Tile_X3Y14_W2BEGb[7] ,
    \Tile_X3Y14_W2BEGb[6] ,
    \Tile_X3Y14_W2BEGb[5] ,
    \Tile_X3Y14_W2BEGb[4] ,
    \Tile_X3Y14_W2BEGb[3] ,
    \Tile_X3Y14_W2BEGb[2] ,
    \Tile_X3Y14_W2BEGb[1] ,
    \Tile_X3Y14_W2BEGb[0] }),
    .W2MID({\Tile_X3Y14_W2BEG[7] ,
    \Tile_X3Y14_W2BEG[6] ,
    \Tile_X3Y14_W2BEG[5] ,
    \Tile_X3Y14_W2BEG[4] ,
    \Tile_X3Y14_W2BEG[3] ,
    \Tile_X3Y14_W2BEG[2] ,
    \Tile_X3Y14_W2BEG[1] ,
    \Tile_X3Y14_W2BEG[0] }),
    .W6BEG({\Tile_X2Y14_W6BEG[11] ,
    \Tile_X2Y14_W6BEG[10] ,
    \Tile_X2Y14_W6BEG[9] ,
    \Tile_X2Y14_W6BEG[8] ,
    \Tile_X2Y14_W6BEG[7] ,
    \Tile_X2Y14_W6BEG[6] ,
    \Tile_X2Y14_W6BEG[5] ,
    \Tile_X2Y14_W6BEG[4] ,
    \Tile_X2Y14_W6BEG[3] ,
    \Tile_X2Y14_W6BEG[2] ,
    \Tile_X2Y14_W6BEG[1] ,
    \Tile_X2Y14_W6BEG[0] }),
    .W6END({\Tile_X3Y14_W6BEG[11] ,
    \Tile_X3Y14_W6BEG[10] ,
    \Tile_X3Y14_W6BEG[9] ,
    \Tile_X3Y14_W6BEG[8] ,
    \Tile_X3Y14_W6BEG[7] ,
    \Tile_X3Y14_W6BEG[6] ,
    \Tile_X3Y14_W6BEG[5] ,
    \Tile_X3Y14_W6BEG[4] ,
    \Tile_X3Y14_W6BEG[3] ,
    \Tile_X3Y14_W6BEG[2] ,
    \Tile_X3Y14_W6BEG[1] ,
    \Tile_X3Y14_W6BEG[0] }),
    .WW4BEG({\Tile_X2Y14_WW4BEG[15] ,
    \Tile_X2Y14_WW4BEG[14] ,
    \Tile_X2Y14_WW4BEG[13] ,
    \Tile_X2Y14_WW4BEG[12] ,
    \Tile_X2Y14_WW4BEG[11] ,
    \Tile_X2Y14_WW4BEG[10] ,
    \Tile_X2Y14_WW4BEG[9] ,
    \Tile_X2Y14_WW4BEG[8] ,
    \Tile_X2Y14_WW4BEG[7] ,
    \Tile_X2Y14_WW4BEG[6] ,
    \Tile_X2Y14_WW4BEG[5] ,
    \Tile_X2Y14_WW4BEG[4] ,
    \Tile_X2Y14_WW4BEG[3] ,
    \Tile_X2Y14_WW4BEG[2] ,
    \Tile_X2Y14_WW4BEG[1] ,
    \Tile_X2Y14_WW4BEG[0] }),
    .WW4END({\Tile_X3Y14_WW4BEG[15] ,
    \Tile_X3Y14_WW4BEG[14] ,
    \Tile_X3Y14_WW4BEG[13] ,
    \Tile_X3Y14_WW4BEG[12] ,
    \Tile_X3Y14_WW4BEG[11] ,
    \Tile_X3Y14_WW4BEG[10] ,
    \Tile_X3Y14_WW4BEG[9] ,
    \Tile_X3Y14_WW4BEG[8] ,
    \Tile_X3Y14_WW4BEG[7] ,
    \Tile_X3Y14_WW4BEG[6] ,
    \Tile_X3Y14_WW4BEG[5] ,
    \Tile_X3Y14_WW4BEG[4] ,
    \Tile_X3Y14_WW4BEG[3] ,
    \Tile_X3Y14_WW4BEG[2] ,
    \Tile_X3Y14_WW4BEG[1] ,
    \Tile_X3Y14_WW4BEG[0] }));
 S_WARMBOOT Tile_X2Y15_S_WARMBOOT (.BOOT_top(Tile_X2Y15_BOOT_top),
    .CONFIGURED_top(Tile_X2Y15_CONFIGURED_top),
    .Co(Tile_X2Y15_Co),
    .RESET_top(Tile_X2Y15_RESET_top),
    .SLOT_top0(Tile_X2Y15_SLOT_top0),
    .SLOT_top1(Tile_X2Y15_SLOT_top1),
    .SLOT_top2(Tile_X2Y15_SLOT_top2),
    .SLOT_top3(Tile_X2Y15_SLOT_top3),
    .UserCLK(UserCLK),
    .UserCLKo(Tile_X2Y15_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .FrameData({\Tile_X1Y15_FrameData_O[31] ,
    \Tile_X1Y15_FrameData_O[30] ,
    \Tile_X1Y15_FrameData_O[29] ,
    \Tile_X1Y15_FrameData_O[28] ,
    \Tile_X1Y15_FrameData_O[27] ,
    \Tile_X1Y15_FrameData_O[26] ,
    \Tile_X1Y15_FrameData_O[25] ,
    \Tile_X1Y15_FrameData_O[24] ,
    \Tile_X1Y15_FrameData_O[23] ,
    \Tile_X1Y15_FrameData_O[22] ,
    \Tile_X1Y15_FrameData_O[21] ,
    \Tile_X1Y15_FrameData_O[20] ,
    \Tile_X1Y15_FrameData_O[19] ,
    \Tile_X1Y15_FrameData_O[18] ,
    \Tile_X1Y15_FrameData_O[17] ,
    \Tile_X1Y15_FrameData_O[16] ,
    \Tile_X1Y15_FrameData_O[15] ,
    \Tile_X1Y15_FrameData_O[14] ,
    \Tile_X1Y15_FrameData_O[13] ,
    \Tile_X1Y15_FrameData_O[12] ,
    \Tile_X1Y15_FrameData_O[11] ,
    \Tile_X1Y15_FrameData_O[10] ,
    \Tile_X1Y15_FrameData_O[9] ,
    \Tile_X1Y15_FrameData_O[8] ,
    \Tile_X1Y15_FrameData_O[7] ,
    \Tile_X1Y15_FrameData_O[6] ,
    \Tile_X1Y15_FrameData_O[5] ,
    \Tile_X1Y15_FrameData_O[4] ,
    \Tile_X1Y15_FrameData_O[3] ,
    \Tile_X1Y15_FrameData_O[2] ,
    \Tile_X1Y15_FrameData_O[1] ,
    \Tile_X1Y15_FrameData_O[0] }),
    .FrameData_O({\Tile_X2Y15_FrameData_O[31] ,
    \Tile_X2Y15_FrameData_O[30] ,
    \Tile_X2Y15_FrameData_O[29] ,
    \Tile_X2Y15_FrameData_O[28] ,
    \Tile_X2Y15_FrameData_O[27] ,
    \Tile_X2Y15_FrameData_O[26] ,
    \Tile_X2Y15_FrameData_O[25] ,
    \Tile_X2Y15_FrameData_O[24] ,
    \Tile_X2Y15_FrameData_O[23] ,
    \Tile_X2Y15_FrameData_O[22] ,
    \Tile_X2Y15_FrameData_O[21] ,
    \Tile_X2Y15_FrameData_O[20] ,
    \Tile_X2Y15_FrameData_O[19] ,
    \Tile_X2Y15_FrameData_O[18] ,
    \Tile_X2Y15_FrameData_O[17] ,
    \Tile_X2Y15_FrameData_O[16] ,
    \Tile_X2Y15_FrameData_O[15] ,
    \Tile_X2Y15_FrameData_O[14] ,
    \Tile_X2Y15_FrameData_O[13] ,
    \Tile_X2Y15_FrameData_O[12] ,
    \Tile_X2Y15_FrameData_O[11] ,
    \Tile_X2Y15_FrameData_O[10] ,
    \Tile_X2Y15_FrameData_O[9] ,
    \Tile_X2Y15_FrameData_O[8] ,
    \Tile_X2Y15_FrameData_O[7] ,
    \Tile_X2Y15_FrameData_O[6] ,
    \Tile_X2Y15_FrameData_O[5] ,
    \Tile_X2Y15_FrameData_O[4] ,
    \Tile_X2Y15_FrameData_O[3] ,
    \Tile_X2Y15_FrameData_O[2] ,
    \Tile_X2Y15_FrameData_O[1] ,
    \Tile_X2Y15_FrameData_O[0] }),
    .FrameStrobe({FrameStrobe[59],
    FrameStrobe[58],
    FrameStrobe[57],
    FrameStrobe[56],
    FrameStrobe[55],
    FrameStrobe[54],
    FrameStrobe[53],
    FrameStrobe[52],
    FrameStrobe[51],
    FrameStrobe[50],
    FrameStrobe[49],
    FrameStrobe[48],
    FrameStrobe[47],
    FrameStrobe[46],
    FrameStrobe[45],
    FrameStrobe[44],
    FrameStrobe[43],
    FrameStrobe[42],
    FrameStrobe[41],
    FrameStrobe[40]}),
    .FrameStrobe_O({\Tile_X2Y15_FrameStrobe_O[19] ,
    \Tile_X2Y15_FrameStrobe_O[18] ,
    \Tile_X2Y15_FrameStrobe_O[17] ,
    \Tile_X2Y15_FrameStrobe_O[16] ,
    \Tile_X2Y15_FrameStrobe_O[15] ,
    \Tile_X2Y15_FrameStrobe_O[14] ,
    \Tile_X2Y15_FrameStrobe_O[13] ,
    \Tile_X2Y15_FrameStrobe_O[12] ,
    \Tile_X2Y15_FrameStrobe_O[11] ,
    \Tile_X2Y15_FrameStrobe_O[10] ,
    \Tile_X2Y15_FrameStrobe_O[9] ,
    \Tile_X2Y15_FrameStrobe_O[8] ,
    \Tile_X2Y15_FrameStrobe_O[7] ,
    \Tile_X2Y15_FrameStrobe_O[6] ,
    \Tile_X2Y15_FrameStrobe_O[5] ,
    \Tile_X2Y15_FrameStrobe_O[4] ,
    \Tile_X2Y15_FrameStrobe_O[3] ,
    \Tile_X2Y15_FrameStrobe_O[2] ,
    \Tile_X2Y15_FrameStrobe_O[1] ,
    \Tile_X2Y15_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X2Y15_N1BEG[3] ,
    \Tile_X2Y15_N1BEG[2] ,
    \Tile_X2Y15_N1BEG[1] ,
    \Tile_X2Y15_N1BEG[0] }),
    .N2BEG({\Tile_X2Y15_N2BEG[7] ,
    \Tile_X2Y15_N2BEG[6] ,
    \Tile_X2Y15_N2BEG[5] ,
    \Tile_X2Y15_N2BEG[4] ,
    \Tile_X2Y15_N2BEG[3] ,
    \Tile_X2Y15_N2BEG[2] ,
    \Tile_X2Y15_N2BEG[1] ,
    \Tile_X2Y15_N2BEG[0] }),
    .N2BEGb({\Tile_X2Y15_N2BEGb[7] ,
    \Tile_X2Y15_N2BEGb[6] ,
    \Tile_X2Y15_N2BEGb[5] ,
    \Tile_X2Y15_N2BEGb[4] ,
    \Tile_X2Y15_N2BEGb[3] ,
    \Tile_X2Y15_N2BEGb[2] ,
    \Tile_X2Y15_N2BEGb[1] ,
    \Tile_X2Y15_N2BEGb[0] }),
    .N4BEG({\Tile_X2Y15_N4BEG[15] ,
    \Tile_X2Y15_N4BEG[14] ,
    \Tile_X2Y15_N4BEG[13] ,
    \Tile_X2Y15_N4BEG[12] ,
    \Tile_X2Y15_N4BEG[11] ,
    \Tile_X2Y15_N4BEG[10] ,
    \Tile_X2Y15_N4BEG[9] ,
    \Tile_X2Y15_N4BEG[8] ,
    \Tile_X2Y15_N4BEG[7] ,
    \Tile_X2Y15_N4BEG[6] ,
    \Tile_X2Y15_N4BEG[5] ,
    \Tile_X2Y15_N4BEG[4] ,
    \Tile_X2Y15_N4BEG[3] ,
    \Tile_X2Y15_N4BEG[2] ,
    \Tile_X2Y15_N4BEG[1] ,
    \Tile_X2Y15_N4BEG[0] }),
    .NN4BEG({\Tile_X2Y15_NN4BEG[15] ,
    \Tile_X2Y15_NN4BEG[14] ,
    \Tile_X2Y15_NN4BEG[13] ,
    \Tile_X2Y15_NN4BEG[12] ,
    \Tile_X2Y15_NN4BEG[11] ,
    \Tile_X2Y15_NN4BEG[10] ,
    \Tile_X2Y15_NN4BEG[9] ,
    \Tile_X2Y15_NN4BEG[8] ,
    \Tile_X2Y15_NN4BEG[7] ,
    \Tile_X2Y15_NN4BEG[6] ,
    \Tile_X2Y15_NN4BEG[5] ,
    \Tile_X2Y15_NN4BEG[4] ,
    \Tile_X2Y15_NN4BEG[3] ,
    \Tile_X2Y15_NN4BEG[2] ,
    \Tile_X2Y15_NN4BEG[1] ,
    \Tile_X2Y15_NN4BEG[0] }),
    .S1END({\Tile_X2Y14_S1BEG[3] ,
    \Tile_X2Y14_S1BEG[2] ,
    \Tile_X2Y14_S1BEG[1] ,
    \Tile_X2Y14_S1BEG[0] }),
    .S2END({\Tile_X2Y14_S2BEGb[7] ,
    \Tile_X2Y14_S2BEGb[6] ,
    \Tile_X2Y14_S2BEGb[5] ,
    \Tile_X2Y14_S2BEGb[4] ,
    \Tile_X2Y14_S2BEGb[3] ,
    \Tile_X2Y14_S2BEGb[2] ,
    \Tile_X2Y14_S2BEGb[1] ,
    \Tile_X2Y14_S2BEGb[0] }),
    .S2MID({\Tile_X2Y14_S2BEG[7] ,
    \Tile_X2Y14_S2BEG[6] ,
    \Tile_X2Y14_S2BEG[5] ,
    \Tile_X2Y14_S2BEG[4] ,
    \Tile_X2Y14_S2BEG[3] ,
    \Tile_X2Y14_S2BEG[2] ,
    \Tile_X2Y14_S2BEG[1] ,
    \Tile_X2Y14_S2BEG[0] }),
    .S4END({\Tile_X2Y14_S4BEG[15] ,
    \Tile_X2Y14_S4BEG[14] ,
    \Tile_X2Y14_S4BEG[13] ,
    \Tile_X2Y14_S4BEG[12] ,
    \Tile_X2Y14_S4BEG[11] ,
    \Tile_X2Y14_S4BEG[10] ,
    \Tile_X2Y14_S4BEG[9] ,
    \Tile_X2Y14_S4BEG[8] ,
    \Tile_X2Y14_S4BEG[7] ,
    \Tile_X2Y14_S4BEG[6] ,
    \Tile_X2Y14_S4BEG[5] ,
    \Tile_X2Y14_S4BEG[4] ,
    \Tile_X2Y14_S4BEG[3] ,
    \Tile_X2Y14_S4BEG[2] ,
    \Tile_X2Y14_S4BEG[1] ,
    \Tile_X2Y14_S4BEG[0] }),
    .SS4END({\Tile_X2Y14_SS4BEG[15] ,
    \Tile_X2Y14_SS4BEG[14] ,
    \Tile_X2Y14_SS4BEG[13] ,
    \Tile_X2Y14_SS4BEG[12] ,
    \Tile_X2Y14_SS4BEG[11] ,
    \Tile_X2Y14_SS4BEG[10] ,
    \Tile_X2Y14_SS4BEG[9] ,
    \Tile_X2Y14_SS4BEG[8] ,
    \Tile_X2Y14_SS4BEG[7] ,
    \Tile_X2Y14_SS4BEG[6] ,
    \Tile_X2Y14_SS4BEG[5] ,
    \Tile_X2Y14_SS4BEG[4] ,
    \Tile_X2Y14_SS4BEG[3] ,
    \Tile_X2Y14_SS4BEG[2] ,
    \Tile_X2Y14_SS4BEG[1] ,
    \Tile_X2Y14_SS4BEG[0] }));
 LUT4AB Tile_X2Y1_LUT4AB (.Ci(Tile_X2Y2_Co),
    .Co(Tile_X2Y1_Co),
    .UserCLK(Tile_X2Y2_UserCLKo),
    .UserCLKo(Tile_X2Y1_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X2Y1_E1BEG[3] ,
    \Tile_X2Y1_E1BEG[2] ,
    \Tile_X2Y1_E1BEG[1] ,
    \Tile_X2Y1_E1BEG[0] }),
    .E1END({\Tile_X1Y1_E1BEG[3] ,
    \Tile_X1Y1_E1BEG[2] ,
    \Tile_X1Y1_E1BEG[1] ,
    \Tile_X1Y1_E1BEG[0] }),
    .E2BEG({\Tile_X2Y1_E2BEG[7] ,
    \Tile_X2Y1_E2BEG[6] ,
    \Tile_X2Y1_E2BEG[5] ,
    \Tile_X2Y1_E2BEG[4] ,
    \Tile_X2Y1_E2BEG[3] ,
    \Tile_X2Y1_E2BEG[2] ,
    \Tile_X2Y1_E2BEG[1] ,
    \Tile_X2Y1_E2BEG[0] }),
    .E2BEGb({\Tile_X2Y1_E2BEGb[7] ,
    \Tile_X2Y1_E2BEGb[6] ,
    \Tile_X2Y1_E2BEGb[5] ,
    \Tile_X2Y1_E2BEGb[4] ,
    \Tile_X2Y1_E2BEGb[3] ,
    \Tile_X2Y1_E2BEGb[2] ,
    \Tile_X2Y1_E2BEGb[1] ,
    \Tile_X2Y1_E2BEGb[0] }),
    .E2END({\Tile_X1Y1_E2BEGb[7] ,
    \Tile_X1Y1_E2BEGb[6] ,
    \Tile_X1Y1_E2BEGb[5] ,
    \Tile_X1Y1_E2BEGb[4] ,
    \Tile_X1Y1_E2BEGb[3] ,
    \Tile_X1Y1_E2BEGb[2] ,
    \Tile_X1Y1_E2BEGb[1] ,
    \Tile_X1Y1_E2BEGb[0] }),
    .E2MID({\Tile_X1Y1_E2BEG[7] ,
    \Tile_X1Y1_E2BEG[6] ,
    \Tile_X1Y1_E2BEG[5] ,
    \Tile_X1Y1_E2BEG[4] ,
    \Tile_X1Y1_E2BEG[3] ,
    \Tile_X1Y1_E2BEG[2] ,
    \Tile_X1Y1_E2BEG[1] ,
    \Tile_X1Y1_E2BEG[0] }),
    .E6BEG({\Tile_X2Y1_E6BEG[11] ,
    \Tile_X2Y1_E6BEG[10] ,
    \Tile_X2Y1_E6BEG[9] ,
    \Tile_X2Y1_E6BEG[8] ,
    \Tile_X2Y1_E6BEG[7] ,
    \Tile_X2Y1_E6BEG[6] ,
    \Tile_X2Y1_E6BEG[5] ,
    \Tile_X2Y1_E6BEG[4] ,
    \Tile_X2Y1_E6BEG[3] ,
    \Tile_X2Y1_E6BEG[2] ,
    \Tile_X2Y1_E6BEG[1] ,
    \Tile_X2Y1_E6BEG[0] }),
    .E6END({\Tile_X1Y1_E6BEG[11] ,
    \Tile_X1Y1_E6BEG[10] ,
    \Tile_X1Y1_E6BEG[9] ,
    \Tile_X1Y1_E6BEG[8] ,
    \Tile_X1Y1_E6BEG[7] ,
    \Tile_X1Y1_E6BEG[6] ,
    \Tile_X1Y1_E6BEG[5] ,
    \Tile_X1Y1_E6BEG[4] ,
    \Tile_X1Y1_E6BEG[3] ,
    \Tile_X1Y1_E6BEG[2] ,
    \Tile_X1Y1_E6BEG[1] ,
    \Tile_X1Y1_E6BEG[0] }),
    .EE4BEG({\Tile_X2Y1_EE4BEG[15] ,
    \Tile_X2Y1_EE4BEG[14] ,
    \Tile_X2Y1_EE4BEG[13] ,
    \Tile_X2Y1_EE4BEG[12] ,
    \Tile_X2Y1_EE4BEG[11] ,
    \Tile_X2Y1_EE4BEG[10] ,
    \Tile_X2Y1_EE4BEG[9] ,
    \Tile_X2Y1_EE4BEG[8] ,
    \Tile_X2Y1_EE4BEG[7] ,
    \Tile_X2Y1_EE4BEG[6] ,
    \Tile_X2Y1_EE4BEG[5] ,
    \Tile_X2Y1_EE4BEG[4] ,
    \Tile_X2Y1_EE4BEG[3] ,
    \Tile_X2Y1_EE4BEG[2] ,
    \Tile_X2Y1_EE4BEG[1] ,
    \Tile_X2Y1_EE4BEG[0] }),
    .EE4END({\Tile_X1Y1_EE4BEG[15] ,
    \Tile_X1Y1_EE4BEG[14] ,
    \Tile_X1Y1_EE4BEG[13] ,
    \Tile_X1Y1_EE4BEG[12] ,
    \Tile_X1Y1_EE4BEG[11] ,
    \Tile_X1Y1_EE4BEG[10] ,
    \Tile_X1Y1_EE4BEG[9] ,
    \Tile_X1Y1_EE4BEG[8] ,
    \Tile_X1Y1_EE4BEG[7] ,
    \Tile_X1Y1_EE4BEG[6] ,
    \Tile_X1Y1_EE4BEG[5] ,
    \Tile_X1Y1_EE4BEG[4] ,
    \Tile_X1Y1_EE4BEG[3] ,
    \Tile_X1Y1_EE4BEG[2] ,
    \Tile_X1Y1_EE4BEG[1] ,
    \Tile_X1Y1_EE4BEG[0] }),
    .FrameData({\Tile_X1Y1_FrameData_O[31] ,
    \Tile_X1Y1_FrameData_O[30] ,
    \Tile_X1Y1_FrameData_O[29] ,
    \Tile_X1Y1_FrameData_O[28] ,
    \Tile_X1Y1_FrameData_O[27] ,
    \Tile_X1Y1_FrameData_O[26] ,
    \Tile_X1Y1_FrameData_O[25] ,
    \Tile_X1Y1_FrameData_O[24] ,
    \Tile_X1Y1_FrameData_O[23] ,
    \Tile_X1Y1_FrameData_O[22] ,
    \Tile_X1Y1_FrameData_O[21] ,
    \Tile_X1Y1_FrameData_O[20] ,
    \Tile_X1Y1_FrameData_O[19] ,
    \Tile_X1Y1_FrameData_O[18] ,
    \Tile_X1Y1_FrameData_O[17] ,
    \Tile_X1Y1_FrameData_O[16] ,
    \Tile_X1Y1_FrameData_O[15] ,
    \Tile_X1Y1_FrameData_O[14] ,
    \Tile_X1Y1_FrameData_O[13] ,
    \Tile_X1Y1_FrameData_O[12] ,
    \Tile_X1Y1_FrameData_O[11] ,
    \Tile_X1Y1_FrameData_O[10] ,
    \Tile_X1Y1_FrameData_O[9] ,
    \Tile_X1Y1_FrameData_O[8] ,
    \Tile_X1Y1_FrameData_O[7] ,
    \Tile_X1Y1_FrameData_O[6] ,
    \Tile_X1Y1_FrameData_O[5] ,
    \Tile_X1Y1_FrameData_O[4] ,
    \Tile_X1Y1_FrameData_O[3] ,
    \Tile_X1Y1_FrameData_O[2] ,
    \Tile_X1Y1_FrameData_O[1] ,
    \Tile_X1Y1_FrameData_O[0] }),
    .FrameData_O({\Tile_X2Y1_FrameData_O[31] ,
    \Tile_X2Y1_FrameData_O[30] ,
    \Tile_X2Y1_FrameData_O[29] ,
    \Tile_X2Y1_FrameData_O[28] ,
    \Tile_X2Y1_FrameData_O[27] ,
    \Tile_X2Y1_FrameData_O[26] ,
    \Tile_X2Y1_FrameData_O[25] ,
    \Tile_X2Y1_FrameData_O[24] ,
    \Tile_X2Y1_FrameData_O[23] ,
    \Tile_X2Y1_FrameData_O[22] ,
    \Tile_X2Y1_FrameData_O[21] ,
    \Tile_X2Y1_FrameData_O[20] ,
    \Tile_X2Y1_FrameData_O[19] ,
    \Tile_X2Y1_FrameData_O[18] ,
    \Tile_X2Y1_FrameData_O[17] ,
    \Tile_X2Y1_FrameData_O[16] ,
    \Tile_X2Y1_FrameData_O[15] ,
    \Tile_X2Y1_FrameData_O[14] ,
    \Tile_X2Y1_FrameData_O[13] ,
    \Tile_X2Y1_FrameData_O[12] ,
    \Tile_X2Y1_FrameData_O[11] ,
    \Tile_X2Y1_FrameData_O[10] ,
    \Tile_X2Y1_FrameData_O[9] ,
    \Tile_X2Y1_FrameData_O[8] ,
    \Tile_X2Y1_FrameData_O[7] ,
    \Tile_X2Y1_FrameData_O[6] ,
    \Tile_X2Y1_FrameData_O[5] ,
    \Tile_X2Y1_FrameData_O[4] ,
    \Tile_X2Y1_FrameData_O[3] ,
    \Tile_X2Y1_FrameData_O[2] ,
    \Tile_X2Y1_FrameData_O[1] ,
    \Tile_X2Y1_FrameData_O[0] }),
    .FrameStrobe({\Tile_X2Y2_FrameStrobe_O[19] ,
    \Tile_X2Y2_FrameStrobe_O[18] ,
    \Tile_X2Y2_FrameStrobe_O[17] ,
    \Tile_X2Y2_FrameStrobe_O[16] ,
    \Tile_X2Y2_FrameStrobe_O[15] ,
    \Tile_X2Y2_FrameStrobe_O[14] ,
    \Tile_X2Y2_FrameStrobe_O[13] ,
    \Tile_X2Y2_FrameStrobe_O[12] ,
    \Tile_X2Y2_FrameStrobe_O[11] ,
    \Tile_X2Y2_FrameStrobe_O[10] ,
    \Tile_X2Y2_FrameStrobe_O[9] ,
    \Tile_X2Y2_FrameStrobe_O[8] ,
    \Tile_X2Y2_FrameStrobe_O[7] ,
    \Tile_X2Y2_FrameStrobe_O[6] ,
    \Tile_X2Y2_FrameStrobe_O[5] ,
    \Tile_X2Y2_FrameStrobe_O[4] ,
    \Tile_X2Y2_FrameStrobe_O[3] ,
    \Tile_X2Y2_FrameStrobe_O[2] ,
    \Tile_X2Y2_FrameStrobe_O[1] ,
    \Tile_X2Y2_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X2Y1_FrameStrobe_O[19] ,
    \Tile_X2Y1_FrameStrobe_O[18] ,
    \Tile_X2Y1_FrameStrobe_O[17] ,
    \Tile_X2Y1_FrameStrobe_O[16] ,
    \Tile_X2Y1_FrameStrobe_O[15] ,
    \Tile_X2Y1_FrameStrobe_O[14] ,
    \Tile_X2Y1_FrameStrobe_O[13] ,
    \Tile_X2Y1_FrameStrobe_O[12] ,
    \Tile_X2Y1_FrameStrobe_O[11] ,
    \Tile_X2Y1_FrameStrobe_O[10] ,
    \Tile_X2Y1_FrameStrobe_O[9] ,
    \Tile_X2Y1_FrameStrobe_O[8] ,
    \Tile_X2Y1_FrameStrobe_O[7] ,
    \Tile_X2Y1_FrameStrobe_O[6] ,
    \Tile_X2Y1_FrameStrobe_O[5] ,
    \Tile_X2Y1_FrameStrobe_O[4] ,
    \Tile_X2Y1_FrameStrobe_O[3] ,
    \Tile_X2Y1_FrameStrobe_O[2] ,
    \Tile_X2Y1_FrameStrobe_O[1] ,
    \Tile_X2Y1_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X2Y1_N1BEG[3] ,
    \Tile_X2Y1_N1BEG[2] ,
    \Tile_X2Y1_N1BEG[1] ,
    \Tile_X2Y1_N1BEG[0] }),
    .N1END({\Tile_X2Y2_N1BEG[3] ,
    \Tile_X2Y2_N1BEG[2] ,
    \Tile_X2Y2_N1BEG[1] ,
    \Tile_X2Y2_N1BEG[0] }),
    .N2BEG({\Tile_X2Y1_N2BEG[7] ,
    \Tile_X2Y1_N2BEG[6] ,
    \Tile_X2Y1_N2BEG[5] ,
    \Tile_X2Y1_N2BEG[4] ,
    \Tile_X2Y1_N2BEG[3] ,
    \Tile_X2Y1_N2BEG[2] ,
    \Tile_X2Y1_N2BEG[1] ,
    \Tile_X2Y1_N2BEG[0] }),
    .N2BEGb({\Tile_X2Y1_N2BEGb[7] ,
    \Tile_X2Y1_N2BEGb[6] ,
    \Tile_X2Y1_N2BEGb[5] ,
    \Tile_X2Y1_N2BEGb[4] ,
    \Tile_X2Y1_N2BEGb[3] ,
    \Tile_X2Y1_N2BEGb[2] ,
    \Tile_X2Y1_N2BEGb[1] ,
    \Tile_X2Y1_N2BEGb[0] }),
    .N2END({\Tile_X2Y2_N2BEGb[7] ,
    \Tile_X2Y2_N2BEGb[6] ,
    \Tile_X2Y2_N2BEGb[5] ,
    \Tile_X2Y2_N2BEGb[4] ,
    \Tile_X2Y2_N2BEGb[3] ,
    \Tile_X2Y2_N2BEGb[2] ,
    \Tile_X2Y2_N2BEGb[1] ,
    \Tile_X2Y2_N2BEGb[0] }),
    .N2MID({\Tile_X2Y2_N2BEG[7] ,
    \Tile_X2Y2_N2BEG[6] ,
    \Tile_X2Y2_N2BEG[5] ,
    \Tile_X2Y2_N2BEG[4] ,
    \Tile_X2Y2_N2BEG[3] ,
    \Tile_X2Y2_N2BEG[2] ,
    \Tile_X2Y2_N2BEG[1] ,
    \Tile_X2Y2_N2BEG[0] }),
    .N4BEG({\Tile_X2Y1_N4BEG[15] ,
    \Tile_X2Y1_N4BEG[14] ,
    \Tile_X2Y1_N4BEG[13] ,
    \Tile_X2Y1_N4BEG[12] ,
    \Tile_X2Y1_N4BEG[11] ,
    \Tile_X2Y1_N4BEG[10] ,
    \Tile_X2Y1_N4BEG[9] ,
    \Tile_X2Y1_N4BEG[8] ,
    \Tile_X2Y1_N4BEG[7] ,
    \Tile_X2Y1_N4BEG[6] ,
    \Tile_X2Y1_N4BEG[5] ,
    \Tile_X2Y1_N4BEG[4] ,
    \Tile_X2Y1_N4BEG[3] ,
    \Tile_X2Y1_N4BEG[2] ,
    \Tile_X2Y1_N4BEG[1] ,
    \Tile_X2Y1_N4BEG[0] }),
    .N4END({\Tile_X2Y2_N4BEG[15] ,
    \Tile_X2Y2_N4BEG[14] ,
    \Tile_X2Y2_N4BEG[13] ,
    \Tile_X2Y2_N4BEG[12] ,
    \Tile_X2Y2_N4BEG[11] ,
    \Tile_X2Y2_N4BEG[10] ,
    \Tile_X2Y2_N4BEG[9] ,
    \Tile_X2Y2_N4BEG[8] ,
    \Tile_X2Y2_N4BEG[7] ,
    \Tile_X2Y2_N4BEG[6] ,
    \Tile_X2Y2_N4BEG[5] ,
    \Tile_X2Y2_N4BEG[4] ,
    \Tile_X2Y2_N4BEG[3] ,
    \Tile_X2Y2_N4BEG[2] ,
    \Tile_X2Y2_N4BEG[1] ,
    \Tile_X2Y2_N4BEG[0] }),
    .NN4BEG({\Tile_X2Y1_NN4BEG[15] ,
    \Tile_X2Y1_NN4BEG[14] ,
    \Tile_X2Y1_NN4BEG[13] ,
    \Tile_X2Y1_NN4BEG[12] ,
    \Tile_X2Y1_NN4BEG[11] ,
    \Tile_X2Y1_NN4BEG[10] ,
    \Tile_X2Y1_NN4BEG[9] ,
    \Tile_X2Y1_NN4BEG[8] ,
    \Tile_X2Y1_NN4BEG[7] ,
    \Tile_X2Y1_NN4BEG[6] ,
    \Tile_X2Y1_NN4BEG[5] ,
    \Tile_X2Y1_NN4BEG[4] ,
    \Tile_X2Y1_NN4BEG[3] ,
    \Tile_X2Y1_NN4BEG[2] ,
    \Tile_X2Y1_NN4BEG[1] ,
    \Tile_X2Y1_NN4BEG[0] }),
    .NN4END({\Tile_X2Y2_NN4BEG[15] ,
    \Tile_X2Y2_NN4BEG[14] ,
    \Tile_X2Y2_NN4BEG[13] ,
    \Tile_X2Y2_NN4BEG[12] ,
    \Tile_X2Y2_NN4BEG[11] ,
    \Tile_X2Y2_NN4BEG[10] ,
    \Tile_X2Y2_NN4BEG[9] ,
    \Tile_X2Y2_NN4BEG[8] ,
    \Tile_X2Y2_NN4BEG[7] ,
    \Tile_X2Y2_NN4BEG[6] ,
    \Tile_X2Y2_NN4BEG[5] ,
    \Tile_X2Y2_NN4BEG[4] ,
    \Tile_X2Y2_NN4BEG[3] ,
    \Tile_X2Y2_NN4BEG[2] ,
    \Tile_X2Y2_NN4BEG[1] ,
    \Tile_X2Y2_NN4BEG[0] }),
    .S1BEG({\Tile_X2Y1_S1BEG[3] ,
    \Tile_X2Y1_S1BEG[2] ,
    \Tile_X2Y1_S1BEG[1] ,
    \Tile_X2Y1_S1BEG[0] }),
    .S1END({\Tile_X2Y0_S1BEG[3] ,
    \Tile_X2Y0_S1BEG[2] ,
    \Tile_X2Y0_S1BEG[1] ,
    \Tile_X2Y0_S1BEG[0] }),
    .S2BEG({\Tile_X2Y1_S2BEG[7] ,
    \Tile_X2Y1_S2BEG[6] ,
    \Tile_X2Y1_S2BEG[5] ,
    \Tile_X2Y1_S2BEG[4] ,
    \Tile_X2Y1_S2BEG[3] ,
    \Tile_X2Y1_S2BEG[2] ,
    \Tile_X2Y1_S2BEG[1] ,
    \Tile_X2Y1_S2BEG[0] }),
    .S2BEGb({\Tile_X2Y1_S2BEGb[7] ,
    \Tile_X2Y1_S2BEGb[6] ,
    \Tile_X2Y1_S2BEGb[5] ,
    \Tile_X2Y1_S2BEGb[4] ,
    \Tile_X2Y1_S2BEGb[3] ,
    \Tile_X2Y1_S2BEGb[2] ,
    \Tile_X2Y1_S2BEGb[1] ,
    \Tile_X2Y1_S2BEGb[0] }),
    .S2END({\Tile_X2Y0_S2BEGb[7] ,
    \Tile_X2Y0_S2BEGb[6] ,
    \Tile_X2Y0_S2BEGb[5] ,
    \Tile_X2Y0_S2BEGb[4] ,
    \Tile_X2Y0_S2BEGb[3] ,
    \Tile_X2Y0_S2BEGb[2] ,
    \Tile_X2Y0_S2BEGb[1] ,
    \Tile_X2Y0_S2BEGb[0] }),
    .S2MID({\Tile_X2Y0_S2BEG[7] ,
    \Tile_X2Y0_S2BEG[6] ,
    \Tile_X2Y0_S2BEG[5] ,
    \Tile_X2Y0_S2BEG[4] ,
    \Tile_X2Y0_S2BEG[3] ,
    \Tile_X2Y0_S2BEG[2] ,
    \Tile_X2Y0_S2BEG[1] ,
    \Tile_X2Y0_S2BEG[0] }),
    .S4BEG({\Tile_X2Y1_S4BEG[15] ,
    \Tile_X2Y1_S4BEG[14] ,
    \Tile_X2Y1_S4BEG[13] ,
    \Tile_X2Y1_S4BEG[12] ,
    \Tile_X2Y1_S4BEG[11] ,
    \Tile_X2Y1_S4BEG[10] ,
    \Tile_X2Y1_S4BEG[9] ,
    \Tile_X2Y1_S4BEG[8] ,
    \Tile_X2Y1_S4BEG[7] ,
    \Tile_X2Y1_S4BEG[6] ,
    \Tile_X2Y1_S4BEG[5] ,
    \Tile_X2Y1_S4BEG[4] ,
    \Tile_X2Y1_S4BEG[3] ,
    \Tile_X2Y1_S4BEG[2] ,
    \Tile_X2Y1_S4BEG[1] ,
    \Tile_X2Y1_S4BEG[0] }),
    .S4END({\Tile_X2Y0_S4BEG[15] ,
    \Tile_X2Y0_S4BEG[14] ,
    \Tile_X2Y0_S4BEG[13] ,
    \Tile_X2Y0_S4BEG[12] ,
    \Tile_X2Y0_S4BEG[11] ,
    \Tile_X2Y0_S4BEG[10] ,
    \Tile_X2Y0_S4BEG[9] ,
    \Tile_X2Y0_S4BEG[8] ,
    \Tile_X2Y0_S4BEG[7] ,
    \Tile_X2Y0_S4BEG[6] ,
    \Tile_X2Y0_S4BEG[5] ,
    \Tile_X2Y0_S4BEG[4] ,
    \Tile_X2Y0_S4BEG[3] ,
    \Tile_X2Y0_S4BEG[2] ,
    \Tile_X2Y0_S4BEG[1] ,
    \Tile_X2Y0_S4BEG[0] }),
    .SS4BEG({\Tile_X2Y1_SS4BEG[15] ,
    \Tile_X2Y1_SS4BEG[14] ,
    \Tile_X2Y1_SS4BEG[13] ,
    \Tile_X2Y1_SS4BEG[12] ,
    \Tile_X2Y1_SS4BEG[11] ,
    \Tile_X2Y1_SS4BEG[10] ,
    \Tile_X2Y1_SS4BEG[9] ,
    \Tile_X2Y1_SS4BEG[8] ,
    \Tile_X2Y1_SS4BEG[7] ,
    \Tile_X2Y1_SS4BEG[6] ,
    \Tile_X2Y1_SS4BEG[5] ,
    \Tile_X2Y1_SS4BEG[4] ,
    \Tile_X2Y1_SS4BEG[3] ,
    \Tile_X2Y1_SS4BEG[2] ,
    \Tile_X2Y1_SS4BEG[1] ,
    \Tile_X2Y1_SS4BEG[0] }),
    .SS4END({\Tile_X2Y0_SS4BEG[15] ,
    \Tile_X2Y0_SS4BEG[14] ,
    \Tile_X2Y0_SS4BEG[13] ,
    \Tile_X2Y0_SS4BEG[12] ,
    \Tile_X2Y0_SS4BEG[11] ,
    \Tile_X2Y0_SS4BEG[10] ,
    \Tile_X2Y0_SS4BEG[9] ,
    \Tile_X2Y0_SS4BEG[8] ,
    \Tile_X2Y0_SS4BEG[7] ,
    \Tile_X2Y0_SS4BEG[6] ,
    \Tile_X2Y0_SS4BEG[5] ,
    \Tile_X2Y0_SS4BEG[4] ,
    \Tile_X2Y0_SS4BEG[3] ,
    \Tile_X2Y0_SS4BEG[2] ,
    \Tile_X2Y0_SS4BEG[1] ,
    \Tile_X2Y0_SS4BEG[0] }),
    .W1BEG({\Tile_X2Y1_W1BEG[3] ,
    \Tile_X2Y1_W1BEG[2] ,
    \Tile_X2Y1_W1BEG[1] ,
    \Tile_X2Y1_W1BEG[0] }),
    .W1END({\Tile_X3Y1_W1BEG[3] ,
    \Tile_X3Y1_W1BEG[2] ,
    \Tile_X3Y1_W1BEG[1] ,
    \Tile_X3Y1_W1BEG[0] }),
    .W2BEG({\Tile_X2Y1_W2BEG[7] ,
    \Tile_X2Y1_W2BEG[6] ,
    \Tile_X2Y1_W2BEG[5] ,
    \Tile_X2Y1_W2BEG[4] ,
    \Tile_X2Y1_W2BEG[3] ,
    \Tile_X2Y1_W2BEG[2] ,
    \Tile_X2Y1_W2BEG[1] ,
    \Tile_X2Y1_W2BEG[0] }),
    .W2BEGb({\Tile_X2Y1_W2BEGb[7] ,
    \Tile_X2Y1_W2BEGb[6] ,
    \Tile_X2Y1_W2BEGb[5] ,
    \Tile_X2Y1_W2BEGb[4] ,
    \Tile_X2Y1_W2BEGb[3] ,
    \Tile_X2Y1_W2BEGb[2] ,
    \Tile_X2Y1_W2BEGb[1] ,
    \Tile_X2Y1_W2BEGb[0] }),
    .W2END({\Tile_X3Y1_W2BEGb[7] ,
    \Tile_X3Y1_W2BEGb[6] ,
    \Tile_X3Y1_W2BEGb[5] ,
    \Tile_X3Y1_W2BEGb[4] ,
    \Tile_X3Y1_W2BEGb[3] ,
    \Tile_X3Y1_W2BEGb[2] ,
    \Tile_X3Y1_W2BEGb[1] ,
    \Tile_X3Y1_W2BEGb[0] }),
    .W2MID({\Tile_X3Y1_W2BEG[7] ,
    \Tile_X3Y1_W2BEG[6] ,
    \Tile_X3Y1_W2BEG[5] ,
    \Tile_X3Y1_W2BEG[4] ,
    \Tile_X3Y1_W2BEG[3] ,
    \Tile_X3Y1_W2BEG[2] ,
    \Tile_X3Y1_W2BEG[1] ,
    \Tile_X3Y1_W2BEG[0] }),
    .W6BEG({\Tile_X2Y1_W6BEG[11] ,
    \Tile_X2Y1_W6BEG[10] ,
    \Tile_X2Y1_W6BEG[9] ,
    \Tile_X2Y1_W6BEG[8] ,
    \Tile_X2Y1_W6BEG[7] ,
    \Tile_X2Y1_W6BEG[6] ,
    \Tile_X2Y1_W6BEG[5] ,
    \Tile_X2Y1_W6BEG[4] ,
    \Tile_X2Y1_W6BEG[3] ,
    \Tile_X2Y1_W6BEG[2] ,
    \Tile_X2Y1_W6BEG[1] ,
    \Tile_X2Y1_W6BEG[0] }),
    .W6END({\Tile_X3Y1_W6BEG[11] ,
    \Tile_X3Y1_W6BEG[10] ,
    \Tile_X3Y1_W6BEG[9] ,
    \Tile_X3Y1_W6BEG[8] ,
    \Tile_X3Y1_W6BEG[7] ,
    \Tile_X3Y1_W6BEG[6] ,
    \Tile_X3Y1_W6BEG[5] ,
    \Tile_X3Y1_W6BEG[4] ,
    \Tile_X3Y1_W6BEG[3] ,
    \Tile_X3Y1_W6BEG[2] ,
    \Tile_X3Y1_W6BEG[1] ,
    \Tile_X3Y1_W6BEG[0] }),
    .WW4BEG({\Tile_X2Y1_WW4BEG[15] ,
    \Tile_X2Y1_WW4BEG[14] ,
    \Tile_X2Y1_WW4BEG[13] ,
    \Tile_X2Y1_WW4BEG[12] ,
    \Tile_X2Y1_WW4BEG[11] ,
    \Tile_X2Y1_WW4BEG[10] ,
    \Tile_X2Y1_WW4BEG[9] ,
    \Tile_X2Y1_WW4BEG[8] ,
    \Tile_X2Y1_WW4BEG[7] ,
    \Tile_X2Y1_WW4BEG[6] ,
    \Tile_X2Y1_WW4BEG[5] ,
    \Tile_X2Y1_WW4BEG[4] ,
    \Tile_X2Y1_WW4BEG[3] ,
    \Tile_X2Y1_WW4BEG[2] ,
    \Tile_X2Y1_WW4BEG[1] ,
    \Tile_X2Y1_WW4BEG[0] }),
    .WW4END({\Tile_X3Y1_WW4BEG[15] ,
    \Tile_X3Y1_WW4BEG[14] ,
    \Tile_X3Y1_WW4BEG[13] ,
    \Tile_X3Y1_WW4BEG[12] ,
    \Tile_X3Y1_WW4BEG[11] ,
    \Tile_X3Y1_WW4BEG[10] ,
    \Tile_X3Y1_WW4BEG[9] ,
    \Tile_X3Y1_WW4BEG[8] ,
    \Tile_X3Y1_WW4BEG[7] ,
    \Tile_X3Y1_WW4BEG[6] ,
    \Tile_X3Y1_WW4BEG[5] ,
    \Tile_X3Y1_WW4BEG[4] ,
    \Tile_X3Y1_WW4BEG[3] ,
    \Tile_X3Y1_WW4BEG[2] ,
    \Tile_X3Y1_WW4BEG[1] ,
    \Tile_X3Y1_WW4BEG[0] }));
 LUT4AB Tile_X2Y2_LUT4AB (.Ci(Tile_X2Y3_Co),
    .Co(Tile_X2Y2_Co),
    .UserCLK(Tile_X2Y3_UserCLKo),
    .UserCLKo(Tile_X2Y2_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X2Y2_E1BEG[3] ,
    \Tile_X2Y2_E1BEG[2] ,
    \Tile_X2Y2_E1BEG[1] ,
    \Tile_X2Y2_E1BEG[0] }),
    .E1END({\Tile_X1Y2_E1BEG[3] ,
    \Tile_X1Y2_E1BEG[2] ,
    \Tile_X1Y2_E1BEG[1] ,
    \Tile_X1Y2_E1BEG[0] }),
    .E2BEG({\Tile_X2Y2_E2BEG[7] ,
    \Tile_X2Y2_E2BEG[6] ,
    \Tile_X2Y2_E2BEG[5] ,
    \Tile_X2Y2_E2BEG[4] ,
    \Tile_X2Y2_E2BEG[3] ,
    \Tile_X2Y2_E2BEG[2] ,
    \Tile_X2Y2_E2BEG[1] ,
    \Tile_X2Y2_E2BEG[0] }),
    .E2BEGb({\Tile_X2Y2_E2BEGb[7] ,
    \Tile_X2Y2_E2BEGb[6] ,
    \Tile_X2Y2_E2BEGb[5] ,
    \Tile_X2Y2_E2BEGb[4] ,
    \Tile_X2Y2_E2BEGb[3] ,
    \Tile_X2Y2_E2BEGb[2] ,
    \Tile_X2Y2_E2BEGb[1] ,
    \Tile_X2Y2_E2BEGb[0] }),
    .E2END({\Tile_X1Y2_E2BEGb[7] ,
    \Tile_X1Y2_E2BEGb[6] ,
    \Tile_X1Y2_E2BEGb[5] ,
    \Tile_X1Y2_E2BEGb[4] ,
    \Tile_X1Y2_E2BEGb[3] ,
    \Tile_X1Y2_E2BEGb[2] ,
    \Tile_X1Y2_E2BEGb[1] ,
    \Tile_X1Y2_E2BEGb[0] }),
    .E2MID({\Tile_X1Y2_E2BEG[7] ,
    \Tile_X1Y2_E2BEG[6] ,
    \Tile_X1Y2_E2BEG[5] ,
    \Tile_X1Y2_E2BEG[4] ,
    \Tile_X1Y2_E2BEG[3] ,
    \Tile_X1Y2_E2BEG[2] ,
    \Tile_X1Y2_E2BEG[1] ,
    \Tile_X1Y2_E2BEG[0] }),
    .E6BEG({\Tile_X2Y2_E6BEG[11] ,
    \Tile_X2Y2_E6BEG[10] ,
    \Tile_X2Y2_E6BEG[9] ,
    \Tile_X2Y2_E6BEG[8] ,
    \Tile_X2Y2_E6BEG[7] ,
    \Tile_X2Y2_E6BEG[6] ,
    \Tile_X2Y2_E6BEG[5] ,
    \Tile_X2Y2_E6BEG[4] ,
    \Tile_X2Y2_E6BEG[3] ,
    \Tile_X2Y2_E6BEG[2] ,
    \Tile_X2Y2_E6BEG[1] ,
    \Tile_X2Y2_E6BEG[0] }),
    .E6END({\Tile_X1Y2_E6BEG[11] ,
    \Tile_X1Y2_E6BEG[10] ,
    \Tile_X1Y2_E6BEG[9] ,
    \Tile_X1Y2_E6BEG[8] ,
    \Tile_X1Y2_E6BEG[7] ,
    \Tile_X1Y2_E6BEG[6] ,
    \Tile_X1Y2_E6BEG[5] ,
    \Tile_X1Y2_E6BEG[4] ,
    \Tile_X1Y2_E6BEG[3] ,
    \Tile_X1Y2_E6BEG[2] ,
    \Tile_X1Y2_E6BEG[1] ,
    \Tile_X1Y2_E6BEG[0] }),
    .EE4BEG({\Tile_X2Y2_EE4BEG[15] ,
    \Tile_X2Y2_EE4BEG[14] ,
    \Tile_X2Y2_EE4BEG[13] ,
    \Tile_X2Y2_EE4BEG[12] ,
    \Tile_X2Y2_EE4BEG[11] ,
    \Tile_X2Y2_EE4BEG[10] ,
    \Tile_X2Y2_EE4BEG[9] ,
    \Tile_X2Y2_EE4BEG[8] ,
    \Tile_X2Y2_EE4BEG[7] ,
    \Tile_X2Y2_EE4BEG[6] ,
    \Tile_X2Y2_EE4BEG[5] ,
    \Tile_X2Y2_EE4BEG[4] ,
    \Tile_X2Y2_EE4BEG[3] ,
    \Tile_X2Y2_EE4BEG[2] ,
    \Tile_X2Y2_EE4BEG[1] ,
    \Tile_X2Y2_EE4BEG[0] }),
    .EE4END({\Tile_X1Y2_EE4BEG[15] ,
    \Tile_X1Y2_EE4BEG[14] ,
    \Tile_X1Y2_EE4BEG[13] ,
    \Tile_X1Y2_EE4BEG[12] ,
    \Tile_X1Y2_EE4BEG[11] ,
    \Tile_X1Y2_EE4BEG[10] ,
    \Tile_X1Y2_EE4BEG[9] ,
    \Tile_X1Y2_EE4BEG[8] ,
    \Tile_X1Y2_EE4BEG[7] ,
    \Tile_X1Y2_EE4BEG[6] ,
    \Tile_X1Y2_EE4BEG[5] ,
    \Tile_X1Y2_EE4BEG[4] ,
    \Tile_X1Y2_EE4BEG[3] ,
    \Tile_X1Y2_EE4BEG[2] ,
    \Tile_X1Y2_EE4BEG[1] ,
    \Tile_X1Y2_EE4BEG[0] }),
    .FrameData({\Tile_X1Y2_FrameData_O[31] ,
    \Tile_X1Y2_FrameData_O[30] ,
    \Tile_X1Y2_FrameData_O[29] ,
    \Tile_X1Y2_FrameData_O[28] ,
    \Tile_X1Y2_FrameData_O[27] ,
    \Tile_X1Y2_FrameData_O[26] ,
    \Tile_X1Y2_FrameData_O[25] ,
    \Tile_X1Y2_FrameData_O[24] ,
    \Tile_X1Y2_FrameData_O[23] ,
    \Tile_X1Y2_FrameData_O[22] ,
    \Tile_X1Y2_FrameData_O[21] ,
    \Tile_X1Y2_FrameData_O[20] ,
    \Tile_X1Y2_FrameData_O[19] ,
    \Tile_X1Y2_FrameData_O[18] ,
    \Tile_X1Y2_FrameData_O[17] ,
    \Tile_X1Y2_FrameData_O[16] ,
    \Tile_X1Y2_FrameData_O[15] ,
    \Tile_X1Y2_FrameData_O[14] ,
    \Tile_X1Y2_FrameData_O[13] ,
    \Tile_X1Y2_FrameData_O[12] ,
    \Tile_X1Y2_FrameData_O[11] ,
    \Tile_X1Y2_FrameData_O[10] ,
    \Tile_X1Y2_FrameData_O[9] ,
    \Tile_X1Y2_FrameData_O[8] ,
    \Tile_X1Y2_FrameData_O[7] ,
    \Tile_X1Y2_FrameData_O[6] ,
    \Tile_X1Y2_FrameData_O[5] ,
    \Tile_X1Y2_FrameData_O[4] ,
    \Tile_X1Y2_FrameData_O[3] ,
    \Tile_X1Y2_FrameData_O[2] ,
    \Tile_X1Y2_FrameData_O[1] ,
    \Tile_X1Y2_FrameData_O[0] }),
    .FrameData_O({\Tile_X2Y2_FrameData_O[31] ,
    \Tile_X2Y2_FrameData_O[30] ,
    \Tile_X2Y2_FrameData_O[29] ,
    \Tile_X2Y2_FrameData_O[28] ,
    \Tile_X2Y2_FrameData_O[27] ,
    \Tile_X2Y2_FrameData_O[26] ,
    \Tile_X2Y2_FrameData_O[25] ,
    \Tile_X2Y2_FrameData_O[24] ,
    \Tile_X2Y2_FrameData_O[23] ,
    \Tile_X2Y2_FrameData_O[22] ,
    \Tile_X2Y2_FrameData_O[21] ,
    \Tile_X2Y2_FrameData_O[20] ,
    \Tile_X2Y2_FrameData_O[19] ,
    \Tile_X2Y2_FrameData_O[18] ,
    \Tile_X2Y2_FrameData_O[17] ,
    \Tile_X2Y2_FrameData_O[16] ,
    \Tile_X2Y2_FrameData_O[15] ,
    \Tile_X2Y2_FrameData_O[14] ,
    \Tile_X2Y2_FrameData_O[13] ,
    \Tile_X2Y2_FrameData_O[12] ,
    \Tile_X2Y2_FrameData_O[11] ,
    \Tile_X2Y2_FrameData_O[10] ,
    \Tile_X2Y2_FrameData_O[9] ,
    \Tile_X2Y2_FrameData_O[8] ,
    \Tile_X2Y2_FrameData_O[7] ,
    \Tile_X2Y2_FrameData_O[6] ,
    \Tile_X2Y2_FrameData_O[5] ,
    \Tile_X2Y2_FrameData_O[4] ,
    \Tile_X2Y2_FrameData_O[3] ,
    \Tile_X2Y2_FrameData_O[2] ,
    \Tile_X2Y2_FrameData_O[1] ,
    \Tile_X2Y2_FrameData_O[0] }),
    .FrameStrobe({\Tile_X2Y3_FrameStrobe_O[19] ,
    \Tile_X2Y3_FrameStrobe_O[18] ,
    \Tile_X2Y3_FrameStrobe_O[17] ,
    \Tile_X2Y3_FrameStrobe_O[16] ,
    \Tile_X2Y3_FrameStrobe_O[15] ,
    \Tile_X2Y3_FrameStrobe_O[14] ,
    \Tile_X2Y3_FrameStrobe_O[13] ,
    \Tile_X2Y3_FrameStrobe_O[12] ,
    \Tile_X2Y3_FrameStrobe_O[11] ,
    \Tile_X2Y3_FrameStrobe_O[10] ,
    \Tile_X2Y3_FrameStrobe_O[9] ,
    \Tile_X2Y3_FrameStrobe_O[8] ,
    \Tile_X2Y3_FrameStrobe_O[7] ,
    \Tile_X2Y3_FrameStrobe_O[6] ,
    \Tile_X2Y3_FrameStrobe_O[5] ,
    \Tile_X2Y3_FrameStrobe_O[4] ,
    \Tile_X2Y3_FrameStrobe_O[3] ,
    \Tile_X2Y3_FrameStrobe_O[2] ,
    \Tile_X2Y3_FrameStrobe_O[1] ,
    \Tile_X2Y3_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X2Y2_FrameStrobe_O[19] ,
    \Tile_X2Y2_FrameStrobe_O[18] ,
    \Tile_X2Y2_FrameStrobe_O[17] ,
    \Tile_X2Y2_FrameStrobe_O[16] ,
    \Tile_X2Y2_FrameStrobe_O[15] ,
    \Tile_X2Y2_FrameStrobe_O[14] ,
    \Tile_X2Y2_FrameStrobe_O[13] ,
    \Tile_X2Y2_FrameStrobe_O[12] ,
    \Tile_X2Y2_FrameStrobe_O[11] ,
    \Tile_X2Y2_FrameStrobe_O[10] ,
    \Tile_X2Y2_FrameStrobe_O[9] ,
    \Tile_X2Y2_FrameStrobe_O[8] ,
    \Tile_X2Y2_FrameStrobe_O[7] ,
    \Tile_X2Y2_FrameStrobe_O[6] ,
    \Tile_X2Y2_FrameStrobe_O[5] ,
    \Tile_X2Y2_FrameStrobe_O[4] ,
    \Tile_X2Y2_FrameStrobe_O[3] ,
    \Tile_X2Y2_FrameStrobe_O[2] ,
    \Tile_X2Y2_FrameStrobe_O[1] ,
    \Tile_X2Y2_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X2Y2_N1BEG[3] ,
    \Tile_X2Y2_N1BEG[2] ,
    \Tile_X2Y2_N1BEG[1] ,
    \Tile_X2Y2_N1BEG[0] }),
    .N1END({\Tile_X2Y3_N1BEG[3] ,
    \Tile_X2Y3_N1BEG[2] ,
    \Tile_X2Y3_N1BEG[1] ,
    \Tile_X2Y3_N1BEG[0] }),
    .N2BEG({\Tile_X2Y2_N2BEG[7] ,
    \Tile_X2Y2_N2BEG[6] ,
    \Tile_X2Y2_N2BEG[5] ,
    \Tile_X2Y2_N2BEG[4] ,
    \Tile_X2Y2_N2BEG[3] ,
    \Tile_X2Y2_N2BEG[2] ,
    \Tile_X2Y2_N2BEG[1] ,
    \Tile_X2Y2_N2BEG[0] }),
    .N2BEGb({\Tile_X2Y2_N2BEGb[7] ,
    \Tile_X2Y2_N2BEGb[6] ,
    \Tile_X2Y2_N2BEGb[5] ,
    \Tile_X2Y2_N2BEGb[4] ,
    \Tile_X2Y2_N2BEGb[3] ,
    \Tile_X2Y2_N2BEGb[2] ,
    \Tile_X2Y2_N2BEGb[1] ,
    \Tile_X2Y2_N2BEGb[0] }),
    .N2END({\Tile_X2Y3_N2BEGb[7] ,
    \Tile_X2Y3_N2BEGb[6] ,
    \Tile_X2Y3_N2BEGb[5] ,
    \Tile_X2Y3_N2BEGb[4] ,
    \Tile_X2Y3_N2BEGb[3] ,
    \Tile_X2Y3_N2BEGb[2] ,
    \Tile_X2Y3_N2BEGb[1] ,
    \Tile_X2Y3_N2BEGb[0] }),
    .N2MID({\Tile_X2Y3_N2BEG[7] ,
    \Tile_X2Y3_N2BEG[6] ,
    \Tile_X2Y3_N2BEG[5] ,
    \Tile_X2Y3_N2BEG[4] ,
    \Tile_X2Y3_N2BEG[3] ,
    \Tile_X2Y3_N2BEG[2] ,
    \Tile_X2Y3_N2BEG[1] ,
    \Tile_X2Y3_N2BEG[0] }),
    .N4BEG({\Tile_X2Y2_N4BEG[15] ,
    \Tile_X2Y2_N4BEG[14] ,
    \Tile_X2Y2_N4BEG[13] ,
    \Tile_X2Y2_N4BEG[12] ,
    \Tile_X2Y2_N4BEG[11] ,
    \Tile_X2Y2_N4BEG[10] ,
    \Tile_X2Y2_N4BEG[9] ,
    \Tile_X2Y2_N4BEG[8] ,
    \Tile_X2Y2_N4BEG[7] ,
    \Tile_X2Y2_N4BEG[6] ,
    \Tile_X2Y2_N4BEG[5] ,
    \Tile_X2Y2_N4BEG[4] ,
    \Tile_X2Y2_N4BEG[3] ,
    \Tile_X2Y2_N4BEG[2] ,
    \Tile_X2Y2_N4BEG[1] ,
    \Tile_X2Y2_N4BEG[0] }),
    .N4END({\Tile_X2Y3_N4BEG[15] ,
    \Tile_X2Y3_N4BEG[14] ,
    \Tile_X2Y3_N4BEG[13] ,
    \Tile_X2Y3_N4BEG[12] ,
    \Tile_X2Y3_N4BEG[11] ,
    \Tile_X2Y3_N4BEG[10] ,
    \Tile_X2Y3_N4BEG[9] ,
    \Tile_X2Y3_N4BEG[8] ,
    \Tile_X2Y3_N4BEG[7] ,
    \Tile_X2Y3_N4BEG[6] ,
    \Tile_X2Y3_N4BEG[5] ,
    \Tile_X2Y3_N4BEG[4] ,
    \Tile_X2Y3_N4BEG[3] ,
    \Tile_X2Y3_N4BEG[2] ,
    \Tile_X2Y3_N4BEG[1] ,
    \Tile_X2Y3_N4BEG[0] }),
    .NN4BEG({\Tile_X2Y2_NN4BEG[15] ,
    \Tile_X2Y2_NN4BEG[14] ,
    \Tile_X2Y2_NN4BEG[13] ,
    \Tile_X2Y2_NN4BEG[12] ,
    \Tile_X2Y2_NN4BEG[11] ,
    \Tile_X2Y2_NN4BEG[10] ,
    \Tile_X2Y2_NN4BEG[9] ,
    \Tile_X2Y2_NN4BEG[8] ,
    \Tile_X2Y2_NN4BEG[7] ,
    \Tile_X2Y2_NN4BEG[6] ,
    \Tile_X2Y2_NN4BEG[5] ,
    \Tile_X2Y2_NN4BEG[4] ,
    \Tile_X2Y2_NN4BEG[3] ,
    \Tile_X2Y2_NN4BEG[2] ,
    \Tile_X2Y2_NN4BEG[1] ,
    \Tile_X2Y2_NN4BEG[0] }),
    .NN4END({\Tile_X2Y3_NN4BEG[15] ,
    \Tile_X2Y3_NN4BEG[14] ,
    \Tile_X2Y3_NN4BEG[13] ,
    \Tile_X2Y3_NN4BEG[12] ,
    \Tile_X2Y3_NN4BEG[11] ,
    \Tile_X2Y3_NN4BEG[10] ,
    \Tile_X2Y3_NN4BEG[9] ,
    \Tile_X2Y3_NN4BEG[8] ,
    \Tile_X2Y3_NN4BEG[7] ,
    \Tile_X2Y3_NN4BEG[6] ,
    \Tile_X2Y3_NN4BEG[5] ,
    \Tile_X2Y3_NN4BEG[4] ,
    \Tile_X2Y3_NN4BEG[3] ,
    \Tile_X2Y3_NN4BEG[2] ,
    \Tile_X2Y3_NN4BEG[1] ,
    \Tile_X2Y3_NN4BEG[0] }),
    .S1BEG({\Tile_X2Y2_S1BEG[3] ,
    \Tile_X2Y2_S1BEG[2] ,
    \Tile_X2Y2_S1BEG[1] ,
    \Tile_X2Y2_S1BEG[0] }),
    .S1END({\Tile_X2Y1_S1BEG[3] ,
    \Tile_X2Y1_S1BEG[2] ,
    \Tile_X2Y1_S1BEG[1] ,
    \Tile_X2Y1_S1BEG[0] }),
    .S2BEG({\Tile_X2Y2_S2BEG[7] ,
    \Tile_X2Y2_S2BEG[6] ,
    \Tile_X2Y2_S2BEG[5] ,
    \Tile_X2Y2_S2BEG[4] ,
    \Tile_X2Y2_S2BEG[3] ,
    \Tile_X2Y2_S2BEG[2] ,
    \Tile_X2Y2_S2BEG[1] ,
    \Tile_X2Y2_S2BEG[0] }),
    .S2BEGb({\Tile_X2Y2_S2BEGb[7] ,
    \Tile_X2Y2_S2BEGb[6] ,
    \Tile_X2Y2_S2BEGb[5] ,
    \Tile_X2Y2_S2BEGb[4] ,
    \Tile_X2Y2_S2BEGb[3] ,
    \Tile_X2Y2_S2BEGb[2] ,
    \Tile_X2Y2_S2BEGb[1] ,
    \Tile_X2Y2_S2BEGb[0] }),
    .S2END({\Tile_X2Y1_S2BEGb[7] ,
    \Tile_X2Y1_S2BEGb[6] ,
    \Tile_X2Y1_S2BEGb[5] ,
    \Tile_X2Y1_S2BEGb[4] ,
    \Tile_X2Y1_S2BEGb[3] ,
    \Tile_X2Y1_S2BEGb[2] ,
    \Tile_X2Y1_S2BEGb[1] ,
    \Tile_X2Y1_S2BEGb[0] }),
    .S2MID({\Tile_X2Y1_S2BEG[7] ,
    \Tile_X2Y1_S2BEG[6] ,
    \Tile_X2Y1_S2BEG[5] ,
    \Tile_X2Y1_S2BEG[4] ,
    \Tile_X2Y1_S2BEG[3] ,
    \Tile_X2Y1_S2BEG[2] ,
    \Tile_X2Y1_S2BEG[1] ,
    \Tile_X2Y1_S2BEG[0] }),
    .S4BEG({\Tile_X2Y2_S4BEG[15] ,
    \Tile_X2Y2_S4BEG[14] ,
    \Tile_X2Y2_S4BEG[13] ,
    \Tile_X2Y2_S4BEG[12] ,
    \Tile_X2Y2_S4BEG[11] ,
    \Tile_X2Y2_S4BEG[10] ,
    \Tile_X2Y2_S4BEG[9] ,
    \Tile_X2Y2_S4BEG[8] ,
    \Tile_X2Y2_S4BEG[7] ,
    \Tile_X2Y2_S4BEG[6] ,
    \Tile_X2Y2_S4BEG[5] ,
    \Tile_X2Y2_S4BEG[4] ,
    \Tile_X2Y2_S4BEG[3] ,
    \Tile_X2Y2_S4BEG[2] ,
    \Tile_X2Y2_S4BEG[1] ,
    \Tile_X2Y2_S4BEG[0] }),
    .S4END({\Tile_X2Y1_S4BEG[15] ,
    \Tile_X2Y1_S4BEG[14] ,
    \Tile_X2Y1_S4BEG[13] ,
    \Tile_X2Y1_S4BEG[12] ,
    \Tile_X2Y1_S4BEG[11] ,
    \Tile_X2Y1_S4BEG[10] ,
    \Tile_X2Y1_S4BEG[9] ,
    \Tile_X2Y1_S4BEG[8] ,
    \Tile_X2Y1_S4BEG[7] ,
    \Tile_X2Y1_S4BEG[6] ,
    \Tile_X2Y1_S4BEG[5] ,
    \Tile_X2Y1_S4BEG[4] ,
    \Tile_X2Y1_S4BEG[3] ,
    \Tile_X2Y1_S4BEG[2] ,
    \Tile_X2Y1_S4BEG[1] ,
    \Tile_X2Y1_S4BEG[0] }),
    .SS4BEG({\Tile_X2Y2_SS4BEG[15] ,
    \Tile_X2Y2_SS4BEG[14] ,
    \Tile_X2Y2_SS4BEG[13] ,
    \Tile_X2Y2_SS4BEG[12] ,
    \Tile_X2Y2_SS4BEG[11] ,
    \Tile_X2Y2_SS4BEG[10] ,
    \Tile_X2Y2_SS4BEG[9] ,
    \Tile_X2Y2_SS4BEG[8] ,
    \Tile_X2Y2_SS4BEG[7] ,
    \Tile_X2Y2_SS4BEG[6] ,
    \Tile_X2Y2_SS4BEG[5] ,
    \Tile_X2Y2_SS4BEG[4] ,
    \Tile_X2Y2_SS4BEG[3] ,
    \Tile_X2Y2_SS4BEG[2] ,
    \Tile_X2Y2_SS4BEG[1] ,
    \Tile_X2Y2_SS4BEG[0] }),
    .SS4END({\Tile_X2Y1_SS4BEG[15] ,
    \Tile_X2Y1_SS4BEG[14] ,
    \Tile_X2Y1_SS4BEG[13] ,
    \Tile_X2Y1_SS4BEG[12] ,
    \Tile_X2Y1_SS4BEG[11] ,
    \Tile_X2Y1_SS4BEG[10] ,
    \Tile_X2Y1_SS4BEG[9] ,
    \Tile_X2Y1_SS4BEG[8] ,
    \Tile_X2Y1_SS4BEG[7] ,
    \Tile_X2Y1_SS4BEG[6] ,
    \Tile_X2Y1_SS4BEG[5] ,
    \Tile_X2Y1_SS4BEG[4] ,
    \Tile_X2Y1_SS4BEG[3] ,
    \Tile_X2Y1_SS4BEG[2] ,
    \Tile_X2Y1_SS4BEG[1] ,
    \Tile_X2Y1_SS4BEG[0] }),
    .W1BEG({\Tile_X2Y2_W1BEG[3] ,
    \Tile_X2Y2_W1BEG[2] ,
    \Tile_X2Y2_W1BEG[1] ,
    \Tile_X2Y2_W1BEG[0] }),
    .W1END({\Tile_X3Y2_W1BEG[3] ,
    \Tile_X3Y2_W1BEG[2] ,
    \Tile_X3Y2_W1BEG[1] ,
    \Tile_X3Y2_W1BEG[0] }),
    .W2BEG({\Tile_X2Y2_W2BEG[7] ,
    \Tile_X2Y2_W2BEG[6] ,
    \Tile_X2Y2_W2BEG[5] ,
    \Tile_X2Y2_W2BEG[4] ,
    \Tile_X2Y2_W2BEG[3] ,
    \Tile_X2Y2_W2BEG[2] ,
    \Tile_X2Y2_W2BEG[1] ,
    \Tile_X2Y2_W2BEG[0] }),
    .W2BEGb({\Tile_X2Y2_W2BEGb[7] ,
    \Tile_X2Y2_W2BEGb[6] ,
    \Tile_X2Y2_W2BEGb[5] ,
    \Tile_X2Y2_W2BEGb[4] ,
    \Tile_X2Y2_W2BEGb[3] ,
    \Tile_X2Y2_W2BEGb[2] ,
    \Tile_X2Y2_W2BEGb[1] ,
    \Tile_X2Y2_W2BEGb[0] }),
    .W2END({\Tile_X3Y2_W2BEGb[7] ,
    \Tile_X3Y2_W2BEGb[6] ,
    \Tile_X3Y2_W2BEGb[5] ,
    \Tile_X3Y2_W2BEGb[4] ,
    \Tile_X3Y2_W2BEGb[3] ,
    \Tile_X3Y2_W2BEGb[2] ,
    \Tile_X3Y2_W2BEGb[1] ,
    \Tile_X3Y2_W2BEGb[0] }),
    .W2MID({\Tile_X3Y2_W2BEG[7] ,
    \Tile_X3Y2_W2BEG[6] ,
    \Tile_X3Y2_W2BEG[5] ,
    \Tile_X3Y2_W2BEG[4] ,
    \Tile_X3Y2_W2BEG[3] ,
    \Tile_X3Y2_W2BEG[2] ,
    \Tile_X3Y2_W2BEG[1] ,
    \Tile_X3Y2_W2BEG[0] }),
    .W6BEG({\Tile_X2Y2_W6BEG[11] ,
    \Tile_X2Y2_W6BEG[10] ,
    \Tile_X2Y2_W6BEG[9] ,
    \Tile_X2Y2_W6BEG[8] ,
    \Tile_X2Y2_W6BEG[7] ,
    \Tile_X2Y2_W6BEG[6] ,
    \Tile_X2Y2_W6BEG[5] ,
    \Tile_X2Y2_W6BEG[4] ,
    \Tile_X2Y2_W6BEG[3] ,
    \Tile_X2Y2_W6BEG[2] ,
    \Tile_X2Y2_W6BEG[1] ,
    \Tile_X2Y2_W6BEG[0] }),
    .W6END({\Tile_X3Y2_W6BEG[11] ,
    \Tile_X3Y2_W6BEG[10] ,
    \Tile_X3Y2_W6BEG[9] ,
    \Tile_X3Y2_W6BEG[8] ,
    \Tile_X3Y2_W6BEG[7] ,
    \Tile_X3Y2_W6BEG[6] ,
    \Tile_X3Y2_W6BEG[5] ,
    \Tile_X3Y2_W6BEG[4] ,
    \Tile_X3Y2_W6BEG[3] ,
    \Tile_X3Y2_W6BEG[2] ,
    \Tile_X3Y2_W6BEG[1] ,
    \Tile_X3Y2_W6BEG[0] }),
    .WW4BEG({\Tile_X2Y2_WW4BEG[15] ,
    \Tile_X2Y2_WW4BEG[14] ,
    \Tile_X2Y2_WW4BEG[13] ,
    \Tile_X2Y2_WW4BEG[12] ,
    \Tile_X2Y2_WW4BEG[11] ,
    \Tile_X2Y2_WW4BEG[10] ,
    \Tile_X2Y2_WW4BEG[9] ,
    \Tile_X2Y2_WW4BEG[8] ,
    \Tile_X2Y2_WW4BEG[7] ,
    \Tile_X2Y2_WW4BEG[6] ,
    \Tile_X2Y2_WW4BEG[5] ,
    \Tile_X2Y2_WW4BEG[4] ,
    \Tile_X2Y2_WW4BEG[3] ,
    \Tile_X2Y2_WW4BEG[2] ,
    \Tile_X2Y2_WW4BEG[1] ,
    \Tile_X2Y2_WW4BEG[0] }),
    .WW4END({\Tile_X3Y2_WW4BEG[15] ,
    \Tile_X3Y2_WW4BEG[14] ,
    \Tile_X3Y2_WW4BEG[13] ,
    \Tile_X3Y2_WW4BEG[12] ,
    \Tile_X3Y2_WW4BEG[11] ,
    \Tile_X3Y2_WW4BEG[10] ,
    \Tile_X3Y2_WW4BEG[9] ,
    \Tile_X3Y2_WW4BEG[8] ,
    \Tile_X3Y2_WW4BEG[7] ,
    \Tile_X3Y2_WW4BEG[6] ,
    \Tile_X3Y2_WW4BEG[5] ,
    \Tile_X3Y2_WW4BEG[4] ,
    \Tile_X3Y2_WW4BEG[3] ,
    \Tile_X3Y2_WW4BEG[2] ,
    \Tile_X3Y2_WW4BEG[1] ,
    \Tile_X3Y2_WW4BEG[0] }));
 LUT4AB Tile_X2Y3_LUT4AB (.Ci(Tile_X2Y4_Co),
    .Co(Tile_X2Y3_Co),
    .UserCLK(Tile_X2Y4_UserCLKo),
    .UserCLKo(Tile_X2Y3_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X2Y3_E1BEG[3] ,
    \Tile_X2Y3_E1BEG[2] ,
    \Tile_X2Y3_E1BEG[1] ,
    \Tile_X2Y3_E1BEG[0] }),
    .E1END({\Tile_X1Y3_E1BEG[3] ,
    \Tile_X1Y3_E1BEG[2] ,
    \Tile_X1Y3_E1BEG[1] ,
    \Tile_X1Y3_E1BEG[0] }),
    .E2BEG({\Tile_X2Y3_E2BEG[7] ,
    \Tile_X2Y3_E2BEG[6] ,
    \Tile_X2Y3_E2BEG[5] ,
    \Tile_X2Y3_E2BEG[4] ,
    \Tile_X2Y3_E2BEG[3] ,
    \Tile_X2Y3_E2BEG[2] ,
    \Tile_X2Y3_E2BEG[1] ,
    \Tile_X2Y3_E2BEG[0] }),
    .E2BEGb({\Tile_X2Y3_E2BEGb[7] ,
    \Tile_X2Y3_E2BEGb[6] ,
    \Tile_X2Y3_E2BEGb[5] ,
    \Tile_X2Y3_E2BEGb[4] ,
    \Tile_X2Y3_E2BEGb[3] ,
    \Tile_X2Y3_E2BEGb[2] ,
    \Tile_X2Y3_E2BEGb[1] ,
    \Tile_X2Y3_E2BEGb[0] }),
    .E2END({\Tile_X1Y3_E2BEGb[7] ,
    \Tile_X1Y3_E2BEGb[6] ,
    \Tile_X1Y3_E2BEGb[5] ,
    \Tile_X1Y3_E2BEGb[4] ,
    \Tile_X1Y3_E2BEGb[3] ,
    \Tile_X1Y3_E2BEGb[2] ,
    \Tile_X1Y3_E2BEGb[1] ,
    \Tile_X1Y3_E2BEGb[0] }),
    .E2MID({\Tile_X1Y3_E2BEG[7] ,
    \Tile_X1Y3_E2BEG[6] ,
    \Tile_X1Y3_E2BEG[5] ,
    \Tile_X1Y3_E2BEG[4] ,
    \Tile_X1Y3_E2BEG[3] ,
    \Tile_X1Y3_E2BEG[2] ,
    \Tile_X1Y3_E2BEG[1] ,
    \Tile_X1Y3_E2BEG[0] }),
    .E6BEG({\Tile_X2Y3_E6BEG[11] ,
    \Tile_X2Y3_E6BEG[10] ,
    \Tile_X2Y3_E6BEG[9] ,
    \Tile_X2Y3_E6BEG[8] ,
    \Tile_X2Y3_E6BEG[7] ,
    \Tile_X2Y3_E6BEG[6] ,
    \Tile_X2Y3_E6BEG[5] ,
    \Tile_X2Y3_E6BEG[4] ,
    \Tile_X2Y3_E6BEG[3] ,
    \Tile_X2Y3_E6BEG[2] ,
    \Tile_X2Y3_E6BEG[1] ,
    \Tile_X2Y3_E6BEG[0] }),
    .E6END({\Tile_X1Y3_E6BEG[11] ,
    \Tile_X1Y3_E6BEG[10] ,
    \Tile_X1Y3_E6BEG[9] ,
    \Tile_X1Y3_E6BEG[8] ,
    \Tile_X1Y3_E6BEG[7] ,
    \Tile_X1Y3_E6BEG[6] ,
    \Tile_X1Y3_E6BEG[5] ,
    \Tile_X1Y3_E6BEG[4] ,
    \Tile_X1Y3_E6BEG[3] ,
    \Tile_X1Y3_E6BEG[2] ,
    \Tile_X1Y3_E6BEG[1] ,
    \Tile_X1Y3_E6BEG[0] }),
    .EE4BEG({\Tile_X2Y3_EE4BEG[15] ,
    \Tile_X2Y3_EE4BEG[14] ,
    \Tile_X2Y3_EE4BEG[13] ,
    \Tile_X2Y3_EE4BEG[12] ,
    \Tile_X2Y3_EE4BEG[11] ,
    \Tile_X2Y3_EE4BEG[10] ,
    \Tile_X2Y3_EE4BEG[9] ,
    \Tile_X2Y3_EE4BEG[8] ,
    \Tile_X2Y3_EE4BEG[7] ,
    \Tile_X2Y3_EE4BEG[6] ,
    \Tile_X2Y3_EE4BEG[5] ,
    \Tile_X2Y3_EE4BEG[4] ,
    \Tile_X2Y3_EE4BEG[3] ,
    \Tile_X2Y3_EE4BEG[2] ,
    \Tile_X2Y3_EE4BEG[1] ,
    \Tile_X2Y3_EE4BEG[0] }),
    .EE4END({\Tile_X1Y3_EE4BEG[15] ,
    \Tile_X1Y3_EE4BEG[14] ,
    \Tile_X1Y3_EE4BEG[13] ,
    \Tile_X1Y3_EE4BEG[12] ,
    \Tile_X1Y3_EE4BEG[11] ,
    \Tile_X1Y3_EE4BEG[10] ,
    \Tile_X1Y3_EE4BEG[9] ,
    \Tile_X1Y3_EE4BEG[8] ,
    \Tile_X1Y3_EE4BEG[7] ,
    \Tile_X1Y3_EE4BEG[6] ,
    \Tile_X1Y3_EE4BEG[5] ,
    \Tile_X1Y3_EE4BEG[4] ,
    \Tile_X1Y3_EE4BEG[3] ,
    \Tile_X1Y3_EE4BEG[2] ,
    \Tile_X1Y3_EE4BEG[1] ,
    \Tile_X1Y3_EE4BEG[0] }),
    .FrameData({\Tile_X1Y3_FrameData_O[31] ,
    \Tile_X1Y3_FrameData_O[30] ,
    \Tile_X1Y3_FrameData_O[29] ,
    \Tile_X1Y3_FrameData_O[28] ,
    \Tile_X1Y3_FrameData_O[27] ,
    \Tile_X1Y3_FrameData_O[26] ,
    \Tile_X1Y3_FrameData_O[25] ,
    \Tile_X1Y3_FrameData_O[24] ,
    \Tile_X1Y3_FrameData_O[23] ,
    \Tile_X1Y3_FrameData_O[22] ,
    \Tile_X1Y3_FrameData_O[21] ,
    \Tile_X1Y3_FrameData_O[20] ,
    \Tile_X1Y3_FrameData_O[19] ,
    \Tile_X1Y3_FrameData_O[18] ,
    \Tile_X1Y3_FrameData_O[17] ,
    \Tile_X1Y3_FrameData_O[16] ,
    \Tile_X1Y3_FrameData_O[15] ,
    \Tile_X1Y3_FrameData_O[14] ,
    \Tile_X1Y3_FrameData_O[13] ,
    \Tile_X1Y3_FrameData_O[12] ,
    \Tile_X1Y3_FrameData_O[11] ,
    \Tile_X1Y3_FrameData_O[10] ,
    \Tile_X1Y3_FrameData_O[9] ,
    \Tile_X1Y3_FrameData_O[8] ,
    \Tile_X1Y3_FrameData_O[7] ,
    \Tile_X1Y3_FrameData_O[6] ,
    \Tile_X1Y3_FrameData_O[5] ,
    \Tile_X1Y3_FrameData_O[4] ,
    \Tile_X1Y3_FrameData_O[3] ,
    \Tile_X1Y3_FrameData_O[2] ,
    \Tile_X1Y3_FrameData_O[1] ,
    \Tile_X1Y3_FrameData_O[0] }),
    .FrameData_O({\Tile_X2Y3_FrameData_O[31] ,
    \Tile_X2Y3_FrameData_O[30] ,
    \Tile_X2Y3_FrameData_O[29] ,
    \Tile_X2Y3_FrameData_O[28] ,
    \Tile_X2Y3_FrameData_O[27] ,
    \Tile_X2Y3_FrameData_O[26] ,
    \Tile_X2Y3_FrameData_O[25] ,
    \Tile_X2Y3_FrameData_O[24] ,
    \Tile_X2Y3_FrameData_O[23] ,
    \Tile_X2Y3_FrameData_O[22] ,
    \Tile_X2Y3_FrameData_O[21] ,
    \Tile_X2Y3_FrameData_O[20] ,
    \Tile_X2Y3_FrameData_O[19] ,
    \Tile_X2Y3_FrameData_O[18] ,
    \Tile_X2Y3_FrameData_O[17] ,
    \Tile_X2Y3_FrameData_O[16] ,
    \Tile_X2Y3_FrameData_O[15] ,
    \Tile_X2Y3_FrameData_O[14] ,
    \Tile_X2Y3_FrameData_O[13] ,
    \Tile_X2Y3_FrameData_O[12] ,
    \Tile_X2Y3_FrameData_O[11] ,
    \Tile_X2Y3_FrameData_O[10] ,
    \Tile_X2Y3_FrameData_O[9] ,
    \Tile_X2Y3_FrameData_O[8] ,
    \Tile_X2Y3_FrameData_O[7] ,
    \Tile_X2Y3_FrameData_O[6] ,
    \Tile_X2Y3_FrameData_O[5] ,
    \Tile_X2Y3_FrameData_O[4] ,
    \Tile_X2Y3_FrameData_O[3] ,
    \Tile_X2Y3_FrameData_O[2] ,
    \Tile_X2Y3_FrameData_O[1] ,
    \Tile_X2Y3_FrameData_O[0] }),
    .FrameStrobe({\Tile_X2Y4_FrameStrobe_O[19] ,
    \Tile_X2Y4_FrameStrobe_O[18] ,
    \Tile_X2Y4_FrameStrobe_O[17] ,
    \Tile_X2Y4_FrameStrobe_O[16] ,
    \Tile_X2Y4_FrameStrobe_O[15] ,
    \Tile_X2Y4_FrameStrobe_O[14] ,
    \Tile_X2Y4_FrameStrobe_O[13] ,
    \Tile_X2Y4_FrameStrobe_O[12] ,
    \Tile_X2Y4_FrameStrobe_O[11] ,
    \Tile_X2Y4_FrameStrobe_O[10] ,
    \Tile_X2Y4_FrameStrobe_O[9] ,
    \Tile_X2Y4_FrameStrobe_O[8] ,
    \Tile_X2Y4_FrameStrobe_O[7] ,
    \Tile_X2Y4_FrameStrobe_O[6] ,
    \Tile_X2Y4_FrameStrobe_O[5] ,
    \Tile_X2Y4_FrameStrobe_O[4] ,
    \Tile_X2Y4_FrameStrobe_O[3] ,
    \Tile_X2Y4_FrameStrobe_O[2] ,
    \Tile_X2Y4_FrameStrobe_O[1] ,
    \Tile_X2Y4_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X2Y3_FrameStrobe_O[19] ,
    \Tile_X2Y3_FrameStrobe_O[18] ,
    \Tile_X2Y3_FrameStrobe_O[17] ,
    \Tile_X2Y3_FrameStrobe_O[16] ,
    \Tile_X2Y3_FrameStrobe_O[15] ,
    \Tile_X2Y3_FrameStrobe_O[14] ,
    \Tile_X2Y3_FrameStrobe_O[13] ,
    \Tile_X2Y3_FrameStrobe_O[12] ,
    \Tile_X2Y3_FrameStrobe_O[11] ,
    \Tile_X2Y3_FrameStrobe_O[10] ,
    \Tile_X2Y3_FrameStrobe_O[9] ,
    \Tile_X2Y3_FrameStrobe_O[8] ,
    \Tile_X2Y3_FrameStrobe_O[7] ,
    \Tile_X2Y3_FrameStrobe_O[6] ,
    \Tile_X2Y3_FrameStrobe_O[5] ,
    \Tile_X2Y3_FrameStrobe_O[4] ,
    \Tile_X2Y3_FrameStrobe_O[3] ,
    \Tile_X2Y3_FrameStrobe_O[2] ,
    \Tile_X2Y3_FrameStrobe_O[1] ,
    \Tile_X2Y3_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X2Y3_N1BEG[3] ,
    \Tile_X2Y3_N1BEG[2] ,
    \Tile_X2Y3_N1BEG[1] ,
    \Tile_X2Y3_N1BEG[0] }),
    .N1END({\Tile_X2Y4_N1BEG[3] ,
    \Tile_X2Y4_N1BEG[2] ,
    \Tile_X2Y4_N1BEG[1] ,
    \Tile_X2Y4_N1BEG[0] }),
    .N2BEG({\Tile_X2Y3_N2BEG[7] ,
    \Tile_X2Y3_N2BEG[6] ,
    \Tile_X2Y3_N2BEG[5] ,
    \Tile_X2Y3_N2BEG[4] ,
    \Tile_X2Y3_N2BEG[3] ,
    \Tile_X2Y3_N2BEG[2] ,
    \Tile_X2Y3_N2BEG[1] ,
    \Tile_X2Y3_N2BEG[0] }),
    .N2BEGb({\Tile_X2Y3_N2BEGb[7] ,
    \Tile_X2Y3_N2BEGb[6] ,
    \Tile_X2Y3_N2BEGb[5] ,
    \Tile_X2Y3_N2BEGb[4] ,
    \Tile_X2Y3_N2BEGb[3] ,
    \Tile_X2Y3_N2BEGb[2] ,
    \Tile_X2Y3_N2BEGb[1] ,
    \Tile_X2Y3_N2BEGb[0] }),
    .N2END({\Tile_X2Y4_N2BEGb[7] ,
    \Tile_X2Y4_N2BEGb[6] ,
    \Tile_X2Y4_N2BEGb[5] ,
    \Tile_X2Y4_N2BEGb[4] ,
    \Tile_X2Y4_N2BEGb[3] ,
    \Tile_X2Y4_N2BEGb[2] ,
    \Tile_X2Y4_N2BEGb[1] ,
    \Tile_X2Y4_N2BEGb[0] }),
    .N2MID({\Tile_X2Y4_N2BEG[7] ,
    \Tile_X2Y4_N2BEG[6] ,
    \Tile_X2Y4_N2BEG[5] ,
    \Tile_X2Y4_N2BEG[4] ,
    \Tile_X2Y4_N2BEG[3] ,
    \Tile_X2Y4_N2BEG[2] ,
    \Tile_X2Y4_N2BEG[1] ,
    \Tile_X2Y4_N2BEG[0] }),
    .N4BEG({\Tile_X2Y3_N4BEG[15] ,
    \Tile_X2Y3_N4BEG[14] ,
    \Tile_X2Y3_N4BEG[13] ,
    \Tile_X2Y3_N4BEG[12] ,
    \Tile_X2Y3_N4BEG[11] ,
    \Tile_X2Y3_N4BEG[10] ,
    \Tile_X2Y3_N4BEG[9] ,
    \Tile_X2Y3_N4BEG[8] ,
    \Tile_X2Y3_N4BEG[7] ,
    \Tile_X2Y3_N4BEG[6] ,
    \Tile_X2Y3_N4BEG[5] ,
    \Tile_X2Y3_N4BEG[4] ,
    \Tile_X2Y3_N4BEG[3] ,
    \Tile_X2Y3_N4BEG[2] ,
    \Tile_X2Y3_N4BEG[1] ,
    \Tile_X2Y3_N4BEG[0] }),
    .N4END({\Tile_X2Y4_N4BEG[15] ,
    \Tile_X2Y4_N4BEG[14] ,
    \Tile_X2Y4_N4BEG[13] ,
    \Tile_X2Y4_N4BEG[12] ,
    \Tile_X2Y4_N4BEG[11] ,
    \Tile_X2Y4_N4BEG[10] ,
    \Tile_X2Y4_N4BEG[9] ,
    \Tile_X2Y4_N4BEG[8] ,
    \Tile_X2Y4_N4BEG[7] ,
    \Tile_X2Y4_N4BEG[6] ,
    \Tile_X2Y4_N4BEG[5] ,
    \Tile_X2Y4_N4BEG[4] ,
    \Tile_X2Y4_N4BEG[3] ,
    \Tile_X2Y4_N4BEG[2] ,
    \Tile_X2Y4_N4BEG[1] ,
    \Tile_X2Y4_N4BEG[0] }),
    .NN4BEG({\Tile_X2Y3_NN4BEG[15] ,
    \Tile_X2Y3_NN4BEG[14] ,
    \Tile_X2Y3_NN4BEG[13] ,
    \Tile_X2Y3_NN4BEG[12] ,
    \Tile_X2Y3_NN4BEG[11] ,
    \Tile_X2Y3_NN4BEG[10] ,
    \Tile_X2Y3_NN4BEG[9] ,
    \Tile_X2Y3_NN4BEG[8] ,
    \Tile_X2Y3_NN4BEG[7] ,
    \Tile_X2Y3_NN4BEG[6] ,
    \Tile_X2Y3_NN4BEG[5] ,
    \Tile_X2Y3_NN4BEG[4] ,
    \Tile_X2Y3_NN4BEG[3] ,
    \Tile_X2Y3_NN4BEG[2] ,
    \Tile_X2Y3_NN4BEG[1] ,
    \Tile_X2Y3_NN4BEG[0] }),
    .NN4END({\Tile_X2Y4_NN4BEG[15] ,
    \Tile_X2Y4_NN4BEG[14] ,
    \Tile_X2Y4_NN4BEG[13] ,
    \Tile_X2Y4_NN4BEG[12] ,
    \Tile_X2Y4_NN4BEG[11] ,
    \Tile_X2Y4_NN4BEG[10] ,
    \Tile_X2Y4_NN4BEG[9] ,
    \Tile_X2Y4_NN4BEG[8] ,
    \Tile_X2Y4_NN4BEG[7] ,
    \Tile_X2Y4_NN4BEG[6] ,
    \Tile_X2Y4_NN4BEG[5] ,
    \Tile_X2Y4_NN4BEG[4] ,
    \Tile_X2Y4_NN4BEG[3] ,
    \Tile_X2Y4_NN4BEG[2] ,
    \Tile_X2Y4_NN4BEG[1] ,
    \Tile_X2Y4_NN4BEG[0] }),
    .S1BEG({\Tile_X2Y3_S1BEG[3] ,
    \Tile_X2Y3_S1BEG[2] ,
    \Tile_X2Y3_S1BEG[1] ,
    \Tile_X2Y3_S1BEG[0] }),
    .S1END({\Tile_X2Y2_S1BEG[3] ,
    \Tile_X2Y2_S1BEG[2] ,
    \Tile_X2Y2_S1BEG[1] ,
    \Tile_X2Y2_S1BEG[0] }),
    .S2BEG({\Tile_X2Y3_S2BEG[7] ,
    \Tile_X2Y3_S2BEG[6] ,
    \Tile_X2Y3_S2BEG[5] ,
    \Tile_X2Y3_S2BEG[4] ,
    \Tile_X2Y3_S2BEG[3] ,
    \Tile_X2Y3_S2BEG[2] ,
    \Tile_X2Y3_S2BEG[1] ,
    \Tile_X2Y3_S2BEG[0] }),
    .S2BEGb({\Tile_X2Y3_S2BEGb[7] ,
    \Tile_X2Y3_S2BEGb[6] ,
    \Tile_X2Y3_S2BEGb[5] ,
    \Tile_X2Y3_S2BEGb[4] ,
    \Tile_X2Y3_S2BEGb[3] ,
    \Tile_X2Y3_S2BEGb[2] ,
    \Tile_X2Y3_S2BEGb[1] ,
    \Tile_X2Y3_S2BEGb[0] }),
    .S2END({\Tile_X2Y2_S2BEGb[7] ,
    \Tile_X2Y2_S2BEGb[6] ,
    \Tile_X2Y2_S2BEGb[5] ,
    \Tile_X2Y2_S2BEGb[4] ,
    \Tile_X2Y2_S2BEGb[3] ,
    \Tile_X2Y2_S2BEGb[2] ,
    \Tile_X2Y2_S2BEGb[1] ,
    \Tile_X2Y2_S2BEGb[0] }),
    .S2MID({\Tile_X2Y2_S2BEG[7] ,
    \Tile_X2Y2_S2BEG[6] ,
    \Tile_X2Y2_S2BEG[5] ,
    \Tile_X2Y2_S2BEG[4] ,
    \Tile_X2Y2_S2BEG[3] ,
    \Tile_X2Y2_S2BEG[2] ,
    \Tile_X2Y2_S2BEG[1] ,
    \Tile_X2Y2_S2BEG[0] }),
    .S4BEG({\Tile_X2Y3_S4BEG[15] ,
    \Tile_X2Y3_S4BEG[14] ,
    \Tile_X2Y3_S4BEG[13] ,
    \Tile_X2Y3_S4BEG[12] ,
    \Tile_X2Y3_S4BEG[11] ,
    \Tile_X2Y3_S4BEG[10] ,
    \Tile_X2Y3_S4BEG[9] ,
    \Tile_X2Y3_S4BEG[8] ,
    \Tile_X2Y3_S4BEG[7] ,
    \Tile_X2Y3_S4BEG[6] ,
    \Tile_X2Y3_S4BEG[5] ,
    \Tile_X2Y3_S4BEG[4] ,
    \Tile_X2Y3_S4BEG[3] ,
    \Tile_X2Y3_S4BEG[2] ,
    \Tile_X2Y3_S4BEG[1] ,
    \Tile_X2Y3_S4BEG[0] }),
    .S4END({\Tile_X2Y2_S4BEG[15] ,
    \Tile_X2Y2_S4BEG[14] ,
    \Tile_X2Y2_S4BEG[13] ,
    \Tile_X2Y2_S4BEG[12] ,
    \Tile_X2Y2_S4BEG[11] ,
    \Tile_X2Y2_S4BEG[10] ,
    \Tile_X2Y2_S4BEG[9] ,
    \Tile_X2Y2_S4BEG[8] ,
    \Tile_X2Y2_S4BEG[7] ,
    \Tile_X2Y2_S4BEG[6] ,
    \Tile_X2Y2_S4BEG[5] ,
    \Tile_X2Y2_S4BEG[4] ,
    \Tile_X2Y2_S4BEG[3] ,
    \Tile_X2Y2_S4BEG[2] ,
    \Tile_X2Y2_S4BEG[1] ,
    \Tile_X2Y2_S4BEG[0] }),
    .SS4BEG({\Tile_X2Y3_SS4BEG[15] ,
    \Tile_X2Y3_SS4BEG[14] ,
    \Tile_X2Y3_SS4BEG[13] ,
    \Tile_X2Y3_SS4BEG[12] ,
    \Tile_X2Y3_SS4BEG[11] ,
    \Tile_X2Y3_SS4BEG[10] ,
    \Tile_X2Y3_SS4BEG[9] ,
    \Tile_X2Y3_SS4BEG[8] ,
    \Tile_X2Y3_SS4BEG[7] ,
    \Tile_X2Y3_SS4BEG[6] ,
    \Tile_X2Y3_SS4BEG[5] ,
    \Tile_X2Y3_SS4BEG[4] ,
    \Tile_X2Y3_SS4BEG[3] ,
    \Tile_X2Y3_SS4BEG[2] ,
    \Tile_X2Y3_SS4BEG[1] ,
    \Tile_X2Y3_SS4BEG[0] }),
    .SS4END({\Tile_X2Y2_SS4BEG[15] ,
    \Tile_X2Y2_SS4BEG[14] ,
    \Tile_X2Y2_SS4BEG[13] ,
    \Tile_X2Y2_SS4BEG[12] ,
    \Tile_X2Y2_SS4BEG[11] ,
    \Tile_X2Y2_SS4BEG[10] ,
    \Tile_X2Y2_SS4BEG[9] ,
    \Tile_X2Y2_SS4BEG[8] ,
    \Tile_X2Y2_SS4BEG[7] ,
    \Tile_X2Y2_SS4BEG[6] ,
    \Tile_X2Y2_SS4BEG[5] ,
    \Tile_X2Y2_SS4BEG[4] ,
    \Tile_X2Y2_SS4BEG[3] ,
    \Tile_X2Y2_SS4BEG[2] ,
    \Tile_X2Y2_SS4BEG[1] ,
    \Tile_X2Y2_SS4BEG[0] }),
    .W1BEG({\Tile_X2Y3_W1BEG[3] ,
    \Tile_X2Y3_W1BEG[2] ,
    \Tile_X2Y3_W1BEG[1] ,
    \Tile_X2Y3_W1BEG[0] }),
    .W1END({\Tile_X3Y3_W1BEG[3] ,
    \Tile_X3Y3_W1BEG[2] ,
    \Tile_X3Y3_W1BEG[1] ,
    \Tile_X3Y3_W1BEG[0] }),
    .W2BEG({\Tile_X2Y3_W2BEG[7] ,
    \Tile_X2Y3_W2BEG[6] ,
    \Tile_X2Y3_W2BEG[5] ,
    \Tile_X2Y3_W2BEG[4] ,
    \Tile_X2Y3_W2BEG[3] ,
    \Tile_X2Y3_W2BEG[2] ,
    \Tile_X2Y3_W2BEG[1] ,
    \Tile_X2Y3_W2BEG[0] }),
    .W2BEGb({\Tile_X2Y3_W2BEGb[7] ,
    \Tile_X2Y3_W2BEGb[6] ,
    \Tile_X2Y3_W2BEGb[5] ,
    \Tile_X2Y3_W2BEGb[4] ,
    \Tile_X2Y3_W2BEGb[3] ,
    \Tile_X2Y3_W2BEGb[2] ,
    \Tile_X2Y3_W2BEGb[1] ,
    \Tile_X2Y3_W2BEGb[0] }),
    .W2END({\Tile_X3Y3_W2BEGb[7] ,
    \Tile_X3Y3_W2BEGb[6] ,
    \Tile_X3Y3_W2BEGb[5] ,
    \Tile_X3Y3_W2BEGb[4] ,
    \Tile_X3Y3_W2BEGb[3] ,
    \Tile_X3Y3_W2BEGb[2] ,
    \Tile_X3Y3_W2BEGb[1] ,
    \Tile_X3Y3_W2BEGb[0] }),
    .W2MID({\Tile_X3Y3_W2BEG[7] ,
    \Tile_X3Y3_W2BEG[6] ,
    \Tile_X3Y3_W2BEG[5] ,
    \Tile_X3Y3_W2BEG[4] ,
    \Tile_X3Y3_W2BEG[3] ,
    \Tile_X3Y3_W2BEG[2] ,
    \Tile_X3Y3_W2BEG[1] ,
    \Tile_X3Y3_W2BEG[0] }),
    .W6BEG({\Tile_X2Y3_W6BEG[11] ,
    \Tile_X2Y3_W6BEG[10] ,
    \Tile_X2Y3_W6BEG[9] ,
    \Tile_X2Y3_W6BEG[8] ,
    \Tile_X2Y3_W6BEG[7] ,
    \Tile_X2Y3_W6BEG[6] ,
    \Tile_X2Y3_W6BEG[5] ,
    \Tile_X2Y3_W6BEG[4] ,
    \Tile_X2Y3_W6BEG[3] ,
    \Tile_X2Y3_W6BEG[2] ,
    \Tile_X2Y3_W6BEG[1] ,
    \Tile_X2Y3_W6BEG[0] }),
    .W6END({\Tile_X3Y3_W6BEG[11] ,
    \Tile_X3Y3_W6BEG[10] ,
    \Tile_X3Y3_W6BEG[9] ,
    \Tile_X3Y3_W6BEG[8] ,
    \Tile_X3Y3_W6BEG[7] ,
    \Tile_X3Y3_W6BEG[6] ,
    \Tile_X3Y3_W6BEG[5] ,
    \Tile_X3Y3_W6BEG[4] ,
    \Tile_X3Y3_W6BEG[3] ,
    \Tile_X3Y3_W6BEG[2] ,
    \Tile_X3Y3_W6BEG[1] ,
    \Tile_X3Y3_W6BEG[0] }),
    .WW4BEG({\Tile_X2Y3_WW4BEG[15] ,
    \Tile_X2Y3_WW4BEG[14] ,
    \Tile_X2Y3_WW4BEG[13] ,
    \Tile_X2Y3_WW4BEG[12] ,
    \Tile_X2Y3_WW4BEG[11] ,
    \Tile_X2Y3_WW4BEG[10] ,
    \Tile_X2Y3_WW4BEG[9] ,
    \Tile_X2Y3_WW4BEG[8] ,
    \Tile_X2Y3_WW4BEG[7] ,
    \Tile_X2Y3_WW4BEG[6] ,
    \Tile_X2Y3_WW4BEG[5] ,
    \Tile_X2Y3_WW4BEG[4] ,
    \Tile_X2Y3_WW4BEG[3] ,
    \Tile_X2Y3_WW4BEG[2] ,
    \Tile_X2Y3_WW4BEG[1] ,
    \Tile_X2Y3_WW4BEG[0] }),
    .WW4END({\Tile_X3Y3_WW4BEG[15] ,
    \Tile_X3Y3_WW4BEG[14] ,
    \Tile_X3Y3_WW4BEG[13] ,
    \Tile_X3Y3_WW4BEG[12] ,
    \Tile_X3Y3_WW4BEG[11] ,
    \Tile_X3Y3_WW4BEG[10] ,
    \Tile_X3Y3_WW4BEG[9] ,
    \Tile_X3Y3_WW4BEG[8] ,
    \Tile_X3Y3_WW4BEG[7] ,
    \Tile_X3Y3_WW4BEG[6] ,
    \Tile_X3Y3_WW4BEG[5] ,
    \Tile_X3Y3_WW4BEG[4] ,
    \Tile_X3Y3_WW4BEG[3] ,
    \Tile_X3Y3_WW4BEG[2] ,
    \Tile_X3Y3_WW4BEG[1] ,
    \Tile_X3Y3_WW4BEG[0] }));
 LUT4AB Tile_X2Y4_LUT4AB (.Ci(Tile_X2Y5_Co),
    .Co(Tile_X2Y4_Co),
    .UserCLK(Tile_X2Y5_UserCLKo),
    .UserCLKo(Tile_X2Y4_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X2Y4_E1BEG[3] ,
    \Tile_X2Y4_E1BEG[2] ,
    \Tile_X2Y4_E1BEG[1] ,
    \Tile_X2Y4_E1BEG[0] }),
    .E1END({\Tile_X1Y4_E1BEG[3] ,
    \Tile_X1Y4_E1BEG[2] ,
    \Tile_X1Y4_E1BEG[1] ,
    \Tile_X1Y4_E1BEG[0] }),
    .E2BEG({\Tile_X2Y4_E2BEG[7] ,
    \Tile_X2Y4_E2BEG[6] ,
    \Tile_X2Y4_E2BEG[5] ,
    \Tile_X2Y4_E2BEG[4] ,
    \Tile_X2Y4_E2BEG[3] ,
    \Tile_X2Y4_E2BEG[2] ,
    \Tile_X2Y4_E2BEG[1] ,
    \Tile_X2Y4_E2BEG[0] }),
    .E2BEGb({\Tile_X2Y4_E2BEGb[7] ,
    \Tile_X2Y4_E2BEGb[6] ,
    \Tile_X2Y4_E2BEGb[5] ,
    \Tile_X2Y4_E2BEGb[4] ,
    \Tile_X2Y4_E2BEGb[3] ,
    \Tile_X2Y4_E2BEGb[2] ,
    \Tile_X2Y4_E2BEGb[1] ,
    \Tile_X2Y4_E2BEGb[0] }),
    .E2END({\Tile_X1Y4_E2BEGb[7] ,
    \Tile_X1Y4_E2BEGb[6] ,
    \Tile_X1Y4_E2BEGb[5] ,
    \Tile_X1Y4_E2BEGb[4] ,
    \Tile_X1Y4_E2BEGb[3] ,
    \Tile_X1Y4_E2BEGb[2] ,
    \Tile_X1Y4_E2BEGb[1] ,
    \Tile_X1Y4_E2BEGb[0] }),
    .E2MID({\Tile_X1Y4_E2BEG[7] ,
    \Tile_X1Y4_E2BEG[6] ,
    \Tile_X1Y4_E2BEG[5] ,
    \Tile_X1Y4_E2BEG[4] ,
    \Tile_X1Y4_E2BEG[3] ,
    \Tile_X1Y4_E2BEG[2] ,
    \Tile_X1Y4_E2BEG[1] ,
    \Tile_X1Y4_E2BEG[0] }),
    .E6BEG({\Tile_X2Y4_E6BEG[11] ,
    \Tile_X2Y4_E6BEG[10] ,
    \Tile_X2Y4_E6BEG[9] ,
    \Tile_X2Y4_E6BEG[8] ,
    \Tile_X2Y4_E6BEG[7] ,
    \Tile_X2Y4_E6BEG[6] ,
    \Tile_X2Y4_E6BEG[5] ,
    \Tile_X2Y4_E6BEG[4] ,
    \Tile_X2Y4_E6BEG[3] ,
    \Tile_X2Y4_E6BEG[2] ,
    \Tile_X2Y4_E6BEG[1] ,
    \Tile_X2Y4_E6BEG[0] }),
    .E6END({\Tile_X1Y4_E6BEG[11] ,
    \Tile_X1Y4_E6BEG[10] ,
    \Tile_X1Y4_E6BEG[9] ,
    \Tile_X1Y4_E6BEG[8] ,
    \Tile_X1Y4_E6BEG[7] ,
    \Tile_X1Y4_E6BEG[6] ,
    \Tile_X1Y4_E6BEG[5] ,
    \Tile_X1Y4_E6BEG[4] ,
    \Tile_X1Y4_E6BEG[3] ,
    \Tile_X1Y4_E6BEG[2] ,
    \Tile_X1Y4_E6BEG[1] ,
    \Tile_X1Y4_E6BEG[0] }),
    .EE4BEG({\Tile_X2Y4_EE4BEG[15] ,
    \Tile_X2Y4_EE4BEG[14] ,
    \Tile_X2Y4_EE4BEG[13] ,
    \Tile_X2Y4_EE4BEG[12] ,
    \Tile_X2Y4_EE4BEG[11] ,
    \Tile_X2Y4_EE4BEG[10] ,
    \Tile_X2Y4_EE4BEG[9] ,
    \Tile_X2Y4_EE4BEG[8] ,
    \Tile_X2Y4_EE4BEG[7] ,
    \Tile_X2Y4_EE4BEG[6] ,
    \Tile_X2Y4_EE4BEG[5] ,
    \Tile_X2Y4_EE4BEG[4] ,
    \Tile_X2Y4_EE4BEG[3] ,
    \Tile_X2Y4_EE4BEG[2] ,
    \Tile_X2Y4_EE4BEG[1] ,
    \Tile_X2Y4_EE4BEG[0] }),
    .EE4END({\Tile_X1Y4_EE4BEG[15] ,
    \Tile_X1Y4_EE4BEG[14] ,
    \Tile_X1Y4_EE4BEG[13] ,
    \Tile_X1Y4_EE4BEG[12] ,
    \Tile_X1Y4_EE4BEG[11] ,
    \Tile_X1Y4_EE4BEG[10] ,
    \Tile_X1Y4_EE4BEG[9] ,
    \Tile_X1Y4_EE4BEG[8] ,
    \Tile_X1Y4_EE4BEG[7] ,
    \Tile_X1Y4_EE4BEG[6] ,
    \Tile_X1Y4_EE4BEG[5] ,
    \Tile_X1Y4_EE4BEG[4] ,
    \Tile_X1Y4_EE4BEG[3] ,
    \Tile_X1Y4_EE4BEG[2] ,
    \Tile_X1Y4_EE4BEG[1] ,
    \Tile_X1Y4_EE4BEG[0] }),
    .FrameData({\Tile_X1Y4_FrameData_O[31] ,
    \Tile_X1Y4_FrameData_O[30] ,
    \Tile_X1Y4_FrameData_O[29] ,
    \Tile_X1Y4_FrameData_O[28] ,
    \Tile_X1Y4_FrameData_O[27] ,
    \Tile_X1Y4_FrameData_O[26] ,
    \Tile_X1Y4_FrameData_O[25] ,
    \Tile_X1Y4_FrameData_O[24] ,
    \Tile_X1Y4_FrameData_O[23] ,
    \Tile_X1Y4_FrameData_O[22] ,
    \Tile_X1Y4_FrameData_O[21] ,
    \Tile_X1Y4_FrameData_O[20] ,
    \Tile_X1Y4_FrameData_O[19] ,
    \Tile_X1Y4_FrameData_O[18] ,
    \Tile_X1Y4_FrameData_O[17] ,
    \Tile_X1Y4_FrameData_O[16] ,
    \Tile_X1Y4_FrameData_O[15] ,
    \Tile_X1Y4_FrameData_O[14] ,
    \Tile_X1Y4_FrameData_O[13] ,
    \Tile_X1Y4_FrameData_O[12] ,
    \Tile_X1Y4_FrameData_O[11] ,
    \Tile_X1Y4_FrameData_O[10] ,
    \Tile_X1Y4_FrameData_O[9] ,
    \Tile_X1Y4_FrameData_O[8] ,
    \Tile_X1Y4_FrameData_O[7] ,
    \Tile_X1Y4_FrameData_O[6] ,
    \Tile_X1Y4_FrameData_O[5] ,
    \Tile_X1Y4_FrameData_O[4] ,
    \Tile_X1Y4_FrameData_O[3] ,
    \Tile_X1Y4_FrameData_O[2] ,
    \Tile_X1Y4_FrameData_O[1] ,
    \Tile_X1Y4_FrameData_O[0] }),
    .FrameData_O({\Tile_X2Y4_FrameData_O[31] ,
    \Tile_X2Y4_FrameData_O[30] ,
    \Tile_X2Y4_FrameData_O[29] ,
    \Tile_X2Y4_FrameData_O[28] ,
    \Tile_X2Y4_FrameData_O[27] ,
    \Tile_X2Y4_FrameData_O[26] ,
    \Tile_X2Y4_FrameData_O[25] ,
    \Tile_X2Y4_FrameData_O[24] ,
    \Tile_X2Y4_FrameData_O[23] ,
    \Tile_X2Y4_FrameData_O[22] ,
    \Tile_X2Y4_FrameData_O[21] ,
    \Tile_X2Y4_FrameData_O[20] ,
    \Tile_X2Y4_FrameData_O[19] ,
    \Tile_X2Y4_FrameData_O[18] ,
    \Tile_X2Y4_FrameData_O[17] ,
    \Tile_X2Y4_FrameData_O[16] ,
    \Tile_X2Y4_FrameData_O[15] ,
    \Tile_X2Y4_FrameData_O[14] ,
    \Tile_X2Y4_FrameData_O[13] ,
    \Tile_X2Y4_FrameData_O[12] ,
    \Tile_X2Y4_FrameData_O[11] ,
    \Tile_X2Y4_FrameData_O[10] ,
    \Tile_X2Y4_FrameData_O[9] ,
    \Tile_X2Y4_FrameData_O[8] ,
    \Tile_X2Y4_FrameData_O[7] ,
    \Tile_X2Y4_FrameData_O[6] ,
    \Tile_X2Y4_FrameData_O[5] ,
    \Tile_X2Y4_FrameData_O[4] ,
    \Tile_X2Y4_FrameData_O[3] ,
    \Tile_X2Y4_FrameData_O[2] ,
    \Tile_X2Y4_FrameData_O[1] ,
    \Tile_X2Y4_FrameData_O[0] }),
    .FrameStrobe({\Tile_X2Y5_FrameStrobe_O[19] ,
    \Tile_X2Y5_FrameStrobe_O[18] ,
    \Tile_X2Y5_FrameStrobe_O[17] ,
    \Tile_X2Y5_FrameStrobe_O[16] ,
    \Tile_X2Y5_FrameStrobe_O[15] ,
    \Tile_X2Y5_FrameStrobe_O[14] ,
    \Tile_X2Y5_FrameStrobe_O[13] ,
    \Tile_X2Y5_FrameStrobe_O[12] ,
    \Tile_X2Y5_FrameStrobe_O[11] ,
    \Tile_X2Y5_FrameStrobe_O[10] ,
    \Tile_X2Y5_FrameStrobe_O[9] ,
    \Tile_X2Y5_FrameStrobe_O[8] ,
    \Tile_X2Y5_FrameStrobe_O[7] ,
    \Tile_X2Y5_FrameStrobe_O[6] ,
    \Tile_X2Y5_FrameStrobe_O[5] ,
    \Tile_X2Y5_FrameStrobe_O[4] ,
    \Tile_X2Y5_FrameStrobe_O[3] ,
    \Tile_X2Y5_FrameStrobe_O[2] ,
    \Tile_X2Y5_FrameStrobe_O[1] ,
    \Tile_X2Y5_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X2Y4_FrameStrobe_O[19] ,
    \Tile_X2Y4_FrameStrobe_O[18] ,
    \Tile_X2Y4_FrameStrobe_O[17] ,
    \Tile_X2Y4_FrameStrobe_O[16] ,
    \Tile_X2Y4_FrameStrobe_O[15] ,
    \Tile_X2Y4_FrameStrobe_O[14] ,
    \Tile_X2Y4_FrameStrobe_O[13] ,
    \Tile_X2Y4_FrameStrobe_O[12] ,
    \Tile_X2Y4_FrameStrobe_O[11] ,
    \Tile_X2Y4_FrameStrobe_O[10] ,
    \Tile_X2Y4_FrameStrobe_O[9] ,
    \Tile_X2Y4_FrameStrobe_O[8] ,
    \Tile_X2Y4_FrameStrobe_O[7] ,
    \Tile_X2Y4_FrameStrobe_O[6] ,
    \Tile_X2Y4_FrameStrobe_O[5] ,
    \Tile_X2Y4_FrameStrobe_O[4] ,
    \Tile_X2Y4_FrameStrobe_O[3] ,
    \Tile_X2Y4_FrameStrobe_O[2] ,
    \Tile_X2Y4_FrameStrobe_O[1] ,
    \Tile_X2Y4_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X2Y4_N1BEG[3] ,
    \Tile_X2Y4_N1BEG[2] ,
    \Tile_X2Y4_N1BEG[1] ,
    \Tile_X2Y4_N1BEG[0] }),
    .N1END({\Tile_X2Y5_N1BEG[3] ,
    \Tile_X2Y5_N1BEG[2] ,
    \Tile_X2Y5_N1BEG[1] ,
    \Tile_X2Y5_N1BEG[0] }),
    .N2BEG({\Tile_X2Y4_N2BEG[7] ,
    \Tile_X2Y4_N2BEG[6] ,
    \Tile_X2Y4_N2BEG[5] ,
    \Tile_X2Y4_N2BEG[4] ,
    \Tile_X2Y4_N2BEG[3] ,
    \Tile_X2Y4_N2BEG[2] ,
    \Tile_X2Y4_N2BEG[1] ,
    \Tile_X2Y4_N2BEG[0] }),
    .N2BEGb({\Tile_X2Y4_N2BEGb[7] ,
    \Tile_X2Y4_N2BEGb[6] ,
    \Tile_X2Y4_N2BEGb[5] ,
    \Tile_X2Y4_N2BEGb[4] ,
    \Tile_X2Y4_N2BEGb[3] ,
    \Tile_X2Y4_N2BEGb[2] ,
    \Tile_X2Y4_N2BEGb[1] ,
    \Tile_X2Y4_N2BEGb[0] }),
    .N2END({\Tile_X2Y5_N2BEGb[7] ,
    \Tile_X2Y5_N2BEGb[6] ,
    \Tile_X2Y5_N2BEGb[5] ,
    \Tile_X2Y5_N2BEGb[4] ,
    \Tile_X2Y5_N2BEGb[3] ,
    \Tile_X2Y5_N2BEGb[2] ,
    \Tile_X2Y5_N2BEGb[1] ,
    \Tile_X2Y5_N2BEGb[0] }),
    .N2MID({\Tile_X2Y5_N2BEG[7] ,
    \Tile_X2Y5_N2BEG[6] ,
    \Tile_X2Y5_N2BEG[5] ,
    \Tile_X2Y5_N2BEG[4] ,
    \Tile_X2Y5_N2BEG[3] ,
    \Tile_X2Y5_N2BEG[2] ,
    \Tile_X2Y5_N2BEG[1] ,
    \Tile_X2Y5_N2BEG[0] }),
    .N4BEG({\Tile_X2Y4_N4BEG[15] ,
    \Tile_X2Y4_N4BEG[14] ,
    \Tile_X2Y4_N4BEG[13] ,
    \Tile_X2Y4_N4BEG[12] ,
    \Tile_X2Y4_N4BEG[11] ,
    \Tile_X2Y4_N4BEG[10] ,
    \Tile_X2Y4_N4BEG[9] ,
    \Tile_X2Y4_N4BEG[8] ,
    \Tile_X2Y4_N4BEG[7] ,
    \Tile_X2Y4_N4BEG[6] ,
    \Tile_X2Y4_N4BEG[5] ,
    \Tile_X2Y4_N4BEG[4] ,
    \Tile_X2Y4_N4BEG[3] ,
    \Tile_X2Y4_N4BEG[2] ,
    \Tile_X2Y4_N4BEG[1] ,
    \Tile_X2Y4_N4BEG[0] }),
    .N4END({\Tile_X2Y5_N4BEG[15] ,
    \Tile_X2Y5_N4BEG[14] ,
    \Tile_X2Y5_N4BEG[13] ,
    \Tile_X2Y5_N4BEG[12] ,
    \Tile_X2Y5_N4BEG[11] ,
    \Tile_X2Y5_N4BEG[10] ,
    \Tile_X2Y5_N4BEG[9] ,
    \Tile_X2Y5_N4BEG[8] ,
    \Tile_X2Y5_N4BEG[7] ,
    \Tile_X2Y5_N4BEG[6] ,
    \Tile_X2Y5_N4BEG[5] ,
    \Tile_X2Y5_N4BEG[4] ,
    \Tile_X2Y5_N4BEG[3] ,
    \Tile_X2Y5_N4BEG[2] ,
    \Tile_X2Y5_N4BEG[1] ,
    \Tile_X2Y5_N4BEG[0] }),
    .NN4BEG({\Tile_X2Y4_NN4BEG[15] ,
    \Tile_X2Y4_NN4BEG[14] ,
    \Tile_X2Y4_NN4BEG[13] ,
    \Tile_X2Y4_NN4BEG[12] ,
    \Tile_X2Y4_NN4BEG[11] ,
    \Tile_X2Y4_NN4BEG[10] ,
    \Tile_X2Y4_NN4BEG[9] ,
    \Tile_X2Y4_NN4BEG[8] ,
    \Tile_X2Y4_NN4BEG[7] ,
    \Tile_X2Y4_NN4BEG[6] ,
    \Tile_X2Y4_NN4BEG[5] ,
    \Tile_X2Y4_NN4BEG[4] ,
    \Tile_X2Y4_NN4BEG[3] ,
    \Tile_X2Y4_NN4BEG[2] ,
    \Tile_X2Y4_NN4BEG[1] ,
    \Tile_X2Y4_NN4BEG[0] }),
    .NN4END({\Tile_X2Y5_NN4BEG[15] ,
    \Tile_X2Y5_NN4BEG[14] ,
    \Tile_X2Y5_NN4BEG[13] ,
    \Tile_X2Y5_NN4BEG[12] ,
    \Tile_X2Y5_NN4BEG[11] ,
    \Tile_X2Y5_NN4BEG[10] ,
    \Tile_X2Y5_NN4BEG[9] ,
    \Tile_X2Y5_NN4BEG[8] ,
    \Tile_X2Y5_NN4BEG[7] ,
    \Tile_X2Y5_NN4BEG[6] ,
    \Tile_X2Y5_NN4BEG[5] ,
    \Tile_X2Y5_NN4BEG[4] ,
    \Tile_X2Y5_NN4BEG[3] ,
    \Tile_X2Y5_NN4BEG[2] ,
    \Tile_X2Y5_NN4BEG[1] ,
    \Tile_X2Y5_NN4BEG[0] }),
    .S1BEG({\Tile_X2Y4_S1BEG[3] ,
    \Tile_X2Y4_S1BEG[2] ,
    \Tile_X2Y4_S1BEG[1] ,
    \Tile_X2Y4_S1BEG[0] }),
    .S1END({\Tile_X2Y3_S1BEG[3] ,
    \Tile_X2Y3_S1BEG[2] ,
    \Tile_X2Y3_S1BEG[1] ,
    \Tile_X2Y3_S1BEG[0] }),
    .S2BEG({\Tile_X2Y4_S2BEG[7] ,
    \Tile_X2Y4_S2BEG[6] ,
    \Tile_X2Y4_S2BEG[5] ,
    \Tile_X2Y4_S2BEG[4] ,
    \Tile_X2Y4_S2BEG[3] ,
    \Tile_X2Y4_S2BEG[2] ,
    \Tile_X2Y4_S2BEG[1] ,
    \Tile_X2Y4_S2BEG[0] }),
    .S2BEGb({\Tile_X2Y4_S2BEGb[7] ,
    \Tile_X2Y4_S2BEGb[6] ,
    \Tile_X2Y4_S2BEGb[5] ,
    \Tile_X2Y4_S2BEGb[4] ,
    \Tile_X2Y4_S2BEGb[3] ,
    \Tile_X2Y4_S2BEGb[2] ,
    \Tile_X2Y4_S2BEGb[1] ,
    \Tile_X2Y4_S2BEGb[0] }),
    .S2END({\Tile_X2Y3_S2BEGb[7] ,
    \Tile_X2Y3_S2BEGb[6] ,
    \Tile_X2Y3_S2BEGb[5] ,
    \Tile_X2Y3_S2BEGb[4] ,
    \Tile_X2Y3_S2BEGb[3] ,
    \Tile_X2Y3_S2BEGb[2] ,
    \Tile_X2Y3_S2BEGb[1] ,
    \Tile_X2Y3_S2BEGb[0] }),
    .S2MID({\Tile_X2Y3_S2BEG[7] ,
    \Tile_X2Y3_S2BEG[6] ,
    \Tile_X2Y3_S2BEG[5] ,
    \Tile_X2Y3_S2BEG[4] ,
    \Tile_X2Y3_S2BEG[3] ,
    \Tile_X2Y3_S2BEG[2] ,
    \Tile_X2Y3_S2BEG[1] ,
    \Tile_X2Y3_S2BEG[0] }),
    .S4BEG({\Tile_X2Y4_S4BEG[15] ,
    \Tile_X2Y4_S4BEG[14] ,
    \Tile_X2Y4_S4BEG[13] ,
    \Tile_X2Y4_S4BEG[12] ,
    \Tile_X2Y4_S4BEG[11] ,
    \Tile_X2Y4_S4BEG[10] ,
    \Tile_X2Y4_S4BEG[9] ,
    \Tile_X2Y4_S4BEG[8] ,
    \Tile_X2Y4_S4BEG[7] ,
    \Tile_X2Y4_S4BEG[6] ,
    \Tile_X2Y4_S4BEG[5] ,
    \Tile_X2Y4_S4BEG[4] ,
    \Tile_X2Y4_S4BEG[3] ,
    \Tile_X2Y4_S4BEG[2] ,
    \Tile_X2Y4_S4BEG[1] ,
    \Tile_X2Y4_S4BEG[0] }),
    .S4END({\Tile_X2Y3_S4BEG[15] ,
    \Tile_X2Y3_S4BEG[14] ,
    \Tile_X2Y3_S4BEG[13] ,
    \Tile_X2Y3_S4BEG[12] ,
    \Tile_X2Y3_S4BEG[11] ,
    \Tile_X2Y3_S4BEG[10] ,
    \Tile_X2Y3_S4BEG[9] ,
    \Tile_X2Y3_S4BEG[8] ,
    \Tile_X2Y3_S4BEG[7] ,
    \Tile_X2Y3_S4BEG[6] ,
    \Tile_X2Y3_S4BEG[5] ,
    \Tile_X2Y3_S4BEG[4] ,
    \Tile_X2Y3_S4BEG[3] ,
    \Tile_X2Y3_S4BEG[2] ,
    \Tile_X2Y3_S4BEG[1] ,
    \Tile_X2Y3_S4BEG[0] }),
    .SS4BEG({\Tile_X2Y4_SS4BEG[15] ,
    \Tile_X2Y4_SS4BEG[14] ,
    \Tile_X2Y4_SS4BEG[13] ,
    \Tile_X2Y4_SS4BEG[12] ,
    \Tile_X2Y4_SS4BEG[11] ,
    \Tile_X2Y4_SS4BEG[10] ,
    \Tile_X2Y4_SS4BEG[9] ,
    \Tile_X2Y4_SS4BEG[8] ,
    \Tile_X2Y4_SS4BEG[7] ,
    \Tile_X2Y4_SS4BEG[6] ,
    \Tile_X2Y4_SS4BEG[5] ,
    \Tile_X2Y4_SS4BEG[4] ,
    \Tile_X2Y4_SS4BEG[3] ,
    \Tile_X2Y4_SS4BEG[2] ,
    \Tile_X2Y4_SS4BEG[1] ,
    \Tile_X2Y4_SS4BEG[0] }),
    .SS4END({\Tile_X2Y3_SS4BEG[15] ,
    \Tile_X2Y3_SS4BEG[14] ,
    \Tile_X2Y3_SS4BEG[13] ,
    \Tile_X2Y3_SS4BEG[12] ,
    \Tile_X2Y3_SS4BEG[11] ,
    \Tile_X2Y3_SS4BEG[10] ,
    \Tile_X2Y3_SS4BEG[9] ,
    \Tile_X2Y3_SS4BEG[8] ,
    \Tile_X2Y3_SS4BEG[7] ,
    \Tile_X2Y3_SS4BEG[6] ,
    \Tile_X2Y3_SS4BEG[5] ,
    \Tile_X2Y3_SS4BEG[4] ,
    \Tile_X2Y3_SS4BEG[3] ,
    \Tile_X2Y3_SS4BEG[2] ,
    \Tile_X2Y3_SS4BEG[1] ,
    \Tile_X2Y3_SS4BEG[0] }),
    .W1BEG({\Tile_X2Y4_W1BEG[3] ,
    \Tile_X2Y4_W1BEG[2] ,
    \Tile_X2Y4_W1BEG[1] ,
    \Tile_X2Y4_W1BEG[0] }),
    .W1END({\Tile_X3Y4_W1BEG[3] ,
    \Tile_X3Y4_W1BEG[2] ,
    \Tile_X3Y4_W1BEG[1] ,
    \Tile_X3Y4_W1BEG[0] }),
    .W2BEG({\Tile_X2Y4_W2BEG[7] ,
    \Tile_X2Y4_W2BEG[6] ,
    \Tile_X2Y4_W2BEG[5] ,
    \Tile_X2Y4_W2BEG[4] ,
    \Tile_X2Y4_W2BEG[3] ,
    \Tile_X2Y4_W2BEG[2] ,
    \Tile_X2Y4_W2BEG[1] ,
    \Tile_X2Y4_W2BEG[0] }),
    .W2BEGb({\Tile_X2Y4_W2BEGb[7] ,
    \Tile_X2Y4_W2BEGb[6] ,
    \Tile_X2Y4_W2BEGb[5] ,
    \Tile_X2Y4_W2BEGb[4] ,
    \Tile_X2Y4_W2BEGb[3] ,
    \Tile_X2Y4_W2BEGb[2] ,
    \Tile_X2Y4_W2BEGb[1] ,
    \Tile_X2Y4_W2BEGb[0] }),
    .W2END({\Tile_X3Y4_W2BEGb[7] ,
    \Tile_X3Y4_W2BEGb[6] ,
    \Tile_X3Y4_W2BEGb[5] ,
    \Tile_X3Y4_W2BEGb[4] ,
    \Tile_X3Y4_W2BEGb[3] ,
    \Tile_X3Y4_W2BEGb[2] ,
    \Tile_X3Y4_W2BEGb[1] ,
    \Tile_X3Y4_W2BEGb[0] }),
    .W2MID({\Tile_X3Y4_W2BEG[7] ,
    \Tile_X3Y4_W2BEG[6] ,
    \Tile_X3Y4_W2BEG[5] ,
    \Tile_X3Y4_W2BEG[4] ,
    \Tile_X3Y4_W2BEG[3] ,
    \Tile_X3Y4_W2BEG[2] ,
    \Tile_X3Y4_W2BEG[1] ,
    \Tile_X3Y4_W2BEG[0] }),
    .W6BEG({\Tile_X2Y4_W6BEG[11] ,
    \Tile_X2Y4_W6BEG[10] ,
    \Tile_X2Y4_W6BEG[9] ,
    \Tile_X2Y4_W6BEG[8] ,
    \Tile_X2Y4_W6BEG[7] ,
    \Tile_X2Y4_W6BEG[6] ,
    \Tile_X2Y4_W6BEG[5] ,
    \Tile_X2Y4_W6BEG[4] ,
    \Tile_X2Y4_W6BEG[3] ,
    \Tile_X2Y4_W6BEG[2] ,
    \Tile_X2Y4_W6BEG[1] ,
    \Tile_X2Y4_W6BEG[0] }),
    .W6END({\Tile_X3Y4_W6BEG[11] ,
    \Tile_X3Y4_W6BEG[10] ,
    \Tile_X3Y4_W6BEG[9] ,
    \Tile_X3Y4_W6BEG[8] ,
    \Tile_X3Y4_W6BEG[7] ,
    \Tile_X3Y4_W6BEG[6] ,
    \Tile_X3Y4_W6BEG[5] ,
    \Tile_X3Y4_W6BEG[4] ,
    \Tile_X3Y4_W6BEG[3] ,
    \Tile_X3Y4_W6BEG[2] ,
    \Tile_X3Y4_W6BEG[1] ,
    \Tile_X3Y4_W6BEG[0] }),
    .WW4BEG({\Tile_X2Y4_WW4BEG[15] ,
    \Tile_X2Y4_WW4BEG[14] ,
    \Tile_X2Y4_WW4BEG[13] ,
    \Tile_X2Y4_WW4BEG[12] ,
    \Tile_X2Y4_WW4BEG[11] ,
    \Tile_X2Y4_WW4BEG[10] ,
    \Tile_X2Y4_WW4BEG[9] ,
    \Tile_X2Y4_WW4BEG[8] ,
    \Tile_X2Y4_WW4BEG[7] ,
    \Tile_X2Y4_WW4BEG[6] ,
    \Tile_X2Y4_WW4BEG[5] ,
    \Tile_X2Y4_WW4BEG[4] ,
    \Tile_X2Y4_WW4BEG[3] ,
    \Tile_X2Y4_WW4BEG[2] ,
    \Tile_X2Y4_WW4BEG[1] ,
    \Tile_X2Y4_WW4BEG[0] }),
    .WW4END({\Tile_X3Y4_WW4BEG[15] ,
    \Tile_X3Y4_WW4BEG[14] ,
    \Tile_X3Y4_WW4BEG[13] ,
    \Tile_X3Y4_WW4BEG[12] ,
    \Tile_X3Y4_WW4BEG[11] ,
    \Tile_X3Y4_WW4BEG[10] ,
    \Tile_X3Y4_WW4BEG[9] ,
    \Tile_X3Y4_WW4BEG[8] ,
    \Tile_X3Y4_WW4BEG[7] ,
    \Tile_X3Y4_WW4BEG[6] ,
    \Tile_X3Y4_WW4BEG[5] ,
    \Tile_X3Y4_WW4BEG[4] ,
    \Tile_X3Y4_WW4BEG[3] ,
    \Tile_X3Y4_WW4BEG[2] ,
    \Tile_X3Y4_WW4BEG[1] ,
    \Tile_X3Y4_WW4BEG[0] }));
 LUT4AB Tile_X2Y5_LUT4AB (.Ci(Tile_X2Y6_Co),
    .Co(Tile_X2Y5_Co),
    .UserCLK(Tile_X2Y6_UserCLKo),
    .UserCLKo(Tile_X2Y5_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X2Y5_E1BEG[3] ,
    \Tile_X2Y5_E1BEG[2] ,
    \Tile_X2Y5_E1BEG[1] ,
    \Tile_X2Y5_E1BEG[0] }),
    .E1END({\Tile_X1Y5_E1BEG[3] ,
    \Tile_X1Y5_E1BEG[2] ,
    \Tile_X1Y5_E1BEG[1] ,
    \Tile_X1Y5_E1BEG[0] }),
    .E2BEG({\Tile_X2Y5_E2BEG[7] ,
    \Tile_X2Y5_E2BEG[6] ,
    \Tile_X2Y5_E2BEG[5] ,
    \Tile_X2Y5_E2BEG[4] ,
    \Tile_X2Y5_E2BEG[3] ,
    \Tile_X2Y5_E2BEG[2] ,
    \Tile_X2Y5_E2BEG[1] ,
    \Tile_X2Y5_E2BEG[0] }),
    .E2BEGb({\Tile_X2Y5_E2BEGb[7] ,
    \Tile_X2Y5_E2BEGb[6] ,
    \Tile_X2Y5_E2BEGb[5] ,
    \Tile_X2Y5_E2BEGb[4] ,
    \Tile_X2Y5_E2BEGb[3] ,
    \Tile_X2Y5_E2BEGb[2] ,
    \Tile_X2Y5_E2BEGb[1] ,
    \Tile_X2Y5_E2BEGb[0] }),
    .E2END({\Tile_X1Y5_E2BEGb[7] ,
    \Tile_X1Y5_E2BEGb[6] ,
    \Tile_X1Y5_E2BEGb[5] ,
    \Tile_X1Y5_E2BEGb[4] ,
    \Tile_X1Y5_E2BEGb[3] ,
    \Tile_X1Y5_E2BEGb[2] ,
    \Tile_X1Y5_E2BEGb[1] ,
    \Tile_X1Y5_E2BEGb[0] }),
    .E2MID({\Tile_X1Y5_E2BEG[7] ,
    \Tile_X1Y5_E2BEG[6] ,
    \Tile_X1Y5_E2BEG[5] ,
    \Tile_X1Y5_E2BEG[4] ,
    \Tile_X1Y5_E2BEG[3] ,
    \Tile_X1Y5_E2BEG[2] ,
    \Tile_X1Y5_E2BEG[1] ,
    \Tile_X1Y5_E2BEG[0] }),
    .E6BEG({\Tile_X2Y5_E6BEG[11] ,
    \Tile_X2Y5_E6BEG[10] ,
    \Tile_X2Y5_E6BEG[9] ,
    \Tile_X2Y5_E6BEG[8] ,
    \Tile_X2Y5_E6BEG[7] ,
    \Tile_X2Y5_E6BEG[6] ,
    \Tile_X2Y5_E6BEG[5] ,
    \Tile_X2Y5_E6BEG[4] ,
    \Tile_X2Y5_E6BEG[3] ,
    \Tile_X2Y5_E6BEG[2] ,
    \Tile_X2Y5_E6BEG[1] ,
    \Tile_X2Y5_E6BEG[0] }),
    .E6END({\Tile_X1Y5_E6BEG[11] ,
    \Tile_X1Y5_E6BEG[10] ,
    \Tile_X1Y5_E6BEG[9] ,
    \Tile_X1Y5_E6BEG[8] ,
    \Tile_X1Y5_E6BEG[7] ,
    \Tile_X1Y5_E6BEG[6] ,
    \Tile_X1Y5_E6BEG[5] ,
    \Tile_X1Y5_E6BEG[4] ,
    \Tile_X1Y5_E6BEG[3] ,
    \Tile_X1Y5_E6BEG[2] ,
    \Tile_X1Y5_E6BEG[1] ,
    \Tile_X1Y5_E6BEG[0] }),
    .EE4BEG({\Tile_X2Y5_EE4BEG[15] ,
    \Tile_X2Y5_EE4BEG[14] ,
    \Tile_X2Y5_EE4BEG[13] ,
    \Tile_X2Y5_EE4BEG[12] ,
    \Tile_X2Y5_EE4BEG[11] ,
    \Tile_X2Y5_EE4BEG[10] ,
    \Tile_X2Y5_EE4BEG[9] ,
    \Tile_X2Y5_EE4BEG[8] ,
    \Tile_X2Y5_EE4BEG[7] ,
    \Tile_X2Y5_EE4BEG[6] ,
    \Tile_X2Y5_EE4BEG[5] ,
    \Tile_X2Y5_EE4BEG[4] ,
    \Tile_X2Y5_EE4BEG[3] ,
    \Tile_X2Y5_EE4BEG[2] ,
    \Tile_X2Y5_EE4BEG[1] ,
    \Tile_X2Y5_EE4BEG[0] }),
    .EE4END({\Tile_X1Y5_EE4BEG[15] ,
    \Tile_X1Y5_EE4BEG[14] ,
    \Tile_X1Y5_EE4BEG[13] ,
    \Tile_X1Y5_EE4BEG[12] ,
    \Tile_X1Y5_EE4BEG[11] ,
    \Tile_X1Y5_EE4BEG[10] ,
    \Tile_X1Y5_EE4BEG[9] ,
    \Tile_X1Y5_EE4BEG[8] ,
    \Tile_X1Y5_EE4BEG[7] ,
    \Tile_X1Y5_EE4BEG[6] ,
    \Tile_X1Y5_EE4BEG[5] ,
    \Tile_X1Y5_EE4BEG[4] ,
    \Tile_X1Y5_EE4BEG[3] ,
    \Tile_X1Y5_EE4BEG[2] ,
    \Tile_X1Y5_EE4BEG[1] ,
    \Tile_X1Y5_EE4BEG[0] }),
    .FrameData({\Tile_X1Y5_FrameData_O[31] ,
    \Tile_X1Y5_FrameData_O[30] ,
    \Tile_X1Y5_FrameData_O[29] ,
    \Tile_X1Y5_FrameData_O[28] ,
    \Tile_X1Y5_FrameData_O[27] ,
    \Tile_X1Y5_FrameData_O[26] ,
    \Tile_X1Y5_FrameData_O[25] ,
    \Tile_X1Y5_FrameData_O[24] ,
    \Tile_X1Y5_FrameData_O[23] ,
    \Tile_X1Y5_FrameData_O[22] ,
    \Tile_X1Y5_FrameData_O[21] ,
    \Tile_X1Y5_FrameData_O[20] ,
    \Tile_X1Y5_FrameData_O[19] ,
    \Tile_X1Y5_FrameData_O[18] ,
    \Tile_X1Y5_FrameData_O[17] ,
    \Tile_X1Y5_FrameData_O[16] ,
    \Tile_X1Y5_FrameData_O[15] ,
    \Tile_X1Y5_FrameData_O[14] ,
    \Tile_X1Y5_FrameData_O[13] ,
    \Tile_X1Y5_FrameData_O[12] ,
    \Tile_X1Y5_FrameData_O[11] ,
    \Tile_X1Y5_FrameData_O[10] ,
    \Tile_X1Y5_FrameData_O[9] ,
    \Tile_X1Y5_FrameData_O[8] ,
    \Tile_X1Y5_FrameData_O[7] ,
    \Tile_X1Y5_FrameData_O[6] ,
    \Tile_X1Y5_FrameData_O[5] ,
    \Tile_X1Y5_FrameData_O[4] ,
    \Tile_X1Y5_FrameData_O[3] ,
    \Tile_X1Y5_FrameData_O[2] ,
    \Tile_X1Y5_FrameData_O[1] ,
    \Tile_X1Y5_FrameData_O[0] }),
    .FrameData_O({\Tile_X2Y5_FrameData_O[31] ,
    \Tile_X2Y5_FrameData_O[30] ,
    \Tile_X2Y5_FrameData_O[29] ,
    \Tile_X2Y5_FrameData_O[28] ,
    \Tile_X2Y5_FrameData_O[27] ,
    \Tile_X2Y5_FrameData_O[26] ,
    \Tile_X2Y5_FrameData_O[25] ,
    \Tile_X2Y5_FrameData_O[24] ,
    \Tile_X2Y5_FrameData_O[23] ,
    \Tile_X2Y5_FrameData_O[22] ,
    \Tile_X2Y5_FrameData_O[21] ,
    \Tile_X2Y5_FrameData_O[20] ,
    \Tile_X2Y5_FrameData_O[19] ,
    \Tile_X2Y5_FrameData_O[18] ,
    \Tile_X2Y5_FrameData_O[17] ,
    \Tile_X2Y5_FrameData_O[16] ,
    \Tile_X2Y5_FrameData_O[15] ,
    \Tile_X2Y5_FrameData_O[14] ,
    \Tile_X2Y5_FrameData_O[13] ,
    \Tile_X2Y5_FrameData_O[12] ,
    \Tile_X2Y5_FrameData_O[11] ,
    \Tile_X2Y5_FrameData_O[10] ,
    \Tile_X2Y5_FrameData_O[9] ,
    \Tile_X2Y5_FrameData_O[8] ,
    \Tile_X2Y5_FrameData_O[7] ,
    \Tile_X2Y5_FrameData_O[6] ,
    \Tile_X2Y5_FrameData_O[5] ,
    \Tile_X2Y5_FrameData_O[4] ,
    \Tile_X2Y5_FrameData_O[3] ,
    \Tile_X2Y5_FrameData_O[2] ,
    \Tile_X2Y5_FrameData_O[1] ,
    \Tile_X2Y5_FrameData_O[0] }),
    .FrameStrobe({\Tile_X2Y6_FrameStrobe_O[19] ,
    \Tile_X2Y6_FrameStrobe_O[18] ,
    \Tile_X2Y6_FrameStrobe_O[17] ,
    \Tile_X2Y6_FrameStrobe_O[16] ,
    \Tile_X2Y6_FrameStrobe_O[15] ,
    \Tile_X2Y6_FrameStrobe_O[14] ,
    \Tile_X2Y6_FrameStrobe_O[13] ,
    \Tile_X2Y6_FrameStrobe_O[12] ,
    \Tile_X2Y6_FrameStrobe_O[11] ,
    \Tile_X2Y6_FrameStrobe_O[10] ,
    \Tile_X2Y6_FrameStrobe_O[9] ,
    \Tile_X2Y6_FrameStrobe_O[8] ,
    \Tile_X2Y6_FrameStrobe_O[7] ,
    \Tile_X2Y6_FrameStrobe_O[6] ,
    \Tile_X2Y6_FrameStrobe_O[5] ,
    \Tile_X2Y6_FrameStrobe_O[4] ,
    \Tile_X2Y6_FrameStrobe_O[3] ,
    \Tile_X2Y6_FrameStrobe_O[2] ,
    \Tile_X2Y6_FrameStrobe_O[1] ,
    \Tile_X2Y6_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X2Y5_FrameStrobe_O[19] ,
    \Tile_X2Y5_FrameStrobe_O[18] ,
    \Tile_X2Y5_FrameStrobe_O[17] ,
    \Tile_X2Y5_FrameStrobe_O[16] ,
    \Tile_X2Y5_FrameStrobe_O[15] ,
    \Tile_X2Y5_FrameStrobe_O[14] ,
    \Tile_X2Y5_FrameStrobe_O[13] ,
    \Tile_X2Y5_FrameStrobe_O[12] ,
    \Tile_X2Y5_FrameStrobe_O[11] ,
    \Tile_X2Y5_FrameStrobe_O[10] ,
    \Tile_X2Y5_FrameStrobe_O[9] ,
    \Tile_X2Y5_FrameStrobe_O[8] ,
    \Tile_X2Y5_FrameStrobe_O[7] ,
    \Tile_X2Y5_FrameStrobe_O[6] ,
    \Tile_X2Y5_FrameStrobe_O[5] ,
    \Tile_X2Y5_FrameStrobe_O[4] ,
    \Tile_X2Y5_FrameStrobe_O[3] ,
    \Tile_X2Y5_FrameStrobe_O[2] ,
    \Tile_X2Y5_FrameStrobe_O[1] ,
    \Tile_X2Y5_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X2Y5_N1BEG[3] ,
    \Tile_X2Y5_N1BEG[2] ,
    \Tile_X2Y5_N1BEG[1] ,
    \Tile_X2Y5_N1BEG[0] }),
    .N1END({\Tile_X2Y6_N1BEG[3] ,
    \Tile_X2Y6_N1BEG[2] ,
    \Tile_X2Y6_N1BEG[1] ,
    \Tile_X2Y6_N1BEG[0] }),
    .N2BEG({\Tile_X2Y5_N2BEG[7] ,
    \Tile_X2Y5_N2BEG[6] ,
    \Tile_X2Y5_N2BEG[5] ,
    \Tile_X2Y5_N2BEG[4] ,
    \Tile_X2Y5_N2BEG[3] ,
    \Tile_X2Y5_N2BEG[2] ,
    \Tile_X2Y5_N2BEG[1] ,
    \Tile_X2Y5_N2BEG[0] }),
    .N2BEGb({\Tile_X2Y5_N2BEGb[7] ,
    \Tile_X2Y5_N2BEGb[6] ,
    \Tile_X2Y5_N2BEGb[5] ,
    \Tile_X2Y5_N2BEGb[4] ,
    \Tile_X2Y5_N2BEGb[3] ,
    \Tile_X2Y5_N2BEGb[2] ,
    \Tile_X2Y5_N2BEGb[1] ,
    \Tile_X2Y5_N2BEGb[0] }),
    .N2END({\Tile_X2Y6_N2BEGb[7] ,
    \Tile_X2Y6_N2BEGb[6] ,
    \Tile_X2Y6_N2BEGb[5] ,
    \Tile_X2Y6_N2BEGb[4] ,
    \Tile_X2Y6_N2BEGb[3] ,
    \Tile_X2Y6_N2BEGb[2] ,
    \Tile_X2Y6_N2BEGb[1] ,
    \Tile_X2Y6_N2BEGb[0] }),
    .N2MID({\Tile_X2Y6_N2BEG[7] ,
    \Tile_X2Y6_N2BEG[6] ,
    \Tile_X2Y6_N2BEG[5] ,
    \Tile_X2Y6_N2BEG[4] ,
    \Tile_X2Y6_N2BEG[3] ,
    \Tile_X2Y6_N2BEG[2] ,
    \Tile_X2Y6_N2BEG[1] ,
    \Tile_X2Y6_N2BEG[0] }),
    .N4BEG({\Tile_X2Y5_N4BEG[15] ,
    \Tile_X2Y5_N4BEG[14] ,
    \Tile_X2Y5_N4BEG[13] ,
    \Tile_X2Y5_N4BEG[12] ,
    \Tile_X2Y5_N4BEG[11] ,
    \Tile_X2Y5_N4BEG[10] ,
    \Tile_X2Y5_N4BEG[9] ,
    \Tile_X2Y5_N4BEG[8] ,
    \Tile_X2Y5_N4BEG[7] ,
    \Tile_X2Y5_N4BEG[6] ,
    \Tile_X2Y5_N4BEG[5] ,
    \Tile_X2Y5_N4BEG[4] ,
    \Tile_X2Y5_N4BEG[3] ,
    \Tile_X2Y5_N4BEG[2] ,
    \Tile_X2Y5_N4BEG[1] ,
    \Tile_X2Y5_N4BEG[0] }),
    .N4END({\Tile_X2Y6_N4BEG[15] ,
    \Tile_X2Y6_N4BEG[14] ,
    \Tile_X2Y6_N4BEG[13] ,
    \Tile_X2Y6_N4BEG[12] ,
    \Tile_X2Y6_N4BEG[11] ,
    \Tile_X2Y6_N4BEG[10] ,
    \Tile_X2Y6_N4BEG[9] ,
    \Tile_X2Y6_N4BEG[8] ,
    \Tile_X2Y6_N4BEG[7] ,
    \Tile_X2Y6_N4BEG[6] ,
    \Tile_X2Y6_N4BEG[5] ,
    \Tile_X2Y6_N4BEG[4] ,
    \Tile_X2Y6_N4BEG[3] ,
    \Tile_X2Y6_N4BEG[2] ,
    \Tile_X2Y6_N4BEG[1] ,
    \Tile_X2Y6_N4BEG[0] }),
    .NN4BEG({\Tile_X2Y5_NN4BEG[15] ,
    \Tile_X2Y5_NN4BEG[14] ,
    \Tile_X2Y5_NN4BEG[13] ,
    \Tile_X2Y5_NN4BEG[12] ,
    \Tile_X2Y5_NN4BEG[11] ,
    \Tile_X2Y5_NN4BEG[10] ,
    \Tile_X2Y5_NN4BEG[9] ,
    \Tile_X2Y5_NN4BEG[8] ,
    \Tile_X2Y5_NN4BEG[7] ,
    \Tile_X2Y5_NN4BEG[6] ,
    \Tile_X2Y5_NN4BEG[5] ,
    \Tile_X2Y5_NN4BEG[4] ,
    \Tile_X2Y5_NN4BEG[3] ,
    \Tile_X2Y5_NN4BEG[2] ,
    \Tile_X2Y5_NN4BEG[1] ,
    \Tile_X2Y5_NN4BEG[0] }),
    .NN4END({\Tile_X2Y6_NN4BEG[15] ,
    \Tile_X2Y6_NN4BEG[14] ,
    \Tile_X2Y6_NN4BEG[13] ,
    \Tile_X2Y6_NN4BEG[12] ,
    \Tile_X2Y6_NN4BEG[11] ,
    \Tile_X2Y6_NN4BEG[10] ,
    \Tile_X2Y6_NN4BEG[9] ,
    \Tile_X2Y6_NN4BEG[8] ,
    \Tile_X2Y6_NN4BEG[7] ,
    \Tile_X2Y6_NN4BEG[6] ,
    \Tile_X2Y6_NN4BEG[5] ,
    \Tile_X2Y6_NN4BEG[4] ,
    \Tile_X2Y6_NN4BEG[3] ,
    \Tile_X2Y6_NN4BEG[2] ,
    \Tile_X2Y6_NN4BEG[1] ,
    \Tile_X2Y6_NN4BEG[0] }),
    .S1BEG({\Tile_X2Y5_S1BEG[3] ,
    \Tile_X2Y5_S1BEG[2] ,
    \Tile_X2Y5_S1BEG[1] ,
    \Tile_X2Y5_S1BEG[0] }),
    .S1END({\Tile_X2Y4_S1BEG[3] ,
    \Tile_X2Y4_S1BEG[2] ,
    \Tile_X2Y4_S1BEG[1] ,
    \Tile_X2Y4_S1BEG[0] }),
    .S2BEG({\Tile_X2Y5_S2BEG[7] ,
    \Tile_X2Y5_S2BEG[6] ,
    \Tile_X2Y5_S2BEG[5] ,
    \Tile_X2Y5_S2BEG[4] ,
    \Tile_X2Y5_S2BEG[3] ,
    \Tile_X2Y5_S2BEG[2] ,
    \Tile_X2Y5_S2BEG[1] ,
    \Tile_X2Y5_S2BEG[0] }),
    .S2BEGb({\Tile_X2Y5_S2BEGb[7] ,
    \Tile_X2Y5_S2BEGb[6] ,
    \Tile_X2Y5_S2BEGb[5] ,
    \Tile_X2Y5_S2BEGb[4] ,
    \Tile_X2Y5_S2BEGb[3] ,
    \Tile_X2Y5_S2BEGb[2] ,
    \Tile_X2Y5_S2BEGb[1] ,
    \Tile_X2Y5_S2BEGb[0] }),
    .S2END({\Tile_X2Y4_S2BEGb[7] ,
    \Tile_X2Y4_S2BEGb[6] ,
    \Tile_X2Y4_S2BEGb[5] ,
    \Tile_X2Y4_S2BEGb[4] ,
    \Tile_X2Y4_S2BEGb[3] ,
    \Tile_X2Y4_S2BEGb[2] ,
    \Tile_X2Y4_S2BEGb[1] ,
    \Tile_X2Y4_S2BEGb[0] }),
    .S2MID({\Tile_X2Y4_S2BEG[7] ,
    \Tile_X2Y4_S2BEG[6] ,
    \Tile_X2Y4_S2BEG[5] ,
    \Tile_X2Y4_S2BEG[4] ,
    \Tile_X2Y4_S2BEG[3] ,
    \Tile_X2Y4_S2BEG[2] ,
    \Tile_X2Y4_S2BEG[1] ,
    \Tile_X2Y4_S2BEG[0] }),
    .S4BEG({\Tile_X2Y5_S4BEG[15] ,
    \Tile_X2Y5_S4BEG[14] ,
    \Tile_X2Y5_S4BEG[13] ,
    \Tile_X2Y5_S4BEG[12] ,
    \Tile_X2Y5_S4BEG[11] ,
    \Tile_X2Y5_S4BEG[10] ,
    \Tile_X2Y5_S4BEG[9] ,
    \Tile_X2Y5_S4BEG[8] ,
    \Tile_X2Y5_S4BEG[7] ,
    \Tile_X2Y5_S4BEG[6] ,
    \Tile_X2Y5_S4BEG[5] ,
    \Tile_X2Y5_S4BEG[4] ,
    \Tile_X2Y5_S4BEG[3] ,
    \Tile_X2Y5_S4BEG[2] ,
    \Tile_X2Y5_S4BEG[1] ,
    \Tile_X2Y5_S4BEG[0] }),
    .S4END({\Tile_X2Y4_S4BEG[15] ,
    \Tile_X2Y4_S4BEG[14] ,
    \Tile_X2Y4_S4BEG[13] ,
    \Tile_X2Y4_S4BEG[12] ,
    \Tile_X2Y4_S4BEG[11] ,
    \Tile_X2Y4_S4BEG[10] ,
    \Tile_X2Y4_S4BEG[9] ,
    \Tile_X2Y4_S4BEG[8] ,
    \Tile_X2Y4_S4BEG[7] ,
    \Tile_X2Y4_S4BEG[6] ,
    \Tile_X2Y4_S4BEG[5] ,
    \Tile_X2Y4_S4BEG[4] ,
    \Tile_X2Y4_S4BEG[3] ,
    \Tile_X2Y4_S4BEG[2] ,
    \Tile_X2Y4_S4BEG[1] ,
    \Tile_X2Y4_S4BEG[0] }),
    .SS4BEG({\Tile_X2Y5_SS4BEG[15] ,
    \Tile_X2Y5_SS4BEG[14] ,
    \Tile_X2Y5_SS4BEG[13] ,
    \Tile_X2Y5_SS4BEG[12] ,
    \Tile_X2Y5_SS4BEG[11] ,
    \Tile_X2Y5_SS4BEG[10] ,
    \Tile_X2Y5_SS4BEG[9] ,
    \Tile_X2Y5_SS4BEG[8] ,
    \Tile_X2Y5_SS4BEG[7] ,
    \Tile_X2Y5_SS4BEG[6] ,
    \Tile_X2Y5_SS4BEG[5] ,
    \Tile_X2Y5_SS4BEG[4] ,
    \Tile_X2Y5_SS4BEG[3] ,
    \Tile_X2Y5_SS4BEG[2] ,
    \Tile_X2Y5_SS4BEG[1] ,
    \Tile_X2Y5_SS4BEG[0] }),
    .SS4END({\Tile_X2Y4_SS4BEG[15] ,
    \Tile_X2Y4_SS4BEG[14] ,
    \Tile_X2Y4_SS4BEG[13] ,
    \Tile_X2Y4_SS4BEG[12] ,
    \Tile_X2Y4_SS4BEG[11] ,
    \Tile_X2Y4_SS4BEG[10] ,
    \Tile_X2Y4_SS4BEG[9] ,
    \Tile_X2Y4_SS4BEG[8] ,
    \Tile_X2Y4_SS4BEG[7] ,
    \Tile_X2Y4_SS4BEG[6] ,
    \Tile_X2Y4_SS4BEG[5] ,
    \Tile_X2Y4_SS4BEG[4] ,
    \Tile_X2Y4_SS4BEG[3] ,
    \Tile_X2Y4_SS4BEG[2] ,
    \Tile_X2Y4_SS4BEG[1] ,
    \Tile_X2Y4_SS4BEG[0] }),
    .W1BEG({\Tile_X2Y5_W1BEG[3] ,
    \Tile_X2Y5_W1BEG[2] ,
    \Tile_X2Y5_W1BEG[1] ,
    \Tile_X2Y5_W1BEG[0] }),
    .W1END({\Tile_X3Y5_W1BEG[3] ,
    \Tile_X3Y5_W1BEG[2] ,
    \Tile_X3Y5_W1BEG[1] ,
    \Tile_X3Y5_W1BEG[0] }),
    .W2BEG({\Tile_X2Y5_W2BEG[7] ,
    \Tile_X2Y5_W2BEG[6] ,
    \Tile_X2Y5_W2BEG[5] ,
    \Tile_X2Y5_W2BEG[4] ,
    \Tile_X2Y5_W2BEG[3] ,
    \Tile_X2Y5_W2BEG[2] ,
    \Tile_X2Y5_W2BEG[1] ,
    \Tile_X2Y5_W2BEG[0] }),
    .W2BEGb({\Tile_X2Y5_W2BEGb[7] ,
    \Tile_X2Y5_W2BEGb[6] ,
    \Tile_X2Y5_W2BEGb[5] ,
    \Tile_X2Y5_W2BEGb[4] ,
    \Tile_X2Y5_W2BEGb[3] ,
    \Tile_X2Y5_W2BEGb[2] ,
    \Tile_X2Y5_W2BEGb[1] ,
    \Tile_X2Y5_W2BEGb[0] }),
    .W2END({\Tile_X3Y5_W2BEGb[7] ,
    \Tile_X3Y5_W2BEGb[6] ,
    \Tile_X3Y5_W2BEGb[5] ,
    \Tile_X3Y5_W2BEGb[4] ,
    \Tile_X3Y5_W2BEGb[3] ,
    \Tile_X3Y5_W2BEGb[2] ,
    \Tile_X3Y5_W2BEGb[1] ,
    \Tile_X3Y5_W2BEGb[0] }),
    .W2MID({\Tile_X3Y5_W2BEG[7] ,
    \Tile_X3Y5_W2BEG[6] ,
    \Tile_X3Y5_W2BEG[5] ,
    \Tile_X3Y5_W2BEG[4] ,
    \Tile_X3Y5_W2BEG[3] ,
    \Tile_X3Y5_W2BEG[2] ,
    \Tile_X3Y5_W2BEG[1] ,
    \Tile_X3Y5_W2BEG[0] }),
    .W6BEG({\Tile_X2Y5_W6BEG[11] ,
    \Tile_X2Y5_W6BEG[10] ,
    \Tile_X2Y5_W6BEG[9] ,
    \Tile_X2Y5_W6BEG[8] ,
    \Tile_X2Y5_W6BEG[7] ,
    \Tile_X2Y5_W6BEG[6] ,
    \Tile_X2Y5_W6BEG[5] ,
    \Tile_X2Y5_W6BEG[4] ,
    \Tile_X2Y5_W6BEG[3] ,
    \Tile_X2Y5_W6BEG[2] ,
    \Tile_X2Y5_W6BEG[1] ,
    \Tile_X2Y5_W6BEG[0] }),
    .W6END({\Tile_X3Y5_W6BEG[11] ,
    \Tile_X3Y5_W6BEG[10] ,
    \Tile_X3Y5_W6BEG[9] ,
    \Tile_X3Y5_W6BEG[8] ,
    \Tile_X3Y5_W6BEG[7] ,
    \Tile_X3Y5_W6BEG[6] ,
    \Tile_X3Y5_W6BEG[5] ,
    \Tile_X3Y5_W6BEG[4] ,
    \Tile_X3Y5_W6BEG[3] ,
    \Tile_X3Y5_W6BEG[2] ,
    \Tile_X3Y5_W6BEG[1] ,
    \Tile_X3Y5_W6BEG[0] }),
    .WW4BEG({\Tile_X2Y5_WW4BEG[15] ,
    \Tile_X2Y5_WW4BEG[14] ,
    \Tile_X2Y5_WW4BEG[13] ,
    \Tile_X2Y5_WW4BEG[12] ,
    \Tile_X2Y5_WW4BEG[11] ,
    \Tile_X2Y5_WW4BEG[10] ,
    \Tile_X2Y5_WW4BEG[9] ,
    \Tile_X2Y5_WW4BEG[8] ,
    \Tile_X2Y5_WW4BEG[7] ,
    \Tile_X2Y5_WW4BEG[6] ,
    \Tile_X2Y5_WW4BEG[5] ,
    \Tile_X2Y5_WW4BEG[4] ,
    \Tile_X2Y5_WW4BEG[3] ,
    \Tile_X2Y5_WW4BEG[2] ,
    \Tile_X2Y5_WW4BEG[1] ,
    \Tile_X2Y5_WW4BEG[0] }),
    .WW4END({\Tile_X3Y5_WW4BEG[15] ,
    \Tile_X3Y5_WW4BEG[14] ,
    \Tile_X3Y5_WW4BEG[13] ,
    \Tile_X3Y5_WW4BEG[12] ,
    \Tile_X3Y5_WW4BEG[11] ,
    \Tile_X3Y5_WW4BEG[10] ,
    \Tile_X3Y5_WW4BEG[9] ,
    \Tile_X3Y5_WW4BEG[8] ,
    \Tile_X3Y5_WW4BEG[7] ,
    \Tile_X3Y5_WW4BEG[6] ,
    \Tile_X3Y5_WW4BEG[5] ,
    \Tile_X3Y5_WW4BEG[4] ,
    \Tile_X3Y5_WW4BEG[3] ,
    \Tile_X3Y5_WW4BEG[2] ,
    \Tile_X3Y5_WW4BEG[1] ,
    \Tile_X3Y5_WW4BEG[0] }));
 LUT4AB Tile_X2Y6_LUT4AB (.Ci(Tile_X2Y7_Co),
    .Co(Tile_X2Y6_Co),
    .UserCLK(Tile_X2Y7_UserCLKo),
    .UserCLKo(Tile_X2Y6_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X2Y6_E1BEG[3] ,
    \Tile_X2Y6_E1BEG[2] ,
    \Tile_X2Y6_E1BEG[1] ,
    \Tile_X2Y6_E1BEG[0] }),
    .E1END({\Tile_X1Y6_E1BEG[3] ,
    \Tile_X1Y6_E1BEG[2] ,
    \Tile_X1Y6_E1BEG[1] ,
    \Tile_X1Y6_E1BEG[0] }),
    .E2BEG({\Tile_X2Y6_E2BEG[7] ,
    \Tile_X2Y6_E2BEG[6] ,
    \Tile_X2Y6_E2BEG[5] ,
    \Tile_X2Y6_E2BEG[4] ,
    \Tile_X2Y6_E2BEG[3] ,
    \Tile_X2Y6_E2BEG[2] ,
    \Tile_X2Y6_E2BEG[1] ,
    \Tile_X2Y6_E2BEG[0] }),
    .E2BEGb({\Tile_X2Y6_E2BEGb[7] ,
    \Tile_X2Y6_E2BEGb[6] ,
    \Tile_X2Y6_E2BEGb[5] ,
    \Tile_X2Y6_E2BEGb[4] ,
    \Tile_X2Y6_E2BEGb[3] ,
    \Tile_X2Y6_E2BEGb[2] ,
    \Tile_X2Y6_E2BEGb[1] ,
    \Tile_X2Y6_E2BEGb[0] }),
    .E2END({\Tile_X1Y6_E2BEGb[7] ,
    \Tile_X1Y6_E2BEGb[6] ,
    \Tile_X1Y6_E2BEGb[5] ,
    \Tile_X1Y6_E2BEGb[4] ,
    \Tile_X1Y6_E2BEGb[3] ,
    \Tile_X1Y6_E2BEGb[2] ,
    \Tile_X1Y6_E2BEGb[1] ,
    \Tile_X1Y6_E2BEGb[0] }),
    .E2MID({\Tile_X1Y6_E2BEG[7] ,
    \Tile_X1Y6_E2BEG[6] ,
    \Tile_X1Y6_E2BEG[5] ,
    \Tile_X1Y6_E2BEG[4] ,
    \Tile_X1Y6_E2BEG[3] ,
    \Tile_X1Y6_E2BEG[2] ,
    \Tile_X1Y6_E2BEG[1] ,
    \Tile_X1Y6_E2BEG[0] }),
    .E6BEG({\Tile_X2Y6_E6BEG[11] ,
    \Tile_X2Y6_E6BEG[10] ,
    \Tile_X2Y6_E6BEG[9] ,
    \Tile_X2Y6_E6BEG[8] ,
    \Tile_X2Y6_E6BEG[7] ,
    \Tile_X2Y6_E6BEG[6] ,
    \Tile_X2Y6_E6BEG[5] ,
    \Tile_X2Y6_E6BEG[4] ,
    \Tile_X2Y6_E6BEG[3] ,
    \Tile_X2Y6_E6BEG[2] ,
    \Tile_X2Y6_E6BEG[1] ,
    \Tile_X2Y6_E6BEG[0] }),
    .E6END({\Tile_X1Y6_E6BEG[11] ,
    \Tile_X1Y6_E6BEG[10] ,
    \Tile_X1Y6_E6BEG[9] ,
    \Tile_X1Y6_E6BEG[8] ,
    \Tile_X1Y6_E6BEG[7] ,
    \Tile_X1Y6_E6BEG[6] ,
    \Tile_X1Y6_E6BEG[5] ,
    \Tile_X1Y6_E6BEG[4] ,
    \Tile_X1Y6_E6BEG[3] ,
    \Tile_X1Y6_E6BEG[2] ,
    \Tile_X1Y6_E6BEG[1] ,
    \Tile_X1Y6_E6BEG[0] }),
    .EE4BEG({\Tile_X2Y6_EE4BEG[15] ,
    \Tile_X2Y6_EE4BEG[14] ,
    \Tile_X2Y6_EE4BEG[13] ,
    \Tile_X2Y6_EE4BEG[12] ,
    \Tile_X2Y6_EE4BEG[11] ,
    \Tile_X2Y6_EE4BEG[10] ,
    \Tile_X2Y6_EE4BEG[9] ,
    \Tile_X2Y6_EE4BEG[8] ,
    \Tile_X2Y6_EE4BEG[7] ,
    \Tile_X2Y6_EE4BEG[6] ,
    \Tile_X2Y6_EE4BEG[5] ,
    \Tile_X2Y6_EE4BEG[4] ,
    \Tile_X2Y6_EE4BEG[3] ,
    \Tile_X2Y6_EE4BEG[2] ,
    \Tile_X2Y6_EE4BEG[1] ,
    \Tile_X2Y6_EE4BEG[0] }),
    .EE4END({\Tile_X1Y6_EE4BEG[15] ,
    \Tile_X1Y6_EE4BEG[14] ,
    \Tile_X1Y6_EE4BEG[13] ,
    \Tile_X1Y6_EE4BEG[12] ,
    \Tile_X1Y6_EE4BEG[11] ,
    \Tile_X1Y6_EE4BEG[10] ,
    \Tile_X1Y6_EE4BEG[9] ,
    \Tile_X1Y6_EE4BEG[8] ,
    \Tile_X1Y6_EE4BEG[7] ,
    \Tile_X1Y6_EE4BEG[6] ,
    \Tile_X1Y6_EE4BEG[5] ,
    \Tile_X1Y6_EE4BEG[4] ,
    \Tile_X1Y6_EE4BEG[3] ,
    \Tile_X1Y6_EE4BEG[2] ,
    \Tile_X1Y6_EE4BEG[1] ,
    \Tile_X1Y6_EE4BEG[0] }),
    .FrameData({\Tile_X1Y6_FrameData_O[31] ,
    \Tile_X1Y6_FrameData_O[30] ,
    \Tile_X1Y6_FrameData_O[29] ,
    \Tile_X1Y6_FrameData_O[28] ,
    \Tile_X1Y6_FrameData_O[27] ,
    \Tile_X1Y6_FrameData_O[26] ,
    \Tile_X1Y6_FrameData_O[25] ,
    \Tile_X1Y6_FrameData_O[24] ,
    \Tile_X1Y6_FrameData_O[23] ,
    \Tile_X1Y6_FrameData_O[22] ,
    \Tile_X1Y6_FrameData_O[21] ,
    \Tile_X1Y6_FrameData_O[20] ,
    \Tile_X1Y6_FrameData_O[19] ,
    \Tile_X1Y6_FrameData_O[18] ,
    \Tile_X1Y6_FrameData_O[17] ,
    \Tile_X1Y6_FrameData_O[16] ,
    \Tile_X1Y6_FrameData_O[15] ,
    \Tile_X1Y6_FrameData_O[14] ,
    \Tile_X1Y6_FrameData_O[13] ,
    \Tile_X1Y6_FrameData_O[12] ,
    \Tile_X1Y6_FrameData_O[11] ,
    \Tile_X1Y6_FrameData_O[10] ,
    \Tile_X1Y6_FrameData_O[9] ,
    \Tile_X1Y6_FrameData_O[8] ,
    \Tile_X1Y6_FrameData_O[7] ,
    \Tile_X1Y6_FrameData_O[6] ,
    \Tile_X1Y6_FrameData_O[5] ,
    \Tile_X1Y6_FrameData_O[4] ,
    \Tile_X1Y6_FrameData_O[3] ,
    \Tile_X1Y6_FrameData_O[2] ,
    \Tile_X1Y6_FrameData_O[1] ,
    \Tile_X1Y6_FrameData_O[0] }),
    .FrameData_O({\Tile_X2Y6_FrameData_O[31] ,
    \Tile_X2Y6_FrameData_O[30] ,
    \Tile_X2Y6_FrameData_O[29] ,
    \Tile_X2Y6_FrameData_O[28] ,
    \Tile_X2Y6_FrameData_O[27] ,
    \Tile_X2Y6_FrameData_O[26] ,
    \Tile_X2Y6_FrameData_O[25] ,
    \Tile_X2Y6_FrameData_O[24] ,
    \Tile_X2Y6_FrameData_O[23] ,
    \Tile_X2Y6_FrameData_O[22] ,
    \Tile_X2Y6_FrameData_O[21] ,
    \Tile_X2Y6_FrameData_O[20] ,
    \Tile_X2Y6_FrameData_O[19] ,
    \Tile_X2Y6_FrameData_O[18] ,
    \Tile_X2Y6_FrameData_O[17] ,
    \Tile_X2Y6_FrameData_O[16] ,
    \Tile_X2Y6_FrameData_O[15] ,
    \Tile_X2Y6_FrameData_O[14] ,
    \Tile_X2Y6_FrameData_O[13] ,
    \Tile_X2Y6_FrameData_O[12] ,
    \Tile_X2Y6_FrameData_O[11] ,
    \Tile_X2Y6_FrameData_O[10] ,
    \Tile_X2Y6_FrameData_O[9] ,
    \Tile_X2Y6_FrameData_O[8] ,
    \Tile_X2Y6_FrameData_O[7] ,
    \Tile_X2Y6_FrameData_O[6] ,
    \Tile_X2Y6_FrameData_O[5] ,
    \Tile_X2Y6_FrameData_O[4] ,
    \Tile_X2Y6_FrameData_O[3] ,
    \Tile_X2Y6_FrameData_O[2] ,
    \Tile_X2Y6_FrameData_O[1] ,
    \Tile_X2Y6_FrameData_O[0] }),
    .FrameStrobe({\Tile_X2Y7_FrameStrobe_O[19] ,
    \Tile_X2Y7_FrameStrobe_O[18] ,
    \Tile_X2Y7_FrameStrobe_O[17] ,
    \Tile_X2Y7_FrameStrobe_O[16] ,
    \Tile_X2Y7_FrameStrobe_O[15] ,
    \Tile_X2Y7_FrameStrobe_O[14] ,
    \Tile_X2Y7_FrameStrobe_O[13] ,
    \Tile_X2Y7_FrameStrobe_O[12] ,
    \Tile_X2Y7_FrameStrobe_O[11] ,
    \Tile_X2Y7_FrameStrobe_O[10] ,
    \Tile_X2Y7_FrameStrobe_O[9] ,
    \Tile_X2Y7_FrameStrobe_O[8] ,
    \Tile_X2Y7_FrameStrobe_O[7] ,
    \Tile_X2Y7_FrameStrobe_O[6] ,
    \Tile_X2Y7_FrameStrobe_O[5] ,
    \Tile_X2Y7_FrameStrobe_O[4] ,
    \Tile_X2Y7_FrameStrobe_O[3] ,
    \Tile_X2Y7_FrameStrobe_O[2] ,
    \Tile_X2Y7_FrameStrobe_O[1] ,
    \Tile_X2Y7_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X2Y6_FrameStrobe_O[19] ,
    \Tile_X2Y6_FrameStrobe_O[18] ,
    \Tile_X2Y6_FrameStrobe_O[17] ,
    \Tile_X2Y6_FrameStrobe_O[16] ,
    \Tile_X2Y6_FrameStrobe_O[15] ,
    \Tile_X2Y6_FrameStrobe_O[14] ,
    \Tile_X2Y6_FrameStrobe_O[13] ,
    \Tile_X2Y6_FrameStrobe_O[12] ,
    \Tile_X2Y6_FrameStrobe_O[11] ,
    \Tile_X2Y6_FrameStrobe_O[10] ,
    \Tile_X2Y6_FrameStrobe_O[9] ,
    \Tile_X2Y6_FrameStrobe_O[8] ,
    \Tile_X2Y6_FrameStrobe_O[7] ,
    \Tile_X2Y6_FrameStrobe_O[6] ,
    \Tile_X2Y6_FrameStrobe_O[5] ,
    \Tile_X2Y6_FrameStrobe_O[4] ,
    \Tile_X2Y6_FrameStrobe_O[3] ,
    \Tile_X2Y6_FrameStrobe_O[2] ,
    \Tile_X2Y6_FrameStrobe_O[1] ,
    \Tile_X2Y6_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X2Y6_N1BEG[3] ,
    \Tile_X2Y6_N1BEG[2] ,
    \Tile_X2Y6_N1BEG[1] ,
    \Tile_X2Y6_N1BEG[0] }),
    .N1END({\Tile_X2Y7_N1BEG[3] ,
    \Tile_X2Y7_N1BEG[2] ,
    \Tile_X2Y7_N1BEG[1] ,
    \Tile_X2Y7_N1BEG[0] }),
    .N2BEG({\Tile_X2Y6_N2BEG[7] ,
    \Tile_X2Y6_N2BEG[6] ,
    \Tile_X2Y6_N2BEG[5] ,
    \Tile_X2Y6_N2BEG[4] ,
    \Tile_X2Y6_N2BEG[3] ,
    \Tile_X2Y6_N2BEG[2] ,
    \Tile_X2Y6_N2BEG[1] ,
    \Tile_X2Y6_N2BEG[0] }),
    .N2BEGb({\Tile_X2Y6_N2BEGb[7] ,
    \Tile_X2Y6_N2BEGb[6] ,
    \Tile_X2Y6_N2BEGb[5] ,
    \Tile_X2Y6_N2BEGb[4] ,
    \Tile_X2Y6_N2BEGb[3] ,
    \Tile_X2Y6_N2BEGb[2] ,
    \Tile_X2Y6_N2BEGb[1] ,
    \Tile_X2Y6_N2BEGb[0] }),
    .N2END({\Tile_X2Y7_N2BEGb[7] ,
    \Tile_X2Y7_N2BEGb[6] ,
    \Tile_X2Y7_N2BEGb[5] ,
    \Tile_X2Y7_N2BEGb[4] ,
    \Tile_X2Y7_N2BEGb[3] ,
    \Tile_X2Y7_N2BEGb[2] ,
    \Tile_X2Y7_N2BEGb[1] ,
    \Tile_X2Y7_N2BEGb[0] }),
    .N2MID({\Tile_X2Y7_N2BEG[7] ,
    \Tile_X2Y7_N2BEG[6] ,
    \Tile_X2Y7_N2BEG[5] ,
    \Tile_X2Y7_N2BEG[4] ,
    \Tile_X2Y7_N2BEG[3] ,
    \Tile_X2Y7_N2BEG[2] ,
    \Tile_X2Y7_N2BEG[1] ,
    \Tile_X2Y7_N2BEG[0] }),
    .N4BEG({\Tile_X2Y6_N4BEG[15] ,
    \Tile_X2Y6_N4BEG[14] ,
    \Tile_X2Y6_N4BEG[13] ,
    \Tile_X2Y6_N4BEG[12] ,
    \Tile_X2Y6_N4BEG[11] ,
    \Tile_X2Y6_N4BEG[10] ,
    \Tile_X2Y6_N4BEG[9] ,
    \Tile_X2Y6_N4BEG[8] ,
    \Tile_X2Y6_N4BEG[7] ,
    \Tile_X2Y6_N4BEG[6] ,
    \Tile_X2Y6_N4BEG[5] ,
    \Tile_X2Y6_N4BEG[4] ,
    \Tile_X2Y6_N4BEG[3] ,
    \Tile_X2Y6_N4BEG[2] ,
    \Tile_X2Y6_N4BEG[1] ,
    \Tile_X2Y6_N4BEG[0] }),
    .N4END({\Tile_X2Y7_N4BEG[15] ,
    \Tile_X2Y7_N4BEG[14] ,
    \Tile_X2Y7_N4BEG[13] ,
    \Tile_X2Y7_N4BEG[12] ,
    \Tile_X2Y7_N4BEG[11] ,
    \Tile_X2Y7_N4BEG[10] ,
    \Tile_X2Y7_N4BEG[9] ,
    \Tile_X2Y7_N4BEG[8] ,
    \Tile_X2Y7_N4BEG[7] ,
    \Tile_X2Y7_N4BEG[6] ,
    \Tile_X2Y7_N4BEG[5] ,
    \Tile_X2Y7_N4BEG[4] ,
    \Tile_X2Y7_N4BEG[3] ,
    \Tile_X2Y7_N4BEG[2] ,
    \Tile_X2Y7_N4BEG[1] ,
    \Tile_X2Y7_N4BEG[0] }),
    .NN4BEG({\Tile_X2Y6_NN4BEG[15] ,
    \Tile_X2Y6_NN4BEG[14] ,
    \Tile_X2Y6_NN4BEG[13] ,
    \Tile_X2Y6_NN4BEG[12] ,
    \Tile_X2Y6_NN4BEG[11] ,
    \Tile_X2Y6_NN4BEG[10] ,
    \Tile_X2Y6_NN4BEG[9] ,
    \Tile_X2Y6_NN4BEG[8] ,
    \Tile_X2Y6_NN4BEG[7] ,
    \Tile_X2Y6_NN4BEG[6] ,
    \Tile_X2Y6_NN4BEG[5] ,
    \Tile_X2Y6_NN4BEG[4] ,
    \Tile_X2Y6_NN4BEG[3] ,
    \Tile_X2Y6_NN4BEG[2] ,
    \Tile_X2Y6_NN4BEG[1] ,
    \Tile_X2Y6_NN4BEG[0] }),
    .NN4END({\Tile_X2Y7_NN4BEG[15] ,
    \Tile_X2Y7_NN4BEG[14] ,
    \Tile_X2Y7_NN4BEG[13] ,
    \Tile_X2Y7_NN4BEG[12] ,
    \Tile_X2Y7_NN4BEG[11] ,
    \Tile_X2Y7_NN4BEG[10] ,
    \Tile_X2Y7_NN4BEG[9] ,
    \Tile_X2Y7_NN4BEG[8] ,
    \Tile_X2Y7_NN4BEG[7] ,
    \Tile_X2Y7_NN4BEG[6] ,
    \Tile_X2Y7_NN4BEG[5] ,
    \Tile_X2Y7_NN4BEG[4] ,
    \Tile_X2Y7_NN4BEG[3] ,
    \Tile_X2Y7_NN4BEG[2] ,
    \Tile_X2Y7_NN4BEG[1] ,
    \Tile_X2Y7_NN4BEG[0] }),
    .S1BEG({\Tile_X2Y6_S1BEG[3] ,
    \Tile_X2Y6_S1BEG[2] ,
    \Tile_X2Y6_S1BEG[1] ,
    \Tile_X2Y6_S1BEG[0] }),
    .S1END({\Tile_X2Y5_S1BEG[3] ,
    \Tile_X2Y5_S1BEG[2] ,
    \Tile_X2Y5_S1BEG[1] ,
    \Tile_X2Y5_S1BEG[0] }),
    .S2BEG({\Tile_X2Y6_S2BEG[7] ,
    \Tile_X2Y6_S2BEG[6] ,
    \Tile_X2Y6_S2BEG[5] ,
    \Tile_X2Y6_S2BEG[4] ,
    \Tile_X2Y6_S2BEG[3] ,
    \Tile_X2Y6_S2BEG[2] ,
    \Tile_X2Y6_S2BEG[1] ,
    \Tile_X2Y6_S2BEG[0] }),
    .S2BEGb({\Tile_X2Y6_S2BEGb[7] ,
    \Tile_X2Y6_S2BEGb[6] ,
    \Tile_X2Y6_S2BEGb[5] ,
    \Tile_X2Y6_S2BEGb[4] ,
    \Tile_X2Y6_S2BEGb[3] ,
    \Tile_X2Y6_S2BEGb[2] ,
    \Tile_X2Y6_S2BEGb[1] ,
    \Tile_X2Y6_S2BEGb[0] }),
    .S2END({\Tile_X2Y5_S2BEGb[7] ,
    \Tile_X2Y5_S2BEGb[6] ,
    \Tile_X2Y5_S2BEGb[5] ,
    \Tile_X2Y5_S2BEGb[4] ,
    \Tile_X2Y5_S2BEGb[3] ,
    \Tile_X2Y5_S2BEGb[2] ,
    \Tile_X2Y5_S2BEGb[1] ,
    \Tile_X2Y5_S2BEGb[0] }),
    .S2MID({\Tile_X2Y5_S2BEG[7] ,
    \Tile_X2Y5_S2BEG[6] ,
    \Tile_X2Y5_S2BEG[5] ,
    \Tile_X2Y5_S2BEG[4] ,
    \Tile_X2Y5_S2BEG[3] ,
    \Tile_X2Y5_S2BEG[2] ,
    \Tile_X2Y5_S2BEG[1] ,
    \Tile_X2Y5_S2BEG[0] }),
    .S4BEG({\Tile_X2Y6_S4BEG[15] ,
    \Tile_X2Y6_S4BEG[14] ,
    \Tile_X2Y6_S4BEG[13] ,
    \Tile_X2Y6_S4BEG[12] ,
    \Tile_X2Y6_S4BEG[11] ,
    \Tile_X2Y6_S4BEG[10] ,
    \Tile_X2Y6_S4BEG[9] ,
    \Tile_X2Y6_S4BEG[8] ,
    \Tile_X2Y6_S4BEG[7] ,
    \Tile_X2Y6_S4BEG[6] ,
    \Tile_X2Y6_S4BEG[5] ,
    \Tile_X2Y6_S4BEG[4] ,
    \Tile_X2Y6_S4BEG[3] ,
    \Tile_X2Y6_S4BEG[2] ,
    \Tile_X2Y6_S4BEG[1] ,
    \Tile_X2Y6_S4BEG[0] }),
    .S4END({\Tile_X2Y5_S4BEG[15] ,
    \Tile_X2Y5_S4BEG[14] ,
    \Tile_X2Y5_S4BEG[13] ,
    \Tile_X2Y5_S4BEG[12] ,
    \Tile_X2Y5_S4BEG[11] ,
    \Tile_X2Y5_S4BEG[10] ,
    \Tile_X2Y5_S4BEG[9] ,
    \Tile_X2Y5_S4BEG[8] ,
    \Tile_X2Y5_S4BEG[7] ,
    \Tile_X2Y5_S4BEG[6] ,
    \Tile_X2Y5_S4BEG[5] ,
    \Tile_X2Y5_S4BEG[4] ,
    \Tile_X2Y5_S4BEG[3] ,
    \Tile_X2Y5_S4BEG[2] ,
    \Tile_X2Y5_S4BEG[1] ,
    \Tile_X2Y5_S4BEG[0] }),
    .SS4BEG({\Tile_X2Y6_SS4BEG[15] ,
    \Tile_X2Y6_SS4BEG[14] ,
    \Tile_X2Y6_SS4BEG[13] ,
    \Tile_X2Y6_SS4BEG[12] ,
    \Tile_X2Y6_SS4BEG[11] ,
    \Tile_X2Y6_SS4BEG[10] ,
    \Tile_X2Y6_SS4BEG[9] ,
    \Tile_X2Y6_SS4BEG[8] ,
    \Tile_X2Y6_SS4BEG[7] ,
    \Tile_X2Y6_SS4BEG[6] ,
    \Tile_X2Y6_SS4BEG[5] ,
    \Tile_X2Y6_SS4BEG[4] ,
    \Tile_X2Y6_SS4BEG[3] ,
    \Tile_X2Y6_SS4BEG[2] ,
    \Tile_X2Y6_SS4BEG[1] ,
    \Tile_X2Y6_SS4BEG[0] }),
    .SS4END({\Tile_X2Y5_SS4BEG[15] ,
    \Tile_X2Y5_SS4BEG[14] ,
    \Tile_X2Y5_SS4BEG[13] ,
    \Tile_X2Y5_SS4BEG[12] ,
    \Tile_X2Y5_SS4BEG[11] ,
    \Tile_X2Y5_SS4BEG[10] ,
    \Tile_X2Y5_SS4BEG[9] ,
    \Tile_X2Y5_SS4BEG[8] ,
    \Tile_X2Y5_SS4BEG[7] ,
    \Tile_X2Y5_SS4BEG[6] ,
    \Tile_X2Y5_SS4BEG[5] ,
    \Tile_X2Y5_SS4BEG[4] ,
    \Tile_X2Y5_SS4BEG[3] ,
    \Tile_X2Y5_SS4BEG[2] ,
    \Tile_X2Y5_SS4BEG[1] ,
    \Tile_X2Y5_SS4BEG[0] }),
    .W1BEG({\Tile_X2Y6_W1BEG[3] ,
    \Tile_X2Y6_W1BEG[2] ,
    \Tile_X2Y6_W1BEG[1] ,
    \Tile_X2Y6_W1BEG[0] }),
    .W1END({\Tile_X3Y6_W1BEG[3] ,
    \Tile_X3Y6_W1BEG[2] ,
    \Tile_X3Y6_W1BEG[1] ,
    \Tile_X3Y6_W1BEG[0] }),
    .W2BEG({\Tile_X2Y6_W2BEG[7] ,
    \Tile_X2Y6_W2BEG[6] ,
    \Tile_X2Y6_W2BEG[5] ,
    \Tile_X2Y6_W2BEG[4] ,
    \Tile_X2Y6_W2BEG[3] ,
    \Tile_X2Y6_W2BEG[2] ,
    \Tile_X2Y6_W2BEG[1] ,
    \Tile_X2Y6_W2BEG[0] }),
    .W2BEGb({\Tile_X2Y6_W2BEGb[7] ,
    \Tile_X2Y6_W2BEGb[6] ,
    \Tile_X2Y6_W2BEGb[5] ,
    \Tile_X2Y6_W2BEGb[4] ,
    \Tile_X2Y6_W2BEGb[3] ,
    \Tile_X2Y6_W2BEGb[2] ,
    \Tile_X2Y6_W2BEGb[1] ,
    \Tile_X2Y6_W2BEGb[0] }),
    .W2END({\Tile_X3Y6_W2BEGb[7] ,
    \Tile_X3Y6_W2BEGb[6] ,
    \Tile_X3Y6_W2BEGb[5] ,
    \Tile_X3Y6_W2BEGb[4] ,
    \Tile_X3Y6_W2BEGb[3] ,
    \Tile_X3Y6_W2BEGb[2] ,
    \Tile_X3Y6_W2BEGb[1] ,
    \Tile_X3Y6_W2BEGb[0] }),
    .W2MID({\Tile_X3Y6_W2BEG[7] ,
    \Tile_X3Y6_W2BEG[6] ,
    \Tile_X3Y6_W2BEG[5] ,
    \Tile_X3Y6_W2BEG[4] ,
    \Tile_X3Y6_W2BEG[3] ,
    \Tile_X3Y6_W2BEG[2] ,
    \Tile_X3Y6_W2BEG[1] ,
    \Tile_X3Y6_W2BEG[0] }),
    .W6BEG({\Tile_X2Y6_W6BEG[11] ,
    \Tile_X2Y6_W6BEG[10] ,
    \Tile_X2Y6_W6BEG[9] ,
    \Tile_X2Y6_W6BEG[8] ,
    \Tile_X2Y6_W6BEG[7] ,
    \Tile_X2Y6_W6BEG[6] ,
    \Tile_X2Y6_W6BEG[5] ,
    \Tile_X2Y6_W6BEG[4] ,
    \Tile_X2Y6_W6BEG[3] ,
    \Tile_X2Y6_W6BEG[2] ,
    \Tile_X2Y6_W6BEG[1] ,
    \Tile_X2Y6_W6BEG[0] }),
    .W6END({\Tile_X3Y6_W6BEG[11] ,
    \Tile_X3Y6_W6BEG[10] ,
    \Tile_X3Y6_W6BEG[9] ,
    \Tile_X3Y6_W6BEG[8] ,
    \Tile_X3Y6_W6BEG[7] ,
    \Tile_X3Y6_W6BEG[6] ,
    \Tile_X3Y6_W6BEG[5] ,
    \Tile_X3Y6_W6BEG[4] ,
    \Tile_X3Y6_W6BEG[3] ,
    \Tile_X3Y6_W6BEG[2] ,
    \Tile_X3Y6_W6BEG[1] ,
    \Tile_X3Y6_W6BEG[0] }),
    .WW4BEG({\Tile_X2Y6_WW4BEG[15] ,
    \Tile_X2Y6_WW4BEG[14] ,
    \Tile_X2Y6_WW4BEG[13] ,
    \Tile_X2Y6_WW4BEG[12] ,
    \Tile_X2Y6_WW4BEG[11] ,
    \Tile_X2Y6_WW4BEG[10] ,
    \Tile_X2Y6_WW4BEG[9] ,
    \Tile_X2Y6_WW4BEG[8] ,
    \Tile_X2Y6_WW4BEG[7] ,
    \Tile_X2Y6_WW4BEG[6] ,
    \Tile_X2Y6_WW4BEG[5] ,
    \Tile_X2Y6_WW4BEG[4] ,
    \Tile_X2Y6_WW4BEG[3] ,
    \Tile_X2Y6_WW4BEG[2] ,
    \Tile_X2Y6_WW4BEG[1] ,
    \Tile_X2Y6_WW4BEG[0] }),
    .WW4END({\Tile_X3Y6_WW4BEG[15] ,
    \Tile_X3Y6_WW4BEG[14] ,
    \Tile_X3Y6_WW4BEG[13] ,
    \Tile_X3Y6_WW4BEG[12] ,
    \Tile_X3Y6_WW4BEG[11] ,
    \Tile_X3Y6_WW4BEG[10] ,
    \Tile_X3Y6_WW4BEG[9] ,
    \Tile_X3Y6_WW4BEG[8] ,
    \Tile_X3Y6_WW4BEG[7] ,
    \Tile_X3Y6_WW4BEG[6] ,
    \Tile_X3Y6_WW4BEG[5] ,
    \Tile_X3Y6_WW4BEG[4] ,
    \Tile_X3Y6_WW4BEG[3] ,
    \Tile_X3Y6_WW4BEG[2] ,
    \Tile_X3Y6_WW4BEG[1] ,
    \Tile_X3Y6_WW4BEG[0] }));
 LUT4AB Tile_X2Y7_LUT4AB (.Ci(Tile_X2Y8_Co),
    .Co(Tile_X2Y7_Co),
    .UserCLK(Tile_X2Y8_UserCLKo),
    .UserCLKo(Tile_X2Y7_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X2Y7_E1BEG[3] ,
    \Tile_X2Y7_E1BEG[2] ,
    \Tile_X2Y7_E1BEG[1] ,
    \Tile_X2Y7_E1BEG[0] }),
    .E1END({\Tile_X1Y7_E1BEG[3] ,
    \Tile_X1Y7_E1BEG[2] ,
    \Tile_X1Y7_E1BEG[1] ,
    \Tile_X1Y7_E1BEG[0] }),
    .E2BEG({\Tile_X2Y7_E2BEG[7] ,
    \Tile_X2Y7_E2BEG[6] ,
    \Tile_X2Y7_E2BEG[5] ,
    \Tile_X2Y7_E2BEG[4] ,
    \Tile_X2Y7_E2BEG[3] ,
    \Tile_X2Y7_E2BEG[2] ,
    \Tile_X2Y7_E2BEG[1] ,
    \Tile_X2Y7_E2BEG[0] }),
    .E2BEGb({\Tile_X2Y7_E2BEGb[7] ,
    \Tile_X2Y7_E2BEGb[6] ,
    \Tile_X2Y7_E2BEGb[5] ,
    \Tile_X2Y7_E2BEGb[4] ,
    \Tile_X2Y7_E2BEGb[3] ,
    \Tile_X2Y7_E2BEGb[2] ,
    \Tile_X2Y7_E2BEGb[1] ,
    \Tile_X2Y7_E2BEGb[0] }),
    .E2END({\Tile_X1Y7_E2BEGb[7] ,
    \Tile_X1Y7_E2BEGb[6] ,
    \Tile_X1Y7_E2BEGb[5] ,
    \Tile_X1Y7_E2BEGb[4] ,
    \Tile_X1Y7_E2BEGb[3] ,
    \Tile_X1Y7_E2BEGb[2] ,
    \Tile_X1Y7_E2BEGb[1] ,
    \Tile_X1Y7_E2BEGb[0] }),
    .E2MID({\Tile_X1Y7_E2BEG[7] ,
    \Tile_X1Y7_E2BEG[6] ,
    \Tile_X1Y7_E2BEG[5] ,
    \Tile_X1Y7_E2BEG[4] ,
    \Tile_X1Y7_E2BEG[3] ,
    \Tile_X1Y7_E2BEG[2] ,
    \Tile_X1Y7_E2BEG[1] ,
    \Tile_X1Y7_E2BEG[0] }),
    .E6BEG({\Tile_X2Y7_E6BEG[11] ,
    \Tile_X2Y7_E6BEG[10] ,
    \Tile_X2Y7_E6BEG[9] ,
    \Tile_X2Y7_E6BEG[8] ,
    \Tile_X2Y7_E6BEG[7] ,
    \Tile_X2Y7_E6BEG[6] ,
    \Tile_X2Y7_E6BEG[5] ,
    \Tile_X2Y7_E6BEG[4] ,
    \Tile_X2Y7_E6BEG[3] ,
    \Tile_X2Y7_E6BEG[2] ,
    \Tile_X2Y7_E6BEG[1] ,
    \Tile_X2Y7_E6BEG[0] }),
    .E6END({\Tile_X1Y7_E6BEG[11] ,
    \Tile_X1Y7_E6BEG[10] ,
    \Tile_X1Y7_E6BEG[9] ,
    \Tile_X1Y7_E6BEG[8] ,
    \Tile_X1Y7_E6BEG[7] ,
    \Tile_X1Y7_E6BEG[6] ,
    \Tile_X1Y7_E6BEG[5] ,
    \Tile_X1Y7_E6BEG[4] ,
    \Tile_X1Y7_E6BEG[3] ,
    \Tile_X1Y7_E6BEG[2] ,
    \Tile_X1Y7_E6BEG[1] ,
    \Tile_X1Y7_E6BEG[0] }),
    .EE4BEG({\Tile_X2Y7_EE4BEG[15] ,
    \Tile_X2Y7_EE4BEG[14] ,
    \Tile_X2Y7_EE4BEG[13] ,
    \Tile_X2Y7_EE4BEG[12] ,
    \Tile_X2Y7_EE4BEG[11] ,
    \Tile_X2Y7_EE4BEG[10] ,
    \Tile_X2Y7_EE4BEG[9] ,
    \Tile_X2Y7_EE4BEG[8] ,
    \Tile_X2Y7_EE4BEG[7] ,
    \Tile_X2Y7_EE4BEG[6] ,
    \Tile_X2Y7_EE4BEG[5] ,
    \Tile_X2Y7_EE4BEG[4] ,
    \Tile_X2Y7_EE4BEG[3] ,
    \Tile_X2Y7_EE4BEG[2] ,
    \Tile_X2Y7_EE4BEG[1] ,
    \Tile_X2Y7_EE4BEG[0] }),
    .EE4END({\Tile_X1Y7_EE4BEG[15] ,
    \Tile_X1Y7_EE4BEG[14] ,
    \Tile_X1Y7_EE4BEG[13] ,
    \Tile_X1Y7_EE4BEG[12] ,
    \Tile_X1Y7_EE4BEG[11] ,
    \Tile_X1Y7_EE4BEG[10] ,
    \Tile_X1Y7_EE4BEG[9] ,
    \Tile_X1Y7_EE4BEG[8] ,
    \Tile_X1Y7_EE4BEG[7] ,
    \Tile_X1Y7_EE4BEG[6] ,
    \Tile_X1Y7_EE4BEG[5] ,
    \Tile_X1Y7_EE4BEG[4] ,
    \Tile_X1Y7_EE4BEG[3] ,
    \Tile_X1Y7_EE4BEG[2] ,
    \Tile_X1Y7_EE4BEG[1] ,
    \Tile_X1Y7_EE4BEG[0] }),
    .FrameData({\Tile_X1Y7_FrameData_O[31] ,
    \Tile_X1Y7_FrameData_O[30] ,
    \Tile_X1Y7_FrameData_O[29] ,
    \Tile_X1Y7_FrameData_O[28] ,
    \Tile_X1Y7_FrameData_O[27] ,
    \Tile_X1Y7_FrameData_O[26] ,
    \Tile_X1Y7_FrameData_O[25] ,
    \Tile_X1Y7_FrameData_O[24] ,
    \Tile_X1Y7_FrameData_O[23] ,
    \Tile_X1Y7_FrameData_O[22] ,
    \Tile_X1Y7_FrameData_O[21] ,
    \Tile_X1Y7_FrameData_O[20] ,
    \Tile_X1Y7_FrameData_O[19] ,
    \Tile_X1Y7_FrameData_O[18] ,
    \Tile_X1Y7_FrameData_O[17] ,
    \Tile_X1Y7_FrameData_O[16] ,
    \Tile_X1Y7_FrameData_O[15] ,
    \Tile_X1Y7_FrameData_O[14] ,
    \Tile_X1Y7_FrameData_O[13] ,
    \Tile_X1Y7_FrameData_O[12] ,
    \Tile_X1Y7_FrameData_O[11] ,
    \Tile_X1Y7_FrameData_O[10] ,
    \Tile_X1Y7_FrameData_O[9] ,
    \Tile_X1Y7_FrameData_O[8] ,
    \Tile_X1Y7_FrameData_O[7] ,
    \Tile_X1Y7_FrameData_O[6] ,
    \Tile_X1Y7_FrameData_O[5] ,
    \Tile_X1Y7_FrameData_O[4] ,
    \Tile_X1Y7_FrameData_O[3] ,
    \Tile_X1Y7_FrameData_O[2] ,
    \Tile_X1Y7_FrameData_O[1] ,
    \Tile_X1Y7_FrameData_O[0] }),
    .FrameData_O({\Tile_X2Y7_FrameData_O[31] ,
    \Tile_X2Y7_FrameData_O[30] ,
    \Tile_X2Y7_FrameData_O[29] ,
    \Tile_X2Y7_FrameData_O[28] ,
    \Tile_X2Y7_FrameData_O[27] ,
    \Tile_X2Y7_FrameData_O[26] ,
    \Tile_X2Y7_FrameData_O[25] ,
    \Tile_X2Y7_FrameData_O[24] ,
    \Tile_X2Y7_FrameData_O[23] ,
    \Tile_X2Y7_FrameData_O[22] ,
    \Tile_X2Y7_FrameData_O[21] ,
    \Tile_X2Y7_FrameData_O[20] ,
    \Tile_X2Y7_FrameData_O[19] ,
    \Tile_X2Y7_FrameData_O[18] ,
    \Tile_X2Y7_FrameData_O[17] ,
    \Tile_X2Y7_FrameData_O[16] ,
    \Tile_X2Y7_FrameData_O[15] ,
    \Tile_X2Y7_FrameData_O[14] ,
    \Tile_X2Y7_FrameData_O[13] ,
    \Tile_X2Y7_FrameData_O[12] ,
    \Tile_X2Y7_FrameData_O[11] ,
    \Tile_X2Y7_FrameData_O[10] ,
    \Tile_X2Y7_FrameData_O[9] ,
    \Tile_X2Y7_FrameData_O[8] ,
    \Tile_X2Y7_FrameData_O[7] ,
    \Tile_X2Y7_FrameData_O[6] ,
    \Tile_X2Y7_FrameData_O[5] ,
    \Tile_X2Y7_FrameData_O[4] ,
    \Tile_X2Y7_FrameData_O[3] ,
    \Tile_X2Y7_FrameData_O[2] ,
    \Tile_X2Y7_FrameData_O[1] ,
    \Tile_X2Y7_FrameData_O[0] }),
    .FrameStrobe({\Tile_X2Y8_FrameStrobe_O[19] ,
    \Tile_X2Y8_FrameStrobe_O[18] ,
    \Tile_X2Y8_FrameStrobe_O[17] ,
    \Tile_X2Y8_FrameStrobe_O[16] ,
    \Tile_X2Y8_FrameStrobe_O[15] ,
    \Tile_X2Y8_FrameStrobe_O[14] ,
    \Tile_X2Y8_FrameStrobe_O[13] ,
    \Tile_X2Y8_FrameStrobe_O[12] ,
    \Tile_X2Y8_FrameStrobe_O[11] ,
    \Tile_X2Y8_FrameStrobe_O[10] ,
    \Tile_X2Y8_FrameStrobe_O[9] ,
    \Tile_X2Y8_FrameStrobe_O[8] ,
    \Tile_X2Y8_FrameStrobe_O[7] ,
    \Tile_X2Y8_FrameStrobe_O[6] ,
    \Tile_X2Y8_FrameStrobe_O[5] ,
    \Tile_X2Y8_FrameStrobe_O[4] ,
    \Tile_X2Y8_FrameStrobe_O[3] ,
    \Tile_X2Y8_FrameStrobe_O[2] ,
    \Tile_X2Y8_FrameStrobe_O[1] ,
    \Tile_X2Y8_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X2Y7_FrameStrobe_O[19] ,
    \Tile_X2Y7_FrameStrobe_O[18] ,
    \Tile_X2Y7_FrameStrobe_O[17] ,
    \Tile_X2Y7_FrameStrobe_O[16] ,
    \Tile_X2Y7_FrameStrobe_O[15] ,
    \Tile_X2Y7_FrameStrobe_O[14] ,
    \Tile_X2Y7_FrameStrobe_O[13] ,
    \Tile_X2Y7_FrameStrobe_O[12] ,
    \Tile_X2Y7_FrameStrobe_O[11] ,
    \Tile_X2Y7_FrameStrobe_O[10] ,
    \Tile_X2Y7_FrameStrobe_O[9] ,
    \Tile_X2Y7_FrameStrobe_O[8] ,
    \Tile_X2Y7_FrameStrobe_O[7] ,
    \Tile_X2Y7_FrameStrobe_O[6] ,
    \Tile_X2Y7_FrameStrobe_O[5] ,
    \Tile_X2Y7_FrameStrobe_O[4] ,
    \Tile_X2Y7_FrameStrobe_O[3] ,
    \Tile_X2Y7_FrameStrobe_O[2] ,
    \Tile_X2Y7_FrameStrobe_O[1] ,
    \Tile_X2Y7_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X2Y7_N1BEG[3] ,
    \Tile_X2Y7_N1BEG[2] ,
    \Tile_X2Y7_N1BEG[1] ,
    \Tile_X2Y7_N1BEG[0] }),
    .N1END({\Tile_X2Y8_N1BEG[3] ,
    \Tile_X2Y8_N1BEG[2] ,
    \Tile_X2Y8_N1BEG[1] ,
    \Tile_X2Y8_N1BEG[0] }),
    .N2BEG({\Tile_X2Y7_N2BEG[7] ,
    \Tile_X2Y7_N2BEG[6] ,
    \Tile_X2Y7_N2BEG[5] ,
    \Tile_X2Y7_N2BEG[4] ,
    \Tile_X2Y7_N2BEG[3] ,
    \Tile_X2Y7_N2BEG[2] ,
    \Tile_X2Y7_N2BEG[1] ,
    \Tile_X2Y7_N2BEG[0] }),
    .N2BEGb({\Tile_X2Y7_N2BEGb[7] ,
    \Tile_X2Y7_N2BEGb[6] ,
    \Tile_X2Y7_N2BEGb[5] ,
    \Tile_X2Y7_N2BEGb[4] ,
    \Tile_X2Y7_N2BEGb[3] ,
    \Tile_X2Y7_N2BEGb[2] ,
    \Tile_X2Y7_N2BEGb[1] ,
    \Tile_X2Y7_N2BEGb[0] }),
    .N2END({\Tile_X2Y8_N2BEGb[7] ,
    \Tile_X2Y8_N2BEGb[6] ,
    \Tile_X2Y8_N2BEGb[5] ,
    \Tile_X2Y8_N2BEGb[4] ,
    \Tile_X2Y8_N2BEGb[3] ,
    \Tile_X2Y8_N2BEGb[2] ,
    \Tile_X2Y8_N2BEGb[1] ,
    \Tile_X2Y8_N2BEGb[0] }),
    .N2MID({\Tile_X2Y8_N2BEG[7] ,
    \Tile_X2Y8_N2BEG[6] ,
    \Tile_X2Y8_N2BEG[5] ,
    \Tile_X2Y8_N2BEG[4] ,
    \Tile_X2Y8_N2BEG[3] ,
    \Tile_X2Y8_N2BEG[2] ,
    \Tile_X2Y8_N2BEG[1] ,
    \Tile_X2Y8_N2BEG[0] }),
    .N4BEG({\Tile_X2Y7_N4BEG[15] ,
    \Tile_X2Y7_N4BEG[14] ,
    \Tile_X2Y7_N4BEG[13] ,
    \Tile_X2Y7_N4BEG[12] ,
    \Tile_X2Y7_N4BEG[11] ,
    \Tile_X2Y7_N4BEG[10] ,
    \Tile_X2Y7_N4BEG[9] ,
    \Tile_X2Y7_N4BEG[8] ,
    \Tile_X2Y7_N4BEG[7] ,
    \Tile_X2Y7_N4BEG[6] ,
    \Tile_X2Y7_N4BEG[5] ,
    \Tile_X2Y7_N4BEG[4] ,
    \Tile_X2Y7_N4BEG[3] ,
    \Tile_X2Y7_N4BEG[2] ,
    \Tile_X2Y7_N4BEG[1] ,
    \Tile_X2Y7_N4BEG[0] }),
    .N4END({\Tile_X2Y8_N4BEG[15] ,
    \Tile_X2Y8_N4BEG[14] ,
    \Tile_X2Y8_N4BEG[13] ,
    \Tile_X2Y8_N4BEG[12] ,
    \Tile_X2Y8_N4BEG[11] ,
    \Tile_X2Y8_N4BEG[10] ,
    \Tile_X2Y8_N4BEG[9] ,
    \Tile_X2Y8_N4BEG[8] ,
    \Tile_X2Y8_N4BEG[7] ,
    \Tile_X2Y8_N4BEG[6] ,
    \Tile_X2Y8_N4BEG[5] ,
    \Tile_X2Y8_N4BEG[4] ,
    \Tile_X2Y8_N4BEG[3] ,
    \Tile_X2Y8_N4BEG[2] ,
    \Tile_X2Y8_N4BEG[1] ,
    \Tile_X2Y8_N4BEG[0] }),
    .NN4BEG({\Tile_X2Y7_NN4BEG[15] ,
    \Tile_X2Y7_NN4BEG[14] ,
    \Tile_X2Y7_NN4BEG[13] ,
    \Tile_X2Y7_NN4BEG[12] ,
    \Tile_X2Y7_NN4BEG[11] ,
    \Tile_X2Y7_NN4BEG[10] ,
    \Tile_X2Y7_NN4BEG[9] ,
    \Tile_X2Y7_NN4BEG[8] ,
    \Tile_X2Y7_NN4BEG[7] ,
    \Tile_X2Y7_NN4BEG[6] ,
    \Tile_X2Y7_NN4BEG[5] ,
    \Tile_X2Y7_NN4BEG[4] ,
    \Tile_X2Y7_NN4BEG[3] ,
    \Tile_X2Y7_NN4BEG[2] ,
    \Tile_X2Y7_NN4BEG[1] ,
    \Tile_X2Y7_NN4BEG[0] }),
    .NN4END({\Tile_X2Y8_NN4BEG[15] ,
    \Tile_X2Y8_NN4BEG[14] ,
    \Tile_X2Y8_NN4BEG[13] ,
    \Tile_X2Y8_NN4BEG[12] ,
    \Tile_X2Y8_NN4BEG[11] ,
    \Tile_X2Y8_NN4BEG[10] ,
    \Tile_X2Y8_NN4BEG[9] ,
    \Tile_X2Y8_NN4BEG[8] ,
    \Tile_X2Y8_NN4BEG[7] ,
    \Tile_X2Y8_NN4BEG[6] ,
    \Tile_X2Y8_NN4BEG[5] ,
    \Tile_X2Y8_NN4BEG[4] ,
    \Tile_X2Y8_NN4BEG[3] ,
    \Tile_X2Y8_NN4BEG[2] ,
    \Tile_X2Y8_NN4BEG[1] ,
    \Tile_X2Y8_NN4BEG[0] }),
    .S1BEG({\Tile_X2Y7_S1BEG[3] ,
    \Tile_X2Y7_S1BEG[2] ,
    \Tile_X2Y7_S1BEG[1] ,
    \Tile_X2Y7_S1BEG[0] }),
    .S1END({\Tile_X2Y6_S1BEG[3] ,
    \Tile_X2Y6_S1BEG[2] ,
    \Tile_X2Y6_S1BEG[1] ,
    \Tile_X2Y6_S1BEG[0] }),
    .S2BEG({\Tile_X2Y7_S2BEG[7] ,
    \Tile_X2Y7_S2BEG[6] ,
    \Tile_X2Y7_S2BEG[5] ,
    \Tile_X2Y7_S2BEG[4] ,
    \Tile_X2Y7_S2BEG[3] ,
    \Tile_X2Y7_S2BEG[2] ,
    \Tile_X2Y7_S2BEG[1] ,
    \Tile_X2Y7_S2BEG[0] }),
    .S2BEGb({\Tile_X2Y7_S2BEGb[7] ,
    \Tile_X2Y7_S2BEGb[6] ,
    \Tile_X2Y7_S2BEGb[5] ,
    \Tile_X2Y7_S2BEGb[4] ,
    \Tile_X2Y7_S2BEGb[3] ,
    \Tile_X2Y7_S2BEGb[2] ,
    \Tile_X2Y7_S2BEGb[1] ,
    \Tile_X2Y7_S2BEGb[0] }),
    .S2END({\Tile_X2Y6_S2BEGb[7] ,
    \Tile_X2Y6_S2BEGb[6] ,
    \Tile_X2Y6_S2BEGb[5] ,
    \Tile_X2Y6_S2BEGb[4] ,
    \Tile_X2Y6_S2BEGb[3] ,
    \Tile_X2Y6_S2BEGb[2] ,
    \Tile_X2Y6_S2BEGb[1] ,
    \Tile_X2Y6_S2BEGb[0] }),
    .S2MID({\Tile_X2Y6_S2BEG[7] ,
    \Tile_X2Y6_S2BEG[6] ,
    \Tile_X2Y6_S2BEG[5] ,
    \Tile_X2Y6_S2BEG[4] ,
    \Tile_X2Y6_S2BEG[3] ,
    \Tile_X2Y6_S2BEG[2] ,
    \Tile_X2Y6_S2BEG[1] ,
    \Tile_X2Y6_S2BEG[0] }),
    .S4BEG({\Tile_X2Y7_S4BEG[15] ,
    \Tile_X2Y7_S4BEG[14] ,
    \Tile_X2Y7_S4BEG[13] ,
    \Tile_X2Y7_S4BEG[12] ,
    \Tile_X2Y7_S4BEG[11] ,
    \Tile_X2Y7_S4BEG[10] ,
    \Tile_X2Y7_S4BEG[9] ,
    \Tile_X2Y7_S4BEG[8] ,
    \Tile_X2Y7_S4BEG[7] ,
    \Tile_X2Y7_S4BEG[6] ,
    \Tile_X2Y7_S4BEG[5] ,
    \Tile_X2Y7_S4BEG[4] ,
    \Tile_X2Y7_S4BEG[3] ,
    \Tile_X2Y7_S4BEG[2] ,
    \Tile_X2Y7_S4BEG[1] ,
    \Tile_X2Y7_S4BEG[0] }),
    .S4END({\Tile_X2Y6_S4BEG[15] ,
    \Tile_X2Y6_S4BEG[14] ,
    \Tile_X2Y6_S4BEG[13] ,
    \Tile_X2Y6_S4BEG[12] ,
    \Tile_X2Y6_S4BEG[11] ,
    \Tile_X2Y6_S4BEG[10] ,
    \Tile_X2Y6_S4BEG[9] ,
    \Tile_X2Y6_S4BEG[8] ,
    \Tile_X2Y6_S4BEG[7] ,
    \Tile_X2Y6_S4BEG[6] ,
    \Tile_X2Y6_S4BEG[5] ,
    \Tile_X2Y6_S4BEG[4] ,
    \Tile_X2Y6_S4BEG[3] ,
    \Tile_X2Y6_S4BEG[2] ,
    \Tile_X2Y6_S4BEG[1] ,
    \Tile_X2Y6_S4BEG[0] }),
    .SS4BEG({\Tile_X2Y7_SS4BEG[15] ,
    \Tile_X2Y7_SS4BEG[14] ,
    \Tile_X2Y7_SS4BEG[13] ,
    \Tile_X2Y7_SS4BEG[12] ,
    \Tile_X2Y7_SS4BEG[11] ,
    \Tile_X2Y7_SS4BEG[10] ,
    \Tile_X2Y7_SS4BEG[9] ,
    \Tile_X2Y7_SS4BEG[8] ,
    \Tile_X2Y7_SS4BEG[7] ,
    \Tile_X2Y7_SS4BEG[6] ,
    \Tile_X2Y7_SS4BEG[5] ,
    \Tile_X2Y7_SS4BEG[4] ,
    \Tile_X2Y7_SS4BEG[3] ,
    \Tile_X2Y7_SS4BEG[2] ,
    \Tile_X2Y7_SS4BEG[1] ,
    \Tile_X2Y7_SS4BEG[0] }),
    .SS4END({\Tile_X2Y6_SS4BEG[15] ,
    \Tile_X2Y6_SS4BEG[14] ,
    \Tile_X2Y6_SS4BEG[13] ,
    \Tile_X2Y6_SS4BEG[12] ,
    \Tile_X2Y6_SS4BEG[11] ,
    \Tile_X2Y6_SS4BEG[10] ,
    \Tile_X2Y6_SS4BEG[9] ,
    \Tile_X2Y6_SS4BEG[8] ,
    \Tile_X2Y6_SS4BEG[7] ,
    \Tile_X2Y6_SS4BEG[6] ,
    \Tile_X2Y6_SS4BEG[5] ,
    \Tile_X2Y6_SS4BEG[4] ,
    \Tile_X2Y6_SS4BEG[3] ,
    \Tile_X2Y6_SS4BEG[2] ,
    \Tile_X2Y6_SS4BEG[1] ,
    \Tile_X2Y6_SS4BEG[0] }),
    .W1BEG({\Tile_X2Y7_W1BEG[3] ,
    \Tile_X2Y7_W1BEG[2] ,
    \Tile_X2Y7_W1BEG[1] ,
    \Tile_X2Y7_W1BEG[0] }),
    .W1END({\Tile_X3Y7_W1BEG[3] ,
    \Tile_X3Y7_W1BEG[2] ,
    \Tile_X3Y7_W1BEG[1] ,
    \Tile_X3Y7_W1BEG[0] }),
    .W2BEG({\Tile_X2Y7_W2BEG[7] ,
    \Tile_X2Y7_W2BEG[6] ,
    \Tile_X2Y7_W2BEG[5] ,
    \Tile_X2Y7_W2BEG[4] ,
    \Tile_X2Y7_W2BEG[3] ,
    \Tile_X2Y7_W2BEG[2] ,
    \Tile_X2Y7_W2BEG[1] ,
    \Tile_X2Y7_W2BEG[0] }),
    .W2BEGb({\Tile_X2Y7_W2BEGb[7] ,
    \Tile_X2Y7_W2BEGb[6] ,
    \Tile_X2Y7_W2BEGb[5] ,
    \Tile_X2Y7_W2BEGb[4] ,
    \Tile_X2Y7_W2BEGb[3] ,
    \Tile_X2Y7_W2BEGb[2] ,
    \Tile_X2Y7_W2BEGb[1] ,
    \Tile_X2Y7_W2BEGb[0] }),
    .W2END({\Tile_X3Y7_W2BEGb[7] ,
    \Tile_X3Y7_W2BEGb[6] ,
    \Tile_X3Y7_W2BEGb[5] ,
    \Tile_X3Y7_W2BEGb[4] ,
    \Tile_X3Y7_W2BEGb[3] ,
    \Tile_X3Y7_W2BEGb[2] ,
    \Tile_X3Y7_W2BEGb[1] ,
    \Tile_X3Y7_W2BEGb[0] }),
    .W2MID({\Tile_X3Y7_W2BEG[7] ,
    \Tile_X3Y7_W2BEG[6] ,
    \Tile_X3Y7_W2BEG[5] ,
    \Tile_X3Y7_W2BEG[4] ,
    \Tile_X3Y7_W2BEG[3] ,
    \Tile_X3Y7_W2BEG[2] ,
    \Tile_X3Y7_W2BEG[1] ,
    \Tile_X3Y7_W2BEG[0] }),
    .W6BEG({\Tile_X2Y7_W6BEG[11] ,
    \Tile_X2Y7_W6BEG[10] ,
    \Tile_X2Y7_W6BEG[9] ,
    \Tile_X2Y7_W6BEG[8] ,
    \Tile_X2Y7_W6BEG[7] ,
    \Tile_X2Y7_W6BEG[6] ,
    \Tile_X2Y7_W6BEG[5] ,
    \Tile_X2Y7_W6BEG[4] ,
    \Tile_X2Y7_W6BEG[3] ,
    \Tile_X2Y7_W6BEG[2] ,
    \Tile_X2Y7_W6BEG[1] ,
    \Tile_X2Y7_W6BEG[0] }),
    .W6END({\Tile_X3Y7_W6BEG[11] ,
    \Tile_X3Y7_W6BEG[10] ,
    \Tile_X3Y7_W6BEG[9] ,
    \Tile_X3Y7_W6BEG[8] ,
    \Tile_X3Y7_W6BEG[7] ,
    \Tile_X3Y7_W6BEG[6] ,
    \Tile_X3Y7_W6BEG[5] ,
    \Tile_X3Y7_W6BEG[4] ,
    \Tile_X3Y7_W6BEG[3] ,
    \Tile_X3Y7_W6BEG[2] ,
    \Tile_X3Y7_W6BEG[1] ,
    \Tile_X3Y7_W6BEG[0] }),
    .WW4BEG({\Tile_X2Y7_WW4BEG[15] ,
    \Tile_X2Y7_WW4BEG[14] ,
    \Tile_X2Y7_WW4BEG[13] ,
    \Tile_X2Y7_WW4BEG[12] ,
    \Tile_X2Y7_WW4BEG[11] ,
    \Tile_X2Y7_WW4BEG[10] ,
    \Tile_X2Y7_WW4BEG[9] ,
    \Tile_X2Y7_WW4BEG[8] ,
    \Tile_X2Y7_WW4BEG[7] ,
    \Tile_X2Y7_WW4BEG[6] ,
    \Tile_X2Y7_WW4BEG[5] ,
    \Tile_X2Y7_WW4BEG[4] ,
    \Tile_X2Y7_WW4BEG[3] ,
    \Tile_X2Y7_WW4BEG[2] ,
    \Tile_X2Y7_WW4BEG[1] ,
    \Tile_X2Y7_WW4BEG[0] }),
    .WW4END({\Tile_X3Y7_WW4BEG[15] ,
    \Tile_X3Y7_WW4BEG[14] ,
    \Tile_X3Y7_WW4BEG[13] ,
    \Tile_X3Y7_WW4BEG[12] ,
    \Tile_X3Y7_WW4BEG[11] ,
    \Tile_X3Y7_WW4BEG[10] ,
    \Tile_X3Y7_WW4BEG[9] ,
    \Tile_X3Y7_WW4BEG[8] ,
    \Tile_X3Y7_WW4BEG[7] ,
    \Tile_X3Y7_WW4BEG[6] ,
    \Tile_X3Y7_WW4BEG[5] ,
    \Tile_X3Y7_WW4BEG[4] ,
    \Tile_X3Y7_WW4BEG[3] ,
    \Tile_X3Y7_WW4BEG[2] ,
    \Tile_X3Y7_WW4BEG[1] ,
    \Tile_X3Y7_WW4BEG[0] }));
 LUT4AB Tile_X2Y8_LUT4AB (.Ci(Tile_X2Y9_Co),
    .Co(Tile_X2Y8_Co),
    .UserCLK(Tile_X2Y9_UserCLKo),
    .UserCLKo(Tile_X2Y8_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X2Y8_E1BEG[3] ,
    \Tile_X2Y8_E1BEG[2] ,
    \Tile_X2Y8_E1BEG[1] ,
    \Tile_X2Y8_E1BEG[0] }),
    .E1END({\Tile_X1Y8_E1BEG[3] ,
    \Tile_X1Y8_E1BEG[2] ,
    \Tile_X1Y8_E1BEG[1] ,
    \Tile_X1Y8_E1BEG[0] }),
    .E2BEG({\Tile_X2Y8_E2BEG[7] ,
    \Tile_X2Y8_E2BEG[6] ,
    \Tile_X2Y8_E2BEG[5] ,
    \Tile_X2Y8_E2BEG[4] ,
    \Tile_X2Y8_E2BEG[3] ,
    \Tile_X2Y8_E2BEG[2] ,
    \Tile_X2Y8_E2BEG[1] ,
    \Tile_X2Y8_E2BEG[0] }),
    .E2BEGb({\Tile_X2Y8_E2BEGb[7] ,
    \Tile_X2Y8_E2BEGb[6] ,
    \Tile_X2Y8_E2BEGb[5] ,
    \Tile_X2Y8_E2BEGb[4] ,
    \Tile_X2Y8_E2BEGb[3] ,
    \Tile_X2Y8_E2BEGb[2] ,
    \Tile_X2Y8_E2BEGb[1] ,
    \Tile_X2Y8_E2BEGb[0] }),
    .E2END({\Tile_X1Y8_E2BEGb[7] ,
    \Tile_X1Y8_E2BEGb[6] ,
    \Tile_X1Y8_E2BEGb[5] ,
    \Tile_X1Y8_E2BEGb[4] ,
    \Tile_X1Y8_E2BEGb[3] ,
    \Tile_X1Y8_E2BEGb[2] ,
    \Tile_X1Y8_E2BEGb[1] ,
    \Tile_X1Y8_E2BEGb[0] }),
    .E2MID({\Tile_X1Y8_E2BEG[7] ,
    \Tile_X1Y8_E2BEG[6] ,
    \Tile_X1Y8_E2BEG[5] ,
    \Tile_X1Y8_E2BEG[4] ,
    \Tile_X1Y8_E2BEG[3] ,
    \Tile_X1Y8_E2BEG[2] ,
    \Tile_X1Y8_E2BEG[1] ,
    \Tile_X1Y8_E2BEG[0] }),
    .E6BEG({\Tile_X2Y8_E6BEG[11] ,
    \Tile_X2Y8_E6BEG[10] ,
    \Tile_X2Y8_E6BEG[9] ,
    \Tile_X2Y8_E6BEG[8] ,
    \Tile_X2Y8_E6BEG[7] ,
    \Tile_X2Y8_E6BEG[6] ,
    \Tile_X2Y8_E6BEG[5] ,
    \Tile_X2Y8_E6BEG[4] ,
    \Tile_X2Y8_E6BEG[3] ,
    \Tile_X2Y8_E6BEG[2] ,
    \Tile_X2Y8_E6BEG[1] ,
    \Tile_X2Y8_E6BEG[0] }),
    .E6END({\Tile_X1Y8_E6BEG[11] ,
    \Tile_X1Y8_E6BEG[10] ,
    \Tile_X1Y8_E6BEG[9] ,
    \Tile_X1Y8_E6BEG[8] ,
    \Tile_X1Y8_E6BEG[7] ,
    \Tile_X1Y8_E6BEG[6] ,
    \Tile_X1Y8_E6BEG[5] ,
    \Tile_X1Y8_E6BEG[4] ,
    \Tile_X1Y8_E6BEG[3] ,
    \Tile_X1Y8_E6BEG[2] ,
    \Tile_X1Y8_E6BEG[1] ,
    \Tile_X1Y8_E6BEG[0] }),
    .EE4BEG({\Tile_X2Y8_EE4BEG[15] ,
    \Tile_X2Y8_EE4BEG[14] ,
    \Tile_X2Y8_EE4BEG[13] ,
    \Tile_X2Y8_EE4BEG[12] ,
    \Tile_X2Y8_EE4BEG[11] ,
    \Tile_X2Y8_EE4BEG[10] ,
    \Tile_X2Y8_EE4BEG[9] ,
    \Tile_X2Y8_EE4BEG[8] ,
    \Tile_X2Y8_EE4BEG[7] ,
    \Tile_X2Y8_EE4BEG[6] ,
    \Tile_X2Y8_EE4BEG[5] ,
    \Tile_X2Y8_EE4BEG[4] ,
    \Tile_X2Y8_EE4BEG[3] ,
    \Tile_X2Y8_EE4BEG[2] ,
    \Tile_X2Y8_EE4BEG[1] ,
    \Tile_X2Y8_EE4BEG[0] }),
    .EE4END({\Tile_X1Y8_EE4BEG[15] ,
    \Tile_X1Y8_EE4BEG[14] ,
    \Tile_X1Y8_EE4BEG[13] ,
    \Tile_X1Y8_EE4BEG[12] ,
    \Tile_X1Y8_EE4BEG[11] ,
    \Tile_X1Y8_EE4BEG[10] ,
    \Tile_X1Y8_EE4BEG[9] ,
    \Tile_X1Y8_EE4BEG[8] ,
    \Tile_X1Y8_EE4BEG[7] ,
    \Tile_X1Y8_EE4BEG[6] ,
    \Tile_X1Y8_EE4BEG[5] ,
    \Tile_X1Y8_EE4BEG[4] ,
    \Tile_X1Y8_EE4BEG[3] ,
    \Tile_X1Y8_EE4BEG[2] ,
    \Tile_X1Y8_EE4BEG[1] ,
    \Tile_X1Y8_EE4BEG[0] }),
    .FrameData({\Tile_X1Y8_FrameData_O[31] ,
    \Tile_X1Y8_FrameData_O[30] ,
    \Tile_X1Y8_FrameData_O[29] ,
    \Tile_X1Y8_FrameData_O[28] ,
    \Tile_X1Y8_FrameData_O[27] ,
    \Tile_X1Y8_FrameData_O[26] ,
    \Tile_X1Y8_FrameData_O[25] ,
    \Tile_X1Y8_FrameData_O[24] ,
    \Tile_X1Y8_FrameData_O[23] ,
    \Tile_X1Y8_FrameData_O[22] ,
    \Tile_X1Y8_FrameData_O[21] ,
    \Tile_X1Y8_FrameData_O[20] ,
    \Tile_X1Y8_FrameData_O[19] ,
    \Tile_X1Y8_FrameData_O[18] ,
    \Tile_X1Y8_FrameData_O[17] ,
    \Tile_X1Y8_FrameData_O[16] ,
    \Tile_X1Y8_FrameData_O[15] ,
    \Tile_X1Y8_FrameData_O[14] ,
    \Tile_X1Y8_FrameData_O[13] ,
    \Tile_X1Y8_FrameData_O[12] ,
    \Tile_X1Y8_FrameData_O[11] ,
    \Tile_X1Y8_FrameData_O[10] ,
    \Tile_X1Y8_FrameData_O[9] ,
    \Tile_X1Y8_FrameData_O[8] ,
    \Tile_X1Y8_FrameData_O[7] ,
    \Tile_X1Y8_FrameData_O[6] ,
    \Tile_X1Y8_FrameData_O[5] ,
    \Tile_X1Y8_FrameData_O[4] ,
    \Tile_X1Y8_FrameData_O[3] ,
    \Tile_X1Y8_FrameData_O[2] ,
    \Tile_X1Y8_FrameData_O[1] ,
    \Tile_X1Y8_FrameData_O[0] }),
    .FrameData_O({\Tile_X2Y8_FrameData_O[31] ,
    \Tile_X2Y8_FrameData_O[30] ,
    \Tile_X2Y8_FrameData_O[29] ,
    \Tile_X2Y8_FrameData_O[28] ,
    \Tile_X2Y8_FrameData_O[27] ,
    \Tile_X2Y8_FrameData_O[26] ,
    \Tile_X2Y8_FrameData_O[25] ,
    \Tile_X2Y8_FrameData_O[24] ,
    \Tile_X2Y8_FrameData_O[23] ,
    \Tile_X2Y8_FrameData_O[22] ,
    \Tile_X2Y8_FrameData_O[21] ,
    \Tile_X2Y8_FrameData_O[20] ,
    \Tile_X2Y8_FrameData_O[19] ,
    \Tile_X2Y8_FrameData_O[18] ,
    \Tile_X2Y8_FrameData_O[17] ,
    \Tile_X2Y8_FrameData_O[16] ,
    \Tile_X2Y8_FrameData_O[15] ,
    \Tile_X2Y8_FrameData_O[14] ,
    \Tile_X2Y8_FrameData_O[13] ,
    \Tile_X2Y8_FrameData_O[12] ,
    \Tile_X2Y8_FrameData_O[11] ,
    \Tile_X2Y8_FrameData_O[10] ,
    \Tile_X2Y8_FrameData_O[9] ,
    \Tile_X2Y8_FrameData_O[8] ,
    \Tile_X2Y8_FrameData_O[7] ,
    \Tile_X2Y8_FrameData_O[6] ,
    \Tile_X2Y8_FrameData_O[5] ,
    \Tile_X2Y8_FrameData_O[4] ,
    \Tile_X2Y8_FrameData_O[3] ,
    \Tile_X2Y8_FrameData_O[2] ,
    \Tile_X2Y8_FrameData_O[1] ,
    \Tile_X2Y8_FrameData_O[0] }),
    .FrameStrobe({\Tile_X2Y9_FrameStrobe_O[19] ,
    \Tile_X2Y9_FrameStrobe_O[18] ,
    \Tile_X2Y9_FrameStrobe_O[17] ,
    \Tile_X2Y9_FrameStrobe_O[16] ,
    \Tile_X2Y9_FrameStrobe_O[15] ,
    \Tile_X2Y9_FrameStrobe_O[14] ,
    \Tile_X2Y9_FrameStrobe_O[13] ,
    \Tile_X2Y9_FrameStrobe_O[12] ,
    \Tile_X2Y9_FrameStrobe_O[11] ,
    \Tile_X2Y9_FrameStrobe_O[10] ,
    \Tile_X2Y9_FrameStrobe_O[9] ,
    \Tile_X2Y9_FrameStrobe_O[8] ,
    \Tile_X2Y9_FrameStrobe_O[7] ,
    \Tile_X2Y9_FrameStrobe_O[6] ,
    \Tile_X2Y9_FrameStrobe_O[5] ,
    \Tile_X2Y9_FrameStrobe_O[4] ,
    \Tile_X2Y9_FrameStrobe_O[3] ,
    \Tile_X2Y9_FrameStrobe_O[2] ,
    \Tile_X2Y9_FrameStrobe_O[1] ,
    \Tile_X2Y9_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X2Y8_FrameStrobe_O[19] ,
    \Tile_X2Y8_FrameStrobe_O[18] ,
    \Tile_X2Y8_FrameStrobe_O[17] ,
    \Tile_X2Y8_FrameStrobe_O[16] ,
    \Tile_X2Y8_FrameStrobe_O[15] ,
    \Tile_X2Y8_FrameStrobe_O[14] ,
    \Tile_X2Y8_FrameStrobe_O[13] ,
    \Tile_X2Y8_FrameStrobe_O[12] ,
    \Tile_X2Y8_FrameStrobe_O[11] ,
    \Tile_X2Y8_FrameStrobe_O[10] ,
    \Tile_X2Y8_FrameStrobe_O[9] ,
    \Tile_X2Y8_FrameStrobe_O[8] ,
    \Tile_X2Y8_FrameStrobe_O[7] ,
    \Tile_X2Y8_FrameStrobe_O[6] ,
    \Tile_X2Y8_FrameStrobe_O[5] ,
    \Tile_X2Y8_FrameStrobe_O[4] ,
    \Tile_X2Y8_FrameStrobe_O[3] ,
    \Tile_X2Y8_FrameStrobe_O[2] ,
    \Tile_X2Y8_FrameStrobe_O[1] ,
    \Tile_X2Y8_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X2Y8_N1BEG[3] ,
    \Tile_X2Y8_N1BEG[2] ,
    \Tile_X2Y8_N1BEG[1] ,
    \Tile_X2Y8_N1BEG[0] }),
    .N1END({\Tile_X2Y9_N1BEG[3] ,
    \Tile_X2Y9_N1BEG[2] ,
    \Tile_X2Y9_N1BEG[1] ,
    \Tile_X2Y9_N1BEG[0] }),
    .N2BEG({\Tile_X2Y8_N2BEG[7] ,
    \Tile_X2Y8_N2BEG[6] ,
    \Tile_X2Y8_N2BEG[5] ,
    \Tile_X2Y8_N2BEG[4] ,
    \Tile_X2Y8_N2BEG[3] ,
    \Tile_X2Y8_N2BEG[2] ,
    \Tile_X2Y8_N2BEG[1] ,
    \Tile_X2Y8_N2BEG[0] }),
    .N2BEGb({\Tile_X2Y8_N2BEGb[7] ,
    \Tile_X2Y8_N2BEGb[6] ,
    \Tile_X2Y8_N2BEGb[5] ,
    \Tile_X2Y8_N2BEGb[4] ,
    \Tile_X2Y8_N2BEGb[3] ,
    \Tile_X2Y8_N2BEGb[2] ,
    \Tile_X2Y8_N2BEGb[1] ,
    \Tile_X2Y8_N2BEGb[0] }),
    .N2END({\Tile_X2Y9_N2BEGb[7] ,
    \Tile_X2Y9_N2BEGb[6] ,
    \Tile_X2Y9_N2BEGb[5] ,
    \Tile_X2Y9_N2BEGb[4] ,
    \Tile_X2Y9_N2BEGb[3] ,
    \Tile_X2Y9_N2BEGb[2] ,
    \Tile_X2Y9_N2BEGb[1] ,
    \Tile_X2Y9_N2BEGb[0] }),
    .N2MID({\Tile_X2Y9_N2BEG[7] ,
    \Tile_X2Y9_N2BEG[6] ,
    \Tile_X2Y9_N2BEG[5] ,
    \Tile_X2Y9_N2BEG[4] ,
    \Tile_X2Y9_N2BEG[3] ,
    \Tile_X2Y9_N2BEG[2] ,
    \Tile_X2Y9_N2BEG[1] ,
    \Tile_X2Y9_N2BEG[0] }),
    .N4BEG({\Tile_X2Y8_N4BEG[15] ,
    \Tile_X2Y8_N4BEG[14] ,
    \Tile_X2Y8_N4BEG[13] ,
    \Tile_X2Y8_N4BEG[12] ,
    \Tile_X2Y8_N4BEG[11] ,
    \Tile_X2Y8_N4BEG[10] ,
    \Tile_X2Y8_N4BEG[9] ,
    \Tile_X2Y8_N4BEG[8] ,
    \Tile_X2Y8_N4BEG[7] ,
    \Tile_X2Y8_N4BEG[6] ,
    \Tile_X2Y8_N4BEG[5] ,
    \Tile_X2Y8_N4BEG[4] ,
    \Tile_X2Y8_N4BEG[3] ,
    \Tile_X2Y8_N4BEG[2] ,
    \Tile_X2Y8_N4BEG[1] ,
    \Tile_X2Y8_N4BEG[0] }),
    .N4END({\Tile_X2Y9_N4BEG[15] ,
    \Tile_X2Y9_N4BEG[14] ,
    \Tile_X2Y9_N4BEG[13] ,
    \Tile_X2Y9_N4BEG[12] ,
    \Tile_X2Y9_N4BEG[11] ,
    \Tile_X2Y9_N4BEG[10] ,
    \Tile_X2Y9_N4BEG[9] ,
    \Tile_X2Y9_N4BEG[8] ,
    \Tile_X2Y9_N4BEG[7] ,
    \Tile_X2Y9_N4BEG[6] ,
    \Tile_X2Y9_N4BEG[5] ,
    \Tile_X2Y9_N4BEG[4] ,
    \Tile_X2Y9_N4BEG[3] ,
    \Tile_X2Y9_N4BEG[2] ,
    \Tile_X2Y9_N4BEG[1] ,
    \Tile_X2Y9_N4BEG[0] }),
    .NN4BEG({\Tile_X2Y8_NN4BEG[15] ,
    \Tile_X2Y8_NN4BEG[14] ,
    \Tile_X2Y8_NN4BEG[13] ,
    \Tile_X2Y8_NN4BEG[12] ,
    \Tile_X2Y8_NN4BEG[11] ,
    \Tile_X2Y8_NN4BEG[10] ,
    \Tile_X2Y8_NN4BEG[9] ,
    \Tile_X2Y8_NN4BEG[8] ,
    \Tile_X2Y8_NN4BEG[7] ,
    \Tile_X2Y8_NN4BEG[6] ,
    \Tile_X2Y8_NN4BEG[5] ,
    \Tile_X2Y8_NN4BEG[4] ,
    \Tile_X2Y8_NN4BEG[3] ,
    \Tile_X2Y8_NN4BEG[2] ,
    \Tile_X2Y8_NN4BEG[1] ,
    \Tile_X2Y8_NN4BEG[0] }),
    .NN4END({\Tile_X2Y9_NN4BEG[15] ,
    \Tile_X2Y9_NN4BEG[14] ,
    \Tile_X2Y9_NN4BEG[13] ,
    \Tile_X2Y9_NN4BEG[12] ,
    \Tile_X2Y9_NN4BEG[11] ,
    \Tile_X2Y9_NN4BEG[10] ,
    \Tile_X2Y9_NN4BEG[9] ,
    \Tile_X2Y9_NN4BEG[8] ,
    \Tile_X2Y9_NN4BEG[7] ,
    \Tile_X2Y9_NN4BEG[6] ,
    \Tile_X2Y9_NN4BEG[5] ,
    \Tile_X2Y9_NN4BEG[4] ,
    \Tile_X2Y9_NN4BEG[3] ,
    \Tile_X2Y9_NN4BEG[2] ,
    \Tile_X2Y9_NN4BEG[1] ,
    \Tile_X2Y9_NN4BEG[0] }),
    .S1BEG({\Tile_X2Y8_S1BEG[3] ,
    \Tile_X2Y8_S1BEG[2] ,
    \Tile_X2Y8_S1BEG[1] ,
    \Tile_X2Y8_S1BEG[0] }),
    .S1END({\Tile_X2Y7_S1BEG[3] ,
    \Tile_X2Y7_S1BEG[2] ,
    \Tile_X2Y7_S1BEG[1] ,
    \Tile_X2Y7_S1BEG[0] }),
    .S2BEG({\Tile_X2Y8_S2BEG[7] ,
    \Tile_X2Y8_S2BEG[6] ,
    \Tile_X2Y8_S2BEG[5] ,
    \Tile_X2Y8_S2BEG[4] ,
    \Tile_X2Y8_S2BEG[3] ,
    \Tile_X2Y8_S2BEG[2] ,
    \Tile_X2Y8_S2BEG[1] ,
    \Tile_X2Y8_S2BEG[0] }),
    .S2BEGb({\Tile_X2Y8_S2BEGb[7] ,
    \Tile_X2Y8_S2BEGb[6] ,
    \Tile_X2Y8_S2BEGb[5] ,
    \Tile_X2Y8_S2BEGb[4] ,
    \Tile_X2Y8_S2BEGb[3] ,
    \Tile_X2Y8_S2BEGb[2] ,
    \Tile_X2Y8_S2BEGb[1] ,
    \Tile_X2Y8_S2BEGb[0] }),
    .S2END({\Tile_X2Y7_S2BEGb[7] ,
    \Tile_X2Y7_S2BEGb[6] ,
    \Tile_X2Y7_S2BEGb[5] ,
    \Tile_X2Y7_S2BEGb[4] ,
    \Tile_X2Y7_S2BEGb[3] ,
    \Tile_X2Y7_S2BEGb[2] ,
    \Tile_X2Y7_S2BEGb[1] ,
    \Tile_X2Y7_S2BEGb[0] }),
    .S2MID({\Tile_X2Y7_S2BEG[7] ,
    \Tile_X2Y7_S2BEG[6] ,
    \Tile_X2Y7_S2BEG[5] ,
    \Tile_X2Y7_S2BEG[4] ,
    \Tile_X2Y7_S2BEG[3] ,
    \Tile_X2Y7_S2BEG[2] ,
    \Tile_X2Y7_S2BEG[1] ,
    \Tile_X2Y7_S2BEG[0] }),
    .S4BEG({\Tile_X2Y8_S4BEG[15] ,
    \Tile_X2Y8_S4BEG[14] ,
    \Tile_X2Y8_S4BEG[13] ,
    \Tile_X2Y8_S4BEG[12] ,
    \Tile_X2Y8_S4BEG[11] ,
    \Tile_X2Y8_S4BEG[10] ,
    \Tile_X2Y8_S4BEG[9] ,
    \Tile_X2Y8_S4BEG[8] ,
    \Tile_X2Y8_S4BEG[7] ,
    \Tile_X2Y8_S4BEG[6] ,
    \Tile_X2Y8_S4BEG[5] ,
    \Tile_X2Y8_S4BEG[4] ,
    \Tile_X2Y8_S4BEG[3] ,
    \Tile_X2Y8_S4BEG[2] ,
    \Tile_X2Y8_S4BEG[1] ,
    \Tile_X2Y8_S4BEG[0] }),
    .S4END({\Tile_X2Y7_S4BEG[15] ,
    \Tile_X2Y7_S4BEG[14] ,
    \Tile_X2Y7_S4BEG[13] ,
    \Tile_X2Y7_S4BEG[12] ,
    \Tile_X2Y7_S4BEG[11] ,
    \Tile_X2Y7_S4BEG[10] ,
    \Tile_X2Y7_S4BEG[9] ,
    \Tile_X2Y7_S4BEG[8] ,
    \Tile_X2Y7_S4BEG[7] ,
    \Tile_X2Y7_S4BEG[6] ,
    \Tile_X2Y7_S4BEG[5] ,
    \Tile_X2Y7_S4BEG[4] ,
    \Tile_X2Y7_S4BEG[3] ,
    \Tile_X2Y7_S4BEG[2] ,
    \Tile_X2Y7_S4BEG[1] ,
    \Tile_X2Y7_S4BEG[0] }),
    .SS4BEG({\Tile_X2Y8_SS4BEG[15] ,
    \Tile_X2Y8_SS4BEG[14] ,
    \Tile_X2Y8_SS4BEG[13] ,
    \Tile_X2Y8_SS4BEG[12] ,
    \Tile_X2Y8_SS4BEG[11] ,
    \Tile_X2Y8_SS4BEG[10] ,
    \Tile_X2Y8_SS4BEG[9] ,
    \Tile_X2Y8_SS4BEG[8] ,
    \Tile_X2Y8_SS4BEG[7] ,
    \Tile_X2Y8_SS4BEG[6] ,
    \Tile_X2Y8_SS4BEG[5] ,
    \Tile_X2Y8_SS4BEG[4] ,
    \Tile_X2Y8_SS4BEG[3] ,
    \Tile_X2Y8_SS4BEG[2] ,
    \Tile_X2Y8_SS4BEG[1] ,
    \Tile_X2Y8_SS4BEG[0] }),
    .SS4END({\Tile_X2Y7_SS4BEG[15] ,
    \Tile_X2Y7_SS4BEG[14] ,
    \Tile_X2Y7_SS4BEG[13] ,
    \Tile_X2Y7_SS4BEG[12] ,
    \Tile_X2Y7_SS4BEG[11] ,
    \Tile_X2Y7_SS4BEG[10] ,
    \Tile_X2Y7_SS4BEG[9] ,
    \Tile_X2Y7_SS4BEG[8] ,
    \Tile_X2Y7_SS4BEG[7] ,
    \Tile_X2Y7_SS4BEG[6] ,
    \Tile_X2Y7_SS4BEG[5] ,
    \Tile_X2Y7_SS4BEG[4] ,
    \Tile_X2Y7_SS4BEG[3] ,
    \Tile_X2Y7_SS4BEG[2] ,
    \Tile_X2Y7_SS4BEG[1] ,
    \Tile_X2Y7_SS4BEG[0] }),
    .W1BEG({\Tile_X2Y8_W1BEG[3] ,
    \Tile_X2Y8_W1BEG[2] ,
    \Tile_X2Y8_W1BEG[1] ,
    \Tile_X2Y8_W1BEG[0] }),
    .W1END({\Tile_X3Y8_W1BEG[3] ,
    \Tile_X3Y8_W1BEG[2] ,
    \Tile_X3Y8_W1BEG[1] ,
    \Tile_X3Y8_W1BEG[0] }),
    .W2BEG({\Tile_X2Y8_W2BEG[7] ,
    \Tile_X2Y8_W2BEG[6] ,
    \Tile_X2Y8_W2BEG[5] ,
    \Tile_X2Y8_W2BEG[4] ,
    \Tile_X2Y8_W2BEG[3] ,
    \Tile_X2Y8_W2BEG[2] ,
    \Tile_X2Y8_W2BEG[1] ,
    \Tile_X2Y8_W2BEG[0] }),
    .W2BEGb({\Tile_X2Y8_W2BEGb[7] ,
    \Tile_X2Y8_W2BEGb[6] ,
    \Tile_X2Y8_W2BEGb[5] ,
    \Tile_X2Y8_W2BEGb[4] ,
    \Tile_X2Y8_W2BEGb[3] ,
    \Tile_X2Y8_W2BEGb[2] ,
    \Tile_X2Y8_W2BEGb[1] ,
    \Tile_X2Y8_W2BEGb[0] }),
    .W2END({\Tile_X3Y8_W2BEGb[7] ,
    \Tile_X3Y8_W2BEGb[6] ,
    \Tile_X3Y8_W2BEGb[5] ,
    \Tile_X3Y8_W2BEGb[4] ,
    \Tile_X3Y8_W2BEGb[3] ,
    \Tile_X3Y8_W2BEGb[2] ,
    \Tile_X3Y8_W2BEGb[1] ,
    \Tile_X3Y8_W2BEGb[0] }),
    .W2MID({\Tile_X3Y8_W2BEG[7] ,
    \Tile_X3Y8_W2BEG[6] ,
    \Tile_X3Y8_W2BEG[5] ,
    \Tile_X3Y8_W2BEG[4] ,
    \Tile_X3Y8_W2BEG[3] ,
    \Tile_X3Y8_W2BEG[2] ,
    \Tile_X3Y8_W2BEG[1] ,
    \Tile_X3Y8_W2BEG[0] }),
    .W6BEG({\Tile_X2Y8_W6BEG[11] ,
    \Tile_X2Y8_W6BEG[10] ,
    \Tile_X2Y8_W6BEG[9] ,
    \Tile_X2Y8_W6BEG[8] ,
    \Tile_X2Y8_W6BEG[7] ,
    \Tile_X2Y8_W6BEG[6] ,
    \Tile_X2Y8_W6BEG[5] ,
    \Tile_X2Y8_W6BEG[4] ,
    \Tile_X2Y8_W6BEG[3] ,
    \Tile_X2Y8_W6BEG[2] ,
    \Tile_X2Y8_W6BEG[1] ,
    \Tile_X2Y8_W6BEG[0] }),
    .W6END({\Tile_X3Y8_W6BEG[11] ,
    \Tile_X3Y8_W6BEG[10] ,
    \Tile_X3Y8_W6BEG[9] ,
    \Tile_X3Y8_W6BEG[8] ,
    \Tile_X3Y8_W6BEG[7] ,
    \Tile_X3Y8_W6BEG[6] ,
    \Tile_X3Y8_W6BEG[5] ,
    \Tile_X3Y8_W6BEG[4] ,
    \Tile_X3Y8_W6BEG[3] ,
    \Tile_X3Y8_W6BEG[2] ,
    \Tile_X3Y8_W6BEG[1] ,
    \Tile_X3Y8_W6BEG[0] }),
    .WW4BEG({\Tile_X2Y8_WW4BEG[15] ,
    \Tile_X2Y8_WW4BEG[14] ,
    \Tile_X2Y8_WW4BEG[13] ,
    \Tile_X2Y8_WW4BEG[12] ,
    \Tile_X2Y8_WW4BEG[11] ,
    \Tile_X2Y8_WW4BEG[10] ,
    \Tile_X2Y8_WW4BEG[9] ,
    \Tile_X2Y8_WW4BEG[8] ,
    \Tile_X2Y8_WW4BEG[7] ,
    \Tile_X2Y8_WW4BEG[6] ,
    \Tile_X2Y8_WW4BEG[5] ,
    \Tile_X2Y8_WW4BEG[4] ,
    \Tile_X2Y8_WW4BEG[3] ,
    \Tile_X2Y8_WW4BEG[2] ,
    \Tile_X2Y8_WW4BEG[1] ,
    \Tile_X2Y8_WW4BEG[0] }),
    .WW4END({\Tile_X3Y8_WW4BEG[15] ,
    \Tile_X3Y8_WW4BEG[14] ,
    \Tile_X3Y8_WW4BEG[13] ,
    \Tile_X3Y8_WW4BEG[12] ,
    \Tile_X3Y8_WW4BEG[11] ,
    \Tile_X3Y8_WW4BEG[10] ,
    \Tile_X3Y8_WW4BEG[9] ,
    \Tile_X3Y8_WW4BEG[8] ,
    \Tile_X3Y8_WW4BEG[7] ,
    \Tile_X3Y8_WW4BEG[6] ,
    \Tile_X3Y8_WW4BEG[5] ,
    \Tile_X3Y8_WW4BEG[4] ,
    \Tile_X3Y8_WW4BEG[3] ,
    \Tile_X3Y8_WW4BEG[2] ,
    \Tile_X3Y8_WW4BEG[1] ,
    \Tile_X3Y8_WW4BEG[0] }));
 LUT4AB Tile_X2Y9_LUT4AB (.Ci(Tile_X2Y10_Co),
    .Co(Tile_X2Y9_Co),
    .UserCLK(Tile_X2Y10_UserCLKo),
    .UserCLKo(Tile_X2Y9_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X2Y9_E1BEG[3] ,
    \Tile_X2Y9_E1BEG[2] ,
    \Tile_X2Y9_E1BEG[1] ,
    \Tile_X2Y9_E1BEG[0] }),
    .E1END({\Tile_X1Y9_E1BEG[3] ,
    \Tile_X1Y9_E1BEG[2] ,
    \Tile_X1Y9_E1BEG[1] ,
    \Tile_X1Y9_E1BEG[0] }),
    .E2BEG({\Tile_X2Y9_E2BEG[7] ,
    \Tile_X2Y9_E2BEG[6] ,
    \Tile_X2Y9_E2BEG[5] ,
    \Tile_X2Y9_E2BEG[4] ,
    \Tile_X2Y9_E2BEG[3] ,
    \Tile_X2Y9_E2BEG[2] ,
    \Tile_X2Y9_E2BEG[1] ,
    \Tile_X2Y9_E2BEG[0] }),
    .E2BEGb({\Tile_X2Y9_E2BEGb[7] ,
    \Tile_X2Y9_E2BEGb[6] ,
    \Tile_X2Y9_E2BEGb[5] ,
    \Tile_X2Y9_E2BEGb[4] ,
    \Tile_X2Y9_E2BEGb[3] ,
    \Tile_X2Y9_E2BEGb[2] ,
    \Tile_X2Y9_E2BEGb[1] ,
    \Tile_X2Y9_E2BEGb[0] }),
    .E2END({\Tile_X1Y9_E2BEGb[7] ,
    \Tile_X1Y9_E2BEGb[6] ,
    \Tile_X1Y9_E2BEGb[5] ,
    \Tile_X1Y9_E2BEGb[4] ,
    \Tile_X1Y9_E2BEGb[3] ,
    \Tile_X1Y9_E2BEGb[2] ,
    \Tile_X1Y9_E2BEGb[1] ,
    \Tile_X1Y9_E2BEGb[0] }),
    .E2MID({\Tile_X1Y9_E2BEG[7] ,
    \Tile_X1Y9_E2BEG[6] ,
    \Tile_X1Y9_E2BEG[5] ,
    \Tile_X1Y9_E2BEG[4] ,
    \Tile_X1Y9_E2BEG[3] ,
    \Tile_X1Y9_E2BEG[2] ,
    \Tile_X1Y9_E2BEG[1] ,
    \Tile_X1Y9_E2BEG[0] }),
    .E6BEG({\Tile_X2Y9_E6BEG[11] ,
    \Tile_X2Y9_E6BEG[10] ,
    \Tile_X2Y9_E6BEG[9] ,
    \Tile_X2Y9_E6BEG[8] ,
    \Tile_X2Y9_E6BEG[7] ,
    \Tile_X2Y9_E6BEG[6] ,
    \Tile_X2Y9_E6BEG[5] ,
    \Tile_X2Y9_E6BEG[4] ,
    \Tile_X2Y9_E6BEG[3] ,
    \Tile_X2Y9_E6BEG[2] ,
    \Tile_X2Y9_E6BEG[1] ,
    \Tile_X2Y9_E6BEG[0] }),
    .E6END({\Tile_X1Y9_E6BEG[11] ,
    \Tile_X1Y9_E6BEG[10] ,
    \Tile_X1Y9_E6BEG[9] ,
    \Tile_X1Y9_E6BEG[8] ,
    \Tile_X1Y9_E6BEG[7] ,
    \Tile_X1Y9_E6BEG[6] ,
    \Tile_X1Y9_E6BEG[5] ,
    \Tile_X1Y9_E6BEG[4] ,
    \Tile_X1Y9_E6BEG[3] ,
    \Tile_X1Y9_E6BEG[2] ,
    \Tile_X1Y9_E6BEG[1] ,
    \Tile_X1Y9_E6BEG[0] }),
    .EE4BEG({\Tile_X2Y9_EE4BEG[15] ,
    \Tile_X2Y9_EE4BEG[14] ,
    \Tile_X2Y9_EE4BEG[13] ,
    \Tile_X2Y9_EE4BEG[12] ,
    \Tile_X2Y9_EE4BEG[11] ,
    \Tile_X2Y9_EE4BEG[10] ,
    \Tile_X2Y9_EE4BEG[9] ,
    \Tile_X2Y9_EE4BEG[8] ,
    \Tile_X2Y9_EE4BEG[7] ,
    \Tile_X2Y9_EE4BEG[6] ,
    \Tile_X2Y9_EE4BEG[5] ,
    \Tile_X2Y9_EE4BEG[4] ,
    \Tile_X2Y9_EE4BEG[3] ,
    \Tile_X2Y9_EE4BEG[2] ,
    \Tile_X2Y9_EE4BEG[1] ,
    \Tile_X2Y9_EE4BEG[0] }),
    .EE4END({\Tile_X1Y9_EE4BEG[15] ,
    \Tile_X1Y9_EE4BEG[14] ,
    \Tile_X1Y9_EE4BEG[13] ,
    \Tile_X1Y9_EE4BEG[12] ,
    \Tile_X1Y9_EE4BEG[11] ,
    \Tile_X1Y9_EE4BEG[10] ,
    \Tile_X1Y9_EE4BEG[9] ,
    \Tile_X1Y9_EE4BEG[8] ,
    \Tile_X1Y9_EE4BEG[7] ,
    \Tile_X1Y9_EE4BEG[6] ,
    \Tile_X1Y9_EE4BEG[5] ,
    \Tile_X1Y9_EE4BEG[4] ,
    \Tile_X1Y9_EE4BEG[3] ,
    \Tile_X1Y9_EE4BEG[2] ,
    \Tile_X1Y9_EE4BEG[1] ,
    \Tile_X1Y9_EE4BEG[0] }),
    .FrameData({\Tile_X1Y9_FrameData_O[31] ,
    \Tile_X1Y9_FrameData_O[30] ,
    \Tile_X1Y9_FrameData_O[29] ,
    \Tile_X1Y9_FrameData_O[28] ,
    \Tile_X1Y9_FrameData_O[27] ,
    \Tile_X1Y9_FrameData_O[26] ,
    \Tile_X1Y9_FrameData_O[25] ,
    \Tile_X1Y9_FrameData_O[24] ,
    \Tile_X1Y9_FrameData_O[23] ,
    \Tile_X1Y9_FrameData_O[22] ,
    \Tile_X1Y9_FrameData_O[21] ,
    \Tile_X1Y9_FrameData_O[20] ,
    \Tile_X1Y9_FrameData_O[19] ,
    \Tile_X1Y9_FrameData_O[18] ,
    \Tile_X1Y9_FrameData_O[17] ,
    \Tile_X1Y9_FrameData_O[16] ,
    \Tile_X1Y9_FrameData_O[15] ,
    \Tile_X1Y9_FrameData_O[14] ,
    \Tile_X1Y9_FrameData_O[13] ,
    \Tile_X1Y9_FrameData_O[12] ,
    \Tile_X1Y9_FrameData_O[11] ,
    \Tile_X1Y9_FrameData_O[10] ,
    \Tile_X1Y9_FrameData_O[9] ,
    \Tile_X1Y9_FrameData_O[8] ,
    \Tile_X1Y9_FrameData_O[7] ,
    \Tile_X1Y9_FrameData_O[6] ,
    \Tile_X1Y9_FrameData_O[5] ,
    \Tile_X1Y9_FrameData_O[4] ,
    \Tile_X1Y9_FrameData_O[3] ,
    \Tile_X1Y9_FrameData_O[2] ,
    \Tile_X1Y9_FrameData_O[1] ,
    \Tile_X1Y9_FrameData_O[0] }),
    .FrameData_O({\Tile_X2Y9_FrameData_O[31] ,
    \Tile_X2Y9_FrameData_O[30] ,
    \Tile_X2Y9_FrameData_O[29] ,
    \Tile_X2Y9_FrameData_O[28] ,
    \Tile_X2Y9_FrameData_O[27] ,
    \Tile_X2Y9_FrameData_O[26] ,
    \Tile_X2Y9_FrameData_O[25] ,
    \Tile_X2Y9_FrameData_O[24] ,
    \Tile_X2Y9_FrameData_O[23] ,
    \Tile_X2Y9_FrameData_O[22] ,
    \Tile_X2Y9_FrameData_O[21] ,
    \Tile_X2Y9_FrameData_O[20] ,
    \Tile_X2Y9_FrameData_O[19] ,
    \Tile_X2Y9_FrameData_O[18] ,
    \Tile_X2Y9_FrameData_O[17] ,
    \Tile_X2Y9_FrameData_O[16] ,
    \Tile_X2Y9_FrameData_O[15] ,
    \Tile_X2Y9_FrameData_O[14] ,
    \Tile_X2Y9_FrameData_O[13] ,
    \Tile_X2Y9_FrameData_O[12] ,
    \Tile_X2Y9_FrameData_O[11] ,
    \Tile_X2Y9_FrameData_O[10] ,
    \Tile_X2Y9_FrameData_O[9] ,
    \Tile_X2Y9_FrameData_O[8] ,
    \Tile_X2Y9_FrameData_O[7] ,
    \Tile_X2Y9_FrameData_O[6] ,
    \Tile_X2Y9_FrameData_O[5] ,
    \Tile_X2Y9_FrameData_O[4] ,
    \Tile_X2Y9_FrameData_O[3] ,
    \Tile_X2Y9_FrameData_O[2] ,
    \Tile_X2Y9_FrameData_O[1] ,
    \Tile_X2Y9_FrameData_O[0] }),
    .FrameStrobe({\Tile_X2Y10_FrameStrobe_O[19] ,
    \Tile_X2Y10_FrameStrobe_O[18] ,
    \Tile_X2Y10_FrameStrobe_O[17] ,
    \Tile_X2Y10_FrameStrobe_O[16] ,
    \Tile_X2Y10_FrameStrobe_O[15] ,
    \Tile_X2Y10_FrameStrobe_O[14] ,
    \Tile_X2Y10_FrameStrobe_O[13] ,
    \Tile_X2Y10_FrameStrobe_O[12] ,
    \Tile_X2Y10_FrameStrobe_O[11] ,
    \Tile_X2Y10_FrameStrobe_O[10] ,
    \Tile_X2Y10_FrameStrobe_O[9] ,
    \Tile_X2Y10_FrameStrobe_O[8] ,
    \Tile_X2Y10_FrameStrobe_O[7] ,
    \Tile_X2Y10_FrameStrobe_O[6] ,
    \Tile_X2Y10_FrameStrobe_O[5] ,
    \Tile_X2Y10_FrameStrobe_O[4] ,
    \Tile_X2Y10_FrameStrobe_O[3] ,
    \Tile_X2Y10_FrameStrobe_O[2] ,
    \Tile_X2Y10_FrameStrobe_O[1] ,
    \Tile_X2Y10_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X2Y9_FrameStrobe_O[19] ,
    \Tile_X2Y9_FrameStrobe_O[18] ,
    \Tile_X2Y9_FrameStrobe_O[17] ,
    \Tile_X2Y9_FrameStrobe_O[16] ,
    \Tile_X2Y9_FrameStrobe_O[15] ,
    \Tile_X2Y9_FrameStrobe_O[14] ,
    \Tile_X2Y9_FrameStrobe_O[13] ,
    \Tile_X2Y9_FrameStrobe_O[12] ,
    \Tile_X2Y9_FrameStrobe_O[11] ,
    \Tile_X2Y9_FrameStrobe_O[10] ,
    \Tile_X2Y9_FrameStrobe_O[9] ,
    \Tile_X2Y9_FrameStrobe_O[8] ,
    \Tile_X2Y9_FrameStrobe_O[7] ,
    \Tile_X2Y9_FrameStrobe_O[6] ,
    \Tile_X2Y9_FrameStrobe_O[5] ,
    \Tile_X2Y9_FrameStrobe_O[4] ,
    \Tile_X2Y9_FrameStrobe_O[3] ,
    \Tile_X2Y9_FrameStrobe_O[2] ,
    \Tile_X2Y9_FrameStrobe_O[1] ,
    \Tile_X2Y9_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X2Y9_N1BEG[3] ,
    \Tile_X2Y9_N1BEG[2] ,
    \Tile_X2Y9_N1BEG[1] ,
    \Tile_X2Y9_N1BEG[0] }),
    .N1END({\Tile_X2Y10_N1BEG[3] ,
    \Tile_X2Y10_N1BEG[2] ,
    \Tile_X2Y10_N1BEG[1] ,
    \Tile_X2Y10_N1BEG[0] }),
    .N2BEG({\Tile_X2Y9_N2BEG[7] ,
    \Tile_X2Y9_N2BEG[6] ,
    \Tile_X2Y9_N2BEG[5] ,
    \Tile_X2Y9_N2BEG[4] ,
    \Tile_X2Y9_N2BEG[3] ,
    \Tile_X2Y9_N2BEG[2] ,
    \Tile_X2Y9_N2BEG[1] ,
    \Tile_X2Y9_N2BEG[0] }),
    .N2BEGb({\Tile_X2Y9_N2BEGb[7] ,
    \Tile_X2Y9_N2BEGb[6] ,
    \Tile_X2Y9_N2BEGb[5] ,
    \Tile_X2Y9_N2BEGb[4] ,
    \Tile_X2Y9_N2BEGb[3] ,
    \Tile_X2Y9_N2BEGb[2] ,
    \Tile_X2Y9_N2BEGb[1] ,
    \Tile_X2Y9_N2BEGb[0] }),
    .N2END({\Tile_X2Y10_N2BEGb[7] ,
    \Tile_X2Y10_N2BEGb[6] ,
    \Tile_X2Y10_N2BEGb[5] ,
    \Tile_X2Y10_N2BEGb[4] ,
    \Tile_X2Y10_N2BEGb[3] ,
    \Tile_X2Y10_N2BEGb[2] ,
    \Tile_X2Y10_N2BEGb[1] ,
    \Tile_X2Y10_N2BEGb[0] }),
    .N2MID({\Tile_X2Y10_N2BEG[7] ,
    \Tile_X2Y10_N2BEG[6] ,
    \Tile_X2Y10_N2BEG[5] ,
    \Tile_X2Y10_N2BEG[4] ,
    \Tile_X2Y10_N2BEG[3] ,
    \Tile_X2Y10_N2BEG[2] ,
    \Tile_X2Y10_N2BEG[1] ,
    \Tile_X2Y10_N2BEG[0] }),
    .N4BEG({\Tile_X2Y9_N4BEG[15] ,
    \Tile_X2Y9_N4BEG[14] ,
    \Tile_X2Y9_N4BEG[13] ,
    \Tile_X2Y9_N4BEG[12] ,
    \Tile_X2Y9_N4BEG[11] ,
    \Tile_X2Y9_N4BEG[10] ,
    \Tile_X2Y9_N4BEG[9] ,
    \Tile_X2Y9_N4BEG[8] ,
    \Tile_X2Y9_N4BEG[7] ,
    \Tile_X2Y9_N4BEG[6] ,
    \Tile_X2Y9_N4BEG[5] ,
    \Tile_X2Y9_N4BEG[4] ,
    \Tile_X2Y9_N4BEG[3] ,
    \Tile_X2Y9_N4BEG[2] ,
    \Tile_X2Y9_N4BEG[1] ,
    \Tile_X2Y9_N4BEG[0] }),
    .N4END({\Tile_X2Y10_N4BEG[15] ,
    \Tile_X2Y10_N4BEG[14] ,
    \Tile_X2Y10_N4BEG[13] ,
    \Tile_X2Y10_N4BEG[12] ,
    \Tile_X2Y10_N4BEG[11] ,
    \Tile_X2Y10_N4BEG[10] ,
    \Tile_X2Y10_N4BEG[9] ,
    \Tile_X2Y10_N4BEG[8] ,
    \Tile_X2Y10_N4BEG[7] ,
    \Tile_X2Y10_N4BEG[6] ,
    \Tile_X2Y10_N4BEG[5] ,
    \Tile_X2Y10_N4BEG[4] ,
    \Tile_X2Y10_N4BEG[3] ,
    \Tile_X2Y10_N4BEG[2] ,
    \Tile_X2Y10_N4BEG[1] ,
    \Tile_X2Y10_N4BEG[0] }),
    .NN4BEG({\Tile_X2Y9_NN4BEG[15] ,
    \Tile_X2Y9_NN4BEG[14] ,
    \Tile_X2Y9_NN4BEG[13] ,
    \Tile_X2Y9_NN4BEG[12] ,
    \Tile_X2Y9_NN4BEG[11] ,
    \Tile_X2Y9_NN4BEG[10] ,
    \Tile_X2Y9_NN4BEG[9] ,
    \Tile_X2Y9_NN4BEG[8] ,
    \Tile_X2Y9_NN4BEG[7] ,
    \Tile_X2Y9_NN4BEG[6] ,
    \Tile_X2Y9_NN4BEG[5] ,
    \Tile_X2Y9_NN4BEG[4] ,
    \Tile_X2Y9_NN4BEG[3] ,
    \Tile_X2Y9_NN4BEG[2] ,
    \Tile_X2Y9_NN4BEG[1] ,
    \Tile_X2Y9_NN4BEG[0] }),
    .NN4END({\Tile_X2Y10_NN4BEG[15] ,
    \Tile_X2Y10_NN4BEG[14] ,
    \Tile_X2Y10_NN4BEG[13] ,
    \Tile_X2Y10_NN4BEG[12] ,
    \Tile_X2Y10_NN4BEG[11] ,
    \Tile_X2Y10_NN4BEG[10] ,
    \Tile_X2Y10_NN4BEG[9] ,
    \Tile_X2Y10_NN4BEG[8] ,
    \Tile_X2Y10_NN4BEG[7] ,
    \Tile_X2Y10_NN4BEG[6] ,
    \Tile_X2Y10_NN4BEG[5] ,
    \Tile_X2Y10_NN4BEG[4] ,
    \Tile_X2Y10_NN4BEG[3] ,
    \Tile_X2Y10_NN4BEG[2] ,
    \Tile_X2Y10_NN4BEG[1] ,
    \Tile_X2Y10_NN4BEG[0] }),
    .S1BEG({\Tile_X2Y9_S1BEG[3] ,
    \Tile_X2Y9_S1BEG[2] ,
    \Tile_X2Y9_S1BEG[1] ,
    \Tile_X2Y9_S1BEG[0] }),
    .S1END({\Tile_X2Y8_S1BEG[3] ,
    \Tile_X2Y8_S1BEG[2] ,
    \Tile_X2Y8_S1BEG[1] ,
    \Tile_X2Y8_S1BEG[0] }),
    .S2BEG({\Tile_X2Y9_S2BEG[7] ,
    \Tile_X2Y9_S2BEG[6] ,
    \Tile_X2Y9_S2BEG[5] ,
    \Tile_X2Y9_S2BEG[4] ,
    \Tile_X2Y9_S2BEG[3] ,
    \Tile_X2Y9_S2BEG[2] ,
    \Tile_X2Y9_S2BEG[1] ,
    \Tile_X2Y9_S2BEG[0] }),
    .S2BEGb({\Tile_X2Y9_S2BEGb[7] ,
    \Tile_X2Y9_S2BEGb[6] ,
    \Tile_X2Y9_S2BEGb[5] ,
    \Tile_X2Y9_S2BEGb[4] ,
    \Tile_X2Y9_S2BEGb[3] ,
    \Tile_X2Y9_S2BEGb[2] ,
    \Tile_X2Y9_S2BEGb[1] ,
    \Tile_X2Y9_S2BEGb[0] }),
    .S2END({\Tile_X2Y8_S2BEGb[7] ,
    \Tile_X2Y8_S2BEGb[6] ,
    \Tile_X2Y8_S2BEGb[5] ,
    \Tile_X2Y8_S2BEGb[4] ,
    \Tile_X2Y8_S2BEGb[3] ,
    \Tile_X2Y8_S2BEGb[2] ,
    \Tile_X2Y8_S2BEGb[1] ,
    \Tile_X2Y8_S2BEGb[0] }),
    .S2MID({\Tile_X2Y8_S2BEG[7] ,
    \Tile_X2Y8_S2BEG[6] ,
    \Tile_X2Y8_S2BEG[5] ,
    \Tile_X2Y8_S2BEG[4] ,
    \Tile_X2Y8_S2BEG[3] ,
    \Tile_X2Y8_S2BEG[2] ,
    \Tile_X2Y8_S2BEG[1] ,
    \Tile_X2Y8_S2BEG[0] }),
    .S4BEG({\Tile_X2Y9_S4BEG[15] ,
    \Tile_X2Y9_S4BEG[14] ,
    \Tile_X2Y9_S4BEG[13] ,
    \Tile_X2Y9_S4BEG[12] ,
    \Tile_X2Y9_S4BEG[11] ,
    \Tile_X2Y9_S4BEG[10] ,
    \Tile_X2Y9_S4BEG[9] ,
    \Tile_X2Y9_S4BEG[8] ,
    \Tile_X2Y9_S4BEG[7] ,
    \Tile_X2Y9_S4BEG[6] ,
    \Tile_X2Y9_S4BEG[5] ,
    \Tile_X2Y9_S4BEG[4] ,
    \Tile_X2Y9_S4BEG[3] ,
    \Tile_X2Y9_S4BEG[2] ,
    \Tile_X2Y9_S4BEG[1] ,
    \Tile_X2Y9_S4BEG[0] }),
    .S4END({\Tile_X2Y8_S4BEG[15] ,
    \Tile_X2Y8_S4BEG[14] ,
    \Tile_X2Y8_S4BEG[13] ,
    \Tile_X2Y8_S4BEG[12] ,
    \Tile_X2Y8_S4BEG[11] ,
    \Tile_X2Y8_S4BEG[10] ,
    \Tile_X2Y8_S4BEG[9] ,
    \Tile_X2Y8_S4BEG[8] ,
    \Tile_X2Y8_S4BEG[7] ,
    \Tile_X2Y8_S4BEG[6] ,
    \Tile_X2Y8_S4BEG[5] ,
    \Tile_X2Y8_S4BEG[4] ,
    \Tile_X2Y8_S4BEG[3] ,
    \Tile_X2Y8_S4BEG[2] ,
    \Tile_X2Y8_S4BEG[1] ,
    \Tile_X2Y8_S4BEG[0] }),
    .SS4BEG({\Tile_X2Y9_SS4BEG[15] ,
    \Tile_X2Y9_SS4BEG[14] ,
    \Tile_X2Y9_SS4BEG[13] ,
    \Tile_X2Y9_SS4BEG[12] ,
    \Tile_X2Y9_SS4BEG[11] ,
    \Tile_X2Y9_SS4BEG[10] ,
    \Tile_X2Y9_SS4BEG[9] ,
    \Tile_X2Y9_SS4BEG[8] ,
    \Tile_X2Y9_SS4BEG[7] ,
    \Tile_X2Y9_SS4BEG[6] ,
    \Tile_X2Y9_SS4BEG[5] ,
    \Tile_X2Y9_SS4BEG[4] ,
    \Tile_X2Y9_SS4BEG[3] ,
    \Tile_X2Y9_SS4BEG[2] ,
    \Tile_X2Y9_SS4BEG[1] ,
    \Tile_X2Y9_SS4BEG[0] }),
    .SS4END({\Tile_X2Y8_SS4BEG[15] ,
    \Tile_X2Y8_SS4BEG[14] ,
    \Tile_X2Y8_SS4BEG[13] ,
    \Tile_X2Y8_SS4BEG[12] ,
    \Tile_X2Y8_SS4BEG[11] ,
    \Tile_X2Y8_SS4BEG[10] ,
    \Tile_X2Y8_SS4BEG[9] ,
    \Tile_X2Y8_SS4BEG[8] ,
    \Tile_X2Y8_SS4BEG[7] ,
    \Tile_X2Y8_SS4BEG[6] ,
    \Tile_X2Y8_SS4BEG[5] ,
    \Tile_X2Y8_SS4BEG[4] ,
    \Tile_X2Y8_SS4BEG[3] ,
    \Tile_X2Y8_SS4BEG[2] ,
    \Tile_X2Y8_SS4BEG[1] ,
    \Tile_X2Y8_SS4BEG[0] }),
    .W1BEG({\Tile_X2Y9_W1BEG[3] ,
    \Tile_X2Y9_W1BEG[2] ,
    \Tile_X2Y9_W1BEG[1] ,
    \Tile_X2Y9_W1BEG[0] }),
    .W1END({\Tile_X3Y9_W1BEG[3] ,
    \Tile_X3Y9_W1BEG[2] ,
    \Tile_X3Y9_W1BEG[1] ,
    \Tile_X3Y9_W1BEG[0] }),
    .W2BEG({\Tile_X2Y9_W2BEG[7] ,
    \Tile_X2Y9_W2BEG[6] ,
    \Tile_X2Y9_W2BEG[5] ,
    \Tile_X2Y9_W2BEG[4] ,
    \Tile_X2Y9_W2BEG[3] ,
    \Tile_X2Y9_W2BEG[2] ,
    \Tile_X2Y9_W2BEG[1] ,
    \Tile_X2Y9_W2BEG[0] }),
    .W2BEGb({\Tile_X2Y9_W2BEGb[7] ,
    \Tile_X2Y9_W2BEGb[6] ,
    \Tile_X2Y9_W2BEGb[5] ,
    \Tile_X2Y9_W2BEGb[4] ,
    \Tile_X2Y9_W2BEGb[3] ,
    \Tile_X2Y9_W2BEGb[2] ,
    \Tile_X2Y9_W2BEGb[1] ,
    \Tile_X2Y9_W2BEGb[0] }),
    .W2END({\Tile_X3Y9_W2BEGb[7] ,
    \Tile_X3Y9_W2BEGb[6] ,
    \Tile_X3Y9_W2BEGb[5] ,
    \Tile_X3Y9_W2BEGb[4] ,
    \Tile_X3Y9_W2BEGb[3] ,
    \Tile_X3Y9_W2BEGb[2] ,
    \Tile_X3Y9_W2BEGb[1] ,
    \Tile_X3Y9_W2BEGb[0] }),
    .W2MID({\Tile_X3Y9_W2BEG[7] ,
    \Tile_X3Y9_W2BEG[6] ,
    \Tile_X3Y9_W2BEG[5] ,
    \Tile_X3Y9_W2BEG[4] ,
    \Tile_X3Y9_W2BEG[3] ,
    \Tile_X3Y9_W2BEG[2] ,
    \Tile_X3Y9_W2BEG[1] ,
    \Tile_X3Y9_W2BEG[0] }),
    .W6BEG({\Tile_X2Y9_W6BEG[11] ,
    \Tile_X2Y9_W6BEG[10] ,
    \Tile_X2Y9_W6BEG[9] ,
    \Tile_X2Y9_W6BEG[8] ,
    \Tile_X2Y9_W6BEG[7] ,
    \Tile_X2Y9_W6BEG[6] ,
    \Tile_X2Y9_W6BEG[5] ,
    \Tile_X2Y9_W6BEG[4] ,
    \Tile_X2Y9_W6BEG[3] ,
    \Tile_X2Y9_W6BEG[2] ,
    \Tile_X2Y9_W6BEG[1] ,
    \Tile_X2Y9_W6BEG[0] }),
    .W6END({\Tile_X3Y9_W6BEG[11] ,
    \Tile_X3Y9_W6BEG[10] ,
    \Tile_X3Y9_W6BEG[9] ,
    \Tile_X3Y9_W6BEG[8] ,
    \Tile_X3Y9_W6BEG[7] ,
    \Tile_X3Y9_W6BEG[6] ,
    \Tile_X3Y9_W6BEG[5] ,
    \Tile_X3Y9_W6BEG[4] ,
    \Tile_X3Y9_W6BEG[3] ,
    \Tile_X3Y9_W6BEG[2] ,
    \Tile_X3Y9_W6BEG[1] ,
    \Tile_X3Y9_W6BEG[0] }),
    .WW4BEG({\Tile_X2Y9_WW4BEG[15] ,
    \Tile_X2Y9_WW4BEG[14] ,
    \Tile_X2Y9_WW4BEG[13] ,
    \Tile_X2Y9_WW4BEG[12] ,
    \Tile_X2Y9_WW4BEG[11] ,
    \Tile_X2Y9_WW4BEG[10] ,
    \Tile_X2Y9_WW4BEG[9] ,
    \Tile_X2Y9_WW4BEG[8] ,
    \Tile_X2Y9_WW4BEG[7] ,
    \Tile_X2Y9_WW4BEG[6] ,
    \Tile_X2Y9_WW4BEG[5] ,
    \Tile_X2Y9_WW4BEG[4] ,
    \Tile_X2Y9_WW4BEG[3] ,
    \Tile_X2Y9_WW4BEG[2] ,
    \Tile_X2Y9_WW4BEG[1] ,
    \Tile_X2Y9_WW4BEG[0] }),
    .WW4END({\Tile_X3Y9_WW4BEG[15] ,
    \Tile_X3Y9_WW4BEG[14] ,
    \Tile_X3Y9_WW4BEG[13] ,
    \Tile_X3Y9_WW4BEG[12] ,
    \Tile_X3Y9_WW4BEG[11] ,
    \Tile_X3Y9_WW4BEG[10] ,
    \Tile_X3Y9_WW4BEG[9] ,
    \Tile_X3Y9_WW4BEG[8] ,
    \Tile_X3Y9_WW4BEG[7] ,
    \Tile_X3Y9_WW4BEG[6] ,
    \Tile_X3Y9_WW4BEG[5] ,
    \Tile_X3Y9_WW4BEG[4] ,
    \Tile_X3Y9_WW4BEG[3] ,
    \Tile_X3Y9_WW4BEG[2] ,
    \Tile_X3Y9_WW4BEG[1] ,
    \Tile_X3Y9_WW4BEG[0] }));
 N_term_single Tile_X3Y0_N_term_single (.Ci(Tile_X3Y1_Co),
    .UserCLK(Tile_X3Y1_UserCLKo),
    .UserCLKo(Tile_X3Y0_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .FrameData({\Tile_X2Y0_FrameData_O[31] ,
    \Tile_X2Y0_FrameData_O[30] ,
    \Tile_X2Y0_FrameData_O[29] ,
    \Tile_X2Y0_FrameData_O[28] ,
    \Tile_X2Y0_FrameData_O[27] ,
    \Tile_X2Y0_FrameData_O[26] ,
    \Tile_X2Y0_FrameData_O[25] ,
    \Tile_X2Y0_FrameData_O[24] ,
    \Tile_X2Y0_FrameData_O[23] ,
    \Tile_X2Y0_FrameData_O[22] ,
    \Tile_X2Y0_FrameData_O[21] ,
    \Tile_X2Y0_FrameData_O[20] ,
    \Tile_X2Y0_FrameData_O[19] ,
    \Tile_X2Y0_FrameData_O[18] ,
    \Tile_X2Y0_FrameData_O[17] ,
    \Tile_X2Y0_FrameData_O[16] ,
    \Tile_X2Y0_FrameData_O[15] ,
    \Tile_X2Y0_FrameData_O[14] ,
    \Tile_X2Y0_FrameData_O[13] ,
    \Tile_X2Y0_FrameData_O[12] ,
    \Tile_X2Y0_FrameData_O[11] ,
    \Tile_X2Y0_FrameData_O[10] ,
    \Tile_X2Y0_FrameData_O[9] ,
    \Tile_X2Y0_FrameData_O[8] ,
    \Tile_X2Y0_FrameData_O[7] ,
    \Tile_X2Y0_FrameData_O[6] ,
    \Tile_X2Y0_FrameData_O[5] ,
    \Tile_X2Y0_FrameData_O[4] ,
    \Tile_X2Y0_FrameData_O[3] ,
    \Tile_X2Y0_FrameData_O[2] ,
    \Tile_X2Y0_FrameData_O[1] ,
    \Tile_X2Y0_FrameData_O[0] }),
    .FrameData_O({\Tile_X3Y0_FrameData_O[31] ,
    \Tile_X3Y0_FrameData_O[30] ,
    \Tile_X3Y0_FrameData_O[29] ,
    \Tile_X3Y0_FrameData_O[28] ,
    \Tile_X3Y0_FrameData_O[27] ,
    \Tile_X3Y0_FrameData_O[26] ,
    \Tile_X3Y0_FrameData_O[25] ,
    \Tile_X3Y0_FrameData_O[24] ,
    \Tile_X3Y0_FrameData_O[23] ,
    \Tile_X3Y0_FrameData_O[22] ,
    \Tile_X3Y0_FrameData_O[21] ,
    \Tile_X3Y0_FrameData_O[20] ,
    \Tile_X3Y0_FrameData_O[19] ,
    \Tile_X3Y0_FrameData_O[18] ,
    \Tile_X3Y0_FrameData_O[17] ,
    \Tile_X3Y0_FrameData_O[16] ,
    \Tile_X3Y0_FrameData_O[15] ,
    \Tile_X3Y0_FrameData_O[14] ,
    \Tile_X3Y0_FrameData_O[13] ,
    \Tile_X3Y0_FrameData_O[12] ,
    \Tile_X3Y0_FrameData_O[11] ,
    \Tile_X3Y0_FrameData_O[10] ,
    \Tile_X3Y0_FrameData_O[9] ,
    \Tile_X3Y0_FrameData_O[8] ,
    \Tile_X3Y0_FrameData_O[7] ,
    \Tile_X3Y0_FrameData_O[6] ,
    \Tile_X3Y0_FrameData_O[5] ,
    \Tile_X3Y0_FrameData_O[4] ,
    \Tile_X3Y0_FrameData_O[3] ,
    \Tile_X3Y0_FrameData_O[2] ,
    \Tile_X3Y0_FrameData_O[1] ,
    \Tile_X3Y0_FrameData_O[0] }),
    .FrameStrobe({\Tile_X3Y1_FrameStrobe_O[19] ,
    \Tile_X3Y1_FrameStrobe_O[18] ,
    \Tile_X3Y1_FrameStrobe_O[17] ,
    \Tile_X3Y1_FrameStrobe_O[16] ,
    \Tile_X3Y1_FrameStrobe_O[15] ,
    \Tile_X3Y1_FrameStrobe_O[14] ,
    \Tile_X3Y1_FrameStrobe_O[13] ,
    \Tile_X3Y1_FrameStrobe_O[12] ,
    \Tile_X3Y1_FrameStrobe_O[11] ,
    \Tile_X3Y1_FrameStrobe_O[10] ,
    \Tile_X3Y1_FrameStrobe_O[9] ,
    \Tile_X3Y1_FrameStrobe_O[8] ,
    \Tile_X3Y1_FrameStrobe_O[7] ,
    \Tile_X3Y1_FrameStrobe_O[6] ,
    \Tile_X3Y1_FrameStrobe_O[5] ,
    \Tile_X3Y1_FrameStrobe_O[4] ,
    \Tile_X3Y1_FrameStrobe_O[3] ,
    \Tile_X3Y1_FrameStrobe_O[2] ,
    \Tile_X3Y1_FrameStrobe_O[1] ,
    \Tile_X3Y1_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X3Y0_FrameStrobe_O[19] ,
    \Tile_X3Y0_FrameStrobe_O[18] ,
    \Tile_X3Y0_FrameStrobe_O[17] ,
    \Tile_X3Y0_FrameStrobe_O[16] ,
    \Tile_X3Y0_FrameStrobe_O[15] ,
    \Tile_X3Y0_FrameStrobe_O[14] ,
    \Tile_X3Y0_FrameStrobe_O[13] ,
    \Tile_X3Y0_FrameStrobe_O[12] ,
    \Tile_X3Y0_FrameStrobe_O[11] ,
    \Tile_X3Y0_FrameStrobe_O[10] ,
    \Tile_X3Y0_FrameStrobe_O[9] ,
    \Tile_X3Y0_FrameStrobe_O[8] ,
    \Tile_X3Y0_FrameStrobe_O[7] ,
    \Tile_X3Y0_FrameStrobe_O[6] ,
    \Tile_X3Y0_FrameStrobe_O[5] ,
    \Tile_X3Y0_FrameStrobe_O[4] ,
    \Tile_X3Y0_FrameStrobe_O[3] ,
    \Tile_X3Y0_FrameStrobe_O[2] ,
    \Tile_X3Y0_FrameStrobe_O[1] ,
    \Tile_X3Y0_FrameStrobe_O[0] }),
    .N1END({\Tile_X3Y1_N1BEG[3] ,
    \Tile_X3Y1_N1BEG[2] ,
    \Tile_X3Y1_N1BEG[1] ,
    \Tile_X3Y1_N1BEG[0] }),
    .N2END({\Tile_X3Y1_N2BEGb[7] ,
    \Tile_X3Y1_N2BEGb[6] ,
    \Tile_X3Y1_N2BEGb[5] ,
    \Tile_X3Y1_N2BEGb[4] ,
    \Tile_X3Y1_N2BEGb[3] ,
    \Tile_X3Y1_N2BEGb[2] ,
    \Tile_X3Y1_N2BEGb[1] ,
    \Tile_X3Y1_N2BEGb[0] }),
    .N2MID({\Tile_X3Y1_N2BEG[7] ,
    \Tile_X3Y1_N2BEG[6] ,
    \Tile_X3Y1_N2BEG[5] ,
    \Tile_X3Y1_N2BEG[4] ,
    \Tile_X3Y1_N2BEG[3] ,
    \Tile_X3Y1_N2BEG[2] ,
    \Tile_X3Y1_N2BEG[1] ,
    \Tile_X3Y1_N2BEG[0] }),
    .N4END({\Tile_X3Y1_N4BEG[15] ,
    \Tile_X3Y1_N4BEG[14] ,
    \Tile_X3Y1_N4BEG[13] ,
    \Tile_X3Y1_N4BEG[12] ,
    \Tile_X3Y1_N4BEG[11] ,
    \Tile_X3Y1_N4BEG[10] ,
    \Tile_X3Y1_N4BEG[9] ,
    \Tile_X3Y1_N4BEG[8] ,
    \Tile_X3Y1_N4BEG[7] ,
    \Tile_X3Y1_N4BEG[6] ,
    \Tile_X3Y1_N4BEG[5] ,
    \Tile_X3Y1_N4BEG[4] ,
    \Tile_X3Y1_N4BEG[3] ,
    \Tile_X3Y1_N4BEG[2] ,
    \Tile_X3Y1_N4BEG[1] ,
    \Tile_X3Y1_N4BEG[0] }),
    .NN4END({\Tile_X3Y1_NN4BEG[15] ,
    \Tile_X3Y1_NN4BEG[14] ,
    \Tile_X3Y1_NN4BEG[13] ,
    \Tile_X3Y1_NN4BEG[12] ,
    \Tile_X3Y1_NN4BEG[11] ,
    \Tile_X3Y1_NN4BEG[10] ,
    \Tile_X3Y1_NN4BEG[9] ,
    \Tile_X3Y1_NN4BEG[8] ,
    \Tile_X3Y1_NN4BEG[7] ,
    \Tile_X3Y1_NN4BEG[6] ,
    \Tile_X3Y1_NN4BEG[5] ,
    \Tile_X3Y1_NN4BEG[4] ,
    \Tile_X3Y1_NN4BEG[3] ,
    \Tile_X3Y1_NN4BEG[2] ,
    \Tile_X3Y1_NN4BEG[1] ,
    \Tile_X3Y1_NN4BEG[0] }),
    .S1BEG({\Tile_X3Y0_S1BEG[3] ,
    \Tile_X3Y0_S1BEG[2] ,
    \Tile_X3Y0_S1BEG[1] ,
    \Tile_X3Y0_S1BEG[0] }),
    .S2BEG({\Tile_X3Y0_S2BEG[7] ,
    \Tile_X3Y0_S2BEG[6] ,
    \Tile_X3Y0_S2BEG[5] ,
    \Tile_X3Y0_S2BEG[4] ,
    \Tile_X3Y0_S2BEG[3] ,
    \Tile_X3Y0_S2BEG[2] ,
    \Tile_X3Y0_S2BEG[1] ,
    \Tile_X3Y0_S2BEG[0] }),
    .S2BEGb({\Tile_X3Y0_S2BEGb[7] ,
    \Tile_X3Y0_S2BEGb[6] ,
    \Tile_X3Y0_S2BEGb[5] ,
    \Tile_X3Y0_S2BEGb[4] ,
    \Tile_X3Y0_S2BEGb[3] ,
    \Tile_X3Y0_S2BEGb[2] ,
    \Tile_X3Y0_S2BEGb[1] ,
    \Tile_X3Y0_S2BEGb[0] }),
    .S4BEG({\Tile_X3Y0_S4BEG[15] ,
    \Tile_X3Y0_S4BEG[14] ,
    \Tile_X3Y0_S4BEG[13] ,
    \Tile_X3Y0_S4BEG[12] ,
    \Tile_X3Y0_S4BEG[11] ,
    \Tile_X3Y0_S4BEG[10] ,
    \Tile_X3Y0_S4BEG[9] ,
    \Tile_X3Y0_S4BEG[8] ,
    \Tile_X3Y0_S4BEG[7] ,
    \Tile_X3Y0_S4BEG[6] ,
    \Tile_X3Y0_S4BEG[5] ,
    \Tile_X3Y0_S4BEG[4] ,
    \Tile_X3Y0_S4BEG[3] ,
    \Tile_X3Y0_S4BEG[2] ,
    \Tile_X3Y0_S4BEG[1] ,
    \Tile_X3Y0_S4BEG[0] }),
    .SS4BEG({\Tile_X3Y0_SS4BEG[15] ,
    \Tile_X3Y0_SS4BEG[14] ,
    \Tile_X3Y0_SS4BEG[13] ,
    \Tile_X3Y0_SS4BEG[12] ,
    \Tile_X3Y0_SS4BEG[11] ,
    \Tile_X3Y0_SS4BEG[10] ,
    \Tile_X3Y0_SS4BEG[9] ,
    \Tile_X3Y0_SS4BEG[8] ,
    \Tile_X3Y0_SS4BEG[7] ,
    \Tile_X3Y0_SS4BEG[6] ,
    \Tile_X3Y0_SS4BEG[5] ,
    \Tile_X3Y0_SS4BEG[4] ,
    \Tile_X3Y0_SS4BEG[3] ,
    \Tile_X3Y0_SS4BEG[2] ,
    \Tile_X3Y0_SS4BEG[1] ,
    \Tile_X3Y0_SS4BEG[0] }));
 LUT4AB Tile_X3Y10_LUT4AB (.Ci(Tile_X3Y11_Co),
    .Co(Tile_X3Y10_Co),
    .UserCLK(Tile_X3Y11_UserCLKo),
    .UserCLKo(Tile_X3Y10_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X3Y10_E1BEG[3] ,
    \Tile_X3Y10_E1BEG[2] ,
    \Tile_X3Y10_E1BEG[1] ,
    \Tile_X3Y10_E1BEG[0] }),
    .E1END({\Tile_X2Y10_E1BEG[3] ,
    \Tile_X2Y10_E1BEG[2] ,
    \Tile_X2Y10_E1BEG[1] ,
    \Tile_X2Y10_E1BEG[0] }),
    .E2BEG({\Tile_X3Y10_E2BEG[7] ,
    \Tile_X3Y10_E2BEG[6] ,
    \Tile_X3Y10_E2BEG[5] ,
    \Tile_X3Y10_E2BEG[4] ,
    \Tile_X3Y10_E2BEG[3] ,
    \Tile_X3Y10_E2BEG[2] ,
    \Tile_X3Y10_E2BEG[1] ,
    \Tile_X3Y10_E2BEG[0] }),
    .E2BEGb({\Tile_X3Y10_E2BEGb[7] ,
    \Tile_X3Y10_E2BEGb[6] ,
    \Tile_X3Y10_E2BEGb[5] ,
    \Tile_X3Y10_E2BEGb[4] ,
    \Tile_X3Y10_E2BEGb[3] ,
    \Tile_X3Y10_E2BEGb[2] ,
    \Tile_X3Y10_E2BEGb[1] ,
    \Tile_X3Y10_E2BEGb[0] }),
    .E2END({\Tile_X2Y10_E2BEGb[7] ,
    \Tile_X2Y10_E2BEGb[6] ,
    \Tile_X2Y10_E2BEGb[5] ,
    \Tile_X2Y10_E2BEGb[4] ,
    \Tile_X2Y10_E2BEGb[3] ,
    \Tile_X2Y10_E2BEGb[2] ,
    \Tile_X2Y10_E2BEGb[1] ,
    \Tile_X2Y10_E2BEGb[0] }),
    .E2MID({\Tile_X2Y10_E2BEG[7] ,
    \Tile_X2Y10_E2BEG[6] ,
    \Tile_X2Y10_E2BEG[5] ,
    \Tile_X2Y10_E2BEG[4] ,
    \Tile_X2Y10_E2BEG[3] ,
    \Tile_X2Y10_E2BEG[2] ,
    \Tile_X2Y10_E2BEG[1] ,
    \Tile_X2Y10_E2BEG[0] }),
    .E6BEG({\Tile_X3Y10_E6BEG[11] ,
    \Tile_X3Y10_E6BEG[10] ,
    \Tile_X3Y10_E6BEG[9] ,
    \Tile_X3Y10_E6BEG[8] ,
    \Tile_X3Y10_E6BEG[7] ,
    \Tile_X3Y10_E6BEG[6] ,
    \Tile_X3Y10_E6BEG[5] ,
    \Tile_X3Y10_E6BEG[4] ,
    \Tile_X3Y10_E6BEG[3] ,
    \Tile_X3Y10_E6BEG[2] ,
    \Tile_X3Y10_E6BEG[1] ,
    \Tile_X3Y10_E6BEG[0] }),
    .E6END({\Tile_X2Y10_E6BEG[11] ,
    \Tile_X2Y10_E6BEG[10] ,
    \Tile_X2Y10_E6BEG[9] ,
    \Tile_X2Y10_E6BEG[8] ,
    \Tile_X2Y10_E6BEG[7] ,
    \Tile_X2Y10_E6BEG[6] ,
    \Tile_X2Y10_E6BEG[5] ,
    \Tile_X2Y10_E6BEG[4] ,
    \Tile_X2Y10_E6BEG[3] ,
    \Tile_X2Y10_E6BEG[2] ,
    \Tile_X2Y10_E6BEG[1] ,
    \Tile_X2Y10_E6BEG[0] }),
    .EE4BEG({\Tile_X3Y10_EE4BEG[15] ,
    \Tile_X3Y10_EE4BEG[14] ,
    \Tile_X3Y10_EE4BEG[13] ,
    \Tile_X3Y10_EE4BEG[12] ,
    \Tile_X3Y10_EE4BEG[11] ,
    \Tile_X3Y10_EE4BEG[10] ,
    \Tile_X3Y10_EE4BEG[9] ,
    \Tile_X3Y10_EE4BEG[8] ,
    \Tile_X3Y10_EE4BEG[7] ,
    \Tile_X3Y10_EE4BEG[6] ,
    \Tile_X3Y10_EE4BEG[5] ,
    \Tile_X3Y10_EE4BEG[4] ,
    \Tile_X3Y10_EE4BEG[3] ,
    \Tile_X3Y10_EE4BEG[2] ,
    \Tile_X3Y10_EE4BEG[1] ,
    \Tile_X3Y10_EE4BEG[0] }),
    .EE4END({\Tile_X2Y10_EE4BEG[15] ,
    \Tile_X2Y10_EE4BEG[14] ,
    \Tile_X2Y10_EE4BEG[13] ,
    \Tile_X2Y10_EE4BEG[12] ,
    \Tile_X2Y10_EE4BEG[11] ,
    \Tile_X2Y10_EE4BEG[10] ,
    \Tile_X2Y10_EE4BEG[9] ,
    \Tile_X2Y10_EE4BEG[8] ,
    \Tile_X2Y10_EE4BEG[7] ,
    \Tile_X2Y10_EE4BEG[6] ,
    \Tile_X2Y10_EE4BEG[5] ,
    \Tile_X2Y10_EE4BEG[4] ,
    \Tile_X2Y10_EE4BEG[3] ,
    \Tile_X2Y10_EE4BEG[2] ,
    \Tile_X2Y10_EE4BEG[1] ,
    \Tile_X2Y10_EE4BEG[0] }),
    .FrameData({\Tile_X2Y10_FrameData_O[31] ,
    \Tile_X2Y10_FrameData_O[30] ,
    \Tile_X2Y10_FrameData_O[29] ,
    \Tile_X2Y10_FrameData_O[28] ,
    \Tile_X2Y10_FrameData_O[27] ,
    \Tile_X2Y10_FrameData_O[26] ,
    \Tile_X2Y10_FrameData_O[25] ,
    \Tile_X2Y10_FrameData_O[24] ,
    \Tile_X2Y10_FrameData_O[23] ,
    \Tile_X2Y10_FrameData_O[22] ,
    \Tile_X2Y10_FrameData_O[21] ,
    \Tile_X2Y10_FrameData_O[20] ,
    \Tile_X2Y10_FrameData_O[19] ,
    \Tile_X2Y10_FrameData_O[18] ,
    \Tile_X2Y10_FrameData_O[17] ,
    \Tile_X2Y10_FrameData_O[16] ,
    \Tile_X2Y10_FrameData_O[15] ,
    \Tile_X2Y10_FrameData_O[14] ,
    \Tile_X2Y10_FrameData_O[13] ,
    \Tile_X2Y10_FrameData_O[12] ,
    \Tile_X2Y10_FrameData_O[11] ,
    \Tile_X2Y10_FrameData_O[10] ,
    \Tile_X2Y10_FrameData_O[9] ,
    \Tile_X2Y10_FrameData_O[8] ,
    \Tile_X2Y10_FrameData_O[7] ,
    \Tile_X2Y10_FrameData_O[6] ,
    \Tile_X2Y10_FrameData_O[5] ,
    \Tile_X2Y10_FrameData_O[4] ,
    \Tile_X2Y10_FrameData_O[3] ,
    \Tile_X2Y10_FrameData_O[2] ,
    \Tile_X2Y10_FrameData_O[1] ,
    \Tile_X2Y10_FrameData_O[0] }),
    .FrameData_O({\Tile_X3Y10_FrameData_O[31] ,
    \Tile_X3Y10_FrameData_O[30] ,
    \Tile_X3Y10_FrameData_O[29] ,
    \Tile_X3Y10_FrameData_O[28] ,
    \Tile_X3Y10_FrameData_O[27] ,
    \Tile_X3Y10_FrameData_O[26] ,
    \Tile_X3Y10_FrameData_O[25] ,
    \Tile_X3Y10_FrameData_O[24] ,
    \Tile_X3Y10_FrameData_O[23] ,
    \Tile_X3Y10_FrameData_O[22] ,
    \Tile_X3Y10_FrameData_O[21] ,
    \Tile_X3Y10_FrameData_O[20] ,
    \Tile_X3Y10_FrameData_O[19] ,
    \Tile_X3Y10_FrameData_O[18] ,
    \Tile_X3Y10_FrameData_O[17] ,
    \Tile_X3Y10_FrameData_O[16] ,
    \Tile_X3Y10_FrameData_O[15] ,
    \Tile_X3Y10_FrameData_O[14] ,
    \Tile_X3Y10_FrameData_O[13] ,
    \Tile_X3Y10_FrameData_O[12] ,
    \Tile_X3Y10_FrameData_O[11] ,
    \Tile_X3Y10_FrameData_O[10] ,
    \Tile_X3Y10_FrameData_O[9] ,
    \Tile_X3Y10_FrameData_O[8] ,
    \Tile_X3Y10_FrameData_O[7] ,
    \Tile_X3Y10_FrameData_O[6] ,
    \Tile_X3Y10_FrameData_O[5] ,
    \Tile_X3Y10_FrameData_O[4] ,
    \Tile_X3Y10_FrameData_O[3] ,
    \Tile_X3Y10_FrameData_O[2] ,
    \Tile_X3Y10_FrameData_O[1] ,
    \Tile_X3Y10_FrameData_O[0] }),
    .FrameStrobe({\Tile_X3Y11_FrameStrobe_O[19] ,
    \Tile_X3Y11_FrameStrobe_O[18] ,
    \Tile_X3Y11_FrameStrobe_O[17] ,
    \Tile_X3Y11_FrameStrobe_O[16] ,
    \Tile_X3Y11_FrameStrobe_O[15] ,
    \Tile_X3Y11_FrameStrobe_O[14] ,
    \Tile_X3Y11_FrameStrobe_O[13] ,
    \Tile_X3Y11_FrameStrobe_O[12] ,
    \Tile_X3Y11_FrameStrobe_O[11] ,
    \Tile_X3Y11_FrameStrobe_O[10] ,
    \Tile_X3Y11_FrameStrobe_O[9] ,
    \Tile_X3Y11_FrameStrobe_O[8] ,
    \Tile_X3Y11_FrameStrobe_O[7] ,
    \Tile_X3Y11_FrameStrobe_O[6] ,
    \Tile_X3Y11_FrameStrobe_O[5] ,
    \Tile_X3Y11_FrameStrobe_O[4] ,
    \Tile_X3Y11_FrameStrobe_O[3] ,
    \Tile_X3Y11_FrameStrobe_O[2] ,
    \Tile_X3Y11_FrameStrobe_O[1] ,
    \Tile_X3Y11_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X3Y10_FrameStrobe_O[19] ,
    \Tile_X3Y10_FrameStrobe_O[18] ,
    \Tile_X3Y10_FrameStrobe_O[17] ,
    \Tile_X3Y10_FrameStrobe_O[16] ,
    \Tile_X3Y10_FrameStrobe_O[15] ,
    \Tile_X3Y10_FrameStrobe_O[14] ,
    \Tile_X3Y10_FrameStrobe_O[13] ,
    \Tile_X3Y10_FrameStrobe_O[12] ,
    \Tile_X3Y10_FrameStrobe_O[11] ,
    \Tile_X3Y10_FrameStrobe_O[10] ,
    \Tile_X3Y10_FrameStrobe_O[9] ,
    \Tile_X3Y10_FrameStrobe_O[8] ,
    \Tile_X3Y10_FrameStrobe_O[7] ,
    \Tile_X3Y10_FrameStrobe_O[6] ,
    \Tile_X3Y10_FrameStrobe_O[5] ,
    \Tile_X3Y10_FrameStrobe_O[4] ,
    \Tile_X3Y10_FrameStrobe_O[3] ,
    \Tile_X3Y10_FrameStrobe_O[2] ,
    \Tile_X3Y10_FrameStrobe_O[1] ,
    \Tile_X3Y10_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X3Y10_N1BEG[3] ,
    \Tile_X3Y10_N1BEG[2] ,
    \Tile_X3Y10_N1BEG[1] ,
    \Tile_X3Y10_N1BEG[0] }),
    .N1END({\Tile_X3Y11_N1BEG[3] ,
    \Tile_X3Y11_N1BEG[2] ,
    \Tile_X3Y11_N1BEG[1] ,
    \Tile_X3Y11_N1BEG[0] }),
    .N2BEG({\Tile_X3Y10_N2BEG[7] ,
    \Tile_X3Y10_N2BEG[6] ,
    \Tile_X3Y10_N2BEG[5] ,
    \Tile_X3Y10_N2BEG[4] ,
    \Tile_X3Y10_N2BEG[3] ,
    \Tile_X3Y10_N2BEG[2] ,
    \Tile_X3Y10_N2BEG[1] ,
    \Tile_X3Y10_N2BEG[0] }),
    .N2BEGb({\Tile_X3Y10_N2BEGb[7] ,
    \Tile_X3Y10_N2BEGb[6] ,
    \Tile_X3Y10_N2BEGb[5] ,
    \Tile_X3Y10_N2BEGb[4] ,
    \Tile_X3Y10_N2BEGb[3] ,
    \Tile_X3Y10_N2BEGb[2] ,
    \Tile_X3Y10_N2BEGb[1] ,
    \Tile_X3Y10_N2BEGb[0] }),
    .N2END({\Tile_X3Y11_N2BEGb[7] ,
    \Tile_X3Y11_N2BEGb[6] ,
    \Tile_X3Y11_N2BEGb[5] ,
    \Tile_X3Y11_N2BEGb[4] ,
    \Tile_X3Y11_N2BEGb[3] ,
    \Tile_X3Y11_N2BEGb[2] ,
    \Tile_X3Y11_N2BEGb[1] ,
    \Tile_X3Y11_N2BEGb[0] }),
    .N2MID({\Tile_X3Y11_N2BEG[7] ,
    \Tile_X3Y11_N2BEG[6] ,
    \Tile_X3Y11_N2BEG[5] ,
    \Tile_X3Y11_N2BEG[4] ,
    \Tile_X3Y11_N2BEG[3] ,
    \Tile_X3Y11_N2BEG[2] ,
    \Tile_X3Y11_N2BEG[1] ,
    \Tile_X3Y11_N2BEG[0] }),
    .N4BEG({\Tile_X3Y10_N4BEG[15] ,
    \Tile_X3Y10_N4BEG[14] ,
    \Tile_X3Y10_N4BEG[13] ,
    \Tile_X3Y10_N4BEG[12] ,
    \Tile_X3Y10_N4BEG[11] ,
    \Tile_X3Y10_N4BEG[10] ,
    \Tile_X3Y10_N4BEG[9] ,
    \Tile_X3Y10_N4BEG[8] ,
    \Tile_X3Y10_N4BEG[7] ,
    \Tile_X3Y10_N4BEG[6] ,
    \Tile_X3Y10_N4BEG[5] ,
    \Tile_X3Y10_N4BEG[4] ,
    \Tile_X3Y10_N4BEG[3] ,
    \Tile_X3Y10_N4BEG[2] ,
    \Tile_X3Y10_N4BEG[1] ,
    \Tile_X3Y10_N4BEG[0] }),
    .N4END({\Tile_X3Y11_N4BEG[15] ,
    \Tile_X3Y11_N4BEG[14] ,
    \Tile_X3Y11_N4BEG[13] ,
    \Tile_X3Y11_N4BEG[12] ,
    \Tile_X3Y11_N4BEG[11] ,
    \Tile_X3Y11_N4BEG[10] ,
    \Tile_X3Y11_N4BEG[9] ,
    \Tile_X3Y11_N4BEG[8] ,
    \Tile_X3Y11_N4BEG[7] ,
    \Tile_X3Y11_N4BEG[6] ,
    \Tile_X3Y11_N4BEG[5] ,
    \Tile_X3Y11_N4BEG[4] ,
    \Tile_X3Y11_N4BEG[3] ,
    \Tile_X3Y11_N4BEG[2] ,
    \Tile_X3Y11_N4BEG[1] ,
    \Tile_X3Y11_N4BEG[0] }),
    .NN4BEG({\Tile_X3Y10_NN4BEG[15] ,
    \Tile_X3Y10_NN4BEG[14] ,
    \Tile_X3Y10_NN4BEG[13] ,
    \Tile_X3Y10_NN4BEG[12] ,
    \Tile_X3Y10_NN4BEG[11] ,
    \Tile_X3Y10_NN4BEG[10] ,
    \Tile_X3Y10_NN4BEG[9] ,
    \Tile_X3Y10_NN4BEG[8] ,
    \Tile_X3Y10_NN4BEG[7] ,
    \Tile_X3Y10_NN4BEG[6] ,
    \Tile_X3Y10_NN4BEG[5] ,
    \Tile_X3Y10_NN4BEG[4] ,
    \Tile_X3Y10_NN4BEG[3] ,
    \Tile_X3Y10_NN4BEG[2] ,
    \Tile_X3Y10_NN4BEG[1] ,
    \Tile_X3Y10_NN4BEG[0] }),
    .NN4END({\Tile_X3Y11_NN4BEG[15] ,
    \Tile_X3Y11_NN4BEG[14] ,
    \Tile_X3Y11_NN4BEG[13] ,
    \Tile_X3Y11_NN4BEG[12] ,
    \Tile_X3Y11_NN4BEG[11] ,
    \Tile_X3Y11_NN4BEG[10] ,
    \Tile_X3Y11_NN4BEG[9] ,
    \Tile_X3Y11_NN4BEG[8] ,
    \Tile_X3Y11_NN4BEG[7] ,
    \Tile_X3Y11_NN4BEG[6] ,
    \Tile_X3Y11_NN4BEG[5] ,
    \Tile_X3Y11_NN4BEG[4] ,
    \Tile_X3Y11_NN4BEG[3] ,
    \Tile_X3Y11_NN4BEG[2] ,
    \Tile_X3Y11_NN4BEG[1] ,
    \Tile_X3Y11_NN4BEG[0] }),
    .S1BEG({\Tile_X3Y10_S1BEG[3] ,
    \Tile_X3Y10_S1BEG[2] ,
    \Tile_X3Y10_S1BEG[1] ,
    \Tile_X3Y10_S1BEG[0] }),
    .S1END({\Tile_X3Y9_S1BEG[3] ,
    \Tile_X3Y9_S1BEG[2] ,
    \Tile_X3Y9_S1BEG[1] ,
    \Tile_X3Y9_S1BEG[0] }),
    .S2BEG({\Tile_X3Y10_S2BEG[7] ,
    \Tile_X3Y10_S2BEG[6] ,
    \Tile_X3Y10_S2BEG[5] ,
    \Tile_X3Y10_S2BEG[4] ,
    \Tile_X3Y10_S2BEG[3] ,
    \Tile_X3Y10_S2BEG[2] ,
    \Tile_X3Y10_S2BEG[1] ,
    \Tile_X3Y10_S2BEG[0] }),
    .S2BEGb({\Tile_X3Y10_S2BEGb[7] ,
    \Tile_X3Y10_S2BEGb[6] ,
    \Tile_X3Y10_S2BEGb[5] ,
    \Tile_X3Y10_S2BEGb[4] ,
    \Tile_X3Y10_S2BEGb[3] ,
    \Tile_X3Y10_S2BEGb[2] ,
    \Tile_X3Y10_S2BEGb[1] ,
    \Tile_X3Y10_S2BEGb[0] }),
    .S2END({\Tile_X3Y9_S2BEGb[7] ,
    \Tile_X3Y9_S2BEGb[6] ,
    \Tile_X3Y9_S2BEGb[5] ,
    \Tile_X3Y9_S2BEGb[4] ,
    \Tile_X3Y9_S2BEGb[3] ,
    \Tile_X3Y9_S2BEGb[2] ,
    \Tile_X3Y9_S2BEGb[1] ,
    \Tile_X3Y9_S2BEGb[0] }),
    .S2MID({\Tile_X3Y9_S2BEG[7] ,
    \Tile_X3Y9_S2BEG[6] ,
    \Tile_X3Y9_S2BEG[5] ,
    \Tile_X3Y9_S2BEG[4] ,
    \Tile_X3Y9_S2BEG[3] ,
    \Tile_X3Y9_S2BEG[2] ,
    \Tile_X3Y9_S2BEG[1] ,
    \Tile_X3Y9_S2BEG[0] }),
    .S4BEG({\Tile_X3Y10_S4BEG[15] ,
    \Tile_X3Y10_S4BEG[14] ,
    \Tile_X3Y10_S4BEG[13] ,
    \Tile_X3Y10_S4BEG[12] ,
    \Tile_X3Y10_S4BEG[11] ,
    \Tile_X3Y10_S4BEG[10] ,
    \Tile_X3Y10_S4BEG[9] ,
    \Tile_X3Y10_S4BEG[8] ,
    \Tile_X3Y10_S4BEG[7] ,
    \Tile_X3Y10_S4BEG[6] ,
    \Tile_X3Y10_S4BEG[5] ,
    \Tile_X3Y10_S4BEG[4] ,
    \Tile_X3Y10_S4BEG[3] ,
    \Tile_X3Y10_S4BEG[2] ,
    \Tile_X3Y10_S4BEG[1] ,
    \Tile_X3Y10_S4BEG[0] }),
    .S4END({\Tile_X3Y9_S4BEG[15] ,
    \Tile_X3Y9_S4BEG[14] ,
    \Tile_X3Y9_S4BEG[13] ,
    \Tile_X3Y9_S4BEG[12] ,
    \Tile_X3Y9_S4BEG[11] ,
    \Tile_X3Y9_S4BEG[10] ,
    \Tile_X3Y9_S4BEG[9] ,
    \Tile_X3Y9_S4BEG[8] ,
    \Tile_X3Y9_S4BEG[7] ,
    \Tile_X3Y9_S4BEG[6] ,
    \Tile_X3Y9_S4BEG[5] ,
    \Tile_X3Y9_S4BEG[4] ,
    \Tile_X3Y9_S4BEG[3] ,
    \Tile_X3Y9_S4BEG[2] ,
    \Tile_X3Y9_S4BEG[1] ,
    \Tile_X3Y9_S4BEG[0] }),
    .SS4BEG({\Tile_X3Y10_SS4BEG[15] ,
    \Tile_X3Y10_SS4BEG[14] ,
    \Tile_X3Y10_SS4BEG[13] ,
    \Tile_X3Y10_SS4BEG[12] ,
    \Tile_X3Y10_SS4BEG[11] ,
    \Tile_X3Y10_SS4BEG[10] ,
    \Tile_X3Y10_SS4BEG[9] ,
    \Tile_X3Y10_SS4BEG[8] ,
    \Tile_X3Y10_SS4BEG[7] ,
    \Tile_X3Y10_SS4BEG[6] ,
    \Tile_X3Y10_SS4BEG[5] ,
    \Tile_X3Y10_SS4BEG[4] ,
    \Tile_X3Y10_SS4BEG[3] ,
    \Tile_X3Y10_SS4BEG[2] ,
    \Tile_X3Y10_SS4BEG[1] ,
    \Tile_X3Y10_SS4BEG[0] }),
    .SS4END({\Tile_X3Y9_SS4BEG[15] ,
    \Tile_X3Y9_SS4BEG[14] ,
    \Tile_X3Y9_SS4BEG[13] ,
    \Tile_X3Y9_SS4BEG[12] ,
    \Tile_X3Y9_SS4BEG[11] ,
    \Tile_X3Y9_SS4BEG[10] ,
    \Tile_X3Y9_SS4BEG[9] ,
    \Tile_X3Y9_SS4BEG[8] ,
    \Tile_X3Y9_SS4BEG[7] ,
    \Tile_X3Y9_SS4BEG[6] ,
    \Tile_X3Y9_SS4BEG[5] ,
    \Tile_X3Y9_SS4BEG[4] ,
    \Tile_X3Y9_SS4BEG[3] ,
    \Tile_X3Y9_SS4BEG[2] ,
    \Tile_X3Y9_SS4BEG[1] ,
    \Tile_X3Y9_SS4BEG[0] }),
    .W1BEG({\Tile_X3Y10_W1BEG[3] ,
    \Tile_X3Y10_W1BEG[2] ,
    \Tile_X3Y10_W1BEG[1] ,
    \Tile_X3Y10_W1BEG[0] }),
    .W1END({\Tile_X4Y10_W1BEG[3] ,
    \Tile_X4Y10_W1BEG[2] ,
    \Tile_X4Y10_W1BEG[1] ,
    \Tile_X4Y10_W1BEG[0] }),
    .W2BEG({\Tile_X3Y10_W2BEG[7] ,
    \Tile_X3Y10_W2BEG[6] ,
    \Tile_X3Y10_W2BEG[5] ,
    \Tile_X3Y10_W2BEG[4] ,
    \Tile_X3Y10_W2BEG[3] ,
    \Tile_X3Y10_W2BEG[2] ,
    \Tile_X3Y10_W2BEG[1] ,
    \Tile_X3Y10_W2BEG[0] }),
    .W2BEGb({\Tile_X3Y10_W2BEGb[7] ,
    \Tile_X3Y10_W2BEGb[6] ,
    \Tile_X3Y10_W2BEGb[5] ,
    \Tile_X3Y10_W2BEGb[4] ,
    \Tile_X3Y10_W2BEGb[3] ,
    \Tile_X3Y10_W2BEGb[2] ,
    \Tile_X3Y10_W2BEGb[1] ,
    \Tile_X3Y10_W2BEGb[0] }),
    .W2END({\Tile_X4Y10_W2BEGb[7] ,
    \Tile_X4Y10_W2BEGb[6] ,
    \Tile_X4Y10_W2BEGb[5] ,
    \Tile_X4Y10_W2BEGb[4] ,
    \Tile_X4Y10_W2BEGb[3] ,
    \Tile_X4Y10_W2BEGb[2] ,
    \Tile_X4Y10_W2BEGb[1] ,
    \Tile_X4Y10_W2BEGb[0] }),
    .W2MID({\Tile_X4Y10_W2BEG[7] ,
    \Tile_X4Y10_W2BEG[6] ,
    \Tile_X4Y10_W2BEG[5] ,
    \Tile_X4Y10_W2BEG[4] ,
    \Tile_X4Y10_W2BEG[3] ,
    \Tile_X4Y10_W2BEG[2] ,
    \Tile_X4Y10_W2BEG[1] ,
    \Tile_X4Y10_W2BEG[0] }),
    .W6BEG({\Tile_X3Y10_W6BEG[11] ,
    \Tile_X3Y10_W6BEG[10] ,
    \Tile_X3Y10_W6BEG[9] ,
    \Tile_X3Y10_W6BEG[8] ,
    \Tile_X3Y10_W6BEG[7] ,
    \Tile_X3Y10_W6BEG[6] ,
    \Tile_X3Y10_W6BEG[5] ,
    \Tile_X3Y10_W6BEG[4] ,
    \Tile_X3Y10_W6BEG[3] ,
    \Tile_X3Y10_W6BEG[2] ,
    \Tile_X3Y10_W6BEG[1] ,
    \Tile_X3Y10_W6BEG[0] }),
    .W6END({\Tile_X4Y10_W6BEG[11] ,
    \Tile_X4Y10_W6BEG[10] ,
    \Tile_X4Y10_W6BEG[9] ,
    \Tile_X4Y10_W6BEG[8] ,
    \Tile_X4Y10_W6BEG[7] ,
    \Tile_X4Y10_W6BEG[6] ,
    \Tile_X4Y10_W6BEG[5] ,
    \Tile_X4Y10_W6BEG[4] ,
    \Tile_X4Y10_W6BEG[3] ,
    \Tile_X4Y10_W6BEG[2] ,
    \Tile_X4Y10_W6BEG[1] ,
    \Tile_X4Y10_W6BEG[0] }),
    .WW4BEG({\Tile_X3Y10_WW4BEG[15] ,
    \Tile_X3Y10_WW4BEG[14] ,
    \Tile_X3Y10_WW4BEG[13] ,
    \Tile_X3Y10_WW4BEG[12] ,
    \Tile_X3Y10_WW4BEG[11] ,
    \Tile_X3Y10_WW4BEG[10] ,
    \Tile_X3Y10_WW4BEG[9] ,
    \Tile_X3Y10_WW4BEG[8] ,
    \Tile_X3Y10_WW4BEG[7] ,
    \Tile_X3Y10_WW4BEG[6] ,
    \Tile_X3Y10_WW4BEG[5] ,
    \Tile_X3Y10_WW4BEG[4] ,
    \Tile_X3Y10_WW4BEG[3] ,
    \Tile_X3Y10_WW4BEG[2] ,
    \Tile_X3Y10_WW4BEG[1] ,
    \Tile_X3Y10_WW4BEG[0] }),
    .WW4END({\Tile_X4Y10_WW4BEG[15] ,
    \Tile_X4Y10_WW4BEG[14] ,
    \Tile_X4Y10_WW4BEG[13] ,
    \Tile_X4Y10_WW4BEG[12] ,
    \Tile_X4Y10_WW4BEG[11] ,
    \Tile_X4Y10_WW4BEG[10] ,
    \Tile_X4Y10_WW4BEG[9] ,
    \Tile_X4Y10_WW4BEG[8] ,
    \Tile_X4Y10_WW4BEG[7] ,
    \Tile_X4Y10_WW4BEG[6] ,
    \Tile_X4Y10_WW4BEG[5] ,
    \Tile_X4Y10_WW4BEG[4] ,
    \Tile_X4Y10_WW4BEG[3] ,
    \Tile_X4Y10_WW4BEG[2] ,
    \Tile_X4Y10_WW4BEG[1] ,
    \Tile_X4Y10_WW4BEG[0] }));
 LUT4AB Tile_X3Y11_LUT4AB (.Ci(Tile_X3Y12_Co),
    .Co(Tile_X3Y11_Co),
    .UserCLK(Tile_X3Y12_UserCLKo),
    .UserCLKo(Tile_X3Y11_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X3Y11_E1BEG[3] ,
    \Tile_X3Y11_E1BEG[2] ,
    \Tile_X3Y11_E1BEG[1] ,
    \Tile_X3Y11_E1BEG[0] }),
    .E1END({\Tile_X2Y11_E1BEG[3] ,
    \Tile_X2Y11_E1BEG[2] ,
    \Tile_X2Y11_E1BEG[1] ,
    \Tile_X2Y11_E1BEG[0] }),
    .E2BEG({\Tile_X3Y11_E2BEG[7] ,
    \Tile_X3Y11_E2BEG[6] ,
    \Tile_X3Y11_E2BEG[5] ,
    \Tile_X3Y11_E2BEG[4] ,
    \Tile_X3Y11_E2BEG[3] ,
    \Tile_X3Y11_E2BEG[2] ,
    \Tile_X3Y11_E2BEG[1] ,
    \Tile_X3Y11_E2BEG[0] }),
    .E2BEGb({\Tile_X3Y11_E2BEGb[7] ,
    \Tile_X3Y11_E2BEGb[6] ,
    \Tile_X3Y11_E2BEGb[5] ,
    \Tile_X3Y11_E2BEGb[4] ,
    \Tile_X3Y11_E2BEGb[3] ,
    \Tile_X3Y11_E2BEGb[2] ,
    \Tile_X3Y11_E2BEGb[1] ,
    \Tile_X3Y11_E2BEGb[0] }),
    .E2END({\Tile_X2Y11_E2BEGb[7] ,
    \Tile_X2Y11_E2BEGb[6] ,
    \Tile_X2Y11_E2BEGb[5] ,
    \Tile_X2Y11_E2BEGb[4] ,
    \Tile_X2Y11_E2BEGb[3] ,
    \Tile_X2Y11_E2BEGb[2] ,
    \Tile_X2Y11_E2BEGb[1] ,
    \Tile_X2Y11_E2BEGb[0] }),
    .E2MID({\Tile_X2Y11_E2BEG[7] ,
    \Tile_X2Y11_E2BEG[6] ,
    \Tile_X2Y11_E2BEG[5] ,
    \Tile_X2Y11_E2BEG[4] ,
    \Tile_X2Y11_E2BEG[3] ,
    \Tile_X2Y11_E2BEG[2] ,
    \Tile_X2Y11_E2BEG[1] ,
    \Tile_X2Y11_E2BEG[0] }),
    .E6BEG({\Tile_X3Y11_E6BEG[11] ,
    \Tile_X3Y11_E6BEG[10] ,
    \Tile_X3Y11_E6BEG[9] ,
    \Tile_X3Y11_E6BEG[8] ,
    \Tile_X3Y11_E6BEG[7] ,
    \Tile_X3Y11_E6BEG[6] ,
    \Tile_X3Y11_E6BEG[5] ,
    \Tile_X3Y11_E6BEG[4] ,
    \Tile_X3Y11_E6BEG[3] ,
    \Tile_X3Y11_E6BEG[2] ,
    \Tile_X3Y11_E6BEG[1] ,
    \Tile_X3Y11_E6BEG[0] }),
    .E6END({\Tile_X2Y11_E6BEG[11] ,
    \Tile_X2Y11_E6BEG[10] ,
    \Tile_X2Y11_E6BEG[9] ,
    \Tile_X2Y11_E6BEG[8] ,
    \Tile_X2Y11_E6BEG[7] ,
    \Tile_X2Y11_E6BEG[6] ,
    \Tile_X2Y11_E6BEG[5] ,
    \Tile_X2Y11_E6BEG[4] ,
    \Tile_X2Y11_E6BEG[3] ,
    \Tile_X2Y11_E6BEG[2] ,
    \Tile_X2Y11_E6BEG[1] ,
    \Tile_X2Y11_E6BEG[0] }),
    .EE4BEG({\Tile_X3Y11_EE4BEG[15] ,
    \Tile_X3Y11_EE4BEG[14] ,
    \Tile_X3Y11_EE4BEG[13] ,
    \Tile_X3Y11_EE4BEG[12] ,
    \Tile_X3Y11_EE4BEG[11] ,
    \Tile_X3Y11_EE4BEG[10] ,
    \Tile_X3Y11_EE4BEG[9] ,
    \Tile_X3Y11_EE4BEG[8] ,
    \Tile_X3Y11_EE4BEG[7] ,
    \Tile_X3Y11_EE4BEG[6] ,
    \Tile_X3Y11_EE4BEG[5] ,
    \Tile_X3Y11_EE4BEG[4] ,
    \Tile_X3Y11_EE4BEG[3] ,
    \Tile_X3Y11_EE4BEG[2] ,
    \Tile_X3Y11_EE4BEG[1] ,
    \Tile_X3Y11_EE4BEG[0] }),
    .EE4END({\Tile_X2Y11_EE4BEG[15] ,
    \Tile_X2Y11_EE4BEG[14] ,
    \Tile_X2Y11_EE4BEG[13] ,
    \Tile_X2Y11_EE4BEG[12] ,
    \Tile_X2Y11_EE4BEG[11] ,
    \Tile_X2Y11_EE4BEG[10] ,
    \Tile_X2Y11_EE4BEG[9] ,
    \Tile_X2Y11_EE4BEG[8] ,
    \Tile_X2Y11_EE4BEG[7] ,
    \Tile_X2Y11_EE4BEG[6] ,
    \Tile_X2Y11_EE4BEG[5] ,
    \Tile_X2Y11_EE4BEG[4] ,
    \Tile_X2Y11_EE4BEG[3] ,
    \Tile_X2Y11_EE4BEG[2] ,
    \Tile_X2Y11_EE4BEG[1] ,
    \Tile_X2Y11_EE4BEG[0] }),
    .FrameData({\Tile_X2Y11_FrameData_O[31] ,
    \Tile_X2Y11_FrameData_O[30] ,
    \Tile_X2Y11_FrameData_O[29] ,
    \Tile_X2Y11_FrameData_O[28] ,
    \Tile_X2Y11_FrameData_O[27] ,
    \Tile_X2Y11_FrameData_O[26] ,
    \Tile_X2Y11_FrameData_O[25] ,
    \Tile_X2Y11_FrameData_O[24] ,
    \Tile_X2Y11_FrameData_O[23] ,
    \Tile_X2Y11_FrameData_O[22] ,
    \Tile_X2Y11_FrameData_O[21] ,
    \Tile_X2Y11_FrameData_O[20] ,
    \Tile_X2Y11_FrameData_O[19] ,
    \Tile_X2Y11_FrameData_O[18] ,
    \Tile_X2Y11_FrameData_O[17] ,
    \Tile_X2Y11_FrameData_O[16] ,
    \Tile_X2Y11_FrameData_O[15] ,
    \Tile_X2Y11_FrameData_O[14] ,
    \Tile_X2Y11_FrameData_O[13] ,
    \Tile_X2Y11_FrameData_O[12] ,
    \Tile_X2Y11_FrameData_O[11] ,
    \Tile_X2Y11_FrameData_O[10] ,
    \Tile_X2Y11_FrameData_O[9] ,
    \Tile_X2Y11_FrameData_O[8] ,
    \Tile_X2Y11_FrameData_O[7] ,
    \Tile_X2Y11_FrameData_O[6] ,
    \Tile_X2Y11_FrameData_O[5] ,
    \Tile_X2Y11_FrameData_O[4] ,
    \Tile_X2Y11_FrameData_O[3] ,
    \Tile_X2Y11_FrameData_O[2] ,
    \Tile_X2Y11_FrameData_O[1] ,
    \Tile_X2Y11_FrameData_O[0] }),
    .FrameData_O({\Tile_X3Y11_FrameData_O[31] ,
    \Tile_X3Y11_FrameData_O[30] ,
    \Tile_X3Y11_FrameData_O[29] ,
    \Tile_X3Y11_FrameData_O[28] ,
    \Tile_X3Y11_FrameData_O[27] ,
    \Tile_X3Y11_FrameData_O[26] ,
    \Tile_X3Y11_FrameData_O[25] ,
    \Tile_X3Y11_FrameData_O[24] ,
    \Tile_X3Y11_FrameData_O[23] ,
    \Tile_X3Y11_FrameData_O[22] ,
    \Tile_X3Y11_FrameData_O[21] ,
    \Tile_X3Y11_FrameData_O[20] ,
    \Tile_X3Y11_FrameData_O[19] ,
    \Tile_X3Y11_FrameData_O[18] ,
    \Tile_X3Y11_FrameData_O[17] ,
    \Tile_X3Y11_FrameData_O[16] ,
    \Tile_X3Y11_FrameData_O[15] ,
    \Tile_X3Y11_FrameData_O[14] ,
    \Tile_X3Y11_FrameData_O[13] ,
    \Tile_X3Y11_FrameData_O[12] ,
    \Tile_X3Y11_FrameData_O[11] ,
    \Tile_X3Y11_FrameData_O[10] ,
    \Tile_X3Y11_FrameData_O[9] ,
    \Tile_X3Y11_FrameData_O[8] ,
    \Tile_X3Y11_FrameData_O[7] ,
    \Tile_X3Y11_FrameData_O[6] ,
    \Tile_X3Y11_FrameData_O[5] ,
    \Tile_X3Y11_FrameData_O[4] ,
    \Tile_X3Y11_FrameData_O[3] ,
    \Tile_X3Y11_FrameData_O[2] ,
    \Tile_X3Y11_FrameData_O[1] ,
    \Tile_X3Y11_FrameData_O[0] }),
    .FrameStrobe({\Tile_X3Y12_FrameStrobe_O[19] ,
    \Tile_X3Y12_FrameStrobe_O[18] ,
    \Tile_X3Y12_FrameStrobe_O[17] ,
    \Tile_X3Y12_FrameStrobe_O[16] ,
    \Tile_X3Y12_FrameStrobe_O[15] ,
    \Tile_X3Y12_FrameStrobe_O[14] ,
    \Tile_X3Y12_FrameStrobe_O[13] ,
    \Tile_X3Y12_FrameStrobe_O[12] ,
    \Tile_X3Y12_FrameStrobe_O[11] ,
    \Tile_X3Y12_FrameStrobe_O[10] ,
    \Tile_X3Y12_FrameStrobe_O[9] ,
    \Tile_X3Y12_FrameStrobe_O[8] ,
    \Tile_X3Y12_FrameStrobe_O[7] ,
    \Tile_X3Y12_FrameStrobe_O[6] ,
    \Tile_X3Y12_FrameStrobe_O[5] ,
    \Tile_X3Y12_FrameStrobe_O[4] ,
    \Tile_X3Y12_FrameStrobe_O[3] ,
    \Tile_X3Y12_FrameStrobe_O[2] ,
    \Tile_X3Y12_FrameStrobe_O[1] ,
    \Tile_X3Y12_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X3Y11_FrameStrobe_O[19] ,
    \Tile_X3Y11_FrameStrobe_O[18] ,
    \Tile_X3Y11_FrameStrobe_O[17] ,
    \Tile_X3Y11_FrameStrobe_O[16] ,
    \Tile_X3Y11_FrameStrobe_O[15] ,
    \Tile_X3Y11_FrameStrobe_O[14] ,
    \Tile_X3Y11_FrameStrobe_O[13] ,
    \Tile_X3Y11_FrameStrobe_O[12] ,
    \Tile_X3Y11_FrameStrobe_O[11] ,
    \Tile_X3Y11_FrameStrobe_O[10] ,
    \Tile_X3Y11_FrameStrobe_O[9] ,
    \Tile_X3Y11_FrameStrobe_O[8] ,
    \Tile_X3Y11_FrameStrobe_O[7] ,
    \Tile_X3Y11_FrameStrobe_O[6] ,
    \Tile_X3Y11_FrameStrobe_O[5] ,
    \Tile_X3Y11_FrameStrobe_O[4] ,
    \Tile_X3Y11_FrameStrobe_O[3] ,
    \Tile_X3Y11_FrameStrobe_O[2] ,
    \Tile_X3Y11_FrameStrobe_O[1] ,
    \Tile_X3Y11_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X3Y11_N1BEG[3] ,
    \Tile_X3Y11_N1BEG[2] ,
    \Tile_X3Y11_N1BEG[1] ,
    \Tile_X3Y11_N1BEG[0] }),
    .N1END({\Tile_X3Y12_N1BEG[3] ,
    \Tile_X3Y12_N1BEG[2] ,
    \Tile_X3Y12_N1BEG[1] ,
    \Tile_X3Y12_N1BEG[0] }),
    .N2BEG({\Tile_X3Y11_N2BEG[7] ,
    \Tile_X3Y11_N2BEG[6] ,
    \Tile_X3Y11_N2BEG[5] ,
    \Tile_X3Y11_N2BEG[4] ,
    \Tile_X3Y11_N2BEG[3] ,
    \Tile_X3Y11_N2BEG[2] ,
    \Tile_X3Y11_N2BEG[1] ,
    \Tile_X3Y11_N2BEG[0] }),
    .N2BEGb({\Tile_X3Y11_N2BEGb[7] ,
    \Tile_X3Y11_N2BEGb[6] ,
    \Tile_X3Y11_N2BEGb[5] ,
    \Tile_X3Y11_N2BEGb[4] ,
    \Tile_X3Y11_N2BEGb[3] ,
    \Tile_X3Y11_N2BEGb[2] ,
    \Tile_X3Y11_N2BEGb[1] ,
    \Tile_X3Y11_N2BEGb[0] }),
    .N2END({\Tile_X3Y12_N2BEGb[7] ,
    \Tile_X3Y12_N2BEGb[6] ,
    \Tile_X3Y12_N2BEGb[5] ,
    \Tile_X3Y12_N2BEGb[4] ,
    \Tile_X3Y12_N2BEGb[3] ,
    \Tile_X3Y12_N2BEGb[2] ,
    \Tile_X3Y12_N2BEGb[1] ,
    \Tile_X3Y12_N2BEGb[0] }),
    .N2MID({\Tile_X3Y12_N2BEG[7] ,
    \Tile_X3Y12_N2BEG[6] ,
    \Tile_X3Y12_N2BEG[5] ,
    \Tile_X3Y12_N2BEG[4] ,
    \Tile_X3Y12_N2BEG[3] ,
    \Tile_X3Y12_N2BEG[2] ,
    \Tile_X3Y12_N2BEG[1] ,
    \Tile_X3Y12_N2BEG[0] }),
    .N4BEG({\Tile_X3Y11_N4BEG[15] ,
    \Tile_X3Y11_N4BEG[14] ,
    \Tile_X3Y11_N4BEG[13] ,
    \Tile_X3Y11_N4BEG[12] ,
    \Tile_X3Y11_N4BEG[11] ,
    \Tile_X3Y11_N4BEG[10] ,
    \Tile_X3Y11_N4BEG[9] ,
    \Tile_X3Y11_N4BEG[8] ,
    \Tile_X3Y11_N4BEG[7] ,
    \Tile_X3Y11_N4BEG[6] ,
    \Tile_X3Y11_N4BEG[5] ,
    \Tile_X3Y11_N4BEG[4] ,
    \Tile_X3Y11_N4BEG[3] ,
    \Tile_X3Y11_N4BEG[2] ,
    \Tile_X3Y11_N4BEG[1] ,
    \Tile_X3Y11_N4BEG[0] }),
    .N4END({\Tile_X3Y12_N4BEG[15] ,
    \Tile_X3Y12_N4BEG[14] ,
    \Tile_X3Y12_N4BEG[13] ,
    \Tile_X3Y12_N4BEG[12] ,
    \Tile_X3Y12_N4BEG[11] ,
    \Tile_X3Y12_N4BEG[10] ,
    \Tile_X3Y12_N4BEG[9] ,
    \Tile_X3Y12_N4BEG[8] ,
    \Tile_X3Y12_N4BEG[7] ,
    \Tile_X3Y12_N4BEG[6] ,
    \Tile_X3Y12_N4BEG[5] ,
    \Tile_X3Y12_N4BEG[4] ,
    \Tile_X3Y12_N4BEG[3] ,
    \Tile_X3Y12_N4BEG[2] ,
    \Tile_X3Y12_N4BEG[1] ,
    \Tile_X3Y12_N4BEG[0] }),
    .NN4BEG({\Tile_X3Y11_NN4BEG[15] ,
    \Tile_X3Y11_NN4BEG[14] ,
    \Tile_X3Y11_NN4BEG[13] ,
    \Tile_X3Y11_NN4BEG[12] ,
    \Tile_X3Y11_NN4BEG[11] ,
    \Tile_X3Y11_NN4BEG[10] ,
    \Tile_X3Y11_NN4BEG[9] ,
    \Tile_X3Y11_NN4BEG[8] ,
    \Tile_X3Y11_NN4BEG[7] ,
    \Tile_X3Y11_NN4BEG[6] ,
    \Tile_X3Y11_NN4BEG[5] ,
    \Tile_X3Y11_NN4BEG[4] ,
    \Tile_X3Y11_NN4BEG[3] ,
    \Tile_X3Y11_NN4BEG[2] ,
    \Tile_X3Y11_NN4BEG[1] ,
    \Tile_X3Y11_NN4BEG[0] }),
    .NN4END({\Tile_X3Y12_NN4BEG[15] ,
    \Tile_X3Y12_NN4BEG[14] ,
    \Tile_X3Y12_NN4BEG[13] ,
    \Tile_X3Y12_NN4BEG[12] ,
    \Tile_X3Y12_NN4BEG[11] ,
    \Tile_X3Y12_NN4BEG[10] ,
    \Tile_X3Y12_NN4BEG[9] ,
    \Tile_X3Y12_NN4BEG[8] ,
    \Tile_X3Y12_NN4BEG[7] ,
    \Tile_X3Y12_NN4BEG[6] ,
    \Tile_X3Y12_NN4BEG[5] ,
    \Tile_X3Y12_NN4BEG[4] ,
    \Tile_X3Y12_NN4BEG[3] ,
    \Tile_X3Y12_NN4BEG[2] ,
    \Tile_X3Y12_NN4BEG[1] ,
    \Tile_X3Y12_NN4BEG[0] }),
    .S1BEG({\Tile_X3Y11_S1BEG[3] ,
    \Tile_X3Y11_S1BEG[2] ,
    \Tile_X3Y11_S1BEG[1] ,
    \Tile_X3Y11_S1BEG[0] }),
    .S1END({\Tile_X3Y10_S1BEG[3] ,
    \Tile_X3Y10_S1BEG[2] ,
    \Tile_X3Y10_S1BEG[1] ,
    \Tile_X3Y10_S1BEG[0] }),
    .S2BEG({\Tile_X3Y11_S2BEG[7] ,
    \Tile_X3Y11_S2BEG[6] ,
    \Tile_X3Y11_S2BEG[5] ,
    \Tile_X3Y11_S2BEG[4] ,
    \Tile_X3Y11_S2BEG[3] ,
    \Tile_X3Y11_S2BEG[2] ,
    \Tile_X3Y11_S2BEG[1] ,
    \Tile_X3Y11_S2BEG[0] }),
    .S2BEGb({\Tile_X3Y11_S2BEGb[7] ,
    \Tile_X3Y11_S2BEGb[6] ,
    \Tile_X3Y11_S2BEGb[5] ,
    \Tile_X3Y11_S2BEGb[4] ,
    \Tile_X3Y11_S2BEGb[3] ,
    \Tile_X3Y11_S2BEGb[2] ,
    \Tile_X3Y11_S2BEGb[1] ,
    \Tile_X3Y11_S2BEGb[0] }),
    .S2END({\Tile_X3Y10_S2BEGb[7] ,
    \Tile_X3Y10_S2BEGb[6] ,
    \Tile_X3Y10_S2BEGb[5] ,
    \Tile_X3Y10_S2BEGb[4] ,
    \Tile_X3Y10_S2BEGb[3] ,
    \Tile_X3Y10_S2BEGb[2] ,
    \Tile_X3Y10_S2BEGb[1] ,
    \Tile_X3Y10_S2BEGb[0] }),
    .S2MID({\Tile_X3Y10_S2BEG[7] ,
    \Tile_X3Y10_S2BEG[6] ,
    \Tile_X3Y10_S2BEG[5] ,
    \Tile_X3Y10_S2BEG[4] ,
    \Tile_X3Y10_S2BEG[3] ,
    \Tile_X3Y10_S2BEG[2] ,
    \Tile_X3Y10_S2BEG[1] ,
    \Tile_X3Y10_S2BEG[0] }),
    .S4BEG({\Tile_X3Y11_S4BEG[15] ,
    \Tile_X3Y11_S4BEG[14] ,
    \Tile_X3Y11_S4BEG[13] ,
    \Tile_X3Y11_S4BEG[12] ,
    \Tile_X3Y11_S4BEG[11] ,
    \Tile_X3Y11_S4BEG[10] ,
    \Tile_X3Y11_S4BEG[9] ,
    \Tile_X3Y11_S4BEG[8] ,
    \Tile_X3Y11_S4BEG[7] ,
    \Tile_X3Y11_S4BEG[6] ,
    \Tile_X3Y11_S4BEG[5] ,
    \Tile_X3Y11_S4BEG[4] ,
    \Tile_X3Y11_S4BEG[3] ,
    \Tile_X3Y11_S4BEG[2] ,
    \Tile_X3Y11_S4BEG[1] ,
    \Tile_X3Y11_S4BEG[0] }),
    .S4END({\Tile_X3Y10_S4BEG[15] ,
    \Tile_X3Y10_S4BEG[14] ,
    \Tile_X3Y10_S4BEG[13] ,
    \Tile_X3Y10_S4BEG[12] ,
    \Tile_X3Y10_S4BEG[11] ,
    \Tile_X3Y10_S4BEG[10] ,
    \Tile_X3Y10_S4BEG[9] ,
    \Tile_X3Y10_S4BEG[8] ,
    \Tile_X3Y10_S4BEG[7] ,
    \Tile_X3Y10_S4BEG[6] ,
    \Tile_X3Y10_S4BEG[5] ,
    \Tile_X3Y10_S4BEG[4] ,
    \Tile_X3Y10_S4BEG[3] ,
    \Tile_X3Y10_S4BEG[2] ,
    \Tile_X3Y10_S4BEG[1] ,
    \Tile_X3Y10_S4BEG[0] }),
    .SS4BEG({\Tile_X3Y11_SS4BEG[15] ,
    \Tile_X3Y11_SS4BEG[14] ,
    \Tile_X3Y11_SS4BEG[13] ,
    \Tile_X3Y11_SS4BEG[12] ,
    \Tile_X3Y11_SS4BEG[11] ,
    \Tile_X3Y11_SS4BEG[10] ,
    \Tile_X3Y11_SS4BEG[9] ,
    \Tile_X3Y11_SS4BEG[8] ,
    \Tile_X3Y11_SS4BEG[7] ,
    \Tile_X3Y11_SS4BEG[6] ,
    \Tile_X3Y11_SS4BEG[5] ,
    \Tile_X3Y11_SS4BEG[4] ,
    \Tile_X3Y11_SS4BEG[3] ,
    \Tile_X3Y11_SS4BEG[2] ,
    \Tile_X3Y11_SS4BEG[1] ,
    \Tile_X3Y11_SS4BEG[0] }),
    .SS4END({\Tile_X3Y10_SS4BEG[15] ,
    \Tile_X3Y10_SS4BEG[14] ,
    \Tile_X3Y10_SS4BEG[13] ,
    \Tile_X3Y10_SS4BEG[12] ,
    \Tile_X3Y10_SS4BEG[11] ,
    \Tile_X3Y10_SS4BEG[10] ,
    \Tile_X3Y10_SS4BEG[9] ,
    \Tile_X3Y10_SS4BEG[8] ,
    \Tile_X3Y10_SS4BEG[7] ,
    \Tile_X3Y10_SS4BEG[6] ,
    \Tile_X3Y10_SS4BEG[5] ,
    \Tile_X3Y10_SS4BEG[4] ,
    \Tile_X3Y10_SS4BEG[3] ,
    \Tile_X3Y10_SS4BEG[2] ,
    \Tile_X3Y10_SS4BEG[1] ,
    \Tile_X3Y10_SS4BEG[0] }),
    .W1BEG({\Tile_X3Y11_W1BEG[3] ,
    \Tile_X3Y11_W1BEG[2] ,
    \Tile_X3Y11_W1BEG[1] ,
    \Tile_X3Y11_W1BEG[0] }),
    .W1END({\Tile_X4Y11_W1BEG[3] ,
    \Tile_X4Y11_W1BEG[2] ,
    \Tile_X4Y11_W1BEG[1] ,
    \Tile_X4Y11_W1BEG[0] }),
    .W2BEG({\Tile_X3Y11_W2BEG[7] ,
    \Tile_X3Y11_W2BEG[6] ,
    \Tile_X3Y11_W2BEG[5] ,
    \Tile_X3Y11_W2BEG[4] ,
    \Tile_X3Y11_W2BEG[3] ,
    \Tile_X3Y11_W2BEG[2] ,
    \Tile_X3Y11_W2BEG[1] ,
    \Tile_X3Y11_W2BEG[0] }),
    .W2BEGb({\Tile_X3Y11_W2BEGb[7] ,
    \Tile_X3Y11_W2BEGb[6] ,
    \Tile_X3Y11_W2BEGb[5] ,
    \Tile_X3Y11_W2BEGb[4] ,
    \Tile_X3Y11_W2BEGb[3] ,
    \Tile_X3Y11_W2BEGb[2] ,
    \Tile_X3Y11_W2BEGb[1] ,
    \Tile_X3Y11_W2BEGb[0] }),
    .W2END({\Tile_X4Y11_W2BEGb[7] ,
    \Tile_X4Y11_W2BEGb[6] ,
    \Tile_X4Y11_W2BEGb[5] ,
    \Tile_X4Y11_W2BEGb[4] ,
    \Tile_X4Y11_W2BEGb[3] ,
    \Tile_X4Y11_W2BEGb[2] ,
    \Tile_X4Y11_W2BEGb[1] ,
    \Tile_X4Y11_W2BEGb[0] }),
    .W2MID({\Tile_X4Y11_W2BEG[7] ,
    \Tile_X4Y11_W2BEG[6] ,
    \Tile_X4Y11_W2BEG[5] ,
    \Tile_X4Y11_W2BEG[4] ,
    \Tile_X4Y11_W2BEG[3] ,
    \Tile_X4Y11_W2BEG[2] ,
    \Tile_X4Y11_W2BEG[1] ,
    \Tile_X4Y11_W2BEG[0] }),
    .W6BEG({\Tile_X3Y11_W6BEG[11] ,
    \Tile_X3Y11_W6BEG[10] ,
    \Tile_X3Y11_W6BEG[9] ,
    \Tile_X3Y11_W6BEG[8] ,
    \Tile_X3Y11_W6BEG[7] ,
    \Tile_X3Y11_W6BEG[6] ,
    \Tile_X3Y11_W6BEG[5] ,
    \Tile_X3Y11_W6BEG[4] ,
    \Tile_X3Y11_W6BEG[3] ,
    \Tile_X3Y11_W6BEG[2] ,
    \Tile_X3Y11_W6BEG[1] ,
    \Tile_X3Y11_W6BEG[0] }),
    .W6END({\Tile_X4Y11_W6BEG[11] ,
    \Tile_X4Y11_W6BEG[10] ,
    \Tile_X4Y11_W6BEG[9] ,
    \Tile_X4Y11_W6BEG[8] ,
    \Tile_X4Y11_W6BEG[7] ,
    \Tile_X4Y11_W6BEG[6] ,
    \Tile_X4Y11_W6BEG[5] ,
    \Tile_X4Y11_W6BEG[4] ,
    \Tile_X4Y11_W6BEG[3] ,
    \Tile_X4Y11_W6BEG[2] ,
    \Tile_X4Y11_W6BEG[1] ,
    \Tile_X4Y11_W6BEG[0] }),
    .WW4BEG({\Tile_X3Y11_WW4BEG[15] ,
    \Tile_X3Y11_WW4BEG[14] ,
    \Tile_X3Y11_WW4BEG[13] ,
    \Tile_X3Y11_WW4BEG[12] ,
    \Tile_X3Y11_WW4BEG[11] ,
    \Tile_X3Y11_WW4BEG[10] ,
    \Tile_X3Y11_WW4BEG[9] ,
    \Tile_X3Y11_WW4BEG[8] ,
    \Tile_X3Y11_WW4BEG[7] ,
    \Tile_X3Y11_WW4BEG[6] ,
    \Tile_X3Y11_WW4BEG[5] ,
    \Tile_X3Y11_WW4BEG[4] ,
    \Tile_X3Y11_WW4BEG[3] ,
    \Tile_X3Y11_WW4BEG[2] ,
    \Tile_X3Y11_WW4BEG[1] ,
    \Tile_X3Y11_WW4BEG[0] }),
    .WW4END({\Tile_X4Y11_WW4BEG[15] ,
    \Tile_X4Y11_WW4BEG[14] ,
    \Tile_X4Y11_WW4BEG[13] ,
    \Tile_X4Y11_WW4BEG[12] ,
    \Tile_X4Y11_WW4BEG[11] ,
    \Tile_X4Y11_WW4BEG[10] ,
    \Tile_X4Y11_WW4BEG[9] ,
    \Tile_X4Y11_WW4BEG[8] ,
    \Tile_X4Y11_WW4BEG[7] ,
    \Tile_X4Y11_WW4BEG[6] ,
    \Tile_X4Y11_WW4BEG[5] ,
    \Tile_X4Y11_WW4BEG[4] ,
    \Tile_X4Y11_WW4BEG[3] ,
    \Tile_X4Y11_WW4BEG[2] ,
    \Tile_X4Y11_WW4BEG[1] ,
    \Tile_X4Y11_WW4BEG[0] }));
 LUT4AB Tile_X3Y12_LUT4AB (.Ci(Tile_X3Y13_Co),
    .Co(Tile_X3Y12_Co),
    .UserCLK(Tile_X3Y13_UserCLKo),
    .UserCLKo(Tile_X3Y12_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X3Y12_E1BEG[3] ,
    \Tile_X3Y12_E1BEG[2] ,
    \Tile_X3Y12_E1BEG[1] ,
    \Tile_X3Y12_E1BEG[0] }),
    .E1END({\Tile_X2Y12_E1BEG[3] ,
    \Tile_X2Y12_E1BEG[2] ,
    \Tile_X2Y12_E1BEG[1] ,
    \Tile_X2Y12_E1BEG[0] }),
    .E2BEG({\Tile_X3Y12_E2BEG[7] ,
    \Tile_X3Y12_E2BEG[6] ,
    \Tile_X3Y12_E2BEG[5] ,
    \Tile_X3Y12_E2BEG[4] ,
    \Tile_X3Y12_E2BEG[3] ,
    \Tile_X3Y12_E2BEG[2] ,
    \Tile_X3Y12_E2BEG[1] ,
    \Tile_X3Y12_E2BEG[0] }),
    .E2BEGb({\Tile_X3Y12_E2BEGb[7] ,
    \Tile_X3Y12_E2BEGb[6] ,
    \Tile_X3Y12_E2BEGb[5] ,
    \Tile_X3Y12_E2BEGb[4] ,
    \Tile_X3Y12_E2BEGb[3] ,
    \Tile_X3Y12_E2BEGb[2] ,
    \Tile_X3Y12_E2BEGb[1] ,
    \Tile_X3Y12_E2BEGb[0] }),
    .E2END({\Tile_X2Y12_E2BEGb[7] ,
    \Tile_X2Y12_E2BEGb[6] ,
    \Tile_X2Y12_E2BEGb[5] ,
    \Tile_X2Y12_E2BEGb[4] ,
    \Tile_X2Y12_E2BEGb[3] ,
    \Tile_X2Y12_E2BEGb[2] ,
    \Tile_X2Y12_E2BEGb[1] ,
    \Tile_X2Y12_E2BEGb[0] }),
    .E2MID({\Tile_X2Y12_E2BEG[7] ,
    \Tile_X2Y12_E2BEG[6] ,
    \Tile_X2Y12_E2BEG[5] ,
    \Tile_X2Y12_E2BEG[4] ,
    \Tile_X2Y12_E2BEG[3] ,
    \Tile_X2Y12_E2BEG[2] ,
    \Tile_X2Y12_E2BEG[1] ,
    \Tile_X2Y12_E2BEG[0] }),
    .E6BEG({\Tile_X3Y12_E6BEG[11] ,
    \Tile_X3Y12_E6BEG[10] ,
    \Tile_X3Y12_E6BEG[9] ,
    \Tile_X3Y12_E6BEG[8] ,
    \Tile_X3Y12_E6BEG[7] ,
    \Tile_X3Y12_E6BEG[6] ,
    \Tile_X3Y12_E6BEG[5] ,
    \Tile_X3Y12_E6BEG[4] ,
    \Tile_X3Y12_E6BEG[3] ,
    \Tile_X3Y12_E6BEG[2] ,
    \Tile_X3Y12_E6BEG[1] ,
    \Tile_X3Y12_E6BEG[0] }),
    .E6END({\Tile_X2Y12_E6BEG[11] ,
    \Tile_X2Y12_E6BEG[10] ,
    \Tile_X2Y12_E6BEG[9] ,
    \Tile_X2Y12_E6BEG[8] ,
    \Tile_X2Y12_E6BEG[7] ,
    \Tile_X2Y12_E6BEG[6] ,
    \Tile_X2Y12_E6BEG[5] ,
    \Tile_X2Y12_E6BEG[4] ,
    \Tile_X2Y12_E6BEG[3] ,
    \Tile_X2Y12_E6BEG[2] ,
    \Tile_X2Y12_E6BEG[1] ,
    \Tile_X2Y12_E6BEG[0] }),
    .EE4BEG({\Tile_X3Y12_EE4BEG[15] ,
    \Tile_X3Y12_EE4BEG[14] ,
    \Tile_X3Y12_EE4BEG[13] ,
    \Tile_X3Y12_EE4BEG[12] ,
    \Tile_X3Y12_EE4BEG[11] ,
    \Tile_X3Y12_EE4BEG[10] ,
    \Tile_X3Y12_EE4BEG[9] ,
    \Tile_X3Y12_EE4BEG[8] ,
    \Tile_X3Y12_EE4BEG[7] ,
    \Tile_X3Y12_EE4BEG[6] ,
    \Tile_X3Y12_EE4BEG[5] ,
    \Tile_X3Y12_EE4BEG[4] ,
    \Tile_X3Y12_EE4BEG[3] ,
    \Tile_X3Y12_EE4BEG[2] ,
    \Tile_X3Y12_EE4BEG[1] ,
    \Tile_X3Y12_EE4BEG[0] }),
    .EE4END({\Tile_X2Y12_EE4BEG[15] ,
    \Tile_X2Y12_EE4BEG[14] ,
    \Tile_X2Y12_EE4BEG[13] ,
    \Tile_X2Y12_EE4BEG[12] ,
    \Tile_X2Y12_EE4BEG[11] ,
    \Tile_X2Y12_EE4BEG[10] ,
    \Tile_X2Y12_EE4BEG[9] ,
    \Tile_X2Y12_EE4BEG[8] ,
    \Tile_X2Y12_EE4BEG[7] ,
    \Tile_X2Y12_EE4BEG[6] ,
    \Tile_X2Y12_EE4BEG[5] ,
    \Tile_X2Y12_EE4BEG[4] ,
    \Tile_X2Y12_EE4BEG[3] ,
    \Tile_X2Y12_EE4BEG[2] ,
    \Tile_X2Y12_EE4BEG[1] ,
    \Tile_X2Y12_EE4BEG[0] }),
    .FrameData({\Tile_X2Y12_FrameData_O[31] ,
    \Tile_X2Y12_FrameData_O[30] ,
    \Tile_X2Y12_FrameData_O[29] ,
    \Tile_X2Y12_FrameData_O[28] ,
    \Tile_X2Y12_FrameData_O[27] ,
    \Tile_X2Y12_FrameData_O[26] ,
    \Tile_X2Y12_FrameData_O[25] ,
    \Tile_X2Y12_FrameData_O[24] ,
    \Tile_X2Y12_FrameData_O[23] ,
    \Tile_X2Y12_FrameData_O[22] ,
    \Tile_X2Y12_FrameData_O[21] ,
    \Tile_X2Y12_FrameData_O[20] ,
    \Tile_X2Y12_FrameData_O[19] ,
    \Tile_X2Y12_FrameData_O[18] ,
    \Tile_X2Y12_FrameData_O[17] ,
    \Tile_X2Y12_FrameData_O[16] ,
    \Tile_X2Y12_FrameData_O[15] ,
    \Tile_X2Y12_FrameData_O[14] ,
    \Tile_X2Y12_FrameData_O[13] ,
    \Tile_X2Y12_FrameData_O[12] ,
    \Tile_X2Y12_FrameData_O[11] ,
    \Tile_X2Y12_FrameData_O[10] ,
    \Tile_X2Y12_FrameData_O[9] ,
    \Tile_X2Y12_FrameData_O[8] ,
    \Tile_X2Y12_FrameData_O[7] ,
    \Tile_X2Y12_FrameData_O[6] ,
    \Tile_X2Y12_FrameData_O[5] ,
    \Tile_X2Y12_FrameData_O[4] ,
    \Tile_X2Y12_FrameData_O[3] ,
    \Tile_X2Y12_FrameData_O[2] ,
    \Tile_X2Y12_FrameData_O[1] ,
    \Tile_X2Y12_FrameData_O[0] }),
    .FrameData_O({\Tile_X3Y12_FrameData_O[31] ,
    \Tile_X3Y12_FrameData_O[30] ,
    \Tile_X3Y12_FrameData_O[29] ,
    \Tile_X3Y12_FrameData_O[28] ,
    \Tile_X3Y12_FrameData_O[27] ,
    \Tile_X3Y12_FrameData_O[26] ,
    \Tile_X3Y12_FrameData_O[25] ,
    \Tile_X3Y12_FrameData_O[24] ,
    \Tile_X3Y12_FrameData_O[23] ,
    \Tile_X3Y12_FrameData_O[22] ,
    \Tile_X3Y12_FrameData_O[21] ,
    \Tile_X3Y12_FrameData_O[20] ,
    \Tile_X3Y12_FrameData_O[19] ,
    \Tile_X3Y12_FrameData_O[18] ,
    \Tile_X3Y12_FrameData_O[17] ,
    \Tile_X3Y12_FrameData_O[16] ,
    \Tile_X3Y12_FrameData_O[15] ,
    \Tile_X3Y12_FrameData_O[14] ,
    \Tile_X3Y12_FrameData_O[13] ,
    \Tile_X3Y12_FrameData_O[12] ,
    \Tile_X3Y12_FrameData_O[11] ,
    \Tile_X3Y12_FrameData_O[10] ,
    \Tile_X3Y12_FrameData_O[9] ,
    \Tile_X3Y12_FrameData_O[8] ,
    \Tile_X3Y12_FrameData_O[7] ,
    \Tile_X3Y12_FrameData_O[6] ,
    \Tile_X3Y12_FrameData_O[5] ,
    \Tile_X3Y12_FrameData_O[4] ,
    \Tile_X3Y12_FrameData_O[3] ,
    \Tile_X3Y12_FrameData_O[2] ,
    \Tile_X3Y12_FrameData_O[1] ,
    \Tile_X3Y12_FrameData_O[0] }),
    .FrameStrobe({\Tile_X3Y13_FrameStrobe_O[19] ,
    \Tile_X3Y13_FrameStrobe_O[18] ,
    \Tile_X3Y13_FrameStrobe_O[17] ,
    \Tile_X3Y13_FrameStrobe_O[16] ,
    \Tile_X3Y13_FrameStrobe_O[15] ,
    \Tile_X3Y13_FrameStrobe_O[14] ,
    \Tile_X3Y13_FrameStrobe_O[13] ,
    \Tile_X3Y13_FrameStrobe_O[12] ,
    \Tile_X3Y13_FrameStrobe_O[11] ,
    \Tile_X3Y13_FrameStrobe_O[10] ,
    \Tile_X3Y13_FrameStrobe_O[9] ,
    \Tile_X3Y13_FrameStrobe_O[8] ,
    \Tile_X3Y13_FrameStrobe_O[7] ,
    \Tile_X3Y13_FrameStrobe_O[6] ,
    \Tile_X3Y13_FrameStrobe_O[5] ,
    \Tile_X3Y13_FrameStrobe_O[4] ,
    \Tile_X3Y13_FrameStrobe_O[3] ,
    \Tile_X3Y13_FrameStrobe_O[2] ,
    \Tile_X3Y13_FrameStrobe_O[1] ,
    \Tile_X3Y13_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X3Y12_FrameStrobe_O[19] ,
    \Tile_X3Y12_FrameStrobe_O[18] ,
    \Tile_X3Y12_FrameStrobe_O[17] ,
    \Tile_X3Y12_FrameStrobe_O[16] ,
    \Tile_X3Y12_FrameStrobe_O[15] ,
    \Tile_X3Y12_FrameStrobe_O[14] ,
    \Tile_X3Y12_FrameStrobe_O[13] ,
    \Tile_X3Y12_FrameStrobe_O[12] ,
    \Tile_X3Y12_FrameStrobe_O[11] ,
    \Tile_X3Y12_FrameStrobe_O[10] ,
    \Tile_X3Y12_FrameStrobe_O[9] ,
    \Tile_X3Y12_FrameStrobe_O[8] ,
    \Tile_X3Y12_FrameStrobe_O[7] ,
    \Tile_X3Y12_FrameStrobe_O[6] ,
    \Tile_X3Y12_FrameStrobe_O[5] ,
    \Tile_X3Y12_FrameStrobe_O[4] ,
    \Tile_X3Y12_FrameStrobe_O[3] ,
    \Tile_X3Y12_FrameStrobe_O[2] ,
    \Tile_X3Y12_FrameStrobe_O[1] ,
    \Tile_X3Y12_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X3Y12_N1BEG[3] ,
    \Tile_X3Y12_N1BEG[2] ,
    \Tile_X3Y12_N1BEG[1] ,
    \Tile_X3Y12_N1BEG[0] }),
    .N1END({\Tile_X3Y13_N1BEG[3] ,
    \Tile_X3Y13_N1BEG[2] ,
    \Tile_X3Y13_N1BEG[1] ,
    \Tile_X3Y13_N1BEG[0] }),
    .N2BEG({\Tile_X3Y12_N2BEG[7] ,
    \Tile_X3Y12_N2BEG[6] ,
    \Tile_X3Y12_N2BEG[5] ,
    \Tile_X3Y12_N2BEG[4] ,
    \Tile_X3Y12_N2BEG[3] ,
    \Tile_X3Y12_N2BEG[2] ,
    \Tile_X3Y12_N2BEG[1] ,
    \Tile_X3Y12_N2BEG[0] }),
    .N2BEGb({\Tile_X3Y12_N2BEGb[7] ,
    \Tile_X3Y12_N2BEGb[6] ,
    \Tile_X3Y12_N2BEGb[5] ,
    \Tile_X3Y12_N2BEGb[4] ,
    \Tile_X3Y12_N2BEGb[3] ,
    \Tile_X3Y12_N2BEGb[2] ,
    \Tile_X3Y12_N2BEGb[1] ,
    \Tile_X3Y12_N2BEGb[0] }),
    .N2END({\Tile_X3Y13_N2BEGb[7] ,
    \Tile_X3Y13_N2BEGb[6] ,
    \Tile_X3Y13_N2BEGb[5] ,
    \Tile_X3Y13_N2BEGb[4] ,
    \Tile_X3Y13_N2BEGb[3] ,
    \Tile_X3Y13_N2BEGb[2] ,
    \Tile_X3Y13_N2BEGb[1] ,
    \Tile_X3Y13_N2BEGb[0] }),
    .N2MID({\Tile_X3Y13_N2BEG[7] ,
    \Tile_X3Y13_N2BEG[6] ,
    \Tile_X3Y13_N2BEG[5] ,
    \Tile_X3Y13_N2BEG[4] ,
    \Tile_X3Y13_N2BEG[3] ,
    \Tile_X3Y13_N2BEG[2] ,
    \Tile_X3Y13_N2BEG[1] ,
    \Tile_X3Y13_N2BEG[0] }),
    .N4BEG({\Tile_X3Y12_N4BEG[15] ,
    \Tile_X3Y12_N4BEG[14] ,
    \Tile_X3Y12_N4BEG[13] ,
    \Tile_X3Y12_N4BEG[12] ,
    \Tile_X3Y12_N4BEG[11] ,
    \Tile_X3Y12_N4BEG[10] ,
    \Tile_X3Y12_N4BEG[9] ,
    \Tile_X3Y12_N4BEG[8] ,
    \Tile_X3Y12_N4BEG[7] ,
    \Tile_X3Y12_N4BEG[6] ,
    \Tile_X3Y12_N4BEG[5] ,
    \Tile_X3Y12_N4BEG[4] ,
    \Tile_X3Y12_N4BEG[3] ,
    \Tile_X3Y12_N4BEG[2] ,
    \Tile_X3Y12_N4BEG[1] ,
    \Tile_X3Y12_N4BEG[0] }),
    .N4END({\Tile_X3Y13_N4BEG[15] ,
    \Tile_X3Y13_N4BEG[14] ,
    \Tile_X3Y13_N4BEG[13] ,
    \Tile_X3Y13_N4BEG[12] ,
    \Tile_X3Y13_N4BEG[11] ,
    \Tile_X3Y13_N4BEG[10] ,
    \Tile_X3Y13_N4BEG[9] ,
    \Tile_X3Y13_N4BEG[8] ,
    \Tile_X3Y13_N4BEG[7] ,
    \Tile_X3Y13_N4BEG[6] ,
    \Tile_X3Y13_N4BEG[5] ,
    \Tile_X3Y13_N4BEG[4] ,
    \Tile_X3Y13_N4BEG[3] ,
    \Tile_X3Y13_N4BEG[2] ,
    \Tile_X3Y13_N4BEG[1] ,
    \Tile_X3Y13_N4BEG[0] }),
    .NN4BEG({\Tile_X3Y12_NN4BEG[15] ,
    \Tile_X3Y12_NN4BEG[14] ,
    \Tile_X3Y12_NN4BEG[13] ,
    \Tile_X3Y12_NN4BEG[12] ,
    \Tile_X3Y12_NN4BEG[11] ,
    \Tile_X3Y12_NN4BEG[10] ,
    \Tile_X3Y12_NN4BEG[9] ,
    \Tile_X3Y12_NN4BEG[8] ,
    \Tile_X3Y12_NN4BEG[7] ,
    \Tile_X3Y12_NN4BEG[6] ,
    \Tile_X3Y12_NN4BEG[5] ,
    \Tile_X3Y12_NN4BEG[4] ,
    \Tile_X3Y12_NN4BEG[3] ,
    \Tile_X3Y12_NN4BEG[2] ,
    \Tile_X3Y12_NN4BEG[1] ,
    \Tile_X3Y12_NN4BEG[0] }),
    .NN4END({\Tile_X3Y13_NN4BEG[15] ,
    \Tile_X3Y13_NN4BEG[14] ,
    \Tile_X3Y13_NN4BEG[13] ,
    \Tile_X3Y13_NN4BEG[12] ,
    \Tile_X3Y13_NN4BEG[11] ,
    \Tile_X3Y13_NN4BEG[10] ,
    \Tile_X3Y13_NN4BEG[9] ,
    \Tile_X3Y13_NN4BEG[8] ,
    \Tile_X3Y13_NN4BEG[7] ,
    \Tile_X3Y13_NN4BEG[6] ,
    \Tile_X3Y13_NN4BEG[5] ,
    \Tile_X3Y13_NN4BEG[4] ,
    \Tile_X3Y13_NN4BEG[3] ,
    \Tile_X3Y13_NN4BEG[2] ,
    \Tile_X3Y13_NN4BEG[1] ,
    \Tile_X3Y13_NN4BEG[0] }),
    .S1BEG({\Tile_X3Y12_S1BEG[3] ,
    \Tile_X3Y12_S1BEG[2] ,
    \Tile_X3Y12_S1BEG[1] ,
    \Tile_X3Y12_S1BEG[0] }),
    .S1END({\Tile_X3Y11_S1BEG[3] ,
    \Tile_X3Y11_S1BEG[2] ,
    \Tile_X3Y11_S1BEG[1] ,
    \Tile_X3Y11_S1BEG[0] }),
    .S2BEG({\Tile_X3Y12_S2BEG[7] ,
    \Tile_X3Y12_S2BEG[6] ,
    \Tile_X3Y12_S2BEG[5] ,
    \Tile_X3Y12_S2BEG[4] ,
    \Tile_X3Y12_S2BEG[3] ,
    \Tile_X3Y12_S2BEG[2] ,
    \Tile_X3Y12_S2BEG[1] ,
    \Tile_X3Y12_S2BEG[0] }),
    .S2BEGb({\Tile_X3Y12_S2BEGb[7] ,
    \Tile_X3Y12_S2BEGb[6] ,
    \Tile_X3Y12_S2BEGb[5] ,
    \Tile_X3Y12_S2BEGb[4] ,
    \Tile_X3Y12_S2BEGb[3] ,
    \Tile_X3Y12_S2BEGb[2] ,
    \Tile_X3Y12_S2BEGb[1] ,
    \Tile_X3Y12_S2BEGb[0] }),
    .S2END({\Tile_X3Y11_S2BEGb[7] ,
    \Tile_X3Y11_S2BEGb[6] ,
    \Tile_X3Y11_S2BEGb[5] ,
    \Tile_X3Y11_S2BEGb[4] ,
    \Tile_X3Y11_S2BEGb[3] ,
    \Tile_X3Y11_S2BEGb[2] ,
    \Tile_X3Y11_S2BEGb[1] ,
    \Tile_X3Y11_S2BEGb[0] }),
    .S2MID({\Tile_X3Y11_S2BEG[7] ,
    \Tile_X3Y11_S2BEG[6] ,
    \Tile_X3Y11_S2BEG[5] ,
    \Tile_X3Y11_S2BEG[4] ,
    \Tile_X3Y11_S2BEG[3] ,
    \Tile_X3Y11_S2BEG[2] ,
    \Tile_X3Y11_S2BEG[1] ,
    \Tile_X3Y11_S2BEG[0] }),
    .S4BEG({\Tile_X3Y12_S4BEG[15] ,
    \Tile_X3Y12_S4BEG[14] ,
    \Tile_X3Y12_S4BEG[13] ,
    \Tile_X3Y12_S4BEG[12] ,
    \Tile_X3Y12_S4BEG[11] ,
    \Tile_X3Y12_S4BEG[10] ,
    \Tile_X3Y12_S4BEG[9] ,
    \Tile_X3Y12_S4BEG[8] ,
    \Tile_X3Y12_S4BEG[7] ,
    \Tile_X3Y12_S4BEG[6] ,
    \Tile_X3Y12_S4BEG[5] ,
    \Tile_X3Y12_S4BEG[4] ,
    \Tile_X3Y12_S4BEG[3] ,
    \Tile_X3Y12_S4BEG[2] ,
    \Tile_X3Y12_S4BEG[1] ,
    \Tile_X3Y12_S4BEG[0] }),
    .S4END({\Tile_X3Y11_S4BEG[15] ,
    \Tile_X3Y11_S4BEG[14] ,
    \Tile_X3Y11_S4BEG[13] ,
    \Tile_X3Y11_S4BEG[12] ,
    \Tile_X3Y11_S4BEG[11] ,
    \Tile_X3Y11_S4BEG[10] ,
    \Tile_X3Y11_S4BEG[9] ,
    \Tile_X3Y11_S4BEG[8] ,
    \Tile_X3Y11_S4BEG[7] ,
    \Tile_X3Y11_S4BEG[6] ,
    \Tile_X3Y11_S4BEG[5] ,
    \Tile_X3Y11_S4BEG[4] ,
    \Tile_X3Y11_S4BEG[3] ,
    \Tile_X3Y11_S4BEG[2] ,
    \Tile_X3Y11_S4BEG[1] ,
    \Tile_X3Y11_S4BEG[0] }),
    .SS4BEG({\Tile_X3Y12_SS4BEG[15] ,
    \Tile_X3Y12_SS4BEG[14] ,
    \Tile_X3Y12_SS4BEG[13] ,
    \Tile_X3Y12_SS4BEG[12] ,
    \Tile_X3Y12_SS4BEG[11] ,
    \Tile_X3Y12_SS4BEG[10] ,
    \Tile_X3Y12_SS4BEG[9] ,
    \Tile_X3Y12_SS4BEG[8] ,
    \Tile_X3Y12_SS4BEG[7] ,
    \Tile_X3Y12_SS4BEG[6] ,
    \Tile_X3Y12_SS4BEG[5] ,
    \Tile_X3Y12_SS4BEG[4] ,
    \Tile_X3Y12_SS4BEG[3] ,
    \Tile_X3Y12_SS4BEG[2] ,
    \Tile_X3Y12_SS4BEG[1] ,
    \Tile_X3Y12_SS4BEG[0] }),
    .SS4END({\Tile_X3Y11_SS4BEG[15] ,
    \Tile_X3Y11_SS4BEG[14] ,
    \Tile_X3Y11_SS4BEG[13] ,
    \Tile_X3Y11_SS4BEG[12] ,
    \Tile_X3Y11_SS4BEG[11] ,
    \Tile_X3Y11_SS4BEG[10] ,
    \Tile_X3Y11_SS4BEG[9] ,
    \Tile_X3Y11_SS4BEG[8] ,
    \Tile_X3Y11_SS4BEG[7] ,
    \Tile_X3Y11_SS4BEG[6] ,
    \Tile_X3Y11_SS4BEG[5] ,
    \Tile_X3Y11_SS4BEG[4] ,
    \Tile_X3Y11_SS4BEG[3] ,
    \Tile_X3Y11_SS4BEG[2] ,
    \Tile_X3Y11_SS4BEG[1] ,
    \Tile_X3Y11_SS4BEG[0] }),
    .W1BEG({\Tile_X3Y12_W1BEG[3] ,
    \Tile_X3Y12_W1BEG[2] ,
    \Tile_X3Y12_W1BEG[1] ,
    \Tile_X3Y12_W1BEG[0] }),
    .W1END({\Tile_X4Y12_W1BEG[3] ,
    \Tile_X4Y12_W1BEG[2] ,
    \Tile_X4Y12_W1BEG[1] ,
    \Tile_X4Y12_W1BEG[0] }),
    .W2BEG({\Tile_X3Y12_W2BEG[7] ,
    \Tile_X3Y12_W2BEG[6] ,
    \Tile_X3Y12_W2BEG[5] ,
    \Tile_X3Y12_W2BEG[4] ,
    \Tile_X3Y12_W2BEG[3] ,
    \Tile_X3Y12_W2BEG[2] ,
    \Tile_X3Y12_W2BEG[1] ,
    \Tile_X3Y12_W2BEG[0] }),
    .W2BEGb({\Tile_X3Y12_W2BEGb[7] ,
    \Tile_X3Y12_W2BEGb[6] ,
    \Tile_X3Y12_W2BEGb[5] ,
    \Tile_X3Y12_W2BEGb[4] ,
    \Tile_X3Y12_W2BEGb[3] ,
    \Tile_X3Y12_W2BEGb[2] ,
    \Tile_X3Y12_W2BEGb[1] ,
    \Tile_X3Y12_W2BEGb[0] }),
    .W2END({\Tile_X4Y12_W2BEGb[7] ,
    \Tile_X4Y12_W2BEGb[6] ,
    \Tile_X4Y12_W2BEGb[5] ,
    \Tile_X4Y12_W2BEGb[4] ,
    \Tile_X4Y12_W2BEGb[3] ,
    \Tile_X4Y12_W2BEGb[2] ,
    \Tile_X4Y12_W2BEGb[1] ,
    \Tile_X4Y12_W2BEGb[0] }),
    .W2MID({\Tile_X4Y12_W2BEG[7] ,
    \Tile_X4Y12_W2BEG[6] ,
    \Tile_X4Y12_W2BEG[5] ,
    \Tile_X4Y12_W2BEG[4] ,
    \Tile_X4Y12_W2BEG[3] ,
    \Tile_X4Y12_W2BEG[2] ,
    \Tile_X4Y12_W2BEG[1] ,
    \Tile_X4Y12_W2BEG[0] }),
    .W6BEG({\Tile_X3Y12_W6BEG[11] ,
    \Tile_X3Y12_W6BEG[10] ,
    \Tile_X3Y12_W6BEG[9] ,
    \Tile_X3Y12_W6BEG[8] ,
    \Tile_X3Y12_W6BEG[7] ,
    \Tile_X3Y12_W6BEG[6] ,
    \Tile_X3Y12_W6BEG[5] ,
    \Tile_X3Y12_W6BEG[4] ,
    \Tile_X3Y12_W6BEG[3] ,
    \Tile_X3Y12_W6BEG[2] ,
    \Tile_X3Y12_W6BEG[1] ,
    \Tile_X3Y12_W6BEG[0] }),
    .W6END({\Tile_X4Y12_W6BEG[11] ,
    \Tile_X4Y12_W6BEG[10] ,
    \Tile_X4Y12_W6BEG[9] ,
    \Tile_X4Y12_W6BEG[8] ,
    \Tile_X4Y12_W6BEG[7] ,
    \Tile_X4Y12_W6BEG[6] ,
    \Tile_X4Y12_W6BEG[5] ,
    \Tile_X4Y12_W6BEG[4] ,
    \Tile_X4Y12_W6BEG[3] ,
    \Tile_X4Y12_W6BEG[2] ,
    \Tile_X4Y12_W6BEG[1] ,
    \Tile_X4Y12_W6BEG[0] }),
    .WW4BEG({\Tile_X3Y12_WW4BEG[15] ,
    \Tile_X3Y12_WW4BEG[14] ,
    \Tile_X3Y12_WW4BEG[13] ,
    \Tile_X3Y12_WW4BEG[12] ,
    \Tile_X3Y12_WW4BEG[11] ,
    \Tile_X3Y12_WW4BEG[10] ,
    \Tile_X3Y12_WW4BEG[9] ,
    \Tile_X3Y12_WW4BEG[8] ,
    \Tile_X3Y12_WW4BEG[7] ,
    \Tile_X3Y12_WW4BEG[6] ,
    \Tile_X3Y12_WW4BEG[5] ,
    \Tile_X3Y12_WW4BEG[4] ,
    \Tile_X3Y12_WW4BEG[3] ,
    \Tile_X3Y12_WW4BEG[2] ,
    \Tile_X3Y12_WW4BEG[1] ,
    \Tile_X3Y12_WW4BEG[0] }),
    .WW4END({\Tile_X4Y12_WW4BEG[15] ,
    \Tile_X4Y12_WW4BEG[14] ,
    \Tile_X4Y12_WW4BEG[13] ,
    \Tile_X4Y12_WW4BEG[12] ,
    \Tile_X4Y12_WW4BEG[11] ,
    \Tile_X4Y12_WW4BEG[10] ,
    \Tile_X4Y12_WW4BEG[9] ,
    \Tile_X4Y12_WW4BEG[8] ,
    \Tile_X4Y12_WW4BEG[7] ,
    \Tile_X4Y12_WW4BEG[6] ,
    \Tile_X4Y12_WW4BEG[5] ,
    \Tile_X4Y12_WW4BEG[4] ,
    \Tile_X4Y12_WW4BEG[3] ,
    \Tile_X4Y12_WW4BEG[2] ,
    \Tile_X4Y12_WW4BEG[1] ,
    \Tile_X4Y12_WW4BEG[0] }));
 LUT4AB Tile_X3Y13_LUT4AB (.Ci(Tile_X3Y14_Co),
    .Co(Tile_X3Y13_Co),
    .UserCLK(Tile_X3Y14_UserCLKo),
    .UserCLKo(Tile_X3Y13_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X3Y13_E1BEG[3] ,
    \Tile_X3Y13_E1BEG[2] ,
    \Tile_X3Y13_E1BEG[1] ,
    \Tile_X3Y13_E1BEG[0] }),
    .E1END({\Tile_X2Y13_E1BEG[3] ,
    \Tile_X2Y13_E1BEG[2] ,
    \Tile_X2Y13_E1BEG[1] ,
    \Tile_X2Y13_E1BEG[0] }),
    .E2BEG({\Tile_X3Y13_E2BEG[7] ,
    \Tile_X3Y13_E2BEG[6] ,
    \Tile_X3Y13_E2BEG[5] ,
    \Tile_X3Y13_E2BEG[4] ,
    \Tile_X3Y13_E2BEG[3] ,
    \Tile_X3Y13_E2BEG[2] ,
    \Tile_X3Y13_E2BEG[1] ,
    \Tile_X3Y13_E2BEG[0] }),
    .E2BEGb({\Tile_X3Y13_E2BEGb[7] ,
    \Tile_X3Y13_E2BEGb[6] ,
    \Tile_X3Y13_E2BEGb[5] ,
    \Tile_X3Y13_E2BEGb[4] ,
    \Tile_X3Y13_E2BEGb[3] ,
    \Tile_X3Y13_E2BEGb[2] ,
    \Tile_X3Y13_E2BEGb[1] ,
    \Tile_X3Y13_E2BEGb[0] }),
    .E2END({\Tile_X2Y13_E2BEGb[7] ,
    \Tile_X2Y13_E2BEGb[6] ,
    \Tile_X2Y13_E2BEGb[5] ,
    \Tile_X2Y13_E2BEGb[4] ,
    \Tile_X2Y13_E2BEGb[3] ,
    \Tile_X2Y13_E2BEGb[2] ,
    \Tile_X2Y13_E2BEGb[1] ,
    \Tile_X2Y13_E2BEGb[0] }),
    .E2MID({\Tile_X2Y13_E2BEG[7] ,
    \Tile_X2Y13_E2BEG[6] ,
    \Tile_X2Y13_E2BEG[5] ,
    \Tile_X2Y13_E2BEG[4] ,
    \Tile_X2Y13_E2BEG[3] ,
    \Tile_X2Y13_E2BEG[2] ,
    \Tile_X2Y13_E2BEG[1] ,
    \Tile_X2Y13_E2BEG[0] }),
    .E6BEG({\Tile_X3Y13_E6BEG[11] ,
    \Tile_X3Y13_E6BEG[10] ,
    \Tile_X3Y13_E6BEG[9] ,
    \Tile_X3Y13_E6BEG[8] ,
    \Tile_X3Y13_E6BEG[7] ,
    \Tile_X3Y13_E6BEG[6] ,
    \Tile_X3Y13_E6BEG[5] ,
    \Tile_X3Y13_E6BEG[4] ,
    \Tile_X3Y13_E6BEG[3] ,
    \Tile_X3Y13_E6BEG[2] ,
    \Tile_X3Y13_E6BEG[1] ,
    \Tile_X3Y13_E6BEG[0] }),
    .E6END({\Tile_X2Y13_E6BEG[11] ,
    \Tile_X2Y13_E6BEG[10] ,
    \Tile_X2Y13_E6BEG[9] ,
    \Tile_X2Y13_E6BEG[8] ,
    \Tile_X2Y13_E6BEG[7] ,
    \Tile_X2Y13_E6BEG[6] ,
    \Tile_X2Y13_E6BEG[5] ,
    \Tile_X2Y13_E6BEG[4] ,
    \Tile_X2Y13_E6BEG[3] ,
    \Tile_X2Y13_E6BEG[2] ,
    \Tile_X2Y13_E6BEG[1] ,
    \Tile_X2Y13_E6BEG[0] }),
    .EE4BEG({\Tile_X3Y13_EE4BEG[15] ,
    \Tile_X3Y13_EE4BEG[14] ,
    \Tile_X3Y13_EE4BEG[13] ,
    \Tile_X3Y13_EE4BEG[12] ,
    \Tile_X3Y13_EE4BEG[11] ,
    \Tile_X3Y13_EE4BEG[10] ,
    \Tile_X3Y13_EE4BEG[9] ,
    \Tile_X3Y13_EE4BEG[8] ,
    \Tile_X3Y13_EE4BEG[7] ,
    \Tile_X3Y13_EE4BEG[6] ,
    \Tile_X3Y13_EE4BEG[5] ,
    \Tile_X3Y13_EE4BEG[4] ,
    \Tile_X3Y13_EE4BEG[3] ,
    \Tile_X3Y13_EE4BEG[2] ,
    \Tile_X3Y13_EE4BEG[1] ,
    \Tile_X3Y13_EE4BEG[0] }),
    .EE4END({\Tile_X2Y13_EE4BEG[15] ,
    \Tile_X2Y13_EE4BEG[14] ,
    \Tile_X2Y13_EE4BEG[13] ,
    \Tile_X2Y13_EE4BEG[12] ,
    \Tile_X2Y13_EE4BEG[11] ,
    \Tile_X2Y13_EE4BEG[10] ,
    \Tile_X2Y13_EE4BEG[9] ,
    \Tile_X2Y13_EE4BEG[8] ,
    \Tile_X2Y13_EE4BEG[7] ,
    \Tile_X2Y13_EE4BEG[6] ,
    \Tile_X2Y13_EE4BEG[5] ,
    \Tile_X2Y13_EE4BEG[4] ,
    \Tile_X2Y13_EE4BEG[3] ,
    \Tile_X2Y13_EE4BEG[2] ,
    \Tile_X2Y13_EE4BEG[1] ,
    \Tile_X2Y13_EE4BEG[0] }),
    .FrameData({\Tile_X2Y13_FrameData_O[31] ,
    \Tile_X2Y13_FrameData_O[30] ,
    \Tile_X2Y13_FrameData_O[29] ,
    \Tile_X2Y13_FrameData_O[28] ,
    \Tile_X2Y13_FrameData_O[27] ,
    \Tile_X2Y13_FrameData_O[26] ,
    \Tile_X2Y13_FrameData_O[25] ,
    \Tile_X2Y13_FrameData_O[24] ,
    \Tile_X2Y13_FrameData_O[23] ,
    \Tile_X2Y13_FrameData_O[22] ,
    \Tile_X2Y13_FrameData_O[21] ,
    \Tile_X2Y13_FrameData_O[20] ,
    \Tile_X2Y13_FrameData_O[19] ,
    \Tile_X2Y13_FrameData_O[18] ,
    \Tile_X2Y13_FrameData_O[17] ,
    \Tile_X2Y13_FrameData_O[16] ,
    \Tile_X2Y13_FrameData_O[15] ,
    \Tile_X2Y13_FrameData_O[14] ,
    \Tile_X2Y13_FrameData_O[13] ,
    \Tile_X2Y13_FrameData_O[12] ,
    \Tile_X2Y13_FrameData_O[11] ,
    \Tile_X2Y13_FrameData_O[10] ,
    \Tile_X2Y13_FrameData_O[9] ,
    \Tile_X2Y13_FrameData_O[8] ,
    \Tile_X2Y13_FrameData_O[7] ,
    \Tile_X2Y13_FrameData_O[6] ,
    \Tile_X2Y13_FrameData_O[5] ,
    \Tile_X2Y13_FrameData_O[4] ,
    \Tile_X2Y13_FrameData_O[3] ,
    \Tile_X2Y13_FrameData_O[2] ,
    \Tile_X2Y13_FrameData_O[1] ,
    \Tile_X2Y13_FrameData_O[0] }),
    .FrameData_O({\Tile_X3Y13_FrameData_O[31] ,
    \Tile_X3Y13_FrameData_O[30] ,
    \Tile_X3Y13_FrameData_O[29] ,
    \Tile_X3Y13_FrameData_O[28] ,
    \Tile_X3Y13_FrameData_O[27] ,
    \Tile_X3Y13_FrameData_O[26] ,
    \Tile_X3Y13_FrameData_O[25] ,
    \Tile_X3Y13_FrameData_O[24] ,
    \Tile_X3Y13_FrameData_O[23] ,
    \Tile_X3Y13_FrameData_O[22] ,
    \Tile_X3Y13_FrameData_O[21] ,
    \Tile_X3Y13_FrameData_O[20] ,
    \Tile_X3Y13_FrameData_O[19] ,
    \Tile_X3Y13_FrameData_O[18] ,
    \Tile_X3Y13_FrameData_O[17] ,
    \Tile_X3Y13_FrameData_O[16] ,
    \Tile_X3Y13_FrameData_O[15] ,
    \Tile_X3Y13_FrameData_O[14] ,
    \Tile_X3Y13_FrameData_O[13] ,
    \Tile_X3Y13_FrameData_O[12] ,
    \Tile_X3Y13_FrameData_O[11] ,
    \Tile_X3Y13_FrameData_O[10] ,
    \Tile_X3Y13_FrameData_O[9] ,
    \Tile_X3Y13_FrameData_O[8] ,
    \Tile_X3Y13_FrameData_O[7] ,
    \Tile_X3Y13_FrameData_O[6] ,
    \Tile_X3Y13_FrameData_O[5] ,
    \Tile_X3Y13_FrameData_O[4] ,
    \Tile_X3Y13_FrameData_O[3] ,
    \Tile_X3Y13_FrameData_O[2] ,
    \Tile_X3Y13_FrameData_O[1] ,
    \Tile_X3Y13_FrameData_O[0] }),
    .FrameStrobe({\Tile_X3Y14_FrameStrobe_O[19] ,
    \Tile_X3Y14_FrameStrobe_O[18] ,
    \Tile_X3Y14_FrameStrobe_O[17] ,
    \Tile_X3Y14_FrameStrobe_O[16] ,
    \Tile_X3Y14_FrameStrobe_O[15] ,
    \Tile_X3Y14_FrameStrobe_O[14] ,
    \Tile_X3Y14_FrameStrobe_O[13] ,
    \Tile_X3Y14_FrameStrobe_O[12] ,
    \Tile_X3Y14_FrameStrobe_O[11] ,
    \Tile_X3Y14_FrameStrobe_O[10] ,
    \Tile_X3Y14_FrameStrobe_O[9] ,
    \Tile_X3Y14_FrameStrobe_O[8] ,
    \Tile_X3Y14_FrameStrobe_O[7] ,
    \Tile_X3Y14_FrameStrobe_O[6] ,
    \Tile_X3Y14_FrameStrobe_O[5] ,
    \Tile_X3Y14_FrameStrobe_O[4] ,
    \Tile_X3Y14_FrameStrobe_O[3] ,
    \Tile_X3Y14_FrameStrobe_O[2] ,
    \Tile_X3Y14_FrameStrobe_O[1] ,
    \Tile_X3Y14_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X3Y13_FrameStrobe_O[19] ,
    \Tile_X3Y13_FrameStrobe_O[18] ,
    \Tile_X3Y13_FrameStrobe_O[17] ,
    \Tile_X3Y13_FrameStrobe_O[16] ,
    \Tile_X3Y13_FrameStrobe_O[15] ,
    \Tile_X3Y13_FrameStrobe_O[14] ,
    \Tile_X3Y13_FrameStrobe_O[13] ,
    \Tile_X3Y13_FrameStrobe_O[12] ,
    \Tile_X3Y13_FrameStrobe_O[11] ,
    \Tile_X3Y13_FrameStrobe_O[10] ,
    \Tile_X3Y13_FrameStrobe_O[9] ,
    \Tile_X3Y13_FrameStrobe_O[8] ,
    \Tile_X3Y13_FrameStrobe_O[7] ,
    \Tile_X3Y13_FrameStrobe_O[6] ,
    \Tile_X3Y13_FrameStrobe_O[5] ,
    \Tile_X3Y13_FrameStrobe_O[4] ,
    \Tile_X3Y13_FrameStrobe_O[3] ,
    \Tile_X3Y13_FrameStrobe_O[2] ,
    \Tile_X3Y13_FrameStrobe_O[1] ,
    \Tile_X3Y13_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X3Y13_N1BEG[3] ,
    \Tile_X3Y13_N1BEG[2] ,
    \Tile_X3Y13_N1BEG[1] ,
    \Tile_X3Y13_N1BEG[0] }),
    .N1END({\Tile_X3Y14_N1BEG[3] ,
    \Tile_X3Y14_N1BEG[2] ,
    \Tile_X3Y14_N1BEG[1] ,
    \Tile_X3Y14_N1BEG[0] }),
    .N2BEG({\Tile_X3Y13_N2BEG[7] ,
    \Tile_X3Y13_N2BEG[6] ,
    \Tile_X3Y13_N2BEG[5] ,
    \Tile_X3Y13_N2BEG[4] ,
    \Tile_X3Y13_N2BEG[3] ,
    \Tile_X3Y13_N2BEG[2] ,
    \Tile_X3Y13_N2BEG[1] ,
    \Tile_X3Y13_N2BEG[0] }),
    .N2BEGb({\Tile_X3Y13_N2BEGb[7] ,
    \Tile_X3Y13_N2BEGb[6] ,
    \Tile_X3Y13_N2BEGb[5] ,
    \Tile_X3Y13_N2BEGb[4] ,
    \Tile_X3Y13_N2BEGb[3] ,
    \Tile_X3Y13_N2BEGb[2] ,
    \Tile_X3Y13_N2BEGb[1] ,
    \Tile_X3Y13_N2BEGb[0] }),
    .N2END({\Tile_X3Y14_N2BEGb[7] ,
    \Tile_X3Y14_N2BEGb[6] ,
    \Tile_X3Y14_N2BEGb[5] ,
    \Tile_X3Y14_N2BEGb[4] ,
    \Tile_X3Y14_N2BEGb[3] ,
    \Tile_X3Y14_N2BEGb[2] ,
    \Tile_X3Y14_N2BEGb[1] ,
    \Tile_X3Y14_N2BEGb[0] }),
    .N2MID({\Tile_X3Y14_N2BEG[7] ,
    \Tile_X3Y14_N2BEG[6] ,
    \Tile_X3Y14_N2BEG[5] ,
    \Tile_X3Y14_N2BEG[4] ,
    \Tile_X3Y14_N2BEG[3] ,
    \Tile_X3Y14_N2BEG[2] ,
    \Tile_X3Y14_N2BEG[1] ,
    \Tile_X3Y14_N2BEG[0] }),
    .N4BEG({\Tile_X3Y13_N4BEG[15] ,
    \Tile_X3Y13_N4BEG[14] ,
    \Tile_X3Y13_N4BEG[13] ,
    \Tile_X3Y13_N4BEG[12] ,
    \Tile_X3Y13_N4BEG[11] ,
    \Tile_X3Y13_N4BEG[10] ,
    \Tile_X3Y13_N4BEG[9] ,
    \Tile_X3Y13_N4BEG[8] ,
    \Tile_X3Y13_N4BEG[7] ,
    \Tile_X3Y13_N4BEG[6] ,
    \Tile_X3Y13_N4BEG[5] ,
    \Tile_X3Y13_N4BEG[4] ,
    \Tile_X3Y13_N4BEG[3] ,
    \Tile_X3Y13_N4BEG[2] ,
    \Tile_X3Y13_N4BEG[1] ,
    \Tile_X3Y13_N4BEG[0] }),
    .N4END({\Tile_X3Y14_N4BEG[15] ,
    \Tile_X3Y14_N4BEG[14] ,
    \Tile_X3Y14_N4BEG[13] ,
    \Tile_X3Y14_N4BEG[12] ,
    \Tile_X3Y14_N4BEG[11] ,
    \Tile_X3Y14_N4BEG[10] ,
    \Tile_X3Y14_N4BEG[9] ,
    \Tile_X3Y14_N4BEG[8] ,
    \Tile_X3Y14_N4BEG[7] ,
    \Tile_X3Y14_N4BEG[6] ,
    \Tile_X3Y14_N4BEG[5] ,
    \Tile_X3Y14_N4BEG[4] ,
    \Tile_X3Y14_N4BEG[3] ,
    \Tile_X3Y14_N4BEG[2] ,
    \Tile_X3Y14_N4BEG[1] ,
    \Tile_X3Y14_N4BEG[0] }),
    .NN4BEG({\Tile_X3Y13_NN4BEG[15] ,
    \Tile_X3Y13_NN4BEG[14] ,
    \Tile_X3Y13_NN4BEG[13] ,
    \Tile_X3Y13_NN4BEG[12] ,
    \Tile_X3Y13_NN4BEG[11] ,
    \Tile_X3Y13_NN4BEG[10] ,
    \Tile_X3Y13_NN4BEG[9] ,
    \Tile_X3Y13_NN4BEG[8] ,
    \Tile_X3Y13_NN4BEG[7] ,
    \Tile_X3Y13_NN4BEG[6] ,
    \Tile_X3Y13_NN4BEG[5] ,
    \Tile_X3Y13_NN4BEG[4] ,
    \Tile_X3Y13_NN4BEG[3] ,
    \Tile_X3Y13_NN4BEG[2] ,
    \Tile_X3Y13_NN4BEG[1] ,
    \Tile_X3Y13_NN4BEG[0] }),
    .NN4END({\Tile_X3Y14_NN4BEG[15] ,
    \Tile_X3Y14_NN4BEG[14] ,
    \Tile_X3Y14_NN4BEG[13] ,
    \Tile_X3Y14_NN4BEG[12] ,
    \Tile_X3Y14_NN4BEG[11] ,
    \Tile_X3Y14_NN4BEG[10] ,
    \Tile_X3Y14_NN4BEG[9] ,
    \Tile_X3Y14_NN4BEG[8] ,
    \Tile_X3Y14_NN4BEG[7] ,
    \Tile_X3Y14_NN4BEG[6] ,
    \Tile_X3Y14_NN4BEG[5] ,
    \Tile_X3Y14_NN4BEG[4] ,
    \Tile_X3Y14_NN4BEG[3] ,
    \Tile_X3Y14_NN4BEG[2] ,
    \Tile_X3Y14_NN4BEG[1] ,
    \Tile_X3Y14_NN4BEG[0] }),
    .S1BEG({\Tile_X3Y13_S1BEG[3] ,
    \Tile_X3Y13_S1BEG[2] ,
    \Tile_X3Y13_S1BEG[1] ,
    \Tile_X3Y13_S1BEG[0] }),
    .S1END({\Tile_X3Y12_S1BEG[3] ,
    \Tile_X3Y12_S1BEG[2] ,
    \Tile_X3Y12_S1BEG[1] ,
    \Tile_X3Y12_S1BEG[0] }),
    .S2BEG({\Tile_X3Y13_S2BEG[7] ,
    \Tile_X3Y13_S2BEG[6] ,
    \Tile_X3Y13_S2BEG[5] ,
    \Tile_X3Y13_S2BEG[4] ,
    \Tile_X3Y13_S2BEG[3] ,
    \Tile_X3Y13_S2BEG[2] ,
    \Tile_X3Y13_S2BEG[1] ,
    \Tile_X3Y13_S2BEG[0] }),
    .S2BEGb({\Tile_X3Y13_S2BEGb[7] ,
    \Tile_X3Y13_S2BEGb[6] ,
    \Tile_X3Y13_S2BEGb[5] ,
    \Tile_X3Y13_S2BEGb[4] ,
    \Tile_X3Y13_S2BEGb[3] ,
    \Tile_X3Y13_S2BEGb[2] ,
    \Tile_X3Y13_S2BEGb[1] ,
    \Tile_X3Y13_S2BEGb[0] }),
    .S2END({\Tile_X3Y12_S2BEGb[7] ,
    \Tile_X3Y12_S2BEGb[6] ,
    \Tile_X3Y12_S2BEGb[5] ,
    \Tile_X3Y12_S2BEGb[4] ,
    \Tile_X3Y12_S2BEGb[3] ,
    \Tile_X3Y12_S2BEGb[2] ,
    \Tile_X3Y12_S2BEGb[1] ,
    \Tile_X3Y12_S2BEGb[0] }),
    .S2MID({\Tile_X3Y12_S2BEG[7] ,
    \Tile_X3Y12_S2BEG[6] ,
    \Tile_X3Y12_S2BEG[5] ,
    \Tile_X3Y12_S2BEG[4] ,
    \Tile_X3Y12_S2BEG[3] ,
    \Tile_X3Y12_S2BEG[2] ,
    \Tile_X3Y12_S2BEG[1] ,
    \Tile_X3Y12_S2BEG[0] }),
    .S4BEG({\Tile_X3Y13_S4BEG[15] ,
    \Tile_X3Y13_S4BEG[14] ,
    \Tile_X3Y13_S4BEG[13] ,
    \Tile_X3Y13_S4BEG[12] ,
    \Tile_X3Y13_S4BEG[11] ,
    \Tile_X3Y13_S4BEG[10] ,
    \Tile_X3Y13_S4BEG[9] ,
    \Tile_X3Y13_S4BEG[8] ,
    \Tile_X3Y13_S4BEG[7] ,
    \Tile_X3Y13_S4BEG[6] ,
    \Tile_X3Y13_S4BEG[5] ,
    \Tile_X3Y13_S4BEG[4] ,
    \Tile_X3Y13_S4BEG[3] ,
    \Tile_X3Y13_S4BEG[2] ,
    \Tile_X3Y13_S4BEG[1] ,
    \Tile_X3Y13_S4BEG[0] }),
    .S4END({\Tile_X3Y12_S4BEG[15] ,
    \Tile_X3Y12_S4BEG[14] ,
    \Tile_X3Y12_S4BEG[13] ,
    \Tile_X3Y12_S4BEG[12] ,
    \Tile_X3Y12_S4BEG[11] ,
    \Tile_X3Y12_S4BEG[10] ,
    \Tile_X3Y12_S4BEG[9] ,
    \Tile_X3Y12_S4BEG[8] ,
    \Tile_X3Y12_S4BEG[7] ,
    \Tile_X3Y12_S4BEG[6] ,
    \Tile_X3Y12_S4BEG[5] ,
    \Tile_X3Y12_S4BEG[4] ,
    \Tile_X3Y12_S4BEG[3] ,
    \Tile_X3Y12_S4BEG[2] ,
    \Tile_X3Y12_S4BEG[1] ,
    \Tile_X3Y12_S4BEG[0] }),
    .SS4BEG({\Tile_X3Y13_SS4BEG[15] ,
    \Tile_X3Y13_SS4BEG[14] ,
    \Tile_X3Y13_SS4BEG[13] ,
    \Tile_X3Y13_SS4BEG[12] ,
    \Tile_X3Y13_SS4BEG[11] ,
    \Tile_X3Y13_SS4BEG[10] ,
    \Tile_X3Y13_SS4BEG[9] ,
    \Tile_X3Y13_SS4BEG[8] ,
    \Tile_X3Y13_SS4BEG[7] ,
    \Tile_X3Y13_SS4BEG[6] ,
    \Tile_X3Y13_SS4BEG[5] ,
    \Tile_X3Y13_SS4BEG[4] ,
    \Tile_X3Y13_SS4BEG[3] ,
    \Tile_X3Y13_SS4BEG[2] ,
    \Tile_X3Y13_SS4BEG[1] ,
    \Tile_X3Y13_SS4BEG[0] }),
    .SS4END({\Tile_X3Y12_SS4BEG[15] ,
    \Tile_X3Y12_SS4BEG[14] ,
    \Tile_X3Y12_SS4BEG[13] ,
    \Tile_X3Y12_SS4BEG[12] ,
    \Tile_X3Y12_SS4BEG[11] ,
    \Tile_X3Y12_SS4BEG[10] ,
    \Tile_X3Y12_SS4BEG[9] ,
    \Tile_X3Y12_SS4BEG[8] ,
    \Tile_X3Y12_SS4BEG[7] ,
    \Tile_X3Y12_SS4BEG[6] ,
    \Tile_X3Y12_SS4BEG[5] ,
    \Tile_X3Y12_SS4BEG[4] ,
    \Tile_X3Y12_SS4BEG[3] ,
    \Tile_X3Y12_SS4BEG[2] ,
    \Tile_X3Y12_SS4BEG[1] ,
    \Tile_X3Y12_SS4BEG[0] }),
    .W1BEG({\Tile_X3Y13_W1BEG[3] ,
    \Tile_X3Y13_W1BEG[2] ,
    \Tile_X3Y13_W1BEG[1] ,
    \Tile_X3Y13_W1BEG[0] }),
    .W1END({\Tile_X4Y13_W1BEG[3] ,
    \Tile_X4Y13_W1BEG[2] ,
    \Tile_X4Y13_W1BEG[1] ,
    \Tile_X4Y13_W1BEG[0] }),
    .W2BEG({\Tile_X3Y13_W2BEG[7] ,
    \Tile_X3Y13_W2BEG[6] ,
    \Tile_X3Y13_W2BEG[5] ,
    \Tile_X3Y13_W2BEG[4] ,
    \Tile_X3Y13_W2BEG[3] ,
    \Tile_X3Y13_W2BEG[2] ,
    \Tile_X3Y13_W2BEG[1] ,
    \Tile_X3Y13_W2BEG[0] }),
    .W2BEGb({\Tile_X3Y13_W2BEGb[7] ,
    \Tile_X3Y13_W2BEGb[6] ,
    \Tile_X3Y13_W2BEGb[5] ,
    \Tile_X3Y13_W2BEGb[4] ,
    \Tile_X3Y13_W2BEGb[3] ,
    \Tile_X3Y13_W2BEGb[2] ,
    \Tile_X3Y13_W2BEGb[1] ,
    \Tile_X3Y13_W2BEGb[0] }),
    .W2END({\Tile_X4Y13_W2BEGb[7] ,
    \Tile_X4Y13_W2BEGb[6] ,
    \Tile_X4Y13_W2BEGb[5] ,
    \Tile_X4Y13_W2BEGb[4] ,
    \Tile_X4Y13_W2BEGb[3] ,
    \Tile_X4Y13_W2BEGb[2] ,
    \Tile_X4Y13_W2BEGb[1] ,
    \Tile_X4Y13_W2BEGb[0] }),
    .W2MID({\Tile_X4Y13_W2BEG[7] ,
    \Tile_X4Y13_W2BEG[6] ,
    \Tile_X4Y13_W2BEG[5] ,
    \Tile_X4Y13_W2BEG[4] ,
    \Tile_X4Y13_W2BEG[3] ,
    \Tile_X4Y13_W2BEG[2] ,
    \Tile_X4Y13_W2BEG[1] ,
    \Tile_X4Y13_W2BEG[0] }),
    .W6BEG({\Tile_X3Y13_W6BEG[11] ,
    \Tile_X3Y13_W6BEG[10] ,
    \Tile_X3Y13_W6BEG[9] ,
    \Tile_X3Y13_W6BEG[8] ,
    \Tile_X3Y13_W6BEG[7] ,
    \Tile_X3Y13_W6BEG[6] ,
    \Tile_X3Y13_W6BEG[5] ,
    \Tile_X3Y13_W6BEG[4] ,
    \Tile_X3Y13_W6BEG[3] ,
    \Tile_X3Y13_W6BEG[2] ,
    \Tile_X3Y13_W6BEG[1] ,
    \Tile_X3Y13_W6BEG[0] }),
    .W6END({\Tile_X4Y13_W6BEG[11] ,
    \Tile_X4Y13_W6BEG[10] ,
    \Tile_X4Y13_W6BEG[9] ,
    \Tile_X4Y13_W6BEG[8] ,
    \Tile_X4Y13_W6BEG[7] ,
    \Tile_X4Y13_W6BEG[6] ,
    \Tile_X4Y13_W6BEG[5] ,
    \Tile_X4Y13_W6BEG[4] ,
    \Tile_X4Y13_W6BEG[3] ,
    \Tile_X4Y13_W6BEG[2] ,
    \Tile_X4Y13_W6BEG[1] ,
    \Tile_X4Y13_W6BEG[0] }),
    .WW4BEG({\Tile_X3Y13_WW4BEG[15] ,
    \Tile_X3Y13_WW4BEG[14] ,
    \Tile_X3Y13_WW4BEG[13] ,
    \Tile_X3Y13_WW4BEG[12] ,
    \Tile_X3Y13_WW4BEG[11] ,
    \Tile_X3Y13_WW4BEG[10] ,
    \Tile_X3Y13_WW4BEG[9] ,
    \Tile_X3Y13_WW4BEG[8] ,
    \Tile_X3Y13_WW4BEG[7] ,
    \Tile_X3Y13_WW4BEG[6] ,
    \Tile_X3Y13_WW4BEG[5] ,
    \Tile_X3Y13_WW4BEG[4] ,
    \Tile_X3Y13_WW4BEG[3] ,
    \Tile_X3Y13_WW4BEG[2] ,
    \Tile_X3Y13_WW4BEG[1] ,
    \Tile_X3Y13_WW4BEG[0] }),
    .WW4END({\Tile_X4Y13_WW4BEG[15] ,
    \Tile_X4Y13_WW4BEG[14] ,
    \Tile_X4Y13_WW4BEG[13] ,
    \Tile_X4Y13_WW4BEG[12] ,
    \Tile_X4Y13_WW4BEG[11] ,
    \Tile_X4Y13_WW4BEG[10] ,
    \Tile_X4Y13_WW4BEG[9] ,
    \Tile_X4Y13_WW4BEG[8] ,
    \Tile_X4Y13_WW4BEG[7] ,
    \Tile_X4Y13_WW4BEG[6] ,
    \Tile_X4Y13_WW4BEG[5] ,
    \Tile_X4Y13_WW4BEG[4] ,
    \Tile_X4Y13_WW4BEG[3] ,
    \Tile_X4Y13_WW4BEG[2] ,
    \Tile_X4Y13_WW4BEG[1] ,
    \Tile_X4Y13_WW4BEG[0] }));
 LUT4AB Tile_X3Y14_LUT4AB (.Ci(Tile_X3Y15_Co),
    .Co(Tile_X3Y14_Co),
    .UserCLK(Tile_X3Y15_UserCLKo),
    .UserCLKo(Tile_X3Y14_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X3Y14_E1BEG[3] ,
    \Tile_X3Y14_E1BEG[2] ,
    \Tile_X3Y14_E1BEG[1] ,
    \Tile_X3Y14_E1BEG[0] }),
    .E1END({\Tile_X2Y14_E1BEG[3] ,
    \Tile_X2Y14_E1BEG[2] ,
    \Tile_X2Y14_E1BEG[1] ,
    \Tile_X2Y14_E1BEG[0] }),
    .E2BEG({\Tile_X3Y14_E2BEG[7] ,
    \Tile_X3Y14_E2BEG[6] ,
    \Tile_X3Y14_E2BEG[5] ,
    \Tile_X3Y14_E2BEG[4] ,
    \Tile_X3Y14_E2BEG[3] ,
    \Tile_X3Y14_E2BEG[2] ,
    \Tile_X3Y14_E2BEG[1] ,
    \Tile_X3Y14_E2BEG[0] }),
    .E2BEGb({\Tile_X3Y14_E2BEGb[7] ,
    \Tile_X3Y14_E2BEGb[6] ,
    \Tile_X3Y14_E2BEGb[5] ,
    \Tile_X3Y14_E2BEGb[4] ,
    \Tile_X3Y14_E2BEGb[3] ,
    \Tile_X3Y14_E2BEGb[2] ,
    \Tile_X3Y14_E2BEGb[1] ,
    \Tile_X3Y14_E2BEGb[0] }),
    .E2END({\Tile_X2Y14_E2BEGb[7] ,
    \Tile_X2Y14_E2BEGb[6] ,
    \Tile_X2Y14_E2BEGb[5] ,
    \Tile_X2Y14_E2BEGb[4] ,
    \Tile_X2Y14_E2BEGb[3] ,
    \Tile_X2Y14_E2BEGb[2] ,
    \Tile_X2Y14_E2BEGb[1] ,
    \Tile_X2Y14_E2BEGb[0] }),
    .E2MID({\Tile_X2Y14_E2BEG[7] ,
    \Tile_X2Y14_E2BEG[6] ,
    \Tile_X2Y14_E2BEG[5] ,
    \Tile_X2Y14_E2BEG[4] ,
    \Tile_X2Y14_E2BEG[3] ,
    \Tile_X2Y14_E2BEG[2] ,
    \Tile_X2Y14_E2BEG[1] ,
    \Tile_X2Y14_E2BEG[0] }),
    .E6BEG({\Tile_X3Y14_E6BEG[11] ,
    \Tile_X3Y14_E6BEG[10] ,
    \Tile_X3Y14_E6BEG[9] ,
    \Tile_X3Y14_E6BEG[8] ,
    \Tile_X3Y14_E6BEG[7] ,
    \Tile_X3Y14_E6BEG[6] ,
    \Tile_X3Y14_E6BEG[5] ,
    \Tile_X3Y14_E6BEG[4] ,
    \Tile_X3Y14_E6BEG[3] ,
    \Tile_X3Y14_E6BEG[2] ,
    \Tile_X3Y14_E6BEG[1] ,
    \Tile_X3Y14_E6BEG[0] }),
    .E6END({\Tile_X2Y14_E6BEG[11] ,
    \Tile_X2Y14_E6BEG[10] ,
    \Tile_X2Y14_E6BEG[9] ,
    \Tile_X2Y14_E6BEG[8] ,
    \Tile_X2Y14_E6BEG[7] ,
    \Tile_X2Y14_E6BEG[6] ,
    \Tile_X2Y14_E6BEG[5] ,
    \Tile_X2Y14_E6BEG[4] ,
    \Tile_X2Y14_E6BEG[3] ,
    \Tile_X2Y14_E6BEG[2] ,
    \Tile_X2Y14_E6BEG[1] ,
    \Tile_X2Y14_E6BEG[0] }),
    .EE4BEG({\Tile_X3Y14_EE4BEG[15] ,
    \Tile_X3Y14_EE4BEG[14] ,
    \Tile_X3Y14_EE4BEG[13] ,
    \Tile_X3Y14_EE4BEG[12] ,
    \Tile_X3Y14_EE4BEG[11] ,
    \Tile_X3Y14_EE4BEG[10] ,
    \Tile_X3Y14_EE4BEG[9] ,
    \Tile_X3Y14_EE4BEG[8] ,
    \Tile_X3Y14_EE4BEG[7] ,
    \Tile_X3Y14_EE4BEG[6] ,
    \Tile_X3Y14_EE4BEG[5] ,
    \Tile_X3Y14_EE4BEG[4] ,
    \Tile_X3Y14_EE4BEG[3] ,
    \Tile_X3Y14_EE4BEG[2] ,
    \Tile_X3Y14_EE4BEG[1] ,
    \Tile_X3Y14_EE4BEG[0] }),
    .EE4END({\Tile_X2Y14_EE4BEG[15] ,
    \Tile_X2Y14_EE4BEG[14] ,
    \Tile_X2Y14_EE4BEG[13] ,
    \Tile_X2Y14_EE4BEG[12] ,
    \Tile_X2Y14_EE4BEG[11] ,
    \Tile_X2Y14_EE4BEG[10] ,
    \Tile_X2Y14_EE4BEG[9] ,
    \Tile_X2Y14_EE4BEG[8] ,
    \Tile_X2Y14_EE4BEG[7] ,
    \Tile_X2Y14_EE4BEG[6] ,
    \Tile_X2Y14_EE4BEG[5] ,
    \Tile_X2Y14_EE4BEG[4] ,
    \Tile_X2Y14_EE4BEG[3] ,
    \Tile_X2Y14_EE4BEG[2] ,
    \Tile_X2Y14_EE4BEG[1] ,
    \Tile_X2Y14_EE4BEG[0] }),
    .FrameData({\Tile_X2Y14_FrameData_O[31] ,
    \Tile_X2Y14_FrameData_O[30] ,
    \Tile_X2Y14_FrameData_O[29] ,
    \Tile_X2Y14_FrameData_O[28] ,
    \Tile_X2Y14_FrameData_O[27] ,
    \Tile_X2Y14_FrameData_O[26] ,
    \Tile_X2Y14_FrameData_O[25] ,
    \Tile_X2Y14_FrameData_O[24] ,
    \Tile_X2Y14_FrameData_O[23] ,
    \Tile_X2Y14_FrameData_O[22] ,
    \Tile_X2Y14_FrameData_O[21] ,
    \Tile_X2Y14_FrameData_O[20] ,
    \Tile_X2Y14_FrameData_O[19] ,
    \Tile_X2Y14_FrameData_O[18] ,
    \Tile_X2Y14_FrameData_O[17] ,
    \Tile_X2Y14_FrameData_O[16] ,
    \Tile_X2Y14_FrameData_O[15] ,
    \Tile_X2Y14_FrameData_O[14] ,
    \Tile_X2Y14_FrameData_O[13] ,
    \Tile_X2Y14_FrameData_O[12] ,
    \Tile_X2Y14_FrameData_O[11] ,
    \Tile_X2Y14_FrameData_O[10] ,
    \Tile_X2Y14_FrameData_O[9] ,
    \Tile_X2Y14_FrameData_O[8] ,
    \Tile_X2Y14_FrameData_O[7] ,
    \Tile_X2Y14_FrameData_O[6] ,
    \Tile_X2Y14_FrameData_O[5] ,
    \Tile_X2Y14_FrameData_O[4] ,
    \Tile_X2Y14_FrameData_O[3] ,
    \Tile_X2Y14_FrameData_O[2] ,
    \Tile_X2Y14_FrameData_O[1] ,
    \Tile_X2Y14_FrameData_O[0] }),
    .FrameData_O({\Tile_X3Y14_FrameData_O[31] ,
    \Tile_X3Y14_FrameData_O[30] ,
    \Tile_X3Y14_FrameData_O[29] ,
    \Tile_X3Y14_FrameData_O[28] ,
    \Tile_X3Y14_FrameData_O[27] ,
    \Tile_X3Y14_FrameData_O[26] ,
    \Tile_X3Y14_FrameData_O[25] ,
    \Tile_X3Y14_FrameData_O[24] ,
    \Tile_X3Y14_FrameData_O[23] ,
    \Tile_X3Y14_FrameData_O[22] ,
    \Tile_X3Y14_FrameData_O[21] ,
    \Tile_X3Y14_FrameData_O[20] ,
    \Tile_X3Y14_FrameData_O[19] ,
    \Tile_X3Y14_FrameData_O[18] ,
    \Tile_X3Y14_FrameData_O[17] ,
    \Tile_X3Y14_FrameData_O[16] ,
    \Tile_X3Y14_FrameData_O[15] ,
    \Tile_X3Y14_FrameData_O[14] ,
    \Tile_X3Y14_FrameData_O[13] ,
    \Tile_X3Y14_FrameData_O[12] ,
    \Tile_X3Y14_FrameData_O[11] ,
    \Tile_X3Y14_FrameData_O[10] ,
    \Tile_X3Y14_FrameData_O[9] ,
    \Tile_X3Y14_FrameData_O[8] ,
    \Tile_X3Y14_FrameData_O[7] ,
    \Tile_X3Y14_FrameData_O[6] ,
    \Tile_X3Y14_FrameData_O[5] ,
    \Tile_X3Y14_FrameData_O[4] ,
    \Tile_X3Y14_FrameData_O[3] ,
    \Tile_X3Y14_FrameData_O[2] ,
    \Tile_X3Y14_FrameData_O[1] ,
    \Tile_X3Y14_FrameData_O[0] }),
    .FrameStrobe({\Tile_X3Y15_FrameStrobe_O[19] ,
    \Tile_X3Y15_FrameStrobe_O[18] ,
    \Tile_X3Y15_FrameStrobe_O[17] ,
    \Tile_X3Y15_FrameStrobe_O[16] ,
    \Tile_X3Y15_FrameStrobe_O[15] ,
    \Tile_X3Y15_FrameStrobe_O[14] ,
    \Tile_X3Y15_FrameStrobe_O[13] ,
    \Tile_X3Y15_FrameStrobe_O[12] ,
    \Tile_X3Y15_FrameStrobe_O[11] ,
    \Tile_X3Y15_FrameStrobe_O[10] ,
    \Tile_X3Y15_FrameStrobe_O[9] ,
    \Tile_X3Y15_FrameStrobe_O[8] ,
    \Tile_X3Y15_FrameStrobe_O[7] ,
    \Tile_X3Y15_FrameStrobe_O[6] ,
    \Tile_X3Y15_FrameStrobe_O[5] ,
    \Tile_X3Y15_FrameStrobe_O[4] ,
    \Tile_X3Y15_FrameStrobe_O[3] ,
    \Tile_X3Y15_FrameStrobe_O[2] ,
    \Tile_X3Y15_FrameStrobe_O[1] ,
    \Tile_X3Y15_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X3Y14_FrameStrobe_O[19] ,
    \Tile_X3Y14_FrameStrobe_O[18] ,
    \Tile_X3Y14_FrameStrobe_O[17] ,
    \Tile_X3Y14_FrameStrobe_O[16] ,
    \Tile_X3Y14_FrameStrobe_O[15] ,
    \Tile_X3Y14_FrameStrobe_O[14] ,
    \Tile_X3Y14_FrameStrobe_O[13] ,
    \Tile_X3Y14_FrameStrobe_O[12] ,
    \Tile_X3Y14_FrameStrobe_O[11] ,
    \Tile_X3Y14_FrameStrobe_O[10] ,
    \Tile_X3Y14_FrameStrobe_O[9] ,
    \Tile_X3Y14_FrameStrobe_O[8] ,
    \Tile_X3Y14_FrameStrobe_O[7] ,
    \Tile_X3Y14_FrameStrobe_O[6] ,
    \Tile_X3Y14_FrameStrobe_O[5] ,
    \Tile_X3Y14_FrameStrobe_O[4] ,
    \Tile_X3Y14_FrameStrobe_O[3] ,
    \Tile_X3Y14_FrameStrobe_O[2] ,
    \Tile_X3Y14_FrameStrobe_O[1] ,
    \Tile_X3Y14_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X3Y14_N1BEG[3] ,
    \Tile_X3Y14_N1BEG[2] ,
    \Tile_X3Y14_N1BEG[1] ,
    \Tile_X3Y14_N1BEG[0] }),
    .N1END({\Tile_X3Y15_N1BEG[3] ,
    \Tile_X3Y15_N1BEG[2] ,
    \Tile_X3Y15_N1BEG[1] ,
    \Tile_X3Y15_N1BEG[0] }),
    .N2BEG({\Tile_X3Y14_N2BEG[7] ,
    \Tile_X3Y14_N2BEG[6] ,
    \Tile_X3Y14_N2BEG[5] ,
    \Tile_X3Y14_N2BEG[4] ,
    \Tile_X3Y14_N2BEG[3] ,
    \Tile_X3Y14_N2BEG[2] ,
    \Tile_X3Y14_N2BEG[1] ,
    \Tile_X3Y14_N2BEG[0] }),
    .N2BEGb({\Tile_X3Y14_N2BEGb[7] ,
    \Tile_X3Y14_N2BEGb[6] ,
    \Tile_X3Y14_N2BEGb[5] ,
    \Tile_X3Y14_N2BEGb[4] ,
    \Tile_X3Y14_N2BEGb[3] ,
    \Tile_X3Y14_N2BEGb[2] ,
    \Tile_X3Y14_N2BEGb[1] ,
    \Tile_X3Y14_N2BEGb[0] }),
    .N2END({\Tile_X3Y15_N2BEGb[7] ,
    \Tile_X3Y15_N2BEGb[6] ,
    \Tile_X3Y15_N2BEGb[5] ,
    \Tile_X3Y15_N2BEGb[4] ,
    \Tile_X3Y15_N2BEGb[3] ,
    \Tile_X3Y15_N2BEGb[2] ,
    \Tile_X3Y15_N2BEGb[1] ,
    \Tile_X3Y15_N2BEGb[0] }),
    .N2MID({\Tile_X3Y15_N2BEG[7] ,
    \Tile_X3Y15_N2BEG[6] ,
    \Tile_X3Y15_N2BEG[5] ,
    \Tile_X3Y15_N2BEG[4] ,
    \Tile_X3Y15_N2BEG[3] ,
    \Tile_X3Y15_N2BEG[2] ,
    \Tile_X3Y15_N2BEG[1] ,
    \Tile_X3Y15_N2BEG[0] }),
    .N4BEG({\Tile_X3Y14_N4BEG[15] ,
    \Tile_X3Y14_N4BEG[14] ,
    \Tile_X3Y14_N4BEG[13] ,
    \Tile_X3Y14_N4BEG[12] ,
    \Tile_X3Y14_N4BEG[11] ,
    \Tile_X3Y14_N4BEG[10] ,
    \Tile_X3Y14_N4BEG[9] ,
    \Tile_X3Y14_N4BEG[8] ,
    \Tile_X3Y14_N4BEG[7] ,
    \Tile_X3Y14_N4BEG[6] ,
    \Tile_X3Y14_N4BEG[5] ,
    \Tile_X3Y14_N4BEG[4] ,
    \Tile_X3Y14_N4BEG[3] ,
    \Tile_X3Y14_N4BEG[2] ,
    \Tile_X3Y14_N4BEG[1] ,
    \Tile_X3Y14_N4BEG[0] }),
    .N4END({\Tile_X3Y15_N4BEG[15] ,
    \Tile_X3Y15_N4BEG[14] ,
    \Tile_X3Y15_N4BEG[13] ,
    \Tile_X3Y15_N4BEG[12] ,
    \Tile_X3Y15_N4BEG[11] ,
    \Tile_X3Y15_N4BEG[10] ,
    \Tile_X3Y15_N4BEG[9] ,
    \Tile_X3Y15_N4BEG[8] ,
    \Tile_X3Y15_N4BEG[7] ,
    \Tile_X3Y15_N4BEG[6] ,
    \Tile_X3Y15_N4BEG[5] ,
    \Tile_X3Y15_N4BEG[4] ,
    \Tile_X3Y15_N4BEG[3] ,
    \Tile_X3Y15_N4BEG[2] ,
    \Tile_X3Y15_N4BEG[1] ,
    \Tile_X3Y15_N4BEG[0] }),
    .NN4BEG({\Tile_X3Y14_NN4BEG[15] ,
    \Tile_X3Y14_NN4BEG[14] ,
    \Tile_X3Y14_NN4BEG[13] ,
    \Tile_X3Y14_NN4BEG[12] ,
    \Tile_X3Y14_NN4BEG[11] ,
    \Tile_X3Y14_NN4BEG[10] ,
    \Tile_X3Y14_NN4BEG[9] ,
    \Tile_X3Y14_NN4BEG[8] ,
    \Tile_X3Y14_NN4BEG[7] ,
    \Tile_X3Y14_NN4BEG[6] ,
    \Tile_X3Y14_NN4BEG[5] ,
    \Tile_X3Y14_NN4BEG[4] ,
    \Tile_X3Y14_NN4BEG[3] ,
    \Tile_X3Y14_NN4BEG[2] ,
    \Tile_X3Y14_NN4BEG[1] ,
    \Tile_X3Y14_NN4BEG[0] }),
    .NN4END({\Tile_X3Y15_NN4BEG[15] ,
    \Tile_X3Y15_NN4BEG[14] ,
    \Tile_X3Y15_NN4BEG[13] ,
    \Tile_X3Y15_NN4BEG[12] ,
    \Tile_X3Y15_NN4BEG[11] ,
    \Tile_X3Y15_NN4BEG[10] ,
    \Tile_X3Y15_NN4BEG[9] ,
    \Tile_X3Y15_NN4BEG[8] ,
    \Tile_X3Y15_NN4BEG[7] ,
    \Tile_X3Y15_NN4BEG[6] ,
    \Tile_X3Y15_NN4BEG[5] ,
    \Tile_X3Y15_NN4BEG[4] ,
    \Tile_X3Y15_NN4BEG[3] ,
    \Tile_X3Y15_NN4BEG[2] ,
    \Tile_X3Y15_NN4BEG[1] ,
    \Tile_X3Y15_NN4BEG[0] }),
    .S1BEG({\Tile_X3Y14_S1BEG[3] ,
    \Tile_X3Y14_S1BEG[2] ,
    \Tile_X3Y14_S1BEG[1] ,
    \Tile_X3Y14_S1BEG[0] }),
    .S1END({\Tile_X3Y13_S1BEG[3] ,
    \Tile_X3Y13_S1BEG[2] ,
    \Tile_X3Y13_S1BEG[1] ,
    \Tile_X3Y13_S1BEG[0] }),
    .S2BEG({\Tile_X3Y14_S2BEG[7] ,
    \Tile_X3Y14_S2BEG[6] ,
    \Tile_X3Y14_S2BEG[5] ,
    \Tile_X3Y14_S2BEG[4] ,
    \Tile_X3Y14_S2BEG[3] ,
    \Tile_X3Y14_S2BEG[2] ,
    \Tile_X3Y14_S2BEG[1] ,
    \Tile_X3Y14_S2BEG[0] }),
    .S2BEGb({\Tile_X3Y14_S2BEGb[7] ,
    \Tile_X3Y14_S2BEGb[6] ,
    \Tile_X3Y14_S2BEGb[5] ,
    \Tile_X3Y14_S2BEGb[4] ,
    \Tile_X3Y14_S2BEGb[3] ,
    \Tile_X3Y14_S2BEGb[2] ,
    \Tile_X3Y14_S2BEGb[1] ,
    \Tile_X3Y14_S2BEGb[0] }),
    .S2END({\Tile_X3Y13_S2BEGb[7] ,
    \Tile_X3Y13_S2BEGb[6] ,
    \Tile_X3Y13_S2BEGb[5] ,
    \Tile_X3Y13_S2BEGb[4] ,
    \Tile_X3Y13_S2BEGb[3] ,
    \Tile_X3Y13_S2BEGb[2] ,
    \Tile_X3Y13_S2BEGb[1] ,
    \Tile_X3Y13_S2BEGb[0] }),
    .S2MID({\Tile_X3Y13_S2BEG[7] ,
    \Tile_X3Y13_S2BEG[6] ,
    \Tile_X3Y13_S2BEG[5] ,
    \Tile_X3Y13_S2BEG[4] ,
    \Tile_X3Y13_S2BEG[3] ,
    \Tile_X3Y13_S2BEG[2] ,
    \Tile_X3Y13_S2BEG[1] ,
    \Tile_X3Y13_S2BEG[0] }),
    .S4BEG({\Tile_X3Y14_S4BEG[15] ,
    \Tile_X3Y14_S4BEG[14] ,
    \Tile_X3Y14_S4BEG[13] ,
    \Tile_X3Y14_S4BEG[12] ,
    \Tile_X3Y14_S4BEG[11] ,
    \Tile_X3Y14_S4BEG[10] ,
    \Tile_X3Y14_S4BEG[9] ,
    \Tile_X3Y14_S4BEG[8] ,
    \Tile_X3Y14_S4BEG[7] ,
    \Tile_X3Y14_S4BEG[6] ,
    \Tile_X3Y14_S4BEG[5] ,
    \Tile_X3Y14_S4BEG[4] ,
    \Tile_X3Y14_S4BEG[3] ,
    \Tile_X3Y14_S4BEG[2] ,
    \Tile_X3Y14_S4BEG[1] ,
    \Tile_X3Y14_S4BEG[0] }),
    .S4END({\Tile_X3Y13_S4BEG[15] ,
    \Tile_X3Y13_S4BEG[14] ,
    \Tile_X3Y13_S4BEG[13] ,
    \Tile_X3Y13_S4BEG[12] ,
    \Tile_X3Y13_S4BEG[11] ,
    \Tile_X3Y13_S4BEG[10] ,
    \Tile_X3Y13_S4BEG[9] ,
    \Tile_X3Y13_S4BEG[8] ,
    \Tile_X3Y13_S4BEG[7] ,
    \Tile_X3Y13_S4BEG[6] ,
    \Tile_X3Y13_S4BEG[5] ,
    \Tile_X3Y13_S4BEG[4] ,
    \Tile_X3Y13_S4BEG[3] ,
    \Tile_X3Y13_S4BEG[2] ,
    \Tile_X3Y13_S4BEG[1] ,
    \Tile_X3Y13_S4BEG[0] }),
    .SS4BEG({\Tile_X3Y14_SS4BEG[15] ,
    \Tile_X3Y14_SS4BEG[14] ,
    \Tile_X3Y14_SS4BEG[13] ,
    \Tile_X3Y14_SS4BEG[12] ,
    \Tile_X3Y14_SS4BEG[11] ,
    \Tile_X3Y14_SS4BEG[10] ,
    \Tile_X3Y14_SS4BEG[9] ,
    \Tile_X3Y14_SS4BEG[8] ,
    \Tile_X3Y14_SS4BEG[7] ,
    \Tile_X3Y14_SS4BEG[6] ,
    \Tile_X3Y14_SS4BEG[5] ,
    \Tile_X3Y14_SS4BEG[4] ,
    \Tile_X3Y14_SS4BEG[3] ,
    \Tile_X3Y14_SS4BEG[2] ,
    \Tile_X3Y14_SS4BEG[1] ,
    \Tile_X3Y14_SS4BEG[0] }),
    .SS4END({\Tile_X3Y13_SS4BEG[15] ,
    \Tile_X3Y13_SS4BEG[14] ,
    \Tile_X3Y13_SS4BEG[13] ,
    \Tile_X3Y13_SS4BEG[12] ,
    \Tile_X3Y13_SS4BEG[11] ,
    \Tile_X3Y13_SS4BEG[10] ,
    \Tile_X3Y13_SS4BEG[9] ,
    \Tile_X3Y13_SS4BEG[8] ,
    \Tile_X3Y13_SS4BEG[7] ,
    \Tile_X3Y13_SS4BEG[6] ,
    \Tile_X3Y13_SS4BEG[5] ,
    \Tile_X3Y13_SS4BEG[4] ,
    \Tile_X3Y13_SS4BEG[3] ,
    \Tile_X3Y13_SS4BEG[2] ,
    \Tile_X3Y13_SS4BEG[1] ,
    \Tile_X3Y13_SS4BEG[0] }),
    .W1BEG({\Tile_X3Y14_W1BEG[3] ,
    \Tile_X3Y14_W1BEG[2] ,
    \Tile_X3Y14_W1BEG[1] ,
    \Tile_X3Y14_W1BEG[0] }),
    .W1END({\Tile_X4Y14_W1BEG[3] ,
    \Tile_X4Y14_W1BEG[2] ,
    \Tile_X4Y14_W1BEG[1] ,
    \Tile_X4Y14_W1BEG[0] }),
    .W2BEG({\Tile_X3Y14_W2BEG[7] ,
    \Tile_X3Y14_W2BEG[6] ,
    \Tile_X3Y14_W2BEG[5] ,
    \Tile_X3Y14_W2BEG[4] ,
    \Tile_X3Y14_W2BEG[3] ,
    \Tile_X3Y14_W2BEG[2] ,
    \Tile_X3Y14_W2BEG[1] ,
    \Tile_X3Y14_W2BEG[0] }),
    .W2BEGb({\Tile_X3Y14_W2BEGb[7] ,
    \Tile_X3Y14_W2BEGb[6] ,
    \Tile_X3Y14_W2BEGb[5] ,
    \Tile_X3Y14_W2BEGb[4] ,
    \Tile_X3Y14_W2BEGb[3] ,
    \Tile_X3Y14_W2BEGb[2] ,
    \Tile_X3Y14_W2BEGb[1] ,
    \Tile_X3Y14_W2BEGb[0] }),
    .W2END({\Tile_X4Y14_W2BEGb[7] ,
    \Tile_X4Y14_W2BEGb[6] ,
    \Tile_X4Y14_W2BEGb[5] ,
    \Tile_X4Y14_W2BEGb[4] ,
    \Tile_X4Y14_W2BEGb[3] ,
    \Tile_X4Y14_W2BEGb[2] ,
    \Tile_X4Y14_W2BEGb[1] ,
    \Tile_X4Y14_W2BEGb[0] }),
    .W2MID({\Tile_X4Y14_W2BEG[7] ,
    \Tile_X4Y14_W2BEG[6] ,
    \Tile_X4Y14_W2BEG[5] ,
    \Tile_X4Y14_W2BEG[4] ,
    \Tile_X4Y14_W2BEG[3] ,
    \Tile_X4Y14_W2BEG[2] ,
    \Tile_X4Y14_W2BEG[1] ,
    \Tile_X4Y14_W2BEG[0] }),
    .W6BEG({\Tile_X3Y14_W6BEG[11] ,
    \Tile_X3Y14_W6BEG[10] ,
    \Tile_X3Y14_W6BEG[9] ,
    \Tile_X3Y14_W6BEG[8] ,
    \Tile_X3Y14_W6BEG[7] ,
    \Tile_X3Y14_W6BEG[6] ,
    \Tile_X3Y14_W6BEG[5] ,
    \Tile_X3Y14_W6BEG[4] ,
    \Tile_X3Y14_W6BEG[3] ,
    \Tile_X3Y14_W6BEG[2] ,
    \Tile_X3Y14_W6BEG[1] ,
    \Tile_X3Y14_W6BEG[0] }),
    .W6END({\Tile_X4Y14_W6BEG[11] ,
    \Tile_X4Y14_W6BEG[10] ,
    \Tile_X4Y14_W6BEG[9] ,
    \Tile_X4Y14_W6BEG[8] ,
    \Tile_X4Y14_W6BEG[7] ,
    \Tile_X4Y14_W6BEG[6] ,
    \Tile_X4Y14_W6BEG[5] ,
    \Tile_X4Y14_W6BEG[4] ,
    \Tile_X4Y14_W6BEG[3] ,
    \Tile_X4Y14_W6BEG[2] ,
    \Tile_X4Y14_W6BEG[1] ,
    \Tile_X4Y14_W6BEG[0] }),
    .WW4BEG({\Tile_X3Y14_WW4BEG[15] ,
    \Tile_X3Y14_WW4BEG[14] ,
    \Tile_X3Y14_WW4BEG[13] ,
    \Tile_X3Y14_WW4BEG[12] ,
    \Tile_X3Y14_WW4BEG[11] ,
    \Tile_X3Y14_WW4BEG[10] ,
    \Tile_X3Y14_WW4BEG[9] ,
    \Tile_X3Y14_WW4BEG[8] ,
    \Tile_X3Y14_WW4BEG[7] ,
    \Tile_X3Y14_WW4BEG[6] ,
    \Tile_X3Y14_WW4BEG[5] ,
    \Tile_X3Y14_WW4BEG[4] ,
    \Tile_X3Y14_WW4BEG[3] ,
    \Tile_X3Y14_WW4BEG[2] ,
    \Tile_X3Y14_WW4BEG[1] ,
    \Tile_X3Y14_WW4BEG[0] }),
    .WW4END({\Tile_X4Y14_WW4BEG[15] ,
    \Tile_X4Y14_WW4BEG[14] ,
    \Tile_X4Y14_WW4BEG[13] ,
    \Tile_X4Y14_WW4BEG[12] ,
    \Tile_X4Y14_WW4BEG[11] ,
    \Tile_X4Y14_WW4BEG[10] ,
    \Tile_X4Y14_WW4BEG[9] ,
    \Tile_X4Y14_WW4BEG[8] ,
    \Tile_X4Y14_WW4BEG[7] ,
    \Tile_X4Y14_WW4BEG[6] ,
    \Tile_X4Y14_WW4BEG[5] ,
    \Tile_X4Y14_WW4BEG[4] ,
    \Tile_X4Y14_WW4BEG[3] ,
    \Tile_X4Y14_WW4BEG[2] ,
    \Tile_X4Y14_WW4BEG[1] ,
    \Tile_X4Y14_WW4BEG[0] }));
 S_CPU_IRQ Tile_X3Y15_S_CPU_IRQ (.CONFIGURED_top(Tile_X3Y15_CONFIGURED_top),
    .Co(Tile_X3Y15_Co),
    .IRQ_top0(Tile_X3Y15_IRQ_top0),
    .IRQ_top1(Tile_X3Y15_IRQ_top1),
    .IRQ_top2(Tile_X3Y15_IRQ_top2),
    .IRQ_top3(Tile_X3Y15_IRQ_top3),
    .UserCLK(UserCLK),
    .UserCLKo(Tile_X3Y15_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .FrameData({\Tile_X2Y15_FrameData_O[31] ,
    \Tile_X2Y15_FrameData_O[30] ,
    \Tile_X2Y15_FrameData_O[29] ,
    \Tile_X2Y15_FrameData_O[28] ,
    \Tile_X2Y15_FrameData_O[27] ,
    \Tile_X2Y15_FrameData_O[26] ,
    \Tile_X2Y15_FrameData_O[25] ,
    \Tile_X2Y15_FrameData_O[24] ,
    \Tile_X2Y15_FrameData_O[23] ,
    \Tile_X2Y15_FrameData_O[22] ,
    \Tile_X2Y15_FrameData_O[21] ,
    \Tile_X2Y15_FrameData_O[20] ,
    \Tile_X2Y15_FrameData_O[19] ,
    \Tile_X2Y15_FrameData_O[18] ,
    \Tile_X2Y15_FrameData_O[17] ,
    \Tile_X2Y15_FrameData_O[16] ,
    \Tile_X2Y15_FrameData_O[15] ,
    \Tile_X2Y15_FrameData_O[14] ,
    \Tile_X2Y15_FrameData_O[13] ,
    \Tile_X2Y15_FrameData_O[12] ,
    \Tile_X2Y15_FrameData_O[11] ,
    \Tile_X2Y15_FrameData_O[10] ,
    \Tile_X2Y15_FrameData_O[9] ,
    \Tile_X2Y15_FrameData_O[8] ,
    \Tile_X2Y15_FrameData_O[7] ,
    \Tile_X2Y15_FrameData_O[6] ,
    \Tile_X2Y15_FrameData_O[5] ,
    \Tile_X2Y15_FrameData_O[4] ,
    \Tile_X2Y15_FrameData_O[3] ,
    \Tile_X2Y15_FrameData_O[2] ,
    \Tile_X2Y15_FrameData_O[1] ,
    \Tile_X2Y15_FrameData_O[0] }),
    .FrameData_O({\Tile_X3Y15_FrameData_O[31] ,
    \Tile_X3Y15_FrameData_O[30] ,
    \Tile_X3Y15_FrameData_O[29] ,
    \Tile_X3Y15_FrameData_O[28] ,
    \Tile_X3Y15_FrameData_O[27] ,
    \Tile_X3Y15_FrameData_O[26] ,
    \Tile_X3Y15_FrameData_O[25] ,
    \Tile_X3Y15_FrameData_O[24] ,
    \Tile_X3Y15_FrameData_O[23] ,
    \Tile_X3Y15_FrameData_O[22] ,
    \Tile_X3Y15_FrameData_O[21] ,
    \Tile_X3Y15_FrameData_O[20] ,
    \Tile_X3Y15_FrameData_O[19] ,
    \Tile_X3Y15_FrameData_O[18] ,
    \Tile_X3Y15_FrameData_O[17] ,
    \Tile_X3Y15_FrameData_O[16] ,
    \Tile_X3Y15_FrameData_O[15] ,
    \Tile_X3Y15_FrameData_O[14] ,
    \Tile_X3Y15_FrameData_O[13] ,
    \Tile_X3Y15_FrameData_O[12] ,
    \Tile_X3Y15_FrameData_O[11] ,
    \Tile_X3Y15_FrameData_O[10] ,
    \Tile_X3Y15_FrameData_O[9] ,
    \Tile_X3Y15_FrameData_O[8] ,
    \Tile_X3Y15_FrameData_O[7] ,
    \Tile_X3Y15_FrameData_O[6] ,
    \Tile_X3Y15_FrameData_O[5] ,
    \Tile_X3Y15_FrameData_O[4] ,
    \Tile_X3Y15_FrameData_O[3] ,
    \Tile_X3Y15_FrameData_O[2] ,
    \Tile_X3Y15_FrameData_O[1] ,
    \Tile_X3Y15_FrameData_O[0] }),
    .FrameStrobe({FrameStrobe[79],
    FrameStrobe[78],
    FrameStrobe[77],
    FrameStrobe[76],
    FrameStrobe[75],
    FrameStrobe[74],
    FrameStrobe[73],
    FrameStrobe[72],
    FrameStrobe[71],
    FrameStrobe[70],
    FrameStrobe[69],
    FrameStrobe[68],
    FrameStrobe[67],
    FrameStrobe[66],
    FrameStrobe[65],
    FrameStrobe[64],
    FrameStrobe[63],
    FrameStrobe[62],
    FrameStrobe[61],
    FrameStrobe[60]}),
    .FrameStrobe_O({\Tile_X3Y15_FrameStrobe_O[19] ,
    \Tile_X3Y15_FrameStrobe_O[18] ,
    \Tile_X3Y15_FrameStrobe_O[17] ,
    \Tile_X3Y15_FrameStrobe_O[16] ,
    \Tile_X3Y15_FrameStrobe_O[15] ,
    \Tile_X3Y15_FrameStrobe_O[14] ,
    \Tile_X3Y15_FrameStrobe_O[13] ,
    \Tile_X3Y15_FrameStrobe_O[12] ,
    \Tile_X3Y15_FrameStrobe_O[11] ,
    \Tile_X3Y15_FrameStrobe_O[10] ,
    \Tile_X3Y15_FrameStrobe_O[9] ,
    \Tile_X3Y15_FrameStrobe_O[8] ,
    \Tile_X3Y15_FrameStrobe_O[7] ,
    \Tile_X3Y15_FrameStrobe_O[6] ,
    \Tile_X3Y15_FrameStrobe_O[5] ,
    \Tile_X3Y15_FrameStrobe_O[4] ,
    \Tile_X3Y15_FrameStrobe_O[3] ,
    \Tile_X3Y15_FrameStrobe_O[2] ,
    \Tile_X3Y15_FrameStrobe_O[1] ,
    \Tile_X3Y15_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X3Y15_N1BEG[3] ,
    \Tile_X3Y15_N1BEG[2] ,
    \Tile_X3Y15_N1BEG[1] ,
    \Tile_X3Y15_N1BEG[0] }),
    .N2BEG({\Tile_X3Y15_N2BEG[7] ,
    \Tile_X3Y15_N2BEG[6] ,
    \Tile_X3Y15_N2BEG[5] ,
    \Tile_X3Y15_N2BEG[4] ,
    \Tile_X3Y15_N2BEG[3] ,
    \Tile_X3Y15_N2BEG[2] ,
    \Tile_X3Y15_N2BEG[1] ,
    \Tile_X3Y15_N2BEG[0] }),
    .N2BEGb({\Tile_X3Y15_N2BEGb[7] ,
    \Tile_X3Y15_N2BEGb[6] ,
    \Tile_X3Y15_N2BEGb[5] ,
    \Tile_X3Y15_N2BEGb[4] ,
    \Tile_X3Y15_N2BEGb[3] ,
    \Tile_X3Y15_N2BEGb[2] ,
    \Tile_X3Y15_N2BEGb[1] ,
    \Tile_X3Y15_N2BEGb[0] }),
    .N4BEG({\Tile_X3Y15_N4BEG[15] ,
    \Tile_X3Y15_N4BEG[14] ,
    \Tile_X3Y15_N4BEG[13] ,
    \Tile_X3Y15_N4BEG[12] ,
    \Tile_X3Y15_N4BEG[11] ,
    \Tile_X3Y15_N4BEG[10] ,
    \Tile_X3Y15_N4BEG[9] ,
    \Tile_X3Y15_N4BEG[8] ,
    \Tile_X3Y15_N4BEG[7] ,
    \Tile_X3Y15_N4BEG[6] ,
    \Tile_X3Y15_N4BEG[5] ,
    \Tile_X3Y15_N4BEG[4] ,
    \Tile_X3Y15_N4BEG[3] ,
    \Tile_X3Y15_N4BEG[2] ,
    \Tile_X3Y15_N4BEG[1] ,
    \Tile_X3Y15_N4BEG[0] }),
    .NN4BEG({\Tile_X3Y15_NN4BEG[15] ,
    \Tile_X3Y15_NN4BEG[14] ,
    \Tile_X3Y15_NN4BEG[13] ,
    \Tile_X3Y15_NN4BEG[12] ,
    \Tile_X3Y15_NN4BEG[11] ,
    \Tile_X3Y15_NN4BEG[10] ,
    \Tile_X3Y15_NN4BEG[9] ,
    \Tile_X3Y15_NN4BEG[8] ,
    \Tile_X3Y15_NN4BEG[7] ,
    \Tile_X3Y15_NN4BEG[6] ,
    \Tile_X3Y15_NN4BEG[5] ,
    \Tile_X3Y15_NN4BEG[4] ,
    \Tile_X3Y15_NN4BEG[3] ,
    \Tile_X3Y15_NN4BEG[2] ,
    \Tile_X3Y15_NN4BEG[1] ,
    \Tile_X3Y15_NN4BEG[0] }),
    .S1END({\Tile_X3Y14_S1BEG[3] ,
    \Tile_X3Y14_S1BEG[2] ,
    \Tile_X3Y14_S1BEG[1] ,
    \Tile_X3Y14_S1BEG[0] }),
    .S2END({\Tile_X3Y14_S2BEGb[7] ,
    \Tile_X3Y14_S2BEGb[6] ,
    \Tile_X3Y14_S2BEGb[5] ,
    \Tile_X3Y14_S2BEGb[4] ,
    \Tile_X3Y14_S2BEGb[3] ,
    \Tile_X3Y14_S2BEGb[2] ,
    \Tile_X3Y14_S2BEGb[1] ,
    \Tile_X3Y14_S2BEGb[0] }),
    .S2MID({\Tile_X3Y14_S2BEG[7] ,
    \Tile_X3Y14_S2BEG[6] ,
    \Tile_X3Y14_S2BEG[5] ,
    \Tile_X3Y14_S2BEG[4] ,
    \Tile_X3Y14_S2BEG[3] ,
    \Tile_X3Y14_S2BEG[2] ,
    \Tile_X3Y14_S2BEG[1] ,
    \Tile_X3Y14_S2BEG[0] }),
    .S4END({\Tile_X3Y14_S4BEG[15] ,
    \Tile_X3Y14_S4BEG[14] ,
    \Tile_X3Y14_S4BEG[13] ,
    \Tile_X3Y14_S4BEG[12] ,
    \Tile_X3Y14_S4BEG[11] ,
    \Tile_X3Y14_S4BEG[10] ,
    \Tile_X3Y14_S4BEG[9] ,
    \Tile_X3Y14_S4BEG[8] ,
    \Tile_X3Y14_S4BEG[7] ,
    \Tile_X3Y14_S4BEG[6] ,
    \Tile_X3Y14_S4BEG[5] ,
    \Tile_X3Y14_S4BEG[4] ,
    \Tile_X3Y14_S4BEG[3] ,
    \Tile_X3Y14_S4BEG[2] ,
    \Tile_X3Y14_S4BEG[1] ,
    \Tile_X3Y14_S4BEG[0] }),
    .SS4END({\Tile_X3Y14_SS4BEG[15] ,
    \Tile_X3Y14_SS4BEG[14] ,
    \Tile_X3Y14_SS4BEG[13] ,
    \Tile_X3Y14_SS4BEG[12] ,
    \Tile_X3Y14_SS4BEG[11] ,
    \Tile_X3Y14_SS4BEG[10] ,
    \Tile_X3Y14_SS4BEG[9] ,
    \Tile_X3Y14_SS4BEG[8] ,
    \Tile_X3Y14_SS4BEG[7] ,
    \Tile_X3Y14_SS4BEG[6] ,
    \Tile_X3Y14_SS4BEG[5] ,
    \Tile_X3Y14_SS4BEG[4] ,
    \Tile_X3Y14_SS4BEG[3] ,
    \Tile_X3Y14_SS4BEG[2] ,
    \Tile_X3Y14_SS4BEG[1] ,
    \Tile_X3Y14_SS4BEG[0] }));
 LUT4AB Tile_X3Y1_LUT4AB (.Ci(Tile_X3Y2_Co),
    .Co(Tile_X3Y1_Co),
    .UserCLK(Tile_X3Y2_UserCLKo),
    .UserCLKo(Tile_X3Y1_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X3Y1_E1BEG[3] ,
    \Tile_X3Y1_E1BEG[2] ,
    \Tile_X3Y1_E1BEG[1] ,
    \Tile_X3Y1_E1BEG[0] }),
    .E1END({\Tile_X2Y1_E1BEG[3] ,
    \Tile_X2Y1_E1BEG[2] ,
    \Tile_X2Y1_E1BEG[1] ,
    \Tile_X2Y1_E1BEG[0] }),
    .E2BEG({\Tile_X3Y1_E2BEG[7] ,
    \Tile_X3Y1_E2BEG[6] ,
    \Tile_X3Y1_E2BEG[5] ,
    \Tile_X3Y1_E2BEG[4] ,
    \Tile_X3Y1_E2BEG[3] ,
    \Tile_X3Y1_E2BEG[2] ,
    \Tile_X3Y1_E2BEG[1] ,
    \Tile_X3Y1_E2BEG[0] }),
    .E2BEGb({\Tile_X3Y1_E2BEGb[7] ,
    \Tile_X3Y1_E2BEGb[6] ,
    \Tile_X3Y1_E2BEGb[5] ,
    \Tile_X3Y1_E2BEGb[4] ,
    \Tile_X3Y1_E2BEGb[3] ,
    \Tile_X3Y1_E2BEGb[2] ,
    \Tile_X3Y1_E2BEGb[1] ,
    \Tile_X3Y1_E2BEGb[0] }),
    .E2END({\Tile_X2Y1_E2BEGb[7] ,
    \Tile_X2Y1_E2BEGb[6] ,
    \Tile_X2Y1_E2BEGb[5] ,
    \Tile_X2Y1_E2BEGb[4] ,
    \Tile_X2Y1_E2BEGb[3] ,
    \Tile_X2Y1_E2BEGb[2] ,
    \Tile_X2Y1_E2BEGb[1] ,
    \Tile_X2Y1_E2BEGb[0] }),
    .E2MID({\Tile_X2Y1_E2BEG[7] ,
    \Tile_X2Y1_E2BEG[6] ,
    \Tile_X2Y1_E2BEG[5] ,
    \Tile_X2Y1_E2BEG[4] ,
    \Tile_X2Y1_E2BEG[3] ,
    \Tile_X2Y1_E2BEG[2] ,
    \Tile_X2Y1_E2BEG[1] ,
    \Tile_X2Y1_E2BEG[0] }),
    .E6BEG({\Tile_X3Y1_E6BEG[11] ,
    \Tile_X3Y1_E6BEG[10] ,
    \Tile_X3Y1_E6BEG[9] ,
    \Tile_X3Y1_E6BEG[8] ,
    \Tile_X3Y1_E6BEG[7] ,
    \Tile_X3Y1_E6BEG[6] ,
    \Tile_X3Y1_E6BEG[5] ,
    \Tile_X3Y1_E6BEG[4] ,
    \Tile_X3Y1_E6BEG[3] ,
    \Tile_X3Y1_E6BEG[2] ,
    \Tile_X3Y1_E6BEG[1] ,
    \Tile_X3Y1_E6BEG[0] }),
    .E6END({\Tile_X2Y1_E6BEG[11] ,
    \Tile_X2Y1_E6BEG[10] ,
    \Tile_X2Y1_E6BEG[9] ,
    \Tile_X2Y1_E6BEG[8] ,
    \Tile_X2Y1_E6BEG[7] ,
    \Tile_X2Y1_E6BEG[6] ,
    \Tile_X2Y1_E6BEG[5] ,
    \Tile_X2Y1_E6BEG[4] ,
    \Tile_X2Y1_E6BEG[3] ,
    \Tile_X2Y1_E6BEG[2] ,
    \Tile_X2Y1_E6BEG[1] ,
    \Tile_X2Y1_E6BEG[0] }),
    .EE4BEG({\Tile_X3Y1_EE4BEG[15] ,
    \Tile_X3Y1_EE4BEG[14] ,
    \Tile_X3Y1_EE4BEG[13] ,
    \Tile_X3Y1_EE4BEG[12] ,
    \Tile_X3Y1_EE4BEG[11] ,
    \Tile_X3Y1_EE4BEG[10] ,
    \Tile_X3Y1_EE4BEG[9] ,
    \Tile_X3Y1_EE4BEG[8] ,
    \Tile_X3Y1_EE4BEG[7] ,
    \Tile_X3Y1_EE4BEG[6] ,
    \Tile_X3Y1_EE4BEG[5] ,
    \Tile_X3Y1_EE4BEG[4] ,
    \Tile_X3Y1_EE4BEG[3] ,
    \Tile_X3Y1_EE4BEG[2] ,
    \Tile_X3Y1_EE4BEG[1] ,
    \Tile_X3Y1_EE4BEG[0] }),
    .EE4END({\Tile_X2Y1_EE4BEG[15] ,
    \Tile_X2Y1_EE4BEG[14] ,
    \Tile_X2Y1_EE4BEG[13] ,
    \Tile_X2Y1_EE4BEG[12] ,
    \Tile_X2Y1_EE4BEG[11] ,
    \Tile_X2Y1_EE4BEG[10] ,
    \Tile_X2Y1_EE4BEG[9] ,
    \Tile_X2Y1_EE4BEG[8] ,
    \Tile_X2Y1_EE4BEG[7] ,
    \Tile_X2Y1_EE4BEG[6] ,
    \Tile_X2Y1_EE4BEG[5] ,
    \Tile_X2Y1_EE4BEG[4] ,
    \Tile_X2Y1_EE4BEG[3] ,
    \Tile_X2Y1_EE4BEG[2] ,
    \Tile_X2Y1_EE4BEG[1] ,
    \Tile_X2Y1_EE4BEG[0] }),
    .FrameData({\Tile_X2Y1_FrameData_O[31] ,
    \Tile_X2Y1_FrameData_O[30] ,
    \Tile_X2Y1_FrameData_O[29] ,
    \Tile_X2Y1_FrameData_O[28] ,
    \Tile_X2Y1_FrameData_O[27] ,
    \Tile_X2Y1_FrameData_O[26] ,
    \Tile_X2Y1_FrameData_O[25] ,
    \Tile_X2Y1_FrameData_O[24] ,
    \Tile_X2Y1_FrameData_O[23] ,
    \Tile_X2Y1_FrameData_O[22] ,
    \Tile_X2Y1_FrameData_O[21] ,
    \Tile_X2Y1_FrameData_O[20] ,
    \Tile_X2Y1_FrameData_O[19] ,
    \Tile_X2Y1_FrameData_O[18] ,
    \Tile_X2Y1_FrameData_O[17] ,
    \Tile_X2Y1_FrameData_O[16] ,
    \Tile_X2Y1_FrameData_O[15] ,
    \Tile_X2Y1_FrameData_O[14] ,
    \Tile_X2Y1_FrameData_O[13] ,
    \Tile_X2Y1_FrameData_O[12] ,
    \Tile_X2Y1_FrameData_O[11] ,
    \Tile_X2Y1_FrameData_O[10] ,
    \Tile_X2Y1_FrameData_O[9] ,
    \Tile_X2Y1_FrameData_O[8] ,
    \Tile_X2Y1_FrameData_O[7] ,
    \Tile_X2Y1_FrameData_O[6] ,
    \Tile_X2Y1_FrameData_O[5] ,
    \Tile_X2Y1_FrameData_O[4] ,
    \Tile_X2Y1_FrameData_O[3] ,
    \Tile_X2Y1_FrameData_O[2] ,
    \Tile_X2Y1_FrameData_O[1] ,
    \Tile_X2Y1_FrameData_O[0] }),
    .FrameData_O({\Tile_X3Y1_FrameData_O[31] ,
    \Tile_X3Y1_FrameData_O[30] ,
    \Tile_X3Y1_FrameData_O[29] ,
    \Tile_X3Y1_FrameData_O[28] ,
    \Tile_X3Y1_FrameData_O[27] ,
    \Tile_X3Y1_FrameData_O[26] ,
    \Tile_X3Y1_FrameData_O[25] ,
    \Tile_X3Y1_FrameData_O[24] ,
    \Tile_X3Y1_FrameData_O[23] ,
    \Tile_X3Y1_FrameData_O[22] ,
    \Tile_X3Y1_FrameData_O[21] ,
    \Tile_X3Y1_FrameData_O[20] ,
    \Tile_X3Y1_FrameData_O[19] ,
    \Tile_X3Y1_FrameData_O[18] ,
    \Tile_X3Y1_FrameData_O[17] ,
    \Tile_X3Y1_FrameData_O[16] ,
    \Tile_X3Y1_FrameData_O[15] ,
    \Tile_X3Y1_FrameData_O[14] ,
    \Tile_X3Y1_FrameData_O[13] ,
    \Tile_X3Y1_FrameData_O[12] ,
    \Tile_X3Y1_FrameData_O[11] ,
    \Tile_X3Y1_FrameData_O[10] ,
    \Tile_X3Y1_FrameData_O[9] ,
    \Tile_X3Y1_FrameData_O[8] ,
    \Tile_X3Y1_FrameData_O[7] ,
    \Tile_X3Y1_FrameData_O[6] ,
    \Tile_X3Y1_FrameData_O[5] ,
    \Tile_X3Y1_FrameData_O[4] ,
    \Tile_X3Y1_FrameData_O[3] ,
    \Tile_X3Y1_FrameData_O[2] ,
    \Tile_X3Y1_FrameData_O[1] ,
    \Tile_X3Y1_FrameData_O[0] }),
    .FrameStrobe({\Tile_X3Y2_FrameStrobe_O[19] ,
    \Tile_X3Y2_FrameStrobe_O[18] ,
    \Tile_X3Y2_FrameStrobe_O[17] ,
    \Tile_X3Y2_FrameStrobe_O[16] ,
    \Tile_X3Y2_FrameStrobe_O[15] ,
    \Tile_X3Y2_FrameStrobe_O[14] ,
    \Tile_X3Y2_FrameStrobe_O[13] ,
    \Tile_X3Y2_FrameStrobe_O[12] ,
    \Tile_X3Y2_FrameStrobe_O[11] ,
    \Tile_X3Y2_FrameStrobe_O[10] ,
    \Tile_X3Y2_FrameStrobe_O[9] ,
    \Tile_X3Y2_FrameStrobe_O[8] ,
    \Tile_X3Y2_FrameStrobe_O[7] ,
    \Tile_X3Y2_FrameStrobe_O[6] ,
    \Tile_X3Y2_FrameStrobe_O[5] ,
    \Tile_X3Y2_FrameStrobe_O[4] ,
    \Tile_X3Y2_FrameStrobe_O[3] ,
    \Tile_X3Y2_FrameStrobe_O[2] ,
    \Tile_X3Y2_FrameStrobe_O[1] ,
    \Tile_X3Y2_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X3Y1_FrameStrobe_O[19] ,
    \Tile_X3Y1_FrameStrobe_O[18] ,
    \Tile_X3Y1_FrameStrobe_O[17] ,
    \Tile_X3Y1_FrameStrobe_O[16] ,
    \Tile_X3Y1_FrameStrobe_O[15] ,
    \Tile_X3Y1_FrameStrobe_O[14] ,
    \Tile_X3Y1_FrameStrobe_O[13] ,
    \Tile_X3Y1_FrameStrobe_O[12] ,
    \Tile_X3Y1_FrameStrobe_O[11] ,
    \Tile_X3Y1_FrameStrobe_O[10] ,
    \Tile_X3Y1_FrameStrobe_O[9] ,
    \Tile_X3Y1_FrameStrobe_O[8] ,
    \Tile_X3Y1_FrameStrobe_O[7] ,
    \Tile_X3Y1_FrameStrobe_O[6] ,
    \Tile_X3Y1_FrameStrobe_O[5] ,
    \Tile_X3Y1_FrameStrobe_O[4] ,
    \Tile_X3Y1_FrameStrobe_O[3] ,
    \Tile_X3Y1_FrameStrobe_O[2] ,
    \Tile_X3Y1_FrameStrobe_O[1] ,
    \Tile_X3Y1_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X3Y1_N1BEG[3] ,
    \Tile_X3Y1_N1BEG[2] ,
    \Tile_X3Y1_N1BEG[1] ,
    \Tile_X3Y1_N1BEG[0] }),
    .N1END({\Tile_X3Y2_N1BEG[3] ,
    \Tile_X3Y2_N1BEG[2] ,
    \Tile_X3Y2_N1BEG[1] ,
    \Tile_X3Y2_N1BEG[0] }),
    .N2BEG({\Tile_X3Y1_N2BEG[7] ,
    \Tile_X3Y1_N2BEG[6] ,
    \Tile_X3Y1_N2BEG[5] ,
    \Tile_X3Y1_N2BEG[4] ,
    \Tile_X3Y1_N2BEG[3] ,
    \Tile_X3Y1_N2BEG[2] ,
    \Tile_X3Y1_N2BEG[1] ,
    \Tile_X3Y1_N2BEG[0] }),
    .N2BEGb({\Tile_X3Y1_N2BEGb[7] ,
    \Tile_X3Y1_N2BEGb[6] ,
    \Tile_X3Y1_N2BEGb[5] ,
    \Tile_X3Y1_N2BEGb[4] ,
    \Tile_X3Y1_N2BEGb[3] ,
    \Tile_X3Y1_N2BEGb[2] ,
    \Tile_X3Y1_N2BEGb[1] ,
    \Tile_X3Y1_N2BEGb[0] }),
    .N2END({\Tile_X3Y2_N2BEGb[7] ,
    \Tile_X3Y2_N2BEGb[6] ,
    \Tile_X3Y2_N2BEGb[5] ,
    \Tile_X3Y2_N2BEGb[4] ,
    \Tile_X3Y2_N2BEGb[3] ,
    \Tile_X3Y2_N2BEGb[2] ,
    \Tile_X3Y2_N2BEGb[1] ,
    \Tile_X3Y2_N2BEGb[0] }),
    .N2MID({\Tile_X3Y2_N2BEG[7] ,
    \Tile_X3Y2_N2BEG[6] ,
    \Tile_X3Y2_N2BEG[5] ,
    \Tile_X3Y2_N2BEG[4] ,
    \Tile_X3Y2_N2BEG[3] ,
    \Tile_X3Y2_N2BEG[2] ,
    \Tile_X3Y2_N2BEG[1] ,
    \Tile_X3Y2_N2BEG[0] }),
    .N4BEG({\Tile_X3Y1_N4BEG[15] ,
    \Tile_X3Y1_N4BEG[14] ,
    \Tile_X3Y1_N4BEG[13] ,
    \Tile_X3Y1_N4BEG[12] ,
    \Tile_X3Y1_N4BEG[11] ,
    \Tile_X3Y1_N4BEG[10] ,
    \Tile_X3Y1_N4BEG[9] ,
    \Tile_X3Y1_N4BEG[8] ,
    \Tile_X3Y1_N4BEG[7] ,
    \Tile_X3Y1_N4BEG[6] ,
    \Tile_X3Y1_N4BEG[5] ,
    \Tile_X3Y1_N4BEG[4] ,
    \Tile_X3Y1_N4BEG[3] ,
    \Tile_X3Y1_N4BEG[2] ,
    \Tile_X3Y1_N4BEG[1] ,
    \Tile_X3Y1_N4BEG[0] }),
    .N4END({\Tile_X3Y2_N4BEG[15] ,
    \Tile_X3Y2_N4BEG[14] ,
    \Tile_X3Y2_N4BEG[13] ,
    \Tile_X3Y2_N4BEG[12] ,
    \Tile_X3Y2_N4BEG[11] ,
    \Tile_X3Y2_N4BEG[10] ,
    \Tile_X3Y2_N4BEG[9] ,
    \Tile_X3Y2_N4BEG[8] ,
    \Tile_X3Y2_N4BEG[7] ,
    \Tile_X3Y2_N4BEG[6] ,
    \Tile_X3Y2_N4BEG[5] ,
    \Tile_X3Y2_N4BEG[4] ,
    \Tile_X3Y2_N4BEG[3] ,
    \Tile_X3Y2_N4BEG[2] ,
    \Tile_X3Y2_N4BEG[1] ,
    \Tile_X3Y2_N4BEG[0] }),
    .NN4BEG({\Tile_X3Y1_NN4BEG[15] ,
    \Tile_X3Y1_NN4BEG[14] ,
    \Tile_X3Y1_NN4BEG[13] ,
    \Tile_X3Y1_NN4BEG[12] ,
    \Tile_X3Y1_NN4BEG[11] ,
    \Tile_X3Y1_NN4BEG[10] ,
    \Tile_X3Y1_NN4BEG[9] ,
    \Tile_X3Y1_NN4BEG[8] ,
    \Tile_X3Y1_NN4BEG[7] ,
    \Tile_X3Y1_NN4BEG[6] ,
    \Tile_X3Y1_NN4BEG[5] ,
    \Tile_X3Y1_NN4BEG[4] ,
    \Tile_X3Y1_NN4BEG[3] ,
    \Tile_X3Y1_NN4BEG[2] ,
    \Tile_X3Y1_NN4BEG[1] ,
    \Tile_X3Y1_NN4BEG[0] }),
    .NN4END({\Tile_X3Y2_NN4BEG[15] ,
    \Tile_X3Y2_NN4BEG[14] ,
    \Tile_X3Y2_NN4BEG[13] ,
    \Tile_X3Y2_NN4BEG[12] ,
    \Tile_X3Y2_NN4BEG[11] ,
    \Tile_X3Y2_NN4BEG[10] ,
    \Tile_X3Y2_NN4BEG[9] ,
    \Tile_X3Y2_NN4BEG[8] ,
    \Tile_X3Y2_NN4BEG[7] ,
    \Tile_X3Y2_NN4BEG[6] ,
    \Tile_X3Y2_NN4BEG[5] ,
    \Tile_X3Y2_NN4BEG[4] ,
    \Tile_X3Y2_NN4BEG[3] ,
    \Tile_X3Y2_NN4BEG[2] ,
    \Tile_X3Y2_NN4BEG[1] ,
    \Tile_X3Y2_NN4BEG[0] }),
    .S1BEG({\Tile_X3Y1_S1BEG[3] ,
    \Tile_X3Y1_S1BEG[2] ,
    \Tile_X3Y1_S1BEG[1] ,
    \Tile_X3Y1_S1BEG[0] }),
    .S1END({\Tile_X3Y0_S1BEG[3] ,
    \Tile_X3Y0_S1BEG[2] ,
    \Tile_X3Y0_S1BEG[1] ,
    \Tile_X3Y0_S1BEG[0] }),
    .S2BEG({\Tile_X3Y1_S2BEG[7] ,
    \Tile_X3Y1_S2BEG[6] ,
    \Tile_X3Y1_S2BEG[5] ,
    \Tile_X3Y1_S2BEG[4] ,
    \Tile_X3Y1_S2BEG[3] ,
    \Tile_X3Y1_S2BEG[2] ,
    \Tile_X3Y1_S2BEG[1] ,
    \Tile_X3Y1_S2BEG[0] }),
    .S2BEGb({\Tile_X3Y1_S2BEGb[7] ,
    \Tile_X3Y1_S2BEGb[6] ,
    \Tile_X3Y1_S2BEGb[5] ,
    \Tile_X3Y1_S2BEGb[4] ,
    \Tile_X3Y1_S2BEGb[3] ,
    \Tile_X3Y1_S2BEGb[2] ,
    \Tile_X3Y1_S2BEGb[1] ,
    \Tile_X3Y1_S2BEGb[0] }),
    .S2END({\Tile_X3Y0_S2BEGb[7] ,
    \Tile_X3Y0_S2BEGb[6] ,
    \Tile_X3Y0_S2BEGb[5] ,
    \Tile_X3Y0_S2BEGb[4] ,
    \Tile_X3Y0_S2BEGb[3] ,
    \Tile_X3Y0_S2BEGb[2] ,
    \Tile_X3Y0_S2BEGb[1] ,
    \Tile_X3Y0_S2BEGb[0] }),
    .S2MID({\Tile_X3Y0_S2BEG[7] ,
    \Tile_X3Y0_S2BEG[6] ,
    \Tile_X3Y0_S2BEG[5] ,
    \Tile_X3Y0_S2BEG[4] ,
    \Tile_X3Y0_S2BEG[3] ,
    \Tile_X3Y0_S2BEG[2] ,
    \Tile_X3Y0_S2BEG[1] ,
    \Tile_X3Y0_S2BEG[0] }),
    .S4BEG({\Tile_X3Y1_S4BEG[15] ,
    \Tile_X3Y1_S4BEG[14] ,
    \Tile_X3Y1_S4BEG[13] ,
    \Tile_X3Y1_S4BEG[12] ,
    \Tile_X3Y1_S4BEG[11] ,
    \Tile_X3Y1_S4BEG[10] ,
    \Tile_X3Y1_S4BEG[9] ,
    \Tile_X3Y1_S4BEG[8] ,
    \Tile_X3Y1_S4BEG[7] ,
    \Tile_X3Y1_S4BEG[6] ,
    \Tile_X3Y1_S4BEG[5] ,
    \Tile_X3Y1_S4BEG[4] ,
    \Tile_X3Y1_S4BEG[3] ,
    \Tile_X3Y1_S4BEG[2] ,
    \Tile_X3Y1_S4BEG[1] ,
    \Tile_X3Y1_S4BEG[0] }),
    .S4END({\Tile_X3Y0_S4BEG[15] ,
    \Tile_X3Y0_S4BEG[14] ,
    \Tile_X3Y0_S4BEG[13] ,
    \Tile_X3Y0_S4BEG[12] ,
    \Tile_X3Y0_S4BEG[11] ,
    \Tile_X3Y0_S4BEG[10] ,
    \Tile_X3Y0_S4BEG[9] ,
    \Tile_X3Y0_S4BEG[8] ,
    \Tile_X3Y0_S4BEG[7] ,
    \Tile_X3Y0_S4BEG[6] ,
    \Tile_X3Y0_S4BEG[5] ,
    \Tile_X3Y0_S4BEG[4] ,
    \Tile_X3Y0_S4BEG[3] ,
    \Tile_X3Y0_S4BEG[2] ,
    \Tile_X3Y0_S4BEG[1] ,
    \Tile_X3Y0_S4BEG[0] }),
    .SS4BEG({\Tile_X3Y1_SS4BEG[15] ,
    \Tile_X3Y1_SS4BEG[14] ,
    \Tile_X3Y1_SS4BEG[13] ,
    \Tile_X3Y1_SS4BEG[12] ,
    \Tile_X3Y1_SS4BEG[11] ,
    \Tile_X3Y1_SS4BEG[10] ,
    \Tile_X3Y1_SS4BEG[9] ,
    \Tile_X3Y1_SS4BEG[8] ,
    \Tile_X3Y1_SS4BEG[7] ,
    \Tile_X3Y1_SS4BEG[6] ,
    \Tile_X3Y1_SS4BEG[5] ,
    \Tile_X3Y1_SS4BEG[4] ,
    \Tile_X3Y1_SS4BEG[3] ,
    \Tile_X3Y1_SS4BEG[2] ,
    \Tile_X3Y1_SS4BEG[1] ,
    \Tile_X3Y1_SS4BEG[0] }),
    .SS4END({\Tile_X3Y0_SS4BEG[15] ,
    \Tile_X3Y0_SS4BEG[14] ,
    \Tile_X3Y0_SS4BEG[13] ,
    \Tile_X3Y0_SS4BEG[12] ,
    \Tile_X3Y0_SS4BEG[11] ,
    \Tile_X3Y0_SS4BEG[10] ,
    \Tile_X3Y0_SS4BEG[9] ,
    \Tile_X3Y0_SS4BEG[8] ,
    \Tile_X3Y0_SS4BEG[7] ,
    \Tile_X3Y0_SS4BEG[6] ,
    \Tile_X3Y0_SS4BEG[5] ,
    \Tile_X3Y0_SS4BEG[4] ,
    \Tile_X3Y0_SS4BEG[3] ,
    \Tile_X3Y0_SS4BEG[2] ,
    \Tile_X3Y0_SS4BEG[1] ,
    \Tile_X3Y0_SS4BEG[0] }),
    .W1BEG({\Tile_X3Y1_W1BEG[3] ,
    \Tile_X3Y1_W1BEG[2] ,
    \Tile_X3Y1_W1BEG[1] ,
    \Tile_X3Y1_W1BEG[0] }),
    .W1END({\Tile_X4Y1_W1BEG[3] ,
    \Tile_X4Y1_W1BEG[2] ,
    \Tile_X4Y1_W1BEG[1] ,
    \Tile_X4Y1_W1BEG[0] }),
    .W2BEG({\Tile_X3Y1_W2BEG[7] ,
    \Tile_X3Y1_W2BEG[6] ,
    \Tile_X3Y1_W2BEG[5] ,
    \Tile_X3Y1_W2BEG[4] ,
    \Tile_X3Y1_W2BEG[3] ,
    \Tile_X3Y1_W2BEG[2] ,
    \Tile_X3Y1_W2BEG[1] ,
    \Tile_X3Y1_W2BEG[0] }),
    .W2BEGb({\Tile_X3Y1_W2BEGb[7] ,
    \Tile_X3Y1_W2BEGb[6] ,
    \Tile_X3Y1_W2BEGb[5] ,
    \Tile_X3Y1_W2BEGb[4] ,
    \Tile_X3Y1_W2BEGb[3] ,
    \Tile_X3Y1_W2BEGb[2] ,
    \Tile_X3Y1_W2BEGb[1] ,
    \Tile_X3Y1_W2BEGb[0] }),
    .W2END({\Tile_X4Y1_W2BEGb[7] ,
    \Tile_X4Y1_W2BEGb[6] ,
    \Tile_X4Y1_W2BEGb[5] ,
    \Tile_X4Y1_W2BEGb[4] ,
    \Tile_X4Y1_W2BEGb[3] ,
    \Tile_X4Y1_W2BEGb[2] ,
    \Tile_X4Y1_W2BEGb[1] ,
    \Tile_X4Y1_W2BEGb[0] }),
    .W2MID({\Tile_X4Y1_W2BEG[7] ,
    \Tile_X4Y1_W2BEG[6] ,
    \Tile_X4Y1_W2BEG[5] ,
    \Tile_X4Y1_W2BEG[4] ,
    \Tile_X4Y1_W2BEG[3] ,
    \Tile_X4Y1_W2BEG[2] ,
    \Tile_X4Y1_W2BEG[1] ,
    \Tile_X4Y1_W2BEG[0] }),
    .W6BEG({\Tile_X3Y1_W6BEG[11] ,
    \Tile_X3Y1_W6BEG[10] ,
    \Tile_X3Y1_W6BEG[9] ,
    \Tile_X3Y1_W6BEG[8] ,
    \Tile_X3Y1_W6BEG[7] ,
    \Tile_X3Y1_W6BEG[6] ,
    \Tile_X3Y1_W6BEG[5] ,
    \Tile_X3Y1_W6BEG[4] ,
    \Tile_X3Y1_W6BEG[3] ,
    \Tile_X3Y1_W6BEG[2] ,
    \Tile_X3Y1_W6BEG[1] ,
    \Tile_X3Y1_W6BEG[0] }),
    .W6END({\Tile_X4Y1_W6BEG[11] ,
    \Tile_X4Y1_W6BEG[10] ,
    \Tile_X4Y1_W6BEG[9] ,
    \Tile_X4Y1_W6BEG[8] ,
    \Tile_X4Y1_W6BEG[7] ,
    \Tile_X4Y1_W6BEG[6] ,
    \Tile_X4Y1_W6BEG[5] ,
    \Tile_X4Y1_W6BEG[4] ,
    \Tile_X4Y1_W6BEG[3] ,
    \Tile_X4Y1_W6BEG[2] ,
    \Tile_X4Y1_W6BEG[1] ,
    \Tile_X4Y1_W6BEG[0] }),
    .WW4BEG({\Tile_X3Y1_WW4BEG[15] ,
    \Tile_X3Y1_WW4BEG[14] ,
    \Tile_X3Y1_WW4BEG[13] ,
    \Tile_X3Y1_WW4BEG[12] ,
    \Tile_X3Y1_WW4BEG[11] ,
    \Tile_X3Y1_WW4BEG[10] ,
    \Tile_X3Y1_WW4BEG[9] ,
    \Tile_X3Y1_WW4BEG[8] ,
    \Tile_X3Y1_WW4BEG[7] ,
    \Tile_X3Y1_WW4BEG[6] ,
    \Tile_X3Y1_WW4BEG[5] ,
    \Tile_X3Y1_WW4BEG[4] ,
    \Tile_X3Y1_WW4BEG[3] ,
    \Tile_X3Y1_WW4BEG[2] ,
    \Tile_X3Y1_WW4BEG[1] ,
    \Tile_X3Y1_WW4BEG[0] }),
    .WW4END({\Tile_X4Y1_WW4BEG[15] ,
    \Tile_X4Y1_WW4BEG[14] ,
    \Tile_X4Y1_WW4BEG[13] ,
    \Tile_X4Y1_WW4BEG[12] ,
    \Tile_X4Y1_WW4BEG[11] ,
    \Tile_X4Y1_WW4BEG[10] ,
    \Tile_X4Y1_WW4BEG[9] ,
    \Tile_X4Y1_WW4BEG[8] ,
    \Tile_X4Y1_WW4BEG[7] ,
    \Tile_X4Y1_WW4BEG[6] ,
    \Tile_X4Y1_WW4BEG[5] ,
    \Tile_X4Y1_WW4BEG[4] ,
    \Tile_X4Y1_WW4BEG[3] ,
    \Tile_X4Y1_WW4BEG[2] ,
    \Tile_X4Y1_WW4BEG[1] ,
    \Tile_X4Y1_WW4BEG[0] }));
 LUT4AB Tile_X3Y2_LUT4AB (.Ci(Tile_X3Y3_Co),
    .Co(Tile_X3Y2_Co),
    .UserCLK(Tile_X3Y3_UserCLKo),
    .UserCLKo(Tile_X3Y2_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X3Y2_E1BEG[3] ,
    \Tile_X3Y2_E1BEG[2] ,
    \Tile_X3Y2_E1BEG[1] ,
    \Tile_X3Y2_E1BEG[0] }),
    .E1END({\Tile_X2Y2_E1BEG[3] ,
    \Tile_X2Y2_E1BEG[2] ,
    \Tile_X2Y2_E1BEG[1] ,
    \Tile_X2Y2_E1BEG[0] }),
    .E2BEG({\Tile_X3Y2_E2BEG[7] ,
    \Tile_X3Y2_E2BEG[6] ,
    \Tile_X3Y2_E2BEG[5] ,
    \Tile_X3Y2_E2BEG[4] ,
    \Tile_X3Y2_E2BEG[3] ,
    \Tile_X3Y2_E2BEG[2] ,
    \Tile_X3Y2_E2BEG[1] ,
    \Tile_X3Y2_E2BEG[0] }),
    .E2BEGb({\Tile_X3Y2_E2BEGb[7] ,
    \Tile_X3Y2_E2BEGb[6] ,
    \Tile_X3Y2_E2BEGb[5] ,
    \Tile_X3Y2_E2BEGb[4] ,
    \Tile_X3Y2_E2BEGb[3] ,
    \Tile_X3Y2_E2BEGb[2] ,
    \Tile_X3Y2_E2BEGb[1] ,
    \Tile_X3Y2_E2BEGb[0] }),
    .E2END({\Tile_X2Y2_E2BEGb[7] ,
    \Tile_X2Y2_E2BEGb[6] ,
    \Tile_X2Y2_E2BEGb[5] ,
    \Tile_X2Y2_E2BEGb[4] ,
    \Tile_X2Y2_E2BEGb[3] ,
    \Tile_X2Y2_E2BEGb[2] ,
    \Tile_X2Y2_E2BEGb[1] ,
    \Tile_X2Y2_E2BEGb[0] }),
    .E2MID({\Tile_X2Y2_E2BEG[7] ,
    \Tile_X2Y2_E2BEG[6] ,
    \Tile_X2Y2_E2BEG[5] ,
    \Tile_X2Y2_E2BEG[4] ,
    \Tile_X2Y2_E2BEG[3] ,
    \Tile_X2Y2_E2BEG[2] ,
    \Tile_X2Y2_E2BEG[1] ,
    \Tile_X2Y2_E2BEG[0] }),
    .E6BEG({\Tile_X3Y2_E6BEG[11] ,
    \Tile_X3Y2_E6BEG[10] ,
    \Tile_X3Y2_E6BEG[9] ,
    \Tile_X3Y2_E6BEG[8] ,
    \Tile_X3Y2_E6BEG[7] ,
    \Tile_X3Y2_E6BEG[6] ,
    \Tile_X3Y2_E6BEG[5] ,
    \Tile_X3Y2_E6BEG[4] ,
    \Tile_X3Y2_E6BEG[3] ,
    \Tile_X3Y2_E6BEG[2] ,
    \Tile_X3Y2_E6BEG[1] ,
    \Tile_X3Y2_E6BEG[0] }),
    .E6END({\Tile_X2Y2_E6BEG[11] ,
    \Tile_X2Y2_E6BEG[10] ,
    \Tile_X2Y2_E6BEG[9] ,
    \Tile_X2Y2_E6BEG[8] ,
    \Tile_X2Y2_E6BEG[7] ,
    \Tile_X2Y2_E6BEG[6] ,
    \Tile_X2Y2_E6BEG[5] ,
    \Tile_X2Y2_E6BEG[4] ,
    \Tile_X2Y2_E6BEG[3] ,
    \Tile_X2Y2_E6BEG[2] ,
    \Tile_X2Y2_E6BEG[1] ,
    \Tile_X2Y2_E6BEG[0] }),
    .EE4BEG({\Tile_X3Y2_EE4BEG[15] ,
    \Tile_X3Y2_EE4BEG[14] ,
    \Tile_X3Y2_EE4BEG[13] ,
    \Tile_X3Y2_EE4BEG[12] ,
    \Tile_X3Y2_EE4BEG[11] ,
    \Tile_X3Y2_EE4BEG[10] ,
    \Tile_X3Y2_EE4BEG[9] ,
    \Tile_X3Y2_EE4BEG[8] ,
    \Tile_X3Y2_EE4BEG[7] ,
    \Tile_X3Y2_EE4BEG[6] ,
    \Tile_X3Y2_EE4BEG[5] ,
    \Tile_X3Y2_EE4BEG[4] ,
    \Tile_X3Y2_EE4BEG[3] ,
    \Tile_X3Y2_EE4BEG[2] ,
    \Tile_X3Y2_EE4BEG[1] ,
    \Tile_X3Y2_EE4BEG[0] }),
    .EE4END({\Tile_X2Y2_EE4BEG[15] ,
    \Tile_X2Y2_EE4BEG[14] ,
    \Tile_X2Y2_EE4BEG[13] ,
    \Tile_X2Y2_EE4BEG[12] ,
    \Tile_X2Y2_EE4BEG[11] ,
    \Tile_X2Y2_EE4BEG[10] ,
    \Tile_X2Y2_EE4BEG[9] ,
    \Tile_X2Y2_EE4BEG[8] ,
    \Tile_X2Y2_EE4BEG[7] ,
    \Tile_X2Y2_EE4BEG[6] ,
    \Tile_X2Y2_EE4BEG[5] ,
    \Tile_X2Y2_EE4BEG[4] ,
    \Tile_X2Y2_EE4BEG[3] ,
    \Tile_X2Y2_EE4BEG[2] ,
    \Tile_X2Y2_EE4BEG[1] ,
    \Tile_X2Y2_EE4BEG[0] }),
    .FrameData({\Tile_X2Y2_FrameData_O[31] ,
    \Tile_X2Y2_FrameData_O[30] ,
    \Tile_X2Y2_FrameData_O[29] ,
    \Tile_X2Y2_FrameData_O[28] ,
    \Tile_X2Y2_FrameData_O[27] ,
    \Tile_X2Y2_FrameData_O[26] ,
    \Tile_X2Y2_FrameData_O[25] ,
    \Tile_X2Y2_FrameData_O[24] ,
    \Tile_X2Y2_FrameData_O[23] ,
    \Tile_X2Y2_FrameData_O[22] ,
    \Tile_X2Y2_FrameData_O[21] ,
    \Tile_X2Y2_FrameData_O[20] ,
    \Tile_X2Y2_FrameData_O[19] ,
    \Tile_X2Y2_FrameData_O[18] ,
    \Tile_X2Y2_FrameData_O[17] ,
    \Tile_X2Y2_FrameData_O[16] ,
    \Tile_X2Y2_FrameData_O[15] ,
    \Tile_X2Y2_FrameData_O[14] ,
    \Tile_X2Y2_FrameData_O[13] ,
    \Tile_X2Y2_FrameData_O[12] ,
    \Tile_X2Y2_FrameData_O[11] ,
    \Tile_X2Y2_FrameData_O[10] ,
    \Tile_X2Y2_FrameData_O[9] ,
    \Tile_X2Y2_FrameData_O[8] ,
    \Tile_X2Y2_FrameData_O[7] ,
    \Tile_X2Y2_FrameData_O[6] ,
    \Tile_X2Y2_FrameData_O[5] ,
    \Tile_X2Y2_FrameData_O[4] ,
    \Tile_X2Y2_FrameData_O[3] ,
    \Tile_X2Y2_FrameData_O[2] ,
    \Tile_X2Y2_FrameData_O[1] ,
    \Tile_X2Y2_FrameData_O[0] }),
    .FrameData_O({\Tile_X3Y2_FrameData_O[31] ,
    \Tile_X3Y2_FrameData_O[30] ,
    \Tile_X3Y2_FrameData_O[29] ,
    \Tile_X3Y2_FrameData_O[28] ,
    \Tile_X3Y2_FrameData_O[27] ,
    \Tile_X3Y2_FrameData_O[26] ,
    \Tile_X3Y2_FrameData_O[25] ,
    \Tile_X3Y2_FrameData_O[24] ,
    \Tile_X3Y2_FrameData_O[23] ,
    \Tile_X3Y2_FrameData_O[22] ,
    \Tile_X3Y2_FrameData_O[21] ,
    \Tile_X3Y2_FrameData_O[20] ,
    \Tile_X3Y2_FrameData_O[19] ,
    \Tile_X3Y2_FrameData_O[18] ,
    \Tile_X3Y2_FrameData_O[17] ,
    \Tile_X3Y2_FrameData_O[16] ,
    \Tile_X3Y2_FrameData_O[15] ,
    \Tile_X3Y2_FrameData_O[14] ,
    \Tile_X3Y2_FrameData_O[13] ,
    \Tile_X3Y2_FrameData_O[12] ,
    \Tile_X3Y2_FrameData_O[11] ,
    \Tile_X3Y2_FrameData_O[10] ,
    \Tile_X3Y2_FrameData_O[9] ,
    \Tile_X3Y2_FrameData_O[8] ,
    \Tile_X3Y2_FrameData_O[7] ,
    \Tile_X3Y2_FrameData_O[6] ,
    \Tile_X3Y2_FrameData_O[5] ,
    \Tile_X3Y2_FrameData_O[4] ,
    \Tile_X3Y2_FrameData_O[3] ,
    \Tile_X3Y2_FrameData_O[2] ,
    \Tile_X3Y2_FrameData_O[1] ,
    \Tile_X3Y2_FrameData_O[0] }),
    .FrameStrobe({\Tile_X3Y3_FrameStrobe_O[19] ,
    \Tile_X3Y3_FrameStrobe_O[18] ,
    \Tile_X3Y3_FrameStrobe_O[17] ,
    \Tile_X3Y3_FrameStrobe_O[16] ,
    \Tile_X3Y3_FrameStrobe_O[15] ,
    \Tile_X3Y3_FrameStrobe_O[14] ,
    \Tile_X3Y3_FrameStrobe_O[13] ,
    \Tile_X3Y3_FrameStrobe_O[12] ,
    \Tile_X3Y3_FrameStrobe_O[11] ,
    \Tile_X3Y3_FrameStrobe_O[10] ,
    \Tile_X3Y3_FrameStrobe_O[9] ,
    \Tile_X3Y3_FrameStrobe_O[8] ,
    \Tile_X3Y3_FrameStrobe_O[7] ,
    \Tile_X3Y3_FrameStrobe_O[6] ,
    \Tile_X3Y3_FrameStrobe_O[5] ,
    \Tile_X3Y3_FrameStrobe_O[4] ,
    \Tile_X3Y3_FrameStrobe_O[3] ,
    \Tile_X3Y3_FrameStrobe_O[2] ,
    \Tile_X3Y3_FrameStrobe_O[1] ,
    \Tile_X3Y3_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X3Y2_FrameStrobe_O[19] ,
    \Tile_X3Y2_FrameStrobe_O[18] ,
    \Tile_X3Y2_FrameStrobe_O[17] ,
    \Tile_X3Y2_FrameStrobe_O[16] ,
    \Tile_X3Y2_FrameStrobe_O[15] ,
    \Tile_X3Y2_FrameStrobe_O[14] ,
    \Tile_X3Y2_FrameStrobe_O[13] ,
    \Tile_X3Y2_FrameStrobe_O[12] ,
    \Tile_X3Y2_FrameStrobe_O[11] ,
    \Tile_X3Y2_FrameStrobe_O[10] ,
    \Tile_X3Y2_FrameStrobe_O[9] ,
    \Tile_X3Y2_FrameStrobe_O[8] ,
    \Tile_X3Y2_FrameStrobe_O[7] ,
    \Tile_X3Y2_FrameStrobe_O[6] ,
    \Tile_X3Y2_FrameStrobe_O[5] ,
    \Tile_X3Y2_FrameStrobe_O[4] ,
    \Tile_X3Y2_FrameStrobe_O[3] ,
    \Tile_X3Y2_FrameStrobe_O[2] ,
    \Tile_X3Y2_FrameStrobe_O[1] ,
    \Tile_X3Y2_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X3Y2_N1BEG[3] ,
    \Tile_X3Y2_N1BEG[2] ,
    \Tile_X3Y2_N1BEG[1] ,
    \Tile_X3Y2_N1BEG[0] }),
    .N1END({\Tile_X3Y3_N1BEG[3] ,
    \Tile_X3Y3_N1BEG[2] ,
    \Tile_X3Y3_N1BEG[1] ,
    \Tile_X3Y3_N1BEG[0] }),
    .N2BEG({\Tile_X3Y2_N2BEG[7] ,
    \Tile_X3Y2_N2BEG[6] ,
    \Tile_X3Y2_N2BEG[5] ,
    \Tile_X3Y2_N2BEG[4] ,
    \Tile_X3Y2_N2BEG[3] ,
    \Tile_X3Y2_N2BEG[2] ,
    \Tile_X3Y2_N2BEG[1] ,
    \Tile_X3Y2_N2BEG[0] }),
    .N2BEGb({\Tile_X3Y2_N2BEGb[7] ,
    \Tile_X3Y2_N2BEGb[6] ,
    \Tile_X3Y2_N2BEGb[5] ,
    \Tile_X3Y2_N2BEGb[4] ,
    \Tile_X3Y2_N2BEGb[3] ,
    \Tile_X3Y2_N2BEGb[2] ,
    \Tile_X3Y2_N2BEGb[1] ,
    \Tile_X3Y2_N2BEGb[0] }),
    .N2END({\Tile_X3Y3_N2BEGb[7] ,
    \Tile_X3Y3_N2BEGb[6] ,
    \Tile_X3Y3_N2BEGb[5] ,
    \Tile_X3Y3_N2BEGb[4] ,
    \Tile_X3Y3_N2BEGb[3] ,
    \Tile_X3Y3_N2BEGb[2] ,
    \Tile_X3Y3_N2BEGb[1] ,
    \Tile_X3Y3_N2BEGb[0] }),
    .N2MID({\Tile_X3Y3_N2BEG[7] ,
    \Tile_X3Y3_N2BEG[6] ,
    \Tile_X3Y3_N2BEG[5] ,
    \Tile_X3Y3_N2BEG[4] ,
    \Tile_X3Y3_N2BEG[3] ,
    \Tile_X3Y3_N2BEG[2] ,
    \Tile_X3Y3_N2BEG[1] ,
    \Tile_X3Y3_N2BEG[0] }),
    .N4BEG({\Tile_X3Y2_N4BEG[15] ,
    \Tile_X3Y2_N4BEG[14] ,
    \Tile_X3Y2_N4BEG[13] ,
    \Tile_X3Y2_N4BEG[12] ,
    \Tile_X3Y2_N4BEG[11] ,
    \Tile_X3Y2_N4BEG[10] ,
    \Tile_X3Y2_N4BEG[9] ,
    \Tile_X3Y2_N4BEG[8] ,
    \Tile_X3Y2_N4BEG[7] ,
    \Tile_X3Y2_N4BEG[6] ,
    \Tile_X3Y2_N4BEG[5] ,
    \Tile_X3Y2_N4BEG[4] ,
    \Tile_X3Y2_N4BEG[3] ,
    \Tile_X3Y2_N4BEG[2] ,
    \Tile_X3Y2_N4BEG[1] ,
    \Tile_X3Y2_N4BEG[0] }),
    .N4END({\Tile_X3Y3_N4BEG[15] ,
    \Tile_X3Y3_N4BEG[14] ,
    \Tile_X3Y3_N4BEG[13] ,
    \Tile_X3Y3_N4BEG[12] ,
    \Tile_X3Y3_N4BEG[11] ,
    \Tile_X3Y3_N4BEG[10] ,
    \Tile_X3Y3_N4BEG[9] ,
    \Tile_X3Y3_N4BEG[8] ,
    \Tile_X3Y3_N4BEG[7] ,
    \Tile_X3Y3_N4BEG[6] ,
    \Tile_X3Y3_N4BEG[5] ,
    \Tile_X3Y3_N4BEG[4] ,
    \Tile_X3Y3_N4BEG[3] ,
    \Tile_X3Y3_N4BEG[2] ,
    \Tile_X3Y3_N4BEG[1] ,
    \Tile_X3Y3_N4BEG[0] }),
    .NN4BEG({\Tile_X3Y2_NN4BEG[15] ,
    \Tile_X3Y2_NN4BEG[14] ,
    \Tile_X3Y2_NN4BEG[13] ,
    \Tile_X3Y2_NN4BEG[12] ,
    \Tile_X3Y2_NN4BEG[11] ,
    \Tile_X3Y2_NN4BEG[10] ,
    \Tile_X3Y2_NN4BEG[9] ,
    \Tile_X3Y2_NN4BEG[8] ,
    \Tile_X3Y2_NN4BEG[7] ,
    \Tile_X3Y2_NN4BEG[6] ,
    \Tile_X3Y2_NN4BEG[5] ,
    \Tile_X3Y2_NN4BEG[4] ,
    \Tile_X3Y2_NN4BEG[3] ,
    \Tile_X3Y2_NN4BEG[2] ,
    \Tile_X3Y2_NN4BEG[1] ,
    \Tile_X3Y2_NN4BEG[0] }),
    .NN4END({\Tile_X3Y3_NN4BEG[15] ,
    \Tile_X3Y3_NN4BEG[14] ,
    \Tile_X3Y3_NN4BEG[13] ,
    \Tile_X3Y3_NN4BEG[12] ,
    \Tile_X3Y3_NN4BEG[11] ,
    \Tile_X3Y3_NN4BEG[10] ,
    \Tile_X3Y3_NN4BEG[9] ,
    \Tile_X3Y3_NN4BEG[8] ,
    \Tile_X3Y3_NN4BEG[7] ,
    \Tile_X3Y3_NN4BEG[6] ,
    \Tile_X3Y3_NN4BEG[5] ,
    \Tile_X3Y3_NN4BEG[4] ,
    \Tile_X3Y3_NN4BEG[3] ,
    \Tile_X3Y3_NN4BEG[2] ,
    \Tile_X3Y3_NN4BEG[1] ,
    \Tile_X3Y3_NN4BEG[0] }),
    .S1BEG({\Tile_X3Y2_S1BEG[3] ,
    \Tile_X3Y2_S1BEG[2] ,
    \Tile_X3Y2_S1BEG[1] ,
    \Tile_X3Y2_S1BEG[0] }),
    .S1END({\Tile_X3Y1_S1BEG[3] ,
    \Tile_X3Y1_S1BEG[2] ,
    \Tile_X3Y1_S1BEG[1] ,
    \Tile_X3Y1_S1BEG[0] }),
    .S2BEG({\Tile_X3Y2_S2BEG[7] ,
    \Tile_X3Y2_S2BEG[6] ,
    \Tile_X3Y2_S2BEG[5] ,
    \Tile_X3Y2_S2BEG[4] ,
    \Tile_X3Y2_S2BEG[3] ,
    \Tile_X3Y2_S2BEG[2] ,
    \Tile_X3Y2_S2BEG[1] ,
    \Tile_X3Y2_S2BEG[0] }),
    .S2BEGb({\Tile_X3Y2_S2BEGb[7] ,
    \Tile_X3Y2_S2BEGb[6] ,
    \Tile_X3Y2_S2BEGb[5] ,
    \Tile_X3Y2_S2BEGb[4] ,
    \Tile_X3Y2_S2BEGb[3] ,
    \Tile_X3Y2_S2BEGb[2] ,
    \Tile_X3Y2_S2BEGb[1] ,
    \Tile_X3Y2_S2BEGb[0] }),
    .S2END({\Tile_X3Y1_S2BEGb[7] ,
    \Tile_X3Y1_S2BEGb[6] ,
    \Tile_X3Y1_S2BEGb[5] ,
    \Tile_X3Y1_S2BEGb[4] ,
    \Tile_X3Y1_S2BEGb[3] ,
    \Tile_X3Y1_S2BEGb[2] ,
    \Tile_X3Y1_S2BEGb[1] ,
    \Tile_X3Y1_S2BEGb[0] }),
    .S2MID({\Tile_X3Y1_S2BEG[7] ,
    \Tile_X3Y1_S2BEG[6] ,
    \Tile_X3Y1_S2BEG[5] ,
    \Tile_X3Y1_S2BEG[4] ,
    \Tile_X3Y1_S2BEG[3] ,
    \Tile_X3Y1_S2BEG[2] ,
    \Tile_X3Y1_S2BEG[1] ,
    \Tile_X3Y1_S2BEG[0] }),
    .S4BEG({\Tile_X3Y2_S4BEG[15] ,
    \Tile_X3Y2_S4BEG[14] ,
    \Tile_X3Y2_S4BEG[13] ,
    \Tile_X3Y2_S4BEG[12] ,
    \Tile_X3Y2_S4BEG[11] ,
    \Tile_X3Y2_S4BEG[10] ,
    \Tile_X3Y2_S4BEG[9] ,
    \Tile_X3Y2_S4BEG[8] ,
    \Tile_X3Y2_S4BEG[7] ,
    \Tile_X3Y2_S4BEG[6] ,
    \Tile_X3Y2_S4BEG[5] ,
    \Tile_X3Y2_S4BEG[4] ,
    \Tile_X3Y2_S4BEG[3] ,
    \Tile_X3Y2_S4BEG[2] ,
    \Tile_X3Y2_S4BEG[1] ,
    \Tile_X3Y2_S4BEG[0] }),
    .S4END({\Tile_X3Y1_S4BEG[15] ,
    \Tile_X3Y1_S4BEG[14] ,
    \Tile_X3Y1_S4BEG[13] ,
    \Tile_X3Y1_S4BEG[12] ,
    \Tile_X3Y1_S4BEG[11] ,
    \Tile_X3Y1_S4BEG[10] ,
    \Tile_X3Y1_S4BEG[9] ,
    \Tile_X3Y1_S4BEG[8] ,
    \Tile_X3Y1_S4BEG[7] ,
    \Tile_X3Y1_S4BEG[6] ,
    \Tile_X3Y1_S4BEG[5] ,
    \Tile_X3Y1_S4BEG[4] ,
    \Tile_X3Y1_S4BEG[3] ,
    \Tile_X3Y1_S4BEG[2] ,
    \Tile_X3Y1_S4BEG[1] ,
    \Tile_X3Y1_S4BEG[0] }),
    .SS4BEG({\Tile_X3Y2_SS4BEG[15] ,
    \Tile_X3Y2_SS4BEG[14] ,
    \Tile_X3Y2_SS4BEG[13] ,
    \Tile_X3Y2_SS4BEG[12] ,
    \Tile_X3Y2_SS4BEG[11] ,
    \Tile_X3Y2_SS4BEG[10] ,
    \Tile_X3Y2_SS4BEG[9] ,
    \Tile_X3Y2_SS4BEG[8] ,
    \Tile_X3Y2_SS4BEG[7] ,
    \Tile_X3Y2_SS4BEG[6] ,
    \Tile_X3Y2_SS4BEG[5] ,
    \Tile_X3Y2_SS4BEG[4] ,
    \Tile_X3Y2_SS4BEG[3] ,
    \Tile_X3Y2_SS4BEG[2] ,
    \Tile_X3Y2_SS4BEG[1] ,
    \Tile_X3Y2_SS4BEG[0] }),
    .SS4END({\Tile_X3Y1_SS4BEG[15] ,
    \Tile_X3Y1_SS4BEG[14] ,
    \Tile_X3Y1_SS4BEG[13] ,
    \Tile_X3Y1_SS4BEG[12] ,
    \Tile_X3Y1_SS4BEG[11] ,
    \Tile_X3Y1_SS4BEG[10] ,
    \Tile_X3Y1_SS4BEG[9] ,
    \Tile_X3Y1_SS4BEG[8] ,
    \Tile_X3Y1_SS4BEG[7] ,
    \Tile_X3Y1_SS4BEG[6] ,
    \Tile_X3Y1_SS4BEG[5] ,
    \Tile_X3Y1_SS4BEG[4] ,
    \Tile_X3Y1_SS4BEG[3] ,
    \Tile_X3Y1_SS4BEG[2] ,
    \Tile_X3Y1_SS4BEG[1] ,
    \Tile_X3Y1_SS4BEG[0] }),
    .W1BEG({\Tile_X3Y2_W1BEG[3] ,
    \Tile_X3Y2_W1BEG[2] ,
    \Tile_X3Y2_W1BEG[1] ,
    \Tile_X3Y2_W1BEG[0] }),
    .W1END({\Tile_X4Y2_W1BEG[3] ,
    \Tile_X4Y2_W1BEG[2] ,
    \Tile_X4Y2_W1BEG[1] ,
    \Tile_X4Y2_W1BEG[0] }),
    .W2BEG({\Tile_X3Y2_W2BEG[7] ,
    \Tile_X3Y2_W2BEG[6] ,
    \Tile_X3Y2_W2BEG[5] ,
    \Tile_X3Y2_W2BEG[4] ,
    \Tile_X3Y2_W2BEG[3] ,
    \Tile_X3Y2_W2BEG[2] ,
    \Tile_X3Y2_W2BEG[1] ,
    \Tile_X3Y2_W2BEG[0] }),
    .W2BEGb({\Tile_X3Y2_W2BEGb[7] ,
    \Tile_X3Y2_W2BEGb[6] ,
    \Tile_X3Y2_W2BEGb[5] ,
    \Tile_X3Y2_W2BEGb[4] ,
    \Tile_X3Y2_W2BEGb[3] ,
    \Tile_X3Y2_W2BEGb[2] ,
    \Tile_X3Y2_W2BEGb[1] ,
    \Tile_X3Y2_W2BEGb[0] }),
    .W2END({\Tile_X4Y2_W2BEGb[7] ,
    \Tile_X4Y2_W2BEGb[6] ,
    \Tile_X4Y2_W2BEGb[5] ,
    \Tile_X4Y2_W2BEGb[4] ,
    \Tile_X4Y2_W2BEGb[3] ,
    \Tile_X4Y2_W2BEGb[2] ,
    \Tile_X4Y2_W2BEGb[1] ,
    \Tile_X4Y2_W2BEGb[0] }),
    .W2MID({\Tile_X4Y2_W2BEG[7] ,
    \Tile_X4Y2_W2BEG[6] ,
    \Tile_X4Y2_W2BEG[5] ,
    \Tile_X4Y2_W2BEG[4] ,
    \Tile_X4Y2_W2BEG[3] ,
    \Tile_X4Y2_W2BEG[2] ,
    \Tile_X4Y2_W2BEG[1] ,
    \Tile_X4Y2_W2BEG[0] }),
    .W6BEG({\Tile_X3Y2_W6BEG[11] ,
    \Tile_X3Y2_W6BEG[10] ,
    \Tile_X3Y2_W6BEG[9] ,
    \Tile_X3Y2_W6BEG[8] ,
    \Tile_X3Y2_W6BEG[7] ,
    \Tile_X3Y2_W6BEG[6] ,
    \Tile_X3Y2_W6BEG[5] ,
    \Tile_X3Y2_W6BEG[4] ,
    \Tile_X3Y2_W6BEG[3] ,
    \Tile_X3Y2_W6BEG[2] ,
    \Tile_X3Y2_W6BEG[1] ,
    \Tile_X3Y2_W6BEG[0] }),
    .W6END({\Tile_X4Y2_W6BEG[11] ,
    \Tile_X4Y2_W6BEG[10] ,
    \Tile_X4Y2_W6BEG[9] ,
    \Tile_X4Y2_W6BEG[8] ,
    \Tile_X4Y2_W6BEG[7] ,
    \Tile_X4Y2_W6BEG[6] ,
    \Tile_X4Y2_W6BEG[5] ,
    \Tile_X4Y2_W6BEG[4] ,
    \Tile_X4Y2_W6BEG[3] ,
    \Tile_X4Y2_W6BEG[2] ,
    \Tile_X4Y2_W6BEG[1] ,
    \Tile_X4Y2_W6BEG[0] }),
    .WW4BEG({\Tile_X3Y2_WW4BEG[15] ,
    \Tile_X3Y2_WW4BEG[14] ,
    \Tile_X3Y2_WW4BEG[13] ,
    \Tile_X3Y2_WW4BEG[12] ,
    \Tile_X3Y2_WW4BEG[11] ,
    \Tile_X3Y2_WW4BEG[10] ,
    \Tile_X3Y2_WW4BEG[9] ,
    \Tile_X3Y2_WW4BEG[8] ,
    \Tile_X3Y2_WW4BEG[7] ,
    \Tile_X3Y2_WW4BEG[6] ,
    \Tile_X3Y2_WW4BEG[5] ,
    \Tile_X3Y2_WW4BEG[4] ,
    \Tile_X3Y2_WW4BEG[3] ,
    \Tile_X3Y2_WW4BEG[2] ,
    \Tile_X3Y2_WW4BEG[1] ,
    \Tile_X3Y2_WW4BEG[0] }),
    .WW4END({\Tile_X4Y2_WW4BEG[15] ,
    \Tile_X4Y2_WW4BEG[14] ,
    \Tile_X4Y2_WW4BEG[13] ,
    \Tile_X4Y2_WW4BEG[12] ,
    \Tile_X4Y2_WW4BEG[11] ,
    \Tile_X4Y2_WW4BEG[10] ,
    \Tile_X4Y2_WW4BEG[9] ,
    \Tile_X4Y2_WW4BEG[8] ,
    \Tile_X4Y2_WW4BEG[7] ,
    \Tile_X4Y2_WW4BEG[6] ,
    \Tile_X4Y2_WW4BEG[5] ,
    \Tile_X4Y2_WW4BEG[4] ,
    \Tile_X4Y2_WW4BEG[3] ,
    \Tile_X4Y2_WW4BEG[2] ,
    \Tile_X4Y2_WW4BEG[1] ,
    \Tile_X4Y2_WW4BEG[0] }));
 LUT4AB Tile_X3Y3_LUT4AB (.Ci(Tile_X3Y4_Co),
    .Co(Tile_X3Y3_Co),
    .UserCLK(Tile_X3Y4_UserCLKo),
    .UserCLKo(Tile_X3Y3_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X3Y3_E1BEG[3] ,
    \Tile_X3Y3_E1BEG[2] ,
    \Tile_X3Y3_E1BEG[1] ,
    \Tile_X3Y3_E1BEG[0] }),
    .E1END({\Tile_X2Y3_E1BEG[3] ,
    \Tile_X2Y3_E1BEG[2] ,
    \Tile_X2Y3_E1BEG[1] ,
    \Tile_X2Y3_E1BEG[0] }),
    .E2BEG({\Tile_X3Y3_E2BEG[7] ,
    \Tile_X3Y3_E2BEG[6] ,
    \Tile_X3Y3_E2BEG[5] ,
    \Tile_X3Y3_E2BEG[4] ,
    \Tile_X3Y3_E2BEG[3] ,
    \Tile_X3Y3_E2BEG[2] ,
    \Tile_X3Y3_E2BEG[1] ,
    \Tile_X3Y3_E2BEG[0] }),
    .E2BEGb({\Tile_X3Y3_E2BEGb[7] ,
    \Tile_X3Y3_E2BEGb[6] ,
    \Tile_X3Y3_E2BEGb[5] ,
    \Tile_X3Y3_E2BEGb[4] ,
    \Tile_X3Y3_E2BEGb[3] ,
    \Tile_X3Y3_E2BEGb[2] ,
    \Tile_X3Y3_E2BEGb[1] ,
    \Tile_X3Y3_E2BEGb[0] }),
    .E2END({\Tile_X2Y3_E2BEGb[7] ,
    \Tile_X2Y3_E2BEGb[6] ,
    \Tile_X2Y3_E2BEGb[5] ,
    \Tile_X2Y3_E2BEGb[4] ,
    \Tile_X2Y3_E2BEGb[3] ,
    \Tile_X2Y3_E2BEGb[2] ,
    \Tile_X2Y3_E2BEGb[1] ,
    \Tile_X2Y3_E2BEGb[0] }),
    .E2MID({\Tile_X2Y3_E2BEG[7] ,
    \Tile_X2Y3_E2BEG[6] ,
    \Tile_X2Y3_E2BEG[5] ,
    \Tile_X2Y3_E2BEG[4] ,
    \Tile_X2Y3_E2BEG[3] ,
    \Tile_X2Y3_E2BEG[2] ,
    \Tile_X2Y3_E2BEG[1] ,
    \Tile_X2Y3_E2BEG[0] }),
    .E6BEG({\Tile_X3Y3_E6BEG[11] ,
    \Tile_X3Y3_E6BEG[10] ,
    \Tile_X3Y3_E6BEG[9] ,
    \Tile_X3Y3_E6BEG[8] ,
    \Tile_X3Y3_E6BEG[7] ,
    \Tile_X3Y3_E6BEG[6] ,
    \Tile_X3Y3_E6BEG[5] ,
    \Tile_X3Y3_E6BEG[4] ,
    \Tile_X3Y3_E6BEG[3] ,
    \Tile_X3Y3_E6BEG[2] ,
    \Tile_X3Y3_E6BEG[1] ,
    \Tile_X3Y3_E6BEG[0] }),
    .E6END({\Tile_X2Y3_E6BEG[11] ,
    \Tile_X2Y3_E6BEG[10] ,
    \Tile_X2Y3_E6BEG[9] ,
    \Tile_X2Y3_E6BEG[8] ,
    \Tile_X2Y3_E6BEG[7] ,
    \Tile_X2Y3_E6BEG[6] ,
    \Tile_X2Y3_E6BEG[5] ,
    \Tile_X2Y3_E6BEG[4] ,
    \Tile_X2Y3_E6BEG[3] ,
    \Tile_X2Y3_E6BEG[2] ,
    \Tile_X2Y3_E6BEG[1] ,
    \Tile_X2Y3_E6BEG[0] }),
    .EE4BEG({\Tile_X3Y3_EE4BEG[15] ,
    \Tile_X3Y3_EE4BEG[14] ,
    \Tile_X3Y3_EE4BEG[13] ,
    \Tile_X3Y3_EE4BEG[12] ,
    \Tile_X3Y3_EE4BEG[11] ,
    \Tile_X3Y3_EE4BEG[10] ,
    \Tile_X3Y3_EE4BEG[9] ,
    \Tile_X3Y3_EE4BEG[8] ,
    \Tile_X3Y3_EE4BEG[7] ,
    \Tile_X3Y3_EE4BEG[6] ,
    \Tile_X3Y3_EE4BEG[5] ,
    \Tile_X3Y3_EE4BEG[4] ,
    \Tile_X3Y3_EE4BEG[3] ,
    \Tile_X3Y3_EE4BEG[2] ,
    \Tile_X3Y3_EE4BEG[1] ,
    \Tile_X3Y3_EE4BEG[0] }),
    .EE4END({\Tile_X2Y3_EE4BEG[15] ,
    \Tile_X2Y3_EE4BEG[14] ,
    \Tile_X2Y3_EE4BEG[13] ,
    \Tile_X2Y3_EE4BEG[12] ,
    \Tile_X2Y3_EE4BEG[11] ,
    \Tile_X2Y3_EE4BEG[10] ,
    \Tile_X2Y3_EE4BEG[9] ,
    \Tile_X2Y3_EE4BEG[8] ,
    \Tile_X2Y3_EE4BEG[7] ,
    \Tile_X2Y3_EE4BEG[6] ,
    \Tile_X2Y3_EE4BEG[5] ,
    \Tile_X2Y3_EE4BEG[4] ,
    \Tile_X2Y3_EE4BEG[3] ,
    \Tile_X2Y3_EE4BEG[2] ,
    \Tile_X2Y3_EE4BEG[1] ,
    \Tile_X2Y3_EE4BEG[0] }),
    .FrameData({\Tile_X2Y3_FrameData_O[31] ,
    \Tile_X2Y3_FrameData_O[30] ,
    \Tile_X2Y3_FrameData_O[29] ,
    \Tile_X2Y3_FrameData_O[28] ,
    \Tile_X2Y3_FrameData_O[27] ,
    \Tile_X2Y3_FrameData_O[26] ,
    \Tile_X2Y3_FrameData_O[25] ,
    \Tile_X2Y3_FrameData_O[24] ,
    \Tile_X2Y3_FrameData_O[23] ,
    \Tile_X2Y3_FrameData_O[22] ,
    \Tile_X2Y3_FrameData_O[21] ,
    \Tile_X2Y3_FrameData_O[20] ,
    \Tile_X2Y3_FrameData_O[19] ,
    \Tile_X2Y3_FrameData_O[18] ,
    \Tile_X2Y3_FrameData_O[17] ,
    \Tile_X2Y3_FrameData_O[16] ,
    \Tile_X2Y3_FrameData_O[15] ,
    \Tile_X2Y3_FrameData_O[14] ,
    \Tile_X2Y3_FrameData_O[13] ,
    \Tile_X2Y3_FrameData_O[12] ,
    \Tile_X2Y3_FrameData_O[11] ,
    \Tile_X2Y3_FrameData_O[10] ,
    \Tile_X2Y3_FrameData_O[9] ,
    \Tile_X2Y3_FrameData_O[8] ,
    \Tile_X2Y3_FrameData_O[7] ,
    \Tile_X2Y3_FrameData_O[6] ,
    \Tile_X2Y3_FrameData_O[5] ,
    \Tile_X2Y3_FrameData_O[4] ,
    \Tile_X2Y3_FrameData_O[3] ,
    \Tile_X2Y3_FrameData_O[2] ,
    \Tile_X2Y3_FrameData_O[1] ,
    \Tile_X2Y3_FrameData_O[0] }),
    .FrameData_O({\Tile_X3Y3_FrameData_O[31] ,
    \Tile_X3Y3_FrameData_O[30] ,
    \Tile_X3Y3_FrameData_O[29] ,
    \Tile_X3Y3_FrameData_O[28] ,
    \Tile_X3Y3_FrameData_O[27] ,
    \Tile_X3Y3_FrameData_O[26] ,
    \Tile_X3Y3_FrameData_O[25] ,
    \Tile_X3Y3_FrameData_O[24] ,
    \Tile_X3Y3_FrameData_O[23] ,
    \Tile_X3Y3_FrameData_O[22] ,
    \Tile_X3Y3_FrameData_O[21] ,
    \Tile_X3Y3_FrameData_O[20] ,
    \Tile_X3Y3_FrameData_O[19] ,
    \Tile_X3Y3_FrameData_O[18] ,
    \Tile_X3Y3_FrameData_O[17] ,
    \Tile_X3Y3_FrameData_O[16] ,
    \Tile_X3Y3_FrameData_O[15] ,
    \Tile_X3Y3_FrameData_O[14] ,
    \Tile_X3Y3_FrameData_O[13] ,
    \Tile_X3Y3_FrameData_O[12] ,
    \Tile_X3Y3_FrameData_O[11] ,
    \Tile_X3Y3_FrameData_O[10] ,
    \Tile_X3Y3_FrameData_O[9] ,
    \Tile_X3Y3_FrameData_O[8] ,
    \Tile_X3Y3_FrameData_O[7] ,
    \Tile_X3Y3_FrameData_O[6] ,
    \Tile_X3Y3_FrameData_O[5] ,
    \Tile_X3Y3_FrameData_O[4] ,
    \Tile_X3Y3_FrameData_O[3] ,
    \Tile_X3Y3_FrameData_O[2] ,
    \Tile_X3Y3_FrameData_O[1] ,
    \Tile_X3Y3_FrameData_O[0] }),
    .FrameStrobe({\Tile_X3Y4_FrameStrobe_O[19] ,
    \Tile_X3Y4_FrameStrobe_O[18] ,
    \Tile_X3Y4_FrameStrobe_O[17] ,
    \Tile_X3Y4_FrameStrobe_O[16] ,
    \Tile_X3Y4_FrameStrobe_O[15] ,
    \Tile_X3Y4_FrameStrobe_O[14] ,
    \Tile_X3Y4_FrameStrobe_O[13] ,
    \Tile_X3Y4_FrameStrobe_O[12] ,
    \Tile_X3Y4_FrameStrobe_O[11] ,
    \Tile_X3Y4_FrameStrobe_O[10] ,
    \Tile_X3Y4_FrameStrobe_O[9] ,
    \Tile_X3Y4_FrameStrobe_O[8] ,
    \Tile_X3Y4_FrameStrobe_O[7] ,
    \Tile_X3Y4_FrameStrobe_O[6] ,
    \Tile_X3Y4_FrameStrobe_O[5] ,
    \Tile_X3Y4_FrameStrobe_O[4] ,
    \Tile_X3Y4_FrameStrobe_O[3] ,
    \Tile_X3Y4_FrameStrobe_O[2] ,
    \Tile_X3Y4_FrameStrobe_O[1] ,
    \Tile_X3Y4_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X3Y3_FrameStrobe_O[19] ,
    \Tile_X3Y3_FrameStrobe_O[18] ,
    \Tile_X3Y3_FrameStrobe_O[17] ,
    \Tile_X3Y3_FrameStrobe_O[16] ,
    \Tile_X3Y3_FrameStrobe_O[15] ,
    \Tile_X3Y3_FrameStrobe_O[14] ,
    \Tile_X3Y3_FrameStrobe_O[13] ,
    \Tile_X3Y3_FrameStrobe_O[12] ,
    \Tile_X3Y3_FrameStrobe_O[11] ,
    \Tile_X3Y3_FrameStrobe_O[10] ,
    \Tile_X3Y3_FrameStrobe_O[9] ,
    \Tile_X3Y3_FrameStrobe_O[8] ,
    \Tile_X3Y3_FrameStrobe_O[7] ,
    \Tile_X3Y3_FrameStrobe_O[6] ,
    \Tile_X3Y3_FrameStrobe_O[5] ,
    \Tile_X3Y3_FrameStrobe_O[4] ,
    \Tile_X3Y3_FrameStrobe_O[3] ,
    \Tile_X3Y3_FrameStrobe_O[2] ,
    \Tile_X3Y3_FrameStrobe_O[1] ,
    \Tile_X3Y3_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X3Y3_N1BEG[3] ,
    \Tile_X3Y3_N1BEG[2] ,
    \Tile_X3Y3_N1BEG[1] ,
    \Tile_X3Y3_N1BEG[0] }),
    .N1END({\Tile_X3Y4_N1BEG[3] ,
    \Tile_X3Y4_N1BEG[2] ,
    \Tile_X3Y4_N1BEG[1] ,
    \Tile_X3Y4_N1BEG[0] }),
    .N2BEG({\Tile_X3Y3_N2BEG[7] ,
    \Tile_X3Y3_N2BEG[6] ,
    \Tile_X3Y3_N2BEG[5] ,
    \Tile_X3Y3_N2BEG[4] ,
    \Tile_X3Y3_N2BEG[3] ,
    \Tile_X3Y3_N2BEG[2] ,
    \Tile_X3Y3_N2BEG[1] ,
    \Tile_X3Y3_N2BEG[0] }),
    .N2BEGb({\Tile_X3Y3_N2BEGb[7] ,
    \Tile_X3Y3_N2BEGb[6] ,
    \Tile_X3Y3_N2BEGb[5] ,
    \Tile_X3Y3_N2BEGb[4] ,
    \Tile_X3Y3_N2BEGb[3] ,
    \Tile_X3Y3_N2BEGb[2] ,
    \Tile_X3Y3_N2BEGb[1] ,
    \Tile_X3Y3_N2BEGb[0] }),
    .N2END({\Tile_X3Y4_N2BEGb[7] ,
    \Tile_X3Y4_N2BEGb[6] ,
    \Tile_X3Y4_N2BEGb[5] ,
    \Tile_X3Y4_N2BEGb[4] ,
    \Tile_X3Y4_N2BEGb[3] ,
    \Tile_X3Y4_N2BEGb[2] ,
    \Tile_X3Y4_N2BEGb[1] ,
    \Tile_X3Y4_N2BEGb[0] }),
    .N2MID({\Tile_X3Y4_N2BEG[7] ,
    \Tile_X3Y4_N2BEG[6] ,
    \Tile_X3Y4_N2BEG[5] ,
    \Tile_X3Y4_N2BEG[4] ,
    \Tile_X3Y4_N2BEG[3] ,
    \Tile_X3Y4_N2BEG[2] ,
    \Tile_X3Y4_N2BEG[1] ,
    \Tile_X3Y4_N2BEG[0] }),
    .N4BEG({\Tile_X3Y3_N4BEG[15] ,
    \Tile_X3Y3_N4BEG[14] ,
    \Tile_X3Y3_N4BEG[13] ,
    \Tile_X3Y3_N4BEG[12] ,
    \Tile_X3Y3_N4BEG[11] ,
    \Tile_X3Y3_N4BEG[10] ,
    \Tile_X3Y3_N4BEG[9] ,
    \Tile_X3Y3_N4BEG[8] ,
    \Tile_X3Y3_N4BEG[7] ,
    \Tile_X3Y3_N4BEG[6] ,
    \Tile_X3Y3_N4BEG[5] ,
    \Tile_X3Y3_N4BEG[4] ,
    \Tile_X3Y3_N4BEG[3] ,
    \Tile_X3Y3_N4BEG[2] ,
    \Tile_X3Y3_N4BEG[1] ,
    \Tile_X3Y3_N4BEG[0] }),
    .N4END({\Tile_X3Y4_N4BEG[15] ,
    \Tile_X3Y4_N4BEG[14] ,
    \Tile_X3Y4_N4BEG[13] ,
    \Tile_X3Y4_N4BEG[12] ,
    \Tile_X3Y4_N4BEG[11] ,
    \Tile_X3Y4_N4BEG[10] ,
    \Tile_X3Y4_N4BEG[9] ,
    \Tile_X3Y4_N4BEG[8] ,
    \Tile_X3Y4_N4BEG[7] ,
    \Tile_X3Y4_N4BEG[6] ,
    \Tile_X3Y4_N4BEG[5] ,
    \Tile_X3Y4_N4BEG[4] ,
    \Tile_X3Y4_N4BEG[3] ,
    \Tile_X3Y4_N4BEG[2] ,
    \Tile_X3Y4_N4BEG[1] ,
    \Tile_X3Y4_N4BEG[0] }),
    .NN4BEG({\Tile_X3Y3_NN4BEG[15] ,
    \Tile_X3Y3_NN4BEG[14] ,
    \Tile_X3Y3_NN4BEG[13] ,
    \Tile_X3Y3_NN4BEG[12] ,
    \Tile_X3Y3_NN4BEG[11] ,
    \Tile_X3Y3_NN4BEG[10] ,
    \Tile_X3Y3_NN4BEG[9] ,
    \Tile_X3Y3_NN4BEG[8] ,
    \Tile_X3Y3_NN4BEG[7] ,
    \Tile_X3Y3_NN4BEG[6] ,
    \Tile_X3Y3_NN4BEG[5] ,
    \Tile_X3Y3_NN4BEG[4] ,
    \Tile_X3Y3_NN4BEG[3] ,
    \Tile_X3Y3_NN4BEG[2] ,
    \Tile_X3Y3_NN4BEG[1] ,
    \Tile_X3Y3_NN4BEG[0] }),
    .NN4END({\Tile_X3Y4_NN4BEG[15] ,
    \Tile_X3Y4_NN4BEG[14] ,
    \Tile_X3Y4_NN4BEG[13] ,
    \Tile_X3Y4_NN4BEG[12] ,
    \Tile_X3Y4_NN4BEG[11] ,
    \Tile_X3Y4_NN4BEG[10] ,
    \Tile_X3Y4_NN4BEG[9] ,
    \Tile_X3Y4_NN4BEG[8] ,
    \Tile_X3Y4_NN4BEG[7] ,
    \Tile_X3Y4_NN4BEG[6] ,
    \Tile_X3Y4_NN4BEG[5] ,
    \Tile_X3Y4_NN4BEG[4] ,
    \Tile_X3Y4_NN4BEG[3] ,
    \Tile_X3Y4_NN4BEG[2] ,
    \Tile_X3Y4_NN4BEG[1] ,
    \Tile_X3Y4_NN4BEG[0] }),
    .S1BEG({\Tile_X3Y3_S1BEG[3] ,
    \Tile_X3Y3_S1BEG[2] ,
    \Tile_X3Y3_S1BEG[1] ,
    \Tile_X3Y3_S1BEG[0] }),
    .S1END({\Tile_X3Y2_S1BEG[3] ,
    \Tile_X3Y2_S1BEG[2] ,
    \Tile_X3Y2_S1BEG[1] ,
    \Tile_X3Y2_S1BEG[0] }),
    .S2BEG({\Tile_X3Y3_S2BEG[7] ,
    \Tile_X3Y3_S2BEG[6] ,
    \Tile_X3Y3_S2BEG[5] ,
    \Tile_X3Y3_S2BEG[4] ,
    \Tile_X3Y3_S2BEG[3] ,
    \Tile_X3Y3_S2BEG[2] ,
    \Tile_X3Y3_S2BEG[1] ,
    \Tile_X3Y3_S2BEG[0] }),
    .S2BEGb({\Tile_X3Y3_S2BEGb[7] ,
    \Tile_X3Y3_S2BEGb[6] ,
    \Tile_X3Y3_S2BEGb[5] ,
    \Tile_X3Y3_S2BEGb[4] ,
    \Tile_X3Y3_S2BEGb[3] ,
    \Tile_X3Y3_S2BEGb[2] ,
    \Tile_X3Y3_S2BEGb[1] ,
    \Tile_X3Y3_S2BEGb[0] }),
    .S2END({\Tile_X3Y2_S2BEGb[7] ,
    \Tile_X3Y2_S2BEGb[6] ,
    \Tile_X3Y2_S2BEGb[5] ,
    \Tile_X3Y2_S2BEGb[4] ,
    \Tile_X3Y2_S2BEGb[3] ,
    \Tile_X3Y2_S2BEGb[2] ,
    \Tile_X3Y2_S2BEGb[1] ,
    \Tile_X3Y2_S2BEGb[0] }),
    .S2MID({\Tile_X3Y2_S2BEG[7] ,
    \Tile_X3Y2_S2BEG[6] ,
    \Tile_X3Y2_S2BEG[5] ,
    \Tile_X3Y2_S2BEG[4] ,
    \Tile_X3Y2_S2BEG[3] ,
    \Tile_X3Y2_S2BEG[2] ,
    \Tile_X3Y2_S2BEG[1] ,
    \Tile_X3Y2_S2BEG[0] }),
    .S4BEG({\Tile_X3Y3_S4BEG[15] ,
    \Tile_X3Y3_S4BEG[14] ,
    \Tile_X3Y3_S4BEG[13] ,
    \Tile_X3Y3_S4BEG[12] ,
    \Tile_X3Y3_S4BEG[11] ,
    \Tile_X3Y3_S4BEG[10] ,
    \Tile_X3Y3_S4BEG[9] ,
    \Tile_X3Y3_S4BEG[8] ,
    \Tile_X3Y3_S4BEG[7] ,
    \Tile_X3Y3_S4BEG[6] ,
    \Tile_X3Y3_S4BEG[5] ,
    \Tile_X3Y3_S4BEG[4] ,
    \Tile_X3Y3_S4BEG[3] ,
    \Tile_X3Y3_S4BEG[2] ,
    \Tile_X3Y3_S4BEG[1] ,
    \Tile_X3Y3_S4BEG[0] }),
    .S4END({\Tile_X3Y2_S4BEG[15] ,
    \Tile_X3Y2_S4BEG[14] ,
    \Tile_X3Y2_S4BEG[13] ,
    \Tile_X3Y2_S4BEG[12] ,
    \Tile_X3Y2_S4BEG[11] ,
    \Tile_X3Y2_S4BEG[10] ,
    \Tile_X3Y2_S4BEG[9] ,
    \Tile_X3Y2_S4BEG[8] ,
    \Tile_X3Y2_S4BEG[7] ,
    \Tile_X3Y2_S4BEG[6] ,
    \Tile_X3Y2_S4BEG[5] ,
    \Tile_X3Y2_S4BEG[4] ,
    \Tile_X3Y2_S4BEG[3] ,
    \Tile_X3Y2_S4BEG[2] ,
    \Tile_X3Y2_S4BEG[1] ,
    \Tile_X3Y2_S4BEG[0] }),
    .SS4BEG({\Tile_X3Y3_SS4BEG[15] ,
    \Tile_X3Y3_SS4BEG[14] ,
    \Tile_X3Y3_SS4BEG[13] ,
    \Tile_X3Y3_SS4BEG[12] ,
    \Tile_X3Y3_SS4BEG[11] ,
    \Tile_X3Y3_SS4BEG[10] ,
    \Tile_X3Y3_SS4BEG[9] ,
    \Tile_X3Y3_SS4BEG[8] ,
    \Tile_X3Y3_SS4BEG[7] ,
    \Tile_X3Y3_SS4BEG[6] ,
    \Tile_X3Y3_SS4BEG[5] ,
    \Tile_X3Y3_SS4BEG[4] ,
    \Tile_X3Y3_SS4BEG[3] ,
    \Tile_X3Y3_SS4BEG[2] ,
    \Tile_X3Y3_SS4BEG[1] ,
    \Tile_X3Y3_SS4BEG[0] }),
    .SS4END({\Tile_X3Y2_SS4BEG[15] ,
    \Tile_X3Y2_SS4BEG[14] ,
    \Tile_X3Y2_SS4BEG[13] ,
    \Tile_X3Y2_SS4BEG[12] ,
    \Tile_X3Y2_SS4BEG[11] ,
    \Tile_X3Y2_SS4BEG[10] ,
    \Tile_X3Y2_SS4BEG[9] ,
    \Tile_X3Y2_SS4BEG[8] ,
    \Tile_X3Y2_SS4BEG[7] ,
    \Tile_X3Y2_SS4BEG[6] ,
    \Tile_X3Y2_SS4BEG[5] ,
    \Tile_X3Y2_SS4BEG[4] ,
    \Tile_X3Y2_SS4BEG[3] ,
    \Tile_X3Y2_SS4BEG[2] ,
    \Tile_X3Y2_SS4BEG[1] ,
    \Tile_X3Y2_SS4BEG[0] }),
    .W1BEG({\Tile_X3Y3_W1BEG[3] ,
    \Tile_X3Y3_W1BEG[2] ,
    \Tile_X3Y3_W1BEG[1] ,
    \Tile_X3Y3_W1BEG[0] }),
    .W1END({\Tile_X4Y3_W1BEG[3] ,
    \Tile_X4Y3_W1BEG[2] ,
    \Tile_X4Y3_W1BEG[1] ,
    \Tile_X4Y3_W1BEG[0] }),
    .W2BEG({\Tile_X3Y3_W2BEG[7] ,
    \Tile_X3Y3_W2BEG[6] ,
    \Tile_X3Y3_W2BEG[5] ,
    \Tile_X3Y3_W2BEG[4] ,
    \Tile_X3Y3_W2BEG[3] ,
    \Tile_X3Y3_W2BEG[2] ,
    \Tile_X3Y3_W2BEG[1] ,
    \Tile_X3Y3_W2BEG[0] }),
    .W2BEGb({\Tile_X3Y3_W2BEGb[7] ,
    \Tile_X3Y3_W2BEGb[6] ,
    \Tile_X3Y3_W2BEGb[5] ,
    \Tile_X3Y3_W2BEGb[4] ,
    \Tile_X3Y3_W2BEGb[3] ,
    \Tile_X3Y3_W2BEGb[2] ,
    \Tile_X3Y3_W2BEGb[1] ,
    \Tile_X3Y3_W2BEGb[0] }),
    .W2END({\Tile_X4Y3_W2BEGb[7] ,
    \Tile_X4Y3_W2BEGb[6] ,
    \Tile_X4Y3_W2BEGb[5] ,
    \Tile_X4Y3_W2BEGb[4] ,
    \Tile_X4Y3_W2BEGb[3] ,
    \Tile_X4Y3_W2BEGb[2] ,
    \Tile_X4Y3_W2BEGb[1] ,
    \Tile_X4Y3_W2BEGb[0] }),
    .W2MID({\Tile_X4Y3_W2BEG[7] ,
    \Tile_X4Y3_W2BEG[6] ,
    \Tile_X4Y3_W2BEG[5] ,
    \Tile_X4Y3_W2BEG[4] ,
    \Tile_X4Y3_W2BEG[3] ,
    \Tile_X4Y3_W2BEG[2] ,
    \Tile_X4Y3_W2BEG[1] ,
    \Tile_X4Y3_W2BEG[0] }),
    .W6BEG({\Tile_X3Y3_W6BEG[11] ,
    \Tile_X3Y3_W6BEG[10] ,
    \Tile_X3Y3_W6BEG[9] ,
    \Tile_X3Y3_W6BEG[8] ,
    \Tile_X3Y3_W6BEG[7] ,
    \Tile_X3Y3_W6BEG[6] ,
    \Tile_X3Y3_W6BEG[5] ,
    \Tile_X3Y3_W6BEG[4] ,
    \Tile_X3Y3_W6BEG[3] ,
    \Tile_X3Y3_W6BEG[2] ,
    \Tile_X3Y3_W6BEG[1] ,
    \Tile_X3Y3_W6BEG[0] }),
    .W6END({\Tile_X4Y3_W6BEG[11] ,
    \Tile_X4Y3_W6BEG[10] ,
    \Tile_X4Y3_W6BEG[9] ,
    \Tile_X4Y3_W6BEG[8] ,
    \Tile_X4Y3_W6BEG[7] ,
    \Tile_X4Y3_W6BEG[6] ,
    \Tile_X4Y3_W6BEG[5] ,
    \Tile_X4Y3_W6BEG[4] ,
    \Tile_X4Y3_W6BEG[3] ,
    \Tile_X4Y3_W6BEG[2] ,
    \Tile_X4Y3_W6BEG[1] ,
    \Tile_X4Y3_W6BEG[0] }),
    .WW4BEG({\Tile_X3Y3_WW4BEG[15] ,
    \Tile_X3Y3_WW4BEG[14] ,
    \Tile_X3Y3_WW4BEG[13] ,
    \Tile_X3Y3_WW4BEG[12] ,
    \Tile_X3Y3_WW4BEG[11] ,
    \Tile_X3Y3_WW4BEG[10] ,
    \Tile_X3Y3_WW4BEG[9] ,
    \Tile_X3Y3_WW4BEG[8] ,
    \Tile_X3Y3_WW4BEG[7] ,
    \Tile_X3Y3_WW4BEG[6] ,
    \Tile_X3Y3_WW4BEG[5] ,
    \Tile_X3Y3_WW4BEG[4] ,
    \Tile_X3Y3_WW4BEG[3] ,
    \Tile_X3Y3_WW4BEG[2] ,
    \Tile_X3Y3_WW4BEG[1] ,
    \Tile_X3Y3_WW4BEG[0] }),
    .WW4END({\Tile_X4Y3_WW4BEG[15] ,
    \Tile_X4Y3_WW4BEG[14] ,
    \Tile_X4Y3_WW4BEG[13] ,
    \Tile_X4Y3_WW4BEG[12] ,
    \Tile_X4Y3_WW4BEG[11] ,
    \Tile_X4Y3_WW4BEG[10] ,
    \Tile_X4Y3_WW4BEG[9] ,
    \Tile_X4Y3_WW4BEG[8] ,
    \Tile_X4Y3_WW4BEG[7] ,
    \Tile_X4Y3_WW4BEG[6] ,
    \Tile_X4Y3_WW4BEG[5] ,
    \Tile_X4Y3_WW4BEG[4] ,
    \Tile_X4Y3_WW4BEG[3] ,
    \Tile_X4Y3_WW4BEG[2] ,
    \Tile_X4Y3_WW4BEG[1] ,
    \Tile_X4Y3_WW4BEG[0] }));
 LUT4AB Tile_X3Y4_LUT4AB (.Ci(Tile_X3Y5_Co),
    .Co(Tile_X3Y4_Co),
    .UserCLK(Tile_X3Y5_UserCLKo),
    .UserCLKo(Tile_X3Y4_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X3Y4_E1BEG[3] ,
    \Tile_X3Y4_E1BEG[2] ,
    \Tile_X3Y4_E1BEG[1] ,
    \Tile_X3Y4_E1BEG[0] }),
    .E1END({\Tile_X2Y4_E1BEG[3] ,
    \Tile_X2Y4_E1BEG[2] ,
    \Tile_X2Y4_E1BEG[1] ,
    \Tile_X2Y4_E1BEG[0] }),
    .E2BEG({\Tile_X3Y4_E2BEG[7] ,
    \Tile_X3Y4_E2BEG[6] ,
    \Tile_X3Y4_E2BEG[5] ,
    \Tile_X3Y4_E2BEG[4] ,
    \Tile_X3Y4_E2BEG[3] ,
    \Tile_X3Y4_E2BEG[2] ,
    \Tile_X3Y4_E2BEG[1] ,
    \Tile_X3Y4_E2BEG[0] }),
    .E2BEGb({\Tile_X3Y4_E2BEGb[7] ,
    \Tile_X3Y4_E2BEGb[6] ,
    \Tile_X3Y4_E2BEGb[5] ,
    \Tile_X3Y4_E2BEGb[4] ,
    \Tile_X3Y4_E2BEGb[3] ,
    \Tile_X3Y4_E2BEGb[2] ,
    \Tile_X3Y4_E2BEGb[1] ,
    \Tile_X3Y4_E2BEGb[0] }),
    .E2END({\Tile_X2Y4_E2BEGb[7] ,
    \Tile_X2Y4_E2BEGb[6] ,
    \Tile_X2Y4_E2BEGb[5] ,
    \Tile_X2Y4_E2BEGb[4] ,
    \Tile_X2Y4_E2BEGb[3] ,
    \Tile_X2Y4_E2BEGb[2] ,
    \Tile_X2Y4_E2BEGb[1] ,
    \Tile_X2Y4_E2BEGb[0] }),
    .E2MID({\Tile_X2Y4_E2BEG[7] ,
    \Tile_X2Y4_E2BEG[6] ,
    \Tile_X2Y4_E2BEG[5] ,
    \Tile_X2Y4_E2BEG[4] ,
    \Tile_X2Y4_E2BEG[3] ,
    \Tile_X2Y4_E2BEG[2] ,
    \Tile_X2Y4_E2BEG[1] ,
    \Tile_X2Y4_E2BEG[0] }),
    .E6BEG({\Tile_X3Y4_E6BEG[11] ,
    \Tile_X3Y4_E6BEG[10] ,
    \Tile_X3Y4_E6BEG[9] ,
    \Tile_X3Y4_E6BEG[8] ,
    \Tile_X3Y4_E6BEG[7] ,
    \Tile_X3Y4_E6BEG[6] ,
    \Tile_X3Y4_E6BEG[5] ,
    \Tile_X3Y4_E6BEG[4] ,
    \Tile_X3Y4_E6BEG[3] ,
    \Tile_X3Y4_E6BEG[2] ,
    \Tile_X3Y4_E6BEG[1] ,
    \Tile_X3Y4_E6BEG[0] }),
    .E6END({\Tile_X2Y4_E6BEG[11] ,
    \Tile_X2Y4_E6BEG[10] ,
    \Tile_X2Y4_E6BEG[9] ,
    \Tile_X2Y4_E6BEG[8] ,
    \Tile_X2Y4_E6BEG[7] ,
    \Tile_X2Y4_E6BEG[6] ,
    \Tile_X2Y4_E6BEG[5] ,
    \Tile_X2Y4_E6BEG[4] ,
    \Tile_X2Y4_E6BEG[3] ,
    \Tile_X2Y4_E6BEG[2] ,
    \Tile_X2Y4_E6BEG[1] ,
    \Tile_X2Y4_E6BEG[0] }),
    .EE4BEG({\Tile_X3Y4_EE4BEG[15] ,
    \Tile_X3Y4_EE4BEG[14] ,
    \Tile_X3Y4_EE4BEG[13] ,
    \Tile_X3Y4_EE4BEG[12] ,
    \Tile_X3Y4_EE4BEG[11] ,
    \Tile_X3Y4_EE4BEG[10] ,
    \Tile_X3Y4_EE4BEG[9] ,
    \Tile_X3Y4_EE4BEG[8] ,
    \Tile_X3Y4_EE4BEG[7] ,
    \Tile_X3Y4_EE4BEG[6] ,
    \Tile_X3Y4_EE4BEG[5] ,
    \Tile_X3Y4_EE4BEG[4] ,
    \Tile_X3Y4_EE4BEG[3] ,
    \Tile_X3Y4_EE4BEG[2] ,
    \Tile_X3Y4_EE4BEG[1] ,
    \Tile_X3Y4_EE4BEG[0] }),
    .EE4END({\Tile_X2Y4_EE4BEG[15] ,
    \Tile_X2Y4_EE4BEG[14] ,
    \Tile_X2Y4_EE4BEG[13] ,
    \Tile_X2Y4_EE4BEG[12] ,
    \Tile_X2Y4_EE4BEG[11] ,
    \Tile_X2Y4_EE4BEG[10] ,
    \Tile_X2Y4_EE4BEG[9] ,
    \Tile_X2Y4_EE4BEG[8] ,
    \Tile_X2Y4_EE4BEG[7] ,
    \Tile_X2Y4_EE4BEG[6] ,
    \Tile_X2Y4_EE4BEG[5] ,
    \Tile_X2Y4_EE4BEG[4] ,
    \Tile_X2Y4_EE4BEG[3] ,
    \Tile_X2Y4_EE4BEG[2] ,
    \Tile_X2Y4_EE4BEG[1] ,
    \Tile_X2Y4_EE4BEG[0] }),
    .FrameData({\Tile_X2Y4_FrameData_O[31] ,
    \Tile_X2Y4_FrameData_O[30] ,
    \Tile_X2Y4_FrameData_O[29] ,
    \Tile_X2Y4_FrameData_O[28] ,
    \Tile_X2Y4_FrameData_O[27] ,
    \Tile_X2Y4_FrameData_O[26] ,
    \Tile_X2Y4_FrameData_O[25] ,
    \Tile_X2Y4_FrameData_O[24] ,
    \Tile_X2Y4_FrameData_O[23] ,
    \Tile_X2Y4_FrameData_O[22] ,
    \Tile_X2Y4_FrameData_O[21] ,
    \Tile_X2Y4_FrameData_O[20] ,
    \Tile_X2Y4_FrameData_O[19] ,
    \Tile_X2Y4_FrameData_O[18] ,
    \Tile_X2Y4_FrameData_O[17] ,
    \Tile_X2Y4_FrameData_O[16] ,
    \Tile_X2Y4_FrameData_O[15] ,
    \Tile_X2Y4_FrameData_O[14] ,
    \Tile_X2Y4_FrameData_O[13] ,
    \Tile_X2Y4_FrameData_O[12] ,
    \Tile_X2Y4_FrameData_O[11] ,
    \Tile_X2Y4_FrameData_O[10] ,
    \Tile_X2Y4_FrameData_O[9] ,
    \Tile_X2Y4_FrameData_O[8] ,
    \Tile_X2Y4_FrameData_O[7] ,
    \Tile_X2Y4_FrameData_O[6] ,
    \Tile_X2Y4_FrameData_O[5] ,
    \Tile_X2Y4_FrameData_O[4] ,
    \Tile_X2Y4_FrameData_O[3] ,
    \Tile_X2Y4_FrameData_O[2] ,
    \Tile_X2Y4_FrameData_O[1] ,
    \Tile_X2Y4_FrameData_O[0] }),
    .FrameData_O({\Tile_X3Y4_FrameData_O[31] ,
    \Tile_X3Y4_FrameData_O[30] ,
    \Tile_X3Y4_FrameData_O[29] ,
    \Tile_X3Y4_FrameData_O[28] ,
    \Tile_X3Y4_FrameData_O[27] ,
    \Tile_X3Y4_FrameData_O[26] ,
    \Tile_X3Y4_FrameData_O[25] ,
    \Tile_X3Y4_FrameData_O[24] ,
    \Tile_X3Y4_FrameData_O[23] ,
    \Tile_X3Y4_FrameData_O[22] ,
    \Tile_X3Y4_FrameData_O[21] ,
    \Tile_X3Y4_FrameData_O[20] ,
    \Tile_X3Y4_FrameData_O[19] ,
    \Tile_X3Y4_FrameData_O[18] ,
    \Tile_X3Y4_FrameData_O[17] ,
    \Tile_X3Y4_FrameData_O[16] ,
    \Tile_X3Y4_FrameData_O[15] ,
    \Tile_X3Y4_FrameData_O[14] ,
    \Tile_X3Y4_FrameData_O[13] ,
    \Tile_X3Y4_FrameData_O[12] ,
    \Tile_X3Y4_FrameData_O[11] ,
    \Tile_X3Y4_FrameData_O[10] ,
    \Tile_X3Y4_FrameData_O[9] ,
    \Tile_X3Y4_FrameData_O[8] ,
    \Tile_X3Y4_FrameData_O[7] ,
    \Tile_X3Y4_FrameData_O[6] ,
    \Tile_X3Y4_FrameData_O[5] ,
    \Tile_X3Y4_FrameData_O[4] ,
    \Tile_X3Y4_FrameData_O[3] ,
    \Tile_X3Y4_FrameData_O[2] ,
    \Tile_X3Y4_FrameData_O[1] ,
    \Tile_X3Y4_FrameData_O[0] }),
    .FrameStrobe({\Tile_X3Y5_FrameStrobe_O[19] ,
    \Tile_X3Y5_FrameStrobe_O[18] ,
    \Tile_X3Y5_FrameStrobe_O[17] ,
    \Tile_X3Y5_FrameStrobe_O[16] ,
    \Tile_X3Y5_FrameStrobe_O[15] ,
    \Tile_X3Y5_FrameStrobe_O[14] ,
    \Tile_X3Y5_FrameStrobe_O[13] ,
    \Tile_X3Y5_FrameStrobe_O[12] ,
    \Tile_X3Y5_FrameStrobe_O[11] ,
    \Tile_X3Y5_FrameStrobe_O[10] ,
    \Tile_X3Y5_FrameStrobe_O[9] ,
    \Tile_X3Y5_FrameStrobe_O[8] ,
    \Tile_X3Y5_FrameStrobe_O[7] ,
    \Tile_X3Y5_FrameStrobe_O[6] ,
    \Tile_X3Y5_FrameStrobe_O[5] ,
    \Tile_X3Y5_FrameStrobe_O[4] ,
    \Tile_X3Y5_FrameStrobe_O[3] ,
    \Tile_X3Y5_FrameStrobe_O[2] ,
    \Tile_X3Y5_FrameStrobe_O[1] ,
    \Tile_X3Y5_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X3Y4_FrameStrobe_O[19] ,
    \Tile_X3Y4_FrameStrobe_O[18] ,
    \Tile_X3Y4_FrameStrobe_O[17] ,
    \Tile_X3Y4_FrameStrobe_O[16] ,
    \Tile_X3Y4_FrameStrobe_O[15] ,
    \Tile_X3Y4_FrameStrobe_O[14] ,
    \Tile_X3Y4_FrameStrobe_O[13] ,
    \Tile_X3Y4_FrameStrobe_O[12] ,
    \Tile_X3Y4_FrameStrobe_O[11] ,
    \Tile_X3Y4_FrameStrobe_O[10] ,
    \Tile_X3Y4_FrameStrobe_O[9] ,
    \Tile_X3Y4_FrameStrobe_O[8] ,
    \Tile_X3Y4_FrameStrobe_O[7] ,
    \Tile_X3Y4_FrameStrobe_O[6] ,
    \Tile_X3Y4_FrameStrobe_O[5] ,
    \Tile_X3Y4_FrameStrobe_O[4] ,
    \Tile_X3Y4_FrameStrobe_O[3] ,
    \Tile_X3Y4_FrameStrobe_O[2] ,
    \Tile_X3Y4_FrameStrobe_O[1] ,
    \Tile_X3Y4_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X3Y4_N1BEG[3] ,
    \Tile_X3Y4_N1BEG[2] ,
    \Tile_X3Y4_N1BEG[1] ,
    \Tile_X3Y4_N1BEG[0] }),
    .N1END({\Tile_X3Y5_N1BEG[3] ,
    \Tile_X3Y5_N1BEG[2] ,
    \Tile_X3Y5_N1BEG[1] ,
    \Tile_X3Y5_N1BEG[0] }),
    .N2BEG({\Tile_X3Y4_N2BEG[7] ,
    \Tile_X3Y4_N2BEG[6] ,
    \Tile_X3Y4_N2BEG[5] ,
    \Tile_X3Y4_N2BEG[4] ,
    \Tile_X3Y4_N2BEG[3] ,
    \Tile_X3Y4_N2BEG[2] ,
    \Tile_X3Y4_N2BEG[1] ,
    \Tile_X3Y4_N2BEG[0] }),
    .N2BEGb({\Tile_X3Y4_N2BEGb[7] ,
    \Tile_X3Y4_N2BEGb[6] ,
    \Tile_X3Y4_N2BEGb[5] ,
    \Tile_X3Y4_N2BEGb[4] ,
    \Tile_X3Y4_N2BEGb[3] ,
    \Tile_X3Y4_N2BEGb[2] ,
    \Tile_X3Y4_N2BEGb[1] ,
    \Tile_X3Y4_N2BEGb[0] }),
    .N2END({\Tile_X3Y5_N2BEGb[7] ,
    \Tile_X3Y5_N2BEGb[6] ,
    \Tile_X3Y5_N2BEGb[5] ,
    \Tile_X3Y5_N2BEGb[4] ,
    \Tile_X3Y5_N2BEGb[3] ,
    \Tile_X3Y5_N2BEGb[2] ,
    \Tile_X3Y5_N2BEGb[1] ,
    \Tile_X3Y5_N2BEGb[0] }),
    .N2MID({\Tile_X3Y5_N2BEG[7] ,
    \Tile_X3Y5_N2BEG[6] ,
    \Tile_X3Y5_N2BEG[5] ,
    \Tile_X3Y5_N2BEG[4] ,
    \Tile_X3Y5_N2BEG[3] ,
    \Tile_X3Y5_N2BEG[2] ,
    \Tile_X3Y5_N2BEG[1] ,
    \Tile_X3Y5_N2BEG[0] }),
    .N4BEG({\Tile_X3Y4_N4BEG[15] ,
    \Tile_X3Y4_N4BEG[14] ,
    \Tile_X3Y4_N4BEG[13] ,
    \Tile_X3Y4_N4BEG[12] ,
    \Tile_X3Y4_N4BEG[11] ,
    \Tile_X3Y4_N4BEG[10] ,
    \Tile_X3Y4_N4BEG[9] ,
    \Tile_X3Y4_N4BEG[8] ,
    \Tile_X3Y4_N4BEG[7] ,
    \Tile_X3Y4_N4BEG[6] ,
    \Tile_X3Y4_N4BEG[5] ,
    \Tile_X3Y4_N4BEG[4] ,
    \Tile_X3Y4_N4BEG[3] ,
    \Tile_X3Y4_N4BEG[2] ,
    \Tile_X3Y4_N4BEG[1] ,
    \Tile_X3Y4_N4BEG[0] }),
    .N4END({\Tile_X3Y5_N4BEG[15] ,
    \Tile_X3Y5_N4BEG[14] ,
    \Tile_X3Y5_N4BEG[13] ,
    \Tile_X3Y5_N4BEG[12] ,
    \Tile_X3Y5_N4BEG[11] ,
    \Tile_X3Y5_N4BEG[10] ,
    \Tile_X3Y5_N4BEG[9] ,
    \Tile_X3Y5_N4BEG[8] ,
    \Tile_X3Y5_N4BEG[7] ,
    \Tile_X3Y5_N4BEG[6] ,
    \Tile_X3Y5_N4BEG[5] ,
    \Tile_X3Y5_N4BEG[4] ,
    \Tile_X3Y5_N4BEG[3] ,
    \Tile_X3Y5_N4BEG[2] ,
    \Tile_X3Y5_N4BEG[1] ,
    \Tile_X3Y5_N4BEG[0] }),
    .NN4BEG({\Tile_X3Y4_NN4BEG[15] ,
    \Tile_X3Y4_NN4BEG[14] ,
    \Tile_X3Y4_NN4BEG[13] ,
    \Tile_X3Y4_NN4BEG[12] ,
    \Tile_X3Y4_NN4BEG[11] ,
    \Tile_X3Y4_NN4BEG[10] ,
    \Tile_X3Y4_NN4BEG[9] ,
    \Tile_X3Y4_NN4BEG[8] ,
    \Tile_X3Y4_NN4BEG[7] ,
    \Tile_X3Y4_NN4BEG[6] ,
    \Tile_X3Y4_NN4BEG[5] ,
    \Tile_X3Y4_NN4BEG[4] ,
    \Tile_X3Y4_NN4BEG[3] ,
    \Tile_X3Y4_NN4BEG[2] ,
    \Tile_X3Y4_NN4BEG[1] ,
    \Tile_X3Y4_NN4BEG[0] }),
    .NN4END({\Tile_X3Y5_NN4BEG[15] ,
    \Tile_X3Y5_NN4BEG[14] ,
    \Tile_X3Y5_NN4BEG[13] ,
    \Tile_X3Y5_NN4BEG[12] ,
    \Tile_X3Y5_NN4BEG[11] ,
    \Tile_X3Y5_NN4BEG[10] ,
    \Tile_X3Y5_NN4BEG[9] ,
    \Tile_X3Y5_NN4BEG[8] ,
    \Tile_X3Y5_NN4BEG[7] ,
    \Tile_X3Y5_NN4BEG[6] ,
    \Tile_X3Y5_NN4BEG[5] ,
    \Tile_X3Y5_NN4BEG[4] ,
    \Tile_X3Y5_NN4BEG[3] ,
    \Tile_X3Y5_NN4BEG[2] ,
    \Tile_X3Y5_NN4BEG[1] ,
    \Tile_X3Y5_NN4BEG[0] }),
    .S1BEG({\Tile_X3Y4_S1BEG[3] ,
    \Tile_X3Y4_S1BEG[2] ,
    \Tile_X3Y4_S1BEG[1] ,
    \Tile_X3Y4_S1BEG[0] }),
    .S1END({\Tile_X3Y3_S1BEG[3] ,
    \Tile_X3Y3_S1BEG[2] ,
    \Tile_X3Y3_S1BEG[1] ,
    \Tile_X3Y3_S1BEG[0] }),
    .S2BEG({\Tile_X3Y4_S2BEG[7] ,
    \Tile_X3Y4_S2BEG[6] ,
    \Tile_X3Y4_S2BEG[5] ,
    \Tile_X3Y4_S2BEG[4] ,
    \Tile_X3Y4_S2BEG[3] ,
    \Tile_X3Y4_S2BEG[2] ,
    \Tile_X3Y4_S2BEG[1] ,
    \Tile_X3Y4_S2BEG[0] }),
    .S2BEGb({\Tile_X3Y4_S2BEGb[7] ,
    \Tile_X3Y4_S2BEGb[6] ,
    \Tile_X3Y4_S2BEGb[5] ,
    \Tile_X3Y4_S2BEGb[4] ,
    \Tile_X3Y4_S2BEGb[3] ,
    \Tile_X3Y4_S2BEGb[2] ,
    \Tile_X3Y4_S2BEGb[1] ,
    \Tile_X3Y4_S2BEGb[0] }),
    .S2END({\Tile_X3Y3_S2BEGb[7] ,
    \Tile_X3Y3_S2BEGb[6] ,
    \Tile_X3Y3_S2BEGb[5] ,
    \Tile_X3Y3_S2BEGb[4] ,
    \Tile_X3Y3_S2BEGb[3] ,
    \Tile_X3Y3_S2BEGb[2] ,
    \Tile_X3Y3_S2BEGb[1] ,
    \Tile_X3Y3_S2BEGb[0] }),
    .S2MID({\Tile_X3Y3_S2BEG[7] ,
    \Tile_X3Y3_S2BEG[6] ,
    \Tile_X3Y3_S2BEG[5] ,
    \Tile_X3Y3_S2BEG[4] ,
    \Tile_X3Y3_S2BEG[3] ,
    \Tile_X3Y3_S2BEG[2] ,
    \Tile_X3Y3_S2BEG[1] ,
    \Tile_X3Y3_S2BEG[0] }),
    .S4BEG({\Tile_X3Y4_S4BEG[15] ,
    \Tile_X3Y4_S4BEG[14] ,
    \Tile_X3Y4_S4BEG[13] ,
    \Tile_X3Y4_S4BEG[12] ,
    \Tile_X3Y4_S4BEG[11] ,
    \Tile_X3Y4_S4BEG[10] ,
    \Tile_X3Y4_S4BEG[9] ,
    \Tile_X3Y4_S4BEG[8] ,
    \Tile_X3Y4_S4BEG[7] ,
    \Tile_X3Y4_S4BEG[6] ,
    \Tile_X3Y4_S4BEG[5] ,
    \Tile_X3Y4_S4BEG[4] ,
    \Tile_X3Y4_S4BEG[3] ,
    \Tile_X3Y4_S4BEG[2] ,
    \Tile_X3Y4_S4BEG[1] ,
    \Tile_X3Y4_S4BEG[0] }),
    .S4END({\Tile_X3Y3_S4BEG[15] ,
    \Tile_X3Y3_S4BEG[14] ,
    \Tile_X3Y3_S4BEG[13] ,
    \Tile_X3Y3_S4BEG[12] ,
    \Tile_X3Y3_S4BEG[11] ,
    \Tile_X3Y3_S4BEG[10] ,
    \Tile_X3Y3_S4BEG[9] ,
    \Tile_X3Y3_S4BEG[8] ,
    \Tile_X3Y3_S4BEG[7] ,
    \Tile_X3Y3_S4BEG[6] ,
    \Tile_X3Y3_S4BEG[5] ,
    \Tile_X3Y3_S4BEG[4] ,
    \Tile_X3Y3_S4BEG[3] ,
    \Tile_X3Y3_S4BEG[2] ,
    \Tile_X3Y3_S4BEG[1] ,
    \Tile_X3Y3_S4BEG[0] }),
    .SS4BEG({\Tile_X3Y4_SS4BEG[15] ,
    \Tile_X3Y4_SS4BEG[14] ,
    \Tile_X3Y4_SS4BEG[13] ,
    \Tile_X3Y4_SS4BEG[12] ,
    \Tile_X3Y4_SS4BEG[11] ,
    \Tile_X3Y4_SS4BEG[10] ,
    \Tile_X3Y4_SS4BEG[9] ,
    \Tile_X3Y4_SS4BEG[8] ,
    \Tile_X3Y4_SS4BEG[7] ,
    \Tile_X3Y4_SS4BEG[6] ,
    \Tile_X3Y4_SS4BEG[5] ,
    \Tile_X3Y4_SS4BEG[4] ,
    \Tile_X3Y4_SS4BEG[3] ,
    \Tile_X3Y4_SS4BEG[2] ,
    \Tile_X3Y4_SS4BEG[1] ,
    \Tile_X3Y4_SS4BEG[0] }),
    .SS4END({\Tile_X3Y3_SS4BEG[15] ,
    \Tile_X3Y3_SS4BEG[14] ,
    \Tile_X3Y3_SS4BEG[13] ,
    \Tile_X3Y3_SS4BEG[12] ,
    \Tile_X3Y3_SS4BEG[11] ,
    \Tile_X3Y3_SS4BEG[10] ,
    \Tile_X3Y3_SS4BEG[9] ,
    \Tile_X3Y3_SS4BEG[8] ,
    \Tile_X3Y3_SS4BEG[7] ,
    \Tile_X3Y3_SS4BEG[6] ,
    \Tile_X3Y3_SS4BEG[5] ,
    \Tile_X3Y3_SS4BEG[4] ,
    \Tile_X3Y3_SS4BEG[3] ,
    \Tile_X3Y3_SS4BEG[2] ,
    \Tile_X3Y3_SS4BEG[1] ,
    \Tile_X3Y3_SS4BEG[0] }),
    .W1BEG({\Tile_X3Y4_W1BEG[3] ,
    \Tile_X3Y4_W1BEG[2] ,
    \Tile_X3Y4_W1BEG[1] ,
    \Tile_X3Y4_W1BEG[0] }),
    .W1END({\Tile_X4Y4_W1BEG[3] ,
    \Tile_X4Y4_W1BEG[2] ,
    \Tile_X4Y4_W1BEG[1] ,
    \Tile_X4Y4_W1BEG[0] }),
    .W2BEG({\Tile_X3Y4_W2BEG[7] ,
    \Tile_X3Y4_W2BEG[6] ,
    \Tile_X3Y4_W2BEG[5] ,
    \Tile_X3Y4_W2BEG[4] ,
    \Tile_X3Y4_W2BEG[3] ,
    \Tile_X3Y4_W2BEG[2] ,
    \Tile_X3Y4_W2BEG[1] ,
    \Tile_X3Y4_W2BEG[0] }),
    .W2BEGb({\Tile_X3Y4_W2BEGb[7] ,
    \Tile_X3Y4_W2BEGb[6] ,
    \Tile_X3Y4_W2BEGb[5] ,
    \Tile_X3Y4_W2BEGb[4] ,
    \Tile_X3Y4_W2BEGb[3] ,
    \Tile_X3Y4_W2BEGb[2] ,
    \Tile_X3Y4_W2BEGb[1] ,
    \Tile_X3Y4_W2BEGb[0] }),
    .W2END({\Tile_X4Y4_W2BEGb[7] ,
    \Tile_X4Y4_W2BEGb[6] ,
    \Tile_X4Y4_W2BEGb[5] ,
    \Tile_X4Y4_W2BEGb[4] ,
    \Tile_X4Y4_W2BEGb[3] ,
    \Tile_X4Y4_W2BEGb[2] ,
    \Tile_X4Y4_W2BEGb[1] ,
    \Tile_X4Y4_W2BEGb[0] }),
    .W2MID({\Tile_X4Y4_W2BEG[7] ,
    \Tile_X4Y4_W2BEG[6] ,
    \Tile_X4Y4_W2BEG[5] ,
    \Tile_X4Y4_W2BEG[4] ,
    \Tile_X4Y4_W2BEG[3] ,
    \Tile_X4Y4_W2BEG[2] ,
    \Tile_X4Y4_W2BEG[1] ,
    \Tile_X4Y4_W2BEG[0] }),
    .W6BEG({\Tile_X3Y4_W6BEG[11] ,
    \Tile_X3Y4_W6BEG[10] ,
    \Tile_X3Y4_W6BEG[9] ,
    \Tile_X3Y4_W6BEG[8] ,
    \Tile_X3Y4_W6BEG[7] ,
    \Tile_X3Y4_W6BEG[6] ,
    \Tile_X3Y4_W6BEG[5] ,
    \Tile_X3Y4_W6BEG[4] ,
    \Tile_X3Y4_W6BEG[3] ,
    \Tile_X3Y4_W6BEG[2] ,
    \Tile_X3Y4_W6BEG[1] ,
    \Tile_X3Y4_W6BEG[0] }),
    .W6END({\Tile_X4Y4_W6BEG[11] ,
    \Tile_X4Y4_W6BEG[10] ,
    \Tile_X4Y4_W6BEG[9] ,
    \Tile_X4Y4_W6BEG[8] ,
    \Tile_X4Y4_W6BEG[7] ,
    \Tile_X4Y4_W6BEG[6] ,
    \Tile_X4Y4_W6BEG[5] ,
    \Tile_X4Y4_W6BEG[4] ,
    \Tile_X4Y4_W6BEG[3] ,
    \Tile_X4Y4_W6BEG[2] ,
    \Tile_X4Y4_W6BEG[1] ,
    \Tile_X4Y4_W6BEG[0] }),
    .WW4BEG({\Tile_X3Y4_WW4BEG[15] ,
    \Tile_X3Y4_WW4BEG[14] ,
    \Tile_X3Y4_WW4BEG[13] ,
    \Tile_X3Y4_WW4BEG[12] ,
    \Tile_X3Y4_WW4BEG[11] ,
    \Tile_X3Y4_WW4BEG[10] ,
    \Tile_X3Y4_WW4BEG[9] ,
    \Tile_X3Y4_WW4BEG[8] ,
    \Tile_X3Y4_WW4BEG[7] ,
    \Tile_X3Y4_WW4BEG[6] ,
    \Tile_X3Y4_WW4BEG[5] ,
    \Tile_X3Y4_WW4BEG[4] ,
    \Tile_X3Y4_WW4BEG[3] ,
    \Tile_X3Y4_WW4BEG[2] ,
    \Tile_X3Y4_WW4BEG[1] ,
    \Tile_X3Y4_WW4BEG[0] }),
    .WW4END({\Tile_X4Y4_WW4BEG[15] ,
    \Tile_X4Y4_WW4BEG[14] ,
    \Tile_X4Y4_WW4BEG[13] ,
    \Tile_X4Y4_WW4BEG[12] ,
    \Tile_X4Y4_WW4BEG[11] ,
    \Tile_X4Y4_WW4BEG[10] ,
    \Tile_X4Y4_WW4BEG[9] ,
    \Tile_X4Y4_WW4BEG[8] ,
    \Tile_X4Y4_WW4BEG[7] ,
    \Tile_X4Y4_WW4BEG[6] ,
    \Tile_X4Y4_WW4BEG[5] ,
    \Tile_X4Y4_WW4BEG[4] ,
    \Tile_X4Y4_WW4BEG[3] ,
    \Tile_X4Y4_WW4BEG[2] ,
    \Tile_X4Y4_WW4BEG[1] ,
    \Tile_X4Y4_WW4BEG[0] }));
 LUT4AB Tile_X3Y5_LUT4AB (.Ci(Tile_X3Y6_Co),
    .Co(Tile_X3Y5_Co),
    .UserCLK(Tile_X3Y6_UserCLKo),
    .UserCLKo(Tile_X3Y5_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X3Y5_E1BEG[3] ,
    \Tile_X3Y5_E1BEG[2] ,
    \Tile_X3Y5_E1BEG[1] ,
    \Tile_X3Y5_E1BEG[0] }),
    .E1END({\Tile_X2Y5_E1BEG[3] ,
    \Tile_X2Y5_E1BEG[2] ,
    \Tile_X2Y5_E1BEG[1] ,
    \Tile_X2Y5_E1BEG[0] }),
    .E2BEG({\Tile_X3Y5_E2BEG[7] ,
    \Tile_X3Y5_E2BEG[6] ,
    \Tile_X3Y5_E2BEG[5] ,
    \Tile_X3Y5_E2BEG[4] ,
    \Tile_X3Y5_E2BEG[3] ,
    \Tile_X3Y5_E2BEG[2] ,
    \Tile_X3Y5_E2BEG[1] ,
    \Tile_X3Y5_E2BEG[0] }),
    .E2BEGb({\Tile_X3Y5_E2BEGb[7] ,
    \Tile_X3Y5_E2BEGb[6] ,
    \Tile_X3Y5_E2BEGb[5] ,
    \Tile_X3Y5_E2BEGb[4] ,
    \Tile_X3Y5_E2BEGb[3] ,
    \Tile_X3Y5_E2BEGb[2] ,
    \Tile_X3Y5_E2BEGb[1] ,
    \Tile_X3Y5_E2BEGb[0] }),
    .E2END({\Tile_X2Y5_E2BEGb[7] ,
    \Tile_X2Y5_E2BEGb[6] ,
    \Tile_X2Y5_E2BEGb[5] ,
    \Tile_X2Y5_E2BEGb[4] ,
    \Tile_X2Y5_E2BEGb[3] ,
    \Tile_X2Y5_E2BEGb[2] ,
    \Tile_X2Y5_E2BEGb[1] ,
    \Tile_X2Y5_E2BEGb[0] }),
    .E2MID({\Tile_X2Y5_E2BEG[7] ,
    \Tile_X2Y5_E2BEG[6] ,
    \Tile_X2Y5_E2BEG[5] ,
    \Tile_X2Y5_E2BEG[4] ,
    \Tile_X2Y5_E2BEG[3] ,
    \Tile_X2Y5_E2BEG[2] ,
    \Tile_X2Y5_E2BEG[1] ,
    \Tile_X2Y5_E2BEG[0] }),
    .E6BEG({\Tile_X3Y5_E6BEG[11] ,
    \Tile_X3Y5_E6BEG[10] ,
    \Tile_X3Y5_E6BEG[9] ,
    \Tile_X3Y5_E6BEG[8] ,
    \Tile_X3Y5_E6BEG[7] ,
    \Tile_X3Y5_E6BEG[6] ,
    \Tile_X3Y5_E6BEG[5] ,
    \Tile_X3Y5_E6BEG[4] ,
    \Tile_X3Y5_E6BEG[3] ,
    \Tile_X3Y5_E6BEG[2] ,
    \Tile_X3Y5_E6BEG[1] ,
    \Tile_X3Y5_E6BEG[0] }),
    .E6END({\Tile_X2Y5_E6BEG[11] ,
    \Tile_X2Y5_E6BEG[10] ,
    \Tile_X2Y5_E6BEG[9] ,
    \Tile_X2Y5_E6BEG[8] ,
    \Tile_X2Y5_E6BEG[7] ,
    \Tile_X2Y5_E6BEG[6] ,
    \Tile_X2Y5_E6BEG[5] ,
    \Tile_X2Y5_E6BEG[4] ,
    \Tile_X2Y5_E6BEG[3] ,
    \Tile_X2Y5_E6BEG[2] ,
    \Tile_X2Y5_E6BEG[1] ,
    \Tile_X2Y5_E6BEG[0] }),
    .EE4BEG({\Tile_X3Y5_EE4BEG[15] ,
    \Tile_X3Y5_EE4BEG[14] ,
    \Tile_X3Y5_EE4BEG[13] ,
    \Tile_X3Y5_EE4BEG[12] ,
    \Tile_X3Y5_EE4BEG[11] ,
    \Tile_X3Y5_EE4BEG[10] ,
    \Tile_X3Y5_EE4BEG[9] ,
    \Tile_X3Y5_EE4BEG[8] ,
    \Tile_X3Y5_EE4BEG[7] ,
    \Tile_X3Y5_EE4BEG[6] ,
    \Tile_X3Y5_EE4BEG[5] ,
    \Tile_X3Y5_EE4BEG[4] ,
    \Tile_X3Y5_EE4BEG[3] ,
    \Tile_X3Y5_EE4BEG[2] ,
    \Tile_X3Y5_EE4BEG[1] ,
    \Tile_X3Y5_EE4BEG[0] }),
    .EE4END({\Tile_X2Y5_EE4BEG[15] ,
    \Tile_X2Y5_EE4BEG[14] ,
    \Tile_X2Y5_EE4BEG[13] ,
    \Tile_X2Y5_EE4BEG[12] ,
    \Tile_X2Y5_EE4BEG[11] ,
    \Tile_X2Y5_EE4BEG[10] ,
    \Tile_X2Y5_EE4BEG[9] ,
    \Tile_X2Y5_EE4BEG[8] ,
    \Tile_X2Y5_EE4BEG[7] ,
    \Tile_X2Y5_EE4BEG[6] ,
    \Tile_X2Y5_EE4BEG[5] ,
    \Tile_X2Y5_EE4BEG[4] ,
    \Tile_X2Y5_EE4BEG[3] ,
    \Tile_X2Y5_EE4BEG[2] ,
    \Tile_X2Y5_EE4BEG[1] ,
    \Tile_X2Y5_EE4BEG[0] }),
    .FrameData({\Tile_X2Y5_FrameData_O[31] ,
    \Tile_X2Y5_FrameData_O[30] ,
    \Tile_X2Y5_FrameData_O[29] ,
    \Tile_X2Y5_FrameData_O[28] ,
    \Tile_X2Y5_FrameData_O[27] ,
    \Tile_X2Y5_FrameData_O[26] ,
    \Tile_X2Y5_FrameData_O[25] ,
    \Tile_X2Y5_FrameData_O[24] ,
    \Tile_X2Y5_FrameData_O[23] ,
    \Tile_X2Y5_FrameData_O[22] ,
    \Tile_X2Y5_FrameData_O[21] ,
    \Tile_X2Y5_FrameData_O[20] ,
    \Tile_X2Y5_FrameData_O[19] ,
    \Tile_X2Y5_FrameData_O[18] ,
    \Tile_X2Y5_FrameData_O[17] ,
    \Tile_X2Y5_FrameData_O[16] ,
    \Tile_X2Y5_FrameData_O[15] ,
    \Tile_X2Y5_FrameData_O[14] ,
    \Tile_X2Y5_FrameData_O[13] ,
    \Tile_X2Y5_FrameData_O[12] ,
    \Tile_X2Y5_FrameData_O[11] ,
    \Tile_X2Y5_FrameData_O[10] ,
    \Tile_X2Y5_FrameData_O[9] ,
    \Tile_X2Y5_FrameData_O[8] ,
    \Tile_X2Y5_FrameData_O[7] ,
    \Tile_X2Y5_FrameData_O[6] ,
    \Tile_X2Y5_FrameData_O[5] ,
    \Tile_X2Y5_FrameData_O[4] ,
    \Tile_X2Y5_FrameData_O[3] ,
    \Tile_X2Y5_FrameData_O[2] ,
    \Tile_X2Y5_FrameData_O[1] ,
    \Tile_X2Y5_FrameData_O[0] }),
    .FrameData_O({\Tile_X3Y5_FrameData_O[31] ,
    \Tile_X3Y5_FrameData_O[30] ,
    \Tile_X3Y5_FrameData_O[29] ,
    \Tile_X3Y5_FrameData_O[28] ,
    \Tile_X3Y5_FrameData_O[27] ,
    \Tile_X3Y5_FrameData_O[26] ,
    \Tile_X3Y5_FrameData_O[25] ,
    \Tile_X3Y5_FrameData_O[24] ,
    \Tile_X3Y5_FrameData_O[23] ,
    \Tile_X3Y5_FrameData_O[22] ,
    \Tile_X3Y5_FrameData_O[21] ,
    \Tile_X3Y5_FrameData_O[20] ,
    \Tile_X3Y5_FrameData_O[19] ,
    \Tile_X3Y5_FrameData_O[18] ,
    \Tile_X3Y5_FrameData_O[17] ,
    \Tile_X3Y5_FrameData_O[16] ,
    \Tile_X3Y5_FrameData_O[15] ,
    \Tile_X3Y5_FrameData_O[14] ,
    \Tile_X3Y5_FrameData_O[13] ,
    \Tile_X3Y5_FrameData_O[12] ,
    \Tile_X3Y5_FrameData_O[11] ,
    \Tile_X3Y5_FrameData_O[10] ,
    \Tile_X3Y5_FrameData_O[9] ,
    \Tile_X3Y5_FrameData_O[8] ,
    \Tile_X3Y5_FrameData_O[7] ,
    \Tile_X3Y5_FrameData_O[6] ,
    \Tile_X3Y5_FrameData_O[5] ,
    \Tile_X3Y5_FrameData_O[4] ,
    \Tile_X3Y5_FrameData_O[3] ,
    \Tile_X3Y5_FrameData_O[2] ,
    \Tile_X3Y5_FrameData_O[1] ,
    \Tile_X3Y5_FrameData_O[0] }),
    .FrameStrobe({\Tile_X3Y6_FrameStrobe_O[19] ,
    \Tile_X3Y6_FrameStrobe_O[18] ,
    \Tile_X3Y6_FrameStrobe_O[17] ,
    \Tile_X3Y6_FrameStrobe_O[16] ,
    \Tile_X3Y6_FrameStrobe_O[15] ,
    \Tile_X3Y6_FrameStrobe_O[14] ,
    \Tile_X3Y6_FrameStrobe_O[13] ,
    \Tile_X3Y6_FrameStrobe_O[12] ,
    \Tile_X3Y6_FrameStrobe_O[11] ,
    \Tile_X3Y6_FrameStrobe_O[10] ,
    \Tile_X3Y6_FrameStrobe_O[9] ,
    \Tile_X3Y6_FrameStrobe_O[8] ,
    \Tile_X3Y6_FrameStrobe_O[7] ,
    \Tile_X3Y6_FrameStrobe_O[6] ,
    \Tile_X3Y6_FrameStrobe_O[5] ,
    \Tile_X3Y6_FrameStrobe_O[4] ,
    \Tile_X3Y6_FrameStrobe_O[3] ,
    \Tile_X3Y6_FrameStrobe_O[2] ,
    \Tile_X3Y6_FrameStrobe_O[1] ,
    \Tile_X3Y6_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X3Y5_FrameStrobe_O[19] ,
    \Tile_X3Y5_FrameStrobe_O[18] ,
    \Tile_X3Y5_FrameStrobe_O[17] ,
    \Tile_X3Y5_FrameStrobe_O[16] ,
    \Tile_X3Y5_FrameStrobe_O[15] ,
    \Tile_X3Y5_FrameStrobe_O[14] ,
    \Tile_X3Y5_FrameStrobe_O[13] ,
    \Tile_X3Y5_FrameStrobe_O[12] ,
    \Tile_X3Y5_FrameStrobe_O[11] ,
    \Tile_X3Y5_FrameStrobe_O[10] ,
    \Tile_X3Y5_FrameStrobe_O[9] ,
    \Tile_X3Y5_FrameStrobe_O[8] ,
    \Tile_X3Y5_FrameStrobe_O[7] ,
    \Tile_X3Y5_FrameStrobe_O[6] ,
    \Tile_X3Y5_FrameStrobe_O[5] ,
    \Tile_X3Y5_FrameStrobe_O[4] ,
    \Tile_X3Y5_FrameStrobe_O[3] ,
    \Tile_X3Y5_FrameStrobe_O[2] ,
    \Tile_X3Y5_FrameStrobe_O[1] ,
    \Tile_X3Y5_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X3Y5_N1BEG[3] ,
    \Tile_X3Y5_N1BEG[2] ,
    \Tile_X3Y5_N1BEG[1] ,
    \Tile_X3Y5_N1BEG[0] }),
    .N1END({\Tile_X3Y6_N1BEG[3] ,
    \Tile_X3Y6_N1BEG[2] ,
    \Tile_X3Y6_N1BEG[1] ,
    \Tile_X3Y6_N1BEG[0] }),
    .N2BEG({\Tile_X3Y5_N2BEG[7] ,
    \Tile_X3Y5_N2BEG[6] ,
    \Tile_X3Y5_N2BEG[5] ,
    \Tile_X3Y5_N2BEG[4] ,
    \Tile_X3Y5_N2BEG[3] ,
    \Tile_X3Y5_N2BEG[2] ,
    \Tile_X3Y5_N2BEG[1] ,
    \Tile_X3Y5_N2BEG[0] }),
    .N2BEGb({\Tile_X3Y5_N2BEGb[7] ,
    \Tile_X3Y5_N2BEGb[6] ,
    \Tile_X3Y5_N2BEGb[5] ,
    \Tile_X3Y5_N2BEGb[4] ,
    \Tile_X3Y5_N2BEGb[3] ,
    \Tile_X3Y5_N2BEGb[2] ,
    \Tile_X3Y5_N2BEGb[1] ,
    \Tile_X3Y5_N2BEGb[0] }),
    .N2END({\Tile_X3Y6_N2BEGb[7] ,
    \Tile_X3Y6_N2BEGb[6] ,
    \Tile_X3Y6_N2BEGb[5] ,
    \Tile_X3Y6_N2BEGb[4] ,
    \Tile_X3Y6_N2BEGb[3] ,
    \Tile_X3Y6_N2BEGb[2] ,
    \Tile_X3Y6_N2BEGb[1] ,
    \Tile_X3Y6_N2BEGb[0] }),
    .N2MID({\Tile_X3Y6_N2BEG[7] ,
    \Tile_X3Y6_N2BEG[6] ,
    \Tile_X3Y6_N2BEG[5] ,
    \Tile_X3Y6_N2BEG[4] ,
    \Tile_X3Y6_N2BEG[3] ,
    \Tile_X3Y6_N2BEG[2] ,
    \Tile_X3Y6_N2BEG[1] ,
    \Tile_X3Y6_N2BEG[0] }),
    .N4BEG({\Tile_X3Y5_N4BEG[15] ,
    \Tile_X3Y5_N4BEG[14] ,
    \Tile_X3Y5_N4BEG[13] ,
    \Tile_X3Y5_N4BEG[12] ,
    \Tile_X3Y5_N4BEG[11] ,
    \Tile_X3Y5_N4BEG[10] ,
    \Tile_X3Y5_N4BEG[9] ,
    \Tile_X3Y5_N4BEG[8] ,
    \Tile_X3Y5_N4BEG[7] ,
    \Tile_X3Y5_N4BEG[6] ,
    \Tile_X3Y5_N4BEG[5] ,
    \Tile_X3Y5_N4BEG[4] ,
    \Tile_X3Y5_N4BEG[3] ,
    \Tile_X3Y5_N4BEG[2] ,
    \Tile_X3Y5_N4BEG[1] ,
    \Tile_X3Y5_N4BEG[0] }),
    .N4END({\Tile_X3Y6_N4BEG[15] ,
    \Tile_X3Y6_N4BEG[14] ,
    \Tile_X3Y6_N4BEG[13] ,
    \Tile_X3Y6_N4BEG[12] ,
    \Tile_X3Y6_N4BEG[11] ,
    \Tile_X3Y6_N4BEG[10] ,
    \Tile_X3Y6_N4BEG[9] ,
    \Tile_X3Y6_N4BEG[8] ,
    \Tile_X3Y6_N4BEG[7] ,
    \Tile_X3Y6_N4BEG[6] ,
    \Tile_X3Y6_N4BEG[5] ,
    \Tile_X3Y6_N4BEG[4] ,
    \Tile_X3Y6_N4BEG[3] ,
    \Tile_X3Y6_N4BEG[2] ,
    \Tile_X3Y6_N4BEG[1] ,
    \Tile_X3Y6_N4BEG[0] }),
    .NN4BEG({\Tile_X3Y5_NN4BEG[15] ,
    \Tile_X3Y5_NN4BEG[14] ,
    \Tile_X3Y5_NN4BEG[13] ,
    \Tile_X3Y5_NN4BEG[12] ,
    \Tile_X3Y5_NN4BEG[11] ,
    \Tile_X3Y5_NN4BEG[10] ,
    \Tile_X3Y5_NN4BEG[9] ,
    \Tile_X3Y5_NN4BEG[8] ,
    \Tile_X3Y5_NN4BEG[7] ,
    \Tile_X3Y5_NN4BEG[6] ,
    \Tile_X3Y5_NN4BEG[5] ,
    \Tile_X3Y5_NN4BEG[4] ,
    \Tile_X3Y5_NN4BEG[3] ,
    \Tile_X3Y5_NN4BEG[2] ,
    \Tile_X3Y5_NN4BEG[1] ,
    \Tile_X3Y5_NN4BEG[0] }),
    .NN4END({\Tile_X3Y6_NN4BEG[15] ,
    \Tile_X3Y6_NN4BEG[14] ,
    \Tile_X3Y6_NN4BEG[13] ,
    \Tile_X3Y6_NN4BEG[12] ,
    \Tile_X3Y6_NN4BEG[11] ,
    \Tile_X3Y6_NN4BEG[10] ,
    \Tile_X3Y6_NN4BEG[9] ,
    \Tile_X3Y6_NN4BEG[8] ,
    \Tile_X3Y6_NN4BEG[7] ,
    \Tile_X3Y6_NN4BEG[6] ,
    \Tile_X3Y6_NN4BEG[5] ,
    \Tile_X3Y6_NN4BEG[4] ,
    \Tile_X3Y6_NN4BEG[3] ,
    \Tile_X3Y6_NN4BEG[2] ,
    \Tile_X3Y6_NN4BEG[1] ,
    \Tile_X3Y6_NN4BEG[0] }),
    .S1BEG({\Tile_X3Y5_S1BEG[3] ,
    \Tile_X3Y5_S1BEG[2] ,
    \Tile_X3Y5_S1BEG[1] ,
    \Tile_X3Y5_S1BEG[0] }),
    .S1END({\Tile_X3Y4_S1BEG[3] ,
    \Tile_X3Y4_S1BEG[2] ,
    \Tile_X3Y4_S1BEG[1] ,
    \Tile_X3Y4_S1BEG[0] }),
    .S2BEG({\Tile_X3Y5_S2BEG[7] ,
    \Tile_X3Y5_S2BEG[6] ,
    \Tile_X3Y5_S2BEG[5] ,
    \Tile_X3Y5_S2BEG[4] ,
    \Tile_X3Y5_S2BEG[3] ,
    \Tile_X3Y5_S2BEG[2] ,
    \Tile_X3Y5_S2BEG[1] ,
    \Tile_X3Y5_S2BEG[0] }),
    .S2BEGb({\Tile_X3Y5_S2BEGb[7] ,
    \Tile_X3Y5_S2BEGb[6] ,
    \Tile_X3Y5_S2BEGb[5] ,
    \Tile_X3Y5_S2BEGb[4] ,
    \Tile_X3Y5_S2BEGb[3] ,
    \Tile_X3Y5_S2BEGb[2] ,
    \Tile_X3Y5_S2BEGb[1] ,
    \Tile_X3Y5_S2BEGb[0] }),
    .S2END({\Tile_X3Y4_S2BEGb[7] ,
    \Tile_X3Y4_S2BEGb[6] ,
    \Tile_X3Y4_S2BEGb[5] ,
    \Tile_X3Y4_S2BEGb[4] ,
    \Tile_X3Y4_S2BEGb[3] ,
    \Tile_X3Y4_S2BEGb[2] ,
    \Tile_X3Y4_S2BEGb[1] ,
    \Tile_X3Y4_S2BEGb[0] }),
    .S2MID({\Tile_X3Y4_S2BEG[7] ,
    \Tile_X3Y4_S2BEG[6] ,
    \Tile_X3Y4_S2BEG[5] ,
    \Tile_X3Y4_S2BEG[4] ,
    \Tile_X3Y4_S2BEG[3] ,
    \Tile_X3Y4_S2BEG[2] ,
    \Tile_X3Y4_S2BEG[1] ,
    \Tile_X3Y4_S2BEG[0] }),
    .S4BEG({\Tile_X3Y5_S4BEG[15] ,
    \Tile_X3Y5_S4BEG[14] ,
    \Tile_X3Y5_S4BEG[13] ,
    \Tile_X3Y5_S4BEG[12] ,
    \Tile_X3Y5_S4BEG[11] ,
    \Tile_X3Y5_S4BEG[10] ,
    \Tile_X3Y5_S4BEG[9] ,
    \Tile_X3Y5_S4BEG[8] ,
    \Tile_X3Y5_S4BEG[7] ,
    \Tile_X3Y5_S4BEG[6] ,
    \Tile_X3Y5_S4BEG[5] ,
    \Tile_X3Y5_S4BEG[4] ,
    \Tile_X3Y5_S4BEG[3] ,
    \Tile_X3Y5_S4BEG[2] ,
    \Tile_X3Y5_S4BEG[1] ,
    \Tile_X3Y5_S4BEG[0] }),
    .S4END({\Tile_X3Y4_S4BEG[15] ,
    \Tile_X3Y4_S4BEG[14] ,
    \Tile_X3Y4_S4BEG[13] ,
    \Tile_X3Y4_S4BEG[12] ,
    \Tile_X3Y4_S4BEG[11] ,
    \Tile_X3Y4_S4BEG[10] ,
    \Tile_X3Y4_S4BEG[9] ,
    \Tile_X3Y4_S4BEG[8] ,
    \Tile_X3Y4_S4BEG[7] ,
    \Tile_X3Y4_S4BEG[6] ,
    \Tile_X3Y4_S4BEG[5] ,
    \Tile_X3Y4_S4BEG[4] ,
    \Tile_X3Y4_S4BEG[3] ,
    \Tile_X3Y4_S4BEG[2] ,
    \Tile_X3Y4_S4BEG[1] ,
    \Tile_X3Y4_S4BEG[0] }),
    .SS4BEG({\Tile_X3Y5_SS4BEG[15] ,
    \Tile_X3Y5_SS4BEG[14] ,
    \Tile_X3Y5_SS4BEG[13] ,
    \Tile_X3Y5_SS4BEG[12] ,
    \Tile_X3Y5_SS4BEG[11] ,
    \Tile_X3Y5_SS4BEG[10] ,
    \Tile_X3Y5_SS4BEG[9] ,
    \Tile_X3Y5_SS4BEG[8] ,
    \Tile_X3Y5_SS4BEG[7] ,
    \Tile_X3Y5_SS4BEG[6] ,
    \Tile_X3Y5_SS4BEG[5] ,
    \Tile_X3Y5_SS4BEG[4] ,
    \Tile_X3Y5_SS4BEG[3] ,
    \Tile_X3Y5_SS4BEG[2] ,
    \Tile_X3Y5_SS4BEG[1] ,
    \Tile_X3Y5_SS4BEG[0] }),
    .SS4END({\Tile_X3Y4_SS4BEG[15] ,
    \Tile_X3Y4_SS4BEG[14] ,
    \Tile_X3Y4_SS4BEG[13] ,
    \Tile_X3Y4_SS4BEG[12] ,
    \Tile_X3Y4_SS4BEG[11] ,
    \Tile_X3Y4_SS4BEG[10] ,
    \Tile_X3Y4_SS4BEG[9] ,
    \Tile_X3Y4_SS4BEG[8] ,
    \Tile_X3Y4_SS4BEG[7] ,
    \Tile_X3Y4_SS4BEG[6] ,
    \Tile_X3Y4_SS4BEG[5] ,
    \Tile_X3Y4_SS4BEG[4] ,
    \Tile_X3Y4_SS4BEG[3] ,
    \Tile_X3Y4_SS4BEG[2] ,
    \Tile_X3Y4_SS4BEG[1] ,
    \Tile_X3Y4_SS4BEG[0] }),
    .W1BEG({\Tile_X3Y5_W1BEG[3] ,
    \Tile_X3Y5_W1BEG[2] ,
    \Tile_X3Y5_W1BEG[1] ,
    \Tile_X3Y5_W1BEG[0] }),
    .W1END({\Tile_X4Y5_W1BEG[3] ,
    \Tile_X4Y5_W1BEG[2] ,
    \Tile_X4Y5_W1BEG[1] ,
    \Tile_X4Y5_W1BEG[0] }),
    .W2BEG({\Tile_X3Y5_W2BEG[7] ,
    \Tile_X3Y5_W2BEG[6] ,
    \Tile_X3Y5_W2BEG[5] ,
    \Tile_X3Y5_W2BEG[4] ,
    \Tile_X3Y5_W2BEG[3] ,
    \Tile_X3Y5_W2BEG[2] ,
    \Tile_X3Y5_W2BEG[1] ,
    \Tile_X3Y5_W2BEG[0] }),
    .W2BEGb({\Tile_X3Y5_W2BEGb[7] ,
    \Tile_X3Y5_W2BEGb[6] ,
    \Tile_X3Y5_W2BEGb[5] ,
    \Tile_X3Y5_W2BEGb[4] ,
    \Tile_X3Y5_W2BEGb[3] ,
    \Tile_X3Y5_W2BEGb[2] ,
    \Tile_X3Y5_W2BEGb[1] ,
    \Tile_X3Y5_W2BEGb[0] }),
    .W2END({\Tile_X4Y5_W2BEGb[7] ,
    \Tile_X4Y5_W2BEGb[6] ,
    \Tile_X4Y5_W2BEGb[5] ,
    \Tile_X4Y5_W2BEGb[4] ,
    \Tile_X4Y5_W2BEGb[3] ,
    \Tile_X4Y5_W2BEGb[2] ,
    \Tile_X4Y5_W2BEGb[1] ,
    \Tile_X4Y5_W2BEGb[0] }),
    .W2MID({\Tile_X4Y5_W2BEG[7] ,
    \Tile_X4Y5_W2BEG[6] ,
    \Tile_X4Y5_W2BEG[5] ,
    \Tile_X4Y5_W2BEG[4] ,
    \Tile_X4Y5_W2BEG[3] ,
    \Tile_X4Y5_W2BEG[2] ,
    \Tile_X4Y5_W2BEG[1] ,
    \Tile_X4Y5_W2BEG[0] }),
    .W6BEG({\Tile_X3Y5_W6BEG[11] ,
    \Tile_X3Y5_W6BEG[10] ,
    \Tile_X3Y5_W6BEG[9] ,
    \Tile_X3Y5_W6BEG[8] ,
    \Tile_X3Y5_W6BEG[7] ,
    \Tile_X3Y5_W6BEG[6] ,
    \Tile_X3Y5_W6BEG[5] ,
    \Tile_X3Y5_W6BEG[4] ,
    \Tile_X3Y5_W6BEG[3] ,
    \Tile_X3Y5_W6BEG[2] ,
    \Tile_X3Y5_W6BEG[1] ,
    \Tile_X3Y5_W6BEG[0] }),
    .W6END({\Tile_X4Y5_W6BEG[11] ,
    \Tile_X4Y5_W6BEG[10] ,
    \Tile_X4Y5_W6BEG[9] ,
    \Tile_X4Y5_W6BEG[8] ,
    \Tile_X4Y5_W6BEG[7] ,
    \Tile_X4Y5_W6BEG[6] ,
    \Tile_X4Y5_W6BEG[5] ,
    \Tile_X4Y5_W6BEG[4] ,
    \Tile_X4Y5_W6BEG[3] ,
    \Tile_X4Y5_W6BEG[2] ,
    \Tile_X4Y5_W6BEG[1] ,
    \Tile_X4Y5_W6BEG[0] }),
    .WW4BEG({\Tile_X3Y5_WW4BEG[15] ,
    \Tile_X3Y5_WW4BEG[14] ,
    \Tile_X3Y5_WW4BEG[13] ,
    \Tile_X3Y5_WW4BEG[12] ,
    \Tile_X3Y5_WW4BEG[11] ,
    \Tile_X3Y5_WW4BEG[10] ,
    \Tile_X3Y5_WW4BEG[9] ,
    \Tile_X3Y5_WW4BEG[8] ,
    \Tile_X3Y5_WW4BEG[7] ,
    \Tile_X3Y5_WW4BEG[6] ,
    \Tile_X3Y5_WW4BEG[5] ,
    \Tile_X3Y5_WW4BEG[4] ,
    \Tile_X3Y5_WW4BEG[3] ,
    \Tile_X3Y5_WW4BEG[2] ,
    \Tile_X3Y5_WW4BEG[1] ,
    \Tile_X3Y5_WW4BEG[0] }),
    .WW4END({\Tile_X4Y5_WW4BEG[15] ,
    \Tile_X4Y5_WW4BEG[14] ,
    \Tile_X4Y5_WW4BEG[13] ,
    \Tile_X4Y5_WW4BEG[12] ,
    \Tile_X4Y5_WW4BEG[11] ,
    \Tile_X4Y5_WW4BEG[10] ,
    \Tile_X4Y5_WW4BEG[9] ,
    \Tile_X4Y5_WW4BEG[8] ,
    \Tile_X4Y5_WW4BEG[7] ,
    \Tile_X4Y5_WW4BEG[6] ,
    \Tile_X4Y5_WW4BEG[5] ,
    \Tile_X4Y5_WW4BEG[4] ,
    \Tile_X4Y5_WW4BEG[3] ,
    \Tile_X4Y5_WW4BEG[2] ,
    \Tile_X4Y5_WW4BEG[1] ,
    \Tile_X4Y5_WW4BEG[0] }));
 LUT4AB Tile_X3Y6_LUT4AB (.Ci(Tile_X3Y7_Co),
    .Co(Tile_X3Y6_Co),
    .UserCLK(Tile_X3Y7_UserCLKo),
    .UserCLKo(Tile_X3Y6_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X3Y6_E1BEG[3] ,
    \Tile_X3Y6_E1BEG[2] ,
    \Tile_X3Y6_E1BEG[1] ,
    \Tile_X3Y6_E1BEG[0] }),
    .E1END({\Tile_X2Y6_E1BEG[3] ,
    \Tile_X2Y6_E1BEG[2] ,
    \Tile_X2Y6_E1BEG[1] ,
    \Tile_X2Y6_E1BEG[0] }),
    .E2BEG({\Tile_X3Y6_E2BEG[7] ,
    \Tile_X3Y6_E2BEG[6] ,
    \Tile_X3Y6_E2BEG[5] ,
    \Tile_X3Y6_E2BEG[4] ,
    \Tile_X3Y6_E2BEG[3] ,
    \Tile_X3Y6_E2BEG[2] ,
    \Tile_X3Y6_E2BEG[1] ,
    \Tile_X3Y6_E2BEG[0] }),
    .E2BEGb({\Tile_X3Y6_E2BEGb[7] ,
    \Tile_X3Y6_E2BEGb[6] ,
    \Tile_X3Y6_E2BEGb[5] ,
    \Tile_X3Y6_E2BEGb[4] ,
    \Tile_X3Y6_E2BEGb[3] ,
    \Tile_X3Y6_E2BEGb[2] ,
    \Tile_X3Y6_E2BEGb[1] ,
    \Tile_X3Y6_E2BEGb[0] }),
    .E2END({\Tile_X2Y6_E2BEGb[7] ,
    \Tile_X2Y6_E2BEGb[6] ,
    \Tile_X2Y6_E2BEGb[5] ,
    \Tile_X2Y6_E2BEGb[4] ,
    \Tile_X2Y6_E2BEGb[3] ,
    \Tile_X2Y6_E2BEGb[2] ,
    \Tile_X2Y6_E2BEGb[1] ,
    \Tile_X2Y6_E2BEGb[0] }),
    .E2MID({\Tile_X2Y6_E2BEG[7] ,
    \Tile_X2Y6_E2BEG[6] ,
    \Tile_X2Y6_E2BEG[5] ,
    \Tile_X2Y6_E2BEG[4] ,
    \Tile_X2Y6_E2BEG[3] ,
    \Tile_X2Y6_E2BEG[2] ,
    \Tile_X2Y6_E2BEG[1] ,
    \Tile_X2Y6_E2BEG[0] }),
    .E6BEG({\Tile_X3Y6_E6BEG[11] ,
    \Tile_X3Y6_E6BEG[10] ,
    \Tile_X3Y6_E6BEG[9] ,
    \Tile_X3Y6_E6BEG[8] ,
    \Tile_X3Y6_E6BEG[7] ,
    \Tile_X3Y6_E6BEG[6] ,
    \Tile_X3Y6_E6BEG[5] ,
    \Tile_X3Y6_E6BEG[4] ,
    \Tile_X3Y6_E6BEG[3] ,
    \Tile_X3Y6_E6BEG[2] ,
    \Tile_X3Y6_E6BEG[1] ,
    \Tile_X3Y6_E6BEG[0] }),
    .E6END({\Tile_X2Y6_E6BEG[11] ,
    \Tile_X2Y6_E6BEG[10] ,
    \Tile_X2Y6_E6BEG[9] ,
    \Tile_X2Y6_E6BEG[8] ,
    \Tile_X2Y6_E6BEG[7] ,
    \Tile_X2Y6_E6BEG[6] ,
    \Tile_X2Y6_E6BEG[5] ,
    \Tile_X2Y6_E6BEG[4] ,
    \Tile_X2Y6_E6BEG[3] ,
    \Tile_X2Y6_E6BEG[2] ,
    \Tile_X2Y6_E6BEG[1] ,
    \Tile_X2Y6_E6BEG[0] }),
    .EE4BEG({\Tile_X3Y6_EE4BEG[15] ,
    \Tile_X3Y6_EE4BEG[14] ,
    \Tile_X3Y6_EE4BEG[13] ,
    \Tile_X3Y6_EE4BEG[12] ,
    \Tile_X3Y6_EE4BEG[11] ,
    \Tile_X3Y6_EE4BEG[10] ,
    \Tile_X3Y6_EE4BEG[9] ,
    \Tile_X3Y6_EE4BEG[8] ,
    \Tile_X3Y6_EE4BEG[7] ,
    \Tile_X3Y6_EE4BEG[6] ,
    \Tile_X3Y6_EE4BEG[5] ,
    \Tile_X3Y6_EE4BEG[4] ,
    \Tile_X3Y6_EE4BEG[3] ,
    \Tile_X3Y6_EE4BEG[2] ,
    \Tile_X3Y6_EE4BEG[1] ,
    \Tile_X3Y6_EE4BEG[0] }),
    .EE4END({\Tile_X2Y6_EE4BEG[15] ,
    \Tile_X2Y6_EE4BEG[14] ,
    \Tile_X2Y6_EE4BEG[13] ,
    \Tile_X2Y6_EE4BEG[12] ,
    \Tile_X2Y6_EE4BEG[11] ,
    \Tile_X2Y6_EE4BEG[10] ,
    \Tile_X2Y6_EE4BEG[9] ,
    \Tile_X2Y6_EE4BEG[8] ,
    \Tile_X2Y6_EE4BEG[7] ,
    \Tile_X2Y6_EE4BEG[6] ,
    \Tile_X2Y6_EE4BEG[5] ,
    \Tile_X2Y6_EE4BEG[4] ,
    \Tile_X2Y6_EE4BEG[3] ,
    \Tile_X2Y6_EE4BEG[2] ,
    \Tile_X2Y6_EE4BEG[1] ,
    \Tile_X2Y6_EE4BEG[0] }),
    .FrameData({\Tile_X2Y6_FrameData_O[31] ,
    \Tile_X2Y6_FrameData_O[30] ,
    \Tile_X2Y6_FrameData_O[29] ,
    \Tile_X2Y6_FrameData_O[28] ,
    \Tile_X2Y6_FrameData_O[27] ,
    \Tile_X2Y6_FrameData_O[26] ,
    \Tile_X2Y6_FrameData_O[25] ,
    \Tile_X2Y6_FrameData_O[24] ,
    \Tile_X2Y6_FrameData_O[23] ,
    \Tile_X2Y6_FrameData_O[22] ,
    \Tile_X2Y6_FrameData_O[21] ,
    \Tile_X2Y6_FrameData_O[20] ,
    \Tile_X2Y6_FrameData_O[19] ,
    \Tile_X2Y6_FrameData_O[18] ,
    \Tile_X2Y6_FrameData_O[17] ,
    \Tile_X2Y6_FrameData_O[16] ,
    \Tile_X2Y6_FrameData_O[15] ,
    \Tile_X2Y6_FrameData_O[14] ,
    \Tile_X2Y6_FrameData_O[13] ,
    \Tile_X2Y6_FrameData_O[12] ,
    \Tile_X2Y6_FrameData_O[11] ,
    \Tile_X2Y6_FrameData_O[10] ,
    \Tile_X2Y6_FrameData_O[9] ,
    \Tile_X2Y6_FrameData_O[8] ,
    \Tile_X2Y6_FrameData_O[7] ,
    \Tile_X2Y6_FrameData_O[6] ,
    \Tile_X2Y6_FrameData_O[5] ,
    \Tile_X2Y6_FrameData_O[4] ,
    \Tile_X2Y6_FrameData_O[3] ,
    \Tile_X2Y6_FrameData_O[2] ,
    \Tile_X2Y6_FrameData_O[1] ,
    \Tile_X2Y6_FrameData_O[0] }),
    .FrameData_O({\Tile_X3Y6_FrameData_O[31] ,
    \Tile_X3Y6_FrameData_O[30] ,
    \Tile_X3Y6_FrameData_O[29] ,
    \Tile_X3Y6_FrameData_O[28] ,
    \Tile_X3Y6_FrameData_O[27] ,
    \Tile_X3Y6_FrameData_O[26] ,
    \Tile_X3Y6_FrameData_O[25] ,
    \Tile_X3Y6_FrameData_O[24] ,
    \Tile_X3Y6_FrameData_O[23] ,
    \Tile_X3Y6_FrameData_O[22] ,
    \Tile_X3Y6_FrameData_O[21] ,
    \Tile_X3Y6_FrameData_O[20] ,
    \Tile_X3Y6_FrameData_O[19] ,
    \Tile_X3Y6_FrameData_O[18] ,
    \Tile_X3Y6_FrameData_O[17] ,
    \Tile_X3Y6_FrameData_O[16] ,
    \Tile_X3Y6_FrameData_O[15] ,
    \Tile_X3Y6_FrameData_O[14] ,
    \Tile_X3Y6_FrameData_O[13] ,
    \Tile_X3Y6_FrameData_O[12] ,
    \Tile_X3Y6_FrameData_O[11] ,
    \Tile_X3Y6_FrameData_O[10] ,
    \Tile_X3Y6_FrameData_O[9] ,
    \Tile_X3Y6_FrameData_O[8] ,
    \Tile_X3Y6_FrameData_O[7] ,
    \Tile_X3Y6_FrameData_O[6] ,
    \Tile_X3Y6_FrameData_O[5] ,
    \Tile_X3Y6_FrameData_O[4] ,
    \Tile_X3Y6_FrameData_O[3] ,
    \Tile_X3Y6_FrameData_O[2] ,
    \Tile_X3Y6_FrameData_O[1] ,
    \Tile_X3Y6_FrameData_O[0] }),
    .FrameStrobe({\Tile_X3Y7_FrameStrobe_O[19] ,
    \Tile_X3Y7_FrameStrobe_O[18] ,
    \Tile_X3Y7_FrameStrobe_O[17] ,
    \Tile_X3Y7_FrameStrobe_O[16] ,
    \Tile_X3Y7_FrameStrobe_O[15] ,
    \Tile_X3Y7_FrameStrobe_O[14] ,
    \Tile_X3Y7_FrameStrobe_O[13] ,
    \Tile_X3Y7_FrameStrobe_O[12] ,
    \Tile_X3Y7_FrameStrobe_O[11] ,
    \Tile_X3Y7_FrameStrobe_O[10] ,
    \Tile_X3Y7_FrameStrobe_O[9] ,
    \Tile_X3Y7_FrameStrobe_O[8] ,
    \Tile_X3Y7_FrameStrobe_O[7] ,
    \Tile_X3Y7_FrameStrobe_O[6] ,
    \Tile_X3Y7_FrameStrobe_O[5] ,
    \Tile_X3Y7_FrameStrobe_O[4] ,
    \Tile_X3Y7_FrameStrobe_O[3] ,
    \Tile_X3Y7_FrameStrobe_O[2] ,
    \Tile_X3Y7_FrameStrobe_O[1] ,
    \Tile_X3Y7_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X3Y6_FrameStrobe_O[19] ,
    \Tile_X3Y6_FrameStrobe_O[18] ,
    \Tile_X3Y6_FrameStrobe_O[17] ,
    \Tile_X3Y6_FrameStrobe_O[16] ,
    \Tile_X3Y6_FrameStrobe_O[15] ,
    \Tile_X3Y6_FrameStrobe_O[14] ,
    \Tile_X3Y6_FrameStrobe_O[13] ,
    \Tile_X3Y6_FrameStrobe_O[12] ,
    \Tile_X3Y6_FrameStrobe_O[11] ,
    \Tile_X3Y6_FrameStrobe_O[10] ,
    \Tile_X3Y6_FrameStrobe_O[9] ,
    \Tile_X3Y6_FrameStrobe_O[8] ,
    \Tile_X3Y6_FrameStrobe_O[7] ,
    \Tile_X3Y6_FrameStrobe_O[6] ,
    \Tile_X3Y6_FrameStrobe_O[5] ,
    \Tile_X3Y6_FrameStrobe_O[4] ,
    \Tile_X3Y6_FrameStrobe_O[3] ,
    \Tile_X3Y6_FrameStrobe_O[2] ,
    \Tile_X3Y6_FrameStrobe_O[1] ,
    \Tile_X3Y6_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X3Y6_N1BEG[3] ,
    \Tile_X3Y6_N1BEG[2] ,
    \Tile_X3Y6_N1BEG[1] ,
    \Tile_X3Y6_N1BEG[0] }),
    .N1END({\Tile_X3Y7_N1BEG[3] ,
    \Tile_X3Y7_N1BEG[2] ,
    \Tile_X3Y7_N1BEG[1] ,
    \Tile_X3Y7_N1BEG[0] }),
    .N2BEG({\Tile_X3Y6_N2BEG[7] ,
    \Tile_X3Y6_N2BEG[6] ,
    \Tile_X3Y6_N2BEG[5] ,
    \Tile_X3Y6_N2BEG[4] ,
    \Tile_X3Y6_N2BEG[3] ,
    \Tile_X3Y6_N2BEG[2] ,
    \Tile_X3Y6_N2BEG[1] ,
    \Tile_X3Y6_N2BEG[0] }),
    .N2BEGb({\Tile_X3Y6_N2BEGb[7] ,
    \Tile_X3Y6_N2BEGb[6] ,
    \Tile_X3Y6_N2BEGb[5] ,
    \Tile_X3Y6_N2BEGb[4] ,
    \Tile_X3Y6_N2BEGb[3] ,
    \Tile_X3Y6_N2BEGb[2] ,
    \Tile_X3Y6_N2BEGb[1] ,
    \Tile_X3Y6_N2BEGb[0] }),
    .N2END({\Tile_X3Y7_N2BEGb[7] ,
    \Tile_X3Y7_N2BEGb[6] ,
    \Tile_X3Y7_N2BEGb[5] ,
    \Tile_X3Y7_N2BEGb[4] ,
    \Tile_X3Y7_N2BEGb[3] ,
    \Tile_X3Y7_N2BEGb[2] ,
    \Tile_X3Y7_N2BEGb[1] ,
    \Tile_X3Y7_N2BEGb[0] }),
    .N2MID({\Tile_X3Y7_N2BEG[7] ,
    \Tile_X3Y7_N2BEG[6] ,
    \Tile_X3Y7_N2BEG[5] ,
    \Tile_X3Y7_N2BEG[4] ,
    \Tile_X3Y7_N2BEG[3] ,
    \Tile_X3Y7_N2BEG[2] ,
    \Tile_X3Y7_N2BEG[1] ,
    \Tile_X3Y7_N2BEG[0] }),
    .N4BEG({\Tile_X3Y6_N4BEG[15] ,
    \Tile_X3Y6_N4BEG[14] ,
    \Tile_X3Y6_N4BEG[13] ,
    \Tile_X3Y6_N4BEG[12] ,
    \Tile_X3Y6_N4BEG[11] ,
    \Tile_X3Y6_N4BEG[10] ,
    \Tile_X3Y6_N4BEG[9] ,
    \Tile_X3Y6_N4BEG[8] ,
    \Tile_X3Y6_N4BEG[7] ,
    \Tile_X3Y6_N4BEG[6] ,
    \Tile_X3Y6_N4BEG[5] ,
    \Tile_X3Y6_N4BEG[4] ,
    \Tile_X3Y6_N4BEG[3] ,
    \Tile_X3Y6_N4BEG[2] ,
    \Tile_X3Y6_N4BEG[1] ,
    \Tile_X3Y6_N4BEG[0] }),
    .N4END({\Tile_X3Y7_N4BEG[15] ,
    \Tile_X3Y7_N4BEG[14] ,
    \Tile_X3Y7_N4BEG[13] ,
    \Tile_X3Y7_N4BEG[12] ,
    \Tile_X3Y7_N4BEG[11] ,
    \Tile_X3Y7_N4BEG[10] ,
    \Tile_X3Y7_N4BEG[9] ,
    \Tile_X3Y7_N4BEG[8] ,
    \Tile_X3Y7_N4BEG[7] ,
    \Tile_X3Y7_N4BEG[6] ,
    \Tile_X3Y7_N4BEG[5] ,
    \Tile_X3Y7_N4BEG[4] ,
    \Tile_X3Y7_N4BEG[3] ,
    \Tile_X3Y7_N4BEG[2] ,
    \Tile_X3Y7_N4BEG[1] ,
    \Tile_X3Y7_N4BEG[0] }),
    .NN4BEG({\Tile_X3Y6_NN4BEG[15] ,
    \Tile_X3Y6_NN4BEG[14] ,
    \Tile_X3Y6_NN4BEG[13] ,
    \Tile_X3Y6_NN4BEG[12] ,
    \Tile_X3Y6_NN4BEG[11] ,
    \Tile_X3Y6_NN4BEG[10] ,
    \Tile_X3Y6_NN4BEG[9] ,
    \Tile_X3Y6_NN4BEG[8] ,
    \Tile_X3Y6_NN4BEG[7] ,
    \Tile_X3Y6_NN4BEG[6] ,
    \Tile_X3Y6_NN4BEG[5] ,
    \Tile_X3Y6_NN4BEG[4] ,
    \Tile_X3Y6_NN4BEG[3] ,
    \Tile_X3Y6_NN4BEG[2] ,
    \Tile_X3Y6_NN4BEG[1] ,
    \Tile_X3Y6_NN4BEG[0] }),
    .NN4END({\Tile_X3Y7_NN4BEG[15] ,
    \Tile_X3Y7_NN4BEG[14] ,
    \Tile_X3Y7_NN4BEG[13] ,
    \Tile_X3Y7_NN4BEG[12] ,
    \Tile_X3Y7_NN4BEG[11] ,
    \Tile_X3Y7_NN4BEG[10] ,
    \Tile_X3Y7_NN4BEG[9] ,
    \Tile_X3Y7_NN4BEG[8] ,
    \Tile_X3Y7_NN4BEG[7] ,
    \Tile_X3Y7_NN4BEG[6] ,
    \Tile_X3Y7_NN4BEG[5] ,
    \Tile_X3Y7_NN4BEG[4] ,
    \Tile_X3Y7_NN4BEG[3] ,
    \Tile_X3Y7_NN4BEG[2] ,
    \Tile_X3Y7_NN4BEG[1] ,
    \Tile_X3Y7_NN4BEG[0] }),
    .S1BEG({\Tile_X3Y6_S1BEG[3] ,
    \Tile_X3Y6_S1BEG[2] ,
    \Tile_X3Y6_S1BEG[1] ,
    \Tile_X3Y6_S1BEG[0] }),
    .S1END({\Tile_X3Y5_S1BEG[3] ,
    \Tile_X3Y5_S1BEG[2] ,
    \Tile_X3Y5_S1BEG[1] ,
    \Tile_X3Y5_S1BEG[0] }),
    .S2BEG({\Tile_X3Y6_S2BEG[7] ,
    \Tile_X3Y6_S2BEG[6] ,
    \Tile_X3Y6_S2BEG[5] ,
    \Tile_X3Y6_S2BEG[4] ,
    \Tile_X3Y6_S2BEG[3] ,
    \Tile_X3Y6_S2BEG[2] ,
    \Tile_X3Y6_S2BEG[1] ,
    \Tile_X3Y6_S2BEG[0] }),
    .S2BEGb({\Tile_X3Y6_S2BEGb[7] ,
    \Tile_X3Y6_S2BEGb[6] ,
    \Tile_X3Y6_S2BEGb[5] ,
    \Tile_X3Y6_S2BEGb[4] ,
    \Tile_X3Y6_S2BEGb[3] ,
    \Tile_X3Y6_S2BEGb[2] ,
    \Tile_X3Y6_S2BEGb[1] ,
    \Tile_X3Y6_S2BEGb[0] }),
    .S2END({\Tile_X3Y5_S2BEGb[7] ,
    \Tile_X3Y5_S2BEGb[6] ,
    \Tile_X3Y5_S2BEGb[5] ,
    \Tile_X3Y5_S2BEGb[4] ,
    \Tile_X3Y5_S2BEGb[3] ,
    \Tile_X3Y5_S2BEGb[2] ,
    \Tile_X3Y5_S2BEGb[1] ,
    \Tile_X3Y5_S2BEGb[0] }),
    .S2MID({\Tile_X3Y5_S2BEG[7] ,
    \Tile_X3Y5_S2BEG[6] ,
    \Tile_X3Y5_S2BEG[5] ,
    \Tile_X3Y5_S2BEG[4] ,
    \Tile_X3Y5_S2BEG[3] ,
    \Tile_X3Y5_S2BEG[2] ,
    \Tile_X3Y5_S2BEG[1] ,
    \Tile_X3Y5_S2BEG[0] }),
    .S4BEG({\Tile_X3Y6_S4BEG[15] ,
    \Tile_X3Y6_S4BEG[14] ,
    \Tile_X3Y6_S4BEG[13] ,
    \Tile_X3Y6_S4BEG[12] ,
    \Tile_X3Y6_S4BEG[11] ,
    \Tile_X3Y6_S4BEG[10] ,
    \Tile_X3Y6_S4BEG[9] ,
    \Tile_X3Y6_S4BEG[8] ,
    \Tile_X3Y6_S4BEG[7] ,
    \Tile_X3Y6_S4BEG[6] ,
    \Tile_X3Y6_S4BEG[5] ,
    \Tile_X3Y6_S4BEG[4] ,
    \Tile_X3Y6_S4BEG[3] ,
    \Tile_X3Y6_S4BEG[2] ,
    \Tile_X3Y6_S4BEG[1] ,
    \Tile_X3Y6_S4BEG[0] }),
    .S4END({\Tile_X3Y5_S4BEG[15] ,
    \Tile_X3Y5_S4BEG[14] ,
    \Tile_X3Y5_S4BEG[13] ,
    \Tile_X3Y5_S4BEG[12] ,
    \Tile_X3Y5_S4BEG[11] ,
    \Tile_X3Y5_S4BEG[10] ,
    \Tile_X3Y5_S4BEG[9] ,
    \Tile_X3Y5_S4BEG[8] ,
    \Tile_X3Y5_S4BEG[7] ,
    \Tile_X3Y5_S4BEG[6] ,
    \Tile_X3Y5_S4BEG[5] ,
    \Tile_X3Y5_S4BEG[4] ,
    \Tile_X3Y5_S4BEG[3] ,
    \Tile_X3Y5_S4BEG[2] ,
    \Tile_X3Y5_S4BEG[1] ,
    \Tile_X3Y5_S4BEG[0] }),
    .SS4BEG({\Tile_X3Y6_SS4BEG[15] ,
    \Tile_X3Y6_SS4BEG[14] ,
    \Tile_X3Y6_SS4BEG[13] ,
    \Tile_X3Y6_SS4BEG[12] ,
    \Tile_X3Y6_SS4BEG[11] ,
    \Tile_X3Y6_SS4BEG[10] ,
    \Tile_X3Y6_SS4BEG[9] ,
    \Tile_X3Y6_SS4BEG[8] ,
    \Tile_X3Y6_SS4BEG[7] ,
    \Tile_X3Y6_SS4BEG[6] ,
    \Tile_X3Y6_SS4BEG[5] ,
    \Tile_X3Y6_SS4BEG[4] ,
    \Tile_X3Y6_SS4BEG[3] ,
    \Tile_X3Y6_SS4BEG[2] ,
    \Tile_X3Y6_SS4BEG[1] ,
    \Tile_X3Y6_SS4BEG[0] }),
    .SS4END({\Tile_X3Y5_SS4BEG[15] ,
    \Tile_X3Y5_SS4BEG[14] ,
    \Tile_X3Y5_SS4BEG[13] ,
    \Tile_X3Y5_SS4BEG[12] ,
    \Tile_X3Y5_SS4BEG[11] ,
    \Tile_X3Y5_SS4BEG[10] ,
    \Tile_X3Y5_SS4BEG[9] ,
    \Tile_X3Y5_SS4BEG[8] ,
    \Tile_X3Y5_SS4BEG[7] ,
    \Tile_X3Y5_SS4BEG[6] ,
    \Tile_X3Y5_SS4BEG[5] ,
    \Tile_X3Y5_SS4BEG[4] ,
    \Tile_X3Y5_SS4BEG[3] ,
    \Tile_X3Y5_SS4BEG[2] ,
    \Tile_X3Y5_SS4BEG[1] ,
    \Tile_X3Y5_SS4BEG[0] }),
    .W1BEG({\Tile_X3Y6_W1BEG[3] ,
    \Tile_X3Y6_W1BEG[2] ,
    \Tile_X3Y6_W1BEG[1] ,
    \Tile_X3Y6_W1BEG[0] }),
    .W1END({\Tile_X4Y6_W1BEG[3] ,
    \Tile_X4Y6_W1BEG[2] ,
    \Tile_X4Y6_W1BEG[1] ,
    \Tile_X4Y6_W1BEG[0] }),
    .W2BEG({\Tile_X3Y6_W2BEG[7] ,
    \Tile_X3Y6_W2BEG[6] ,
    \Tile_X3Y6_W2BEG[5] ,
    \Tile_X3Y6_W2BEG[4] ,
    \Tile_X3Y6_W2BEG[3] ,
    \Tile_X3Y6_W2BEG[2] ,
    \Tile_X3Y6_W2BEG[1] ,
    \Tile_X3Y6_W2BEG[0] }),
    .W2BEGb({\Tile_X3Y6_W2BEGb[7] ,
    \Tile_X3Y6_W2BEGb[6] ,
    \Tile_X3Y6_W2BEGb[5] ,
    \Tile_X3Y6_W2BEGb[4] ,
    \Tile_X3Y6_W2BEGb[3] ,
    \Tile_X3Y6_W2BEGb[2] ,
    \Tile_X3Y6_W2BEGb[1] ,
    \Tile_X3Y6_W2BEGb[0] }),
    .W2END({\Tile_X4Y6_W2BEGb[7] ,
    \Tile_X4Y6_W2BEGb[6] ,
    \Tile_X4Y6_W2BEGb[5] ,
    \Tile_X4Y6_W2BEGb[4] ,
    \Tile_X4Y6_W2BEGb[3] ,
    \Tile_X4Y6_W2BEGb[2] ,
    \Tile_X4Y6_W2BEGb[1] ,
    \Tile_X4Y6_W2BEGb[0] }),
    .W2MID({\Tile_X4Y6_W2BEG[7] ,
    \Tile_X4Y6_W2BEG[6] ,
    \Tile_X4Y6_W2BEG[5] ,
    \Tile_X4Y6_W2BEG[4] ,
    \Tile_X4Y6_W2BEG[3] ,
    \Tile_X4Y6_W2BEG[2] ,
    \Tile_X4Y6_W2BEG[1] ,
    \Tile_X4Y6_W2BEG[0] }),
    .W6BEG({\Tile_X3Y6_W6BEG[11] ,
    \Tile_X3Y6_W6BEG[10] ,
    \Tile_X3Y6_W6BEG[9] ,
    \Tile_X3Y6_W6BEG[8] ,
    \Tile_X3Y6_W6BEG[7] ,
    \Tile_X3Y6_W6BEG[6] ,
    \Tile_X3Y6_W6BEG[5] ,
    \Tile_X3Y6_W6BEG[4] ,
    \Tile_X3Y6_W6BEG[3] ,
    \Tile_X3Y6_W6BEG[2] ,
    \Tile_X3Y6_W6BEG[1] ,
    \Tile_X3Y6_W6BEG[0] }),
    .W6END({\Tile_X4Y6_W6BEG[11] ,
    \Tile_X4Y6_W6BEG[10] ,
    \Tile_X4Y6_W6BEG[9] ,
    \Tile_X4Y6_W6BEG[8] ,
    \Tile_X4Y6_W6BEG[7] ,
    \Tile_X4Y6_W6BEG[6] ,
    \Tile_X4Y6_W6BEG[5] ,
    \Tile_X4Y6_W6BEG[4] ,
    \Tile_X4Y6_W6BEG[3] ,
    \Tile_X4Y6_W6BEG[2] ,
    \Tile_X4Y6_W6BEG[1] ,
    \Tile_X4Y6_W6BEG[0] }),
    .WW4BEG({\Tile_X3Y6_WW4BEG[15] ,
    \Tile_X3Y6_WW4BEG[14] ,
    \Tile_X3Y6_WW4BEG[13] ,
    \Tile_X3Y6_WW4BEG[12] ,
    \Tile_X3Y6_WW4BEG[11] ,
    \Tile_X3Y6_WW4BEG[10] ,
    \Tile_X3Y6_WW4BEG[9] ,
    \Tile_X3Y6_WW4BEG[8] ,
    \Tile_X3Y6_WW4BEG[7] ,
    \Tile_X3Y6_WW4BEG[6] ,
    \Tile_X3Y6_WW4BEG[5] ,
    \Tile_X3Y6_WW4BEG[4] ,
    \Tile_X3Y6_WW4BEG[3] ,
    \Tile_X3Y6_WW4BEG[2] ,
    \Tile_X3Y6_WW4BEG[1] ,
    \Tile_X3Y6_WW4BEG[0] }),
    .WW4END({\Tile_X4Y6_WW4BEG[15] ,
    \Tile_X4Y6_WW4BEG[14] ,
    \Tile_X4Y6_WW4BEG[13] ,
    \Tile_X4Y6_WW4BEG[12] ,
    \Tile_X4Y6_WW4BEG[11] ,
    \Tile_X4Y6_WW4BEG[10] ,
    \Tile_X4Y6_WW4BEG[9] ,
    \Tile_X4Y6_WW4BEG[8] ,
    \Tile_X4Y6_WW4BEG[7] ,
    \Tile_X4Y6_WW4BEG[6] ,
    \Tile_X4Y6_WW4BEG[5] ,
    \Tile_X4Y6_WW4BEG[4] ,
    \Tile_X4Y6_WW4BEG[3] ,
    \Tile_X4Y6_WW4BEG[2] ,
    \Tile_X4Y6_WW4BEG[1] ,
    \Tile_X4Y6_WW4BEG[0] }));
 LUT4AB Tile_X3Y7_LUT4AB (.Ci(Tile_X3Y8_Co),
    .Co(Tile_X3Y7_Co),
    .UserCLK(Tile_X3Y8_UserCLKo),
    .UserCLKo(Tile_X3Y7_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X3Y7_E1BEG[3] ,
    \Tile_X3Y7_E1BEG[2] ,
    \Tile_X3Y7_E1BEG[1] ,
    \Tile_X3Y7_E1BEG[0] }),
    .E1END({\Tile_X2Y7_E1BEG[3] ,
    \Tile_X2Y7_E1BEG[2] ,
    \Tile_X2Y7_E1BEG[1] ,
    \Tile_X2Y7_E1BEG[0] }),
    .E2BEG({\Tile_X3Y7_E2BEG[7] ,
    \Tile_X3Y7_E2BEG[6] ,
    \Tile_X3Y7_E2BEG[5] ,
    \Tile_X3Y7_E2BEG[4] ,
    \Tile_X3Y7_E2BEG[3] ,
    \Tile_X3Y7_E2BEG[2] ,
    \Tile_X3Y7_E2BEG[1] ,
    \Tile_X3Y7_E2BEG[0] }),
    .E2BEGb({\Tile_X3Y7_E2BEGb[7] ,
    \Tile_X3Y7_E2BEGb[6] ,
    \Tile_X3Y7_E2BEGb[5] ,
    \Tile_X3Y7_E2BEGb[4] ,
    \Tile_X3Y7_E2BEGb[3] ,
    \Tile_X3Y7_E2BEGb[2] ,
    \Tile_X3Y7_E2BEGb[1] ,
    \Tile_X3Y7_E2BEGb[0] }),
    .E2END({\Tile_X2Y7_E2BEGb[7] ,
    \Tile_X2Y7_E2BEGb[6] ,
    \Tile_X2Y7_E2BEGb[5] ,
    \Tile_X2Y7_E2BEGb[4] ,
    \Tile_X2Y7_E2BEGb[3] ,
    \Tile_X2Y7_E2BEGb[2] ,
    \Tile_X2Y7_E2BEGb[1] ,
    \Tile_X2Y7_E2BEGb[0] }),
    .E2MID({\Tile_X2Y7_E2BEG[7] ,
    \Tile_X2Y7_E2BEG[6] ,
    \Tile_X2Y7_E2BEG[5] ,
    \Tile_X2Y7_E2BEG[4] ,
    \Tile_X2Y7_E2BEG[3] ,
    \Tile_X2Y7_E2BEG[2] ,
    \Tile_X2Y7_E2BEG[1] ,
    \Tile_X2Y7_E2BEG[0] }),
    .E6BEG({\Tile_X3Y7_E6BEG[11] ,
    \Tile_X3Y7_E6BEG[10] ,
    \Tile_X3Y7_E6BEG[9] ,
    \Tile_X3Y7_E6BEG[8] ,
    \Tile_X3Y7_E6BEG[7] ,
    \Tile_X3Y7_E6BEG[6] ,
    \Tile_X3Y7_E6BEG[5] ,
    \Tile_X3Y7_E6BEG[4] ,
    \Tile_X3Y7_E6BEG[3] ,
    \Tile_X3Y7_E6BEG[2] ,
    \Tile_X3Y7_E6BEG[1] ,
    \Tile_X3Y7_E6BEG[0] }),
    .E6END({\Tile_X2Y7_E6BEG[11] ,
    \Tile_X2Y7_E6BEG[10] ,
    \Tile_X2Y7_E6BEG[9] ,
    \Tile_X2Y7_E6BEG[8] ,
    \Tile_X2Y7_E6BEG[7] ,
    \Tile_X2Y7_E6BEG[6] ,
    \Tile_X2Y7_E6BEG[5] ,
    \Tile_X2Y7_E6BEG[4] ,
    \Tile_X2Y7_E6BEG[3] ,
    \Tile_X2Y7_E6BEG[2] ,
    \Tile_X2Y7_E6BEG[1] ,
    \Tile_X2Y7_E6BEG[0] }),
    .EE4BEG({\Tile_X3Y7_EE4BEG[15] ,
    \Tile_X3Y7_EE4BEG[14] ,
    \Tile_X3Y7_EE4BEG[13] ,
    \Tile_X3Y7_EE4BEG[12] ,
    \Tile_X3Y7_EE4BEG[11] ,
    \Tile_X3Y7_EE4BEG[10] ,
    \Tile_X3Y7_EE4BEG[9] ,
    \Tile_X3Y7_EE4BEG[8] ,
    \Tile_X3Y7_EE4BEG[7] ,
    \Tile_X3Y7_EE4BEG[6] ,
    \Tile_X3Y7_EE4BEG[5] ,
    \Tile_X3Y7_EE4BEG[4] ,
    \Tile_X3Y7_EE4BEG[3] ,
    \Tile_X3Y7_EE4BEG[2] ,
    \Tile_X3Y7_EE4BEG[1] ,
    \Tile_X3Y7_EE4BEG[0] }),
    .EE4END({\Tile_X2Y7_EE4BEG[15] ,
    \Tile_X2Y7_EE4BEG[14] ,
    \Tile_X2Y7_EE4BEG[13] ,
    \Tile_X2Y7_EE4BEG[12] ,
    \Tile_X2Y7_EE4BEG[11] ,
    \Tile_X2Y7_EE4BEG[10] ,
    \Tile_X2Y7_EE4BEG[9] ,
    \Tile_X2Y7_EE4BEG[8] ,
    \Tile_X2Y7_EE4BEG[7] ,
    \Tile_X2Y7_EE4BEG[6] ,
    \Tile_X2Y7_EE4BEG[5] ,
    \Tile_X2Y7_EE4BEG[4] ,
    \Tile_X2Y7_EE4BEG[3] ,
    \Tile_X2Y7_EE4BEG[2] ,
    \Tile_X2Y7_EE4BEG[1] ,
    \Tile_X2Y7_EE4BEG[0] }),
    .FrameData({\Tile_X2Y7_FrameData_O[31] ,
    \Tile_X2Y7_FrameData_O[30] ,
    \Tile_X2Y7_FrameData_O[29] ,
    \Tile_X2Y7_FrameData_O[28] ,
    \Tile_X2Y7_FrameData_O[27] ,
    \Tile_X2Y7_FrameData_O[26] ,
    \Tile_X2Y7_FrameData_O[25] ,
    \Tile_X2Y7_FrameData_O[24] ,
    \Tile_X2Y7_FrameData_O[23] ,
    \Tile_X2Y7_FrameData_O[22] ,
    \Tile_X2Y7_FrameData_O[21] ,
    \Tile_X2Y7_FrameData_O[20] ,
    \Tile_X2Y7_FrameData_O[19] ,
    \Tile_X2Y7_FrameData_O[18] ,
    \Tile_X2Y7_FrameData_O[17] ,
    \Tile_X2Y7_FrameData_O[16] ,
    \Tile_X2Y7_FrameData_O[15] ,
    \Tile_X2Y7_FrameData_O[14] ,
    \Tile_X2Y7_FrameData_O[13] ,
    \Tile_X2Y7_FrameData_O[12] ,
    \Tile_X2Y7_FrameData_O[11] ,
    \Tile_X2Y7_FrameData_O[10] ,
    \Tile_X2Y7_FrameData_O[9] ,
    \Tile_X2Y7_FrameData_O[8] ,
    \Tile_X2Y7_FrameData_O[7] ,
    \Tile_X2Y7_FrameData_O[6] ,
    \Tile_X2Y7_FrameData_O[5] ,
    \Tile_X2Y7_FrameData_O[4] ,
    \Tile_X2Y7_FrameData_O[3] ,
    \Tile_X2Y7_FrameData_O[2] ,
    \Tile_X2Y7_FrameData_O[1] ,
    \Tile_X2Y7_FrameData_O[0] }),
    .FrameData_O({\Tile_X3Y7_FrameData_O[31] ,
    \Tile_X3Y7_FrameData_O[30] ,
    \Tile_X3Y7_FrameData_O[29] ,
    \Tile_X3Y7_FrameData_O[28] ,
    \Tile_X3Y7_FrameData_O[27] ,
    \Tile_X3Y7_FrameData_O[26] ,
    \Tile_X3Y7_FrameData_O[25] ,
    \Tile_X3Y7_FrameData_O[24] ,
    \Tile_X3Y7_FrameData_O[23] ,
    \Tile_X3Y7_FrameData_O[22] ,
    \Tile_X3Y7_FrameData_O[21] ,
    \Tile_X3Y7_FrameData_O[20] ,
    \Tile_X3Y7_FrameData_O[19] ,
    \Tile_X3Y7_FrameData_O[18] ,
    \Tile_X3Y7_FrameData_O[17] ,
    \Tile_X3Y7_FrameData_O[16] ,
    \Tile_X3Y7_FrameData_O[15] ,
    \Tile_X3Y7_FrameData_O[14] ,
    \Tile_X3Y7_FrameData_O[13] ,
    \Tile_X3Y7_FrameData_O[12] ,
    \Tile_X3Y7_FrameData_O[11] ,
    \Tile_X3Y7_FrameData_O[10] ,
    \Tile_X3Y7_FrameData_O[9] ,
    \Tile_X3Y7_FrameData_O[8] ,
    \Tile_X3Y7_FrameData_O[7] ,
    \Tile_X3Y7_FrameData_O[6] ,
    \Tile_X3Y7_FrameData_O[5] ,
    \Tile_X3Y7_FrameData_O[4] ,
    \Tile_X3Y7_FrameData_O[3] ,
    \Tile_X3Y7_FrameData_O[2] ,
    \Tile_X3Y7_FrameData_O[1] ,
    \Tile_X3Y7_FrameData_O[0] }),
    .FrameStrobe({\Tile_X3Y8_FrameStrobe_O[19] ,
    \Tile_X3Y8_FrameStrobe_O[18] ,
    \Tile_X3Y8_FrameStrobe_O[17] ,
    \Tile_X3Y8_FrameStrobe_O[16] ,
    \Tile_X3Y8_FrameStrobe_O[15] ,
    \Tile_X3Y8_FrameStrobe_O[14] ,
    \Tile_X3Y8_FrameStrobe_O[13] ,
    \Tile_X3Y8_FrameStrobe_O[12] ,
    \Tile_X3Y8_FrameStrobe_O[11] ,
    \Tile_X3Y8_FrameStrobe_O[10] ,
    \Tile_X3Y8_FrameStrobe_O[9] ,
    \Tile_X3Y8_FrameStrobe_O[8] ,
    \Tile_X3Y8_FrameStrobe_O[7] ,
    \Tile_X3Y8_FrameStrobe_O[6] ,
    \Tile_X3Y8_FrameStrobe_O[5] ,
    \Tile_X3Y8_FrameStrobe_O[4] ,
    \Tile_X3Y8_FrameStrobe_O[3] ,
    \Tile_X3Y8_FrameStrobe_O[2] ,
    \Tile_X3Y8_FrameStrobe_O[1] ,
    \Tile_X3Y8_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X3Y7_FrameStrobe_O[19] ,
    \Tile_X3Y7_FrameStrobe_O[18] ,
    \Tile_X3Y7_FrameStrobe_O[17] ,
    \Tile_X3Y7_FrameStrobe_O[16] ,
    \Tile_X3Y7_FrameStrobe_O[15] ,
    \Tile_X3Y7_FrameStrobe_O[14] ,
    \Tile_X3Y7_FrameStrobe_O[13] ,
    \Tile_X3Y7_FrameStrobe_O[12] ,
    \Tile_X3Y7_FrameStrobe_O[11] ,
    \Tile_X3Y7_FrameStrobe_O[10] ,
    \Tile_X3Y7_FrameStrobe_O[9] ,
    \Tile_X3Y7_FrameStrobe_O[8] ,
    \Tile_X3Y7_FrameStrobe_O[7] ,
    \Tile_X3Y7_FrameStrobe_O[6] ,
    \Tile_X3Y7_FrameStrobe_O[5] ,
    \Tile_X3Y7_FrameStrobe_O[4] ,
    \Tile_X3Y7_FrameStrobe_O[3] ,
    \Tile_X3Y7_FrameStrobe_O[2] ,
    \Tile_X3Y7_FrameStrobe_O[1] ,
    \Tile_X3Y7_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X3Y7_N1BEG[3] ,
    \Tile_X3Y7_N1BEG[2] ,
    \Tile_X3Y7_N1BEG[1] ,
    \Tile_X3Y7_N1BEG[0] }),
    .N1END({\Tile_X3Y8_N1BEG[3] ,
    \Tile_X3Y8_N1BEG[2] ,
    \Tile_X3Y8_N1BEG[1] ,
    \Tile_X3Y8_N1BEG[0] }),
    .N2BEG({\Tile_X3Y7_N2BEG[7] ,
    \Tile_X3Y7_N2BEG[6] ,
    \Tile_X3Y7_N2BEG[5] ,
    \Tile_X3Y7_N2BEG[4] ,
    \Tile_X3Y7_N2BEG[3] ,
    \Tile_X3Y7_N2BEG[2] ,
    \Tile_X3Y7_N2BEG[1] ,
    \Tile_X3Y7_N2BEG[0] }),
    .N2BEGb({\Tile_X3Y7_N2BEGb[7] ,
    \Tile_X3Y7_N2BEGb[6] ,
    \Tile_X3Y7_N2BEGb[5] ,
    \Tile_X3Y7_N2BEGb[4] ,
    \Tile_X3Y7_N2BEGb[3] ,
    \Tile_X3Y7_N2BEGb[2] ,
    \Tile_X3Y7_N2BEGb[1] ,
    \Tile_X3Y7_N2BEGb[0] }),
    .N2END({\Tile_X3Y8_N2BEGb[7] ,
    \Tile_X3Y8_N2BEGb[6] ,
    \Tile_X3Y8_N2BEGb[5] ,
    \Tile_X3Y8_N2BEGb[4] ,
    \Tile_X3Y8_N2BEGb[3] ,
    \Tile_X3Y8_N2BEGb[2] ,
    \Tile_X3Y8_N2BEGb[1] ,
    \Tile_X3Y8_N2BEGb[0] }),
    .N2MID({\Tile_X3Y8_N2BEG[7] ,
    \Tile_X3Y8_N2BEG[6] ,
    \Tile_X3Y8_N2BEG[5] ,
    \Tile_X3Y8_N2BEG[4] ,
    \Tile_X3Y8_N2BEG[3] ,
    \Tile_X3Y8_N2BEG[2] ,
    \Tile_X3Y8_N2BEG[1] ,
    \Tile_X3Y8_N2BEG[0] }),
    .N4BEG({\Tile_X3Y7_N4BEG[15] ,
    \Tile_X3Y7_N4BEG[14] ,
    \Tile_X3Y7_N4BEG[13] ,
    \Tile_X3Y7_N4BEG[12] ,
    \Tile_X3Y7_N4BEG[11] ,
    \Tile_X3Y7_N4BEG[10] ,
    \Tile_X3Y7_N4BEG[9] ,
    \Tile_X3Y7_N4BEG[8] ,
    \Tile_X3Y7_N4BEG[7] ,
    \Tile_X3Y7_N4BEG[6] ,
    \Tile_X3Y7_N4BEG[5] ,
    \Tile_X3Y7_N4BEG[4] ,
    \Tile_X3Y7_N4BEG[3] ,
    \Tile_X3Y7_N4BEG[2] ,
    \Tile_X3Y7_N4BEG[1] ,
    \Tile_X3Y7_N4BEG[0] }),
    .N4END({\Tile_X3Y8_N4BEG[15] ,
    \Tile_X3Y8_N4BEG[14] ,
    \Tile_X3Y8_N4BEG[13] ,
    \Tile_X3Y8_N4BEG[12] ,
    \Tile_X3Y8_N4BEG[11] ,
    \Tile_X3Y8_N4BEG[10] ,
    \Tile_X3Y8_N4BEG[9] ,
    \Tile_X3Y8_N4BEG[8] ,
    \Tile_X3Y8_N4BEG[7] ,
    \Tile_X3Y8_N4BEG[6] ,
    \Tile_X3Y8_N4BEG[5] ,
    \Tile_X3Y8_N4BEG[4] ,
    \Tile_X3Y8_N4BEG[3] ,
    \Tile_X3Y8_N4BEG[2] ,
    \Tile_X3Y8_N4BEG[1] ,
    \Tile_X3Y8_N4BEG[0] }),
    .NN4BEG({\Tile_X3Y7_NN4BEG[15] ,
    \Tile_X3Y7_NN4BEG[14] ,
    \Tile_X3Y7_NN4BEG[13] ,
    \Tile_X3Y7_NN4BEG[12] ,
    \Tile_X3Y7_NN4BEG[11] ,
    \Tile_X3Y7_NN4BEG[10] ,
    \Tile_X3Y7_NN4BEG[9] ,
    \Tile_X3Y7_NN4BEG[8] ,
    \Tile_X3Y7_NN4BEG[7] ,
    \Tile_X3Y7_NN4BEG[6] ,
    \Tile_X3Y7_NN4BEG[5] ,
    \Tile_X3Y7_NN4BEG[4] ,
    \Tile_X3Y7_NN4BEG[3] ,
    \Tile_X3Y7_NN4BEG[2] ,
    \Tile_X3Y7_NN4BEG[1] ,
    \Tile_X3Y7_NN4BEG[0] }),
    .NN4END({\Tile_X3Y8_NN4BEG[15] ,
    \Tile_X3Y8_NN4BEG[14] ,
    \Tile_X3Y8_NN4BEG[13] ,
    \Tile_X3Y8_NN4BEG[12] ,
    \Tile_X3Y8_NN4BEG[11] ,
    \Tile_X3Y8_NN4BEG[10] ,
    \Tile_X3Y8_NN4BEG[9] ,
    \Tile_X3Y8_NN4BEG[8] ,
    \Tile_X3Y8_NN4BEG[7] ,
    \Tile_X3Y8_NN4BEG[6] ,
    \Tile_X3Y8_NN4BEG[5] ,
    \Tile_X3Y8_NN4BEG[4] ,
    \Tile_X3Y8_NN4BEG[3] ,
    \Tile_X3Y8_NN4BEG[2] ,
    \Tile_X3Y8_NN4BEG[1] ,
    \Tile_X3Y8_NN4BEG[0] }),
    .S1BEG({\Tile_X3Y7_S1BEG[3] ,
    \Tile_X3Y7_S1BEG[2] ,
    \Tile_X3Y7_S1BEG[1] ,
    \Tile_X3Y7_S1BEG[0] }),
    .S1END({\Tile_X3Y6_S1BEG[3] ,
    \Tile_X3Y6_S1BEG[2] ,
    \Tile_X3Y6_S1BEG[1] ,
    \Tile_X3Y6_S1BEG[0] }),
    .S2BEG({\Tile_X3Y7_S2BEG[7] ,
    \Tile_X3Y7_S2BEG[6] ,
    \Tile_X3Y7_S2BEG[5] ,
    \Tile_X3Y7_S2BEG[4] ,
    \Tile_X3Y7_S2BEG[3] ,
    \Tile_X3Y7_S2BEG[2] ,
    \Tile_X3Y7_S2BEG[1] ,
    \Tile_X3Y7_S2BEG[0] }),
    .S2BEGb({\Tile_X3Y7_S2BEGb[7] ,
    \Tile_X3Y7_S2BEGb[6] ,
    \Tile_X3Y7_S2BEGb[5] ,
    \Tile_X3Y7_S2BEGb[4] ,
    \Tile_X3Y7_S2BEGb[3] ,
    \Tile_X3Y7_S2BEGb[2] ,
    \Tile_X3Y7_S2BEGb[1] ,
    \Tile_X3Y7_S2BEGb[0] }),
    .S2END({\Tile_X3Y6_S2BEGb[7] ,
    \Tile_X3Y6_S2BEGb[6] ,
    \Tile_X3Y6_S2BEGb[5] ,
    \Tile_X3Y6_S2BEGb[4] ,
    \Tile_X3Y6_S2BEGb[3] ,
    \Tile_X3Y6_S2BEGb[2] ,
    \Tile_X3Y6_S2BEGb[1] ,
    \Tile_X3Y6_S2BEGb[0] }),
    .S2MID({\Tile_X3Y6_S2BEG[7] ,
    \Tile_X3Y6_S2BEG[6] ,
    \Tile_X3Y6_S2BEG[5] ,
    \Tile_X3Y6_S2BEG[4] ,
    \Tile_X3Y6_S2BEG[3] ,
    \Tile_X3Y6_S2BEG[2] ,
    \Tile_X3Y6_S2BEG[1] ,
    \Tile_X3Y6_S2BEG[0] }),
    .S4BEG({\Tile_X3Y7_S4BEG[15] ,
    \Tile_X3Y7_S4BEG[14] ,
    \Tile_X3Y7_S4BEG[13] ,
    \Tile_X3Y7_S4BEG[12] ,
    \Tile_X3Y7_S4BEG[11] ,
    \Tile_X3Y7_S4BEG[10] ,
    \Tile_X3Y7_S4BEG[9] ,
    \Tile_X3Y7_S4BEG[8] ,
    \Tile_X3Y7_S4BEG[7] ,
    \Tile_X3Y7_S4BEG[6] ,
    \Tile_X3Y7_S4BEG[5] ,
    \Tile_X3Y7_S4BEG[4] ,
    \Tile_X3Y7_S4BEG[3] ,
    \Tile_X3Y7_S4BEG[2] ,
    \Tile_X3Y7_S4BEG[1] ,
    \Tile_X3Y7_S4BEG[0] }),
    .S4END({\Tile_X3Y6_S4BEG[15] ,
    \Tile_X3Y6_S4BEG[14] ,
    \Tile_X3Y6_S4BEG[13] ,
    \Tile_X3Y6_S4BEG[12] ,
    \Tile_X3Y6_S4BEG[11] ,
    \Tile_X3Y6_S4BEG[10] ,
    \Tile_X3Y6_S4BEG[9] ,
    \Tile_X3Y6_S4BEG[8] ,
    \Tile_X3Y6_S4BEG[7] ,
    \Tile_X3Y6_S4BEG[6] ,
    \Tile_X3Y6_S4BEG[5] ,
    \Tile_X3Y6_S4BEG[4] ,
    \Tile_X3Y6_S4BEG[3] ,
    \Tile_X3Y6_S4BEG[2] ,
    \Tile_X3Y6_S4BEG[1] ,
    \Tile_X3Y6_S4BEG[0] }),
    .SS4BEG({\Tile_X3Y7_SS4BEG[15] ,
    \Tile_X3Y7_SS4BEG[14] ,
    \Tile_X3Y7_SS4BEG[13] ,
    \Tile_X3Y7_SS4BEG[12] ,
    \Tile_X3Y7_SS4BEG[11] ,
    \Tile_X3Y7_SS4BEG[10] ,
    \Tile_X3Y7_SS4BEG[9] ,
    \Tile_X3Y7_SS4BEG[8] ,
    \Tile_X3Y7_SS4BEG[7] ,
    \Tile_X3Y7_SS4BEG[6] ,
    \Tile_X3Y7_SS4BEG[5] ,
    \Tile_X3Y7_SS4BEG[4] ,
    \Tile_X3Y7_SS4BEG[3] ,
    \Tile_X3Y7_SS4BEG[2] ,
    \Tile_X3Y7_SS4BEG[1] ,
    \Tile_X3Y7_SS4BEG[0] }),
    .SS4END({\Tile_X3Y6_SS4BEG[15] ,
    \Tile_X3Y6_SS4BEG[14] ,
    \Tile_X3Y6_SS4BEG[13] ,
    \Tile_X3Y6_SS4BEG[12] ,
    \Tile_X3Y6_SS4BEG[11] ,
    \Tile_X3Y6_SS4BEG[10] ,
    \Tile_X3Y6_SS4BEG[9] ,
    \Tile_X3Y6_SS4BEG[8] ,
    \Tile_X3Y6_SS4BEG[7] ,
    \Tile_X3Y6_SS4BEG[6] ,
    \Tile_X3Y6_SS4BEG[5] ,
    \Tile_X3Y6_SS4BEG[4] ,
    \Tile_X3Y6_SS4BEG[3] ,
    \Tile_X3Y6_SS4BEG[2] ,
    \Tile_X3Y6_SS4BEG[1] ,
    \Tile_X3Y6_SS4BEG[0] }),
    .W1BEG({\Tile_X3Y7_W1BEG[3] ,
    \Tile_X3Y7_W1BEG[2] ,
    \Tile_X3Y7_W1BEG[1] ,
    \Tile_X3Y7_W1BEG[0] }),
    .W1END({\Tile_X4Y7_W1BEG[3] ,
    \Tile_X4Y7_W1BEG[2] ,
    \Tile_X4Y7_W1BEG[1] ,
    \Tile_X4Y7_W1BEG[0] }),
    .W2BEG({\Tile_X3Y7_W2BEG[7] ,
    \Tile_X3Y7_W2BEG[6] ,
    \Tile_X3Y7_W2BEG[5] ,
    \Tile_X3Y7_W2BEG[4] ,
    \Tile_X3Y7_W2BEG[3] ,
    \Tile_X3Y7_W2BEG[2] ,
    \Tile_X3Y7_W2BEG[1] ,
    \Tile_X3Y7_W2BEG[0] }),
    .W2BEGb({\Tile_X3Y7_W2BEGb[7] ,
    \Tile_X3Y7_W2BEGb[6] ,
    \Tile_X3Y7_W2BEGb[5] ,
    \Tile_X3Y7_W2BEGb[4] ,
    \Tile_X3Y7_W2BEGb[3] ,
    \Tile_X3Y7_W2BEGb[2] ,
    \Tile_X3Y7_W2BEGb[1] ,
    \Tile_X3Y7_W2BEGb[0] }),
    .W2END({\Tile_X4Y7_W2BEGb[7] ,
    \Tile_X4Y7_W2BEGb[6] ,
    \Tile_X4Y7_W2BEGb[5] ,
    \Tile_X4Y7_W2BEGb[4] ,
    \Tile_X4Y7_W2BEGb[3] ,
    \Tile_X4Y7_W2BEGb[2] ,
    \Tile_X4Y7_W2BEGb[1] ,
    \Tile_X4Y7_W2BEGb[0] }),
    .W2MID({\Tile_X4Y7_W2BEG[7] ,
    \Tile_X4Y7_W2BEG[6] ,
    \Tile_X4Y7_W2BEG[5] ,
    \Tile_X4Y7_W2BEG[4] ,
    \Tile_X4Y7_W2BEG[3] ,
    \Tile_X4Y7_W2BEG[2] ,
    \Tile_X4Y7_W2BEG[1] ,
    \Tile_X4Y7_W2BEG[0] }),
    .W6BEG({\Tile_X3Y7_W6BEG[11] ,
    \Tile_X3Y7_W6BEG[10] ,
    \Tile_X3Y7_W6BEG[9] ,
    \Tile_X3Y7_W6BEG[8] ,
    \Tile_X3Y7_W6BEG[7] ,
    \Tile_X3Y7_W6BEG[6] ,
    \Tile_X3Y7_W6BEG[5] ,
    \Tile_X3Y7_W6BEG[4] ,
    \Tile_X3Y7_W6BEG[3] ,
    \Tile_X3Y7_W6BEG[2] ,
    \Tile_X3Y7_W6BEG[1] ,
    \Tile_X3Y7_W6BEG[0] }),
    .W6END({\Tile_X4Y7_W6BEG[11] ,
    \Tile_X4Y7_W6BEG[10] ,
    \Tile_X4Y7_W6BEG[9] ,
    \Tile_X4Y7_W6BEG[8] ,
    \Tile_X4Y7_W6BEG[7] ,
    \Tile_X4Y7_W6BEG[6] ,
    \Tile_X4Y7_W6BEG[5] ,
    \Tile_X4Y7_W6BEG[4] ,
    \Tile_X4Y7_W6BEG[3] ,
    \Tile_X4Y7_W6BEG[2] ,
    \Tile_X4Y7_W6BEG[1] ,
    \Tile_X4Y7_W6BEG[0] }),
    .WW4BEG({\Tile_X3Y7_WW4BEG[15] ,
    \Tile_X3Y7_WW4BEG[14] ,
    \Tile_X3Y7_WW4BEG[13] ,
    \Tile_X3Y7_WW4BEG[12] ,
    \Tile_X3Y7_WW4BEG[11] ,
    \Tile_X3Y7_WW4BEG[10] ,
    \Tile_X3Y7_WW4BEG[9] ,
    \Tile_X3Y7_WW4BEG[8] ,
    \Tile_X3Y7_WW4BEG[7] ,
    \Tile_X3Y7_WW4BEG[6] ,
    \Tile_X3Y7_WW4BEG[5] ,
    \Tile_X3Y7_WW4BEG[4] ,
    \Tile_X3Y7_WW4BEG[3] ,
    \Tile_X3Y7_WW4BEG[2] ,
    \Tile_X3Y7_WW4BEG[1] ,
    \Tile_X3Y7_WW4BEG[0] }),
    .WW4END({\Tile_X4Y7_WW4BEG[15] ,
    \Tile_X4Y7_WW4BEG[14] ,
    \Tile_X4Y7_WW4BEG[13] ,
    \Tile_X4Y7_WW4BEG[12] ,
    \Tile_X4Y7_WW4BEG[11] ,
    \Tile_X4Y7_WW4BEG[10] ,
    \Tile_X4Y7_WW4BEG[9] ,
    \Tile_X4Y7_WW4BEG[8] ,
    \Tile_X4Y7_WW4BEG[7] ,
    \Tile_X4Y7_WW4BEG[6] ,
    \Tile_X4Y7_WW4BEG[5] ,
    \Tile_X4Y7_WW4BEG[4] ,
    \Tile_X4Y7_WW4BEG[3] ,
    \Tile_X4Y7_WW4BEG[2] ,
    \Tile_X4Y7_WW4BEG[1] ,
    \Tile_X4Y7_WW4BEG[0] }));
 LUT4AB Tile_X3Y8_LUT4AB (.Ci(Tile_X3Y9_Co),
    .Co(Tile_X3Y8_Co),
    .UserCLK(Tile_X3Y9_UserCLKo),
    .UserCLKo(Tile_X3Y8_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X3Y8_E1BEG[3] ,
    \Tile_X3Y8_E1BEG[2] ,
    \Tile_X3Y8_E1BEG[1] ,
    \Tile_X3Y8_E1BEG[0] }),
    .E1END({\Tile_X2Y8_E1BEG[3] ,
    \Tile_X2Y8_E1BEG[2] ,
    \Tile_X2Y8_E1BEG[1] ,
    \Tile_X2Y8_E1BEG[0] }),
    .E2BEG({\Tile_X3Y8_E2BEG[7] ,
    \Tile_X3Y8_E2BEG[6] ,
    \Tile_X3Y8_E2BEG[5] ,
    \Tile_X3Y8_E2BEG[4] ,
    \Tile_X3Y8_E2BEG[3] ,
    \Tile_X3Y8_E2BEG[2] ,
    \Tile_X3Y8_E2BEG[1] ,
    \Tile_X3Y8_E2BEG[0] }),
    .E2BEGb({\Tile_X3Y8_E2BEGb[7] ,
    \Tile_X3Y8_E2BEGb[6] ,
    \Tile_X3Y8_E2BEGb[5] ,
    \Tile_X3Y8_E2BEGb[4] ,
    \Tile_X3Y8_E2BEGb[3] ,
    \Tile_X3Y8_E2BEGb[2] ,
    \Tile_X3Y8_E2BEGb[1] ,
    \Tile_X3Y8_E2BEGb[0] }),
    .E2END({\Tile_X2Y8_E2BEGb[7] ,
    \Tile_X2Y8_E2BEGb[6] ,
    \Tile_X2Y8_E2BEGb[5] ,
    \Tile_X2Y8_E2BEGb[4] ,
    \Tile_X2Y8_E2BEGb[3] ,
    \Tile_X2Y8_E2BEGb[2] ,
    \Tile_X2Y8_E2BEGb[1] ,
    \Tile_X2Y8_E2BEGb[0] }),
    .E2MID({\Tile_X2Y8_E2BEG[7] ,
    \Tile_X2Y8_E2BEG[6] ,
    \Tile_X2Y8_E2BEG[5] ,
    \Tile_X2Y8_E2BEG[4] ,
    \Tile_X2Y8_E2BEG[3] ,
    \Tile_X2Y8_E2BEG[2] ,
    \Tile_X2Y8_E2BEG[1] ,
    \Tile_X2Y8_E2BEG[0] }),
    .E6BEG({\Tile_X3Y8_E6BEG[11] ,
    \Tile_X3Y8_E6BEG[10] ,
    \Tile_X3Y8_E6BEG[9] ,
    \Tile_X3Y8_E6BEG[8] ,
    \Tile_X3Y8_E6BEG[7] ,
    \Tile_X3Y8_E6BEG[6] ,
    \Tile_X3Y8_E6BEG[5] ,
    \Tile_X3Y8_E6BEG[4] ,
    \Tile_X3Y8_E6BEG[3] ,
    \Tile_X3Y8_E6BEG[2] ,
    \Tile_X3Y8_E6BEG[1] ,
    \Tile_X3Y8_E6BEG[0] }),
    .E6END({\Tile_X2Y8_E6BEG[11] ,
    \Tile_X2Y8_E6BEG[10] ,
    \Tile_X2Y8_E6BEG[9] ,
    \Tile_X2Y8_E6BEG[8] ,
    \Tile_X2Y8_E6BEG[7] ,
    \Tile_X2Y8_E6BEG[6] ,
    \Tile_X2Y8_E6BEG[5] ,
    \Tile_X2Y8_E6BEG[4] ,
    \Tile_X2Y8_E6BEG[3] ,
    \Tile_X2Y8_E6BEG[2] ,
    \Tile_X2Y8_E6BEG[1] ,
    \Tile_X2Y8_E6BEG[0] }),
    .EE4BEG({\Tile_X3Y8_EE4BEG[15] ,
    \Tile_X3Y8_EE4BEG[14] ,
    \Tile_X3Y8_EE4BEG[13] ,
    \Tile_X3Y8_EE4BEG[12] ,
    \Tile_X3Y8_EE4BEG[11] ,
    \Tile_X3Y8_EE4BEG[10] ,
    \Tile_X3Y8_EE4BEG[9] ,
    \Tile_X3Y8_EE4BEG[8] ,
    \Tile_X3Y8_EE4BEG[7] ,
    \Tile_X3Y8_EE4BEG[6] ,
    \Tile_X3Y8_EE4BEG[5] ,
    \Tile_X3Y8_EE4BEG[4] ,
    \Tile_X3Y8_EE4BEG[3] ,
    \Tile_X3Y8_EE4BEG[2] ,
    \Tile_X3Y8_EE4BEG[1] ,
    \Tile_X3Y8_EE4BEG[0] }),
    .EE4END({\Tile_X2Y8_EE4BEG[15] ,
    \Tile_X2Y8_EE4BEG[14] ,
    \Tile_X2Y8_EE4BEG[13] ,
    \Tile_X2Y8_EE4BEG[12] ,
    \Tile_X2Y8_EE4BEG[11] ,
    \Tile_X2Y8_EE4BEG[10] ,
    \Tile_X2Y8_EE4BEG[9] ,
    \Tile_X2Y8_EE4BEG[8] ,
    \Tile_X2Y8_EE4BEG[7] ,
    \Tile_X2Y8_EE4BEG[6] ,
    \Tile_X2Y8_EE4BEG[5] ,
    \Tile_X2Y8_EE4BEG[4] ,
    \Tile_X2Y8_EE4BEG[3] ,
    \Tile_X2Y8_EE4BEG[2] ,
    \Tile_X2Y8_EE4BEG[1] ,
    \Tile_X2Y8_EE4BEG[0] }),
    .FrameData({\Tile_X2Y8_FrameData_O[31] ,
    \Tile_X2Y8_FrameData_O[30] ,
    \Tile_X2Y8_FrameData_O[29] ,
    \Tile_X2Y8_FrameData_O[28] ,
    \Tile_X2Y8_FrameData_O[27] ,
    \Tile_X2Y8_FrameData_O[26] ,
    \Tile_X2Y8_FrameData_O[25] ,
    \Tile_X2Y8_FrameData_O[24] ,
    \Tile_X2Y8_FrameData_O[23] ,
    \Tile_X2Y8_FrameData_O[22] ,
    \Tile_X2Y8_FrameData_O[21] ,
    \Tile_X2Y8_FrameData_O[20] ,
    \Tile_X2Y8_FrameData_O[19] ,
    \Tile_X2Y8_FrameData_O[18] ,
    \Tile_X2Y8_FrameData_O[17] ,
    \Tile_X2Y8_FrameData_O[16] ,
    \Tile_X2Y8_FrameData_O[15] ,
    \Tile_X2Y8_FrameData_O[14] ,
    \Tile_X2Y8_FrameData_O[13] ,
    \Tile_X2Y8_FrameData_O[12] ,
    \Tile_X2Y8_FrameData_O[11] ,
    \Tile_X2Y8_FrameData_O[10] ,
    \Tile_X2Y8_FrameData_O[9] ,
    \Tile_X2Y8_FrameData_O[8] ,
    \Tile_X2Y8_FrameData_O[7] ,
    \Tile_X2Y8_FrameData_O[6] ,
    \Tile_X2Y8_FrameData_O[5] ,
    \Tile_X2Y8_FrameData_O[4] ,
    \Tile_X2Y8_FrameData_O[3] ,
    \Tile_X2Y8_FrameData_O[2] ,
    \Tile_X2Y8_FrameData_O[1] ,
    \Tile_X2Y8_FrameData_O[0] }),
    .FrameData_O({\Tile_X3Y8_FrameData_O[31] ,
    \Tile_X3Y8_FrameData_O[30] ,
    \Tile_X3Y8_FrameData_O[29] ,
    \Tile_X3Y8_FrameData_O[28] ,
    \Tile_X3Y8_FrameData_O[27] ,
    \Tile_X3Y8_FrameData_O[26] ,
    \Tile_X3Y8_FrameData_O[25] ,
    \Tile_X3Y8_FrameData_O[24] ,
    \Tile_X3Y8_FrameData_O[23] ,
    \Tile_X3Y8_FrameData_O[22] ,
    \Tile_X3Y8_FrameData_O[21] ,
    \Tile_X3Y8_FrameData_O[20] ,
    \Tile_X3Y8_FrameData_O[19] ,
    \Tile_X3Y8_FrameData_O[18] ,
    \Tile_X3Y8_FrameData_O[17] ,
    \Tile_X3Y8_FrameData_O[16] ,
    \Tile_X3Y8_FrameData_O[15] ,
    \Tile_X3Y8_FrameData_O[14] ,
    \Tile_X3Y8_FrameData_O[13] ,
    \Tile_X3Y8_FrameData_O[12] ,
    \Tile_X3Y8_FrameData_O[11] ,
    \Tile_X3Y8_FrameData_O[10] ,
    \Tile_X3Y8_FrameData_O[9] ,
    \Tile_X3Y8_FrameData_O[8] ,
    \Tile_X3Y8_FrameData_O[7] ,
    \Tile_X3Y8_FrameData_O[6] ,
    \Tile_X3Y8_FrameData_O[5] ,
    \Tile_X3Y8_FrameData_O[4] ,
    \Tile_X3Y8_FrameData_O[3] ,
    \Tile_X3Y8_FrameData_O[2] ,
    \Tile_X3Y8_FrameData_O[1] ,
    \Tile_X3Y8_FrameData_O[0] }),
    .FrameStrobe({\Tile_X3Y9_FrameStrobe_O[19] ,
    \Tile_X3Y9_FrameStrobe_O[18] ,
    \Tile_X3Y9_FrameStrobe_O[17] ,
    \Tile_X3Y9_FrameStrobe_O[16] ,
    \Tile_X3Y9_FrameStrobe_O[15] ,
    \Tile_X3Y9_FrameStrobe_O[14] ,
    \Tile_X3Y9_FrameStrobe_O[13] ,
    \Tile_X3Y9_FrameStrobe_O[12] ,
    \Tile_X3Y9_FrameStrobe_O[11] ,
    \Tile_X3Y9_FrameStrobe_O[10] ,
    \Tile_X3Y9_FrameStrobe_O[9] ,
    \Tile_X3Y9_FrameStrobe_O[8] ,
    \Tile_X3Y9_FrameStrobe_O[7] ,
    \Tile_X3Y9_FrameStrobe_O[6] ,
    \Tile_X3Y9_FrameStrobe_O[5] ,
    \Tile_X3Y9_FrameStrobe_O[4] ,
    \Tile_X3Y9_FrameStrobe_O[3] ,
    \Tile_X3Y9_FrameStrobe_O[2] ,
    \Tile_X3Y9_FrameStrobe_O[1] ,
    \Tile_X3Y9_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X3Y8_FrameStrobe_O[19] ,
    \Tile_X3Y8_FrameStrobe_O[18] ,
    \Tile_X3Y8_FrameStrobe_O[17] ,
    \Tile_X3Y8_FrameStrobe_O[16] ,
    \Tile_X3Y8_FrameStrobe_O[15] ,
    \Tile_X3Y8_FrameStrobe_O[14] ,
    \Tile_X3Y8_FrameStrobe_O[13] ,
    \Tile_X3Y8_FrameStrobe_O[12] ,
    \Tile_X3Y8_FrameStrobe_O[11] ,
    \Tile_X3Y8_FrameStrobe_O[10] ,
    \Tile_X3Y8_FrameStrobe_O[9] ,
    \Tile_X3Y8_FrameStrobe_O[8] ,
    \Tile_X3Y8_FrameStrobe_O[7] ,
    \Tile_X3Y8_FrameStrobe_O[6] ,
    \Tile_X3Y8_FrameStrobe_O[5] ,
    \Tile_X3Y8_FrameStrobe_O[4] ,
    \Tile_X3Y8_FrameStrobe_O[3] ,
    \Tile_X3Y8_FrameStrobe_O[2] ,
    \Tile_X3Y8_FrameStrobe_O[1] ,
    \Tile_X3Y8_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X3Y8_N1BEG[3] ,
    \Tile_X3Y8_N1BEG[2] ,
    \Tile_X3Y8_N1BEG[1] ,
    \Tile_X3Y8_N1BEG[0] }),
    .N1END({\Tile_X3Y9_N1BEG[3] ,
    \Tile_X3Y9_N1BEG[2] ,
    \Tile_X3Y9_N1BEG[1] ,
    \Tile_X3Y9_N1BEG[0] }),
    .N2BEG({\Tile_X3Y8_N2BEG[7] ,
    \Tile_X3Y8_N2BEG[6] ,
    \Tile_X3Y8_N2BEG[5] ,
    \Tile_X3Y8_N2BEG[4] ,
    \Tile_X3Y8_N2BEG[3] ,
    \Tile_X3Y8_N2BEG[2] ,
    \Tile_X3Y8_N2BEG[1] ,
    \Tile_X3Y8_N2BEG[0] }),
    .N2BEGb({\Tile_X3Y8_N2BEGb[7] ,
    \Tile_X3Y8_N2BEGb[6] ,
    \Tile_X3Y8_N2BEGb[5] ,
    \Tile_X3Y8_N2BEGb[4] ,
    \Tile_X3Y8_N2BEGb[3] ,
    \Tile_X3Y8_N2BEGb[2] ,
    \Tile_X3Y8_N2BEGb[1] ,
    \Tile_X3Y8_N2BEGb[0] }),
    .N2END({\Tile_X3Y9_N2BEGb[7] ,
    \Tile_X3Y9_N2BEGb[6] ,
    \Tile_X3Y9_N2BEGb[5] ,
    \Tile_X3Y9_N2BEGb[4] ,
    \Tile_X3Y9_N2BEGb[3] ,
    \Tile_X3Y9_N2BEGb[2] ,
    \Tile_X3Y9_N2BEGb[1] ,
    \Tile_X3Y9_N2BEGb[0] }),
    .N2MID({\Tile_X3Y9_N2BEG[7] ,
    \Tile_X3Y9_N2BEG[6] ,
    \Tile_X3Y9_N2BEG[5] ,
    \Tile_X3Y9_N2BEG[4] ,
    \Tile_X3Y9_N2BEG[3] ,
    \Tile_X3Y9_N2BEG[2] ,
    \Tile_X3Y9_N2BEG[1] ,
    \Tile_X3Y9_N2BEG[0] }),
    .N4BEG({\Tile_X3Y8_N4BEG[15] ,
    \Tile_X3Y8_N4BEG[14] ,
    \Tile_X3Y8_N4BEG[13] ,
    \Tile_X3Y8_N4BEG[12] ,
    \Tile_X3Y8_N4BEG[11] ,
    \Tile_X3Y8_N4BEG[10] ,
    \Tile_X3Y8_N4BEG[9] ,
    \Tile_X3Y8_N4BEG[8] ,
    \Tile_X3Y8_N4BEG[7] ,
    \Tile_X3Y8_N4BEG[6] ,
    \Tile_X3Y8_N4BEG[5] ,
    \Tile_X3Y8_N4BEG[4] ,
    \Tile_X3Y8_N4BEG[3] ,
    \Tile_X3Y8_N4BEG[2] ,
    \Tile_X3Y8_N4BEG[1] ,
    \Tile_X3Y8_N4BEG[0] }),
    .N4END({\Tile_X3Y9_N4BEG[15] ,
    \Tile_X3Y9_N4BEG[14] ,
    \Tile_X3Y9_N4BEG[13] ,
    \Tile_X3Y9_N4BEG[12] ,
    \Tile_X3Y9_N4BEG[11] ,
    \Tile_X3Y9_N4BEG[10] ,
    \Tile_X3Y9_N4BEG[9] ,
    \Tile_X3Y9_N4BEG[8] ,
    \Tile_X3Y9_N4BEG[7] ,
    \Tile_X3Y9_N4BEG[6] ,
    \Tile_X3Y9_N4BEG[5] ,
    \Tile_X3Y9_N4BEG[4] ,
    \Tile_X3Y9_N4BEG[3] ,
    \Tile_X3Y9_N4BEG[2] ,
    \Tile_X3Y9_N4BEG[1] ,
    \Tile_X3Y9_N4BEG[0] }),
    .NN4BEG({\Tile_X3Y8_NN4BEG[15] ,
    \Tile_X3Y8_NN4BEG[14] ,
    \Tile_X3Y8_NN4BEG[13] ,
    \Tile_X3Y8_NN4BEG[12] ,
    \Tile_X3Y8_NN4BEG[11] ,
    \Tile_X3Y8_NN4BEG[10] ,
    \Tile_X3Y8_NN4BEG[9] ,
    \Tile_X3Y8_NN4BEG[8] ,
    \Tile_X3Y8_NN4BEG[7] ,
    \Tile_X3Y8_NN4BEG[6] ,
    \Tile_X3Y8_NN4BEG[5] ,
    \Tile_X3Y8_NN4BEG[4] ,
    \Tile_X3Y8_NN4BEG[3] ,
    \Tile_X3Y8_NN4BEG[2] ,
    \Tile_X3Y8_NN4BEG[1] ,
    \Tile_X3Y8_NN4BEG[0] }),
    .NN4END({\Tile_X3Y9_NN4BEG[15] ,
    \Tile_X3Y9_NN4BEG[14] ,
    \Tile_X3Y9_NN4BEG[13] ,
    \Tile_X3Y9_NN4BEG[12] ,
    \Tile_X3Y9_NN4BEG[11] ,
    \Tile_X3Y9_NN4BEG[10] ,
    \Tile_X3Y9_NN4BEG[9] ,
    \Tile_X3Y9_NN4BEG[8] ,
    \Tile_X3Y9_NN4BEG[7] ,
    \Tile_X3Y9_NN4BEG[6] ,
    \Tile_X3Y9_NN4BEG[5] ,
    \Tile_X3Y9_NN4BEG[4] ,
    \Tile_X3Y9_NN4BEG[3] ,
    \Tile_X3Y9_NN4BEG[2] ,
    \Tile_X3Y9_NN4BEG[1] ,
    \Tile_X3Y9_NN4BEG[0] }),
    .S1BEG({\Tile_X3Y8_S1BEG[3] ,
    \Tile_X3Y8_S1BEG[2] ,
    \Tile_X3Y8_S1BEG[1] ,
    \Tile_X3Y8_S1BEG[0] }),
    .S1END({\Tile_X3Y7_S1BEG[3] ,
    \Tile_X3Y7_S1BEG[2] ,
    \Tile_X3Y7_S1BEG[1] ,
    \Tile_X3Y7_S1BEG[0] }),
    .S2BEG({\Tile_X3Y8_S2BEG[7] ,
    \Tile_X3Y8_S2BEG[6] ,
    \Tile_X3Y8_S2BEG[5] ,
    \Tile_X3Y8_S2BEG[4] ,
    \Tile_X3Y8_S2BEG[3] ,
    \Tile_X3Y8_S2BEG[2] ,
    \Tile_X3Y8_S2BEG[1] ,
    \Tile_X3Y8_S2BEG[0] }),
    .S2BEGb({\Tile_X3Y8_S2BEGb[7] ,
    \Tile_X3Y8_S2BEGb[6] ,
    \Tile_X3Y8_S2BEGb[5] ,
    \Tile_X3Y8_S2BEGb[4] ,
    \Tile_X3Y8_S2BEGb[3] ,
    \Tile_X3Y8_S2BEGb[2] ,
    \Tile_X3Y8_S2BEGb[1] ,
    \Tile_X3Y8_S2BEGb[0] }),
    .S2END({\Tile_X3Y7_S2BEGb[7] ,
    \Tile_X3Y7_S2BEGb[6] ,
    \Tile_X3Y7_S2BEGb[5] ,
    \Tile_X3Y7_S2BEGb[4] ,
    \Tile_X3Y7_S2BEGb[3] ,
    \Tile_X3Y7_S2BEGb[2] ,
    \Tile_X3Y7_S2BEGb[1] ,
    \Tile_X3Y7_S2BEGb[0] }),
    .S2MID({\Tile_X3Y7_S2BEG[7] ,
    \Tile_X3Y7_S2BEG[6] ,
    \Tile_X3Y7_S2BEG[5] ,
    \Tile_X3Y7_S2BEG[4] ,
    \Tile_X3Y7_S2BEG[3] ,
    \Tile_X3Y7_S2BEG[2] ,
    \Tile_X3Y7_S2BEG[1] ,
    \Tile_X3Y7_S2BEG[0] }),
    .S4BEG({\Tile_X3Y8_S4BEG[15] ,
    \Tile_X3Y8_S4BEG[14] ,
    \Tile_X3Y8_S4BEG[13] ,
    \Tile_X3Y8_S4BEG[12] ,
    \Tile_X3Y8_S4BEG[11] ,
    \Tile_X3Y8_S4BEG[10] ,
    \Tile_X3Y8_S4BEG[9] ,
    \Tile_X3Y8_S4BEG[8] ,
    \Tile_X3Y8_S4BEG[7] ,
    \Tile_X3Y8_S4BEG[6] ,
    \Tile_X3Y8_S4BEG[5] ,
    \Tile_X3Y8_S4BEG[4] ,
    \Tile_X3Y8_S4BEG[3] ,
    \Tile_X3Y8_S4BEG[2] ,
    \Tile_X3Y8_S4BEG[1] ,
    \Tile_X3Y8_S4BEG[0] }),
    .S4END({\Tile_X3Y7_S4BEG[15] ,
    \Tile_X3Y7_S4BEG[14] ,
    \Tile_X3Y7_S4BEG[13] ,
    \Tile_X3Y7_S4BEG[12] ,
    \Tile_X3Y7_S4BEG[11] ,
    \Tile_X3Y7_S4BEG[10] ,
    \Tile_X3Y7_S4BEG[9] ,
    \Tile_X3Y7_S4BEG[8] ,
    \Tile_X3Y7_S4BEG[7] ,
    \Tile_X3Y7_S4BEG[6] ,
    \Tile_X3Y7_S4BEG[5] ,
    \Tile_X3Y7_S4BEG[4] ,
    \Tile_X3Y7_S4BEG[3] ,
    \Tile_X3Y7_S4BEG[2] ,
    \Tile_X3Y7_S4BEG[1] ,
    \Tile_X3Y7_S4BEG[0] }),
    .SS4BEG({\Tile_X3Y8_SS4BEG[15] ,
    \Tile_X3Y8_SS4BEG[14] ,
    \Tile_X3Y8_SS4BEG[13] ,
    \Tile_X3Y8_SS4BEG[12] ,
    \Tile_X3Y8_SS4BEG[11] ,
    \Tile_X3Y8_SS4BEG[10] ,
    \Tile_X3Y8_SS4BEG[9] ,
    \Tile_X3Y8_SS4BEG[8] ,
    \Tile_X3Y8_SS4BEG[7] ,
    \Tile_X3Y8_SS4BEG[6] ,
    \Tile_X3Y8_SS4BEG[5] ,
    \Tile_X3Y8_SS4BEG[4] ,
    \Tile_X3Y8_SS4BEG[3] ,
    \Tile_X3Y8_SS4BEG[2] ,
    \Tile_X3Y8_SS4BEG[1] ,
    \Tile_X3Y8_SS4BEG[0] }),
    .SS4END({\Tile_X3Y7_SS4BEG[15] ,
    \Tile_X3Y7_SS4BEG[14] ,
    \Tile_X3Y7_SS4BEG[13] ,
    \Tile_X3Y7_SS4BEG[12] ,
    \Tile_X3Y7_SS4BEG[11] ,
    \Tile_X3Y7_SS4BEG[10] ,
    \Tile_X3Y7_SS4BEG[9] ,
    \Tile_X3Y7_SS4BEG[8] ,
    \Tile_X3Y7_SS4BEG[7] ,
    \Tile_X3Y7_SS4BEG[6] ,
    \Tile_X3Y7_SS4BEG[5] ,
    \Tile_X3Y7_SS4BEG[4] ,
    \Tile_X3Y7_SS4BEG[3] ,
    \Tile_X3Y7_SS4BEG[2] ,
    \Tile_X3Y7_SS4BEG[1] ,
    \Tile_X3Y7_SS4BEG[0] }),
    .W1BEG({\Tile_X3Y8_W1BEG[3] ,
    \Tile_X3Y8_W1BEG[2] ,
    \Tile_X3Y8_W1BEG[1] ,
    \Tile_X3Y8_W1BEG[0] }),
    .W1END({\Tile_X4Y8_W1BEG[3] ,
    \Tile_X4Y8_W1BEG[2] ,
    \Tile_X4Y8_W1BEG[1] ,
    \Tile_X4Y8_W1BEG[0] }),
    .W2BEG({\Tile_X3Y8_W2BEG[7] ,
    \Tile_X3Y8_W2BEG[6] ,
    \Tile_X3Y8_W2BEG[5] ,
    \Tile_X3Y8_W2BEG[4] ,
    \Tile_X3Y8_W2BEG[3] ,
    \Tile_X3Y8_W2BEG[2] ,
    \Tile_X3Y8_W2BEG[1] ,
    \Tile_X3Y8_W2BEG[0] }),
    .W2BEGb({\Tile_X3Y8_W2BEGb[7] ,
    \Tile_X3Y8_W2BEGb[6] ,
    \Tile_X3Y8_W2BEGb[5] ,
    \Tile_X3Y8_W2BEGb[4] ,
    \Tile_X3Y8_W2BEGb[3] ,
    \Tile_X3Y8_W2BEGb[2] ,
    \Tile_X3Y8_W2BEGb[1] ,
    \Tile_X3Y8_W2BEGb[0] }),
    .W2END({\Tile_X4Y8_W2BEGb[7] ,
    \Tile_X4Y8_W2BEGb[6] ,
    \Tile_X4Y8_W2BEGb[5] ,
    \Tile_X4Y8_W2BEGb[4] ,
    \Tile_X4Y8_W2BEGb[3] ,
    \Tile_X4Y8_W2BEGb[2] ,
    \Tile_X4Y8_W2BEGb[1] ,
    \Tile_X4Y8_W2BEGb[0] }),
    .W2MID({\Tile_X4Y8_W2BEG[7] ,
    \Tile_X4Y8_W2BEG[6] ,
    \Tile_X4Y8_W2BEG[5] ,
    \Tile_X4Y8_W2BEG[4] ,
    \Tile_X4Y8_W2BEG[3] ,
    \Tile_X4Y8_W2BEG[2] ,
    \Tile_X4Y8_W2BEG[1] ,
    \Tile_X4Y8_W2BEG[0] }),
    .W6BEG({\Tile_X3Y8_W6BEG[11] ,
    \Tile_X3Y8_W6BEG[10] ,
    \Tile_X3Y8_W6BEG[9] ,
    \Tile_X3Y8_W6BEG[8] ,
    \Tile_X3Y8_W6BEG[7] ,
    \Tile_X3Y8_W6BEG[6] ,
    \Tile_X3Y8_W6BEG[5] ,
    \Tile_X3Y8_W6BEG[4] ,
    \Tile_X3Y8_W6BEG[3] ,
    \Tile_X3Y8_W6BEG[2] ,
    \Tile_X3Y8_W6BEG[1] ,
    \Tile_X3Y8_W6BEG[0] }),
    .W6END({\Tile_X4Y8_W6BEG[11] ,
    \Tile_X4Y8_W6BEG[10] ,
    \Tile_X4Y8_W6BEG[9] ,
    \Tile_X4Y8_W6BEG[8] ,
    \Tile_X4Y8_W6BEG[7] ,
    \Tile_X4Y8_W6BEG[6] ,
    \Tile_X4Y8_W6BEG[5] ,
    \Tile_X4Y8_W6BEG[4] ,
    \Tile_X4Y8_W6BEG[3] ,
    \Tile_X4Y8_W6BEG[2] ,
    \Tile_X4Y8_W6BEG[1] ,
    \Tile_X4Y8_W6BEG[0] }),
    .WW4BEG({\Tile_X3Y8_WW4BEG[15] ,
    \Tile_X3Y8_WW4BEG[14] ,
    \Tile_X3Y8_WW4BEG[13] ,
    \Tile_X3Y8_WW4BEG[12] ,
    \Tile_X3Y8_WW4BEG[11] ,
    \Tile_X3Y8_WW4BEG[10] ,
    \Tile_X3Y8_WW4BEG[9] ,
    \Tile_X3Y8_WW4BEG[8] ,
    \Tile_X3Y8_WW4BEG[7] ,
    \Tile_X3Y8_WW4BEG[6] ,
    \Tile_X3Y8_WW4BEG[5] ,
    \Tile_X3Y8_WW4BEG[4] ,
    \Tile_X3Y8_WW4BEG[3] ,
    \Tile_X3Y8_WW4BEG[2] ,
    \Tile_X3Y8_WW4BEG[1] ,
    \Tile_X3Y8_WW4BEG[0] }),
    .WW4END({\Tile_X4Y8_WW4BEG[15] ,
    \Tile_X4Y8_WW4BEG[14] ,
    \Tile_X4Y8_WW4BEG[13] ,
    \Tile_X4Y8_WW4BEG[12] ,
    \Tile_X4Y8_WW4BEG[11] ,
    \Tile_X4Y8_WW4BEG[10] ,
    \Tile_X4Y8_WW4BEG[9] ,
    \Tile_X4Y8_WW4BEG[8] ,
    \Tile_X4Y8_WW4BEG[7] ,
    \Tile_X4Y8_WW4BEG[6] ,
    \Tile_X4Y8_WW4BEG[5] ,
    \Tile_X4Y8_WW4BEG[4] ,
    \Tile_X4Y8_WW4BEG[3] ,
    \Tile_X4Y8_WW4BEG[2] ,
    \Tile_X4Y8_WW4BEG[1] ,
    \Tile_X4Y8_WW4BEG[0] }));
 LUT4AB Tile_X3Y9_LUT4AB (.Ci(Tile_X3Y10_Co),
    .Co(Tile_X3Y9_Co),
    .UserCLK(Tile_X3Y10_UserCLKo),
    .UserCLKo(Tile_X3Y9_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X3Y9_E1BEG[3] ,
    \Tile_X3Y9_E1BEG[2] ,
    \Tile_X3Y9_E1BEG[1] ,
    \Tile_X3Y9_E1BEG[0] }),
    .E1END({\Tile_X2Y9_E1BEG[3] ,
    \Tile_X2Y9_E1BEG[2] ,
    \Tile_X2Y9_E1BEG[1] ,
    \Tile_X2Y9_E1BEG[0] }),
    .E2BEG({\Tile_X3Y9_E2BEG[7] ,
    \Tile_X3Y9_E2BEG[6] ,
    \Tile_X3Y9_E2BEG[5] ,
    \Tile_X3Y9_E2BEG[4] ,
    \Tile_X3Y9_E2BEG[3] ,
    \Tile_X3Y9_E2BEG[2] ,
    \Tile_X3Y9_E2BEG[1] ,
    \Tile_X3Y9_E2BEG[0] }),
    .E2BEGb({\Tile_X3Y9_E2BEGb[7] ,
    \Tile_X3Y9_E2BEGb[6] ,
    \Tile_X3Y9_E2BEGb[5] ,
    \Tile_X3Y9_E2BEGb[4] ,
    \Tile_X3Y9_E2BEGb[3] ,
    \Tile_X3Y9_E2BEGb[2] ,
    \Tile_X3Y9_E2BEGb[1] ,
    \Tile_X3Y9_E2BEGb[0] }),
    .E2END({\Tile_X2Y9_E2BEGb[7] ,
    \Tile_X2Y9_E2BEGb[6] ,
    \Tile_X2Y9_E2BEGb[5] ,
    \Tile_X2Y9_E2BEGb[4] ,
    \Tile_X2Y9_E2BEGb[3] ,
    \Tile_X2Y9_E2BEGb[2] ,
    \Tile_X2Y9_E2BEGb[1] ,
    \Tile_X2Y9_E2BEGb[0] }),
    .E2MID({\Tile_X2Y9_E2BEG[7] ,
    \Tile_X2Y9_E2BEG[6] ,
    \Tile_X2Y9_E2BEG[5] ,
    \Tile_X2Y9_E2BEG[4] ,
    \Tile_X2Y9_E2BEG[3] ,
    \Tile_X2Y9_E2BEG[2] ,
    \Tile_X2Y9_E2BEG[1] ,
    \Tile_X2Y9_E2BEG[0] }),
    .E6BEG({\Tile_X3Y9_E6BEG[11] ,
    \Tile_X3Y9_E6BEG[10] ,
    \Tile_X3Y9_E6BEG[9] ,
    \Tile_X3Y9_E6BEG[8] ,
    \Tile_X3Y9_E6BEG[7] ,
    \Tile_X3Y9_E6BEG[6] ,
    \Tile_X3Y9_E6BEG[5] ,
    \Tile_X3Y9_E6BEG[4] ,
    \Tile_X3Y9_E6BEG[3] ,
    \Tile_X3Y9_E6BEG[2] ,
    \Tile_X3Y9_E6BEG[1] ,
    \Tile_X3Y9_E6BEG[0] }),
    .E6END({\Tile_X2Y9_E6BEG[11] ,
    \Tile_X2Y9_E6BEG[10] ,
    \Tile_X2Y9_E6BEG[9] ,
    \Tile_X2Y9_E6BEG[8] ,
    \Tile_X2Y9_E6BEG[7] ,
    \Tile_X2Y9_E6BEG[6] ,
    \Tile_X2Y9_E6BEG[5] ,
    \Tile_X2Y9_E6BEG[4] ,
    \Tile_X2Y9_E6BEG[3] ,
    \Tile_X2Y9_E6BEG[2] ,
    \Tile_X2Y9_E6BEG[1] ,
    \Tile_X2Y9_E6BEG[0] }),
    .EE4BEG({\Tile_X3Y9_EE4BEG[15] ,
    \Tile_X3Y9_EE4BEG[14] ,
    \Tile_X3Y9_EE4BEG[13] ,
    \Tile_X3Y9_EE4BEG[12] ,
    \Tile_X3Y9_EE4BEG[11] ,
    \Tile_X3Y9_EE4BEG[10] ,
    \Tile_X3Y9_EE4BEG[9] ,
    \Tile_X3Y9_EE4BEG[8] ,
    \Tile_X3Y9_EE4BEG[7] ,
    \Tile_X3Y9_EE4BEG[6] ,
    \Tile_X3Y9_EE4BEG[5] ,
    \Tile_X3Y9_EE4BEG[4] ,
    \Tile_X3Y9_EE4BEG[3] ,
    \Tile_X3Y9_EE4BEG[2] ,
    \Tile_X3Y9_EE4BEG[1] ,
    \Tile_X3Y9_EE4BEG[0] }),
    .EE4END({\Tile_X2Y9_EE4BEG[15] ,
    \Tile_X2Y9_EE4BEG[14] ,
    \Tile_X2Y9_EE4BEG[13] ,
    \Tile_X2Y9_EE4BEG[12] ,
    \Tile_X2Y9_EE4BEG[11] ,
    \Tile_X2Y9_EE4BEG[10] ,
    \Tile_X2Y9_EE4BEG[9] ,
    \Tile_X2Y9_EE4BEG[8] ,
    \Tile_X2Y9_EE4BEG[7] ,
    \Tile_X2Y9_EE4BEG[6] ,
    \Tile_X2Y9_EE4BEG[5] ,
    \Tile_X2Y9_EE4BEG[4] ,
    \Tile_X2Y9_EE4BEG[3] ,
    \Tile_X2Y9_EE4BEG[2] ,
    \Tile_X2Y9_EE4BEG[1] ,
    \Tile_X2Y9_EE4BEG[0] }),
    .FrameData({\Tile_X2Y9_FrameData_O[31] ,
    \Tile_X2Y9_FrameData_O[30] ,
    \Tile_X2Y9_FrameData_O[29] ,
    \Tile_X2Y9_FrameData_O[28] ,
    \Tile_X2Y9_FrameData_O[27] ,
    \Tile_X2Y9_FrameData_O[26] ,
    \Tile_X2Y9_FrameData_O[25] ,
    \Tile_X2Y9_FrameData_O[24] ,
    \Tile_X2Y9_FrameData_O[23] ,
    \Tile_X2Y9_FrameData_O[22] ,
    \Tile_X2Y9_FrameData_O[21] ,
    \Tile_X2Y9_FrameData_O[20] ,
    \Tile_X2Y9_FrameData_O[19] ,
    \Tile_X2Y9_FrameData_O[18] ,
    \Tile_X2Y9_FrameData_O[17] ,
    \Tile_X2Y9_FrameData_O[16] ,
    \Tile_X2Y9_FrameData_O[15] ,
    \Tile_X2Y9_FrameData_O[14] ,
    \Tile_X2Y9_FrameData_O[13] ,
    \Tile_X2Y9_FrameData_O[12] ,
    \Tile_X2Y9_FrameData_O[11] ,
    \Tile_X2Y9_FrameData_O[10] ,
    \Tile_X2Y9_FrameData_O[9] ,
    \Tile_X2Y9_FrameData_O[8] ,
    \Tile_X2Y9_FrameData_O[7] ,
    \Tile_X2Y9_FrameData_O[6] ,
    \Tile_X2Y9_FrameData_O[5] ,
    \Tile_X2Y9_FrameData_O[4] ,
    \Tile_X2Y9_FrameData_O[3] ,
    \Tile_X2Y9_FrameData_O[2] ,
    \Tile_X2Y9_FrameData_O[1] ,
    \Tile_X2Y9_FrameData_O[0] }),
    .FrameData_O({\Tile_X3Y9_FrameData_O[31] ,
    \Tile_X3Y9_FrameData_O[30] ,
    \Tile_X3Y9_FrameData_O[29] ,
    \Tile_X3Y9_FrameData_O[28] ,
    \Tile_X3Y9_FrameData_O[27] ,
    \Tile_X3Y9_FrameData_O[26] ,
    \Tile_X3Y9_FrameData_O[25] ,
    \Tile_X3Y9_FrameData_O[24] ,
    \Tile_X3Y9_FrameData_O[23] ,
    \Tile_X3Y9_FrameData_O[22] ,
    \Tile_X3Y9_FrameData_O[21] ,
    \Tile_X3Y9_FrameData_O[20] ,
    \Tile_X3Y9_FrameData_O[19] ,
    \Tile_X3Y9_FrameData_O[18] ,
    \Tile_X3Y9_FrameData_O[17] ,
    \Tile_X3Y9_FrameData_O[16] ,
    \Tile_X3Y9_FrameData_O[15] ,
    \Tile_X3Y9_FrameData_O[14] ,
    \Tile_X3Y9_FrameData_O[13] ,
    \Tile_X3Y9_FrameData_O[12] ,
    \Tile_X3Y9_FrameData_O[11] ,
    \Tile_X3Y9_FrameData_O[10] ,
    \Tile_X3Y9_FrameData_O[9] ,
    \Tile_X3Y9_FrameData_O[8] ,
    \Tile_X3Y9_FrameData_O[7] ,
    \Tile_X3Y9_FrameData_O[6] ,
    \Tile_X3Y9_FrameData_O[5] ,
    \Tile_X3Y9_FrameData_O[4] ,
    \Tile_X3Y9_FrameData_O[3] ,
    \Tile_X3Y9_FrameData_O[2] ,
    \Tile_X3Y9_FrameData_O[1] ,
    \Tile_X3Y9_FrameData_O[0] }),
    .FrameStrobe({\Tile_X3Y10_FrameStrobe_O[19] ,
    \Tile_X3Y10_FrameStrobe_O[18] ,
    \Tile_X3Y10_FrameStrobe_O[17] ,
    \Tile_X3Y10_FrameStrobe_O[16] ,
    \Tile_X3Y10_FrameStrobe_O[15] ,
    \Tile_X3Y10_FrameStrobe_O[14] ,
    \Tile_X3Y10_FrameStrobe_O[13] ,
    \Tile_X3Y10_FrameStrobe_O[12] ,
    \Tile_X3Y10_FrameStrobe_O[11] ,
    \Tile_X3Y10_FrameStrobe_O[10] ,
    \Tile_X3Y10_FrameStrobe_O[9] ,
    \Tile_X3Y10_FrameStrobe_O[8] ,
    \Tile_X3Y10_FrameStrobe_O[7] ,
    \Tile_X3Y10_FrameStrobe_O[6] ,
    \Tile_X3Y10_FrameStrobe_O[5] ,
    \Tile_X3Y10_FrameStrobe_O[4] ,
    \Tile_X3Y10_FrameStrobe_O[3] ,
    \Tile_X3Y10_FrameStrobe_O[2] ,
    \Tile_X3Y10_FrameStrobe_O[1] ,
    \Tile_X3Y10_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X3Y9_FrameStrobe_O[19] ,
    \Tile_X3Y9_FrameStrobe_O[18] ,
    \Tile_X3Y9_FrameStrobe_O[17] ,
    \Tile_X3Y9_FrameStrobe_O[16] ,
    \Tile_X3Y9_FrameStrobe_O[15] ,
    \Tile_X3Y9_FrameStrobe_O[14] ,
    \Tile_X3Y9_FrameStrobe_O[13] ,
    \Tile_X3Y9_FrameStrobe_O[12] ,
    \Tile_X3Y9_FrameStrobe_O[11] ,
    \Tile_X3Y9_FrameStrobe_O[10] ,
    \Tile_X3Y9_FrameStrobe_O[9] ,
    \Tile_X3Y9_FrameStrobe_O[8] ,
    \Tile_X3Y9_FrameStrobe_O[7] ,
    \Tile_X3Y9_FrameStrobe_O[6] ,
    \Tile_X3Y9_FrameStrobe_O[5] ,
    \Tile_X3Y9_FrameStrobe_O[4] ,
    \Tile_X3Y9_FrameStrobe_O[3] ,
    \Tile_X3Y9_FrameStrobe_O[2] ,
    \Tile_X3Y9_FrameStrobe_O[1] ,
    \Tile_X3Y9_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X3Y9_N1BEG[3] ,
    \Tile_X3Y9_N1BEG[2] ,
    \Tile_X3Y9_N1BEG[1] ,
    \Tile_X3Y9_N1BEG[0] }),
    .N1END({\Tile_X3Y10_N1BEG[3] ,
    \Tile_X3Y10_N1BEG[2] ,
    \Tile_X3Y10_N1BEG[1] ,
    \Tile_X3Y10_N1BEG[0] }),
    .N2BEG({\Tile_X3Y9_N2BEG[7] ,
    \Tile_X3Y9_N2BEG[6] ,
    \Tile_X3Y9_N2BEG[5] ,
    \Tile_X3Y9_N2BEG[4] ,
    \Tile_X3Y9_N2BEG[3] ,
    \Tile_X3Y9_N2BEG[2] ,
    \Tile_X3Y9_N2BEG[1] ,
    \Tile_X3Y9_N2BEG[0] }),
    .N2BEGb({\Tile_X3Y9_N2BEGb[7] ,
    \Tile_X3Y9_N2BEGb[6] ,
    \Tile_X3Y9_N2BEGb[5] ,
    \Tile_X3Y9_N2BEGb[4] ,
    \Tile_X3Y9_N2BEGb[3] ,
    \Tile_X3Y9_N2BEGb[2] ,
    \Tile_X3Y9_N2BEGb[1] ,
    \Tile_X3Y9_N2BEGb[0] }),
    .N2END({\Tile_X3Y10_N2BEGb[7] ,
    \Tile_X3Y10_N2BEGb[6] ,
    \Tile_X3Y10_N2BEGb[5] ,
    \Tile_X3Y10_N2BEGb[4] ,
    \Tile_X3Y10_N2BEGb[3] ,
    \Tile_X3Y10_N2BEGb[2] ,
    \Tile_X3Y10_N2BEGb[1] ,
    \Tile_X3Y10_N2BEGb[0] }),
    .N2MID({\Tile_X3Y10_N2BEG[7] ,
    \Tile_X3Y10_N2BEG[6] ,
    \Tile_X3Y10_N2BEG[5] ,
    \Tile_X3Y10_N2BEG[4] ,
    \Tile_X3Y10_N2BEG[3] ,
    \Tile_X3Y10_N2BEG[2] ,
    \Tile_X3Y10_N2BEG[1] ,
    \Tile_X3Y10_N2BEG[0] }),
    .N4BEG({\Tile_X3Y9_N4BEG[15] ,
    \Tile_X3Y9_N4BEG[14] ,
    \Tile_X3Y9_N4BEG[13] ,
    \Tile_X3Y9_N4BEG[12] ,
    \Tile_X3Y9_N4BEG[11] ,
    \Tile_X3Y9_N4BEG[10] ,
    \Tile_X3Y9_N4BEG[9] ,
    \Tile_X3Y9_N4BEG[8] ,
    \Tile_X3Y9_N4BEG[7] ,
    \Tile_X3Y9_N4BEG[6] ,
    \Tile_X3Y9_N4BEG[5] ,
    \Tile_X3Y9_N4BEG[4] ,
    \Tile_X3Y9_N4BEG[3] ,
    \Tile_X3Y9_N4BEG[2] ,
    \Tile_X3Y9_N4BEG[1] ,
    \Tile_X3Y9_N4BEG[0] }),
    .N4END({\Tile_X3Y10_N4BEG[15] ,
    \Tile_X3Y10_N4BEG[14] ,
    \Tile_X3Y10_N4BEG[13] ,
    \Tile_X3Y10_N4BEG[12] ,
    \Tile_X3Y10_N4BEG[11] ,
    \Tile_X3Y10_N4BEG[10] ,
    \Tile_X3Y10_N4BEG[9] ,
    \Tile_X3Y10_N4BEG[8] ,
    \Tile_X3Y10_N4BEG[7] ,
    \Tile_X3Y10_N4BEG[6] ,
    \Tile_X3Y10_N4BEG[5] ,
    \Tile_X3Y10_N4BEG[4] ,
    \Tile_X3Y10_N4BEG[3] ,
    \Tile_X3Y10_N4BEG[2] ,
    \Tile_X3Y10_N4BEG[1] ,
    \Tile_X3Y10_N4BEG[0] }),
    .NN4BEG({\Tile_X3Y9_NN4BEG[15] ,
    \Tile_X3Y9_NN4BEG[14] ,
    \Tile_X3Y9_NN4BEG[13] ,
    \Tile_X3Y9_NN4BEG[12] ,
    \Tile_X3Y9_NN4BEG[11] ,
    \Tile_X3Y9_NN4BEG[10] ,
    \Tile_X3Y9_NN4BEG[9] ,
    \Tile_X3Y9_NN4BEG[8] ,
    \Tile_X3Y9_NN4BEG[7] ,
    \Tile_X3Y9_NN4BEG[6] ,
    \Tile_X3Y9_NN4BEG[5] ,
    \Tile_X3Y9_NN4BEG[4] ,
    \Tile_X3Y9_NN4BEG[3] ,
    \Tile_X3Y9_NN4BEG[2] ,
    \Tile_X3Y9_NN4BEG[1] ,
    \Tile_X3Y9_NN4BEG[0] }),
    .NN4END({\Tile_X3Y10_NN4BEG[15] ,
    \Tile_X3Y10_NN4BEG[14] ,
    \Tile_X3Y10_NN4BEG[13] ,
    \Tile_X3Y10_NN4BEG[12] ,
    \Tile_X3Y10_NN4BEG[11] ,
    \Tile_X3Y10_NN4BEG[10] ,
    \Tile_X3Y10_NN4BEG[9] ,
    \Tile_X3Y10_NN4BEG[8] ,
    \Tile_X3Y10_NN4BEG[7] ,
    \Tile_X3Y10_NN4BEG[6] ,
    \Tile_X3Y10_NN4BEG[5] ,
    \Tile_X3Y10_NN4BEG[4] ,
    \Tile_X3Y10_NN4BEG[3] ,
    \Tile_X3Y10_NN4BEG[2] ,
    \Tile_X3Y10_NN4BEG[1] ,
    \Tile_X3Y10_NN4BEG[0] }),
    .S1BEG({\Tile_X3Y9_S1BEG[3] ,
    \Tile_X3Y9_S1BEG[2] ,
    \Tile_X3Y9_S1BEG[1] ,
    \Tile_X3Y9_S1BEG[0] }),
    .S1END({\Tile_X3Y8_S1BEG[3] ,
    \Tile_X3Y8_S1BEG[2] ,
    \Tile_X3Y8_S1BEG[1] ,
    \Tile_X3Y8_S1BEG[0] }),
    .S2BEG({\Tile_X3Y9_S2BEG[7] ,
    \Tile_X3Y9_S2BEG[6] ,
    \Tile_X3Y9_S2BEG[5] ,
    \Tile_X3Y9_S2BEG[4] ,
    \Tile_X3Y9_S2BEG[3] ,
    \Tile_X3Y9_S2BEG[2] ,
    \Tile_X3Y9_S2BEG[1] ,
    \Tile_X3Y9_S2BEG[0] }),
    .S2BEGb({\Tile_X3Y9_S2BEGb[7] ,
    \Tile_X3Y9_S2BEGb[6] ,
    \Tile_X3Y9_S2BEGb[5] ,
    \Tile_X3Y9_S2BEGb[4] ,
    \Tile_X3Y9_S2BEGb[3] ,
    \Tile_X3Y9_S2BEGb[2] ,
    \Tile_X3Y9_S2BEGb[1] ,
    \Tile_X3Y9_S2BEGb[0] }),
    .S2END({\Tile_X3Y8_S2BEGb[7] ,
    \Tile_X3Y8_S2BEGb[6] ,
    \Tile_X3Y8_S2BEGb[5] ,
    \Tile_X3Y8_S2BEGb[4] ,
    \Tile_X3Y8_S2BEGb[3] ,
    \Tile_X3Y8_S2BEGb[2] ,
    \Tile_X3Y8_S2BEGb[1] ,
    \Tile_X3Y8_S2BEGb[0] }),
    .S2MID({\Tile_X3Y8_S2BEG[7] ,
    \Tile_X3Y8_S2BEG[6] ,
    \Tile_X3Y8_S2BEG[5] ,
    \Tile_X3Y8_S2BEG[4] ,
    \Tile_X3Y8_S2BEG[3] ,
    \Tile_X3Y8_S2BEG[2] ,
    \Tile_X3Y8_S2BEG[1] ,
    \Tile_X3Y8_S2BEG[0] }),
    .S4BEG({\Tile_X3Y9_S4BEG[15] ,
    \Tile_X3Y9_S4BEG[14] ,
    \Tile_X3Y9_S4BEG[13] ,
    \Tile_X3Y9_S4BEG[12] ,
    \Tile_X3Y9_S4BEG[11] ,
    \Tile_X3Y9_S4BEG[10] ,
    \Tile_X3Y9_S4BEG[9] ,
    \Tile_X3Y9_S4BEG[8] ,
    \Tile_X3Y9_S4BEG[7] ,
    \Tile_X3Y9_S4BEG[6] ,
    \Tile_X3Y9_S4BEG[5] ,
    \Tile_X3Y9_S4BEG[4] ,
    \Tile_X3Y9_S4BEG[3] ,
    \Tile_X3Y9_S4BEG[2] ,
    \Tile_X3Y9_S4BEG[1] ,
    \Tile_X3Y9_S4BEG[0] }),
    .S4END({\Tile_X3Y8_S4BEG[15] ,
    \Tile_X3Y8_S4BEG[14] ,
    \Tile_X3Y8_S4BEG[13] ,
    \Tile_X3Y8_S4BEG[12] ,
    \Tile_X3Y8_S4BEG[11] ,
    \Tile_X3Y8_S4BEG[10] ,
    \Tile_X3Y8_S4BEG[9] ,
    \Tile_X3Y8_S4BEG[8] ,
    \Tile_X3Y8_S4BEG[7] ,
    \Tile_X3Y8_S4BEG[6] ,
    \Tile_X3Y8_S4BEG[5] ,
    \Tile_X3Y8_S4BEG[4] ,
    \Tile_X3Y8_S4BEG[3] ,
    \Tile_X3Y8_S4BEG[2] ,
    \Tile_X3Y8_S4BEG[1] ,
    \Tile_X3Y8_S4BEG[0] }),
    .SS4BEG({\Tile_X3Y9_SS4BEG[15] ,
    \Tile_X3Y9_SS4BEG[14] ,
    \Tile_X3Y9_SS4BEG[13] ,
    \Tile_X3Y9_SS4BEG[12] ,
    \Tile_X3Y9_SS4BEG[11] ,
    \Tile_X3Y9_SS4BEG[10] ,
    \Tile_X3Y9_SS4BEG[9] ,
    \Tile_X3Y9_SS4BEG[8] ,
    \Tile_X3Y9_SS4BEG[7] ,
    \Tile_X3Y9_SS4BEG[6] ,
    \Tile_X3Y9_SS4BEG[5] ,
    \Tile_X3Y9_SS4BEG[4] ,
    \Tile_X3Y9_SS4BEG[3] ,
    \Tile_X3Y9_SS4BEG[2] ,
    \Tile_X3Y9_SS4BEG[1] ,
    \Tile_X3Y9_SS4BEG[0] }),
    .SS4END({\Tile_X3Y8_SS4BEG[15] ,
    \Tile_X3Y8_SS4BEG[14] ,
    \Tile_X3Y8_SS4BEG[13] ,
    \Tile_X3Y8_SS4BEG[12] ,
    \Tile_X3Y8_SS4BEG[11] ,
    \Tile_X3Y8_SS4BEG[10] ,
    \Tile_X3Y8_SS4BEG[9] ,
    \Tile_X3Y8_SS4BEG[8] ,
    \Tile_X3Y8_SS4BEG[7] ,
    \Tile_X3Y8_SS4BEG[6] ,
    \Tile_X3Y8_SS4BEG[5] ,
    \Tile_X3Y8_SS4BEG[4] ,
    \Tile_X3Y8_SS4BEG[3] ,
    \Tile_X3Y8_SS4BEG[2] ,
    \Tile_X3Y8_SS4BEG[1] ,
    \Tile_X3Y8_SS4BEG[0] }),
    .W1BEG({\Tile_X3Y9_W1BEG[3] ,
    \Tile_X3Y9_W1BEG[2] ,
    \Tile_X3Y9_W1BEG[1] ,
    \Tile_X3Y9_W1BEG[0] }),
    .W1END({\Tile_X4Y9_W1BEG[3] ,
    \Tile_X4Y9_W1BEG[2] ,
    \Tile_X4Y9_W1BEG[1] ,
    \Tile_X4Y9_W1BEG[0] }),
    .W2BEG({\Tile_X3Y9_W2BEG[7] ,
    \Tile_X3Y9_W2BEG[6] ,
    \Tile_X3Y9_W2BEG[5] ,
    \Tile_X3Y9_W2BEG[4] ,
    \Tile_X3Y9_W2BEG[3] ,
    \Tile_X3Y9_W2BEG[2] ,
    \Tile_X3Y9_W2BEG[1] ,
    \Tile_X3Y9_W2BEG[0] }),
    .W2BEGb({\Tile_X3Y9_W2BEGb[7] ,
    \Tile_X3Y9_W2BEGb[6] ,
    \Tile_X3Y9_W2BEGb[5] ,
    \Tile_X3Y9_W2BEGb[4] ,
    \Tile_X3Y9_W2BEGb[3] ,
    \Tile_X3Y9_W2BEGb[2] ,
    \Tile_X3Y9_W2BEGb[1] ,
    \Tile_X3Y9_W2BEGb[0] }),
    .W2END({\Tile_X4Y9_W2BEGb[7] ,
    \Tile_X4Y9_W2BEGb[6] ,
    \Tile_X4Y9_W2BEGb[5] ,
    \Tile_X4Y9_W2BEGb[4] ,
    \Tile_X4Y9_W2BEGb[3] ,
    \Tile_X4Y9_W2BEGb[2] ,
    \Tile_X4Y9_W2BEGb[1] ,
    \Tile_X4Y9_W2BEGb[0] }),
    .W2MID({\Tile_X4Y9_W2BEG[7] ,
    \Tile_X4Y9_W2BEG[6] ,
    \Tile_X4Y9_W2BEG[5] ,
    \Tile_X4Y9_W2BEG[4] ,
    \Tile_X4Y9_W2BEG[3] ,
    \Tile_X4Y9_W2BEG[2] ,
    \Tile_X4Y9_W2BEG[1] ,
    \Tile_X4Y9_W2BEG[0] }),
    .W6BEG({\Tile_X3Y9_W6BEG[11] ,
    \Tile_X3Y9_W6BEG[10] ,
    \Tile_X3Y9_W6BEG[9] ,
    \Tile_X3Y9_W6BEG[8] ,
    \Tile_X3Y9_W6BEG[7] ,
    \Tile_X3Y9_W6BEG[6] ,
    \Tile_X3Y9_W6BEG[5] ,
    \Tile_X3Y9_W6BEG[4] ,
    \Tile_X3Y9_W6BEG[3] ,
    \Tile_X3Y9_W6BEG[2] ,
    \Tile_X3Y9_W6BEG[1] ,
    \Tile_X3Y9_W6BEG[0] }),
    .W6END({\Tile_X4Y9_W6BEG[11] ,
    \Tile_X4Y9_W6BEG[10] ,
    \Tile_X4Y9_W6BEG[9] ,
    \Tile_X4Y9_W6BEG[8] ,
    \Tile_X4Y9_W6BEG[7] ,
    \Tile_X4Y9_W6BEG[6] ,
    \Tile_X4Y9_W6BEG[5] ,
    \Tile_X4Y9_W6BEG[4] ,
    \Tile_X4Y9_W6BEG[3] ,
    \Tile_X4Y9_W6BEG[2] ,
    \Tile_X4Y9_W6BEG[1] ,
    \Tile_X4Y9_W6BEG[0] }),
    .WW4BEG({\Tile_X3Y9_WW4BEG[15] ,
    \Tile_X3Y9_WW4BEG[14] ,
    \Tile_X3Y9_WW4BEG[13] ,
    \Tile_X3Y9_WW4BEG[12] ,
    \Tile_X3Y9_WW4BEG[11] ,
    \Tile_X3Y9_WW4BEG[10] ,
    \Tile_X3Y9_WW4BEG[9] ,
    \Tile_X3Y9_WW4BEG[8] ,
    \Tile_X3Y9_WW4BEG[7] ,
    \Tile_X3Y9_WW4BEG[6] ,
    \Tile_X3Y9_WW4BEG[5] ,
    \Tile_X3Y9_WW4BEG[4] ,
    \Tile_X3Y9_WW4BEG[3] ,
    \Tile_X3Y9_WW4BEG[2] ,
    \Tile_X3Y9_WW4BEG[1] ,
    \Tile_X3Y9_WW4BEG[0] }),
    .WW4END({\Tile_X4Y9_WW4BEG[15] ,
    \Tile_X4Y9_WW4BEG[14] ,
    \Tile_X4Y9_WW4BEG[13] ,
    \Tile_X4Y9_WW4BEG[12] ,
    \Tile_X4Y9_WW4BEG[11] ,
    \Tile_X4Y9_WW4BEG[10] ,
    \Tile_X4Y9_WW4BEG[9] ,
    \Tile_X4Y9_WW4BEG[8] ,
    \Tile_X4Y9_WW4BEG[7] ,
    \Tile_X4Y9_WW4BEG[6] ,
    \Tile_X4Y9_WW4BEG[5] ,
    \Tile_X4Y9_WW4BEG[4] ,
    \Tile_X4Y9_WW4BEG[3] ,
    \Tile_X4Y9_WW4BEG[2] ,
    \Tile_X4Y9_WW4BEG[1] ,
    \Tile_X4Y9_WW4BEG[0] }));
 N_term_single2 Tile_X4Y0_N_term_single2 (.UserCLK(Tile_X4Y1_UserCLKo),
    .UserCLKo(Tile_X4Y0_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .FrameData({\Tile_X3Y0_FrameData_O[31] ,
    \Tile_X3Y0_FrameData_O[30] ,
    \Tile_X3Y0_FrameData_O[29] ,
    \Tile_X3Y0_FrameData_O[28] ,
    \Tile_X3Y0_FrameData_O[27] ,
    \Tile_X3Y0_FrameData_O[26] ,
    \Tile_X3Y0_FrameData_O[25] ,
    \Tile_X3Y0_FrameData_O[24] ,
    \Tile_X3Y0_FrameData_O[23] ,
    \Tile_X3Y0_FrameData_O[22] ,
    \Tile_X3Y0_FrameData_O[21] ,
    \Tile_X3Y0_FrameData_O[20] ,
    \Tile_X3Y0_FrameData_O[19] ,
    \Tile_X3Y0_FrameData_O[18] ,
    \Tile_X3Y0_FrameData_O[17] ,
    \Tile_X3Y0_FrameData_O[16] ,
    \Tile_X3Y0_FrameData_O[15] ,
    \Tile_X3Y0_FrameData_O[14] ,
    \Tile_X3Y0_FrameData_O[13] ,
    \Tile_X3Y0_FrameData_O[12] ,
    \Tile_X3Y0_FrameData_O[11] ,
    \Tile_X3Y0_FrameData_O[10] ,
    \Tile_X3Y0_FrameData_O[9] ,
    \Tile_X3Y0_FrameData_O[8] ,
    \Tile_X3Y0_FrameData_O[7] ,
    \Tile_X3Y0_FrameData_O[6] ,
    \Tile_X3Y0_FrameData_O[5] ,
    \Tile_X3Y0_FrameData_O[4] ,
    \Tile_X3Y0_FrameData_O[3] ,
    \Tile_X3Y0_FrameData_O[2] ,
    \Tile_X3Y0_FrameData_O[1] ,
    \Tile_X3Y0_FrameData_O[0] }),
    .FrameData_O({\Tile_X4Y0_FrameData_O[31] ,
    \Tile_X4Y0_FrameData_O[30] ,
    \Tile_X4Y0_FrameData_O[29] ,
    \Tile_X4Y0_FrameData_O[28] ,
    \Tile_X4Y0_FrameData_O[27] ,
    \Tile_X4Y0_FrameData_O[26] ,
    \Tile_X4Y0_FrameData_O[25] ,
    \Tile_X4Y0_FrameData_O[24] ,
    \Tile_X4Y0_FrameData_O[23] ,
    \Tile_X4Y0_FrameData_O[22] ,
    \Tile_X4Y0_FrameData_O[21] ,
    \Tile_X4Y0_FrameData_O[20] ,
    \Tile_X4Y0_FrameData_O[19] ,
    \Tile_X4Y0_FrameData_O[18] ,
    \Tile_X4Y0_FrameData_O[17] ,
    \Tile_X4Y0_FrameData_O[16] ,
    \Tile_X4Y0_FrameData_O[15] ,
    \Tile_X4Y0_FrameData_O[14] ,
    \Tile_X4Y0_FrameData_O[13] ,
    \Tile_X4Y0_FrameData_O[12] ,
    \Tile_X4Y0_FrameData_O[11] ,
    \Tile_X4Y0_FrameData_O[10] ,
    \Tile_X4Y0_FrameData_O[9] ,
    \Tile_X4Y0_FrameData_O[8] ,
    \Tile_X4Y0_FrameData_O[7] ,
    \Tile_X4Y0_FrameData_O[6] ,
    \Tile_X4Y0_FrameData_O[5] ,
    \Tile_X4Y0_FrameData_O[4] ,
    \Tile_X4Y0_FrameData_O[3] ,
    \Tile_X4Y0_FrameData_O[2] ,
    \Tile_X4Y0_FrameData_O[1] ,
    \Tile_X4Y0_FrameData_O[0] }),
    .FrameStrobe({\Tile_X4Y1_FrameStrobe_O[19] ,
    \Tile_X4Y1_FrameStrobe_O[18] ,
    \Tile_X4Y1_FrameStrobe_O[17] ,
    \Tile_X4Y1_FrameStrobe_O[16] ,
    \Tile_X4Y1_FrameStrobe_O[15] ,
    \Tile_X4Y1_FrameStrobe_O[14] ,
    \Tile_X4Y1_FrameStrobe_O[13] ,
    \Tile_X4Y1_FrameStrobe_O[12] ,
    \Tile_X4Y1_FrameStrobe_O[11] ,
    \Tile_X4Y1_FrameStrobe_O[10] ,
    \Tile_X4Y1_FrameStrobe_O[9] ,
    \Tile_X4Y1_FrameStrobe_O[8] ,
    \Tile_X4Y1_FrameStrobe_O[7] ,
    \Tile_X4Y1_FrameStrobe_O[6] ,
    \Tile_X4Y1_FrameStrobe_O[5] ,
    \Tile_X4Y1_FrameStrobe_O[4] ,
    \Tile_X4Y1_FrameStrobe_O[3] ,
    \Tile_X4Y1_FrameStrobe_O[2] ,
    \Tile_X4Y1_FrameStrobe_O[1] ,
    \Tile_X4Y1_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X4Y0_FrameStrobe_O[19] ,
    \Tile_X4Y0_FrameStrobe_O[18] ,
    \Tile_X4Y0_FrameStrobe_O[17] ,
    \Tile_X4Y0_FrameStrobe_O[16] ,
    \Tile_X4Y0_FrameStrobe_O[15] ,
    \Tile_X4Y0_FrameStrobe_O[14] ,
    \Tile_X4Y0_FrameStrobe_O[13] ,
    \Tile_X4Y0_FrameStrobe_O[12] ,
    \Tile_X4Y0_FrameStrobe_O[11] ,
    \Tile_X4Y0_FrameStrobe_O[10] ,
    \Tile_X4Y0_FrameStrobe_O[9] ,
    \Tile_X4Y0_FrameStrobe_O[8] ,
    \Tile_X4Y0_FrameStrobe_O[7] ,
    \Tile_X4Y0_FrameStrobe_O[6] ,
    \Tile_X4Y0_FrameStrobe_O[5] ,
    \Tile_X4Y0_FrameStrobe_O[4] ,
    \Tile_X4Y0_FrameStrobe_O[3] ,
    \Tile_X4Y0_FrameStrobe_O[2] ,
    \Tile_X4Y0_FrameStrobe_O[1] ,
    \Tile_X4Y0_FrameStrobe_O[0] }),
    .N1END({\Tile_X4Y1_N1BEG[3] ,
    \Tile_X4Y1_N1BEG[2] ,
    \Tile_X4Y1_N1BEG[1] ,
    \Tile_X4Y1_N1BEG[0] }),
    .N2END({\Tile_X4Y1_N2BEGb[7] ,
    \Tile_X4Y1_N2BEGb[6] ,
    \Tile_X4Y1_N2BEGb[5] ,
    \Tile_X4Y1_N2BEGb[4] ,
    \Tile_X4Y1_N2BEGb[3] ,
    \Tile_X4Y1_N2BEGb[2] ,
    \Tile_X4Y1_N2BEGb[1] ,
    \Tile_X4Y1_N2BEGb[0] }),
    .N2MID({\Tile_X4Y1_N2BEG[7] ,
    \Tile_X4Y1_N2BEG[6] ,
    \Tile_X4Y1_N2BEG[5] ,
    \Tile_X4Y1_N2BEG[4] ,
    \Tile_X4Y1_N2BEG[3] ,
    \Tile_X4Y1_N2BEG[2] ,
    \Tile_X4Y1_N2BEG[1] ,
    \Tile_X4Y1_N2BEG[0] }),
    .N4END({\Tile_X4Y1_N4BEG[15] ,
    \Tile_X4Y1_N4BEG[14] ,
    \Tile_X4Y1_N4BEG[13] ,
    \Tile_X4Y1_N4BEG[12] ,
    \Tile_X4Y1_N4BEG[11] ,
    \Tile_X4Y1_N4BEG[10] ,
    \Tile_X4Y1_N4BEG[9] ,
    \Tile_X4Y1_N4BEG[8] ,
    \Tile_X4Y1_N4BEG[7] ,
    \Tile_X4Y1_N4BEG[6] ,
    \Tile_X4Y1_N4BEG[5] ,
    \Tile_X4Y1_N4BEG[4] ,
    \Tile_X4Y1_N4BEG[3] ,
    \Tile_X4Y1_N4BEG[2] ,
    \Tile_X4Y1_N4BEG[1] ,
    \Tile_X4Y1_N4BEG[0] }),
    .NN4END({\Tile_X4Y1_NN4BEG[15] ,
    \Tile_X4Y1_NN4BEG[14] ,
    \Tile_X4Y1_NN4BEG[13] ,
    \Tile_X4Y1_NN4BEG[12] ,
    \Tile_X4Y1_NN4BEG[11] ,
    \Tile_X4Y1_NN4BEG[10] ,
    \Tile_X4Y1_NN4BEG[9] ,
    \Tile_X4Y1_NN4BEG[8] ,
    \Tile_X4Y1_NN4BEG[7] ,
    \Tile_X4Y1_NN4BEG[6] ,
    \Tile_X4Y1_NN4BEG[5] ,
    \Tile_X4Y1_NN4BEG[4] ,
    \Tile_X4Y1_NN4BEG[3] ,
    \Tile_X4Y1_NN4BEG[2] ,
    \Tile_X4Y1_NN4BEG[1] ,
    \Tile_X4Y1_NN4BEG[0] }),
    .S1BEG({\Tile_X4Y0_S1BEG[3] ,
    \Tile_X4Y0_S1BEG[2] ,
    \Tile_X4Y0_S1BEG[1] ,
    \Tile_X4Y0_S1BEG[0] }),
    .S2BEG({\Tile_X4Y0_S2BEG[7] ,
    \Tile_X4Y0_S2BEG[6] ,
    \Tile_X4Y0_S2BEG[5] ,
    \Tile_X4Y0_S2BEG[4] ,
    \Tile_X4Y0_S2BEG[3] ,
    \Tile_X4Y0_S2BEG[2] ,
    \Tile_X4Y0_S2BEG[1] ,
    \Tile_X4Y0_S2BEG[0] }),
    .S2BEGb({\Tile_X4Y0_S2BEGb[7] ,
    \Tile_X4Y0_S2BEGb[6] ,
    \Tile_X4Y0_S2BEGb[5] ,
    \Tile_X4Y0_S2BEGb[4] ,
    \Tile_X4Y0_S2BEGb[3] ,
    \Tile_X4Y0_S2BEGb[2] ,
    \Tile_X4Y0_S2BEGb[1] ,
    \Tile_X4Y0_S2BEGb[0] }),
    .S4BEG({\Tile_X4Y0_S4BEG[15] ,
    \Tile_X4Y0_S4BEG[14] ,
    \Tile_X4Y0_S4BEG[13] ,
    \Tile_X4Y0_S4BEG[12] ,
    \Tile_X4Y0_S4BEG[11] ,
    \Tile_X4Y0_S4BEG[10] ,
    \Tile_X4Y0_S4BEG[9] ,
    \Tile_X4Y0_S4BEG[8] ,
    \Tile_X4Y0_S4BEG[7] ,
    \Tile_X4Y0_S4BEG[6] ,
    \Tile_X4Y0_S4BEG[5] ,
    \Tile_X4Y0_S4BEG[4] ,
    \Tile_X4Y0_S4BEG[3] ,
    \Tile_X4Y0_S4BEG[2] ,
    \Tile_X4Y0_S4BEG[1] ,
    \Tile_X4Y0_S4BEG[0] }),
    .SS4BEG({\Tile_X4Y0_SS4BEG[15] ,
    \Tile_X4Y0_SS4BEG[14] ,
    \Tile_X4Y0_SS4BEG[13] ,
    \Tile_X4Y0_SS4BEG[12] ,
    \Tile_X4Y0_SS4BEG[11] ,
    \Tile_X4Y0_SS4BEG[10] ,
    \Tile_X4Y0_SS4BEG[9] ,
    \Tile_X4Y0_SS4BEG[8] ,
    \Tile_X4Y0_SS4BEG[7] ,
    \Tile_X4Y0_SS4BEG[6] ,
    \Tile_X4Y0_SS4BEG[5] ,
    \Tile_X4Y0_SS4BEG[4] ,
    \Tile_X4Y0_SS4BEG[3] ,
    \Tile_X4Y0_SS4BEG[2] ,
    \Tile_X4Y0_SS4BEG[1] ,
    \Tile_X4Y0_SS4BEG[0] }));
 RegFile Tile_X4Y10_RegFile (.UserCLK(Tile_X4Y11_UserCLKo),
    .UserCLKo(Tile_X4Y10_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X4Y10_E1BEG[3] ,
    \Tile_X4Y10_E1BEG[2] ,
    \Tile_X4Y10_E1BEG[1] ,
    \Tile_X4Y10_E1BEG[0] }),
    .E1END({\Tile_X3Y10_E1BEG[3] ,
    \Tile_X3Y10_E1BEG[2] ,
    \Tile_X3Y10_E1BEG[1] ,
    \Tile_X3Y10_E1BEG[0] }),
    .E2BEG({\Tile_X4Y10_E2BEG[7] ,
    \Tile_X4Y10_E2BEG[6] ,
    \Tile_X4Y10_E2BEG[5] ,
    \Tile_X4Y10_E2BEG[4] ,
    \Tile_X4Y10_E2BEG[3] ,
    \Tile_X4Y10_E2BEG[2] ,
    \Tile_X4Y10_E2BEG[1] ,
    \Tile_X4Y10_E2BEG[0] }),
    .E2BEGb({\Tile_X4Y10_E2BEGb[7] ,
    \Tile_X4Y10_E2BEGb[6] ,
    \Tile_X4Y10_E2BEGb[5] ,
    \Tile_X4Y10_E2BEGb[4] ,
    \Tile_X4Y10_E2BEGb[3] ,
    \Tile_X4Y10_E2BEGb[2] ,
    \Tile_X4Y10_E2BEGb[1] ,
    \Tile_X4Y10_E2BEGb[0] }),
    .E2END({\Tile_X3Y10_E2BEGb[7] ,
    \Tile_X3Y10_E2BEGb[6] ,
    \Tile_X3Y10_E2BEGb[5] ,
    \Tile_X3Y10_E2BEGb[4] ,
    \Tile_X3Y10_E2BEGb[3] ,
    \Tile_X3Y10_E2BEGb[2] ,
    \Tile_X3Y10_E2BEGb[1] ,
    \Tile_X3Y10_E2BEGb[0] }),
    .E2MID({\Tile_X3Y10_E2BEG[7] ,
    \Tile_X3Y10_E2BEG[6] ,
    \Tile_X3Y10_E2BEG[5] ,
    \Tile_X3Y10_E2BEG[4] ,
    \Tile_X3Y10_E2BEG[3] ,
    \Tile_X3Y10_E2BEG[2] ,
    \Tile_X3Y10_E2BEG[1] ,
    \Tile_X3Y10_E2BEG[0] }),
    .E6BEG({\Tile_X4Y10_E6BEG[11] ,
    \Tile_X4Y10_E6BEG[10] ,
    \Tile_X4Y10_E6BEG[9] ,
    \Tile_X4Y10_E6BEG[8] ,
    \Tile_X4Y10_E6BEG[7] ,
    \Tile_X4Y10_E6BEG[6] ,
    \Tile_X4Y10_E6BEG[5] ,
    \Tile_X4Y10_E6BEG[4] ,
    \Tile_X4Y10_E6BEG[3] ,
    \Tile_X4Y10_E6BEG[2] ,
    \Tile_X4Y10_E6BEG[1] ,
    \Tile_X4Y10_E6BEG[0] }),
    .E6END({\Tile_X3Y10_E6BEG[11] ,
    \Tile_X3Y10_E6BEG[10] ,
    \Tile_X3Y10_E6BEG[9] ,
    \Tile_X3Y10_E6BEG[8] ,
    \Tile_X3Y10_E6BEG[7] ,
    \Tile_X3Y10_E6BEG[6] ,
    \Tile_X3Y10_E6BEG[5] ,
    \Tile_X3Y10_E6BEG[4] ,
    \Tile_X3Y10_E6BEG[3] ,
    \Tile_X3Y10_E6BEG[2] ,
    \Tile_X3Y10_E6BEG[1] ,
    \Tile_X3Y10_E6BEG[0] }),
    .EE4BEG({\Tile_X4Y10_EE4BEG[15] ,
    \Tile_X4Y10_EE4BEG[14] ,
    \Tile_X4Y10_EE4BEG[13] ,
    \Tile_X4Y10_EE4BEG[12] ,
    \Tile_X4Y10_EE4BEG[11] ,
    \Tile_X4Y10_EE4BEG[10] ,
    \Tile_X4Y10_EE4BEG[9] ,
    \Tile_X4Y10_EE4BEG[8] ,
    \Tile_X4Y10_EE4BEG[7] ,
    \Tile_X4Y10_EE4BEG[6] ,
    \Tile_X4Y10_EE4BEG[5] ,
    \Tile_X4Y10_EE4BEG[4] ,
    \Tile_X4Y10_EE4BEG[3] ,
    \Tile_X4Y10_EE4BEG[2] ,
    \Tile_X4Y10_EE4BEG[1] ,
    \Tile_X4Y10_EE4BEG[0] }),
    .EE4END({\Tile_X3Y10_EE4BEG[15] ,
    \Tile_X3Y10_EE4BEG[14] ,
    \Tile_X3Y10_EE4BEG[13] ,
    \Tile_X3Y10_EE4BEG[12] ,
    \Tile_X3Y10_EE4BEG[11] ,
    \Tile_X3Y10_EE4BEG[10] ,
    \Tile_X3Y10_EE4BEG[9] ,
    \Tile_X3Y10_EE4BEG[8] ,
    \Tile_X3Y10_EE4BEG[7] ,
    \Tile_X3Y10_EE4BEG[6] ,
    \Tile_X3Y10_EE4BEG[5] ,
    \Tile_X3Y10_EE4BEG[4] ,
    \Tile_X3Y10_EE4BEG[3] ,
    \Tile_X3Y10_EE4BEG[2] ,
    \Tile_X3Y10_EE4BEG[1] ,
    \Tile_X3Y10_EE4BEG[0] }),
    .FrameData({\Tile_X3Y10_FrameData_O[31] ,
    \Tile_X3Y10_FrameData_O[30] ,
    \Tile_X3Y10_FrameData_O[29] ,
    \Tile_X3Y10_FrameData_O[28] ,
    \Tile_X3Y10_FrameData_O[27] ,
    \Tile_X3Y10_FrameData_O[26] ,
    \Tile_X3Y10_FrameData_O[25] ,
    \Tile_X3Y10_FrameData_O[24] ,
    \Tile_X3Y10_FrameData_O[23] ,
    \Tile_X3Y10_FrameData_O[22] ,
    \Tile_X3Y10_FrameData_O[21] ,
    \Tile_X3Y10_FrameData_O[20] ,
    \Tile_X3Y10_FrameData_O[19] ,
    \Tile_X3Y10_FrameData_O[18] ,
    \Tile_X3Y10_FrameData_O[17] ,
    \Tile_X3Y10_FrameData_O[16] ,
    \Tile_X3Y10_FrameData_O[15] ,
    \Tile_X3Y10_FrameData_O[14] ,
    \Tile_X3Y10_FrameData_O[13] ,
    \Tile_X3Y10_FrameData_O[12] ,
    \Tile_X3Y10_FrameData_O[11] ,
    \Tile_X3Y10_FrameData_O[10] ,
    \Tile_X3Y10_FrameData_O[9] ,
    \Tile_X3Y10_FrameData_O[8] ,
    \Tile_X3Y10_FrameData_O[7] ,
    \Tile_X3Y10_FrameData_O[6] ,
    \Tile_X3Y10_FrameData_O[5] ,
    \Tile_X3Y10_FrameData_O[4] ,
    \Tile_X3Y10_FrameData_O[3] ,
    \Tile_X3Y10_FrameData_O[2] ,
    \Tile_X3Y10_FrameData_O[1] ,
    \Tile_X3Y10_FrameData_O[0] }),
    .FrameData_O({\Tile_X4Y10_FrameData_O[31] ,
    \Tile_X4Y10_FrameData_O[30] ,
    \Tile_X4Y10_FrameData_O[29] ,
    \Tile_X4Y10_FrameData_O[28] ,
    \Tile_X4Y10_FrameData_O[27] ,
    \Tile_X4Y10_FrameData_O[26] ,
    \Tile_X4Y10_FrameData_O[25] ,
    \Tile_X4Y10_FrameData_O[24] ,
    \Tile_X4Y10_FrameData_O[23] ,
    \Tile_X4Y10_FrameData_O[22] ,
    \Tile_X4Y10_FrameData_O[21] ,
    \Tile_X4Y10_FrameData_O[20] ,
    \Tile_X4Y10_FrameData_O[19] ,
    \Tile_X4Y10_FrameData_O[18] ,
    \Tile_X4Y10_FrameData_O[17] ,
    \Tile_X4Y10_FrameData_O[16] ,
    \Tile_X4Y10_FrameData_O[15] ,
    \Tile_X4Y10_FrameData_O[14] ,
    \Tile_X4Y10_FrameData_O[13] ,
    \Tile_X4Y10_FrameData_O[12] ,
    \Tile_X4Y10_FrameData_O[11] ,
    \Tile_X4Y10_FrameData_O[10] ,
    \Tile_X4Y10_FrameData_O[9] ,
    \Tile_X4Y10_FrameData_O[8] ,
    \Tile_X4Y10_FrameData_O[7] ,
    \Tile_X4Y10_FrameData_O[6] ,
    \Tile_X4Y10_FrameData_O[5] ,
    \Tile_X4Y10_FrameData_O[4] ,
    \Tile_X4Y10_FrameData_O[3] ,
    \Tile_X4Y10_FrameData_O[2] ,
    \Tile_X4Y10_FrameData_O[1] ,
    \Tile_X4Y10_FrameData_O[0] }),
    .FrameStrobe({\Tile_X4Y11_FrameStrobe_O[19] ,
    \Tile_X4Y11_FrameStrobe_O[18] ,
    \Tile_X4Y11_FrameStrobe_O[17] ,
    \Tile_X4Y11_FrameStrobe_O[16] ,
    \Tile_X4Y11_FrameStrobe_O[15] ,
    \Tile_X4Y11_FrameStrobe_O[14] ,
    \Tile_X4Y11_FrameStrobe_O[13] ,
    \Tile_X4Y11_FrameStrobe_O[12] ,
    \Tile_X4Y11_FrameStrobe_O[11] ,
    \Tile_X4Y11_FrameStrobe_O[10] ,
    \Tile_X4Y11_FrameStrobe_O[9] ,
    \Tile_X4Y11_FrameStrobe_O[8] ,
    \Tile_X4Y11_FrameStrobe_O[7] ,
    \Tile_X4Y11_FrameStrobe_O[6] ,
    \Tile_X4Y11_FrameStrobe_O[5] ,
    \Tile_X4Y11_FrameStrobe_O[4] ,
    \Tile_X4Y11_FrameStrobe_O[3] ,
    \Tile_X4Y11_FrameStrobe_O[2] ,
    \Tile_X4Y11_FrameStrobe_O[1] ,
    \Tile_X4Y11_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X4Y10_FrameStrobe_O[19] ,
    \Tile_X4Y10_FrameStrobe_O[18] ,
    \Tile_X4Y10_FrameStrobe_O[17] ,
    \Tile_X4Y10_FrameStrobe_O[16] ,
    \Tile_X4Y10_FrameStrobe_O[15] ,
    \Tile_X4Y10_FrameStrobe_O[14] ,
    \Tile_X4Y10_FrameStrobe_O[13] ,
    \Tile_X4Y10_FrameStrobe_O[12] ,
    \Tile_X4Y10_FrameStrobe_O[11] ,
    \Tile_X4Y10_FrameStrobe_O[10] ,
    \Tile_X4Y10_FrameStrobe_O[9] ,
    \Tile_X4Y10_FrameStrobe_O[8] ,
    \Tile_X4Y10_FrameStrobe_O[7] ,
    \Tile_X4Y10_FrameStrobe_O[6] ,
    \Tile_X4Y10_FrameStrobe_O[5] ,
    \Tile_X4Y10_FrameStrobe_O[4] ,
    \Tile_X4Y10_FrameStrobe_O[3] ,
    \Tile_X4Y10_FrameStrobe_O[2] ,
    \Tile_X4Y10_FrameStrobe_O[1] ,
    \Tile_X4Y10_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X4Y10_N1BEG[3] ,
    \Tile_X4Y10_N1BEG[2] ,
    \Tile_X4Y10_N1BEG[1] ,
    \Tile_X4Y10_N1BEG[0] }),
    .N1END({\Tile_X4Y11_N1BEG[3] ,
    \Tile_X4Y11_N1BEG[2] ,
    \Tile_X4Y11_N1BEG[1] ,
    \Tile_X4Y11_N1BEG[0] }),
    .N2BEG({\Tile_X4Y10_N2BEG[7] ,
    \Tile_X4Y10_N2BEG[6] ,
    \Tile_X4Y10_N2BEG[5] ,
    \Tile_X4Y10_N2BEG[4] ,
    \Tile_X4Y10_N2BEG[3] ,
    \Tile_X4Y10_N2BEG[2] ,
    \Tile_X4Y10_N2BEG[1] ,
    \Tile_X4Y10_N2BEG[0] }),
    .N2BEGb({\Tile_X4Y10_N2BEGb[7] ,
    \Tile_X4Y10_N2BEGb[6] ,
    \Tile_X4Y10_N2BEGb[5] ,
    \Tile_X4Y10_N2BEGb[4] ,
    \Tile_X4Y10_N2BEGb[3] ,
    \Tile_X4Y10_N2BEGb[2] ,
    \Tile_X4Y10_N2BEGb[1] ,
    \Tile_X4Y10_N2BEGb[0] }),
    .N2END({\Tile_X4Y11_N2BEGb[7] ,
    \Tile_X4Y11_N2BEGb[6] ,
    \Tile_X4Y11_N2BEGb[5] ,
    \Tile_X4Y11_N2BEGb[4] ,
    \Tile_X4Y11_N2BEGb[3] ,
    \Tile_X4Y11_N2BEGb[2] ,
    \Tile_X4Y11_N2BEGb[1] ,
    \Tile_X4Y11_N2BEGb[0] }),
    .N2MID({\Tile_X4Y11_N2BEG[7] ,
    \Tile_X4Y11_N2BEG[6] ,
    \Tile_X4Y11_N2BEG[5] ,
    \Tile_X4Y11_N2BEG[4] ,
    \Tile_X4Y11_N2BEG[3] ,
    \Tile_X4Y11_N2BEG[2] ,
    \Tile_X4Y11_N2BEG[1] ,
    \Tile_X4Y11_N2BEG[0] }),
    .N4BEG({\Tile_X4Y10_N4BEG[15] ,
    \Tile_X4Y10_N4BEG[14] ,
    \Tile_X4Y10_N4BEG[13] ,
    \Tile_X4Y10_N4BEG[12] ,
    \Tile_X4Y10_N4BEG[11] ,
    \Tile_X4Y10_N4BEG[10] ,
    \Tile_X4Y10_N4BEG[9] ,
    \Tile_X4Y10_N4BEG[8] ,
    \Tile_X4Y10_N4BEG[7] ,
    \Tile_X4Y10_N4BEG[6] ,
    \Tile_X4Y10_N4BEG[5] ,
    \Tile_X4Y10_N4BEG[4] ,
    \Tile_X4Y10_N4BEG[3] ,
    \Tile_X4Y10_N4BEG[2] ,
    \Tile_X4Y10_N4BEG[1] ,
    \Tile_X4Y10_N4BEG[0] }),
    .N4END({\Tile_X4Y11_N4BEG[15] ,
    \Tile_X4Y11_N4BEG[14] ,
    \Tile_X4Y11_N4BEG[13] ,
    \Tile_X4Y11_N4BEG[12] ,
    \Tile_X4Y11_N4BEG[11] ,
    \Tile_X4Y11_N4BEG[10] ,
    \Tile_X4Y11_N4BEG[9] ,
    \Tile_X4Y11_N4BEG[8] ,
    \Tile_X4Y11_N4BEG[7] ,
    \Tile_X4Y11_N4BEG[6] ,
    \Tile_X4Y11_N4BEG[5] ,
    \Tile_X4Y11_N4BEG[4] ,
    \Tile_X4Y11_N4BEG[3] ,
    \Tile_X4Y11_N4BEG[2] ,
    \Tile_X4Y11_N4BEG[1] ,
    \Tile_X4Y11_N4BEG[0] }),
    .NN4BEG({\Tile_X4Y10_NN4BEG[15] ,
    \Tile_X4Y10_NN4BEG[14] ,
    \Tile_X4Y10_NN4BEG[13] ,
    \Tile_X4Y10_NN4BEG[12] ,
    \Tile_X4Y10_NN4BEG[11] ,
    \Tile_X4Y10_NN4BEG[10] ,
    \Tile_X4Y10_NN4BEG[9] ,
    \Tile_X4Y10_NN4BEG[8] ,
    \Tile_X4Y10_NN4BEG[7] ,
    \Tile_X4Y10_NN4BEG[6] ,
    \Tile_X4Y10_NN4BEG[5] ,
    \Tile_X4Y10_NN4BEG[4] ,
    \Tile_X4Y10_NN4BEG[3] ,
    \Tile_X4Y10_NN4BEG[2] ,
    \Tile_X4Y10_NN4BEG[1] ,
    \Tile_X4Y10_NN4BEG[0] }),
    .NN4END({\Tile_X4Y11_NN4BEG[15] ,
    \Tile_X4Y11_NN4BEG[14] ,
    \Tile_X4Y11_NN4BEG[13] ,
    \Tile_X4Y11_NN4BEG[12] ,
    \Tile_X4Y11_NN4BEG[11] ,
    \Tile_X4Y11_NN4BEG[10] ,
    \Tile_X4Y11_NN4BEG[9] ,
    \Tile_X4Y11_NN4BEG[8] ,
    \Tile_X4Y11_NN4BEG[7] ,
    \Tile_X4Y11_NN4BEG[6] ,
    \Tile_X4Y11_NN4BEG[5] ,
    \Tile_X4Y11_NN4BEG[4] ,
    \Tile_X4Y11_NN4BEG[3] ,
    \Tile_X4Y11_NN4BEG[2] ,
    \Tile_X4Y11_NN4BEG[1] ,
    \Tile_X4Y11_NN4BEG[0] }),
    .S1BEG({\Tile_X4Y10_S1BEG[3] ,
    \Tile_X4Y10_S1BEG[2] ,
    \Tile_X4Y10_S1BEG[1] ,
    \Tile_X4Y10_S1BEG[0] }),
    .S1END({\Tile_X4Y9_S1BEG[3] ,
    \Tile_X4Y9_S1BEG[2] ,
    \Tile_X4Y9_S1BEG[1] ,
    \Tile_X4Y9_S1BEG[0] }),
    .S2BEG({\Tile_X4Y10_S2BEG[7] ,
    \Tile_X4Y10_S2BEG[6] ,
    \Tile_X4Y10_S2BEG[5] ,
    \Tile_X4Y10_S2BEG[4] ,
    \Tile_X4Y10_S2BEG[3] ,
    \Tile_X4Y10_S2BEG[2] ,
    \Tile_X4Y10_S2BEG[1] ,
    \Tile_X4Y10_S2BEG[0] }),
    .S2BEGb({\Tile_X4Y10_S2BEGb[7] ,
    \Tile_X4Y10_S2BEGb[6] ,
    \Tile_X4Y10_S2BEGb[5] ,
    \Tile_X4Y10_S2BEGb[4] ,
    \Tile_X4Y10_S2BEGb[3] ,
    \Tile_X4Y10_S2BEGb[2] ,
    \Tile_X4Y10_S2BEGb[1] ,
    \Tile_X4Y10_S2BEGb[0] }),
    .S2END({\Tile_X4Y9_S2BEGb[7] ,
    \Tile_X4Y9_S2BEGb[6] ,
    \Tile_X4Y9_S2BEGb[5] ,
    \Tile_X4Y9_S2BEGb[4] ,
    \Tile_X4Y9_S2BEGb[3] ,
    \Tile_X4Y9_S2BEGb[2] ,
    \Tile_X4Y9_S2BEGb[1] ,
    \Tile_X4Y9_S2BEGb[0] }),
    .S2MID({\Tile_X4Y9_S2BEG[7] ,
    \Tile_X4Y9_S2BEG[6] ,
    \Tile_X4Y9_S2BEG[5] ,
    \Tile_X4Y9_S2BEG[4] ,
    \Tile_X4Y9_S2BEG[3] ,
    \Tile_X4Y9_S2BEG[2] ,
    \Tile_X4Y9_S2BEG[1] ,
    \Tile_X4Y9_S2BEG[0] }),
    .S4BEG({\Tile_X4Y10_S4BEG[15] ,
    \Tile_X4Y10_S4BEG[14] ,
    \Tile_X4Y10_S4BEG[13] ,
    \Tile_X4Y10_S4BEG[12] ,
    \Tile_X4Y10_S4BEG[11] ,
    \Tile_X4Y10_S4BEG[10] ,
    \Tile_X4Y10_S4BEG[9] ,
    \Tile_X4Y10_S4BEG[8] ,
    \Tile_X4Y10_S4BEG[7] ,
    \Tile_X4Y10_S4BEG[6] ,
    \Tile_X4Y10_S4BEG[5] ,
    \Tile_X4Y10_S4BEG[4] ,
    \Tile_X4Y10_S4BEG[3] ,
    \Tile_X4Y10_S4BEG[2] ,
    \Tile_X4Y10_S4BEG[1] ,
    \Tile_X4Y10_S4BEG[0] }),
    .S4END({\Tile_X4Y9_S4BEG[15] ,
    \Tile_X4Y9_S4BEG[14] ,
    \Tile_X4Y9_S4BEG[13] ,
    \Tile_X4Y9_S4BEG[12] ,
    \Tile_X4Y9_S4BEG[11] ,
    \Tile_X4Y9_S4BEG[10] ,
    \Tile_X4Y9_S4BEG[9] ,
    \Tile_X4Y9_S4BEG[8] ,
    \Tile_X4Y9_S4BEG[7] ,
    \Tile_X4Y9_S4BEG[6] ,
    \Tile_X4Y9_S4BEG[5] ,
    \Tile_X4Y9_S4BEG[4] ,
    \Tile_X4Y9_S4BEG[3] ,
    \Tile_X4Y9_S4BEG[2] ,
    \Tile_X4Y9_S4BEG[1] ,
    \Tile_X4Y9_S4BEG[0] }),
    .SS4BEG({\Tile_X4Y10_SS4BEG[15] ,
    \Tile_X4Y10_SS4BEG[14] ,
    \Tile_X4Y10_SS4BEG[13] ,
    \Tile_X4Y10_SS4BEG[12] ,
    \Tile_X4Y10_SS4BEG[11] ,
    \Tile_X4Y10_SS4BEG[10] ,
    \Tile_X4Y10_SS4BEG[9] ,
    \Tile_X4Y10_SS4BEG[8] ,
    \Tile_X4Y10_SS4BEG[7] ,
    \Tile_X4Y10_SS4BEG[6] ,
    \Tile_X4Y10_SS4BEG[5] ,
    \Tile_X4Y10_SS4BEG[4] ,
    \Tile_X4Y10_SS4BEG[3] ,
    \Tile_X4Y10_SS4BEG[2] ,
    \Tile_X4Y10_SS4BEG[1] ,
    \Tile_X4Y10_SS4BEG[0] }),
    .SS4END({\Tile_X4Y9_SS4BEG[15] ,
    \Tile_X4Y9_SS4BEG[14] ,
    \Tile_X4Y9_SS4BEG[13] ,
    \Tile_X4Y9_SS4BEG[12] ,
    \Tile_X4Y9_SS4BEG[11] ,
    \Tile_X4Y9_SS4BEG[10] ,
    \Tile_X4Y9_SS4BEG[9] ,
    \Tile_X4Y9_SS4BEG[8] ,
    \Tile_X4Y9_SS4BEG[7] ,
    \Tile_X4Y9_SS4BEG[6] ,
    \Tile_X4Y9_SS4BEG[5] ,
    \Tile_X4Y9_SS4BEG[4] ,
    \Tile_X4Y9_SS4BEG[3] ,
    \Tile_X4Y9_SS4BEG[2] ,
    \Tile_X4Y9_SS4BEG[1] ,
    \Tile_X4Y9_SS4BEG[0] }),
    .W1BEG({\Tile_X4Y10_W1BEG[3] ,
    \Tile_X4Y10_W1BEG[2] ,
    \Tile_X4Y10_W1BEG[1] ,
    \Tile_X4Y10_W1BEG[0] }),
    .W1END({\Tile_X5Y10_W1BEG[3] ,
    \Tile_X5Y10_W1BEG[2] ,
    \Tile_X5Y10_W1BEG[1] ,
    \Tile_X5Y10_W1BEG[0] }),
    .W2BEG({\Tile_X4Y10_W2BEG[7] ,
    \Tile_X4Y10_W2BEG[6] ,
    \Tile_X4Y10_W2BEG[5] ,
    \Tile_X4Y10_W2BEG[4] ,
    \Tile_X4Y10_W2BEG[3] ,
    \Tile_X4Y10_W2BEG[2] ,
    \Tile_X4Y10_W2BEG[1] ,
    \Tile_X4Y10_W2BEG[0] }),
    .W2BEGb({\Tile_X4Y10_W2BEGb[7] ,
    \Tile_X4Y10_W2BEGb[6] ,
    \Tile_X4Y10_W2BEGb[5] ,
    \Tile_X4Y10_W2BEGb[4] ,
    \Tile_X4Y10_W2BEGb[3] ,
    \Tile_X4Y10_W2BEGb[2] ,
    \Tile_X4Y10_W2BEGb[1] ,
    \Tile_X4Y10_W2BEGb[0] }),
    .W2END({\Tile_X5Y10_W2BEGb[7] ,
    \Tile_X5Y10_W2BEGb[6] ,
    \Tile_X5Y10_W2BEGb[5] ,
    \Tile_X5Y10_W2BEGb[4] ,
    \Tile_X5Y10_W2BEGb[3] ,
    \Tile_X5Y10_W2BEGb[2] ,
    \Tile_X5Y10_W2BEGb[1] ,
    \Tile_X5Y10_W2BEGb[0] }),
    .W2MID({\Tile_X5Y10_W2BEG[7] ,
    \Tile_X5Y10_W2BEG[6] ,
    \Tile_X5Y10_W2BEG[5] ,
    \Tile_X5Y10_W2BEG[4] ,
    \Tile_X5Y10_W2BEG[3] ,
    \Tile_X5Y10_W2BEG[2] ,
    \Tile_X5Y10_W2BEG[1] ,
    \Tile_X5Y10_W2BEG[0] }),
    .W6BEG({\Tile_X4Y10_W6BEG[11] ,
    \Tile_X4Y10_W6BEG[10] ,
    \Tile_X4Y10_W6BEG[9] ,
    \Tile_X4Y10_W6BEG[8] ,
    \Tile_X4Y10_W6BEG[7] ,
    \Tile_X4Y10_W6BEG[6] ,
    \Tile_X4Y10_W6BEG[5] ,
    \Tile_X4Y10_W6BEG[4] ,
    \Tile_X4Y10_W6BEG[3] ,
    \Tile_X4Y10_W6BEG[2] ,
    \Tile_X4Y10_W6BEG[1] ,
    \Tile_X4Y10_W6BEG[0] }),
    .W6END({\Tile_X5Y10_W6BEG[11] ,
    \Tile_X5Y10_W6BEG[10] ,
    \Tile_X5Y10_W6BEG[9] ,
    \Tile_X5Y10_W6BEG[8] ,
    \Tile_X5Y10_W6BEG[7] ,
    \Tile_X5Y10_W6BEG[6] ,
    \Tile_X5Y10_W6BEG[5] ,
    \Tile_X5Y10_W6BEG[4] ,
    \Tile_X5Y10_W6BEG[3] ,
    \Tile_X5Y10_W6BEG[2] ,
    \Tile_X5Y10_W6BEG[1] ,
    \Tile_X5Y10_W6BEG[0] }),
    .WW4BEG({\Tile_X4Y10_WW4BEG[15] ,
    \Tile_X4Y10_WW4BEG[14] ,
    \Tile_X4Y10_WW4BEG[13] ,
    \Tile_X4Y10_WW4BEG[12] ,
    \Tile_X4Y10_WW4BEG[11] ,
    \Tile_X4Y10_WW4BEG[10] ,
    \Tile_X4Y10_WW4BEG[9] ,
    \Tile_X4Y10_WW4BEG[8] ,
    \Tile_X4Y10_WW4BEG[7] ,
    \Tile_X4Y10_WW4BEG[6] ,
    \Tile_X4Y10_WW4BEG[5] ,
    \Tile_X4Y10_WW4BEG[4] ,
    \Tile_X4Y10_WW4BEG[3] ,
    \Tile_X4Y10_WW4BEG[2] ,
    \Tile_X4Y10_WW4BEG[1] ,
    \Tile_X4Y10_WW4BEG[0] }),
    .WW4END({\Tile_X5Y10_WW4BEG[15] ,
    \Tile_X5Y10_WW4BEG[14] ,
    \Tile_X5Y10_WW4BEG[13] ,
    \Tile_X5Y10_WW4BEG[12] ,
    \Tile_X5Y10_WW4BEG[11] ,
    \Tile_X5Y10_WW4BEG[10] ,
    \Tile_X5Y10_WW4BEG[9] ,
    \Tile_X5Y10_WW4BEG[8] ,
    \Tile_X5Y10_WW4BEG[7] ,
    \Tile_X5Y10_WW4BEG[6] ,
    \Tile_X5Y10_WW4BEG[5] ,
    \Tile_X5Y10_WW4BEG[4] ,
    \Tile_X5Y10_WW4BEG[3] ,
    \Tile_X5Y10_WW4BEG[2] ,
    \Tile_X5Y10_WW4BEG[1] ,
    \Tile_X5Y10_WW4BEG[0] }));
 RegFile Tile_X4Y11_RegFile (.UserCLK(Tile_X4Y12_UserCLKo),
    .UserCLKo(Tile_X4Y11_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X4Y11_E1BEG[3] ,
    \Tile_X4Y11_E1BEG[2] ,
    \Tile_X4Y11_E1BEG[1] ,
    \Tile_X4Y11_E1BEG[0] }),
    .E1END({\Tile_X3Y11_E1BEG[3] ,
    \Tile_X3Y11_E1BEG[2] ,
    \Tile_X3Y11_E1BEG[1] ,
    \Tile_X3Y11_E1BEG[0] }),
    .E2BEG({\Tile_X4Y11_E2BEG[7] ,
    \Tile_X4Y11_E2BEG[6] ,
    \Tile_X4Y11_E2BEG[5] ,
    \Tile_X4Y11_E2BEG[4] ,
    \Tile_X4Y11_E2BEG[3] ,
    \Tile_X4Y11_E2BEG[2] ,
    \Tile_X4Y11_E2BEG[1] ,
    \Tile_X4Y11_E2BEG[0] }),
    .E2BEGb({\Tile_X4Y11_E2BEGb[7] ,
    \Tile_X4Y11_E2BEGb[6] ,
    \Tile_X4Y11_E2BEGb[5] ,
    \Tile_X4Y11_E2BEGb[4] ,
    \Tile_X4Y11_E2BEGb[3] ,
    \Tile_X4Y11_E2BEGb[2] ,
    \Tile_X4Y11_E2BEGb[1] ,
    \Tile_X4Y11_E2BEGb[0] }),
    .E2END({\Tile_X3Y11_E2BEGb[7] ,
    \Tile_X3Y11_E2BEGb[6] ,
    \Tile_X3Y11_E2BEGb[5] ,
    \Tile_X3Y11_E2BEGb[4] ,
    \Tile_X3Y11_E2BEGb[3] ,
    \Tile_X3Y11_E2BEGb[2] ,
    \Tile_X3Y11_E2BEGb[1] ,
    \Tile_X3Y11_E2BEGb[0] }),
    .E2MID({\Tile_X3Y11_E2BEG[7] ,
    \Tile_X3Y11_E2BEG[6] ,
    \Tile_X3Y11_E2BEG[5] ,
    \Tile_X3Y11_E2BEG[4] ,
    \Tile_X3Y11_E2BEG[3] ,
    \Tile_X3Y11_E2BEG[2] ,
    \Tile_X3Y11_E2BEG[1] ,
    \Tile_X3Y11_E2BEG[0] }),
    .E6BEG({\Tile_X4Y11_E6BEG[11] ,
    \Tile_X4Y11_E6BEG[10] ,
    \Tile_X4Y11_E6BEG[9] ,
    \Tile_X4Y11_E6BEG[8] ,
    \Tile_X4Y11_E6BEG[7] ,
    \Tile_X4Y11_E6BEG[6] ,
    \Tile_X4Y11_E6BEG[5] ,
    \Tile_X4Y11_E6BEG[4] ,
    \Tile_X4Y11_E6BEG[3] ,
    \Tile_X4Y11_E6BEG[2] ,
    \Tile_X4Y11_E6BEG[1] ,
    \Tile_X4Y11_E6BEG[0] }),
    .E6END({\Tile_X3Y11_E6BEG[11] ,
    \Tile_X3Y11_E6BEG[10] ,
    \Tile_X3Y11_E6BEG[9] ,
    \Tile_X3Y11_E6BEG[8] ,
    \Tile_X3Y11_E6BEG[7] ,
    \Tile_X3Y11_E6BEG[6] ,
    \Tile_X3Y11_E6BEG[5] ,
    \Tile_X3Y11_E6BEG[4] ,
    \Tile_X3Y11_E6BEG[3] ,
    \Tile_X3Y11_E6BEG[2] ,
    \Tile_X3Y11_E6BEG[1] ,
    \Tile_X3Y11_E6BEG[0] }),
    .EE4BEG({\Tile_X4Y11_EE4BEG[15] ,
    \Tile_X4Y11_EE4BEG[14] ,
    \Tile_X4Y11_EE4BEG[13] ,
    \Tile_X4Y11_EE4BEG[12] ,
    \Tile_X4Y11_EE4BEG[11] ,
    \Tile_X4Y11_EE4BEG[10] ,
    \Tile_X4Y11_EE4BEG[9] ,
    \Tile_X4Y11_EE4BEG[8] ,
    \Tile_X4Y11_EE4BEG[7] ,
    \Tile_X4Y11_EE4BEG[6] ,
    \Tile_X4Y11_EE4BEG[5] ,
    \Tile_X4Y11_EE4BEG[4] ,
    \Tile_X4Y11_EE4BEG[3] ,
    \Tile_X4Y11_EE4BEG[2] ,
    \Tile_X4Y11_EE4BEG[1] ,
    \Tile_X4Y11_EE4BEG[0] }),
    .EE4END({\Tile_X3Y11_EE4BEG[15] ,
    \Tile_X3Y11_EE4BEG[14] ,
    \Tile_X3Y11_EE4BEG[13] ,
    \Tile_X3Y11_EE4BEG[12] ,
    \Tile_X3Y11_EE4BEG[11] ,
    \Tile_X3Y11_EE4BEG[10] ,
    \Tile_X3Y11_EE4BEG[9] ,
    \Tile_X3Y11_EE4BEG[8] ,
    \Tile_X3Y11_EE4BEG[7] ,
    \Tile_X3Y11_EE4BEG[6] ,
    \Tile_X3Y11_EE4BEG[5] ,
    \Tile_X3Y11_EE4BEG[4] ,
    \Tile_X3Y11_EE4BEG[3] ,
    \Tile_X3Y11_EE4BEG[2] ,
    \Tile_X3Y11_EE4BEG[1] ,
    \Tile_X3Y11_EE4BEG[0] }),
    .FrameData({\Tile_X3Y11_FrameData_O[31] ,
    \Tile_X3Y11_FrameData_O[30] ,
    \Tile_X3Y11_FrameData_O[29] ,
    \Tile_X3Y11_FrameData_O[28] ,
    \Tile_X3Y11_FrameData_O[27] ,
    \Tile_X3Y11_FrameData_O[26] ,
    \Tile_X3Y11_FrameData_O[25] ,
    \Tile_X3Y11_FrameData_O[24] ,
    \Tile_X3Y11_FrameData_O[23] ,
    \Tile_X3Y11_FrameData_O[22] ,
    \Tile_X3Y11_FrameData_O[21] ,
    \Tile_X3Y11_FrameData_O[20] ,
    \Tile_X3Y11_FrameData_O[19] ,
    \Tile_X3Y11_FrameData_O[18] ,
    \Tile_X3Y11_FrameData_O[17] ,
    \Tile_X3Y11_FrameData_O[16] ,
    \Tile_X3Y11_FrameData_O[15] ,
    \Tile_X3Y11_FrameData_O[14] ,
    \Tile_X3Y11_FrameData_O[13] ,
    \Tile_X3Y11_FrameData_O[12] ,
    \Tile_X3Y11_FrameData_O[11] ,
    \Tile_X3Y11_FrameData_O[10] ,
    \Tile_X3Y11_FrameData_O[9] ,
    \Tile_X3Y11_FrameData_O[8] ,
    \Tile_X3Y11_FrameData_O[7] ,
    \Tile_X3Y11_FrameData_O[6] ,
    \Tile_X3Y11_FrameData_O[5] ,
    \Tile_X3Y11_FrameData_O[4] ,
    \Tile_X3Y11_FrameData_O[3] ,
    \Tile_X3Y11_FrameData_O[2] ,
    \Tile_X3Y11_FrameData_O[1] ,
    \Tile_X3Y11_FrameData_O[0] }),
    .FrameData_O({\Tile_X4Y11_FrameData_O[31] ,
    \Tile_X4Y11_FrameData_O[30] ,
    \Tile_X4Y11_FrameData_O[29] ,
    \Tile_X4Y11_FrameData_O[28] ,
    \Tile_X4Y11_FrameData_O[27] ,
    \Tile_X4Y11_FrameData_O[26] ,
    \Tile_X4Y11_FrameData_O[25] ,
    \Tile_X4Y11_FrameData_O[24] ,
    \Tile_X4Y11_FrameData_O[23] ,
    \Tile_X4Y11_FrameData_O[22] ,
    \Tile_X4Y11_FrameData_O[21] ,
    \Tile_X4Y11_FrameData_O[20] ,
    \Tile_X4Y11_FrameData_O[19] ,
    \Tile_X4Y11_FrameData_O[18] ,
    \Tile_X4Y11_FrameData_O[17] ,
    \Tile_X4Y11_FrameData_O[16] ,
    \Tile_X4Y11_FrameData_O[15] ,
    \Tile_X4Y11_FrameData_O[14] ,
    \Tile_X4Y11_FrameData_O[13] ,
    \Tile_X4Y11_FrameData_O[12] ,
    \Tile_X4Y11_FrameData_O[11] ,
    \Tile_X4Y11_FrameData_O[10] ,
    \Tile_X4Y11_FrameData_O[9] ,
    \Tile_X4Y11_FrameData_O[8] ,
    \Tile_X4Y11_FrameData_O[7] ,
    \Tile_X4Y11_FrameData_O[6] ,
    \Tile_X4Y11_FrameData_O[5] ,
    \Tile_X4Y11_FrameData_O[4] ,
    \Tile_X4Y11_FrameData_O[3] ,
    \Tile_X4Y11_FrameData_O[2] ,
    \Tile_X4Y11_FrameData_O[1] ,
    \Tile_X4Y11_FrameData_O[0] }),
    .FrameStrobe({\Tile_X4Y12_FrameStrobe_O[19] ,
    \Tile_X4Y12_FrameStrobe_O[18] ,
    \Tile_X4Y12_FrameStrobe_O[17] ,
    \Tile_X4Y12_FrameStrobe_O[16] ,
    \Tile_X4Y12_FrameStrobe_O[15] ,
    \Tile_X4Y12_FrameStrobe_O[14] ,
    \Tile_X4Y12_FrameStrobe_O[13] ,
    \Tile_X4Y12_FrameStrobe_O[12] ,
    \Tile_X4Y12_FrameStrobe_O[11] ,
    \Tile_X4Y12_FrameStrobe_O[10] ,
    \Tile_X4Y12_FrameStrobe_O[9] ,
    \Tile_X4Y12_FrameStrobe_O[8] ,
    \Tile_X4Y12_FrameStrobe_O[7] ,
    \Tile_X4Y12_FrameStrobe_O[6] ,
    \Tile_X4Y12_FrameStrobe_O[5] ,
    \Tile_X4Y12_FrameStrobe_O[4] ,
    \Tile_X4Y12_FrameStrobe_O[3] ,
    \Tile_X4Y12_FrameStrobe_O[2] ,
    \Tile_X4Y12_FrameStrobe_O[1] ,
    \Tile_X4Y12_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X4Y11_FrameStrobe_O[19] ,
    \Tile_X4Y11_FrameStrobe_O[18] ,
    \Tile_X4Y11_FrameStrobe_O[17] ,
    \Tile_X4Y11_FrameStrobe_O[16] ,
    \Tile_X4Y11_FrameStrobe_O[15] ,
    \Tile_X4Y11_FrameStrobe_O[14] ,
    \Tile_X4Y11_FrameStrobe_O[13] ,
    \Tile_X4Y11_FrameStrobe_O[12] ,
    \Tile_X4Y11_FrameStrobe_O[11] ,
    \Tile_X4Y11_FrameStrobe_O[10] ,
    \Tile_X4Y11_FrameStrobe_O[9] ,
    \Tile_X4Y11_FrameStrobe_O[8] ,
    \Tile_X4Y11_FrameStrobe_O[7] ,
    \Tile_X4Y11_FrameStrobe_O[6] ,
    \Tile_X4Y11_FrameStrobe_O[5] ,
    \Tile_X4Y11_FrameStrobe_O[4] ,
    \Tile_X4Y11_FrameStrobe_O[3] ,
    \Tile_X4Y11_FrameStrobe_O[2] ,
    \Tile_X4Y11_FrameStrobe_O[1] ,
    \Tile_X4Y11_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X4Y11_N1BEG[3] ,
    \Tile_X4Y11_N1BEG[2] ,
    \Tile_X4Y11_N1BEG[1] ,
    \Tile_X4Y11_N1BEG[0] }),
    .N1END({\Tile_X4Y12_N1BEG[3] ,
    \Tile_X4Y12_N1BEG[2] ,
    \Tile_X4Y12_N1BEG[1] ,
    \Tile_X4Y12_N1BEG[0] }),
    .N2BEG({\Tile_X4Y11_N2BEG[7] ,
    \Tile_X4Y11_N2BEG[6] ,
    \Tile_X4Y11_N2BEG[5] ,
    \Tile_X4Y11_N2BEG[4] ,
    \Tile_X4Y11_N2BEG[3] ,
    \Tile_X4Y11_N2BEG[2] ,
    \Tile_X4Y11_N2BEG[1] ,
    \Tile_X4Y11_N2BEG[0] }),
    .N2BEGb({\Tile_X4Y11_N2BEGb[7] ,
    \Tile_X4Y11_N2BEGb[6] ,
    \Tile_X4Y11_N2BEGb[5] ,
    \Tile_X4Y11_N2BEGb[4] ,
    \Tile_X4Y11_N2BEGb[3] ,
    \Tile_X4Y11_N2BEGb[2] ,
    \Tile_X4Y11_N2BEGb[1] ,
    \Tile_X4Y11_N2BEGb[0] }),
    .N2END({\Tile_X4Y12_N2BEGb[7] ,
    \Tile_X4Y12_N2BEGb[6] ,
    \Tile_X4Y12_N2BEGb[5] ,
    \Tile_X4Y12_N2BEGb[4] ,
    \Tile_X4Y12_N2BEGb[3] ,
    \Tile_X4Y12_N2BEGb[2] ,
    \Tile_X4Y12_N2BEGb[1] ,
    \Tile_X4Y12_N2BEGb[0] }),
    .N2MID({\Tile_X4Y12_N2BEG[7] ,
    \Tile_X4Y12_N2BEG[6] ,
    \Tile_X4Y12_N2BEG[5] ,
    \Tile_X4Y12_N2BEG[4] ,
    \Tile_X4Y12_N2BEG[3] ,
    \Tile_X4Y12_N2BEG[2] ,
    \Tile_X4Y12_N2BEG[1] ,
    \Tile_X4Y12_N2BEG[0] }),
    .N4BEG({\Tile_X4Y11_N4BEG[15] ,
    \Tile_X4Y11_N4BEG[14] ,
    \Tile_X4Y11_N4BEG[13] ,
    \Tile_X4Y11_N4BEG[12] ,
    \Tile_X4Y11_N4BEG[11] ,
    \Tile_X4Y11_N4BEG[10] ,
    \Tile_X4Y11_N4BEG[9] ,
    \Tile_X4Y11_N4BEG[8] ,
    \Tile_X4Y11_N4BEG[7] ,
    \Tile_X4Y11_N4BEG[6] ,
    \Tile_X4Y11_N4BEG[5] ,
    \Tile_X4Y11_N4BEG[4] ,
    \Tile_X4Y11_N4BEG[3] ,
    \Tile_X4Y11_N4BEG[2] ,
    \Tile_X4Y11_N4BEG[1] ,
    \Tile_X4Y11_N4BEG[0] }),
    .N4END({\Tile_X4Y12_N4BEG[15] ,
    \Tile_X4Y12_N4BEG[14] ,
    \Tile_X4Y12_N4BEG[13] ,
    \Tile_X4Y12_N4BEG[12] ,
    \Tile_X4Y12_N4BEG[11] ,
    \Tile_X4Y12_N4BEG[10] ,
    \Tile_X4Y12_N4BEG[9] ,
    \Tile_X4Y12_N4BEG[8] ,
    \Tile_X4Y12_N4BEG[7] ,
    \Tile_X4Y12_N4BEG[6] ,
    \Tile_X4Y12_N4BEG[5] ,
    \Tile_X4Y12_N4BEG[4] ,
    \Tile_X4Y12_N4BEG[3] ,
    \Tile_X4Y12_N4BEG[2] ,
    \Tile_X4Y12_N4BEG[1] ,
    \Tile_X4Y12_N4BEG[0] }),
    .NN4BEG({\Tile_X4Y11_NN4BEG[15] ,
    \Tile_X4Y11_NN4BEG[14] ,
    \Tile_X4Y11_NN4BEG[13] ,
    \Tile_X4Y11_NN4BEG[12] ,
    \Tile_X4Y11_NN4BEG[11] ,
    \Tile_X4Y11_NN4BEG[10] ,
    \Tile_X4Y11_NN4BEG[9] ,
    \Tile_X4Y11_NN4BEG[8] ,
    \Tile_X4Y11_NN4BEG[7] ,
    \Tile_X4Y11_NN4BEG[6] ,
    \Tile_X4Y11_NN4BEG[5] ,
    \Tile_X4Y11_NN4BEG[4] ,
    \Tile_X4Y11_NN4BEG[3] ,
    \Tile_X4Y11_NN4BEG[2] ,
    \Tile_X4Y11_NN4BEG[1] ,
    \Tile_X4Y11_NN4BEG[0] }),
    .NN4END({\Tile_X4Y12_NN4BEG[15] ,
    \Tile_X4Y12_NN4BEG[14] ,
    \Tile_X4Y12_NN4BEG[13] ,
    \Tile_X4Y12_NN4BEG[12] ,
    \Tile_X4Y12_NN4BEG[11] ,
    \Tile_X4Y12_NN4BEG[10] ,
    \Tile_X4Y12_NN4BEG[9] ,
    \Tile_X4Y12_NN4BEG[8] ,
    \Tile_X4Y12_NN4BEG[7] ,
    \Tile_X4Y12_NN4BEG[6] ,
    \Tile_X4Y12_NN4BEG[5] ,
    \Tile_X4Y12_NN4BEG[4] ,
    \Tile_X4Y12_NN4BEG[3] ,
    \Tile_X4Y12_NN4BEG[2] ,
    \Tile_X4Y12_NN4BEG[1] ,
    \Tile_X4Y12_NN4BEG[0] }),
    .S1BEG({\Tile_X4Y11_S1BEG[3] ,
    \Tile_X4Y11_S1BEG[2] ,
    \Tile_X4Y11_S1BEG[1] ,
    \Tile_X4Y11_S1BEG[0] }),
    .S1END({\Tile_X4Y10_S1BEG[3] ,
    \Tile_X4Y10_S1BEG[2] ,
    \Tile_X4Y10_S1BEG[1] ,
    \Tile_X4Y10_S1BEG[0] }),
    .S2BEG({\Tile_X4Y11_S2BEG[7] ,
    \Tile_X4Y11_S2BEG[6] ,
    \Tile_X4Y11_S2BEG[5] ,
    \Tile_X4Y11_S2BEG[4] ,
    \Tile_X4Y11_S2BEG[3] ,
    \Tile_X4Y11_S2BEG[2] ,
    \Tile_X4Y11_S2BEG[1] ,
    \Tile_X4Y11_S2BEG[0] }),
    .S2BEGb({\Tile_X4Y11_S2BEGb[7] ,
    \Tile_X4Y11_S2BEGb[6] ,
    \Tile_X4Y11_S2BEGb[5] ,
    \Tile_X4Y11_S2BEGb[4] ,
    \Tile_X4Y11_S2BEGb[3] ,
    \Tile_X4Y11_S2BEGb[2] ,
    \Tile_X4Y11_S2BEGb[1] ,
    \Tile_X4Y11_S2BEGb[0] }),
    .S2END({\Tile_X4Y10_S2BEGb[7] ,
    \Tile_X4Y10_S2BEGb[6] ,
    \Tile_X4Y10_S2BEGb[5] ,
    \Tile_X4Y10_S2BEGb[4] ,
    \Tile_X4Y10_S2BEGb[3] ,
    \Tile_X4Y10_S2BEGb[2] ,
    \Tile_X4Y10_S2BEGb[1] ,
    \Tile_X4Y10_S2BEGb[0] }),
    .S2MID({\Tile_X4Y10_S2BEG[7] ,
    \Tile_X4Y10_S2BEG[6] ,
    \Tile_X4Y10_S2BEG[5] ,
    \Tile_X4Y10_S2BEG[4] ,
    \Tile_X4Y10_S2BEG[3] ,
    \Tile_X4Y10_S2BEG[2] ,
    \Tile_X4Y10_S2BEG[1] ,
    \Tile_X4Y10_S2BEG[0] }),
    .S4BEG({\Tile_X4Y11_S4BEG[15] ,
    \Tile_X4Y11_S4BEG[14] ,
    \Tile_X4Y11_S4BEG[13] ,
    \Tile_X4Y11_S4BEG[12] ,
    \Tile_X4Y11_S4BEG[11] ,
    \Tile_X4Y11_S4BEG[10] ,
    \Tile_X4Y11_S4BEG[9] ,
    \Tile_X4Y11_S4BEG[8] ,
    \Tile_X4Y11_S4BEG[7] ,
    \Tile_X4Y11_S4BEG[6] ,
    \Tile_X4Y11_S4BEG[5] ,
    \Tile_X4Y11_S4BEG[4] ,
    \Tile_X4Y11_S4BEG[3] ,
    \Tile_X4Y11_S4BEG[2] ,
    \Tile_X4Y11_S4BEG[1] ,
    \Tile_X4Y11_S4BEG[0] }),
    .S4END({\Tile_X4Y10_S4BEG[15] ,
    \Tile_X4Y10_S4BEG[14] ,
    \Tile_X4Y10_S4BEG[13] ,
    \Tile_X4Y10_S4BEG[12] ,
    \Tile_X4Y10_S4BEG[11] ,
    \Tile_X4Y10_S4BEG[10] ,
    \Tile_X4Y10_S4BEG[9] ,
    \Tile_X4Y10_S4BEG[8] ,
    \Tile_X4Y10_S4BEG[7] ,
    \Tile_X4Y10_S4BEG[6] ,
    \Tile_X4Y10_S4BEG[5] ,
    \Tile_X4Y10_S4BEG[4] ,
    \Tile_X4Y10_S4BEG[3] ,
    \Tile_X4Y10_S4BEG[2] ,
    \Tile_X4Y10_S4BEG[1] ,
    \Tile_X4Y10_S4BEG[0] }),
    .SS4BEG({\Tile_X4Y11_SS4BEG[15] ,
    \Tile_X4Y11_SS4BEG[14] ,
    \Tile_X4Y11_SS4BEG[13] ,
    \Tile_X4Y11_SS4BEG[12] ,
    \Tile_X4Y11_SS4BEG[11] ,
    \Tile_X4Y11_SS4BEG[10] ,
    \Tile_X4Y11_SS4BEG[9] ,
    \Tile_X4Y11_SS4BEG[8] ,
    \Tile_X4Y11_SS4BEG[7] ,
    \Tile_X4Y11_SS4BEG[6] ,
    \Tile_X4Y11_SS4BEG[5] ,
    \Tile_X4Y11_SS4BEG[4] ,
    \Tile_X4Y11_SS4BEG[3] ,
    \Tile_X4Y11_SS4BEG[2] ,
    \Tile_X4Y11_SS4BEG[1] ,
    \Tile_X4Y11_SS4BEG[0] }),
    .SS4END({\Tile_X4Y10_SS4BEG[15] ,
    \Tile_X4Y10_SS4BEG[14] ,
    \Tile_X4Y10_SS4BEG[13] ,
    \Tile_X4Y10_SS4BEG[12] ,
    \Tile_X4Y10_SS4BEG[11] ,
    \Tile_X4Y10_SS4BEG[10] ,
    \Tile_X4Y10_SS4BEG[9] ,
    \Tile_X4Y10_SS4BEG[8] ,
    \Tile_X4Y10_SS4BEG[7] ,
    \Tile_X4Y10_SS4BEG[6] ,
    \Tile_X4Y10_SS4BEG[5] ,
    \Tile_X4Y10_SS4BEG[4] ,
    \Tile_X4Y10_SS4BEG[3] ,
    \Tile_X4Y10_SS4BEG[2] ,
    \Tile_X4Y10_SS4BEG[1] ,
    \Tile_X4Y10_SS4BEG[0] }),
    .W1BEG({\Tile_X4Y11_W1BEG[3] ,
    \Tile_X4Y11_W1BEG[2] ,
    \Tile_X4Y11_W1BEG[1] ,
    \Tile_X4Y11_W1BEG[0] }),
    .W1END({\Tile_X5Y11_W1BEG[3] ,
    \Tile_X5Y11_W1BEG[2] ,
    \Tile_X5Y11_W1BEG[1] ,
    \Tile_X5Y11_W1BEG[0] }),
    .W2BEG({\Tile_X4Y11_W2BEG[7] ,
    \Tile_X4Y11_W2BEG[6] ,
    \Tile_X4Y11_W2BEG[5] ,
    \Tile_X4Y11_W2BEG[4] ,
    \Tile_X4Y11_W2BEG[3] ,
    \Tile_X4Y11_W2BEG[2] ,
    \Tile_X4Y11_W2BEG[1] ,
    \Tile_X4Y11_W2BEG[0] }),
    .W2BEGb({\Tile_X4Y11_W2BEGb[7] ,
    \Tile_X4Y11_W2BEGb[6] ,
    \Tile_X4Y11_W2BEGb[5] ,
    \Tile_X4Y11_W2BEGb[4] ,
    \Tile_X4Y11_W2BEGb[3] ,
    \Tile_X4Y11_W2BEGb[2] ,
    \Tile_X4Y11_W2BEGb[1] ,
    \Tile_X4Y11_W2BEGb[0] }),
    .W2END({\Tile_X5Y11_W2BEGb[7] ,
    \Tile_X5Y11_W2BEGb[6] ,
    \Tile_X5Y11_W2BEGb[5] ,
    \Tile_X5Y11_W2BEGb[4] ,
    \Tile_X5Y11_W2BEGb[3] ,
    \Tile_X5Y11_W2BEGb[2] ,
    \Tile_X5Y11_W2BEGb[1] ,
    \Tile_X5Y11_W2BEGb[0] }),
    .W2MID({\Tile_X5Y11_W2BEG[7] ,
    \Tile_X5Y11_W2BEG[6] ,
    \Tile_X5Y11_W2BEG[5] ,
    \Tile_X5Y11_W2BEG[4] ,
    \Tile_X5Y11_W2BEG[3] ,
    \Tile_X5Y11_W2BEG[2] ,
    \Tile_X5Y11_W2BEG[1] ,
    \Tile_X5Y11_W2BEG[0] }),
    .W6BEG({\Tile_X4Y11_W6BEG[11] ,
    \Tile_X4Y11_W6BEG[10] ,
    \Tile_X4Y11_W6BEG[9] ,
    \Tile_X4Y11_W6BEG[8] ,
    \Tile_X4Y11_W6BEG[7] ,
    \Tile_X4Y11_W6BEG[6] ,
    \Tile_X4Y11_W6BEG[5] ,
    \Tile_X4Y11_W6BEG[4] ,
    \Tile_X4Y11_W6BEG[3] ,
    \Tile_X4Y11_W6BEG[2] ,
    \Tile_X4Y11_W6BEG[1] ,
    \Tile_X4Y11_W6BEG[0] }),
    .W6END({\Tile_X5Y11_W6BEG[11] ,
    \Tile_X5Y11_W6BEG[10] ,
    \Tile_X5Y11_W6BEG[9] ,
    \Tile_X5Y11_W6BEG[8] ,
    \Tile_X5Y11_W6BEG[7] ,
    \Tile_X5Y11_W6BEG[6] ,
    \Tile_X5Y11_W6BEG[5] ,
    \Tile_X5Y11_W6BEG[4] ,
    \Tile_X5Y11_W6BEG[3] ,
    \Tile_X5Y11_W6BEG[2] ,
    \Tile_X5Y11_W6BEG[1] ,
    \Tile_X5Y11_W6BEG[0] }),
    .WW4BEG({\Tile_X4Y11_WW4BEG[15] ,
    \Tile_X4Y11_WW4BEG[14] ,
    \Tile_X4Y11_WW4BEG[13] ,
    \Tile_X4Y11_WW4BEG[12] ,
    \Tile_X4Y11_WW4BEG[11] ,
    \Tile_X4Y11_WW4BEG[10] ,
    \Tile_X4Y11_WW4BEG[9] ,
    \Tile_X4Y11_WW4BEG[8] ,
    \Tile_X4Y11_WW4BEG[7] ,
    \Tile_X4Y11_WW4BEG[6] ,
    \Tile_X4Y11_WW4BEG[5] ,
    \Tile_X4Y11_WW4BEG[4] ,
    \Tile_X4Y11_WW4BEG[3] ,
    \Tile_X4Y11_WW4BEG[2] ,
    \Tile_X4Y11_WW4BEG[1] ,
    \Tile_X4Y11_WW4BEG[0] }),
    .WW4END({\Tile_X5Y11_WW4BEG[15] ,
    \Tile_X5Y11_WW4BEG[14] ,
    \Tile_X5Y11_WW4BEG[13] ,
    \Tile_X5Y11_WW4BEG[12] ,
    \Tile_X5Y11_WW4BEG[11] ,
    \Tile_X5Y11_WW4BEG[10] ,
    \Tile_X5Y11_WW4BEG[9] ,
    \Tile_X5Y11_WW4BEG[8] ,
    \Tile_X5Y11_WW4BEG[7] ,
    \Tile_X5Y11_WW4BEG[6] ,
    \Tile_X5Y11_WW4BEG[5] ,
    \Tile_X5Y11_WW4BEG[4] ,
    \Tile_X5Y11_WW4BEG[3] ,
    \Tile_X5Y11_WW4BEG[2] ,
    \Tile_X5Y11_WW4BEG[1] ,
    \Tile_X5Y11_WW4BEG[0] }));
 RegFile Tile_X4Y12_RegFile (.UserCLK(Tile_X4Y13_UserCLKo),
    .UserCLKo(Tile_X4Y12_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X4Y12_E1BEG[3] ,
    \Tile_X4Y12_E1BEG[2] ,
    \Tile_X4Y12_E1BEG[1] ,
    \Tile_X4Y12_E1BEG[0] }),
    .E1END({\Tile_X3Y12_E1BEG[3] ,
    \Tile_X3Y12_E1BEG[2] ,
    \Tile_X3Y12_E1BEG[1] ,
    \Tile_X3Y12_E1BEG[0] }),
    .E2BEG({\Tile_X4Y12_E2BEG[7] ,
    \Tile_X4Y12_E2BEG[6] ,
    \Tile_X4Y12_E2BEG[5] ,
    \Tile_X4Y12_E2BEG[4] ,
    \Tile_X4Y12_E2BEG[3] ,
    \Tile_X4Y12_E2BEG[2] ,
    \Tile_X4Y12_E2BEG[1] ,
    \Tile_X4Y12_E2BEG[0] }),
    .E2BEGb({\Tile_X4Y12_E2BEGb[7] ,
    \Tile_X4Y12_E2BEGb[6] ,
    \Tile_X4Y12_E2BEGb[5] ,
    \Tile_X4Y12_E2BEGb[4] ,
    \Tile_X4Y12_E2BEGb[3] ,
    \Tile_X4Y12_E2BEGb[2] ,
    \Tile_X4Y12_E2BEGb[1] ,
    \Tile_X4Y12_E2BEGb[0] }),
    .E2END({\Tile_X3Y12_E2BEGb[7] ,
    \Tile_X3Y12_E2BEGb[6] ,
    \Tile_X3Y12_E2BEGb[5] ,
    \Tile_X3Y12_E2BEGb[4] ,
    \Tile_X3Y12_E2BEGb[3] ,
    \Tile_X3Y12_E2BEGb[2] ,
    \Tile_X3Y12_E2BEGb[1] ,
    \Tile_X3Y12_E2BEGb[0] }),
    .E2MID({\Tile_X3Y12_E2BEG[7] ,
    \Tile_X3Y12_E2BEG[6] ,
    \Tile_X3Y12_E2BEG[5] ,
    \Tile_X3Y12_E2BEG[4] ,
    \Tile_X3Y12_E2BEG[3] ,
    \Tile_X3Y12_E2BEG[2] ,
    \Tile_X3Y12_E2BEG[1] ,
    \Tile_X3Y12_E2BEG[0] }),
    .E6BEG({\Tile_X4Y12_E6BEG[11] ,
    \Tile_X4Y12_E6BEG[10] ,
    \Tile_X4Y12_E6BEG[9] ,
    \Tile_X4Y12_E6BEG[8] ,
    \Tile_X4Y12_E6BEG[7] ,
    \Tile_X4Y12_E6BEG[6] ,
    \Tile_X4Y12_E6BEG[5] ,
    \Tile_X4Y12_E6BEG[4] ,
    \Tile_X4Y12_E6BEG[3] ,
    \Tile_X4Y12_E6BEG[2] ,
    \Tile_X4Y12_E6BEG[1] ,
    \Tile_X4Y12_E6BEG[0] }),
    .E6END({\Tile_X3Y12_E6BEG[11] ,
    \Tile_X3Y12_E6BEG[10] ,
    \Tile_X3Y12_E6BEG[9] ,
    \Tile_X3Y12_E6BEG[8] ,
    \Tile_X3Y12_E6BEG[7] ,
    \Tile_X3Y12_E6BEG[6] ,
    \Tile_X3Y12_E6BEG[5] ,
    \Tile_X3Y12_E6BEG[4] ,
    \Tile_X3Y12_E6BEG[3] ,
    \Tile_X3Y12_E6BEG[2] ,
    \Tile_X3Y12_E6BEG[1] ,
    \Tile_X3Y12_E6BEG[0] }),
    .EE4BEG({\Tile_X4Y12_EE4BEG[15] ,
    \Tile_X4Y12_EE4BEG[14] ,
    \Tile_X4Y12_EE4BEG[13] ,
    \Tile_X4Y12_EE4BEG[12] ,
    \Tile_X4Y12_EE4BEG[11] ,
    \Tile_X4Y12_EE4BEG[10] ,
    \Tile_X4Y12_EE4BEG[9] ,
    \Tile_X4Y12_EE4BEG[8] ,
    \Tile_X4Y12_EE4BEG[7] ,
    \Tile_X4Y12_EE4BEG[6] ,
    \Tile_X4Y12_EE4BEG[5] ,
    \Tile_X4Y12_EE4BEG[4] ,
    \Tile_X4Y12_EE4BEG[3] ,
    \Tile_X4Y12_EE4BEG[2] ,
    \Tile_X4Y12_EE4BEG[1] ,
    \Tile_X4Y12_EE4BEG[0] }),
    .EE4END({\Tile_X3Y12_EE4BEG[15] ,
    \Tile_X3Y12_EE4BEG[14] ,
    \Tile_X3Y12_EE4BEG[13] ,
    \Tile_X3Y12_EE4BEG[12] ,
    \Tile_X3Y12_EE4BEG[11] ,
    \Tile_X3Y12_EE4BEG[10] ,
    \Tile_X3Y12_EE4BEG[9] ,
    \Tile_X3Y12_EE4BEG[8] ,
    \Tile_X3Y12_EE4BEG[7] ,
    \Tile_X3Y12_EE4BEG[6] ,
    \Tile_X3Y12_EE4BEG[5] ,
    \Tile_X3Y12_EE4BEG[4] ,
    \Tile_X3Y12_EE4BEG[3] ,
    \Tile_X3Y12_EE4BEG[2] ,
    \Tile_X3Y12_EE4BEG[1] ,
    \Tile_X3Y12_EE4BEG[0] }),
    .FrameData({\Tile_X3Y12_FrameData_O[31] ,
    \Tile_X3Y12_FrameData_O[30] ,
    \Tile_X3Y12_FrameData_O[29] ,
    \Tile_X3Y12_FrameData_O[28] ,
    \Tile_X3Y12_FrameData_O[27] ,
    \Tile_X3Y12_FrameData_O[26] ,
    \Tile_X3Y12_FrameData_O[25] ,
    \Tile_X3Y12_FrameData_O[24] ,
    \Tile_X3Y12_FrameData_O[23] ,
    \Tile_X3Y12_FrameData_O[22] ,
    \Tile_X3Y12_FrameData_O[21] ,
    \Tile_X3Y12_FrameData_O[20] ,
    \Tile_X3Y12_FrameData_O[19] ,
    \Tile_X3Y12_FrameData_O[18] ,
    \Tile_X3Y12_FrameData_O[17] ,
    \Tile_X3Y12_FrameData_O[16] ,
    \Tile_X3Y12_FrameData_O[15] ,
    \Tile_X3Y12_FrameData_O[14] ,
    \Tile_X3Y12_FrameData_O[13] ,
    \Tile_X3Y12_FrameData_O[12] ,
    \Tile_X3Y12_FrameData_O[11] ,
    \Tile_X3Y12_FrameData_O[10] ,
    \Tile_X3Y12_FrameData_O[9] ,
    \Tile_X3Y12_FrameData_O[8] ,
    \Tile_X3Y12_FrameData_O[7] ,
    \Tile_X3Y12_FrameData_O[6] ,
    \Tile_X3Y12_FrameData_O[5] ,
    \Tile_X3Y12_FrameData_O[4] ,
    \Tile_X3Y12_FrameData_O[3] ,
    \Tile_X3Y12_FrameData_O[2] ,
    \Tile_X3Y12_FrameData_O[1] ,
    \Tile_X3Y12_FrameData_O[0] }),
    .FrameData_O({\Tile_X4Y12_FrameData_O[31] ,
    \Tile_X4Y12_FrameData_O[30] ,
    \Tile_X4Y12_FrameData_O[29] ,
    \Tile_X4Y12_FrameData_O[28] ,
    \Tile_X4Y12_FrameData_O[27] ,
    \Tile_X4Y12_FrameData_O[26] ,
    \Tile_X4Y12_FrameData_O[25] ,
    \Tile_X4Y12_FrameData_O[24] ,
    \Tile_X4Y12_FrameData_O[23] ,
    \Tile_X4Y12_FrameData_O[22] ,
    \Tile_X4Y12_FrameData_O[21] ,
    \Tile_X4Y12_FrameData_O[20] ,
    \Tile_X4Y12_FrameData_O[19] ,
    \Tile_X4Y12_FrameData_O[18] ,
    \Tile_X4Y12_FrameData_O[17] ,
    \Tile_X4Y12_FrameData_O[16] ,
    \Tile_X4Y12_FrameData_O[15] ,
    \Tile_X4Y12_FrameData_O[14] ,
    \Tile_X4Y12_FrameData_O[13] ,
    \Tile_X4Y12_FrameData_O[12] ,
    \Tile_X4Y12_FrameData_O[11] ,
    \Tile_X4Y12_FrameData_O[10] ,
    \Tile_X4Y12_FrameData_O[9] ,
    \Tile_X4Y12_FrameData_O[8] ,
    \Tile_X4Y12_FrameData_O[7] ,
    \Tile_X4Y12_FrameData_O[6] ,
    \Tile_X4Y12_FrameData_O[5] ,
    \Tile_X4Y12_FrameData_O[4] ,
    \Tile_X4Y12_FrameData_O[3] ,
    \Tile_X4Y12_FrameData_O[2] ,
    \Tile_X4Y12_FrameData_O[1] ,
    \Tile_X4Y12_FrameData_O[0] }),
    .FrameStrobe({\Tile_X4Y13_FrameStrobe_O[19] ,
    \Tile_X4Y13_FrameStrobe_O[18] ,
    \Tile_X4Y13_FrameStrobe_O[17] ,
    \Tile_X4Y13_FrameStrobe_O[16] ,
    \Tile_X4Y13_FrameStrobe_O[15] ,
    \Tile_X4Y13_FrameStrobe_O[14] ,
    \Tile_X4Y13_FrameStrobe_O[13] ,
    \Tile_X4Y13_FrameStrobe_O[12] ,
    \Tile_X4Y13_FrameStrobe_O[11] ,
    \Tile_X4Y13_FrameStrobe_O[10] ,
    \Tile_X4Y13_FrameStrobe_O[9] ,
    \Tile_X4Y13_FrameStrobe_O[8] ,
    \Tile_X4Y13_FrameStrobe_O[7] ,
    \Tile_X4Y13_FrameStrobe_O[6] ,
    \Tile_X4Y13_FrameStrobe_O[5] ,
    \Tile_X4Y13_FrameStrobe_O[4] ,
    \Tile_X4Y13_FrameStrobe_O[3] ,
    \Tile_X4Y13_FrameStrobe_O[2] ,
    \Tile_X4Y13_FrameStrobe_O[1] ,
    \Tile_X4Y13_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X4Y12_FrameStrobe_O[19] ,
    \Tile_X4Y12_FrameStrobe_O[18] ,
    \Tile_X4Y12_FrameStrobe_O[17] ,
    \Tile_X4Y12_FrameStrobe_O[16] ,
    \Tile_X4Y12_FrameStrobe_O[15] ,
    \Tile_X4Y12_FrameStrobe_O[14] ,
    \Tile_X4Y12_FrameStrobe_O[13] ,
    \Tile_X4Y12_FrameStrobe_O[12] ,
    \Tile_X4Y12_FrameStrobe_O[11] ,
    \Tile_X4Y12_FrameStrobe_O[10] ,
    \Tile_X4Y12_FrameStrobe_O[9] ,
    \Tile_X4Y12_FrameStrobe_O[8] ,
    \Tile_X4Y12_FrameStrobe_O[7] ,
    \Tile_X4Y12_FrameStrobe_O[6] ,
    \Tile_X4Y12_FrameStrobe_O[5] ,
    \Tile_X4Y12_FrameStrobe_O[4] ,
    \Tile_X4Y12_FrameStrobe_O[3] ,
    \Tile_X4Y12_FrameStrobe_O[2] ,
    \Tile_X4Y12_FrameStrobe_O[1] ,
    \Tile_X4Y12_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X4Y12_N1BEG[3] ,
    \Tile_X4Y12_N1BEG[2] ,
    \Tile_X4Y12_N1BEG[1] ,
    \Tile_X4Y12_N1BEG[0] }),
    .N1END({\Tile_X4Y13_N1BEG[3] ,
    \Tile_X4Y13_N1BEG[2] ,
    \Tile_X4Y13_N1BEG[1] ,
    \Tile_X4Y13_N1BEG[0] }),
    .N2BEG({\Tile_X4Y12_N2BEG[7] ,
    \Tile_X4Y12_N2BEG[6] ,
    \Tile_X4Y12_N2BEG[5] ,
    \Tile_X4Y12_N2BEG[4] ,
    \Tile_X4Y12_N2BEG[3] ,
    \Tile_X4Y12_N2BEG[2] ,
    \Tile_X4Y12_N2BEG[1] ,
    \Tile_X4Y12_N2BEG[0] }),
    .N2BEGb({\Tile_X4Y12_N2BEGb[7] ,
    \Tile_X4Y12_N2BEGb[6] ,
    \Tile_X4Y12_N2BEGb[5] ,
    \Tile_X4Y12_N2BEGb[4] ,
    \Tile_X4Y12_N2BEGb[3] ,
    \Tile_X4Y12_N2BEGb[2] ,
    \Tile_X4Y12_N2BEGb[1] ,
    \Tile_X4Y12_N2BEGb[0] }),
    .N2END({\Tile_X4Y13_N2BEGb[7] ,
    \Tile_X4Y13_N2BEGb[6] ,
    \Tile_X4Y13_N2BEGb[5] ,
    \Tile_X4Y13_N2BEGb[4] ,
    \Tile_X4Y13_N2BEGb[3] ,
    \Tile_X4Y13_N2BEGb[2] ,
    \Tile_X4Y13_N2BEGb[1] ,
    \Tile_X4Y13_N2BEGb[0] }),
    .N2MID({\Tile_X4Y13_N2BEG[7] ,
    \Tile_X4Y13_N2BEG[6] ,
    \Tile_X4Y13_N2BEG[5] ,
    \Tile_X4Y13_N2BEG[4] ,
    \Tile_X4Y13_N2BEG[3] ,
    \Tile_X4Y13_N2BEG[2] ,
    \Tile_X4Y13_N2BEG[1] ,
    \Tile_X4Y13_N2BEG[0] }),
    .N4BEG({\Tile_X4Y12_N4BEG[15] ,
    \Tile_X4Y12_N4BEG[14] ,
    \Tile_X4Y12_N4BEG[13] ,
    \Tile_X4Y12_N4BEG[12] ,
    \Tile_X4Y12_N4BEG[11] ,
    \Tile_X4Y12_N4BEG[10] ,
    \Tile_X4Y12_N4BEG[9] ,
    \Tile_X4Y12_N4BEG[8] ,
    \Tile_X4Y12_N4BEG[7] ,
    \Tile_X4Y12_N4BEG[6] ,
    \Tile_X4Y12_N4BEG[5] ,
    \Tile_X4Y12_N4BEG[4] ,
    \Tile_X4Y12_N4BEG[3] ,
    \Tile_X4Y12_N4BEG[2] ,
    \Tile_X4Y12_N4BEG[1] ,
    \Tile_X4Y12_N4BEG[0] }),
    .N4END({\Tile_X4Y13_N4BEG[15] ,
    \Tile_X4Y13_N4BEG[14] ,
    \Tile_X4Y13_N4BEG[13] ,
    \Tile_X4Y13_N4BEG[12] ,
    \Tile_X4Y13_N4BEG[11] ,
    \Tile_X4Y13_N4BEG[10] ,
    \Tile_X4Y13_N4BEG[9] ,
    \Tile_X4Y13_N4BEG[8] ,
    \Tile_X4Y13_N4BEG[7] ,
    \Tile_X4Y13_N4BEG[6] ,
    \Tile_X4Y13_N4BEG[5] ,
    \Tile_X4Y13_N4BEG[4] ,
    \Tile_X4Y13_N4BEG[3] ,
    \Tile_X4Y13_N4BEG[2] ,
    \Tile_X4Y13_N4BEG[1] ,
    \Tile_X4Y13_N4BEG[0] }),
    .NN4BEG({\Tile_X4Y12_NN4BEG[15] ,
    \Tile_X4Y12_NN4BEG[14] ,
    \Tile_X4Y12_NN4BEG[13] ,
    \Tile_X4Y12_NN4BEG[12] ,
    \Tile_X4Y12_NN4BEG[11] ,
    \Tile_X4Y12_NN4BEG[10] ,
    \Tile_X4Y12_NN4BEG[9] ,
    \Tile_X4Y12_NN4BEG[8] ,
    \Tile_X4Y12_NN4BEG[7] ,
    \Tile_X4Y12_NN4BEG[6] ,
    \Tile_X4Y12_NN4BEG[5] ,
    \Tile_X4Y12_NN4BEG[4] ,
    \Tile_X4Y12_NN4BEG[3] ,
    \Tile_X4Y12_NN4BEG[2] ,
    \Tile_X4Y12_NN4BEG[1] ,
    \Tile_X4Y12_NN4BEG[0] }),
    .NN4END({\Tile_X4Y13_NN4BEG[15] ,
    \Tile_X4Y13_NN4BEG[14] ,
    \Tile_X4Y13_NN4BEG[13] ,
    \Tile_X4Y13_NN4BEG[12] ,
    \Tile_X4Y13_NN4BEG[11] ,
    \Tile_X4Y13_NN4BEG[10] ,
    \Tile_X4Y13_NN4BEG[9] ,
    \Tile_X4Y13_NN4BEG[8] ,
    \Tile_X4Y13_NN4BEG[7] ,
    \Tile_X4Y13_NN4BEG[6] ,
    \Tile_X4Y13_NN4BEG[5] ,
    \Tile_X4Y13_NN4BEG[4] ,
    \Tile_X4Y13_NN4BEG[3] ,
    \Tile_X4Y13_NN4BEG[2] ,
    \Tile_X4Y13_NN4BEG[1] ,
    \Tile_X4Y13_NN4BEG[0] }),
    .S1BEG({\Tile_X4Y12_S1BEG[3] ,
    \Tile_X4Y12_S1BEG[2] ,
    \Tile_X4Y12_S1BEG[1] ,
    \Tile_X4Y12_S1BEG[0] }),
    .S1END({\Tile_X4Y11_S1BEG[3] ,
    \Tile_X4Y11_S1BEG[2] ,
    \Tile_X4Y11_S1BEG[1] ,
    \Tile_X4Y11_S1BEG[0] }),
    .S2BEG({\Tile_X4Y12_S2BEG[7] ,
    \Tile_X4Y12_S2BEG[6] ,
    \Tile_X4Y12_S2BEG[5] ,
    \Tile_X4Y12_S2BEG[4] ,
    \Tile_X4Y12_S2BEG[3] ,
    \Tile_X4Y12_S2BEG[2] ,
    \Tile_X4Y12_S2BEG[1] ,
    \Tile_X4Y12_S2BEG[0] }),
    .S2BEGb({\Tile_X4Y12_S2BEGb[7] ,
    \Tile_X4Y12_S2BEGb[6] ,
    \Tile_X4Y12_S2BEGb[5] ,
    \Tile_X4Y12_S2BEGb[4] ,
    \Tile_X4Y12_S2BEGb[3] ,
    \Tile_X4Y12_S2BEGb[2] ,
    \Tile_X4Y12_S2BEGb[1] ,
    \Tile_X4Y12_S2BEGb[0] }),
    .S2END({\Tile_X4Y11_S2BEGb[7] ,
    \Tile_X4Y11_S2BEGb[6] ,
    \Tile_X4Y11_S2BEGb[5] ,
    \Tile_X4Y11_S2BEGb[4] ,
    \Tile_X4Y11_S2BEGb[3] ,
    \Tile_X4Y11_S2BEGb[2] ,
    \Tile_X4Y11_S2BEGb[1] ,
    \Tile_X4Y11_S2BEGb[0] }),
    .S2MID({\Tile_X4Y11_S2BEG[7] ,
    \Tile_X4Y11_S2BEG[6] ,
    \Tile_X4Y11_S2BEG[5] ,
    \Tile_X4Y11_S2BEG[4] ,
    \Tile_X4Y11_S2BEG[3] ,
    \Tile_X4Y11_S2BEG[2] ,
    \Tile_X4Y11_S2BEG[1] ,
    \Tile_X4Y11_S2BEG[0] }),
    .S4BEG({\Tile_X4Y12_S4BEG[15] ,
    \Tile_X4Y12_S4BEG[14] ,
    \Tile_X4Y12_S4BEG[13] ,
    \Tile_X4Y12_S4BEG[12] ,
    \Tile_X4Y12_S4BEG[11] ,
    \Tile_X4Y12_S4BEG[10] ,
    \Tile_X4Y12_S4BEG[9] ,
    \Tile_X4Y12_S4BEG[8] ,
    \Tile_X4Y12_S4BEG[7] ,
    \Tile_X4Y12_S4BEG[6] ,
    \Tile_X4Y12_S4BEG[5] ,
    \Tile_X4Y12_S4BEG[4] ,
    \Tile_X4Y12_S4BEG[3] ,
    \Tile_X4Y12_S4BEG[2] ,
    \Tile_X4Y12_S4BEG[1] ,
    \Tile_X4Y12_S4BEG[0] }),
    .S4END({\Tile_X4Y11_S4BEG[15] ,
    \Tile_X4Y11_S4BEG[14] ,
    \Tile_X4Y11_S4BEG[13] ,
    \Tile_X4Y11_S4BEG[12] ,
    \Tile_X4Y11_S4BEG[11] ,
    \Tile_X4Y11_S4BEG[10] ,
    \Tile_X4Y11_S4BEG[9] ,
    \Tile_X4Y11_S4BEG[8] ,
    \Tile_X4Y11_S4BEG[7] ,
    \Tile_X4Y11_S4BEG[6] ,
    \Tile_X4Y11_S4BEG[5] ,
    \Tile_X4Y11_S4BEG[4] ,
    \Tile_X4Y11_S4BEG[3] ,
    \Tile_X4Y11_S4BEG[2] ,
    \Tile_X4Y11_S4BEG[1] ,
    \Tile_X4Y11_S4BEG[0] }),
    .SS4BEG({\Tile_X4Y12_SS4BEG[15] ,
    \Tile_X4Y12_SS4BEG[14] ,
    \Tile_X4Y12_SS4BEG[13] ,
    \Tile_X4Y12_SS4BEG[12] ,
    \Tile_X4Y12_SS4BEG[11] ,
    \Tile_X4Y12_SS4BEG[10] ,
    \Tile_X4Y12_SS4BEG[9] ,
    \Tile_X4Y12_SS4BEG[8] ,
    \Tile_X4Y12_SS4BEG[7] ,
    \Tile_X4Y12_SS4BEG[6] ,
    \Tile_X4Y12_SS4BEG[5] ,
    \Tile_X4Y12_SS4BEG[4] ,
    \Tile_X4Y12_SS4BEG[3] ,
    \Tile_X4Y12_SS4BEG[2] ,
    \Tile_X4Y12_SS4BEG[1] ,
    \Tile_X4Y12_SS4BEG[0] }),
    .SS4END({\Tile_X4Y11_SS4BEG[15] ,
    \Tile_X4Y11_SS4BEG[14] ,
    \Tile_X4Y11_SS4BEG[13] ,
    \Tile_X4Y11_SS4BEG[12] ,
    \Tile_X4Y11_SS4BEG[11] ,
    \Tile_X4Y11_SS4BEG[10] ,
    \Tile_X4Y11_SS4BEG[9] ,
    \Tile_X4Y11_SS4BEG[8] ,
    \Tile_X4Y11_SS4BEG[7] ,
    \Tile_X4Y11_SS4BEG[6] ,
    \Tile_X4Y11_SS4BEG[5] ,
    \Tile_X4Y11_SS4BEG[4] ,
    \Tile_X4Y11_SS4BEG[3] ,
    \Tile_X4Y11_SS4BEG[2] ,
    \Tile_X4Y11_SS4BEG[1] ,
    \Tile_X4Y11_SS4BEG[0] }),
    .W1BEG({\Tile_X4Y12_W1BEG[3] ,
    \Tile_X4Y12_W1BEG[2] ,
    \Tile_X4Y12_W1BEG[1] ,
    \Tile_X4Y12_W1BEG[0] }),
    .W1END({\Tile_X5Y12_W1BEG[3] ,
    \Tile_X5Y12_W1BEG[2] ,
    \Tile_X5Y12_W1BEG[1] ,
    \Tile_X5Y12_W1BEG[0] }),
    .W2BEG({\Tile_X4Y12_W2BEG[7] ,
    \Tile_X4Y12_W2BEG[6] ,
    \Tile_X4Y12_W2BEG[5] ,
    \Tile_X4Y12_W2BEG[4] ,
    \Tile_X4Y12_W2BEG[3] ,
    \Tile_X4Y12_W2BEG[2] ,
    \Tile_X4Y12_W2BEG[1] ,
    \Tile_X4Y12_W2BEG[0] }),
    .W2BEGb({\Tile_X4Y12_W2BEGb[7] ,
    \Tile_X4Y12_W2BEGb[6] ,
    \Tile_X4Y12_W2BEGb[5] ,
    \Tile_X4Y12_W2BEGb[4] ,
    \Tile_X4Y12_W2BEGb[3] ,
    \Tile_X4Y12_W2BEGb[2] ,
    \Tile_X4Y12_W2BEGb[1] ,
    \Tile_X4Y12_W2BEGb[0] }),
    .W2END({\Tile_X5Y12_W2BEGb[7] ,
    \Tile_X5Y12_W2BEGb[6] ,
    \Tile_X5Y12_W2BEGb[5] ,
    \Tile_X5Y12_W2BEGb[4] ,
    \Tile_X5Y12_W2BEGb[3] ,
    \Tile_X5Y12_W2BEGb[2] ,
    \Tile_X5Y12_W2BEGb[1] ,
    \Tile_X5Y12_W2BEGb[0] }),
    .W2MID({\Tile_X5Y12_W2BEG[7] ,
    \Tile_X5Y12_W2BEG[6] ,
    \Tile_X5Y12_W2BEG[5] ,
    \Tile_X5Y12_W2BEG[4] ,
    \Tile_X5Y12_W2BEG[3] ,
    \Tile_X5Y12_W2BEG[2] ,
    \Tile_X5Y12_W2BEG[1] ,
    \Tile_X5Y12_W2BEG[0] }),
    .W6BEG({\Tile_X4Y12_W6BEG[11] ,
    \Tile_X4Y12_W6BEG[10] ,
    \Tile_X4Y12_W6BEG[9] ,
    \Tile_X4Y12_W6BEG[8] ,
    \Tile_X4Y12_W6BEG[7] ,
    \Tile_X4Y12_W6BEG[6] ,
    \Tile_X4Y12_W6BEG[5] ,
    \Tile_X4Y12_W6BEG[4] ,
    \Tile_X4Y12_W6BEG[3] ,
    \Tile_X4Y12_W6BEG[2] ,
    \Tile_X4Y12_W6BEG[1] ,
    \Tile_X4Y12_W6BEG[0] }),
    .W6END({\Tile_X5Y12_W6BEG[11] ,
    \Tile_X5Y12_W6BEG[10] ,
    \Tile_X5Y12_W6BEG[9] ,
    \Tile_X5Y12_W6BEG[8] ,
    \Tile_X5Y12_W6BEG[7] ,
    \Tile_X5Y12_W6BEG[6] ,
    \Tile_X5Y12_W6BEG[5] ,
    \Tile_X5Y12_W6BEG[4] ,
    \Tile_X5Y12_W6BEG[3] ,
    \Tile_X5Y12_W6BEG[2] ,
    \Tile_X5Y12_W6BEG[1] ,
    \Tile_X5Y12_W6BEG[0] }),
    .WW4BEG({\Tile_X4Y12_WW4BEG[15] ,
    \Tile_X4Y12_WW4BEG[14] ,
    \Tile_X4Y12_WW4BEG[13] ,
    \Tile_X4Y12_WW4BEG[12] ,
    \Tile_X4Y12_WW4BEG[11] ,
    \Tile_X4Y12_WW4BEG[10] ,
    \Tile_X4Y12_WW4BEG[9] ,
    \Tile_X4Y12_WW4BEG[8] ,
    \Tile_X4Y12_WW4BEG[7] ,
    \Tile_X4Y12_WW4BEG[6] ,
    \Tile_X4Y12_WW4BEG[5] ,
    \Tile_X4Y12_WW4BEG[4] ,
    \Tile_X4Y12_WW4BEG[3] ,
    \Tile_X4Y12_WW4BEG[2] ,
    \Tile_X4Y12_WW4BEG[1] ,
    \Tile_X4Y12_WW4BEG[0] }),
    .WW4END({\Tile_X5Y12_WW4BEG[15] ,
    \Tile_X5Y12_WW4BEG[14] ,
    \Tile_X5Y12_WW4BEG[13] ,
    \Tile_X5Y12_WW4BEG[12] ,
    \Tile_X5Y12_WW4BEG[11] ,
    \Tile_X5Y12_WW4BEG[10] ,
    \Tile_X5Y12_WW4BEG[9] ,
    \Tile_X5Y12_WW4BEG[8] ,
    \Tile_X5Y12_WW4BEG[7] ,
    \Tile_X5Y12_WW4BEG[6] ,
    \Tile_X5Y12_WW4BEG[5] ,
    \Tile_X5Y12_WW4BEG[4] ,
    \Tile_X5Y12_WW4BEG[3] ,
    \Tile_X5Y12_WW4BEG[2] ,
    \Tile_X5Y12_WW4BEG[1] ,
    \Tile_X5Y12_WW4BEG[0] }));
 RegFile Tile_X4Y13_RegFile (.UserCLK(Tile_X4Y14_UserCLKo),
    .UserCLKo(Tile_X4Y13_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X4Y13_E1BEG[3] ,
    \Tile_X4Y13_E1BEG[2] ,
    \Tile_X4Y13_E1BEG[1] ,
    \Tile_X4Y13_E1BEG[0] }),
    .E1END({\Tile_X3Y13_E1BEG[3] ,
    \Tile_X3Y13_E1BEG[2] ,
    \Tile_X3Y13_E1BEG[1] ,
    \Tile_X3Y13_E1BEG[0] }),
    .E2BEG({\Tile_X4Y13_E2BEG[7] ,
    \Tile_X4Y13_E2BEG[6] ,
    \Tile_X4Y13_E2BEG[5] ,
    \Tile_X4Y13_E2BEG[4] ,
    \Tile_X4Y13_E2BEG[3] ,
    \Tile_X4Y13_E2BEG[2] ,
    \Tile_X4Y13_E2BEG[1] ,
    \Tile_X4Y13_E2BEG[0] }),
    .E2BEGb({\Tile_X4Y13_E2BEGb[7] ,
    \Tile_X4Y13_E2BEGb[6] ,
    \Tile_X4Y13_E2BEGb[5] ,
    \Tile_X4Y13_E2BEGb[4] ,
    \Tile_X4Y13_E2BEGb[3] ,
    \Tile_X4Y13_E2BEGb[2] ,
    \Tile_X4Y13_E2BEGb[1] ,
    \Tile_X4Y13_E2BEGb[0] }),
    .E2END({\Tile_X3Y13_E2BEGb[7] ,
    \Tile_X3Y13_E2BEGb[6] ,
    \Tile_X3Y13_E2BEGb[5] ,
    \Tile_X3Y13_E2BEGb[4] ,
    \Tile_X3Y13_E2BEGb[3] ,
    \Tile_X3Y13_E2BEGb[2] ,
    \Tile_X3Y13_E2BEGb[1] ,
    \Tile_X3Y13_E2BEGb[0] }),
    .E2MID({\Tile_X3Y13_E2BEG[7] ,
    \Tile_X3Y13_E2BEG[6] ,
    \Tile_X3Y13_E2BEG[5] ,
    \Tile_X3Y13_E2BEG[4] ,
    \Tile_X3Y13_E2BEG[3] ,
    \Tile_X3Y13_E2BEG[2] ,
    \Tile_X3Y13_E2BEG[1] ,
    \Tile_X3Y13_E2BEG[0] }),
    .E6BEG({\Tile_X4Y13_E6BEG[11] ,
    \Tile_X4Y13_E6BEG[10] ,
    \Tile_X4Y13_E6BEG[9] ,
    \Tile_X4Y13_E6BEG[8] ,
    \Tile_X4Y13_E6BEG[7] ,
    \Tile_X4Y13_E6BEG[6] ,
    \Tile_X4Y13_E6BEG[5] ,
    \Tile_X4Y13_E6BEG[4] ,
    \Tile_X4Y13_E6BEG[3] ,
    \Tile_X4Y13_E6BEG[2] ,
    \Tile_X4Y13_E6BEG[1] ,
    \Tile_X4Y13_E6BEG[0] }),
    .E6END({\Tile_X3Y13_E6BEG[11] ,
    \Tile_X3Y13_E6BEG[10] ,
    \Tile_X3Y13_E6BEG[9] ,
    \Tile_X3Y13_E6BEG[8] ,
    \Tile_X3Y13_E6BEG[7] ,
    \Tile_X3Y13_E6BEG[6] ,
    \Tile_X3Y13_E6BEG[5] ,
    \Tile_X3Y13_E6BEG[4] ,
    \Tile_X3Y13_E6BEG[3] ,
    \Tile_X3Y13_E6BEG[2] ,
    \Tile_X3Y13_E6BEG[1] ,
    \Tile_X3Y13_E6BEG[0] }),
    .EE4BEG({\Tile_X4Y13_EE4BEG[15] ,
    \Tile_X4Y13_EE4BEG[14] ,
    \Tile_X4Y13_EE4BEG[13] ,
    \Tile_X4Y13_EE4BEG[12] ,
    \Tile_X4Y13_EE4BEG[11] ,
    \Tile_X4Y13_EE4BEG[10] ,
    \Tile_X4Y13_EE4BEG[9] ,
    \Tile_X4Y13_EE4BEG[8] ,
    \Tile_X4Y13_EE4BEG[7] ,
    \Tile_X4Y13_EE4BEG[6] ,
    \Tile_X4Y13_EE4BEG[5] ,
    \Tile_X4Y13_EE4BEG[4] ,
    \Tile_X4Y13_EE4BEG[3] ,
    \Tile_X4Y13_EE4BEG[2] ,
    \Tile_X4Y13_EE4BEG[1] ,
    \Tile_X4Y13_EE4BEG[0] }),
    .EE4END({\Tile_X3Y13_EE4BEG[15] ,
    \Tile_X3Y13_EE4BEG[14] ,
    \Tile_X3Y13_EE4BEG[13] ,
    \Tile_X3Y13_EE4BEG[12] ,
    \Tile_X3Y13_EE4BEG[11] ,
    \Tile_X3Y13_EE4BEG[10] ,
    \Tile_X3Y13_EE4BEG[9] ,
    \Tile_X3Y13_EE4BEG[8] ,
    \Tile_X3Y13_EE4BEG[7] ,
    \Tile_X3Y13_EE4BEG[6] ,
    \Tile_X3Y13_EE4BEG[5] ,
    \Tile_X3Y13_EE4BEG[4] ,
    \Tile_X3Y13_EE4BEG[3] ,
    \Tile_X3Y13_EE4BEG[2] ,
    \Tile_X3Y13_EE4BEG[1] ,
    \Tile_X3Y13_EE4BEG[0] }),
    .FrameData({\Tile_X3Y13_FrameData_O[31] ,
    \Tile_X3Y13_FrameData_O[30] ,
    \Tile_X3Y13_FrameData_O[29] ,
    \Tile_X3Y13_FrameData_O[28] ,
    \Tile_X3Y13_FrameData_O[27] ,
    \Tile_X3Y13_FrameData_O[26] ,
    \Tile_X3Y13_FrameData_O[25] ,
    \Tile_X3Y13_FrameData_O[24] ,
    \Tile_X3Y13_FrameData_O[23] ,
    \Tile_X3Y13_FrameData_O[22] ,
    \Tile_X3Y13_FrameData_O[21] ,
    \Tile_X3Y13_FrameData_O[20] ,
    \Tile_X3Y13_FrameData_O[19] ,
    \Tile_X3Y13_FrameData_O[18] ,
    \Tile_X3Y13_FrameData_O[17] ,
    \Tile_X3Y13_FrameData_O[16] ,
    \Tile_X3Y13_FrameData_O[15] ,
    \Tile_X3Y13_FrameData_O[14] ,
    \Tile_X3Y13_FrameData_O[13] ,
    \Tile_X3Y13_FrameData_O[12] ,
    \Tile_X3Y13_FrameData_O[11] ,
    \Tile_X3Y13_FrameData_O[10] ,
    \Tile_X3Y13_FrameData_O[9] ,
    \Tile_X3Y13_FrameData_O[8] ,
    \Tile_X3Y13_FrameData_O[7] ,
    \Tile_X3Y13_FrameData_O[6] ,
    \Tile_X3Y13_FrameData_O[5] ,
    \Tile_X3Y13_FrameData_O[4] ,
    \Tile_X3Y13_FrameData_O[3] ,
    \Tile_X3Y13_FrameData_O[2] ,
    \Tile_X3Y13_FrameData_O[1] ,
    \Tile_X3Y13_FrameData_O[0] }),
    .FrameData_O({\Tile_X4Y13_FrameData_O[31] ,
    \Tile_X4Y13_FrameData_O[30] ,
    \Tile_X4Y13_FrameData_O[29] ,
    \Tile_X4Y13_FrameData_O[28] ,
    \Tile_X4Y13_FrameData_O[27] ,
    \Tile_X4Y13_FrameData_O[26] ,
    \Tile_X4Y13_FrameData_O[25] ,
    \Tile_X4Y13_FrameData_O[24] ,
    \Tile_X4Y13_FrameData_O[23] ,
    \Tile_X4Y13_FrameData_O[22] ,
    \Tile_X4Y13_FrameData_O[21] ,
    \Tile_X4Y13_FrameData_O[20] ,
    \Tile_X4Y13_FrameData_O[19] ,
    \Tile_X4Y13_FrameData_O[18] ,
    \Tile_X4Y13_FrameData_O[17] ,
    \Tile_X4Y13_FrameData_O[16] ,
    \Tile_X4Y13_FrameData_O[15] ,
    \Tile_X4Y13_FrameData_O[14] ,
    \Tile_X4Y13_FrameData_O[13] ,
    \Tile_X4Y13_FrameData_O[12] ,
    \Tile_X4Y13_FrameData_O[11] ,
    \Tile_X4Y13_FrameData_O[10] ,
    \Tile_X4Y13_FrameData_O[9] ,
    \Tile_X4Y13_FrameData_O[8] ,
    \Tile_X4Y13_FrameData_O[7] ,
    \Tile_X4Y13_FrameData_O[6] ,
    \Tile_X4Y13_FrameData_O[5] ,
    \Tile_X4Y13_FrameData_O[4] ,
    \Tile_X4Y13_FrameData_O[3] ,
    \Tile_X4Y13_FrameData_O[2] ,
    \Tile_X4Y13_FrameData_O[1] ,
    \Tile_X4Y13_FrameData_O[0] }),
    .FrameStrobe({\Tile_X4Y14_FrameStrobe_O[19] ,
    \Tile_X4Y14_FrameStrobe_O[18] ,
    \Tile_X4Y14_FrameStrobe_O[17] ,
    \Tile_X4Y14_FrameStrobe_O[16] ,
    \Tile_X4Y14_FrameStrobe_O[15] ,
    \Tile_X4Y14_FrameStrobe_O[14] ,
    \Tile_X4Y14_FrameStrobe_O[13] ,
    \Tile_X4Y14_FrameStrobe_O[12] ,
    \Tile_X4Y14_FrameStrobe_O[11] ,
    \Tile_X4Y14_FrameStrobe_O[10] ,
    \Tile_X4Y14_FrameStrobe_O[9] ,
    \Tile_X4Y14_FrameStrobe_O[8] ,
    \Tile_X4Y14_FrameStrobe_O[7] ,
    \Tile_X4Y14_FrameStrobe_O[6] ,
    \Tile_X4Y14_FrameStrobe_O[5] ,
    \Tile_X4Y14_FrameStrobe_O[4] ,
    \Tile_X4Y14_FrameStrobe_O[3] ,
    \Tile_X4Y14_FrameStrobe_O[2] ,
    \Tile_X4Y14_FrameStrobe_O[1] ,
    \Tile_X4Y14_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X4Y13_FrameStrobe_O[19] ,
    \Tile_X4Y13_FrameStrobe_O[18] ,
    \Tile_X4Y13_FrameStrobe_O[17] ,
    \Tile_X4Y13_FrameStrobe_O[16] ,
    \Tile_X4Y13_FrameStrobe_O[15] ,
    \Tile_X4Y13_FrameStrobe_O[14] ,
    \Tile_X4Y13_FrameStrobe_O[13] ,
    \Tile_X4Y13_FrameStrobe_O[12] ,
    \Tile_X4Y13_FrameStrobe_O[11] ,
    \Tile_X4Y13_FrameStrobe_O[10] ,
    \Tile_X4Y13_FrameStrobe_O[9] ,
    \Tile_X4Y13_FrameStrobe_O[8] ,
    \Tile_X4Y13_FrameStrobe_O[7] ,
    \Tile_X4Y13_FrameStrobe_O[6] ,
    \Tile_X4Y13_FrameStrobe_O[5] ,
    \Tile_X4Y13_FrameStrobe_O[4] ,
    \Tile_X4Y13_FrameStrobe_O[3] ,
    \Tile_X4Y13_FrameStrobe_O[2] ,
    \Tile_X4Y13_FrameStrobe_O[1] ,
    \Tile_X4Y13_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X4Y13_N1BEG[3] ,
    \Tile_X4Y13_N1BEG[2] ,
    \Tile_X4Y13_N1BEG[1] ,
    \Tile_X4Y13_N1BEG[0] }),
    .N1END({\Tile_X4Y14_N1BEG[3] ,
    \Tile_X4Y14_N1BEG[2] ,
    \Tile_X4Y14_N1BEG[1] ,
    \Tile_X4Y14_N1BEG[0] }),
    .N2BEG({\Tile_X4Y13_N2BEG[7] ,
    \Tile_X4Y13_N2BEG[6] ,
    \Tile_X4Y13_N2BEG[5] ,
    \Tile_X4Y13_N2BEG[4] ,
    \Tile_X4Y13_N2BEG[3] ,
    \Tile_X4Y13_N2BEG[2] ,
    \Tile_X4Y13_N2BEG[1] ,
    \Tile_X4Y13_N2BEG[0] }),
    .N2BEGb({\Tile_X4Y13_N2BEGb[7] ,
    \Tile_X4Y13_N2BEGb[6] ,
    \Tile_X4Y13_N2BEGb[5] ,
    \Tile_X4Y13_N2BEGb[4] ,
    \Tile_X4Y13_N2BEGb[3] ,
    \Tile_X4Y13_N2BEGb[2] ,
    \Tile_X4Y13_N2BEGb[1] ,
    \Tile_X4Y13_N2BEGb[0] }),
    .N2END({\Tile_X4Y14_N2BEGb[7] ,
    \Tile_X4Y14_N2BEGb[6] ,
    \Tile_X4Y14_N2BEGb[5] ,
    \Tile_X4Y14_N2BEGb[4] ,
    \Tile_X4Y14_N2BEGb[3] ,
    \Tile_X4Y14_N2BEGb[2] ,
    \Tile_X4Y14_N2BEGb[1] ,
    \Tile_X4Y14_N2BEGb[0] }),
    .N2MID({\Tile_X4Y14_N2BEG[7] ,
    \Tile_X4Y14_N2BEG[6] ,
    \Tile_X4Y14_N2BEG[5] ,
    \Tile_X4Y14_N2BEG[4] ,
    \Tile_X4Y14_N2BEG[3] ,
    \Tile_X4Y14_N2BEG[2] ,
    \Tile_X4Y14_N2BEG[1] ,
    \Tile_X4Y14_N2BEG[0] }),
    .N4BEG({\Tile_X4Y13_N4BEG[15] ,
    \Tile_X4Y13_N4BEG[14] ,
    \Tile_X4Y13_N4BEG[13] ,
    \Tile_X4Y13_N4BEG[12] ,
    \Tile_X4Y13_N4BEG[11] ,
    \Tile_X4Y13_N4BEG[10] ,
    \Tile_X4Y13_N4BEG[9] ,
    \Tile_X4Y13_N4BEG[8] ,
    \Tile_X4Y13_N4BEG[7] ,
    \Tile_X4Y13_N4BEG[6] ,
    \Tile_X4Y13_N4BEG[5] ,
    \Tile_X4Y13_N4BEG[4] ,
    \Tile_X4Y13_N4BEG[3] ,
    \Tile_X4Y13_N4BEG[2] ,
    \Tile_X4Y13_N4BEG[1] ,
    \Tile_X4Y13_N4BEG[0] }),
    .N4END({\Tile_X4Y14_N4BEG[15] ,
    \Tile_X4Y14_N4BEG[14] ,
    \Tile_X4Y14_N4BEG[13] ,
    \Tile_X4Y14_N4BEG[12] ,
    \Tile_X4Y14_N4BEG[11] ,
    \Tile_X4Y14_N4BEG[10] ,
    \Tile_X4Y14_N4BEG[9] ,
    \Tile_X4Y14_N4BEG[8] ,
    \Tile_X4Y14_N4BEG[7] ,
    \Tile_X4Y14_N4BEG[6] ,
    \Tile_X4Y14_N4BEG[5] ,
    \Tile_X4Y14_N4BEG[4] ,
    \Tile_X4Y14_N4BEG[3] ,
    \Tile_X4Y14_N4BEG[2] ,
    \Tile_X4Y14_N4BEG[1] ,
    \Tile_X4Y14_N4BEG[0] }),
    .NN4BEG({\Tile_X4Y13_NN4BEG[15] ,
    \Tile_X4Y13_NN4BEG[14] ,
    \Tile_X4Y13_NN4BEG[13] ,
    \Tile_X4Y13_NN4BEG[12] ,
    \Tile_X4Y13_NN4BEG[11] ,
    \Tile_X4Y13_NN4BEG[10] ,
    \Tile_X4Y13_NN4BEG[9] ,
    \Tile_X4Y13_NN4BEG[8] ,
    \Tile_X4Y13_NN4BEG[7] ,
    \Tile_X4Y13_NN4BEG[6] ,
    \Tile_X4Y13_NN4BEG[5] ,
    \Tile_X4Y13_NN4BEG[4] ,
    \Tile_X4Y13_NN4BEG[3] ,
    \Tile_X4Y13_NN4BEG[2] ,
    \Tile_X4Y13_NN4BEG[1] ,
    \Tile_X4Y13_NN4BEG[0] }),
    .NN4END({\Tile_X4Y14_NN4BEG[15] ,
    \Tile_X4Y14_NN4BEG[14] ,
    \Tile_X4Y14_NN4BEG[13] ,
    \Tile_X4Y14_NN4BEG[12] ,
    \Tile_X4Y14_NN4BEG[11] ,
    \Tile_X4Y14_NN4BEG[10] ,
    \Tile_X4Y14_NN4BEG[9] ,
    \Tile_X4Y14_NN4BEG[8] ,
    \Tile_X4Y14_NN4BEG[7] ,
    \Tile_X4Y14_NN4BEG[6] ,
    \Tile_X4Y14_NN4BEG[5] ,
    \Tile_X4Y14_NN4BEG[4] ,
    \Tile_X4Y14_NN4BEG[3] ,
    \Tile_X4Y14_NN4BEG[2] ,
    \Tile_X4Y14_NN4BEG[1] ,
    \Tile_X4Y14_NN4BEG[0] }),
    .S1BEG({\Tile_X4Y13_S1BEG[3] ,
    \Tile_X4Y13_S1BEG[2] ,
    \Tile_X4Y13_S1BEG[1] ,
    \Tile_X4Y13_S1BEG[0] }),
    .S1END({\Tile_X4Y12_S1BEG[3] ,
    \Tile_X4Y12_S1BEG[2] ,
    \Tile_X4Y12_S1BEG[1] ,
    \Tile_X4Y12_S1BEG[0] }),
    .S2BEG({\Tile_X4Y13_S2BEG[7] ,
    \Tile_X4Y13_S2BEG[6] ,
    \Tile_X4Y13_S2BEG[5] ,
    \Tile_X4Y13_S2BEG[4] ,
    \Tile_X4Y13_S2BEG[3] ,
    \Tile_X4Y13_S2BEG[2] ,
    \Tile_X4Y13_S2BEG[1] ,
    \Tile_X4Y13_S2BEG[0] }),
    .S2BEGb({\Tile_X4Y13_S2BEGb[7] ,
    \Tile_X4Y13_S2BEGb[6] ,
    \Tile_X4Y13_S2BEGb[5] ,
    \Tile_X4Y13_S2BEGb[4] ,
    \Tile_X4Y13_S2BEGb[3] ,
    \Tile_X4Y13_S2BEGb[2] ,
    \Tile_X4Y13_S2BEGb[1] ,
    \Tile_X4Y13_S2BEGb[0] }),
    .S2END({\Tile_X4Y12_S2BEGb[7] ,
    \Tile_X4Y12_S2BEGb[6] ,
    \Tile_X4Y12_S2BEGb[5] ,
    \Tile_X4Y12_S2BEGb[4] ,
    \Tile_X4Y12_S2BEGb[3] ,
    \Tile_X4Y12_S2BEGb[2] ,
    \Tile_X4Y12_S2BEGb[1] ,
    \Tile_X4Y12_S2BEGb[0] }),
    .S2MID({\Tile_X4Y12_S2BEG[7] ,
    \Tile_X4Y12_S2BEG[6] ,
    \Tile_X4Y12_S2BEG[5] ,
    \Tile_X4Y12_S2BEG[4] ,
    \Tile_X4Y12_S2BEG[3] ,
    \Tile_X4Y12_S2BEG[2] ,
    \Tile_X4Y12_S2BEG[1] ,
    \Tile_X4Y12_S2BEG[0] }),
    .S4BEG({\Tile_X4Y13_S4BEG[15] ,
    \Tile_X4Y13_S4BEG[14] ,
    \Tile_X4Y13_S4BEG[13] ,
    \Tile_X4Y13_S4BEG[12] ,
    \Tile_X4Y13_S4BEG[11] ,
    \Tile_X4Y13_S4BEG[10] ,
    \Tile_X4Y13_S4BEG[9] ,
    \Tile_X4Y13_S4BEG[8] ,
    \Tile_X4Y13_S4BEG[7] ,
    \Tile_X4Y13_S4BEG[6] ,
    \Tile_X4Y13_S4BEG[5] ,
    \Tile_X4Y13_S4BEG[4] ,
    \Tile_X4Y13_S4BEG[3] ,
    \Tile_X4Y13_S4BEG[2] ,
    \Tile_X4Y13_S4BEG[1] ,
    \Tile_X4Y13_S4BEG[0] }),
    .S4END({\Tile_X4Y12_S4BEG[15] ,
    \Tile_X4Y12_S4BEG[14] ,
    \Tile_X4Y12_S4BEG[13] ,
    \Tile_X4Y12_S4BEG[12] ,
    \Tile_X4Y12_S4BEG[11] ,
    \Tile_X4Y12_S4BEG[10] ,
    \Tile_X4Y12_S4BEG[9] ,
    \Tile_X4Y12_S4BEG[8] ,
    \Tile_X4Y12_S4BEG[7] ,
    \Tile_X4Y12_S4BEG[6] ,
    \Tile_X4Y12_S4BEG[5] ,
    \Tile_X4Y12_S4BEG[4] ,
    \Tile_X4Y12_S4BEG[3] ,
    \Tile_X4Y12_S4BEG[2] ,
    \Tile_X4Y12_S4BEG[1] ,
    \Tile_X4Y12_S4BEG[0] }),
    .SS4BEG({\Tile_X4Y13_SS4BEG[15] ,
    \Tile_X4Y13_SS4BEG[14] ,
    \Tile_X4Y13_SS4BEG[13] ,
    \Tile_X4Y13_SS4BEG[12] ,
    \Tile_X4Y13_SS4BEG[11] ,
    \Tile_X4Y13_SS4BEG[10] ,
    \Tile_X4Y13_SS4BEG[9] ,
    \Tile_X4Y13_SS4BEG[8] ,
    \Tile_X4Y13_SS4BEG[7] ,
    \Tile_X4Y13_SS4BEG[6] ,
    \Tile_X4Y13_SS4BEG[5] ,
    \Tile_X4Y13_SS4BEG[4] ,
    \Tile_X4Y13_SS4BEG[3] ,
    \Tile_X4Y13_SS4BEG[2] ,
    \Tile_X4Y13_SS4BEG[1] ,
    \Tile_X4Y13_SS4BEG[0] }),
    .SS4END({\Tile_X4Y12_SS4BEG[15] ,
    \Tile_X4Y12_SS4BEG[14] ,
    \Tile_X4Y12_SS4BEG[13] ,
    \Tile_X4Y12_SS4BEG[12] ,
    \Tile_X4Y12_SS4BEG[11] ,
    \Tile_X4Y12_SS4BEG[10] ,
    \Tile_X4Y12_SS4BEG[9] ,
    \Tile_X4Y12_SS4BEG[8] ,
    \Tile_X4Y12_SS4BEG[7] ,
    \Tile_X4Y12_SS4BEG[6] ,
    \Tile_X4Y12_SS4BEG[5] ,
    \Tile_X4Y12_SS4BEG[4] ,
    \Tile_X4Y12_SS4BEG[3] ,
    \Tile_X4Y12_SS4BEG[2] ,
    \Tile_X4Y12_SS4BEG[1] ,
    \Tile_X4Y12_SS4BEG[0] }),
    .W1BEG({\Tile_X4Y13_W1BEG[3] ,
    \Tile_X4Y13_W1BEG[2] ,
    \Tile_X4Y13_W1BEG[1] ,
    \Tile_X4Y13_W1BEG[0] }),
    .W1END({\Tile_X5Y13_W1BEG[3] ,
    \Tile_X5Y13_W1BEG[2] ,
    \Tile_X5Y13_W1BEG[1] ,
    \Tile_X5Y13_W1BEG[0] }),
    .W2BEG({\Tile_X4Y13_W2BEG[7] ,
    \Tile_X4Y13_W2BEG[6] ,
    \Tile_X4Y13_W2BEG[5] ,
    \Tile_X4Y13_W2BEG[4] ,
    \Tile_X4Y13_W2BEG[3] ,
    \Tile_X4Y13_W2BEG[2] ,
    \Tile_X4Y13_W2BEG[1] ,
    \Tile_X4Y13_W2BEG[0] }),
    .W2BEGb({\Tile_X4Y13_W2BEGb[7] ,
    \Tile_X4Y13_W2BEGb[6] ,
    \Tile_X4Y13_W2BEGb[5] ,
    \Tile_X4Y13_W2BEGb[4] ,
    \Tile_X4Y13_W2BEGb[3] ,
    \Tile_X4Y13_W2BEGb[2] ,
    \Tile_X4Y13_W2BEGb[1] ,
    \Tile_X4Y13_W2BEGb[0] }),
    .W2END({\Tile_X5Y13_W2BEGb[7] ,
    \Tile_X5Y13_W2BEGb[6] ,
    \Tile_X5Y13_W2BEGb[5] ,
    \Tile_X5Y13_W2BEGb[4] ,
    \Tile_X5Y13_W2BEGb[3] ,
    \Tile_X5Y13_W2BEGb[2] ,
    \Tile_X5Y13_W2BEGb[1] ,
    \Tile_X5Y13_W2BEGb[0] }),
    .W2MID({\Tile_X5Y13_W2BEG[7] ,
    \Tile_X5Y13_W2BEG[6] ,
    \Tile_X5Y13_W2BEG[5] ,
    \Tile_X5Y13_W2BEG[4] ,
    \Tile_X5Y13_W2BEG[3] ,
    \Tile_X5Y13_W2BEG[2] ,
    \Tile_X5Y13_W2BEG[1] ,
    \Tile_X5Y13_W2BEG[0] }),
    .W6BEG({\Tile_X4Y13_W6BEG[11] ,
    \Tile_X4Y13_W6BEG[10] ,
    \Tile_X4Y13_W6BEG[9] ,
    \Tile_X4Y13_W6BEG[8] ,
    \Tile_X4Y13_W6BEG[7] ,
    \Tile_X4Y13_W6BEG[6] ,
    \Tile_X4Y13_W6BEG[5] ,
    \Tile_X4Y13_W6BEG[4] ,
    \Tile_X4Y13_W6BEG[3] ,
    \Tile_X4Y13_W6BEG[2] ,
    \Tile_X4Y13_W6BEG[1] ,
    \Tile_X4Y13_W6BEG[0] }),
    .W6END({\Tile_X5Y13_W6BEG[11] ,
    \Tile_X5Y13_W6BEG[10] ,
    \Tile_X5Y13_W6BEG[9] ,
    \Tile_X5Y13_W6BEG[8] ,
    \Tile_X5Y13_W6BEG[7] ,
    \Tile_X5Y13_W6BEG[6] ,
    \Tile_X5Y13_W6BEG[5] ,
    \Tile_X5Y13_W6BEG[4] ,
    \Tile_X5Y13_W6BEG[3] ,
    \Tile_X5Y13_W6BEG[2] ,
    \Tile_X5Y13_W6BEG[1] ,
    \Tile_X5Y13_W6BEG[0] }),
    .WW4BEG({\Tile_X4Y13_WW4BEG[15] ,
    \Tile_X4Y13_WW4BEG[14] ,
    \Tile_X4Y13_WW4BEG[13] ,
    \Tile_X4Y13_WW4BEG[12] ,
    \Tile_X4Y13_WW4BEG[11] ,
    \Tile_X4Y13_WW4BEG[10] ,
    \Tile_X4Y13_WW4BEG[9] ,
    \Tile_X4Y13_WW4BEG[8] ,
    \Tile_X4Y13_WW4BEG[7] ,
    \Tile_X4Y13_WW4BEG[6] ,
    \Tile_X4Y13_WW4BEG[5] ,
    \Tile_X4Y13_WW4BEG[4] ,
    \Tile_X4Y13_WW4BEG[3] ,
    \Tile_X4Y13_WW4BEG[2] ,
    \Tile_X4Y13_WW4BEG[1] ,
    \Tile_X4Y13_WW4BEG[0] }),
    .WW4END({\Tile_X5Y13_WW4BEG[15] ,
    \Tile_X5Y13_WW4BEG[14] ,
    \Tile_X5Y13_WW4BEG[13] ,
    \Tile_X5Y13_WW4BEG[12] ,
    \Tile_X5Y13_WW4BEG[11] ,
    \Tile_X5Y13_WW4BEG[10] ,
    \Tile_X5Y13_WW4BEG[9] ,
    \Tile_X5Y13_WW4BEG[8] ,
    \Tile_X5Y13_WW4BEG[7] ,
    \Tile_X5Y13_WW4BEG[6] ,
    \Tile_X5Y13_WW4BEG[5] ,
    \Tile_X5Y13_WW4BEG[4] ,
    \Tile_X5Y13_WW4BEG[3] ,
    \Tile_X5Y13_WW4BEG[2] ,
    \Tile_X5Y13_WW4BEG[1] ,
    \Tile_X5Y13_WW4BEG[0] }));
 RegFile Tile_X4Y14_RegFile (.UserCLK(Tile_X4Y15_UserCLKo),
    .UserCLKo(Tile_X4Y14_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X4Y14_E1BEG[3] ,
    \Tile_X4Y14_E1BEG[2] ,
    \Tile_X4Y14_E1BEG[1] ,
    \Tile_X4Y14_E1BEG[0] }),
    .E1END({\Tile_X3Y14_E1BEG[3] ,
    \Tile_X3Y14_E1BEG[2] ,
    \Tile_X3Y14_E1BEG[1] ,
    \Tile_X3Y14_E1BEG[0] }),
    .E2BEG({\Tile_X4Y14_E2BEG[7] ,
    \Tile_X4Y14_E2BEG[6] ,
    \Tile_X4Y14_E2BEG[5] ,
    \Tile_X4Y14_E2BEG[4] ,
    \Tile_X4Y14_E2BEG[3] ,
    \Tile_X4Y14_E2BEG[2] ,
    \Tile_X4Y14_E2BEG[1] ,
    \Tile_X4Y14_E2BEG[0] }),
    .E2BEGb({\Tile_X4Y14_E2BEGb[7] ,
    \Tile_X4Y14_E2BEGb[6] ,
    \Tile_X4Y14_E2BEGb[5] ,
    \Tile_X4Y14_E2BEGb[4] ,
    \Tile_X4Y14_E2BEGb[3] ,
    \Tile_X4Y14_E2BEGb[2] ,
    \Tile_X4Y14_E2BEGb[1] ,
    \Tile_X4Y14_E2BEGb[0] }),
    .E2END({\Tile_X3Y14_E2BEGb[7] ,
    \Tile_X3Y14_E2BEGb[6] ,
    \Tile_X3Y14_E2BEGb[5] ,
    \Tile_X3Y14_E2BEGb[4] ,
    \Tile_X3Y14_E2BEGb[3] ,
    \Tile_X3Y14_E2BEGb[2] ,
    \Tile_X3Y14_E2BEGb[1] ,
    \Tile_X3Y14_E2BEGb[0] }),
    .E2MID({\Tile_X3Y14_E2BEG[7] ,
    \Tile_X3Y14_E2BEG[6] ,
    \Tile_X3Y14_E2BEG[5] ,
    \Tile_X3Y14_E2BEG[4] ,
    \Tile_X3Y14_E2BEG[3] ,
    \Tile_X3Y14_E2BEG[2] ,
    \Tile_X3Y14_E2BEG[1] ,
    \Tile_X3Y14_E2BEG[0] }),
    .E6BEG({\Tile_X4Y14_E6BEG[11] ,
    \Tile_X4Y14_E6BEG[10] ,
    \Tile_X4Y14_E6BEG[9] ,
    \Tile_X4Y14_E6BEG[8] ,
    \Tile_X4Y14_E6BEG[7] ,
    \Tile_X4Y14_E6BEG[6] ,
    \Tile_X4Y14_E6BEG[5] ,
    \Tile_X4Y14_E6BEG[4] ,
    \Tile_X4Y14_E6BEG[3] ,
    \Tile_X4Y14_E6BEG[2] ,
    \Tile_X4Y14_E6BEG[1] ,
    \Tile_X4Y14_E6BEG[0] }),
    .E6END({\Tile_X3Y14_E6BEG[11] ,
    \Tile_X3Y14_E6BEG[10] ,
    \Tile_X3Y14_E6BEG[9] ,
    \Tile_X3Y14_E6BEG[8] ,
    \Tile_X3Y14_E6BEG[7] ,
    \Tile_X3Y14_E6BEG[6] ,
    \Tile_X3Y14_E6BEG[5] ,
    \Tile_X3Y14_E6BEG[4] ,
    \Tile_X3Y14_E6BEG[3] ,
    \Tile_X3Y14_E6BEG[2] ,
    \Tile_X3Y14_E6BEG[1] ,
    \Tile_X3Y14_E6BEG[0] }),
    .EE4BEG({\Tile_X4Y14_EE4BEG[15] ,
    \Tile_X4Y14_EE4BEG[14] ,
    \Tile_X4Y14_EE4BEG[13] ,
    \Tile_X4Y14_EE4BEG[12] ,
    \Tile_X4Y14_EE4BEG[11] ,
    \Tile_X4Y14_EE4BEG[10] ,
    \Tile_X4Y14_EE4BEG[9] ,
    \Tile_X4Y14_EE4BEG[8] ,
    \Tile_X4Y14_EE4BEG[7] ,
    \Tile_X4Y14_EE4BEG[6] ,
    \Tile_X4Y14_EE4BEG[5] ,
    \Tile_X4Y14_EE4BEG[4] ,
    \Tile_X4Y14_EE4BEG[3] ,
    \Tile_X4Y14_EE4BEG[2] ,
    \Tile_X4Y14_EE4BEG[1] ,
    \Tile_X4Y14_EE4BEG[0] }),
    .EE4END({\Tile_X3Y14_EE4BEG[15] ,
    \Tile_X3Y14_EE4BEG[14] ,
    \Tile_X3Y14_EE4BEG[13] ,
    \Tile_X3Y14_EE4BEG[12] ,
    \Tile_X3Y14_EE4BEG[11] ,
    \Tile_X3Y14_EE4BEG[10] ,
    \Tile_X3Y14_EE4BEG[9] ,
    \Tile_X3Y14_EE4BEG[8] ,
    \Tile_X3Y14_EE4BEG[7] ,
    \Tile_X3Y14_EE4BEG[6] ,
    \Tile_X3Y14_EE4BEG[5] ,
    \Tile_X3Y14_EE4BEG[4] ,
    \Tile_X3Y14_EE4BEG[3] ,
    \Tile_X3Y14_EE4BEG[2] ,
    \Tile_X3Y14_EE4BEG[1] ,
    \Tile_X3Y14_EE4BEG[0] }),
    .FrameData({\Tile_X3Y14_FrameData_O[31] ,
    \Tile_X3Y14_FrameData_O[30] ,
    \Tile_X3Y14_FrameData_O[29] ,
    \Tile_X3Y14_FrameData_O[28] ,
    \Tile_X3Y14_FrameData_O[27] ,
    \Tile_X3Y14_FrameData_O[26] ,
    \Tile_X3Y14_FrameData_O[25] ,
    \Tile_X3Y14_FrameData_O[24] ,
    \Tile_X3Y14_FrameData_O[23] ,
    \Tile_X3Y14_FrameData_O[22] ,
    \Tile_X3Y14_FrameData_O[21] ,
    \Tile_X3Y14_FrameData_O[20] ,
    \Tile_X3Y14_FrameData_O[19] ,
    \Tile_X3Y14_FrameData_O[18] ,
    \Tile_X3Y14_FrameData_O[17] ,
    \Tile_X3Y14_FrameData_O[16] ,
    \Tile_X3Y14_FrameData_O[15] ,
    \Tile_X3Y14_FrameData_O[14] ,
    \Tile_X3Y14_FrameData_O[13] ,
    \Tile_X3Y14_FrameData_O[12] ,
    \Tile_X3Y14_FrameData_O[11] ,
    \Tile_X3Y14_FrameData_O[10] ,
    \Tile_X3Y14_FrameData_O[9] ,
    \Tile_X3Y14_FrameData_O[8] ,
    \Tile_X3Y14_FrameData_O[7] ,
    \Tile_X3Y14_FrameData_O[6] ,
    \Tile_X3Y14_FrameData_O[5] ,
    \Tile_X3Y14_FrameData_O[4] ,
    \Tile_X3Y14_FrameData_O[3] ,
    \Tile_X3Y14_FrameData_O[2] ,
    \Tile_X3Y14_FrameData_O[1] ,
    \Tile_X3Y14_FrameData_O[0] }),
    .FrameData_O({\Tile_X4Y14_FrameData_O[31] ,
    \Tile_X4Y14_FrameData_O[30] ,
    \Tile_X4Y14_FrameData_O[29] ,
    \Tile_X4Y14_FrameData_O[28] ,
    \Tile_X4Y14_FrameData_O[27] ,
    \Tile_X4Y14_FrameData_O[26] ,
    \Tile_X4Y14_FrameData_O[25] ,
    \Tile_X4Y14_FrameData_O[24] ,
    \Tile_X4Y14_FrameData_O[23] ,
    \Tile_X4Y14_FrameData_O[22] ,
    \Tile_X4Y14_FrameData_O[21] ,
    \Tile_X4Y14_FrameData_O[20] ,
    \Tile_X4Y14_FrameData_O[19] ,
    \Tile_X4Y14_FrameData_O[18] ,
    \Tile_X4Y14_FrameData_O[17] ,
    \Tile_X4Y14_FrameData_O[16] ,
    \Tile_X4Y14_FrameData_O[15] ,
    \Tile_X4Y14_FrameData_O[14] ,
    \Tile_X4Y14_FrameData_O[13] ,
    \Tile_X4Y14_FrameData_O[12] ,
    \Tile_X4Y14_FrameData_O[11] ,
    \Tile_X4Y14_FrameData_O[10] ,
    \Tile_X4Y14_FrameData_O[9] ,
    \Tile_X4Y14_FrameData_O[8] ,
    \Tile_X4Y14_FrameData_O[7] ,
    \Tile_X4Y14_FrameData_O[6] ,
    \Tile_X4Y14_FrameData_O[5] ,
    \Tile_X4Y14_FrameData_O[4] ,
    \Tile_X4Y14_FrameData_O[3] ,
    \Tile_X4Y14_FrameData_O[2] ,
    \Tile_X4Y14_FrameData_O[1] ,
    \Tile_X4Y14_FrameData_O[0] }),
    .FrameStrobe({\Tile_X4Y15_FrameStrobe_O[19] ,
    \Tile_X4Y15_FrameStrobe_O[18] ,
    \Tile_X4Y15_FrameStrobe_O[17] ,
    \Tile_X4Y15_FrameStrobe_O[16] ,
    \Tile_X4Y15_FrameStrobe_O[15] ,
    \Tile_X4Y15_FrameStrobe_O[14] ,
    \Tile_X4Y15_FrameStrobe_O[13] ,
    \Tile_X4Y15_FrameStrobe_O[12] ,
    \Tile_X4Y15_FrameStrobe_O[11] ,
    \Tile_X4Y15_FrameStrobe_O[10] ,
    \Tile_X4Y15_FrameStrobe_O[9] ,
    \Tile_X4Y15_FrameStrobe_O[8] ,
    \Tile_X4Y15_FrameStrobe_O[7] ,
    \Tile_X4Y15_FrameStrobe_O[6] ,
    \Tile_X4Y15_FrameStrobe_O[5] ,
    \Tile_X4Y15_FrameStrobe_O[4] ,
    \Tile_X4Y15_FrameStrobe_O[3] ,
    \Tile_X4Y15_FrameStrobe_O[2] ,
    \Tile_X4Y15_FrameStrobe_O[1] ,
    \Tile_X4Y15_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X4Y14_FrameStrobe_O[19] ,
    \Tile_X4Y14_FrameStrobe_O[18] ,
    \Tile_X4Y14_FrameStrobe_O[17] ,
    \Tile_X4Y14_FrameStrobe_O[16] ,
    \Tile_X4Y14_FrameStrobe_O[15] ,
    \Tile_X4Y14_FrameStrobe_O[14] ,
    \Tile_X4Y14_FrameStrobe_O[13] ,
    \Tile_X4Y14_FrameStrobe_O[12] ,
    \Tile_X4Y14_FrameStrobe_O[11] ,
    \Tile_X4Y14_FrameStrobe_O[10] ,
    \Tile_X4Y14_FrameStrobe_O[9] ,
    \Tile_X4Y14_FrameStrobe_O[8] ,
    \Tile_X4Y14_FrameStrobe_O[7] ,
    \Tile_X4Y14_FrameStrobe_O[6] ,
    \Tile_X4Y14_FrameStrobe_O[5] ,
    \Tile_X4Y14_FrameStrobe_O[4] ,
    \Tile_X4Y14_FrameStrobe_O[3] ,
    \Tile_X4Y14_FrameStrobe_O[2] ,
    \Tile_X4Y14_FrameStrobe_O[1] ,
    \Tile_X4Y14_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X4Y14_N1BEG[3] ,
    \Tile_X4Y14_N1BEG[2] ,
    \Tile_X4Y14_N1BEG[1] ,
    \Tile_X4Y14_N1BEG[0] }),
    .N1END({\Tile_X4Y15_N1BEG[3] ,
    \Tile_X4Y15_N1BEG[2] ,
    \Tile_X4Y15_N1BEG[1] ,
    \Tile_X4Y15_N1BEG[0] }),
    .N2BEG({\Tile_X4Y14_N2BEG[7] ,
    \Tile_X4Y14_N2BEG[6] ,
    \Tile_X4Y14_N2BEG[5] ,
    \Tile_X4Y14_N2BEG[4] ,
    \Tile_X4Y14_N2BEG[3] ,
    \Tile_X4Y14_N2BEG[2] ,
    \Tile_X4Y14_N2BEG[1] ,
    \Tile_X4Y14_N2BEG[0] }),
    .N2BEGb({\Tile_X4Y14_N2BEGb[7] ,
    \Tile_X4Y14_N2BEGb[6] ,
    \Tile_X4Y14_N2BEGb[5] ,
    \Tile_X4Y14_N2BEGb[4] ,
    \Tile_X4Y14_N2BEGb[3] ,
    \Tile_X4Y14_N2BEGb[2] ,
    \Tile_X4Y14_N2BEGb[1] ,
    \Tile_X4Y14_N2BEGb[0] }),
    .N2END({\Tile_X4Y15_N2BEGb[7] ,
    \Tile_X4Y15_N2BEGb[6] ,
    \Tile_X4Y15_N2BEGb[5] ,
    \Tile_X4Y15_N2BEGb[4] ,
    \Tile_X4Y15_N2BEGb[3] ,
    \Tile_X4Y15_N2BEGb[2] ,
    \Tile_X4Y15_N2BEGb[1] ,
    \Tile_X4Y15_N2BEGb[0] }),
    .N2MID({\Tile_X4Y15_N2BEG[7] ,
    \Tile_X4Y15_N2BEG[6] ,
    \Tile_X4Y15_N2BEG[5] ,
    \Tile_X4Y15_N2BEG[4] ,
    \Tile_X4Y15_N2BEG[3] ,
    \Tile_X4Y15_N2BEG[2] ,
    \Tile_X4Y15_N2BEG[1] ,
    \Tile_X4Y15_N2BEG[0] }),
    .N4BEG({\Tile_X4Y14_N4BEG[15] ,
    \Tile_X4Y14_N4BEG[14] ,
    \Tile_X4Y14_N4BEG[13] ,
    \Tile_X4Y14_N4BEG[12] ,
    \Tile_X4Y14_N4BEG[11] ,
    \Tile_X4Y14_N4BEG[10] ,
    \Tile_X4Y14_N4BEG[9] ,
    \Tile_X4Y14_N4BEG[8] ,
    \Tile_X4Y14_N4BEG[7] ,
    \Tile_X4Y14_N4BEG[6] ,
    \Tile_X4Y14_N4BEG[5] ,
    \Tile_X4Y14_N4BEG[4] ,
    \Tile_X4Y14_N4BEG[3] ,
    \Tile_X4Y14_N4BEG[2] ,
    \Tile_X4Y14_N4BEG[1] ,
    \Tile_X4Y14_N4BEG[0] }),
    .N4END({\Tile_X4Y15_N4BEG[15] ,
    \Tile_X4Y15_N4BEG[14] ,
    \Tile_X4Y15_N4BEG[13] ,
    \Tile_X4Y15_N4BEG[12] ,
    \Tile_X4Y15_N4BEG[11] ,
    \Tile_X4Y15_N4BEG[10] ,
    \Tile_X4Y15_N4BEG[9] ,
    \Tile_X4Y15_N4BEG[8] ,
    \Tile_X4Y15_N4BEG[7] ,
    \Tile_X4Y15_N4BEG[6] ,
    \Tile_X4Y15_N4BEG[5] ,
    \Tile_X4Y15_N4BEG[4] ,
    \Tile_X4Y15_N4BEG[3] ,
    \Tile_X4Y15_N4BEG[2] ,
    \Tile_X4Y15_N4BEG[1] ,
    \Tile_X4Y15_N4BEG[0] }),
    .NN4BEG({\Tile_X4Y14_NN4BEG[15] ,
    \Tile_X4Y14_NN4BEG[14] ,
    \Tile_X4Y14_NN4BEG[13] ,
    \Tile_X4Y14_NN4BEG[12] ,
    \Tile_X4Y14_NN4BEG[11] ,
    \Tile_X4Y14_NN4BEG[10] ,
    \Tile_X4Y14_NN4BEG[9] ,
    \Tile_X4Y14_NN4BEG[8] ,
    \Tile_X4Y14_NN4BEG[7] ,
    \Tile_X4Y14_NN4BEG[6] ,
    \Tile_X4Y14_NN4BEG[5] ,
    \Tile_X4Y14_NN4BEG[4] ,
    \Tile_X4Y14_NN4BEG[3] ,
    \Tile_X4Y14_NN4BEG[2] ,
    \Tile_X4Y14_NN4BEG[1] ,
    \Tile_X4Y14_NN4BEG[0] }),
    .NN4END({\Tile_X4Y15_NN4BEG[15] ,
    \Tile_X4Y15_NN4BEG[14] ,
    \Tile_X4Y15_NN4BEG[13] ,
    \Tile_X4Y15_NN4BEG[12] ,
    \Tile_X4Y15_NN4BEG[11] ,
    \Tile_X4Y15_NN4BEG[10] ,
    \Tile_X4Y15_NN4BEG[9] ,
    \Tile_X4Y15_NN4BEG[8] ,
    \Tile_X4Y15_NN4BEG[7] ,
    \Tile_X4Y15_NN4BEG[6] ,
    \Tile_X4Y15_NN4BEG[5] ,
    \Tile_X4Y15_NN4BEG[4] ,
    \Tile_X4Y15_NN4BEG[3] ,
    \Tile_X4Y15_NN4BEG[2] ,
    \Tile_X4Y15_NN4BEG[1] ,
    \Tile_X4Y15_NN4BEG[0] }),
    .S1BEG({\Tile_X4Y14_S1BEG[3] ,
    \Tile_X4Y14_S1BEG[2] ,
    \Tile_X4Y14_S1BEG[1] ,
    \Tile_X4Y14_S1BEG[0] }),
    .S1END({\Tile_X4Y13_S1BEG[3] ,
    \Tile_X4Y13_S1BEG[2] ,
    \Tile_X4Y13_S1BEG[1] ,
    \Tile_X4Y13_S1BEG[0] }),
    .S2BEG({\Tile_X4Y14_S2BEG[7] ,
    \Tile_X4Y14_S2BEG[6] ,
    \Tile_X4Y14_S2BEG[5] ,
    \Tile_X4Y14_S2BEG[4] ,
    \Tile_X4Y14_S2BEG[3] ,
    \Tile_X4Y14_S2BEG[2] ,
    \Tile_X4Y14_S2BEG[1] ,
    \Tile_X4Y14_S2BEG[0] }),
    .S2BEGb({\Tile_X4Y14_S2BEGb[7] ,
    \Tile_X4Y14_S2BEGb[6] ,
    \Tile_X4Y14_S2BEGb[5] ,
    \Tile_X4Y14_S2BEGb[4] ,
    \Tile_X4Y14_S2BEGb[3] ,
    \Tile_X4Y14_S2BEGb[2] ,
    \Tile_X4Y14_S2BEGb[1] ,
    \Tile_X4Y14_S2BEGb[0] }),
    .S2END({\Tile_X4Y13_S2BEGb[7] ,
    \Tile_X4Y13_S2BEGb[6] ,
    \Tile_X4Y13_S2BEGb[5] ,
    \Tile_X4Y13_S2BEGb[4] ,
    \Tile_X4Y13_S2BEGb[3] ,
    \Tile_X4Y13_S2BEGb[2] ,
    \Tile_X4Y13_S2BEGb[1] ,
    \Tile_X4Y13_S2BEGb[0] }),
    .S2MID({\Tile_X4Y13_S2BEG[7] ,
    \Tile_X4Y13_S2BEG[6] ,
    \Tile_X4Y13_S2BEG[5] ,
    \Tile_X4Y13_S2BEG[4] ,
    \Tile_X4Y13_S2BEG[3] ,
    \Tile_X4Y13_S2BEG[2] ,
    \Tile_X4Y13_S2BEG[1] ,
    \Tile_X4Y13_S2BEG[0] }),
    .S4BEG({\Tile_X4Y14_S4BEG[15] ,
    \Tile_X4Y14_S4BEG[14] ,
    \Tile_X4Y14_S4BEG[13] ,
    \Tile_X4Y14_S4BEG[12] ,
    \Tile_X4Y14_S4BEG[11] ,
    \Tile_X4Y14_S4BEG[10] ,
    \Tile_X4Y14_S4BEG[9] ,
    \Tile_X4Y14_S4BEG[8] ,
    \Tile_X4Y14_S4BEG[7] ,
    \Tile_X4Y14_S4BEG[6] ,
    \Tile_X4Y14_S4BEG[5] ,
    \Tile_X4Y14_S4BEG[4] ,
    \Tile_X4Y14_S4BEG[3] ,
    \Tile_X4Y14_S4BEG[2] ,
    \Tile_X4Y14_S4BEG[1] ,
    \Tile_X4Y14_S4BEG[0] }),
    .S4END({\Tile_X4Y13_S4BEG[15] ,
    \Tile_X4Y13_S4BEG[14] ,
    \Tile_X4Y13_S4BEG[13] ,
    \Tile_X4Y13_S4BEG[12] ,
    \Tile_X4Y13_S4BEG[11] ,
    \Tile_X4Y13_S4BEG[10] ,
    \Tile_X4Y13_S4BEG[9] ,
    \Tile_X4Y13_S4BEG[8] ,
    \Tile_X4Y13_S4BEG[7] ,
    \Tile_X4Y13_S4BEG[6] ,
    \Tile_X4Y13_S4BEG[5] ,
    \Tile_X4Y13_S4BEG[4] ,
    \Tile_X4Y13_S4BEG[3] ,
    \Tile_X4Y13_S4BEG[2] ,
    \Tile_X4Y13_S4BEG[1] ,
    \Tile_X4Y13_S4BEG[0] }),
    .SS4BEG({\Tile_X4Y14_SS4BEG[15] ,
    \Tile_X4Y14_SS4BEG[14] ,
    \Tile_X4Y14_SS4BEG[13] ,
    \Tile_X4Y14_SS4BEG[12] ,
    \Tile_X4Y14_SS4BEG[11] ,
    \Tile_X4Y14_SS4BEG[10] ,
    \Tile_X4Y14_SS4BEG[9] ,
    \Tile_X4Y14_SS4BEG[8] ,
    \Tile_X4Y14_SS4BEG[7] ,
    \Tile_X4Y14_SS4BEG[6] ,
    \Tile_X4Y14_SS4BEG[5] ,
    \Tile_X4Y14_SS4BEG[4] ,
    \Tile_X4Y14_SS4BEG[3] ,
    \Tile_X4Y14_SS4BEG[2] ,
    \Tile_X4Y14_SS4BEG[1] ,
    \Tile_X4Y14_SS4BEG[0] }),
    .SS4END({\Tile_X4Y13_SS4BEG[15] ,
    \Tile_X4Y13_SS4BEG[14] ,
    \Tile_X4Y13_SS4BEG[13] ,
    \Tile_X4Y13_SS4BEG[12] ,
    \Tile_X4Y13_SS4BEG[11] ,
    \Tile_X4Y13_SS4BEG[10] ,
    \Tile_X4Y13_SS4BEG[9] ,
    \Tile_X4Y13_SS4BEG[8] ,
    \Tile_X4Y13_SS4BEG[7] ,
    \Tile_X4Y13_SS4BEG[6] ,
    \Tile_X4Y13_SS4BEG[5] ,
    \Tile_X4Y13_SS4BEG[4] ,
    \Tile_X4Y13_SS4BEG[3] ,
    \Tile_X4Y13_SS4BEG[2] ,
    \Tile_X4Y13_SS4BEG[1] ,
    \Tile_X4Y13_SS4BEG[0] }),
    .W1BEG({\Tile_X4Y14_W1BEG[3] ,
    \Tile_X4Y14_W1BEG[2] ,
    \Tile_X4Y14_W1BEG[1] ,
    \Tile_X4Y14_W1BEG[0] }),
    .W1END({\Tile_X5Y14_W1BEG[3] ,
    \Tile_X5Y14_W1BEG[2] ,
    \Tile_X5Y14_W1BEG[1] ,
    \Tile_X5Y14_W1BEG[0] }),
    .W2BEG({\Tile_X4Y14_W2BEG[7] ,
    \Tile_X4Y14_W2BEG[6] ,
    \Tile_X4Y14_W2BEG[5] ,
    \Tile_X4Y14_W2BEG[4] ,
    \Tile_X4Y14_W2BEG[3] ,
    \Tile_X4Y14_W2BEG[2] ,
    \Tile_X4Y14_W2BEG[1] ,
    \Tile_X4Y14_W2BEG[0] }),
    .W2BEGb({\Tile_X4Y14_W2BEGb[7] ,
    \Tile_X4Y14_W2BEGb[6] ,
    \Tile_X4Y14_W2BEGb[5] ,
    \Tile_X4Y14_W2BEGb[4] ,
    \Tile_X4Y14_W2BEGb[3] ,
    \Tile_X4Y14_W2BEGb[2] ,
    \Tile_X4Y14_W2BEGb[1] ,
    \Tile_X4Y14_W2BEGb[0] }),
    .W2END({\Tile_X5Y14_W2BEGb[7] ,
    \Tile_X5Y14_W2BEGb[6] ,
    \Tile_X5Y14_W2BEGb[5] ,
    \Tile_X5Y14_W2BEGb[4] ,
    \Tile_X5Y14_W2BEGb[3] ,
    \Tile_X5Y14_W2BEGb[2] ,
    \Tile_X5Y14_W2BEGb[1] ,
    \Tile_X5Y14_W2BEGb[0] }),
    .W2MID({\Tile_X5Y14_W2BEG[7] ,
    \Tile_X5Y14_W2BEG[6] ,
    \Tile_X5Y14_W2BEG[5] ,
    \Tile_X5Y14_W2BEG[4] ,
    \Tile_X5Y14_W2BEG[3] ,
    \Tile_X5Y14_W2BEG[2] ,
    \Tile_X5Y14_W2BEG[1] ,
    \Tile_X5Y14_W2BEG[0] }),
    .W6BEG({\Tile_X4Y14_W6BEG[11] ,
    \Tile_X4Y14_W6BEG[10] ,
    \Tile_X4Y14_W6BEG[9] ,
    \Tile_X4Y14_W6BEG[8] ,
    \Tile_X4Y14_W6BEG[7] ,
    \Tile_X4Y14_W6BEG[6] ,
    \Tile_X4Y14_W6BEG[5] ,
    \Tile_X4Y14_W6BEG[4] ,
    \Tile_X4Y14_W6BEG[3] ,
    \Tile_X4Y14_W6BEG[2] ,
    \Tile_X4Y14_W6BEG[1] ,
    \Tile_X4Y14_W6BEG[0] }),
    .W6END({\Tile_X5Y14_W6BEG[11] ,
    \Tile_X5Y14_W6BEG[10] ,
    \Tile_X5Y14_W6BEG[9] ,
    \Tile_X5Y14_W6BEG[8] ,
    \Tile_X5Y14_W6BEG[7] ,
    \Tile_X5Y14_W6BEG[6] ,
    \Tile_X5Y14_W6BEG[5] ,
    \Tile_X5Y14_W6BEG[4] ,
    \Tile_X5Y14_W6BEG[3] ,
    \Tile_X5Y14_W6BEG[2] ,
    \Tile_X5Y14_W6BEG[1] ,
    \Tile_X5Y14_W6BEG[0] }),
    .WW4BEG({\Tile_X4Y14_WW4BEG[15] ,
    \Tile_X4Y14_WW4BEG[14] ,
    \Tile_X4Y14_WW4BEG[13] ,
    \Tile_X4Y14_WW4BEG[12] ,
    \Tile_X4Y14_WW4BEG[11] ,
    \Tile_X4Y14_WW4BEG[10] ,
    \Tile_X4Y14_WW4BEG[9] ,
    \Tile_X4Y14_WW4BEG[8] ,
    \Tile_X4Y14_WW4BEG[7] ,
    \Tile_X4Y14_WW4BEG[6] ,
    \Tile_X4Y14_WW4BEG[5] ,
    \Tile_X4Y14_WW4BEG[4] ,
    \Tile_X4Y14_WW4BEG[3] ,
    \Tile_X4Y14_WW4BEG[2] ,
    \Tile_X4Y14_WW4BEG[1] ,
    \Tile_X4Y14_WW4BEG[0] }),
    .WW4END({\Tile_X5Y14_WW4BEG[15] ,
    \Tile_X5Y14_WW4BEG[14] ,
    \Tile_X5Y14_WW4BEG[13] ,
    \Tile_X5Y14_WW4BEG[12] ,
    \Tile_X5Y14_WW4BEG[11] ,
    \Tile_X5Y14_WW4BEG[10] ,
    \Tile_X5Y14_WW4BEG[9] ,
    \Tile_X5Y14_WW4BEG[8] ,
    \Tile_X5Y14_WW4BEG[7] ,
    \Tile_X5Y14_WW4BEG[6] ,
    \Tile_X5Y14_WW4BEG[5] ,
    \Tile_X5Y14_WW4BEG[4] ,
    \Tile_X5Y14_WW4BEG[3] ,
    \Tile_X5Y14_WW4BEG[2] ,
    \Tile_X5Y14_WW4BEG[1] ,
    \Tile_X5Y14_WW4BEG[0] }));
 S_term_single2 Tile_X4Y15_S_term_single2 (.UserCLK(UserCLK),
    .UserCLKo(Tile_X4Y15_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .FrameData({\Tile_X3Y15_FrameData_O[31] ,
    \Tile_X3Y15_FrameData_O[30] ,
    \Tile_X3Y15_FrameData_O[29] ,
    \Tile_X3Y15_FrameData_O[28] ,
    \Tile_X3Y15_FrameData_O[27] ,
    \Tile_X3Y15_FrameData_O[26] ,
    \Tile_X3Y15_FrameData_O[25] ,
    \Tile_X3Y15_FrameData_O[24] ,
    \Tile_X3Y15_FrameData_O[23] ,
    \Tile_X3Y15_FrameData_O[22] ,
    \Tile_X3Y15_FrameData_O[21] ,
    \Tile_X3Y15_FrameData_O[20] ,
    \Tile_X3Y15_FrameData_O[19] ,
    \Tile_X3Y15_FrameData_O[18] ,
    \Tile_X3Y15_FrameData_O[17] ,
    \Tile_X3Y15_FrameData_O[16] ,
    \Tile_X3Y15_FrameData_O[15] ,
    \Tile_X3Y15_FrameData_O[14] ,
    \Tile_X3Y15_FrameData_O[13] ,
    \Tile_X3Y15_FrameData_O[12] ,
    \Tile_X3Y15_FrameData_O[11] ,
    \Tile_X3Y15_FrameData_O[10] ,
    \Tile_X3Y15_FrameData_O[9] ,
    \Tile_X3Y15_FrameData_O[8] ,
    \Tile_X3Y15_FrameData_O[7] ,
    \Tile_X3Y15_FrameData_O[6] ,
    \Tile_X3Y15_FrameData_O[5] ,
    \Tile_X3Y15_FrameData_O[4] ,
    \Tile_X3Y15_FrameData_O[3] ,
    \Tile_X3Y15_FrameData_O[2] ,
    \Tile_X3Y15_FrameData_O[1] ,
    \Tile_X3Y15_FrameData_O[0] }),
    .FrameData_O({\Tile_X4Y15_FrameData_O[31] ,
    \Tile_X4Y15_FrameData_O[30] ,
    \Tile_X4Y15_FrameData_O[29] ,
    \Tile_X4Y15_FrameData_O[28] ,
    \Tile_X4Y15_FrameData_O[27] ,
    \Tile_X4Y15_FrameData_O[26] ,
    \Tile_X4Y15_FrameData_O[25] ,
    \Tile_X4Y15_FrameData_O[24] ,
    \Tile_X4Y15_FrameData_O[23] ,
    \Tile_X4Y15_FrameData_O[22] ,
    \Tile_X4Y15_FrameData_O[21] ,
    \Tile_X4Y15_FrameData_O[20] ,
    \Tile_X4Y15_FrameData_O[19] ,
    \Tile_X4Y15_FrameData_O[18] ,
    \Tile_X4Y15_FrameData_O[17] ,
    \Tile_X4Y15_FrameData_O[16] ,
    \Tile_X4Y15_FrameData_O[15] ,
    \Tile_X4Y15_FrameData_O[14] ,
    \Tile_X4Y15_FrameData_O[13] ,
    \Tile_X4Y15_FrameData_O[12] ,
    \Tile_X4Y15_FrameData_O[11] ,
    \Tile_X4Y15_FrameData_O[10] ,
    \Tile_X4Y15_FrameData_O[9] ,
    \Tile_X4Y15_FrameData_O[8] ,
    \Tile_X4Y15_FrameData_O[7] ,
    \Tile_X4Y15_FrameData_O[6] ,
    \Tile_X4Y15_FrameData_O[5] ,
    \Tile_X4Y15_FrameData_O[4] ,
    \Tile_X4Y15_FrameData_O[3] ,
    \Tile_X4Y15_FrameData_O[2] ,
    \Tile_X4Y15_FrameData_O[1] ,
    \Tile_X4Y15_FrameData_O[0] }),
    .FrameStrobe({FrameStrobe[99],
    FrameStrobe[98],
    FrameStrobe[97],
    FrameStrobe[96],
    FrameStrobe[95],
    FrameStrobe[94],
    FrameStrobe[93],
    FrameStrobe[92],
    FrameStrobe[91],
    FrameStrobe[90],
    FrameStrobe[89],
    FrameStrobe[88],
    FrameStrobe[87],
    FrameStrobe[86],
    FrameStrobe[85],
    FrameStrobe[84],
    FrameStrobe[83],
    FrameStrobe[82],
    FrameStrobe[81],
    FrameStrobe[80]}),
    .FrameStrobe_O({\Tile_X4Y15_FrameStrobe_O[19] ,
    \Tile_X4Y15_FrameStrobe_O[18] ,
    \Tile_X4Y15_FrameStrobe_O[17] ,
    \Tile_X4Y15_FrameStrobe_O[16] ,
    \Tile_X4Y15_FrameStrobe_O[15] ,
    \Tile_X4Y15_FrameStrobe_O[14] ,
    \Tile_X4Y15_FrameStrobe_O[13] ,
    \Tile_X4Y15_FrameStrobe_O[12] ,
    \Tile_X4Y15_FrameStrobe_O[11] ,
    \Tile_X4Y15_FrameStrobe_O[10] ,
    \Tile_X4Y15_FrameStrobe_O[9] ,
    \Tile_X4Y15_FrameStrobe_O[8] ,
    \Tile_X4Y15_FrameStrobe_O[7] ,
    \Tile_X4Y15_FrameStrobe_O[6] ,
    \Tile_X4Y15_FrameStrobe_O[5] ,
    \Tile_X4Y15_FrameStrobe_O[4] ,
    \Tile_X4Y15_FrameStrobe_O[3] ,
    \Tile_X4Y15_FrameStrobe_O[2] ,
    \Tile_X4Y15_FrameStrobe_O[1] ,
    \Tile_X4Y15_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X4Y15_N1BEG[3] ,
    \Tile_X4Y15_N1BEG[2] ,
    \Tile_X4Y15_N1BEG[1] ,
    \Tile_X4Y15_N1BEG[0] }),
    .N2BEG({\Tile_X4Y15_N2BEG[7] ,
    \Tile_X4Y15_N2BEG[6] ,
    \Tile_X4Y15_N2BEG[5] ,
    \Tile_X4Y15_N2BEG[4] ,
    \Tile_X4Y15_N2BEG[3] ,
    \Tile_X4Y15_N2BEG[2] ,
    \Tile_X4Y15_N2BEG[1] ,
    \Tile_X4Y15_N2BEG[0] }),
    .N2BEGb({\Tile_X4Y15_N2BEGb[7] ,
    \Tile_X4Y15_N2BEGb[6] ,
    \Tile_X4Y15_N2BEGb[5] ,
    \Tile_X4Y15_N2BEGb[4] ,
    \Tile_X4Y15_N2BEGb[3] ,
    \Tile_X4Y15_N2BEGb[2] ,
    \Tile_X4Y15_N2BEGb[1] ,
    \Tile_X4Y15_N2BEGb[0] }),
    .N4BEG({\Tile_X4Y15_N4BEG[15] ,
    \Tile_X4Y15_N4BEG[14] ,
    \Tile_X4Y15_N4BEG[13] ,
    \Tile_X4Y15_N4BEG[12] ,
    \Tile_X4Y15_N4BEG[11] ,
    \Tile_X4Y15_N4BEG[10] ,
    \Tile_X4Y15_N4BEG[9] ,
    \Tile_X4Y15_N4BEG[8] ,
    \Tile_X4Y15_N4BEG[7] ,
    \Tile_X4Y15_N4BEG[6] ,
    \Tile_X4Y15_N4BEG[5] ,
    \Tile_X4Y15_N4BEG[4] ,
    \Tile_X4Y15_N4BEG[3] ,
    \Tile_X4Y15_N4BEG[2] ,
    \Tile_X4Y15_N4BEG[1] ,
    \Tile_X4Y15_N4BEG[0] }),
    .NN4BEG({\Tile_X4Y15_NN4BEG[15] ,
    \Tile_X4Y15_NN4BEG[14] ,
    \Tile_X4Y15_NN4BEG[13] ,
    \Tile_X4Y15_NN4BEG[12] ,
    \Tile_X4Y15_NN4BEG[11] ,
    \Tile_X4Y15_NN4BEG[10] ,
    \Tile_X4Y15_NN4BEG[9] ,
    \Tile_X4Y15_NN4BEG[8] ,
    \Tile_X4Y15_NN4BEG[7] ,
    \Tile_X4Y15_NN4BEG[6] ,
    \Tile_X4Y15_NN4BEG[5] ,
    \Tile_X4Y15_NN4BEG[4] ,
    \Tile_X4Y15_NN4BEG[3] ,
    \Tile_X4Y15_NN4BEG[2] ,
    \Tile_X4Y15_NN4BEG[1] ,
    \Tile_X4Y15_NN4BEG[0] }),
    .S1END({\Tile_X4Y14_S1BEG[3] ,
    \Tile_X4Y14_S1BEG[2] ,
    \Tile_X4Y14_S1BEG[1] ,
    \Tile_X4Y14_S1BEG[0] }),
    .S2END({\Tile_X4Y14_S2BEGb[7] ,
    \Tile_X4Y14_S2BEGb[6] ,
    \Tile_X4Y14_S2BEGb[5] ,
    \Tile_X4Y14_S2BEGb[4] ,
    \Tile_X4Y14_S2BEGb[3] ,
    \Tile_X4Y14_S2BEGb[2] ,
    \Tile_X4Y14_S2BEGb[1] ,
    \Tile_X4Y14_S2BEGb[0] }),
    .S2MID({\Tile_X4Y14_S2BEG[7] ,
    \Tile_X4Y14_S2BEG[6] ,
    \Tile_X4Y14_S2BEG[5] ,
    \Tile_X4Y14_S2BEG[4] ,
    \Tile_X4Y14_S2BEG[3] ,
    \Tile_X4Y14_S2BEG[2] ,
    \Tile_X4Y14_S2BEG[1] ,
    \Tile_X4Y14_S2BEG[0] }),
    .S4END({\Tile_X4Y14_S4BEG[15] ,
    \Tile_X4Y14_S4BEG[14] ,
    \Tile_X4Y14_S4BEG[13] ,
    \Tile_X4Y14_S4BEG[12] ,
    \Tile_X4Y14_S4BEG[11] ,
    \Tile_X4Y14_S4BEG[10] ,
    \Tile_X4Y14_S4BEG[9] ,
    \Tile_X4Y14_S4BEG[8] ,
    \Tile_X4Y14_S4BEG[7] ,
    \Tile_X4Y14_S4BEG[6] ,
    \Tile_X4Y14_S4BEG[5] ,
    \Tile_X4Y14_S4BEG[4] ,
    \Tile_X4Y14_S4BEG[3] ,
    \Tile_X4Y14_S4BEG[2] ,
    \Tile_X4Y14_S4BEG[1] ,
    \Tile_X4Y14_S4BEG[0] }),
    .SS4END({\Tile_X4Y14_SS4BEG[15] ,
    \Tile_X4Y14_SS4BEG[14] ,
    \Tile_X4Y14_SS4BEG[13] ,
    \Tile_X4Y14_SS4BEG[12] ,
    \Tile_X4Y14_SS4BEG[11] ,
    \Tile_X4Y14_SS4BEG[10] ,
    \Tile_X4Y14_SS4BEG[9] ,
    \Tile_X4Y14_SS4BEG[8] ,
    \Tile_X4Y14_SS4BEG[7] ,
    \Tile_X4Y14_SS4BEG[6] ,
    \Tile_X4Y14_SS4BEG[5] ,
    \Tile_X4Y14_SS4BEG[4] ,
    \Tile_X4Y14_SS4BEG[3] ,
    \Tile_X4Y14_SS4BEG[2] ,
    \Tile_X4Y14_SS4BEG[1] ,
    \Tile_X4Y14_SS4BEG[0] }));
 RegFile Tile_X4Y1_RegFile (.UserCLK(Tile_X4Y2_UserCLKo),
    .UserCLKo(Tile_X4Y1_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X4Y1_E1BEG[3] ,
    \Tile_X4Y1_E1BEG[2] ,
    \Tile_X4Y1_E1BEG[1] ,
    \Tile_X4Y1_E1BEG[0] }),
    .E1END({\Tile_X3Y1_E1BEG[3] ,
    \Tile_X3Y1_E1BEG[2] ,
    \Tile_X3Y1_E1BEG[1] ,
    \Tile_X3Y1_E1BEG[0] }),
    .E2BEG({\Tile_X4Y1_E2BEG[7] ,
    \Tile_X4Y1_E2BEG[6] ,
    \Tile_X4Y1_E2BEG[5] ,
    \Tile_X4Y1_E2BEG[4] ,
    \Tile_X4Y1_E2BEG[3] ,
    \Tile_X4Y1_E2BEG[2] ,
    \Tile_X4Y1_E2BEG[1] ,
    \Tile_X4Y1_E2BEG[0] }),
    .E2BEGb({\Tile_X4Y1_E2BEGb[7] ,
    \Tile_X4Y1_E2BEGb[6] ,
    \Tile_X4Y1_E2BEGb[5] ,
    \Tile_X4Y1_E2BEGb[4] ,
    \Tile_X4Y1_E2BEGb[3] ,
    \Tile_X4Y1_E2BEGb[2] ,
    \Tile_X4Y1_E2BEGb[1] ,
    \Tile_X4Y1_E2BEGb[0] }),
    .E2END({\Tile_X3Y1_E2BEGb[7] ,
    \Tile_X3Y1_E2BEGb[6] ,
    \Tile_X3Y1_E2BEGb[5] ,
    \Tile_X3Y1_E2BEGb[4] ,
    \Tile_X3Y1_E2BEGb[3] ,
    \Tile_X3Y1_E2BEGb[2] ,
    \Tile_X3Y1_E2BEGb[1] ,
    \Tile_X3Y1_E2BEGb[0] }),
    .E2MID({\Tile_X3Y1_E2BEG[7] ,
    \Tile_X3Y1_E2BEG[6] ,
    \Tile_X3Y1_E2BEG[5] ,
    \Tile_X3Y1_E2BEG[4] ,
    \Tile_X3Y1_E2BEG[3] ,
    \Tile_X3Y1_E2BEG[2] ,
    \Tile_X3Y1_E2BEG[1] ,
    \Tile_X3Y1_E2BEG[0] }),
    .E6BEG({\Tile_X4Y1_E6BEG[11] ,
    \Tile_X4Y1_E6BEG[10] ,
    \Tile_X4Y1_E6BEG[9] ,
    \Tile_X4Y1_E6BEG[8] ,
    \Tile_X4Y1_E6BEG[7] ,
    \Tile_X4Y1_E6BEG[6] ,
    \Tile_X4Y1_E6BEG[5] ,
    \Tile_X4Y1_E6BEG[4] ,
    \Tile_X4Y1_E6BEG[3] ,
    \Tile_X4Y1_E6BEG[2] ,
    \Tile_X4Y1_E6BEG[1] ,
    \Tile_X4Y1_E6BEG[0] }),
    .E6END({\Tile_X3Y1_E6BEG[11] ,
    \Tile_X3Y1_E6BEG[10] ,
    \Tile_X3Y1_E6BEG[9] ,
    \Tile_X3Y1_E6BEG[8] ,
    \Tile_X3Y1_E6BEG[7] ,
    \Tile_X3Y1_E6BEG[6] ,
    \Tile_X3Y1_E6BEG[5] ,
    \Tile_X3Y1_E6BEG[4] ,
    \Tile_X3Y1_E6BEG[3] ,
    \Tile_X3Y1_E6BEG[2] ,
    \Tile_X3Y1_E6BEG[1] ,
    \Tile_X3Y1_E6BEG[0] }),
    .EE4BEG({\Tile_X4Y1_EE4BEG[15] ,
    \Tile_X4Y1_EE4BEG[14] ,
    \Tile_X4Y1_EE4BEG[13] ,
    \Tile_X4Y1_EE4BEG[12] ,
    \Tile_X4Y1_EE4BEG[11] ,
    \Tile_X4Y1_EE4BEG[10] ,
    \Tile_X4Y1_EE4BEG[9] ,
    \Tile_X4Y1_EE4BEG[8] ,
    \Tile_X4Y1_EE4BEG[7] ,
    \Tile_X4Y1_EE4BEG[6] ,
    \Tile_X4Y1_EE4BEG[5] ,
    \Tile_X4Y1_EE4BEG[4] ,
    \Tile_X4Y1_EE4BEG[3] ,
    \Tile_X4Y1_EE4BEG[2] ,
    \Tile_X4Y1_EE4BEG[1] ,
    \Tile_X4Y1_EE4BEG[0] }),
    .EE4END({\Tile_X3Y1_EE4BEG[15] ,
    \Tile_X3Y1_EE4BEG[14] ,
    \Tile_X3Y1_EE4BEG[13] ,
    \Tile_X3Y1_EE4BEG[12] ,
    \Tile_X3Y1_EE4BEG[11] ,
    \Tile_X3Y1_EE4BEG[10] ,
    \Tile_X3Y1_EE4BEG[9] ,
    \Tile_X3Y1_EE4BEG[8] ,
    \Tile_X3Y1_EE4BEG[7] ,
    \Tile_X3Y1_EE4BEG[6] ,
    \Tile_X3Y1_EE4BEG[5] ,
    \Tile_X3Y1_EE4BEG[4] ,
    \Tile_X3Y1_EE4BEG[3] ,
    \Tile_X3Y1_EE4BEG[2] ,
    \Tile_X3Y1_EE4BEG[1] ,
    \Tile_X3Y1_EE4BEG[0] }),
    .FrameData({\Tile_X3Y1_FrameData_O[31] ,
    \Tile_X3Y1_FrameData_O[30] ,
    \Tile_X3Y1_FrameData_O[29] ,
    \Tile_X3Y1_FrameData_O[28] ,
    \Tile_X3Y1_FrameData_O[27] ,
    \Tile_X3Y1_FrameData_O[26] ,
    \Tile_X3Y1_FrameData_O[25] ,
    \Tile_X3Y1_FrameData_O[24] ,
    \Tile_X3Y1_FrameData_O[23] ,
    \Tile_X3Y1_FrameData_O[22] ,
    \Tile_X3Y1_FrameData_O[21] ,
    \Tile_X3Y1_FrameData_O[20] ,
    \Tile_X3Y1_FrameData_O[19] ,
    \Tile_X3Y1_FrameData_O[18] ,
    \Tile_X3Y1_FrameData_O[17] ,
    \Tile_X3Y1_FrameData_O[16] ,
    \Tile_X3Y1_FrameData_O[15] ,
    \Tile_X3Y1_FrameData_O[14] ,
    \Tile_X3Y1_FrameData_O[13] ,
    \Tile_X3Y1_FrameData_O[12] ,
    \Tile_X3Y1_FrameData_O[11] ,
    \Tile_X3Y1_FrameData_O[10] ,
    \Tile_X3Y1_FrameData_O[9] ,
    \Tile_X3Y1_FrameData_O[8] ,
    \Tile_X3Y1_FrameData_O[7] ,
    \Tile_X3Y1_FrameData_O[6] ,
    \Tile_X3Y1_FrameData_O[5] ,
    \Tile_X3Y1_FrameData_O[4] ,
    \Tile_X3Y1_FrameData_O[3] ,
    \Tile_X3Y1_FrameData_O[2] ,
    \Tile_X3Y1_FrameData_O[1] ,
    \Tile_X3Y1_FrameData_O[0] }),
    .FrameData_O({\Tile_X4Y1_FrameData_O[31] ,
    \Tile_X4Y1_FrameData_O[30] ,
    \Tile_X4Y1_FrameData_O[29] ,
    \Tile_X4Y1_FrameData_O[28] ,
    \Tile_X4Y1_FrameData_O[27] ,
    \Tile_X4Y1_FrameData_O[26] ,
    \Tile_X4Y1_FrameData_O[25] ,
    \Tile_X4Y1_FrameData_O[24] ,
    \Tile_X4Y1_FrameData_O[23] ,
    \Tile_X4Y1_FrameData_O[22] ,
    \Tile_X4Y1_FrameData_O[21] ,
    \Tile_X4Y1_FrameData_O[20] ,
    \Tile_X4Y1_FrameData_O[19] ,
    \Tile_X4Y1_FrameData_O[18] ,
    \Tile_X4Y1_FrameData_O[17] ,
    \Tile_X4Y1_FrameData_O[16] ,
    \Tile_X4Y1_FrameData_O[15] ,
    \Tile_X4Y1_FrameData_O[14] ,
    \Tile_X4Y1_FrameData_O[13] ,
    \Tile_X4Y1_FrameData_O[12] ,
    \Tile_X4Y1_FrameData_O[11] ,
    \Tile_X4Y1_FrameData_O[10] ,
    \Tile_X4Y1_FrameData_O[9] ,
    \Tile_X4Y1_FrameData_O[8] ,
    \Tile_X4Y1_FrameData_O[7] ,
    \Tile_X4Y1_FrameData_O[6] ,
    \Tile_X4Y1_FrameData_O[5] ,
    \Tile_X4Y1_FrameData_O[4] ,
    \Tile_X4Y1_FrameData_O[3] ,
    \Tile_X4Y1_FrameData_O[2] ,
    \Tile_X4Y1_FrameData_O[1] ,
    \Tile_X4Y1_FrameData_O[0] }),
    .FrameStrobe({\Tile_X4Y2_FrameStrobe_O[19] ,
    \Tile_X4Y2_FrameStrobe_O[18] ,
    \Tile_X4Y2_FrameStrobe_O[17] ,
    \Tile_X4Y2_FrameStrobe_O[16] ,
    \Tile_X4Y2_FrameStrobe_O[15] ,
    \Tile_X4Y2_FrameStrobe_O[14] ,
    \Tile_X4Y2_FrameStrobe_O[13] ,
    \Tile_X4Y2_FrameStrobe_O[12] ,
    \Tile_X4Y2_FrameStrobe_O[11] ,
    \Tile_X4Y2_FrameStrobe_O[10] ,
    \Tile_X4Y2_FrameStrobe_O[9] ,
    \Tile_X4Y2_FrameStrobe_O[8] ,
    \Tile_X4Y2_FrameStrobe_O[7] ,
    \Tile_X4Y2_FrameStrobe_O[6] ,
    \Tile_X4Y2_FrameStrobe_O[5] ,
    \Tile_X4Y2_FrameStrobe_O[4] ,
    \Tile_X4Y2_FrameStrobe_O[3] ,
    \Tile_X4Y2_FrameStrobe_O[2] ,
    \Tile_X4Y2_FrameStrobe_O[1] ,
    \Tile_X4Y2_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X4Y1_FrameStrobe_O[19] ,
    \Tile_X4Y1_FrameStrobe_O[18] ,
    \Tile_X4Y1_FrameStrobe_O[17] ,
    \Tile_X4Y1_FrameStrobe_O[16] ,
    \Tile_X4Y1_FrameStrobe_O[15] ,
    \Tile_X4Y1_FrameStrobe_O[14] ,
    \Tile_X4Y1_FrameStrobe_O[13] ,
    \Tile_X4Y1_FrameStrobe_O[12] ,
    \Tile_X4Y1_FrameStrobe_O[11] ,
    \Tile_X4Y1_FrameStrobe_O[10] ,
    \Tile_X4Y1_FrameStrobe_O[9] ,
    \Tile_X4Y1_FrameStrobe_O[8] ,
    \Tile_X4Y1_FrameStrobe_O[7] ,
    \Tile_X4Y1_FrameStrobe_O[6] ,
    \Tile_X4Y1_FrameStrobe_O[5] ,
    \Tile_X4Y1_FrameStrobe_O[4] ,
    \Tile_X4Y1_FrameStrobe_O[3] ,
    \Tile_X4Y1_FrameStrobe_O[2] ,
    \Tile_X4Y1_FrameStrobe_O[1] ,
    \Tile_X4Y1_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X4Y1_N1BEG[3] ,
    \Tile_X4Y1_N1BEG[2] ,
    \Tile_X4Y1_N1BEG[1] ,
    \Tile_X4Y1_N1BEG[0] }),
    .N1END({\Tile_X4Y2_N1BEG[3] ,
    \Tile_X4Y2_N1BEG[2] ,
    \Tile_X4Y2_N1BEG[1] ,
    \Tile_X4Y2_N1BEG[0] }),
    .N2BEG({\Tile_X4Y1_N2BEG[7] ,
    \Tile_X4Y1_N2BEG[6] ,
    \Tile_X4Y1_N2BEG[5] ,
    \Tile_X4Y1_N2BEG[4] ,
    \Tile_X4Y1_N2BEG[3] ,
    \Tile_X4Y1_N2BEG[2] ,
    \Tile_X4Y1_N2BEG[1] ,
    \Tile_X4Y1_N2BEG[0] }),
    .N2BEGb({\Tile_X4Y1_N2BEGb[7] ,
    \Tile_X4Y1_N2BEGb[6] ,
    \Tile_X4Y1_N2BEGb[5] ,
    \Tile_X4Y1_N2BEGb[4] ,
    \Tile_X4Y1_N2BEGb[3] ,
    \Tile_X4Y1_N2BEGb[2] ,
    \Tile_X4Y1_N2BEGb[1] ,
    \Tile_X4Y1_N2BEGb[0] }),
    .N2END({\Tile_X4Y2_N2BEGb[7] ,
    \Tile_X4Y2_N2BEGb[6] ,
    \Tile_X4Y2_N2BEGb[5] ,
    \Tile_X4Y2_N2BEGb[4] ,
    \Tile_X4Y2_N2BEGb[3] ,
    \Tile_X4Y2_N2BEGb[2] ,
    \Tile_X4Y2_N2BEGb[1] ,
    \Tile_X4Y2_N2BEGb[0] }),
    .N2MID({\Tile_X4Y2_N2BEG[7] ,
    \Tile_X4Y2_N2BEG[6] ,
    \Tile_X4Y2_N2BEG[5] ,
    \Tile_X4Y2_N2BEG[4] ,
    \Tile_X4Y2_N2BEG[3] ,
    \Tile_X4Y2_N2BEG[2] ,
    \Tile_X4Y2_N2BEG[1] ,
    \Tile_X4Y2_N2BEG[0] }),
    .N4BEG({\Tile_X4Y1_N4BEG[15] ,
    \Tile_X4Y1_N4BEG[14] ,
    \Tile_X4Y1_N4BEG[13] ,
    \Tile_X4Y1_N4BEG[12] ,
    \Tile_X4Y1_N4BEG[11] ,
    \Tile_X4Y1_N4BEG[10] ,
    \Tile_X4Y1_N4BEG[9] ,
    \Tile_X4Y1_N4BEG[8] ,
    \Tile_X4Y1_N4BEG[7] ,
    \Tile_X4Y1_N4BEG[6] ,
    \Tile_X4Y1_N4BEG[5] ,
    \Tile_X4Y1_N4BEG[4] ,
    \Tile_X4Y1_N4BEG[3] ,
    \Tile_X4Y1_N4BEG[2] ,
    \Tile_X4Y1_N4BEG[1] ,
    \Tile_X4Y1_N4BEG[0] }),
    .N4END({\Tile_X4Y2_N4BEG[15] ,
    \Tile_X4Y2_N4BEG[14] ,
    \Tile_X4Y2_N4BEG[13] ,
    \Tile_X4Y2_N4BEG[12] ,
    \Tile_X4Y2_N4BEG[11] ,
    \Tile_X4Y2_N4BEG[10] ,
    \Tile_X4Y2_N4BEG[9] ,
    \Tile_X4Y2_N4BEG[8] ,
    \Tile_X4Y2_N4BEG[7] ,
    \Tile_X4Y2_N4BEG[6] ,
    \Tile_X4Y2_N4BEG[5] ,
    \Tile_X4Y2_N4BEG[4] ,
    \Tile_X4Y2_N4BEG[3] ,
    \Tile_X4Y2_N4BEG[2] ,
    \Tile_X4Y2_N4BEG[1] ,
    \Tile_X4Y2_N4BEG[0] }),
    .NN4BEG({\Tile_X4Y1_NN4BEG[15] ,
    \Tile_X4Y1_NN4BEG[14] ,
    \Tile_X4Y1_NN4BEG[13] ,
    \Tile_X4Y1_NN4BEG[12] ,
    \Tile_X4Y1_NN4BEG[11] ,
    \Tile_X4Y1_NN4BEG[10] ,
    \Tile_X4Y1_NN4BEG[9] ,
    \Tile_X4Y1_NN4BEG[8] ,
    \Tile_X4Y1_NN4BEG[7] ,
    \Tile_X4Y1_NN4BEG[6] ,
    \Tile_X4Y1_NN4BEG[5] ,
    \Tile_X4Y1_NN4BEG[4] ,
    \Tile_X4Y1_NN4BEG[3] ,
    \Tile_X4Y1_NN4BEG[2] ,
    \Tile_X4Y1_NN4BEG[1] ,
    \Tile_X4Y1_NN4BEG[0] }),
    .NN4END({\Tile_X4Y2_NN4BEG[15] ,
    \Tile_X4Y2_NN4BEG[14] ,
    \Tile_X4Y2_NN4BEG[13] ,
    \Tile_X4Y2_NN4BEG[12] ,
    \Tile_X4Y2_NN4BEG[11] ,
    \Tile_X4Y2_NN4BEG[10] ,
    \Tile_X4Y2_NN4BEG[9] ,
    \Tile_X4Y2_NN4BEG[8] ,
    \Tile_X4Y2_NN4BEG[7] ,
    \Tile_X4Y2_NN4BEG[6] ,
    \Tile_X4Y2_NN4BEG[5] ,
    \Tile_X4Y2_NN4BEG[4] ,
    \Tile_X4Y2_NN4BEG[3] ,
    \Tile_X4Y2_NN4BEG[2] ,
    \Tile_X4Y2_NN4BEG[1] ,
    \Tile_X4Y2_NN4BEG[0] }),
    .S1BEG({\Tile_X4Y1_S1BEG[3] ,
    \Tile_X4Y1_S1BEG[2] ,
    \Tile_X4Y1_S1BEG[1] ,
    \Tile_X4Y1_S1BEG[0] }),
    .S1END({\Tile_X4Y0_S1BEG[3] ,
    \Tile_X4Y0_S1BEG[2] ,
    \Tile_X4Y0_S1BEG[1] ,
    \Tile_X4Y0_S1BEG[0] }),
    .S2BEG({\Tile_X4Y1_S2BEG[7] ,
    \Tile_X4Y1_S2BEG[6] ,
    \Tile_X4Y1_S2BEG[5] ,
    \Tile_X4Y1_S2BEG[4] ,
    \Tile_X4Y1_S2BEG[3] ,
    \Tile_X4Y1_S2BEG[2] ,
    \Tile_X4Y1_S2BEG[1] ,
    \Tile_X4Y1_S2BEG[0] }),
    .S2BEGb({\Tile_X4Y1_S2BEGb[7] ,
    \Tile_X4Y1_S2BEGb[6] ,
    \Tile_X4Y1_S2BEGb[5] ,
    \Tile_X4Y1_S2BEGb[4] ,
    \Tile_X4Y1_S2BEGb[3] ,
    \Tile_X4Y1_S2BEGb[2] ,
    \Tile_X4Y1_S2BEGb[1] ,
    \Tile_X4Y1_S2BEGb[0] }),
    .S2END({\Tile_X4Y0_S2BEGb[7] ,
    \Tile_X4Y0_S2BEGb[6] ,
    \Tile_X4Y0_S2BEGb[5] ,
    \Tile_X4Y0_S2BEGb[4] ,
    \Tile_X4Y0_S2BEGb[3] ,
    \Tile_X4Y0_S2BEGb[2] ,
    \Tile_X4Y0_S2BEGb[1] ,
    \Tile_X4Y0_S2BEGb[0] }),
    .S2MID({\Tile_X4Y0_S2BEG[7] ,
    \Tile_X4Y0_S2BEG[6] ,
    \Tile_X4Y0_S2BEG[5] ,
    \Tile_X4Y0_S2BEG[4] ,
    \Tile_X4Y0_S2BEG[3] ,
    \Tile_X4Y0_S2BEG[2] ,
    \Tile_X4Y0_S2BEG[1] ,
    \Tile_X4Y0_S2BEG[0] }),
    .S4BEG({\Tile_X4Y1_S4BEG[15] ,
    \Tile_X4Y1_S4BEG[14] ,
    \Tile_X4Y1_S4BEG[13] ,
    \Tile_X4Y1_S4BEG[12] ,
    \Tile_X4Y1_S4BEG[11] ,
    \Tile_X4Y1_S4BEG[10] ,
    \Tile_X4Y1_S4BEG[9] ,
    \Tile_X4Y1_S4BEG[8] ,
    \Tile_X4Y1_S4BEG[7] ,
    \Tile_X4Y1_S4BEG[6] ,
    \Tile_X4Y1_S4BEG[5] ,
    \Tile_X4Y1_S4BEG[4] ,
    \Tile_X4Y1_S4BEG[3] ,
    \Tile_X4Y1_S4BEG[2] ,
    \Tile_X4Y1_S4BEG[1] ,
    \Tile_X4Y1_S4BEG[0] }),
    .S4END({\Tile_X4Y0_S4BEG[15] ,
    \Tile_X4Y0_S4BEG[14] ,
    \Tile_X4Y0_S4BEG[13] ,
    \Tile_X4Y0_S4BEG[12] ,
    \Tile_X4Y0_S4BEG[11] ,
    \Tile_X4Y0_S4BEG[10] ,
    \Tile_X4Y0_S4BEG[9] ,
    \Tile_X4Y0_S4BEG[8] ,
    \Tile_X4Y0_S4BEG[7] ,
    \Tile_X4Y0_S4BEG[6] ,
    \Tile_X4Y0_S4BEG[5] ,
    \Tile_X4Y0_S4BEG[4] ,
    \Tile_X4Y0_S4BEG[3] ,
    \Tile_X4Y0_S4BEG[2] ,
    \Tile_X4Y0_S4BEG[1] ,
    \Tile_X4Y0_S4BEG[0] }),
    .SS4BEG({\Tile_X4Y1_SS4BEG[15] ,
    \Tile_X4Y1_SS4BEG[14] ,
    \Tile_X4Y1_SS4BEG[13] ,
    \Tile_X4Y1_SS4BEG[12] ,
    \Tile_X4Y1_SS4BEG[11] ,
    \Tile_X4Y1_SS4BEG[10] ,
    \Tile_X4Y1_SS4BEG[9] ,
    \Tile_X4Y1_SS4BEG[8] ,
    \Tile_X4Y1_SS4BEG[7] ,
    \Tile_X4Y1_SS4BEG[6] ,
    \Tile_X4Y1_SS4BEG[5] ,
    \Tile_X4Y1_SS4BEG[4] ,
    \Tile_X4Y1_SS4BEG[3] ,
    \Tile_X4Y1_SS4BEG[2] ,
    \Tile_X4Y1_SS4BEG[1] ,
    \Tile_X4Y1_SS4BEG[0] }),
    .SS4END({\Tile_X4Y0_SS4BEG[15] ,
    \Tile_X4Y0_SS4BEG[14] ,
    \Tile_X4Y0_SS4BEG[13] ,
    \Tile_X4Y0_SS4BEG[12] ,
    \Tile_X4Y0_SS4BEG[11] ,
    \Tile_X4Y0_SS4BEG[10] ,
    \Tile_X4Y0_SS4BEG[9] ,
    \Tile_X4Y0_SS4BEG[8] ,
    \Tile_X4Y0_SS4BEG[7] ,
    \Tile_X4Y0_SS4BEG[6] ,
    \Tile_X4Y0_SS4BEG[5] ,
    \Tile_X4Y0_SS4BEG[4] ,
    \Tile_X4Y0_SS4BEG[3] ,
    \Tile_X4Y0_SS4BEG[2] ,
    \Tile_X4Y0_SS4BEG[1] ,
    \Tile_X4Y0_SS4BEG[0] }),
    .W1BEG({\Tile_X4Y1_W1BEG[3] ,
    \Tile_X4Y1_W1BEG[2] ,
    \Tile_X4Y1_W1BEG[1] ,
    \Tile_X4Y1_W1BEG[0] }),
    .W1END({\Tile_X5Y1_W1BEG[3] ,
    \Tile_X5Y1_W1BEG[2] ,
    \Tile_X5Y1_W1BEG[1] ,
    \Tile_X5Y1_W1BEG[0] }),
    .W2BEG({\Tile_X4Y1_W2BEG[7] ,
    \Tile_X4Y1_W2BEG[6] ,
    \Tile_X4Y1_W2BEG[5] ,
    \Tile_X4Y1_W2BEG[4] ,
    \Tile_X4Y1_W2BEG[3] ,
    \Tile_X4Y1_W2BEG[2] ,
    \Tile_X4Y1_W2BEG[1] ,
    \Tile_X4Y1_W2BEG[0] }),
    .W2BEGb({\Tile_X4Y1_W2BEGb[7] ,
    \Tile_X4Y1_W2BEGb[6] ,
    \Tile_X4Y1_W2BEGb[5] ,
    \Tile_X4Y1_W2BEGb[4] ,
    \Tile_X4Y1_W2BEGb[3] ,
    \Tile_X4Y1_W2BEGb[2] ,
    \Tile_X4Y1_W2BEGb[1] ,
    \Tile_X4Y1_W2BEGb[0] }),
    .W2END({\Tile_X5Y1_W2BEGb[7] ,
    \Tile_X5Y1_W2BEGb[6] ,
    \Tile_X5Y1_W2BEGb[5] ,
    \Tile_X5Y1_W2BEGb[4] ,
    \Tile_X5Y1_W2BEGb[3] ,
    \Tile_X5Y1_W2BEGb[2] ,
    \Tile_X5Y1_W2BEGb[1] ,
    \Tile_X5Y1_W2BEGb[0] }),
    .W2MID({\Tile_X5Y1_W2BEG[7] ,
    \Tile_X5Y1_W2BEG[6] ,
    \Tile_X5Y1_W2BEG[5] ,
    \Tile_X5Y1_W2BEG[4] ,
    \Tile_X5Y1_W2BEG[3] ,
    \Tile_X5Y1_W2BEG[2] ,
    \Tile_X5Y1_W2BEG[1] ,
    \Tile_X5Y1_W2BEG[0] }),
    .W6BEG({\Tile_X4Y1_W6BEG[11] ,
    \Tile_X4Y1_W6BEG[10] ,
    \Tile_X4Y1_W6BEG[9] ,
    \Tile_X4Y1_W6BEG[8] ,
    \Tile_X4Y1_W6BEG[7] ,
    \Tile_X4Y1_W6BEG[6] ,
    \Tile_X4Y1_W6BEG[5] ,
    \Tile_X4Y1_W6BEG[4] ,
    \Tile_X4Y1_W6BEG[3] ,
    \Tile_X4Y1_W6BEG[2] ,
    \Tile_X4Y1_W6BEG[1] ,
    \Tile_X4Y1_W6BEG[0] }),
    .W6END({\Tile_X5Y1_W6BEG[11] ,
    \Tile_X5Y1_W6BEG[10] ,
    \Tile_X5Y1_W6BEG[9] ,
    \Tile_X5Y1_W6BEG[8] ,
    \Tile_X5Y1_W6BEG[7] ,
    \Tile_X5Y1_W6BEG[6] ,
    \Tile_X5Y1_W6BEG[5] ,
    \Tile_X5Y1_W6BEG[4] ,
    \Tile_X5Y1_W6BEG[3] ,
    \Tile_X5Y1_W6BEG[2] ,
    \Tile_X5Y1_W6BEG[1] ,
    \Tile_X5Y1_W6BEG[0] }),
    .WW4BEG({\Tile_X4Y1_WW4BEG[15] ,
    \Tile_X4Y1_WW4BEG[14] ,
    \Tile_X4Y1_WW4BEG[13] ,
    \Tile_X4Y1_WW4BEG[12] ,
    \Tile_X4Y1_WW4BEG[11] ,
    \Tile_X4Y1_WW4BEG[10] ,
    \Tile_X4Y1_WW4BEG[9] ,
    \Tile_X4Y1_WW4BEG[8] ,
    \Tile_X4Y1_WW4BEG[7] ,
    \Tile_X4Y1_WW4BEG[6] ,
    \Tile_X4Y1_WW4BEG[5] ,
    \Tile_X4Y1_WW4BEG[4] ,
    \Tile_X4Y1_WW4BEG[3] ,
    \Tile_X4Y1_WW4BEG[2] ,
    \Tile_X4Y1_WW4BEG[1] ,
    \Tile_X4Y1_WW4BEG[0] }),
    .WW4END({\Tile_X5Y1_WW4BEG[15] ,
    \Tile_X5Y1_WW4BEG[14] ,
    \Tile_X5Y1_WW4BEG[13] ,
    \Tile_X5Y1_WW4BEG[12] ,
    \Tile_X5Y1_WW4BEG[11] ,
    \Tile_X5Y1_WW4BEG[10] ,
    \Tile_X5Y1_WW4BEG[9] ,
    \Tile_X5Y1_WW4BEG[8] ,
    \Tile_X5Y1_WW4BEG[7] ,
    \Tile_X5Y1_WW4BEG[6] ,
    \Tile_X5Y1_WW4BEG[5] ,
    \Tile_X5Y1_WW4BEG[4] ,
    \Tile_X5Y1_WW4BEG[3] ,
    \Tile_X5Y1_WW4BEG[2] ,
    \Tile_X5Y1_WW4BEG[1] ,
    \Tile_X5Y1_WW4BEG[0] }));
 RegFile Tile_X4Y2_RegFile (.UserCLK(Tile_X4Y3_UserCLKo),
    .UserCLKo(Tile_X4Y2_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X4Y2_E1BEG[3] ,
    \Tile_X4Y2_E1BEG[2] ,
    \Tile_X4Y2_E1BEG[1] ,
    \Tile_X4Y2_E1BEG[0] }),
    .E1END({\Tile_X3Y2_E1BEG[3] ,
    \Tile_X3Y2_E1BEG[2] ,
    \Tile_X3Y2_E1BEG[1] ,
    \Tile_X3Y2_E1BEG[0] }),
    .E2BEG({\Tile_X4Y2_E2BEG[7] ,
    \Tile_X4Y2_E2BEG[6] ,
    \Tile_X4Y2_E2BEG[5] ,
    \Tile_X4Y2_E2BEG[4] ,
    \Tile_X4Y2_E2BEG[3] ,
    \Tile_X4Y2_E2BEG[2] ,
    \Tile_X4Y2_E2BEG[1] ,
    \Tile_X4Y2_E2BEG[0] }),
    .E2BEGb({\Tile_X4Y2_E2BEGb[7] ,
    \Tile_X4Y2_E2BEGb[6] ,
    \Tile_X4Y2_E2BEGb[5] ,
    \Tile_X4Y2_E2BEGb[4] ,
    \Tile_X4Y2_E2BEGb[3] ,
    \Tile_X4Y2_E2BEGb[2] ,
    \Tile_X4Y2_E2BEGb[1] ,
    \Tile_X4Y2_E2BEGb[0] }),
    .E2END({\Tile_X3Y2_E2BEGb[7] ,
    \Tile_X3Y2_E2BEGb[6] ,
    \Tile_X3Y2_E2BEGb[5] ,
    \Tile_X3Y2_E2BEGb[4] ,
    \Tile_X3Y2_E2BEGb[3] ,
    \Tile_X3Y2_E2BEGb[2] ,
    \Tile_X3Y2_E2BEGb[1] ,
    \Tile_X3Y2_E2BEGb[0] }),
    .E2MID({\Tile_X3Y2_E2BEG[7] ,
    \Tile_X3Y2_E2BEG[6] ,
    \Tile_X3Y2_E2BEG[5] ,
    \Tile_X3Y2_E2BEG[4] ,
    \Tile_X3Y2_E2BEG[3] ,
    \Tile_X3Y2_E2BEG[2] ,
    \Tile_X3Y2_E2BEG[1] ,
    \Tile_X3Y2_E2BEG[0] }),
    .E6BEG({\Tile_X4Y2_E6BEG[11] ,
    \Tile_X4Y2_E6BEG[10] ,
    \Tile_X4Y2_E6BEG[9] ,
    \Tile_X4Y2_E6BEG[8] ,
    \Tile_X4Y2_E6BEG[7] ,
    \Tile_X4Y2_E6BEG[6] ,
    \Tile_X4Y2_E6BEG[5] ,
    \Tile_X4Y2_E6BEG[4] ,
    \Tile_X4Y2_E6BEG[3] ,
    \Tile_X4Y2_E6BEG[2] ,
    \Tile_X4Y2_E6BEG[1] ,
    \Tile_X4Y2_E6BEG[0] }),
    .E6END({\Tile_X3Y2_E6BEG[11] ,
    \Tile_X3Y2_E6BEG[10] ,
    \Tile_X3Y2_E6BEG[9] ,
    \Tile_X3Y2_E6BEG[8] ,
    \Tile_X3Y2_E6BEG[7] ,
    \Tile_X3Y2_E6BEG[6] ,
    \Tile_X3Y2_E6BEG[5] ,
    \Tile_X3Y2_E6BEG[4] ,
    \Tile_X3Y2_E6BEG[3] ,
    \Tile_X3Y2_E6BEG[2] ,
    \Tile_X3Y2_E6BEG[1] ,
    \Tile_X3Y2_E6BEG[0] }),
    .EE4BEG({\Tile_X4Y2_EE4BEG[15] ,
    \Tile_X4Y2_EE4BEG[14] ,
    \Tile_X4Y2_EE4BEG[13] ,
    \Tile_X4Y2_EE4BEG[12] ,
    \Tile_X4Y2_EE4BEG[11] ,
    \Tile_X4Y2_EE4BEG[10] ,
    \Tile_X4Y2_EE4BEG[9] ,
    \Tile_X4Y2_EE4BEG[8] ,
    \Tile_X4Y2_EE4BEG[7] ,
    \Tile_X4Y2_EE4BEG[6] ,
    \Tile_X4Y2_EE4BEG[5] ,
    \Tile_X4Y2_EE4BEG[4] ,
    \Tile_X4Y2_EE4BEG[3] ,
    \Tile_X4Y2_EE4BEG[2] ,
    \Tile_X4Y2_EE4BEG[1] ,
    \Tile_X4Y2_EE4BEG[0] }),
    .EE4END({\Tile_X3Y2_EE4BEG[15] ,
    \Tile_X3Y2_EE4BEG[14] ,
    \Tile_X3Y2_EE4BEG[13] ,
    \Tile_X3Y2_EE4BEG[12] ,
    \Tile_X3Y2_EE4BEG[11] ,
    \Tile_X3Y2_EE4BEG[10] ,
    \Tile_X3Y2_EE4BEG[9] ,
    \Tile_X3Y2_EE4BEG[8] ,
    \Tile_X3Y2_EE4BEG[7] ,
    \Tile_X3Y2_EE4BEG[6] ,
    \Tile_X3Y2_EE4BEG[5] ,
    \Tile_X3Y2_EE4BEG[4] ,
    \Tile_X3Y2_EE4BEG[3] ,
    \Tile_X3Y2_EE4BEG[2] ,
    \Tile_X3Y2_EE4BEG[1] ,
    \Tile_X3Y2_EE4BEG[0] }),
    .FrameData({\Tile_X3Y2_FrameData_O[31] ,
    \Tile_X3Y2_FrameData_O[30] ,
    \Tile_X3Y2_FrameData_O[29] ,
    \Tile_X3Y2_FrameData_O[28] ,
    \Tile_X3Y2_FrameData_O[27] ,
    \Tile_X3Y2_FrameData_O[26] ,
    \Tile_X3Y2_FrameData_O[25] ,
    \Tile_X3Y2_FrameData_O[24] ,
    \Tile_X3Y2_FrameData_O[23] ,
    \Tile_X3Y2_FrameData_O[22] ,
    \Tile_X3Y2_FrameData_O[21] ,
    \Tile_X3Y2_FrameData_O[20] ,
    \Tile_X3Y2_FrameData_O[19] ,
    \Tile_X3Y2_FrameData_O[18] ,
    \Tile_X3Y2_FrameData_O[17] ,
    \Tile_X3Y2_FrameData_O[16] ,
    \Tile_X3Y2_FrameData_O[15] ,
    \Tile_X3Y2_FrameData_O[14] ,
    \Tile_X3Y2_FrameData_O[13] ,
    \Tile_X3Y2_FrameData_O[12] ,
    \Tile_X3Y2_FrameData_O[11] ,
    \Tile_X3Y2_FrameData_O[10] ,
    \Tile_X3Y2_FrameData_O[9] ,
    \Tile_X3Y2_FrameData_O[8] ,
    \Tile_X3Y2_FrameData_O[7] ,
    \Tile_X3Y2_FrameData_O[6] ,
    \Tile_X3Y2_FrameData_O[5] ,
    \Tile_X3Y2_FrameData_O[4] ,
    \Tile_X3Y2_FrameData_O[3] ,
    \Tile_X3Y2_FrameData_O[2] ,
    \Tile_X3Y2_FrameData_O[1] ,
    \Tile_X3Y2_FrameData_O[0] }),
    .FrameData_O({\Tile_X4Y2_FrameData_O[31] ,
    \Tile_X4Y2_FrameData_O[30] ,
    \Tile_X4Y2_FrameData_O[29] ,
    \Tile_X4Y2_FrameData_O[28] ,
    \Tile_X4Y2_FrameData_O[27] ,
    \Tile_X4Y2_FrameData_O[26] ,
    \Tile_X4Y2_FrameData_O[25] ,
    \Tile_X4Y2_FrameData_O[24] ,
    \Tile_X4Y2_FrameData_O[23] ,
    \Tile_X4Y2_FrameData_O[22] ,
    \Tile_X4Y2_FrameData_O[21] ,
    \Tile_X4Y2_FrameData_O[20] ,
    \Tile_X4Y2_FrameData_O[19] ,
    \Tile_X4Y2_FrameData_O[18] ,
    \Tile_X4Y2_FrameData_O[17] ,
    \Tile_X4Y2_FrameData_O[16] ,
    \Tile_X4Y2_FrameData_O[15] ,
    \Tile_X4Y2_FrameData_O[14] ,
    \Tile_X4Y2_FrameData_O[13] ,
    \Tile_X4Y2_FrameData_O[12] ,
    \Tile_X4Y2_FrameData_O[11] ,
    \Tile_X4Y2_FrameData_O[10] ,
    \Tile_X4Y2_FrameData_O[9] ,
    \Tile_X4Y2_FrameData_O[8] ,
    \Tile_X4Y2_FrameData_O[7] ,
    \Tile_X4Y2_FrameData_O[6] ,
    \Tile_X4Y2_FrameData_O[5] ,
    \Tile_X4Y2_FrameData_O[4] ,
    \Tile_X4Y2_FrameData_O[3] ,
    \Tile_X4Y2_FrameData_O[2] ,
    \Tile_X4Y2_FrameData_O[1] ,
    \Tile_X4Y2_FrameData_O[0] }),
    .FrameStrobe({\Tile_X4Y3_FrameStrobe_O[19] ,
    \Tile_X4Y3_FrameStrobe_O[18] ,
    \Tile_X4Y3_FrameStrobe_O[17] ,
    \Tile_X4Y3_FrameStrobe_O[16] ,
    \Tile_X4Y3_FrameStrobe_O[15] ,
    \Tile_X4Y3_FrameStrobe_O[14] ,
    \Tile_X4Y3_FrameStrobe_O[13] ,
    \Tile_X4Y3_FrameStrobe_O[12] ,
    \Tile_X4Y3_FrameStrobe_O[11] ,
    \Tile_X4Y3_FrameStrobe_O[10] ,
    \Tile_X4Y3_FrameStrobe_O[9] ,
    \Tile_X4Y3_FrameStrobe_O[8] ,
    \Tile_X4Y3_FrameStrobe_O[7] ,
    \Tile_X4Y3_FrameStrobe_O[6] ,
    \Tile_X4Y3_FrameStrobe_O[5] ,
    \Tile_X4Y3_FrameStrobe_O[4] ,
    \Tile_X4Y3_FrameStrobe_O[3] ,
    \Tile_X4Y3_FrameStrobe_O[2] ,
    \Tile_X4Y3_FrameStrobe_O[1] ,
    \Tile_X4Y3_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X4Y2_FrameStrobe_O[19] ,
    \Tile_X4Y2_FrameStrobe_O[18] ,
    \Tile_X4Y2_FrameStrobe_O[17] ,
    \Tile_X4Y2_FrameStrobe_O[16] ,
    \Tile_X4Y2_FrameStrobe_O[15] ,
    \Tile_X4Y2_FrameStrobe_O[14] ,
    \Tile_X4Y2_FrameStrobe_O[13] ,
    \Tile_X4Y2_FrameStrobe_O[12] ,
    \Tile_X4Y2_FrameStrobe_O[11] ,
    \Tile_X4Y2_FrameStrobe_O[10] ,
    \Tile_X4Y2_FrameStrobe_O[9] ,
    \Tile_X4Y2_FrameStrobe_O[8] ,
    \Tile_X4Y2_FrameStrobe_O[7] ,
    \Tile_X4Y2_FrameStrobe_O[6] ,
    \Tile_X4Y2_FrameStrobe_O[5] ,
    \Tile_X4Y2_FrameStrobe_O[4] ,
    \Tile_X4Y2_FrameStrobe_O[3] ,
    \Tile_X4Y2_FrameStrobe_O[2] ,
    \Tile_X4Y2_FrameStrobe_O[1] ,
    \Tile_X4Y2_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X4Y2_N1BEG[3] ,
    \Tile_X4Y2_N1BEG[2] ,
    \Tile_X4Y2_N1BEG[1] ,
    \Tile_X4Y2_N1BEG[0] }),
    .N1END({\Tile_X4Y3_N1BEG[3] ,
    \Tile_X4Y3_N1BEG[2] ,
    \Tile_X4Y3_N1BEG[1] ,
    \Tile_X4Y3_N1BEG[0] }),
    .N2BEG({\Tile_X4Y2_N2BEG[7] ,
    \Tile_X4Y2_N2BEG[6] ,
    \Tile_X4Y2_N2BEG[5] ,
    \Tile_X4Y2_N2BEG[4] ,
    \Tile_X4Y2_N2BEG[3] ,
    \Tile_X4Y2_N2BEG[2] ,
    \Tile_X4Y2_N2BEG[1] ,
    \Tile_X4Y2_N2BEG[0] }),
    .N2BEGb({\Tile_X4Y2_N2BEGb[7] ,
    \Tile_X4Y2_N2BEGb[6] ,
    \Tile_X4Y2_N2BEGb[5] ,
    \Tile_X4Y2_N2BEGb[4] ,
    \Tile_X4Y2_N2BEGb[3] ,
    \Tile_X4Y2_N2BEGb[2] ,
    \Tile_X4Y2_N2BEGb[1] ,
    \Tile_X4Y2_N2BEGb[0] }),
    .N2END({\Tile_X4Y3_N2BEGb[7] ,
    \Tile_X4Y3_N2BEGb[6] ,
    \Tile_X4Y3_N2BEGb[5] ,
    \Tile_X4Y3_N2BEGb[4] ,
    \Tile_X4Y3_N2BEGb[3] ,
    \Tile_X4Y3_N2BEGb[2] ,
    \Tile_X4Y3_N2BEGb[1] ,
    \Tile_X4Y3_N2BEGb[0] }),
    .N2MID({\Tile_X4Y3_N2BEG[7] ,
    \Tile_X4Y3_N2BEG[6] ,
    \Tile_X4Y3_N2BEG[5] ,
    \Tile_X4Y3_N2BEG[4] ,
    \Tile_X4Y3_N2BEG[3] ,
    \Tile_X4Y3_N2BEG[2] ,
    \Tile_X4Y3_N2BEG[1] ,
    \Tile_X4Y3_N2BEG[0] }),
    .N4BEG({\Tile_X4Y2_N4BEG[15] ,
    \Tile_X4Y2_N4BEG[14] ,
    \Tile_X4Y2_N4BEG[13] ,
    \Tile_X4Y2_N4BEG[12] ,
    \Tile_X4Y2_N4BEG[11] ,
    \Tile_X4Y2_N4BEG[10] ,
    \Tile_X4Y2_N4BEG[9] ,
    \Tile_X4Y2_N4BEG[8] ,
    \Tile_X4Y2_N4BEG[7] ,
    \Tile_X4Y2_N4BEG[6] ,
    \Tile_X4Y2_N4BEG[5] ,
    \Tile_X4Y2_N4BEG[4] ,
    \Tile_X4Y2_N4BEG[3] ,
    \Tile_X4Y2_N4BEG[2] ,
    \Tile_X4Y2_N4BEG[1] ,
    \Tile_X4Y2_N4BEG[0] }),
    .N4END({\Tile_X4Y3_N4BEG[15] ,
    \Tile_X4Y3_N4BEG[14] ,
    \Tile_X4Y3_N4BEG[13] ,
    \Tile_X4Y3_N4BEG[12] ,
    \Tile_X4Y3_N4BEG[11] ,
    \Tile_X4Y3_N4BEG[10] ,
    \Tile_X4Y3_N4BEG[9] ,
    \Tile_X4Y3_N4BEG[8] ,
    \Tile_X4Y3_N4BEG[7] ,
    \Tile_X4Y3_N4BEG[6] ,
    \Tile_X4Y3_N4BEG[5] ,
    \Tile_X4Y3_N4BEG[4] ,
    \Tile_X4Y3_N4BEG[3] ,
    \Tile_X4Y3_N4BEG[2] ,
    \Tile_X4Y3_N4BEG[1] ,
    \Tile_X4Y3_N4BEG[0] }),
    .NN4BEG({\Tile_X4Y2_NN4BEG[15] ,
    \Tile_X4Y2_NN4BEG[14] ,
    \Tile_X4Y2_NN4BEG[13] ,
    \Tile_X4Y2_NN4BEG[12] ,
    \Tile_X4Y2_NN4BEG[11] ,
    \Tile_X4Y2_NN4BEG[10] ,
    \Tile_X4Y2_NN4BEG[9] ,
    \Tile_X4Y2_NN4BEG[8] ,
    \Tile_X4Y2_NN4BEG[7] ,
    \Tile_X4Y2_NN4BEG[6] ,
    \Tile_X4Y2_NN4BEG[5] ,
    \Tile_X4Y2_NN4BEG[4] ,
    \Tile_X4Y2_NN4BEG[3] ,
    \Tile_X4Y2_NN4BEG[2] ,
    \Tile_X4Y2_NN4BEG[1] ,
    \Tile_X4Y2_NN4BEG[0] }),
    .NN4END({\Tile_X4Y3_NN4BEG[15] ,
    \Tile_X4Y3_NN4BEG[14] ,
    \Tile_X4Y3_NN4BEG[13] ,
    \Tile_X4Y3_NN4BEG[12] ,
    \Tile_X4Y3_NN4BEG[11] ,
    \Tile_X4Y3_NN4BEG[10] ,
    \Tile_X4Y3_NN4BEG[9] ,
    \Tile_X4Y3_NN4BEG[8] ,
    \Tile_X4Y3_NN4BEG[7] ,
    \Tile_X4Y3_NN4BEG[6] ,
    \Tile_X4Y3_NN4BEG[5] ,
    \Tile_X4Y3_NN4BEG[4] ,
    \Tile_X4Y3_NN4BEG[3] ,
    \Tile_X4Y3_NN4BEG[2] ,
    \Tile_X4Y3_NN4BEG[1] ,
    \Tile_X4Y3_NN4BEG[0] }),
    .S1BEG({\Tile_X4Y2_S1BEG[3] ,
    \Tile_X4Y2_S1BEG[2] ,
    \Tile_X4Y2_S1BEG[1] ,
    \Tile_X4Y2_S1BEG[0] }),
    .S1END({\Tile_X4Y1_S1BEG[3] ,
    \Tile_X4Y1_S1BEG[2] ,
    \Tile_X4Y1_S1BEG[1] ,
    \Tile_X4Y1_S1BEG[0] }),
    .S2BEG({\Tile_X4Y2_S2BEG[7] ,
    \Tile_X4Y2_S2BEG[6] ,
    \Tile_X4Y2_S2BEG[5] ,
    \Tile_X4Y2_S2BEG[4] ,
    \Tile_X4Y2_S2BEG[3] ,
    \Tile_X4Y2_S2BEG[2] ,
    \Tile_X4Y2_S2BEG[1] ,
    \Tile_X4Y2_S2BEG[0] }),
    .S2BEGb({\Tile_X4Y2_S2BEGb[7] ,
    \Tile_X4Y2_S2BEGb[6] ,
    \Tile_X4Y2_S2BEGb[5] ,
    \Tile_X4Y2_S2BEGb[4] ,
    \Tile_X4Y2_S2BEGb[3] ,
    \Tile_X4Y2_S2BEGb[2] ,
    \Tile_X4Y2_S2BEGb[1] ,
    \Tile_X4Y2_S2BEGb[0] }),
    .S2END({\Tile_X4Y1_S2BEGb[7] ,
    \Tile_X4Y1_S2BEGb[6] ,
    \Tile_X4Y1_S2BEGb[5] ,
    \Tile_X4Y1_S2BEGb[4] ,
    \Tile_X4Y1_S2BEGb[3] ,
    \Tile_X4Y1_S2BEGb[2] ,
    \Tile_X4Y1_S2BEGb[1] ,
    \Tile_X4Y1_S2BEGb[0] }),
    .S2MID({\Tile_X4Y1_S2BEG[7] ,
    \Tile_X4Y1_S2BEG[6] ,
    \Tile_X4Y1_S2BEG[5] ,
    \Tile_X4Y1_S2BEG[4] ,
    \Tile_X4Y1_S2BEG[3] ,
    \Tile_X4Y1_S2BEG[2] ,
    \Tile_X4Y1_S2BEG[1] ,
    \Tile_X4Y1_S2BEG[0] }),
    .S4BEG({\Tile_X4Y2_S4BEG[15] ,
    \Tile_X4Y2_S4BEG[14] ,
    \Tile_X4Y2_S4BEG[13] ,
    \Tile_X4Y2_S4BEG[12] ,
    \Tile_X4Y2_S4BEG[11] ,
    \Tile_X4Y2_S4BEG[10] ,
    \Tile_X4Y2_S4BEG[9] ,
    \Tile_X4Y2_S4BEG[8] ,
    \Tile_X4Y2_S4BEG[7] ,
    \Tile_X4Y2_S4BEG[6] ,
    \Tile_X4Y2_S4BEG[5] ,
    \Tile_X4Y2_S4BEG[4] ,
    \Tile_X4Y2_S4BEG[3] ,
    \Tile_X4Y2_S4BEG[2] ,
    \Tile_X4Y2_S4BEG[1] ,
    \Tile_X4Y2_S4BEG[0] }),
    .S4END({\Tile_X4Y1_S4BEG[15] ,
    \Tile_X4Y1_S4BEG[14] ,
    \Tile_X4Y1_S4BEG[13] ,
    \Tile_X4Y1_S4BEG[12] ,
    \Tile_X4Y1_S4BEG[11] ,
    \Tile_X4Y1_S4BEG[10] ,
    \Tile_X4Y1_S4BEG[9] ,
    \Tile_X4Y1_S4BEG[8] ,
    \Tile_X4Y1_S4BEG[7] ,
    \Tile_X4Y1_S4BEG[6] ,
    \Tile_X4Y1_S4BEG[5] ,
    \Tile_X4Y1_S4BEG[4] ,
    \Tile_X4Y1_S4BEG[3] ,
    \Tile_X4Y1_S4BEG[2] ,
    \Tile_X4Y1_S4BEG[1] ,
    \Tile_X4Y1_S4BEG[0] }),
    .SS4BEG({\Tile_X4Y2_SS4BEG[15] ,
    \Tile_X4Y2_SS4BEG[14] ,
    \Tile_X4Y2_SS4BEG[13] ,
    \Tile_X4Y2_SS4BEG[12] ,
    \Tile_X4Y2_SS4BEG[11] ,
    \Tile_X4Y2_SS4BEG[10] ,
    \Tile_X4Y2_SS4BEG[9] ,
    \Tile_X4Y2_SS4BEG[8] ,
    \Tile_X4Y2_SS4BEG[7] ,
    \Tile_X4Y2_SS4BEG[6] ,
    \Tile_X4Y2_SS4BEG[5] ,
    \Tile_X4Y2_SS4BEG[4] ,
    \Tile_X4Y2_SS4BEG[3] ,
    \Tile_X4Y2_SS4BEG[2] ,
    \Tile_X4Y2_SS4BEG[1] ,
    \Tile_X4Y2_SS4BEG[0] }),
    .SS4END({\Tile_X4Y1_SS4BEG[15] ,
    \Tile_X4Y1_SS4BEG[14] ,
    \Tile_X4Y1_SS4BEG[13] ,
    \Tile_X4Y1_SS4BEG[12] ,
    \Tile_X4Y1_SS4BEG[11] ,
    \Tile_X4Y1_SS4BEG[10] ,
    \Tile_X4Y1_SS4BEG[9] ,
    \Tile_X4Y1_SS4BEG[8] ,
    \Tile_X4Y1_SS4BEG[7] ,
    \Tile_X4Y1_SS4BEG[6] ,
    \Tile_X4Y1_SS4BEG[5] ,
    \Tile_X4Y1_SS4BEG[4] ,
    \Tile_X4Y1_SS4BEG[3] ,
    \Tile_X4Y1_SS4BEG[2] ,
    \Tile_X4Y1_SS4BEG[1] ,
    \Tile_X4Y1_SS4BEG[0] }),
    .W1BEG({\Tile_X4Y2_W1BEG[3] ,
    \Tile_X4Y2_W1BEG[2] ,
    \Tile_X4Y2_W1BEG[1] ,
    \Tile_X4Y2_W1BEG[0] }),
    .W1END({\Tile_X5Y2_W1BEG[3] ,
    \Tile_X5Y2_W1BEG[2] ,
    \Tile_X5Y2_W1BEG[1] ,
    \Tile_X5Y2_W1BEG[0] }),
    .W2BEG({\Tile_X4Y2_W2BEG[7] ,
    \Tile_X4Y2_W2BEG[6] ,
    \Tile_X4Y2_W2BEG[5] ,
    \Tile_X4Y2_W2BEG[4] ,
    \Tile_X4Y2_W2BEG[3] ,
    \Tile_X4Y2_W2BEG[2] ,
    \Tile_X4Y2_W2BEG[1] ,
    \Tile_X4Y2_W2BEG[0] }),
    .W2BEGb({\Tile_X4Y2_W2BEGb[7] ,
    \Tile_X4Y2_W2BEGb[6] ,
    \Tile_X4Y2_W2BEGb[5] ,
    \Tile_X4Y2_W2BEGb[4] ,
    \Tile_X4Y2_W2BEGb[3] ,
    \Tile_X4Y2_W2BEGb[2] ,
    \Tile_X4Y2_W2BEGb[1] ,
    \Tile_X4Y2_W2BEGb[0] }),
    .W2END({\Tile_X5Y2_W2BEGb[7] ,
    \Tile_X5Y2_W2BEGb[6] ,
    \Tile_X5Y2_W2BEGb[5] ,
    \Tile_X5Y2_W2BEGb[4] ,
    \Tile_X5Y2_W2BEGb[3] ,
    \Tile_X5Y2_W2BEGb[2] ,
    \Tile_X5Y2_W2BEGb[1] ,
    \Tile_X5Y2_W2BEGb[0] }),
    .W2MID({\Tile_X5Y2_W2BEG[7] ,
    \Tile_X5Y2_W2BEG[6] ,
    \Tile_X5Y2_W2BEG[5] ,
    \Tile_X5Y2_W2BEG[4] ,
    \Tile_X5Y2_W2BEG[3] ,
    \Tile_X5Y2_W2BEG[2] ,
    \Tile_X5Y2_W2BEG[1] ,
    \Tile_X5Y2_W2BEG[0] }),
    .W6BEG({\Tile_X4Y2_W6BEG[11] ,
    \Tile_X4Y2_W6BEG[10] ,
    \Tile_X4Y2_W6BEG[9] ,
    \Tile_X4Y2_W6BEG[8] ,
    \Tile_X4Y2_W6BEG[7] ,
    \Tile_X4Y2_W6BEG[6] ,
    \Tile_X4Y2_W6BEG[5] ,
    \Tile_X4Y2_W6BEG[4] ,
    \Tile_X4Y2_W6BEG[3] ,
    \Tile_X4Y2_W6BEG[2] ,
    \Tile_X4Y2_W6BEG[1] ,
    \Tile_X4Y2_W6BEG[0] }),
    .W6END({\Tile_X5Y2_W6BEG[11] ,
    \Tile_X5Y2_W6BEG[10] ,
    \Tile_X5Y2_W6BEG[9] ,
    \Tile_X5Y2_W6BEG[8] ,
    \Tile_X5Y2_W6BEG[7] ,
    \Tile_X5Y2_W6BEG[6] ,
    \Tile_X5Y2_W6BEG[5] ,
    \Tile_X5Y2_W6BEG[4] ,
    \Tile_X5Y2_W6BEG[3] ,
    \Tile_X5Y2_W6BEG[2] ,
    \Tile_X5Y2_W6BEG[1] ,
    \Tile_X5Y2_W6BEG[0] }),
    .WW4BEG({\Tile_X4Y2_WW4BEG[15] ,
    \Tile_X4Y2_WW4BEG[14] ,
    \Tile_X4Y2_WW4BEG[13] ,
    \Tile_X4Y2_WW4BEG[12] ,
    \Tile_X4Y2_WW4BEG[11] ,
    \Tile_X4Y2_WW4BEG[10] ,
    \Tile_X4Y2_WW4BEG[9] ,
    \Tile_X4Y2_WW4BEG[8] ,
    \Tile_X4Y2_WW4BEG[7] ,
    \Tile_X4Y2_WW4BEG[6] ,
    \Tile_X4Y2_WW4BEG[5] ,
    \Tile_X4Y2_WW4BEG[4] ,
    \Tile_X4Y2_WW4BEG[3] ,
    \Tile_X4Y2_WW4BEG[2] ,
    \Tile_X4Y2_WW4BEG[1] ,
    \Tile_X4Y2_WW4BEG[0] }),
    .WW4END({\Tile_X5Y2_WW4BEG[15] ,
    \Tile_X5Y2_WW4BEG[14] ,
    \Tile_X5Y2_WW4BEG[13] ,
    \Tile_X5Y2_WW4BEG[12] ,
    \Tile_X5Y2_WW4BEG[11] ,
    \Tile_X5Y2_WW4BEG[10] ,
    \Tile_X5Y2_WW4BEG[9] ,
    \Tile_X5Y2_WW4BEG[8] ,
    \Tile_X5Y2_WW4BEG[7] ,
    \Tile_X5Y2_WW4BEG[6] ,
    \Tile_X5Y2_WW4BEG[5] ,
    \Tile_X5Y2_WW4BEG[4] ,
    \Tile_X5Y2_WW4BEG[3] ,
    \Tile_X5Y2_WW4BEG[2] ,
    \Tile_X5Y2_WW4BEG[1] ,
    \Tile_X5Y2_WW4BEG[0] }));
 RegFile Tile_X4Y3_RegFile (.UserCLK(Tile_X4Y4_UserCLKo),
    .UserCLKo(Tile_X4Y3_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X4Y3_E1BEG[3] ,
    \Tile_X4Y3_E1BEG[2] ,
    \Tile_X4Y3_E1BEG[1] ,
    \Tile_X4Y3_E1BEG[0] }),
    .E1END({\Tile_X3Y3_E1BEG[3] ,
    \Tile_X3Y3_E1BEG[2] ,
    \Tile_X3Y3_E1BEG[1] ,
    \Tile_X3Y3_E1BEG[0] }),
    .E2BEG({\Tile_X4Y3_E2BEG[7] ,
    \Tile_X4Y3_E2BEG[6] ,
    \Tile_X4Y3_E2BEG[5] ,
    \Tile_X4Y3_E2BEG[4] ,
    \Tile_X4Y3_E2BEG[3] ,
    \Tile_X4Y3_E2BEG[2] ,
    \Tile_X4Y3_E2BEG[1] ,
    \Tile_X4Y3_E2BEG[0] }),
    .E2BEGb({\Tile_X4Y3_E2BEGb[7] ,
    \Tile_X4Y3_E2BEGb[6] ,
    \Tile_X4Y3_E2BEGb[5] ,
    \Tile_X4Y3_E2BEGb[4] ,
    \Tile_X4Y3_E2BEGb[3] ,
    \Tile_X4Y3_E2BEGb[2] ,
    \Tile_X4Y3_E2BEGb[1] ,
    \Tile_X4Y3_E2BEGb[0] }),
    .E2END({\Tile_X3Y3_E2BEGb[7] ,
    \Tile_X3Y3_E2BEGb[6] ,
    \Tile_X3Y3_E2BEGb[5] ,
    \Tile_X3Y3_E2BEGb[4] ,
    \Tile_X3Y3_E2BEGb[3] ,
    \Tile_X3Y3_E2BEGb[2] ,
    \Tile_X3Y3_E2BEGb[1] ,
    \Tile_X3Y3_E2BEGb[0] }),
    .E2MID({\Tile_X3Y3_E2BEG[7] ,
    \Tile_X3Y3_E2BEG[6] ,
    \Tile_X3Y3_E2BEG[5] ,
    \Tile_X3Y3_E2BEG[4] ,
    \Tile_X3Y3_E2BEG[3] ,
    \Tile_X3Y3_E2BEG[2] ,
    \Tile_X3Y3_E2BEG[1] ,
    \Tile_X3Y3_E2BEG[0] }),
    .E6BEG({\Tile_X4Y3_E6BEG[11] ,
    \Tile_X4Y3_E6BEG[10] ,
    \Tile_X4Y3_E6BEG[9] ,
    \Tile_X4Y3_E6BEG[8] ,
    \Tile_X4Y3_E6BEG[7] ,
    \Tile_X4Y3_E6BEG[6] ,
    \Tile_X4Y3_E6BEG[5] ,
    \Tile_X4Y3_E6BEG[4] ,
    \Tile_X4Y3_E6BEG[3] ,
    \Tile_X4Y3_E6BEG[2] ,
    \Tile_X4Y3_E6BEG[1] ,
    \Tile_X4Y3_E6BEG[0] }),
    .E6END({\Tile_X3Y3_E6BEG[11] ,
    \Tile_X3Y3_E6BEG[10] ,
    \Tile_X3Y3_E6BEG[9] ,
    \Tile_X3Y3_E6BEG[8] ,
    \Tile_X3Y3_E6BEG[7] ,
    \Tile_X3Y3_E6BEG[6] ,
    \Tile_X3Y3_E6BEG[5] ,
    \Tile_X3Y3_E6BEG[4] ,
    \Tile_X3Y3_E6BEG[3] ,
    \Tile_X3Y3_E6BEG[2] ,
    \Tile_X3Y3_E6BEG[1] ,
    \Tile_X3Y3_E6BEG[0] }),
    .EE4BEG({\Tile_X4Y3_EE4BEG[15] ,
    \Tile_X4Y3_EE4BEG[14] ,
    \Tile_X4Y3_EE4BEG[13] ,
    \Tile_X4Y3_EE4BEG[12] ,
    \Tile_X4Y3_EE4BEG[11] ,
    \Tile_X4Y3_EE4BEG[10] ,
    \Tile_X4Y3_EE4BEG[9] ,
    \Tile_X4Y3_EE4BEG[8] ,
    \Tile_X4Y3_EE4BEG[7] ,
    \Tile_X4Y3_EE4BEG[6] ,
    \Tile_X4Y3_EE4BEG[5] ,
    \Tile_X4Y3_EE4BEG[4] ,
    \Tile_X4Y3_EE4BEG[3] ,
    \Tile_X4Y3_EE4BEG[2] ,
    \Tile_X4Y3_EE4BEG[1] ,
    \Tile_X4Y3_EE4BEG[0] }),
    .EE4END({\Tile_X3Y3_EE4BEG[15] ,
    \Tile_X3Y3_EE4BEG[14] ,
    \Tile_X3Y3_EE4BEG[13] ,
    \Tile_X3Y3_EE4BEG[12] ,
    \Tile_X3Y3_EE4BEG[11] ,
    \Tile_X3Y3_EE4BEG[10] ,
    \Tile_X3Y3_EE4BEG[9] ,
    \Tile_X3Y3_EE4BEG[8] ,
    \Tile_X3Y3_EE4BEG[7] ,
    \Tile_X3Y3_EE4BEG[6] ,
    \Tile_X3Y3_EE4BEG[5] ,
    \Tile_X3Y3_EE4BEG[4] ,
    \Tile_X3Y3_EE4BEG[3] ,
    \Tile_X3Y3_EE4BEG[2] ,
    \Tile_X3Y3_EE4BEG[1] ,
    \Tile_X3Y3_EE4BEG[0] }),
    .FrameData({\Tile_X3Y3_FrameData_O[31] ,
    \Tile_X3Y3_FrameData_O[30] ,
    \Tile_X3Y3_FrameData_O[29] ,
    \Tile_X3Y3_FrameData_O[28] ,
    \Tile_X3Y3_FrameData_O[27] ,
    \Tile_X3Y3_FrameData_O[26] ,
    \Tile_X3Y3_FrameData_O[25] ,
    \Tile_X3Y3_FrameData_O[24] ,
    \Tile_X3Y3_FrameData_O[23] ,
    \Tile_X3Y3_FrameData_O[22] ,
    \Tile_X3Y3_FrameData_O[21] ,
    \Tile_X3Y3_FrameData_O[20] ,
    \Tile_X3Y3_FrameData_O[19] ,
    \Tile_X3Y3_FrameData_O[18] ,
    \Tile_X3Y3_FrameData_O[17] ,
    \Tile_X3Y3_FrameData_O[16] ,
    \Tile_X3Y3_FrameData_O[15] ,
    \Tile_X3Y3_FrameData_O[14] ,
    \Tile_X3Y3_FrameData_O[13] ,
    \Tile_X3Y3_FrameData_O[12] ,
    \Tile_X3Y3_FrameData_O[11] ,
    \Tile_X3Y3_FrameData_O[10] ,
    \Tile_X3Y3_FrameData_O[9] ,
    \Tile_X3Y3_FrameData_O[8] ,
    \Tile_X3Y3_FrameData_O[7] ,
    \Tile_X3Y3_FrameData_O[6] ,
    \Tile_X3Y3_FrameData_O[5] ,
    \Tile_X3Y3_FrameData_O[4] ,
    \Tile_X3Y3_FrameData_O[3] ,
    \Tile_X3Y3_FrameData_O[2] ,
    \Tile_X3Y3_FrameData_O[1] ,
    \Tile_X3Y3_FrameData_O[0] }),
    .FrameData_O({\Tile_X4Y3_FrameData_O[31] ,
    \Tile_X4Y3_FrameData_O[30] ,
    \Tile_X4Y3_FrameData_O[29] ,
    \Tile_X4Y3_FrameData_O[28] ,
    \Tile_X4Y3_FrameData_O[27] ,
    \Tile_X4Y3_FrameData_O[26] ,
    \Tile_X4Y3_FrameData_O[25] ,
    \Tile_X4Y3_FrameData_O[24] ,
    \Tile_X4Y3_FrameData_O[23] ,
    \Tile_X4Y3_FrameData_O[22] ,
    \Tile_X4Y3_FrameData_O[21] ,
    \Tile_X4Y3_FrameData_O[20] ,
    \Tile_X4Y3_FrameData_O[19] ,
    \Tile_X4Y3_FrameData_O[18] ,
    \Tile_X4Y3_FrameData_O[17] ,
    \Tile_X4Y3_FrameData_O[16] ,
    \Tile_X4Y3_FrameData_O[15] ,
    \Tile_X4Y3_FrameData_O[14] ,
    \Tile_X4Y3_FrameData_O[13] ,
    \Tile_X4Y3_FrameData_O[12] ,
    \Tile_X4Y3_FrameData_O[11] ,
    \Tile_X4Y3_FrameData_O[10] ,
    \Tile_X4Y3_FrameData_O[9] ,
    \Tile_X4Y3_FrameData_O[8] ,
    \Tile_X4Y3_FrameData_O[7] ,
    \Tile_X4Y3_FrameData_O[6] ,
    \Tile_X4Y3_FrameData_O[5] ,
    \Tile_X4Y3_FrameData_O[4] ,
    \Tile_X4Y3_FrameData_O[3] ,
    \Tile_X4Y3_FrameData_O[2] ,
    \Tile_X4Y3_FrameData_O[1] ,
    \Tile_X4Y3_FrameData_O[0] }),
    .FrameStrobe({\Tile_X4Y4_FrameStrobe_O[19] ,
    \Tile_X4Y4_FrameStrobe_O[18] ,
    \Tile_X4Y4_FrameStrobe_O[17] ,
    \Tile_X4Y4_FrameStrobe_O[16] ,
    \Tile_X4Y4_FrameStrobe_O[15] ,
    \Tile_X4Y4_FrameStrobe_O[14] ,
    \Tile_X4Y4_FrameStrobe_O[13] ,
    \Tile_X4Y4_FrameStrobe_O[12] ,
    \Tile_X4Y4_FrameStrobe_O[11] ,
    \Tile_X4Y4_FrameStrobe_O[10] ,
    \Tile_X4Y4_FrameStrobe_O[9] ,
    \Tile_X4Y4_FrameStrobe_O[8] ,
    \Tile_X4Y4_FrameStrobe_O[7] ,
    \Tile_X4Y4_FrameStrobe_O[6] ,
    \Tile_X4Y4_FrameStrobe_O[5] ,
    \Tile_X4Y4_FrameStrobe_O[4] ,
    \Tile_X4Y4_FrameStrobe_O[3] ,
    \Tile_X4Y4_FrameStrobe_O[2] ,
    \Tile_X4Y4_FrameStrobe_O[1] ,
    \Tile_X4Y4_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X4Y3_FrameStrobe_O[19] ,
    \Tile_X4Y3_FrameStrobe_O[18] ,
    \Tile_X4Y3_FrameStrobe_O[17] ,
    \Tile_X4Y3_FrameStrobe_O[16] ,
    \Tile_X4Y3_FrameStrobe_O[15] ,
    \Tile_X4Y3_FrameStrobe_O[14] ,
    \Tile_X4Y3_FrameStrobe_O[13] ,
    \Tile_X4Y3_FrameStrobe_O[12] ,
    \Tile_X4Y3_FrameStrobe_O[11] ,
    \Tile_X4Y3_FrameStrobe_O[10] ,
    \Tile_X4Y3_FrameStrobe_O[9] ,
    \Tile_X4Y3_FrameStrobe_O[8] ,
    \Tile_X4Y3_FrameStrobe_O[7] ,
    \Tile_X4Y3_FrameStrobe_O[6] ,
    \Tile_X4Y3_FrameStrobe_O[5] ,
    \Tile_X4Y3_FrameStrobe_O[4] ,
    \Tile_X4Y3_FrameStrobe_O[3] ,
    \Tile_X4Y3_FrameStrobe_O[2] ,
    \Tile_X4Y3_FrameStrobe_O[1] ,
    \Tile_X4Y3_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X4Y3_N1BEG[3] ,
    \Tile_X4Y3_N1BEG[2] ,
    \Tile_X4Y3_N1BEG[1] ,
    \Tile_X4Y3_N1BEG[0] }),
    .N1END({\Tile_X4Y4_N1BEG[3] ,
    \Tile_X4Y4_N1BEG[2] ,
    \Tile_X4Y4_N1BEG[1] ,
    \Tile_X4Y4_N1BEG[0] }),
    .N2BEG({\Tile_X4Y3_N2BEG[7] ,
    \Tile_X4Y3_N2BEG[6] ,
    \Tile_X4Y3_N2BEG[5] ,
    \Tile_X4Y3_N2BEG[4] ,
    \Tile_X4Y3_N2BEG[3] ,
    \Tile_X4Y3_N2BEG[2] ,
    \Tile_X4Y3_N2BEG[1] ,
    \Tile_X4Y3_N2BEG[0] }),
    .N2BEGb({\Tile_X4Y3_N2BEGb[7] ,
    \Tile_X4Y3_N2BEGb[6] ,
    \Tile_X4Y3_N2BEGb[5] ,
    \Tile_X4Y3_N2BEGb[4] ,
    \Tile_X4Y3_N2BEGb[3] ,
    \Tile_X4Y3_N2BEGb[2] ,
    \Tile_X4Y3_N2BEGb[1] ,
    \Tile_X4Y3_N2BEGb[0] }),
    .N2END({\Tile_X4Y4_N2BEGb[7] ,
    \Tile_X4Y4_N2BEGb[6] ,
    \Tile_X4Y4_N2BEGb[5] ,
    \Tile_X4Y4_N2BEGb[4] ,
    \Tile_X4Y4_N2BEGb[3] ,
    \Tile_X4Y4_N2BEGb[2] ,
    \Tile_X4Y4_N2BEGb[1] ,
    \Tile_X4Y4_N2BEGb[0] }),
    .N2MID({\Tile_X4Y4_N2BEG[7] ,
    \Tile_X4Y4_N2BEG[6] ,
    \Tile_X4Y4_N2BEG[5] ,
    \Tile_X4Y4_N2BEG[4] ,
    \Tile_X4Y4_N2BEG[3] ,
    \Tile_X4Y4_N2BEG[2] ,
    \Tile_X4Y4_N2BEG[1] ,
    \Tile_X4Y4_N2BEG[0] }),
    .N4BEG({\Tile_X4Y3_N4BEG[15] ,
    \Tile_X4Y3_N4BEG[14] ,
    \Tile_X4Y3_N4BEG[13] ,
    \Tile_X4Y3_N4BEG[12] ,
    \Tile_X4Y3_N4BEG[11] ,
    \Tile_X4Y3_N4BEG[10] ,
    \Tile_X4Y3_N4BEG[9] ,
    \Tile_X4Y3_N4BEG[8] ,
    \Tile_X4Y3_N4BEG[7] ,
    \Tile_X4Y3_N4BEG[6] ,
    \Tile_X4Y3_N4BEG[5] ,
    \Tile_X4Y3_N4BEG[4] ,
    \Tile_X4Y3_N4BEG[3] ,
    \Tile_X4Y3_N4BEG[2] ,
    \Tile_X4Y3_N4BEG[1] ,
    \Tile_X4Y3_N4BEG[0] }),
    .N4END({\Tile_X4Y4_N4BEG[15] ,
    \Tile_X4Y4_N4BEG[14] ,
    \Tile_X4Y4_N4BEG[13] ,
    \Tile_X4Y4_N4BEG[12] ,
    \Tile_X4Y4_N4BEG[11] ,
    \Tile_X4Y4_N4BEG[10] ,
    \Tile_X4Y4_N4BEG[9] ,
    \Tile_X4Y4_N4BEG[8] ,
    \Tile_X4Y4_N4BEG[7] ,
    \Tile_X4Y4_N4BEG[6] ,
    \Tile_X4Y4_N4BEG[5] ,
    \Tile_X4Y4_N4BEG[4] ,
    \Tile_X4Y4_N4BEG[3] ,
    \Tile_X4Y4_N4BEG[2] ,
    \Tile_X4Y4_N4BEG[1] ,
    \Tile_X4Y4_N4BEG[0] }),
    .NN4BEG({\Tile_X4Y3_NN4BEG[15] ,
    \Tile_X4Y3_NN4BEG[14] ,
    \Tile_X4Y3_NN4BEG[13] ,
    \Tile_X4Y3_NN4BEG[12] ,
    \Tile_X4Y3_NN4BEG[11] ,
    \Tile_X4Y3_NN4BEG[10] ,
    \Tile_X4Y3_NN4BEG[9] ,
    \Tile_X4Y3_NN4BEG[8] ,
    \Tile_X4Y3_NN4BEG[7] ,
    \Tile_X4Y3_NN4BEG[6] ,
    \Tile_X4Y3_NN4BEG[5] ,
    \Tile_X4Y3_NN4BEG[4] ,
    \Tile_X4Y3_NN4BEG[3] ,
    \Tile_X4Y3_NN4BEG[2] ,
    \Tile_X4Y3_NN4BEG[1] ,
    \Tile_X4Y3_NN4BEG[0] }),
    .NN4END({\Tile_X4Y4_NN4BEG[15] ,
    \Tile_X4Y4_NN4BEG[14] ,
    \Tile_X4Y4_NN4BEG[13] ,
    \Tile_X4Y4_NN4BEG[12] ,
    \Tile_X4Y4_NN4BEG[11] ,
    \Tile_X4Y4_NN4BEG[10] ,
    \Tile_X4Y4_NN4BEG[9] ,
    \Tile_X4Y4_NN4BEG[8] ,
    \Tile_X4Y4_NN4BEG[7] ,
    \Tile_X4Y4_NN4BEG[6] ,
    \Tile_X4Y4_NN4BEG[5] ,
    \Tile_X4Y4_NN4BEG[4] ,
    \Tile_X4Y4_NN4BEG[3] ,
    \Tile_X4Y4_NN4BEG[2] ,
    \Tile_X4Y4_NN4BEG[1] ,
    \Tile_X4Y4_NN4BEG[0] }),
    .S1BEG({\Tile_X4Y3_S1BEG[3] ,
    \Tile_X4Y3_S1BEG[2] ,
    \Tile_X4Y3_S1BEG[1] ,
    \Tile_X4Y3_S1BEG[0] }),
    .S1END({\Tile_X4Y2_S1BEG[3] ,
    \Tile_X4Y2_S1BEG[2] ,
    \Tile_X4Y2_S1BEG[1] ,
    \Tile_X4Y2_S1BEG[0] }),
    .S2BEG({\Tile_X4Y3_S2BEG[7] ,
    \Tile_X4Y3_S2BEG[6] ,
    \Tile_X4Y3_S2BEG[5] ,
    \Tile_X4Y3_S2BEG[4] ,
    \Tile_X4Y3_S2BEG[3] ,
    \Tile_X4Y3_S2BEG[2] ,
    \Tile_X4Y3_S2BEG[1] ,
    \Tile_X4Y3_S2BEG[0] }),
    .S2BEGb({\Tile_X4Y3_S2BEGb[7] ,
    \Tile_X4Y3_S2BEGb[6] ,
    \Tile_X4Y3_S2BEGb[5] ,
    \Tile_X4Y3_S2BEGb[4] ,
    \Tile_X4Y3_S2BEGb[3] ,
    \Tile_X4Y3_S2BEGb[2] ,
    \Tile_X4Y3_S2BEGb[1] ,
    \Tile_X4Y3_S2BEGb[0] }),
    .S2END({\Tile_X4Y2_S2BEGb[7] ,
    \Tile_X4Y2_S2BEGb[6] ,
    \Tile_X4Y2_S2BEGb[5] ,
    \Tile_X4Y2_S2BEGb[4] ,
    \Tile_X4Y2_S2BEGb[3] ,
    \Tile_X4Y2_S2BEGb[2] ,
    \Tile_X4Y2_S2BEGb[1] ,
    \Tile_X4Y2_S2BEGb[0] }),
    .S2MID({\Tile_X4Y2_S2BEG[7] ,
    \Tile_X4Y2_S2BEG[6] ,
    \Tile_X4Y2_S2BEG[5] ,
    \Tile_X4Y2_S2BEG[4] ,
    \Tile_X4Y2_S2BEG[3] ,
    \Tile_X4Y2_S2BEG[2] ,
    \Tile_X4Y2_S2BEG[1] ,
    \Tile_X4Y2_S2BEG[0] }),
    .S4BEG({\Tile_X4Y3_S4BEG[15] ,
    \Tile_X4Y3_S4BEG[14] ,
    \Tile_X4Y3_S4BEG[13] ,
    \Tile_X4Y3_S4BEG[12] ,
    \Tile_X4Y3_S4BEG[11] ,
    \Tile_X4Y3_S4BEG[10] ,
    \Tile_X4Y3_S4BEG[9] ,
    \Tile_X4Y3_S4BEG[8] ,
    \Tile_X4Y3_S4BEG[7] ,
    \Tile_X4Y3_S4BEG[6] ,
    \Tile_X4Y3_S4BEG[5] ,
    \Tile_X4Y3_S4BEG[4] ,
    \Tile_X4Y3_S4BEG[3] ,
    \Tile_X4Y3_S4BEG[2] ,
    \Tile_X4Y3_S4BEG[1] ,
    \Tile_X4Y3_S4BEG[0] }),
    .S4END({\Tile_X4Y2_S4BEG[15] ,
    \Tile_X4Y2_S4BEG[14] ,
    \Tile_X4Y2_S4BEG[13] ,
    \Tile_X4Y2_S4BEG[12] ,
    \Tile_X4Y2_S4BEG[11] ,
    \Tile_X4Y2_S4BEG[10] ,
    \Tile_X4Y2_S4BEG[9] ,
    \Tile_X4Y2_S4BEG[8] ,
    \Tile_X4Y2_S4BEG[7] ,
    \Tile_X4Y2_S4BEG[6] ,
    \Tile_X4Y2_S4BEG[5] ,
    \Tile_X4Y2_S4BEG[4] ,
    \Tile_X4Y2_S4BEG[3] ,
    \Tile_X4Y2_S4BEG[2] ,
    \Tile_X4Y2_S4BEG[1] ,
    \Tile_X4Y2_S4BEG[0] }),
    .SS4BEG({\Tile_X4Y3_SS4BEG[15] ,
    \Tile_X4Y3_SS4BEG[14] ,
    \Tile_X4Y3_SS4BEG[13] ,
    \Tile_X4Y3_SS4BEG[12] ,
    \Tile_X4Y3_SS4BEG[11] ,
    \Tile_X4Y3_SS4BEG[10] ,
    \Tile_X4Y3_SS4BEG[9] ,
    \Tile_X4Y3_SS4BEG[8] ,
    \Tile_X4Y3_SS4BEG[7] ,
    \Tile_X4Y3_SS4BEG[6] ,
    \Tile_X4Y3_SS4BEG[5] ,
    \Tile_X4Y3_SS4BEG[4] ,
    \Tile_X4Y3_SS4BEG[3] ,
    \Tile_X4Y3_SS4BEG[2] ,
    \Tile_X4Y3_SS4BEG[1] ,
    \Tile_X4Y3_SS4BEG[0] }),
    .SS4END({\Tile_X4Y2_SS4BEG[15] ,
    \Tile_X4Y2_SS4BEG[14] ,
    \Tile_X4Y2_SS4BEG[13] ,
    \Tile_X4Y2_SS4BEG[12] ,
    \Tile_X4Y2_SS4BEG[11] ,
    \Tile_X4Y2_SS4BEG[10] ,
    \Tile_X4Y2_SS4BEG[9] ,
    \Tile_X4Y2_SS4BEG[8] ,
    \Tile_X4Y2_SS4BEG[7] ,
    \Tile_X4Y2_SS4BEG[6] ,
    \Tile_X4Y2_SS4BEG[5] ,
    \Tile_X4Y2_SS4BEG[4] ,
    \Tile_X4Y2_SS4BEG[3] ,
    \Tile_X4Y2_SS4BEG[2] ,
    \Tile_X4Y2_SS4BEG[1] ,
    \Tile_X4Y2_SS4BEG[0] }),
    .W1BEG({\Tile_X4Y3_W1BEG[3] ,
    \Tile_X4Y3_W1BEG[2] ,
    \Tile_X4Y3_W1BEG[1] ,
    \Tile_X4Y3_W1BEG[0] }),
    .W1END({\Tile_X5Y3_W1BEG[3] ,
    \Tile_X5Y3_W1BEG[2] ,
    \Tile_X5Y3_W1BEG[1] ,
    \Tile_X5Y3_W1BEG[0] }),
    .W2BEG({\Tile_X4Y3_W2BEG[7] ,
    \Tile_X4Y3_W2BEG[6] ,
    \Tile_X4Y3_W2BEG[5] ,
    \Tile_X4Y3_W2BEG[4] ,
    \Tile_X4Y3_W2BEG[3] ,
    \Tile_X4Y3_W2BEG[2] ,
    \Tile_X4Y3_W2BEG[1] ,
    \Tile_X4Y3_W2BEG[0] }),
    .W2BEGb({\Tile_X4Y3_W2BEGb[7] ,
    \Tile_X4Y3_W2BEGb[6] ,
    \Tile_X4Y3_W2BEGb[5] ,
    \Tile_X4Y3_W2BEGb[4] ,
    \Tile_X4Y3_W2BEGb[3] ,
    \Tile_X4Y3_W2BEGb[2] ,
    \Tile_X4Y3_W2BEGb[1] ,
    \Tile_X4Y3_W2BEGb[0] }),
    .W2END({\Tile_X5Y3_W2BEGb[7] ,
    \Tile_X5Y3_W2BEGb[6] ,
    \Tile_X5Y3_W2BEGb[5] ,
    \Tile_X5Y3_W2BEGb[4] ,
    \Tile_X5Y3_W2BEGb[3] ,
    \Tile_X5Y3_W2BEGb[2] ,
    \Tile_X5Y3_W2BEGb[1] ,
    \Tile_X5Y3_W2BEGb[0] }),
    .W2MID({\Tile_X5Y3_W2BEG[7] ,
    \Tile_X5Y3_W2BEG[6] ,
    \Tile_X5Y3_W2BEG[5] ,
    \Tile_X5Y3_W2BEG[4] ,
    \Tile_X5Y3_W2BEG[3] ,
    \Tile_X5Y3_W2BEG[2] ,
    \Tile_X5Y3_W2BEG[1] ,
    \Tile_X5Y3_W2BEG[0] }),
    .W6BEG({\Tile_X4Y3_W6BEG[11] ,
    \Tile_X4Y3_W6BEG[10] ,
    \Tile_X4Y3_W6BEG[9] ,
    \Tile_X4Y3_W6BEG[8] ,
    \Tile_X4Y3_W6BEG[7] ,
    \Tile_X4Y3_W6BEG[6] ,
    \Tile_X4Y3_W6BEG[5] ,
    \Tile_X4Y3_W6BEG[4] ,
    \Tile_X4Y3_W6BEG[3] ,
    \Tile_X4Y3_W6BEG[2] ,
    \Tile_X4Y3_W6BEG[1] ,
    \Tile_X4Y3_W6BEG[0] }),
    .W6END({\Tile_X5Y3_W6BEG[11] ,
    \Tile_X5Y3_W6BEG[10] ,
    \Tile_X5Y3_W6BEG[9] ,
    \Tile_X5Y3_W6BEG[8] ,
    \Tile_X5Y3_W6BEG[7] ,
    \Tile_X5Y3_W6BEG[6] ,
    \Tile_X5Y3_W6BEG[5] ,
    \Tile_X5Y3_W6BEG[4] ,
    \Tile_X5Y3_W6BEG[3] ,
    \Tile_X5Y3_W6BEG[2] ,
    \Tile_X5Y3_W6BEG[1] ,
    \Tile_X5Y3_W6BEG[0] }),
    .WW4BEG({\Tile_X4Y3_WW4BEG[15] ,
    \Tile_X4Y3_WW4BEG[14] ,
    \Tile_X4Y3_WW4BEG[13] ,
    \Tile_X4Y3_WW4BEG[12] ,
    \Tile_X4Y3_WW4BEG[11] ,
    \Tile_X4Y3_WW4BEG[10] ,
    \Tile_X4Y3_WW4BEG[9] ,
    \Tile_X4Y3_WW4BEG[8] ,
    \Tile_X4Y3_WW4BEG[7] ,
    \Tile_X4Y3_WW4BEG[6] ,
    \Tile_X4Y3_WW4BEG[5] ,
    \Tile_X4Y3_WW4BEG[4] ,
    \Tile_X4Y3_WW4BEG[3] ,
    \Tile_X4Y3_WW4BEG[2] ,
    \Tile_X4Y3_WW4BEG[1] ,
    \Tile_X4Y3_WW4BEG[0] }),
    .WW4END({\Tile_X5Y3_WW4BEG[15] ,
    \Tile_X5Y3_WW4BEG[14] ,
    \Tile_X5Y3_WW4BEG[13] ,
    \Tile_X5Y3_WW4BEG[12] ,
    \Tile_X5Y3_WW4BEG[11] ,
    \Tile_X5Y3_WW4BEG[10] ,
    \Tile_X5Y3_WW4BEG[9] ,
    \Tile_X5Y3_WW4BEG[8] ,
    \Tile_X5Y3_WW4BEG[7] ,
    \Tile_X5Y3_WW4BEG[6] ,
    \Tile_X5Y3_WW4BEG[5] ,
    \Tile_X5Y3_WW4BEG[4] ,
    \Tile_X5Y3_WW4BEG[3] ,
    \Tile_X5Y3_WW4BEG[2] ,
    \Tile_X5Y3_WW4BEG[1] ,
    \Tile_X5Y3_WW4BEG[0] }));
 RegFile Tile_X4Y4_RegFile (.UserCLK(Tile_X4Y5_UserCLKo),
    .UserCLKo(Tile_X4Y4_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X4Y4_E1BEG[3] ,
    \Tile_X4Y4_E1BEG[2] ,
    \Tile_X4Y4_E1BEG[1] ,
    \Tile_X4Y4_E1BEG[0] }),
    .E1END({\Tile_X3Y4_E1BEG[3] ,
    \Tile_X3Y4_E1BEG[2] ,
    \Tile_X3Y4_E1BEG[1] ,
    \Tile_X3Y4_E1BEG[0] }),
    .E2BEG({\Tile_X4Y4_E2BEG[7] ,
    \Tile_X4Y4_E2BEG[6] ,
    \Tile_X4Y4_E2BEG[5] ,
    \Tile_X4Y4_E2BEG[4] ,
    \Tile_X4Y4_E2BEG[3] ,
    \Tile_X4Y4_E2BEG[2] ,
    \Tile_X4Y4_E2BEG[1] ,
    \Tile_X4Y4_E2BEG[0] }),
    .E2BEGb({\Tile_X4Y4_E2BEGb[7] ,
    \Tile_X4Y4_E2BEGb[6] ,
    \Tile_X4Y4_E2BEGb[5] ,
    \Tile_X4Y4_E2BEGb[4] ,
    \Tile_X4Y4_E2BEGb[3] ,
    \Tile_X4Y4_E2BEGb[2] ,
    \Tile_X4Y4_E2BEGb[1] ,
    \Tile_X4Y4_E2BEGb[0] }),
    .E2END({\Tile_X3Y4_E2BEGb[7] ,
    \Tile_X3Y4_E2BEGb[6] ,
    \Tile_X3Y4_E2BEGb[5] ,
    \Tile_X3Y4_E2BEGb[4] ,
    \Tile_X3Y4_E2BEGb[3] ,
    \Tile_X3Y4_E2BEGb[2] ,
    \Tile_X3Y4_E2BEGb[1] ,
    \Tile_X3Y4_E2BEGb[0] }),
    .E2MID({\Tile_X3Y4_E2BEG[7] ,
    \Tile_X3Y4_E2BEG[6] ,
    \Tile_X3Y4_E2BEG[5] ,
    \Tile_X3Y4_E2BEG[4] ,
    \Tile_X3Y4_E2BEG[3] ,
    \Tile_X3Y4_E2BEG[2] ,
    \Tile_X3Y4_E2BEG[1] ,
    \Tile_X3Y4_E2BEG[0] }),
    .E6BEG({\Tile_X4Y4_E6BEG[11] ,
    \Tile_X4Y4_E6BEG[10] ,
    \Tile_X4Y4_E6BEG[9] ,
    \Tile_X4Y4_E6BEG[8] ,
    \Tile_X4Y4_E6BEG[7] ,
    \Tile_X4Y4_E6BEG[6] ,
    \Tile_X4Y4_E6BEG[5] ,
    \Tile_X4Y4_E6BEG[4] ,
    \Tile_X4Y4_E6BEG[3] ,
    \Tile_X4Y4_E6BEG[2] ,
    \Tile_X4Y4_E6BEG[1] ,
    \Tile_X4Y4_E6BEG[0] }),
    .E6END({\Tile_X3Y4_E6BEG[11] ,
    \Tile_X3Y4_E6BEG[10] ,
    \Tile_X3Y4_E6BEG[9] ,
    \Tile_X3Y4_E6BEG[8] ,
    \Tile_X3Y4_E6BEG[7] ,
    \Tile_X3Y4_E6BEG[6] ,
    \Tile_X3Y4_E6BEG[5] ,
    \Tile_X3Y4_E6BEG[4] ,
    \Tile_X3Y4_E6BEG[3] ,
    \Tile_X3Y4_E6BEG[2] ,
    \Tile_X3Y4_E6BEG[1] ,
    \Tile_X3Y4_E6BEG[0] }),
    .EE4BEG({\Tile_X4Y4_EE4BEG[15] ,
    \Tile_X4Y4_EE4BEG[14] ,
    \Tile_X4Y4_EE4BEG[13] ,
    \Tile_X4Y4_EE4BEG[12] ,
    \Tile_X4Y4_EE4BEG[11] ,
    \Tile_X4Y4_EE4BEG[10] ,
    \Tile_X4Y4_EE4BEG[9] ,
    \Tile_X4Y4_EE4BEG[8] ,
    \Tile_X4Y4_EE4BEG[7] ,
    \Tile_X4Y4_EE4BEG[6] ,
    \Tile_X4Y4_EE4BEG[5] ,
    \Tile_X4Y4_EE4BEG[4] ,
    \Tile_X4Y4_EE4BEG[3] ,
    \Tile_X4Y4_EE4BEG[2] ,
    \Tile_X4Y4_EE4BEG[1] ,
    \Tile_X4Y4_EE4BEG[0] }),
    .EE4END({\Tile_X3Y4_EE4BEG[15] ,
    \Tile_X3Y4_EE4BEG[14] ,
    \Tile_X3Y4_EE4BEG[13] ,
    \Tile_X3Y4_EE4BEG[12] ,
    \Tile_X3Y4_EE4BEG[11] ,
    \Tile_X3Y4_EE4BEG[10] ,
    \Tile_X3Y4_EE4BEG[9] ,
    \Tile_X3Y4_EE4BEG[8] ,
    \Tile_X3Y4_EE4BEG[7] ,
    \Tile_X3Y4_EE4BEG[6] ,
    \Tile_X3Y4_EE4BEG[5] ,
    \Tile_X3Y4_EE4BEG[4] ,
    \Tile_X3Y4_EE4BEG[3] ,
    \Tile_X3Y4_EE4BEG[2] ,
    \Tile_X3Y4_EE4BEG[1] ,
    \Tile_X3Y4_EE4BEG[0] }),
    .FrameData({\Tile_X3Y4_FrameData_O[31] ,
    \Tile_X3Y4_FrameData_O[30] ,
    \Tile_X3Y4_FrameData_O[29] ,
    \Tile_X3Y4_FrameData_O[28] ,
    \Tile_X3Y4_FrameData_O[27] ,
    \Tile_X3Y4_FrameData_O[26] ,
    \Tile_X3Y4_FrameData_O[25] ,
    \Tile_X3Y4_FrameData_O[24] ,
    \Tile_X3Y4_FrameData_O[23] ,
    \Tile_X3Y4_FrameData_O[22] ,
    \Tile_X3Y4_FrameData_O[21] ,
    \Tile_X3Y4_FrameData_O[20] ,
    \Tile_X3Y4_FrameData_O[19] ,
    \Tile_X3Y4_FrameData_O[18] ,
    \Tile_X3Y4_FrameData_O[17] ,
    \Tile_X3Y4_FrameData_O[16] ,
    \Tile_X3Y4_FrameData_O[15] ,
    \Tile_X3Y4_FrameData_O[14] ,
    \Tile_X3Y4_FrameData_O[13] ,
    \Tile_X3Y4_FrameData_O[12] ,
    \Tile_X3Y4_FrameData_O[11] ,
    \Tile_X3Y4_FrameData_O[10] ,
    \Tile_X3Y4_FrameData_O[9] ,
    \Tile_X3Y4_FrameData_O[8] ,
    \Tile_X3Y4_FrameData_O[7] ,
    \Tile_X3Y4_FrameData_O[6] ,
    \Tile_X3Y4_FrameData_O[5] ,
    \Tile_X3Y4_FrameData_O[4] ,
    \Tile_X3Y4_FrameData_O[3] ,
    \Tile_X3Y4_FrameData_O[2] ,
    \Tile_X3Y4_FrameData_O[1] ,
    \Tile_X3Y4_FrameData_O[0] }),
    .FrameData_O({\Tile_X4Y4_FrameData_O[31] ,
    \Tile_X4Y4_FrameData_O[30] ,
    \Tile_X4Y4_FrameData_O[29] ,
    \Tile_X4Y4_FrameData_O[28] ,
    \Tile_X4Y4_FrameData_O[27] ,
    \Tile_X4Y4_FrameData_O[26] ,
    \Tile_X4Y4_FrameData_O[25] ,
    \Tile_X4Y4_FrameData_O[24] ,
    \Tile_X4Y4_FrameData_O[23] ,
    \Tile_X4Y4_FrameData_O[22] ,
    \Tile_X4Y4_FrameData_O[21] ,
    \Tile_X4Y4_FrameData_O[20] ,
    \Tile_X4Y4_FrameData_O[19] ,
    \Tile_X4Y4_FrameData_O[18] ,
    \Tile_X4Y4_FrameData_O[17] ,
    \Tile_X4Y4_FrameData_O[16] ,
    \Tile_X4Y4_FrameData_O[15] ,
    \Tile_X4Y4_FrameData_O[14] ,
    \Tile_X4Y4_FrameData_O[13] ,
    \Tile_X4Y4_FrameData_O[12] ,
    \Tile_X4Y4_FrameData_O[11] ,
    \Tile_X4Y4_FrameData_O[10] ,
    \Tile_X4Y4_FrameData_O[9] ,
    \Tile_X4Y4_FrameData_O[8] ,
    \Tile_X4Y4_FrameData_O[7] ,
    \Tile_X4Y4_FrameData_O[6] ,
    \Tile_X4Y4_FrameData_O[5] ,
    \Tile_X4Y4_FrameData_O[4] ,
    \Tile_X4Y4_FrameData_O[3] ,
    \Tile_X4Y4_FrameData_O[2] ,
    \Tile_X4Y4_FrameData_O[1] ,
    \Tile_X4Y4_FrameData_O[0] }),
    .FrameStrobe({\Tile_X4Y5_FrameStrobe_O[19] ,
    \Tile_X4Y5_FrameStrobe_O[18] ,
    \Tile_X4Y5_FrameStrobe_O[17] ,
    \Tile_X4Y5_FrameStrobe_O[16] ,
    \Tile_X4Y5_FrameStrobe_O[15] ,
    \Tile_X4Y5_FrameStrobe_O[14] ,
    \Tile_X4Y5_FrameStrobe_O[13] ,
    \Tile_X4Y5_FrameStrobe_O[12] ,
    \Tile_X4Y5_FrameStrobe_O[11] ,
    \Tile_X4Y5_FrameStrobe_O[10] ,
    \Tile_X4Y5_FrameStrobe_O[9] ,
    \Tile_X4Y5_FrameStrobe_O[8] ,
    \Tile_X4Y5_FrameStrobe_O[7] ,
    \Tile_X4Y5_FrameStrobe_O[6] ,
    \Tile_X4Y5_FrameStrobe_O[5] ,
    \Tile_X4Y5_FrameStrobe_O[4] ,
    \Tile_X4Y5_FrameStrobe_O[3] ,
    \Tile_X4Y5_FrameStrobe_O[2] ,
    \Tile_X4Y5_FrameStrobe_O[1] ,
    \Tile_X4Y5_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X4Y4_FrameStrobe_O[19] ,
    \Tile_X4Y4_FrameStrobe_O[18] ,
    \Tile_X4Y4_FrameStrobe_O[17] ,
    \Tile_X4Y4_FrameStrobe_O[16] ,
    \Tile_X4Y4_FrameStrobe_O[15] ,
    \Tile_X4Y4_FrameStrobe_O[14] ,
    \Tile_X4Y4_FrameStrobe_O[13] ,
    \Tile_X4Y4_FrameStrobe_O[12] ,
    \Tile_X4Y4_FrameStrobe_O[11] ,
    \Tile_X4Y4_FrameStrobe_O[10] ,
    \Tile_X4Y4_FrameStrobe_O[9] ,
    \Tile_X4Y4_FrameStrobe_O[8] ,
    \Tile_X4Y4_FrameStrobe_O[7] ,
    \Tile_X4Y4_FrameStrobe_O[6] ,
    \Tile_X4Y4_FrameStrobe_O[5] ,
    \Tile_X4Y4_FrameStrobe_O[4] ,
    \Tile_X4Y4_FrameStrobe_O[3] ,
    \Tile_X4Y4_FrameStrobe_O[2] ,
    \Tile_X4Y4_FrameStrobe_O[1] ,
    \Tile_X4Y4_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X4Y4_N1BEG[3] ,
    \Tile_X4Y4_N1BEG[2] ,
    \Tile_X4Y4_N1BEG[1] ,
    \Tile_X4Y4_N1BEG[0] }),
    .N1END({\Tile_X4Y5_N1BEG[3] ,
    \Tile_X4Y5_N1BEG[2] ,
    \Tile_X4Y5_N1BEG[1] ,
    \Tile_X4Y5_N1BEG[0] }),
    .N2BEG({\Tile_X4Y4_N2BEG[7] ,
    \Tile_X4Y4_N2BEG[6] ,
    \Tile_X4Y4_N2BEG[5] ,
    \Tile_X4Y4_N2BEG[4] ,
    \Tile_X4Y4_N2BEG[3] ,
    \Tile_X4Y4_N2BEG[2] ,
    \Tile_X4Y4_N2BEG[1] ,
    \Tile_X4Y4_N2BEG[0] }),
    .N2BEGb({\Tile_X4Y4_N2BEGb[7] ,
    \Tile_X4Y4_N2BEGb[6] ,
    \Tile_X4Y4_N2BEGb[5] ,
    \Tile_X4Y4_N2BEGb[4] ,
    \Tile_X4Y4_N2BEGb[3] ,
    \Tile_X4Y4_N2BEGb[2] ,
    \Tile_X4Y4_N2BEGb[1] ,
    \Tile_X4Y4_N2BEGb[0] }),
    .N2END({\Tile_X4Y5_N2BEGb[7] ,
    \Tile_X4Y5_N2BEGb[6] ,
    \Tile_X4Y5_N2BEGb[5] ,
    \Tile_X4Y5_N2BEGb[4] ,
    \Tile_X4Y5_N2BEGb[3] ,
    \Tile_X4Y5_N2BEGb[2] ,
    \Tile_X4Y5_N2BEGb[1] ,
    \Tile_X4Y5_N2BEGb[0] }),
    .N2MID({\Tile_X4Y5_N2BEG[7] ,
    \Tile_X4Y5_N2BEG[6] ,
    \Tile_X4Y5_N2BEG[5] ,
    \Tile_X4Y5_N2BEG[4] ,
    \Tile_X4Y5_N2BEG[3] ,
    \Tile_X4Y5_N2BEG[2] ,
    \Tile_X4Y5_N2BEG[1] ,
    \Tile_X4Y5_N2BEG[0] }),
    .N4BEG({\Tile_X4Y4_N4BEG[15] ,
    \Tile_X4Y4_N4BEG[14] ,
    \Tile_X4Y4_N4BEG[13] ,
    \Tile_X4Y4_N4BEG[12] ,
    \Tile_X4Y4_N4BEG[11] ,
    \Tile_X4Y4_N4BEG[10] ,
    \Tile_X4Y4_N4BEG[9] ,
    \Tile_X4Y4_N4BEG[8] ,
    \Tile_X4Y4_N4BEG[7] ,
    \Tile_X4Y4_N4BEG[6] ,
    \Tile_X4Y4_N4BEG[5] ,
    \Tile_X4Y4_N4BEG[4] ,
    \Tile_X4Y4_N4BEG[3] ,
    \Tile_X4Y4_N4BEG[2] ,
    \Tile_X4Y4_N4BEG[1] ,
    \Tile_X4Y4_N4BEG[0] }),
    .N4END({\Tile_X4Y5_N4BEG[15] ,
    \Tile_X4Y5_N4BEG[14] ,
    \Tile_X4Y5_N4BEG[13] ,
    \Tile_X4Y5_N4BEG[12] ,
    \Tile_X4Y5_N4BEG[11] ,
    \Tile_X4Y5_N4BEG[10] ,
    \Tile_X4Y5_N4BEG[9] ,
    \Tile_X4Y5_N4BEG[8] ,
    \Tile_X4Y5_N4BEG[7] ,
    \Tile_X4Y5_N4BEG[6] ,
    \Tile_X4Y5_N4BEG[5] ,
    \Tile_X4Y5_N4BEG[4] ,
    \Tile_X4Y5_N4BEG[3] ,
    \Tile_X4Y5_N4BEG[2] ,
    \Tile_X4Y5_N4BEG[1] ,
    \Tile_X4Y5_N4BEG[0] }),
    .NN4BEG({\Tile_X4Y4_NN4BEG[15] ,
    \Tile_X4Y4_NN4BEG[14] ,
    \Tile_X4Y4_NN4BEG[13] ,
    \Tile_X4Y4_NN4BEG[12] ,
    \Tile_X4Y4_NN4BEG[11] ,
    \Tile_X4Y4_NN4BEG[10] ,
    \Tile_X4Y4_NN4BEG[9] ,
    \Tile_X4Y4_NN4BEG[8] ,
    \Tile_X4Y4_NN4BEG[7] ,
    \Tile_X4Y4_NN4BEG[6] ,
    \Tile_X4Y4_NN4BEG[5] ,
    \Tile_X4Y4_NN4BEG[4] ,
    \Tile_X4Y4_NN4BEG[3] ,
    \Tile_X4Y4_NN4BEG[2] ,
    \Tile_X4Y4_NN4BEG[1] ,
    \Tile_X4Y4_NN4BEG[0] }),
    .NN4END({\Tile_X4Y5_NN4BEG[15] ,
    \Tile_X4Y5_NN4BEG[14] ,
    \Tile_X4Y5_NN4BEG[13] ,
    \Tile_X4Y5_NN4BEG[12] ,
    \Tile_X4Y5_NN4BEG[11] ,
    \Tile_X4Y5_NN4BEG[10] ,
    \Tile_X4Y5_NN4BEG[9] ,
    \Tile_X4Y5_NN4BEG[8] ,
    \Tile_X4Y5_NN4BEG[7] ,
    \Tile_X4Y5_NN4BEG[6] ,
    \Tile_X4Y5_NN4BEG[5] ,
    \Tile_X4Y5_NN4BEG[4] ,
    \Tile_X4Y5_NN4BEG[3] ,
    \Tile_X4Y5_NN4BEG[2] ,
    \Tile_X4Y5_NN4BEG[1] ,
    \Tile_X4Y5_NN4BEG[0] }),
    .S1BEG({\Tile_X4Y4_S1BEG[3] ,
    \Tile_X4Y4_S1BEG[2] ,
    \Tile_X4Y4_S1BEG[1] ,
    \Tile_X4Y4_S1BEG[0] }),
    .S1END({\Tile_X4Y3_S1BEG[3] ,
    \Tile_X4Y3_S1BEG[2] ,
    \Tile_X4Y3_S1BEG[1] ,
    \Tile_X4Y3_S1BEG[0] }),
    .S2BEG({\Tile_X4Y4_S2BEG[7] ,
    \Tile_X4Y4_S2BEG[6] ,
    \Tile_X4Y4_S2BEG[5] ,
    \Tile_X4Y4_S2BEG[4] ,
    \Tile_X4Y4_S2BEG[3] ,
    \Tile_X4Y4_S2BEG[2] ,
    \Tile_X4Y4_S2BEG[1] ,
    \Tile_X4Y4_S2BEG[0] }),
    .S2BEGb({\Tile_X4Y4_S2BEGb[7] ,
    \Tile_X4Y4_S2BEGb[6] ,
    \Tile_X4Y4_S2BEGb[5] ,
    \Tile_X4Y4_S2BEGb[4] ,
    \Tile_X4Y4_S2BEGb[3] ,
    \Tile_X4Y4_S2BEGb[2] ,
    \Tile_X4Y4_S2BEGb[1] ,
    \Tile_X4Y4_S2BEGb[0] }),
    .S2END({\Tile_X4Y3_S2BEGb[7] ,
    \Tile_X4Y3_S2BEGb[6] ,
    \Tile_X4Y3_S2BEGb[5] ,
    \Tile_X4Y3_S2BEGb[4] ,
    \Tile_X4Y3_S2BEGb[3] ,
    \Tile_X4Y3_S2BEGb[2] ,
    \Tile_X4Y3_S2BEGb[1] ,
    \Tile_X4Y3_S2BEGb[0] }),
    .S2MID({\Tile_X4Y3_S2BEG[7] ,
    \Tile_X4Y3_S2BEG[6] ,
    \Tile_X4Y3_S2BEG[5] ,
    \Tile_X4Y3_S2BEG[4] ,
    \Tile_X4Y3_S2BEG[3] ,
    \Tile_X4Y3_S2BEG[2] ,
    \Tile_X4Y3_S2BEG[1] ,
    \Tile_X4Y3_S2BEG[0] }),
    .S4BEG({\Tile_X4Y4_S4BEG[15] ,
    \Tile_X4Y4_S4BEG[14] ,
    \Tile_X4Y4_S4BEG[13] ,
    \Tile_X4Y4_S4BEG[12] ,
    \Tile_X4Y4_S4BEG[11] ,
    \Tile_X4Y4_S4BEG[10] ,
    \Tile_X4Y4_S4BEG[9] ,
    \Tile_X4Y4_S4BEG[8] ,
    \Tile_X4Y4_S4BEG[7] ,
    \Tile_X4Y4_S4BEG[6] ,
    \Tile_X4Y4_S4BEG[5] ,
    \Tile_X4Y4_S4BEG[4] ,
    \Tile_X4Y4_S4BEG[3] ,
    \Tile_X4Y4_S4BEG[2] ,
    \Tile_X4Y4_S4BEG[1] ,
    \Tile_X4Y4_S4BEG[0] }),
    .S4END({\Tile_X4Y3_S4BEG[15] ,
    \Tile_X4Y3_S4BEG[14] ,
    \Tile_X4Y3_S4BEG[13] ,
    \Tile_X4Y3_S4BEG[12] ,
    \Tile_X4Y3_S4BEG[11] ,
    \Tile_X4Y3_S4BEG[10] ,
    \Tile_X4Y3_S4BEG[9] ,
    \Tile_X4Y3_S4BEG[8] ,
    \Tile_X4Y3_S4BEG[7] ,
    \Tile_X4Y3_S4BEG[6] ,
    \Tile_X4Y3_S4BEG[5] ,
    \Tile_X4Y3_S4BEG[4] ,
    \Tile_X4Y3_S4BEG[3] ,
    \Tile_X4Y3_S4BEG[2] ,
    \Tile_X4Y3_S4BEG[1] ,
    \Tile_X4Y3_S4BEG[0] }),
    .SS4BEG({\Tile_X4Y4_SS4BEG[15] ,
    \Tile_X4Y4_SS4BEG[14] ,
    \Tile_X4Y4_SS4BEG[13] ,
    \Tile_X4Y4_SS4BEG[12] ,
    \Tile_X4Y4_SS4BEG[11] ,
    \Tile_X4Y4_SS4BEG[10] ,
    \Tile_X4Y4_SS4BEG[9] ,
    \Tile_X4Y4_SS4BEG[8] ,
    \Tile_X4Y4_SS4BEG[7] ,
    \Tile_X4Y4_SS4BEG[6] ,
    \Tile_X4Y4_SS4BEG[5] ,
    \Tile_X4Y4_SS4BEG[4] ,
    \Tile_X4Y4_SS4BEG[3] ,
    \Tile_X4Y4_SS4BEG[2] ,
    \Tile_X4Y4_SS4BEG[1] ,
    \Tile_X4Y4_SS4BEG[0] }),
    .SS4END({\Tile_X4Y3_SS4BEG[15] ,
    \Tile_X4Y3_SS4BEG[14] ,
    \Tile_X4Y3_SS4BEG[13] ,
    \Tile_X4Y3_SS4BEG[12] ,
    \Tile_X4Y3_SS4BEG[11] ,
    \Tile_X4Y3_SS4BEG[10] ,
    \Tile_X4Y3_SS4BEG[9] ,
    \Tile_X4Y3_SS4BEG[8] ,
    \Tile_X4Y3_SS4BEG[7] ,
    \Tile_X4Y3_SS4BEG[6] ,
    \Tile_X4Y3_SS4BEG[5] ,
    \Tile_X4Y3_SS4BEG[4] ,
    \Tile_X4Y3_SS4BEG[3] ,
    \Tile_X4Y3_SS4BEG[2] ,
    \Tile_X4Y3_SS4BEG[1] ,
    \Tile_X4Y3_SS4BEG[0] }),
    .W1BEG({\Tile_X4Y4_W1BEG[3] ,
    \Tile_X4Y4_W1BEG[2] ,
    \Tile_X4Y4_W1BEG[1] ,
    \Tile_X4Y4_W1BEG[0] }),
    .W1END({\Tile_X5Y4_W1BEG[3] ,
    \Tile_X5Y4_W1BEG[2] ,
    \Tile_X5Y4_W1BEG[1] ,
    \Tile_X5Y4_W1BEG[0] }),
    .W2BEG({\Tile_X4Y4_W2BEG[7] ,
    \Tile_X4Y4_W2BEG[6] ,
    \Tile_X4Y4_W2BEG[5] ,
    \Tile_X4Y4_W2BEG[4] ,
    \Tile_X4Y4_W2BEG[3] ,
    \Tile_X4Y4_W2BEG[2] ,
    \Tile_X4Y4_W2BEG[1] ,
    \Tile_X4Y4_W2BEG[0] }),
    .W2BEGb({\Tile_X4Y4_W2BEGb[7] ,
    \Tile_X4Y4_W2BEGb[6] ,
    \Tile_X4Y4_W2BEGb[5] ,
    \Tile_X4Y4_W2BEGb[4] ,
    \Tile_X4Y4_W2BEGb[3] ,
    \Tile_X4Y4_W2BEGb[2] ,
    \Tile_X4Y4_W2BEGb[1] ,
    \Tile_X4Y4_W2BEGb[0] }),
    .W2END({\Tile_X5Y4_W2BEGb[7] ,
    \Tile_X5Y4_W2BEGb[6] ,
    \Tile_X5Y4_W2BEGb[5] ,
    \Tile_X5Y4_W2BEGb[4] ,
    \Tile_X5Y4_W2BEGb[3] ,
    \Tile_X5Y4_W2BEGb[2] ,
    \Tile_X5Y4_W2BEGb[1] ,
    \Tile_X5Y4_W2BEGb[0] }),
    .W2MID({\Tile_X5Y4_W2BEG[7] ,
    \Tile_X5Y4_W2BEG[6] ,
    \Tile_X5Y4_W2BEG[5] ,
    \Tile_X5Y4_W2BEG[4] ,
    \Tile_X5Y4_W2BEG[3] ,
    \Tile_X5Y4_W2BEG[2] ,
    \Tile_X5Y4_W2BEG[1] ,
    \Tile_X5Y4_W2BEG[0] }),
    .W6BEG({\Tile_X4Y4_W6BEG[11] ,
    \Tile_X4Y4_W6BEG[10] ,
    \Tile_X4Y4_W6BEG[9] ,
    \Tile_X4Y4_W6BEG[8] ,
    \Tile_X4Y4_W6BEG[7] ,
    \Tile_X4Y4_W6BEG[6] ,
    \Tile_X4Y4_W6BEG[5] ,
    \Tile_X4Y4_W6BEG[4] ,
    \Tile_X4Y4_W6BEG[3] ,
    \Tile_X4Y4_W6BEG[2] ,
    \Tile_X4Y4_W6BEG[1] ,
    \Tile_X4Y4_W6BEG[0] }),
    .W6END({\Tile_X5Y4_W6BEG[11] ,
    \Tile_X5Y4_W6BEG[10] ,
    \Tile_X5Y4_W6BEG[9] ,
    \Tile_X5Y4_W6BEG[8] ,
    \Tile_X5Y4_W6BEG[7] ,
    \Tile_X5Y4_W6BEG[6] ,
    \Tile_X5Y4_W6BEG[5] ,
    \Tile_X5Y4_W6BEG[4] ,
    \Tile_X5Y4_W6BEG[3] ,
    \Tile_X5Y4_W6BEG[2] ,
    \Tile_X5Y4_W6BEG[1] ,
    \Tile_X5Y4_W6BEG[0] }),
    .WW4BEG({\Tile_X4Y4_WW4BEG[15] ,
    \Tile_X4Y4_WW4BEG[14] ,
    \Tile_X4Y4_WW4BEG[13] ,
    \Tile_X4Y4_WW4BEG[12] ,
    \Tile_X4Y4_WW4BEG[11] ,
    \Tile_X4Y4_WW4BEG[10] ,
    \Tile_X4Y4_WW4BEG[9] ,
    \Tile_X4Y4_WW4BEG[8] ,
    \Tile_X4Y4_WW4BEG[7] ,
    \Tile_X4Y4_WW4BEG[6] ,
    \Tile_X4Y4_WW4BEG[5] ,
    \Tile_X4Y4_WW4BEG[4] ,
    \Tile_X4Y4_WW4BEG[3] ,
    \Tile_X4Y4_WW4BEG[2] ,
    \Tile_X4Y4_WW4BEG[1] ,
    \Tile_X4Y4_WW4BEG[0] }),
    .WW4END({\Tile_X5Y4_WW4BEG[15] ,
    \Tile_X5Y4_WW4BEG[14] ,
    \Tile_X5Y4_WW4BEG[13] ,
    \Tile_X5Y4_WW4BEG[12] ,
    \Tile_X5Y4_WW4BEG[11] ,
    \Tile_X5Y4_WW4BEG[10] ,
    \Tile_X5Y4_WW4BEG[9] ,
    \Tile_X5Y4_WW4BEG[8] ,
    \Tile_X5Y4_WW4BEG[7] ,
    \Tile_X5Y4_WW4BEG[6] ,
    \Tile_X5Y4_WW4BEG[5] ,
    \Tile_X5Y4_WW4BEG[4] ,
    \Tile_X5Y4_WW4BEG[3] ,
    \Tile_X5Y4_WW4BEG[2] ,
    \Tile_X5Y4_WW4BEG[1] ,
    \Tile_X5Y4_WW4BEG[0] }));
 RegFile Tile_X4Y5_RegFile (.UserCLK(Tile_X4Y6_UserCLKo),
    .UserCLKo(Tile_X4Y5_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X4Y5_E1BEG[3] ,
    \Tile_X4Y5_E1BEG[2] ,
    \Tile_X4Y5_E1BEG[1] ,
    \Tile_X4Y5_E1BEG[0] }),
    .E1END({\Tile_X3Y5_E1BEG[3] ,
    \Tile_X3Y5_E1BEG[2] ,
    \Tile_X3Y5_E1BEG[1] ,
    \Tile_X3Y5_E1BEG[0] }),
    .E2BEG({\Tile_X4Y5_E2BEG[7] ,
    \Tile_X4Y5_E2BEG[6] ,
    \Tile_X4Y5_E2BEG[5] ,
    \Tile_X4Y5_E2BEG[4] ,
    \Tile_X4Y5_E2BEG[3] ,
    \Tile_X4Y5_E2BEG[2] ,
    \Tile_X4Y5_E2BEG[1] ,
    \Tile_X4Y5_E2BEG[0] }),
    .E2BEGb({\Tile_X4Y5_E2BEGb[7] ,
    \Tile_X4Y5_E2BEGb[6] ,
    \Tile_X4Y5_E2BEGb[5] ,
    \Tile_X4Y5_E2BEGb[4] ,
    \Tile_X4Y5_E2BEGb[3] ,
    \Tile_X4Y5_E2BEGb[2] ,
    \Tile_X4Y5_E2BEGb[1] ,
    \Tile_X4Y5_E2BEGb[0] }),
    .E2END({\Tile_X3Y5_E2BEGb[7] ,
    \Tile_X3Y5_E2BEGb[6] ,
    \Tile_X3Y5_E2BEGb[5] ,
    \Tile_X3Y5_E2BEGb[4] ,
    \Tile_X3Y5_E2BEGb[3] ,
    \Tile_X3Y5_E2BEGb[2] ,
    \Tile_X3Y5_E2BEGb[1] ,
    \Tile_X3Y5_E2BEGb[0] }),
    .E2MID({\Tile_X3Y5_E2BEG[7] ,
    \Tile_X3Y5_E2BEG[6] ,
    \Tile_X3Y5_E2BEG[5] ,
    \Tile_X3Y5_E2BEG[4] ,
    \Tile_X3Y5_E2BEG[3] ,
    \Tile_X3Y5_E2BEG[2] ,
    \Tile_X3Y5_E2BEG[1] ,
    \Tile_X3Y5_E2BEG[0] }),
    .E6BEG({\Tile_X4Y5_E6BEG[11] ,
    \Tile_X4Y5_E6BEG[10] ,
    \Tile_X4Y5_E6BEG[9] ,
    \Tile_X4Y5_E6BEG[8] ,
    \Tile_X4Y5_E6BEG[7] ,
    \Tile_X4Y5_E6BEG[6] ,
    \Tile_X4Y5_E6BEG[5] ,
    \Tile_X4Y5_E6BEG[4] ,
    \Tile_X4Y5_E6BEG[3] ,
    \Tile_X4Y5_E6BEG[2] ,
    \Tile_X4Y5_E6BEG[1] ,
    \Tile_X4Y5_E6BEG[0] }),
    .E6END({\Tile_X3Y5_E6BEG[11] ,
    \Tile_X3Y5_E6BEG[10] ,
    \Tile_X3Y5_E6BEG[9] ,
    \Tile_X3Y5_E6BEG[8] ,
    \Tile_X3Y5_E6BEG[7] ,
    \Tile_X3Y5_E6BEG[6] ,
    \Tile_X3Y5_E6BEG[5] ,
    \Tile_X3Y5_E6BEG[4] ,
    \Tile_X3Y5_E6BEG[3] ,
    \Tile_X3Y5_E6BEG[2] ,
    \Tile_X3Y5_E6BEG[1] ,
    \Tile_X3Y5_E6BEG[0] }),
    .EE4BEG({\Tile_X4Y5_EE4BEG[15] ,
    \Tile_X4Y5_EE4BEG[14] ,
    \Tile_X4Y5_EE4BEG[13] ,
    \Tile_X4Y5_EE4BEG[12] ,
    \Tile_X4Y5_EE4BEG[11] ,
    \Tile_X4Y5_EE4BEG[10] ,
    \Tile_X4Y5_EE4BEG[9] ,
    \Tile_X4Y5_EE4BEG[8] ,
    \Tile_X4Y5_EE4BEG[7] ,
    \Tile_X4Y5_EE4BEG[6] ,
    \Tile_X4Y5_EE4BEG[5] ,
    \Tile_X4Y5_EE4BEG[4] ,
    \Tile_X4Y5_EE4BEG[3] ,
    \Tile_X4Y5_EE4BEG[2] ,
    \Tile_X4Y5_EE4BEG[1] ,
    \Tile_X4Y5_EE4BEG[0] }),
    .EE4END({\Tile_X3Y5_EE4BEG[15] ,
    \Tile_X3Y5_EE4BEG[14] ,
    \Tile_X3Y5_EE4BEG[13] ,
    \Tile_X3Y5_EE4BEG[12] ,
    \Tile_X3Y5_EE4BEG[11] ,
    \Tile_X3Y5_EE4BEG[10] ,
    \Tile_X3Y5_EE4BEG[9] ,
    \Tile_X3Y5_EE4BEG[8] ,
    \Tile_X3Y5_EE4BEG[7] ,
    \Tile_X3Y5_EE4BEG[6] ,
    \Tile_X3Y5_EE4BEG[5] ,
    \Tile_X3Y5_EE4BEG[4] ,
    \Tile_X3Y5_EE4BEG[3] ,
    \Tile_X3Y5_EE4BEG[2] ,
    \Tile_X3Y5_EE4BEG[1] ,
    \Tile_X3Y5_EE4BEG[0] }),
    .FrameData({\Tile_X3Y5_FrameData_O[31] ,
    \Tile_X3Y5_FrameData_O[30] ,
    \Tile_X3Y5_FrameData_O[29] ,
    \Tile_X3Y5_FrameData_O[28] ,
    \Tile_X3Y5_FrameData_O[27] ,
    \Tile_X3Y5_FrameData_O[26] ,
    \Tile_X3Y5_FrameData_O[25] ,
    \Tile_X3Y5_FrameData_O[24] ,
    \Tile_X3Y5_FrameData_O[23] ,
    \Tile_X3Y5_FrameData_O[22] ,
    \Tile_X3Y5_FrameData_O[21] ,
    \Tile_X3Y5_FrameData_O[20] ,
    \Tile_X3Y5_FrameData_O[19] ,
    \Tile_X3Y5_FrameData_O[18] ,
    \Tile_X3Y5_FrameData_O[17] ,
    \Tile_X3Y5_FrameData_O[16] ,
    \Tile_X3Y5_FrameData_O[15] ,
    \Tile_X3Y5_FrameData_O[14] ,
    \Tile_X3Y5_FrameData_O[13] ,
    \Tile_X3Y5_FrameData_O[12] ,
    \Tile_X3Y5_FrameData_O[11] ,
    \Tile_X3Y5_FrameData_O[10] ,
    \Tile_X3Y5_FrameData_O[9] ,
    \Tile_X3Y5_FrameData_O[8] ,
    \Tile_X3Y5_FrameData_O[7] ,
    \Tile_X3Y5_FrameData_O[6] ,
    \Tile_X3Y5_FrameData_O[5] ,
    \Tile_X3Y5_FrameData_O[4] ,
    \Tile_X3Y5_FrameData_O[3] ,
    \Tile_X3Y5_FrameData_O[2] ,
    \Tile_X3Y5_FrameData_O[1] ,
    \Tile_X3Y5_FrameData_O[0] }),
    .FrameData_O({\Tile_X4Y5_FrameData_O[31] ,
    \Tile_X4Y5_FrameData_O[30] ,
    \Tile_X4Y5_FrameData_O[29] ,
    \Tile_X4Y5_FrameData_O[28] ,
    \Tile_X4Y5_FrameData_O[27] ,
    \Tile_X4Y5_FrameData_O[26] ,
    \Tile_X4Y5_FrameData_O[25] ,
    \Tile_X4Y5_FrameData_O[24] ,
    \Tile_X4Y5_FrameData_O[23] ,
    \Tile_X4Y5_FrameData_O[22] ,
    \Tile_X4Y5_FrameData_O[21] ,
    \Tile_X4Y5_FrameData_O[20] ,
    \Tile_X4Y5_FrameData_O[19] ,
    \Tile_X4Y5_FrameData_O[18] ,
    \Tile_X4Y5_FrameData_O[17] ,
    \Tile_X4Y5_FrameData_O[16] ,
    \Tile_X4Y5_FrameData_O[15] ,
    \Tile_X4Y5_FrameData_O[14] ,
    \Tile_X4Y5_FrameData_O[13] ,
    \Tile_X4Y5_FrameData_O[12] ,
    \Tile_X4Y5_FrameData_O[11] ,
    \Tile_X4Y5_FrameData_O[10] ,
    \Tile_X4Y5_FrameData_O[9] ,
    \Tile_X4Y5_FrameData_O[8] ,
    \Tile_X4Y5_FrameData_O[7] ,
    \Tile_X4Y5_FrameData_O[6] ,
    \Tile_X4Y5_FrameData_O[5] ,
    \Tile_X4Y5_FrameData_O[4] ,
    \Tile_X4Y5_FrameData_O[3] ,
    \Tile_X4Y5_FrameData_O[2] ,
    \Tile_X4Y5_FrameData_O[1] ,
    \Tile_X4Y5_FrameData_O[0] }),
    .FrameStrobe({\Tile_X4Y6_FrameStrobe_O[19] ,
    \Tile_X4Y6_FrameStrobe_O[18] ,
    \Tile_X4Y6_FrameStrobe_O[17] ,
    \Tile_X4Y6_FrameStrobe_O[16] ,
    \Tile_X4Y6_FrameStrobe_O[15] ,
    \Tile_X4Y6_FrameStrobe_O[14] ,
    \Tile_X4Y6_FrameStrobe_O[13] ,
    \Tile_X4Y6_FrameStrobe_O[12] ,
    \Tile_X4Y6_FrameStrobe_O[11] ,
    \Tile_X4Y6_FrameStrobe_O[10] ,
    \Tile_X4Y6_FrameStrobe_O[9] ,
    \Tile_X4Y6_FrameStrobe_O[8] ,
    \Tile_X4Y6_FrameStrobe_O[7] ,
    \Tile_X4Y6_FrameStrobe_O[6] ,
    \Tile_X4Y6_FrameStrobe_O[5] ,
    \Tile_X4Y6_FrameStrobe_O[4] ,
    \Tile_X4Y6_FrameStrobe_O[3] ,
    \Tile_X4Y6_FrameStrobe_O[2] ,
    \Tile_X4Y6_FrameStrobe_O[1] ,
    \Tile_X4Y6_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X4Y5_FrameStrobe_O[19] ,
    \Tile_X4Y5_FrameStrobe_O[18] ,
    \Tile_X4Y5_FrameStrobe_O[17] ,
    \Tile_X4Y5_FrameStrobe_O[16] ,
    \Tile_X4Y5_FrameStrobe_O[15] ,
    \Tile_X4Y5_FrameStrobe_O[14] ,
    \Tile_X4Y5_FrameStrobe_O[13] ,
    \Tile_X4Y5_FrameStrobe_O[12] ,
    \Tile_X4Y5_FrameStrobe_O[11] ,
    \Tile_X4Y5_FrameStrobe_O[10] ,
    \Tile_X4Y5_FrameStrobe_O[9] ,
    \Tile_X4Y5_FrameStrobe_O[8] ,
    \Tile_X4Y5_FrameStrobe_O[7] ,
    \Tile_X4Y5_FrameStrobe_O[6] ,
    \Tile_X4Y5_FrameStrobe_O[5] ,
    \Tile_X4Y5_FrameStrobe_O[4] ,
    \Tile_X4Y5_FrameStrobe_O[3] ,
    \Tile_X4Y5_FrameStrobe_O[2] ,
    \Tile_X4Y5_FrameStrobe_O[1] ,
    \Tile_X4Y5_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X4Y5_N1BEG[3] ,
    \Tile_X4Y5_N1BEG[2] ,
    \Tile_X4Y5_N1BEG[1] ,
    \Tile_X4Y5_N1BEG[0] }),
    .N1END({\Tile_X4Y6_N1BEG[3] ,
    \Tile_X4Y6_N1BEG[2] ,
    \Tile_X4Y6_N1BEG[1] ,
    \Tile_X4Y6_N1BEG[0] }),
    .N2BEG({\Tile_X4Y5_N2BEG[7] ,
    \Tile_X4Y5_N2BEG[6] ,
    \Tile_X4Y5_N2BEG[5] ,
    \Tile_X4Y5_N2BEG[4] ,
    \Tile_X4Y5_N2BEG[3] ,
    \Tile_X4Y5_N2BEG[2] ,
    \Tile_X4Y5_N2BEG[1] ,
    \Tile_X4Y5_N2BEG[0] }),
    .N2BEGb({\Tile_X4Y5_N2BEGb[7] ,
    \Tile_X4Y5_N2BEGb[6] ,
    \Tile_X4Y5_N2BEGb[5] ,
    \Tile_X4Y5_N2BEGb[4] ,
    \Tile_X4Y5_N2BEGb[3] ,
    \Tile_X4Y5_N2BEGb[2] ,
    \Tile_X4Y5_N2BEGb[1] ,
    \Tile_X4Y5_N2BEGb[0] }),
    .N2END({\Tile_X4Y6_N2BEGb[7] ,
    \Tile_X4Y6_N2BEGb[6] ,
    \Tile_X4Y6_N2BEGb[5] ,
    \Tile_X4Y6_N2BEGb[4] ,
    \Tile_X4Y6_N2BEGb[3] ,
    \Tile_X4Y6_N2BEGb[2] ,
    \Tile_X4Y6_N2BEGb[1] ,
    \Tile_X4Y6_N2BEGb[0] }),
    .N2MID({\Tile_X4Y6_N2BEG[7] ,
    \Tile_X4Y6_N2BEG[6] ,
    \Tile_X4Y6_N2BEG[5] ,
    \Tile_X4Y6_N2BEG[4] ,
    \Tile_X4Y6_N2BEG[3] ,
    \Tile_X4Y6_N2BEG[2] ,
    \Tile_X4Y6_N2BEG[1] ,
    \Tile_X4Y6_N2BEG[0] }),
    .N4BEG({\Tile_X4Y5_N4BEG[15] ,
    \Tile_X4Y5_N4BEG[14] ,
    \Tile_X4Y5_N4BEG[13] ,
    \Tile_X4Y5_N4BEG[12] ,
    \Tile_X4Y5_N4BEG[11] ,
    \Tile_X4Y5_N4BEG[10] ,
    \Tile_X4Y5_N4BEG[9] ,
    \Tile_X4Y5_N4BEG[8] ,
    \Tile_X4Y5_N4BEG[7] ,
    \Tile_X4Y5_N4BEG[6] ,
    \Tile_X4Y5_N4BEG[5] ,
    \Tile_X4Y5_N4BEG[4] ,
    \Tile_X4Y5_N4BEG[3] ,
    \Tile_X4Y5_N4BEG[2] ,
    \Tile_X4Y5_N4BEG[1] ,
    \Tile_X4Y5_N4BEG[0] }),
    .N4END({\Tile_X4Y6_N4BEG[15] ,
    \Tile_X4Y6_N4BEG[14] ,
    \Tile_X4Y6_N4BEG[13] ,
    \Tile_X4Y6_N4BEG[12] ,
    \Tile_X4Y6_N4BEG[11] ,
    \Tile_X4Y6_N4BEG[10] ,
    \Tile_X4Y6_N4BEG[9] ,
    \Tile_X4Y6_N4BEG[8] ,
    \Tile_X4Y6_N4BEG[7] ,
    \Tile_X4Y6_N4BEG[6] ,
    \Tile_X4Y6_N4BEG[5] ,
    \Tile_X4Y6_N4BEG[4] ,
    \Tile_X4Y6_N4BEG[3] ,
    \Tile_X4Y6_N4BEG[2] ,
    \Tile_X4Y6_N4BEG[1] ,
    \Tile_X4Y6_N4BEG[0] }),
    .NN4BEG({\Tile_X4Y5_NN4BEG[15] ,
    \Tile_X4Y5_NN4BEG[14] ,
    \Tile_X4Y5_NN4BEG[13] ,
    \Tile_X4Y5_NN4BEG[12] ,
    \Tile_X4Y5_NN4BEG[11] ,
    \Tile_X4Y5_NN4BEG[10] ,
    \Tile_X4Y5_NN4BEG[9] ,
    \Tile_X4Y5_NN4BEG[8] ,
    \Tile_X4Y5_NN4BEG[7] ,
    \Tile_X4Y5_NN4BEG[6] ,
    \Tile_X4Y5_NN4BEG[5] ,
    \Tile_X4Y5_NN4BEG[4] ,
    \Tile_X4Y5_NN4BEG[3] ,
    \Tile_X4Y5_NN4BEG[2] ,
    \Tile_X4Y5_NN4BEG[1] ,
    \Tile_X4Y5_NN4BEG[0] }),
    .NN4END({\Tile_X4Y6_NN4BEG[15] ,
    \Tile_X4Y6_NN4BEG[14] ,
    \Tile_X4Y6_NN4BEG[13] ,
    \Tile_X4Y6_NN4BEG[12] ,
    \Tile_X4Y6_NN4BEG[11] ,
    \Tile_X4Y6_NN4BEG[10] ,
    \Tile_X4Y6_NN4BEG[9] ,
    \Tile_X4Y6_NN4BEG[8] ,
    \Tile_X4Y6_NN4BEG[7] ,
    \Tile_X4Y6_NN4BEG[6] ,
    \Tile_X4Y6_NN4BEG[5] ,
    \Tile_X4Y6_NN4BEG[4] ,
    \Tile_X4Y6_NN4BEG[3] ,
    \Tile_X4Y6_NN4BEG[2] ,
    \Tile_X4Y6_NN4BEG[1] ,
    \Tile_X4Y6_NN4BEG[0] }),
    .S1BEG({\Tile_X4Y5_S1BEG[3] ,
    \Tile_X4Y5_S1BEG[2] ,
    \Tile_X4Y5_S1BEG[1] ,
    \Tile_X4Y5_S1BEG[0] }),
    .S1END({\Tile_X4Y4_S1BEG[3] ,
    \Tile_X4Y4_S1BEG[2] ,
    \Tile_X4Y4_S1BEG[1] ,
    \Tile_X4Y4_S1BEG[0] }),
    .S2BEG({\Tile_X4Y5_S2BEG[7] ,
    \Tile_X4Y5_S2BEG[6] ,
    \Tile_X4Y5_S2BEG[5] ,
    \Tile_X4Y5_S2BEG[4] ,
    \Tile_X4Y5_S2BEG[3] ,
    \Tile_X4Y5_S2BEG[2] ,
    \Tile_X4Y5_S2BEG[1] ,
    \Tile_X4Y5_S2BEG[0] }),
    .S2BEGb({\Tile_X4Y5_S2BEGb[7] ,
    \Tile_X4Y5_S2BEGb[6] ,
    \Tile_X4Y5_S2BEGb[5] ,
    \Tile_X4Y5_S2BEGb[4] ,
    \Tile_X4Y5_S2BEGb[3] ,
    \Tile_X4Y5_S2BEGb[2] ,
    \Tile_X4Y5_S2BEGb[1] ,
    \Tile_X4Y5_S2BEGb[0] }),
    .S2END({\Tile_X4Y4_S2BEGb[7] ,
    \Tile_X4Y4_S2BEGb[6] ,
    \Tile_X4Y4_S2BEGb[5] ,
    \Tile_X4Y4_S2BEGb[4] ,
    \Tile_X4Y4_S2BEGb[3] ,
    \Tile_X4Y4_S2BEGb[2] ,
    \Tile_X4Y4_S2BEGb[1] ,
    \Tile_X4Y4_S2BEGb[0] }),
    .S2MID({\Tile_X4Y4_S2BEG[7] ,
    \Tile_X4Y4_S2BEG[6] ,
    \Tile_X4Y4_S2BEG[5] ,
    \Tile_X4Y4_S2BEG[4] ,
    \Tile_X4Y4_S2BEG[3] ,
    \Tile_X4Y4_S2BEG[2] ,
    \Tile_X4Y4_S2BEG[1] ,
    \Tile_X4Y4_S2BEG[0] }),
    .S4BEG({\Tile_X4Y5_S4BEG[15] ,
    \Tile_X4Y5_S4BEG[14] ,
    \Tile_X4Y5_S4BEG[13] ,
    \Tile_X4Y5_S4BEG[12] ,
    \Tile_X4Y5_S4BEG[11] ,
    \Tile_X4Y5_S4BEG[10] ,
    \Tile_X4Y5_S4BEG[9] ,
    \Tile_X4Y5_S4BEG[8] ,
    \Tile_X4Y5_S4BEG[7] ,
    \Tile_X4Y5_S4BEG[6] ,
    \Tile_X4Y5_S4BEG[5] ,
    \Tile_X4Y5_S4BEG[4] ,
    \Tile_X4Y5_S4BEG[3] ,
    \Tile_X4Y5_S4BEG[2] ,
    \Tile_X4Y5_S4BEG[1] ,
    \Tile_X4Y5_S4BEG[0] }),
    .S4END({\Tile_X4Y4_S4BEG[15] ,
    \Tile_X4Y4_S4BEG[14] ,
    \Tile_X4Y4_S4BEG[13] ,
    \Tile_X4Y4_S4BEG[12] ,
    \Tile_X4Y4_S4BEG[11] ,
    \Tile_X4Y4_S4BEG[10] ,
    \Tile_X4Y4_S4BEG[9] ,
    \Tile_X4Y4_S4BEG[8] ,
    \Tile_X4Y4_S4BEG[7] ,
    \Tile_X4Y4_S4BEG[6] ,
    \Tile_X4Y4_S4BEG[5] ,
    \Tile_X4Y4_S4BEG[4] ,
    \Tile_X4Y4_S4BEG[3] ,
    \Tile_X4Y4_S4BEG[2] ,
    \Tile_X4Y4_S4BEG[1] ,
    \Tile_X4Y4_S4BEG[0] }),
    .SS4BEG({\Tile_X4Y5_SS4BEG[15] ,
    \Tile_X4Y5_SS4BEG[14] ,
    \Tile_X4Y5_SS4BEG[13] ,
    \Tile_X4Y5_SS4BEG[12] ,
    \Tile_X4Y5_SS4BEG[11] ,
    \Tile_X4Y5_SS4BEG[10] ,
    \Tile_X4Y5_SS4BEG[9] ,
    \Tile_X4Y5_SS4BEG[8] ,
    \Tile_X4Y5_SS4BEG[7] ,
    \Tile_X4Y5_SS4BEG[6] ,
    \Tile_X4Y5_SS4BEG[5] ,
    \Tile_X4Y5_SS4BEG[4] ,
    \Tile_X4Y5_SS4BEG[3] ,
    \Tile_X4Y5_SS4BEG[2] ,
    \Tile_X4Y5_SS4BEG[1] ,
    \Tile_X4Y5_SS4BEG[0] }),
    .SS4END({\Tile_X4Y4_SS4BEG[15] ,
    \Tile_X4Y4_SS4BEG[14] ,
    \Tile_X4Y4_SS4BEG[13] ,
    \Tile_X4Y4_SS4BEG[12] ,
    \Tile_X4Y4_SS4BEG[11] ,
    \Tile_X4Y4_SS4BEG[10] ,
    \Tile_X4Y4_SS4BEG[9] ,
    \Tile_X4Y4_SS4BEG[8] ,
    \Tile_X4Y4_SS4BEG[7] ,
    \Tile_X4Y4_SS4BEG[6] ,
    \Tile_X4Y4_SS4BEG[5] ,
    \Tile_X4Y4_SS4BEG[4] ,
    \Tile_X4Y4_SS4BEG[3] ,
    \Tile_X4Y4_SS4BEG[2] ,
    \Tile_X4Y4_SS4BEG[1] ,
    \Tile_X4Y4_SS4BEG[0] }),
    .W1BEG({\Tile_X4Y5_W1BEG[3] ,
    \Tile_X4Y5_W1BEG[2] ,
    \Tile_X4Y5_W1BEG[1] ,
    \Tile_X4Y5_W1BEG[0] }),
    .W1END({\Tile_X5Y5_W1BEG[3] ,
    \Tile_X5Y5_W1BEG[2] ,
    \Tile_X5Y5_W1BEG[1] ,
    \Tile_X5Y5_W1BEG[0] }),
    .W2BEG({\Tile_X4Y5_W2BEG[7] ,
    \Tile_X4Y5_W2BEG[6] ,
    \Tile_X4Y5_W2BEG[5] ,
    \Tile_X4Y5_W2BEG[4] ,
    \Tile_X4Y5_W2BEG[3] ,
    \Tile_X4Y5_W2BEG[2] ,
    \Tile_X4Y5_W2BEG[1] ,
    \Tile_X4Y5_W2BEG[0] }),
    .W2BEGb({\Tile_X4Y5_W2BEGb[7] ,
    \Tile_X4Y5_W2BEGb[6] ,
    \Tile_X4Y5_W2BEGb[5] ,
    \Tile_X4Y5_W2BEGb[4] ,
    \Tile_X4Y5_W2BEGb[3] ,
    \Tile_X4Y5_W2BEGb[2] ,
    \Tile_X4Y5_W2BEGb[1] ,
    \Tile_X4Y5_W2BEGb[0] }),
    .W2END({\Tile_X5Y5_W2BEGb[7] ,
    \Tile_X5Y5_W2BEGb[6] ,
    \Tile_X5Y5_W2BEGb[5] ,
    \Tile_X5Y5_W2BEGb[4] ,
    \Tile_X5Y5_W2BEGb[3] ,
    \Tile_X5Y5_W2BEGb[2] ,
    \Tile_X5Y5_W2BEGb[1] ,
    \Tile_X5Y5_W2BEGb[0] }),
    .W2MID({\Tile_X5Y5_W2BEG[7] ,
    \Tile_X5Y5_W2BEG[6] ,
    \Tile_X5Y5_W2BEG[5] ,
    \Tile_X5Y5_W2BEG[4] ,
    \Tile_X5Y5_W2BEG[3] ,
    \Tile_X5Y5_W2BEG[2] ,
    \Tile_X5Y5_W2BEG[1] ,
    \Tile_X5Y5_W2BEG[0] }),
    .W6BEG({\Tile_X4Y5_W6BEG[11] ,
    \Tile_X4Y5_W6BEG[10] ,
    \Tile_X4Y5_W6BEG[9] ,
    \Tile_X4Y5_W6BEG[8] ,
    \Tile_X4Y5_W6BEG[7] ,
    \Tile_X4Y5_W6BEG[6] ,
    \Tile_X4Y5_W6BEG[5] ,
    \Tile_X4Y5_W6BEG[4] ,
    \Tile_X4Y5_W6BEG[3] ,
    \Tile_X4Y5_W6BEG[2] ,
    \Tile_X4Y5_W6BEG[1] ,
    \Tile_X4Y5_W6BEG[0] }),
    .W6END({\Tile_X5Y5_W6BEG[11] ,
    \Tile_X5Y5_W6BEG[10] ,
    \Tile_X5Y5_W6BEG[9] ,
    \Tile_X5Y5_W6BEG[8] ,
    \Tile_X5Y5_W6BEG[7] ,
    \Tile_X5Y5_W6BEG[6] ,
    \Tile_X5Y5_W6BEG[5] ,
    \Tile_X5Y5_W6BEG[4] ,
    \Tile_X5Y5_W6BEG[3] ,
    \Tile_X5Y5_W6BEG[2] ,
    \Tile_X5Y5_W6BEG[1] ,
    \Tile_X5Y5_W6BEG[0] }),
    .WW4BEG({\Tile_X4Y5_WW4BEG[15] ,
    \Tile_X4Y5_WW4BEG[14] ,
    \Tile_X4Y5_WW4BEG[13] ,
    \Tile_X4Y5_WW4BEG[12] ,
    \Tile_X4Y5_WW4BEG[11] ,
    \Tile_X4Y5_WW4BEG[10] ,
    \Tile_X4Y5_WW4BEG[9] ,
    \Tile_X4Y5_WW4BEG[8] ,
    \Tile_X4Y5_WW4BEG[7] ,
    \Tile_X4Y5_WW4BEG[6] ,
    \Tile_X4Y5_WW4BEG[5] ,
    \Tile_X4Y5_WW4BEG[4] ,
    \Tile_X4Y5_WW4BEG[3] ,
    \Tile_X4Y5_WW4BEG[2] ,
    \Tile_X4Y5_WW4BEG[1] ,
    \Tile_X4Y5_WW4BEG[0] }),
    .WW4END({\Tile_X5Y5_WW4BEG[15] ,
    \Tile_X5Y5_WW4BEG[14] ,
    \Tile_X5Y5_WW4BEG[13] ,
    \Tile_X5Y5_WW4BEG[12] ,
    \Tile_X5Y5_WW4BEG[11] ,
    \Tile_X5Y5_WW4BEG[10] ,
    \Tile_X5Y5_WW4BEG[9] ,
    \Tile_X5Y5_WW4BEG[8] ,
    \Tile_X5Y5_WW4BEG[7] ,
    \Tile_X5Y5_WW4BEG[6] ,
    \Tile_X5Y5_WW4BEG[5] ,
    \Tile_X5Y5_WW4BEG[4] ,
    \Tile_X5Y5_WW4BEG[3] ,
    \Tile_X5Y5_WW4BEG[2] ,
    \Tile_X5Y5_WW4BEG[1] ,
    \Tile_X5Y5_WW4BEG[0] }));
 RegFile Tile_X4Y6_RegFile (.UserCLK(Tile_X4Y7_UserCLKo),
    .UserCLKo(Tile_X4Y6_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X4Y6_E1BEG[3] ,
    \Tile_X4Y6_E1BEG[2] ,
    \Tile_X4Y6_E1BEG[1] ,
    \Tile_X4Y6_E1BEG[0] }),
    .E1END({\Tile_X3Y6_E1BEG[3] ,
    \Tile_X3Y6_E1BEG[2] ,
    \Tile_X3Y6_E1BEG[1] ,
    \Tile_X3Y6_E1BEG[0] }),
    .E2BEG({\Tile_X4Y6_E2BEG[7] ,
    \Tile_X4Y6_E2BEG[6] ,
    \Tile_X4Y6_E2BEG[5] ,
    \Tile_X4Y6_E2BEG[4] ,
    \Tile_X4Y6_E2BEG[3] ,
    \Tile_X4Y6_E2BEG[2] ,
    \Tile_X4Y6_E2BEG[1] ,
    \Tile_X4Y6_E2BEG[0] }),
    .E2BEGb({\Tile_X4Y6_E2BEGb[7] ,
    \Tile_X4Y6_E2BEGb[6] ,
    \Tile_X4Y6_E2BEGb[5] ,
    \Tile_X4Y6_E2BEGb[4] ,
    \Tile_X4Y6_E2BEGb[3] ,
    \Tile_X4Y6_E2BEGb[2] ,
    \Tile_X4Y6_E2BEGb[1] ,
    \Tile_X4Y6_E2BEGb[0] }),
    .E2END({\Tile_X3Y6_E2BEGb[7] ,
    \Tile_X3Y6_E2BEGb[6] ,
    \Tile_X3Y6_E2BEGb[5] ,
    \Tile_X3Y6_E2BEGb[4] ,
    \Tile_X3Y6_E2BEGb[3] ,
    \Tile_X3Y6_E2BEGb[2] ,
    \Tile_X3Y6_E2BEGb[1] ,
    \Tile_X3Y6_E2BEGb[0] }),
    .E2MID({\Tile_X3Y6_E2BEG[7] ,
    \Tile_X3Y6_E2BEG[6] ,
    \Tile_X3Y6_E2BEG[5] ,
    \Tile_X3Y6_E2BEG[4] ,
    \Tile_X3Y6_E2BEG[3] ,
    \Tile_X3Y6_E2BEG[2] ,
    \Tile_X3Y6_E2BEG[1] ,
    \Tile_X3Y6_E2BEG[0] }),
    .E6BEG({\Tile_X4Y6_E6BEG[11] ,
    \Tile_X4Y6_E6BEG[10] ,
    \Tile_X4Y6_E6BEG[9] ,
    \Tile_X4Y6_E6BEG[8] ,
    \Tile_X4Y6_E6BEG[7] ,
    \Tile_X4Y6_E6BEG[6] ,
    \Tile_X4Y6_E6BEG[5] ,
    \Tile_X4Y6_E6BEG[4] ,
    \Tile_X4Y6_E6BEG[3] ,
    \Tile_X4Y6_E6BEG[2] ,
    \Tile_X4Y6_E6BEG[1] ,
    \Tile_X4Y6_E6BEG[0] }),
    .E6END({\Tile_X3Y6_E6BEG[11] ,
    \Tile_X3Y6_E6BEG[10] ,
    \Tile_X3Y6_E6BEG[9] ,
    \Tile_X3Y6_E6BEG[8] ,
    \Tile_X3Y6_E6BEG[7] ,
    \Tile_X3Y6_E6BEG[6] ,
    \Tile_X3Y6_E6BEG[5] ,
    \Tile_X3Y6_E6BEG[4] ,
    \Tile_X3Y6_E6BEG[3] ,
    \Tile_X3Y6_E6BEG[2] ,
    \Tile_X3Y6_E6BEG[1] ,
    \Tile_X3Y6_E6BEG[0] }),
    .EE4BEG({\Tile_X4Y6_EE4BEG[15] ,
    \Tile_X4Y6_EE4BEG[14] ,
    \Tile_X4Y6_EE4BEG[13] ,
    \Tile_X4Y6_EE4BEG[12] ,
    \Tile_X4Y6_EE4BEG[11] ,
    \Tile_X4Y6_EE4BEG[10] ,
    \Tile_X4Y6_EE4BEG[9] ,
    \Tile_X4Y6_EE4BEG[8] ,
    \Tile_X4Y6_EE4BEG[7] ,
    \Tile_X4Y6_EE4BEG[6] ,
    \Tile_X4Y6_EE4BEG[5] ,
    \Tile_X4Y6_EE4BEG[4] ,
    \Tile_X4Y6_EE4BEG[3] ,
    \Tile_X4Y6_EE4BEG[2] ,
    \Tile_X4Y6_EE4BEG[1] ,
    \Tile_X4Y6_EE4BEG[0] }),
    .EE4END({\Tile_X3Y6_EE4BEG[15] ,
    \Tile_X3Y6_EE4BEG[14] ,
    \Tile_X3Y6_EE4BEG[13] ,
    \Tile_X3Y6_EE4BEG[12] ,
    \Tile_X3Y6_EE4BEG[11] ,
    \Tile_X3Y6_EE4BEG[10] ,
    \Tile_X3Y6_EE4BEG[9] ,
    \Tile_X3Y6_EE4BEG[8] ,
    \Tile_X3Y6_EE4BEG[7] ,
    \Tile_X3Y6_EE4BEG[6] ,
    \Tile_X3Y6_EE4BEG[5] ,
    \Tile_X3Y6_EE4BEG[4] ,
    \Tile_X3Y6_EE4BEG[3] ,
    \Tile_X3Y6_EE4BEG[2] ,
    \Tile_X3Y6_EE4BEG[1] ,
    \Tile_X3Y6_EE4BEG[0] }),
    .FrameData({\Tile_X3Y6_FrameData_O[31] ,
    \Tile_X3Y6_FrameData_O[30] ,
    \Tile_X3Y6_FrameData_O[29] ,
    \Tile_X3Y6_FrameData_O[28] ,
    \Tile_X3Y6_FrameData_O[27] ,
    \Tile_X3Y6_FrameData_O[26] ,
    \Tile_X3Y6_FrameData_O[25] ,
    \Tile_X3Y6_FrameData_O[24] ,
    \Tile_X3Y6_FrameData_O[23] ,
    \Tile_X3Y6_FrameData_O[22] ,
    \Tile_X3Y6_FrameData_O[21] ,
    \Tile_X3Y6_FrameData_O[20] ,
    \Tile_X3Y6_FrameData_O[19] ,
    \Tile_X3Y6_FrameData_O[18] ,
    \Tile_X3Y6_FrameData_O[17] ,
    \Tile_X3Y6_FrameData_O[16] ,
    \Tile_X3Y6_FrameData_O[15] ,
    \Tile_X3Y6_FrameData_O[14] ,
    \Tile_X3Y6_FrameData_O[13] ,
    \Tile_X3Y6_FrameData_O[12] ,
    \Tile_X3Y6_FrameData_O[11] ,
    \Tile_X3Y6_FrameData_O[10] ,
    \Tile_X3Y6_FrameData_O[9] ,
    \Tile_X3Y6_FrameData_O[8] ,
    \Tile_X3Y6_FrameData_O[7] ,
    \Tile_X3Y6_FrameData_O[6] ,
    \Tile_X3Y6_FrameData_O[5] ,
    \Tile_X3Y6_FrameData_O[4] ,
    \Tile_X3Y6_FrameData_O[3] ,
    \Tile_X3Y6_FrameData_O[2] ,
    \Tile_X3Y6_FrameData_O[1] ,
    \Tile_X3Y6_FrameData_O[0] }),
    .FrameData_O({\Tile_X4Y6_FrameData_O[31] ,
    \Tile_X4Y6_FrameData_O[30] ,
    \Tile_X4Y6_FrameData_O[29] ,
    \Tile_X4Y6_FrameData_O[28] ,
    \Tile_X4Y6_FrameData_O[27] ,
    \Tile_X4Y6_FrameData_O[26] ,
    \Tile_X4Y6_FrameData_O[25] ,
    \Tile_X4Y6_FrameData_O[24] ,
    \Tile_X4Y6_FrameData_O[23] ,
    \Tile_X4Y6_FrameData_O[22] ,
    \Tile_X4Y6_FrameData_O[21] ,
    \Tile_X4Y6_FrameData_O[20] ,
    \Tile_X4Y6_FrameData_O[19] ,
    \Tile_X4Y6_FrameData_O[18] ,
    \Tile_X4Y6_FrameData_O[17] ,
    \Tile_X4Y6_FrameData_O[16] ,
    \Tile_X4Y6_FrameData_O[15] ,
    \Tile_X4Y6_FrameData_O[14] ,
    \Tile_X4Y6_FrameData_O[13] ,
    \Tile_X4Y6_FrameData_O[12] ,
    \Tile_X4Y6_FrameData_O[11] ,
    \Tile_X4Y6_FrameData_O[10] ,
    \Tile_X4Y6_FrameData_O[9] ,
    \Tile_X4Y6_FrameData_O[8] ,
    \Tile_X4Y6_FrameData_O[7] ,
    \Tile_X4Y6_FrameData_O[6] ,
    \Tile_X4Y6_FrameData_O[5] ,
    \Tile_X4Y6_FrameData_O[4] ,
    \Tile_X4Y6_FrameData_O[3] ,
    \Tile_X4Y6_FrameData_O[2] ,
    \Tile_X4Y6_FrameData_O[1] ,
    \Tile_X4Y6_FrameData_O[0] }),
    .FrameStrobe({\Tile_X4Y7_FrameStrobe_O[19] ,
    \Tile_X4Y7_FrameStrobe_O[18] ,
    \Tile_X4Y7_FrameStrobe_O[17] ,
    \Tile_X4Y7_FrameStrobe_O[16] ,
    \Tile_X4Y7_FrameStrobe_O[15] ,
    \Tile_X4Y7_FrameStrobe_O[14] ,
    \Tile_X4Y7_FrameStrobe_O[13] ,
    \Tile_X4Y7_FrameStrobe_O[12] ,
    \Tile_X4Y7_FrameStrobe_O[11] ,
    \Tile_X4Y7_FrameStrobe_O[10] ,
    \Tile_X4Y7_FrameStrobe_O[9] ,
    \Tile_X4Y7_FrameStrobe_O[8] ,
    \Tile_X4Y7_FrameStrobe_O[7] ,
    \Tile_X4Y7_FrameStrobe_O[6] ,
    \Tile_X4Y7_FrameStrobe_O[5] ,
    \Tile_X4Y7_FrameStrobe_O[4] ,
    \Tile_X4Y7_FrameStrobe_O[3] ,
    \Tile_X4Y7_FrameStrobe_O[2] ,
    \Tile_X4Y7_FrameStrobe_O[1] ,
    \Tile_X4Y7_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X4Y6_FrameStrobe_O[19] ,
    \Tile_X4Y6_FrameStrobe_O[18] ,
    \Tile_X4Y6_FrameStrobe_O[17] ,
    \Tile_X4Y6_FrameStrobe_O[16] ,
    \Tile_X4Y6_FrameStrobe_O[15] ,
    \Tile_X4Y6_FrameStrobe_O[14] ,
    \Tile_X4Y6_FrameStrobe_O[13] ,
    \Tile_X4Y6_FrameStrobe_O[12] ,
    \Tile_X4Y6_FrameStrobe_O[11] ,
    \Tile_X4Y6_FrameStrobe_O[10] ,
    \Tile_X4Y6_FrameStrobe_O[9] ,
    \Tile_X4Y6_FrameStrobe_O[8] ,
    \Tile_X4Y6_FrameStrobe_O[7] ,
    \Tile_X4Y6_FrameStrobe_O[6] ,
    \Tile_X4Y6_FrameStrobe_O[5] ,
    \Tile_X4Y6_FrameStrobe_O[4] ,
    \Tile_X4Y6_FrameStrobe_O[3] ,
    \Tile_X4Y6_FrameStrobe_O[2] ,
    \Tile_X4Y6_FrameStrobe_O[1] ,
    \Tile_X4Y6_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X4Y6_N1BEG[3] ,
    \Tile_X4Y6_N1BEG[2] ,
    \Tile_X4Y6_N1BEG[1] ,
    \Tile_X4Y6_N1BEG[0] }),
    .N1END({\Tile_X4Y7_N1BEG[3] ,
    \Tile_X4Y7_N1BEG[2] ,
    \Tile_X4Y7_N1BEG[1] ,
    \Tile_X4Y7_N1BEG[0] }),
    .N2BEG({\Tile_X4Y6_N2BEG[7] ,
    \Tile_X4Y6_N2BEG[6] ,
    \Tile_X4Y6_N2BEG[5] ,
    \Tile_X4Y6_N2BEG[4] ,
    \Tile_X4Y6_N2BEG[3] ,
    \Tile_X4Y6_N2BEG[2] ,
    \Tile_X4Y6_N2BEG[1] ,
    \Tile_X4Y6_N2BEG[0] }),
    .N2BEGb({\Tile_X4Y6_N2BEGb[7] ,
    \Tile_X4Y6_N2BEGb[6] ,
    \Tile_X4Y6_N2BEGb[5] ,
    \Tile_X4Y6_N2BEGb[4] ,
    \Tile_X4Y6_N2BEGb[3] ,
    \Tile_X4Y6_N2BEGb[2] ,
    \Tile_X4Y6_N2BEGb[1] ,
    \Tile_X4Y6_N2BEGb[0] }),
    .N2END({\Tile_X4Y7_N2BEGb[7] ,
    \Tile_X4Y7_N2BEGb[6] ,
    \Tile_X4Y7_N2BEGb[5] ,
    \Tile_X4Y7_N2BEGb[4] ,
    \Tile_X4Y7_N2BEGb[3] ,
    \Tile_X4Y7_N2BEGb[2] ,
    \Tile_X4Y7_N2BEGb[1] ,
    \Tile_X4Y7_N2BEGb[0] }),
    .N2MID({\Tile_X4Y7_N2BEG[7] ,
    \Tile_X4Y7_N2BEG[6] ,
    \Tile_X4Y7_N2BEG[5] ,
    \Tile_X4Y7_N2BEG[4] ,
    \Tile_X4Y7_N2BEG[3] ,
    \Tile_X4Y7_N2BEG[2] ,
    \Tile_X4Y7_N2BEG[1] ,
    \Tile_X4Y7_N2BEG[0] }),
    .N4BEG({\Tile_X4Y6_N4BEG[15] ,
    \Tile_X4Y6_N4BEG[14] ,
    \Tile_X4Y6_N4BEG[13] ,
    \Tile_X4Y6_N4BEG[12] ,
    \Tile_X4Y6_N4BEG[11] ,
    \Tile_X4Y6_N4BEG[10] ,
    \Tile_X4Y6_N4BEG[9] ,
    \Tile_X4Y6_N4BEG[8] ,
    \Tile_X4Y6_N4BEG[7] ,
    \Tile_X4Y6_N4BEG[6] ,
    \Tile_X4Y6_N4BEG[5] ,
    \Tile_X4Y6_N4BEG[4] ,
    \Tile_X4Y6_N4BEG[3] ,
    \Tile_X4Y6_N4BEG[2] ,
    \Tile_X4Y6_N4BEG[1] ,
    \Tile_X4Y6_N4BEG[0] }),
    .N4END({\Tile_X4Y7_N4BEG[15] ,
    \Tile_X4Y7_N4BEG[14] ,
    \Tile_X4Y7_N4BEG[13] ,
    \Tile_X4Y7_N4BEG[12] ,
    \Tile_X4Y7_N4BEG[11] ,
    \Tile_X4Y7_N4BEG[10] ,
    \Tile_X4Y7_N4BEG[9] ,
    \Tile_X4Y7_N4BEG[8] ,
    \Tile_X4Y7_N4BEG[7] ,
    \Tile_X4Y7_N4BEG[6] ,
    \Tile_X4Y7_N4BEG[5] ,
    \Tile_X4Y7_N4BEG[4] ,
    \Tile_X4Y7_N4BEG[3] ,
    \Tile_X4Y7_N4BEG[2] ,
    \Tile_X4Y7_N4BEG[1] ,
    \Tile_X4Y7_N4BEG[0] }),
    .NN4BEG({\Tile_X4Y6_NN4BEG[15] ,
    \Tile_X4Y6_NN4BEG[14] ,
    \Tile_X4Y6_NN4BEG[13] ,
    \Tile_X4Y6_NN4BEG[12] ,
    \Tile_X4Y6_NN4BEG[11] ,
    \Tile_X4Y6_NN4BEG[10] ,
    \Tile_X4Y6_NN4BEG[9] ,
    \Tile_X4Y6_NN4BEG[8] ,
    \Tile_X4Y6_NN4BEG[7] ,
    \Tile_X4Y6_NN4BEG[6] ,
    \Tile_X4Y6_NN4BEG[5] ,
    \Tile_X4Y6_NN4BEG[4] ,
    \Tile_X4Y6_NN4BEG[3] ,
    \Tile_X4Y6_NN4BEG[2] ,
    \Tile_X4Y6_NN4BEG[1] ,
    \Tile_X4Y6_NN4BEG[0] }),
    .NN4END({\Tile_X4Y7_NN4BEG[15] ,
    \Tile_X4Y7_NN4BEG[14] ,
    \Tile_X4Y7_NN4BEG[13] ,
    \Tile_X4Y7_NN4BEG[12] ,
    \Tile_X4Y7_NN4BEG[11] ,
    \Tile_X4Y7_NN4BEG[10] ,
    \Tile_X4Y7_NN4BEG[9] ,
    \Tile_X4Y7_NN4BEG[8] ,
    \Tile_X4Y7_NN4BEG[7] ,
    \Tile_X4Y7_NN4BEG[6] ,
    \Tile_X4Y7_NN4BEG[5] ,
    \Tile_X4Y7_NN4BEG[4] ,
    \Tile_X4Y7_NN4BEG[3] ,
    \Tile_X4Y7_NN4BEG[2] ,
    \Tile_X4Y7_NN4BEG[1] ,
    \Tile_X4Y7_NN4BEG[0] }),
    .S1BEG({\Tile_X4Y6_S1BEG[3] ,
    \Tile_X4Y6_S1BEG[2] ,
    \Tile_X4Y6_S1BEG[1] ,
    \Tile_X4Y6_S1BEG[0] }),
    .S1END({\Tile_X4Y5_S1BEG[3] ,
    \Tile_X4Y5_S1BEG[2] ,
    \Tile_X4Y5_S1BEG[1] ,
    \Tile_X4Y5_S1BEG[0] }),
    .S2BEG({\Tile_X4Y6_S2BEG[7] ,
    \Tile_X4Y6_S2BEG[6] ,
    \Tile_X4Y6_S2BEG[5] ,
    \Tile_X4Y6_S2BEG[4] ,
    \Tile_X4Y6_S2BEG[3] ,
    \Tile_X4Y6_S2BEG[2] ,
    \Tile_X4Y6_S2BEG[1] ,
    \Tile_X4Y6_S2BEG[0] }),
    .S2BEGb({\Tile_X4Y6_S2BEGb[7] ,
    \Tile_X4Y6_S2BEGb[6] ,
    \Tile_X4Y6_S2BEGb[5] ,
    \Tile_X4Y6_S2BEGb[4] ,
    \Tile_X4Y6_S2BEGb[3] ,
    \Tile_X4Y6_S2BEGb[2] ,
    \Tile_X4Y6_S2BEGb[1] ,
    \Tile_X4Y6_S2BEGb[0] }),
    .S2END({\Tile_X4Y5_S2BEGb[7] ,
    \Tile_X4Y5_S2BEGb[6] ,
    \Tile_X4Y5_S2BEGb[5] ,
    \Tile_X4Y5_S2BEGb[4] ,
    \Tile_X4Y5_S2BEGb[3] ,
    \Tile_X4Y5_S2BEGb[2] ,
    \Tile_X4Y5_S2BEGb[1] ,
    \Tile_X4Y5_S2BEGb[0] }),
    .S2MID({\Tile_X4Y5_S2BEG[7] ,
    \Tile_X4Y5_S2BEG[6] ,
    \Tile_X4Y5_S2BEG[5] ,
    \Tile_X4Y5_S2BEG[4] ,
    \Tile_X4Y5_S2BEG[3] ,
    \Tile_X4Y5_S2BEG[2] ,
    \Tile_X4Y5_S2BEG[1] ,
    \Tile_X4Y5_S2BEG[0] }),
    .S4BEG({\Tile_X4Y6_S4BEG[15] ,
    \Tile_X4Y6_S4BEG[14] ,
    \Tile_X4Y6_S4BEG[13] ,
    \Tile_X4Y6_S4BEG[12] ,
    \Tile_X4Y6_S4BEG[11] ,
    \Tile_X4Y6_S4BEG[10] ,
    \Tile_X4Y6_S4BEG[9] ,
    \Tile_X4Y6_S4BEG[8] ,
    \Tile_X4Y6_S4BEG[7] ,
    \Tile_X4Y6_S4BEG[6] ,
    \Tile_X4Y6_S4BEG[5] ,
    \Tile_X4Y6_S4BEG[4] ,
    \Tile_X4Y6_S4BEG[3] ,
    \Tile_X4Y6_S4BEG[2] ,
    \Tile_X4Y6_S4BEG[1] ,
    \Tile_X4Y6_S4BEG[0] }),
    .S4END({\Tile_X4Y5_S4BEG[15] ,
    \Tile_X4Y5_S4BEG[14] ,
    \Tile_X4Y5_S4BEG[13] ,
    \Tile_X4Y5_S4BEG[12] ,
    \Tile_X4Y5_S4BEG[11] ,
    \Tile_X4Y5_S4BEG[10] ,
    \Tile_X4Y5_S4BEG[9] ,
    \Tile_X4Y5_S4BEG[8] ,
    \Tile_X4Y5_S4BEG[7] ,
    \Tile_X4Y5_S4BEG[6] ,
    \Tile_X4Y5_S4BEG[5] ,
    \Tile_X4Y5_S4BEG[4] ,
    \Tile_X4Y5_S4BEG[3] ,
    \Tile_X4Y5_S4BEG[2] ,
    \Tile_X4Y5_S4BEG[1] ,
    \Tile_X4Y5_S4BEG[0] }),
    .SS4BEG({\Tile_X4Y6_SS4BEG[15] ,
    \Tile_X4Y6_SS4BEG[14] ,
    \Tile_X4Y6_SS4BEG[13] ,
    \Tile_X4Y6_SS4BEG[12] ,
    \Tile_X4Y6_SS4BEG[11] ,
    \Tile_X4Y6_SS4BEG[10] ,
    \Tile_X4Y6_SS4BEG[9] ,
    \Tile_X4Y6_SS4BEG[8] ,
    \Tile_X4Y6_SS4BEG[7] ,
    \Tile_X4Y6_SS4BEG[6] ,
    \Tile_X4Y6_SS4BEG[5] ,
    \Tile_X4Y6_SS4BEG[4] ,
    \Tile_X4Y6_SS4BEG[3] ,
    \Tile_X4Y6_SS4BEG[2] ,
    \Tile_X4Y6_SS4BEG[1] ,
    \Tile_X4Y6_SS4BEG[0] }),
    .SS4END({\Tile_X4Y5_SS4BEG[15] ,
    \Tile_X4Y5_SS4BEG[14] ,
    \Tile_X4Y5_SS4BEG[13] ,
    \Tile_X4Y5_SS4BEG[12] ,
    \Tile_X4Y5_SS4BEG[11] ,
    \Tile_X4Y5_SS4BEG[10] ,
    \Tile_X4Y5_SS4BEG[9] ,
    \Tile_X4Y5_SS4BEG[8] ,
    \Tile_X4Y5_SS4BEG[7] ,
    \Tile_X4Y5_SS4BEG[6] ,
    \Tile_X4Y5_SS4BEG[5] ,
    \Tile_X4Y5_SS4BEG[4] ,
    \Tile_X4Y5_SS4BEG[3] ,
    \Tile_X4Y5_SS4BEG[2] ,
    \Tile_X4Y5_SS4BEG[1] ,
    \Tile_X4Y5_SS4BEG[0] }),
    .W1BEG({\Tile_X4Y6_W1BEG[3] ,
    \Tile_X4Y6_W1BEG[2] ,
    \Tile_X4Y6_W1BEG[1] ,
    \Tile_X4Y6_W1BEG[0] }),
    .W1END({\Tile_X5Y6_W1BEG[3] ,
    \Tile_X5Y6_W1BEG[2] ,
    \Tile_X5Y6_W1BEG[1] ,
    \Tile_X5Y6_W1BEG[0] }),
    .W2BEG({\Tile_X4Y6_W2BEG[7] ,
    \Tile_X4Y6_W2BEG[6] ,
    \Tile_X4Y6_W2BEG[5] ,
    \Tile_X4Y6_W2BEG[4] ,
    \Tile_X4Y6_W2BEG[3] ,
    \Tile_X4Y6_W2BEG[2] ,
    \Tile_X4Y6_W2BEG[1] ,
    \Tile_X4Y6_W2BEG[0] }),
    .W2BEGb({\Tile_X4Y6_W2BEGb[7] ,
    \Tile_X4Y6_W2BEGb[6] ,
    \Tile_X4Y6_W2BEGb[5] ,
    \Tile_X4Y6_W2BEGb[4] ,
    \Tile_X4Y6_W2BEGb[3] ,
    \Tile_X4Y6_W2BEGb[2] ,
    \Tile_X4Y6_W2BEGb[1] ,
    \Tile_X4Y6_W2BEGb[0] }),
    .W2END({\Tile_X5Y6_W2BEGb[7] ,
    \Tile_X5Y6_W2BEGb[6] ,
    \Tile_X5Y6_W2BEGb[5] ,
    \Tile_X5Y6_W2BEGb[4] ,
    \Tile_X5Y6_W2BEGb[3] ,
    \Tile_X5Y6_W2BEGb[2] ,
    \Tile_X5Y6_W2BEGb[1] ,
    \Tile_X5Y6_W2BEGb[0] }),
    .W2MID({\Tile_X5Y6_W2BEG[7] ,
    \Tile_X5Y6_W2BEG[6] ,
    \Tile_X5Y6_W2BEG[5] ,
    \Tile_X5Y6_W2BEG[4] ,
    \Tile_X5Y6_W2BEG[3] ,
    \Tile_X5Y6_W2BEG[2] ,
    \Tile_X5Y6_W2BEG[1] ,
    \Tile_X5Y6_W2BEG[0] }),
    .W6BEG({\Tile_X4Y6_W6BEG[11] ,
    \Tile_X4Y6_W6BEG[10] ,
    \Tile_X4Y6_W6BEG[9] ,
    \Tile_X4Y6_W6BEG[8] ,
    \Tile_X4Y6_W6BEG[7] ,
    \Tile_X4Y6_W6BEG[6] ,
    \Tile_X4Y6_W6BEG[5] ,
    \Tile_X4Y6_W6BEG[4] ,
    \Tile_X4Y6_W6BEG[3] ,
    \Tile_X4Y6_W6BEG[2] ,
    \Tile_X4Y6_W6BEG[1] ,
    \Tile_X4Y6_W6BEG[0] }),
    .W6END({\Tile_X5Y6_W6BEG[11] ,
    \Tile_X5Y6_W6BEG[10] ,
    \Tile_X5Y6_W6BEG[9] ,
    \Tile_X5Y6_W6BEG[8] ,
    \Tile_X5Y6_W6BEG[7] ,
    \Tile_X5Y6_W6BEG[6] ,
    \Tile_X5Y6_W6BEG[5] ,
    \Tile_X5Y6_W6BEG[4] ,
    \Tile_X5Y6_W6BEG[3] ,
    \Tile_X5Y6_W6BEG[2] ,
    \Tile_X5Y6_W6BEG[1] ,
    \Tile_X5Y6_W6BEG[0] }),
    .WW4BEG({\Tile_X4Y6_WW4BEG[15] ,
    \Tile_X4Y6_WW4BEG[14] ,
    \Tile_X4Y6_WW4BEG[13] ,
    \Tile_X4Y6_WW4BEG[12] ,
    \Tile_X4Y6_WW4BEG[11] ,
    \Tile_X4Y6_WW4BEG[10] ,
    \Tile_X4Y6_WW4BEG[9] ,
    \Tile_X4Y6_WW4BEG[8] ,
    \Tile_X4Y6_WW4BEG[7] ,
    \Tile_X4Y6_WW4BEG[6] ,
    \Tile_X4Y6_WW4BEG[5] ,
    \Tile_X4Y6_WW4BEG[4] ,
    \Tile_X4Y6_WW4BEG[3] ,
    \Tile_X4Y6_WW4BEG[2] ,
    \Tile_X4Y6_WW4BEG[1] ,
    \Tile_X4Y6_WW4BEG[0] }),
    .WW4END({\Tile_X5Y6_WW4BEG[15] ,
    \Tile_X5Y6_WW4BEG[14] ,
    \Tile_X5Y6_WW4BEG[13] ,
    \Tile_X5Y6_WW4BEG[12] ,
    \Tile_X5Y6_WW4BEG[11] ,
    \Tile_X5Y6_WW4BEG[10] ,
    \Tile_X5Y6_WW4BEG[9] ,
    \Tile_X5Y6_WW4BEG[8] ,
    \Tile_X5Y6_WW4BEG[7] ,
    \Tile_X5Y6_WW4BEG[6] ,
    \Tile_X5Y6_WW4BEG[5] ,
    \Tile_X5Y6_WW4BEG[4] ,
    \Tile_X5Y6_WW4BEG[3] ,
    \Tile_X5Y6_WW4BEG[2] ,
    \Tile_X5Y6_WW4BEG[1] ,
    \Tile_X5Y6_WW4BEG[0] }));
 RegFile Tile_X4Y7_RegFile (.UserCLK(Tile_X4Y8_UserCLKo),
    .UserCLKo(Tile_X4Y7_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X4Y7_E1BEG[3] ,
    \Tile_X4Y7_E1BEG[2] ,
    \Tile_X4Y7_E1BEG[1] ,
    \Tile_X4Y7_E1BEG[0] }),
    .E1END({\Tile_X3Y7_E1BEG[3] ,
    \Tile_X3Y7_E1BEG[2] ,
    \Tile_X3Y7_E1BEG[1] ,
    \Tile_X3Y7_E1BEG[0] }),
    .E2BEG({\Tile_X4Y7_E2BEG[7] ,
    \Tile_X4Y7_E2BEG[6] ,
    \Tile_X4Y7_E2BEG[5] ,
    \Tile_X4Y7_E2BEG[4] ,
    \Tile_X4Y7_E2BEG[3] ,
    \Tile_X4Y7_E2BEG[2] ,
    \Tile_X4Y7_E2BEG[1] ,
    \Tile_X4Y7_E2BEG[0] }),
    .E2BEGb({\Tile_X4Y7_E2BEGb[7] ,
    \Tile_X4Y7_E2BEGb[6] ,
    \Tile_X4Y7_E2BEGb[5] ,
    \Tile_X4Y7_E2BEGb[4] ,
    \Tile_X4Y7_E2BEGb[3] ,
    \Tile_X4Y7_E2BEGb[2] ,
    \Tile_X4Y7_E2BEGb[1] ,
    \Tile_X4Y7_E2BEGb[0] }),
    .E2END({\Tile_X3Y7_E2BEGb[7] ,
    \Tile_X3Y7_E2BEGb[6] ,
    \Tile_X3Y7_E2BEGb[5] ,
    \Tile_X3Y7_E2BEGb[4] ,
    \Tile_X3Y7_E2BEGb[3] ,
    \Tile_X3Y7_E2BEGb[2] ,
    \Tile_X3Y7_E2BEGb[1] ,
    \Tile_X3Y7_E2BEGb[0] }),
    .E2MID({\Tile_X3Y7_E2BEG[7] ,
    \Tile_X3Y7_E2BEG[6] ,
    \Tile_X3Y7_E2BEG[5] ,
    \Tile_X3Y7_E2BEG[4] ,
    \Tile_X3Y7_E2BEG[3] ,
    \Tile_X3Y7_E2BEG[2] ,
    \Tile_X3Y7_E2BEG[1] ,
    \Tile_X3Y7_E2BEG[0] }),
    .E6BEG({\Tile_X4Y7_E6BEG[11] ,
    \Tile_X4Y7_E6BEG[10] ,
    \Tile_X4Y7_E6BEG[9] ,
    \Tile_X4Y7_E6BEG[8] ,
    \Tile_X4Y7_E6BEG[7] ,
    \Tile_X4Y7_E6BEG[6] ,
    \Tile_X4Y7_E6BEG[5] ,
    \Tile_X4Y7_E6BEG[4] ,
    \Tile_X4Y7_E6BEG[3] ,
    \Tile_X4Y7_E6BEG[2] ,
    \Tile_X4Y7_E6BEG[1] ,
    \Tile_X4Y7_E6BEG[0] }),
    .E6END({\Tile_X3Y7_E6BEG[11] ,
    \Tile_X3Y7_E6BEG[10] ,
    \Tile_X3Y7_E6BEG[9] ,
    \Tile_X3Y7_E6BEG[8] ,
    \Tile_X3Y7_E6BEG[7] ,
    \Tile_X3Y7_E6BEG[6] ,
    \Tile_X3Y7_E6BEG[5] ,
    \Tile_X3Y7_E6BEG[4] ,
    \Tile_X3Y7_E6BEG[3] ,
    \Tile_X3Y7_E6BEG[2] ,
    \Tile_X3Y7_E6BEG[1] ,
    \Tile_X3Y7_E6BEG[0] }),
    .EE4BEG({\Tile_X4Y7_EE4BEG[15] ,
    \Tile_X4Y7_EE4BEG[14] ,
    \Tile_X4Y7_EE4BEG[13] ,
    \Tile_X4Y7_EE4BEG[12] ,
    \Tile_X4Y7_EE4BEG[11] ,
    \Tile_X4Y7_EE4BEG[10] ,
    \Tile_X4Y7_EE4BEG[9] ,
    \Tile_X4Y7_EE4BEG[8] ,
    \Tile_X4Y7_EE4BEG[7] ,
    \Tile_X4Y7_EE4BEG[6] ,
    \Tile_X4Y7_EE4BEG[5] ,
    \Tile_X4Y7_EE4BEG[4] ,
    \Tile_X4Y7_EE4BEG[3] ,
    \Tile_X4Y7_EE4BEG[2] ,
    \Tile_X4Y7_EE4BEG[1] ,
    \Tile_X4Y7_EE4BEG[0] }),
    .EE4END({\Tile_X3Y7_EE4BEG[15] ,
    \Tile_X3Y7_EE4BEG[14] ,
    \Tile_X3Y7_EE4BEG[13] ,
    \Tile_X3Y7_EE4BEG[12] ,
    \Tile_X3Y7_EE4BEG[11] ,
    \Tile_X3Y7_EE4BEG[10] ,
    \Tile_X3Y7_EE4BEG[9] ,
    \Tile_X3Y7_EE4BEG[8] ,
    \Tile_X3Y7_EE4BEG[7] ,
    \Tile_X3Y7_EE4BEG[6] ,
    \Tile_X3Y7_EE4BEG[5] ,
    \Tile_X3Y7_EE4BEG[4] ,
    \Tile_X3Y7_EE4BEG[3] ,
    \Tile_X3Y7_EE4BEG[2] ,
    \Tile_X3Y7_EE4BEG[1] ,
    \Tile_X3Y7_EE4BEG[0] }),
    .FrameData({\Tile_X3Y7_FrameData_O[31] ,
    \Tile_X3Y7_FrameData_O[30] ,
    \Tile_X3Y7_FrameData_O[29] ,
    \Tile_X3Y7_FrameData_O[28] ,
    \Tile_X3Y7_FrameData_O[27] ,
    \Tile_X3Y7_FrameData_O[26] ,
    \Tile_X3Y7_FrameData_O[25] ,
    \Tile_X3Y7_FrameData_O[24] ,
    \Tile_X3Y7_FrameData_O[23] ,
    \Tile_X3Y7_FrameData_O[22] ,
    \Tile_X3Y7_FrameData_O[21] ,
    \Tile_X3Y7_FrameData_O[20] ,
    \Tile_X3Y7_FrameData_O[19] ,
    \Tile_X3Y7_FrameData_O[18] ,
    \Tile_X3Y7_FrameData_O[17] ,
    \Tile_X3Y7_FrameData_O[16] ,
    \Tile_X3Y7_FrameData_O[15] ,
    \Tile_X3Y7_FrameData_O[14] ,
    \Tile_X3Y7_FrameData_O[13] ,
    \Tile_X3Y7_FrameData_O[12] ,
    \Tile_X3Y7_FrameData_O[11] ,
    \Tile_X3Y7_FrameData_O[10] ,
    \Tile_X3Y7_FrameData_O[9] ,
    \Tile_X3Y7_FrameData_O[8] ,
    \Tile_X3Y7_FrameData_O[7] ,
    \Tile_X3Y7_FrameData_O[6] ,
    \Tile_X3Y7_FrameData_O[5] ,
    \Tile_X3Y7_FrameData_O[4] ,
    \Tile_X3Y7_FrameData_O[3] ,
    \Tile_X3Y7_FrameData_O[2] ,
    \Tile_X3Y7_FrameData_O[1] ,
    \Tile_X3Y7_FrameData_O[0] }),
    .FrameData_O({\Tile_X4Y7_FrameData_O[31] ,
    \Tile_X4Y7_FrameData_O[30] ,
    \Tile_X4Y7_FrameData_O[29] ,
    \Tile_X4Y7_FrameData_O[28] ,
    \Tile_X4Y7_FrameData_O[27] ,
    \Tile_X4Y7_FrameData_O[26] ,
    \Tile_X4Y7_FrameData_O[25] ,
    \Tile_X4Y7_FrameData_O[24] ,
    \Tile_X4Y7_FrameData_O[23] ,
    \Tile_X4Y7_FrameData_O[22] ,
    \Tile_X4Y7_FrameData_O[21] ,
    \Tile_X4Y7_FrameData_O[20] ,
    \Tile_X4Y7_FrameData_O[19] ,
    \Tile_X4Y7_FrameData_O[18] ,
    \Tile_X4Y7_FrameData_O[17] ,
    \Tile_X4Y7_FrameData_O[16] ,
    \Tile_X4Y7_FrameData_O[15] ,
    \Tile_X4Y7_FrameData_O[14] ,
    \Tile_X4Y7_FrameData_O[13] ,
    \Tile_X4Y7_FrameData_O[12] ,
    \Tile_X4Y7_FrameData_O[11] ,
    \Tile_X4Y7_FrameData_O[10] ,
    \Tile_X4Y7_FrameData_O[9] ,
    \Tile_X4Y7_FrameData_O[8] ,
    \Tile_X4Y7_FrameData_O[7] ,
    \Tile_X4Y7_FrameData_O[6] ,
    \Tile_X4Y7_FrameData_O[5] ,
    \Tile_X4Y7_FrameData_O[4] ,
    \Tile_X4Y7_FrameData_O[3] ,
    \Tile_X4Y7_FrameData_O[2] ,
    \Tile_X4Y7_FrameData_O[1] ,
    \Tile_X4Y7_FrameData_O[0] }),
    .FrameStrobe({\Tile_X4Y8_FrameStrobe_O[19] ,
    \Tile_X4Y8_FrameStrobe_O[18] ,
    \Tile_X4Y8_FrameStrobe_O[17] ,
    \Tile_X4Y8_FrameStrobe_O[16] ,
    \Tile_X4Y8_FrameStrobe_O[15] ,
    \Tile_X4Y8_FrameStrobe_O[14] ,
    \Tile_X4Y8_FrameStrobe_O[13] ,
    \Tile_X4Y8_FrameStrobe_O[12] ,
    \Tile_X4Y8_FrameStrobe_O[11] ,
    \Tile_X4Y8_FrameStrobe_O[10] ,
    \Tile_X4Y8_FrameStrobe_O[9] ,
    \Tile_X4Y8_FrameStrobe_O[8] ,
    \Tile_X4Y8_FrameStrobe_O[7] ,
    \Tile_X4Y8_FrameStrobe_O[6] ,
    \Tile_X4Y8_FrameStrobe_O[5] ,
    \Tile_X4Y8_FrameStrobe_O[4] ,
    \Tile_X4Y8_FrameStrobe_O[3] ,
    \Tile_X4Y8_FrameStrobe_O[2] ,
    \Tile_X4Y8_FrameStrobe_O[1] ,
    \Tile_X4Y8_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X4Y7_FrameStrobe_O[19] ,
    \Tile_X4Y7_FrameStrobe_O[18] ,
    \Tile_X4Y7_FrameStrobe_O[17] ,
    \Tile_X4Y7_FrameStrobe_O[16] ,
    \Tile_X4Y7_FrameStrobe_O[15] ,
    \Tile_X4Y7_FrameStrobe_O[14] ,
    \Tile_X4Y7_FrameStrobe_O[13] ,
    \Tile_X4Y7_FrameStrobe_O[12] ,
    \Tile_X4Y7_FrameStrobe_O[11] ,
    \Tile_X4Y7_FrameStrobe_O[10] ,
    \Tile_X4Y7_FrameStrobe_O[9] ,
    \Tile_X4Y7_FrameStrobe_O[8] ,
    \Tile_X4Y7_FrameStrobe_O[7] ,
    \Tile_X4Y7_FrameStrobe_O[6] ,
    \Tile_X4Y7_FrameStrobe_O[5] ,
    \Tile_X4Y7_FrameStrobe_O[4] ,
    \Tile_X4Y7_FrameStrobe_O[3] ,
    \Tile_X4Y7_FrameStrobe_O[2] ,
    \Tile_X4Y7_FrameStrobe_O[1] ,
    \Tile_X4Y7_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X4Y7_N1BEG[3] ,
    \Tile_X4Y7_N1BEG[2] ,
    \Tile_X4Y7_N1BEG[1] ,
    \Tile_X4Y7_N1BEG[0] }),
    .N1END({\Tile_X4Y8_N1BEG[3] ,
    \Tile_X4Y8_N1BEG[2] ,
    \Tile_X4Y8_N1BEG[1] ,
    \Tile_X4Y8_N1BEG[0] }),
    .N2BEG({\Tile_X4Y7_N2BEG[7] ,
    \Tile_X4Y7_N2BEG[6] ,
    \Tile_X4Y7_N2BEG[5] ,
    \Tile_X4Y7_N2BEG[4] ,
    \Tile_X4Y7_N2BEG[3] ,
    \Tile_X4Y7_N2BEG[2] ,
    \Tile_X4Y7_N2BEG[1] ,
    \Tile_X4Y7_N2BEG[0] }),
    .N2BEGb({\Tile_X4Y7_N2BEGb[7] ,
    \Tile_X4Y7_N2BEGb[6] ,
    \Tile_X4Y7_N2BEGb[5] ,
    \Tile_X4Y7_N2BEGb[4] ,
    \Tile_X4Y7_N2BEGb[3] ,
    \Tile_X4Y7_N2BEGb[2] ,
    \Tile_X4Y7_N2BEGb[1] ,
    \Tile_X4Y7_N2BEGb[0] }),
    .N2END({\Tile_X4Y8_N2BEGb[7] ,
    \Tile_X4Y8_N2BEGb[6] ,
    \Tile_X4Y8_N2BEGb[5] ,
    \Tile_X4Y8_N2BEGb[4] ,
    \Tile_X4Y8_N2BEGb[3] ,
    \Tile_X4Y8_N2BEGb[2] ,
    \Tile_X4Y8_N2BEGb[1] ,
    \Tile_X4Y8_N2BEGb[0] }),
    .N2MID({\Tile_X4Y8_N2BEG[7] ,
    \Tile_X4Y8_N2BEG[6] ,
    \Tile_X4Y8_N2BEG[5] ,
    \Tile_X4Y8_N2BEG[4] ,
    \Tile_X4Y8_N2BEG[3] ,
    \Tile_X4Y8_N2BEG[2] ,
    \Tile_X4Y8_N2BEG[1] ,
    \Tile_X4Y8_N2BEG[0] }),
    .N4BEG({\Tile_X4Y7_N4BEG[15] ,
    \Tile_X4Y7_N4BEG[14] ,
    \Tile_X4Y7_N4BEG[13] ,
    \Tile_X4Y7_N4BEG[12] ,
    \Tile_X4Y7_N4BEG[11] ,
    \Tile_X4Y7_N4BEG[10] ,
    \Tile_X4Y7_N4BEG[9] ,
    \Tile_X4Y7_N4BEG[8] ,
    \Tile_X4Y7_N4BEG[7] ,
    \Tile_X4Y7_N4BEG[6] ,
    \Tile_X4Y7_N4BEG[5] ,
    \Tile_X4Y7_N4BEG[4] ,
    \Tile_X4Y7_N4BEG[3] ,
    \Tile_X4Y7_N4BEG[2] ,
    \Tile_X4Y7_N4BEG[1] ,
    \Tile_X4Y7_N4BEG[0] }),
    .N4END({\Tile_X4Y8_N4BEG[15] ,
    \Tile_X4Y8_N4BEG[14] ,
    \Tile_X4Y8_N4BEG[13] ,
    \Tile_X4Y8_N4BEG[12] ,
    \Tile_X4Y8_N4BEG[11] ,
    \Tile_X4Y8_N4BEG[10] ,
    \Tile_X4Y8_N4BEG[9] ,
    \Tile_X4Y8_N4BEG[8] ,
    \Tile_X4Y8_N4BEG[7] ,
    \Tile_X4Y8_N4BEG[6] ,
    \Tile_X4Y8_N4BEG[5] ,
    \Tile_X4Y8_N4BEG[4] ,
    \Tile_X4Y8_N4BEG[3] ,
    \Tile_X4Y8_N4BEG[2] ,
    \Tile_X4Y8_N4BEG[1] ,
    \Tile_X4Y8_N4BEG[0] }),
    .NN4BEG({\Tile_X4Y7_NN4BEG[15] ,
    \Tile_X4Y7_NN4BEG[14] ,
    \Tile_X4Y7_NN4BEG[13] ,
    \Tile_X4Y7_NN4BEG[12] ,
    \Tile_X4Y7_NN4BEG[11] ,
    \Tile_X4Y7_NN4BEG[10] ,
    \Tile_X4Y7_NN4BEG[9] ,
    \Tile_X4Y7_NN4BEG[8] ,
    \Tile_X4Y7_NN4BEG[7] ,
    \Tile_X4Y7_NN4BEG[6] ,
    \Tile_X4Y7_NN4BEG[5] ,
    \Tile_X4Y7_NN4BEG[4] ,
    \Tile_X4Y7_NN4BEG[3] ,
    \Tile_X4Y7_NN4BEG[2] ,
    \Tile_X4Y7_NN4BEG[1] ,
    \Tile_X4Y7_NN4BEG[0] }),
    .NN4END({\Tile_X4Y8_NN4BEG[15] ,
    \Tile_X4Y8_NN4BEG[14] ,
    \Tile_X4Y8_NN4BEG[13] ,
    \Tile_X4Y8_NN4BEG[12] ,
    \Tile_X4Y8_NN4BEG[11] ,
    \Tile_X4Y8_NN4BEG[10] ,
    \Tile_X4Y8_NN4BEG[9] ,
    \Tile_X4Y8_NN4BEG[8] ,
    \Tile_X4Y8_NN4BEG[7] ,
    \Tile_X4Y8_NN4BEG[6] ,
    \Tile_X4Y8_NN4BEG[5] ,
    \Tile_X4Y8_NN4BEG[4] ,
    \Tile_X4Y8_NN4BEG[3] ,
    \Tile_X4Y8_NN4BEG[2] ,
    \Tile_X4Y8_NN4BEG[1] ,
    \Tile_X4Y8_NN4BEG[0] }),
    .S1BEG({\Tile_X4Y7_S1BEG[3] ,
    \Tile_X4Y7_S1BEG[2] ,
    \Tile_X4Y7_S1BEG[1] ,
    \Tile_X4Y7_S1BEG[0] }),
    .S1END({\Tile_X4Y6_S1BEG[3] ,
    \Tile_X4Y6_S1BEG[2] ,
    \Tile_X4Y6_S1BEG[1] ,
    \Tile_X4Y6_S1BEG[0] }),
    .S2BEG({\Tile_X4Y7_S2BEG[7] ,
    \Tile_X4Y7_S2BEG[6] ,
    \Tile_X4Y7_S2BEG[5] ,
    \Tile_X4Y7_S2BEG[4] ,
    \Tile_X4Y7_S2BEG[3] ,
    \Tile_X4Y7_S2BEG[2] ,
    \Tile_X4Y7_S2BEG[1] ,
    \Tile_X4Y7_S2BEG[0] }),
    .S2BEGb({\Tile_X4Y7_S2BEGb[7] ,
    \Tile_X4Y7_S2BEGb[6] ,
    \Tile_X4Y7_S2BEGb[5] ,
    \Tile_X4Y7_S2BEGb[4] ,
    \Tile_X4Y7_S2BEGb[3] ,
    \Tile_X4Y7_S2BEGb[2] ,
    \Tile_X4Y7_S2BEGb[1] ,
    \Tile_X4Y7_S2BEGb[0] }),
    .S2END({\Tile_X4Y6_S2BEGb[7] ,
    \Tile_X4Y6_S2BEGb[6] ,
    \Tile_X4Y6_S2BEGb[5] ,
    \Tile_X4Y6_S2BEGb[4] ,
    \Tile_X4Y6_S2BEGb[3] ,
    \Tile_X4Y6_S2BEGb[2] ,
    \Tile_X4Y6_S2BEGb[1] ,
    \Tile_X4Y6_S2BEGb[0] }),
    .S2MID({\Tile_X4Y6_S2BEG[7] ,
    \Tile_X4Y6_S2BEG[6] ,
    \Tile_X4Y6_S2BEG[5] ,
    \Tile_X4Y6_S2BEG[4] ,
    \Tile_X4Y6_S2BEG[3] ,
    \Tile_X4Y6_S2BEG[2] ,
    \Tile_X4Y6_S2BEG[1] ,
    \Tile_X4Y6_S2BEG[0] }),
    .S4BEG({\Tile_X4Y7_S4BEG[15] ,
    \Tile_X4Y7_S4BEG[14] ,
    \Tile_X4Y7_S4BEG[13] ,
    \Tile_X4Y7_S4BEG[12] ,
    \Tile_X4Y7_S4BEG[11] ,
    \Tile_X4Y7_S4BEG[10] ,
    \Tile_X4Y7_S4BEG[9] ,
    \Tile_X4Y7_S4BEG[8] ,
    \Tile_X4Y7_S4BEG[7] ,
    \Tile_X4Y7_S4BEG[6] ,
    \Tile_X4Y7_S4BEG[5] ,
    \Tile_X4Y7_S4BEG[4] ,
    \Tile_X4Y7_S4BEG[3] ,
    \Tile_X4Y7_S4BEG[2] ,
    \Tile_X4Y7_S4BEG[1] ,
    \Tile_X4Y7_S4BEG[0] }),
    .S4END({\Tile_X4Y6_S4BEG[15] ,
    \Tile_X4Y6_S4BEG[14] ,
    \Tile_X4Y6_S4BEG[13] ,
    \Tile_X4Y6_S4BEG[12] ,
    \Tile_X4Y6_S4BEG[11] ,
    \Tile_X4Y6_S4BEG[10] ,
    \Tile_X4Y6_S4BEG[9] ,
    \Tile_X4Y6_S4BEG[8] ,
    \Tile_X4Y6_S4BEG[7] ,
    \Tile_X4Y6_S4BEG[6] ,
    \Tile_X4Y6_S4BEG[5] ,
    \Tile_X4Y6_S4BEG[4] ,
    \Tile_X4Y6_S4BEG[3] ,
    \Tile_X4Y6_S4BEG[2] ,
    \Tile_X4Y6_S4BEG[1] ,
    \Tile_X4Y6_S4BEG[0] }),
    .SS4BEG({\Tile_X4Y7_SS4BEG[15] ,
    \Tile_X4Y7_SS4BEG[14] ,
    \Tile_X4Y7_SS4BEG[13] ,
    \Tile_X4Y7_SS4BEG[12] ,
    \Tile_X4Y7_SS4BEG[11] ,
    \Tile_X4Y7_SS4BEG[10] ,
    \Tile_X4Y7_SS4BEG[9] ,
    \Tile_X4Y7_SS4BEG[8] ,
    \Tile_X4Y7_SS4BEG[7] ,
    \Tile_X4Y7_SS4BEG[6] ,
    \Tile_X4Y7_SS4BEG[5] ,
    \Tile_X4Y7_SS4BEG[4] ,
    \Tile_X4Y7_SS4BEG[3] ,
    \Tile_X4Y7_SS4BEG[2] ,
    \Tile_X4Y7_SS4BEG[1] ,
    \Tile_X4Y7_SS4BEG[0] }),
    .SS4END({\Tile_X4Y6_SS4BEG[15] ,
    \Tile_X4Y6_SS4BEG[14] ,
    \Tile_X4Y6_SS4BEG[13] ,
    \Tile_X4Y6_SS4BEG[12] ,
    \Tile_X4Y6_SS4BEG[11] ,
    \Tile_X4Y6_SS4BEG[10] ,
    \Tile_X4Y6_SS4BEG[9] ,
    \Tile_X4Y6_SS4BEG[8] ,
    \Tile_X4Y6_SS4BEG[7] ,
    \Tile_X4Y6_SS4BEG[6] ,
    \Tile_X4Y6_SS4BEG[5] ,
    \Tile_X4Y6_SS4BEG[4] ,
    \Tile_X4Y6_SS4BEG[3] ,
    \Tile_X4Y6_SS4BEG[2] ,
    \Tile_X4Y6_SS4BEG[1] ,
    \Tile_X4Y6_SS4BEG[0] }),
    .W1BEG({\Tile_X4Y7_W1BEG[3] ,
    \Tile_X4Y7_W1BEG[2] ,
    \Tile_X4Y7_W1BEG[1] ,
    \Tile_X4Y7_W1BEG[0] }),
    .W1END({\Tile_X5Y7_W1BEG[3] ,
    \Tile_X5Y7_W1BEG[2] ,
    \Tile_X5Y7_W1BEG[1] ,
    \Tile_X5Y7_W1BEG[0] }),
    .W2BEG({\Tile_X4Y7_W2BEG[7] ,
    \Tile_X4Y7_W2BEG[6] ,
    \Tile_X4Y7_W2BEG[5] ,
    \Tile_X4Y7_W2BEG[4] ,
    \Tile_X4Y7_W2BEG[3] ,
    \Tile_X4Y7_W2BEG[2] ,
    \Tile_X4Y7_W2BEG[1] ,
    \Tile_X4Y7_W2BEG[0] }),
    .W2BEGb({\Tile_X4Y7_W2BEGb[7] ,
    \Tile_X4Y7_W2BEGb[6] ,
    \Tile_X4Y7_W2BEGb[5] ,
    \Tile_X4Y7_W2BEGb[4] ,
    \Tile_X4Y7_W2BEGb[3] ,
    \Tile_X4Y7_W2BEGb[2] ,
    \Tile_X4Y7_W2BEGb[1] ,
    \Tile_X4Y7_W2BEGb[0] }),
    .W2END({\Tile_X5Y7_W2BEGb[7] ,
    \Tile_X5Y7_W2BEGb[6] ,
    \Tile_X5Y7_W2BEGb[5] ,
    \Tile_X5Y7_W2BEGb[4] ,
    \Tile_X5Y7_W2BEGb[3] ,
    \Tile_X5Y7_W2BEGb[2] ,
    \Tile_X5Y7_W2BEGb[1] ,
    \Tile_X5Y7_W2BEGb[0] }),
    .W2MID({\Tile_X5Y7_W2BEG[7] ,
    \Tile_X5Y7_W2BEG[6] ,
    \Tile_X5Y7_W2BEG[5] ,
    \Tile_X5Y7_W2BEG[4] ,
    \Tile_X5Y7_W2BEG[3] ,
    \Tile_X5Y7_W2BEG[2] ,
    \Tile_X5Y7_W2BEG[1] ,
    \Tile_X5Y7_W2BEG[0] }),
    .W6BEG({\Tile_X4Y7_W6BEG[11] ,
    \Tile_X4Y7_W6BEG[10] ,
    \Tile_X4Y7_W6BEG[9] ,
    \Tile_X4Y7_W6BEG[8] ,
    \Tile_X4Y7_W6BEG[7] ,
    \Tile_X4Y7_W6BEG[6] ,
    \Tile_X4Y7_W6BEG[5] ,
    \Tile_X4Y7_W6BEG[4] ,
    \Tile_X4Y7_W6BEG[3] ,
    \Tile_X4Y7_W6BEG[2] ,
    \Tile_X4Y7_W6BEG[1] ,
    \Tile_X4Y7_W6BEG[0] }),
    .W6END({\Tile_X5Y7_W6BEG[11] ,
    \Tile_X5Y7_W6BEG[10] ,
    \Tile_X5Y7_W6BEG[9] ,
    \Tile_X5Y7_W6BEG[8] ,
    \Tile_X5Y7_W6BEG[7] ,
    \Tile_X5Y7_W6BEG[6] ,
    \Tile_X5Y7_W6BEG[5] ,
    \Tile_X5Y7_W6BEG[4] ,
    \Tile_X5Y7_W6BEG[3] ,
    \Tile_X5Y7_W6BEG[2] ,
    \Tile_X5Y7_W6BEG[1] ,
    \Tile_X5Y7_W6BEG[0] }),
    .WW4BEG({\Tile_X4Y7_WW4BEG[15] ,
    \Tile_X4Y7_WW4BEG[14] ,
    \Tile_X4Y7_WW4BEG[13] ,
    \Tile_X4Y7_WW4BEG[12] ,
    \Tile_X4Y7_WW4BEG[11] ,
    \Tile_X4Y7_WW4BEG[10] ,
    \Tile_X4Y7_WW4BEG[9] ,
    \Tile_X4Y7_WW4BEG[8] ,
    \Tile_X4Y7_WW4BEG[7] ,
    \Tile_X4Y7_WW4BEG[6] ,
    \Tile_X4Y7_WW4BEG[5] ,
    \Tile_X4Y7_WW4BEG[4] ,
    \Tile_X4Y7_WW4BEG[3] ,
    \Tile_X4Y7_WW4BEG[2] ,
    \Tile_X4Y7_WW4BEG[1] ,
    \Tile_X4Y7_WW4BEG[0] }),
    .WW4END({\Tile_X5Y7_WW4BEG[15] ,
    \Tile_X5Y7_WW4BEG[14] ,
    \Tile_X5Y7_WW4BEG[13] ,
    \Tile_X5Y7_WW4BEG[12] ,
    \Tile_X5Y7_WW4BEG[11] ,
    \Tile_X5Y7_WW4BEG[10] ,
    \Tile_X5Y7_WW4BEG[9] ,
    \Tile_X5Y7_WW4BEG[8] ,
    \Tile_X5Y7_WW4BEG[7] ,
    \Tile_X5Y7_WW4BEG[6] ,
    \Tile_X5Y7_WW4BEG[5] ,
    \Tile_X5Y7_WW4BEG[4] ,
    \Tile_X5Y7_WW4BEG[3] ,
    \Tile_X5Y7_WW4BEG[2] ,
    \Tile_X5Y7_WW4BEG[1] ,
    \Tile_X5Y7_WW4BEG[0] }));
 RegFile Tile_X4Y8_RegFile (.UserCLK(Tile_X4Y9_UserCLKo),
    .UserCLKo(Tile_X4Y8_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X4Y8_E1BEG[3] ,
    \Tile_X4Y8_E1BEG[2] ,
    \Tile_X4Y8_E1BEG[1] ,
    \Tile_X4Y8_E1BEG[0] }),
    .E1END({\Tile_X3Y8_E1BEG[3] ,
    \Tile_X3Y8_E1BEG[2] ,
    \Tile_X3Y8_E1BEG[1] ,
    \Tile_X3Y8_E1BEG[0] }),
    .E2BEG({\Tile_X4Y8_E2BEG[7] ,
    \Tile_X4Y8_E2BEG[6] ,
    \Tile_X4Y8_E2BEG[5] ,
    \Tile_X4Y8_E2BEG[4] ,
    \Tile_X4Y8_E2BEG[3] ,
    \Tile_X4Y8_E2BEG[2] ,
    \Tile_X4Y8_E2BEG[1] ,
    \Tile_X4Y8_E2BEG[0] }),
    .E2BEGb({\Tile_X4Y8_E2BEGb[7] ,
    \Tile_X4Y8_E2BEGb[6] ,
    \Tile_X4Y8_E2BEGb[5] ,
    \Tile_X4Y8_E2BEGb[4] ,
    \Tile_X4Y8_E2BEGb[3] ,
    \Tile_X4Y8_E2BEGb[2] ,
    \Tile_X4Y8_E2BEGb[1] ,
    \Tile_X4Y8_E2BEGb[0] }),
    .E2END({\Tile_X3Y8_E2BEGb[7] ,
    \Tile_X3Y8_E2BEGb[6] ,
    \Tile_X3Y8_E2BEGb[5] ,
    \Tile_X3Y8_E2BEGb[4] ,
    \Tile_X3Y8_E2BEGb[3] ,
    \Tile_X3Y8_E2BEGb[2] ,
    \Tile_X3Y8_E2BEGb[1] ,
    \Tile_X3Y8_E2BEGb[0] }),
    .E2MID({\Tile_X3Y8_E2BEG[7] ,
    \Tile_X3Y8_E2BEG[6] ,
    \Tile_X3Y8_E2BEG[5] ,
    \Tile_X3Y8_E2BEG[4] ,
    \Tile_X3Y8_E2BEG[3] ,
    \Tile_X3Y8_E2BEG[2] ,
    \Tile_X3Y8_E2BEG[1] ,
    \Tile_X3Y8_E2BEG[0] }),
    .E6BEG({\Tile_X4Y8_E6BEG[11] ,
    \Tile_X4Y8_E6BEG[10] ,
    \Tile_X4Y8_E6BEG[9] ,
    \Tile_X4Y8_E6BEG[8] ,
    \Tile_X4Y8_E6BEG[7] ,
    \Tile_X4Y8_E6BEG[6] ,
    \Tile_X4Y8_E6BEG[5] ,
    \Tile_X4Y8_E6BEG[4] ,
    \Tile_X4Y8_E6BEG[3] ,
    \Tile_X4Y8_E6BEG[2] ,
    \Tile_X4Y8_E6BEG[1] ,
    \Tile_X4Y8_E6BEG[0] }),
    .E6END({\Tile_X3Y8_E6BEG[11] ,
    \Tile_X3Y8_E6BEG[10] ,
    \Tile_X3Y8_E6BEG[9] ,
    \Tile_X3Y8_E6BEG[8] ,
    \Tile_X3Y8_E6BEG[7] ,
    \Tile_X3Y8_E6BEG[6] ,
    \Tile_X3Y8_E6BEG[5] ,
    \Tile_X3Y8_E6BEG[4] ,
    \Tile_X3Y8_E6BEG[3] ,
    \Tile_X3Y8_E6BEG[2] ,
    \Tile_X3Y8_E6BEG[1] ,
    \Tile_X3Y8_E6BEG[0] }),
    .EE4BEG({\Tile_X4Y8_EE4BEG[15] ,
    \Tile_X4Y8_EE4BEG[14] ,
    \Tile_X4Y8_EE4BEG[13] ,
    \Tile_X4Y8_EE4BEG[12] ,
    \Tile_X4Y8_EE4BEG[11] ,
    \Tile_X4Y8_EE4BEG[10] ,
    \Tile_X4Y8_EE4BEG[9] ,
    \Tile_X4Y8_EE4BEG[8] ,
    \Tile_X4Y8_EE4BEG[7] ,
    \Tile_X4Y8_EE4BEG[6] ,
    \Tile_X4Y8_EE4BEG[5] ,
    \Tile_X4Y8_EE4BEG[4] ,
    \Tile_X4Y8_EE4BEG[3] ,
    \Tile_X4Y8_EE4BEG[2] ,
    \Tile_X4Y8_EE4BEG[1] ,
    \Tile_X4Y8_EE4BEG[0] }),
    .EE4END({\Tile_X3Y8_EE4BEG[15] ,
    \Tile_X3Y8_EE4BEG[14] ,
    \Tile_X3Y8_EE4BEG[13] ,
    \Tile_X3Y8_EE4BEG[12] ,
    \Tile_X3Y8_EE4BEG[11] ,
    \Tile_X3Y8_EE4BEG[10] ,
    \Tile_X3Y8_EE4BEG[9] ,
    \Tile_X3Y8_EE4BEG[8] ,
    \Tile_X3Y8_EE4BEG[7] ,
    \Tile_X3Y8_EE4BEG[6] ,
    \Tile_X3Y8_EE4BEG[5] ,
    \Tile_X3Y8_EE4BEG[4] ,
    \Tile_X3Y8_EE4BEG[3] ,
    \Tile_X3Y8_EE4BEG[2] ,
    \Tile_X3Y8_EE4BEG[1] ,
    \Tile_X3Y8_EE4BEG[0] }),
    .FrameData({\Tile_X3Y8_FrameData_O[31] ,
    \Tile_X3Y8_FrameData_O[30] ,
    \Tile_X3Y8_FrameData_O[29] ,
    \Tile_X3Y8_FrameData_O[28] ,
    \Tile_X3Y8_FrameData_O[27] ,
    \Tile_X3Y8_FrameData_O[26] ,
    \Tile_X3Y8_FrameData_O[25] ,
    \Tile_X3Y8_FrameData_O[24] ,
    \Tile_X3Y8_FrameData_O[23] ,
    \Tile_X3Y8_FrameData_O[22] ,
    \Tile_X3Y8_FrameData_O[21] ,
    \Tile_X3Y8_FrameData_O[20] ,
    \Tile_X3Y8_FrameData_O[19] ,
    \Tile_X3Y8_FrameData_O[18] ,
    \Tile_X3Y8_FrameData_O[17] ,
    \Tile_X3Y8_FrameData_O[16] ,
    \Tile_X3Y8_FrameData_O[15] ,
    \Tile_X3Y8_FrameData_O[14] ,
    \Tile_X3Y8_FrameData_O[13] ,
    \Tile_X3Y8_FrameData_O[12] ,
    \Tile_X3Y8_FrameData_O[11] ,
    \Tile_X3Y8_FrameData_O[10] ,
    \Tile_X3Y8_FrameData_O[9] ,
    \Tile_X3Y8_FrameData_O[8] ,
    \Tile_X3Y8_FrameData_O[7] ,
    \Tile_X3Y8_FrameData_O[6] ,
    \Tile_X3Y8_FrameData_O[5] ,
    \Tile_X3Y8_FrameData_O[4] ,
    \Tile_X3Y8_FrameData_O[3] ,
    \Tile_X3Y8_FrameData_O[2] ,
    \Tile_X3Y8_FrameData_O[1] ,
    \Tile_X3Y8_FrameData_O[0] }),
    .FrameData_O({\Tile_X4Y8_FrameData_O[31] ,
    \Tile_X4Y8_FrameData_O[30] ,
    \Tile_X4Y8_FrameData_O[29] ,
    \Tile_X4Y8_FrameData_O[28] ,
    \Tile_X4Y8_FrameData_O[27] ,
    \Tile_X4Y8_FrameData_O[26] ,
    \Tile_X4Y8_FrameData_O[25] ,
    \Tile_X4Y8_FrameData_O[24] ,
    \Tile_X4Y8_FrameData_O[23] ,
    \Tile_X4Y8_FrameData_O[22] ,
    \Tile_X4Y8_FrameData_O[21] ,
    \Tile_X4Y8_FrameData_O[20] ,
    \Tile_X4Y8_FrameData_O[19] ,
    \Tile_X4Y8_FrameData_O[18] ,
    \Tile_X4Y8_FrameData_O[17] ,
    \Tile_X4Y8_FrameData_O[16] ,
    \Tile_X4Y8_FrameData_O[15] ,
    \Tile_X4Y8_FrameData_O[14] ,
    \Tile_X4Y8_FrameData_O[13] ,
    \Tile_X4Y8_FrameData_O[12] ,
    \Tile_X4Y8_FrameData_O[11] ,
    \Tile_X4Y8_FrameData_O[10] ,
    \Tile_X4Y8_FrameData_O[9] ,
    \Tile_X4Y8_FrameData_O[8] ,
    \Tile_X4Y8_FrameData_O[7] ,
    \Tile_X4Y8_FrameData_O[6] ,
    \Tile_X4Y8_FrameData_O[5] ,
    \Tile_X4Y8_FrameData_O[4] ,
    \Tile_X4Y8_FrameData_O[3] ,
    \Tile_X4Y8_FrameData_O[2] ,
    \Tile_X4Y8_FrameData_O[1] ,
    \Tile_X4Y8_FrameData_O[0] }),
    .FrameStrobe({\Tile_X4Y9_FrameStrobe_O[19] ,
    \Tile_X4Y9_FrameStrobe_O[18] ,
    \Tile_X4Y9_FrameStrobe_O[17] ,
    \Tile_X4Y9_FrameStrobe_O[16] ,
    \Tile_X4Y9_FrameStrobe_O[15] ,
    \Tile_X4Y9_FrameStrobe_O[14] ,
    \Tile_X4Y9_FrameStrobe_O[13] ,
    \Tile_X4Y9_FrameStrobe_O[12] ,
    \Tile_X4Y9_FrameStrobe_O[11] ,
    \Tile_X4Y9_FrameStrobe_O[10] ,
    \Tile_X4Y9_FrameStrobe_O[9] ,
    \Tile_X4Y9_FrameStrobe_O[8] ,
    \Tile_X4Y9_FrameStrobe_O[7] ,
    \Tile_X4Y9_FrameStrobe_O[6] ,
    \Tile_X4Y9_FrameStrobe_O[5] ,
    \Tile_X4Y9_FrameStrobe_O[4] ,
    \Tile_X4Y9_FrameStrobe_O[3] ,
    \Tile_X4Y9_FrameStrobe_O[2] ,
    \Tile_X4Y9_FrameStrobe_O[1] ,
    \Tile_X4Y9_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X4Y8_FrameStrobe_O[19] ,
    \Tile_X4Y8_FrameStrobe_O[18] ,
    \Tile_X4Y8_FrameStrobe_O[17] ,
    \Tile_X4Y8_FrameStrobe_O[16] ,
    \Tile_X4Y8_FrameStrobe_O[15] ,
    \Tile_X4Y8_FrameStrobe_O[14] ,
    \Tile_X4Y8_FrameStrobe_O[13] ,
    \Tile_X4Y8_FrameStrobe_O[12] ,
    \Tile_X4Y8_FrameStrobe_O[11] ,
    \Tile_X4Y8_FrameStrobe_O[10] ,
    \Tile_X4Y8_FrameStrobe_O[9] ,
    \Tile_X4Y8_FrameStrobe_O[8] ,
    \Tile_X4Y8_FrameStrobe_O[7] ,
    \Tile_X4Y8_FrameStrobe_O[6] ,
    \Tile_X4Y8_FrameStrobe_O[5] ,
    \Tile_X4Y8_FrameStrobe_O[4] ,
    \Tile_X4Y8_FrameStrobe_O[3] ,
    \Tile_X4Y8_FrameStrobe_O[2] ,
    \Tile_X4Y8_FrameStrobe_O[1] ,
    \Tile_X4Y8_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X4Y8_N1BEG[3] ,
    \Tile_X4Y8_N1BEG[2] ,
    \Tile_X4Y8_N1BEG[1] ,
    \Tile_X4Y8_N1BEG[0] }),
    .N1END({\Tile_X4Y9_N1BEG[3] ,
    \Tile_X4Y9_N1BEG[2] ,
    \Tile_X4Y9_N1BEG[1] ,
    \Tile_X4Y9_N1BEG[0] }),
    .N2BEG({\Tile_X4Y8_N2BEG[7] ,
    \Tile_X4Y8_N2BEG[6] ,
    \Tile_X4Y8_N2BEG[5] ,
    \Tile_X4Y8_N2BEG[4] ,
    \Tile_X4Y8_N2BEG[3] ,
    \Tile_X4Y8_N2BEG[2] ,
    \Tile_X4Y8_N2BEG[1] ,
    \Tile_X4Y8_N2BEG[0] }),
    .N2BEGb({\Tile_X4Y8_N2BEGb[7] ,
    \Tile_X4Y8_N2BEGb[6] ,
    \Tile_X4Y8_N2BEGb[5] ,
    \Tile_X4Y8_N2BEGb[4] ,
    \Tile_X4Y8_N2BEGb[3] ,
    \Tile_X4Y8_N2BEGb[2] ,
    \Tile_X4Y8_N2BEGb[1] ,
    \Tile_X4Y8_N2BEGb[0] }),
    .N2END({\Tile_X4Y9_N2BEGb[7] ,
    \Tile_X4Y9_N2BEGb[6] ,
    \Tile_X4Y9_N2BEGb[5] ,
    \Tile_X4Y9_N2BEGb[4] ,
    \Tile_X4Y9_N2BEGb[3] ,
    \Tile_X4Y9_N2BEGb[2] ,
    \Tile_X4Y9_N2BEGb[1] ,
    \Tile_X4Y9_N2BEGb[0] }),
    .N2MID({\Tile_X4Y9_N2BEG[7] ,
    \Tile_X4Y9_N2BEG[6] ,
    \Tile_X4Y9_N2BEG[5] ,
    \Tile_X4Y9_N2BEG[4] ,
    \Tile_X4Y9_N2BEG[3] ,
    \Tile_X4Y9_N2BEG[2] ,
    \Tile_X4Y9_N2BEG[1] ,
    \Tile_X4Y9_N2BEG[0] }),
    .N4BEG({\Tile_X4Y8_N4BEG[15] ,
    \Tile_X4Y8_N4BEG[14] ,
    \Tile_X4Y8_N4BEG[13] ,
    \Tile_X4Y8_N4BEG[12] ,
    \Tile_X4Y8_N4BEG[11] ,
    \Tile_X4Y8_N4BEG[10] ,
    \Tile_X4Y8_N4BEG[9] ,
    \Tile_X4Y8_N4BEG[8] ,
    \Tile_X4Y8_N4BEG[7] ,
    \Tile_X4Y8_N4BEG[6] ,
    \Tile_X4Y8_N4BEG[5] ,
    \Tile_X4Y8_N4BEG[4] ,
    \Tile_X4Y8_N4BEG[3] ,
    \Tile_X4Y8_N4BEG[2] ,
    \Tile_X4Y8_N4BEG[1] ,
    \Tile_X4Y8_N4BEG[0] }),
    .N4END({\Tile_X4Y9_N4BEG[15] ,
    \Tile_X4Y9_N4BEG[14] ,
    \Tile_X4Y9_N4BEG[13] ,
    \Tile_X4Y9_N4BEG[12] ,
    \Tile_X4Y9_N4BEG[11] ,
    \Tile_X4Y9_N4BEG[10] ,
    \Tile_X4Y9_N4BEG[9] ,
    \Tile_X4Y9_N4BEG[8] ,
    \Tile_X4Y9_N4BEG[7] ,
    \Tile_X4Y9_N4BEG[6] ,
    \Tile_X4Y9_N4BEG[5] ,
    \Tile_X4Y9_N4BEG[4] ,
    \Tile_X4Y9_N4BEG[3] ,
    \Tile_X4Y9_N4BEG[2] ,
    \Tile_X4Y9_N4BEG[1] ,
    \Tile_X4Y9_N4BEG[0] }),
    .NN4BEG({\Tile_X4Y8_NN4BEG[15] ,
    \Tile_X4Y8_NN4BEG[14] ,
    \Tile_X4Y8_NN4BEG[13] ,
    \Tile_X4Y8_NN4BEG[12] ,
    \Tile_X4Y8_NN4BEG[11] ,
    \Tile_X4Y8_NN4BEG[10] ,
    \Tile_X4Y8_NN4BEG[9] ,
    \Tile_X4Y8_NN4BEG[8] ,
    \Tile_X4Y8_NN4BEG[7] ,
    \Tile_X4Y8_NN4BEG[6] ,
    \Tile_X4Y8_NN4BEG[5] ,
    \Tile_X4Y8_NN4BEG[4] ,
    \Tile_X4Y8_NN4BEG[3] ,
    \Tile_X4Y8_NN4BEG[2] ,
    \Tile_X4Y8_NN4BEG[1] ,
    \Tile_X4Y8_NN4BEG[0] }),
    .NN4END({\Tile_X4Y9_NN4BEG[15] ,
    \Tile_X4Y9_NN4BEG[14] ,
    \Tile_X4Y9_NN4BEG[13] ,
    \Tile_X4Y9_NN4BEG[12] ,
    \Tile_X4Y9_NN4BEG[11] ,
    \Tile_X4Y9_NN4BEG[10] ,
    \Tile_X4Y9_NN4BEG[9] ,
    \Tile_X4Y9_NN4BEG[8] ,
    \Tile_X4Y9_NN4BEG[7] ,
    \Tile_X4Y9_NN4BEG[6] ,
    \Tile_X4Y9_NN4BEG[5] ,
    \Tile_X4Y9_NN4BEG[4] ,
    \Tile_X4Y9_NN4BEG[3] ,
    \Tile_X4Y9_NN4BEG[2] ,
    \Tile_X4Y9_NN4BEG[1] ,
    \Tile_X4Y9_NN4BEG[0] }),
    .S1BEG({\Tile_X4Y8_S1BEG[3] ,
    \Tile_X4Y8_S1BEG[2] ,
    \Tile_X4Y8_S1BEG[1] ,
    \Tile_X4Y8_S1BEG[0] }),
    .S1END({\Tile_X4Y7_S1BEG[3] ,
    \Tile_X4Y7_S1BEG[2] ,
    \Tile_X4Y7_S1BEG[1] ,
    \Tile_X4Y7_S1BEG[0] }),
    .S2BEG({\Tile_X4Y8_S2BEG[7] ,
    \Tile_X4Y8_S2BEG[6] ,
    \Tile_X4Y8_S2BEG[5] ,
    \Tile_X4Y8_S2BEG[4] ,
    \Tile_X4Y8_S2BEG[3] ,
    \Tile_X4Y8_S2BEG[2] ,
    \Tile_X4Y8_S2BEG[1] ,
    \Tile_X4Y8_S2BEG[0] }),
    .S2BEGb({\Tile_X4Y8_S2BEGb[7] ,
    \Tile_X4Y8_S2BEGb[6] ,
    \Tile_X4Y8_S2BEGb[5] ,
    \Tile_X4Y8_S2BEGb[4] ,
    \Tile_X4Y8_S2BEGb[3] ,
    \Tile_X4Y8_S2BEGb[2] ,
    \Tile_X4Y8_S2BEGb[1] ,
    \Tile_X4Y8_S2BEGb[0] }),
    .S2END({\Tile_X4Y7_S2BEGb[7] ,
    \Tile_X4Y7_S2BEGb[6] ,
    \Tile_X4Y7_S2BEGb[5] ,
    \Tile_X4Y7_S2BEGb[4] ,
    \Tile_X4Y7_S2BEGb[3] ,
    \Tile_X4Y7_S2BEGb[2] ,
    \Tile_X4Y7_S2BEGb[1] ,
    \Tile_X4Y7_S2BEGb[0] }),
    .S2MID({\Tile_X4Y7_S2BEG[7] ,
    \Tile_X4Y7_S2BEG[6] ,
    \Tile_X4Y7_S2BEG[5] ,
    \Tile_X4Y7_S2BEG[4] ,
    \Tile_X4Y7_S2BEG[3] ,
    \Tile_X4Y7_S2BEG[2] ,
    \Tile_X4Y7_S2BEG[1] ,
    \Tile_X4Y7_S2BEG[0] }),
    .S4BEG({\Tile_X4Y8_S4BEG[15] ,
    \Tile_X4Y8_S4BEG[14] ,
    \Tile_X4Y8_S4BEG[13] ,
    \Tile_X4Y8_S4BEG[12] ,
    \Tile_X4Y8_S4BEG[11] ,
    \Tile_X4Y8_S4BEG[10] ,
    \Tile_X4Y8_S4BEG[9] ,
    \Tile_X4Y8_S4BEG[8] ,
    \Tile_X4Y8_S4BEG[7] ,
    \Tile_X4Y8_S4BEG[6] ,
    \Tile_X4Y8_S4BEG[5] ,
    \Tile_X4Y8_S4BEG[4] ,
    \Tile_X4Y8_S4BEG[3] ,
    \Tile_X4Y8_S4BEG[2] ,
    \Tile_X4Y8_S4BEG[1] ,
    \Tile_X4Y8_S4BEG[0] }),
    .S4END({\Tile_X4Y7_S4BEG[15] ,
    \Tile_X4Y7_S4BEG[14] ,
    \Tile_X4Y7_S4BEG[13] ,
    \Tile_X4Y7_S4BEG[12] ,
    \Tile_X4Y7_S4BEG[11] ,
    \Tile_X4Y7_S4BEG[10] ,
    \Tile_X4Y7_S4BEG[9] ,
    \Tile_X4Y7_S4BEG[8] ,
    \Tile_X4Y7_S4BEG[7] ,
    \Tile_X4Y7_S4BEG[6] ,
    \Tile_X4Y7_S4BEG[5] ,
    \Tile_X4Y7_S4BEG[4] ,
    \Tile_X4Y7_S4BEG[3] ,
    \Tile_X4Y7_S4BEG[2] ,
    \Tile_X4Y7_S4BEG[1] ,
    \Tile_X4Y7_S4BEG[0] }),
    .SS4BEG({\Tile_X4Y8_SS4BEG[15] ,
    \Tile_X4Y8_SS4BEG[14] ,
    \Tile_X4Y8_SS4BEG[13] ,
    \Tile_X4Y8_SS4BEG[12] ,
    \Tile_X4Y8_SS4BEG[11] ,
    \Tile_X4Y8_SS4BEG[10] ,
    \Tile_X4Y8_SS4BEG[9] ,
    \Tile_X4Y8_SS4BEG[8] ,
    \Tile_X4Y8_SS4BEG[7] ,
    \Tile_X4Y8_SS4BEG[6] ,
    \Tile_X4Y8_SS4BEG[5] ,
    \Tile_X4Y8_SS4BEG[4] ,
    \Tile_X4Y8_SS4BEG[3] ,
    \Tile_X4Y8_SS4BEG[2] ,
    \Tile_X4Y8_SS4BEG[1] ,
    \Tile_X4Y8_SS4BEG[0] }),
    .SS4END({\Tile_X4Y7_SS4BEG[15] ,
    \Tile_X4Y7_SS4BEG[14] ,
    \Tile_X4Y7_SS4BEG[13] ,
    \Tile_X4Y7_SS4BEG[12] ,
    \Tile_X4Y7_SS4BEG[11] ,
    \Tile_X4Y7_SS4BEG[10] ,
    \Tile_X4Y7_SS4BEG[9] ,
    \Tile_X4Y7_SS4BEG[8] ,
    \Tile_X4Y7_SS4BEG[7] ,
    \Tile_X4Y7_SS4BEG[6] ,
    \Tile_X4Y7_SS4BEG[5] ,
    \Tile_X4Y7_SS4BEG[4] ,
    \Tile_X4Y7_SS4BEG[3] ,
    \Tile_X4Y7_SS4BEG[2] ,
    \Tile_X4Y7_SS4BEG[1] ,
    \Tile_X4Y7_SS4BEG[0] }),
    .W1BEG({\Tile_X4Y8_W1BEG[3] ,
    \Tile_X4Y8_W1BEG[2] ,
    \Tile_X4Y8_W1BEG[1] ,
    \Tile_X4Y8_W1BEG[0] }),
    .W1END({\Tile_X5Y8_W1BEG[3] ,
    \Tile_X5Y8_W1BEG[2] ,
    \Tile_X5Y8_W1BEG[1] ,
    \Tile_X5Y8_W1BEG[0] }),
    .W2BEG({\Tile_X4Y8_W2BEG[7] ,
    \Tile_X4Y8_W2BEG[6] ,
    \Tile_X4Y8_W2BEG[5] ,
    \Tile_X4Y8_W2BEG[4] ,
    \Tile_X4Y8_W2BEG[3] ,
    \Tile_X4Y8_W2BEG[2] ,
    \Tile_X4Y8_W2BEG[1] ,
    \Tile_X4Y8_W2BEG[0] }),
    .W2BEGb({\Tile_X4Y8_W2BEGb[7] ,
    \Tile_X4Y8_W2BEGb[6] ,
    \Tile_X4Y8_W2BEGb[5] ,
    \Tile_X4Y8_W2BEGb[4] ,
    \Tile_X4Y8_W2BEGb[3] ,
    \Tile_X4Y8_W2BEGb[2] ,
    \Tile_X4Y8_W2BEGb[1] ,
    \Tile_X4Y8_W2BEGb[0] }),
    .W2END({\Tile_X5Y8_W2BEGb[7] ,
    \Tile_X5Y8_W2BEGb[6] ,
    \Tile_X5Y8_W2BEGb[5] ,
    \Tile_X5Y8_W2BEGb[4] ,
    \Tile_X5Y8_W2BEGb[3] ,
    \Tile_X5Y8_W2BEGb[2] ,
    \Tile_X5Y8_W2BEGb[1] ,
    \Tile_X5Y8_W2BEGb[0] }),
    .W2MID({\Tile_X5Y8_W2BEG[7] ,
    \Tile_X5Y8_W2BEG[6] ,
    \Tile_X5Y8_W2BEG[5] ,
    \Tile_X5Y8_W2BEG[4] ,
    \Tile_X5Y8_W2BEG[3] ,
    \Tile_X5Y8_W2BEG[2] ,
    \Tile_X5Y8_W2BEG[1] ,
    \Tile_X5Y8_W2BEG[0] }),
    .W6BEG({\Tile_X4Y8_W6BEG[11] ,
    \Tile_X4Y8_W6BEG[10] ,
    \Tile_X4Y8_W6BEG[9] ,
    \Tile_X4Y8_W6BEG[8] ,
    \Tile_X4Y8_W6BEG[7] ,
    \Tile_X4Y8_W6BEG[6] ,
    \Tile_X4Y8_W6BEG[5] ,
    \Tile_X4Y8_W6BEG[4] ,
    \Tile_X4Y8_W6BEG[3] ,
    \Tile_X4Y8_W6BEG[2] ,
    \Tile_X4Y8_W6BEG[1] ,
    \Tile_X4Y8_W6BEG[0] }),
    .W6END({\Tile_X5Y8_W6BEG[11] ,
    \Tile_X5Y8_W6BEG[10] ,
    \Tile_X5Y8_W6BEG[9] ,
    \Tile_X5Y8_W6BEG[8] ,
    \Tile_X5Y8_W6BEG[7] ,
    \Tile_X5Y8_W6BEG[6] ,
    \Tile_X5Y8_W6BEG[5] ,
    \Tile_X5Y8_W6BEG[4] ,
    \Tile_X5Y8_W6BEG[3] ,
    \Tile_X5Y8_W6BEG[2] ,
    \Tile_X5Y8_W6BEG[1] ,
    \Tile_X5Y8_W6BEG[0] }),
    .WW4BEG({\Tile_X4Y8_WW4BEG[15] ,
    \Tile_X4Y8_WW4BEG[14] ,
    \Tile_X4Y8_WW4BEG[13] ,
    \Tile_X4Y8_WW4BEG[12] ,
    \Tile_X4Y8_WW4BEG[11] ,
    \Tile_X4Y8_WW4BEG[10] ,
    \Tile_X4Y8_WW4BEG[9] ,
    \Tile_X4Y8_WW4BEG[8] ,
    \Tile_X4Y8_WW4BEG[7] ,
    \Tile_X4Y8_WW4BEG[6] ,
    \Tile_X4Y8_WW4BEG[5] ,
    \Tile_X4Y8_WW4BEG[4] ,
    \Tile_X4Y8_WW4BEG[3] ,
    \Tile_X4Y8_WW4BEG[2] ,
    \Tile_X4Y8_WW4BEG[1] ,
    \Tile_X4Y8_WW4BEG[0] }),
    .WW4END({\Tile_X5Y8_WW4BEG[15] ,
    \Tile_X5Y8_WW4BEG[14] ,
    \Tile_X5Y8_WW4BEG[13] ,
    \Tile_X5Y8_WW4BEG[12] ,
    \Tile_X5Y8_WW4BEG[11] ,
    \Tile_X5Y8_WW4BEG[10] ,
    \Tile_X5Y8_WW4BEG[9] ,
    \Tile_X5Y8_WW4BEG[8] ,
    \Tile_X5Y8_WW4BEG[7] ,
    \Tile_X5Y8_WW4BEG[6] ,
    \Tile_X5Y8_WW4BEG[5] ,
    \Tile_X5Y8_WW4BEG[4] ,
    \Tile_X5Y8_WW4BEG[3] ,
    \Tile_X5Y8_WW4BEG[2] ,
    \Tile_X5Y8_WW4BEG[1] ,
    \Tile_X5Y8_WW4BEG[0] }));
 RegFile Tile_X4Y9_RegFile (.UserCLK(Tile_X4Y10_UserCLKo),
    .UserCLKo(Tile_X4Y9_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X4Y9_E1BEG[3] ,
    \Tile_X4Y9_E1BEG[2] ,
    \Tile_X4Y9_E1BEG[1] ,
    \Tile_X4Y9_E1BEG[0] }),
    .E1END({\Tile_X3Y9_E1BEG[3] ,
    \Tile_X3Y9_E1BEG[2] ,
    \Tile_X3Y9_E1BEG[1] ,
    \Tile_X3Y9_E1BEG[0] }),
    .E2BEG({\Tile_X4Y9_E2BEG[7] ,
    \Tile_X4Y9_E2BEG[6] ,
    \Tile_X4Y9_E2BEG[5] ,
    \Tile_X4Y9_E2BEG[4] ,
    \Tile_X4Y9_E2BEG[3] ,
    \Tile_X4Y9_E2BEG[2] ,
    \Tile_X4Y9_E2BEG[1] ,
    \Tile_X4Y9_E2BEG[0] }),
    .E2BEGb({\Tile_X4Y9_E2BEGb[7] ,
    \Tile_X4Y9_E2BEGb[6] ,
    \Tile_X4Y9_E2BEGb[5] ,
    \Tile_X4Y9_E2BEGb[4] ,
    \Tile_X4Y9_E2BEGb[3] ,
    \Tile_X4Y9_E2BEGb[2] ,
    \Tile_X4Y9_E2BEGb[1] ,
    \Tile_X4Y9_E2BEGb[0] }),
    .E2END({\Tile_X3Y9_E2BEGb[7] ,
    \Tile_X3Y9_E2BEGb[6] ,
    \Tile_X3Y9_E2BEGb[5] ,
    \Tile_X3Y9_E2BEGb[4] ,
    \Tile_X3Y9_E2BEGb[3] ,
    \Tile_X3Y9_E2BEGb[2] ,
    \Tile_X3Y9_E2BEGb[1] ,
    \Tile_X3Y9_E2BEGb[0] }),
    .E2MID({\Tile_X3Y9_E2BEG[7] ,
    \Tile_X3Y9_E2BEG[6] ,
    \Tile_X3Y9_E2BEG[5] ,
    \Tile_X3Y9_E2BEG[4] ,
    \Tile_X3Y9_E2BEG[3] ,
    \Tile_X3Y9_E2BEG[2] ,
    \Tile_X3Y9_E2BEG[1] ,
    \Tile_X3Y9_E2BEG[0] }),
    .E6BEG({\Tile_X4Y9_E6BEG[11] ,
    \Tile_X4Y9_E6BEG[10] ,
    \Tile_X4Y9_E6BEG[9] ,
    \Tile_X4Y9_E6BEG[8] ,
    \Tile_X4Y9_E6BEG[7] ,
    \Tile_X4Y9_E6BEG[6] ,
    \Tile_X4Y9_E6BEG[5] ,
    \Tile_X4Y9_E6BEG[4] ,
    \Tile_X4Y9_E6BEG[3] ,
    \Tile_X4Y9_E6BEG[2] ,
    \Tile_X4Y9_E6BEG[1] ,
    \Tile_X4Y9_E6BEG[0] }),
    .E6END({\Tile_X3Y9_E6BEG[11] ,
    \Tile_X3Y9_E6BEG[10] ,
    \Tile_X3Y9_E6BEG[9] ,
    \Tile_X3Y9_E6BEG[8] ,
    \Tile_X3Y9_E6BEG[7] ,
    \Tile_X3Y9_E6BEG[6] ,
    \Tile_X3Y9_E6BEG[5] ,
    \Tile_X3Y9_E6BEG[4] ,
    \Tile_X3Y9_E6BEG[3] ,
    \Tile_X3Y9_E6BEG[2] ,
    \Tile_X3Y9_E6BEG[1] ,
    \Tile_X3Y9_E6BEG[0] }),
    .EE4BEG({\Tile_X4Y9_EE4BEG[15] ,
    \Tile_X4Y9_EE4BEG[14] ,
    \Tile_X4Y9_EE4BEG[13] ,
    \Tile_X4Y9_EE4BEG[12] ,
    \Tile_X4Y9_EE4BEG[11] ,
    \Tile_X4Y9_EE4BEG[10] ,
    \Tile_X4Y9_EE4BEG[9] ,
    \Tile_X4Y9_EE4BEG[8] ,
    \Tile_X4Y9_EE4BEG[7] ,
    \Tile_X4Y9_EE4BEG[6] ,
    \Tile_X4Y9_EE4BEG[5] ,
    \Tile_X4Y9_EE4BEG[4] ,
    \Tile_X4Y9_EE4BEG[3] ,
    \Tile_X4Y9_EE4BEG[2] ,
    \Tile_X4Y9_EE4BEG[1] ,
    \Tile_X4Y9_EE4BEG[0] }),
    .EE4END({\Tile_X3Y9_EE4BEG[15] ,
    \Tile_X3Y9_EE4BEG[14] ,
    \Tile_X3Y9_EE4BEG[13] ,
    \Tile_X3Y9_EE4BEG[12] ,
    \Tile_X3Y9_EE4BEG[11] ,
    \Tile_X3Y9_EE4BEG[10] ,
    \Tile_X3Y9_EE4BEG[9] ,
    \Tile_X3Y9_EE4BEG[8] ,
    \Tile_X3Y9_EE4BEG[7] ,
    \Tile_X3Y9_EE4BEG[6] ,
    \Tile_X3Y9_EE4BEG[5] ,
    \Tile_X3Y9_EE4BEG[4] ,
    \Tile_X3Y9_EE4BEG[3] ,
    \Tile_X3Y9_EE4BEG[2] ,
    \Tile_X3Y9_EE4BEG[1] ,
    \Tile_X3Y9_EE4BEG[0] }),
    .FrameData({\Tile_X3Y9_FrameData_O[31] ,
    \Tile_X3Y9_FrameData_O[30] ,
    \Tile_X3Y9_FrameData_O[29] ,
    \Tile_X3Y9_FrameData_O[28] ,
    \Tile_X3Y9_FrameData_O[27] ,
    \Tile_X3Y9_FrameData_O[26] ,
    \Tile_X3Y9_FrameData_O[25] ,
    \Tile_X3Y9_FrameData_O[24] ,
    \Tile_X3Y9_FrameData_O[23] ,
    \Tile_X3Y9_FrameData_O[22] ,
    \Tile_X3Y9_FrameData_O[21] ,
    \Tile_X3Y9_FrameData_O[20] ,
    \Tile_X3Y9_FrameData_O[19] ,
    \Tile_X3Y9_FrameData_O[18] ,
    \Tile_X3Y9_FrameData_O[17] ,
    \Tile_X3Y9_FrameData_O[16] ,
    \Tile_X3Y9_FrameData_O[15] ,
    \Tile_X3Y9_FrameData_O[14] ,
    \Tile_X3Y9_FrameData_O[13] ,
    \Tile_X3Y9_FrameData_O[12] ,
    \Tile_X3Y9_FrameData_O[11] ,
    \Tile_X3Y9_FrameData_O[10] ,
    \Tile_X3Y9_FrameData_O[9] ,
    \Tile_X3Y9_FrameData_O[8] ,
    \Tile_X3Y9_FrameData_O[7] ,
    \Tile_X3Y9_FrameData_O[6] ,
    \Tile_X3Y9_FrameData_O[5] ,
    \Tile_X3Y9_FrameData_O[4] ,
    \Tile_X3Y9_FrameData_O[3] ,
    \Tile_X3Y9_FrameData_O[2] ,
    \Tile_X3Y9_FrameData_O[1] ,
    \Tile_X3Y9_FrameData_O[0] }),
    .FrameData_O({\Tile_X4Y9_FrameData_O[31] ,
    \Tile_X4Y9_FrameData_O[30] ,
    \Tile_X4Y9_FrameData_O[29] ,
    \Tile_X4Y9_FrameData_O[28] ,
    \Tile_X4Y9_FrameData_O[27] ,
    \Tile_X4Y9_FrameData_O[26] ,
    \Tile_X4Y9_FrameData_O[25] ,
    \Tile_X4Y9_FrameData_O[24] ,
    \Tile_X4Y9_FrameData_O[23] ,
    \Tile_X4Y9_FrameData_O[22] ,
    \Tile_X4Y9_FrameData_O[21] ,
    \Tile_X4Y9_FrameData_O[20] ,
    \Tile_X4Y9_FrameData_O[19] ,
    \Tile_X4Y9_FrameData_O[18] ,
    \Tile_X4Y9_FrameData_O[17] ,
    \Tile_X4Y9_FrameData_O[16] ,
    \Tile_X4Y9_FrameData_O[15] ,
    \Tile_X4Y9_FrameData_O[14] ,
    \Tile_X4Y9_FrameData_O[13] ,
    \Tile_X4Y9_FrameData_O[12] ,
    \Tile_X4Y9_FrameData_O[11] ,
    \Tile_X4Y9_FrameData_O[10] ,
    \Tile_X4Y9_FrameData_O[9] ,
    \Tile_X4Y9_FrameData_O[8] ,
    \Tile_X4Y9_FrameData_O[7] ,
    \Tile_X4Y9_FrameData_O[6] ,
    \Tile_X4Y9_FrameData_O[5] ,
    \Tile_X4Y9_FrameData_O[4] ,
    \Tile_X4Y9_FrameData_O[3] ,
    \Tile_X4Y9_FrameData_O[2] ,
    \Tile_X4Y9_FrameData_O[1] ,
    \Tile_X4Y9_FrameData_O[0] }),
    .FrameStrobe({\Tile_X4Y10_FrameStrobe_O[19] ,
    \Tile_X4Y10_FrameStrobe_O[18] ,
    \Tile_X4Y10_FrameStrobe_O[17] ,
    \Tile_X4Y10_FrameStrobe_O[16] ,
    \Tile_X4Y10_FrameStrobe_O[15] ,
    \Tile_X4Y10_FrameStrobe_O[14] ,
    \Tile_X4Y10_FrameStrobe_O[13] ,
    \Tile_X4Y10_FrameStrobe_O[12] ,
    \Tile_X4Y10_FrameStrobe_O[11] ,
    \Tile_X4Y10_FrameStrobe_O[10] ,
    \Tile_X4Y10_FrameStrobe_O[9] ,
    \Tile_X4Y10_FrameStrobe_O[8] ,
    \Tile_X4Y10_FrameStrobe_O[7] ,
    \Tile_X4Y10_FrameStrobe_O[6] ,
    \Tile_X4Y10_FrameStrobe_O[5] ,
    \Tile_X4Y10_FrameStrobe_O[4] ,
    \Tile_X4Y10_FrameStrobe_O[3] ,
    \Tile_X4Y10_FrameStrobe_O[2] ,
    \Tile_X4Y10_FrameStrobe_O[1] ,
    \Tile_X4Y10_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X4Y9_FrameStrobe_O[19] ,
    \Tile_X4Y9_FrameStrobe_O[18] ,
    \Tile_X4Y9_FrameStrobe_O[17] ,
    \Tile_X4Y9_FrameStrobe_O[16] ,
    \Tile_X4Y9_FrameStrobe_O[15] ,
    \Tile_X4Y9_FrameStrobe_O[14] ,
    \Tile_X4Y9_FrameStrobe_O[13] ,
    \Tile_X4Y9_FrameStrobe_O[12] ,
    \Tile_X4Y9_FrameStrobe_O[11] ,
    \Tile_X4Y9_FrameStrobe_O[10] ,
    \Tile_X4Y9_FrameStrobe_O[9] ,
    \Tile_X4Y9_FrameStrobe_O[8] ,
    \Tile_X4Y9_FrameStrobe_O[7] ,
    \Tile_X4Y9_FrameStrobe_O[6] ,
    \Tile_X4Y9_FrameStrobe_O[5] ,
    \Tile_X4Y9_FrameStrobe_O[4] ,
    \Tile_X4Y9_FrameStrobe_O[3] ,
    \Tile_X4Y9_FrameStrobe_O[2] ,
    \Tile_X4Y9_FrameStrobe_O[1] ,
    \Tile_X4Y9_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X4Y9_N1BEG[3] ,
    \Tile_X4Y9_N1BEG[2] ,
    \Tile_X4Y9_N1BEG[1] ,
    \Tile_X4Y9_N1BEG[0] }),
    .N1END({\Tile_X4Y10_N1BEG[3] ,
    \Tile_X4Y10_N1BEG[2] ,
    \Tile_X4Y10_N1BEG[1] ,
    \Tile_X4Y10_N1BEG[0] }),
    .N2BEG({\Tile_X4Y9_N2BEG[7] ,
    \Tile_X4Y9_N2BEG[6] ,
    \Tile_X4Y9_N2BEG[5] ,
    \Tile_X4Y9_N2BEG[4] ,
    \Tile_X4Y9_N2BEG[3] ,
    \Tile_X4Y9_N2BEG[2] ,
    \Tile_X4Y9_N2BEG[1] ,
    \Tile_X4Y9_N2BEG[0] }),
    .N2BEGb({\Tile_X4Y9_N2BEGb[7] ,
    \Tile_X4Y9_N2BEGb[6] ,
    \Tile_X4Y9_N2BEGb[5] ,
    \Tile_X4Y9_N2BEGb[4] ,
    \Tile_X4Y9_N2BEGb[3] ,
    \Tile_X4Y9_N2BEGb[2] ,
    \Tile_X4Y9_N2BEGb[1] ,
    \Tile_X4Y9_N2BEGb[0] }),
    .N2END({\Tile_X4Y10_N2BEGb[7] ,
    \Tile_X4Y10_N2BEGb[6] ,
    \Tile_X4Y10_N2BEGb[5] ,
    \Tile_X4Y10_N2BEGb[4] ,
    \Tile_X4Y10_N2BEGb[3] ,
    \Tile_X4Y10_N2BEGb[2] ,
    \Tile_X4Y10_N2BEGb[1] ,
    \Tile_X4Y10_N2BEGb[0] }),
    .N2MID({\Tile_X4Y10_N2BEG[7] ,
    \Tile_X4Y10_N2BEG[6] ,
    \Tile_X4Y10_N2BEG[5] ,
    \Tile_X4Y10_N2BEG[4] ,
    \Tile_X4Y10_N2BEG[3] ,
    \Tile_X4Y10_N2BEG[2] ,
    \Tile_X4Y10_N2BEG[1] ,
    \Tile_X4Y10_N2BEG[0] }),
    .N4BEG({\Tile_X4Y9_N4BEG[15] ,
    \Tile_X4Y9_N4BEG[14] ,
    \Tile_X4Y9_N4BEG[13] ,
    \Tile_X4Y9_N4BEG[12] ,
    \Tile_X4Y9_N4BEG[11] ,
    \Tile_X4Y9_N4BEG[10] ,
    \Tile_X4Y9_N4BEG[9] ,
    \Tile_X4Y9_N4BEG[8] ,
    \Tile_X4Y9_N4BEG[7] ,
    \Tile_X4Y9_N4BEG[6] ,
    \Tile_X4Y9_N4BEG[5] ,
    \Tile_X4Y9_N4BEG[4] ,
    \Tile_X4Y9_N4BEG[3] ,
    \Tile_X4Y9_N4BEG[2] ,
    \Tile_X4Y9_N4BEG[1] ,
    \Tile_X4Y9_N4BEG[0] }),
    .N4END({\Tile_X4Y10_N4BEG[15] ,
    \Tile_X4Y10_N4BEG[14] ,
    \Tile_X4Y10_N4BEG[13] ,
    \Tile_X4Y10_N4BEG[12] ,
    \Tile_X4Y10_N4BEG[11] ,
    \Tile_X4Y10_N4BEG[10] ,
    \Tile_X4Y10_N4BEG[9] ,
    \Tile_X4Y10_N4BEG[8] ,
    \Tile_X4Y10_N4BEG[7] ,
    \Tile_X4Y10_N4BEG[6] ,
    \Tile_X4Y10_N4BEG[5] ,
    \Tile_X4Y10_N4BEG[4] ,
    \Tile_X4Y10_N4BEG[3] ,
    \Tile_X4Y10_N4BEG[2] ,
    \Tile_X4Y10_N4BEG[1] ,
    \Tile_X4Y10_N4BEG[0] }),
    .NN4BEG({\Tile_X4Y9_NN4BEG[15] ,
    \Tile_X4Y9_NN4BEG[14] ,
    \Tile_X4Y9_NN4BEG[13] ,
    \Tile_X4Y9_NN4BEG[12] ,
    \Tile_X4Y9_NN4BEG[11] ,
    \Tile_X4Y9_NN4BEG[10] ,
    \Tile_X4Y9_NN4BEG[9] ,
    \Tile_X4Y9_NN4BEG[8] ,
    \Tile_X4Y9_NN4BEG[7] ,
    \Tile_X4Y9_NN4BEG[6] ,
    \Tile_X4Y9_NN4BEG[5] ,
    \Tile_X4Y9_NN4BEG[4] ,
    \Tile_X4Y9_NN4BEG[3] ,
    \Tile_X4Y9_NN4BEG[2] ,
    \Tile_X4Y9_NN4BEG[1] ,
    \Tile_X4Y9_NN4BEG[0] }),
    .NN4END({\Tile_X4Y10_NN4BEG[15] ,
    \Tile_X4Y10_NN4BEG[14] ,
    \Tile_X4Y10_NN4BEG[13] ,
    \Tile_X4Y10_NN4BEG[12] ,
    \Tile_X4Y10_NN4BEG[11] ,
    \Tile_X4Y10_NN4BEG[10] ,
    \Tile_X4Y10_NN4BEG[9] ,
    \Tile_X4Y10_NN4BEG[8] ,
    \Tile_X4Y10_NN4BEG[7] ,
    \Tile_X4Y10_NN4BEG[6] ,
    \Tile_X4Y10_NN4BEG[5] ,
    \Tile_X4Y10_NN4BEG[4] ,
    \Tile_X4Y10_NN4BEG[3] ,
    \Tile_X4Y10_NN4BEG[2] ,
    \Tile_X4Y10_NN4BEG[1] ,
    \Tile_X4Y10_NN4BEG[0] }),
    .S1BEG({\Tile_X4Y9_S1BEG[3] ,
    \Tile_X4Y9_S1BEG[2] ,
    \Tile_X4Y9_S1BEG[1] ,
    \Tile_X4Y9_S1BEG[0] }),
    .S1END({\Tile_X4Y8_S1BEG[3] ,
    \Tile_X4Y8_S1BEG[2] ,
    \Tile_X4Y8_S1BEG[1] ,
    \Tile_X4Y8_S1BEG[0] }),
    .S2BEG({\Tile_X4Y9_S2BEG[7] ,
    \Tile_X4Y9_S2BEG[6] ,
    \Tile_X4Y9_S2BEG[5] ,
    \Tile_X4Y9_S2BEG[4] ,
    \Tile_X4Y9_S2BEG[3] ,
    \Tile_X4Y9_S2BEG[2] ,
    \Tile_X4Y9_S2BEG[1] ,
    \Tile_X4Y9_S2BEG[0] }),
    .S2BEGb({\Tile_X4Y9_S2BEGb[7] ,
    \Tile_X4Y9_S2BEGb[6] ,
    \Tile_X4Y9_S2BEGb[5] ,
    \Tile_X4Y9_S2BEGb[4] ,
    \Tile_X4Y9_S2BEGb[3] ,
    \Tile_X4Y9_S2BEGb[2] ,
    \Tile_X4Y9_S2BEGb[1] ,
    \Tile_X4Y9_S2BEGb[0] }),
    .S2END({\Tile_X4Y8_S2BEGb[7] ,
    \Tile_X4Y8_S2BEGb[6] ,
    \Tile_X4Y8_S2BEGb[5] ,
    \Tile_X4Y8_S2BEGb[4] ,
    \Tile_X4Y8_S2BEGb[3] ,
    \Tile_X4Y8_S2BEGb[2] ,
    \Tile_X4Y8_S2BEGb[1] ,
    \Tile_X4Y8_S2BEGb[0] }),
    .S2MID({\Tile_X4Y8_S2BEG[7] ,
    \Tile_X4Y8_S2BEG[6] ,
    \Tile_X4Y8_S2BEG[5] ,
    \Tile_X4Y8_S2BEG[4] ,
    \Tile_X4Y8_S2BEG[3] ,
    \Tile_X4Y8_S2BEG[2] ,
    \Tile_X4Y8_S2BEG[1] ,
    \Tile_X4Y8_S2BEG[0] }),
    .S4BEG({\Tile_X4Y9_S4BEG[15] ,
    \Tile_X4Y9_S4BEG[14] ,
    \Tile_X4Y9_S4BEG[13] ,
    \Tile_X4Y9_S4BEG[12] ,
    \Tile_X4Y9_S4BEG[11] ,
    \Tile_X4Y9_S4BEG[10] ,
    \Tile_X4Y9_S4BEG[9] ,
    \Tile_X4Y9_S4BEG[8] ,
    \Tile_X4Y9_S4BEG[7] ,
    \Tile_X4Y9_S4BEG[6] ,
    \Tile_X4Y9_S4BEG[5] ,
    \Tile_X4Y9_S4BEG[4] ,
    \Tile_X4Y9_S4BEG[3] ,
    \Tile_X4Y9_S4BEG[2] ,
    \Tile_X4Y9_S4BEG[1] ,
    \Tile_X4Y9_S4BEG[0] }),
    .S4END({\Tile_X4Y8_S4BEG[15] ,
    \Tile_X4Y8_S4BEG[14] ,
    \Tile_X4Y8_S4BEG[13] ,
    \Tile_X4Y8_S4BEG[12] ,
    \Tile_X4Y8_S4BEG[11] ,
    \Tile_X4Y8_S4BEG[10] ,
    \Tile_X4Y8_S4BEG[9] ,
    \Tile_X4Y8_S4BEG[8] ,
    \Tile_X4Y8_S4BEG[7] ,
    \Tile_X4Y8_S4BEG[6] ,
    \Tile_X4Y8_S4BEG[5] ,
    \Tile_X4Y8_S4BEG[4] ,
    \Tile_X4Y8_S4BEG[3] ,
    \Tile_X4Y8_S4BEG[2] ,
    \Tile_X4Y8_S4BEG[1] ,
    \Tile_X4Y8_S4BEG[0] }),
    .SS4BEG({\Tile_X4Y9_SS4BEG[15] ,
    \Tile_X4Y9_SS4BEG[14] ,
    \Tile_X4Y9_SS4BEG[13] ,
    \Tile_X4Y9_SS4BEG[12] ,
    \Tile_X4Y9_SS4BEG[11] ,
    \Tile_X4Y9_SS4BEG[10] ,
    \Tile_X4Y9_SS4BEG[9] ,
    \Tile_X4Y9_SS4BEG[8] ,
    \Tile_X4Y9_SS4BEG[7] ,
    \Tile_X4Y9_SS4BEG[6] ,
    \Tile_X4Y9_SS4BEG[5] ,
    \Tile_X4Y9_SS4BEG[4] ,
    \Tile_X4Y9_SS4BEG[3] ,
    \Tile_X4Y9_SS4BEG[2] ,
    \Tile_X4Y9_SS4BEG[1] ,
    \Tile_X4Y9_SS4BEG[0] }),
    .SS4END({\Tile_X4Y8_SS4BEG[15] ,
    \Tile_X4Y8_SS4BEG[14] ,
    \Tile_X4Y8_SS4BEG[13] ,
    \Tile_X4Y8_SS4BEG[12] ,
    \Tile_X4Y8_SS4BEG[11] ,
    \Tile_X4Y8_SS4BEG[10] ,
    \Tile_X4Y8_SS4BEG[9] ,
    \Tile_X4Y8_SS4BEG[8] ,
    \Tile_X4Y8_SS4BEG[7] ,
    \Tile_X4Y8_SS4BEG[6] ,
    \Tile_X4Y8_SS4BEG[5] ,
    \Tile_X4Y8_SS4BEG[4] ,
    \Tile_X4Y8_SS4BEG[3] ,
    \Tile_X4Y8_SS4BEG[2] ,
    \Tile_X4Y8_SS4BEG[1] ,
    \Tile_X4Y8_SS4BEG[0] }),
    .W1BEG({\Tile_X4Y9_W1BEG[3] ,
    \Tile_X4Y9_W1BEG[2] ,
    \Tile_X4Y9_W1BEG[1] ,
    \Tile_X4Y9_W1BEG[0] }),
    .W1END({\Tile_X5Y9_W1BEG[3] ,
    \Tile_X5Y9_W1BEG[2] ,
    \Tile_X5Y9_W1BEG[1] ,
    \Tile_X5Y9_W1BEG[0] }),
    .W2BEG({\Tile_X4Y9_W2BEG[7] ,
    \Tile_X4Y9_W2BEG[6] ,
    \Tile_X4Y9_W2BEG[5] ,
    \Tile_X4Y9_W2BEG[4] ,
    \Tile_X4Y9_W2BEG[3] ,
    \Tile_X4Y9_W2BEG[2] ,
    \Tile_X4Y9_W2BEG[1] ,
    \Tile_X4Y9_W2BEG[0] }),
    .W2BEGb({\Tile_X4Y9_W2BEGb[7] ,
    \Tile_X4Y9_W2BEGb[6] ,
    \Tile_X4Y9_W2BEGb[5] ,
    \Tile_X4Y9_W2BEGb[4] ,
    \Tile_X4Y9_W2BEGb[3] ,
    \Tile_X4Y9_W2BEGb[2] ,
    \Tile_X4Y9_W2BEGb[1] ,
    \Tile_X4Y9_W2BEGb[0] }),
    .W2END({\Tile_X5Y9_W2BEGb[7] ,
    \Tile_X5Y9_W2BEGb[6] ,
    \Tile_X5Y9_W2BEGb[5] ,
    \Tile_X5Y9_W2BEGb[4] ,
    \Tile_X5Y9_W2BEGb[3] ,
    \Tile_X5Y9_W2BEGb[2] ,
    \Tile_X5Y9_W2BEGb[1] ,
    \Tile_X5Y9_W2BEGb[0] }),
    .W2MID({\Tile_X5Y9_W2BEG[7] ,
    \Tile_X5Y9_W2BEG[6] ,
    \Tile_X5Y9_W2BEG[5] ,
    \Tile_X5Y9_W2BEG[4] ,
    \Tile_X5Y9_W2BEG[3] ,
    \Tile_X5Y9_W2BEG[2] ,
    \Tile_X5Y9_W2BEG[1] ,
    \Tile_X5Y9_W2BEG[0] }),
    .W6BEG({\Tile_X4Y9_W6BEG[11] ,
    \Tile_X4Y9_W6BEG[10] ,
    \Tile_X4Y9_W6BEG[9] ,
    \Tile_X4Y9_W6BEG[8] ,
    \Tile_X4Y9_W6BEG[7] ,
    \Tile_X4Y9_W6BEG[6] ,
    \Tile_X4Y9_W6BEG[5] ,
    \Tile_X4Y9_W6BEG[4] ,
    \Tile_X4Y9_W6BEG[3] ,
    \Tile_X4Y9_W6BEG[2] ,
    \Tile_X4Y9_W6BEG[1] ,
    \Tile_X4Y9_W6BEG[0] }),
    .W6END({\Tile_X5Y9_W6BEG[11] ,
    \Tile_X5Y9_W6BEG[10] ,
    \Tile_X5Y9_W6BEG[9] ,
    \Tile_X5Y9_W6BEG[8] ,
    \Tile_X5Y9_W6BEG[7] ,
    \Tile_X5Y9_W6BEG[6] ,
    \Tile_X5Y9_W6BEG[5] ,
    \Tile_X5Y9_W6BEG[4] ,
    \Tile_X5Y9_W6BEG[3] ,
    \Tile_X5Y9_W6BEG[2] ,
    \Tile_X5Y9_W6BEG[1] ,
    \Tile_X5Y9_W6BEG[0] }),
    .WW4BEG({\Tile_X4Y9_WW4BEG[15] ,
    \Tile_X4Y9_WW4BEG[14] ,
    \Tile_X4Y9_WW4BEG[13] ,
    \Tile_X4Y9_WW4BEG[12] ,
    \Tile_X4Y9_WW4BEG[11] ,
    \Tile_X4Y9_WW4BEG[10] ,
    \Tile_X4Y9_WW4BEG[9] ,
    \Tile_X4Y9_WW4BEG[8] ,
    \Tile_X4Y9_WW4BEG[7] ,
    \Tile_X4Y9_WW4BEG[6] ,
    \Tile_X4Y9_WW4BEG[5] ,
    \Tile_X4Y9_WW4BEG[4] ,
    \Tile_X4Y9_WW4BEG[3] ,
    \Tile_X4Y9_WW4BEG[2] ,
    \Tile_X4Y9_WW4BEG[1] ,
    \Tile_X4Y9_WW4BEG[0] }),
    .WW4END({\Tile_X5Y9_WW4BEG[15] ,
    \Tile_X5Y9_WW4BEG[14] ,
    \Tile_X5Y9_WW4BEG[13] ,
    \Tile_X5Y9_WW4BEG[12] ,
    \Tile_X5Y9_WW4BEG[11] ,
    \Tile_X5Y9_WW4BEG[10] ,
    \Tile_X5Y9_WW4BEG[9] ,
    \Tile_X5Y9_WW4BEG[8] ,
    \Tile_X5Y9_WW4BEG[7] ,
    \Tile_X5Y9_WW4BEG[6] ,
    \Tile_X5Y9_WW4BEG[5] ,
    \Tile_X5Y9_WW4BEG[4] ,
    \Tile_X5Y9_WW4BEG[3] ,
    \Tile_X5Y9_WW4BEG[2] ,
    \Tile_X5Y9_WW4BEG[1] ,
    \Tile_X5Y9_WW4BEG[0] }));
 N_term_single Tile_X5Y0_N_term_single (.Ci(Tile_X5Y1_Co),
    .UserCLK(Tile_X5Y1_UserCLKo),
    .UserCLKo(Tile_X5Y0_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .FrameData({\Tile_X4Y0_FrameData_O[31] ,
    \Tile_X4Y0_FrameData_O[30] ,
    \Tile_X4Y0_FrameData_O[29] ,
    \Tile_X4Y0_FrameData_O[28] ,
    \Tile_X4Y0_FrameData_O[27] ,
    \Tile_X4Y0_FrameData_O[26] ,
    \Tile_X4Y0_FrameData_O[25] ,
    \Tile_X4Y0_FrameData_O[24] ,
    \Tile_X4Y0_FrameData_O[23] ,
    \Tile_X4Y0_FrameData_O[22] ,
    \Tile_X4Y0_FrameData_O[21] ,
    \Tile_X4Y0_FrameData_O[20] ,
    \Tile_X4Y0_FrameData_O[19] ,
    \Tile_X4Y0_FrameData_O[18] ,
    \Tile_X4Y0_FrameData_O[17] ,
    \Tile_X4Y0_FrameData_O[16] ,
    \Tile_X4Y0_FrameData_O[15] ,
    \Tile_X4Y0_FrameData_O[14] ,
    \Tile_X4Y0_FrameData_O[13] ,
    \Tile_X4Y0_FrameData_O[12] ,
    \Tile_X4Y0_FrameData_O[11] ,
    \Tile_X4Y0_FrameData_O[10] ,
    \Tile_X4Y0_FrameData_O[9] ,
    \Tile_X4Y0_FrameData_O[8] ,
    \Tile_X4Y0_FrameData_O[7] ,
    \Tile_X4Y0_FrameData_O[6] ,
    \Tile_X4Y0_FrameData_O[5] ,
    \Tile_X4Y0_FrameData_O[4] ,
    \Tile_X4Y0_FrameData_O[3] ,
    \Tile_X4Y0_FrameData_O[2] ,
    \Tile_X4Y0_FrameData_O[1] ,
    \Tile_X4Y0_FrameData_O[0] }),
    .FrameData_O({\Tile_X5Y0_FrameData_O[31] ,
    \Tile_X5Y0_FrameData_O[30] ,
    \Tile_X5Y0_FrameData_O[29] ,
    \Tile_X5Y0_FrameData_O[28] ,
    \Tile_X5Y0_FrameData_O[27] ,
    \Tile_X5Y0_FrameData_O[26] ,
    \Tile_X5Y0_FrameData_O[25] ,
    \Tile_X5Y0_FrameData_O[24] ,
    \Tile_X5Y0_FrameData_O[23] ,
    \Tile_X5Y0_FrameData_O[22] ,
    \Tile_X5Y0_FrameData_O[21] ,
    \Tile_X5Y0_FrameData_O[20] ,
    \Tile_X5Y0_FrameData_O[19] ,
    \Tile_X5Y0_FrameData_O[18] ,
    \Tile_X5Y0_FrameData_O[17] ,
    \Tile_X5Y0_FrameData_O[16] ,
    \Tile_X5Y0_FrameData_O[15] ,
    \Tile_X5Y0_FrameData_O[14] ,
    \Tile_X5Y0_FrameData_O[13] ,
    \Tile_X5Y0_FrameData_O[12] ,
    \Tile_X5Y0_FrameData_O[11] ,
    \Tile_X5Y0_FrameData_O[10] ,
    \Tile_X5Y0_FrameData_O[9] ,
    \Tile_X5Y0_FrameData_O[8] ,
    \Tile_X5Y0_FrameData_O[7] ,
    \Tile_X5Y0_FrameData_O[6] ,
    \Tile_X5Y0_FrameData_O[5] ,
    \Tile_X5Y0_FrameData_O[4] ,
    \Tile_X5Y0_FrameData_O[3] ,
    \Tile_X5Y0_FrameData_O[2] ,
    \Tile_X5Y0_FrameData_O[1] ,
    \Tile_X5Y0_FrameData_O[0] }),
    .FrameStrobe({\Tile_X5Y1_FrameStrobe_O[19] ,
    \Tile_X5Y1_FrameStrobe_O[18] ,
    \Tile_X5Y1_FrameStrobe_O[17] ,
    \Tile_X5Y1_FrameStrobe_O[16] ,
    \Tile_X5Y1_FrameStrobe_O[15] ,
    \Tile_X5Y1_FrameStrobe_O[14] ,
    \Tile_X5Y1_FrameStrobe_O[13] ,
    \Tile_X5Y1_FrameStrobe_O[12] ,
    \Tile_X5Y1_FrameStrobe_O[11] ,
    \Tile_X5Y1_FrameStrobe_O[10] ,
    \Tile_X5Y1_FrameStrobe_O[9] ,
    \Tile_X5Y1_FrameStrobe_O[8] ,
    \Tile_X5Y1_FrameStrobe_O[7] ,
    \Tile_X5Y1_FrameStrobe_O[6] ,
    \Tile_X5Y1_FrameStrobe_O[5] ,
    \Tile_X5Y1_FrameStrobe_O[4] ,
    \Tile_X5Y1_FrameStrobe_O[3] ,
    \Tile_X5Y1_FrameStrobe_O[2] ,
    \Tile_X5Y1_FrameStrobe_O[1] ,
    \Tile_X5Y1_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X5Y0_FrameStrobe_O[19] ,
    \Tile_X5Y0_FrameStrobe_O[18] ,
    \Tile_X5Y0_FrameStrobe_O[17] ,
    \Tile_X5Y0_FrameStrobe_O[16] ,
    \Tile_X5Y0_FrameStrobe_O[15] ,
    \Tile_X5Y0_FrameStrobe_O[14] ,
    \Tile_X5Y0_FrameStrobe_O[13] ,
    \Tile_X5Y0_FrameStrobe_O[12] ,
    \Tile_X5Y0_FrameStrobe_O[11] ,
    \Tile_X5Y0_FrameStrobe_O[10] ,
    \Tile_X5Y0_FrameStrobe_O[9] ,
    \Tile_X5Y0_FrameStrobe_O[8] ,
    \Tile_X5Y0_FrameStrobe_O[7] ,
    \Tile_X5Y0_FrameStrobe_O[6] ,
    \Tile_X5Y0_FrameStrobe_O[5] ,
    \Tile_X5Y0_FrameStrobe_O[4] ,
    \Tile_X5Y0_FrameStrobe_O[3] ,
    \Tile_X5Y0_FrameStrobe_O[2] ,
    \Tile_X5Y0_FrameStrobe_O[1] ,
    \Tile_X5Y0_FrameStrobe_O[0] }),
    .N1END({\Tile_X5Y1_N1BEG[3] ,
    \Tile_X5Y1_N1BEG[2] ,
    \Tile_X5Y1_N1BEG[1] ,
    \Tile_X5Y1_N1BEG[0] }),
    .N2END({\Tile_X5Y1_N2BEGb[7] ,
    \Tile_X5Y1_N2BEGb[6] ,
    \Tile_X5Y1_N2BEGb[5] ,
    \Tile_X5Y1_N2BEGb[4] ,
    \Tile_X5Y1_N2BEGb[3] ,
    \Tile_X5Y1_N2BEGb[2] ,
    \Tile_X5Y1_N2BEGb[1] ,
    \Tile_X5Y1_N2BEGb[0] }),
    .N2MID({\Tile_X5Y1_N2BEG[7] ,
    \Tile_X5Y1_N2BEG[6] ,
    \Tile_X5Y1_N2BEG[5] ,
    \Tile_X5Y1_N2BEG[4] ,
    \Tile_X5Y1_N2BEG[3] ,
    \Tile_X5Y1_N2BEG[2] ,
    \Tile_X5Y1_N2BEG[1] ,
    \Tile_X5Y1_N2BEG[0] }),
    .N4END({\Tile_X5Y1_N4BEG[15] ,
    \Tile_X5Y1_N4BEG[14] ,
    \Tile_X5Y1_N4BEG[13] ,
    \Tile_X5Y1_N4BEG[12] ,
    \Tile_X5Y1_N4BEG[11] ,
    \Tile_X5Y1_N4BEG[10] ,
    \Tile_X5Y1_N4BEG[9] ,
    \Tile_X5Y1_N4BEG[8] ,
    \Tile_X5Y1_N4BEG[7] ,
    \Tile_X5Y1_N4BEG[6] ,
    \Tile_X5Y1_N4BEG[5] ,
    \Tile_X5Y1_N4BEG[4] ,
    \Tile_X5Y1_N4BEG[3] ,
    \Tile_X5Y1_N4BEG[2] ,
    \Tile_X5Y1_N4BEG[1] ,
    \Tile_X5Y1_N4BEG[0] }),
    .NN4END({\Tile_X5Y1_NN4BEG[15] ,
    \Tile_X5Y1_NN4BEG[14] ,
    \Tile_X5Y1_NN4BEG[13] ,
    \Tile_X5Y1_NN4BEG[12] ,
    \Tile_X5Y1_NN4BEG[11] ,
    \Tile_X5Y1_NN4BEG[10] ,
    \Tile_X5Y1_NN4BEG[9] ,
    \Tile_X5Y1_NN4BEG[8] ,
    \Tile_X5Y1_NN4BEG[7] ,
    \Tile_X5Y1_NN4BEG[6] ,
    \Tile_X5Y1_NN4BEG[5] ,
    \Tile_X5Y1_NN4BEG[4] ,
    \Tile_X5Y1_NN4BEG[3] ,
    \Tile_X5Y1_NN4BEG[2] ,
    \Tile_X5Y1_NN4BEG[1] ,
    \Tile_X5Y1_NN4BEG[0] }),
    .S1BEG({\Tile_X5Y0_S1BEG[3] ,
    \Tile_X5Y0_S1BEG[2] ,
    \Tile_X5Y0_S1BEG[1] ,
    \Tile_X5Y0_S1BEG[0] }),
    .S2BEG({\Tile_X5Y0_S2BEG[7] ,
    \Tile_X5Y0_S2BEG[6] ,
    \Tile_X5Y0_S2BEG[5] ,
    \Tile_X5Y0_S2BEG[4] ,
    \Tile_X5Y0_S2BEG[3] ,
    \Tile_X5Y0_S2BEG[2] ,
    \Tile_X5Y0_S2BEG[1] ,
    \Tile_X5Y0_S2BEG[0] }),
    .S2BEGb({\Tile_X5Y0_S2BEGb[7] ,
    \Tile_X5Y0_S2BEGb[6] ,
    \Tile_X5Y0_S2BEGb[5] ,
    \Tile_X5Y0_S2BEGb[4] ,
    \Tile_X5Y0_S2BEGb[3] ,
    \Tile_X5Y0_S2BEGb[2] ,
    \Tile_X5Y0_S2BEGb[1] ,
    \Tile_X5Y0_S2BEGb[0] }),
    .S4BEG({\Tile_X5Y0_S4BEG[15] ,
    \Tile_X5Y0_S4BEG[14] ,
    \Tile_X5Y0_S4BEG[13] ,
    \Tile_X5Y0_S4BEG[12] ,
    \Tile_X5Y0_S4BEG[11] ,
    \Tile_X5Y0_S4BEG[10] ,
    \Tile_X5Y0_S4BEG[9] ,
    \Tile_X5Y0_S4BEG[8] ,
    \Tile_X5Y0_S4BEG[7] ,
    \Tile_X5Y0_S4BEG[6] ,
    \Tile_X5Y0_S4BEG[5] ,
    \Tile_X5Y0_S4BEG[4] ,
    \Tile_X5Y0_S4BEG[3] ,
    \Tile_X5Y0_S4BEG[2] ,
    \Tile_X5Y0_S4BEG[1] ,
    \Tile_X5Y0_S4BEG[0] }),
    .SS4BEG({\Tile_X5Y0_SS4BEG[15] ,
    \Tile_X5Y0_SS4BEG[14] ,
    \Tile_X5Y0_SS4BEG[13] ,
    \Tile_X5Y0_SS4BEG[12] ,
    \Tile_X5Y0_SS4BEG[11] ,
    \Tile_X5Y0_SS4BEG[10] ,
    \Tile_X5Y0_SS4BEG[9] ,
    \Tile_X5Y0_SS4BEG[8] ,
    \Tile_X5Y0_SS4BEG[7] ,
    \Tile_X5Y0_SS4BEG[6] ,
    \Tile_X5Y0_SS4BEG[5] ,
    \Tile_X5Y0_SS4BEG[4] ,
    \Tile_X5Y0_SS4BEG[3] ,
    \Tile_X5Y0_SS4BEG[2] ,
    \Tile_X5Y0_SS4BEG[1] ,
    \Tile_X5Y0_SS4BEG[0] }));
 LUT4AB Tile_X5Y10_LUT4AB (.Ci(Tile_X5Y11_Co),
    .Co(Tile_X5Y10_Co),
    .UserCLK(Tile_X5Y11_UserCLKo),
    .UserCLKo(Tile_X5Y10_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X5Y10_E1BEG[3] ,
    \Tile_X5Y10_E1BEG[2] ,
    \Tile_X5Y10_E1BEG[1] ,
    \Tile_X5Y10_E1BEG[0] }),
    .E1END({\Tile_X4Y10_E1BEG[3] ,
    \Tile_X4Y10_E1BEG[2] ,
    \Tile_X4Y10_E1BEG[1] ,
    \Tile_X4Y10_E1BEG[0] }),
    .E2BEG({\Tile_X5Y10_E2BEG[7] ,
    \Tile_X5Y10_E2BEG[6] ,
    \Tile_X5Y10_E2BEG[5] ,
    \Tile_X5Y10_E2BEG[4] ,
    \Tile_X5Y10_E2BEG[3] ,
    \Tile_X5Y10_E2BEG[2] ,
    \Tile_X5Y10_E2BEG[1] ,
    \Tile_X5Y10_E2BEG[0] }),
    .E2BEGb({\Tile_X5Y10_E2BEGb[7] ,
    \Tile_X5Y10_E2BEGb[6] ,
    \Tile_X5Y10_E2BEGb[5] ,
    \Tile_X5Y10_E2BEGb[4] ,
    \Tile_X5Y10_E2BEGb[3] ,
    \Tile_X5Y10_E2BEGb[2] ,
    \Tile_X5Y10_E2BEGb[1] ,
    \Tile_X5Y10_E2BEGb[0] }),
    .E2END({\Tile_X4Y10_E2BEGb[7] ,
    \Tile_X4Y10_E2BEGb[6] ,
    \Tile_X4Y10_E2BEGb[5] ,
    \Tile_X4Y10_E2BEGb[4] ,
    \Tile_X4Y10_E2BEGb[3] ,
    \Tile_X4Y10_E2BEGb[2] ,
    \Tile_X4Y10_E2BEGb[1] ,
    \Tile_X4Y10_E2BEGb[0] }),
    .E2MID({\Tile_X4Y10_E2BEG[7] ,
    \Tile_X4Y10_E2BEG[6] ,
    \Tile_X4Y10_E2BEG[5] ,
    \Tile_X4Y10_E2BEG[4] ,
    \Tile_X4Y10_E2BEG[3] ,
    \Tile_X4Y10_E2BEG[2] ,
    \Tile_X4Y10_E2BEG[1] ,
    \Tile_X4Y10_E2BEG[0] }),
    .E6BEG({\Tile_X5Y10_E6BEG[11] ,
    \Tile_X5Y10_E6BEG[10] ,
    \Tile_X5Y10_E6BEG[9] ,
    \Tile_X5Y10_E6BEG[8] ,
    \Tile_X5Y10_E6BEG[7] ,
    \Tile_X5Y10_E6BEG[6] ,
    \Tile_X5Y10_E6BEG[5] ,
    \Tile_X5Y10_E6BEG[4] ,
    \Tile_X5Y10_E6BEG[3] ,
    \Tile_X5Y10_E6BEG[2] ,
    \Tile_X5Y10_E6BEG[1] ,
    \Tile_X5Y10_E6BEG[0] }),
    .E6END({\Tile_X4Y10_E6BEG[11] ,
    \Tile_X4Y10_E6BEG[10] ,
    \Tile_X4Y10_E6BEG[9] ,
    \Tile_X4Y10_E6BEG[8] ,
    \Tile_X4Y10_E6BEG[7] ,
    \Tile_X4Y10_E6BEG[6] ,
    \Tile_X4Y10_E6BEG[5] ,
    \Tile_X4Y10_E6BEG[4] ,
    \Tile_X4Y10_E6BEG[3] ,
    \Tile_X4Y10_E6BEG[2] ,
    \Tile_X4Y10_E6BEG[1] ,
    \Tile_X4Y10_E6BEG[0] }),
    .EE4BEG({\Tile_X5Y10_EE4BEG[15] ,
    \Tile_X5Y10_EE4BEG[14] ,
    \Tile_X5Y10_EE4BEG[13] ,
    \Tile_X5Y10_EE4BEG[12] ,
    \Tile_X5Y10_EE4BEG[11] ,
    \Tile_X5Y10_EE4BEG[10] ,
    \Tile_X5Y10_EE4BEG[9] ,
    \Tile_X5Y10_EE4BEG[8] ,
    \Tile_X5Y10_EE4BEG[7] ,
    \Tile_X5Y10_EE4BEG[6] ,
    \Tile_X5Y10_EE4BEG[5] ,
    \Tile_X5Y10_EE4BEG[4] ,
    \Tile_X5Y10_EE4BEG[3] ,
    \Tile_X5Y10_EE4BEG[2] ,
    \Tile_X5Y10_EE4BEG[1] ,
    \Tile_X5Y10_EE4BEG[0] }),
    .EE4END({\Tile_X4Y10_EE4BEG[15] ,
    \Tile_X4Y10_EE4BEG[14] ,
    \Tile_X4Y10_EE4BEG[13] ,
    \Tile_X4Y10_EE4BEG[12] ,
    \Tile_X4Y10_EE4BEG[11] ,
    \Tile_X4Y10_EE4BEG[10] ,
    \Tile_X4Y10_EE4BEG[9] ,
    \Tile_X4Y10_EE4BEG[8] ,
    \Tile_X4Y10_EE4BEG[7] ,
    \Tile_X4Y10_EE4BEG[6] ,
    \Tile_X4Y10_EE4BEG[5] ,
    \Tile_X4Y10_EE4BEG[4] ,
    \Tile_X4Y10_EE4BEG[3] ,
    \Tile_X4Y10_EE4BEG[2] ,
    \Tile_X4Y10_EE4BEG[1] ,
    \Tile_X4Y10_EE4BEG[0] }),
    .FrameData({\Tile_X4Y10_FrameData_O[31] ,
    \Tile_X4Y10_FrameData_O[30] ,
    \Tile_X4Y10_FrameData_O[29] ,
    \Tile_X4Y10_FrameData_O[28] ,
    \Tile_X4Y10_FrameData_O[27] ,
    \Tile_X4Y10_FrameData_O[26] ,
    \Tile_X4Y10_FrameData_O[25] ,
    \Tile_X4Y10_FrameData_O[24] ,
    \Tile_X4Y10_FrameData_O[23] ,
    \Tile_X4Y10_FrameData_O[22] ,
    \Tile_X4Y10_FrameData_O[21] ,
    \Tile_X4Y10_FrameData_O[20] ,
    \Tile_X4Y10_FrameData_O[19] ,
    \Tile_X4Y10_FrameData_O[18] ,
    \Tile_X4Y10_FrameData_O[17] ,
    \Tile_X4Y10_FrameData_O[16] ,
    \Tile_X4Y10_FrameData_O[15] ,
    \Tile_X4Y10_FrameData_O[14] ,
    \Tile_X4Y10_FrameData_O[13] ,
    \Tile_X4Y10_FrameData_O[12] ,
    \Tile_X4Y10_FrameData_O[11] ,
    \Tile_X4Y10_FrameData_O[10] ,
    \Tile_X4Y10_FrameData_O[9] ,
    \Tile_X4Y10_FrameData_O[8] ,
    \Tile_X4Y10_FrameData_O[7] ,
    \Tile_X4Y10_FrameData_O[6] ,
    \Tile_X4Y10_FrameData_O[5] ,
    \Tile_X4Y10_FrameData_O[4] ,
    \Tile_X4Y10_FrameData_O[3] ,
    \Tile_X4Y10_FrameData_O[2] ,
    \Tile_X4Y10_FrameData_O[1] ,
    \Tile_X4Y10_FrameData_O[0] }),
    .FrameData_O({\Tile_X5Y10_FrameData_O[31] ,
    \Tile_X5Y10_FrameData_O[30] ,
    \Tile_X5Y10_FrameData_O[29] ,
    \Tile_X5Y10_FrameData_O[28] ,
    \Tile_X5Y10_FrameData_O[27] ,
    \Tile_X5Y10_FrameData_O[26] ,
    \Tile_X5Y10_FrameData_O[25] ,
    \Tile_X5Y10_FrameData_O[24] ,
    \Tile_X5Y10_FrameData_O[23] ,
    \Tile_X5Y10_FrameData_O[22] ,
    \Tile_X5Y10_FrameData_O[21] ,
    \Tile_X5Y10_FrameData_O[20] ,
    \Tile_X5Y10_FrameData_O[19] ,
    \Tile_X5Y10_FrameData_O[18] ,
    \Tile_X5Y10_FrameData_O[17] ,
    \Tile_X5Y10_FrameData_O[16] ,
    \Tile_X5Y10_FrameData_O[15] ,
    \Tile_X5Y10_FrameData_O[14] ,
    \Tile_X5Y10_FrameData_O[13] ,
    \Tile_X5Y10_FrameData_O[12] ,
    \Tile_X5Y10_FrameData_O[11] ,
    \Tile_X5Y10_FrameData_O[10] ,
    \Tile_X5Y10_FrameData_O[9] ,
    \Tile_X5Y10_FrameData_O[8] ,
    \Tile_X5Y10_FrameData_O[7] ,
    \Tile_X5Y10_FrameData_O[6] ,
    \Tile_X5Y10_FrameData_O[5] ,
    \Tile_X5Y10_FrameData_O[4] ,
    \Tile_X5Y10_FrameData_O[3] ,
    \Tile_X5Y10_FrameData_O[2] ,
    \Tile_X5Y10_FrameData_O[1] ,
    \Tile_X5Y10_FrameData_O[0] }),
    .FrameStrobe({\Tile_X5Y11_FrameStrobe_O[19] ,
    \Tile_X5Y11_FrameStrobe_O[18] ,
    \Tile_X5Y11_FrameStrobe_O[17] ,
    \Tile_X5Y11_FrameStrobe_O[16] ,
    \Tile_X5Y11_FrameStrobe_O[15] ,
    \Tile_X5Y11_FrameStrobe_O[14] ,
    \Tile_X5Y11_FrameStrobe_O[13] ,
    \Tile_X5Y11_FrameStrobe_O[12] ,
    \Tile_X5Y11_FrameStrobe_O[11] ,
    \Tile_X5Y11_FrameStrobe_O[10] ,
    \Tile_X5Y11_FrameStrobe_O[9] ,
    \Tile_X5Y11_FrameStrobe_O[8] ,
    \Tile_X5Y11_FrameStrobe_O[7] ,
    \Tile_X5Y11_FrameStrobe_O[6] ,
    \Tile_X5Y11_FrameStrobe_O[5] ,
    \Tile_X5Y11_FrameStrobe_O[4] ,
    \Tile_X5Y11_FrameStrobe_O[3] ,
    \Tile_X5Y11_FrameStrobe_O[2] ,
    \Tile_X5Y11_FrameStrobe_O[1] ,
    \Tile_X5Y11_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X5Y10_FrameStrobe_O[19] ,
    \Tile_X5Y10_FrameStrobe_O[18] ,
    \Tile_X5Y10_FrameStrobe_O[17] ,
    \Tile_X5Y10_FrameStrobe_O[16] ,
    \Tile_X5Y10_FrameStrobe_O[15] ,
    \Tile_X5Y10_FrameStrobe_O[14] ,
    \Tile_X5Y10_FrameStrobe_O[13] ,
    \Tile_X5Y10_FrameStrobe_O[12] ,
    \Tile_X5Y10_FrameStrobe_O[11] ,
    \Tile_X5Y10_FrameStrobe_O[10] ,
    \Tile_X5Y10_FrameStrobe_O[9] ,
    \Tile_X5Y10_FrameStrobe_O[8] ,
    \Tile_X5Y10_FrameStrobe_O[7] ,
    \Tile_X5Y10_FrameStrobe_O[6] ,
    \Tile_X5Y10_FrameStrobe_O[5] ,
    \Tile_X5Y10_FrameStrobe_O[4] ,
    \Tile_X5Y10_FrameStrobe_O[3] ,
    \Tile_X5Y10_FrameStrobe_O[2] ,
    \Tile_X5Y10_FrameStrobe_O[1] ,
    \Tile_X5Y10_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X5Y10_N1BEG[3] ,
    \Tile_X5Y10_N1BEG[2] ,
    \Tile_X5Y10_N1BEG[1] ,
    \Tile_X5Y10_N1BEG[0] }),
    .N1END({\Tile_X5Y11_N1BEG[3] ,
    \Tile_X5Y11_N1BEG[2] ,
    \Tile_X5Y11_N1BEG[1] ,
    \Tile_X5Y11_N1BEG[0] }),
    .N2BEG({\Tile_X5Y10_N2BEG[7] ,
    \Tile_X5Y10_N2BEG[6] ,
    \Tile_X5Y10_N2BEG[5] ,
    \Tile_X5Y10_N2BEG[4] ,
    \Tile_X5Y10_N2BEG[3] ,
    \Tile_X5Y10_N2BEG[2] ,
    \Tile_X5Y10_N2BEG[1] ,
    \Tile_X5Y10_N2BEG[0] }),
    .N2BEGb({\Tile_X5Y10_N2BEGb[7] ,
    \Tile_X5Y10_N2BEGb[6] ,
    \Tile_X5Y10_N2BEGb[5] ,
    \Tile_X5Y10_N2BEGb[4] ,
    \Tile_X5Y10_N2BEGb[3] ,
    \Tile_X5Y10_N2BEGb[2] ,
    \Tile_X5Y10_N2BEGb[1] ,
    \Tile_X5Y10_N2BEGb[0] }),
    .N2END({\Tile_X5Y11_N2BEGb[7] ,
    \Tile_X5Y11_N2BEGb[6] ,
    \Tile_X5Y11_N2BEGb[5] ,
    \Tile_X5Y11_N2BEGb[4] ,
    \Tile_X5Y11_N2BEGb[3] ,
    \Tile_X5Y11_N2BEGb[2] ,
    \Tile_X5Y11_N2BEGb[1] ,
    \Tile_X5Y11_N2BEGb[0] }),
    .N2MID({\Tile_X5Y11_N2BEG[7] ,
    \Tile_X5Y11_N2BEG[6] ,
    \Tile_X5Y11_N2BEG[5] ,
    \Tile_X5Y11_N2BEG[4] ,
    \Tile_X5Y11_N2BEG[3] ,
    \Tile_X5Y11_N2BEG[2] ,
    \Tile_X5Y11_N2BEG[1] ,
    \Tile_X5Y11_N2BEG[0] }),
    .N4BEG({\Tile_X5Y10_N4BEG[15] ,
    \Tile_X5Y10_N4BEG[14] ,
    \Tile_X5Y10_N4BEG[13] ,
    \Tile_X5Y10_N4BEG[12] ,
    \Tile_X5Y10_N4BEG[11] ,
    \Tile_X5Y10_N4BEG[10] ,
    \Tile_X5Y10_N4BEG[9] ,
    \Tile_X5Y10_N4BEG[8] ,
    \Tile_X5Y10_N4BEG[7] ,
    \Tile_X5Y10_N4BEG[6] ,
    \Tile_X5Y10_N4BEG[5] ,
    \Tile_X5Y10_N4BEG[4] ,
    \Tile_X5Y10_N4BEG[3] ,
    \Tile_X5Y10_N4BEG[2] ,
    \Tile_X5Y10_N4BEG[1] ,
    \Tile_X5Y10_N4BEG[0] }),
    .N4END({\Tile_X5Y11_N4BEG[15] ,
    \Tile_X5Y11_N4BEG[14] ,
    \Tile_X5Y11_N4BEG[13] ,
    \Tile_X5Y11_N4BEG[12] ,
    \Tile_X5Y11_N4BEG[11] ,
    \Tile_X5Y11_N4BEG[10] ,
    \Tile_X5Y11_N4BEG[9] ,
    \Tile_X5Y11_N4BEG[8] ,
    \Tile_X5Y11_N4BEG[7] ,
    \Tile_X5Y11_N4BEG[6] ,
    \Tile_X5Y11_N4BEG[5] ,
    \Tile_X5Y11_N4BEG[4] ,
    \Tile_X5Y11_N4BEG[3] ,
    \Tile_X5Y11_N4BEG[2] ,
    \Tile_X5Y11_N4BEG[1] ,
    \Tile_X5Y11_N4BEG[0] }),
    .NN4BEG({\Tile_X5Y10_NN4BEG[15] ,
    \Tile_X5Y10_NN4BEG[14] ,
    \Tile_X5Y10_NN4BEG[13] ,
    \Tile_X5Y10_NN4BEG[12] ,
    \Tile_X5Y10_NN4BEG[11] ,
    \Tile_X5Y10_NN4BEG[10] ,
    \Tile_X5Y10_NN4BEG[9] ,
    \Tile_X5Y10_NN4BEG[8] ,
    \Tile_X5Y10_NN4BEG[7] ,
    \Tile_X5Y10_NN4BEG[6] ,
    \Tile_X5Y10_NN4BEG[5] ,
    \Tile_X5Y10_NN4BEG[4] ,
    \Tile_X5Y10_NN4BEG[3] ,
    \Tile_X5Y10_NN4BEG[2] ,
    \Tile_X5Y10_NN4BEG[1] ,
    \Tile_X5Y10_NN4BEG[0] }),
    .NN4END({\Tile_X5Y11_NN4BEG[15] ,
    \Tile_X5Y11_NN4BEG[14] ,
    \Tile_X5Y11_NN4BEG[13] ,
    \Tile_X5Y11_NN4BEG[12] ,
    \Tile_X5Y11_NN4BEG[11] ,
    \Tile_X5Y11_NN4BEG[10] ,
    \Tile_X5Y11_NN4BEG[9] ,
    \Tile_X5Y11_NN4BEG[8] ,
    \Tile_X5Y11_NN4BEG[7] ,
    \Tile_X5Y11_NN4BEG[6] ,
    \Tile_X5Y11_NN4BEG[5] ,
    \Tile_X5Y11_NN4BEG[4] ,
    \Tile_X5Y11_NN4BEG[3] ,
    \Tile_X5Y11_NN4BEG[2] ,
    \Tile_X5Y11_NN4BEG[1] ,
    \Tile_X5Y11_NN4BEG[0] }),
    .S1BEG({\Tile_X5Y10_S1BEG[3] ,
    \Tile_X5Y10_S1BEG[2] ,
    \Tile_X5Y10_S1BEG[1] ,
    \Tile_X5Y10_S1BEG[0] }),
    .S1END({\Tile_X5Y9_S1BEG[3] ,
    \Tile_X5Y9_S1BEG[2] ,
    \Tile_X5Y9_S1BEG[1] ,
    \Tile_X5Y9_S1BEG[0] }),
    .S2BEG({\Tile_X5Y10_S2BEG[7] ,
    \Tile_X5Y10_S2BEG[6] ,
    \Tile_X5Y10_S2BEG[5] ,
    \Tile_X5Y10_S2BEG[4] ,
    \Tile_X5Y10_S2BEG[3] ,
    \Tile_X5Y10_S2BEG[2] ,
    \Tile_X5Y10_S2BEG[1] ,
    \Tile_X5Y10_S2BEG[0] }),
    .S2BEGb({\Tile_X5Y10_S2BEGb[7] ,
    \Tile_X5Y10_S2BEGb[6] ,
    \Tile_X5Y10_S2BEGb[5] ,
    \Tile_X5Y10_S2BEGb[4] ,
    \Tile_X5Y10_S2BEGb[3] ,
    \Tile_X5Y10_S2BEGb[2] ,
    \Tile_X5Y10_S2BEGb[1] ,
    \Tile_X5Y10_S2BEGb[0] }),
    .S2END({\Tile_X5Y9_S2BEGb[7] ,
    \Tile_X5Y9_S2BEGb[6] ,
    \Tile_X5Y9_S2BEGb[5] ,
    \Tile_X5Y9_S2BEGb[4] ,
    \Tile_X5Y9_S2BEGb[3] ,
    \Tile_X5Y9_S2BEGb[2] ,
    \Tile_X5Y9_S2BEGb[1] ,
    \Tile_X5Y9_S2BEGb[0] }),
    .S2MID({\Tile_X5Y9_S2BEG[7] ,
    \Tile_X5Y9_S2BEG[6] ,
    \Tile_X5Y9_S2BEG[5] ,
    \Tile_X5Y9_S2BEG[4] ,
    \Tile_X5Y9_S2BEG[3] ,
    \Tile_X5Y9_S2BEG[2] ,
    \Tile_X5Y9_S2BEG[1] ,
    \Tile_X5Y9_S2BEG[0] }),
    .S4BEG({\Tile_X5Y10_S4BEG[15] ,
    \Tile_X5Y10_S4BEG[14] ,
    \Tile_X5Y10_S4BEG[13] ,
    \Tile_X5Y10_S4BEG[12] ,
    \Tile_X5Y10_S4BEG[11] ,
    \Tile_X5Y10_S4BEG[10] ,
    \Tile_X5Y10_S4BEG[9] ,
    \Tile_X5Y10_S4BEG[8] ,
    \Tile_X5Y10_S4BEG[7] ,
    \Tile_X5Y10_S4BEG[6] ,
    \Tile_X5Y10_S4BEG[5] ,
    \Tile_X5Y10_S4BEG[4] ,
    \Tile_X5Y10_S4BEG[3] ,
    \Tile_X5Y10_S4BEG[2] ,
    \Tile_X5Y10_S4BEG[1] ,
    \Tile_X5Y10_S4BEG[0] }),
    .S4END({\Tile_X5Y9_S4BEG[15] ,
    \Tile_X5Y9_S4BEG[14] ,
    \Tile_X5Y9_S4BEG[13] ,
    \Tile_X5Y9_S4BEG[12] ,
    \Tile_X5Y9_S4BEG[11] ,
    \Tile_X5Y9_S4BEG[10] ,
    \Tile_X5Y9_S4BEG[9] ,
    \Tile_X5Y9_S4BEG[8] ,
    \Tile_X5Y9_S4BEG[7] ,
    \Tile_X5Y9_S4BEG[6] ,
    \Tile_X5Y9_S4BEG[5] ,
    \Tile_X5Y9_S4BEG[4] ,
    \Tile_X5Y9_S4BEG[3] ,
    \Tile_X5Y9_S4BEG[2] ,
    \Tile_X5Y9_S4BEG[1] ,
    \Tile_X5Y9_S4BEG[0] }),
    .SS4BEG({\Tile_X5Y10_SS4BEG[15] ,
    \Tile_X5Y10_SS4BEG[14] ,
    \Tile_X5Y10_SS4BEG[13] ,
    \Tile_X5Y10_SS4BEG[12] ,
    \Tile_X5Y10_SS4BEG[11] ,
    \Tile_X5Y10_SS4BEG[10] ,
    \Tile_X5Y10_SS4BEG[9] ,
    \Tile_X5Y10_SS4BEG[8] ,
    \Tile_X5Y10_SS4BEG[7] ,
    \Tile_X5Y10_SS4BEG[6] ,
    \Tile_X5Y10_SS4BEG[5] ,
    \Tile_X5Y10_SS4BEG[4] ,
    \Tile_X5Y10_SS4BEG[3] ,
    \Tile_X5Y10_SS4BEG[2] ,
    \Tile_X5Y10_SS4BEG[1] ,
    \Tile_X5Y10_SS4BEG[0] }),
    .SS4END({\Tile_X5Y9_SS4BEG[15] ,
    \Tile_X5Y9_SS4BEG[14] ,
    \Tile_X5Y9_SS4BEG[13] ,
    \Tile_X5Y9_SS4BEG[12] ,
    \Tile_X5Y9_SS4BEG[11] ,
    \Tile_X5Y9_SS4BEG[10] ,
    \Tile_X5Y9_SS4BEG[9] ,
    \Tile_X5Y9_SS4BEG[8] ,
    \Tile_X5Y9_SS4BEG[7] ,
    \Tile_X5Y9_SS4BEG[6] ,
    \Tile_X5Y9_SS4BEG[5] ,
    \Tile_X5Y9_SS4BEG[4] ,
    \Tile_X5Y9_SS4BEG[3] ,
    \Tile_X5Y9_SS4BEG[2] ,
    \Tile_X5Y9_SS4BEG[1] ,
    \Tile_X5Y9_SS4BEG[0] }),
    .W1BEG({\Tile_X5Y10_W1BEG[3] ,
    \Tile_X5Y10_W1BEG[2] ,
    \Tile_X5Y10_W1BEG[1] ,
    \Tile_X5Y10_W1BEG[0] }),
    .W1END({\Tile_X6Y10_W1BEG[3] ,
    \Tile_X6Y10_W1BEG[2] ,
    \Tile_X6Y10_W1BEG[1] ,
    \Tile_X6Y10_W1BEG[0] }),
    .W2BEG({\Tile_X5Y10_W2BEG[7] ,
    \Tile_X5Y10_W2BEG[6] ,
    \Tile_X5Y10_W2BEG[5] ,
    \Tile_X5Y10_W2BEG[4] ,
    \Tile_X5Y10_W2BEG[3] ,
    \Tile_X5Y10_W2BEG[2] ,
    \Tile_X5Y10_W2BEG[1] ,
    \Tile_X5Y10_W2BEG[0] }),
    .W2BEGb({\Tile_X5Y10_W2BEGb[7] ,
    \Tile_X5Y10_W2BEGb[6] ,
    \Tile_X5Y10_W2BEGb[5] ,
    \Tile_X5Y10_W2BEGb[4] ,
    \Tile_X5Y10_W2BEGb[3] ,
    \Tile_X5Y10_W2BEGb[2] ,
    \Tile_X5Y10_W2BEGb[1] ,
    \Tile_X5Y10_W2BEGb[0] }),
    .W2END({\Tile_X6Y10_W2BEGb[7] ,
    \Tile_X6Y10_W2BEGb[6] ,
    \Tile_X6Y10_W2BEGb[5] ,
    \Tile_X6Y10_W2BEGb[4] ,
    \Tile_X6Y10_W2BEGb[3] ,
    \Tile_X6Y10_W2BEGb[2] ,
    \Tile_X6Y10_W2BEGb[1] ,
    \Tile_X6Y10_W2BEGb[0] }),
    .W2MID({\Tile_X6Y10_W2BEG[7] ,
    \Tile_X6Y10_W2BEG[6] ,
    \Tile_X6Y10_W2BEG[5] ,
    \Tile_X6Y10_W2BEG[4] ,
    \Tile_X6Y10_W2BEG[3] ,
    \Tile_X6Y10_W2BEG[2] ,
    \Tile_X6Y10_W2BEG[1] ,
    \Tile_X6Y10_W2BEG[0] }),
    .W6BEG({\Tile_X5Y10_W6BEG[11] ,
    \Tile_X5Y10_W6BEG[10] ,
    \Tile_X5Y10_W6BEG[9] ,
    \Tile_X5Y10_W6BEG[8] ,
    \Tile_X5Y10_W6BEG[7] ,
    \Tile_X5Y10_W6BEG[6] ,
    \Tile_X5Y10_W6BEG[5] ,
    \Tile_X5Y10_W6BEG[4] ,
    \Tile_X5Y10_W6BEG[3] ,
    \Tile_X5Y10_W6BEG[2] ,
    \Tile_X5Y10_W6BEG[1] ,
    \Tile_X5Y10_W6BEG[0] }),
    .W6END({\Tile_X6Y10_W6BEG[11] ,
    \Tile_X6Y10_W6BEG[10] ,
    \Tile_X6Y10_W6BEG[9] ,
    \Tile_X6Y10_W6BEG[8] ,
    \Tile_X6Y10_W6BEG[7] ,
    \Tile_X6Y10_W6BEG[6] ,
    \Tile_X6Y10_W6BEG[5] ,
    \Tile_X6Y10_W6BEG[4] ,
    \Tile_X6Y10_W6BEG[3] ,
    \Tile_X6Y10_W6BEG[2] ,
    \Tile_X6Y10_W6BEG[1] ,
    \Tile_X6Y10_W6BEG[0] }),
    .WW4BEG({\Tile_X5Y10_WW4BEG[15] ,
    \Tile_X5Y10_WW4BEG[14] ,
    \Tile_X5Y10_WW4BEG[13] ,
    \Tile_X5Y10_WW4BEG[12] ,
    \Tile_X5Y10_WW4BEG[11] ,
    \Tile_X5Y10_WW4BEG[10] ,
    \Tile_X5Y10_WW4BEG[9] ,
    \Tile_X5Y10_WW4BEG[8] ,
    \Tile_X5Y10_WW4BEG[7] ,
    \Tile_X5Y10_WW4BEG[6] ,
    \Tile_X5Y10_WW4BEG[5] ,
    \Tile_X5Y10_WW4BEG[4] ,
    \Tile_X5Y10_WW4BEG[3] ,
    \Tile_X5Y10_WW4BEG[2] ,
    \Tile_X5Y10_WW4BEG[1] ,
    \Tile_X5Y10_WW4BEG[0] }),
    .WW4END({\Tile_X6Y10_WW4BEG[15] ,
    \Tile_X6Y10_WW4BEG[14] ,
    \Tile_X6Y10_WW4BEG[13] ,
    \Tile_X6Y10_WW4BEG[12] ,
    \Tile_X6Y10_WW4BEG[11] ,
    \Tile_X6Y10_WW4BEG[10] ,
    \Tile_X6Y10_WW4BEG[9] ,
    \Tile_X6Y10_WW4BEG[8] ,
    \Tile_X6Y10_WW4BEG[7] ,
    \Tile_X6Y10_WW4BEG[6] ,
    \Tile_X6Y10_WW4BEG[5] ,
    \Tile_X6Y10_WW4BEG[4] ,
    \Tile_X6Y10_WW4BEG[3] ,
    \Tile_X6Y10_WW4BEG[2] ,
    \Tile_X6Y10_WW4BEG[1] ,
    \Tile_X6Y10_WW4BEG[0] }));
 LUT4AB Tile_X5Y11_LUT4AB (.Ci(Tile_X5Y12_Co),
    .Co(Tile_X5Y11_Co),
    .UserCLK(Tile_X5Y12_UserCLKo),
    .UserCLKo(Tile_X5Y11_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X5Y11_E1BEG[3] ,
    \Tile_X5Y11_E1BEG[2] ,
    \Tile_X5Y11_E1BEG[1] ,
    \Tile_X5Y11_E1BEG[0] }),
    .E1END({\Tile_X4Y11_E1BEG[3] ,
    \Tile_X4Y11_E1BEG[2] ,
    \Tile_X4Y11_E1BEG[1] ,
    \Tile_X4Y11_E1BEG[0] }),
    .E2BEG({\Tile_X5Y11_E2BEG[7] ,
    \Tile_X5Y11_E2BEG[6] ,
    \Tile_X5Y11_E2BEG[5] ,
    \Tile_X5Y11_E2BEG[4] ,
    \Tile_X5Y11_E2BEG[3] ,
    \Tile_X5Y11_E2BEG[2] ,
    \Tile_X5Y11_E2BEG[1] ,
    \Tile_X5Y11_E2BEG[0] }),
    .E2BEGb({\Tile_X5Y11_E2BEGb[7] ,
    \Tile_X5Y11_E2BEGb[6] ,
    \Tile_X5Y11_E2BEGb[5] ,
    \Tile_X5Y11_E2BEGb[4] ,
    \Tile_X5Y11_E2BEGb[3] ,
    \Tile_X5Y11_E2BEGb[2] ,
    \Tile_X5Y11_E2BEGb[1] ,
    \Tile_X5Y11_E2BEGb[0] }),
    .E2END({\Tile_X4Y11_E2BEGb[7] ,
    \Tile_X4Y11_E2BEGb[6] ,
    \Tile_X4Y11_E2BEGb[5] ,
    \Tile_X4Y11_E2BEGb[4] ,
    \Tile_X4Y11_E2BEGb[3] ,
    \Tile_X4Y11_E2BEGb[2] ,
    \Tile_X4Y11_E2BEGb[1] ,
    \Tile_X4Y11_E2BEGb[0] }),
    .E2MID({\Tile_X4Y11_E2BEG[7] ,
    \Tile_X4Y11_E2BEG[6] ,
    \Tile_X4Y11_E2BEG[5] ,
    \Tile_X4Y11_E2BEG[4] ,
    \Tile_X4Y11_E2BEG[3] ,
    \Tile_X4Y11_E2BEG[2] ,
    \Tile_X4Y11_E2BEG[1] ,
    \Tile_X4Y11_E2BEG[0] }),
    .E6BEG({\Tile_X5Y11_E6BEG[11] ,
    \Tile_X5Y11_E6BEG[10] ,
    \Tile_X5Y11_E6BEG[9] ,
    \Tile_X5Y11_E6BEG[8] ,
    \Tile_X5Y11_E6BEG[7] ,
    \Tile_X5Y11_E6BEG[6] ,
    \Tile_X5Y11_E6BEG[5] ,
    \Tile_X5Y11_E6BEG[4] ,
    \Tile_X5Y11_E6BEG[3] ,
    \Tile_X5Y11_E6BEG[2] ,
    \Tile_X5Y11_E6BEG[1] ,
    \Tile_X5Y11_E6BEG[0] }),
    .E6END({\Tile_X4Y11_E6BEG[11] ,
    \Tile_X4Y11_E6BEG[10] ,
    \Tile_X4Y11_E6BEG[9] ,
    \Tile_X4Y11_E6BEG[8] ,
    \Tile_X4Y11_E6BEG[7] ,
    \Tile_X4Y11_E6BEG[6] ,
    \Tile_X4Y11_E6BEG[5] ,
    \Tile_X4Y11_E6BEG[4] ,
    \Tile_X4Y11_E6BEG[3] ,
    \Tile_X4Y11_E6BEG[2] ,
    \Tile_X4Y11_E6BEG[1] ,
    \Tile_X4Y11_E6BEG[0] }),
    .EE4BEG({\Tile_X5Y11_EE4BEG[15] ,
    \Tile_X5Y11_EE4BEG[14] ,
    \Tile_X5Y11_EE4BEG[13] ,
    \Tile_X5Y11_EE4BEG[12] ,
    \Tile_X5Y11_EE4BEG[11] ,
    \Tile_X5Y11_EE4BEG[10] ,
    \Tile_X5Y11_EE4BEG[9] ,
    \Tile_X5Y11_EE4BEG[8] ,
    \Tile_X5Y11_EE4BEG[7] ,
    \Tile_X5Y11_EE4BEG[6] ,
    \Tile_X5Y11_EE4BEG[5] ,
    \Tile_X5Y11_EE4BEG[4] ,
    \Tile_X5Y11_EE4BEG[3] ,
    \Tile_X5Y11_EE4BEG[2] ,
    \Tile_X5Y11_EE4BEG[1] ,
    \Tile_X5Y11_EE4BEG[0] }),
    .EE4END({\Tile_X4Y11_EE4BEG[15] ,
    \Tile_X4Y11_EE4BEG[14] ,
    \Tile_X4Y11_EE4BEG[13] ,
    \Tile_X4Y11_EE4BEG[12] ,
    \Tile_X4Y11_EE4BEG[11] ,
    \Tile_X4Y11_EE4BEG[10] ,
    \Tile_X4Y11_EE4BEG[9] ,
    \Tile_X4Y11_EE4BEG[8] ,
    \Tile_X4Y11_EE4BEG[7] ,
    \Tile_X4Y11_EE4BEG[6] ,
    \Tile_X4Y11_EE4BEG[5] ,
    \Tile_X4Y11_EE4BEG[4] ,
    \Tile_X4Y11_EE4BEG[3] ,
    \Tile_X4Y11_EE4BEG[2] ,
    \Tile_X4Y11_EE4BEG[1] ,
    \Tile_X4Y11_EE4BEG[0] }),
    .FrameData({\Tile_X4Y11_FrameData_O[31] ,
    \Tile_X4Y11_FrameData_O[30] ,
    \Tile_X4Y11_FrameData_O[29] ,
    \Tile_X4Y11_FrameData_O[28] ,
    \Tile_X4Y11_FrameData_O[27] ,
    \Tile_X4Y11_FrameData_O[26] ,
    \Tile_X4Y11_FrameData_O[25] ,
    \Tile_X4Y11_FrameData_O[24] ,
    \Tile_X4Y11_FrameData_O[23] ,
    \Tile_X4Y11_FrameData_O[22] ,
    \Tile_X4Y11_FrameData_O[21] ,
    \Tile_X4Y11_FrameData_O[20] ,
    \Tile_X4Y11_FrameData_O[19] ,
    \Tile_X4Y11_FrameData_O[18] ,
    \Tile_X4Y11_FrameData_O[17] ,
    \Tile_X4Y11_FrameData_O[16] ,
    \Tile_X4Y11_FrameData_O[15] ,
    \Tile_X4Y11_FrameData_O[14] ,
    \Tile_X4Y11_FrameData_O[13] ,
    \Tile_X4Y11_FrameData_O[12] ,
    \Tile_X4Y11_FrameData_O[11] ,
    \Tile_X4Y11_FrameData_O[10] ,
    \Tile_X4Y11_FrameData_O[9] ,
    \Tile_X4Y11_FrameData_O[8] ,
    \Tile_X4Y11_FrameData_O[7] ,
    \Tile_X4Y11_FrameData_O[6] ,
    \Tile_X4Y11_FrameData_O[5] ,
    \Tile_X4Y11_FrameData_O[4] ,
    \Tile_X4Y11_FrameData_O[3] ,
    \Tile_X4Y11_FrameData_O[2] ,
    \Tile_X4Y11_FrameData_O[1] ,
    \Tile_X4Y11_FrameData_O[0] }),
    .FrameData_O({\Tile_X5Y11_FrameData_O[31] ,
    \Tile_X5Y11_FrameData_O[30] ,
    \Tile_X5Y11_FrameData_O[29] ,
    \Tile_X5Y11_FrameData_O[28] ,
    \Tile_X5Y11_FrameData_O[27] ,
    \Tile_X5Y11_FrameData_O[26] ,
    \Tile_X5Y11_FrameData_O[25] ,
    \Tile_X5Y11_FrameData_O[24] ,
    \Tile_X5Y11_FrameData_O[23] ,
    \Tile_X5Y11_FrameData_O[22] ,
    \Tile_X5Y11_FrameData_O[21] ,
    \Tile_X5Y11_FrameData_O[20] ,
    \Tile_X5Y11_FrameData_O[19] ,
    \Tile_X5Y11_FrameData_O[18] ,
    \Tile_X5Y11_FrameData_O[17] ,
    \Tile_X5Y11_FrameData_O[16] ,
    \Tile_X5Y11_FrameData_O[15] ,
    \Tile_X5Y11_FrameData_O[14] ,
    \Tile_X5Y11_FrameData_O[13] ,
    \Tile_X5Y11_FrameData_O[12] ,
    \Tile_X5Y11_FrameData_O[11] ,
    \Tile_X5Y11_FrameData_O[10] ,
    \Tile_X5Y11_FrameData_O[9] ,
    \Tile_X5Y11_FrameData_O[8] ,
    \Tile_X5Y11_FrameData_O[7] ,
    \Tile_X5Y11_FrameData_O[6] ,
    \Tile_X5Y11_FrameData_O[5] ,
    \Tile_X5Y11_FrameData_O[4] ,
    \Tile_X5Y11_FrameData_O[3] ,
    \Tile_X5Y11_FrameData_O[2] ,
    \Tile_X5Y11_FrameData_O[1] ,
    \Tile_X5Y11_FrameData_O[0] }),
    .FrameStrobe({\Tile_X5Y12_FrameStrobe_O[19] ,
    \Tile_X5Y12_FrameStrobe_O[18] ,
    \Tile_X5Y12_FrameStrobe_O[17] ,
    \Tile_X5Y12_FrameStrobe_O[16] ,
    \Tile_X5Y12_FrameStrobe_O[15] ,
    \Tile_X5Y12_FrameStrobe_O[14] ,
    \Tile_X5Y12_FrameStrobe_O[13] ,
    \Tile_X5Y12_FrameStrobe_O[12] ,
    \Tile_X5Y12_FrameStrobe_O[11] ,
    \Tile_X5Y12_FrameStrobe_O[10] ,
    \Tile_X5Y12_FrameStrobe_O[9] ,
    \Tile_X5Y12_FrameStrobe_O[8] ,
    \Tile_X5Y12_FrameStrobe_O[7] ,
    \Tile_X5Y12_FrameStrobe_O[6] ,
    \Tile_X5Y12_FrameStrobe_O[5] ,
    \Tile_X5Y12_FrameStrobe_O[4] ,
    \Tile_X5Y12_FrameStrobe_O[3] ,
    \Tile_X5Y12_FrameStrobe_O[2] ,
    \Tile_X5Y12_FrameStrobe_O[1] ,
    \Tile_X5Y12_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X5Y11_FrameStrobe_O[19] ,
    \Tile_X5Y11_FrameStrobe_O[18] ,
    \Tile_X5Y11_FrameStrobe_O[17] ,
    \Tile_X5Y11_FrameStrobe_O[16] ,
    \Tile_X5Y11_FrameStrobe_O[15] ,
    \Tile_X5Y11_FrameStrobe_O[14] ,
    \Tile_X5Y11_FrameStrobe_O[13] ,
    \Tile_X5Y11_FrameStrobe_O[12] ,
    \Tile_X5Y11_FrameStrobe_O[11] ,
    \Tile_X5Y11_FrameStrobe_O[10] ,
    \Tile_X5Y11_FrameStrobe_O[9] ,
    \Tile_X5Y11_FrameStrobe_O[8] ,
    \Tile_X5Y11_FrameStrobe_O[7] ,
    \Tile_X5Y11_FrameStrobe_O[6] ,
    \Tile_X5Y11_FrameStrobe_O[5] ,
    \Tile_X5Y11_FrameStrobe_O[4] ,
    \Tile_X5Y11_FrameStrobe_O[3] ,
    \Tile_X5Y11_FrameStrobe_O[2] ,
    \Tile_X5Y11_FrameStrobe_O[1] ,
    \Tile_X5Y11_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X5Y11_N1BEG[3] ,
    \Tile_X5Y11_N1BEG[2] ,
    \Tile_X5Y11_N1BEG[1] ,
    \Tile_X5Y11_N1BEG[0] }),
    .N1END({\Tile_X5Y12_N1BEG[3] ,
    \Tile_X5Y12_N1BEG[2] ,
    \Tile_X5Y12_N1BEG[1] ,
    \Tile_X5Y12_N1BEG[0] }),
    .N2BEG({\Tile_X5Y11_N2BEG[7] ,
    \Tile_X5Y11_N2BEG[6] ,
    \Tile_X5Y11_N2BEG[5] ,
    \Tile_X5Y11_N2BEG[4] ,
    \Tile_X5Y11_N2BEG[3] ,
    \Tile_X5Y11_N2BEG[2] ,
    \Tile_X5Y11_N2BEG[1] ,
    \Tile_X5Y11_N2BEG[0] }),
    .N2BEGb({\Tile_X5Y11_N2BEGb[7] ,
    \Tile_X5Y11_N2BEGb[6] ,
    \Tile_X5Y11_N2BEGb[5] ,
    \Tile_X5Y11_N2BEGb[4] ,
    \Tile_X5Y11_N2BEGb[3] ,
    \Tile_X5Y11_N2BEGb[2] ,
    \Tile_X5Y11_N2BEGb[1] ,
    \Tile_X5Y11_N2BEGb[0] }),
    .N2END({\Tile_X5Y12_N2BEGb[7] ,
    \Tile_X5Y12_N2BEGb[6] ,
    \Tile_X5Y12_N2BEGb[5] ,
    \Tile_X5Y12_N2BEGb[4] ,
    \Tile_X5Y12_N2BEGb[3] ,
    \Tile_X5Y12_N2BEGb[2] ,
    \Tile_X5Y12_N2BEGb[1] ,
    \Tile_X5Y12_N2BEGb[0] }),
    .N2MID({\Tile_X5Y12_N2BEG[7] ,
    \Tile_X5Y12_N2BEG[6] ,
    \Tile_X5Y12_N2BEG[5] ,
    \Tile_X5Y12_N2BEG[4] ,
    \Tile_X5Y12_N2BEG[3] ,
    \Tile_X5Y12_N2BEG[2] ,
    \Tile_X5Y12_N2BEG[1] ,
    \Tile_X5Y12_N2BEG[0] }),
    .N4BEG({\Tile_X5Y11_N4BEG[15] ,
    \Tile_X5Y11_N4BEG[14] ,
    \Tile_X5Y11_N4BEG[13] ,
    \Tile_X5Y11_N4BEG[12] ,
    \Tile_X5Y11_N4BEG[11] ,
    \Tile_X5Y11_N4BEG[10] ,
    \Tile_X5Y11_N4BEG[9] ,
    \Tile_X5Y11_N4BEG[8] ,
    \Tile_X5Y11_N4BEG[7] ,
    \Tile_X5Y11_N4BEG[6] ,
    \Tile_X5Y11_N4BEG[5] ,
    \Tile_X5Y11_N4BEG[4] ,
    \Tile_X5Y11_N4BEG[3] ,
    \Tile_X5Y11_N4BEG[2] ,
    \Tile_X5Y11_N4BEG[1] ,
    \Tile_X5Y11_N4BEG[0] }),
    .N4END({\Tile_X5Y12_N4BEG[15] ,
    \Tile_X5Y12_N4BEG[14] ,
    \Tile_X5Y12_N4BEG[13] ,
    \Tile_X5Y12_N4BEG[12] ,
    \Tile_X5Y12_N4BEG[11] ,
    \Tile_X5Y12_N4BEG[10] ,
    \Tile_X5Y12_N4BEG[9] ,
    \Tile_X5Y12_N4BEG[8] ,
    \Tile_X5Y12_N4BEG[7] ,
    \Tile_X5Y12_N4BEG[6] ,
    \Tile_X5Y12_N4BEG[5] ,
    \Tile_X5Y12_N4BEG[4] ,
    \Tile_X5Y12_N4BEG[3] ,
    \Tile_X5Y12_N4BEG[2] ,
    \Tile_X5Y12_N4BEG[1] ,
    \Tile_X5Y12_N4BEG[0] }),
    .NN4BEG({\Tile_X5Y11_NN4BEG[15] ,
    \Tile_X5Y11_NN4BEG[14] ,
    \Tile_X5Y11_NN4BEG[13] ,
    \Tile_X5Y11_NN4BEG[12] ,
    \Tile_X5Y11_NN4BEG[11] ,
    \Tile_X5Y11_NN4BEG[10] ,
    \Tile_X5Y11_NN4BEG[9] ,
    \Tile_X5Y11_NN4BEG[8] ,
    \Tile_X5Y11_NN4BEG[7] ,
    \Tile_X5Y11_NN4BEG[6] ,
    \Tile_X5Y11_NN4BEG[5] ,
    \Tile_X5Y11_NN4BEG[4] ,
    \Tile_X5Y11_NN4BEG[3] ,
    \Tile_X5Y11_NN4BEG[2] ,
    \Tile_X5Y11_NN4BEG[1] ,
    \Tile_X5Y11_NN4BEG[0] }),
    .NN4END({\Tile_X5Y12_NN4BEG[15] ,
    \Tile_X5Y12_NN4BEG[14] ,
    \Tile_X5Y12_NN4BEG[13] ,
    \Tile_X5Y12_NN4BEG[12] ,
    \Tile_X5Y12_NN4BEG[11] ,
    \Tile_X5Y12_NN4BEG[10] ,
    \Tile_X5Y12_NN4BEG[9] ,
    \Tile_X5Y12_NN4BEG[8] ,
    \Tile_X5Y12_NN4BEG[7] ,
    \Tile_X5Y12_NN4BEG[6] ,
    \Tile_X5Y12_NN4BEG[5] ,
    \Tile_X5Y12_NN4BEG[4] ,
    \Tile_X5Y12_NN4BEG[3] ,
    \Tile_X5Y12_NN4BEG[2] ,
    \Tile_X5Y12_NN4BEG[1] ,
    \Tile_X5Y12_NN4BEG[0] }),
    .S1BEG({\Tile_X5Y11_S1BEG[3] ,
    \Tile_X5Y11_S1BEG[2] ,
    \Tile_X5Y11_S1BEG[1] ,
    \Tile_X5Y11_S1BEG[0] }),
    .S1END({\Tile_X5Y10_S1BEG[3] ,
    \Tile_X5Y10_S1BEG[2] ,
    \Tile_X5Y10_S1BEG[1] ,
    \Tile_X5Y10_S1BEG[0] }),
    .S2BEG({\Tile_X5Y11_S2BEG[7] ,
    \Tile_X5Y11_S2BEG[6] ,
    \Tile_X5Y11_S2BEG[5] ,
    \Tile_X5Y11_S2BEG[4] ,
    \Tile_X5Y11_S2BEG[3] ,
    \Tile_X5Y11_S2BEG[2] ,
    \Tile_X5Y11_S2BEG[1] ,
    \Tile_X5Y11_S2BEG[0] }),
    .S2BEGb({\Tile_X5Y11_S2BEGb[7] ,
    \Tile_X5Y11_S2BEGb[6] ,
    \Tile_X5Y11_S2BEGb[5] ,
    \Tile_X5Y11_S2BEGb[4] ,
    \Tile_X5Y11_S2BEGb[3] ,
    \Tile_X5Y11_S2BEGb[2] ,
    \Tile_X5Y11_S2BEGb[1] ,
    \Tile_X5Y11_S2BEGb[0] }),
    .S2END({\Tile_X5Y10_S2BEGb[7] ,
    \Tile_X5Y10_S2BEGb[6] ,
    \Tile_X5Y10_S2BEGb[5] ,
    \Tile_X5Y10_S2BEGb[4] ,
    \Tile_X5Y10_S2BEGb[3] ,
    \Tile_X5Y10_S2BEGb[2] ,
    \Tile_X5Y10_S2BEGb[1] ,
    \Tile_X5Y10_S2BEGb[0] }),
    .S2MID({\Tile_X5Y10_S2BEG[7] ,
    \Tile_X5Y10_S2BEG[6] ,
    \Tile_X5Y10_S2BEG[5] ,
    \Tile_X5Y10_S2BEG[4] ,
    \Tile_X5Y10_S2BEG[3] ,
    \Tile_X5Y10_S2BEG[2] ,
    \Tile_X5Y10_S2BEG[1] ,
    \Tile_X5Y10_S2BEG[0] }),
    .S4BEG({\Tile_X5Y11_S4BEG[15] ,
    \Tile_X5Y11_S4BEG[14] ,
    \Tile_X5Y11_S4BEG[13] ,
    \Tile_X5Y11_S4BEG[12] ,
    \Tile_X5Y11_S4BEG[11] ,
    \Tile_X5Y11_S4BEG[10] ,
    \Tile_X5Y11_S4BEG[9] ,
    \Tile_X5Y11_S4BEG[8] ,
    \Tile_X5Y11_S4BEG[7] ,
    \Tile_X5Y11_S4BEG[6] ,
    \Tile_X5Y11_S4BEG[5] ,
    \Tile_X5Y11_S4BEG[4] ,
    \Tile_X5Y11_S4BEG[3] ,
    \Tile_X5Y11_S4BEG[2] ,
    \Tile_X5Y11_S4BEG[1] ,
    \Tile_X5Y11_S4BEG[0] }),
    .S4END({\Tile_X5Y10_S4BEG[15] ,
    \Tile_X5Y10_S4BEG[14] ,
    \Tile_X5Y10_S4BEG[13] ,
    \Tile_X5Y10_S4BEG[12] ,
    \Tile_X5Y10_S4BEG[11] ,
    \Tile_X5Y10_S4BEG[10] ,
    \Tile_X5Y10_S4BEG[9] ,
    \Tile_X5Y10_S4BEG[8] ,
    \Tile_X5Y10_S4BEG[7] ,
    \Tile_X5Y10_S4BEG[6] ,
    \Tile_X5Y10_S4BEG[5] ,
    \Tile_X5Y10_S4BEG[4] ,
    \Tile_X5Y10_S4BEG[3] ,
    \Tile_X5Y10_S4BEG[2] ,
    \Tile_X5Y10_S4BEG[1] ,
    \Tile_X5Y10_S4BEG[0] }),
    .SS4BEG({\Tile_X5Y11_SS4BEG[15] ,
    \Tile_X5Y11_SS4BEG[14] ,
    \Tile_X5Y11_SS4BEG[13] ,
    \Tile_X5Y11_SS4BEG[12] ,
    \Tile_X5Y11_SS4BEG[11] ,
    \Tile_X5Y11_SS4BEG[10] ,
    \Tile_X5Y11_SS4BEG[9] ,
    \Tile_X5Y11_SS4BEG[8] ,
    \Tile_X5Y11_SS4BEG[7] ,
    \Tile_X5Y11_SS4BEG[6] ,
    \Tile_X5Y11_SS4BEG[5] ,
    \Tile_X5Y11_SS4BEG[4] ,
    \Tile_X5Y11_SS4BEG[3] ,
    \Tile_X5Y11_SS4BEG[2] ,
    \Tile_X5Y11_SS4BEG[1] ,
    \Tile_X5Y11_SS4BEG[0] }),
    .SS4END({\Tile_X5Y10_SS4BEG[15] ,
    \Tile_X5Y10_SS4BEG[14] ,
    \Tile_X5Y10_SS4BEG[13] ,
    \Tile_X5Y10_SS4BEG[12] ,
    \Tile_X5Y10_SS4BEG[11] ,
    \Tile_X5Y10_SS4BEG[10] ,
    \Tile_X5Y10_SS4BEG[9] ,
    \Tile_X5Y10_SS4BEG[8] ,
    \Tile_X5Y10_SS4BEG[7] ,
    \Tile_X5Y10_SS4BEG[6] ,
    \Tile_X5Y10_SS4BEG[5] ,
    \Tile_X5Y10_SS4BEG[4] ,
    \Tile_X5Y10_SS4BEG[3] ,
    \Tile_X5Y10_SS4BEG[2] ,
    \Tile_X5Y10_SS4BEG[1] ,
    \Tile_X5Y10_SS4BEG[0] }),
    .W1BEG({\Tile_X5Y11_W1BEG[3] ,
    \Tile_X5Y11_W1BEG[2] ,
    \Tile_X5Y11_W1BEG[1] ,
    \Tile_X5Y11_W1BEG[0] }),
    .W1END({\Tile_X6Y11_W1BEG[3] ,
    \Tile_X6Y11_W1BEG[2] ,
    \Tile_X6Y11_W1BEG[1] ,
    \Tile_X6Y11_W1BEG[0] }),
    .W2BEG({\Tile_X5Y11_W2BEG[7] ,
    \Tile_X5Y11_W2BEG[6] ,
    \Tile_X5Y11_W2BEG[5] ,
    \Tile_X5Y11_W2BEG[4] ,
    \Tile_X5Y11_W2BEG[3] ,
    \Tile_X5Y11_W2BEG[2] ,
    \Tile_X5Y11_W2BEG[1] ,
    \Tile_X5Y11_W2BEG[0] }),
    .W2BEGb({\Tile_X5Y11_W2BEGb[7] ,
    \Tile_X5Y11_W2BEGb[6] ,
    \Tile_X5Y11_W2BEGb[5] ,
    \Tile_X5Y11_W2BEGb[4] ,
    \Tile_X5Y11_W2BEGb[3] ,
    \Tile_X5Y11_W2BEGb[2] ,
    \Tile_X5Y11_W2BEGb[1] ,
    \Tile_X5Y11_W2BEGb[0] }),
    .W2END({\Tile_X6Y11_W2BEGb[7] ,
    \Tile_X6Y11_W2BEGb[6] ,
    \Tile_X6Y11_W2BEGb[5] ,
    \Tile_X6Y11_W2BEGb[4] ,
    \Tile_X6Y11_W2BEGb[3] ,
    \Tile_X6Y11_W2BEGb[2] ,
    \Tile_X6Y11_W2BEGb[1] ,
    \Tile_X6Y11_W2BEGb[0] }),
    .W2MID({\Tile_X6Y11_W2BEG[7] ,
    \Tile_X6Y11_W2BEG[6] ,
    \Tile_X6Y11_W2BEG[5] ,
    \Tile_X6Y11_W2BEG[4] ,
    \Tile_X6Y11_W2BEG[3] ,
    \Tile_X6Y11_W2BEG[2] ,
    \Tile_X6Y11_W2BEG[1] ,
    \Tile_X6Y11_W2BEG[0] }),
    .W6BEG({\Tile_X5Y11_W6BEG[11] ,
    \Tile_X5Y11_W6BEG[10] ,
    \Tile_X5Y11_W6BEG[9] ,
    \Tile_X5Y11_W6BEG[8] ,
    \Tile_X5Y11_W6BEG[7] ,
    \Tile_X5Y11_W6BEG[6] ,
    \Tile_X5Y11_W6BEG[5] ,
    \Tile_X5Y11_W6BEG[4] ,
    \Tile_X5Y11_W6BEG[3] ,
    \Tile_X5Y11_W6BEG[2] ,
    \Tile_X5Y11_W6BEG[1] ,
    \Tile_X5Y11_W6BEG[0] }),
    .W6END({\Tile_X6Y11_W6BEG[11] ,
    \Tile_X6Y11_W6BEG[10] ,
    \Tile_X6Y11_W6BEG[9] ,
    \Tile_X6Y11_W6BEG[8] ,
    \Tile_X6Y11_W6BEG[7] ,
    \Tile_X6Y11_W6BEG[6] ,
    \Tile_X6Y11_W6BEG[5] ,
    \Tile_X6Y11_W6BEG[4] ,
    \Tile_X6Y11_W6BEG[3] ,
    \Tile_X6Y11_W6BEG[2] ,
    \Tile_X6Y11_W6BEG[1] ,
    \Tile_X6Y11_W6BEG[0] }),
    .WW4BEG({\Tile_X5Y11_WW4BEG[15] ,
    \Tile_X5Y11_WW4BEG[14] ,
    \Tile_X5Y11_WW4BEG[13] ,
    \Tile_X5Y11_WW4BEG[12] ,
    \Tile_X5Y11_WW4BEG[11] ,
    \Tile_X5Y11_WW4BEG[10] ,
    \Tile_X5Y11_WW4BEG[9] ,
    \Tile_X5Y11_WW4BEG[8] ,
    \Tile_X5Y11_WW4BEG[7] ,
    \Tile_X5Y11_WW4BEG[6] ,
    \Tile_X5Y11_WW4BEG[5] ,
    \Tile_X5Y11_WW4BEG[4] ,
    \Tile_X5Y11_WW4BEG[3] ,
    \Tile_X5Y11_WW4BEG[2] ,
    \Tile_X5Y11_WW4BEG[1] ,
    \Tile_X5Y11_WW4BEG[0] }),
    .WW4END({\Tile_X6Y11_WW4BEG[15] ,
    \Tile_X6Y11_WW4BEG[14] ,
    \Tile_X6Y11_WW4BEG[13] ,
    \Tile_X6Y11_WW4BEG[12] ,
    \Tile_X6Y11_WW4BEG[11] ,
    \Tile_X6Y11_WW4BEG[10] ,
    \Tile_X6Y11_WW4BEG[9] ,
    \Tile_X6Y11_WW4BEG[8] ,
    \Tile_X6Y11_WW4BEG[7] ,
    \Tile_X6Y11_WW4BEG[6] ,
    \Tile_X6Y11_WW4BEG[5] ,
    \Tile_X6Y11_WW4BEG[4] ,
    \Tile_X6Y11_WW4BEG[3] ,
    \Tile_X6Y11_WW4BEG[2] ,
    \Tile_X6Y11_WW4BEG[1] ,
    \Tile_X6Y11_WW4BEG[0] }));
 LUT4AB Tile_X5Y12_LUT4AB (.Ci(Tile_X5Y13_Co),
    .Co(Tile_X5Y12_Co),
    .UserCLK(Tile_X5Y13_UserCLKo),
    .UserCLKo(Tile_X5Y12_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X5Y12_E1BEG[3] ,
    \Tile_X5Y12_E1BEG[2] ,
    \Tile_X5Y12_E1BEG[1] ,
    \Tile_X5Y12_E1BEG[0] }),
    .E1END({\Tile_X4Y12_E1BEG[3] ,
    \Tile_X4Y12_E1BEG[2] ,
    \Tile_X4Y12_E1BEG[1] ,
    \Tile_X4Y12_E1BEG[0] }),
    .E2BEG({\Tile_X5Y12_E2BEG[7] ,
    \Tile_X5Y12_E2BEG[6] ,
    \Tile_X5Y12_E2BEG[5] ,
    \Tile_X5Y12_E2BEG[4] ,
    \Tile_X5Y12_E2BEG[3] ,
    \Tile_X5Y12_E2BEG[2] ,
    \Tile_X5Y12_E2BEG[1] ,
    \Tile_X5Y12_E2BEG[0] }),
    .E2BEGb({\Tile_X5Y12_E2BEGb[7] ,
    \Tile_X5Y12_E2BEGb[6] ,
    \Tile_X5Y12_E2BEGb[5] ,
    \Tile_X5Y12_E2BEGb[4] ,
    \Tile_X5Y12_E2BEGb[3] ,
    \Tile_X5Y12_E2BEGb[2] ,
    \Tile_X5Y12_E2BEGb[1] ,
    \Tile_X5Y12_E2BEGb[0] }),
    .E2END({\Tile_X4Y12_E2BEGb[7] ,
    \Tile_X4Y12_E2BEGb[6] ,
    \Tile_X4Y12_E2BEGb[5] ,
    \Tile_X4Y12_E2BEGb[4] ,
    \Tile_X4Y12_E2BEGb[3] ,
    \Tile_X4Y12_E2BEGb[2] ,
    \Tile_X4Y12_E2BEGb[1] ,
    \Tile_X4Y12_E2BEGb[0] }),
    .E2MID({\Tile_X4Y12_E2BEG[7] ,
    \Tile_X4Y12_E2BEG[6] ,
    \Tile_X4Y12_E2BEG[5] ,
    \Tile_X4Y12_E2BEG[4] ,
    \Tile_X4Y12_E2BEG[3] ,
    \Tile_X4Y12_E2BEG[2] ,
    \Tile_X4Y12_E2BEG[1] ,
    \Tile_X4Y12_E2BEG[0] }),
    .E6BEG({\Tile_X5Y12_E6BEG[11] ,
    \Tile_X5Y12_E6BEG[10] ,
    \Tile_X5Y12_E6BEG[9] ,
    \Tile_X5Y12_E6BEG[8] ,
    \Tile_X5Y12_E6BEG[7] ,
    \Tile_X5Y12_E6BEG[6] ,
    \Tile_X5Y12_E6BEG[5] ,
    \Tile_X5Y12_E6BEG[4] ,
    \Tile_X5Y12_E6BEG[3] ,
    \Tile_X5Y12_E6BEG[2] ,
    \Tile_X5Y12_E6BEG[1] ,
    \Tile_X5Y12_E6BEG[0] }),
    .E6END({\Tile_X4Y12_E6BEG[11] ,
    \Tile_X4Y12_E6BEG[10] ,
    \Tile_X4Y12_E6BEG[9] ,
    \Tile_X4Y12_E6BEG[8] ,
    \Tile_X4Y12_E6BEG[7] ,
    \Tile_X4Y12_E6BEG[6] ,
    \Tile_X4Y12_E6BEG[5] ,
    \Tile_X4Y12_E6BEG[4] ,
    \Tile_X4Y12_E6BEG[3] ,
    \Tile_X4Y12_E6BEG[2] ,
    \Tile_X4Y12_E6BEG[1] ,
    \Tile_X4Y12_E6BEG[0] }),
    .EE4BEG({\Tile_X5Y12_EE4BEG[15] ,
    \Tile_X5Y12_EE4BEG[14] ,
    \Tile_X5Y12_EE4BEG[13] ,
    \Tile_X5Y12_EE4BEG[12] ,
    \Tile_X5Y12_EE4BEG[11] ,
    \Tile_X5Y12_EE4BEG[10] ,
    \Tile_X5Y12_EE4BEG[9] ,
    \Tile_X5Y12_EE4BEG[8] ,
    \Tile_X5Y12_EE4BEG[7] ,
    \Tile_X5Y12_EE4BEG[6] ,
    \Tile_X5Y12_EE4BEG[5] ,
    \Tile_X5Y12_EE4BEG[4] ,
    \Tile_X5Y12_EE4BEG[3] ,
    \Tile_X5Y12_EE4BEG[2] ,
    \Tile_X5Y12_EE4BEG[1] ,
    \Tile_X5Y12_EE4BEG[0] }),
    .EE4END({\Tile_X4Y12_EE4BEG[15] ,
    \Tile_X4Y12_EE4BEG[14] ,
    \Tile_X4Y12_EE4BEG[13] ,
    \Tile_X4Y12_EE4BEG[12] ,
    \Tile_X4Y12_EE4BEG[11] ,
    \Tile_X4Y12_EE4BEG[10] ,
    \Tile_X4Y12_EE4BEG[9] ,
    \Tile_X4Y12_EE4BEG[8] ,
    \Tile_X4Y12_EE4BEG[7] ,
    \Tile_X4Y12_EE4BEG[6] ,
    \Tile_X4Y12_EE4BEG[5] ,
    \Tile_X4Y12_EE4BEG[4] ,
    \Tile_X4Y12_EE4BEG[3] ,
    \Tile_X4Y12_EE4BEG[2] ,
    \Tile_X4Y12_EE4BEG[1] ,
    \Tile_X4Y12_EE4BEG[0] }),
    .FrameData({\Tile_X4Y12_FrameData_O[31] ,
    \Tile_X4Y12_FrameData_O[30] ,
    \Tile_X4Y12_FrameData_O[29] ,
    \Tile_X4Y12_FrameData_O[28] ,
    \Tile_X4Y12_FrameData_O[27] ,
    \Tile_X4Y12_FrameData_O[26] ,
    \Tile_X4Y12_FrameData_O[25] ,
    \Tile_X4Y12_FrameData_O[24] ,
    \Tile_X4Y12_FrameData_O[23] ,
    \Tile_X4Y12_FrameData_O[22] ,
    \Tile_X4Y12_FrameData_O[21] ,
    \Tile_X4Y12_FrameData_O[20] ,
    \Tile_X4Y12_FrameData_O[19] ,
    \Tile_X4Y12_FrameData_O[18] ,
    \Tile_X4Y12_FrameData_O[17] ,
    \Tile_X4Y12_FrameData_O[16] ,
    \Tile_X4Y12_FrameData_O[15] ,
    \Tile_X4Y12_FrameData_O[14] ,
    \Tile_X4Y12_FrameData_O[13] ,
    \Tile_X4Y12_FrameData_O[12] ,
    \Tile_X4Y12_FrameData_O[11] ,
    \Tile_X4Y12_FrameData_O[10] ,
    \Tile_X4Y12_FrameData_O[9] ,
    \Tile_X4Y12_FrameData_O[8] ,
    \Tile_X4Y12_FrameData_O[7] ,
    \Tile_X4Y12_FrameData_O[6] ,
    \Tile_X4Y12_FrameData_O[5] ,
    \Tile_X4Y12_FrameData_O[4] ,
    \Tile_X4Y12_FrameData_O[3] ,
    \Tile_X4Y12_FrameData_O[2] ,
    \Tile_X4Y12_FrameData_O[1] ,
    \Tile_X4Y12_FrameData_O[0] }),
    .FrameData_O({\Tile_X5Y12_FrameData_O[31] ,
    \Tile_X5Y12_FrameData_O[30] ,
    \Tile_X5Y12_FrameData_O[29] ,
    \Tile_X5Y12_FrameData_O[28] ,
    \Tile_X5Y12_FrameData_O[27] ,
    \Tile_X5Y12_FrameData_O[26] ,
    \Tile_X5Y12_FrameData_O[25] ,
    \Tile_X5Y12_FrameData_O[24] ,
    \Tile_X5Y12_FrameData_O[23] ,
    \Tile_X5Y12_FrameData_O[22] ,
    \Tile_X5Y12_FrameData_O[21] ,
    \Tile_X5Y12_FrameData_O[20] ,
    \Tile_X5Y12_FrameData_O[19] ,
    \Tile_X5Y12_FrameData_O[18] ,
    \Tile_X5Y12_FrameData_O[17] ,
    \Tile_X5Y12_FrameData_O[16] ,
    \Tile_X5Y12_FrameData_O[15] ,
    \Tile_X5Y12_FrameData_O[14] ,
    \Tile_X5Y12_FrameData_O[13] ,
    \Tile_X5Y12_FrameData_O[12] ,
    \Tile_X5Y12_FrameData_O[11] ,
    \Tile_X5Y12_FrameData_O[10] ,
    \Tile_X5Y12_FrameData_O[9] ,
    \Tile_X5Y12_FrameData_O[8] ,
    \Tile_X5Y12_FrameData_O[7] ,
    \Tile_X5Y12_FrameData_O[6] ,
    \Tile_X5Y12_FrameData_O[5] ,
    \Tile_X5Y12_FrameData_O[4] ,
    \Tile_X5Y12_FrameData_O[3] ,
    \Tile_X5Y12_FrameData_O[2] ,
    \Tile_X5Y12_FrameData_O[1] ,
    \Tile_X5Y12_FrameData_O[0] }),
    .FrameStrobe({\Tile_X5Y13_FrameStrobe_O[19] ,
    \Tile_X5Y13_FrameStrobe_O[18] ,
    \Tile_X5Y13_FrameStrobe_O[17] ,
    \Tile_X5Y13_FrameStrobe_O[16] ,
    \Tile_X5Y13_FrameStrobe_O[15] ,
    \Tile_X5Y13_FrameStrobe_O[14] ,
    \Tile_X5Y13_FrameStrobe_O[13] ,
    \Tile_X5Y13_FrameStrobe_O[12] ,
    \Tile_X5Y13_FrameStrobe_O[11] ,
    \Tile_X5Y13_FrameStrobe_O[10] ,
    \Tile_X5Y13_FrameStrobe_O[9] ,
    \Tile_X5Y13_FrameStrobe_O[8] ,
    \Tile_X5Y13_FrameStrobe_O[7] ,
    \Tile_X5Y13_FrameStrobe_O[6] ,
    \Tile_X5Y13_FrameStrobe_O[5] ,
    \Tile_X5Y13_FrameStrobe_O[4] ,
    \Tile_X5Y13_FrameStrobe_O[3] ,
    \Tile_X5Y13_FrameStrobe_O[2] ,
    \Tile_X5Y13_FrameStrobe_O[1] ,
    \Tile_X5Y13_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X5Y12_FrameStrobe_O[19] ,
    \Tile_X5Y12_FrameStrobe_O[18] ,
    \Tile_X5Y12_FrameStrobe_O[17] ,
    \Tile_X5Y12_FrameStrobe_O[16] ,
    \Tile_X5Y12_FrameStrobe_O[15] ,
    \Tile_X5Y12_FrameStrobe_O[14] ,
    \Tile_X5Y12_FrameStrobe_O[13] ,
    \Tile_X5Y12_FrameStrobe_O[12] ,
    \Tile_X5Y12_FrameStrobe_O[11] ,
    \Tile_X5Y12_FrameStrobe_O[10] ,
    \Tile_X5Y12_FrameStrobe_O[9] ,
    \Tile_X5Y12_FrameStrobe_O[8] ,
    \Tile_X5Y12_FrameStrobe_O[7] ,
    \Tile_X5Y12_FrameStrobe_O[6] ,
    \Tile_X5Y12_FrameStrobe_O[5] ,
    \Tile_X5Y12_FrameStrobe_O[4] ,
    \Tile_X5Y12_FrameStrobe_O[3] ,
    \Tile_X5Y12_FrameStrobe_O[2] ,
    \Tile_X5Y12_FrameStrobe_O[1] ,
    \Tile_X5Y12_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X5Y12_N1BEG[3] ,
    \Tile_X5Y12_N1BEG[2] ,
    \Tile_X5Y12_N1BEG[1] ,
    \Tile_X5Y12_N1BEG[0] }),
    .N1END({\Tile_X5Y13_N1BEG[3] ,
    \Tile_X5Y13_N1BEG[2] ,
    \Tile_X5Y13_N1BEG[1] ,
    \Tile_X5Y13_N1BEG[0] }),
    .N2BEG({\Tile_X5Y12_N2BEG[7] ,
    \Tile_X5Y12_N2BEG[6] ,
    \Tile_X5Y12_N2BEG[5] ,
    \Tile_X5Y12_N2BEG[4] ,
    \Tile_X5Y12_N2BEG[3] ,
    \Tile_X5Y12_N2BEG[2] ,
    \Tile_X5Y12_N2BEG[1] ,
    \Tile_X5Y12_N2BEG[0] }),
    .N2BEGb({\Tile_X5Y12_N2BEGb[7] ,
    \Tile_X5Y12_N2BEGb[6] ,
    \Tile_X5Y12_N2BEGb[5] ,
    \Tile_X5Y12_N2BEGb[4] ,
    \Tile_X5Y12_N2BEGb[3] ,
    \Tile_X5Y12_N2BEGb[2] ,
    \Tile_X5Y12_N2BEGb[1] ,
    \Tile_X5Y12_N2BEGb[0] }),
    .N2END({\Tile_X5Y13_N2BEGb[7] ,
    \Tile_X5Y13_N2BEGb[6] ,
    \Tile_X5Y13_N2BEGb[5] ,
    \Tile_X5Y13_N2BEGb[4] ,
    \Tile_X5Y13_N2BEGb[3] ,
    \Tile_X5Y13_N2BEGb[2] ,
    \Tile_X5Y13_N2BEGb[1] ,
    \Tile_X5Y13_N2BEGb[0] }),
    .N2MID({\Tile_X5Y13_N2BEG[7] ,
    \Tile_X5Y13_N2BEG[6] ,
    \Tile_X5Y13_N2BEG[5] ,
    \Tile_X5Y13_N2BEG[4] ,
    \Tile_X5Y13_N2BEG[3] ,
    \Tile_X5Y13_N2BEG[2] ,
    \Tile_X5Y13_N2BEG[1] ,
    \Tile_X5Y13_N2BEG[0] }),
    .N4BEG({\Tile_X5Y12_N4BEG[15] ,
    \Tile_X5Y12_N4BEG[14] ,
    \Tile_X5Y12_N4BEG[13] ,
    \Tile_X5Y12_N4BEG[12] ,
    \Tile_X5Y12_N4BEG[11] ,
    \Tile_X5Y12_N4BEG[10] ,
    \Tile_X5Y12_N4BEG[9] ,
    \Tile_X5Y12_N4BEG[8] ,
    \Tile_X5Y12_N4BEG[7] ,
    \Tile_X5Y12_N4BEG[6] ,
    \Tile_X5Y12_N4BEG[5] ,
    \Tile_X5Y12_N4BEG[4] ,
    \Tile_X5Y12_N4BEG[3] ,
    \Tile_X5Y12_N4BEG[2] ,
    \Tile_X5Y12_N4BEG[1] ,
    \Tile_X5Y12_N4BEG[0] }),
    .N4END({\Tile_X5Y13_N4BEG[15] ,
    \Tile_X5Y13_N4BEG[14] ,
    \Tile_X5Y13_N4BEG[13] ,
    \Tile_X5Y13_N4BEG[12] ,
    \Tile_X5Y13_N4BEG[11] ,
    \Tile_X5Y13_N4BEG[10] ,
    \Tile_X5Y13_N4BEG[9] ,
    \Tile_X5Y13_N4BEG[8] ,
    \Tile_X5Y13_N4BEG[7] ,
    \Tile_X5Y13_N4BEG[6] ,
    \Tile_X5Y13_N4BEG[5] ,
    \Tile_X5Y13_N4BEG[4] ,
    \Tile_X5Y13_N4BEG[3] ,
    \Tile_X5Y13_N4BEG[2] ,
    \Tile_X5Y13_N4BEG[1] ,
    \Tile_X5Y13_N4BEG[0] }),
    .NN4BEG({\Tile_X5Y12_NN4BEG[15] ,
    \Tile_X5Y12_NN4BEG[14] ,
    \Tile_X5Y12_NN4BEG[13] ,
    \Tile_X5Y12_NN4BEG[12] ,
    \Tile_X5Y12_NN4BEG[11] ,
    \Tile_X5Y12_NN4BEG[10] ,
    \Tile_X5Y12_NN4BEG[9] ,
    \Tile_X5Y12_NN4BEG[8] ,
    \Tile_X5Y12_NN4BEG[7] ,
    \Tile_X5Y12_NN4BEG[6] ,
    \Tile_X5Y12_NN4BEG[5] ,
    \Tile_X5Y12_NN4BEG[4] ,
    \Tile_X5Y12_NN4BEG[3] ,
    \Tile_X5Y12_NN4BEG[2] ,
    \Tile_X5Y12_NN4BEG[1] ,
    \Tile_X5Y12_NN4BEG[0] }),
    .NN4END({\Tile_X5Y13_NN4BEG[15] ,
    \Tile_X5Y13_NN4BEG[14] ,
    \Tile_X5Y13_NN4BEG[13] ,
    \Tile_X5Y13_NN4BEG[12] ,
    \Tile_X5Y13_NN4BEG[11] ,
    \Tile_X5Y13_NN4BEG[10] ,
    \Tile_X5Y13_NN4BEG[9] ,
    \Tile_X5Y13_NN4BEG[8] ,
    \Tile_X5Y13_NN4BEG[7] ,
    \Tile_X5Y13_NN4BEG[6] ,
    \Tile_X5Y13_NN4BEG[5] ,
    \Tile_X5Y13_NN4BEG[4] ,
    \Tile_X5Y13_NN4BEG[3] ,
    \Tile_X5Y13_NN4BEG[2] ,
    \Tile_X5Y13_NN4BEG[1] ,
    \Tile_X5Y13_NN4BEG[0] }),
    .S1BEG({\Tile_X5Y12_S1BEG[3] ,
    \Tile_X5Y12_S1BEG[2] ,
    \Tile_X5Y12_S1BEG[1] ,
    \Tile_X5Y12_S1BEG[0] }),
    .S1END({\Tile_X5Y11_S1BEG[3] ,
    \Tile_X5Y11_S1BEG[2] ,
    \Tile_X5Y11_S1BEG[1] ,
    \Tile_X5Y11_S1BEG[0] }),
    .S2BEG({\Tile_X5Y12_S2BEG[7] ,
    \Tile_X5Y12_S2BEG[6] ,
    \Tile_X5Y12_S2BEG[5] ,
    \Tile_X5Y12_S2BEG[4] ,
    \Tile_X5Y12_S2BEG[3] ,
    \Tile_X5Y12_S2BEG[2] ,
    \Tile_X5Y12_S2BEG[1] ,
    \Tile_X5Y12_S2BEG[0] }),
    .S2BEGb({\Tile_X5Y12_S2BEGb[7] ,
    \Tile_X5Y12_S2BEGb[6] ,
    \Tile_X5Y12_S2BEGb[5] ,
    \Tile_X5Y12_S2BEGb[4] ,
    \Tile_X5Y12_S2BEGb[3] ,
    \Tile_X5Y12_S2BEGb[2] ,
    \Tile_X5Y12_S2BEGb[1] ,
    \Tile_X5Y12_S2BEGb[0] }),
    .S2END({\Tile_X5Y11_S2BEGb[7] ,
    \Tile_X5Y11_S2BEGb[6] ,
    \Tile_X5Y11_S2BEGb[5] ,
    \Tile_X5Y11_S2BEGb[4] ,
    \Tile_X5Y11_S2BEGb[3] ,
    \Tile_X5Y11_S2BEGb[2] ,
    \Tile_X5Y11_S2BEGb[1] ,
    \Tile_X5Y11_S2BEGb[0] }),
    .S2MID({\Tile_X5Y11_S2BEG[7] ,
    \Tile_X5Y11_S2BEG[6] ,
    \Tile_X5Y11_S2BEG[5] ,
    \Tile_X5Y11_S2BEG[4] ,
    \Tile_X5Y11_S2BEG[3] ,
    \Tile_X5Y11_S2BEG[2] ,
    \Tile_X5Y11_S2BEG[1] ,
    \Tile_X5Y11_S2BEG[0] }),
    .S4BEG({\Tile_X5Y12_S4BEG[15] ,
    \Tile_X5Y12_S4BEG[14] ,
    \Tile_X5Y12_S4BEG[13] ,
    \Tile_X5Y12_S4BEG[12] ,
    \Tile_X5Y12_S4BEG[11] ,
    \Tile_X5Y12_S4BEG[10] ,
    \Tile_X5Y12_S4BEG[9] ,
    \Tile_X5Y12_S4BEG[8] ,
    \Tile_X5Y12_S4BEG[7] ,
    \Tile_X5Y12_S4BEG[6] ,
    \Tile_X5Y12_S4BEG[5] ,
    \Tile_X5Y12_S4BEG[4] ,
    \Tile_X5Y12_S4BEG[3] ,
    \Tile_X5Y12_S4BEG[2] ,
    \Tile_X5Y12_S4BEG[1] ,
    \Tile_X5Y12_S4BEG[0] }),
    .S4END({\Tile_X5Y11_S4BEG[15] ,
    \Tile_X5Y11_S4BEG[14] ,
    \Tile_X5Y11_S4BEG[13] ,
    \Tile_X5Y11_S4BEG[12] ,
    \Tile_X5Y11_S4BEG[11] ,
    \Tile_X5Y11_S4BEG[10] ,
    \Tile_X5Y11_S4BEG[9] ,
    \Tile_X5Y11_S4BEG[8] ,
    \Tile_X5Y11_S4BEG[7] ,
    \Tile_X5Y11_S4BEG[6] ,
    \Tile_X5Y11_S4BEG[5] ,
    \Tile_X5Y11_S4BEG[4] ,
    \Tile_X5Y11_S4BEG[3] ,
    \Tile_X5Y11_S4BEG[2] ,
    \Tile_X5Y11_S4BEG[1] ,
    \Tile_X5Y11_S4BEG[0] }),
    .SS4BEG({\Tile_X5Y12_SS4BEG[15] ,
    \Tile_X5Y12_SS4BEG[14] ,
    \Tile_X5Y12_SS4BEG[13] ,
    \Tile_X5Y12_SS4BEG[12] ,
    \Tile_X5Y12_SS4BEG[11] ,
    \Tile_X5Y12_SS4BEG[10] ,
    \Tile_X5Y12_SS4BEG[9] ,
    \Tile_X5Y12_SS4BEG[8] ,
    \Tile_X5Y12_SS4BEG[7] ,
    \Tile_X5Y12_SS4BEG[6] ,
    \Tile_X5Y12_SS4BEG[5] ,
    \Tile_X5Y12_SS4BEG[4] ,
    \Tile_X5Y12_SS4BEG[3] ,
    \Tile_X5Y12_SS4BEG[2] ,
    \Tile_X5Y12_SS4BEG[1] ,
    \Tile_X5Y12_SS4BEG[0] }),
    .SS4END({\Tile_X5Y11_SS4BEG[15] ,
    \Tile_X5Y11_SS4BEG[14] ,
    \Tile_X5Y11_SS4BEG[13] ,
    \Tile_X5Y11_SS4BEG[12] ,
    \Tile_X5Y11_SS4BEG[11] ,
    \Tile_X5Y11_SS4BEG[10] ,
    \Tile_X5Y11_SS4BEG[9] ,
    \Tile_X5Y11_SS4BEG[8] ,
    \Tile_X5Y11_SS4BEG[7] ,
    \Tile_X5Y11_SS4BEG[6] ,
    \Tile_X5Y11_SS4BEG[5] ,
    \Tile_X5Y11_SS4BEG[4] ,
    \Tile_X5Y11_SS4BEG[3] ,
    \Tile_X5Y11_SS4BEG[2] ,
    \Tile_X5Y11_SS4BEG[1] ,
    \Tile_X5Y11_SS4BEG[0] }),
    .W1BEG({\Tile_X5Y12_W1BEG[3] ,
    \Tile_X5Y12_W1BEG[2] ,
    \Tile_X5Y12_W1BEG[1] ,
    \Tile_X5Y12_W1BEG[0] }),
    .W1END({\Tile_X6Y12_W1BEG[3] ,
    \Tile_X6Y12_W1BEG[2] ,
    \Tile_X6Y12_W1BEG[1] ,
    \Tile_X6Y12_W1BEG[0] }),
    .W2BEG({\Tile_X5Y12_W2BEG[7] ,
    \Tile_X5Y12_W2BEG[6] ,
    \Tile_X5Y12_W2BEG[5] ,
    \Tile_X5Y12_W2BEG[4] ,
    \Tile_X5Y12_W2BEG[3] ,
    \Tile_X5Y12_W2BEG[2] ,
    \Tile_X5Y12_W2BEG[1] ,
    \Tile_X5Y12_W2BEG[0] }),
    .W2BEGb({\Tile_X5Y12_W2BEGb[7] ,
    \Tile_X5Y12_W2BEGb[6] ,
    \Tile_X5Y12_W2BEGb[5] ,
    \Tile_X5Y12_W2BEGb[4] ,
    \Tile_X5Y12_W2BEGb[3] ,
    \Tile_X5Y12_W2BEGb[2] ,
    \Tile_X5Y12_W2BEGb[1] ,
    \Tile_X5Y12_W2BEGb[0] }),
    .W2END({\Tile_X6Y12_W2BEGb[7] ,
    \Tile_X6Y12_W2BEGb[6] ,
    \Tile_X6Y12_W2BEGb[5] ,
    \Tile_X6Y12_W2BEGb[4] ,
    \Tile_X6Y12_W2BEGb[3] ,
    \Tile_X6Y12_W2BEGb[2] ,
    \Tile_X6Y12_W2BEGb[1] ,
    \Tile_X6Y12_W2BEGb[0] }),
    .W2MID({\Tile_X6Y12_W2BEG[7] ,
    \Tile_X6Y12_W2BEG[6] ,
    \Tile_X6Y12_W2BEG[5] ,
    \Tile_X6Y12_W2BEG[4] ,
    \Tile_X6Y12_W2BEG[3] ,
    \Tile_X6Y12_W2BEG[2] ,
    \Tile_X6Y12_W2BEG[1] ,
    \Tile_X6Y12_W2BEG[0] }),
    .W6BEG({\Tile_X5Y12_W6BEG[11] ,
    \Tile_X5Y12_W6BEG[10] ,
    \Tile_X5Y12_W6BEG[9] ,
    \Tile_X5Y12_W6BEG[8] ,
    \Tile_X5Y12_W6BEG[7] ,
    \Tile_X5Y12_W6BEG[6] ,
    \Tile_X5Y12_W6BEG[5] ,
    \Tile_X5Y12_W6BEG[4] ,
    \Tile_X5Y12_W6BEG[3] ,
    \Tile_X5Y12_W6BEG[2] ,
    \Tile_X5Y12_W6BEG[1] ,
    \Tile_X5Y12_W6BEG[0] }),
    .W6END({\Tile_X6Y12_W6BEG[11] ,
    \Tile_X6Y12_W6BEG[10] ,
    \Tile_X6Y12_W6BEG[9] ,
    \Tile_X6Y12_W6BEG[8] ,
    \Tile_X6Y12_W6BEG[7] ,
    \Tile_X6Y12_W6BEG[6] ,
    \Tile_X6Y12_W6BEG[5] ,
    \Tile_X6Y12_W6BEG[4] ,
    \Tile_X6Y12_W6BEG[3] ,
    \Tile_X6Y12_W6BEG[2] ,
    \Tile_X6Y12_W6BEG[1] ,
    \Tile_X6Y12_W6BEG[0] }),
    .WW4BEG({\Tile_X5Y12_WW4BEG[15] ,
    \Tile_X5Y12_WW4BEG[14] ,
    \Tile_X5Y12_WW4BEG[13] ,
    \Tile_X5Y12_WW4BEG[12] ,
    \Tile_X5Y12_WW4BEG[11] ,
    \Tile_X5Y12_WW4BEG[10] ,
    \Tile_X5Y12_WW4BEG[9] ,
    \Tile_X5Y12_WW4BEG[8] ,
    \Tile_X5Y12_WW4BEG[7] ,
    \Tile_X5Y12_WW4BEG[6] ,
    \Tile_X5Y12_WW4BEG[5] ,
    \Tile_X5Y12_WW4BEG[4] ,
    \Tile_X5Y12_WW4BEG[3] ,
    \Tile_X5Y12_WW4BEG[2] ,
    \Tile_X5Y12_WW4BEG[1] ,
    \Tile_X5Y12_WW4BEG[0] }),
    .WW4END({\Tile_X6Y12_WW4BEG[15] ,
    \Tile_X6Y12_WW4BEG[14] ,
    \Tile_X6Y12_WW4BEG[13] ,
    \Tile_X6Y12_WW4BEG[12] ,
    \Tile_X6Y12_WW4BEG[11] ,
    \Tile_X6Y12_WW4BEG[10] ,
    \Tile_X6Y12_WW4BEG[9] ,
    \Tile_X6Y12_WW4BEG[8] ,
    \Tile_X6Y12_WW4BEG[7] ,
    \Tile_X6Y12_WW4BEG[6] ,
    \Tile_X6Y12_WW4BEG[5] ,
    \Tile_X6Y12_WW4BEG[4] ,
    \Tile_X6Y12_WW4BEG[3] ,
    \Tile_X6Y12_WW4BEG[2] ,
    \Tile_X6Y12_WW4BEG[1] ,
    \Tile_X6Y12_WW4BEG[0] }));
 LUT4AB Tile_X5Y13_LUT4AB (.Ci(Tile_X5Y14_Co),
    .Co(Tile_X5Y13_Co),
    .UserCLK(Tile_X5Y14_UserCLKo),
    .UserCLKo(Tile_X5Y13_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X5Y13_E1BEG[3] ,
    \Tile_X5Y13_E1BEG[2] ,
    \Tile_X5Y13_E1BEG[1] ,
    \Tile_X5Y13_E1BEG[0] }),
    .E1END({\Tile_X4Y13_E1BEG[3] ,
    \Tile_X4Y13_E1BEG[2] ,
    \Tile_X4Y13_E1BEG[1] ,
    \Tile_X4Y13_E1BEG[0] }),
    .E2BEG({\Tile_X5Y13_E2BEG[7] ,
    \Tile_X5Y13_E2BEG[6] ,
    \Tile_X5Y13_E2BEG[5] ,
    \Tile_X5Y13_E2BEG[4] ,
    \Tile_X5Y13_E2BEG[3] ,
    \Tile_X5Y13_E2BEG[2] ,
    \Tile_X5Y13_E2BEG[1] ,
    \Tile_X5Y13_E2BEG[0] }),
    .E2BEGb({\Tile_X5Y13_E2BEGb[7] ,
    \Tile_X5Y13_E2BEGb[6] ,
    \Tile_X5Y13_E2BEGb[5] ,
    \Tile_X5Y13_E2BEGb[4] ,
    \Tile_X5Y13_E2BEGb[3] ,
    \Tile_X5Y13_E2BEGb[2] ,
    \Tile_X5Y13_E2BEGb[1] ,
    \Tile_X5Y13_E2BEGb[0] }),
    .E2END({\Tile_X4Y13_E2BEGb[7] ,
    \Tile_X4Y13_E2BEGb[6] ,
    \Tile_X4Y13_E2BEGb[5] ,
    \Tile_X4Y13_E2BEGb[4] ,
    \Tile_X4Y13_E2BEGb[3] ,
    \Tile_X4Y13_E2BEGb[2] ,
    \Tile_X4Y13_E2BEGb[1] ,
    \Tile_X4Y13_E2BEGb[0] }),
    .E2MID({\Tile_X4Y13_E2BEG[7] ,
    \Tile_X4Y13_E2BEG[6] ,
    \Tile_X4Y13_E2BEG[5] ,
    \Tile_X4Y13_E2BEG[4] ,
    \Tile_X4Y13_E2BEG[3] ,
    \Tile_X4Y13_E2BEG[2] ,
    \Tile_X4Y13_E2BEG[1] ,
    \Tile_X4Y13_E2BEG[0] }),
    .E6BEG({\Tile_X5Y13_E6BEG[11] ,
    \Tile_X5Y13_E6BEG[10] ,
    \Tile_X5Y13_E6BEG[9] ,
    \Tile_X5Y13_E6BEG[8] ,
    \Tile_X5Y13_E6BEG[7] ,
    \Tile_X5Y13_E6BEG[6] ,
    \Tile_X5Y13_E6BEG[5] ,
    \Tile_X5Y13_E6BEG[4] ,
    \Tile_X5Y13_E6BEG[3] ,
    \Tile_X5Y13_E6BEG[2] ,
    \Tile_X5Y13_E6BEG[1] ,
    \Tile_X5Y13_E6BEG[0] }),
    .E6END({\Tile_X4Y13_E6BEG[11] ,
    \Tile_X4Y13_E6BEG[10] ,
    \Tile_X4Y13_E6BEG[9] ,
    \Tile_X4Y13_E6BEG[8] ,
    \Tile_X4Y13_E6BEG[7] ,
    \Tile_X4Y13_E6BEG[6] ,
    \Tile_X4Y13_E6BEG[5] ,
    \Tile_X4Y13_E6BEG[4] ,
    \Tile_X4Y13_E6BEG[3] ,
    \Tile_X4Y13_E6BEG[2] ,
    \Tile_X4Y13_E6BEG[1] ,
    \Tile_X4Y13_E6BEG[0] }),
    .EE4BEG({\Tile_X5Y13_EE4BEG[15] ,
    \Tile_X5Y13_EE4BEG[14] ,
    \Tile_X5Y13_EE4BEG[13] ,
    \Tile_X5Y13_EE4BEG[12] ,
    \Tile_X5Y13_EE4BEG[11] ,
    \Tile_X5Y13_EE4BEG[10] ,
    \Tile_X5Y13_EE4BEG[9] ,
    \Tile_X5Y13_EE4BEG[8] ,
    \Tile_X5Y13_EE4BEG[7] ,
    \Tile_X5Y13_EE4BEG[6] ,
    \Tile_X5Y13_EE4BEG[5] ,
    \Tile_X5Y13_EE4BEG[4] ,
    \Tile_X5Y13_EE4BEG[3] ,
    \Tile_X5Y13_EE4BEG[2] ,
    \Tile_X5Y13_EE4BEG[1] ,
    \Tile_X5Y13_EE4BEG[0] }),
    .EE4END({\Tile_X4Y13_EE4BEG[15] ,
    \Tile_X4Y13_EE4BEG[14] ,
    \Tile_X4Y13_EE4BEG[13] ,
    \Tile_X4Y13_EE4BEG[12] ,
    \Tile_X4Y13_EE4BEG[11] ,
    \Tile_X4Y13_EE4BEG[10] ,
    \Tile_X4Y13_EE4BEG[9] ,
    \Tile_X4Y13_EE4BEG[8] ,
    \Tile_X4Y13_EE4BEG[7] ,
    \Tile_X4Y13_EE4BEG[6] ,
    \Tile_X4Y13_EE4BEG[5] ,
    \Tile_X4Y13_EE4BEG[4] ,
    \Tile_X4Y13_EE4BEG[3] ,
    \Tile_X4Y13_EE4BEG[2] ,
    \Tile_X4Y13_EE4BEG[1] ,
    \Tile_X4Y13_EE4BEG[0] }),
    .FrameData({\Tile_X4Y13_FrameData_O[31] ,
    \Tile_X4Y13_FrameData_O[30] ,
    \Tile_X4Y13_FrameData_O[29] ,
    \Tile_X4Y13_FrameData_O[28] ,
    \Tile_X4Y13_FrameData_O[27] ,
    \Tile_X4Y13_FrameData_O[26] ,
    \Tile_X4Y13_FrameData_O[25] ,
    \Tile_X4Y13_FrameData_O[24] ,
    \Tile_X4Y13_FrameData_O[23] ,
    \Tile_X4Y13_FrameData_O[22] ,
    \Tile_X4Y13_FrameData_O[21] ,
    \Tile_X4Y13_FrameData_O[20] ,
    \Tile_X4Y13_FrameData_O[19] ,
    \Tile_X4Y13_FrameData_O[18] ,
    \Tile_X4Y13_FrameData_O[17] ,
    \Tile_X4Y13_FrameData_O[16] ,
    \Tile_X4Y13_FrameData_O[15] ,
    \Tile_X4Y13_FrameData_O[14] ,
    \Tile_X4Y13_FrameData_O[13] ,
    \Tile_X4Y13_FrameData_O[12] ,
    \Tile_X4Y13_FrameData_O[11] ,
    \Tile_X4Y13_FrameData_O[10] ,
    \Tile_X4Y13_FrameData_O[9] ,
    \Tile_X4Y13_FrameData_O[8] ,
    \Tile_X4Y13_FrameData_O[7] ,
    \Tile_X4Y13_FrameData_O[6] ,
    \Tile_X4Y13_FrameData_O[5] ,
    \Tile_X4Y13_FrameData_O[4] ,
    \Tile_X4Y13_FrameData_O[3] ,
    \Tile_X4Y13_FrameData_O[2] ,
    \Tile_X4Y13_FrameData_O[1] ,
    \Tile_X4Y13_FrameData_O[0] }),
    .FrameData_O({\Tile_X5Y13_FrameData_O[31] ,
    \Tile_X5Y13_FrameData_O[30] ,
    \Tile_X5Y13_FrameData_O[29] ,
    \Tile_X5Y13_FrameData_O[28] ,
    \Tile_X5Y13_FrameData_O[27] ,
    \Tile_X5Y13_FrameData_O[26] ,
    \Tile_X5Y13_FrameData_O[25] ,
    \Tile_X5Y13_FrameData_O[24] ,
    \Tile_X5Y13_FrameData_O[23] ,
    \Tile_X5Y13_FrameData_O[22] ,
    \Tile_X5Y13_FrameData_O[21] ,
    \Tile_X5Y13_FrameData_O[20] ,
    \Tile_X5Y13_FrameData_O[19] ,
    \Tile_X5Y13_FrameData_O[18] ,
    \Tile_X5Y13_FrameData_O[17] ,
    \Tile_X5Y13_FrameData_O[16] ,
    \Tile_X5Y13_FrameData_O[15] ,
    \Tile_X5Y13_FrameData_O[14] ,
    \Tile_X5Y13_FrameData_O[13] ,
    \Tile_X5Y13_FrameData_O[12] ,
    \Tile_X5Y13_FrameData_O[11] ,
    \Tile_X5Y13_FrameData_O[10] ,
    \Tile_X5Y13_FrameData_O[9] ,
    \Tile_X5Y13_FrameData_O[8] ,
    \Tile_X5Y13_FrameData_O[7] ,
    \Tile_X5Y13_FrameData_O[6] ,
    \Tile_X5Y13_FrameData_O[5] ,
    \Tile_X5Y13_FrameData_O[4] ,
    \Tile_X5Y13_FrameData_O[3] ,
    \Tile_X5Y13_FrameData_O[2] ,
    \Tile_X5Y13_FrameData_O[1] ,
    \Tile_X5Y13_FrameData_O[0] }),
    .FrameStrobe({\Tile_X5Y14_FrameStrobe_O[19] ,
    \Tile_X5Y14_FrameStrobe_O[18] ,
    \Tile_X5Y14_FrameStrobe_O[17] ,
    \Tile_X5Y14_FrameStrobe_O[16] ,
    \Tile_X5Y14_FrameStrobe_O[15] ,
    \Tile_X5Y14_FrameStrobe_O[14] ,
    \Tile_X5Y14_FrameStrobe_O[13] ,
    \Tile_X5Y14_FrameStrobe_O[12] ,
    \Tile_X5Y14_FrameStrobe_O[11] ,
    \Tile_X5Y14_FrameStrobe_O[10] ,
    \Tile_X5Y14_FrameStrobe_O[9] ,
    \Tile_X5Y14_FrameStrobe_O[8] ,
    \Tile_X5Y14_FrameStrobe_O[7] ,
    \Tile_X5Y14_FrameStrobe_O[6] ,
    \Tile_X5Y14_FrameStrobe_O[5] ,
    \Tile_X5Y14_FrameStrobe_O[4] ,
    \Tile_X5Y14_FrameStrobe_O[3] ,
    \Tile_X5Y14_FrameStrobe_O[2] ,
    \Tile_X5Y14_FrameStrobe_O[1] ,
    \Tile_X5Y14_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X5Y13_FrameStrobe_O[19] ,
    \Tile_X5Y13_FrameStrobe_O[18] ,
    \Tile_X5Y13_FrameStrobe_O[17] ,
    \Tile_X5Y13_FrameStrobe_O[16] ,
    \Tile_X5Y13_FrameStrobe_O[15] ,
    \Tile_X5Y13_FrameStrobe_O[14] ,
    \Tile_X5Y13_FrameStrobe_O[13] ,
    \Tile_X5Y13_FrameStrobe_O[12] ,
    \Tile_X5Y13_FrameStrobe_O[11] ,
    \Tile_X5Y13_FrameStrobe_O[10] ,
    \Tile_X5Y13_FrameStrobe_O[9] ,
    \Tile_X5Y13_FrameStrobe_O[8] ,
    \Tile_X5Y13_FrameStrobe_O[7] ,
    \Tile_X5Y13_FrameStrobe_O[6] ,
    \Tile_X5Y13_FrameStrobe_O[5] ,
    \Tile_X5Y13_FrameStrobe_O[4] ,
    \Tile_X5Y13_FrameStrobe_O[3] ,
    \Tile_X5Y13_FrameStrobe_O[2] ,
    \Tile_X5Y13_FrameStrobe_O[1] ,
    \Tile_X5Y13_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X5Y13_N1BEG[3] ,
    \Tile_X5Y13_N1BEG[2] ,
    \Tile_X5Y13_N1BEG[1] ,
    \Tile_X5Y13_N1BEG[0] }),
    .N1END({\Tile_X5Y14_N1BEG[3] ,
    \Tile_X5Y14_N1BEG[2] ,
    \Tile_X5Y14_N1BEG[1] ,
    \Tile_X5Y14_N1BEG[0] }),
    .N2BEG({\Tile_X5Y13_N2BEG[7] ,
    \Tile_X5Y13_N2BEG[6] ,
    \Tile_X5Y13_N2BEG[5] ,
    \Tile_X5Y13_N2BEG[4] ,
    \Tile_X5Y13_N2BEG[3] ,
    \Tile_X5Y13_N2BEG[2] ,
    \Tile_X5Y13_N2BEG[1] ,
    \Tile_X5Y13_N2BEG[0] }),
    .N2BEGb({\Tile_X5Y13_N2BEGb[7] ,
    \Tile_X5Y13_N2BEGb[6] ,
    \Tile_X5Y13_N2BEGb[5] ,
    \Tile_X5Y13_N2BEGb[4] ,
    \Tile_X5Y13_N2BEGb[3] ,
    \Tile_X5Y13_N2BEGb[2] ,
    \Tile_X5Y13_N2BEGb[1] ,
    \Tile_X5Y13_N2BEGb[0] }),
    .N2END({\Tile_X5Y14_N2BEGb[7] ,
    \Tile_X5Y14_N2BEGb[6] ,
    \Tile_X5Y14_N2BEGb[5] ,
    \Tile_X5Y14_N2BEGb[4] ,
    \Tile_X5Y14_N2BEGb[3] ,
    \Tile_X5Y14_N2BEGb[2] ,
    \Tile_X5Y14_N2BEGb[1] ,
    \Tile_X5Y14_N2BEGb[0] }),
    .N2MID({\Tile_X5Y14_N2BEG[7] ,
    \Tile_X5Y14_N2BEG[6] ,
    \Tile_X5Y14_N2BEG[5] ,
    \Tile_X5Y14_N2BEG[4] ,
    \Tile_X5Y14_N2BEG[3] ,
    \Tile_X5Y14_N2BEG[2] ,
    \Tile_X5Y14_N2BEG[1] ,
    \Tile_X5Y14_N2BEG[0] }),
    .N4BEG({\Tile_X5Y13_N4BEG[15] ,
    \Tile_X5Y13_N4BEG[14] ,
    \Tile_X5Y13_N4BEG[13] ,
    \Tile_X5Y13_N4BEG[12] ,
    \Tile_X5Y13_N4BEG[11] ,
    \Tile_X5Y13_N4BEG[10] ,
    \Tile_X5Y13_N4BEG[9] ,
    \Tile_X5Y13_N4BEG[8] ,
    \Tile_X5Y13_N4BEG[7] ,
    \Tile_X5Y13_N4BEG[6] ,
    \Tile_X5Y13_N4BEG[5] ,
    \Tile_X5Y13_N4BEG[4] ,
    \Tile_X5Y13_N4BEG[3] ,
    \Tile_X5Y13_N4BEG[2] ,
    \Tile_X5Y13_N4BEG[1] ,
    \Tile_X5Y13_N4BEG[0] }),
    .N4END({\Tile_X5Y14_N4BEG[15] ,
    \Tile_X5Y14_N4BEG[14] ,
    \Tile_X5Y14_N4BEG[13] ,
    \Tile_X5Y14_N4BEG[12] ,
    \Tile_X5Y14_N4BEG[11] ,
    \Tile_X5Y14_N4BEG[10] ,
    \Tile_X5Y14_N4BEG[9] ,
    \Tile_X5Y14_N4BEG[8] ,
    \Tile_X5Y14_N4BEG[7] ,
    \Tile_X5Y14_N4BEG[6] ,
    \Tile_X5Y14_N4BEG[5] ,
    \Tile_X5Y14_N4BEG[4] ,
    \Tile_X5Y14_N4BEG[3] ,
    \Tile_X5Y14_N4BEG[2] ,
    \Tile_X5Y14_N4BEG[1] ,
    \Tile_X5Y14_N4BEG[0] }),
    .NN4BEG({\Tile_X5Y13_NN4BEG[15] ,
    \Tile_X5Y13_NN4BEG[14] ,
    \Tile_X5Y13_NN4BEG[13] ,
    \Tile_X5Y13_NN4BEG[12] ,
    \Tile_X5Y13_NN4BEG[11] ,
    \Tile_X5Y13_NN4BEG[10] ,
    \Tile_X5Y13_NN4BEG[9] ,
    \Tile_X5Y13_NN4BEG[8] ,
    \Tile_X5Y13_NN4BEG[7] ,
    \Tile_X5Y13_NN4BEG[6] ,
    \Tile_X5Y13_NN4BEG[5] ,
    \Tile_X5Y13_NN4BEG[4] ,
    \Tile_X5Y13_NN4BEG[3] ,
    \Tile_X5Y13_NN4BEG[2] ,
    \Tile_X5Y13_NN4BEG[1] ,
    \Tile_X5Y13_NN4BEG[0] }),
    .NN4END({\Tile_X5Y14_NN4BEG[15] ,
    \Tile_X5Y14_NN4BEG[14] ,
    \Tile_X5Y14_NN4BEG[13] ,
    \Tile_X5Y14_NN4BEG[12] ,
    \Tile_X5Y14_NN4BEG[11] ,
    \Tile_X5Y14_NN4BEG[10] ,
    \Tile_X5Y14_NN4BEG[9] ,
    \Tile_X5Y14_NN4BEG[8] ,
    \Tile_X5Y14_NN4BEG[7] ,
    \Tile_X5Y14_NN4BEG[6] ,
    \Tile_X5Y14_NN4BEG[5] ,
    \Tile_X5Y14_NN4BEG[4] ,
    \Tile_X5Y14_NN4BEG[3] ,
    \Tile_X5Y14_NN4BEG[2] ,
    \Tile_X5Y14_NN4BEG[1] ,
    \Tile_X5Y14_NN4BEG[0] }),
    .S1BEG({\Tile_X5Y13_S1BEG[3] ,
    \Tile_X5Y13_S1BEG[2] ,
    \Tile_X5Y13_S1BEG[1] ,
    \Tile_X5Y13_S1BEG[0] }),
    .S1END({\Tile_X5Y12_S1BEG[3] ,
    \Tile_X5Y12_S1BEG[2] ,
    \Tile_X5Y12_S1BEG[1] ,
    \Tile_X5Y12_S1BEG[0] }),
    .S2BEG({\Tile_X5Y13_S2BEG[7] ,
    \Tile_X5Y13_S2BEG[6] ,
    \Tile_X5Y13_S2BEG[5] ,
    \Tile_X5Y13_S2BEG[4] ,
    \Tile_X5Y13_S2BEG[3] ,
    \Tile_X5Y13_S2BEG[2] ,
    \Tile_X5Y13_S2BEG[1] ,
    \Tile_X5Y13_S2BEG[0] }),
    .S2BEGb({\Tile_X5Y13_S2BEGb[7] ,
    \Tile_X5Y13_S2BEGb[6] ,
    \Tile_X5Y13_S2BEGb[5] ,
    \Tile_X5Y13_S2BEGb[4] ,
    \Tile_X5Y13_S2BEGb[3] ,
    \Tile_X5Y13_S2BEGb[2] ,
    \Tile_X5Y13_S2BEGb[1] ,
    \Tile_X5Y13_S2BEGb[0] }),
    .S2END({\Tile_X5Y12_S2BEGb[7] ,
    \Tile_X5Y12_S2BEGb[6] ,
    \Tile_X5Y12_S2BEGb[5] ,
    \Tile_X5Y12_S2BEGb[4] ,
    \Tile_X5Y12_S2BEGb[3] ,
    \Tile_X5Y12_S2BEGb[2] ,
    \Tile_X5Y12_S2BEGb[1] ,
    \Tile_X5Y12_S2BEGb[0] }),
    .S2MID({\Tile_X5Y12_S2BEG[7] ,
    \Tile_X5Y12_S2BEG[6] ,
    \Tile_X5Y12_S2BEG[5] ,
    \Tile_X5Y12_S2BEG[4] ,
    \Tile_X5Y12_S2BEG[3] ,
    \Tile_X5Y12_S2BEG[2] ,
    \Tile_X5Y12_S2BEG[1] ,
    \Tile_X5Y12_S2BEG[0] }),
    .S4BEG({\Tile_X5Y13_S4BEG[15] ,
    \Tile_X5Y13_S4BEG[14] ,
    \Tile_X5Y13_S4BEG[13] ,
    \Tile_X5Y13_S4BEG[12] ,
    \Tile_X5Y13_S4BEG[11] ,
    \Tile_X5Y13_S4BEG[10] ,
    \Tile_X5Y13_S4BEG[9] ,
    \Tile_X5Y13_S4BEG[8] ,
    \Tile_X5Y13_S4BEG[7] ,
    \Tile_X5Y13_S4BEG[6] ,
    \Tile_X5Y13_S4BEG[5] ,
    \Tile_X5Y13_S4BEG[4] ,
    \Tile_X5Y13_S4BEG[3] ,
    \Tile_X5Y13_S4BEG[2] ,
    \Tile_X5Y13_S4BEG[1] ,
    \Tile_X5Y13_S4BEG[0] }),
    .S4END({\Tile_X5Y12_S4BEG[15] ,
    \Tile_X5Y12_S4BEG[14] ,
    \Tile_X5Y12_S4BEG[13] ,
    \Tile_X5Y12_S4BEG[12] ,
    \Tile_X5Y12_S4BEG[11] ,
    \Tile_X5Y12_S4BEG[10] ,
    \Tile_X5Y12_S4BEG[9] ,
    \Tile_X5Y12_S4BEG[8] ,
    \Tile_X5Y12_S4BEG[7] ,
    \Tile_X5Y12_S4BEG[6] ,
    \Tile_X5Y12_S4BEG[5] ,
    \Tile_X5Y12_S4BEG[4] ,
    \Tile_X5Y12_S4BEG[3] ,
    \Tile_X5Y12_S4BEG[2] ,
    \Tile_X5Y12_S4BEG[1] ,
    \Tile_X5Y12_S4BEG[0] }),
    .SS4BEG({\Tile_X5Y13_SS4BEG[15] ,
    \Tile_X5Y13_SS4BEG[14] ,
    \Tile_X5Y13_SS4BEG[13] ,
    \Tile_X5Y13_SS4BEG[12] ,
    \Tile_X5Y13_SS4BEG[11] ,
    \Tile_X5Y13_SS4BEG[10] ,
    \Tile_X5Y13_SS4BEG[9] ,
    \Tile_X5Y13_SS4BEG[8] ,
    \Tile_X5Y13_SS4BEG[7] ,
    \Tile_X5Y13_SS4BEG[6] ,
    \Tile_X5Y13_SS4BEG[5] ,
    \Tile_X5Y13_SS4BEG[4] ,
    \Tile_X5Y13_SS4BEG[3] ,
    \Tile_X5Y13_SS4BEG[2] ,
    \Tile_X5Y13_SS4BEG[1] ,
    \Tile_X5Y13_SS4BEG[0] }),
    .SS4END({\Tile_X5Y12_SS4BEG[15] ,
    \Tile_X5Y12_SS4BEG[14] ,
    \Tile_X5Y12_SS4BEG[13] ,
    \Tile_X5Y12_SS4BEG[12] ,
    \Tile_X5Y12_SS4BEG[11] ,
    \Tile_X5Y12_SS4BEG[10] ,
    \Tile_X5Y12_SS4BEG[9] ,
    \Tile_X5Y12_SS4BEG[8] ,
    \Tile_X5Y12_SS4BEG[7] ,
    \Tile_X5Y12_SS4BEG[6] ,
    \Tile_X5Y12_SS4BEG[5] ,
    \Tile_X5Y12_SS4BEG[4] ,
    \Tile_X5Y12_SS4BEG[3] ,
    \Tile_X5Y12_SS4BEG[2] ,
    \Tile_X5Y12_SS4BEG[1] ,
    \Tile_X5Y12_SS4BEG[0] }),
    .W1BEG({\Tile_X5Y13_W1BEG[3] ,
    \Tile_X5Y13_W1BEG[2] ,
    \Tile_X5Y13_W1BEG[1] ,
    \Tile_X5Y13_W1BEG[0] }),
    .W1END({\Tile_X6Y13_W1BEG[3] ,
    \Tile_X6Y13_W1BEG[2] ,
    \Tile_X6Y13_W1BEG[1] ,
    \Tile_X6Y13_W1BEG[0] }),
    .W2BEG({\Tile_X5Y13_W2BEG[7] ,
    \Tile_X5Y13_W2BEG[6] ,
    \Tile_X5Y13_W2BEG[5] ,
    \Tile_X5Y13_W2BEG[4] ,
    \Tile_X5Y13_W2BEG[3] ,
    \Tile_X5Y13_W2BEG[2] ,
    \Tile_X5Y13_W2BEG[1] ,
    \Tile_X5Y13_W2BEG[0] }),
    .W2BEGb({\Tile_X5Y13_W2BEGb[7] ,
    \Tile_X5Y13_W2BEGb[6] ,
    \Tile_X5Y13_W2BEGb[5] ,
    \Tile_X5Y13_W2BEGb[4] ,
    \Tile_X5Y13_W2BEGb[3] ,
    \Tile_X5Y13_W2BEGb[2] ,
    \Tile_X5Y13_W2BEGb[1] ,
    \Tile_X5Y13_W2BEGb[0] }),
    .W2END({\Tile_X6Y13_W2BEGb[7] ,
    \Tile_X6Y13_W2BEGb[6] ,
    \Tile_X6Y13_W2BEGb[5] ,
    \Tile_X6Y13_W2BEGb[4] ,
    \Tile_X6Y13_W2BEGb[3] ,
    \Tile_X6Y13_W2BEGb[2] ,
    \Tile_X6Y13_W2BEGb[1] ,
    \Tile_X6Y13_W2BEGb[0] }),
    .W2MID({\Tile_X6Y13_W2BEG[7] ,
    \Tile_X6Y13_W2BEG[6] ,
    \Tile_X6Y13_W2BEG[5] ,
    \Tile_X6Y13_W2BEG[4] ,
    \Tile_X6Y13_W2BEG[3] ,
    \Tile_X6Y13_W2BEG[2] ,
    \Tile_X6Y13_W2BEG[1] ,
    \Tile_X6Y13_W2BEG[0] }),
    .W6BEG({\Tile_X5Y13_W6BEG[11] ,
    \Tile_X5Y13_W6BEG[10] ,
    \Tile_X5Y13_W6BEG[9] ,
    \Tile_X5Y13_W6BEG[8] ,
    \Tile_X5Y13_W6BEG[7] ,
    \Tile_X5Y13_W6BEG[6] ,
    \Tile_X5Y13_W6BEG[5] ,
    \Tile_X5Y13_W6BEG[4] ,
    \Tile_X5Y13_W6BEG[3] ,
    \Tile_X5Y13_W6BEG[2] ,
    \Tile_X5Y13_W6BEG[1] ,
    \Tile_X5Y13_W6BEG[0] }),
    .W6END({\Tile_X6Y13_W6BEG[11] ,
    \Tile_X6Y13_W6BEG[10] ,
    \Tile_X6Y13_W6BEG[9] ,
    \Tile_X6Y13_W6BEG[8] ,
    \Tile_X6Y13_W6BEG[7] ,
    \Tile_X6Y13_W6BEG[6] ,
    \Tile_X6Y13_W6BEG[5] ,
    \Tile_X6Y13_W6BEG[4] ,
    \Tile_X6Y13_W6BEG[3] ,
    \Tile_X6Y13_W6BEG[2] ,
    \Tile_X6Y13_W6BEG[1] ,
    \Tile_X6Y13_W6BEG[0] }),
    .WW4BEG({\Tile_X5Y13_WW4BEG[15] ,
    \Tile_X5Y13_WW4BEG[14] ,
    \Tile_X5Y13_WW4BEG[13] ,
    \Tile_X5Y13_WW4BEG[12] ,
    \Tile_X5Y13_WW4BEG[11] ,
    \Tile_X5Y13_WW4BEG[10] ,
    \Tile_X5Y13_WW4BEG[9] ,
    \Tile_X5Y13_WW4BEG[8] ,
    \Tile_X5Y13_WW4BEG[7] ,
    \Tile_X5Y13_WW4BEG[6] ,
    \Tile_X5Y13_WW4BEG[5] ,
    \Tile_X5Y13_WW4BEG[4] ,
    \Tile_X5Y13_WW4BEG[3] ,
    \Tile_X5Y13_WW4BEG[2] ,
    \Tile_X5Y13_WW4BEG[1] ,
    \Tile_X5Y13_WW4BEG[0] }),
    .WW4END({\Tile_X6Y13_WW4BEG[15] ,
    \Tile_X6Y13_WW4BEG[14] ,
    \Tile_X6Y13_WW4BEG[13] ,
    \Tile_X6Y13_WW4BEG[12] ,
    \Tile_X6Y13_WW4BEG[11] ,
    \Tile_X6Y13_WW4BEG[10] ,
    \Tile_X6Y13_WW4BEG[9] ,
    \Tile_X6Y13_WW4BEG[8] ,
    \Tile_X6Y13_WW4BEG[7] ,
    \Tile_X6Y13_WW4BEG[6] ,
    \Tile_X6Y13_WW4BEG[5] ,
    \Tile_X6Y13_WW4BEG[4] ,
    \Tile_X6Y13_WW4BEG[3] ,
    \Tile_X6Y13_WW4BEG[2] ,
    \Tile_X6Y13_WW4BEG[1] ,
    \Tile_X6Y13_WW4BEG[0] }));
 LUT4AB Tile_X5Y14_LUT4AB (.Ci(Tile_X5Y15_Co),
    .Co(Tile_X5Y14_Co),
    .UserCLK(Tile_X5Y15_UserCLKo),
    .UserCLKo(Tile_X5Y14_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X5Y14_E1BEG[3] ,
    \Tile_X5Y14_E1BEG[2] ,
    \Tile_X5Y14_E1BEG[1] ,
    \Tile_X5Y14_E1BEG[0] }),
    .E1END({\Tile_X4Y14_E1BEG[3] ,
    \Tile_X4Y14_E1BEG[2] ,
    \Tile_X4Y14_E1BEG[1] ,
    \Tile_X4Y14_E1BEG[0] }),
    .E2BEG({\Tile_X5Y14_E2BEG[7] ,
    \Tile_X5Y14_E2BEG[6] ,
    \Tile_X5Y14_E2BEG[5] ,
    \Tile_X5Y14_E2BEG[4] ,
    \Tile_X5Y14_E2BEG[3] ,
    \Tile_X5Y14_E2BEG[2] ,
    \Tile_X5Y14_E2BEG[1] ,
    \Tile_X5Y14_E2BEG[0] }),
    .E2BEGb({\Tile_X5Y14_E2BEGb[7] ,
    \Tile_X5Y14_E2BEGb[6] ,
    \Tile_X5Y14_E2BEGb[5] ,
    \Tile_X5Y14_E2BEGb[4] ,
    \Tile_X5Y14_E2BEGb[3] ,
    \Tile_X5Y14_E2BEGb[2] ,
    \Tile_X5Y14_E2BEGb[1] ,
    \Tile_X5Y14_E2BEGb[0] }),
    .E2END({\Tile_X4Y14_E2BEGb[7] ,
    \Tile_X4Y14_E2BEGb[6] ,
    \Tile_X4Y14_E2BEGb[5] ,
    \Tile_X4Y14_E2BEGb[4] ,
    \Tile_X4Y14_E2BEGb[3] ,
    \Tile_X4Y14_E2BEGb[2] ,
    \Tile_X4Y14_E2BEGb[1] ,
    \Tile_X4Y14_E2BEGb[0] }),
    .E2MID({\Tile_X4Y14_E2BEG[7] ,
    \Tile_X4Y14_E2BEG[6] ,
    \Tile_X4Y14_E2BEG[5] ,
    \Tile_X4Y14_E2BEG[4] ,
    \Tile_X4Y14_E2BEG[3] ,
    \Tile_X4Y14_E2BEG[2] ,
    \Tile_X4Y14_E2BEG[1] ,
    \Tile_X4Y14_E2BEG[0] }),
    .E6BEG({\Tile_X5Y14_E6BEG[11] ,
    \Tile_X5Y14_E6BEG[10] ,
    \Tile_X5Y14_E6BEG[9] ,
    \Tile_X5Y14_E6BEG[8] ,
    \Tile_X5Y14_E6BEG[7] ,
    \Tile_X5Y14_E6BEG[6] ,
    \Tile_X5Y14_E6BEG[5] ,
    \Tile_X5Y14_E6BEG[4] ,
    \Tile_X5Y14_E6BEG[3] ,
    \Tile_X5Y14_E6BEG[2] ,
    \Tile_X5Y14_E6BEG[1] ,
    \Tile_X5Y14_E6BEG[0] }),
    .E6END({\Tile_X4Y14_E6BEG[11] ,
    \Tile_X4Y14_E6BEG[10] ,
    \Tile_X4Y14_E6BEG[9] ,
    \Tile_X4Y14_E6BEG[8] ,
    \Tile_X4Y14_E6BEG[7] ,
    \Tile_X4Y14_E6BEG[6] ,
    \Tile_X4Y14_E6BEG[5] ,
    \Tile_X4Y14_E6BEG[4] ,
    \Tile_X4Y14_E6BEG[3] ,
    \Tile_X4Y14_E6BEG[2] ,
    \Tile_X4Y14_E6BEG[1] ,
    \Tile_X4Y14_E6BEG[0] }),
    .EE4BEG({\Tile_X5Y14_EE4BEG[15] ,
    \Tile_X5Y14_EE4BEG[14] ,
    \Tile_X5Y14_EE4BEG[13] ,
    \Tile_X5Y14_EE4BEG[12] ,
    \Tile_X5Y14_EE4BEG[11] ,
    \Tile_X5Y14_EE4BEG[10] ,
    \Tile_X5Y14_EE4BEG[9] ,
    \Tile_X5Y14_EE4BEG[8] ,
    \Tile_X5Y14_EE4BEG[7] ,
    \Tile_X5Y14_EE4BEG[6] ,
    \Tile_X5Y14_EE4BEG[5] ,
    \Tile_X5Y14_EE4BEG[4] ,
    \Tile_X5Y14_EE4BEG[3] ,
    \Tile_X5Y14_EE4BEG[2] ,
    \Tile_X5Y14_EE4BEG[1] ,
    \Tile_X5Y14_EE4BEG[0] }),
    .EE4END({\Tile_X4Y14_EE4BEG[15] ,
    \Tile_X4Y14_EE4BEG[14] ,
    \Tile_X4Y14_EE4BEG[13] ,
    \Tile_X4Y14_EE4BEG[12] ,
    \Tile_X4Y14_EE4BEG[11] ,
    \Tile_X4Y14_EE4BEG[10] ,
    \Tile_X4Y14_EE4BEG[9] ,
    \Tile_X4Y14_EE4BEG[8] ,
    \Tile_X4Y14_EE4BEG[7] ,
    \Tile_X4Y14_EE4BEG[6] ,
    \Tile_X4Y14_EE4BEG[5] ,
    \Tile_X4Y14_EE4BEG[4] ,
    \Tile_X4Y14_EE4BEG[3] ,
    \Tile_X4Y14_EE4BEG[2] ,
    \Tile_X4Y14_EE4BEG[1] ,
    \Tile_X4Y14_EE4BEG[0] }),
    .FrameData({\Tile_X4Y14_FrameData_O[31] ,
    \Tile_X4Y14_FrameData_O[30] ,
    \Tile_X4Y14_FrameData_O[29] ,
    \Tile_X4Y14_FrameData_O[28] ,
    \Tile_X4Y14_FrameData_O[27] ,
    \Tile_X4Y14_FrameData_O[26] ,
    \Tile_X4Y14_FrameData_O[25] ,
    \Tile_X4Y14_FrameData_O[24] ,
    \Tile_X4Y14_FrameData_O[23] ,
    \Tile_X4Y14_FrameData_O[22] ,
    \Tile_X4Y14_FrameData_O[21] ,
    \Tile_X4Y14_FrameData_O[20] ,
    \Tile_X4Y14_FrameData_O[19] ,
    \Tile_X4Y14_FrameData_O[18] ,
    \Tile_X4Y14_FrameData_O[17] ,
    \Tile_X4Y14_FrameData_O[16] ,
    \Tile_X4Y14_FrameData_O[15] ,
    \Tile_X4Y14_FrameData_O[14] ,
    \Tile_X4Y14_FrameData_O[13] ,
    \Tile_X4Y14_FrameData_O[12] ,
    \Tile_X4Y14_FrameData_O[11] ,
    \Tile_X4Y14_FrameData_O[10] ,
    \Tile_X4Y14_FrameData_O[9] ,
    \Tile_X4Y14_FrameData_O[8] ,
    \Tile_X4Y14_FrameData_O[7] ,
    \Tile_X4Y14_FrameData_O[6] ,
    \Tile_X4Y14_FrameData_O[5] ,
    \Tile_X4Y14_FrameData_O[4] ,
    \Tile_X4Y14_FrameData_O[3] ,
    \Tile_X4Y14_FrameData_O[2] ,
    \Tile_X4Y14_FrameData_O[1] ,
    \Tile_X4Y14_FrameData_O[0] }),
    .FrameData_O({\Tile_X5Y14_FrameData_O[31] ,
    \Tile_X5Y14_FrameData_O[30] ,
    \Tile_X5Y14_FrameData_O[29] ,
    \Tile_X5Y14_FrameData_O[28] ,
    \Tile_X5Y14_FrameData_O[27] ,
    \Tile_X5Y14_FrameData_O[26] ,
    \Tile_X5Y14_FrameData_O[25] ,
    \Tile_X5Y14_FrameData_O[24] ,
    \Tile_X5Y14_FrameData_O[23] ,
    \Tile_X5Y14_FrameData_O[22] ,
    \Tile_X5Y14_FrameData_O[21] ,
    \Tile_X5Y14_FrameData_O[20] ,
    \Tile_X5Y14_FrameData_O[19] ,
    \Tile_X5Y14_FrameData_O[18] ,
    \Tile_X5Y14_FrameData_O[17] ,
    \Tile_X5Y14_FrameData_O[16] ,
    \Tile_X5Y14_FrameData_O[15] ,
    \Tile_X5Y14_FrameData_O[14] ,
    \Tile_X5Y14_FrameData_O[13] ,
    \Tile_X5Y14_FrameData_O[12] ,
    \Tile_X5Y14_FrameData_O[11] ,
    \Tile_X5Y14_FrameData_O[10] ,
    \Tile_X5Y14_FrameData_O[9] ,
    \Tile_X5Y14_FrameData_O[8] ,
    \Tile_X5Y14_FrameData_O[7] ,
    \Tile_X5Y14_FrameData_O[6] ,
    \Tile_X5Y14_FrameData_O[5] ,
    \Tile_X5Y14_FrameData_O[4] ,
    \Tile_X5Y14_FrameData_O[3] ,
    \Tile_X5Y14_FrameData_O[2] ,
    \Tile_X5Y14_FrameData_O[1] ,
    \Tile_X5Y14_FrameData_O[0] }),
    .FrameStrobe({\Tile_X5Y15_FrameStrobe_O[19] ,
    \Tile_X5Y15_FrameStrobe_O[18] ,
    \Tile_X5Y15_FrameStrobe_O[17] ,
    \Tile_X5Y15_FrameStrobe_O[16] ,
    \Tile_X5Y15_FrameStrobe_O[15] ,
    \Tile_X5Y15_FrameStrobe_O[14] ,
    \Tile_X5Y15_FrameStrobe_O[13] ,
    \Tile_X5Y15_FrameStrobe_O[12] ,
    \Tile_X5Y15_FrameStrobe_O[11] ,
    \Tile_X5Y15_FrameStrobe_O[10] ,
    \Tile_X5Y15_FrameStrobe_O[9] ,
    \Tile_X5Y15_FrameStrobe_O[8] ,
    \Tile_X5Y15_FrameStrobe_O[7] ,
    \Tile_X5Y15_FrameStrobe_O[6] ,
    \Tile_X5Y15_FrameStrobe_O[5] ,
    \Tile_X5Y15_FrameStrobe_O[4] ,
    \Tile_X5Y15_FrameStrobe_O[3] ,
    \Tile_X5Y15_FrameStrobe_O[2] ,
    \Tile_X5Y15_FrameStrobe_O[1] ,
    \Tile_X5Y15_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X5Y14_FrameStrobe_O[19] ,
    \Tile_X5Y14_FrameStrobe_O[18] ,
    \Tile_X5Y14_FrameStrobe_O[17] ,
    \Tile_X5Y14_FrameStrobe_O[16] ,
    \Tile_X5Y14_FrameStrobe_O[15] ,
    \Tile_X5Y14_FrameStrobe_O[14] ,
    \Tile_X5Y14_FrameStrobe_O[13] ,
    \Tile_X5Y14_FrameStrobe_O[12] ,
    \Tile_X5Y14_FrameStrobe_O[11] ,
    \Tile_X5Y14_FrameStrobe_O[10] ,
    \Tile_X5Y14_FrameStrobe_O[9] ,
    \Tile_X5Y14_FrameStrobe_O[8] ,
    \Tile_X5Y14_FrameStrobe_O[7] ,
    \Tile_X5Y14_FrameStrobe_O[6] ,
    \Tile_X5Y14_FrameStrobe_O[5] ,
    \Tile_X5Y14_FrameStrobe_O[4] ,
    \Tile_X5Y14_FrameStrobe_O[3] ,
    \Tile_X5Y14_FrameStrobe_O[2] ,
    \Tile_X5Y14_FrameStrobe_O[1] ,
    \Tile_X5Y14_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X5Y14_N1BEG[3] ,
    \Tile_X5Y14_N1BEG[2] ,
    \Tile_X5Y14_N1BEG[1] ,
    \Tile_X5Y14_N1BEG[0] }),
    .N1END({\Tile_X5Y15_N1BEG[3] ,
    \Tile_X5Y15_N1BEG[2] ,
    \Tile_X5Y15_N1BEG[1] ,
    \Tile_X5Y15_N1BEG[0] }),
    .N2BEG({\Tile_X5Y14_N2BEG[7] ,
    \Tile_X5Y14_N2BEG[6] ,
    \Tile_X5Y14_N2BEG[5] ,
    \Tile_X5Y14_N2BEG[4] ,
    \Tile_X5Y14_N2BEG[3] ,
    \Tile_X5Y14_N2BEG[2] ,
    \Tile_X5Y14_N2BEG[1] ,
    \Tile_X5Y14_N2BEG[0] }),
    .N2BEGb({\Tile_X5Y14_N2BEGb[7] ,
    \Tile_X5Y14_N2BEGb[6] ,
    \Tile_X5Y14_N2BEGb[5] ,
    \Tile_X5Y14_N2BEGb[4] ,
    \Tile_X5Y14_N2BEGb[3] ,
    \Tile_X5Y14_N2BEGb[2] ,
    \Tile_X5Y14_N2BEGb[1] ,
    \Tile_X5Y14_N2BEGb[0] }),
    .N2END({\Tile_X5Y15_N2BEGb[7] ,
    \Tile_X5Y15_N2BEGb[6] ,
    \Tile_X5Y15_N2BEGb[5] ,
    \Tile_X5Y15_N2BEGb[4] ,
    \Tile_X5Y15_N2BEGb[3] ,
    \Tile_X5Y15_N2BEGb[2] ,
    \Tile_X5Y15_N2BEGb[1] ,
    \Tile_X5Y15_N2BEGb[0] }),
    .N2MID({\Tile_X5Y15_N2BEG[7] ,
    \Tile_X5Y15_N2BEG[6] ,
    \Tile_X5Y15_N2BEG[5] ,
    \Tile_X5Y15_N2BEG[4] ,
    \Tile_X5Y15_N2BEG[3] ,
    \Tile_X5Y15_N2BEG[2] ,
    \Tile_X5Y15_N2BEG[1] ,
    \Tile_X5Y15_N2BEG[0] }),
    .N4BEG({\Tile_X5Y14_N4BEG[15] ,
    \Tile_X5Y14_N4BEG[14] ,
    \Tile_X5Y14_N4BEG[13] ,
    \Tile_X5Y14_N4BEG[12] ,
    \Tile_X5Y14_N4BEG[11] ,
    \Tile_X5Y14_N4BEG[10] ,
    \Tile_X5Y14_N4BEG[9] ,
    \Tile_X5Y14_N4BEG[8] ,
    \Tile_X5Y14_N4BEG[7] ,
    \Tile_X5Y14_N4BEG[6] ,
    \Tile_X5Y14_N4BEG[5] ,
    \Tile_X5Y14_N4BEG[4] ,
    \Tile_X5Y14_N4BEG[3] ,
    \Tile_X5Y14_N4BEG[2] ,
    \Tile_X5Y14_N4BEG[1] ,
    \Tile_X5Y14_N4BEG[0] }),
    .N4END({\Tile_X5Y15_N4BEG[15] ,
    \Tile_X5Y15_N4BEG[14] ,
    \Tile_X5Y15_N4BEG[13] ,
    \Tile_X5Y15_N4BEG[12] ,
    \Tile_X5Y15_N4BEG[11] ,
    \Tile_X5Y15_N4BEG[10] ,
    \Tile_X5Y15_N4BEG[9] ,
    \Tile_X5Y15_N4BEG[8] ,
    \Tile_X5Y15_N4BEG[7] ,
    \Tile_X5Y15_N4BEG[6] ,
    \Tile_X5Y15_N4BEG[5] ,
    \Tile_X5Y15_N4BEG[4] ,
    \Tile_X5Y15_N4BEG[3] ,
    \Tile_X5Y15_N4BEG[2] ,
    \Tile_X5Y15_N4BEG[1] ,
    \Tile_X5Y15_N4BEG[0] }),
    .NN4BEG({\Tile_X5Y14_NN4BEG[15] ,
    \Tile_X5Y14_NN4BEG[14] ,
    \Tile_X5Y14_NN4BEG[13] ,
    \Tile_X5Y14_NN4BEG[12] ,
    \Tile_X5Y14_NN4BEG[11] ,
    \Tile_X5Y14_NN4BEG[10] ,
    \Tile_X5Y14_NN4BEG[9] ,
    \Tile_X5Y14_NN4BEG[8] ,
    \Tile_X5Y14_NN4BEG[7] ,
    \Tile_X5Y14_NN4BEG[6] ,
    \Tile_X5Y14_NN4BEG[5] ,
    \Tile_X5Y14_NN4BEG[4] ,
    \Tile_X5Y14_NN4BEG[3] ,
    \Tile_X5Y14_NN4BEG[2] ,
    \Tile_X5Y14_NN4BEG[1] ,
    \Tile_X5Y14_NN4BEG[0] }),
    .NN4END({\Tile_X5Y15_NN4BEG[15] ,
    \Tile_X5Y15_NN4BEG[14] ,
    \Tile_X5Y15_NN4BEG[13] ,
    \Tile_X5Y15_NN4BEG[12] ,
    \Tile_X5Y15_NN4BEG[11] ,
    \Tile_X5Y15_NN4BEG[10] ,
    \Tile_X5Y15_NN4BEG[9] ,
    \Tile_X5Y15_NN4BEG[8] ,
    \Tile_X5Y15_NN4BEG[7] ,
    \Tile_X5Y15_NN4BEG[6] ,
    \Tile_X5Y15_NN4BEG[5] ,
    \Tile_X5Y15_NN4BEG[4] ,
    \Tile_X5Y15_NN4BEG[3] ,
    \Tile_X5Y15_NN4BEG[2] ,
    \Tile_X5Y15_NN4BEG[1] ,
    \Tile_X5Y15_NN4BEG[0] }),
    .S1BEG({\Tile_X5Y14_S1BEG[3] ,
    \Tile_X5Y14_S1BEG[2] ,
    \Tile_X5Y14_S1BEG[1] ,
    \Tile_X5Y14_S1BEG[0] }),
    .S1END({\Tile_X5Y13_S1BEG[3] ,
    \Tile_X5Y13_S1BEG[2] ,
    \Tile_X5Y13_S1BEG[1] ,
    \Tile_X5Y13_S1BEG[0] }),
    .S2BEG({\Tile_X5Y14_S2BEG[7] ,
    \Tile_X5Y14_S2BEG[6] ,
    \Tile_X5Y14_S2BEG[5] ,
    \Tile_X5Y14_S2BEG[4] ,
    \Tile_X5Y14_S2BEG[3] ,
    \Tile_X5Y14_S2BEG[2] ,
    \Tile_X5Y14_S2BEG[1] ,
    \Tile_X5Y14_S2BEG[0] }),
    .S2BEGb({\Tile_X5Y14_S2BEGb[7] ,
    \Tile_X5Y14_S2BEGb[6] ,
    \Tile_X5Y14_S2BEGb[5] ,
    \Tile_X5Y14_S2BEGb[4] ,
    \Tile_X5Y14_S2BEGb[3] ,
    \Tile_X5Y14_S2BEGb[2] ,
    \Tile_X5Y14_S2BEGb[1] ,
    \Tile_X5Y14_S2BEGb[0] }),
    .S2END({\Tile_X5Y13_S2BEGb[7] ,
    \Tile_X5Y13_S2BEGb[6] ,
    \Tile_X5Y13_S2BEGb[5] ,
    \Tile_X5Y13_S2BEGb[4] ,
    \Tile_X5Y13_S2BEGb[3] ,
    \Tile_X5Y13_S2BEGb[2] ,
    \Tile_X5Y13_S2BEGb[1] ,
    \Tile_X5Y13_S2BEGb[0] }),
    .S2MID({\Tile_X5Y13_S2BEG[7] ,
    \Tile_X5Y13_S2BEG[6] ,
    \Tile_X5Y13_S2BEG[5] ,
    \Tile_X5Y13_S2BEG[4] ,
    \Tile_X5Y13_S2BEG[3] ,
    \Tile_X5Y13_S2BEG[2] ,
    \Tile_X5Y13_S2BEG[1] ,
    \Tile_X5Y13_S2BEG[0] }),
    .S4BEG({\Tile_X5Y14_S4BEG[15] ,
    \Tile_X5Y14_S4BEG[14] ,
    \Tile_X5Y14_S4BEG[13] ,
    \Tile_X5Y14_S4BEG[12] ,
    \Tile_X5Y14_S4BEG[11] ,
    \Tile_X5Y14_S4BEG[10] ,
    \Tile_X5Y14_S4BEG[9] ,
    \Tile_X5Y14_S4BEG[8] ,
    \Tile_X5Y14_S4BEG[7] ,
    \Tile_X5Y14_S4BEG[6] ,
    \Tile_X5Y14_S4BEG[5] ,
    \Tile_X5Y14_S4BEG[4] ,
    \Tile_X5Y14_S4BEG[3] ,
    \Tile_X5Y14_S4BEG[2] ,
    \Tile_X5Y14_S4BEG[1] ,
    \Tile_X5Y14_S4BEG[0] }),
    .S4END({\Tile_X5Y13_S4BEG[15] ,
    \Tile_X5Y13_S4BEG[14] ,
    \Tile_X5Y13_S4BEG[13] ,
    \Tile_X5Y13_S4BEG[12] ,
    \Tile_X5Y13_S4BEG[11] ,
    \Tile_X5Y13_S4BEG[10] ,
    \Tile_X5Y13_S4BEG[9] ,
    \Tile_X5Y13_S4BEG[8] ,
    \Tile_X5Y13_S4BEG[7] ,
    \Tile_X5Y13_S4BEG[6] ,
    \Tile_X5Y13_S4BEG[5] ,
    \Tile_X5Y13_S4BEG[4] ,
    \Tile_X5Y13_S4BEG[3] ,
    \Tile_X5Y13_S4BEG[2] ,
    \Tile_X5Y13_S4BEG[1] ,
    \Tile_X5Y13_S4BEG[0] }),
    .SS4BEG({\Tile_X5Y14_SS4BEG[15] ,
    \Tile_X5Y14_SS4BEG[14] ,
    \Tile_X5Y14_SS4BEG[13] ,
    \Tile_X5Y14_SS4BEG[12] ,
    \Tile_X5Y14_SS4BEG[11] ,
    \Tile_X5Y14_SS4BEG[10] ,
    \Tile_X5Y14_SS4BEG[9] ,
    \Tile_X5Y14_SS4BEG[8] ,
    \Tile_X5Y14_SS4BEG[7] ,
    \Tile_X5Y14_SS4BEG[6] ,
    \Tile_X5Y14_SS4BEG[5] ,
    \Tile_X5Y14_SS4BEG[4] ,
    \Tile_X5Y14_SS4BEG[3] ,
    \Tile_X5Y14_SS4BEG[2] ,
    \Tile_X5Y14_SS4BEG[1] ,
    \Tile_X5Y14_SS4BEG[0] }),
    .SS4END({\Tile_X5Y13_SS4BEG[15] ,
    \Tile_X5Y13_SS4BEG[14] ,
    \Tile_X5Y13_SS4BEG[13] ,
    \Tile_X5Y13_SS4BEG[12] ,
    \Tile_X5Y13_SS4BEG[11] ,
    \Tile_X5Y13_SS4BEG[10] ,
    \Tile_X5Y13_SS4BEG[9] ,
    \Tile_X5Y13_SS4BEG[8] ,
    \Tile_X5Y13_SS4BEG[7] ,
    \Tile_X5Y13_SS4BEG[6] ,
    \Tile_X5Y13_SS4BEG[5] ,
    \Tile_X5Y13_SS4BEG[4] ,
    \Tile_X5Y13_SS4BEG[3] ,
    \Tile_X5Y13_SS4BEG[2] ,
    \Tile_X5Y13_SS4BEG[1] ,
    \Tile_X5Y13_SS4BEG[0] }),
    .W1BEG({\Tile_X5Y14_W1BEG[3] ,
    \Tile_X5Y14_W1BEG[2] ,
    \Tile_X5Y14_W1BEG[1] ,
    \Tile_X5Y14_W1BEG[0] }),
    .W1END({\Tile_X6Y14_W1BEG[3] ,
    \Tile_X6Y14_W1BEG[2] ,
    \Tile_X6Y14_W1BEG[1] ,
    \Tile_X6Y14_W1BEG[0] }),
    .W2BEG({\Tile_X5Y14_W2BEG[7] ,
    \Tile_X5Y14_W2BEG[6] ,
    \Tile_X5Y14_W2BEG[5] ,
    \Tile_X5Y14_W2BEG[4] ,
    \Tile_X5Y14_W2BEG[3] ,
    \Tile_X5Y14_W2BEG[2] ,
    \Tile_X5Y14_W2BEG[1] ,
    \Tile_X5Y14_W2BEG[0] }),
    .W2BEGb({\Tile_X5Y14_W2BEGb[7] ,
    \Tile_X5Y14_W2BEGb[6] ,
    \Tile_X5Y14_W2BEGb[5] ,
    \Tile_X5Y14_W2BEGb[4] ,
    \Tile_X5Y14_W2BEGb[3] ,
    \Tile_X5Y14_W2BEGb[2] ,
    \Tile_X5Y14_W2BEGb[1] ,
    \Tile_X5Y14_W2BEGb[0] }),
    .W2END({\Tile_X6Y14_W2BEGb[7] ,
    \Tile_X6Y14_W2BEGb[6] ,
    \Tile_X6Y14_W2BEGb[5] ,
    \Tile_X6Y14_W2BEGb[4] ,
    \Tile_X6Y14_W2BEGb[3] ,
    \Tile_X6Y14_W2BEGb[2] ,
    \Tile_X6Y14_W2BEGb[1] ,
    \Tile_X6Y14_W2BEGb[0] }),
    .W2MID({\Tile_X6Y14_W2BEG[7] ,
    \Tile_X6Y14_W2BEG[6] ,
    \Tile_X6Y14_W2BEG[5] ,
    \Tile_X6Y14_W2BEG[4] ,
    \Tile_X6Y14_W2BEG[3] ,
    \Tile_X6Y14_W2BEG[2] ,
    \Tile_X6Y14_W2BEG[1] ,
    \Tile_X6Y14_W2BEG[0] }),
    .W6BEG({\Tile_X5Y14_W6BEG[11] ,
    \Tile_X5Y14_W6BEG[10] ,
    \Tile_X5Y14_W6BEG[9] ,
    \Tile_X5Y14_W6BEG[8] ,
    \Tile_X5Y14_W6BEG[7] ,
    \Tile_X5Y14_W6BEG[6] ,
    \Tile_X5Y14_W6BEG[5] ,
    \Tile_X5Y14_W6BEG[4] ,
    \Tile_X5Y14_W6BEG[3] ,
    \Tile_X5Y14_W6BEG[2] ,
    \Tile_X5Y14_W6BEG[1] ,
    \Tile_X5Y14_W6BEG[0] }),
    .W6END({\Tile_X6Y14_W6BEG[11] ,
    \Tile_X6Y14_W6BEG[10] ,
    \Tile_X6Y14_W6BEG[9] ,
    \Tile_X6Y14_W6BEG[8] ,
    \Tile_X6Y14_W6BEG[7] ,
    \Tile_X6Y14_W6BEG[6] ,
    \Tile_X6Y14_W6BEG[5] ,
    \Tile_X6Y14_W6BEG[4] ,
    \Tile_X6Y14_W6BEG[3] ,
    \Tile_X6Y14_W6BEG[2] ,
    \Tile_X6Y14_W6BEG[1] ,
    \Tile_X6Y14_W6BEG[0] }),
    .WW4BEG({\Tile_X5Y14_WW4BEG[15] ,
    \Tile_X5Y14_WW4BEG[14] ,
    \Tile_X5Y14_WW4BEG[13] ,
    \Tile_X5Y14_WW4BEG[12] ,
    \Tile_X5Y14_WW4BEG[11] ,
    \Tile_X5Y14_WW4BEG[10] ,
    \Tile_X5Y14_WW4BEG[9] ,
    \Tile_X5Y14_WW4BEG[8] ,
    \Tile_X5Y14_WW4BEG[7] ,
    \Tile_X5Y14_WW4BEG[6] ,
    \Tile_X5Y14_WW4BEG[5] ,
    \Tile_X5Y14_WW4BEG[4] ,
    \Tile_X5Y14_WW4BEG[3] ,
    \Tile_X5Y14_WW4BEG[2] ,
    \Tile_X5Y14_WW4BEG[1] ,
    \Tile_X5Y14_WW4BEG[0] }),
    .WW4END({\Tile_X6Y14_WW4BEG[15] ,
    \Tile_X6Y14_WW4BEG[14] ,
    \Tile_X6Y14_WW4BEG[13] ,
    \Tile_X6Y14_WW4BEG[12] ,
    \Tile_X6Y14_WW4BEG[11] ,
    \Tile_X6Y14_WW4BEG[10] ,
    \Tile_X6Y14_WW4BEG[9] ,
    \Tile_X6Y14_WW4BEG[8] ,
    \Tile_X6Y14_WW4BEG[7] ,
    \Tile_X6Y14_WW4BEG[6] ,
    \Tile_X6Y14_WW4BEG[5] ,
    \Tile_X6Y14_WW4BEG[4] ,
    \Tile_X6Y14_WW4BEG[3] ,
    \Tile_X6Y14_WW4BEG[2] ,
    \Tile_X6Y14_WW4BEG[1] ,
    \Tile_X6Y14_WW4BEG[0] }));
 S_CPU_IF Tile_X5Y15_S_CPU_IF (.Co(Tile_X5Y15_Co),
    .I_top0(Tile_X5Y15_I_top0),
    .I_top1(Tile_X5Y15_I_top1),
    .I_top10(Tile_X5Y15_I_top10),
    .I_top11(Tile_X5Y15_I_top11),
    .I_top12(Tile_X5Y15_I_top12),
    .I_top13(Tile_X5Y15_I_top13),
    .I_top14(Tile_X5Y15_I_top14),
    .I_top15(Tile_X5Y15_I_top15),
    .I_top2(Tile_X5Y15_I_top2),
    .I_top3(Tile_X5Y15_I_top3),
    .I_top4(Tile_X5Y15_I_top4),
    .I_top5(Tile_X5Y15_I_top5),
    .I_top6(Tile_X5Y15_I_top6),
    .I_top7(Tile_X5Y15_I_top7),
    .I_top8(Tile_X5Y15_I_top8),
    .I_top9(Tile_X5Y15_I_top9),
    .O_top0(Tile_X5Y15_O_top0),
    .O_top1(Tile_X5Y15_O_top1),
    .O_top10(Tile_X5Y15_O_top10),
    .O_top11(Tile_X5Y15_O_top11),
    .O_top12(Tile_X5Y15_O_top12),
    .O_top13(Tile_X5Y15_O_top13),
    .O_top14(Tile_X5Y15_O_top14),
    .O_top15(Tile_X5Y15_O_top15),
    .O_top2(Tile_X5Y15_O_top2),
    .O_top3(Tile_X5Y15_O_top3),
    .O_top4(Tile_X5Y15_O_top4),
    .O_top5(Tile_X5Y15_O_top5),
    .O_top6(Tile_X5Y15_O_top6),
    .O_top7(Tile_X5Y15_O_top7),
    .O_top8(Tile_X5Y15_O_top8),
    .O_top9(Tile_X5Y15_O_top9),
    .UserCLK(UserCLK),
    .UserCLKo(Tile_X5Y15_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .FrameData({\Tile_X4Y15_FrameData_O[31] ,
    \Tile_X4Y15_FrameData_O[30] ,
    \Tile_X4Y15_FrameData_O[29] ,
    \Tile_X4Y15_FrameData_O[28] ,
    \Tile_X4Y15_FrameData_O[27] ,
    \Tile_X4Y15_FrameData_O[26] ,
    \Tile_X4Y15_FrameData_O[25] ,
    \Tile_X4Y15_FrameData_O[24] ,
    \Tile_X4Y15_FrameData_O[23] ,
    \Tile_X4Y15_FrameData_O[22] ,
    \Tile_X4Y15_FrameData_O[21] ,
    \Tile_X4Y15_FrameData_O[20] ,
    \Tile_X4Y15_FrameData_O[19] ,
    \Tile_X4Y15_FrameData_O[18] ,
    \Tile_X4Y15_FrameData_O[17] ,
    \Tile_X4Y15_FrameData_O[16] ,
    \Tile_X4Y15_FrameData_O[15] ,
    \Tile_X4Y15_FrameData_O[14] ,
    \Tile_X4Y15_FrameData_O[13] ,
    \Tile_X4Y15_FrameData_O[12] ,
    \Tile_X4Y15_FrameData_O[11] ,
    \Tile_X4Y15_FrameData_O[10] ,
    \Tile_X4Y15_FrameData_O[9] ,
    \Tile_X4Y15_FrameData_O[8] ,
    \Tile_X4Y15_FrameData_O[7] ,
    \Tile_X4Y15_FrameData_O[6] ,
    \Tile_X4Y15_FrameData_O[5] ,
    \Tile_X4Y15_FrameData_O[4] ,
    \Tile_X4Y15_FrameData_O[3] ,
    \Tile_X4Y15_FrameData_O[2] ,
    \Tile_X4Y15_FrameData_O[1] ,
    \Tile_X4Y15_FrameData_O[0] }),
    .FrameData_O({\Tile_X5Y15_FrameData_O[31] ,
    \Tile_X5Y15_FrameData_O[30] ,
    \Tile_X5Y15_FrameData_O[29] ,
    \Tile_X5Y15_FrameData_O[28] ,
    \Tile_X5Y15_FrameData_O[27] ,
    \Tile_X5Y15_FrameData_O[26] ,
    \Tile_X5Y15_FrameData_O[25] ,
    \Tile_X5Y15_FrameData_O[24] ,
    \Tile_X5Y15_FrameData_O[23] ,
    \Tile_X5Y15_FrameData_O[22] ,
    \Tile_X5Y15_FrameData_O[21] ,
    \Tile_X5Y15_FrameData_O[20] ,
    \Tile_X5Y15_FrameData_O[19] ,
    \Tile_X5Y15_FrameData_O[18] ,
    \Tile_X5Y15_FrameData_O[17] ,
    \Tile_X5Y15_FrameData_O[16] ,
    \Tile_X5Y15_FrameData_O[15] ,
    \Tile_X5Y15_FrameData_O[14] ,
    \Tile_X5Y15_FrameData_O[13] ,
    \Tile_X5Y15_FrameData_O[12] ,
    \Tile_X5Y15_FrameData_O[11] ,
    \Tile_X5Y15_FrameData_O[10] ,
    \Tile_X5Y15_FrameData_O[9] ,
    \Tile_X5Y15_FrameData_O[8] ,
    \Tile_X5Y15_FrameData_O[7] ,
    \Tile_X5Y15_FrameData_O[6] ,
    \Tile_X5Y15_FrameData_O[5] ,
    \Tile_X5Y15_FrameData_O[4] ,
    \Tile_X5Y15_FrameData_O[3] ,
    \Tile_X5Y15_FrameData_O[2] ,
    \Tile_X5Y15_FrameData_O[1] ,
    \Tile_X5Y15_FrameData_O[0] }),
    .FrameStrobe({FrameStrobe[119],
    FrameStrobe[118],
    FrameStrobe[117],
    FrameStrobe[116],
    FrameStrobe[115],
    FrameStrobe[114],
    FrameStrobe[113],
    FrameStrobe[112],
    FrameStrobe[111],
    FrameStrobe[110],
    FrameStrobe[109],
    FrameStrobe[108],
    FrameStrobe[107],
    FrameStrobe[106],
    FrameStrobe[105],
    FrameStrobe[104],
    FrameStrobe[103],
    FrameStrobe[102],
    FrameStrobe[101],
    FrameStrobe[100]}),
    .FrameStrobe_O({\Tile_X5Y15_FrameStrobe_O[19] ,
    \Tile_X5Y15_FrameStrobe_O[18] ,
    \Tile_X5Y15_FrameStrobe_O[17] ,
    \Tile_X5Y15_FrameStrobe_O[16] ,
    \Tile_X5Y15_FrameStrobe_O[15] ,
    \Tile_X5Y15_FrameStrobe_O[14] ,
    \Tile_X5Y15_FrameStrobe_O[13] ,
    \Tile_X5Y15_FrameStrobe_O[12] ,
    \Tile_X5Y15_FrameStrobe_O[11] ,
    \Tile_X5Y15_FrameStrobe_O[10] ,
    \Tile_X5Y15_FrameStrobe_O[9] ,
    \Tile_X5Y15_FrameStrobe_O[8] ,
    \Tile_X5Y15_FrameStrobe_O[7] ,
    \Tile_X5Y15_FrameStrobe_O[6] ,
    \Tile_X5Y15_FrameStrobe_O[5] ,
    \Tile_X5Y15_FrameStrobe_O[4] ,
    \Tile_X5Y15_FrameStrobe_O[3] ,
    \Tile_X5Y15_FrameStrobe_O[2] ,
    \Tile_X5Y15_FrameStrobe_O[1] ,
    \Tile_X5Y15_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X5Y15_N1BEG[3] ,
    \Tile_X5Y15_N1BEG[2] ,
    \Tile_X5Y15_N1BEG[1] ,
    \Tile_X5Y15_N1BEG[0] }),
    .N2BEG({\Tile_X5Y15_N2BEG[7] ,
    \Tile_X5Y15_N2BEG[6] ,
    \Tile_X5Y15_N2BEG[5] ,
    \Tile_X5Y15_N2BEG[4] ,
    \Tile_X5Y15_N2BEG[3] ,
    \Tile_X5Y15_N2BEG[2] ,
    \Tile_X5Y15_N2BEG[1] ,
    \Tile_X5Y15_N2BEG[0] }),
    .N2BEGb({\Tile_X5Y15_N2BEGb[7] ,
    \Tile_X5Y15_N2BEGb[6] ,
    \Tile_X5Y15_N2BEGb[5] ,
    \Tile_X5Y15_N2BEGb[4] ,
    \Tile_X5Y15_N2BEGb[3] ,
    \Tile_X5Y15_N2BEGb[2] ,
    \Tile_X5Y15_N2BEGb[1] ,
    \Tile_X5Y15_N2BEGb[0] }),
    .N4BEG({\Tile_X5Y15_N4BEG[15] ,
    \Tile_X5Y15_N4BEG[14] ,
    \Tile_X5Y15_N4BEG[13] ,
    \Tile_X5Y15_N4BEG[12] ,
    \Tile_X5Y15_N4BEG[11] ,
    \Tile_X5Y15_N4BEG[10] ,
    \Tile_X5Y15_N4BEG[9] ,
    \Tile_X5Y15_N4BEG[8] ,
    \Tile_X5Y15_N4BEG[7] ,
    \Tile_X5Y15_N4BEG[6] ,
    \Tile_X5Y15_N4BEG[5] ,
    \Tile_X5Y15_N4BEG[4] ,
    \Tile_X5Y15_N4BEG[3] ,
    \Tile_X5Y15_N4BEG[2] ,
    \Tile_X5Y15_N4BEG[1] ,
    \Tile_X5Y15_N4BEG[0] }),
    .NN4BEG({\Tile_X5Y15_NN4BEG[15] ,
    \Tile_X5Y15_NN4BEG[14] ,
    \Tile_X5Y15_NN4BEG[13] ,
    \Tile_X5Y15_NN4BEG[12] ,
    \Tile_X5Y15_NN4BEG[11] ,
    \Tile_X5Y15_NN4BEG[10] ,
    \Tile_X5Y15_NN4BEG[9] ,
    \Tile_X5Y15_NN4BEG[8] ,
    \Tile_X5Y15_NN4BEG[7] ,
    \Tile_X5Y15_NN4BEG[6] ,
    \Tile_X5Y15_NN4BEG[5] ,
    \Tile_X5Y15_NN4BEG[4] ,
    \Tile_X5Y15_NN4BEG[3] ,
    \Tile_X5Y15_NN4BEG[2] ,
    \Tile_X5Y15_NN4BEG[1] ,
    \Tile_X5Y15_NN4BEG[0] }),
    .S1END({\Tile_X5Y14_S1BEG[3] ,
    \Tile_X5Y14_S1BEG[2] ,
    \Tile_X5Y14_S1BEG[1] ,
    \Tile_X5Y14_S1BEG[0] }),
    .S2END({\Tile_X5Y14_S2BEGb[7] ,
    \Tile_X5Y14_S2BEGb[6] ,
    \Tile_X5Y14_S2BEGb[5] ,
    \Tile_X5Y14_S2BEGb[4] ,
    \Tile_X5Y14_S2BEGb[3] ,
    \Tile_X5Y14_S2BEGb[2] ,
    \Tile_X5Y14_S2BEGb[1] ,
    \Tile_X5Y14_S2BEGb[0] }),
    .S2MID({\Tile_X5Y14_S2BEG[7] ,
    \Tile_X5Y14_S2BEG[6] ,
    \Tile_X5Y14_S2BEG[5] ,
    \Tile_X5Y14_S2BEG[4] ,
    \Tile_X5Y14_S2BEG[3] ,
    \Tile_X5Y14_S2BEG[2] ,
    \Tile_X5Y14_S2BEG[1] ,
    \Tile_X5Y14_S2BEG[0] }),
    .S4END({\Tile_X5Y14_S4BEG[15] ,
    \Tile_X5Y14_S4BEG[14] ,
    \Tile_X5Y14_S4BEG[13] ,
    \Tile_X5Y14_S4BEG[12] ,
    \Tile_X5Y14_S4BEG[11] ,
    \Tile_X5Y14_S4BEG[10] ,
    \Tile_X5Y14_S4BEG[9] ,
    \Tile_X5Y14_S4BEG[8] ,
    \Tile_X5Y14_S4BEG[7] ,
    \Tile_X5Y14_S4BEG[6] ,
    \Tile_X5Y14_S4BEG[5] ,
    \Tile_X5Y14_S4BEG[4] ,
    \Tile_X5Y14_S4BEG[3] ,
    \Tile_X5Y14_S4BEG[2] ,
    \Tile_X5Y14_S4BEG[1] ,
    \Tile_X5Y14_S4BEG[0] }),
    .SS4END({\Tile_X5Y14_SS4BEG[15] ,
    \Tile_X5Y14_SS4BEG[14] ,
    \Tile_X5Y14_SS4BEG[13] ,
    \Tile_X5Y14_SS4BEG[12] ,
    \Tile_X5Y14_SS4BEG[11] ,
    \Tile_X5Y14_SS4BEG[10] ,
    \Tile_X5Y14_SS4BEG[9] ,
    \Tile_X5Y14_SS4BEG[8] ,
    \Tile_X5Y14_SS4BEG[7] ,
    \Tile_X5Y14_SS4BEG[6] ,
    \Tile_X5Y14_SS4BEG[5] ,
    \Tile_X5Y14_SS4BEG[4] ,
    \Tile_X5Y14_SS4BEG[3] ,
    \Tile_X5Y14_SS4BEG[2] ,
    \Tile_X5Y14_SS4BEG[1] ,
    \Tile_X5Y14_SS4BEG[0] }));
 LUT4AB Tile_X5Y1_LUT4AB (.Ci(Tile_X5Y2_Co),
    .Co(Tile_X5Y1_Co),
    .UserCLK(Tile_X5Y2_UserCLKo),
    .UserCLKo(Tile_X5Y1_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X5Y1_E1BEG[3] ,
    \Tile_X5Y1_E1BEG[2] ,
    \Tile_X5Y1_E1BEG[1] ,
    \Tile_X5Y1_E1BEG[0] }),
    .E1END({\Tile_X4Y1_E1BEG[3] ,
    \Tile_X4Y1_E1BEG[2] ,
    \Tile_X4Y1_E1BEG[1] ,
    \Tile_X4Y1_E1BEG[0] }),
    .E2BEG({\Tile_X5Y1_E2BEG[7] ,
    \Tile_X5Y1_E2BEG[6] ,
    \Tile_X5Y1_E2BEG[5] ,
    \Tile_X5Y1_E2BEG[4] ,
    \Tile_X5Y1_E2BEG[3] ,
    \Tile_X5Y1_E2BEG[2] ,
    \Tile_X5Y1_E2BEG[1] ,
    \Tile_X5Y1_E2BEG[0] }),
    .E2BEGb({\Tile_X5Y1_E2BEGb[7] ,
    \Tile_X5Y1_E2BEGb[6] ,
    \Tile_X5Y1_E2BEGb[5] ,
    \Tile_X5Y1_E2BEGb[4] ,
    \Tile_X5Y1_E2BEGb[3] ,
    \Tile_X5Y1_E2BEGb[2] ,
    \Tile_X5Y1_E2BEGb[1] ,
    \Tile_X5Y1_E2BEGb[0] }),
    .E2END({\Tile_X4Y1_E2BEGb[7] ,
    \Tile_X4Y1_E2BEGb[6] ,
    \Tile_X4Y1_E2BEGb[5] ,
    \Tile_X4Y1_E2BEGb[4] ,
    \Tile_X4Y1_E2BEGb[3] ,
    \Tile_X4Y1_E2BEGb[2] ,
    \Tile_X4Y1_E2BEGb[1] ,
    \Tile_X4Y1_E2BEGb[0] }),
    .E2MID({\Tile_X4Y1_E2BEG[7] ,
    \Tile_X4Y1_E2BEG[6] ,
    \Tile_X4Y1_E2BEG[5] ,
    \Tile_X4Y1_E2BEG[4] ,
    \Tile_X4Y1_E2BEG[3] ,
    \Tile_X4Y1_E2BEG[2] ,
    \Tile_X4Y1_E2BEG[1] ,
    \Tile_X4Y1_E2BEG[0] }),
    .E6BEG({\Tile_X5Y1_E6BEG[11] ,
    \Tile_X5Y1_E6BEG[10] ,
    \Tile_X5Y1_E6BEG[9] ,
    \Tile_X5Y1_E6BEG[8] ,
    \Tile_X5Y1_E6BEG[7] ,
    \Tile_X5Y1_E6BEG[6] ,
    \Tile_X5Y1_E6BEG[5] ,
    \Tile_X5Y1_E6BEG[4] ,
    \Tile_X5Y1_E6BEG[3] ,
    \Tile_X5Y1_E6BEG[2] ,
    \Tile_X5Y1_E6BEG[1] ,
    \Tile_X5Y1_E6BEG[0] }),
    .E6END({\Tile_X4Y1_E6BEG[11] ,
    \Tile_X4Y1_E6BEG[10] ,
    \Tile_X4Y1_E6BEG[9] ,
    \Tile_X4Y1_E6BEG[8] ,
    \Tile_X4Y1_E6BEG[7] ,
    \Tile_X4Y1_E6BEG[6] ,
    \Tile_X4Y1_E6BEG[5] ,
    \Tile_X4Y1_E6BEG[4] ,
    \Tile_X4Y1_E6BEG[3] ,
    \Tile_X4Y1_E6BEG[2] ,
    \Tile_X4Y1_E6BEG[1] ,
    \Tile_X4Y1_E6BEG[0] }),
    .EE4BEG({\Tile_X5Y1_EE4BEG[15] ,
    \Tile_X5Y1_EE4BEG[14] ,
    \Tile_X5Y1_EE4BEG[13] ,
    \Tile_X5Y1_EE4BEG[12] ,
    \Tile_X5Y1_EE4BEG[11] ,
    \Tile_X5Y1_EE4BEG[10] ,
    \Tile_X5Y1_EE4BEG[9] ,
    \Tile_X5Y1_EE4BEG[8] ,
    \Tile_X5Y1_EE4BEG[7] ,
    \Tile_X5Y1_EE4BEG[6] ,
    \Tile_X5Y1_EE4BEG[5] ,
    \Tile_X5Y1_EE4BEG[4] ,
    \Tile_X5Y1_EE4BEG[3] ,
    \Tile_X5Y1_EE4BEG[2] ,
    \Tile_X5Y1_EE4BEG[1] ,
    \Tile_X5Y1_EE4BEG[0] }),
    .EE4END({\Tile_X4Y1_EE4BEG[15] ,
    \Tile_X4Y1_EE4BEG[14] ,
    \Tile_X4Y1_EE4BEG[13] ,
    \Tile_X4Y1_EE4BEG[12] ,
    \Tile_X4Y1_EE4BEG[11] ,
    \Tile_X4Y1_EE4BEG[10] ,
    \Tile_X4Y1_EE4BEG[9] ,
    \Tile_X4Y1_EE4BEG[8] ,
    \Tile_X4Y1_EE4BEG[7] ,
    \Tile_X4Y1_EE4BEG[6] ,
    \Tile_X4Y1_EE4BEG[5] ,
    \Tile_X4Y1_EE4BEG[4] ,
    \Tile_X4Y1_EE4BEG[3] ,
    \Tile_X4Y1_EE4BEG[2] ,
    \Tile_X4Y1_EE4BEG[1] ,
    \Tile_X4Y1_EE4BEG[0] }),
    .FrameData({\Tile_X4Y1_FrameData_O[31] ,
    \Tile_X4Y1_FrameData_O[30] ,
    \Tile_X4Y1_FrameData_O[29] ,
    \Tile_X4Y1_FrameData_O[28] ,
    \Tile_X4Y1_FrameData_O[27] ,
    \Tile_X4Y1_FrameData_O[26] ,
    \Tile_X4Y1_FrameData_O[25] ,
    \Tile_X4Y1_FrameData_O[24] ,
    \Tile_X4Y1_FrameData_O[23] ,
    \Tile_X4Y1_FrameData_O[22] ,
    \Tile_X4Y1_FrameData_O[21] ,
    \Tile_X4Y1_FrameData_O[20] ,
    \Tile_X4Y1_FrameData_O[19] ,
    \Tile_X4Y1_FrameData_O[18] ,
    \Tile_X4Y1_FrameData_O[17] ,
    \Tile_X4Y1_FrameData_O[16] ,
    \Tile_X4Y1_FrameData_O[15] ,
    \Tile_X4Y1_FrameData_O[14] ,
    \Tile_X4Y1_FrameData_O[13] ,
    \Tile_X4Y1_FrameData_O[12] ,
    \Tile_X4Y1_FrameData_O[11] ,
    \Tile_X4Y1_FrameData_O[10] ,
    \Tile_X4Y1_FrameData_O[9] ,
    \Tile_X4Y1_FrameData_O[8] ,
    \Tile_X4Y1_FrameData_O[7] ,
    \Tile_X4Y1_FrameData_O[6] ,
    \Tile_X4Y1_FrameData_O[5] ,
    \Tile_X4Y1_FrameData_O[4] ,
    \Tile_X4Y1_FrameData_O[3] ,
    \Tile_X4Y1_FrameData_O[2] ,
    \Tile_X4Y1_FrameData_O[1] ,
    \Tile_X4Y1_FrameData_O[0] }),
    .FrameData_O({\Tile_X5Y1_FrameData_O[31] ,
    \Tile_X5Y1_FrameData_O[30] ,
    \Tile_X5Y1_FrameData_O[29] ,
    \Tile_X5Y1_FrameData_O[28] ,
    \Tile_X5Y1_FrameData_O[27] ,
    \Tile_X5Y1_FrameData_O[26] ,
    \Tile_X5Y1_FrameData_O[25] ,
    \Tile_X5Y1_FrameData_O[24] ,
    \Tile_X5Y1_FrameData_O[23] ,
    \Tile_X5Y1_FrameData_O[22] ,
    \Tile_X5Y1_FrameData_O[21] ,
    \Tile_X5Y1_FrameData_O[20] ,
    \Tile_X5Y1_FrameData_O[19] ,
    \Tile_X5Y1_FrameData_O[18] ,
    \Tile_X5Y1_FrameData_O[17] ,
    \Tile_X5Y1_FrameData_O[16] ,
    \Tile_X5Y1_FrameData_O[15] ,
    \Tile_X5Y1_FrameData_O[14] ,
    \Tile_X5Y1_FrameData_O[13] ,
    \Tile_X5Y1_FrameData_O[12] ,
    \Tile_X5Y1_FrameData_O[11] ,
    \Tile_X5Y1_FrameData_O[10] ,
    \Tile_X5Y1_FrameData_O[9] ,
    \Tile_X5Y1_FrameData_O[8] ,
    \Tile_X5Y1_FrameData_O[7] ,
    \Tile_X5Y1_FrameData_O[6] ,
    \Tile_X5Y1_FrameData_O[5] ,
    \Tile_X5Y1_FrameData_O[4] ,
    \Tile_X5Y1_FrameData_O[3] ,
    \Tile_X5Y1_FrameData_O[2] ,
    \Tile_X5Y1_FrameData_O[1] ,
    \Tile_X5Y1_FrameData_O[0] }),
    .FrameStrobe({\Tile_X5Y2_FrameStrobe_O[19] ,
    \Tile_X5Y2_FrameStrobe_O[18] ,
    \Tile_X5Y2_FrameStrobe_O[17] ,
    \Tile_X5Y2_FrameStrobe_O[16] ,
    \Tile_X5Y2_FrameStrobe_O[15] ,
    \Tile_X5Y2_FrameStrobe_O[14] ,
    \Tile_X5Y2_FrameStrobe_O[13] ,
    \Tile_X5Y2_FrameStrobe_O[12] ,
    \Tile_X5Y2_FrameStrobe_O[11] ,
    \Tile_X5Y2_FrameStrobe_O[10] ,
    \Tile_X5Y2_FrameStrobe_O[9] ,
    \Tile_X5Y2_FrameStrobe_O[8] ,
    \Tile_X5Y2_FrameStrobe_O[7] ,
    \Tile_X5Y2_FrameStrobe_O[6] ,
    \Tile_X5Y2_FrameStrobe_O[5] ,
    \Tile_X5Y2_FrameStrobe_O[4] ,
    \Tile_X5Y2_FrameStrobe_O[3] ,
    \Tile_X5Y2_FrameStrobe_O[2] ,
    \Tile_X5Y2_FrameStrobe_O[1] ,
    \Tile_X5Y2_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X5Y1_FrameStrobe_O[19] ,
    \Tile_X5Y1_FrameStrobe_O[18] ,
    \Tile_X5Y1_FrameStrobe_O[17] ,
    \Tile_X5Y1_FrameStrobe_O[16] ,
    \Tile_X5Y1_FrameStrobe_O[15] ,
    \Tile_X5Y1_FrameStrobe_O[14] ,
    \Tile_X5Y1_FrameStrobe_O[13] ,
    \Tile_X5Y1_FrameStrobe_O[12] ,
    \Tile_X5Y1_FrameStrobe_O[11] ,
    \Tile_X5Y1_FrameStrobe_O[10] ,
    \Tile_X5Y1_FrameStrobe_O[9] ,
    \Tile_X5Y1_FrameStrobe_O[8] ,
    \Tile_X5Y1_FrameStrobe_O[7] ,
    \Tile_X5Y1_FrameStrobe_O[6] ,
    \Tile_X5Y1_FrameStrobe_O[5] ,
    \Tile_X5Y1_FrameStrobe_O[4] ,
    \Tile_X5Y1_FrameStrobe_O[3] ,
    \Tile_X5Y1_FrameStrobe_O[2] ,
    \Tile_X5Y1_FrameStrobe_O[1] ,
    \Tile_X5Y1_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X5Y1_N1BEG[3] ,
    \Tile_X5Y1_N1BEG[2] ,
    \Tile_X5Y1_N1BEG[1] ,
    \Tile_X5Y1_N1BEG[0] }),
    .N1END({\Tile_X5Y2_N1BEG[3] ,
    \Tile_X5Y2_N1BEG[2] ,
    \Tile_X5Y2_N1BEG[1] ,
    \Tile_X5Y2_N1BEG[0] }),
    .N2BEG({\Tile_X5Y1_N2BEG[7] ,
    \Tile_X5Y1_N2BEG[6] ,
    \Tile_X5Y1_N2BEG[5] ,
    \Tile_X5Y1_N2BEG[4] ,
    \Tile_X5Y1_N2BEG[3] ,
    \Tile_X5Y1_N2BEG[2] ,
    \Tile_X5Y1_N2BEG[1] ,
    \Tile_X5Y1_N2BEG[0] }),
    .N2BEGb({\Tile_X5Y1_N2BEGb[7] ,
    \Tile_X5Y1_N2BEGb[6] ,
    \Tile_X5Y1_N2BEGb[5] ,
    \Tile_X5Y1_N2BEGb[4] ,
    \Tile_X5Y1_N2BEGb[3] ,
    \Tile_X5Y1_N2BEGb[2] ,
    \Tile_X5Y1_N2BEGb[1] ,
    \Tile_X5Y1_N2BEGb[0] }),
    .N2END({\Tile_X5Y2_N2BEGb[7] ,
    \Tile_X5Y2_N2BEGb[6] ,
    \Tile_X5Y2_N2BEGb[5] ,
    \Tile_X5Y2_N2BEGb[4] ,
    \Tile_X5Y2_N2BEGb[3] ,
    \Tile_X5Y2_N2BEGb[2] ,
    \Tile_X5Y2_N2BEGb[1] ,
    \Tile_X5Y2_N2BEGb[0] }),
    .N2MID({\Tile_X5Y2_N2BEG[7] ,
    \Tile_X5Y2_N2BEG[6] ,
    \Tile_X5Y2_N2BEG[5] ,
    \Tile_X5Y2_N2BEG[4] ,
    \Tile_X5Y2_N2BEG[3] ,
    \Tile_X5Y2_N2BEG[2] ,
    \Tile_X5Y2_N2BEG[1] ,
    \Tile_X5Y2_N2BEG[0] }),
    .N4BEG({\Tile_X5Y1_N4BEG[15] ,
    \Tile_X5Y1_N4BEG[14] ,
    \Tile_X5Y1_N4BEG[13] ,
    \Tile_X5Y1_N4BEG[12] ,
    \Tile_X5Y1_N4BEG[11] ,
    \Tile_X5Y1_N4BEG[10] ,
    \Tile_X5Y1_N4BEG[9] ,
    \Tile_X5Y1_N4BEG[8] ,
    \Tile_X5Y1_N4BEG[7] ,
    \Tile_X5Y1_N4BEG[6] ,
    \Tile_X5Y1_N4BEG[5] ,
    \Tile_X5Y1_N4BEG[4] ,
    \Tile_X5Y1_N4BEG[3] ,
    \Tile_X5Y1_N4BEG[2] ,
    \Tile_X5Y1_N4BEG[1] ,
    \Tile_X5Y1_N4BEG[0] }),
    .N4END({\Tile_X5Y2_N4BEG[15] ,
    \Tile_X5Y2_N4BEG[14] ,
    \Tile_X5Y2_N4BEG[13] ,
    \Tile_X5Y2_N4BEG[12] ,
    \Tile_X5Y2_N4BEG[11] ,
    \Tile_X5Y2_N4BEG[10] ,
    \Tile_X5Y2_N4BEG[9] ,
    \Tile_X5Y2_N4BEG[8] ,
    \Tile_X5Y2_N4BEG[7] ,
    \Tile_X5Y2_N4BEG[6] ,
    \Tile_X5Y2_N4BEG[5] ,
    \Tile_X5Y2_N4BEG[4] ,
    \Tile_X5Y2_N4BEG[3] ,
    \Tile_X5Y2_N4BEG[2] ,
    \Tile_X5Y2_N4BEG[1] ,
    \Tile_X5Y2_N4BEG[0] }),
    .NN4BEG({\Tile_X5Y1_NN4BEG[15] ,
    \Tile_X5Y1_NN4BEG[14] ,
    \Tile_X5Y1_NN4BEG[13] ,
    \Tile_X5Y1_NN4BEG[12] ,
    \Tile_X5Y1_NN4BEG[11] ,
    \Tile_X5Y1_NN4BEG[10] ,
    \Tile_X5Y1_NN4BEG[9] ,
    \Tile_X5Y1_NN4BEG[8] ,
    \Tile_X5Y1_NN4BEG[7] ,
    \Tile_X5Y1_NN4BEG[6] ,
    \Tile_X5Y1_NN4BEG[5] ,
    \Tile_X5Y1_NN4BEG[4] ,
    \Tile_X5Y1_NN4BEG[3] ,
    \Tile_X5Y1_NN4BEG[2] ,
    \Tile_X5Y1_NN4BEG[1] ,
    \Tile_X5Y1_NN4BEG[0] }),
    .NN4END({\Tile_X5Y2_NN4BEG[15] ,
    \Tile_X5Y2_NN4BEG[14] ,
    \Tile_X5Y2_NN4BEG[13] ,
    \Tile_X5Y2_NN4BEG[12] ,
    \Tile_X5Y2_NN4BEG[11] ,
    \Tile_X5Y2_NN4BEG[10] ,
    \Tile_X5Y2_NN4BEG[9] ,
    \Tile_X5Y2_NN4BEG[8] ,
    \Tile_X5Y2_NN4BEG[7] ,
    \Tile_X5Y2_NN4BEG[6] ,
    \Tile_X5Y2_NN4BEG[5] ,
    \Tile_X5Y2_NN4BEG[4] ,
    \Tile_X5Y2_NN4BEG[3] ,
    \Tile_X5Y2_NN4BEG[2] ,
    \Tile_X5Y2_NN4BEG[1] ,
    \Tile_X5Y2_NN4BEG[0] }),
    .S1BEG({\Tile_X5Y1_S1BEG[3] ,
    \Tile_X5Y1_S1BEG[2] ,
    \Tile_X5Y1_S1BEG[1] ,
    \Tile_X5Y1_S1BEG[0] }),
    .S1END({\Tile_X5Y0_S1BEG[3] ,
    \Tile_X5Y0_S1BEG[2] ,
    \Tile_X5Y0_S1BEG[1] ,
    \Tile_X5Y0_S1BEG[0] }),
    .S2BEG({\Tile_X5Y1_S2BEG[7] ,
    \Tile_X5Y1_S2BEG[6] ,
    \Tile_X5Y1_S2BEG[5] ,
    \Tile_X5Y1_S2BEG[4] ,
    \Tile_X5Y1_S2BEG[3] ,
    \Tile_X5Y1_S2BEG[2] ,
    \Tile_X5Y1_S2BEG[1] ,
    \Tile_X5Y1_S2BEG[0] }),
    .S2BEGb({\Tile_X5Y1_S2BEGb[7] ,
    \Tile_X5Y1_S2BEGb[6] ,
    \Tile_X5Y1_S2BEGb[5] ,
    \Tile_X5Y1_S2BEGb[4] ,
    \Tile_X5Y1_S2BEGb[3] ,
    \Tile_X5Y1_S2BEGb[2] ,
    \Tile_X5Y1_S2BEGb[1] ,
    \Tile_X5Y1_S2BEGb[0] }),
    .S2END({\Tile_X5Y0_S2BEGb[7] ,
    \Tile_X5Y0_S2BEGb[6] ,
    \Tile_X5Y0_S2BEGb[5] ,
    \Tile_X5Y0_S2BEGb[4] ,
    \Tile_X5Y0_S2BEGb[3] ,
    \Tile_X5Y0_S2BEGb[2] ,
    \Tile_X5Y0_S2BEGb[1] ,
    \Tile_X5Y0_S2BEGb[0] }),
    .S2MID({\Tile_X5Y0_S2BEG[7] ,
    \Tile_X5Y0_S2BEG[6] ,
    \Tile_X5Y0_S2BEG[5] ,
    \Tile_X5Y0_S2BEG[4] ,
    \Tile_X5Y0_S2BEG[3] ,
    \Tile_X5Y0_S2BEG[2] ,
    \Tile_X5Y0_S2BEG[1] ,
    \Tile_X5Y0_S2BEG[0] }),
    .S4BEG({\Tile_X5Y1_S4BEG[15] ,
    \Tile_X5Y1_S4BEG[14] ,
    \Tile_X5Y1_S4BEG[13] ,
    \Tile_X5Y1_S4BEG[12] ,
    \Tile_X5Y1_S4BEG[11] ,
    \Tile_X5Y1_S4BEG[10] ,
    \Tile_X5Y1_S4BEG[9] ,
    \Tile_X5Y1_S4BEG[8] ,
    \Tile_X5Y1_S4BEG[7] ,
    \Tile_X5Y1_S4BEG[6] ,
    \Tile_X5Y1_S4BEG[5] ,
    \Tile_X5Y1_S4BEG[4] ,
    \Tile_X5Y1_S4BEG[3] ,
    \Tile_X5Y1_S4BEG[2] ,
    \Tile_X5Y1_S4BEG[1] ,
    \Tile_X5Y1_S4BEG[0] }),
    .S4END({\Tile_X5Y0_S4BEG[15] ,
    \Tile_X5Y0_S4BEG[14] ,
    \Tile_X5Y0_S4BEG[13] ,
    \Tile_X5Y0_S4BEG[12] ,
    \Tile_X5Y0_S4BEG[11] ,
    \Tile_X5Y0_S4BEG[10] ,
    \Tile_X5Y0_S4BEG[9] ,
    \Tile_X5Y0_S4BEG[8] ,
    \Tile_X5Y0_S4BEG[7] ,
    \Tile_X5Y0_S4BEG[6] ,
    \Tile_X5Y0_S4BEG[5] ,
    \Tile_X5Y0_S4BEG[4] ,
    \Tile_X5Y0_S4BEG[3] ,
    \Tile_X5Y0_S4BEG[2] ,
    \Tile_X5Y0_S4BEG[1] ,
    \Tile_X5Y0_S4BEG[0] }),
    .SS4BEG({\Tile_X5Y1_SS4BEG[15] ,
    \Tile_X5Y1_SS4BEG[14] ,
    \Tile_X5Y1_SS4BEG[13] ,
    \Tile_X5Y1_SS4BEG[12] ,
    \Tile_X5Y1_SS4BEG[11] ,
    \Tile_X5Y1_SS4BEG[10] ,
    \Tile_X5Y1_SS4BEG[9] ,
    \Tile_X5Y1_SS4BEG[8] ,
    \Tile_X5Y1_SS4BEG[7] ,
    \Tile_X5Y1_SS4BEG[6] ,
    \Tile_X5Y1_SS4BEG[5] ,
    \Tile_X5Y1_SS4BEG[4] ,
    \Tile_X5Y1_SS4BEG[3] ,
    \Tile_X5Y1_SS4BEG[2] ,
    \Tile_X5Y1_SS4BEG[1] ,
    \Tile_X5Y1_SS4BEG[0] }),
    .SS4END({\Tile_X5Y0_SS4BEG[15] ,
    \Tile_X5Y0_SS4BEG[14] ,
    \Tile_X5Y0_SS4BEG[13] ,
    \Tile_X5Y0_SS4BEG[12] ,
    \Tile_X5Y0_SS4BEG[11] ,
    \Tile_X5Y0_SS4BEG[10] ,
    \Tile_X5Y0_SS4BEG[9] ,
    \Tile_X5Y0_SS4BEG[8] ,
    \Tile_X5Y0_SS4BEG[7] ,
    \Tile_X5Y0_SS4BEG[6] ,
    \Tile_X5Y0_SS4BEG[5] ,
    \Tile_X5Y0_SS4BEG[4] ,
    \Tile_X5Y0_SS4BEG[3] ,
    \Tile_X5Y0_SS4BEG[2] ,
    \Tile_X5Y0_SS4BEG[1] ,
    \Tile_X5Y0_SS4BEG[0] }),
    .W1BEG({\Tile_X5Y1_W1BEG[3] ,
    \Tile_X5Y1_W1BEG[2] ,
    \Tile_X5Y1_W1BEG[1] ,
    \Tile_X5Y1_W1BEG[0] }),
    .W1END({\Tile_X6Y1_W1BEG[3] ,
    \Tile_X6Y1_W1BEG[2] ,
    \Tile_X6Y1_W1BEG[1] ,
    \Tile_X6Y1_W1BEG[0] }),
    .W2BEG({\Tile_X5Y1_W2BEG[7] ,
    \Tile_X5Y1_W2BEG[6] ,
    \Tile_X5Y1_W2BEG[5] ,
    \Tile_X5Y1_W2BEG[4] ,
    \Tile_X5Y1_W2BEG[3] ,
    \Tile_X5Y1_W2BEG[2] ,
    \Tile_X5Y1_W2BEG[1] ,
    \Tile_X5Y1_W2BEG[0] }),
    .W2BEGb({\Tile_X5Y1_W2BEGb[7] ,
    \Tile_X5Y1_W2BEGb[6] ,
    \Tile_X5Y1_W2BEGb[5] ,
    \Tile_X5Y1_W2BEGb[4] ,
    \Tile_X5Y1_W2BEGb[3] ,
    \Tile_X5Y1_W2BEGb[2] ,
    \Tile_X5Y1_W2BEGb[1] ,
    \Tile_X5Y1_W2BEGb[0] }),
    .W2END({\Tile_X6Y1_W2BEGb[7] ,
    \Tile_X6Y1_W2BEGb[6] ,
    \Tile_X6Y1_W2BEGb[5] ,
    \Tile_X6Y1_W2BEGb[4] ,
    \Tile_X6Y1_W2BEGb[3] ,
    \Tile_X6Y1_W2BEGb[2] ,
    \Tile_X6Y1_W2BEGb[1] ,
    \Tile_X6Y1_W2BEGb[0] }),
    .W2MID({\Tile_X6Y1_W2BEG[7] ,
    \Tile_X6Y1_W2BEG[6] ,
    \Tile_X6Y1_W2BEG[5] ,
    \Tile_X6Y1_W2BEG[4] ,
    \Tile_X6Y1_W2BEG[3] ,
    \Tile_X6Y1_W2BEG[2] ,
    \Tile_X6Y1_W2BEG[1] ,
    \Tile_X6Y1_W2BEG[0] }),
    .W6BEG({\Tile_X5Y1_W6BEG[11] ,
    \Tile_X5Y1_W6BEG[10] ,
    \Tile_X5Y1_W6BEG[9] ,
    \Tile_X5Y1_W6BEG[8] ,
    \Tile_X5Y1_W6BEG[7] ,
    \Tile_X5Y1_W6BEG[6] ,
    \Tile_X5Y1_W6BEG[5] ,
    \Tile_X5Y1_W6BEG[4] ,
    \Tile_X5Y1_W6BEG[3] ,
    \Tile_X5Y1_W6BEG[2] ,
    \Tile_X5Y1_W6BEG[1] ,
    \Tile_X5Y1_W6BEG[0] }),
    .W6END({\Tile_X6Y1_W6BEG[11] ,
    \Tile_X6Y1_W6BEG[10] ,
    \Tile_X6Y1_W6BEG[9] ,
    \Tile_X6Y1_W6BEG[8] ,
    \Tile_X6Y1_W6BEG[7] ,
    \Tile_X6Y1_W6BEG[6] ,
    \Tile_X6Y1_W6BEG[5] ,
    \Tile_X6Y1_W6BEG[4] ,
    \Tile_X6Y1_W6BEG[3] ,
    \Tile_X6Y1_W6BEG[2] ,
    \Tile_X6Y1_W6BEG[1] ,
    \Tile_X6Y1_W6BEG[0] }),
    .WW4BEG({\Tile_X5Y1_WW4BEG[15] ,
    \Tile_X5Y1_WW4BEG[14] ,
    \Tile_X5Y1_WW4BEG[13] ,
    \Tile_X5Y1_WW4BEG[12] ,
    \Tile_X5Y1_WW4BEG[11] ,
    \Tile_X5Y1_WW4BEG[10] ,
    \Tile_X5Y1_WW4BEG[9] ,
    \Tile_X5Y1_WW4BEG[8] ,
    \Tile_X5Y1_WW4BEG[7] ,
    \Tile_X5Y1_WW4BEG[6] ,
    \Tile_X5Y1_WW4BEG[5] ,
    \Tile_X5Y1_WW4BEG[4] ,
    \Tile_X5Y1_WW4BEG[3] ,
    \Tile_X5Y1_WW4BEG[2] ,
    \Tile_X5Y1_WW4BEG[1] ,
    \Tile_X5Y1_WW4BEG[0] }),
    .WW4END({\Tile_X6Y1_WW4BEG[15] ,
    \Tile_X6Y1_WW4BEG[14] ,
    \Tile_X6Y1_WW4BEG[13] ,
    \Tile_X6Y1_WW4BEG[12] ,
    \Tile_X6Y1_WW4BEG[11] ,
    \Tile_X6Y1_WW4BEG[10] ,
    \Tile_X6Y1_WW4BEG[9] ,
    \Tile_X6Y1_WW4BEG[8] ,
    \Tile_X6Y1_WW4BEG[7] ,
    \Tile_X6Y1_WW4BEG[6] ,
    \Tile_X6Y1_WW4BEG[5] ,
    \Tile_X6Y1_WW4BEG[4] ,
    \Tile_X6Y1_WW4BEG[3] ,
    \Tile_X6Y1_WW4BEG[2] ,
    \Tile_X6Y1_WW4BEG[1] ,
    \Tile_X6Y1_WW4BEG[0] }));
 LUT4AB Tile_X5Y2_LUT4AB (.Ci(Tile_X5Y3_Co),
    .Co(Tile_X5Y2_Co),
    .UserCLK(Tile_X5Y3_UserCLKo),
    .UserCLKo(Tile_X5Y2_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X5Y2_E1BEG[3] ,
    \Tile_X5Y2_E1BEG[2] ,
    \Tile_X5Y2_E1BEG[1] ,
    \Tile_X5Y2_E1BEG[0] }),
    .E1END({\Tile_X4Y2_E1BEG[3] ,
    \Tile_X4Y2_E1BEG[2] ,
    \Tile_X4Y2_E1BEG[1] ,
    \Tile_X4Y2_E1BEG[0] }),
    .E2BEG({\Tile_X5Y2_E2BEG[7] ,
    \Tile_X5Y2_E2BEG[6] ,
    \Tile_X5Y2_E2BEG[5] ,
    \Tile_X5Y2_E2BEG[4] ,
    \Tile_X5Y2_E2BEG[3] ,
    \Tile_X5Y2_E2BEG[2] ,
    \Tile_X5Y2_E2BEG[1] ,
    \Tile_X5Y2_E2BEG[0] }),
    .E2BEGb({\Tile_X5Y2_E2BEGb[7] ,
    \Tile_X5Y2_E2BEGb[6] ,
    \Tile_X5Y2_E2BEGb[5] ,
    \Tile_X5Y2_E2BEGb[4] ,
    \Tile_X5Y2_E2BEGb[3] ,
    \Tile_X5Y2_E2BEGb[2] ,
    \Tile_X5Y2_E2BEGb[1] ,
    \Tile_X5Y2_E2BEGb[0] }),
    .E2END({\Tile_X4Y2_E2BEGb[7] ,
    \Tile_X4Y2_E2BEGb[6] ,
    \Tile_X4Y2_E2BEGb[5] ,
    \Tile_X4Y2_E2BEGb[4] ,
    \Tile_X4Y2_E2BEGb[3] ,
    \Tile_X4Y2_E2BEGb[2] ,
    \Tile_X4Y2_E2BEGb[1] ,
    \Tile_X4Y2_E2BEGb[0] }),
    .E2MID({\Tile_X4Y2_E2BEG[7] ,
    \Tile_X4Y2_E2BEG[6] ,
    \Tile_X4Y2_E2BEG[5] ,
    \Tile_X4Y2_E2BEG[4] ,
    \Tile_X4Y2_E2BEG[3] ,
    \Tile_X4Y2_E2BEG[2] ,
    \Tile_X4Y2_E2BEG[1] ,
    \Tile_X4Y2_E2BEG[0] }),
    .E6BEG({\Tile_X5Y2_E6BEG[11] ,
    \Tile_X5Y2_E6BEG[10] ,
    \Tile_X5Y2_E6BEG[9] ,
    \Tile_X5Y2_E6BEG[8] ,
    \Tile_X5Y2_E6BEG[7] ,
    \Tile_X5Y2_E6BEG[6] ,
    \Tile_X5Y2_E6BEG[5] ,
    \Tile_X5Y2_E6BEG[4] ,
    \Tile_X5Y2_E6BEG[3] ,
    \Tile_X5Y2_E6BEG[2] ,
    \Tile_X5Y2_E6BEG[1] ,
    \Tile_X5Y2_E6BEG[0] }),
    .E6END({\Tile_X4Y2_E6BEG[11] ,
    \Tile_X4Y2_E6BEG[10] ,
    \Tile_X4Y2_E6BEG[9] ,
    \Tile_X4Y2_E6BEG[8] ,
    \Tile_X4Y2_E6BEG[7] ,
    \Tile_X4Y2_E6BEG[6] ,
    \Tile_X4Y2_E6BEG[5] ,
    \Tile_X4Y2_E6BEG[4] ,
    \Tile_X4Y2_E6BEG[3] ,
    \Tile_X4Y2_E6BEG[2] ,
    \Tile_X4Y2_E6BEG[1] ,
    \Tile_X4Y2_E6BEG[0] }),
    .EE4BEG({\Tile_X5Y2_EE4BEG[15] ,
    \Tile_X5Y2_EE4BEG[14] ,
    \Tile_X5Y2_EE4BEG[13] ,
    \Tile_X5Y2_EE4BEG[12] ,
    \Tile_X5Y2_EE4BEG[11] ,
    \Tile_X5Y2_EE4BEG[10] ,
    \Tile_X5Y2_EE4BEG[9] ,
    \Tile_X5Y2_EE4BEG[8] ,
    \Tile_X5Y2_EE4BEG[7] ,
    \Tile_X5Y2_EE4BEG[6] ,
    \Tile_X5Y2_EE4BEG[5] ,
    \Tile_X5Y2_EE4BEG[4] ,
    \Tile_X5Y2_EE4BEG[3] ,
    \Tile_X5Y2_EE4BEG[2] ,
    \Tile_X5Y2_EE4BEG[1] ,
    \Tile_X5Y2_EE4BEG[0] }),
    .EE4END({\Tile_X4Y2_EE4BEG[15] ,
    \Tile_X4Y2_EE4BEG[14] ,
    \Tile_X4Y2_EE4BEG[13] ,
    \Tile_X4Y2_EE4BEG[12] ,
    \Tile_X4Y2_EE4BEG[11] ,
    \Tile_X4Y2_EE4BEG[10] ,
    \Tile_X4Y2_EE4BEG[9] ,
    \Tile_X4Y2_EE4BEG[8] ,
    \Tile_X4Y2_EE4BEG[7] ,
    \Tile_X4Y2_EE4BEG[6] ,
    \Tile_X4Y2_EE4BEG[5] ,
    \Tile_X4Y2_EE4BEG[4] ,
    \Tile_X4Y2_EE4BEG[3] ,
    \Tile_X4Y2_EE4BEG[2] ,
    \Tile_X4Y2_EE4BEG[1] ,
    \Tile_X4Y2_EE4BEG[0] }),
    .FrameData({\Tile_X4Y2_FrameData_O[31] ,
    \Tile_X4Y2_FrameData_O[30] ,
    \Tile_X4Y2_FrameData_O[29] ,
    \Tile_X4Y2_FrameData_O[28] ,
    \Tile_X4Y2_FrameData_O[27] ,
    \Tile_X4Y2_FrameData_O[26] ,
    \Tile_X4Y2_FrameData_O[25] ,
    \Tile_X4Y2_FrameData_O[24] ,
    \Tile_X4Y2_FrameData_O[23] ,
    \Tile_X4Y2_FrameData_O[22] ,
    \Tile_X4Y2_FrameData_O[21] ,
    \Tile_X4Y2_FrameData_O[20] ,
    \Tile_X4Y2_FrameData_O[19] ,
    \Tile_X4Y2_FrameData_O[18] ,
    \Tile_X4Y2_FrameData_O[17] ,
    \Tile_X4Y2_FrameData_O[16] ,
    \Tile_X4Y2_FrameData_O[15] ,
    \Tile_X4Y2_FrameData_O[14] ,
    \Tile_X4Y2_FrameData_O[13] ,
    \Tile_X4Y2_FrameData_O[12] ,
    \Tile_X4Y2_FrameData_O[11] ,
    \Tile_X4Y2_FrameData_O[10] ,
    \Tile_X4Y2_FrameData_O[9] ,
    \Tile_X4Y2_FrameData_O[8] ,
    \Tile_X4Y2_FrameData_O[7] ,
    \Tile_X4Y2_FrameData_O[6] ,
    \Tile_X4Y2_FrameData_O[5] ,
    \Tile_X4Y2_FrameData_O[4] ,
    \Tile_X4Y2_FrameData_O[3] ,
    \Tile_X4Y2_FrameData_O[2] ,
    \Tile_X4Y2_FrameData_O[1] ,
    \Tile_X4Y2_FrameData_O[0] }),
    .FrameData_O({\Tile_X5Y2_FrameData_O[31] ,
    \Tile_X5Y2_FrameData_O[30] ,
    \Tile_X5Y2_FrameData_O[29] ,
    \Tile_X5Y2_FrameData_O[28] ,
    \Tile_X5Y2_FrameData_O[27] ,
    \Tile_X5Y2_FrameData_O[26] ,
    \Tile_X5Y2_FrameData_O[25] ,
    \Tile_X5Y2_FrameData_O[24] ,
    \Tile_X5Y2_FrameData_O[23] ,
    \Tile_X5Y2_FrameData_O[22] ,
    \Tile_X5Y2_FrameData_O[21] ,
    \Tile_X5Y2_FrameData_O[20] ,
    \Tile_X5Y2_FrameData_O[19] ,
    \Tile_X5Y2_FrameData_O[18] ,
    \Tile_X5Y2_FrameData_O[17] ,
    \Tile_X5Y2_FrameData_O[16] ,
    \Tile_X5Y2_FrameData_O[15] ,
    \Tile_X5Y2_FrameData_O[14] ,
    \Tile_X5Y2_FrameData_O[13] ,
    \Tile_X5Y2_FrameData_O[12] ,
    \Tile_X5Y2_FrameData_O[11] ,
    \Tile_X5Y2_FrameData_O[10] ,
    \Tile_X5Y2_FrameData_O[9] ,
    \Tile_X5Y2_FrameData_O[8] ,
    \Tile_X5Y2_FrameData_O[7] ,
    \Tile_X5Y2_FrameData_O[6] ,
    \Tile_X5Y2_FrameData_O[5] ,
    \Tile_X5Y2_FrameData_O[4] ,
    \Tile_X5Y2_FrameData_O[3] ,
    \Tile_X5Y2_FrameData_O[2] ,
    \Tile_X5Y2_FrameData_O[1] ,
    \Tile_X5Y2_FrameData_O[0] }),
    .FrameStrobe({\Tile_X5Y3_FrameStrobe_O[19] ,
    \Tile_X5Y3_FrameStrobe_O[18] ,
    \Tile_X5Y3_FrameStrobe_O[17] ,
    \Tile_X5Y3_FrameStrobe_O[16] ,
    \Tile_X5Y3_FrameStrobe_O[15] ,
    \Tile_X5Y3_FrameStrobe_O[14] ,
    \Tile_X5Y3_FrameStrobe_O[13] ,
    \Tile_X5Y3_FrameStrobe_O[12] ,
    \Tile_X5Y3_FrameStrobe_O[11] ,
    \Tile_X5Y3_FrameStrobe_O[10] ,
    \Tile_X5Y3_FrameStrobe_O[9] ,
    \Tile_X5Y3_FrameStrobe_O[8] ,
    \Tile_X5Y3_FrameStrobe_O[7] ,
    \Tile_X5Y3_FrameStrobe_O[6] ,
    \Tile_X5Y3_FrameStrobe_O[5] ,
    \Tile_X5Y3_FrameStrobe_O[4] ,
    \Tile_X5Y3_FrameStrobe_O[3] ,
    \Tile_X5Y3_FrameStrobe_O[2] ,
    \Tile_X5Y3_FrameStrobe_O[1] ,
    \Tile_X5Y3_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X5Y2_FrameStrobe_O[19] ,
    \Tile_X5Y2_FrameStrobe_O[18] ,
    \Tile_X5Y2_FrameStrobe_O[17] ,
    \Tile_X5Y2_FrameStrobe_O[16] ,
    \Tile_X5Y2_FrameStrobe_O[15] ,
    \Tile_X5Y2_FrameStrobe_O[14] ,
    \Tile_X5Y2_FrameStrobe_O[13] ,
    \Tile_X5Y2_FrameStrobe_O[12] ,
    \Tile_X5Y2_FrameStrobe_O[11] ,
    \Tile_X5Y2_FrameStrobe_O[10] ,
    \Tile_X5Y2_FrameStrobe_O[9] ,
    \Tile_X5Y2_FrameStrobe_O[8] ,
    \Tile_X5Y2_FrameStrobe_O[7] ,
    \Tile_X5Y2_FrameStrobe_O[6] ,
    \Tile_X5Y2_FrameStrobe_O[5] ,
    \Tile_X5Y2_FrameStrobe_O[4] ,
    \Tile_X5Y2_FrameStrobe_O[3] ,
    \Tile_X5Y2_FrameStrobe_O[2] ,
    \Tile_X5Y2_FrameStrobe_O[1] ,
    \Tile_X5Y2_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X5Y2_N1BEG[3] ,
    \Tile_X5Y2_N1BEG[2] ,
    \Tile_X5Y2_N1BEG[1] ,
    \Tile_X5Y2_N1BEG[0] }),
    .N1END({\Tile_X5Y3_N1BEG[3] ,
    \Tile_X5Y3_N1BEG[2] ,
    \Tile_X5Y3_N1BEG[1] ,
    \Tile_X5Y3_N1BEG[0] }),
    .N2BEG({\Tile_X5Y2_N2BEG[7] ,
    \Tile_X5Y2_N2BEG[6] ,
    \Tile_X5Y2_N2BEG[5] ,
    \Tile_X5Y2_N2BEG[4] ,
    \Tile_X5Y2_N2BEG[3] ,
    \Tile_X5Y2_N2BEG[2] ,
    \Tile_X5Y2_N2BEG[1] ,
    \Tile_X5Y2_N2BEG[0] }),
    .N2BEGb({\Tile_X5Y2_N2BEGb[7] ,
    \Tile_X5Y2_N2BEGb[6] ,
    \Tile_X5Y2_N2BEGb[5] ,
    \Tile_X5Y2_N2BEGb[4] ,
    \Tile_X5Y2_N2BEGb[3] ,
    \Tile_X5Y2_N2BEGb[2] ,
    \Tile_X5Y2_N2BEGb[1] ,
    \Tile_X5Y2_N2BEGb[0] }),
    .N2END({\Tile_X5Y3_N2BEGb[7] ,
    \Tile_X5Y3_N2BEGb[6] ,
    \Tile_X5Y3_N2BEGb[5] ,
    \Tile_X5Y3_N2BEGb[4] ,
    \Tile_X5Y3_N2BEGb[3] ,
    \Tile_X5Y3_N2BEGb[2] ,
    \Tile_X5Y3_N2BEGb[1] ,
    \Tile_X5Y3_N2BEGb[0] }),
    .N2MID({\Tile_X5Y3_N2BEG[7] ,
    \Tile_X5Y3_N2BEG[6] ,
    \Tile_X5Y3_N2BEG[5] ,
    \Tile_X5Y3_N2BEG[4] ,
    \Tile_X5Y3_N2BEG[3] ,
    \Tile_X5Y3_N2BEG[2] ,
    \Tile_X5Y3_N2BEG[1] ,
    \Tile_X5Y3_N2BEG[0] }),
    .N4BEG({\Tile_X5Y2_N4BEG[15] ,
    \Tile_X5Y2_N4BEG[14] ,
    \Tile_X5Y2_N4BEG[13] ,
    \Tile_X5Y2_N4BEG[12] ,
    \Tile_X5Y2_N4BEG[11] ,
    \Tile_X5Y2_N4BEG[10] ,
    \Tile_X5Y2_N4BEG[9] ,
    \Tile_X5Y2_N4BEG[8] ,
    \Tile_X5Y2_N4BEG[7] ,
    \Tile_X5Y2_N4BEG[6] ,
    \Tile_X5Y2_N4BEG[5] ,
    \Tile_X5Y2_N4BEG[4] ,
    \Tile_X5Y2_N4BEG[3] ,
    \Tile_X5Y2_N4BEG[2] ,
    \Tile_X5Y2_N4BEG[1] ,
    \Tile_X5Y2_N4BEG[0] }),
    .N4END({\Tile_X5Y3_N4BEG[15] ,
    \Tile_X5Y3_N4BEG[14] ,
    \Tile_X5Y3_N4BEG[13] ,
    \Tile_X5Y3_N4BEG[12] ,
    \Tile_X5Y3_N4BEG[11] ,
    \Tile_X5Y3_N4BEG[10] ,
    \Tile_X5Y3_N4BEG[9] ,
    \Tile_X5Y3_N4BEG[8] ,
    \Tile_X5Y3_N4BEG[7] ,
    \Tile_X5Y3_N4BEG[6] ,
    \Tile_X5Y3_N4BEG[5] ,
    \Tile_X5Y3_N4BEG[4] ,
    \Tile_X5Y3_N4BEG[3] ,
    \Tile_X5Y3_N4BEG[2] ,
    \Tile_X5Y3_N4BEG[1] ,
    \Tile_X5Y3_N4BEG[0] }),
    .NN4BEG({\Tile_X5Y2_NN4BEG[15] ,
    \Tile_X5Y2_NN4BEG[14] ,
    \Tile_X5Y2_NN4BEG[13] ,
    \Tile_X5Y2_NN4BEG[12] ,
    \Tile_X5Y2_NN4BEG[11] ,
    \Tile_X5Y2_NN4BEG[10] ,
    \Tile_X5Y2_NN4BEG[9] ,
    \Tile_X5Y2_NN4BEG[8] ,
    \Tile_X5Y2_NN4BEG[7] ,
    \Tile_X5Y2_NN4BEG[6] ,
    \Tile_X5Y2_NN4BEG[5] ,
    \Tile_X5Y2_NN4BEG[4] ,
    \Tile_X5Y2_NN4BEG[3] ,
    \Tile_X5Y2_NN4BEG[2] ,
    \Tile_X5Y2_NN4BEG[1] ,
    \Tile_X5Y2_NN4BEG[0] }),
    .NN4END({\Tile_X5Y3_NN4BEG[15] ,
    \Tile_X5Y3_NN4BEG[14] ,
    \Tile_X5Y3_NN4BEG[13] ,
    \Tile_X5Y3_NN4BEG[12] ,
    \Tile_X5Y3_NN4BEG[11] ,
    \Tile_X5Y3_NN4BEG[10] ,
    \Tile_X5Y3_NN4BEG[9] ,
    \Tile_X5Y3_NN4BEG[8] ,
    \Tile_X5Y3_NN4BEG[7] ,
    \Tile_X5Y3_NN4BEG[6] ,
    \Tile_X5Y3_NN4BEG[5] ,
    \Tile_X5Y3_NN4BEG[4] ,
    \Tile_X5Y3_NN4BEG[3] ,
    \Tile_X5Y3_NN4BEG[2] ,
    \Tile_X5Y3_NN4BEG[1] ,
    \Tile_X5Y3_NN4BEG[0] }),
    .S1BEG({\Tile_X5Y2_S1BEG[3] ,
    \Tile_X5Y2_S1BEG[2] ,
    \Tile_X5Y2_S1BEG[1] ,
    \Tile_X5Y2_S1BEG[0] }),
    .S1END({\Tile_X5Y1_S1BEG[3] ,
    \Tile_X5Y1_S1BEG[2] ,
    \Tile_X5Y1_S1BEG[1] ,
    \Tile_X5Y1_S1BEG[0] }),
    .S2BEG({\Tile_X5Y2_S2BEG[7] ,
    \Tile_X5Y2_S2BEG[6] ,
    \Tile_X5Y2_S2BEG[5] ,
    \Tile_X5Y2_S2BEG[4] ,
    \Tile_X5Y2_S2BEG[3] ,
    \Tile_X5Y2_S2BEG[2] ,
    \Tile_X5Y2_S2BEG[1] ,
    \Tile_X5Y2_S2BEG[0] }),
    .S2BEGb({\Tile_X5Y2_S2BEGb[7] ,
    \Tile_X5Y2_S2BEGb[6] ,
    \Tile_X5Y2_S2BEGb[5] ,
    \Tile_X5Y2_S2BEGb[4] ,
    \Tile_X5Y2_S2BEGb[3] ,
    \Tile_X5Y2_S2BEGb[2] ,
    \Tile_X5Y2_S2BEGb[1] ,
    \Tile_X5Y2_S2BEGb[0] }),
    .S2END({\Tile_X5Y1_S2BEGb[7] ,
    \Tile_X5Y1_S2BEGb[6] ,
    \Tile_X5Y1_S2BEGb[5] ,
    \Tile_X5Y1_S2BEGb[4] ,
    \Tile_X5Y1_S2BEGb[3] ,
    \Tile_X5Y1_S2BEGb[2] ,
    \Tile_X5Y1_S2BEGb[1] ,
    \Tile_X5Y1_S2BEGb[0] }),
    .S2MID({\Tile_X5Y1_S2BEG[7] ,
    \Tile_X5Y1_S2BEG[6] ,
    \Tile_X5Y1_S2BEG[5] ,
    \Tile_X5Y1_S2BEG[4] ,
    \Tile_X5Y1_S2BEG[3] ,
    \Tile_X5Y1_S2BEG[2] ,
    \Tile_X5Y1_S2BEG[1] ,
    \Tile_X5Y1_S2BEG[0] }),
    .S4BEG({\Tile_X5Y2_S4BEG[15] ,
    \Tile_X5Y2_S4BEG[14] ,
    \Tile_X5Y2_S4BEG[13] ,
    \Tile_X5Y2_S4BEG[12] ,
    \Tile_X5Y2_S4BEG[11] ,
    \Tile_X5Y2_S4BEG[10] ,
    \Tile_X5Y2_S4BEG[9] ,
    \Tile_X5Y2_S4BEG[8] ,
    \Tile_X5Y2_S4BEG[7] ,
    \Tile_X5Y2_S4BEG[6] ,
    \Tile_X5Y2_S4BEG[5] ,
    \Tile_X5Y2_S4BEG[4] ,
    \Tile_X5Y2_S4BEG[3] ,
    \Tile_X5Y2_S4BEG[2] ,
    \Tile_X5Y2_S4BEG[1] ,
    \Tile_X5Y2_S4BEG[0] }),
    .S4END({\Tile_X5Y1_S4BEG[15] ,
    \Tile_X5Y1_S4BEG[14] ,
    \Tile_X5Y1_S4BEG[13] ,
    \Tile_X5Y1_S4BEG[12] ,
    \Tile_X5Y1_S4BEG[11] ,
    \Tile_X5Y1_S4BEG[10] ,
    \Tile_X5Y1_S4BEG[9] ,
    \Tile_X5Y1_S4BEG[8] ,
    \Tile_X5Y1_S4BEG[7] ,
    \Tile_X5Y1_S4BEG[6] ,
    \Tile_X5Y1_S4BEG[5] ,
    \Tile_X5Y1_S4BEG[4] ,
    \Tile_X5Y1_S4BEG[3] ,
    \Tile_X5Y1_S4BEG[2] ,
    \Tile_X5Y1_S4BEG[1] ,
    \Tile_X5Y1_S4BEG[0] }),
    .SS4BEG({\Tile_X5Y2_SS4BEG[15] ,
    \Tile_X5Y2_SS4BEG[14] ,
    \Tile_X5Y2_SS4BEG[13] ,
    \Tile_X5Y2_SS4BEG[12] ,
    \Tile_X5Y2_SS4BEG[11] ,
    \Tile_X5Y2_SS4BEG[10] ,
    \Tile_X5Y2_SS4BEG[9] ,
    \Tile_X5Y2_SS4BEG[8] ,
    \Tile_X5Y2_SS4BEG[7] ,
    \Tile_X5Y2_SS4BEG[6] ,
    \Tile_X5Y2_SS4BEG[5] ,
    \Tile_X5Y2_SS4BEG[4] ,
    \Tile_X5Y2_SS4BEG[3] ,
    \Tile_X5Y2_SS4BEG[2] ,
    \Tile_X5Y2_SS4BEG[1] ,
    \Tile_X5Y2_SS4BEG[0] }),
    .SS4END({\Tile_X5Y1_SS4BEG[15] ,
    \Tile_X5Y1_SS4BEG[14] ,
    \Tile_X5Y1_SS4BEG[13] ,
    \Tile_X5Y1_SS4BEG[12] ,
    \Tile_X5Y1_SS4BEG[11] ,
    \Tile_X5Y1_SS4BEG[10] ,
    \Tile_X5Y1_SS4BEG[9] ,
    \Tile_X5Y1_SS4BEG[8] ,
    \Tile_X5Y1_SS4BEG[7] ,
    \Tile_X5Y1_SS4BEG[6] ,
    \Tile_X5Y1_SS4BEG[5] ,
    \Tile_X5Y1_SS4BEG[4] ,
    \Tile_X5Y1_SS4BEG[3] ,
    \Tile_X5Y1_SS4BEG[2] ,
    \Tile_X5Y1_SS4BEG[1] ,
    \Tile_X5Y1_SS4BEG[0] }),
    .W1BEG({\Tile_X5Y2_W1BEG[3] ,
    \Tile_X5Y2_W1BEG[2] ,
    \Tile_X5Y2_W1BEG[1] ,
    \Tile_X5Y2_W1BEG[0] }),
    .W1END({\Tile_X6Y2_W1BEG[3] ,
    \Tile_X6Y2_W1BEG[2] ,
    \Tile_X6Y2_W1BEG[1] ,
    \Tile_X6Y2_W1BEG[0] }),
    .W2BEG({\Tile_X5Y2_W2BEG[7] ,
    \Tile_X5Y2_W2BEG[6] ,
    \Tile_X5Y2_W2BEG[5] ,
    \Tile_X5Y2_W2BEG[4] ,
    \Tile_X5Y2_W2BEG[3] ,
    \Tile_X5Y2_W2BEG[2] ,
    \Tile_X5Y2_W2BEG[1] ,
    \Tile_X5Y2_W2BEG[0] }),
    .W2BEGb({\Tile_X5Y2_W2BEGb[7] ,
    \Tile_X5Y2_W2BEGb[6] ,
    \Tile_X5Y2_W2BEGb[5] ,
    \Tile_X5Y2_W2BEGb[4] ,
    \Tile_X5Y2_W2BEGb[3] ,
    \Tile_X5Y2_W2BEGb[2] ,
    \Tile_X5Y2_W2BEGb[1] ,
    \Tile_X5Y2_W2BEGb[0] }),
    .W2END({\Tile_X6Y2_W2BEGb[7] ,
    \Tile_X6Y2_W2BEGb[6] ,
    \Tile_X6Y2_W2BEGb[5] ,
    \Tile_X6Y2_W2BEGb[4] ,
    \Tile_X6Y2_W2BEGb[3] ,
    \Tile_X6Y2_W2BEGb[2] ,
    \Tile_X6Y2_W2BEGb[1] ,
    \Tile_X6Y2_W2BEGb[0] }),
    .W2MID({\Tile_X6Y2_W2BEG[7] ,
    \Tile_X6Y2_W2BEG[6] ,
    \Tile_X6Y2_W2BEG[5] ,
    \Tile_X6Y2_W2BEG[4] ,
    \Tile_X6Y2_W2BEG[3] ,
    \Tile_X6Y2_W2BEG[2] ,
    \Tile_X6Y2_W2BEG[1] ,
    \Tile_X6Y2_W2BEG[0] }),
    .W6BEG({\Tile_X5Y2_W6BEG[11] ,
    \Tile_X5Y2_W6BEG[10] ,
    \Tile_X5Y2_W6BEG[9] ,
    \Tile_X5Y2_W6BEG[8] ,
    \Tile_X5Y2_W6BEG[7] ,
    \Tile_X5Y2_W6BEG[6] ,
    \Tile_X5Y2_W6BEG[5] ,
    \Tile_X5Y2_W6BEG[4] ,
    \Tile_X5Y2_W6BEG[3] ,
    \Tile_X5Y2_W6BEG[2] ,
    \Tile_X5Y2_W6BEG[1] ,
    \Tile_X5Y2_W6BEG[0] }),
    .W6END({\Tile_X6Y2_W6BEG[11] ,
    \Tile_X6Y2_W6BEG[10] ,
    \Tile_X6Y2_W6BEG[9] ,
    \Tile_X6Y2_W6BEG[8] ,
    \Tile_X6Y2_W6BEG[7] ,
    \Tile_X6Y2_W6BEG[6] ,
    \Tile_X6Y2_W6BEG[5] ,
    \Tile_X6Y2_W6BEG[4] ,
    \Tile_X6Y2_W6BEG[3] ,
    \Tile_X6Y2_W6BEG[2] ,
    \Tile_X6Y2_W6BEG[1] ,
    \Tile_X6Y2_W6BEG[0] }),
    .WW4BEG({\Tile_X5Y2_WW4BEG[15] ,
    \Tile_X5Y2_WW4BEG[14] ,
    \Tile_X5Y2_WW4BEG[13] ,
    \Tile_X5Y2_WW4BEG[12] ,
    \Tile_X5Y2_WW4BEG[11] ,
    \Tile_X5Y2_WW4BEG[10] ,
    \Tile_X5Y2_WW4BEG[9] ,
    \Tile_X5Y2_WW4BEG[8] ,
    \Tile_X5Y2_WW4BEG[7] ,
    \Tile_X5Y2_WW4BEG[6] ,
    \Tile_X5Y2_WW4BEG[5] ,
    \Tile_X5Y2_WW4BEG[4] ,
    \Tile_X5Y2_WW4BEG[3] ,
    \Tile_X5Y2_WW4BEG[2] ,
    \Tile_X5Y2_WW4BEG[1] ,
    \Tile_X5Y2_WW4BEG[0] }),
    .WW4END({\Tile_X6Y2_WW4BEG[15] ,
    \Tile_X6Y2_WW4BEG[14] ,
    \Tile_X6Y2_WW4BEG[13] ,
    \Tile_X6Y2_WW4BEG[12] ,
    \Tile_X6Y2_WW4BEG[11] ,
    \Tile_X6Y2_WW4BEG[10] ,
    \Tile_X6Y2_WW4BEG[9] ,
    \Tile_X6Y2_WW4BEG[8] ,
    \Tile_X6Y2_WW4BEG[7] ,
    \Tile_X6Y2_WW4BEG[6] ,
    \Tile_X6Y2_WW4BEG[5] ,
    \Tile_X6Y2_WW4BEG[4] ,
    \Tile_X6Y2_WW4BEG[3] ,
    \Tile_X6Y2_WW4BEG[2] ,
    \Tile_X6Y2_WW4BEG[1] ,
    \Tile_X6Y2_WW4BEG[0] }));
 LUT4AB Tile_X5Y3_LUT4AB (.Ci(Tile_X5Y4_Co),
    .Co(Tile_X5Y3_Co),
    .UserCLK(Tile_X5Y4_UserCLKo),
    .UserCLKo(Tile_X5Y3_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X5Y3_E1BEG[3] ,
    \Tile_X5Y3_E1BEG[2] ,
    \Tile_X5Y3_E1BEG[1] ,
    \Tile_X5Y3_E1BEG[0] }),
    .E1END({\Tile_X4Y3_E1BEG[3] ,
    \Tile_X4Y3_E1BEG[2] ,
    \Tile_X4Y3_E1BEG[1] ,
    \Tile_X4Y3_E1BEG[0] }),
    .E2BEG({\Tile_X5Y3_E2BEG[7] ,
    \Tile_X5Y3_E2BEG[6] ,
    \Tile_X5Y3_E2BEG[5] ,
    \Tile_X5Y3_E2BEG[4] ,
    \Tile_X5Y3_E2BEG[3] ,
    \Tile_X5Y3_E2BEG[2] ,
    \Tile_X5Y3_E2BEG[1] ,
    \Tile_X5Y3_E2BEG[0] }),
    .E2BEGb({\Tile_X5Y3_E2BEGb[7] ,
    \Tile_X5Y3_E2BEGb[6] ,
    \Tile_X5Y3_E2BEGb[5] ,
    \Tile_X5Y3_E2BEGb[4] ,
    \Tile_X5Y3_E2BEGb[3] ,
    \Tile_X5Y3_E2BEGb[2] ,
    \Tile_X5Y3_E2BEGb[1] ,
    \Tile_X5Y3_E2BEGb[0] }),
    .E2END({\Tile_X4Y3_E2BEGb[7] ,
    \Tile_X4Y3_E2BEGb[6] ,
    \Tile_X4Y3_E2BEGb[5] ,
    \Tile_X4Y3_E2BEGb[4] ,
    \Tile_X4Y3_E2BEGb[3] ,
    \Tile_X4Y3_E2BEGb[2] ,
    \Tile_X4Y3_E2BEGb[1] ,
    \Tile_X4Y3_E2BEGb[0] }),
    .E2MID({\Tile_X4Y3_E2BEG[7] ,
    \Tile_X4Y3_E2BEG[6] ,
    \Tile_X4Y3_E2BEG[5] ,
    \Tile_X4Y3_E2BEG[4] ,
    \Tile_X4Y3_E2BEG[3] ,
    \Tile_X4Y3_E2BEG[2] ,
    \Tile_X4Y3_E2BEG[1] ,
    \Tile_X4Y3_E2BEG[0] }),
    .E6BEG({\Tile_X5Y3_E6BEG[11] ,
    \Tile_X5Y3_E6BEG[10] ,
    \Tile_X5Y3_E6BEG[9] ,
    \Tile_X5Y3_E6BEG[8] ,
    \Tile_X5Y3_E6BEG[7] ,
    \Tile_X5Y3_E6BEG[6] ,
    \Tile_X5Y3_E6BEG[5] ,
    \Tile_X5Y3_E6BEG[4] ,
    \Tile_X5Y3_E6BEG[3] ,
    \Tile_X5Y3_E6BEG[2] ,
    \Tile_X5Y3_E6BEG[1] ,
    \Tile_X5Y3_E6BEG[0] }),
    .E6END({\Tile_X4Y3_E6BEG[11] ,
    \Tile_X4Y3_E6BEG[10] ,
    \Tile_X4Y3_E6BEG[9] ,
    \Tile_X4Y3_E6BEG[8] ,
    \Tile_X4Y3_E6BEG[7] ,
    \Tile_X4Y3_E6BEG[6] ,
    \Tile_X4Y3_E6BEG[5] ,
    \Tile_X4Y3_E6BEG[4] ,
    \Tile_X4Y3_E6BEG[3] ,
    \Tile_X4Y3_E6BEG[2] ,
    \Tile_X4Y3_E6BEG[1] ,
    \Tile_X4Y3_E6BEG[0] }),
    .EE4BEG({\Tile_X5Y3_EE4BEG[15] ,
    \Tile_X5Y3_EE4BEG[14] ,
    \Tile_X5Y3_EE4BEG[13] ,
    \Tile_X5Y3_EE4BEG[12] ,
    \Tile_X5Y3_EE4BEG[11] ,
    \Tile_X5Y3_EE4BEG[10] ,
    \Tile_X5Y3_EE4BEG[9] ,
    \Tile_X5Y3_EE4BEG[8] ,
    \Tile_X5Y3_EE4BEG[7] ,
    \Tile_X5Y3_EE4BEG[6] ,
    \Tile_X5Y3_EE4BEG[5] ,
    \Tile_X5Y3_EE4BEG[4] ,
    \Tile_X5Y3_EE4BEG[3] ,
    \Tile_X5Y3_EE4BEG[2] ,
    \Tile_X5Y3_EE4BEG[1] ,
    \Tile_X5Y3_EE4BEG[0] }),
    .EE4END({\Tile_X4Y3_EE4BEG[15] ,
    \Tile_X4Y3_EE4BEG[14] ,
    \Tile_X4Y3_EE4BEG[13] ,
    \Tile_X4Y3_EE4BEG[12] ,
    \Tile_X4Y3_EE4BEG[11] ,
    \Tile_X4Y3_EE4BEG[10] ,
    \Tile_X4Y3_EE4BEG[9] ,
    \Tile_X4Y3_EE4BEG[8] ,
    \Tile_X4Y3_EE4BEG[7] ,
    \Tile_X4Y3_EE4BEG[6] ,
    \Tile_X4Y3_EE4BEG[5] ,
    \Tile_X4Y3_EE4BEG[4] ,
    \Tile_X4Y3_EE4BEG[3] ,
    \Tile_X4Y3_EE4BEG[2] ,
    \Tile_X4Y3_EE4BEG[1] ,
    \Tile_X4Y3_EE4BEG[0] }),
    .FrameData({\Tile_X4Y3_FrameData_O[31] ,
    \Tile_X4Y3_FrameData_O[30] ,
    \Tile_X4Y3_FrameData_O[29] ,
    \Tile_X4Y3_FrameData_O[28] ,
    \Tile_X4Y3_FrameData_O[27] ,
    \Tile_X4Y3_FrameData_O[26] ,
    \Tile_X4Y3_FrameData_O[25] ,
    \Tile_X4Y3_FrameData_O[24] ,
    \Tile_X4Y3_FrameData_O[23] ,
    \Tile_X4Y3_FrameData_O[22] ,
    \Tile_X4Y3_FrameData_O[21] ,
    \Tile_X4Y3_FrameData_O[20] ,
    \Tile_X4Y3_FrameData_O[19] ,
    \Tile_X4Y3_FrameData_O[18] ,
    \Tile_X4Y3_FrameData_O[17] ,
    \Tile_X4Y3_FrameData_O[16] ,
    \Tile_X4Y3_FrameData_O[15] ,
    \Tile_X4Y3_FrameData_O[14] ,
    \Tile_X4Y3_FrameData_O[13] ,
    \Tile_X4Y3_FrameData_O[12] ,
    \Tile_X4Y3_FrameData_O[11] ,
    \Tile_X4Y3_FrameData_O[10] ,
    \Tile_X4Y3_FrameData_O[9] ,
    \Tile_X4Y3_FrameData_O[8] ,
    \Tile_X4Y3_FrameData_O[7] ,
    \Tile_X4Y3_FrameData_O[6] ,
    \Tile_X4Y3_FrameData_O[5] ,
    \Tile_X4Y3_FrameData_O[4] ,
    \Tile_X4Y3_FrameData_O[3] ,
    \Tile_X4Y3_FrameData_O[2] ,
    \Tile_X4Y3_FrameData_O[1] ,
    \Tile_X4Y3_FrameData_O[0] }),
    .FrameData_O({\Tile_X5Y3_FrameData_O[31] ,
    \Tile_X5Y3_FrameData_O[30] ,
    \Tile_X5Y3_FrameData_O[29] ,
    \Tile_X5Y3_FrameData_O[28] ,
    \Tile_X5Y3_FrameData_O[27] ,
    \Tile_X5Y3_FrameData_O[26] ,
    \Tile_X5Y3_FrameData_O[25] ,
    \Tile_X5Y3_FrameData_O[24] ,
    \Tile_X5Y3_FrameData_O[23] ,
    \Tile_X5Y3_FrameData_O[22] ,
    \Tile_X5Y3_FrameData_O[21] ,
    \Tile_X5Y3_FrameData_O[20] ,
    \Tile_X5Y3_FrameData_O[19] ,
    \Tile_X5Y3_FrameData_O[18] ,
    \Tile_X5Y3_FrameData_O[17] ,
    \Tile_X5Y3_FrameData_O[16] ,
    \Tile_X5Y3_FrameData_O[15] ,
    \Tile_X5Y3_FrameData_O[14] ,
    \Tile_X5Y3_FrameData_O[13] ,
    \Tile_X5Y3_FrameData_O[12] ,
    \Tile_X5Y3_FrameData_O[11] ,
    \Tile_X5Y3_FrameData_O[10] ,
    \Tile_X5Y3_FrameData_O[9] ,
    \Tile_X5Y3_FrameData_O[8] ,
    \Tile_X5Y3_FrameData_O[7] ,
    \Tile_X5Y3_FrameData_O[6] ,
    \Tile_X5Y3_FrameData_O[5] ,
    \Tile_X5Y3_FrameData_O[4] ,
    \Tile_X5Y3_FrameData_O[3] ,
    \Tile_X5Y3_FrameData_O[2] ,
    \Tile_X5Y3_FrameData_O[1] ,
    \Tile_X5Y3_FrameData_O[0] }),
    .FrameStrobe({\Tile_X5Y4_FrameStrobe_O[19] ,
    \Tile_X5Y4_FrameStrobe_O[18] ,
    \Tile_X5Y4_FrameStrobe_O[17] ,
    \Tile_X5Y4_FrameStrobe_O[16] ,
    \Tile_X5Y4_FrameStrobe_O[15] ,
    \Tile_X5Y4_FrameStrobe_O[14] ,
    \Tile_X5Y4_FrameStrobe_O[13] ,
    \Tile_X5Y4_FrameStrobe_O[12] ,
    \Tile_X5Y4_FrameStrobe_O[11] ,
    \Tile_X5Y4_FrameStrobe_O[10] ,
    \Tile_X5Y4_FrameStrobe_O[9] ,
    \Tile_X5Y4_FrameStrobe_O[8] ,
    \Tile_X5Y4_FrameStrobe_O[7] ,
    \Tile_X5Y4_FrameStrobe_O[6] ,
    \Tile_X5Y4_FrameStrobe_O[5] ,
    \Tile_X5Y4_FrameStrobe_O[4] ,
    \Tile_X5Y4_FrameStrobe_O[3] ,
    \Tile_X5Y4_FrameStrobe_O[2] ,
    \Tile_X5Y4_FrameStrobe_O[1] ,
    \Tile_X5Y4_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X5Y3_FrameStrobe_O[19] ,
    \Tile_X5Y3_FrameStrobe_O[18] ,
    \Tile_X5Y3_FrameStrobe_O[17] ,
    \Tile_X5Y3_FrameStrobe_O[16] ,
    \Tile_X5Y3_FrameStrobe_O[15] ,
    \Tile_X5Y3_FrameStrobe_O[14] ,
    \Tile_X5Y3_FrameStrobe_O[13] ,
    \Tile_X5Y3_FrameStrobe_O[12] ,
    \Tile_X5Y3_FrameStrobe_O[11] ,
    \Tile_X5Y3_FrameStrobe_O[10] ,
    \Tile_X5Y3_FrameStrobe_O[9] ,
    \Tile_X5Y3_FrameStrobe_O[8] ,
    \Tile_X5Y3_FrameStrobe_O[7] ,
    \Tile_X5Y3_FrameStrobe_O[6] ,
    \Tile_X5Y3_FrameStrobe_O[5] ,
    \Tile_X5Y3_FrameStrobe_O[4] ,
    \Tile_X5Y3_FrameStrobe_O[3] ,
    \Tile_X5Y3_FrameStrobe_O[2] ,
    \Tile_X5Y3_FrameStrobe_O[1] ,
    \Tile_X5Y3_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X5Y3_N1BEG[3] ,
    \Tile_X5Y3_N1BEG[2] ,
    \Tile_X5Y3_N1BEG[1] ,
    \Tile_X5Y3_N1BEG[0] }),
    .N1END({\Tile_X5Y4_N1BEG[3] ,
    \Tile_X5Y4_N1BEG[2] ,
    \Tile_X5Y4_N1BEG[1] ,
    \Tile_X5Y4_N1BEG[0] }),
    .N2BEG({\Tile_X5Y3_N2BEG[7] ,
    \Tile_X5Y3_N2BEG[6] ,
    \Tile_X5Y3_N2BEG[5] ,
    \Tile_X5Y3_N2BEG[4] ,
    \Tile_X5Y3_N2BEG[3] ,
    \Tile_X5Y3_N2BEG[2] ,
    \Tile_X5Y3_N2BEG[1] ,
    \Tile_X5Y3_N2BEG[0] }),
    .N2BEGb({\Tile_X5Y3_N2BEGb[7] ,
    \Tile_X5Y3_N2BEGb[6] ,
    \Tile_X5Y3_N2BEGb[5] ,
    \Tile_X5Y3_N2BEGb[4] ,
    \Tile_X5Y3_N2BEGb[3] ,
    \Tile_X5Y3_N2BEGb[2] ,
    \Tile_X5Y3_N2BEGb[1] ,
    \Tile_X5Y3_N2BEGb[0] }),
    .N2END({\Tile_X5Y4_N2BEGb[7] ,
    \Tile_X5Y4_N2BEGb[6] ,
    \Tile_X5Y4_N2BEGb[5] ,
    \Tile_X5Y4_N2BEGb[4] ,
    \Tile_X5Y4_N2BEGb[3] ,
    \Tile_X5Y4_N2BEGb[2] ,
    \Tile_X5Y4_N2BEGb[1] ,
    \Tile_X5Y4_N2BEGb[0] }),
    .N2MID({\Tile_X5Y4_N2BEG[7] ,
    \Tile_X5Y4_N2BEG[6] ,
    \Tile_X5Y4_N2BEG[5] ,
    \Tile_X5Y4_N2BEG[4] ,
    \Tile_X5Y4_N2BEG[3] ,
    \Tile_X5Y4_N2BEG[2] ,
    \Tile_X5Y4_N2BEG[1] ,
    \Tile_X5Y4_N2BEG[0] }),
    .N4BEG({\Tile_X5Y3_N4BEG[15] ,
    \Tile_X5Y3_N4BEG[14] ,
    \Tile_X5Y3_N4BEG[13] ,
    \Tile_X5Y3_N4BEG[12] ,
    \Tile_X5Y3_N4BEG[11] ,
    \Tile_X5Y3_N4BEG[10] ,
    \Tile_X5Y3_N4BEG[9] ,
    \Tile_X5Y3_N4BEG[8] ,
    \Tile_X5Y3_N4BEG[7] ,
    \Tile_X5Y3_N4BEG[6] ,
    \Tile_X5Y3_N4BEG[5] ,
    \Tile_X5Y3_N4BEG[4] ,
    \Tile_X5Y3_N4BEG[3] ,
    \Tile_X5Y3_N4BEG[2] ,
    \Tile_X5Y3_N4BEG[1] ,
    \Tile_X5Y3_N4BEG[0] }),
    .N4END({\Tile_X5Y4_N4BEG[15] ,
    \Tile_X5Y4_N4BEG[14] ,
    \Tile_X5Y4_N4BEG[13] ,
    \Tile_X5Y4_N4BEG[12] ,
    \Tile_X5Y4_N4BEG[11] ,
    \Tile_X5Y4_N4BEG[10] ,
    \Tile_X5Y4_N4BEG[9] ,
    \Tile_X5Y4_N4BEG[8] ,
    \Tile_X5Y4_N4BEG[7] ,
    \Tile_X5Y4_N4BEG[6] ,
    \Tile_X5Y4_N4BEG[5] ,
    \Tile_X5Y4_N4BEG[4] ,
    \Tile_X5Y4_N4BEG[3] ,
    \Tile_X5Y4_N4BEG[2] ,
    \Tile_X5Y4_N4BEG[1] ,
    \Tile_X5Y4_N4BEG[0] }),
    .NN4BEG({\Tile_X5Y3_NN4BEG[15] ,
    \Tile_X5Y3_NN4BEG[14] ,
    \Tile_X5Y3_NN4BEG[13] ,
    \Tile_X5Y3_NN4BEG[12] ,
    \Tile_X5Y3_NN4BEG[11] ,
    \Tile_X5Y3_NN4BEG[10] ,
    \Tile_X5Y3_NN4BEG[9] ,
    \Tile_X5Y3_NN4BEG[8] ,
    \Tile_X5Y3_NN4BEG[7] ,
    \Tile_X5Y3_NN4BEG[6] ,
    \Tile_X5Y3_NN4BEG[5] ,
    \Tile_X5Y3_NN4BEG[4] ,
    \Tile_X5Y3_NN4BEG[3] ,
    \Tile_X5Y3_NN4BEG[2] ,
    \Tile_X5Y3_NN4BEG[1] ,
    \Tile_X5Y3_NN4BEG[0] }),
    .NN4END({\Tile_X5Y4_NN4BEG[15] ,
    \Tile_X5Y4_NN4BEG[14] ,
    \Tile_X5Y4_NN4BEG[13] ,
    \Tile_X5Y4_NN4BEG[12] ,
    \Tile_X5Y4_NN4BEG[11] ,
    \Tile_X5Y4_NN4BEG[10] ,
    \Tile_X5Y4_NN4BEG[9] ,
    \Tile_X5Y4_NN4BEG[8] ,
    \Tile_X5Y4_NN4BEG[7] ,
    \Tile_X5Y4_NN4BEG[6] ,
    \Tile_X5Y4_NN4BEG[5] ,
    \Tile_X5Y4_NN4BEG[4] ,
    \Tile_X5Y4_NN4BEG[3] ,
    \Tile_X5Y4_NN4BEG[2] ,
    \Tile_X5Y4_NN4BEG[1] ,
    \Tile_X5Y4_NN4BEG[0] }),
    .S1BEG({\Tile_X5Y3_S1BEG[3] ,
    \Tile_X5Y3_S1BEG[2] ,
    \Tile_X5Y3_S1BEG[1] ,
    \Tile_X5Y3_S1BEG[0] }),
    .S1END({\Tile_X5Y2_S1BEG[3] ,
    \Tile_X5Y2_S1BEG[2] ,
    \Tile_X5Y2_S1BEG[1] ,
    \Tile_X5Y2_S1BEG[0] }),
    .S2BEG({\Tile_X5Y3_S2BEG[7] ,
    \Tile_X5Y3_S2BEG[6] ,
    \Tile_X5Y3_S2BEG[5] ,
    \Tile_X5Y3_S2BEG[4] ,
    \Tile_X5Y3_S2BEG[3] ,
    \Tile_X5Y3_S2BEG[2] ,
    \Tile_X5Y3_S2BEG[1] ,
    \Tile_X5Y3_S2BEG[0] }),
    .S2BEGb({\Tile_X5Y3_S2BEGb[7] ,
    \Tile_X5Y3_S2BEGb[6] ,
    \Tile_X5Y3_S2BEGb[5] ,
    \Tile_X5Y3_S2BEGb[4] ,
    \Tile_X5Y3_S2BEGb[3] ,
    \Tile_X5Y3_S2BEGb[2] ,
    \Tile_X5Y3_S2BEGb[1] ,
    \Tile_X5Y3_S2BEGb[0] }),
    .S2END({\Tile_X5Y2_S2BEGb[7] ,
    \Tile_X5Y2_S2BEGb[6] ,
    \Tile_X5Y2_S2BEGb[5] ,
    \Tile_X5Y2_S2BEGb[4] ,
    \Tile_X5Y2_S2BEGb[3] ,
    \Tile_X5Y2_S2BEGb[2] ,
    \Tile_X5Y2_S2BEGb[1] ,
    \Tile_X5Y2_S2BEGb[0] }),
    .S2MID({\Tile_X5Y2_S2BEG[7] ,
    \Tile_X5Y2_S2BEG[6] ,
    \Tile_X5Y2_S2BEG[5] ,
    \Tile_X5Y2_S2BEG[4] ,
    \Tile_X5Y2_S2BEG[3] ,
    \Tile_X5Y2_S2BEG[2] ,
    \Tile_X5Y2_S2BEG[1] ,
    \Tile_X5Y2_S2BEG[0] }),
    .S4BEG({\Tile_X5Y3_S4BEG[15] ,
    \Tile_X5Y3_S4BEG[14] ,
    \Tile_X5Y3_S4BEG[13] ,
    \Tile_X5Y3_S4BEG[12] ,
    \Tile_X5Y3_S4BEG[11] ,
    \Tile_X5Y3_S4BEG[10] ,
    \Tile_X5Y3_S4BEG[9] ,
    \Tile_X5Y3_S4BEG[8] ,
    \Tile_X5Y3_S4BEG[7] ,
    \Tile_X5Y3_S4BEG[6] ,
    \Tile_X5Y3_S4BEG[5] ,
    \Tile_X5Y3_S4BEG[4] ,
    \Tile_X5Y3_S4BEG[3] ,
    \Tile_X5Y3_S4BEG[2] ,
    \Tile_X5Y3_S4BEG[1] ,
    \Tile_X5Y3_S4BEG[0] }),
    .S4END({\Tile_X5Y2_S4BEG[15] ,
    \Tile_X5Y2_S4BEG[14] ,
    \Tile_X5Y2_S4BEG[13] ,
    \Tile_X5Y2_S4BEG[12] ,
    \Tile_X5Y2_S4BEG[11] ,
    \Tile_X5Y2_S4BEG[10] ,
    \Tile_X5Y2_S4BEG[9] ,
    \Tile_X5Y2_S4BEG[8] ,
    \Tile_X5Y2_S4BEG[7] ,
    \Tile_X5Y2_S4BEG[6] ,
    \Tile_X5Y2_S4BEG[5] ,
    \Tile_X5Y2_S4BEG[4] ,
    \Tile_X5Y2_S4BEG[3] ,
    \Tile_X5Y2_S4BEG[2] ,
    \Tile_X5Y2_S4BEG[1] ,
    \Tile_X5Y2_S4BEG[0] }),
    .SS4BEG({\Tile_X5Y3_SS4BEG[15] ,
    \Tile_X5Y3_SS4BEG[14] ,
    \Tile_X5Y3_SS4BEG[13] ,
    \Tile_X5Y3_SS4BEG[12] ,
    \Tile_X5Y3_SS4BEG[11] ,
    \Tile_X5Y3_SS4BEG[10] ,
    \Tile_X5Y3_SS4BEG[9] ,
    \Tile_X5Y3_SS4BEG[8] ,
    \Tile_X5Y3_SS4BEG[7] ,
    \Tile_X5Y3_SS4BEG[6] ,
    \Tile_X5Y3_SS4BEG[5] ,
    \Tile_X5Y3_SS4BEG[4] ,
    \Tile_X5Y3_SS4BEG[3] ,
    \Tile_X5Y3_SS4BEG[2] ,
    \Tile_X5Y3_SS4BEG[1] ,
    \Tile_X5Y3_SS4BEG[0] }),
    .SS4END({\Tile_X5Y2_SS4BEG[15] ,
    \Tile_X5Y2_SS4BEG[14] ,
    \Tile_X5Y2_SS4BEG[13] ,
    \Tile_X5Y2_SS4BEG[12] ,
    \Tile_X5Y2_SS4BEG[11] ,
    \Tile_X5Y2_SS4BEG[10] ,
    \Tile_X5Y2_SS4BEG[9] ,
    \Tile_X5Y2_SS4BEG[8] ,
    \Tile_X5Y2_SS4BEG[7] ,
    \Tile_X5Y2_SS4BEG[6] ,
    \Tile_X5Y2_SS4BEG[5] ,
    \Tile_X5Y2_SS4BEG[4] ,
    \Tile_X5Y2_SS4BEG[3] ,
    \Tile_X5Y2_SS4BEG[2] ,
    \Tile_X5Y2_SS4BEG[1] ,
    \Tile_X5Y2_SS4BEG[0] }),
    .W1BEG({\Tile_X5Y3_W1BEG[3] ,
    \Tile_X5Y3_W1BEG[2] ,
    \Tile_X5Y3_W1BEG[1] ,
    \Tile_X5Y3_W1BEG[0] }),
    .W1END({\Tile_X6Y3_W1BEG[3] ,
    \Tile_X6Y3_W1BEG[2] ,
    \Tile_X6Y3_W1BEG[1] ,
    \Tile_X6Y3_W1BEG[0] }),
    .W2BEG({\Tile_X5Y3_W2BEG[7] ,
    \Tile_X5Y3_W2BEG[6] ,
    \Tile_X5Y3_W2BEG[5] ,
    \Tile_X5Y3_W2BEG[4] ,
    \Tile_X5Y3_W2BEG[3] ,
    \Tile_X5Y3_W2BEG[2] ,
    \Tile_X5Y3_W2BEG[1] ,
    \Tile_X5Y3_W2BEG[0] }),
    .W2BEGb({\Tile_X5Y3_W2BEGb[7] ,
    \Tile_X5Y3_W2BEGb[6] ,
    \Tile_X5Y3_W2BEGb[5] ,
    \Tile_X5Y3_W2BEGb[4] ,
    \Tile_X5Y3_W2BEGb[3] ,
    \Tile_X5Y3_W2BEGb[2] ,
    \Tile_X5Y3_W2BEGb[1] ,
    \Tile_X5Y3_W2BEGb[0] }),
    .W2END({\Tile_X6Y3_W2BEGb[7] ,
    \Tile_X6Y3_W2BEGb[6] ,
    \Tile_X6Y3_W2BEGb[5] ,
    \Tile_X6Y3_W2BEGb[4] ,
    \Tile_X6Y3_W2BEGb[3] ,
    \Tile_X6Y3_W2BEGb[2] ,
    \Tile_X6Y3_W2BEGb[1] ,
    \Tile_X6Y3_W2BEGb[0] }),
    .W2MID({\Tile_X6Y3_W2BEG[7] ,
    \Tile_X6Y3_W2BEG[6] ,
    \Tile_X6Y3_W2BEG[5] ,
    \Tile_X6Y3_W2BEG[4] ,
    \Tile_X6Y3_W2BEG[3] ,
    \Tile_X6Y3_W2BEG[2] ,
    \Tile_X6Y3_W2BEG[1] ,
    \Tile_X6Y3_W2BEG[0] }),
    .W6BEG({\Tile_X5Y3_W6BEG[11] ,
    \Tile_X5Y3_W6BEG[10] ,
    \Tile_X5Y3_W6BEG[9] ,
    \Tile_X5Y3_W6BEG[8] ,
    \Tile_X5Y3_W6BEG[7] ,
    \Tile_X5Y3_W6BEG[6] ,
    \Tile_X5Y3_W6BEG[5] ,
    \Tile_X5Y3_W6BEG[4] ,
    \Tile_X5Y3_W6BEG[3] ,
    \Tile_X5Y3_W6BEG[2] ,
    \Tile_X5Y3_W6BEG[1] ,
    \Tile_X5Y3_W6BEG[0] }),
    .W6END({\Tile_X6Y3_W6BEG[11] ,
    \Tile_X6Y3_W6BEG[10] ,
    \Tile_X6Y3_W6BEG[9] ,
    \Tile_X6Y3_W6BEG[8] ,
    \Tile_X6Y3_W6BEG[7] ,
    \Tile_X6Y3_W6BEG[6] ,
    \Tile_X6Y3_W6BEG[5] ,
    \Tile_X6Y3_W6BEG[4] ,
    \Tile_X6Y3_W6BEG[3] ,
    \Tile_X6Y3_W6BEG[2] ,
    \Tile_X6Y3_W6BEG[1] ,
    \Tile_X6Y3_W6BEG[0] }),
    .WW4BEG({\Tile_X5Y3_WW4BEG[15] ,
    \Tile_X5Y3_WW4BEG[14] ,
    \Tile_X5Y3_WW4BEG[13] ,
    \Tile_X5Y3_WW4BEG[12] ,
    \Tile_X5Y3_WW4BEG[11] ,
    \Tile_X5Y3_WW4BEG[10] ,
    \Tile_X5Y3_WW4BEG[9] ,
    \Tile_X5Y3_WW4BEG[8] ,
    \Tile_X5Y3_WW4BEG[7] ,
    \Tile_X5Y3_WW4BEG[6] ,
    \Tile_X5Y3_WW4BEG[5] ,
    \Tile_X5Y3_WW4BEG[4] ,
    \Tile_X5Y3_WW4BEG[3] ,
    \Tile_X5Y3_WW4BEG[2] ,
    \Tile_X5Y3_WW4BEG[1] ,
    \Tile_X5Y3_WW4BEG[0] }),
    .WW4END({\Tile_X6Y3_WW4BEG[15] ,
    \Tile_X6Y3_WW4BEG[14] ,
    \Tile_X6Y3_WW4BEG[13] ,
    \Tile_X6Y3_WW4BEG[12] ,
    \Tile_X6Y3_WW4BEG[11] ,
    \Tile_X6Y3_WW4BEG[10] ,
    \Tile_X6Y3_WW4BEG[9] ,
    \Tile_X6Y3_WW4BEG[8] ,
    \Tile_X6Y3_WW4BEG[7] ,
    \Tile_X6Y3_WW4BEG[6] ,
    \Tile_X6Y3_WW4BEG[5] ,
    \Tile_X6Y3_WW4BEG[4] ,
    \Tile_X6Y3_WW4BEG[3] ,
    \Tile_X6Y3_WW4BEG[2] ,
    \Tile_X6Y3_WW4BEG[1] ,
    \Tile_X6Y3_WW4BEG[0] }));
 LUT4AB Tile_X5Y4_LUT4AB (.Ci(Tile_X5Y5_Co),
    .Co(Tile_X5Y4_Co),
    .UserCLK(Tile_X5Y5_UserCLKo),
    .UserCLKo(Tile_X5Y4_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X5Y4_E1BEG[3] ,
    \Tile_X5Y4_E1BEG[2] ,
    \Tile_X5Y4_E1BEG[1] ,
    \Tile_X5Y4_E1BEG[0] }),
    .E1END({\Tile_X4Y4_E1BEG[3] ,
    \Tile_X4Y4_E1BEG[2] ,
    \Tile_X4Y4_E1BEG[1] ,
    \Tile_X4Y4_E1BEG[0] }),
    .E2BEG({\Tile_X5Y4_E2BEG[7] ,
    \Tile_X5Y4_E2BEG[6] ,
    \Tile_X5Y4_E2BEG[5] ,
    \Tile_X5Y4_E2BEG[4] ,
    \Tile_X5Y4_E2BEG[3] ,
    \Tile_X5Y4_E2BEG[2] ,
    \Tile_X5Y4_E2BEG[1] ,
    \Tile_X5Y4_E2BEG[0] }),
    .E2BEGb({\Tile_X5Y4_E2BEGb[7] ,
    \Tile_X5Y4_E2BEGb[6] ,
    \Tile_X5Y4_E2BEGb[5] ,
    \Tile_X5Y4_E2BEGb[4] ,
    \Tile_X5Y4_E2BEGb[3] ,
    \Tile_X5Y4_E2BEGb[2] ,
    \Tile_X5Y4_E2BEGb[1] ,
    \Tile_X5Y4_E2BEGb[0] }),
    .E2END({\Tile_X4Y4_E2BEGb[7] ,
    \Tile_X4Y4_E2BEGb[6] ,
    \Tile_X4Y4_E2BEGb[5] ,
    \Tile_X4Y4_E2BEGb[4] ,
    \Tile_X4Y4_E2BEGb[3] ,
    \Tile_X4Y4_E2BEGb[2] ,
    \Tile_X4Y4_E2BEGb[1] ,
    \Tile_X4Y4_E2BEGb[0] }),
    .E2MID({\Tile_X4Y4_E2BEG[7] ,
    \Tile_X4Y4_E2BEG[6] ,
    \Tile_X4Y4_E2BEG[5] ,
    \Tile_X4Y4_E2BEG[4] ,
    \Tile_X4Y4_E2BEG[3] ,
    \Tile_X4Y4_E2BEG[2] ,
    \Tile_X4Y4_E2BEG[1] ,
    \Tile_X4Y4_E2BEG[0] }),
    .E6BEG({\Tile_X5Y4_E6BEG[11] ,
    \Tile_X5Y4_E6BEG[10] ,
    \Tile_X5Y4_E6BEG[9] ,
    \Tile_X5Y4_E6BEG[8] ,
    \Tile_X5Y4_E6BEG[7] ,
    \Tile_X5Y4_E6BEG[6] ,
    \Tile_X5Y4_E6BEG[5] ,
    \Tile_X5Y4_E6BEG[4] ,
    \Tile_X5Y4_E6BEG[3] ,
    \Tile_X5Y4_E6BEG[2] ,
    \Tile_X5Y4_E6BEG[1] ,
    \Tile_X5Y4_E6BEG[0] }),
    .E6END({\Tile_X4Y4_E6BEG[11] ,
    \Tile_X4Y4_E6BEG[10] ,
    \Tile_X4Y4_E6BEG[9] ,
    \Tile_X4Y4_E6BEG[8] ,
    \Tile_X4Y4_E6BEG[7] ,
    \Tile_X4Y4_E6BEG[6] ,
    \Tile_X4Y4_E6BEG[5] ,
    \Tile_X4Y4_E6BEG[4] ,
    \Tile_X4Y4_E6BEG[3] ,
    \Tile_X4Y4_E6BEG[2] ,
    \Tile_X4Y4_E6BEG[1] ,
    \Tile_X4Y4_E6BEG[0] }),
    .EE4BEG({\Tile_X5Y4_EE4BEG[15] ,
    \Tile_X5Y4_EE4BEG[14] ,
    \Tile_X5Y4_EE4BEG[13] ,
    \Tile_X5Y4_EE4BEG[12] ,
    \Tile_X5Y4_EE4BEG[11] ,
    \Tile_X5Y4_EE4BEG[10] ,
    \Tile_X5Y4_EE4BEG[9] ,
    \Tile_X5Y4_EE4BEG[8] ,
    \Tile_X5Y4_EE4BEG[7] ,
    \Tile_X5Y4_EE4BEG[6] ,
    \Tile_X5Y4_EE4BEG[5] ,
    \Tile_X5Y4_EE4BEG[4] ,
    \Tile_X5Y4_EE4BEG[3] ,
    \Tile_X5Y4_EE4BEG[2] ,
    \Tile_X5Y4_EE4BEG[1] ,
    \Tile_X5Y4_EE4BEG[0] }),
    .EE4END({\Tile_X4Y4_EE4BEG[15] ,
    \Tile_X4Y4_EE4BEG[14] ,
    \Tile_X4Y4_EE4BEG[13] ,
    \Tile_X4Y4_EE4BEG[12] ,
    \Tile_X4Y4_EE4BEG[11] ,
    \Tile_X4Y4_EE4BEG[10] ,
    \Tile_X4Y4_EE4BEG[9] ,
    \Tile_X4Y4_EE4BEG[8] ,
    \Tile_X4Y4_EE4BEG[7] ,
    \Tile_X4Y4_EE4BEG[6] ,
    \Tile_X4Y4_EE4BEG[5] ,
    \Tile_X4Y4_EE4BEG[4] ,
    \Tile_X4Y4_EE4BEG[3] ,
    \Tile_X4Y4_EE4BEG[2] ,
    \Tile_X4Y4_EE4BEG[1] ,
    \Tile_X4Y4_EE4BEG[0] }),
    .FrameData({\Tile_X4Y4_FrameData_O[31] ,
    \Tile_X4Y4_FrameData_O[30] ,
    \Tile_X4Y4_FrameData_O[29] ,
    \Tile_X4Y4_FrameData_O[28] ,
    \Tile_X4Y4_FrameData_O[27] ,
    \Tile_X4Y4_FrameData_O[26] ,
    \Tile_X4Y4_FrameData_O[25] ,
    \Tile_X4Y4_FrameData_O[24] ,
    \Tile_X4Y4_FrameData_O[23] ,
    \Tile_X4Y4_FrameData_O[22] ,
    \Tile_X4Y4_FrameData_O[21] ,
    \Tile_X4Y4_FrameData_O[20] ,
    \Tile_X4Y4_FrameData_O[19] ,
    \Tile_X4Y4_FrameData_O[18] ,
    \Tile_X4Y4_FrameData_O[17] ,
    \Tile_X4Y4_FrameData_O[16] ,
    \Tile_X4Y4_FrameData_O[15] ,
    \Tile_X4Y4_FrameData_O[14] ,
    \Tile_X4Y4_FrameData_O[13] ,
    \Tile_X4Y4_FrameData_O[12] ,
    \Tile_X4Y4_FrameData_O[11] ,
    \Tile_X4Y4_FrameData_O[10] ,
    \Tile_X4Y4_FrameData_O[9] ,
    \Tile_X4Y4_FrameData_O[8] ,
    \Tile_X4Y4_FrameData_O[7] ,
    \Tile_X4Y4_FrameData_O[6] ,
    \Tile_X4Y4_FrameData_O[5] ,
    \Tile_X4Y4_FrameData_O[4] ,
    \Tile_X4Y4_FrameData_O[3] ,
    \Tile_X4Y4_FrameData_O[2] ,
    \Tile_X4Y4_FrameData_O[1] ,
    \Tile_X4Y4_FrameData_O[0] }),
    .FrameData_O({\Tile_X5Y4_FrameData_O[31] ,
    \Tile_X5Y4_FrameData_O[30] ,
    \Tile_X5Y4_FrameData_O[29] ,
    \Tile_X5Y4_FrameData_O[28] ,
    \Tile_X5Y4_FrameData_O[27] ,
    \Tile_X5Y4_FrameData_O[26] ,
    \Tile_X5Y4_FrameData_O[25] ,
    \Tile_X5Y4_FrameData_O[24] ,
    \Tile_X5Y4_FrameData_O[23] ,
    \Tile_X5Y4_FrameData_O[22] ,
    \Tile_X5Y4_FrameData_O[21] ,
    \Tile_X5Y4_FrameData_O[20] ,
    \Tile_X5Y4_FrameData_O[19] ,
    \Tile_X5Y4_FrameData_O[18] ,
    \Tile_X5Y4_FrameData_O[17] ,
    \Tile_X5Y4_FrameData_O[16] ,
    \Tile_X5Y4_FrameData_O[15] ,
    \Tile_X5Y4_FrameData_O[14] ,
    \Tile_X5Y4_FrameData_O[13] ,
    \Tile_X5Y4_FrameData_O[12] ,
    \Tile_X5Y4_FrameData_O[11] ,
    \Tile_X5Y4_FrameData_O[10] ,
    \Tile_X5Y4_FrameData_O[9] ,
    \Tile_X5Y4_FrameData_O[8] ,
    \Tile_X5Y4_FrameData_O[7] ,
    \Tile_X5Y4_FrameData_O[6] ,
    \Tile_X5Y4_FrameData_O[5] ,
    \Tile_X5Y4_FrameData_O[4] ,
    \Tile_X5Y4_FrameData_O[3] ,
    \Tile_X5Y4_FrameData_O[2] ,
    \Tile_X5Y4_FrameData_O[1] ,
    \Tile_X5Y4_FrameData_O[0] }),
    .FrameStrobe({\Tile_X5Y5_FrameStrobe_O[19] ,
    \Tile_X5Y5_FrameStrobe_O[18] ,
    \Tile_X5Y5_FrameStrobe_O[17] ,
    \Tile_X5Y5_FrameStrobe_O[16] ,
    \Tile_X5Y5_FrameStrobe_O[15] ,
    \Tile_X5Y5_FrameStrobe_O[14] ,
    \Tile_X5Y5_FrameStrobe_O[13] ,
    \Tile_X5Y5_FrameStrobe_O[12] ,
    \Tile_X5Y5_FrameStrobe_O[11] ,
    \Tile_X5Y5_FrameStrobe_O[10] ,
    \Tile_X5Y5_FrameStrobe_O[9] ,
    \Tile_X5Y5_FrameStrobe_O[8] ,
    \Tile_X5Y5_FrameStrobe_O[7] ,
    \Tile_X5Y5_FrameStrobe_O[6] ,
    \Tile_X5Y5_FrameStrobe_O[5] ,
    \Tile_X5Y5_FrameStrobe_O[4] ,
    \Tile_X5Y5_FrameStrobe_O[3] ,
    \Tile_X5Y5_FrameStrobe_O[2] ,
    \Tile_X5Y5_FrameStrobe_O[1] ,
    \Tile_X5Y5_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X5Y4_FrameStrobe_O[19] ,
    \Tile_X5Y4_FrameStrobe_O[18] ,
    \Tile_X5Y4_FrameStrobe_O[17] ,
    \Tile_X5Y4_FrameStrobe_O[16] ,
    \Tile_X5Y4_FrameStrobe_O[15] ,
    \Tile_X5Y4_FrameStrobe_O[14] ,
    \Tile_X5Y4_FrameStrobe_O[13] ,
    \Tile_X5Y4_FrameStrobe_O[12] ,
    \Tile_X5Y4_FrameStrobe_O[11] ,
    \Tile_X5Y4_FrameStrobe_O[10] ,
    \Tile_X5Y4_FrameStrobe_O[9] ,
    \Tile_X5Y4_FrameStrobe_O[8] ,
    \Tile_X5Y4_FrameStrobe_O[7] ,
    \Tile_X5Y4_FrameStrobe_O[6] ,
    \Tile_X5Y4_FrameStrobe_O[5] ,
    \Tile_X5Y4_FrameStrobe_O[4] ,
    \Tile_X5Y4_FrameStrobe_O[3] ,
    \Tile_X5Y4_FrameStrobe_O[2] ,
    \Tile_X5Y4_FrameStrobe_O[1] ,
    \Tile_X5Y4_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X5Y4_N1BEG[3] ,
    \Tile_X5Y4_N1BEG[2] ,
    \Tile_X5Y4_N1BEG[1] ,
    \Tile_X5Y4_N1BEG[0] }),
    .N1END({\Tile_X5Y5_N1BEG[3] ,
    \Tile_X5Y5_N1BEG[2] ,
    \Tile_X5Y5_N1BEG[1] ,
    \Tile_X5Y5_N1BEG[0] }),
    .N2BEG({\Tile_X5Y4_N2BEG[7] ,
    \Tile_X5Y4_N2BEG[6] ,
    \Tile_X5Y4_N2BEG[5] ,
    \Tile_X5Y4_N2BEG[4] ,
    \Tile_X5Y4_N2BEG[3] ,
    \Tile_X5Y4_N2BEG[2] ,
    \Tile_X5Y4_N2BEG[1] ,
    \Tile_X5Y4_N2BEG[0] }),
    .N2BEGb({\Tile_X5Y4_N2BEGb[7] ,
    \Tile_X5Y4_N2BEGb[6] ,
    \Tile_X5Y4_N2BEGb[5] ,
    \Tile_X5Y4_N2BEGb[4] ,
    \Tile_X5Y4_N2BEGb[3] ,
    \Tile_X5Y4_N2BEGb[2] ,
    \Tile_X5Y4_N2BEGb[1] ,
    \Tile_X5Y4_N2BEGb[0] }),
    .N2END({\Tile_X5Y5_N2BEGb[7] ,
    \Tile_X5Y5_N2BEGb[6] ,
    \Tile_X5Y5_N2BEGb[5] ,
    \Tile_X5Y5_N2BEGb[4] ,
    \Tile_X5Y5_N2BEGb[3] ,
    \Tile_X5Y5_N2BEGb[2] ,
    \Tile_X5Y5_N2BEGb[1] ,
    \Tile_X5Y5_N2BEGb[0] }),
    .N2MID({\Tile_X5Y5_N2BEG[7] ,
    \Tile_X5Y5_N2BEG[6] ,
    \Tile_X5Y5_N2BEG[5] ,
    \Tile_X5Y5_N2BEG[4] ,
    \Tile_X5Y5_N2BEG[3] ,
    \Tile_X5Y5_N2BEG[2] ,
    \Tile_X5Y5_N2BEG[1] ,
    \Tile_X5Y5_N2BEG[0] }),
    .N4BEG({\Tile_X5Y4_N4BEG[15] ,
    \Tile_X5Y4_N4BEG[14] ,
    \Tile_X5Y4_N4BEG[13] ,
    \Tile_X5Y4_N4BEG[12] ,
    \Tile_X5Y4_N4BEG[11] ,
    \Tile_X5Y4_N4BEG[10] ,
    \Tile_X5Y4_N4BEG[9] ,
    \Tile_X5Y4_N4BEG[8] ,
    \Tile_X5Y4_N4BEG[7] ,
    \Tile_X5Y4_N4BEG[6] ,
    \Tile_X5Y4_N4BEG[5] ,
    \Tile_X5Y4_N4BEG[4] ,
    \Tile_X5Y4_N4BEG[3] ,
    \Tile_X5Y4_N4BEG[2] ,
    \Tile_X5Y4_N4BEG[1] ,
    \Tile_X5Y4_N4BEG[0] }),
    .N4END({\Tile_X5Y5_N4BEG[15] ,
    \Tile_X5Y5_N4BEG[14] ,
    \Tile_X5Y5_N4BEG[13] ,
    \Tile_X5Y5_N4BEG[12] ,
    \Tile_X5Y5_N4BEG[11] ,
    \Tile_X5Y5_N4BEG[10] ,
    \Tile_X5Y5_N4BEG[9] ,
    \Tile_X5Y5_N4BEG[8] ,
    \Tile_X5Y5_N4BEG[7] ,
    \Tile_X5Y5_N4BEG[6] ,
    \Tile_X5Y5_N4BEG[5] ,
    \Tile_X5Y5_N4BEG[4] ,
    \Tile_X5Y5_N4BEG[3] ,
    \Tile_X5Y5_N4BEG[2] ,
    \Tile_X5Y5_N4BEG[1] ,
    \Tile_X5Y5_N4BEG[0] }),
    .NN4BEG({\Tile_X5Y4_NN4BEG[15] ,
    \Tile_X5Y4_NN4BEG[14] ,
    \Tile_X5Y4_NN4BEG[13] ,
    \Tile_X5Y4_NN4BEG[12] ,
    \Tile_X5Y4_NN4BEG[11] ,
    \Tile_X5Y4_NN4BEG[10] ,
    \Tile_X5Y4_NN4BEG[9] ,
    \Tile_X5Y4_NN4BEG[8] ,
    \Tile_X5Y4_NN4BEG[7] ,
    \Tile_X5Y4_NN4BEG[6] ,
    \Tile_X5Y4_NN4BEG[5] ,
    \Tile_X5Y4_NN4BEG[4] ,
    \Tile_X5Y4_NN4BEG[3] ,
    \Tile_X5Y4_NN4BEG[2] ,
    \Tile_X5Y4_NN4BEG[1] ,
    \Tile_X5Y4_NN4BEG[0] }),
    .NN4END({\Tile_X5Y5_NN4BEG[15] ,
    \Tile_X5Y5_NN4BEG[14] ,
    \Tile_X5Y5_NN4BEG[13] ,
    \Tile_X5Y5_NN4BEG[12] ,
    \Tile_X5Y5_NN4BEG[11] ,
    \Tile_X5Y5_NN4BEG[10] ,
    \Tile_X5Y5_NN4BEG[9] ,
    \Tile_X5Y5_NN4BEG[8] ,
    \Tile_X5Y5_NN4BEG[7] ,
    \Tile_X5Y5_NN4BEG[6] ,
    \Tile_X5Y5_NN4BEG[5] ,
    \Tile_X5Y5_NN4BEG[4] ,
    \Tile_X5Y5_NN4BEG[3] ,
    \Tile_X5Y5_NN4BEG[2] ,
    \Tile_X5Y5_NN4BEG[1] ,
    \Tile_X5Y5_NN4BEG[0] }),
    .S1BEG({\Tile_X5Y4_S1BEG[3] ,
    \Tile_X5Y4_S1BEG[2] ,
    \Tile_X5Y4_S1BEG[1] ,
    \Tile_X5Y4_S1BEG[0] }),
    .S1END({\Tile_X5Y3_S1BEG[3] ,
    \Tile_X5Y3_S1BEG[2] ,
    \Tile_X5Y3_S1BEG[1] ,
    \Tile_X5Y3_S1BEG[0] }),
    .S2BEG({\Tile_X5Y4_S2BEG[7] ,
    \Tile_X5Y4_S2BEG[6] ,
    \Tile_X5Y4_S2BEG[5] ,
    \Tile_X5Y4_S2BEG[4] ,
    \Tile_X5Y4_S2BEG[3] ,
    \Tile_X5Y4_S2BEG[2] ,
    \Tile_X5Y4_S2BEG[1] ,
    \Tile_X5Y4_S2BEG[0] }),
    .S2BEGb({\Tile_X5Y4_S2BEGb[7] ,
    \Tile_X5Y4_S2BEGb[6] ,
    \Tile_X5Y4_S2BEGb[5] ,
    \Tile_X5Y4_S2BEGb[4] ,
    \Tile_X5Y4_S2BEGb[3] ,
    \Tile_X5Y4_S2BEGb[2] ,
    \Tile_X5Y4_S2BEGb[1] ,
    \Tile_X5Y4_S2BEGb[0] }),
    .S2END({\Tile_X5Y3_S2BEGb[7] ,
    \Tile_X5Y3_S2BEGb[6] ,
    \Tile_X5Y3_S2BEGb[5] ,
    \Tile_X5Y3_S2BEGb[4] ,
    \Tile_X5Y3_S2BEGb[3] ,
    \Tile_X5Y3_S2BEGb[2] ,
    \Tile_X5Y3_S2BEGb[1] ,
    \Tile_X5Y3_S2BEGb[0] }),
    .S2MID({\Tile_X5Y3_S2BEG[7] ,
    \Tile_X5Y3_S2BEG[6] ,
    \Tile_X5Y3_S2BEG[5] ,
    \Tile_X5Y3_S2BEG[4] ,
    \Tile_X5Y3_S2BEG[3] ,
    \Tile_X5Y3_S2BEG[2] ,
    \Tile_X5Y3_S2BEG[1] ,
    \Tile_X5Y3_S2BEG[0] }),
    .S4BEG({\Tile_X5Y4_S4BEG[15] ,
    \Tile_X5Y4_S4BEG[14] ,
    \Tile_X5Y4_S4BEG[13] ,
    \Tile_X5Y4_S4BEG[12] ,
    \Tile_X5Y4_S4BEG[11] ,
    \Tile_X5Y4_S4BEG[10] ,
    \Tile_X5Y4_S4BEG[9] ,
    \Tile_X5Y4_S4BEG[8] ,
    \Tile_X5Y4_S4BEG[7] ,
    \Tile_X5Y4_S4BEG[6] ,
    \Tile_X5Y4_S4BEG[5] ,
    \Tile_X5Y4_S4BEG[4] ,
    \Tile_X5Y4_S4BEG[3] ,
    \Tile_X5Y4_S4BEG[2] ,
    \Tile_X5Y4_S4BEG[1] ,
    \Tile_X5Y4_S4BEG[0] }),
    .S4END({\Tile_X5Y3_S4BEG[15] ,
    \Tile_X5Y3_S4BEG[14] ,
    \Tile_X5Y3_S4BEG[13] ,
    \Tile_X5Y3_S4BEG[12] ,
    \Tile_X5Y3_S4BEG[11] ,
    \Tile_X5Y3_S4BEG[10] ,
    \Tile_X5Y3_S4BEG[9] ,
    \Tile_X5Y3_S4BEG[8] ,
    \Tile_X5Y3_S4BEG[7] ,
    \Tile_X5Y3_S4BEG[6] ,
    \Tile_X5Y3_S4BEG[5] ,
    \Tile_X5Y3_S4BEG[4] ,
    \Tile_X5Y3_S4BEG[3] ,
    \Tile_X5Y3_S4BEG[2] ,
    \Tile_X5Y3_S4BEG[1] ,
    \Tile_X5Y3_S4BEG[0] }),
    .SS4BEG({\Tile_X5Y4_SS4BEG[15] ,
    \Tile_X5Y4_SS4BEG[14] ,
    \Tile_X5Y4_SS4BEG[13] ,
    \Tile_X5Y4_SS4BEG[12] ,
    \Tile_X5Y4_SS4BEG[11] ,
    \Tile_X5Y4_SS4BEG[10] ,
    \Tile_X5Y4_SS4BEG[9] ,
    \Tile_X5Y4_SS4BEG[8] ,
    \Tile_X5Y4_SS4BEG[7] ,
    \Tile_X5Y4_SS4BEG[6] ,
    \Tile_X5Y4_SS4BEG[5] ,
    \Tile_X5Y4_SS4BEG[4] ,
    \Tile_X5Y4_SS4BEG[3] ,
    \Tile_X5Y4_SS4BEG[2] ,
    \Tile_X5Y4_SS4BEG[1] ,
    \Tile_X5Y4_SS4BEG[0] }),
    .SS4END({\Tile_X5Y3_SS4BEG[15] ,
    \Tile_X5Y3_SS4BEG[14] ,
    \Tile_X5Y3_SS4BEG[13] ,
    \Tile_X5Y3_SS4BEG[12] ,
    \Tile_X5Y3_SS4BEG[11] ,
    \Tile_X5Y3_SS4BEG[10] ,
    \Tile_X5Y3_SS4BEG[9] ,
    \Tile_X5Y3_SS4BEG[8] ,
    \Tile_X5Y3_SS4BEG[7] ,
    \Tile_X5Y3_SS4BEG[6] ,
    \Tile_X5Y3_SS4BEG[5] ,
    \Tile_X5Y3_SS4BEG[4] ,
    \Tile_X5Y3_SS4BEG[3] ,
    \Tile_X5Y3_SS4BEG[2] ,
    \Tile_X5Y3_SS4BEG[1] ,
    \Tile_X5Y3_SS4BEG[0] }),
    .W1BEG({\Tile_X5Y4_W1BEG[3] ,
    \Tile_X5Y4_W1BEG[2] ,
    \Tile_X5Y4_W1BEG[1] ,
    \Tile_X5Y4_W1BEG[0] }),
    .W1END({\Tile_X6Y4_W1BEG[3] ,
    \Tile_X6Y4_W1BEG[2] ,
    \Tile_X6Y4_W1BEG[1] ,
    \Tile_X6Y4_W1BEG[0] }),
    .W2BEG({\Tile_X5Y4_W2BEG[7] ,
    \Tile_X5Y4_W2BEG[6] ,
    \Tile_X5Y4_W2BEG[5] ,
    \Tile_X5Y4_W2BEG[4] ,
    \Tile_X5Y4_W2BEG[3] ,
    \Tile_X5Y4_W2BEG[2] ,
    \Tile_X5Y4_W2BEG[1] ,
    \Tile_X5Y4_W2BEG[0] }),
    .W2BEGb({\Tile_X5Y4_W2BEGb[7] ,
    \Tile_X5Y4_W2BEGb[6] ,
    \Tile_X5Y4_W2BEGb[5] ,
    \Tile_X5Y4_W2BEGb[4] ,
    \Tile_X5Y4_W2BEGb[3] ,
    \Tile_X5Y4_W2BEGb[2] ,
    \Tile_X5Y4_W2BEGb[1] ,
    \Tile_X5Y4_W2BEGb[0] }),
    .W2END({\Tile_X6Y4_W2BEGb[7] ,
    \Tile_X6Y4_W2BEGb[6] ,
    \Tile_X6Y4_W2BEGb[5] ,
    \Tile_X6Y4_W2BEGb[4] ,
    \Tile_X6Y4_W2BEGb[3] ,
    \Tile_X6Y4_W2BEGb[2] ,
    \Tile_X6Y4_W2BEGb[1] ,
    \Tile_X6Y4_W2BEGb[0] }),
    .W2MID({\Tile_X6Y4_W2BEG[7] ,
    \Tile_X6Y4_W2BEG[6] ,
    \Tile_X6Y4_W2BEG[5] ,
    \Tile_X6Y4_W2BEG[4] ,
    \Tile_X6Y4_W2BEG[3] ,
    \Tile_X6Y4_W2BEG[2] ,
    \Tile_X6Y4_W2BEG[1] ,
    \Tile_X6Y4_W2BEG[0] }),
    .W6BEG({\Tile_X5Y4_W6BEG[11] ,
    \Tile_X5Y4_W6BEG[10] ,
    \Tile_X5Y4_W6BEG[9] ,
    \Tile_X5Y4_W6BEG[8] ,
    \Tile_X5Y4_W6BEG[7] ,
    \Tile_X5Y4_W6BEG[6] ,
    \Tile_X5Y4_W6BEG[5] ,
    \Tile_X5Y4_W6BEG[4] ,
    \Tile_X5Y4_W6BEG[3] ,
    \Tile_X5Y4_W6BEG[2] ,
    \Tile_X5Y4_W6BEG[1] ,
    \Tile_X5Y4_W6BEG[0] }),
    .W6END({\Tile_X6Y4_W6BEG[11] ,
    \Tile_X6Y4_W6BEG[10] ,
    \Tile_X6Y4_W6BEG[9] ,
    \Tile_X6Y4_W6BEG[8] ,
    \Tile_X6Y4_W6BEG[7] ,
    \Tile_X6Y4_W6BEG[6] ,
    \Tile_X6Y4_W6BEG[5] ,
    \Tile_X6Y4_W6BEG[4] ,
    \Tile_X6Y4_W6BEG[3] ,
    \Tile_X6Y4_W6BEG[2] ,
    \Tile_X6Y4_W6BEG[1] ,
    \Tile_X6Y4_W6BEG[0] }),
    .WW4BEG({\Tile_X5Y4_WW4BEG[15] ,
    \Tile_X5Y4_WW4BEG[14] ,
    \Tile_X5Y4_WW4BEG[13] ,
    \Tile_X5Y4_WW4BEG[12] ,
    \Tile_X5Y4_WW4BEG[11] ,
    \Tile_X5Y4_WW4BEG[10] ,
    \Tile_X5Y4_WW4BEG[9] ,
    \Tile_X5Y4_WW4BEG[8] ,
    \Tile_X5Y4_WW4BEG[7] ,
    \Tile_X5Y4_WW4BEG[6] ,
    \Tile_X5Y4_WW4BEG[5] ,
    \Tile_X5Y4_WW4BEG[4] ,
    \Tile_X5Y4_WW4BEG[3] ,
    \Tile_X5Y4_WW4BEG[2] ,
    \Tile_X5Y4_WW4BEG[1] ,
    \Tile_X5Y4_WW4BEG[0] }),
    .WW4END({\Tile_X6Y4_WW4BEG[15] ,
    \Tile_X6Y4_WW4BEG[14] ,
    \Tile_X6Y4_WW4BEG[13] ,
    \Tile_X6Y4_WW4BEG[12] ,
    \Tile_X6Y4_WW4BEG[11] ,
    \Tile_X6Y4_WW4BEG[10] ,
    \Tile_X6Y4_WW4BEG[9] ,
    \Tile_X6Y4_WW4BEG[8] ,
    \Tile_X6Y4_WW4BEG[7] ,
    \Tile_X6Y4_WW4BEG[6] ,
    \Tile_X6Y4_WW4BEG[5] ,
    \Tile_X6Y4_WW4BEG[4] ,
    \Tile_X6Y4_WW4BEG[3] ,
    \Tile_X6Y4_WW4BEG[2] ,
    \Tile_X6Y4_WW4BEG[1] ,
    \Tile_X6Y4_WW4BEG[0] }));
 LUT4AB Tile_X5Y5_LUT4AB (.Ci(Tile_X5Y6_Co),
    .Co(Tile_X5Y5_Co),
    .UserCLK(Tile_X5Y6_UserCLKo),
    .UserCLKo(Tile_X5Y5_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X5Y5_E1BEG[3] ,
    \Tile_X5Y5_E1BEG[2] ,
    \Tile_X5Y5_E1BEG[1] ,
    \Tile_X5Y5_E1BEG[0] }),
    .E1END({\Tile_X4Y5_E1BEG[3] ,
    \Tile_X4Y5_E1BEG[2] ,
    \Tile_X4Y5_E1BEG[1] ,
    \Tile_X4Y5_E1BEG[0] }),
    .E2BEG({\Tile_X5Y5_E2BEG[7] ,
    \Tile_X5Y5_E2BEG[6] ,
    \Tile_X5Y5_E2BEG[5] ,
    \Tile_X5Y5_E2BEG[4] ,
    \Tile_X5Y5_E2BEG[3] ,
    \Tile_X5Y5_E2BEG[2] ,
    \Tile_X5Y5_E2BEG[1] ,
    \Tile_X5Y5_E2BEG[0] }),
    .E2BEGb({\Tile_X5Y5_E2BEGb[7] ,
    \Tile_X5Y5_E2BEGb[6] ,
    \Tile_X5Y5_E2BEGb[5] ,
    \Tile_X5Y5_E2BEGb[4] ,
    \Tile_X5Y5_E2BEGb[3] ,
    \Tile_X5Y5_E2BEGb[2] ,
    \Tile_X5Y5_E2BEGb[1] ,
    \Tile_X5Y5_E2BEGb[0] }),
    .E2END({\Tile_X4Y5_E2BEGb[7] ,
    \Tile_X4Y5_E2BEGb[6] ,
    \Tile_X4Y5_E2BEGb[5] ,
    \Tile_X4Y5_E2BEGb[4] ,
    \Tile_X4Y5_E2BEGb[3] ,
    \Tile_X4Y5_E2BEGb[2] ,
    \Tile_X4Y5_E2BEGb[1] ,
    \Tile_X4Y5_E2BEGb[0] }),
    .E2MID({\Tile_X4Y5_E2BEG[7] ,
    \Tile_X4Y5_E2BEG[6] ,
    \Tile_X4Y5_E2BEG[5] ,
    \Tile_X4Y5_E2BEG[4] ,
    \Tile_X4Y5_E2BEG[3] ,
    \Tile_X4Y5_E2BEG[2] ,
    \Tile_X4Y5_E2BEG[1] ,
    \Tile_X4Y5_E2BEG[0] }),
    .E6BEG({\Tile_X5Y5_E6BEG[11] ,
    \Tile_X5Y5_E6BEG[10] ,
    \Tile_X5Y5_E6BEG[9] ,
    \Tile_X5Y5_E6BEG[8] ,
    \Tile_X5Y5_E6BEG[7] ,
    \Tile_X5Y5_E6BEG[6] ,
    \Tile_X5Y5_E6BEG[5] ,
    \Tile_X5Y5_E6BEG[4] ,
    \Tile_X5Y5_E6BEG[3] ,
    \Tile_X5Y5_E6BEG[2] ,
    \Tile_X5Y5_E6BEG[1] ,
    \Tile_X5Y5_E6BEG[0] }),
    .E6END({\Tile_X4Y5_E6BEG[11] ,
    \Tile_X4Y5_E6BEG[10] ,
    \Tile_X4Y5_E6BEG[9] ,
    \Tile_X4Y5_E6BEG[8] ,
    \Tile_X4Y5_E6BEG[7] ,
    \Tile_X4Y5_E6BEG[6] ,
    \Tile_X4Y5_E6BEG[5] ,
    \Tile_X4Y5_E6BEG[4] ,
    \Tile_X4Y5_E6BEG[3] ,
    \Tile_X4Y5_E6BEG[2] ,
    \Tile_X4Y5_E6BEG[1] ,
    \Tile_X4Y5_E6BEG[0] }),
    .EE4BEG({\Tile_X5Y5_EE4BEG[15] ,
    \Tile_X5Y5_EE4BEG[14] ,
    \Tile_X5Y5_EE4BEG[13] ,
    \Tile_X5Y5_EE4BEG[12] ,
    \Tile_X5Y5_EE4BEG[11] ,
    \Tile_X5Y5_EE4BEG[10] ,
    \Tile_X5Y5_EE4BEG[9] ,
    \Tile_X5Y5_EE4BEG[8] ,
    \Tile_X5Y5_EE4BEG[7] ,
    \Tile_X5Y5_EE4BEG[6] ,
    \Tile_X5Y5_EE4BEG[5] ,
    \Tile_X5Y5_EE4BEG[4] ,
    \Tile_X5Y5_EE4BEG[3] ,
    \Tile_X5Y5_EE4BEG[2] ,
    \Tile_X5Y5_EE4BEG[1] ,
    \Tile_X5Y5_EE4BEG[0] }),
    .EE4END({\Tile_X4Y5_EE4BEG[15] ,
    \Tile_X4Y5_EE4BEG[14] ,
    \Tile_X4Y5_EE4BEG[13] ,
    \Tile_X4Y5_EE4BEG[12] ,
    \Tile_X4Y5_EE4BEG[11] ,
    \Tile_X4Y5_EE4BEG[10] ,
    \Tile_X4Y5_EE4BEG[9] ,
    \Tile_X4Y5_EE4BEG[8] ,
    \Tile_X4Y5_EE4BEG[7] ,
    \Tile_X4Y5_EE4BEG[6] ,
    \Tile_X4Y5_EE4BEG[5] ,
    \Tile_X4Y5_EE4BEG[4] ,
    \Tile_X4Y5_EE4BEG[3] ,
    \Tile_X4Y5_EE4BEG[2] ,
    \Tile_X4Y5_EE4BEG[1] ,
    \Tile_X4Y5_EE4BEG[0] }),
    .FrameData({\Tile_X4Y5_FrameData_O[31] ,
    \Tile_X4Y5_FrameData_O[30] ,
    \Tile_X4Y5_FrameData_O[29] ,
    \Tile_X4Y5_FrameData_O[28] ,
    \Tile_X4Y5_FrameData_O[27] ,
    \Tile_X4Y5_FrameData_O[26] ,
    \Tile_X4Y5_FrameData_O[25] ,
    \Tile_X4Y5_FrameData_O[24] ,
    \Tile_X4Y5_FrameData_O[23] ,
    \Tile_X4Y5_FrameData_O[22] ,
    \Tile_X4Y5_FrameData_O[21] ,
    \Tile_X4Y5_FrameData_O[20] ,
    \Tile_X4Y5_FrameData_O[19] ,
    \Tile_X4Y5_FrameData_O[18] ,
    \Tile_X4Y5_FrameData_O[17] ,
    \Tile_X4Y5_FrameData_O[16] ,
    \Tile_X4Y5_FrameData_O[15] ,
    \Tile_X4Y5_FrameData_O[14] ,
    \Tile_X4Y5_FrameData_O[13] ,
    \Tile_X4Y5_FrameData_O[12] ,
    \Tile_X4Y5_FrameData_O[11] ,
    \Tile_X4Y5_FrameData_O[10] ,
    \Tile_X4Y5_FrameData_O[9] ,
    \Tile_X4Y5_FrameData_O[8] ,
    \Tile_X4Y5_FrameData_O[7] ,
    \Tile_X4Y5_FrameData_O[6] ,
    \Tile_X4Y5_FrameData_O[5] ,
    \Tile_X4Y5_FrameData_O[4] ,
    \Tile_X4Y5_FrameData_O[3] ,
    \Tile_X4Y5_FrameData_O[2] ,
    \Tile_X4Y5_FrameData_O[1] ,
    \Tile_X4Y5_FrameData_O[0] }),
    .FrameData_O({\Tile_X5Y5_FrameData_O[31] ,
    \Tile_X5Y5_FrameData_O[30] ,
    \Tile_X5Y5_FrameData_O[29] ,
    \Tile_X5Y5_FrameData_O[28] ,
    \Tile_X5Y5_FrameData_O[27] ,
    \Tile_X5Y5_FrameData_O[26] ,
    \Tile_X5Y5_FrameData_O[25] ,
    \Tile_X5Y5_FrameData_O[24] ,
    \Tile_X5Y5_FrameData_O[23] ,
    \Tile_X5Y5_FrameData_O[22] ,
    \Tile_X5Y5_FrameData_O[21] ,
    \Tile_X5Y5_FrameData_O[20] ,
    \Tile_X5Y5_FrameData_O[19] ,
    \Tile_X5Y5_FrameData_O[18] ,
    \Tile_X5Y5_FrameData_O[17] ,
    \Tile_X5Y5_FrameData_O[16] ,
    \Tile_X5Y5_FrameData_O[15] ,
    \Tile_X5Y5_FrameData_O[14] ,
    \Tile_X5Y5_FrameData_O[13] ,
    \Tile_X5Y5_FrameData_O[12] ,
    \Tile_X5Y5_FrameData_O[11] ,
    \Tile_X5Y5_FrameData_O[10] ,
    \Tile_X5Y5_FrameData_O[9] ,
    \Tile_X5Y5_FrameData_O[8] ,
    \Tile_X5Y5_FrameData_O[7] ,
    \Tile_X5Y5_FrameData_O[6] ,
    \Tile_X5Y5_FrameData_O[5] ,
    \Tile_X5Y5_FrameData_O[4] ,
    \Tile_X5Y5_FrameData_O[3] ,
    \Tile_X5Y5_FrameData_O[2] ,
    \Tile_X5Y5_FrameData_O[1] ,
    \Tile_X5Y5_FrameData_O[0] }),
    .FrameStrobe({\Tile_X5Y6_FrameStrobe_O[19] ,
    \Tile_X5Y6_FrameStrobe_O[18] ,
    \Tile_X5Y6_FrameStrobe_O[17] ,
    \Tile_X5Y6_FrameStrobe_O[16] ,
    \Tile_X5Y6_FrameStrobe_O[15] ,
    \Tile_X5Y6_FrameStrobe_O[14] ,
    \Tile_X5Y6_FrameStrobe_O[13] ,
    \Tile_X5Y6_FrameStrobe_O[12] ,
    \Tile_X5Y6_FrameStrobe_O[11] ,
    \Tile_X5Y6_FrameStrobe_O[10] ,
    \Tile_X5Y6_FrameStrobe_O[9] ,
    \Tile_X5Y6_FrameStrobe_O[8] ,
    \Tile_X5Y6_FrameStrobe_O[7] ,
    \Tile_X5Y6_FrameStrobe_O[6] ,
    \Tile_X5Y6_FrameStrobe_O[5] ,
    \Tile_X5Y6_FrameStrobe_O[4] ,
    \Tile_X5Y6_FrameStrobe_O[3] ,
    \Tile_X5Y6_FrameStrobe_O[2] ,
    \Tile_X5Y6_FrameStrobe_O[1] ,
    \Tile_X5Y6_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X5Y5_FrameStrobe_O[19] ,
    \Tile_X5Y5_FrameStrobe_O[18] ,
    \Tile_X5Y5_FrameStrobe_O[17] ,
    \Tile_X5Y5_FrameStrobe_O[16] ,
    \Tile_X5Y5_FrameStrobe_O[15] ,
    \Tile_X5Y5_FrameStrobe_O[14] ,
    \Tile_X5Y5_FrameStrobe_O[13] ,
    \Tile_X5Y5_FrameStrobe_O[12] ,
    \Tile_X5Y5_FrameStrobe_O[11] ,
    \Tile_X5Y5_FrameStrobe_O[10] ,
    \Tile_X5Y5_FrameStrobe_O[9] ,
    \Tile_X5Y5_FrameStrobe_O[8] ,
    \Tile_X5Y5_FrameStrobe_O[7] ,
    \Tile_X5Y5_FrameStrobe_O[6] ,
    \Tile_X5Y5_FrameStrobe_O[5] ,
    \Tile_X5Y5_FrameStrobe_O[4] ,
    \Tile_X5Y5_FrameStrobe_O[3] ,
    \Tile_X5Y5_FrameStrobe_O[2] ,
    \Tile_X5Y5_FrameStrobe_O[1] ,
    \Tile_X5Y5_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X5Y5_N1BEG[3] ,
    \Tile_X5Y5_N1BEG[2] ,
    \Tile_X5Y5_N1BEG[1] ,
    \Tile_X5Y5_N1BEG[0] }),
    .N1END({\Tile_X5Y6_N1BEG[3] ,
    \Tile_X5Y6_N1BEG[2] ,
    \Tile_X5Y6_N1BEG[1] ,
    \Tile_X5Y6_N1BEG[0] }),
    .N2BEG({\Tile_X5Y5_N2BEG[7] ,
    \Tile_X5Y5_N2BEG[6] ,
    \Tile_X5Y5_N2BEG[5] ,
    \Tile_X5Y5_N2BEG[4] ,
    \Tile_X5Y5_N2BEG[3] ,
    \Tile_X5Y5_N2BEG[2] ,
    \Tile_X5Y5_N2BEG[1] ,
    \Tile_X5Y5_N2BEG[0] }),
    .N2BEGb({\Tile_X5Y5_N2BEGb[7] ,
    \Tile_X5Y5_N2BEGb[6] ,
    \Tile_X5Y5_N2BEGb[5] ,
    \Tile_X5Y5_N2BEGb[4] ,
    \Tile_X5Y5_N2BEGb[3] ,
    \Tile_X5Y5_N2BEGb[2] ,
    \Tile_X5Y5_N2BEGb[1] ,
    \Tile_X5Y5_N2BEGb[0] }),
    .N2END({\Tile_X5Y6_N2BEGb[7] ,
    \Tile_X5Y6_N2BEGb[6] ,
    \Tile_X5Y6_N2BEGb[5] ,
    \Tile_X5Y6_N2BEGb[4] ,
    \Tile_X5Y6_N2BEGb[3] ,
    \Tile_X5Y6_N2BEGb[2] ,
    \Tile_X5Y6_N2BEGb[1] ,
    \Tile_X5Y6_N2BEGb[0] }),
    .N2MID({\Tile_X5Y6_N2BEG[7] ,
    \Tile_X5Y6_N2BEG[6] ,
    \Tile_X5Y6_N2BEG[5] ,
    \Tile_X5Y6_N2BEG[4] ,
    \Tile_X5Y6_N2BEG[3] ,
    \Tile_X5Y6_N2BEG[2] ,
    \Tile_X5Y6_N2BEG[1] ,
    \Tile_X5Y6_N2BEG[0] }),
    .N4BEG({\Tile_X5Y5_N4BEG[15] ,
    \Tile_X5Y5_N4BEG[14] ,
    \Tile_X5Y5_N4BEG[13] ,
    \Tile_X5Y5_N4BEG[12] ,
    \Tile_X5Y5_N4BEG[11] ,
    \Tile_X5Y5_N4BEG[10] ,
    \Tile_X5Y5_N4BEG[9] ,
    \Tile_X5Y5_N4BEG[8] ,
    \Tile_X5Y5_N4BEG[7] ,
    \Tile_X5Y5_N4BEG[6] ,
    \Tile_X5Y5_N4BEG[5] ,
    \Tile_X5Y5_N4BEG[4] ,
    \Tile_X5Y5_N4BEG[3] ,
    \Tile_X5Y5_N4BEG[2] ,
    \Tile_X5Y5_N4BEG[1] ,
    \Tile_X5Y5_N4BEG[0] }),
    .N4END({\Tile_X5Y6_N4BEG[15] ,
    \Tile_X5Y6_N4BEG[14] ,
    \Tile_X5Y6_N4BEG[13] ,
    \Tile_X5Y6_N4BEG[12] ,
    \Tile_X5Y6_N4BEG[11] ,
    \Tile_X5Y6_N4BEG[10] ,
    \Tile_X5Y6_N4BEG[9] ,
    \Tile_X5Y6_N4BEG[8] ,
    \Tile_X5Y6_N4BEG[7] ,
    \Tile_X5Y6_N4BEG[6] ,
    \Tile_X5Y6_N4BEG[5] ,
    \Tile_X5Y6_N4BEG[4] ,
    \Tile_X5Y6_N4BEG[3] ,
    \Tile_X5Y6_N4BEG[2] ,
    \Tile_X5Y6_N4BEG[1] ,
    \Tile_X5Y6_N4BEG[0] }),
    .NN4BEG({\Tile_X5Y5_NN4BEG[15] ,
    \Tile_X5Y5_NN4BEG[14] ,
    \Tile_X5Y5_NN4BEG[13] ,
    \Tile_X5Y5_NN4BEG[12] ,
    \Tile_X5Y5_NN4BEG[11] ,
    \Tile_X5Y5_NN4BEG[10] ,
    \Tile_X5Y5_NN4BEG[9] ,
    \Tile_X5Y5_NN4BEG[8] ,
    \Tile_X5Y5_NN4BEG[7] ,
    \Tile_X5Y5_NN4BEG[6] ,
    \Tile_X5Y5_NN4BEG[5] ,
    \Tile_X5Y5_NN4BEG[4] ,
    \Tile_X5Y5_NN4BEG[3] ,
    \Tile_X5Y5_NN4BEG[2] ,
    \Tile_X5Y5_NN4BEG[1] ,
    \Tile_X5Y5_NN4BEG[0] }),
    .NN4END({\Tile_X5Y6_NN4BEG[15] ,
    \Tile_X5Y6_NN4BEG[14] ,
    \Tile_X5Y6_NN4BEG[13] ,
    \Tile_X5Y6_NN4BEG[12] ,
    \Tile_X5Y6_NN4BEG[11] ,
    \Tile_X5Y6_NN4BEG[10] ,
    \Tile_X5Y6_NN4BEG[9] ,
    \Tile_X5Y6_NN4BEG[8] ,
    \Tile_X5Y6_NN4BEG[7] ,
    \Tile_X5Y6_NN4BEG[6] ,
    \Tile_X5Y6_NN4BEG[5] ,
    \Tile_X5Y6_NN4BEG[4] ,
    \Tile_X5Y6_NN4BEG[3] ,
    \Tile_X5Y6_NN4BEG[2] ,
    \Tile_X5Y6_NN4BEG[1] ,
    \Tile_X5Y6_NN4BEG[0] }),
    .S1BEG({\Tile_X5Y5_S1BEG[3] ,
    \Tile_X5Y5_S1BEG[2] ,
    \Tile_X5Y5_S1BEG[1] ,
    \Tile_X5Y5_S1BEG[0] }),
    .S1END({\Tile_X5Y4_S1BEG[3] ,
    \Tile_X5Y4_S1BEG[2] ,
    \Tile_X5Y4_S1BEG[1] ,
    \Tile_X5Y4_S1BEG[0] }),
    .S2BEG({\Tile_X5Y5_S2BEG[7] ,
    \Tile_X5Y5_S2BEG[6] ,
    \Tile_X5Y5_S2BEG[5] ,
    \Tile_X5Y5_S2BEG[4] ,
    \Tile_X5Y5_S2BEG[3] ,
    \Tile_X5Y5_S2BEG[2] ,
    \Tile_X5Y5_S2BEG[1] ,
    \Tile_X5Y5_S2BEG[0] }),
    .S2BEGb({\Tile_X5Y5_S2BEGb[7] ,
    \Tile_X5Y5_S2BEGb[6] ,
    \Tile_X5Y5_S2BEGb[5] ,
    \Tile_X5Y5_S2BEGb[4] ,
    \Tile_X5Y5_S2BEGb[3] ,
    \Tile_X5Y5_S2BEGb[2] ,
    \Tile_X5Y5_S2BEGb[1] ,
    \Tile_X5Y5_S2BEGb[0] }),
    .S2END({\Tile_X5Y4_S2BEGb[7] ,
    \Tile_X5Y4_S2BEGb[6] ,
    \Tile_X5Y4_S2BEGb[5] ,
    \Tile_X5Y4_S2BEGb[4] ,
    \Tile_X5Y4_S2BEGb[3] ,
    \Tile_X5Y4_S2BEGb[2] ,
    \Tile_X5Y4_S2BEGb[1] ,
    \Tile_X5Y4_S2BEGb[0] }),
    .S2MID({\Tile_X5Y4_S2BEG[7] ,
    \Tile_X5Y4_S2BEG[6] ,
    \Tile_X5Y4_S2BEG[5] ,
    \Tile_X5Y4_S2BEG[4] ,
    \Tile_X5Y4_S2BEG[3] ,
    \Tile_X5Y4_S2BEG[2] ,
    \Tile_X5Y4_S2BEG[1] ,
    \Tile_X5Y4_S2BEG[0] }),
    .S4BEG({\Tile_X5Y5_S4BEG[15] ,
    \Tile_X5Y5_S4BEG[14] ,
    \Tile_X5Y5_S4BEG[13] ,
    \Tile_X5Y5_S4BEG[12] ,
    \Tile_X5Y5_S4BEG[11] ,
    \Tile_X5Y5_S4BEG[10] ,
    \Tile_X5Y5_S4BEG[9] ,
    \Tile_X5Y5_S4BEG[8] ,
    \Tile_X5Y5_S4BEG[7] ,
    \Tile_X5Y5_S4BEG[6] ,
    \Tile_X5Y5_S4BEG[5] ,
    \Tile_X5Y5_S4BEG[4] ,
    \Tile_X5Y5_S4BEG[3] ,
    \Tile_X5Y5_S4BEG[2] ,
    \Tile_X5Y5_S4BEG[1] ,
    \Tile_X5Y5_S4BEG[0] }),
    .S4END({\Tile_X5Y4_S4BEG[15] ,
    \Tile_X5Y4_S4BEG[14] ,
    \Tile_X5Y4_S4BEG[13] ,
    \Tile_X5Y4_S4BEG[12] ,
    \Tile_X5Y4_S4BEG[11] ,
    \Tile_X5Y4_S4BEG[10] ,
    \Tile_X5Y4_S4BEG[9] ,
    \Tile_X5Y4_S4BEG[8] ,
    \Tile_X5Y4_S4BEG[7] ,
    \Tile_X5Y4_S4BEG[6] ,
    \Tile_X5Y4_S4BEG[5] ,
    \Tile_X5Y4_S4BEG[4] ,
    \Tile_X5Y4_S4BEG[3] ,
    \Tile_X5Y4_S4BEG[2] ,
    \Tile_X5Y4_S4BEG[1] ,
    \Tile_X5Y4_S4BEG[0] }),
    .SS4BEG({\Tile_X5Y5_SS4BEG[15] ,
    \Tile_X5Y5_SS4BEG[14] ,
    \Tile_X5Y5_SS4BEG[13] ,
    \Tile_X5Y5_SS4BEG[12] ,
    \Tile_X5Y5_SS4BEG[11] ,
    \Tile_X5Y5_SS4BEG[10] ,
    \Tile_X5Y5_SS4BEG[9] ,
    \Tile_X5Y5_SS4BEG[8] ,
    \Tile_X5Y5_SS4BEG[7] ,
    \Tile_X5Y5_SS4BEG[6] ,
    \Tile_X5Y5_SS4BEG[5] ,
    \Tile_X5Y5_SS4BEG[4] ,
    \Tile_X5Y5_SS4BEG[3] ,
    \Tile_X5Y5_SS4BEG[2] ,
    \Tile_X5Y5_SS4BEG[1] ,
    \Tile_X5Y5_SS4BEG[0] }),
    .SS4END({\Tile_X5Y4_SS4BEG[15] ,
    \Tile_X5Y4_SS4BEG[14] ,
    \Tile_X5Y4_SS4BEG[13] ,
    \Tile_X5Y4_SS4BEG[12] ,
    \Tile_X5Y4_SS4BEG[11] ,
    \Tile_X5Y4_SS4BEG[10] ,
    \Tile_X5Y4_SS4BEG[9] ,
    \Tile_X5Y4_SS4BEG[8] ,
    \Tile_X5Y4_SS4BEG[7] ,
    \Tile_X5Y4_SS4BEG[6] ,
    \Tile_X5Y4_SS4BEG[5] ,
    \Tile_X5Y4_SS4BEG[4] ,
    \Tile_X5Y4_SS4BEG[3] ,
    \Tile_X5Y4_SS4BEG[2] ,
    \Tile_X5Y4_SS4BEG[1] ,
    \Tile_X5Y4_SS4BEG[0] }),
    .W1BEG({\Tile_X5Y5_W1BEG[3] ,
    \Tile_X5Y5_W1BEG[2] ,
    \Tile_X5Y5_W1BEG[1] ,
    \Tile_X5Y5_W1BEG[0] }),
    .W1END({\Tile_X6Y5_W1BEG[3] ,
    \Tile_X6Y5_W1BEG[2] ,
    \Tile_X6Y5_W1BEG[1] ,
    \Tile_X6Y5_W1BEG[0] }),
    .W2BEG({\Tile_X5Y5_W2BEG[7] ,
    \Tile_X5Y5_W2BEG[6] ,
    \Tile_X5Y5_W2BEG[5] ,
    \Tile_X5Y5_W2BEG[4] ,
    \Tile_X5Y5_W2BEG[3] ,
    \Tile_X5Y5_W2BEG[2] ,
    \Tile_X5Y5_W2BEG[1] ,
    \Tile_X5Y5_W2BEG[0] }),
    .W2BEGb({\Tile_X5Y5_W2BEGb[7] ,
    \Tile_X5Y5_W2BEGb[6] ,
    \Tile_X5Y5_W2BEGb[5] ,
    \Tile_X5Y5_W2BEGb[4] ,
    \Tile_X5Y5_W2BEGb[3] ,
    \Tile_X5Y5_W2BEGb[2] ,
    \Tile_X5Y5_W2BEGb[1] ,
    \Tile_X5Y5_W2BEGb[0] }),
    .W2END({\Tile_X6Y5_W2BEGb[7] ,
    \Tile_X6Y5_W2BEGb[6] ,
    \Tile_X6Y5_W2BEGb[5] ,
    \Tile_X6Y5_W2BEGb[4] ,
    \Tile_X6Y5_W2BEGb[3] ,
    \Tile_X6Y5_W2BEGb[2] ,
    \Tile_X6Y5_W2BEGb[1] ,
    \Tile_X6Y5_W2BEGb[0] }),
    .W2MID({\Tile_X6Y5_W2BEG[7] ,
    \Tile_X6Y5_W2BEG[6] ,
    \Tile_X6Y5_W2BEG[5] ,
    \Tile_X6Y5_W2BEG[4] ,
    \Tile_X6Y5_W2BEG[3] ,
    \Tile_X6Y5_W2BEG[2] ,
    \Tile_X6Y5_W2BEG[1] ,
    \Tile_X6Y5_W2BEG[0] }),
    .W6BEG({\Tile_X5Y5_W6BEG[11] ,
    \Tile_X5Y5_W6BEG[10] ,
    \Tile_X5Y5_W6BEG[9] ,
    \Tile_X5Y5_W6BEG[8] ,
    \Tile_X5Y5_W6BEG[7] ,
    \Tile_X5Y5_W6BEG[6] ,
    \Tile_X5Y5_W6BEG[5] ,
    \Tile_X5Y5_W6BEG[4] ,
    \Tile_X5Y5_W6BEG[3] ,
    \Tile_X5Y5_W6BEG[2] ,
    \Tile_X5Y5_W6BEG[1] ,
    \Tile_X5Y5_W6BEG[0] }),
    .W6END({\Tile_X6Y5_W6BEG[11] ,
    \Tile_X6Y5_W6BEG[10] ,
    \Tile_X6Y5_W6BEG[9] ,
    \Tile_X6Y5_W6BEG[8] ,
    \Tile_X6Y5_W6BEG[7] ,
    \Tile_X6Y5_W6BEG[6] ,
    \Tile_X6Y5_W6BEG[5] ,
    \Tile_X6Y5_W6BEG[4] ,
    \Tile_X6Y5_W6BEG[3] ,
    \Tile_X6Y5_W6BEG[2] ,
    \Tile_X6Y5_W6BEG[1] ,
    \Tile_X6Y5_W6BEG[0] }),
    .WW4BEG({\Tile_X5Y5_WW4BEG[15] ,
    \Tile_X5Y5_WW4BEG[14] ,
    \Tile_X5Y5_WW4BEG[13] ,
    \Tile_X5Y5_WW4BEG[12] ,
    \Tile_X5Y5_WW4BEG[11] ,
    \Tile_X5Y5_WW4BEG[10] ,
    \Tile_X5Y5_WW4BEG[9] ,
    \Tile_X5Y5_WW4BEG[8] ,
    \Tile_X5Y5_WW4BEG[7] ,
    \Tile_X5Y5_WW4BEG[6] ,
    \Tile_X5Y5_WW4BEG[5] ,
    \Tile_X5Y5_WW4BEG[4] ,
    \Tile_X5Y5_WW4BEG[3] ,
    \Tile_X5Y5_WW4BEG[2] ,
    \Tile_X5Y5_WW4BEG[1] ,
    \Tile_X5Y5_WW4BEG[0] }),
    .WW4END({\Tile_X6Y5_WW4BEG[15] ,
    \Tile_X6Y5_WW4BEG[14] ,
    \Tile_X6Y5_WW4BEG[13] ,
    \Tile_X6Y5_WW4BEG[12] ,
    \Tile_X6Y5_WW4BEG[11] ,
    \Tile_X6Y5_WW4BEG[10] ,
    \Tile_X6Y5_WW4BEG[9] ,
    \Tile_X6Y5_WW4BEG[8] ,
    \Tile_X6Y5_WW4BEG[7] ,
    \Tile_X6Y5_WW4BEG[6] ,
    \Tile_X6Y5_WW4BEG[5] ,
    \Tile_X6Y5_WW4BEG[4] ,
    \Tile_X6Y5_WW4BEG[3] ,
    \Tile_X6Y5_WW4BEG[2] ,
    \Tile_X6Y5_WW4BEG[1] ,
    \Tile_X6Y5_WW4BEG[0] }));
 LUT4AB Tile_X5Y6_LUT4AB (.Ci(Tile_X5Y7_Co),
    .Co(Tile_X5Y6_Co),
    .UserCLK(Tile_X5Y7_UserCLKo),
    .UserCLKo(Tile_X5Y6_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X5Y6_E1BEG[3] ,
    \Tile_X5Y6_E1BEG[2] ,
    \Tile_X5Y6_E1BEG[1] ,
    \Tile_X5Y6_E1BEG[0] }),
    .E1END({\Tile_X4Y6_E1BEG[3] ,
    \Tile_X4Y6_E1BEG[2] ,
    \Tile_X4Y6_E1BEG[1] ,
    \Tile_X4Y6_E1BEG[0] }),
    .E2BEG({\Tile_X5Y6_E2BEG[7] ,
    \Tile_X5Y6_E2BEG[6] ,
    \Tile_X5Y6_E2BEG[5] ,
    \Tile_X5Y6_E2BEG[4] ,
    \Tile_X5Y6_E2BEG[3] ,
    \Tile_X5Y6_E2BEG[2] ,
    \Tile_X5Y6_E2BEG[1] ,
    \Tile_X5Y6_E2BEG[0] }),
    .E2BEGb({\Tile_X5Y6_E2BEGb[7] ,
    \Tile_X5Y6_E2BEGb[6] ,
    \Tile_X5Y6_E2BEGb[5] ,
    \Tile_X5Y6_E2BEGb[4] ,
    \Tile_X5Y6_E2BEGb[3] ,
    \Tile_X5Y6_E2BEGb[2] ,
    \Tile_X5Y6_E2BEGb[1] ,
    \Tile_X5Y6_E2BEGb[0] }),
    .E2END({\Tile_X4Y6_E2BEGb[7] ,
    \Tile_X4Y6_E2BEGb[6] ,
    \Tile_X4Y6_E2BEGb[5] ,
    \Tile_X4Y6_E2BEGb[4] ,
    \Tile_X4Y6_E2BEGb[3] ,
    \Tile_X4Y6_E2BEGb[2] ,
    \Tile_X4Y6_E2BEGb[1] ,
    \Tile_X4Y6_E2BEGb[0] }),
    .E2MID({\Tile_X4Y6_E2BEG[7] ,
    \Tile_X4Y6_E2BEG[6] ,
    \Tile_X4Y6_E2BEG[5] ,
    \Tile_X4Y6_E2BEG[4] ,
    \Tile_X4Y6_E2BEG[3] ,
    \Tile_X4Y6_E2BEG[2] ,
    \Tile_X4Y6_E2BEG[1] ,
    \Tile_X4Y6_E2BEG[0] }),
    .E6BEG({\Tile_X5Y6_E6BEG[11] ,
    \Tile_X5Y6_E6BEG[10] ,
    \Tile_X5Y6_E6BEG[9] ,
    \Tile_X5Y6_E6BEG[8] ,
    \Tile_X5Y6_E6BEG[7] ,
    \Tile_X5Y6_E6BEG[6] ,
    \Tile_X5Y6_E6BEG[5] ,
    \Tile_X5Y6_E6BEG[4] ,
    \Tile_X5Y6_E6BEG[3] ,
    \Tile_X5Y6_E6BEG[2] ,
    \Tile_X5Y6_E6BEG[1] ,
    \Tile_X5Y6_E6BEG[0] }),
    .E6END({\Tile_X4Y6_E6BEG[11] ,
    \Tile_X4Y6_E6BEG[10] ,
    \Tile_X4Y6_E6BEG[9] ,
    \Tile_X4Y6_E6BEG[8] ,
    \Tile_X4Y6_E6BEG[7] ,
    \Tile_X4Y6_E6BEG[6] ,
    \Tile_X4Y6_E6BEG[5] ,
    \Tile_X4Y6_E6BEG[4] ,
    \Tile_X4Y6_E6BEG[3] ,
    \Tile_X4Y6_E6BEG[2] ,
    \Tile_X4Y6_E6BEG[1] ,
    \Tile_X4Y6_E6BEG[0] }),
    .EE4BEG({\Tile_X5Y6_EE4BEG[15] ,
    \Tile_X5Y6_EE4BEG[14] ,
    \Tile_X5Y6_EE4BEG[13] ,
    \Tile_X5Y6_EE4BEG[12] ,
    \Tile_X5Y6_EE4BEG[11] ,
    \Tile_X5Y6_EE4BEG[10] ,
    \Tile_X5Y6_EE4BEG[9] ,
    \Tile_X5Y6_EE4BEG[8] ,
    \Tile_X5Y6_EE4BEG[7] ,
    \Tile_X5Y6_EE4BEG[6] ,
    \Tile_X5Y6_EE4BEG[5] ,
    \Tile_X5Y6_EE4BEG[4] ,
    \Tile_X5Y6_EE4BEG[3] ,
    \Tile_X5Y6_EE4BEG[2] ,
    \Tile_X5Y6_EE4BEG[1] ,
    \Tile_X5Y6_EE4BEG[0] }),
    .EE4END({\Tile_X4Y6_EE4BEG[15] ,
    \Tile_X4Y6_EE4BEG[14] ,
    \Tile_X4Y6_EE4BEG[13] ,
    \Tile_X4Y6_EE4BEG[12] ,
    \Tile_X4Y6_EE4BEG[11] ,
    \Tile_X4Y6_EE4BEG[10] ,
    \Tile_X4Y6_EE4BEG[9] ,
    \Tile_X4Y6_EE4BEG[8] ,
    \Tile_X4Y6_EE4BEG[7] ,
    \Tile_X4Y6_EE4BEG[6] ,
    \Tile_X4Y6_EE4BEG[5] ,
    \Tile_X4Y6_EE4BEG[4] ,
    \Tile_X4Y6_EE4BEG[3] ,
    \Tile_X4Y6_EE4BEG[2] ,
    \Tile_X4Y6_EE4BEG[1] ,
    \Tile_X4Y6_EE4BEG[0] }),
    .FrameData({\Tile_X4Y6_FrameData_O[31] ,
    \Tile_X4Y6_FrameData_O[30] ,
    \Tile_X4Y6_FrameData_O[29] ,
    \Tile_X4Y6_FrameData_O[28] ,
    \Tile_X4Y6_FrameData_O[27] ,
    \Tile_X4Y6_FrameData_O[26] ,
    \Tile_X4Y6_FrameData_O[25] ,
    \Tile_X4Y6_FrameData_O[24] ,
    \Tile_X4Y6_FrameData_O[23] ,
    \Tile_X4Y6_FrameData_O[22] ,
    \Tile_X4Y6_FrameData_O[21] ,
    \Tile_X4Y6_FrameData_O[20] ,
    \Tile_X4Y6_FrameData_O[19] ,
    \Tile_X4Y6_FrameData_O[18] ,
    \Tile_X4Y6_FrameData_O[17] ,
    \Tile_X4Y6_FrameData_O[16] ,
    \Tile_X4Y6_FrameData_O[15] ,
    \Tile_X4Y6_FrameData_O[14] ,
    \Tile_X4Y6_FrameData_O[13] ,
    \Tile_X4Y6_FrameData_O[12] ,
    \Tile_X4Y6_FrameData_O[11] ,
    \Tile_X4Y6_FrameData_O[10] ,
    \Tile_X4Y6_FrameData_O[9] ,
    \Tile_X4Y6_FrameData_O[8] ,
    \Tile_X4Y6_FrameData_O[7] ,
    \Tile_X4Y6_FrameData_O[6] ,
    \Tile_X4Y6_FrameData_O[5] ,
    \Tile_X4Y6_FrameData_O[4] ,
    \Tile_X4Y6_FrameData_O[3] ,
    \Tile_X4Y6_FrameData_O[2] ,
    \Tile_X4Y6_FrameData_O[1] ,
    \Tile_X4Y6_FrameData_O[0] }),
    .FrameData_O({\Tile_X5Y6_FrameData_O[31] ,
    \Tile_X5Y6_FrameData_O[30] ,
    \Tile_X5Y6_FrameData_O[29] ,
    \Tile_X5Y6_FrameData_O[28] ,
    \Tile_X5Y6_FrameData_O[27] ,
    \Tile_X5Y6_FrameData_O[26] ,
    \Tile_X5Y6_FrameData_O[25] ,
    \Tile_X5Y6_FrameData_O[24] ,
    \Tile_X5Y6_FrameData_O[23] ,
    \Tile_X5Y6_FrameData_O[22] ,
    \Tile_X5Y6_FrameData_O[21] ,
    \Tile_X5Y6_FrameData_O[20] ,
    \Tile_X5Y6_FrameData_O[19] ,
    \Tile_X5Y6_FrameData_O[18] ,
    \Tile_X5Y6_FrameData_O[17] ,
    \Tile_X5Y6_FrameData_O[16] ,
    \Tile_X5Y6_FrameData_O[15] ,
    \Tile_X5Y6_FrameData_O[14] ,
    \Tile_X5Y6_FrameData_O[13] ,
    \Tile_X5Y6_FrameData_O[12] ,
    \Tile_X5Y6_FrameData_O[11] ,
    \Tile_X5Y6_FrameData_O[10] ,
    \Tile_X5Y6_FrameData_O[9] ,
    \Tile_X5Y6_FrameData_O[8] ,
    \Tile_X5Y6_FrameData_O[7] ,
    \Tile_X5Y6_FrameData_O[6] ,
    \Tile_X5Y6_FrameData_O[5] ,
    \Tile_X5Y6_FrameData_O[4] ,
    \Tile_X5Y6_FrameData_O[3] ,
    \Tile_X5Y6_FrameData_O[2] ,
    \Tile_X5Y6_FrameData_O[1] ,
    \Tile_X5Y6_FrameData_O[0] }),
    .FrameStrobe({\Tile_X5Y7_FrameStrobe_O[19] ,
    \Tile_X5Y7_FrameStrobe_O[18] ,
    \Tile_X5Y7_FrameStrobe_O[17] ,
    \Tile_X5Y7_FrameStrobe_O[16] ,
    \Tile_X5Y7_FrameStrobe_O[15] ,
    \Tile_X5Y7_FrameStrobe_O[14] ,
    \Tile_X5Y7_FrameStrobe_O[13] ,
    \Tile_X5Y7_FrameStrobe_O[12] ,
    \Tile_X5Y7_FrameStrobe_O[11] ,
    \Tile_X5Y7_FrameStrobe_O[10] ,
    \Tile_X5Y7_FrameStrobe_O[9] ,
    \Tile_X5Y7_FrameStrobe_O[8] ,
    \Tile_X5Y7_FrameStrobe_O[7] ,
    \Tile_X5Y7_FrameStrobe_O[6] ,
    \Tile_X5Y7_FrameStrobe_O[5] ,
    \Tile_X5Y7_FrameStrobe_O[4] ,
    \Tile_X5Y7_FrameStrobe_O[3] ,
    \Tile_X5Y7_FrameStrobe_O[2] ,
    \Tile_X5Y7_FrameStrobe_O[1] ,
    \Tile_X5Y7_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X5Y6_FrameStrobe_O[19] ,
    \Tile_X5Y6_FrameStrobe_O[18] ,
    \Tile_X5Y6_FrameStrobe_O[17] ,
    \Tile_X5Y6_FrameStrobe_O[16] ,
    \Tile_X5Y6_FrameStrobe_O[15] ,
    \Tile_X5Y6_FrameStrobe_O[14] ,
    \Tile_X5Y6_FrameStrobe_O[13] ,
    \Tile_X5Y6_FrameStrobe_O[12] ,
    \Tile_X5Y6_FrameStrobe_O[11] ,
    \Tile_X5Y6_FrameStrobe_O[10] ,
    \Tile_X5Y6_FrameStrobe_O[9] ,
    \Tile_X5Y6_FrameStrobe_O[8] ,
    \Tile_X5Y6_FrameStrobe_O[7] ,
    \Tile_X5Y6_FrameStrobe_O[6] ,
    \Tile_X5Y6_FrameStrobe_O[5] ,
    \Tile_X5Y6_FrameStrobe_O[4] ,
    \Tile_X5Y6_FrameStrobe_O[3] ,
    \Tile_X5Y6_FrameStrobe_O[2] ,
    \Tile_X5Y6_FrameStrobe_O[1] ,
    \Tile_X5Y6_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X5Y6_N1BEG[3] ,
    \Tile_X5Y6_N1BEG[2] ,
    \Tile_X5Y6_N1BEG[1] ,
    \Tile_X5Y6_N1BEG[0] }),
    .N1END({\Tile_X5Y7_N1BEG[3] ,
    \Tile_X5Y7_N1BEG[2] ,
    \Tile_X5Y7_N1BEG[1] ,
    \Tile_X5Y7_N1BEG[0] }),
    .N2BEG({\Tile_X5Y6_N2BEG[7] ,
    \Tile_X5Y6_N2BEG[6] ,
    \Tile_X5Y6_N2BEG[5] ,
    \Tile_X5Y6_N2BEG[4] ,
    \Tile_X5Y6_N2BEG[3] ,
    \Tile_X5Y6_N2BEG[2] ,
    \Tile_X5Y6_N2BEG[1] ,
    \Tile_X5Y6_N2BEG[0] }),
    .N2BEGb({\Tile_X5Y6_N2BEGb[7] ,
    \Tile_X5Y6_N2BEGb[6] ,
    \Tile_X5Y6_N2BEGb[5] ,
    \Tile_X5Y6_N2BEGb[4] ,
    \Tile_X5Y6_N2BEGb[3] ,
    \Tile_X5Y6_N2BEGb[2] ,
    \Tile_X5Y6_N2BEGb[1] ,
    \Tile_X5Y6_N2BEGb[0] }),
    .N2END({\Tile_X5Y7_N2BEGb[7] ,
    \Tile_X5Y7_N2BEGb[6] ,
    \Tile_X5Y7_N2BEGb[5] ,
    \Tile_X5Y7_N2BEGb[4] ,
    \Tile_X5Y7_N2BEGb[3] ,
    \Tile_X5Y7_N2BEGb[2] ,
    \Tile_X5Y7_N2BEGb[1] ,
    \Tile_X5Y7_N2BEGb[0] }),
    .N2MID({\Tile_X5Y7_N2BEG[7] ,
    \Tile_X5Y7_N2BEG[6] ,
    \Tile_X5Y7_N2BEG[5] ,
    \Tile_X5Y7_N2BEG[4] ,
    \Tile_X5Y7_N2BEG[3] ,
    \Tile_X5Y7_N2BEG[2] ,
    \Tile_X5Y7_N2BEG[1] ,
    \Tile_X5Y7_N2BEG[0] }),
    .N4BEG({\Tile_X5Y6_N4BEG[15] ,
    \Tile_X5Y6_N4BEG[14] ,
    \Tile_X5Y6_N4BEG[13] ,
    \Tile_X5Y6_N4BEG[12] ,
    \Tile_X5Y6_N4BEG[11] ,
    \Tile_X5Y6_N4BEG[10] ,
    \Tile_X5Y6_N4BEG[9] ,
    \Tile_X5Y6_N4BEG[8] ,
    \Tile_X5Y6_N4BEG[7] ,
    \Tile_X5Y6_N4BEG[6] ,
    \Tile_X5Y6_N4BEG[5] ,
    \Tile_X5Y6_N4BEG[4] ,
    \Tile_X5Y6_N4BEG[3] ,
    \Tile_X5Y6_N4BEG[2] ,
    \Tile_X5Y6_N4BEG[1] ,
    \Tile_X5Y6_N4BEG[0] }),
    .N4END({\Tile_X5Y7_N4BEG[15] ,
    \Tile_X5Y7_N4BEG[14] ,
    \Tile_X5Y7_N4BEG[13] ,
    \Tile_X5Y7_N4BEG[12] ,
    \Tile_X5Y7_N4BEG[11] ,
    \Tile_X5Y7_N4BEG[10] ,
    \Tile_X5Y7_N4BEG[9] ,
    \Tile_X5Y7_N4BEG[8] ,
    \Tile_X5Y7_N4BEG[7] ,
    \Tile_X5Y7_N4BEG[6] ,
    \Tile_X5Y7_N4BEG[5] ,
    \Tile_X5Y7_N4BEG[4] ,
    \Tile_X5Y7_N4BEG[3] ,
    \Tile_X5Y7_N4BEG[2] ,
    \Tile_X5Y7_N4BEG[1] ,
    \Tile_X5Y7_N4BEG[0] }),
    .NN4BEG({\Tile_X5Y6_NN4BEG[15] ,
    \Tile_X5Y6_NN4BEG[14] ,
    \Tile_X5Y6_NN4BEG[13] ,
    \Tile_X5Y6_NN4BEG[12] ,
    \Tile_X5Y6_NN4BEG[11] ,
    \Tile_X5Y6_NN4BEG[10] ,
    \Tile_X5Y6_NN4BEG[9] ,
    \Tile_X5Y6_NN4BEG[8] ,
    \Tile_X5Y6_NN4BEG[7] ,
    \Tile_X5Y6_NN4BEG[6] ,
    \Tile_X5Y6_NN4BEG[5] ,
    \Tile_X5Y6_NN4BEG[4] ,
    \Tile_X5Y6_NN4BEG[3] ,
    \Tile_X5Y6_NN4BEG[2] ,
    \Tile_X5Y6_NN4BEG[1] ,
    \Tile_X5Y6_NN4BEG[0] }),
    .NN4END({\Tile_X5Y7_NN4BEG[15] ,
    \Tile_X5Y7_NN4BEG[14] ,
    \Tile_X5Y7_NN4BEG[13] ,
    \Tile_X5Y7_NN4BEG[12] ,
    \Tile_X5Y7_NN4BEG[11] ,
    \Tile_X5Y7_NN4BEG[10] ,
    \Tile_X5Y7_NN4BEG[9] ,
    \Tile_X5Y7_NN4BEG[8] ,
    \Tile_X5Y7_NN4BEG[7] ,
    \Tile_X5Y7_NN4BEG[6] ,
    \Tile_X5Y7_NN4BEG[5] ,
    \Tile_X5Y7_NN4BEG[4] ,
    \Tile_X5Y7_NN4BEG[3] ,
    \Tile_X5Y7_NN4BEG[2] ,
    \Tile_X5Y7_NN4BEG[1] ,
    \Tile_X5Y7_NN4BEG[0] }),
    .S1BEG({\Tile_X5Y6_S1BEG[3] ,
    \Tile_X5Y6_S1BEG[2] ,
    \Tile_X5Y6_S1BEG[1] ,
    \Tile_X5Y6_S1BEG[0] }),
    .S1END({\Tile_X5Y5_S1BEG[3] ,
    \Tile_X5Y5_S1BEG[2] ,
    \Tile_X5Y5_S1BEG[1] ,
    \Tile_X5Y5_S1BEG[0] }),
    .S2BEG({\Tile_X5Y6_S2BEG[7] ,
    \Tile_X5Y6_S2BEG[6] ,
    \Tile_X5Y6_S2BEG[5] ,
    \Tile_X5Y6_S2BEG[4] ,
    \Tile_X5Y6_S2BEG[3] ,
    \Tile_X5Y6_S2BEG[2] ,
    \Tile_X5Y6_S2BEG[1] ,
    \Tile_X5Y6_S2BEG[0] }),
    .S2BEGb({\Tile_X5Y6_S2BEGb[7] ,
    \Tile_X5Y6_S2BEGb[6] ,
    \Tile_X5Y6_S2BEGb[5] ,
    \Tile_X5Y6_S2BEGb[4] ,
    \Tile_X5Y6_S2BEGb[3] ,
    \Tile_X5Y6_S2BEGb[2] ,
    \Tile_X5Y6_S2BEGb[1] ,
    \Tile_X5Y6_S2BEGb[0] }),
    .S2END({\Tile_X5Y5_S2BEGb[7] ,
    \Tile_X5Y5_S2BEGb[6] ,
    \Tile_X5Y5_S2BEGb[5] ,
    \Tile_X5Y5_S2BEGb[4] ,
    \Tile_X5Y5_S2BEGb[3] ,
    \Tile_X5Y5_S2BEGb[2] ,
    \Tile_X5Y5_S2BEGb[1] ,
    \Tile_X5Y5_S2BEGb[0] }),
    .S2MID({\Tile_X5Y5_S2BEG[7] ,
    \Tile_X5Y5_S2BEG[6] ,
    \Tile_X5Y5_S2BEG[5] ,
    \Tile_X5Y5_S2BEG[4] ,
    \Tile_X5Y5_S2BEG[3] ,
    \Tile_X5Y5_S2BEG[2] ,
    \Tile_X5Y5_S2BEG[1] ,
    \Tile_X5Y5_S2BEG[0] }),
    .S4BEG({\Tile_X5Y6_S4BEG[15] ,
    \Tile_X5Y6_S4BEG[14] ,
    \Tile_X5Y6_S4BEG[13] ,
    \Tile_X5Y6_S4BEG[12] ,
    \Tile_X5Y6_S4BEG[11] ,
    \Tile_X5Y6_S4BEG[10] ,
    \Tile_X5Y6_S4BEG[9] ,
    \Tile_X5Y6_S4BEG[8] ,
    \Tile_X5Y6_S4BEG[7] ,
    \Tile_X5Y6_S4BEG[6] ,
    \Tile_X5Y6_S4BEG[5] ,
    \Tile_X5Y6_S4BEG[4] ,
    \Tile_X5Y6_S4BEG[3] ,
    \Tile_X5Y6_S4BEG[2] ,
    \Tile_X5Y6_S4BEG[1] ,
    \Tile_X5Y6_S4BEG[0] }),
    .S4END({\Tile_X5Y5_S4BEG[15] ,
    \Tile_X5Y5_S4BEG[14] ,
    \Tile_X5Y5_S4BEG[13] ,
    \Tile_X5Y5_S4BEG[12] ,
    \Tile_X5Y5_S4BEG[11] ,
    \Tile_X5Y5_S4BEG[10] ,
    \Tile_X5Y5_S4BEG[9] ,
    \Tile_X5Y5_S4BEG[8] ,
    \Tile_X5Y5_S4BEG[7] ,
    \Tile_X5Y5_S4BEG[6] ,
    \Tile_X5Y5_S4BEG[5] ,
    \Tile_X5Y5_S4BEG[4] ,
    \Tile_X5Y5_S4BEG[3] ,
    \Tile_X5Y5_S4BEG[2] ,
    \Tile_X5Y5_S4BEG[1] ,
    \Tile_X5Y5_S4BEG[0] }),
    .SS4BEG({\Tile_X5Y6_SS4BEG[15] ,
    \Tile_X5Y6_SS4BEG[14] ,
    \Tile_X5Y6_SS4BEG[13] ,
    \Tile_X5Y6_SS4BEG[12] ,
    \Tile_X5Y6_SS4BEG[11] ,
    \Tile_X5Y6_SS4BEG[10] ,
    \Tile_X5Y6_SS4BEG[9] ,
    \Tile_X5Y6_SS4BEG[8] ,
    \Tile_X5Y6_SS4BEG[7] ,
    \Tile_X5Y6_SS4BEG[6] ,
    \Tile_X5Y6_SS4BEG[5] ,
    \Tile_X5Y6_SS4BEG[4] ,
    \Tile_X5Y6_SS4BEG[3] ,
    \Tile_X5Y6_SS4BEG[2] ,
    \Tile_X5Y6_SS4BEG[1] ,
    \Tile_X5Y6_SS4BEG[0] }),
    .SS4END({\Tile_X5Y5_SS4BEG[15] ,
    \Tile_X5Y5_SS4BEG[14] ,
    \Tile_X5Y5_SS4BEG[13] ,
    \Tile_X5Y5_SS4BEG[12] ,
    \Tile_X5Y5_SS4BEG[11] ,
    \Tile_X5Y5_SS4BEG[10] ,
    \Tile_X5Y5_SS4BEG[9] ,
    \Tile_X5Y5_SS4BEG[8] ,
    \Tile_X5Y5_SS4BEG[7] ,
    \Tile_X5Y5_SS4BEG[6] ,
    \Tile_X5Y5_SS4BEG[5] ,
    \Tile_X5Y5_SS4BEG[4] ,
    \Tile_X5Y5_SS4BEG[3] ,
    \Tile_X5Y5_SS4BEG[2] ,
    \Tile_X5Y5_SS4BEG[1] ,
    \Tile_X5Y5_SS4BEG[0] }),
    .W1BEG({\Tile_X5Y6_W1BEG[3] ,
    \Tile_X5Y6_W1BEG[2] ,
    \Tile_X5Y6_W1BEG[1] ,
    \Tile_X5Y6_W1BEG[0] }),
    .W1END({\Tile_X6Y6_W1BEG[3] ,
    \Tile_X6Y6_W1BEG[2] ,
    \Tile_X6Y6_W1BEG[1] ,
    \Tile_X6Y6_W1BEG[0] }),
    .W2BEG({\Tile_X5Y6_W2BEG[7] ,
    \Tile_X5Y6_W2BEG[6] ,
    \Tile_X5Y6_W2BEG[5] ,
    \Tile_X5Y6_W2BEG[4] ,
    \Tile_X5Y6_W2BEG[3] ,
    \Tile_X5Y6_W2BEG[2] ,
    \Tile_X5Y6_W2BEG[1] ,
    \Tile_X5Y6_W2BEG[0] }),
    .W2BEGb({\Tile_X5Y6_W2BEGb[7] ,
    \Tile_X5Y6_W2BEGb[6] ,
    \Tile_X5Y6_W2BEGb[5] ,
    \Tile_X5Y6_W2BEGb[4] ,
    \Tile_X5Y6_W2BEGb[3] ,
    \Tile_X5Y6_W2BEGb[2] ,
    \Tile_X5Y6_W2BEGb[1] ,
    \Tile_X5Y6_W2BEGb[0] }),
    .W2END({\Tile_X6Y6_W2BEGb[7] ,
    \Tile_X6Y6_W2BEGb[6] ,
    \Tile_X6Y6_W2BEGb[5] ,
    \Tile_X6Y6_W2BEGb[4] ,
    \Tile_X6Y6_W2BEGb[3] ,
    \Tile_X6Y6_W2BEGb[2] ,
    \Tile_X6Y6_W2BEGb[1] ,
    \Tile_X6Y6_W2BEGb[0] }),
    .W2MID({\Tile_X6Y6_W2BEG[7] ,
    \Tile_X6Y6_W2BEG[6] ,
    \Tile_X6Y6_W2BEG[5] ,
    \Tile_X6Y6_W2BEG[4] ,
    \Tile_X6Y6_W2BEG[3] ,
    \Tile_X6Y6_W2BEG[2] ,
    \Tile_X6Y6_W2BEG[1] ,
    \Tile_X6Y6_W2BEG[0] }),
    .W6BEG({\Tile_X5Y6_W6BEG[11] ,
    \Tile_X5Y6_W6BEG[10] ,
    \Tile_X5Y6_W6BEG[9] ,
    \Tile_X5Y6_W6BEG[8] ,
    \Tile_X5Y6_W6BEG[7] ,
    \Tile_X5Y6_W6BEG[6] ,
    \Tile_X5Y6_W6BEG[5] ,
    \Tile_X5Y6_W6BEG[4] ,
    \Tile_X5Y6_W6BEG[3] ,
    \Tile_X5Y6_W6BEG[2] ,
    \Tile_X5Y6_W6BEG[1] ,
    \Tile_X5Y6_W6BEG[0] }),
    .W6END({\Tile_X6Y6_W6BEG[11] ,
    \Tile_X6Y6_W6BEG[10] ,
    \Tile_X6Y6_W6BEG[9] ,
    \Tile_X6Y6_W6BEG[8] ,
    \Tile_X6Y6_W6BEG[7] ,
    \Tile_X6Y6_W6BEG[6] ,
    \Tile_X6Y6_W6BEG[5] ,
    \Tile_X6Y6_W6BEG[4] ,
    \Tile_X6Y6_W6BEG[3] ,
    \Tile_X6Y6_W6BEG[2] ,
    \Tile_X6Y6_W6BEG[1] ,
    \Tile_X6Y6_W6BEG[0] }),
    .WW4BEG({\Tile_X5Y6_WW4BEG[15] ,
    \Tile_X5Y6_WW4BEG[14] ,
    \Tile_X5Y6_WW4BEG[13] ,
    \Tile_X5Y6_WW4BEG[12] ,
    \Tile_X5Y6_WW4BEG[11] ,
    \Tile_X5Y6_WW4BEG[10] ,
    \Tile_X5Y6_WW4BEG[9] ,
    \Tile_X5Y6_WW4BEG[8] ,
    \Tile_X5Y6_WW4BEG[7] ,
    \Tile_X5Y6_WW4BEG[6] ,
    \Tile_X5Y6_WW4BEG[5] ,
    \Tile_X5Y6_WW4BEG[4] ,
    \Tile_X5Y6_WW4BEG[3] ,
    \Tile_X5Y6_WW4BEG[2] ,
    \Tile_X5Y6_WW4BEG[1] ,
    \Tile_X5Y6_WW4BEG[0] }),
    .WW4END({\Tile_X6Y6_WW4BEG[15] ,
    \Tile_X6Y6_WW4BEG[14] ,
    \Tile_X6Y6_WW4BEG[13] ,
    \Tile_X6Y6_WW4BEG[12] ,
    \Tile_X6Y6_WW4BEG[11] ,
    \Tile_X6Y6_WW4BEG[10] ,
    \Tile_X6Y6_WW4BEG[9] ,
    \Tile_X6Y6_WW4BEG[8] ,
    \Tile_X6Y6_WW4BEG[7] ,
    \Tile_X6Y6_WW4BEG[6] ,
    \Tile_X6Y6_WW4BEG[5] ,
    \Tile_X6Y6_WW4BEG[4] ,
    \Tile_X6Y6_WW4BEG[3] ,
    \Tile_X6Y6_WW4BEG[2] ,
    \Tile_X6Y6_WW4BEG[1] ,
    \Tile_X6Y6_WW4BEG[0] }));
 LUT4AB Tile_X5Y7_LUT4AB (.Ci(Tile_X5Y8_Co),
    .Co(Tile_X5Y7_Co),
    .UserCLK(Tile_X5Y8_UserCLKo),
    .UserCLKo(Tile_X5Y7_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X5Y7_E1BEG[3] ,
    \Tile_X5Y7_E1BEG[2] ,
    \Tile_X5Y7_E1BEG[1] ,
    \Tile_X5Y7_E1BEG[0] }),
    .E1END({\Tile_X4Y7_E1BEG[3] ,
    \Tile_X4Y7_E1BEG[2] ,
    \Tile_X4Y7_E1BEG[1] ,
    \Tile_X4Y7_E1BEG[0] }),
    .E2BEG({\Tile_X5Y7_E2BEG[7] ,
    \Tile_X5Y7_E2BEG[6] ,
    \Tile_X5Y7_E2BEG[5] ,
    \Tile_X5Y7_E2BEG[4] ,
    \Tile_X5Y7_E2BEG[3] ,
    \Tile_X5Y7_E2BEG[2] ,
    \Tile_X5Y7_E2BEG[1] ,
    \Tile_X5Y7_E2BEG[0] }),
    .E2BEGb({\Tile_X5Y7_E2BEGb[7] ,
    \Tile_X5Y7_E2BEGb[6] ,
    \Tile_X5Y7_E2BEGb[5] ,
    \Tile_X5Y7_E2BEGb[4] ,
    \Tile_X5Y7_E2BEGb[3] ,
    \Tile_X5Y7_E2BEGb[2] ,
    \Tile_X5Y7_E2BEGb[1] ,
    \Tile_X5Y7_E2BEGb[0] }),
    .E2END({\Tile_X4Y7_E2BEGb[7] ,
    \Tile_X4Y7_E2BEGb[6] ,
    \Tile_X4Y7_E2BEGb[5] ,
    \Tile_X4Y7_E2BEGb[4] ,
    \Tile_X4Y7_E2BEGb[3] ,
    \Tile_X4Y7_E2BEGb[2] ,
    \Tile_X4Y7_E2BEGb[1] ,
    \Tile_X4Y7_E2BEGb[0] }),
    .E2MID({\Tile_X4Y7_E2BEG[7] ,
    \Tile_X4Y7_E2BEG[6] ,
    \Tile_X4Y7_E2BEG[5] ,
    \Tile_X4Y7_E2BEG[4] ,
    \Tile_X4Y7_E2BEG[3] ,
    \Tile_X4Y7_E2BEG[2] ,
    \Tile_X4Y7_E2BEG[1] ,
    \Tile_X4Y7_E2BEG[0] }),
    .E6BEG({\Tile_X5Y7_E6BEG[11] ,
    \Tile_X5Y7_E6BEG[10] ,
    \Tile_X5Y7_E6BEG[9] ,
    \Tile_X5Y7_E6BEG[8] ,
    \Tile_X5Y7_E6BEG[7] ,
    \Tile_X5Y7_E6BEG[6] ,
    \Tile_X5Y7_E6BEG[5] ,
    \Tile_X5Y7_E6BEG[4] ,
    \Tile_X5Y7_E6BEG[3] ,
    \Tile_X5Y7_E6BEG[2] ,
    \Tile_X5Y7_E6BEG[1] ,
    \Tile_X5Y7_E6BEG[0] }),
    .E6END({\Tile_X4Y7_E6BEG[11] ,
    \Tile_X4Y7_E6BEG[10] ,
    \Tile_X4Y7_E6BEG[9] ,
    \Tile_X4Y7_E6BEG[8] ,
    \Tile_X4Y7_E6BEG[7] ,
    \Tile_X4Y7_E6BEG[6] ,
    \Tile_X4Y7_E6BEG[5] ,
    \Tile_X4Y7_E6BEG[4] ,
    \Tile_X4Y7_E6BEG[3] ,
    \Tile_X4Y7_E6BEG[2] ,
    \Tile_X4Y7_E6BEG[1] ,
    \Tile_X4Y7_E6BEG[0] }),
    .EE4BEG({\Tile_X5Y7_EE4BEG[15] ,
    \Tile_X5Y7_EE4BEG[14] ,
    \Tile_X5Y7_EE4BEG[13] ,
    \Tile_X5Y7_EE4BEG[12] ,
    \Tile_X5Y7_EE4BEG[11] ,
    \Tile_X5Y7_EE4BEG[10] ,
    \Tile_X5Y7_EE4BEG[9] ,
    \Tile_X5Y7_EE4BEG[8] ,
    \Tile_X5Y7_EE4BEG[7] ,
    \Tile_X5Y7_EE4BEG[6] ,
    \Tile_X5Y7_EE4BEG[5] ,
    \Tile_X5Y7_EE4BEG[4] ,
    \Tile_X5Y7_EE4BEG[3] ,
    \Tile_X5Y7_EE4BEG[2] ,
    \Tile_X5Y7_EE4BEG[1] ,
    \Tile_X5Y7_EE4BEG[0] }),
    .EE4END({\Tile_X4Y7_EE4BEG[15] ,
    \Tile_X4Y7_EE4BEG[14] ,
    \Tile_X4Y7_EE4BEG[13] ,
    \Tile_X4Y7_EE4BEG[12] ,
    \Tile_X4Y7_EE4BEG[11] ,
    \Tile_X4Y7_EE4BEG[10] ,
    \Tile_X4Y7_EE4BEG[9] ,
    \Tile_X4Y7_EE4BEG[8] ,
    \Tile_X4Y7_EE4BEG[7] ,
    \Tile_X4Y7_EE4BEG[6] ,
    \Tile_X4Y7_EE4BEG[5] ,
    \Tile_X4Y7_EE4BEG[4] ,
    \Tile_X4Y7_EE4BEG[3] ,
    \Tile_X4Y7_EE4BEG[2] ,
    \Tile_X4Y7_EE4BEG[1] ,
    \Tile_X4Y7_EE4BEG[0] }),
    .FrameData({\Tile_X4Y7_FrameData_O[31] ,
    \Tile_X4Y7_FrameData_O[30] ,
    \Tile_X4Y7_FrameData_O[29] ,
    \Tile_X4Y7_FrameData_O[28] ,
    \Tile_X4Y7_FrameData_O[27] ,
    \Tile_X4Y7_FrameData_O[26] ,
    \Tile_X4Y7_FrameData_O[25] ,
    \Tile_X4Y7_FrameData_O[24] ,
    \Tile_X4Y7_FrameData_O[23] ,
    \Tile_X4Y7_FrameData_O[22] ,
    \Tile_X4Y7_FrameData_O[21] ,
    \Tile_X4Y7_FrameData_O[20] ,
    \Tile_X4Y7_FrameData_O[19] ,
    \Tile_X4Y7_FrameData_O[18] ,
    \Tile_X4Y7_FrameData_O[17] ,
    \Tile_X4Y7_FrameData_O[16] ,
    \Tile_X4Y7_FrameData_O[15] ,
    \Tile_X4Y7_FrameData_O[14] ,
    \Tile_X4Y7_FrameData_O[13] ,
    \Tile_X4Y7_FrameData_O[12] ,
    \Tile_X4Y7_FrameData_O[11] ,
    \Tile_X4Y7_FrameData_O[10] ,
    \Tile_X4Y7_FrameData_O[9] ,
    \Tile_X4Y7_FrameData_O[8] ,
    \Tile_X4Y7_FrameData_O[7] ,
    \Tile_X4Y7_FrameData_O[6] ,
    \Tile_X4Y7_FrameData_O[5] ,
    \Tile_X4Y7_FrameData_O[4] ,
    \Tile_X4Y7_FrameData_O[3] ,
    \Tile_X4Y7_FrameData_O[2] ,
    \Tile_X4Y7_FrameData_O[1] ,
    \Tile_X4Y7_FrameData_O[0] }),
    .FrameData_O({\Tile_X5Y7_FrameData_O[31] ,
    \Tile_X5Y7_FrameData_O[30] ,
    \Tile_X5Y7_FrameData_O[29] ,
    \Tile_X5Y7_FrameData_O[28] ,
    \Tile_X5Y7_FrameData_O[27] ,
    \Tile_X5Y7_FrameData_O[26] ,
    \Tile_X5Y7_FrameData_O[25] ,
    \Tile_X5Y7_FrameData_O[24] ,
    \Tile_X5Y7_FrameData_O[23] ,
    \Tile_X5Y7_FrameData_O[22] ,
    \Tile_X5Y7_FrameData_O[21] ,
    \Tile_X5Y7_FrameData_O[20] ,
    \Tile_X5Y7_FrameData_O[19] ,
    \Tile_X5Y7_FrameData_O[18] ,
    \Tile_X5Y7_FrameData_O[17] ,
    \Tile_X5Y7_FrameData_O[16] ,
    \Tile_X5Y7_FrameData_O[15] ,
    \Tile_X5Y7_FrameData_O[14] ,
    \Tile_X5Y7_FrameData_O[13] ,
    \Tile_X5Y7_FrameData_O[12] ,
    \Tile_X5Y7_FrameData_O[11] ,
    \Tile_X5Y7_FrameData_O[10] ,
    \Tile_X5Y7_FrameData_O[9] ,
    \Tile_X5Y7_FrameData_O[8] ,
    \Tile_X5Y7_FrameData_O[7] ,
    \Tile_X5Y7_FrameData_O[6] ,
    \Tile_X5Y7_FrameData_O[5] ,
    \Tile_X5Y7_FrameData_O[4] ,
    \Tile_X5Y7_FrameData_O[3] ,
    \Tile_X5Y7_FrameData_O[2] ,
    \Tile_X5Y7_FrameData_O[1] ,
    \Tile_X5Y7_FrameData_O[0] }),
    .FrameStrobe({\Tile_X5Y8_FrameStrobe_O[19] ,
    \Tile_X5Y8_FrameStrobe_O[18] ,
    \Tile_X5Y8_FrameStrobe_O[17] ,
    \Tile_X5Y8_FrameStrobe_O[16] ,
    \Tile_X5Y8_FrameStrobe_O[15] ,
    \Tile_X5Y8_FrameStrobe_O[14] ,
    \Tile_X5Y8_FrameStrobe_O[13] ,
    \Tile_X5Y8_FrameStrobe_O[12] ,
    \Tile_X5Y8_FrameStrobe_O[11] ,
    \Tile_X5Y8_FrameStrobe_O[10] ,
    \Tile_X5Y8_FrameStrobe_O[9] ,
    \Tile_X5Y8_FrameStrobe_O[8] ,
    \Tile_X5Y8_FrameStrobe_O[7] ,
    \Tile_X5Y8_FrameStrobe_O[6] ,
    \Tile_X5Y8_FrameStrobe_O[5] ,
    \Tile_X5Y8_FrameStrobe_O[4] ,
    \Tile_X5Y8_FrameStrobe_O[3] ,
    \Tile_X5Y8_FrameStrobe_O[2] ,
    \Tile_X5Y8_FrameStrobe_O[1] ,
    \Tile_X5Y8_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X5Y7_FrameStrobe_O[19] ,
    \Tile_X5Y7_FrameStrobe_O[18] ,
    \Tile_X5Y7_FrameStrobe_O[17] ,
    \Tile_X5Y7_FrameStrobe_O[16] ,
    \Tile_X5Y7_FrameStrobe_O[15] ,
    \Tile_X5Y7_FrameStrobe_O[14] ,
    \Tile_X5Y7_FrameStrobe_O[13] ,
    \Tile_X5Y7_FrameStrobe_O[12] ,
    \Tile_X5Y7_FrameStrobe_O[11] ,
    \Tile_X5Y7_FrameStrobe_O[10] ,
    \Tile_X5Y7_FrameStrobe_O[9] ,
    \Tile_X5Y7_FrameStrobe_O[8] ,
    \Tile_X5Y7_FrameStrobe_O[7] ,
    \Tile_X5Y7_FrameStrobe_O[6] ,
    \Tile_X5Y7_FrameStrobe_O[5] ,
    \Tile_X5Y7_FrameStrobe_O[4] ,
    \Tile_X5Y7_FrameStrobe_O[3] ,
    \Tile_X5Y7_FrameStrobe_O[2] ,
    \Tile_X5Y7_FrameStrobe_O[1] ,
    \Tile_X5Y7_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X5Y7_N1BEG[3] ,
    \Tile_X5Y7_N1BEG[2] ,
    \Tile_X5Y7_N1BEG[1] ,
    \Tile_X5Y7_N1BEG[0] }),
    .N1END({\Tile_X5Y8_N1BEG[3] ,
    \Tile_X5Y8_N1BEG[2] ,
    \Tile_X5Y8_N1BEG[1] ,
    \Tile_X5Y8_N1BEG[0] }),
    .N2BEG({\Tile_X5Y7_N2BEG[7] ,
    \Tile_X5Y7_N2BEG[6] ,
    \Tile_X5Y7_N2BEG[5] ,
    \Tile_X5Y7_N2BEG[4] ,
    \Tile_X5Y7_N2BEG[3] ,
    \Tile_X5Y7_N2BEG[2] ,
    \Tile_X5Y7_N2BEG[1] ,
    \Tile_X5Y7_N2BEG[0] }),
    .N2BEGb({\Tile_X5Y7_N2BEGb[7] ,
    \Tile_X5Y7_N2BEGb[6] ,
    \Tile_X5Y7_N2BEGb[5] ,
    \Tile_X5Y7_N2BEGb[4] ,
    \Tile_X5Y7_N2BEGb[3] ,
    \Tile_X5Y7_N2BEGb[2] ,
    \Tile_X5Y7_N2BEGb[1] ,
    \Tile_X5Y7_N2BEGb[0] }),
    .N2END({\Tile_X5Y8_N2BEGb[7] ,
    \Tile_X5Y8_N2BEGb[6] ,
    \Tile_X5Y8_N2BEGb[5] ,
    \Tile_X5Y8_N2BEGb[4] ,
    \Tile_X5Y8_N2BEGb[3] ,
    \Tile_X5Y8_N2BEGb[2] ,
    \Tile_X5Y8_N2BEGb[1] ,
    \Tile_X5Y8_N2BEGb[0] }),
    .N2MID({\Tile_X5Y8_N2BEG[7] ,
    \Tile_X5Y8_N2BEG[6] ,
    \Tile_X5Y8_N2BEG[5] ,
    \Tile_X5Y8_N2BEG[4] ,
    \Tile_X5Y8_N2BEG[3] ,
    \Tile_X5Y8_N2BEG[2] ,
    \Tile_X5Y8_N2BEG[1] ,
    \Tile_X5Y8_N2BEG[0] }),
    .N4BEG({\Tile_X5Y7_N4BEG[15] ,
    \Tile_X5Y7_N4BEG[14] ,
    \Tile_X5Y7_N4BEG[13] ,
    \Tile_X5Y7_N4BEG[12] ,
    \Tile_X5Y7_N4BEG[11] ,
    \Tile_X5Y7_N4BEG[10] ,
    \Tile_X5Y7_N4BEG[9] ,
    \Tile_X5Y7_N4BEG[8] ,
    \Tile_X5Y7_N4BEG[7] ,
    \Tile_X5Y7_N4BEG[6] ,
    \Tile_X5Y7_N4BEG[5] ,
    \Tile_X5Y7_N4BEG[4] ,
    \Tile_X5Y7_N4BEG[3] ,
    \Tile_X5Y7_N4BEG[2] ,
    \Tile_X5Y7_N4BEG[1] ,
    \Tile_X5Y7_N4BEG[0] }),
    .N4END({\Tile_X5Y8_N4BEG[15] ,
    \Tile_X5Y8_N4BEG[14] ,
    \Tile_X5Y8_N4BEG[13] ,
    \Tile_X5Y8_N4BEG[12] ,
    \Tile_X5Y8_N4BEG[11] ,
    \Tile_X5Y8_N4BEG[10] ,
    \Tile_X5Y8_N4BEG[9] ,
    \Tile_X5Y8_N4BEG[8] ,
    \Tile_X5Y8_N4BEG[7] ,
    \Tile_X5Y8_N4BEG[6] ,
    \Tile_X5Y8_N4BEG[5] ,
    \Tile_X5Y8_N4BEG[4] ,
    \Tile_X5Y8_N4BEG[3] ,
    \Tile_X5Y8_N4BEG[2] ,
    \Tile_X5Y8_N4BEG[1] ,
    \Tile_X5Y8_N4BEG[0] }),
    .NN4BEG({\Tile_X5Y7_NN4BEG[15] ,
    \Tile_X5Y7_NN4BEG[14] ,
    \Tile_X5Y7_NN4BEG[13] ,
    \Tile_X5Y7_NN4BEG[12] ,
    \Tile_X5Y7_NN4BEG[11] ,
    \Tile_X5Y7_NN4BEG[10] ,
    \Tile_X5Y7_NN4BEG[9] ,
    \Tile_X5Y7_NN4BEG[8] ,
    \Tile_X5Y7_NN4BEG[7] ,
    \Tile_X5Y7_NN4BEG[6] ,
    \Tile_X5Y7_NN4BEG[5] ,
    \Tile_X5Y7_NN4BEG[4] ,
    \Tile_X5Y7_NN4BEG[3] ,
    \Tile_X5Y7_NN4BEG[2] ,
    \Tile_X5Y7_NN4BEG[1] ,
    \Tile_X5Y7_NN4BEG[0] }),
    .NN4END({\Tile_X5Y8_NN4BEG[15] ,
    \Tile_X5Y8_NN4BEG[14] ,
    \Tile_X5Y8_NN4BEG[13] ,
    \Tile_X5Y8_NN4BEG[12] ,
    \Tile_X5Y8_NN4BEG[11] ,
    \Tile_X5Y8_NN4BEG[10] ,
    \Tile_X5Y8_NN4BEG[9] ,
    \Tile_X5Y8_NN4BEG[8] ,
    \Tile_X5Y8_NN4BEG[7] ,
    \Tile_X5Y8_NN4BEG[6] ,
    \Tile_X5Y8_NN4BEG[5] ,
    \Tile_X5Y8_NN4BEG[4] ,
    \Tile_X5Y8_NN4BEG[3] ,
    \Tile_X5Y8_NN4BEG[2] ,
    \Tile_X5Y8_NN4BEG[1] ,
    \Tile_X5Y8_NN4BEG[0] }),
    .S1BEG({\Tile_X5Y7_S1BEG[3] ,
    \Tile_X5Y7_S1BEG[2] ,
    \Tile_X5Y7_S1BEG[1] ,
    \Tile_X5Y7_S1BEG[0] }),
    .S1END({\Tile_X5Y6_S1BEG[3] ,
    \Tile_X5Y6_S1BEG[2] ,
    \Tile_X5Y6_S1BEG[1] ,
    \Tile_X5Y6_S1BEG[0] }),
    .S2BEG({\Tile_X5Y7_S2BEG[7] ,
    \Tile_X5Y7_S2BEG[6] ,
    \Tile_X5Y7_S2BEG[5] ,
    \Tile_X5Y7_S2BEG[4] ,
    \Tile_X5Y7_S2BEG[3] ,
    \Tile_X5Y7_S2BEG[2] ,
    \Tile_X5Y7_S2BEG[1] ,
    \Tile_X5Y7_S2BEG[0] }),
    .S2BEGb({\Tile_X5Y7_S2BEGb[7] ,
    \Tile_X5Y7_S2BEGb[6] ,
    \Tile_X5Y7_S2BEGb[5] ,
    \Tile_X5Y7_S2BEGb[4] ,
    \Tile_X5Y7_S2BEGb[3] ,
    \Tile_X5Y7_S2BEGb[2] ,
    \Tile_X5Y7_S2BEGb[1] ,
    \Tile_X5Y7_S2BEGb[0] }),
    .S2END({\Tile_X5Y6_S2BEGb[7] ,
    \Tile_X5Y6_S2BEGb[6] ,
    \Tile_X5Y6_S2BEGb[5] ,
    \Tile_X5Y6_S2BEGb[4] ,
    \Tile_X5Y6_S2BEGb[3] ,
    \Tile_X5Y6_S2BEGb[2] ,
    \Tile_X5Y6_S2BEGb[1] ,
    \Tile_X5Y6_S2BEGb[0] }),
    .S2MID({\Tile_X5Y6_S2BEG[7] ,
    \Tile_X5Y6_S2BEG[6] ,
    \Tile_X5Y6_S2BEG[5] ,
    \Tile_X5Y6_S2BEG[4] ,
    \Tile_X5Y6_S2BEG[3] ,
    \Tile_X5Y6_S2BEG[2] ,
    \Tile_X5Y6_S2BEG[1] ,
    \Tile_X5Y6_S2BEG[0] }),
    .S4BEG({\Tile_X5Y7_S4BEG[15] ,
    \Tile_X5Y7_S4BEG[14] ,
    \Tile_X5Y7_S4BEG[13] ,
    \Tile_X5Y7_S4BEG[12] ,
    \Tile_X5Y7_S4BEG[11] ,
    \Tile_X5Y7_S4BEG[10] ,
    \Tile_X5Y7_S4BEG[9] ,
    \Tile_X5Y7_S4BEG[8] ,
    \Tile_X5Y7_S4BEG[7] ,
    \Tile_X5Y7_S4BEG[6] ,
    \Tile_X5Y7_S4BEG[5] ,
    \Tile_X5Y7_S4BEG[4] ,
    \Tile_X5Y7_S4BEG[3] ,
    \Tile_X5Y7_S4BEG[2] ,
    \Tile_X5Y7_S4BEG[1] ,
    \Tile_X5Y7_S4BEG[0] }),
    .S4END({\Tile_X5Y6_S4BEG[15] ,
    \Tile_X5Y6_S4BEG[14] ,
    \Tile_X5Y6_S4BEG[13] ,
    \Tile_X5Y6_S4BEG[12] ,
    \Tile_X5Y6_S4BEG[11] ,
    \Tile_X5Y6_S4BEG[10] ,
    \Tile_X5Y6_S4BEG[9] ,
    \Tile_X5Y6_S4BEG[8] ,
    \Tile_X5Y6_S4BEG[7] ,
    \Tile_X5Y6_S4BEG[6] ,
    \Tile_X5Y6_S4BEG[5] ,
    \Tile_X5Y6_S4BEG[4] ,
    \Tile_X5Y6_S4BEG[3] ,
    \Tile_X5Y6_S4BEG[2] ,
    \Tile_X5Y6_S4BEG[1] ,
    \Tile_X5Y6_S4BEG[0] }),
    .SS4BEG({\Tile_X5Y7_SS4BEG[15] ,
    \Tile_X5Y7_SS4BEG[14] ,
    \Tile_X5Y7_SS4BEG[13] ,
    \Tile_X5Y7_SS4BEG[12] ,
    \Tile_X5Y7_SS4BEG[11] ,
    \Tile_X5Y7_SS4BEG[10] ,
    \Tile_X5Y7_SS4BEG[9] ,
    \Tile_X5Y7_SS4BEG[8] ,
    \Tile_X5Y7_SS4BEG[7] ,
    \Tile_X5Y7_SS4BEG[6] ,
    \Tile_X5Y7_SS4BEG[5] ,
    \Tile_X5Y7_SS4BEG[4] ,
    \Tile_X5Y7_SS4BEG[3] ,
    \Tile_X5Y7_SS4BEG[2] ,
    \Tile_X5Y7_SS4BEG[1] ,
    \Tile_X5Y7_SS4BEG[0] }),
    .SS4END({\Tile_X5Y6_SS4BEG[15] ,
    \Tile_X5Y6_SS4BEG[14] ,
    \Tile_X5Y6_SS4BEG[13] ,
    \Tile_X5Y6_SS4BEG[12] ,
    \Tile_X5Y6_SS4BEG[11] ,
    \Tile_X5Y6_SS4BEG[10] ,
    \Tile_X5Y6_SS4BEG[9] ,
    \Tile_X5Y6_SS4BEG[8] ,
    \Tile_X5Y6_SS4BEG[7] ,
    \Tile_X5Y6_SS4BEG[6] ,
    \Tile_X5Y6_SS4BEG[5] ,
    \Tile_X5Y6_SS4BEG[4] ,
    \Tile_X5Y6_SS4BEG[3] ,
    \Tile_X5Y6_SS4BEG[2] ,
    \Tile_X5Y6_SS4BEG[1] ,
    \Tile_X5Y6_SS4BEG[0] }),
    .W1BEG({\Tile_X5Y7_W1BEG[3] ,
    \Tile_X5Y7_W1BEG[2] ,
    \Tile_X5Y7_W1BEG[1] ,
    \Tile_X5Y7_W1BEG[0] }),
    .W1END({\Tile_X6Y7_W1BEG[3] ,
    \Tile_X6Y7_W1BEG[2] ,
    \Tile_X6Y7_W1BEG[1] ,
    \Tile_X6Y7_W1BEG[0] }),
    .W2BEG({\Tile_X5Y7_W2BEG[7] ,
    \Tile_X5Y7_W2BEG[6] ,
    \Tile_X5Y7_W2BEG[5] ,
    \Tile_X5Y7_W2BEG[4] ,
    \Tile_X5Y7_W2BEG[3] ,
    \Tile_X5Y7_W2BEG[2] ,
    \Tile_X5Y7_W2BEG[1] ,
    \Tile_X5Y7_W2BEG[0] }),
    .W2BEGb({\Tile_X5Y7_W2BEGb[7] ,
    \Tile_X5Y7_W2BEGb[6] ,
    \Tile_X5Y7_W2BEGb[5] ,
    \Tile_X5Y7_W2BEGb[4] ,
    \Tile_X5Y7_W2BEGb[3] ,
    \Tile_X5Y7_W2BEGb[2] ,
    \Tile_X5Y7_W2BEGb[1] ,
    \Tile_X5Y7_W2BEGb[0] }),
    .W2END({\Tile_X6Y7_W2BEGb[7] ,
    \Tile_X6Y7_W2BEGb[6] ,
    \Tile_X6Y7_W2BEGb[5] ,
    \Tile_X6Y7_W2BEGb[4] ,
    \Tile_X6Y7_W2BEGb[3] ,
    \Tile_X6Y7_W2BEGb[2] ,
    \Tile_X6Y7_W2BEGb[1] ,
    \Tile_X6Y7_W2BEGb[0] }),
    .W2MID({\Tile_X6Y7_W2BEG[7] ,
    \Tile_X6Y7_W2BEG[6] ,
    \Tile_X6Y7_W2BEG[5] ,
    \Tile_X6Y7_W2BEG[4] ,
    \Tile_X6Y7_W2BEG[3] ,
    \Tile_X6Y7_W2BEG[2] ,
    \Tile_X6Y7_W2BEG[1] ,
    \Tile_X6Y7_W2BEG[0] }),
    .W6BEG({\Tile_X5Y7_W6BEG[11] ,
    \Tile_X5Y7_W6BEG[10] ,
    \Tile_X5Y7_W6BEG[9] ,
    \Tile_X5Y7_W6BEG[8] ,
    \Tile_X5Y7_W6BEG[7] ,
    \Tile_X5Y7_W6BEG[6] ,
    \Tile_X5Y7_W6BEG[5] ,
    \Tile_X5Y7_W6BEG[4] ,
    \Tile_X5Y7_W6BEG[3] ,
    \Tile_X5Y7_W6BEG[2] ,
    \Tile_X5Y7_W6BEG[1] ,
    \Tile_X5Y7_W6BEG[0] }),
    .W6END({\Tile_X6Y7_W6BEG[11] ,
    \Tile_X6Y7_W6BEG[10] ,
    \Tile_X6Y7_W6BEG[9] ,
    \Tile_X6Y7_W6BEG[8] ,
    \Tile_X6Y7_W6BEG[7] ,
    \Tile_X6Y7_W6BEG[6] ,
    \Tile_X6Y7_W6BEG[5] ,
    \Tile_X6Y7_W6BEG[4] ,
    \Tile_X6Y7_W6BEG[3] ,
    \Tile_X6Y7_W6BEG[2] ,
    \Tile_X6Y7_W6BEG[1] ,
    \Tile_X6Y7_W6BEG[0] }),
    .WW4BEG({\Tile_X5Y7_WW4BEG[15] ,
    \Tile_X5Y7_WW4BEG[14] ,
    \Tile_X5Y7_WW4BEG[13] ,
    \Tile_X5Y7_WW4BEG[12] ,
    \Tile_X5Y7_WW4BEG[11] ,
    \Tile_X5Y7_WW4BEG[10] ,
    \Tile_X5Y7_WW4BEG[9] ,
    \Tile_X5Y7_WW4BEG[8] ,
    \Tile_X5Y7_WW4BEG[7] ,
    \Tile_X5Y7_WW4BEG[6] ,
    \Tile_X5Y7_WW4BEG[5] ,
    \Tile_X5Y7_WW4BEG[4] ,
    \Tile_X5Y7_WW4BEG[3] ,
    \Tile_X5Y7_WW4BEG[2] ,
    \Tile_X5Y7_WW4BEG[1] ,
    \Tile_X5Y7_WW4BEG[0] }),
    .WW4END({\Tile_X6Y7_WW4BEG[15] ,
    \Tile_X6Y7_WW4BEG[14] ,
    \Tile_X6Y7_WW4BEG[13] ,
    \Tile_X6Y7_WW4BEG[12] ,
    \Tile_X6Y7_WW4BEG[11] ,
    \Tile_X6Y7_WW4BEG[10] ,
    \Tile_X6Y7_WW4BEG[9] ,
    \Tile_X6Y7_WW4BEG[8] ,
    \Tile_X6Y7_WW4BEG[7] ,
    \Tile_X6Y7_WW4BEG[6] ,
    \Tile_X6Y7_WW4BEG[5] ,
    \Tile_X6Y7_WW4BEG[4] ,
    \Tile_X6Y7_WW4BEG[3] ,
    \Tile_X6Y7_WW4BEG[2] ,
    \Tile_X6Y7_WW4BEG[1] ,
    \Tile_X6Y7_WW4BEG[0] }));
 LUT4AB Tile_X5Y8_LUT4AB (.Ci(Tile_X5Y9_Co),
    .Co(Tile_X5Y8_Co),
    .UserCLK(Tile_X5Y9_UserCLKo),
    .UserCLKo(Tile_X5Y8_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X5Y8_E1BEG[3] ,
    \Tile_X5Y8_E1BEG[2] ,
    \Tile_X5Y8_E1BEG[1] ,
    \Tile_X5Y8_E1BEG[0] }),
    .E1END({\Tile_X4Y8_E1BEG[3] ,
    \Tile_X4Y8_E1BEG[2] ,
    \Tile_X4Y8_E1BEG[1] ,
    \Tile_X4Y8_E1BEG[0] }),
    .E2BEG({\Tile_X5Y8_E2BEG[7] ,
    \Tile_X5Y8_E2BEG[6] ,
    \Tile_X5Y8_E2BEG[5] ,
    \Tile_X5Y8_E2BEG[4] ,
    \Tile_X5Y8_E2BEG[3] ,
    \Tile_X5Y8_E2BEG[2] ,
    \Tile_X5Y8_E2BEG[1] ,
    \Tile_X5Y8_E2BEG[0] }),
    .E2BEGb({\Tile_X5Y8_E2BEGb[7] ,
    \Tile_X5Y8_E2BEGb[6] ,
    \Tile_X5Y8_E2BEGb[5] ,
    \Tile_X5Y8_E2BEGb[4] ,
    \Tile_X5Y8_E2BEGb[3] ,
    \Tile_X5Y8_E2BEGb[2] ,
    \Tile_X5Y8_E2BEGb[1] ,
    \Tile_X5Y8_E2BEGb[0] }),
    .E2END({\Tile_X4Y8_E2BEGb[7] ,
    \Tile_X4Y8_E2BEGb[6] ,
    \Tile_X4Y8_E2BEGb[5] ,
    \Tile_X4Y8_E2BEGb[4] ,
    \Tile_X4Y8_E2BEGb[3] ,
    \Tile_X4Y8_E2BEGb[2] ,
    \Tile_X4Y8_E2BEGb[1] ,
    \Tile_X4Y8_E2BEGb[0] }),
    .E2MID({\Tile_X4Y8_E2BEG[7] ,
    \Tile_X4Y8_E2BEG[6] ,
    \Tile_X4Y8_E2BEG[5] ,
    \Tile_X4Y8_E2BEG[4] ,
    \Tile_X4Y8_E2BEG[3] ,
    \Tile_X4Y8_E2BEG[2] ,
    \Tile_X4Y8_E2BEG[1] ,
    \Tile_X4Y8_E2BEG[0] }),
    .E6BEG({\Tile_X5Y8_E6BEG[11] ,
    \Tile_X5Y8_E6BEG[10] ,
    \Tile_X5Y8_E6BEG[9] ,
    \Tile_X5Y8_E6BEG[8] ,
    \Tile_X5Y8_E6BEG[7] ,
    \Tile_X5Y8_E6BEG[6] ,
    \Tile_X5Y8_E6BEG[5] ,
    \Tile_X5Y8_E6BEG[4] ,
    \Tile_X5Y8_E6BEG[3] ,
    \Tile_X5Y8_E6BEG[2] ,
    \Tile_X5Y8_E6BEG[1] ,
    \Tile_X5Y8_E6BEG[0] }),
    .E6END({\Tile_X4Y8_E6BEG[11] ,
    \Tile_X4Y8_E6BEG[10] ,
    \Tile_X4Y8_E6BEG[9] ,
    \Tile_X4Y8_E6BEG[8] ,
    \Tile_X4Y8_E6BEG[7] ,
    \Tile_X4Y8_E6BEG[6] ,
    \Tile_X4Y8_E6BEG[5] ,
    \Tile_X4Y8_E6BEG[4] ,
    \Tile_X4Y8_E6BEG[3] ,
    \Tile_X4Y8_E6BEG[2] ,
    \Tile_X4Y8_E6BEG[1] ,
    \Tile_X4Y8_E6BEG[0] }),
    .EE4BEG({\Tile_X5Y8_EE4BEG[15] ,
    \Tile_X5Y8_EE4BEG[14] ,
    \Tile_X5Y8_EE4BEG[13] ,
    \Tile_X5Y8_EE4BEG[12] ,
    \Tile_X5Y8_EE4BEG[11] ,
    \Tile_X5Y8_EE4BEG[10] ,
    \Tile_X5Y8_EE4BEG[9] ,
    \Tile_X5Y8_EE4BEG[8] ,
    \Tile_X5Y8_EE4BEG[7] ,
    \Tile_X5Y8_EE4BEG[6] ,
    \Tile_X5Y8_EE4BEG[5] ,
    \Tile_X5Y8_EE4BEG[4] ,
    \Tile_X5Y8_EE4BEG[3] ,
    \Tile_X5Y8_EE4BEG[2] ,
    \Tile_X5Y8_EE4BEG[1] ,
    \Tile_X5Y8_EE4BEG[0] }),
    .EE4END({\Tile_X4Y8_EE4BEG[15] ,
    \Tile_X4Y8_EE4BEG[14] ,
    \Tile_X4Y8_EE4BEG[13] ,
    \Tile_X4Y8_EE4BEG[12] ,
    \Tile_X4Y8_EE4BEG[11] ,
    \Tile_X4Y8_EE4BEG[10] ,
    \Tile_X4Y8_EE4BEG[9] ,
    \Tile_X4Y8_EE4BEG[8] ,
    \Tile_X4Y8_EE4BEG[7] ,
    \Tile_X4Y8_EE4BEG[6] ,
    \Tile_X4Y8_EE4BEG[5] ,
    \Tile_X4Y8_EE4BEG[4] ,
    \Tile_X4Y8_EE4BEG[3] ,
    \Tile_X4Y8_EE4BEG[2] ,
    \Tile_X4Y8_EE4BEG[1] ,
    \Tile_X4Y8_EE4BEG[0] }),
    .FrameData({\Tile_X4Y8_FrameData_O[31] ,
    \Tile_X4Y8_FrameData_O[30] ,
    \Tile_X4Y8_FrameData_O[29] ,
    \Tile_X4Y8_FrameData_O[28] ,
    \Tile_X4Y8_FrameData_O[27] ,
    \Tile_X4Y8_FrameData_O[26] ,
    \Tile_X4Y8_FrameData_O[25] ,
    \Tile_X4Y8_FrameData_O[24] ,
    \Tile_X4Y8_FrameData_O[23] ,
    \Tile_X4Y8_FrameData_O[22] ,
    \Tile_X4Y8_FrameData_O[21] ,
    \Tile_X4Y8_FrameData_O[20] ,
    \Tile_X4Y8_FrameData_O[19] ,
    \Tile_X4Y8_FrameData_O[18] ,
    \Tile_X4Y8_FrameData_O[17] ,
    \Tile_X4Y8_FrameData_O[16] ,
    \Tile_X4Y8_FrameData_O[15] ,
    \Tile_X4Y8_FrameData_O[14] ,
    \Tile_X4Y8_FrameData_O[13] ,
    \Tile_X4Y8_FrameData_O[12] ,
    \Tile_X4Y8_FrameData_O[11] ,
    \Tile_X4Y8_FrameData_O[10] ,
    \Tile_X4Y8_FrameData_O[9] ,
    \Tile_X4Y8_FrameData_O[8] ,
    \Tile_X4Y8_FrameData_O[7] ,
    \Tile_X4Y8_FrameData_O[6] ,
    \Tile_X4Y8_FrameData_O[5] ,
    \Tile_X4Y8_FrameData_O[4] ,
    \Tile_X4Y8_FrameData_O[3] ,
    \Tile_X4Y8_FrameData_O[2] ,
    \Tile_X4Y8_FrameData_O[1] ,
    \Tile_X4Y8_FrameData_O[0] }),
    .FrameData_O({\Tile_X5Y8_FrameData_O[31] ,
    \Tile_X5Y8_FrameData_O[30] ,
    \Tile_X5Y8_FrameData_O[29] ,
    \Tile_X5Y8_FrameData_O[28] ,
    \Tile_X5Y8_FrameData_O[27] ,
    \Tile_X5Y8_FrameData_O[26] ,
    \Tile_X5Y8_FrameData_O[25] ,
    \Tile_X5Y8_FrameData_O[24] ,
    \Tile_X5Y8_FrameData_O[23] ,
    \Tile_X5Y8_FrameData_O[22] ,
    \Tile_X5Y8_FrameData_O[21] ,
    \Tile_X5Y8_FrameData_O[20] ,
    \Tile_X5Y8_FrameData_O[19] ,
    \Tile_X5Y8_FrameData_O[18] ,
    \Tile_X5Y8_FrameData_O[17] ,
    \Tile_X5Y8_FrameData_O[16] ,
    \Tile_X5Y8_FrameData_O[15] ,
    \Tile_X5Y8_FrameData_O[14] ,
    \Tile_X5Y8_FrameData_O[13] ,
    \Tile_X5Y8_FrameData_O[12] ,
    \Tile_X5Y8_FrameData_O[11] ,
    \Tile_X5Y8_FrameData_O[10] ,
    \Tile_X5Y8_FrameData_O[9] ,
    \Tile_X5Y8_FrameData_O[8] ,
    \Tile_X5Y8_FrameData_O[7] ,
    \Tile_X5Y8_FrameData_O[6] ,
    \Tile_X5Y8_FrameData_O[5] ,
    \Tile_X5Y8_FrameData_O[4] ,
    \Tile_X5Y8_FrameData_O[3] ,
    \Tile_X5Y8_FrameData_O[2] ,
    \Tile_X5Y8_FrameData_O[1] ,
    \Tile_X5Y8_FrameData_O[0] }),
    .FrameStrobe({\Tile_X5Y9_FrameStrobe_O[19] ,
    \Tile_X5Y9_FrameStrobe_O[18] ,
    \Tile_X5Y9_FrameStrobe_O[17] ,
    \Tile_X5Y9_FrameStrobe_O[16] ,
    \Tile_X5Y9_FrameStrobe_O[15] ,
    \Tile_X5Y9_FrameStrobe_O[14] ,
    \Tile_X5Y9_FrameStrobe_O[13] ,
    \Tile_X5Y9_FrameStrobe_O[12] ,
    \Tile_X5Y9_FrameStrobe_O[11] ,
    \Tile_X5Y9_FrameStrobe_O[10] ,
    \Tile_X5Y9_FrameStrobe_O[9] ,
    \Tile_X5Y9_FrameStrobe_O[8] ,
    \Tile_X5Y9_FrameStrobe_O[7] ,
    \Tile_X5Y9_FrameStrobe_O[6] ,
    \Tile_X5Y9_FrameStrobe_O[5] ,
    \Tile_X5Y9_FrameStrobe_O[4] ,
    \Tile_X5Y9_FrameStrobe_O[3] ,
    \Tile_X5Y9_FrameStrobe_O[2] ,
    \Tile_X5Y9_FrameStrobe_O[1] ,
    \Tile_X5Y9_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X5Y8_FrameStrobe_O[19] ,
    \Tile_X5Y8_FrameStrobe_O[18] ,
    \Tile_X5Y8_FrameStrobe_O[17] ,
    \Tile_X5Y8_FrameStrobe_O[16] ,
    \Tile_X5Y8_FrameStrobe_O[15] ,
    \Tile_X5Y8_FrameStrobe_O[14] ,
    \Tile_X5Y8_FrameStrobe_O[13] ,
    \Tile_X5Y8_FrameStrobe_O[12] ,
    \Tile_X5Y8_FrameStrobe_O[11] ,
    \Tile_X5Y8_FrameStrobe_O[10] ,
    \Tile_X5Y8_FrameStrobe_O[9] ,
    \Tile_X5Y8_FrameStrobe_O[8] ,
    \Tile_X5Y8_FrameStrobe_O[7] ,
    \Tile_X5Y8_FrameStrobe_O[6] ,
    \Tile_X5Y8_FrameStrobe_O[5] ,
    \Tile_X5Y8_FrameStrobe_O[4] ,
    \Tile_X5Y8_FrameStrobe_O[3] ,
    \Tile_X5Y8_FrameStrobe_O[2] ,
    \Tile_X5Y8_FrameStrobe_O[1] ,
    \Tile_X5Y8_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X5Y8_N1BEG[3] ,
    \Tile_X5Y8_N1BEG[2] ,
    \Tile_X5Y8_N1BEG[1] ,
    \Tile_X5Y8_N1BEG[0] }),
    .N1END({\Tile_X5Y9_N1BEG[3] ,
    \Tile_X5Y9_N1BEG[2] ,
    \Tile_X5Y9_N1BEG[1] ,
    \Tile_X5Y9_N1BEG[0] }),
    .N2BEG({\Tile_X5Y8_N2BEG[7] ,
    \Tile_X5Y8_N2BEG[6] ,
    \Tile_X5Y8_N2BEG[5] ,
    \Tile_X5Y8_N2BEG[4] ,
    \Tile_X5Y8_N2BEG[3] ,
    \Tile_X5Y8_N2BEG[2] ,
    \Tile_X5Y8_N2BEG[1] ,
    \Tile_X5Y8_N2BEG[0] }),
    .N2BEGb({\Tile_X5Y8_N2BEGb[7] ,
    \Tile_X5Y8_N2BEGb[6] ,
    \Tile_X5Y8_N2BEGb[5] ,
    \Tile_X5Y8_N2BEGb[4] ,
    \Tile_X5Y8_N2BEGb[3] ,
    \Tile_X5Y8_N2BEGb[2] ,
    \Tile_X5Y8_N2BEGb[1] ,
    \Tile_X5Y8_N2BEGb[0] }),
    .N2END({\Tile_X5Y9_N2BEGb[7] ,
    \Tile_X5Y9_N2BEGb[6] ,
    \Tile_X5Y9_N2BEGb[5] ,
    \Tile_X5Y9_N2BEGb[4] ,
    \Tile_X5Y9_N2BEGb[3] ,
    \Tile_X5Y9_N2BEGb[2] ,
    \Tile_X5Y9_N2BEGb[1] ,
    \Tile_X5Y9_N2BEGb[0] }),
    .N2MID({\Tile_X5Y9_N2BEG[7] ,
    \Tile_X5Y9_N2BEG[6] ,
    \Tile_X5Y9_N2BEG[5] ,
    \Tile_X5Y9_N2BEG[4] ,
    \Tile_X5Y9_N2BEG[3] ,
    \Tile_X5Y9_N2BEG[2] ,
    \Tile_X5Y9_N2BEG[1] ,
    \Tile_X5Y9_N2BEG[0] }),
    .N4BEG({\Tile_X5Y8_N4BEG[15] ,
    \Tile_X5Y8_N4BEG[14] ,
    \Tile_X5Y8_N4BEG[13] ,
    \Tile_X5Y8_N4BEG[12] ,
    \Tile_X5Y8_N4BEG[11] ,
    \Tile_X5Y8_N4BEG[10] ,
    \Tile_X5Y8_N4BEG[9] ,
    \Tile_X5Y8_N4BEG[8] ,
    \Tile_X5Y8_N4BEG[7] ,
    \Tile_X5Y8_N4BEG[6] ,
    \Tile_X5Y8_N4BEG[5] ,
    \Tile_X5Y8_N4BEG[4] ,
    \Tile_X5Y8_N4BEG[3] ,
    \Tile_X5Y8_N4BEG[2] ,
    \Tile_X5Y8_N4BEG[1] ,
    \Tile_X5Y8_N4BEG[0] }),
    .N4END({\Tile_X5Y9_N4BEG[15] ,
    \Tile_X5Y9_N4BEG[14] ,
    \Tile_X5Y9_N4BEG[13] ,
    \Tile_X5Y9_N4BEG[12] ,
    \Tile_X5Y9_N4BEG[11] ,
    \Tile_X5Y9_N4BEG[10] ,
    \Tile_X5Y9_N4BEG[9] ,
    \Tile_X5Y9_N4BEG[8] ,
    \Tile_X5Y9_N4BEG[7] ,
    \Tile_X5Y9_N4BEG[6] ,
    \Tile_X5Y9_N4BEG[5] ,
    \Tile_X5Y9_N4BEG[4] ,
    \Tile_X5Y9_N4BEG[3] ,
    \Tile_X5Y9_N4BEG[2] ,
    \Tile_X5Y9_N4BEG[1] ,
    \Tile_X5Y9_N4BEG[0] }),
    .NN4BEG({\Tile_X5Y8_NN4BEG[15] ,
    \Tile_X5Y8_NN4BEG[14] ,
    \Tile_X5Y8_NN4BEG[13] ,
    \Tile_X5Y8_NN4BEG[12] ,
    \Tile_X5Y8_NN4BEG[11] ,
    \Tile_X5Y8_NN4BEG[10] ,
    \Tile_X5Y8_NN4BEG[9] ,
    \Tile_X5Y8_NN4BEG[8] ,
    \Tile_X5Y8_NN4BEG[7] ,
    \Tile_X5Y8_NN4BEG[6] ,
    \Tile_X5Y8_NN4BEG[5] ,
    \Tile_X5Y8_NN4BEG[4] ,
    \Tile_X5Y8_NN4BEG[3] ,
    \Tile_X5Y8_NN4BEG[2] ,
    \Tile_X5Y8_NN4BEG[1] ,
    \Tile_X5Y8_NN4BEG[0] }),
    .NN4END({\Tile_X5Y9_NN4BEG[15] ,
    \Tile_X5Y9_NN4BEG[14] ,
    \Tile_X5Y9_NN4BEG[13] ,
    \Tile_X5Y9_NN4BEG[12] ,
    \Tile_X5Y9_NN4BEG[11] ,
    \Tile_X5Y9_NN4BEG[10] ,
    \Tile_X5Y9_NN4BEG[9] ,
    \Tile_X5Y9_NN4BEG[8] ,
    \Tile_X5Y9_NN4BEG[7] ,
    \Tile_X5Y9_NN4BEG[6] ,
    \Tile_X5Y9_NN4BEG[5] ,
    \Tile_X5Y9_NN4BEG[4] ,
    \Tile_X5Y9_NN4BEG[3] ,
    \Tile_X5Y9_NN4BEG[2] ,
    \Tile_X5Y9_NN4BEG[1] ,
    \Tile_X5Y9_NN4BEG[0] }),
    .S1BEG({\Tile_X5Y8_S1BEG[3] ,
    \Tile_X5Y8_S1BEG[2] ,
    \Tile_X5Y8_S1BEG[1] ,
    \Tile_X5Y8_S1BEG[0] }),
    .S1END({\Tile_X5Y7_S1BEG[3] ,
    \Tile_X5Y7_S1BEG[2] ,
    \Tile_X5Y7_S1BEG[1] ,
    \Tile_X5Y7_S1BEG[0] }),
    .S2BEG({\Tile_X5Y8_S2BEG[7] ,
    \Tile_X5Y8_S2BEG[6] ,
    \Tile_X5Y8_S2BEG[5] ,
    \Tile_X5Y8_S2BEG[4] ,
    \Tile_X5Y8_S2BEG[3] ,
    \Tile_X5Y8_S2BEG[2] ,
    \Tile_X5Y8_S2BEG[1] ,
    \Tile_X5Y8_S2BEG[0] }),
    .S2BEGb({\Tile_X5Y8_S2BEGb[7] ,
    \Tile_X5Y8_S2BEGb[6] ,
    \Tile_X5Y8_S2BEGb[5] ,
    \Tile_X5Y8_S2BEGb[4] ,
    \Tile_X5Y8_S2BEGb[3] ,
    \Tile_X5Y8_S2BEGb[2] ,
    \Tile_X5Y8_S2BEGb[1] ,
    \Tile_X5Y8_S2BEGb[0] }),
    .S2END({\Tile_X5Y7_S2BEGb[7] ,
    \Tile_X5Y7_S2BEGb[6] ,
    \Tile_X5Y7_S2BEGb[5] ,
    \Tile_X5Y7_S2BEGb[4] ,
    \Tile_X5Y7_S2BEGb[3] ,
    \Tile_X5Y7_S2BEGb[2] ,
    \Tile_X5Y7_S2BEGb[1] ,
    \Tile_X5Y7_S2BEGb[0] }),
    .S2MID({\Tile_X5Y7_S2BEG[7] ,
    \Tile_X5Y7_S2BEG[6] ,
    \Tile_X5Y7_S2BEG[5] ,
    \Tile_X5Y7_S2BEG[4] ,
    \Tile_X5Y7_S2BEG[3] ,
    \Tile_X5Y7_S2BEG[2] ,
    \Tile_X5Y7_S2BEG[1] ,
    \Tile_X5Y7_S2BEG[0] }),
    .S4BEG({\Tile_X5Y8_S4BEG[15] ,
    \Tile_X5Y8_S4BEG[14] ,
    \Tile_X5Y8_S4BEG[13] ,
    \Tile_X5Y8_S4BEG[12] ,
    \Tile_X5Y8_S4BEG[11] ,
    \Tile_X5Y8_S4BEG[10] ,
    \Tile_X5Y8_S4BEG[9] ,
    \Tile_X5Y8_S4BEG[8] ,
    \Tile_X5Y8_S4BEG[7] ,
    \Tile_X5Y8_S4BEG[6] ,
    \Tile_X5Y8_S4BEG[5] ,
    \Tile_X5Y8_S4BEG[4] ,
    \Tile_X5Y8_S4BEG[3] ,
    \Tile_X5Y8_S4BEG[2] ,
    \Tile_X5Y8_S4BEG[1] ,
    \Tile_X5Y8_S4BEG[0] }),
    .S4END({\Tile_X5Y7_S4BEG[15] ,
    \Tile_X5Y7_S4BEG[14] ,
    \Tile_X5Y7_S4BEG[13] ,
    \Tile_X5Y7_S4BEG[12] ,
    \Tile_X5Y7_S4BEG[11] ,
    \Tile_X5Y7_S4BEG[10] ,
    \Tile_X5Y7_S4BEG[9] ,
    \Tile_X5Y7_S4BEG[8] ,
    \Tile_X5Y7_S4BEG[7] ,
    \Tile_X5Y7_S4BEG[6] ,
    \Tile_X5Y7_S4BEG[5] ,
    \Tile_X5Y7_S4BEG[4] ,
    \Tile_X5Y7_S4BEG[3] ,
    \Tile_X5Y7_S4BEG[2] ,
    \Tile_X5Y7_S4BEG[1] ,
    \Tile_X5Y7_S4BEG[0] }),
    .SS4BEG({\Tile_X5Y8_SS4BEG[15] ,
    \Tile_X5Y8_SS4BEG[14] ,
    \Tile_X5Y8_SS4BEG[13] ,
    \Tile_X5Y8_SS4BEG[12] ,
    \Tile_X5Y8_SS4BEG[11] ,
    \Tile_X5Y8_SS4BEG[10] ,
    \Tile_X5Y8_SS4BEG[9] ,
    \Tile_X5Y8_SS4BEG[8] ,
    \Tile_X5Y8_SS4BEG[7] ,
    \Tile_X5Y8_SS4BEG[6] ,
    \Tile_X5Y8_SS4BEG[5] ,
    \Tile_X5Y8_SS4BEG[4] ,
    \Tile_X5Y8_SS4BEG[3] ,
    \Tile_X5Y8_SS4BEG[2] ,
    \Tile_X5Y8_SS4BEG[1] ,
    \Tile_X5Y8_SS4BEG[0] }),
    .SS4END({\Tile_X5Y7_SS4BEG[15] ,
    \Tile_X5Y7_SS4BEG[14] ,
    \Tile_X5Y7_SS4BEG[13] ,
    \Tile_X5Y7_SS4BEG[12] ,
    \Tile_X5Y7_SS4BEG[11] ,
    \Tile_X5Y7_SS4BEG[10] ,
    \Tile_X5Y7_SS4BEG[9] ,
    \Tile_X5Y7_SS4BEG[8] ,
    \Tile_X5Y7_SS4BEG[7] ,
    \Tile_X5Y7_SS4BEG[6] ,
    \Tile_X5Y7_SS4BEG[5] ,
    \Tile_X5Y7_SS4BEG[4] ,
    \Tile_X5Y7_SS4BEG[3] ,
    \Tile_X5Y7_SS4BEG[2] ,
    \Tile_X5Y7_SS4BEG[1] ,
    \Tile_X5Y7_SS4BEG[0] }),
    .W1BEG({\Tile_X5Y8_W1BEG[3] ,
    \Tile_X5Y8_W1BEG[2] ,
    \Tile_X5Y8_W1BEG[1] ,
    \Tile_X5Y8_W1BEG[0] }),
    .W1END({\Tile_X6Y8_W1BEG[3] ,
    \Tile_X6Y8_W1BEG[2] ,
    \Tile_X6Y8_W1BEG[1] ,
    \Tile_X6Y8_W1BEG[0] }),
    .W2BEG({\Tile_X5Y8_W2BEG[7] ,
    \Tile_X5Y8_W2BEG[6] ,
    \Tile_X5Y8_W2BEG[5] ,
    \Tile_X5Y8_W2BEG[4] ,
    \Tile_X5Y8_W2BEG[3] ,
    \Tile_X5Y8_W2BEG[2] ,
    \Tile_X5Y8_W2BEG[1] ,
    \Tile_X5Y8_W2BEG[0] }),
    .W2BEGb({\Tile_X5Y8_W2BEGb[7] ,
    \Tile_X5Y8_W2BEGb[6] ,
    \Tile_X5Y8_W2BEGb[5] ,
    \Tile_X5Y8_W2BEGb[4] ,
    \Tile_X5Y8_W2BEGb[3] ,
    \Tile_X5Y8_W2BEGb[2] ,
    \Tile_X5Y8_W2BEGb[1] ,
    \Tile_X5Y8_W2BEGb[0] }),
    .W2END({\Tile_X6Y8_W2BEGb[7] ,
    \Tile_X6Y8_W2BEGb[6] ,
    \Tile_X6Y8_W2BEGb[5] ,
    \Tile_X6Y8_W2BEGb[4] ,
    \Tile_X6Y8_W2BEGb[3] ,
    \Tile_X6Y8_W2BEGb[2] ,
    \Tile_X6Y8_W2BEGb[1] ,
    \Tile_X6Y8_W2BEGb[0] }),
    .W2MID({\Tile_X6Y8_W2BEG[7] ,
    \Tile_X6Y8_W2BEG[6] ,
    \Tile_X6Y8_W2BEG[5] ,
    \Tile_X6Y8_W2BEG[4] ,
    \Tile_X6Y8_W2BEG[3] ,
    \Tile_X6Y8_W2BEG[2] ,
    \Tile_X6Y8_W2BEG[1] ,
    \Tile_X6Y8_W2BEG[0] }),
    .W6BEG({\Tile_X5Y8_W6BEG[11] ,
    \Tile_X5Y8_W6BEG[10] ,
    \Tile_X5Y8_W6BEG[9] ,
    \Tile_X5Y8_W6BEG[8] ,
    \Tile_X5Y8_W6BEG[7] ,
    \Tile_X5Y8_W6BEG[6] ,
    \Tile_X5Y8_W6BEG[5] ,
    \Tile_X5Y8_W6BEG[4] ,
    \Tile_X5Y8_W6BEG[3] ,
    \Tile_X5Y8_W6BEG[2] ,
    \Tile_X5Y8_W6BEG[1] ,
    \Tile_X5Y8_W6BEG[0] }),
    .W6END({\Tile_X6Y8_W6BEG[11] ,
    \Tile_X6Y8_W6BEG[10] ,
    \Tile_X6Y8_W6BEG[9] ,
    \Tile_X6Y8_W6BEG[8] ,
    \Tile_X6Y8_W6BEG[7] ,
    \Tile_X6Y8_W6BEG[6] ,
    \Tile_X6Y8_W6BEG[5] ,
    \Tile_X6Y8_W6BEG[4] ,
    \Tile_X6Y8_W6BEG[3] ,
    \Tile_X6Y8_W6BEG[2] ,
    \Tile_X6Y8_W6BEG[1] ,
    \Tile_X6Y8_W6BEG[0] }),
    .WW4BEG({\Tile_X5Y8_WW4BEG[15] ,
    \Tile_X5Y8_WW4BEG[14] ,
    \Tile_X5Y8_WW4BEG[13] ,
    \Tile_X5Y8_WW4BEG[12] ,
    \Tile_X5Y8_WW4BEG[11] ,
    \Tile_X5Y8_WW4BEG[10] ,
    \Tile_X5Y8_WW4BEG[9] ,
    \Tile_X5Y8_WW4BEG[8] ,
    \Tile_X5Y8_WW4BEG[7] ,
    \Tile_X5Y8_WW4BEG[6] ,
    \Tile_X5Y8_WW4BEG[5] ,
    \Tile_X5Y8_WW4BEG[4] ,
    \Tile_X5Y8_WW4BEG[3] ,
    \Tile_X5Y8_WW4BEG[2] ,
    \Tile_X5Y8_WW4BEG[1] ,
    \Tile_X5Y8_WW4BEG[0] }),
    .WW4END({\Tile_X6Y8_WW4BEG[15] ,
    \Tile_X6Y8_WW4BEG[14] ,
    \Tile_X6Y8_WW4BEG[13] ,
    \Tile_X6Y8_WW4BEG[12] ,
    \Tile_X6Y8_WW4BEG[11] ,
    \Tile_X6Y8_WW4BEG[10] ,
    \Tile_X6Y8_WW4BEG[9] ,
    \Tile_X6Y8_WW4BEG[8] ,
    \Tile_X6Y8_WW4BEG[7] ,
    \Tile_X6Y8_WW4BEG[6] ,
    \Tile_X6Y8_WW4BEG[5] ,
    \Tile_X6Y8_WW4BEG[4] ,
    \Tile_X6Y8_WW4BEG[3] ,
    \Tile_X6Y8_WW4BEG[2] ,
    \Tile_X6Y8_WW4BEG[1] ,
    \Tile_X6Y8_WW4BEG[0] }));
 LUT4AB Tile_X5Y9_LUT4AB (.Ci(Tile_X5Y10_Co),
    .Co(Tile_X5Y9_Co),
    .UserCLK(Tile_X5Y10_UserCLKo),
    .UserCLKo(Tile_X5Y9_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X5Y9_E1BEG[3] ,
    \Tile_X5Y9_E1BEG[2] ,
    \Tile_X5Y9_E1BEG[1] ,
    \Tile_X5Y9_E1BEG[0] }),
    .E1END({\Tile_X4Y9_E1BEG[3] ,
    \Tile_X4Y9_E1BEG[2] ,
    \Tile_X4Y9_E1BEG[1] ,
    \Tile_X4Y9_E1BEG[0] }),
    .E2BEG({\Tile_X5Y9_E2BEG[7] ,
    \Tile_X5Y9_E2BEG[6] ,
    \Tile_X5Y9_E2BEG[5] ,
    \Tile_X5Y9_E2BEG[4] ,
    \Tile_X5Y9_E2BEG[3] ,
    \Tile_X5Y9_E2BEG[2] ,
    \Tile_X5Y9_E2BEG[1] ,
    \Tile_X5Y9_E2BEG[0] }),
    .E2BEGb({\Tile_X5Y9_E2BEGb[7] ,
    \Tile_X5Y9_E2BEGb[6] ,
    \Tile_X5Y9_E2BEGb[5] ,
    \Tile_X5Y9_E2BEGb[4] ,
    \Tile_X5Y9_E2BEGb[3] ,
    \Tile_X5Y9_E2BEGb[2] ,
    \Tile_X5Y9_E2BEGb[1] ,
    \Tile_X5Y9_E2BEGb[0] }),
    .E2END({\Tile_X4Y9_E2BEGb[7] ,
    \Tile_X4Y9_E2BEGb[6] ,
    \Tile_X4Y9_E2BEGb[5] ,
    \Tile_X4Y9_E2BEGb[4] ,
    \Tile_X4Y9_E2BEGb[3] ,
    \Tile_X4Y9_E2BEGb[2] ,
    \Tile_X4Y9_E2BEGb[1] ,
    \Tile_X4Y9_E2BEGb[0] }),
    .E2MID({\Tile_X4Y9_E2BEG[7] ,
    \Tile_X4Y9_E2BEG[6] ,
    \Tile_X4Y9_E2BEG[5] ,
    \Tile_X4Y9_E2BEG[4] ,
    \Tile_X4Y9_E2BEG[3] ,
    \Tile_X4Y9_E2BEG[2] ,
    \Tile_X4Y9_E2BEG[1] ,
    \Tile_X4Y9_E2BEG[0] }),
    .E6BEG({\Tile_X5Y9_E6BEG[11] ,
    \Tile_X5Y9_E6BEG[10] ,
    \Tile_X5Y9_E6BEG[9] ,
    \Tile_X5Y9_E6BEG[8] ,
    \Tile_X5Y9_E6BEG[7] ,
    \Tile_X5Y9_E6BEG[6] ,
    \Tile_X5Y9_E6BEG[5] ,
    \Tile_X5Y9_E6BEG[4] ,
    \Tile_X5Y9_E6BEG[3] ,
    \Tile_X5Y9_E6BEG[2] ,
    \Tile_X5Y9_E6BEG[1] ,
    \Tile_X5Y9_E6BEG[0] }),
    .E6END({\Tile_X4Y9_E6BEG[11] ,
    \Tile_X4Y9_E6BEG[10] ,
    \Tile_X4Y9_E6BEG[9] ,
    \Tile_X4Y9_E6BEG[8] ,
    \Tile_X4Y9_E6BEG[7] ,
    \Tile_X4Y9_E6BEG[6] ,
    \Tile_X4Y9_E6BEG[5] ,
    \Tile_X4Y9_E6BEG[4] ,
    \Tile_X4Y9_E6BEG[3] ,
    \Tile_X4Y9_E6BEG[2] ,
    \Tile_X4Y9_E6BEG[1] ,
    \Tile_X4Y9_E6BEG[0] }),
    .EE4BEG({\Tile_X5Y9_EE4BEG[15] ,
    \Tile_X5Y9_EE4BEG[14] ,
    \Tile_X5Y9_EE4BEG[13] ,
    \Tile_X5Y9_EE4BEG[12] ,
    \Tile_X5Y9_EE4BEG[11] ,
    \Tile_X5Y9_EE4BEG[10] ,
    \Tile_X5Y9_EE4BEG[9] ,
    \Tile_X5Y9_EE4BEG[8] ,
    \Tile_X5Y9_EE4BEG[7] ,
    \Tile_X5Y9_EE4BEG[6] ,
    \Tile_X5Y9_EE4BEG[5] ,
    \Tile_X5Y9_EE4BEG[4] ,
    \Tile_X5Y9_EE4BEG[3] ,
    \Tile_X5Y9_EE4BEG[2] ,
    \Tile_X5Y9_EE4BEG[1] ,
    \Tile_X5Y9_EE4BEG[0] }),
    .EE4END({\Tile_X4Y9_EE4BEG[15] ,
    \Tile_X4Y9_EE4BEG[14] ,
    \Tile_X4Y9_EE4BEG[13] ,
    \Tile_X4Y9_EE4BEG[12] ,
    \Tile_X4Y9_EE4BEG[11] ,
    \Tile_X4Y9_EE4BEG[10] ,
    \Tile_X4Y9_EE4BEG[9] ,
    \Tile_X4Y9_EE4BEG[8] ,
    \Tile_X4Y9_EE4BEG[7] ,
    \Tile_X4Y9_EE4BEG[6] ,
    \Tile_X4Y9_EE4BEG[5] ,
    \Tile_X4Y9_EE4BEG[4] ,
    \Tile_X4Y9_EE4BEG[3] ,
    \Tile_X4Y9_EE4BEG[2] ,
    \Tile_X4Y9_EE4BEG[1] ,
    \Tile_X4Y9_EE4BEG[0] }),
    .FrameData({\Tile_X4Y9_FrameData_O[31] ,
    \Tile_X4Y9_FrameData_O[30] ,
    \Tile_X4Y9_FrameData_O[29] ,
    \Tile_X4Y9_FrameData_O[28] ,
    \Tile_X4Y9_FrameData_O[27] ,
    \Tile_X4Y9_FrameData_O[26] ,
    \Tile_X4Y9_FrameData_O[25] ,
    \Tile_X4Y9_FrameData_O[24] ,
    \Tile_X4Y9_FrameData_O[23] ,
    \Tile_X4Y9_FrameData_O[22] ,
    \Tile_X4Y9_FrameData_O[21] ,
    \Tile_X4Y9_FrameData_O[20] ,
    \Tile_X4Y9_FrameData_O[19] ,
    \Tile_X4Y9_FrameData_O[18] ,
    \Tile_X4Y9_FrameData_O[17] ,
    \Tile_X4Y9_FrameData_O[16] ,
    \Tile_X4Y9_FrameData_O[15] ,
    \Tile_X4Y9_FrameData_O[14] ,
    \Tile_X4Y9_FrameData_O[13] ,
    \Tile_X4Y9_FrameData_O[12] ,
    \Tile_X4Y9_FrameData_O[11] ,
    \Tile_X4Y9_FrameData_O[10] ,
    \Tile_X4Y9_FrameData_O[9] ,
    \Tile_X4Y9_FrameData_O[8] ,
    \Tile_X4Y9_FrameData_O[7] ,
    \Tile_X4Y9_FrameData_O[6] ,
    \Tile_X4Y9_FrameData_O[5] ,
    \Tile_X4Y9_FrameData_O[4] ,
    \Tile_X4Y9_FrameData_O[3] ,
    \Tile_X4Y9_FrameData_O[2] ,
    \Tile_X4Y9_FrameData_O[1] ,
    \Tile_X4Y9_FrameData_O[0] }),
    .FrameData_O({\Tile_X5Y9_FrameData_O[31] ,
    \Tile_X5Y9_FrameData_O[30] ,
    \Tile_X5Y9_FrameData_O[29] ,
    \Tile_X5Y9_FrameData_O[28] ,
    \Tile_X5Y9_FrameData_O[27] ,
    \Tile_X5Y9_FrameData_O[26] ,
    \Tile_X5Y9_FrameData_O[25] ,
    \Tile_X5Y9_FrameData_O[24] ,
    \Tile_X5Y9_FrameData_O[23] ,
    \Tile_X5Y9_FrameData_O[22] ,
    \Tile_X5Y9_FrameData_O[21] ,
    \Tile_X5Y9_FrameData_O[20] ,
    \Tile_X5Y9_FrameData_O[19] ,
    \Tile_X5Y9_FrameData_O[18] ,
    \Tile_X5Y9_FrameData_O[17] ,
    \Tile_X5Y9_FrameData_O[16] ,
    \Tile_X5Y9_FrameData_O[15] ,
    \Tile_X5Y9_FrameData_O[14] ,
    \Tile_X5Y9_FrameData_O[13] ,
    \Tile_X5Y9_FrameData_O[12] ,
    \Tile_X5Y9_FrameData_O[11] ,
    \Tile_X5Y9_FrameData_O[10] ,
    \Tile_X5Y9_FrameData_O[9] ,
    \Tile_X5Y9_FrameData_O[8] ,
    \Tile_X5Y9_FrameData_O[7] ,
    \Tile_X5Y9_FrameData_O[6] ,
    \Tile_X5Y9_FrameData_O[5] ,
    \Tile_X5Y9_FrameData_O[4] ,
    \Tile_X5Y9_FrameData_O[3] ,
    \Tile_X5Y9_FrameData_O[2] ,
    \Tile_X5Y9_FrameData_O[1] ,
    \Tile_X5Y9_FrameData_O[0] }),
    .FrameStrobe({\Tile_X5Y10_FrameStrobe_O[19] ,
    \Tile_X5Y10_FrameStrobe_O[18] ,
    \Tile_X5Y10_FrameStrobe_O[17] ,
    \Tile_X5Y10_FrameStrobe_O[16] ,
    \Tile_X5Y10_FrameStrobe_O[15] ,
    \Tile_X5Y10_FrameStrobe_O[14] ,
    \Tile_X5Y10_FrameStrobe_O[13] ,
    \Tile_X5Y10_FrameStrobe_O[12] ,
    \Tile_X5Y10_FrameStrobe_O[11] ,
    \Tile_X5Y10_FrameStrobe_O[10] ,
    \Tile_X5Y10_FrameStrobe_O[9] ,
    \Tile_X5Y10_FrameStrobe_O[8] ,
    \Tile_X5Y10_FrameStrobe_O[7] ,
    \Tile_X5Y10_FrameStrobe_O[6] ,
    \Tile_X5Y10_FrameStrobe_O[5] ,
    \Tile_X5Y10_FrameStrobe_O[4] ,
    \Tile_X5Y10_FrameStrobe_O[3] ,
    \Tile_X5Y10_FrameStrobe_O[2] ,
    \Tile_X5Y10_FrameStrobe_O[1] ,
    \Tile_X5Y10_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X5Y9_FrameStrobe_O[19] ,
    \Tile_X5Y9_FrameStrobe_O[18] ,
    \Tile_X5Y9_FrameStrobe_O[17] ,
    \Tile_X5Y9_FrameStrobe_O[16] ,
    \Tile_X5Y9_FrameStrobe_O[15] ,
    \Tile_X5Y9_FrameStrobe_O[14] ,
    \Tile_X5Y9_FrameStrobe_O[13] ,
    \Tile_X5Y9_FrameStrobe_O[12] ,
    \Tile_X5Y9_FrameStrobe_O[11] ,
    \Tile_X5Y9_FrameStrobe_O[10] ,
    \Tile_X5Y9_FrameStrobe_O[9] ,
    \Tile_X5Y9_FrameStrobe_O[8] ,
    \Tile_X5Y9_FrameStrobe_O[7] ,
    \Tile_X5Y9_FrameStrobe_O[6] ,
    \Tile_X5Y9_FrameStrobe_O[5] ,
    \Tile_X5Y9_FrameStrobe_O[4] ,
    \Tile_X5Y9_FrameStrobe_O[3] ,
    \Tile_X5Y9_FrameStrobe_O[2] ,
    \Tile_X5Y9_FrameStrobe_O[1] ,
    \Tile_X5Y9_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X5Y9_N1BEG[3] ,
    \Tile_X5Y9_N1BEG[2] ,
    \Tile_X5Y9_N1BEG[1] ,
    \Tile_X5Y9_N1BEG[0] }),
    .N1END({\Tile_X5Y10_N1BEG[3] ,
    \Tile_X5Y10_N1BEG[2] ,
    \Tile_X5Y10_N1BEG[1] ,
    \Tile_X5Y10_N1BEG[0] }),
    .N2BEG({\Tile_X5Y9_N2BEG[7] ,
    \Tile_X5Y9_N2BEG[6] ,
    \Tile_X5Y9_N2BEG[5] ,
    \Tile_X5Y9_N2BEG[4] ,
    \Tile_X5Y9_N2BEG[3] ,
    \Tile_X5Y9_N2BEG[2] ,
    \Tile_X5Y9_N2BEG[1] ,
    \Tile_X5Y9_N2BEG[0] }),
    .N2BEGb({\Tile_X5Y9_N2BEGb[7] ,
    \Tile_X5Y9_N2BEGb[6] ,
    \Tile_X5Y9_N2BEGb[5] ,
    \Tile_X5Y9_N2BEGb[4] ,
    \Tile_X5Y9_N2BEGb[3] ,
    \Tile_X5Y9_N2BEGb[2] ,
    \Tile_X5Y9_N2BEGb[1] ,
    \Tile_X5Y9_N2BEGb[0] }),
    .N2END({\Tile_X5Y10_N2BEGb[7] ,
    \Tile_X5Y10_N2BEGb[6] ,
    \Tile_X5Y10_N2BEGb[5] ,
    \Tile_X5Y10_N2BEGb[4] ,
    \Tile_X5Y10_N2BEGb[3] ,
    \Tile_X5Y10_N2BEGb[2] ,
    \Tile_X5Y10_N2BEGb[1] ,
    \Tile_X5Y10_N2BEGb[0] }),
    .N2MID({\Tile_X5Y10_N2BEG[7] ,
    \Tile_X5Y10_N2BEG[6] ,
    \Tile_X5Y10_N2BEG[5] ,
    \Tile_X5Y10_N2BEG[4] ,
    \Tile_X5Y10_N2BEG[3] ,
    \Tile_X5Y10_N2BEG[2] ,
    \Tile_X5Y10_N2BEG[1] ,
    \Tile_X5Y10_N2BEG[0] }),
    .N4BEG({\Tile_X5Y9_N4BEG[15] ,
    \Tile_X5Y9_N4BEG[14] ,
    \Tile_X5Y9_N4BEG[13] ,
    \Tile_X5Y9_N4BEG[12] ,
    \Tile_X5Y9_N4BEG[11] ,
    \Tile_X5Y9_N4BEG[10] ,
    \Tile_X5Y9_N4BEG[9] ,
    \Tile_X5Y9_N4BEG[8] ,
    \Tile_X5Y9_N4BEG[7] ,
    \Tile_X5Y9_N4BEG[6] ,
    \Tile_X5Y9_N4BEG[5] ,
    \Tile_X5Y9_N4BEG[4] ,
    \Tile_X5Y9_N4BEG[3] ,
    \Tile_X5Y9_N4BEG[2] ,
    \Tile_X5Y9_N4BEG[1] ,
    \Tile_X5Y9_N4BEG[0] }),
    .N4END({\Tile_X5Y10_N4BEG[15] ,
    \Tile_X5Y10_N4BEG[14] ,
    \Tile_X5Y10_N4BEG[13] ,
    \Tile_X5Y10_N4BEG[12] ,
    \Tile_X5Y10_N4BEG[11] ,
    \Tile_X5Y10_N4BEG[10] ,
    \Tile_X5Y10_N4BEG[9] ,
    \Tile_X5Y10_N4BEG[8] ,
    \Tile_X5Y10_N4BEG[7] ,
    \Tile_X5Y10_N4BEG[6] ,
    \Tile_X5Y10_N4BEG[5] ,
    \Tile_X5Y10_N4BEG[4] ,
    \Tile_X5Y10_N4BEG[3] ,
    \Tile_X5Y10_N4BEG[2] ,
    \Tile_X5Y10_N4BEG[1] ,
    \Tile_X5Y10_N4BEG[0] }),
    .NN4BEG({\Tile_X5Y9_NN4BEG[15] ,
    \Tile_X5Y9_NN4BEG[14] ,
    \Tile_X5Y9_NN4BEG[13] ,
    \Tile_X5Y9_NN4BEG[12] ,
    \Tile_X5Y9_NN4BEG[11] ,
    \Tile_X5Y9_NN4BEG[10] ,
    \Tile_X5Y9_NN4BEG[9] ,
    \Tile_X5Y9_NN4BEG[8] ,
    \Tile_X5Y9_NN4BEG[7] ,
    \Tile_X5Y9_NN4BEG[6] ,
    \Tile_X5Y9_NN4BEG[5] ,
    \Tile_X5Y9_NN4BEG[4] ,
    \Tile_X5Y9_NN4BEG[3] ,
    \Tile_X5Y9_NN4BEG[2] ,
    \Tile_X5Y9_NN4BEG[1] ,
    \Tile_X5Y9_NN4BEG[0] }),
    .NN4END({\Tile_X5Y10_NN4BEG[15] ,
    \Tile_X5Y10_NN4BEG[14] ,
    \Tile_X5Y10_NN4BEG[13] ,
    \Tile_X5Y10_NN4BEG[12] ,
    \Tile_X5Y10_NN4BEG[11] ,
    \Tile_X5Y10_NN4BEG[10] ,
    \Tile_X5Y10_NN4BEG[9] ,
    \Tile_X5Y10_NN4BEG[8] ,
    \Tile_X5Y10_NN4BEG[7] ,
    \Tile_X5Y10_NN4BEG[6] ,
    \Tile_X5Y10_NN4BEG[5] ,
    \Tile_X5Y10_NN4BEG[4] ,
    \Tile_X5Y10_NN4BEG[3] ,
    \Tile_X5Y10_NN4BEG[2] ,
    \Tile_X5Y10_NN4BEG[1] ,
    \Tile_X5Y10_NN4BEG[0] }),
    .S1BEG({\Tile_X5Y9_S1BEG[3] ,
    \Tile_X5Y9_S1BEG[2] ,
    \Tile_X5Y9_S1BEG[1] ,
    \Tile_X5Y9_S1BEG[0] }),
    .S1END({\Tile_X5Y8_S1BEG[3] ,
    \Tile_X5Y8_S1BEG[2] ,
    \Tile_X5Y8_S1BEG[1] ,
    \Tile_X5Y8_S1BEG[0] }),
    .S2BEG({\Tile_X5Y9_S2BEG[7] ,
    \Tile_X5Y9_S2BEG[6] ,
    \Tile_X5Y9_S2BEG[5] ,
    \Tile_X5Y9_S2BEG[4] ,
    \Tile_X5Y9_S2BEG[3] ,
    \Tile_X5Y9_S2BEG[2] ,
    \Tile_X5Y9_S2BEG[1] ,
    \Tile_X5Y9_S2BEG[0] }),
    .S2BEGb({\Tile_X5Y9_S2BEGb[7] ,
    \Tile_X5Y9_S2BEGb[6] ,
    \Tile_X5Y9_S2BEGb[5] ,
    \Tile_X5Y9_S2BEGb[4] ,
    \Tile_X5Y9_S2BEGb[3] ,
    \Tile_X5Y9_S2BEGb[2] ,
    \Tile_X5Y9_S2BEGb[1] ,
    \Tile_X5Y9_S2BEGb[0] }),
    .S2END({\Tile_X5Y8_S2BEGb[7] ,
    \Tile_X5Y8_S2BEGb[6] ,
    \Tile_X5Y8_S2BEGb[5] ,
    \Tile_X5Y8_S2BEGb[4] ,
    \Tile_X5Y8_S2BEGb[3] ,
    \Tile_X5Y8_S2BEGb[2] ,
    \Tile_X5Y8_S2BEGb[1] ,
    \Tile_X5Y8_S2BEGb[0] }),
    .S2MID({\Tile_X5Y8_S2BEG[7] ,
    \Tile_X5Y8_S2BEG[6] ,
    \Tile_X5Y8_S2BEG[5] ,
    \Tile_X5Y8_S2BEG[4] ,
    \Tile_X5Y8_S2BEG[3] ,
    \Tile_X5Y8_S2BEG[2] ,
    \Tile_X5Y8_S2BEG[1] ,
    \Tile_X5Y8_S2BEG[0] }),
    .S4BEG({\Tile_X5Y9_S4BEG[15] ,
    \Tile_X5Y9_S4BEG[14] ,
    \Tile_X5Y9_S4BEG[13] ,
    \Tile_X5Y9_S4BEG[12] ,
    \Tile_X5Y9_S4BEG[11] ,
    \Tile_X5Y9_S4BEG[10] ,
    \Tile_X5Y9_S4BEG[9] ,
    \Tile_X5Y9_S4BEG[8] ,
    \Tile_X5Y9_S4BEG[7] ,
    \Tile_X5Y9_S4BEG[6] ,
    \Tile_X5Y9_S4BEG[5] ,
    \Tile_X5Y9_S4BEG[4] ,
    \Tile_X5Y9_S4BEG[3] ,
    \Tile_X5Y9_S4BEG[2] ,
    \Tile_X5Y9_S4BEG[1] ,
    \Tile_X5Y9_S4BEG[0] }),
    .S4END({\Tile_X5Y8_S4BEG[15] ,
    \Tile_X5Y8_S4BEG[14] ,
    \Tile_X5Y8_S4BEG[13] ,
    \Tile_X5Y8_S4BEG[12] ,
    \Tile_X5Y8_S4BEG[11] ,
    \Tile_X5Y8_S4BEG[10] ,
    \Tile_X5Y8_S4BEG[9] ,
    \Tile_X5Y8_S4BEG[8] ,
    \Tile_X5Y8_S4BEG[7] ,
    \Tile_X5Y8_S4BEG[6] ,
    \Tile_X5Y8_S4BEG[5] ,
    \Tile_X5Y8_S4BEG[4] ,
    \Tile_X5Y8_S4BEG[3] ,
    \Tile_X5Y8_S4BEG[2] ,
    \Tile_X5Y8_S4BEG[1] ,
    \Tile_X5Y8_S4BEG[0] }),
    .SS4BEG({\Tile_X5Y9_SS4BEG[15] ,
    \Tile_X5Y9_SS4BEG[14] ,
    \Tile_X5Y9_SS4BEG[13] ,
    \Tile_X5Y9_SS4BEG[12] ,
    \Tile_X5Y9_SS4BEG[11] ,
    \Tile_X5Y9_SS4BEG[10] ,
    \Tile_X5Y9_SS4BEG[9] ,
    \Tile_X5Y9_SS4BEG[8] ,
    \Tile_X5Y9_SS4BEG[7] ,
    \Tile_X5Y9_SS4BEG[6] ,
    \Tile_X5Y9_SS4BEG[5] ,
    \Tile_X5Y9_SS4BEG[4] ,
    \Tile_X5Y9_SS4BEG[3] ,
    \Tile_X5Y9_SS4BEG[2] ,
    \Tile_X5Y9_SS4BEG[1] ,
    \Tile_X5Y9_SS4BEG[0] }),
    .SS4END({\Tile_X5Y8_SS4BEG[15] ,
    \Tile_X5Y8_SS4BEG[14] ,
    \Tile_X5Y8_SS4BEG[13] ,
    \Tile_X5Y8_SS4BEG[12] ,
    \Tile_X5Y8_SS4BEG[11] ,
    \Tile_X5Y8_SS4BEG[10] ,
    \Tile_X5Y8_SS4BEG[9] ,
    \Tile_X5Y8_SS4BEG[8] ,
    \Tile_X5Y8_SS4BEG[7] ,
    \Tile_X5Y8_SS4BEG[6] ,
    \Tile_X5Y8_SS4BEG[5] ,
    \Tile_X5Y8_SS4BEG[4] ,
    \Tile_X5Y8_SS4BEG[3] ,
    \Tile_X5Y8_SS4BEG[2] ,
    \Tile_X5Y8_SS4BEG[1] ,
    \Tile_X5Y8_SS4BEG[0] }),
    .W1BEG({\Tile_X5Y9_W1BEG[3] ,
    \Tile_X5Y9_W1BEG[2] ,
    \Tile_X5Y9_W1BEG[1] ,
    \Tile_X5Y9_W1BEG[0] }),
    .W1END({\Tile_X6Y9_W1BEG[3] ,
    \Tile_X6Y9_W1BEG[2] ,
    \Tile_X6Y9_W1BEG[1] ,
    \Tile_X6Y9_W1BEG[0] }),
    .W2BEG({\Tile_X5Y9_W2BEG[7] ,
    \Tile_X5Y9_W2BEG[6] ,
    \Tile_X5Y9_W2BEG[5] ,
    \Tile_X5Y9_W2BEG[4] ,
    \Tile_X5Y9_W2BEG[3] ,
    \Tile_X5Y9_W2BEG[2] ,
    \Tile_X5Y9_W2BEG[1] ,
    \Tile_X5Y9_W2BEG[0] }),
    .W2BEGb({\Tile_X5Y9_W2BEGb[7] ,
    \Tile_X5Y9_W2BEGb[6] ,
    \Tile_X5Y9_W2BEGb[5] ,
    \Tile_X5Y9_W2BEGb[4] ,
    \Tile_X5Y9_W2BEGb[3] ,
    \Tile_X5Y9_W2BEGb[2] ,
    \Tile_X5Y9_W2BEGb[1] ,
    \Tile_X5Y9_W2BEGb[0] }),
    .W2END({\Tile_X6Y9_W2BEGb[7] ,
    \Tile_X6Y9_W2BEGb[6] ,
    \Tile_X6Y9_W2BEGb[5] ,
    \Tile_X6Y9_W2BEGb[4] ,
    \Tile_X6Y9_W2BEGb[3] ,
    \Tile_X6Y9_W2BEGb[2] ,
    \Tile_X6Y9_W2BEGb[1] ,
    \Tile_X6Y9_W2BEGb[0] }),
    .W2MID({\Tile_X6Y9_W2BEG[7] ,
    \Tile_X6Y9_W2BEG[6] ,
    \Tile_X6Y9_W2BEG[5] ,
    \Tile_X6Y9_W2BEG[4] ,
    \Tile_X6Y9_W2BEG[3] ,
    \Tile_X6Y9_W2BEG[2] ,
    \Tile_X6Y9_W2BEG[1] ,
    \Tile_X6Y9_W2BEG[0] }),
    .W6BEG({\Tile_X5Y9_W6BEG[11] ,
    \Tile_X5Y9_W6BEG[10] ,
    \Tile_X5Y9_W6BEG[9] ,
    \Tile_X5Y9_W6BEG[8] ,
    \Tile_X5Y9_W6BEG[7] ,
    \Tile_X5Y9_W6BEG[6] ,
    \Tile_X5Y9_W6BEG[5] ,
    \Tile_X5Y9_W6BEG[4] ,
    \Tile_X5Y9_W6BEG[3] ,
    \Tile_X5Y9_W6BEG[2] ,
    \Tile_X5Y9_W6BEG[1] ,
    \Tile_X5Y9_W6BEG[0] }),
    .W6END({\Tile_X6Y9_W6BEG[11] ,
    \Tile_X6Y9_W6BEG[10] ,
    \Tile_X6Y9_W6BEG[9] ,
    \Tile_X6Y9_W6BEG[8] ,
    \Tile_X6Y9_W6BEG[7] ,
    \Tile_X6Y9_W6BEG[6] ,
    \Tile_X6Y9_W6BEG[5] ,
    \Tile_X6Y9_W6BEG[4] ,
    \Tile_X6Y9_W6BEG[3] ,
    \Tile_X6Y9_W6BEG[2] ,
    \Tile_X6Y9_W6BEG[1] ,
    \Tile_X6Y9_W6BEG[0] }),
    .WW4BEG({\Tile_X5Y9_WW4BEG[15] ,
    \Tile_X5Y9_WW4BEG[14] ,
    \Tile_X5Y9_WW4BEG[13] ,
    \Tile_X5Y9_WW4BEG[12] ,
    \Tile_X5Y9_WW4BEG[11] ,
    \Tile_X5Y9_WW4BEG[10] ,
    \Tile_X5Y9_WW4BEG[9] ,
    \Tile_X5Y9_WW4BEG[8] ,
    \Tile_X5Y9_WW4BEG[7] ,
    \Tile_X5Y9_WW4BEG[6] ,
    \Tile_X5Y9_WW4BEG[5] ,
    \Tile_X5Y9_WW4BEG[4] ,
    \Tile_X5Y9_WW4BEG[3] ,
    \Tile_X5Y9_WW4BEG[2] ,
    \Tile_X5Y9_WW4BEG[1] ,
    \Tile_X5Y9_WW4BEG[0] }),
    .WW4END({\Tile_X6Y9_WW4BEG[15] ,
    \Tile_X6Y9_WW4BEG[14] ,
    \Tile_X6Y9_WW4BEG[13] ,
    \Tile_X6Y9_WW4BEG[12] ,
    \Tile_X6Y9_WW4BEG[11] ,
    \Tile_X6Y9_WW4BEG[10] ,
    \Tile_X6Y9_WW4BEG[9] ,
    \Tile_X6Y9_WW4BEG[8] ,
    \Tile_X6Y9_WW4BEG[7] ,
    \Tile_X6Y9_WW4BEG[6] ,
    \Tile_X6Y9_WW4BEG[5] ,
    \Tile_X6Y9_WW4BEG[4] ,
    \Tile_X6Y9_WW4BEG[3] ,
    \Tile_X6Y9_WW4BEG[2] ,
    \Tile_X6Y9_WW4BEG[1] ,
    \Tile_X6Y9_WW4BEG[0] }));
 N_term_single Tile_X6Y0_N_term_single (.Ci(Tile_X6Y1_Co),
    .UserCLK(Tile_X6Y1_UserCLKo),
    .UserCLKo(Tile_X6Y0_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .FrameData({\Tile_X5Y0_FrameData_O[31] ,
    \Tile_X5Y0_FrameData_O[30] ,
    \Tile_X5Y0_FrameData_O[29] ,
    \Tile_X5Y0_FrameData_O[28] ,
    \Tile_X5Y0_FrameData_O[27] ,
    \Tile_X5Y0_FrameData_O[26] ,
    \Tile_X5Y0_FrameData_O[25] ,
    \Tile_X5Y0_FrameData_O[24] ,
    \Tile_X5Y0_FrameData_O[23] ,
    \Tile_X5Y0_FrameData_O[22] ,
    \Tile_X5Y0_FrameData_O[21] ,
    \Tile_X5Y0_FrameData_O[20] ,
    \Tile_X5Y0_FrameData_O[19] ,
    \Tile_X5Y0_FrameData_O[18] ,
    \Tile_X5Y0_FrameData_O[17] ,
    \Tile_X5Y0_FrameData_O[16] ,
    \Tile_X5Y0_FrameData_O[15] ,
    \Tile_X5Y0_FrameData_O[14] ,
    \Tile_X5Y0_FrameData_O[13] ,
    \Tile_X5Y0_FrameData_O[12] ,
    \Tile_X5Y0_FrameData_O[11] ,
    \Tile_X5Y0_FrameData_O[10] ,
    \Tile_X5Y0_FrameData_O[9] ,
    \Tile_X5Y0_FrameData_O[8] ,
    \Tile_X5Y0_FrameData_O[7] ,
    \Tile_X5Y0_FrameData_O[6] ,
    \Tile_X5Y0_FrameData_O[5] ,
    \Tile_X5Y0_FrameData_O[4] ,
    \Tile_X5Y0_FrameData_O[3] ,
    \Tile_X5Y0_FrameData_O[2] ,
    \Tile_X5Y0_FrameData_O[1] ,
    \Tile_X5Y0_FrameData_O[0] }),
    .FrameData_O({\Tile_X6Y0_FrameData_O[31] ,
    \Tile_X6Y0_FrameData_O[30] ,
    \Tile_X6Y0_FrameData_O[29] ,
    \Tile_X6Y0_FrameData_O[28] ,
    \Tile_X6Y0_FrameData_O[27] ,
    \Tile_X6Y0_FrameData_O[26] ,
    \Tile_X6Y0_FrameData_O[25] ,
    \Tile_X6Y0_FrameData_O[24] ,
    \Tile_X6Y0_FrameData_O[23] ,
    \Tile_X6Y0_FrameData_O[22] ,
    \Tile_X6Y0_FrameData_O[21] ,
    \Tile_X6Y0_FrameData_O[20] ,
    \Tile_X6Y0_FrameData_O[19] ,
    \Tile_X6Y0_FrameData_O[18] ,
    \Tile_X6Y0_FrameData_O[17] ,
    \Tile_X6Y0_FrameData_O[16] ,
    \Tile_X6Y0_FrameData_O[15] ,
    \Tile_X6Y0_FrameData_O[14] ,
    \Tile_X6Y0_FrameData_O[13] ,
    \Tile_X6Y0_FrameData_O[12] ,
    \Tile_X6Y0_FrameData_O[11] ,
    \Tile_X6Y0_FrameData_O[10] ,
    \Tile_X6Y0_FrameData_O[9] ,
    \Tile_X6Y0_FrameData_O[8] ,
    \Tile_X6Y0_FrameData_O[7] ,
    \Tile_X6Y0_FrameData_O[6] ,
    \Tile_X6Y0_FrameData_O[5] ,
    \Tile_X6Y0_FrameData_O[4] ,
    \Tile_X6Y0_FrameData_O[3] ,
    \Tile_X6Y0_FrameData_O[2] ,
    \Tile_X6Y0_FrameData_O[1] ,
    \Tile_X6Y0_FrameData_O[0] }),
    .FrameStrobe({\Tile_X6Y1_FrameStrobe_O[19] ,
    \Tile_X6Y1_FrameStrobe_O[18] ,
    \Tile_X6Y1_FrameStrobe_O[17] ,
    \Tile_X6Y1_FrameStrobe_O[16] ,
    \Tile_X6Y1_FrameStrobe_O[15] ,
    \Tile_X6Y1_FrameStrobe_O[14] ,
    \Tile_X6Y1_FrameStrobe_O[13] ,
    \Tile_X6Y1_FrameStrobe_O[12] ,
    \Tile_X6Y1_FrameStrobe_O[11] ,
    \Tile_X6Y1_FrameStrobe_O[10] ,
    \Tile_X6Y1_FrameStrobe_O[9] ,
    \Tile_X6Y1_FrameStrobe_O[8] ,
    \Tile_X6Y1_FrameStrobe_O[7] ,
    \Tile_X6Y1_FrameStrobe_O[6] ,
    \Tile_X6Y1_FrameStrobe_O[5] ,
    \Tile_X6Y1_FrameStrobe_O[4] ,
    \Tile_X6Y1_FrameStrobe_O[3] ,
    \Tile_X6Y1_FrameStrobe_O[2] ,
    \Tile_X6Y1_FrameStrobe_O[1] ,
    \Tile_X6Y1_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X6Y0_FrameStrobe_O[19] ,
    \Tile_X6Y0_FrameStrobe_O[18] ,
    \Tile_X6Y0_FrameStrobe_O[17] ,
    \Tile_X6Y0_FrameStrobe_O[16] ,
    \Tile_X6Y0_FrameStrobe_O[15] ,
    \Tile_X6Y0_FrameStrobe_O[14] ,
    \Tile_X6Y0_FrameStrobe_O[13] ,
    \Tile_X6Y0_FrameStrobe_O[12] ,
    \Tile_X6Y0_FrameStrobe_O[11] ,
    \Tile_X6Y0_FrameStrobe_O[10] ,
    \Tile_X6Y0_FrameStrobe_O[9] ,
    \Tile_X6Y0_FrameStrobe_O[8] ,
    \Tile_X6Y0_FrameStrobe_O[7] ,
    \Tile_X6Y0_FrameStrobe_O[6] ,
    \Tile_X6Y0_FrameStrobe_O[5] ,
    \Tile_X6Y0_FrameStrobe_O[4] ,
    \Tile_X6Y0_FrameStrobe_O[3] ,
    \Tile_X6Y0_FrameStrobe_O[2] ,
    \Tile_X6Y0_FrameStrobe_O[1] ,
    \Tile_X6Y0_FrameStrobe_O[0] }),
    .N1END({\Tile_X6Y1_N1BEG[3] ,
    \Tile_X6Y1_N1BEG[2] ,
    \Tile_X6Y1_N1BEG[1] ,
    \Tile_X6Y1_N1BEG[0] }),
    .N2END({\Tile_X6Y1_N2BEGb[7] ,
    \Tile_X6Y1_N2BEGb[6] ,
    \Tile_X6Y1_N2BEGb[5] ,
    \Tile_X6Y1_N2BEGb[4] ,
    \Tile_X6Y1_N2BEGb[3] ,
    \Tile_X6Y1_N2BEGb[2] ,
    \Tile_X6Y1_N2BEGb[1] ,
    \Tile_X6Y1_N2BEGb[0] }),
    .N2MID({\Tile_X6Y1_N2BEG[7] ,
    \Tile_X6Y1_N2BEG[6] ,
    \Tile_X6Y1_N2BEG[5] ,
    \Tile_X6Y1_N2BEG[4] ,
    \Tile_X6Y1_N2BEG[3] ,
    \Tile_X6Y1_N2BEG[2] ,
    \Tile_X6Y1_N2BEG[1] ,
    \Tile_X6Y1_N2BEG[0] }),
    .N4END({\Tile_X6Y1_N4BEG[15] ,
    \Tile_X6Y1_N4BEG[14] ,
    \Tile_X6Y1_N4BEG[13] ,
    \Tile_X6Y1_N4BEG[12] ,
    \Tile_X6Y1_N4BEG[11] ,
    \Tile_X6Y1_N4BEG[10] ,
    \Tile_X6Y1_N4BEG[9] ,
    \Tile_X6Y1_N4BEG[8] ,
    \Tile_X6Y1_N4BEG[7] ,
    \Tile_X6Y1_N4BEG[6] ,
    \Tile_X6Y1_N4BEG[5] ,
    \Tile_X6Y1_N4BEG[4] ,
    \Tile_X6Y1_N4BEG[3] ,
    \Tile_X6Y1_N4BEG[2] ,
    \Tile_X6Y1_N4BEG[1] ,
    \Tile_X6Y1_N4BEG[0] }),
    .NN4END({\Tile_X6Y1_NN4BEG[15] ,
    \Tile_X6Y1_NN4BEG[14] ,
    \Tile_X6Y1_NN4BEG[13] ,
    \Tile_X6Y1_NN4BEG[12] ,
    \Tile_X6Y1_NN4BEG[11] ,
    \Tile_X6Y1_NN4BEG[10] ,
    \Tile_X6Y1_NN4BEG[9] ,
    \Tile_X6Y1_NN4BEG[8] ,
    \Tile_X6Y1_NN4BEG[7] ,
    \Tile_X6Y1_NN4BEG[6] ,
    \Tile_X6Y1_NN4BEG[5] ,
    \Tile_X6Y1_NN4BEG[4] ,
    \Tile_X6Y1_NN4BEG[3] ,
    \Tile_X6Y1_NN4BEG[2] ,
    \Tile_X6Y1_NN4BEG[1] ,
    \Tile_X6Y1_NN4BEG[0] }),
    .S1BEG({\Tile_X6Y0_S1BEG[3] ,
    \Tile_X6Y0_S1BEG[2] ,
    \Tile_X6Y0_S1BEG[1] ,
    \Tile_X6Y0_S1BEG[0] }),
    .S2BEG({\Tile_X6Y0_S2BEG[7] ,
    \Tile_X6Y0_S2BEG[6] ,
    \Tile_X6Y0_S2BEG[5] ,
    \Tile_X6Y0_S2BEG[4] ,
    \Tile_X6Y0_S2BEG[3] ,
    \Tile_X6Y0_S2BEG[2] ,
    \Tile_X6Y0_S2BEG[1] ,
    \Tile_X6Y0_S2BEG[0] }),
    .S2BEGb({\Tile_X6Y0_S2BEGb[7] ,
    \Tile_X6Y0_S2BEGb[6] ,
    \Tile_X6Y0_S2BEGb[5] ,
    \Tile_X6Y0_S2BEGb[4] ,
    \Tile_X6Y0_S2BEGb[3] ,
    \Tile_X6Y0_S2BEGb[2] ,
    \Tile_X6Y0_S2BEGb[1] ,
    \Tile_X6Y0_S2BEGb[0] }),
    .S4BEG({\Tile_X6Y0_S4BEG[15] ,
    \Tile_X6Y0_S4BEG[14] ,
    \Tile_X6Y0_S4BEG[13] ,
    \Tile_X6Y0_S4BEG[12] ,
    \Tile_X6Y0_S4BEG[11] ,
    \Tile_X6Y0_S4BEG[10] ,
    \Tile_X6Y0_S4BEG[9] ,
    \Tile_X6Y0_S4BEG[8] ,
    \Tile_X6Y0_S4BEG[7] ,
    \Tile_X6Y0_S4BEG[6] ,
    \Tile_X6Y0_S4BEG[5] ,
    \Tile_X6Y0_S4BEG[4] ,
    \Tile_X6Y0_S4BEG[3] ,
    \Tile_X6Y0_S4BEG[2] ,
    \Tile_X6Y0_S4BEG[1] ,
    \Tile_X6Y0_S4BEG[0] }),
    .SS4BEG({\Tile_X6Y0_SS4BEG[15] ,
    \Tile_X6Y0_SS4BEG[14] ,
    \Tile_X6Y0_SS4BEG[13] ,
    \Tile_X6Y0_SS4BEG[12] ,
    \Tile_X6Y0_SS4BEG[11] ,
    \Tile_X6Y0_SS4BEG[10] ,
    \Tile_X6Y0_SS4BEG[9] ,
    \Tile_X6Y0_SS4BEG[8] ,
    \Tile_X6Y0_SS4BEG[7] ,
    \Tile_X6Y0_SS4BEG[6] ,
    \Tile_X6Y0_SS4BEG[5] ,
    \Tile_X6Y0_SS4BEG[4] ,
    \Tile_X6Y0_SS4BEG[3] ,
    \Tile_X6Y0_SS4BEG[2] ,
    \Tile_X6Y0_SS4BEG[1] ,
    \Tile_X6Y0_SS4BEG[0] }));
 LUT4AB Tile_X6Y10_LUT4AB (.Ci(Tile_X6Y11_Co),
    .Co(Tile_X6Y10_Co),
    .UserCLK(Tile_X6Y11_UserCLKo),
    .UserCLKo(Tile_X6Y10_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X6Y10_E1BEG[3] ,
    \Tile_X6Y10_E1BEG[2] ,
    \Tile_X6Y10_E1BEG[1] ,
    \Tile_X6Y10_E1BEG[0] }),
    .E1END({\Tile_X5Y10_E1BEG[3] ,
    \Tile_X5Y10_E1BEG[2] ,
    \Tile_X5Y10_E1BEG[1] ,
    \Tile_X5Y10_E1BEG[0] }),
    .E2BEG({\Tile_X6Y10_E2BEG[7] ,
    \Tile_X6Y10_E2BEG[6] ,
    \Tile_X6Y10_E2BEG[5] ,
    \Tile_X6Y10_E2BEG[4] ,
    \Tile_X6Y10_E2BEG[3] ,
    \Tile_X6Y10_E2BEG[2] ,
    \Tile_X6Y10_E2BEG[1] ,
    \Tile_X6Y10_E2BEG[0] }),
    .E2BEGb({\Tile_X6Y10_E2BEGb[7] ,
    \Tile_X6Y10_E2BEGb[6] ,
    \Tile_X6Y10_E2BEGb[5] ,
    \Tile_X6Y10_E2BEGb[4] ,
    \Tile_X6Y10_E2BEGb[3] ,
    \Tile_X6Y10_E2BEGb[2] ,
    \Tile_X6Y10_E2BEGb[1] ,
    \Tile_X6Y10_E2BEGb[0] }),
    .E2END({\Tile_X5Y10_E2BEGb[7] ,
    \Tile_X5Y10_E2BEGb[6] ,
    \Tile_X5Y10_E2BEGb[5] ,
    \Tile_X5Y10_E2BEGb[4] ,
    \Tile_X5Y10_E2BEGb[3] ,
    \Tile_X5Y10_E2BEGb[2] ,
    \Tile_X5Y10_E2BEGb[1] ,
    \Tile_X5Y10_E2BEGb[0] }),
    .E2MID({\Tile_X5Y10_E2BEG[7] ,
    \Tile_X5Y10_E2BEG[6] ,
    \Tile_X5Y10_E2BEG[5] ,
    \Tile_X5Y10_E2BEG[4] ,
    \Tile_X5Y10_E2BEG[3] ,
    \Tile_X5Y10_E2BEG[2] ,
    \Tile_X5Y10_E2BEG[1] ,
    \Tile_X5Y10_E2BEG[0] }),
    .E6BEG({\Tile_X6Y10_E6BEG[11] ,
    \Tile_X6Y10_E6BEG[10] ,
    \Tile_X6Y10_E6BEG[9] ,
    \Tile_X6Y10_E6BEG[8] ,
    \Tile_X6Y10_E6BEG[7] ,
    \Tile_X6Y10_E6BEG[6] ,
    \Tile_X6Y10_E6BEG[5] ,
    \Tile_X6Y10_E6BEG[4] ,
    \Tile_X6Y10_E6BEG[3] ,
    \Tile_X6Y10_E6BEG[2] ,
    \Tile_X6Y10_E6BEG[1] ,
    \Tile_X6Y10_E6BEG[0] }),
    .E6END({\Tile_X5Y10_E6BEG[11] ,
    \Tile_X5Y10_E6BEG[10] ,
    \Tile_X5Y10_E6BEG[9] ,
    \Tile_X5Y10_E6BEG[8] ,
    \Tile_X5Y10_E6BEG[7] ,
    \Tile_X5Y10_E6BEG[6] ,
    \Tile_X5Y10_E6BEG[5] ,
    \Tile_X5Y10_E6BEG[4] ,
    \Tile_X5Y10_E6BEG[3] ,
    \Tile_X5Y10_E6BEG[2] ,
    \Tile_X5Y10_E6BEG[1] ,
    \Tile_X5Y10_E6BEG[0] }),
    .EE4BEG({\Tile_X6Y10_EE4BEG[15] ,
    \Tile_X6Y10_EE4BEG[14] ,
    \Tile_X6Y10_EE4BEG[13] ,
    \Tile_X6Y10_EE4BEG[12] ,
    \Tile_X6Y10_EE4BEG[11] ,
    \Tile_X6Y10_EE4BEG[10] ,
    \Tile_X6Y10_EE4BEG[9] ,
    \Tile_X6Y10_EE4BEG[8] ,
    \Tile_X6Y10_EE4BEG[7] ,
    \Tile_X6Y10_EE4BEG[6] ,
    \Tile_X6Y10_EE4BEG[5] ,
    \Tile_X6Y10_EE4BEG[4] ,
    \Tile_X6Y10_EE4BEG[3] ,
    \Tile_X6Y10_EE4BEG[2] ,
    \Tile_X6Y10_EE4BEG[1] ,
    \Tile_X6Y10_EE4BEG[0] }),
    .EE4END({\Tile_X5Y10_EE4BEG[15] ,
    \Tile_X5Y10_EE4BEG[14] ,
    \Tile_X5Y10_EE4BEG[13] ,
    \Tile_X5Y10_EE4BEG[12] ,
    \Tile_X5Y10_EE4BEG[11] ,
    \Tile_X5Y10_EE4BEG[10] ,
    \Tile_X5Y10_EE4BEG[9] ,
    \Tile_X5Y10_EE4BEG[8] ,
    \Tile_X5Y10_EE4BEG[7] ,
    \Tile_X5Y10_EE4BEG[6] ,
    \Tile_X5Y10_EE4BEG[5] ,
    \Tile_X5Y10_EE4BEG[4] ,
    \Tile_X5Y10_EE4BEG[3] ,
    \Tile_X5Y10_EE4BEG[2] ,
    \Tile_X5Y10_EE4BEG[1] ,
    \Tile_X5Y10_EE4BEG[0] }),
    .FrameData({\Tile_X5Y10_FrameData_O[31] ,
    \Tile_X5Y10_FrameData_O[30] ,
    \Tile_X5Y10_FrameData_O[29] ,
    \Tile_X5Y10_FrameData_O[28] ,
    \Tile_X5Y10_FrameData_O[27] ,
    \Tile_X5Y10_FrameData_O[26] ,
    \Tile_X5Y10_FrameData_O[25] ,
    \Tile_X5Y10_FrameData_O[24] ,
    \Tile_X5Y10_FrameData_O[23] ,
    \Tile_X5Y10_FrameData_O[22] ,
    \Tile_X5Y10_FrameData_O[21] ,
    \Tile_X5Y10_FrameData_O[20] ,
    \Tile_X5Y10_FrameData_O[19] ,
    \Tile_X5Y10_FrameData_O[18] ,
    \Tile_X5Y10_FrameData_O[17] ,
    \Tile_X5Y10_FrameData_O[16] ,
    \Tile_X5Y10_FrameData_O[15] ,
    \Tile_X5Y10_FrameData_O[14] ,
    \Tile_X5Y10_FrameData_O[13] ,
    \Tile_X5Y10_FrameData_O[12] ,
    \Tile_X5Y10_FrameData_O[11] ,
    \Tile_X5Y10_FrameData_O[10] ,
    \Tile_X5Y10_FrameData_O[9] ,
    \Tile_X5Y10_FrameData_O[8] ,
    \Tile_X5Y10_FrameData_O[7] ,
    \Tile_X5Y10_FrameData_O[6] ,
    \Tile_X5Y10_FrameData_O[5] ,
    \Tile_X5Y10_FrameData_O[4] ,
    \Tile_X5Y10_FrameData_O[3] ,
    \Tile_X5Y10_FrameData_O[2] ,
    \Tile_X5Y10_FrameData_O[1] ,
    \Tile_X5Y10_FrameData_O[0] }),
    .FrameData_O({\Tile_X6Y10_FrameData_O[31] ,
    \Tile_X6Y10_FrameData_O[30] ,
    \Tile_X6Y10_FrameData_O[29] ,
    \Tile_X6Y10_FrameData_O[28] ,
    \Tile_X6Y10_FrameData_O[27] ,
    \Tile_X6Y10_FrameData_O[26] ,
    \Tile_X6Y10_FrameData_O[25] ,
    \Tile_X6Y10_FrameData_O[24] ,
    \Tile_X6Y10_FrameData_O[23] ,
    \Tile_X6Y10_FrameData_O[22] ,
    \Tile_X6Y10_FrameData_O[21] ,
    \Tile_X6Y10_FrameData_O[20] ,
    \Tile_X6Y10_FrameData_O[19] ,
    \Tile_X6Y10_FrameData_O[18] ,
    \Tile_X6Y10_FrameData_O[17] ,
    \Tile_X6Y10_FrameData_O[16] ,
    \Tile_X6Y10_FrameData_O[15] ,
    \Tile_X6Y10_FrameData_O[14] ,
    \Tile_X6Y10_FrameData_O[13] ,
    \Tile_X6Y10_FrameData_O[12] ,
    \Tile_X6Y10_FrameData_O[11] ,
    \Tile_X6Y10_FrameData_O[10] ,
    \Tile_X6Y10_FrameData_O[9] ,
    \Tile_X6Y10_FrameData_O[8] ,
    \Tile_X6Y10_FrameData_O[7] ,
    \Tile_X6Y10_FrameData_O[6] ,
    \Tile_X6Y10_FrameData_O[5] ,
    \Tile_X6Y10_FrameData_O[4] ,
    \Tile_X6Y10_FrameData_O[3] ,
    \Tile_X6Y10_FrameData_O[2] ,
    \Tile_X6Y10_FrameData_O[1] ,
    \Tile_X6Y10_FrameData_O[0] }),
    .FrameStrobe({\Tile_X6Y11_FrameStrobe_O[19] ,
    \Tile_X6Y11_FrameStrobe_O[18] ,
    \Tile_X6Y11_FrameStrobe_O[17] ,
    \Tile_X6Y11_FrameStrobe_O[16] ,
    \Tile_X6Y11_FrameStrobe_O[15] ,
    \Tile_X6Y11_FrameStrobe_O[14] ,
    \Tile_X6Y11_FrameStrobe_O[13] ,
    \Tile_X6Y11_FrameStrobe_O[12] ,
    \Tile_X6Y11_FrameStrobe_O[11] ,
    \Tile_X6Y11_FrameStrobe_O[10] ,
    \Tile_X6Y11_FrameStrobe_O[9] ,
    \Tile_X6Y11_FrameStrobe_O[8] ,
    \Tile_X6Y11_FrameStrobe_O[7] ,
    \Tile_X6Y11_FrameStrobe_O[6] ,
    \Tile_X6Y11_FrameStrobe_O[5] ,
    \Tile_X6Y11_FrameStrobe_O[4] ,
    \Tile_X6Y11_FrameStrobe_O[3] ,
    \Tile_X6Y11_FrameStrobe_O[2] ,
    \Tile_X6Y11_FrameStrobe_O[1] ,
    \Tile_X6Y11_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X6Y10_FrameStrobe_O[19] ,
    \Tile_X6Y10_FrameStrobe_O[18] ,
    \Tile_X6Y10_FrameStrobe_O[17] ,
    \Tile_X6Y10_FrameStrobe_O[16] ,
    \Tile_X6Y10_FrameStrobe_O[15] ,
    \Tile_X6Y10_FrameStrobe_O[14] ,
    \Tile_X6Y10_FrameStrobe_O[13] ,
    \Tile_X6Y10_FrameStrobe_O[12] ,
    \Tile_X6Y10_FrameStrobe_O[11] ,
    \Tile_X6Y10_FrameStrobe_O[10] ,
    \Tile_X6Y10_FrameStrobe_O[9] ,
    \Tile_X6Y10_FrameStrobe_O[8] ,
    \Tile_X6Y10_FrameStrobe_O[7] ,
    \Tile_X6Y10_FrameStrobe_O[6] ,
    \Tile_X6Y10_FrameStrobe_O[5] ,
    \Tile_X6Y10_FrameStrobe_O[4] ,
    \Tile_X6Y10_FrameStrobe_O[3] ,
    \Tile_X6Y10_FrameStrobe_O[2] ,
    \Tile_X6Y10_FrameStrobe_O[1] ,
    \Tile_X6Y10_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X6Y10_N1BEG[3] ,
    \Tile_X6Y10_N1BEG[2] ,
    \Tile_X6Y10_N1BEG[1] ,
    \Tile_X6Y10_N1BEG[0] }),
    .N1END({\Tile_X6Y11_N1BEG[3] ,
    \Tile_X6Y11_N1BEG[2] ,
    \Tile_X6Y11_N1BEG[1] ,
    \Tile_X6Y11_N1BEG[0] }),
    .N2BEG({\Tile_X6Y10_N2BEG[7] ,
    \Tile_X6Y10_N2BEG[6] ,
    \Tile_X6Y10_N2BEG[5] ,
    \Tile_X6Y10_N2BEG[4] ,
    \Tile_X6Y10_N2BEG[3] ,
    \Tile_X6Y10_N2BEG[2] ,
    \Tile_X6Y10_N2BEG[1] ,
    \Tile_X6Y10_N2BEG[0] }),
    .N2BEGb({\Tile_X6Y10_N2BEGb[7] ,
    \Tile_X6Y10_N2BEGb[6] ,
    \Tile_X6Y10_N2BEGb[5] ,
    \Tile_X6Y10_N2BEGb[4] ,
    \Tile_X6Y10_N2BEGb[3] ,
    \Tile_X6Y10_N2BEGb[2] ,
    \Tile_X6Y10_N2BEGb[1] ,
    \Tile_X6Y10_N2BEGb[0] }),
    .N2END({\Tile_X6Y11_N2BEGb[7] ,
    \Tile_X6Y11_N2BEGb[6] ,
    \Tile_X6Y11_N2BEGb[5] ,
    \Tile_X6Y11_N2BEGb[4] ,
    \Tile_X6Y11_N2BEGb[3] ,
    \Tile_X6Y11_N2BEGb[2] ,
    \Tile_X6Y11_N2BEGb[1] ,
    \Tile_X6Y11_N2BEGb[0] }),
    .N2MID({\Tile_X6Y11_N2BEG[7] ,
    \Tile_X6Y11_N2BEG[6] ,
    \Tile_X6Y11_N2BEG[5] ,
    \Tile_X6Y11_N2BEG[4] ,
    \Tile_X6Y11_N2BEG[3] ,
    \Tile_X6Y11_N2BEG[2] ,
    \Tile_X6Y11_N2BEG[1] ,
    \Tile_X6Y11_N2BEG[0] }),
    .N4BEG({\Tile_X6Y10_N4BEG[15] ,
    \Tile_X6Y10_N4BEG[14] ,
    \Tile_X6Y10_N4BEG[13] ,
    \Tile_X6Y10_N4BEG[12] ,
    \Tile_X6Y10_N4BEG[11] ,
    \Tile_X6Y10_N4BEG[10] ,
    \Tile_X6Y10_N4BEG[9] ,
    \Tile_X6Y10_N4BEG[8] ,
    \Tile_X6Y10_N4BEG[7] ,
    \Tile_X6Y10_N4BEG[6] ,
    \Tile_X6Y10_N4BEG[5] ,
    \Tile_X6Y10_N4BEG[4] ,
    \Tile_X6Y10_N4BEG[3] ,
    \Tile_X6Y10_N4BEG[2] ,
    \Tile_X6Y10_N4BEG[1] ,
    \Tile_X6Y10_N4BEG[0] }),
    .N4END({\Tile_X6Y11_N4BEG[15] ,
    \Tile_X6Y11_N4BEG[14] ,
    \Tile_X6Y11_N4BEG[13] ,
    \Tile_X6Y11_N4BEG[12] ,
    \Tile_X6Y11_N4BEG[11] ,
    \Tile_X6Y11_N4BEG[10] ,
    \Tile_X6Y11_N4BEG[9] ,
    \Tile_X6Y11_N4BEG[8] ,
    \Tile_X6Y11_N4BEG[7] ,
    \Tile_X6Y11_N4BEG[6] ,
    \Tile_X6Y11_N4BEG[5] ,
    \Tile_X6Y11_N4BEG[4] ,
    \Tile_X6Y11_N4BEG[3] ,
    \Tile_X6Y11_N4BEG[2] ,
    \Tile_X6Y11_N4BEG[1] ,
    \Tile_X6Y11_N4BEG[0] }),
    .NN4BEG({\Tile_X6Y10_NN4BEG[15] ,
    \Tile_X6Y10_NN4BEG[14] ,
    \Tile_X6Y10_NN4BEG[13] ,
    \Tile_X6Y10_NN4BEG[12] ,
    \Tile_X6Y10_NN4BEG[11] ,
    \Tile_X6Y10_NN4BEG[10] ,
    \Tile_X6Y10_NN4BEG[9] ,
    \Tile_X6Y10_NN4BEG[8] ,
    \Tile_X6Y10_NN4BEG[7] ,
    \Tile_X6Y10_NN4BEG[6] ,
    \Tile_X6Y10_NN4BEG[5] ,
    \Tile_X6Y10_NN4BEG[4] ,
    \Tile_X6Y10_NN4BEG[3] ,
    \Tile_X6Y10_NN4BEG[2] ,
    \Tile_X6Y10_NN4BEG[1] ,
    \Tile_X6Y10_NN4BEG[0] }),
    .NN4END({\Tile_X6Y11_NN4BEG[15] ,
    \Tile_X6Y11_NN4BEG[14] ,
    \Tile_X6Y11_NN4BEG[13] ,
    \Tile_X6Y11_NN4BEG[12] ,
    \Tile_X6Y11_NN4BEG[11] ,
    \Tile_X6Y11_NN4BEG[10] ,
    \Tile_X6Y11_NN4BEG[9] ,
    \Tile_X6Y11_NN4BEG[8] ,
    \Tile_X6Y11_NN4BEG[7] ,
    \Tile_X6Y11_NN4BEG[6] ,
    \Tile_X6Y11_NN4BEG[5] ,
    \Tile_X6Y11_NN4BEG[4] ,
    \Tile_X6Y11_NN4BEG[3] ,
    \Tile_X6Y11_NN4BEG[2] ,
    \Tile_X6Y11_NN4BEG[1] ,
    \Tile_X6Y11_NN4BEG[0] }),
    .S1BEG({\Tile_X6Y10_S1BEG[3] ,
    \Tile_X6Y10_S1BEG[2] ,
    \Tile_X6Y10_S1BEG[1] ,
    \Tile_X6Y10_S1BEG[0] }),
    .S1END({\Tile_X6Y9_S1BEG[3] ,
    \Tile_X6Y9_S1BEG[2] ,
    \Tile_X6Y9_S1BEG[1] ,
    \Tile_X6Y9_S1BEG[0] }),
    .S2BEG({\Tile_X6Y10_S2BEG[7] ,
    \Tile_X6Y10_S2BEG[6] ,
    \Tile_X6Y10_S2BEG[5] ,
    \Tile_X6Y10_S2BEG[4] ,
    \Tile_X6Y10_S2BEG[3] ,
    \Tile_X6Y10_S2BEG[2] ,
    \Tile_X6Y10_S2BEG[1] ,
    \Tile_X6Y10_S2BEG[0] }),
    .S2BEGb({\Tile_X6Y10_S2BEGb[7] ,
    \Tile_X6Y10_S2BEGb[6] ,
    \Tile_X6Y10_S2BEGb[5] ,
    \Tile_X6Y10_S2BEGb[4] ,
    \Tile_X6Y10_S2BEGb[3] ,
    \Tile_X6Y10_S2BEGb[2] ,
    \Tile_X6Y10_S2BEGb[1] ,
    \Tile_X6Y10_S2BEGb[0] }),
    .S2END({\Tile_X6Y9_S2BEGb[7] ,
    \Tile_X6Y9_S2BEGb[6] ,
    \Tile_X6Y9_S2BEGb[5] ,
    \Tile_X6Y9_S2BEGb[4] ,
    \Tile_X6Y9_S2BEGb[3] ,
    \Tile_X6Y9_S2BEGb[2] ,
    \Tile_X6Y9_S2BEGb[1] ,
    \Tile_X6Y9_S2BEGb[0] }),
    .S2MID({\Tile_X6Y9_S2BEG[7] ,
    \Tile_X6Y9_S2BEG[6] ,
    \Tile_X6Y9_S2BEG[5] ,
    \Tile_X6Y9_S2BEG[4] ,
    \Tile_X6Y9_S2BEG[3] ,
    \Tile_X6Y9_S2BEG[2] ,
    \Tile_X6Y9_S2BEG[1] ,
    \Tile_X6Y9_S2BEG[0] }),
    .S4BEG({\Tile_X6Y10_S4BEG[15] ,
    \Tile_X6Y10_S4BEG[14] ,
    \Tile_X6Y10_S4BEG[13] ,
    \Tile_X6Y10_S4BEG[12] ,
    \Tile_X6Y10_S4BEG[11] ,
    \Tile_X6Y10_S4BEG[10] ,
    \Tile_X6Y10_S4BEG[9] ,
    \Tile_X6Y10_S4BEG[8] ,
    \Tile_X6Y10_S4BEG[7] ,
    \Tile_X6Y10_S4BEG[6] ,
    \Tile_X6Y10_S4BEG[5] ,
    \Tile_X6Y10_S4BEG[4] ,
    \Tile_X6Y10_S4BEG[3] ,
    \Tile_X6Y10_S4BEG[2] ,
    \Tile_X6Y10_S4BEG[1] ,
    \Tile_X6Y10_S4BEG[0] }),
    .S4END({\Tile_X6Y9_S4BEG[15] ,
    \Tile_X6Y9_S4BEG[14] ,
    \Tile_X6Y9_S4BEG[13] ,
    \Tile_X6Y9_S4BEG[12] ,
    \Tile_X6Y9_S4BEG[11] ,
    \Tile_X6Y9_S4BEG[10] ,
    \Tile_X6Y9_S4BEG[9] ,
    \Tile_X6Y9_S4BEG[8] ,
    \Tile_X6Y9_S4BEG[7] ,
    \Tile_X6Y9_S4BEG[6] ,
    \Tile_X6Y9_S4BEG[5] ,
    \Tile_X6Y9_S4BEG[4] ,
    \Tile_X6Y9_S4BEG[3] ,
    \Tile_X6Y9_S4BEG[2] ,
    \Tile_X6Y9_S4BEG[1] ,
    \Tile_X6Y9_S4BEG[0] }),
    .SS4BEG({\Tile_X6Y10_SS4BEG[15] ,
    \Tile_X6Y10_SS4BEG[14] ,
    \Tile_X6Y10_SS4BEG[13] ,
    \Tile_X6Y10_SS4BEG[12] ,
    \Tile_X6Y10_SS4BEG[11] ,
    \Tile_X6Y10_SS4BEG[10] ,
    \Tile_X6Y10_SS4BEG[9] ,
    \Tile_X6Y10_SS4BEG[8] ,
    \Tile_X6Y10_SS4BEG[7] ,
    \Tile_X6Y10_SS4BEG[6] ,
    \Tile_X6Y10_SS4BEG[5] ,
    \Tile_X6Y10_SS4BEG[4] ,
    \Tile_X6Y10_SS4BEG[3] ,
    \Tile_X6Y10_SS4BEG[2] ,
    \Tile_X6Y10_SS4BEG[1] ,
    \Tile_X6Y10_SS4BEG[0] }),
    .SS4END({\Tile_X6Y9_SS4BEG[15] ,
    \Tile_X6Y9_SS4BEG[14] ,
    \Tile_X6Y9_SS4BEG[13] ,
    \Tile_X6Y9_SS4BEG[12] ,
    \Tile_X6Y9_SS4BEG[11] ,
    \Tile_X6Y9_SS4BEG[10] ,
    \Tile_X6Y9_SS4BEG[9] ,
    \Tile_X6Y9_SS4BEG[8] ,
    \Tile_X6Y9_SS4BEG[7] ,
    \Tile_X6Y9_SS4BEG[6] ,
    \Tile_X6Y9_SS4BEG[5] ,
    \Tile_X6Y9_SS4BEG[4] ,
    \Tile_X6Y9_SS4BEG[3] ,
    \Tile_X6Y9_SS4BEG[2] ,
    \Tile_X6Y9_SS4BEG[1] ,
    \Tile_X6Y9_SS4BEG[0] }),
    .W1BEG({\Tile_X6Y10_W1BEG[3] ,
    \Tile_X6Y10_W1BEG[2] ,
    \Tile_X6Y10_W1BEG[1] ,
    \Tile_X6Y10_W1BEG[0] }),
    .W1END({\Tile_X7Y10_W1BEG[3] ,
    \Tile_X7Y10_W1BEG[2] ,
    \Tile_X7Y10_W1BEG[1] ,
    \Tile_X7Y10_W1BEG[0] }),
    .W2BEG({\Tile_X6Y10_W2BEG[7] ,
    \Tile_X6Y10_W2BEG[6] ,
    \Tile_X6Y10_W2BEG[5] ,
    \Tile_X6Y10_W2BEG[4] ,
    \Tile_X6Y10_W2BEG[3] ,
    \Tile_X6Y10_W2BEG[2] ,
    \Tile_X6Y10_W2BEG[1] ,
    \Tile_X6Y10_W2BEG[0] }),
    .W2BEGb({\Tile_X6Y10_W2BEGb[7] ,
    \Tile_X6Y10_W2BEGb[6] ,
    \Tile_X6Y10_W2BEGb[5] ,
    \Tile_X6Y10_W2BEGb[4] ,
    \Tile_X6Y10_W2BEGb[3] ,
    \Tile_X6Y10_W2BEGb[2] ,
    \Tile_X6Y10_W2BEGb[1] ,
    \Tile_X6Y10_W2BEGb[0] }),
    .W2END({\Tile_X7Y10_W2BEGb[7] ,
    \Tile_X7Y10_W2BEGb[6] ,
    \Tile_X7Y10_W2BEGb[5] ,
    \Tile_X7Y10_W2BEGb[4] ,
    \Tile_X7Y10_W2BEGb[3] ,
    \Tile_X7Y10_W2BEGb[2] ,
    \Tile_X7Y10_W2BEGb[1] ,
    \Tile_X7Y10_W2BEGb[0] }),
    .W2MID({\Tile_X7Y10_W2BEG[7] ,
    \Tile_X7Y10_W2BEG[6] ,
    \Tile_X7Y10_W2BEG[5] ,
    \Tile_X7Y10_W2BEG[4] ,
    \Tile_X7Y10_W2BEG[3] ,
    \Tile_X7Y10_W2BEG[2] ,
    \Tile_X7Y10_W2BEG[1] ,
    \Tile_X7Y10_W2BEG[0] }),
    .W6BEG({\Tile_X6Y10_W6BEG[11] ,
    \Tile_X6Y10_W6BEG[10] ,
    \Tile_X6Y10_W6BEG[9] ,
    \Tile_X6Y10_W6BEG[8] ,
    \Tile_X6Y10_W6BEG[7] ,
    \Tile_X6Y10_W6BEG[6] ,
    \Tile_X6Y10_W6BEG[5] ,
    \Tile_X6Y10_W6BEG[4] ,
    \Tile_X6Y10_W6BEG[3] ,
    \Tile_X6Y10_W6BEG[2] ,
    \Tile_X6Y10_W6BEG[1] ,
    \Tile_X6Y10_W6BEG[0] }),
    .W6END({\Tile_X7Y10_W6BEG[11] ,
    \Tile_X7Y10_W6BEG[10] ,
    \Tile_X7Y10_W6BEG[9] ,
    \Tile_X7Y10_W6BEG[8] ,
    \Tile_X7Y10_W6BEG[7] ,
    \Tile_X7Y10_W6BEG[6] ,
    \Tile_X7Y10_W6BEG[5] ,
    \Tile_X7Y10_W6BEG[4] ,
    \Tile_X7Y10_W6BEG[3] ,
    \Tile_X7Y10_W6BEG[2] ,
    \Tile_X7Y10_W6BEG[1] ,
    \Tile_X7Y10_W6BEG[0] }),
    .WW4BEG({\Tile_X6Y10_WW4BEG[15] ,
    \Tile_X6Y10_WW4BEG[14] ,
    \Tile_X6Y10_WW4BEG[13] ,
    \Tile_X6Y10_WW4BEG[12] ,
    \Tile_X6Y10_WW4BEG[11] ,
    \Tile_X6Y10_WW4BEG[10] ,
    \Tile_X6Y10_WW4BEG[9] ,
    \Tile_X6Y10_WW4BEG[8] ,
    \Tile_X6Y10_WW4BEG[7] ,
    \Tile_X6Y10_WW4BEG[6] ,
    \Tile_X6Y10_WW4BEG[5] ,
    \Tile_X6Y10_WW4BEG[4] ,
    \Tile_X6Y10_WW4BEG[3] ,
    \Tile_X6Y10_WW4BEG[2] ,
    \Tile_X6Y10_WW4BEG[1] ,
    \Tile_X6Y10_WW4BEG[0] }),
    .WW4END({\Tile_X7Y10_WW4BEG[15] ,
    \Tile_X7Y10_WW4BEG[14] ,
    \Tile_X7Y10_WW4BEG[13] ,
    \Tile_X7Y10_WW4BEG[12] ,
    \Tile_X7Y10_WW4BEG[11] ,
    \Tile_X7Y10_WW4BEG[10] ,
    \Tile_X7Y10_WW4BEG[9] ,
    \Tile_X7Y10_WW4BEG[8] ,
    \Tile_X7Y10_WW4BEG[7] ,
    \Tile_X7Y10_WW4BEG[6] ,
    \Tile_X7Y10_WW4BEG[5] ,
    \Tile_X7Y10_WW4BEG[4] ,
    \Tile_X7Y10_WW4BEG[3] ,
    \Tile_X7Y10_WW4BEG[2] ,
    \Tile_X7Y10_WW4BEG[1] ,
    \Tile_X7Y10_WW4BEG[0] }));
 LUT4AB Tile_X6Y11_LUT4AB (.Ci(Tile_X6Y12_Co),
    .Co(Tile_X6Y11_Co),
    .UserCLK(Tile_X6Y12_UserCLKo),
    .UserCLKo(Tile_X6Y11_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X6Y11_E1BEG[3] ,
    \Tile_X6Y11_E1BEG[2] ,
    \Tile_X6Y11_E1BEG[1] ,
    \Tile_X6Y11_E1BEG[0] }),
    .E1END({\Tile_X5Y11_E1BEG[3] ,
    \Tile_X5Y11_E1BEG[2] ,
    \Tile_X5Y11_E1BEG[1] ,
    \Tile_X5Y11_E1BEG[0] }),
    .E2BEG({\Tile_X6Y11_E2BEG[7] ,
    \Tile_X6Y11_E2BEG[6] ,
    \Tile_X6Y11_E2BEG[5] ,
    \Tile_X6Y11_E2BEG[4] ,
    \Tile_X6Y11_E2BEG[3] ,
    \Tile_X6Y11_E2BEG[2] ,
    \Tile_X6Y11_E2BEG[1] ,
    \Tile_X6Y11_E2BEG[0] }),
    .E2BEGb({\Tile_X6Y11_E2BEGb[7] ,
    \Tile_X6Y11_E2BEGb[6] ,
    \Tile_X6Y11_E2BEGb[5] ,
    \Tile_X6Y11_E2BEGb[4] ,
    \Tile_X6Y11_E2BEGb[3] ,
    \Tile_X6Y11_E2BEGb[2] ,
    \Tile_X6Y11_E2BEGb[1] ,
    \Tile_X6Y11_E2BEGb[0] }),
    .E2END({\Tile_X5Y11_E2BEGb[7] ,
    \Tile_X5Y11_E2BEGb[6] ,
    \Tile_X5Y11_E2BEGb[5] ,
    \Tile_X5Y11_E2BEGb[4] ,
    \Tile_X5Y11_E2BEGb[3] ,
    \Tile_X5Y11_E2BEGb[2] ,
    \Tile_X5Y11_E2BEGb[1] ,
    \Tile_X5Y11_E2BEGb[0] }),
    .E2MID({\Tile_X5Y11_E2BEG[7] ,
    \Tile_X5Y11_E2BEG[6] ,
    \Tile_X5Y11_E2BEG[5] ,
    \Tile_X5Y11_E2BEG[4] ,
    \Tile_X5Y11_E2BEG[3] ,
    \Tile_X5Y11_E2BEG[2] ,
    \Tile_X5Y11_E2BEG[1] ,
    \Tile_X5Y11_E2BEG[0] }),
    .E6BEG({\Tile_X6Y11_E6BEG[11] ,
    \Tile_X6Y11_E6BEG[10] ,
    \Tile_X6Y11_E6BEG[9] ,
    \Tile_X6Y11_E6BEG[8] ,
    \Tile_X6Y11_E6BEG[7] ,
    \Tile_X6Y11_E6BEG[6] ,
    \Tile_X6Y11_E6BEG[5] ,
    \Tile_X6Y11_E6BEG[4] ,
    \Tile_X6Y11_E6BEG[3] ,
    \Tile_X6Y11_E6BEG[2] ,
    \Tile_X6Y11_E6BEG[1] ,
    \Tile_X6Y11_E6BEG[0] }),
    .E6END({\Tile_X5Y11_E6BEG[11] ,
    \Tile_X5Y11_E6BEG[10] ,
    \Tile_X5Y11_E6BEG[9] ,
    \Tile_X5Y11_E6BEG[8] ,
    \Tile_X5Y11_E6BEG[7] ,
    \Tile_X5Y11_E6BEG[6] ,
    \Tile_X5Y11_E6BEG[5] ,
    \Tile_X5Y11_E6BEG[4] ,
    \Tile_X5Y11_E6BEG[3] ,
    \Tile_X5Y11_E6BEG[2] ,
    \Tile_X5Y11_E6BEG[1] ,
    \Tile_X5Y11_E6BEG[0] }),
    .EE4BEG({\Tile_X6Y11_EE4BEG[15] ,
    \Tile_X6Y11_EE4BEG[14] ,
    \Tile_X6Y11_EE4BEG[13] ,
    \Tile_X6Y11_EE4BEG[12] ,
    \Tile_X6Y11_EE4BEG[11] ,
    \Tile_X6Y11_EE4BEG[10] ,
    \Tile_X6Y11_EE4BEG[9] ,
    \Tile_X6Y11_EE4BEG[8] ,
    \Tile_X6Y11_EE4BEG[7] ,
    \Tile_X6Y11_EE4BEG[6] ,
    \Tile_X6Y11_EE4BEG[5] ,
    \Tile_X6Y11_EE4BEG[4] ,
    \Tile_X6Y11_EE4BEG[3] ,
    \Tile_X6Y11_EE4BEG[2] ,
    \Tile_X6Y11_EE4BEG[1] ,
    \Tile_X6Y11_EE4BEG[0] }),
    .EE4END({\Tile_X5Y11_EE4BEG[15] ,
    \Tile_X5Y11_EE4BEG[14] ,
    \Tile_X5Y11_EE4BEG[13] ,
    \Tile_X5Y11_EE4BEG[12] ,
    \Tile_X5Y11_EE4BEG[11] ,
    \Tile_X5Y11_EE4BEG[10] ,
    \Tile_X5Y11_EE4BEG[9] ,
    \Tile_X5Y11_EE4BEG[8] ,
    \Tile_X5Y11_EE4BEG[7] ,
    \Tile_X5Y11_EE4BEG[6] ,
    \Tile_X5Y11_EE4BEG[5] ,
    \Tile_X5Y11_EE4BEG[4] ,
    \Tile_X5Y11_EE4BEG[3] ,
    \Tile_X5Y11_EE4BEG[2] ,
    \Tile_X5Y11_EE4BEG[1] ,
    \Tile_X5Y11_EE4BEG[0] }),
    .FrameData({\Tile_X5Y11_FrameData_O[31] ,
    \Tile_X5Y11_FrameData_O[30] ,
    \Tile_X5Y11_FrameData_O[29] ,
    \Tile_X5Y11_FrameData_O[28] ,
    \Tile_X5Y11_FrameData_O[27] ,
    \Tile_X5Y11_FrameData_O[26] ,
    \Tile_X5Y11_FrameData_O[25] ,
    \Tile_X5Y11_FrameData_O[24] ,
    \Tile_X5Y11_FrameData_O[23] ,
    \Tile_X5Y11_FrameData_O[22] ,
    \Tile_X5Y11_FrameData_O[21] ,
    \Tile_X5Y11_FrameData_O[20] ,
    \Tile_X5Y11_FrameData_O[19] ,
    \Tile_X5Y11_FrameData_O[18] ,
    \Tile_X5Y11_FrameData_O[17] ,
    \Tile_X5Y11_FrameData_O[16] ,
    \Tile_X5Y11_FrameData_O[15] ,
    \Tile_X5Y11_FrameData_O[14] ,
    \Tile_X5Y11_FrameData_O[13] ,
    \Tile_X5Y11_FrameData_O[12] ,
    \Tile_X5Y11_FrameData_O[11] ,
    \Tile_X5Y11_FrameData_O[10] ,
    \Tile_X5Y11_FrameData_O[9] ,
    \Tile_X5Y11_FrameData_O[8] ,
    \Tile_X5Y11_FrameData_O[7] ,
    \Tile_X5Y11_FrameData_O[6] ,
    \Tile_X5Y11_FrameData_O[5] ,
    \Tile_X5Y11_FrameData_O[4] ,
    \Tile_X5Y11_FrameData_O[3] ,
    \Tile_X5Y11_FrameData_O[2] ,
    \Tile_X5Y11_FrameData_O[1] ,
    \Tile_X5Y11_FrameData_O[0] }),
    .FrameData_O({\Tile_X6Y11_FrameData_O[31] ,
    \Tile_X6Y11_FrameData_O[30] ,
    \Tile_X6Y11_FrameData_O[29] ,
    \Tile_X6Y11_FrameData_O[28] ,
    \Tile_X6Y11_FrameData_O[27] ,
    \Tile_X6Y11_FrameData_O[26] ,
    \Tile_X6Y11_FrameData_O[25] ,
    \Tile_X6Y11_FrameData_O[24] ,
    \Tile_X6Y11_FrameData_O[23] ,
    \Tile_X6Y11_FrameData_O[22] ,
    \Tile_X6Y11_FrameData_O[21] ,
    \Tile_X6Y11_FrameData_O[20] ,
    \Tile_X6Y11_FrameData_O[19] ,
    \Tile_X6Y11_FrameData_O[18] ,
    \Tile_X6Y11_FrameData_O[17] ,
    \Tile_X6Y11_FrameData_O[16] ,
    \Tile_X6Y11_FrameData_O[15] ,
    \Tile_X6Y11_FrameData_O[14] ,
    \Tile_X6Y11_FrameData_O[13] ,
    \Tile_X6Y11_FrameData_O[12] ,
    \Tile_X6Y11_FrameData_O[11] ,
    \Tile_X6Y11_FrameData_O[10] ,
    \Tile_X6Y11_FrameData_O[9] ,
    \Tile_X6Y11_FrameData_O[8] ,
    \Tile_X6Y11_FrameData_O[7] ,
    \Tile_X6Y11_FrameData_O[6] ,
    \Tile_X6Y11_FrameData_O[5] ,
    \Tile_X6Y11_FrameData_O[4] ,
    \Tile_X6Y11_FrameData_O[3] ,
    \Tile_X6Y11_FrameData_O[2] ,
    \Tile_X6Y11_FrameData_O[1] ,
    \Tile_X6Y11_FrameData_O[0] }),
    .FrameStrobe({\Tile_X6Y12_FrameStrobe_O[19] ,
    \Tile_X6Y12_FrameStrobe_O[18] ,
    \Tile_X6Y12_FrameStrobe_O[17] ,
    \Tile_X6Y12_FrameStrobe_O[16] ,
    \Tile_X6Y12_FrameStrobe_O[15] ,
    \Tile_X6Y12_FrameStrobe_O[14] ,
    \Tile_X6Y12_FrameStrobe_O[13] ,
    \Tile_X6Y12_FrameStrobe_O[12] ,
    \Tile_X6Y12_FrameStrobe_O[11] ,
    \Tile_X6Y12_FrameStrobe_O[10] ,
    \Tile_X6Y12_FrameStrobe_O[9] ,
    \Tile_X6Y12_FrameStrobe_O[8] ,
    \Tile_X6Y12_FrameStrobe_O[7] ,
    \Tile_X6Y12_FrameStrobe_O[6] ,
    \Tile_X6Y12_FrameStrobe_O[5] ,
    \Tile_X6Y12_FrameStrobe_O[4] ,
    \Tile_X6Y12_FrameStrobe_O[3] ,
    \Tile_X6Y12_FrameStrobe_O[2] ,
    \Tile_X6Y12_FrameStrobe_O[1] ,
    \Tile_X6Y12_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X6Y11_FrameStrobe_O[19] ,
    \Tile_X6Y11_FrameStrobe_O[18] ,
    \Tile_X6Y11_FrameStrobe_O[17] ,
    \Tile_X6Y11_FrameStrobe_O[16] ,
    \Tile_X6Y11_FrameStrobe_O[15] ,
    \Tile_X6Y11_FrameStrobe_O[14] ,
    \Tile_X6Y11_FrameStrobe_O[13] ,
    \Tile_X6Y11_FrameStrobe_O[12] ,
    \Tile_X6Y11_FrameStrobe_O[11] ,
    \Tile_X6Y11_FrameStrobe_O[10] ,
    \Tile_X6Y11_FrameStrobe_O[9] ,
    \Tile_X6Y11_FrameStrobe_O[8] ,
    \Tile_X6Y11_FrameStrobe_O[7] ,
    \Tile_X6Y11_FrameStrobe_O[6] ,
    \Tile_X6Y11_FrameStrobe_O[5] ,
    \Tile_X6Y11_FrameStrobe_O[4] ,
    \Tile_X6Y11_FrameStrobe_O[3] ,
    \Tile_X6Y11_FrameStrobe_O[2] ,
    \Tile_X6Y11_FrameStrobe_O[1] ,
    \Tile_X6Y11_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X6Y11_N1BEG[3] ,
    \Tile_X6Y11_N1BEG[2] ,
    \Tile_X6Y11_N1BEG[1] ,
    \Tile_X6Y11_N1BEG[0] }),
    .N1END({\Tile_X6Y12_N1BEG[3] ,
    \Tile_X6Y12_N1BEG[2] ,
    \Tile_X6Y12_N1BEG[1] ,
    \Tile_X6Y12_N1BEG[0] }),
    .N2BEG({\Tile_X6Y11_N2BEG[7] ,
    \Tile_X6Y11_N2BEG[6] ,
    \Tile_X6Y11_N2BEG[5] ,
    \Tile_X6Y11_N2BEG[4] ,
    \Tile_X6Y11_N2BEG[3] ,
    \Tile_X6Y11_N2BEG[2] ,
    \Tile_X6Y11_N2BEG[1] ,
    \Tile_X6Y11_N2BEG[0] }),
    .N2BEGb({\Tile_X6Y11_N2BEGb[7] ,
    \Tile_X6Y11_N2BEGb[6] ,
    \Tile_X6Y11_N2BEGb[5] ,
    \Tile_X6Y11_N2BEGb[4] ,
    \Tile_X6Y11_N2BEGb[3] ,
    \Tile_X6Y11_N2BEGb[2] ,
    \Tile_X6Y11_N2BEGb[1] ,
    \Tile_X6Y11_N2BEGb[0] }),
    .N2END({\Tile_X6Y12_N2BEGb[7] ,
    \Tile_X6Y12_N2BEGb[6] ,
    \Tile_X6Y12_N2BEGb[5] ,
    \Tile_X6Y12_N2BEGb[4] ,
    \Tile_X6Y12_N2BEGb[3] ,
    \Tile_X6Y12_N2BEGb[2] ,
    \Tile_X6Y12_N2BEGb[1] ,
    \Tile_X6Y12_N2BEGb[0] }),
    .N2MID({\Tile_X6Y12_N2BEG[7] ,
    \Tile_X6Y12_N2BEG[6] ,
    \Tile_X6Y12_N2BEG[5] ,
    \Tile_X6Y12_N2BEG[4] ,
    \Tile_X6Y12_N2BEG[3] ,
    \Tile_X6Y12_N2BEG[2] ,
    \Tile_X6Y12_N2BEG[1] ,
    \Tile_X6Y12_N2BEG[0] }),
    .N4BEG({\Tile_X6Y11_N4BEG[15] ,
    \Tile_X6Y11_N4BEG[14] ,
    \Tile_X6Y11_N4BEG[13] ,
    \Tile_X6Y11_N4BEG[12] ,
    \Tile_X6Y11_N4BEG[11] ,
    \Tile_X6Y11_N4BEG[10] ,
    \Tile_X6Y11_N4BEG[9] ,
    \Tile_X6Y11_N4BEG[8] ,
    \Tile_X6Y11_N4BEG[7] ,
    \Tile_X6Y11_N4BEG[6] ,
    \Tile_X6Y11_N4BEG[5] ,
    \Tile_X6Y11_N4BEG[4] ,
    \Tile_X6Y11_N4BEG[3] ,
    \Tile_X6Y11_N4BEG[2] ,
    \Tile_X6Y11_N4BEG[1] ,
    \Tile_X6Y11_N4BEG[0] }),
    .N4END({\Tile_X6Y12_N4BEG[15] ,
    \Tile_X6Y12_N4BEG[14] ,
    \Tile_X6Y12_N4BEG[13] ,
    \Tile_X6Y12_N4BEG[12] ,
    \Tile_X6Y12_N4BEG[11] ,
    \Tile_X6Y12_N4BEG[10] ,
    \Tile_X6Y12_N4BEG[9] ,
    \Tile_X6Y12_N4BEG[8] ,
    \Tile_X6Y12_N4BEG[7] ,
    \Tile_X6Y12_N4BEG[6] ,
    \Tile_X6Y12_N4BEG[5] ,
    \Tile_X6Y12_N4BEG[4] ,
    \Tile_X6Y12_N4BEG[3] ,
    \Tile_X6Y12_N4BEG[2] ,
    \Tile_X6Y12_N4BEG[1] ,
    \Tile_X6Y12_N4BEG[0] }),
    .NN4BEG({\Tile_X6Y11_NN4BEG[15] ,
    \Tile_X6Y11_NN4BEG[14] ,
    \Tile_X6Y11_NN4BEG[13] ,
    \Tile_X6Y11_NN4BEG[12] ,
    \Tile_X6Y11_NN4BEG[11] ,
    \Tile_X6Y11_NN4BEG[10] ,
    \Tile_X6Y11_NN4BEG[9] ,
    \Tile_X6Y11_NN4BEG[8] ,
    \Tile_X6Y11_NN4BEG[7] ,
    \Tile_X6Y11_NN4BEG[6] ,
    \Tile_X6Y11_NN4BEG[5] ,
    \Tile_X6Y11_NN4BEG[4] ,
    \Tile_X6Y11_NN4BEG[3] ,
    \Tile_X6Y11_NN4BEG[2] ,
    \Tile_X6Y11_NN4BEG[1] ,
    \Tile_X6Y11_NN4BEG[0] }),
    .NN4END({\Tile_X6Y12_NN4BEG[15] ,
    \Tile_X6Y12_NN4BEG[14] ,
    \Tile_X6Y12_NN4BEG[13] ,
    \Tile_X6Y12_NN4BEG[12] ,
    \Tile_X6Y12_NN4BEG[11] ,
    \Tile_X6Y12_NN4BEG[10] ,
    \Tile_X6Y12_NN4BEG[9] ,
    \Tile_X6Y12_NN4BEG[8] ,
    \Tile_X6Y12_NN4BEG[7] ,
    \Tile_X6Y12_NN4BEG[6] ,
    \Tile_X6Y12_NN4BEG[5] ,
    \Tile_X6Y12_NN4BEG[4] ,
    \Tile_X6Y12_NN4BEG[3] ,
    \Tile_X6Y12_NN4BEG[2] ,
    \Tile_X6Y12_NN4BEG[1] ,
    \Tile_X6Y12_NN4BEG[0] }),
    .S1BEG({\Tile_X6Y11_S1BEG[3] ,
    \Tile_X6Y11_S1BEG[2] ,
    \Tile_X6Y11_S1BEG[1] ,
    \Tile_X6Y11_S1BEG[0] }),
    .S1END({\Tile_X6Y10_S1BEG[3] ,
    \Tile_X6Y10_S1BEG[2] ,
    \Tile_X6Y10_S1BEG[1] ,
    \Tile_X6Y10_S1BEG[0] }),
    .S2BEG({\Tile_X6Y11_S2BEG[7] ,
    \Tile_X6Y11_S2BEG[6] ,
    \Tile_X6Y11_S2BEG[5] ,
    \Tile_X6Y11_S2BEG[4] ,
    \Tile_X6Y11_S2BEG[3] ,
    \Tile_X6Y11_S2BEG[2] ,
    \Tile_X6Y11_S2BEG[1] ,
    \Tile_X6Y11_S2BEG[0] }),
    .S2BEGb({\Tile_X6Y11_S2BEGb[7] ,
    \Tile_X6Y11_S2BEGb[6] ,
    \Tile_X6Y11_S2BEGb[5] ,
    \Tile_X6Y11_S2BEGb[4] ,
    \Tile_X6Y11_S2BEGb[3] ,
    \Tile_X6Y11_S2BEGb[2] ,
    \Tile_X6Y11_S2BEGb[1] ,
    \Tile_X6Y11_S2BEGb[0] }),
    .S2END({\Tile_X6Y10_S2BEGb[7] ,
    \Tile_X6Y10_S2BEGb[6] ,
    \Tile_X6Y10_S2BEGb[5] ,
    \Tile_X6Y10_S2BEGb[4] ,
    \Tile_X6Y10_S2BEGb[3] ,
    \Tile_X6Y10_S2BEGb[2] ,
    \Tile_X6Y10_S2BEGb[1] ,
    \Tile_X6Y10_S2BEGb[0] }),
    .S2MID({\Tile_X6Y10_S2BEG[7] ,
    \Tile_X6Y10_S2BEG[6] ,
    \Tile_X6Y10_S2BEG[5] ,
    \Tile_X6Y10_S2BEG[4] ,
    \Tile_X6Y10_S2BEG[3] ,
    \Tile_X6Y10_S2BEG[2] ,
    \Tile_X6Y10_S2BEG[1] ,
    \Tile_X6Y10_S2BEG[0] }),
    .S4BEG({\Tile_X6Y11_S4BEG[15] ,
    \Tile_X6Y11_S4BEG[14] ,
    \Tile_X6Y11_S4BEG[13] ,
    \Tile_X6Y11_S4BEG[12] ,
    \Tile_X6Y11_S4BEG[11] ,
    \Tile_X6Y11_S4BEG[10] ,
    \Tile_X6Y11_S4BEG[9] ,
    \Tile_X6Y11_S4BEG[8] ,
    \Tile_X6Y11_S4BEG[7] ,
    \Tile_X6Y11_S4BEG[6] ,
    \Tile_X6Y11_S4BEG[5] ,
    \Tile_X6Y11_S4BEG[4] ,
    \Tile_X6Y11_S4BEG[3] ,
    \Tile_X6Y11_S4BEG[2] ,
    \Tile_X6Y11_S4BEG[1] ,
    \Tile_X6Y11_S4BEG[0] }),
    .S4END({\Tile_X6Y10_S4BEG[15] ,
    \Tile_X6Y10_S4BEG[14] ,
    \Tile_X6Y10_S4BEG[13] ,
    \Tile_X6Y10_S4BEG[12] ,
    \Tile_X6Y10_S4BEG[11] ,
    \Tile_X6Y10_S4BEG[10] ,
    \Tile_X6Y10_S4BEG[9] ,
    \Tile_X6Y10_S4BEG[8] ,
    \Tile_X6Y10_S4BEG[7] ,
    \Tile_X6Y10_S4BEG[6] ,
    \Tile_X6Y10_S4BEG[5] ,
    \Tile_X6Y10_S4BEG[4] ,
    \Tile_X6Y10_S4BEG[3] ,
    \Tile_X6Y10_S4BEG[2] ,
    \Tile_X6Y10_S4BEG[1] ,
    \Tile_X6Y10_S4BEG[0] }),
    .SS4BEG({\Tile_X6Y11_SS4BEG[15] ,
    \Tile_X6Y11_SS4BEG[14] ,
    \Tile_X6Y11_SS4BEG[13] ,
    \Tile_X6Y11_SS4BEG[12] ,
    \Tile_X6Y11_SS4BEG[11] ,
    \Tile_X6Y11_SS4BEG[10] ,
    \Tile_X6Y11_SS4BEG[9] ,
    \Tile_X6Y11_SS4BEG[8] ,
    \Tile_X6Y11_SS4BEG[7] ,
    \Tile_X6Y11_SS4BEG[6] ,
    \Tile_X6Y11_SS4BEG[5] ,
    \Tile_X6Y11_SS4BEG[4] ,
    \Tile_X6Y11_SS4BEG[3] ,
    \Tile_X6Y11_SS4BEG[2] ,
    \Tile_X6Y11_SS4BEG[1] ,
    \Tile_X6Y11_SS4BEG[0] }),
    .SS4END({\Tile_X6Y10_SS4BEG[15] ,
    \Tile_X6Y10_SS4BEG[14] ,
    \Tile_X6Y10_SS4BEG[13] ,
    \Tile_X6Y10_SS4BEG[12] ,
    \Tile_X6Y10_SS4BEG[11] ,
    \Tile_X6Y10_SS4BEG[10] ,
    \Tile_X6Y10_SS4BEG[9] ,
    \Tile_X6Y10_SS4BEG[8] ,
    \Tile_X6Y10_SS4BEG[7] ,
    \Tile_X6Y10_SS4BEG[6] ,
    \Tile_X6Y10_SS4BEG[5] ,
    \Tile_X6Y10_SS4BEG[4] ,
    \Tile_X6Y10_SS4BEG[3] ,
    \Tile_X6Y10_SS4BEG[2] ,
    \Tile_X6Y10_SS4BEG[1] ,
    \Tile_X6Y10_SS4BEG[0] }),
    .W1BEG({\Tile_X6Y11_W1BEG[3] ,
    \Tile_X6Y11_W1BEG[2] ,
    \Tile_X6Y11_W1BEG[1] ,
    \Tile_X6Y11_W1BEG[0] }),
    .W1END({\Tile_X7Y11_W1BEG[3] ,
    \Tile_X7Y11_W1BEG[2] ,
    \Tile_X7Y11_W1BEG[1] ,
    \Tile_X7Y11_W1BEG[0] }),
    .W2BEG({\Tile_X6Y11_W2BEG[7] ,
    \Tile_X6Y11_W2BEG[6] ,
    \Tile_X6Y11_W2BEG[5] ,
    \Tile_X6Y11_W2BEG[4] ,
    \Tile_X6Y11_W2BEG[3] ,
    \Tile_X6Y11_W2BEG[2] ,
    \Tile_X6Y11_W2BEG[1] ,
    \Tile_X6Y11_W2BEG[0] }),
    .W2BEGb({\Tile_X6Y11_W2BEGb[7] ,
    \Tile_X6Y11_W2BEGb[6] ,
    \Tile_X6Y11_W2BEGb[5] ,
    \Tile_X6Y11_W2BEGb[4] ,
    \Tile_X6Y11_W2BEGb[3] ,
    \Tile_X6Y11_W2BEGb[2] ,
    \Tile_X6Y11_W2BEGb[1] ,
    \Tile_X6Y11_W2BEGb[0] }),
    .W2END({\Tile_X7Y11_W2BEGb[7] ,
    \Tile_X7Y11_W2BEGb[6] ,
    \Tile_X7Y11_W2BEGb[5] ,
    \Tile_X7Y11_W2BEGb[4] ,
    \Tile_X7Y11_W2BEGb[3] ,
    \Tile_X7Y11_W2BEGb[2] ,
    \Tile_X7Y11_W2BEGb[1] ,
    \Tile_X7Y11_W2BEGb[0] }),
    .W2MID({\Tile_X7Y11_W2BEG[7] ,
    \Tile_X7Y11_W2BEG[6] ,
    \Tile_X7Y11_W2BEG[5] ,
    \Tile_X7Y11_W2BEG[4] ,
    \Tile_X7Y11_W2BEG[3] ,
    \Tile_X7Y11_W2BEG[2] ,
    \Tile_X7Y11_W2BEG[1] ,
    \Tile_X7Y11_W2BEG[0] }),
    .W6BEG({\Tile_X6Y11_W6BEG[11] ,
    \Tile_X6Y11_W6BEG[10] ,
    \Tile_X6Y11_W6BEG[9] ,
    \Tile_X6Y11_W6BEG[8] ,
    \Tile_X6Y11_W6BEG[7] ,
    \Tile_X6Y11_W6BEG[6] ,
    \Tile_X6Y11_W6BEG[5] ,
    \Tile_X6Y11_W6BEG[4] ,
    \Tile_X6Y11_W6BEG[3] ,
    \Tile_X6Y11_W6BEG[2] ,
    \Tile_X6Y11_W6BEG[1] ,
    \Tile_X6Y11_W6BEG[0] }),
    .W6END({\Tile_X7Y11_W6BEG[11] ,
    \Tile_X7Y11_W6BEG[10] ,
    \Tile_X7Y11_W6BEG[9] ,
    \Tile_X7Y11_W6BEG[8] ,
    \Tile_X7Y11_W6BEG[7] ,
    \Tile_X7Y11_W6BEG[6] ,
    \Tile_X7Y11_W6BEG[5] ,
    \Tile_X7Y11_W6BEG[4] ,
    \Tile_X7Y11_W6BEG[3] ,
    \Tile_X7Y11_W6BEG[2] ,
    \Tile_X7Y11_W6BEG[1] ,
    \Tile_X7Y11_W6BEG[0] }),
    .WW4BEG({\Tile_X6Y11_WW4BEG[15] ,
    \Tile_X6Y11_WW4BEG[14] ,
    \Tile_X6Y11_WW4BEG[13] ,
    \Tile_X6Y11_WW4BEG[12] ,
    \Tile_X6Y11_WW4BEG[11] ,
    \Tile_X6Y11_WW4BEG[10] ,
    \Tile_X6Y11_WW4BEG[9] ,
    \Tile_X6Y11_WW4BEG[8] ,
    \Tile_X6Y11_WW4BEG[7] ,
    \Tile_X6Y11_WW4BEG[6] ,
    \Tile_X6Y11_WW4BEG[5] ,
    \Tile_X6Y11_WW4BEG[4] ,
    \Tile_X6Y11_WW4BEG[3] ,
    \Tile_X6Y11_WW4BEG[2] ,
    \Tile_X6Y11_WW4BEG[1] ,
    \Tile_X6Y11_WW4BEG[0] }),
    .WW4END({\Tile_X7Y11_WW4BEG[15] ,
    \Tile_X7Y11_WW4BEG[14] ,
    \Tile_X7Y11_WW4BEG[13] ,
    \Tile_X7Y11_WW4BEG[12] ,
    \Tile_X7Y11_WW4BEG[11] ,
    \Tile_X7Y11_WW4BEG[10] ,
    \Tile_X7Y11_WW4BEG[9] ,
    \Tile_X7Y11_WW4BEG[8] ,
    \Tile_X7Y11_WW4BEG[7] ,
    \Tile_X7Y11_WW4BEG[6] ,
    \Tile_X7Y11_WW4BEG[5] ,
    \Tile_X7Y11_WW4BEG[4] ,
    \Tile_X7Y11_WW4BEG[3] ,
    \Tile_X7Y11_WW4BEG[2] ,
    \Tile_X7Y11_WW4BEG[1] ,
    \Tile_X7Y11_WW4BEG[0] }));
 LUT4AB Tile_X6Y12_LUT4AB (.Ci(Tile_X6Y13_Co),
    .Co(Tile_X6Y12_Co),
    .UserCLK(Tile_X6Y13_UserCLKo),
    .UserCLKo(Tile_X6Y12_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X6Y12_E1BEG[3] ,
    \Tile_X6Y12_E1BEG[2] ,
    \Tile_X6Y12_E1BEG[1] ,
    \Tile_X6Y12_E1BEG[0] }),
    .E1END({\Tile_X5Y12_E1BEG[3] ,
    \Tile_X5Y12_E1BEG[2] ,
    \Tile_X5Y12_E1BEG[1] ,
    \Tile_X5Y12_E1BEG[0] }),
    .E2BEG({\Tile_X6Y12_E2BEG[7] ,
    \Tile_X6Y12_E2BEG[6] ,
    \Tile_X6Y12_E2BEG[5] ,
    \Tile_X6Y12_E2BEG[4] ,
    \Tile_X6Y12_E2BEG[3] ,
    \Tile_X6Y12_E2BEG[2] ,
    \Tile_X6Y12_E2BEG[1] ,
    \Tile_X6Y12_E2BEG[0] }),
    .E2BEGb({\Tile_X6Y12_E2BEGb[7] ,
    \Tile_X6Y12_E2BEGb[6] ,
    \Tile_X6Y12_E2BEGb[5] ,
    \Tile_X6Y12_E2BEGb[4] ,
    \Tile_X6Y12_E2BEGb[3] ,
    \Tile_X6Y12_E2BEGb[2] ,
    \Tile_X6Y12_E2BEGb[1] ,
    \Tile_X6Y12_E2BEGb[0] }),
    .E2END({\Tile_X5Y12_E2BEGb[7] ,
    \Tile_X5Y12_E2BEGb[6] ,
    \Tile_X5Y12_E2BEGb[5] ,
    \Tile_X5Y12_E2BEGb[4] ,
    \Tile_X5Y12_E2BEGb[3] ,
    \Tile_X5Y12_E2BEGb[2] ,
    \Tile_X5Y12_E2BEGb[1] ,
    \Tile_X5Y12_E2BEGb[0] }),
    .E2MID({\Tile_X5Y12_E2BEG[7] ,
    \Tile_X5Y12_E2BEG[6] ,
    \Tile_X5Y12_E2BEG[5] ,
    \Tile_X5Y12_E2BEG[4] ,
    \Tile_X5Y12_E2BEG[3] ,
    \Tile_X5Y12_E2BEG[2] ,
    \Tile_X5Y12_E2BEG[1] ,
    \Tile_X5Y12_E2BEG[0] }),
    .E6BEG({\Tile_X6Y12_E6BEG[11] ,
    \Tile_X6Y12_E6BEG[10] ,
    \Tile_X6Y12_E6BEG[9] ,
    \Tile_X6Y12_E6BEG[8] ,
    \Tile_X6Y12_E6BEG[7] ,
    \Tile_X6Y12_E6BEG[6] ,
    \Tile_X6Y12_E6BEG[5] ,
    \Tile_X6Y12_E6BEG[4] ,
    \Tile_X6Y12_E6BEG[3] ,
    \Tile_X6Y12_E6BEG[2] ,
    \Tile_X6Y12_E6BEG[1] ,
    \Tile_X6Y12_E6BEG[0] }),
    .E6END({\Tile_X5Y12_E6BEG[11] ,
    \Tile_X5Y12_E6BEG[10] ,
    \Tile_X5Y12_E6BEG[9] ,
    \Tile_X5Y12_E6BEG[8] ,
    \Tile_X5Y12_E6BEG[7] ,
    \Tile_X5Y12_E6BEG[6] ,
    \Tile_X5Y12_E6BEG[5] ,
    \Tile_X5Y12_E6BEG[4] ,
    \Tile_X5Y12_E6BEG[3] ,
    \Tile_X5Y12_E6BEG[2] ,
    \Tile_X5Y12_E6BEG[1] ,
    \Tile_X5Y12_E6BEG[0] }),
    .EE4BEG({\Tile_X6Y12_EE4BEG[15] ,
    \Tile_X6Y12_EE4BEG[14] ,
    \Tile_X6Y12_EE4BEG[13] ,
    \Tile_X6Y12_EE4BEG[12] ,
    \Tile_X6Y12_EE4BEG[11] ,
    \Tile_X6Y12_EE4BEG[10] ,
    \Tile_X6Y12_EE4BEG[9] ,
    \Tile_X6Y12_EE4BEG[8] ,
    \Tile_X6Y12_EE4BEG[7] ,
    \Tile_X6Y12_EE4BEG[6] ,
    \Tile_X6Y12_EE4BEG[5] ,
    \Tile_X6Y12_EE4BEG[4] ,
    \Tile_X6Y12_EE4BEG[3] ,
    \Tile_X6Y12_EE4BEG[2] ,
    \Tile_X6Y12_EE4BEG[1] ,
    \Tile_X6Y12_EE4BEG[0] }),
    .EE4END({\Tile_X5Y12_EE4BEG[15] ,
    \Tile_X5Y12_EE4BEG[14] ,
    \Tile_X5Y12_EE4BEG[13] ,
    \Tile_X5Y12_EE4BEG[12] ,
    \Tile_X5Y12_EE4BEG[11] ,
    \Tile_X5Y12_EE4BEG[10] ,
    \Tile_X5Y12_EE4BEG[9] ,
    \Tile_X5Y12_EE4BEG[8] ,
    \Tile_X5Y12_EE4BEG[7] ,
    \Tile_X5Y12_EE4BEG[6] ,
    \Tile_X5Y12_EE4BEG[5] ,
    \Tile_X5Y12_EE4BEG[4] ,
    \Tile_X5Y12_EE4BEG[3] ,
    \Tile_X5Y12_EE4BEG[2] ,
    \Tile_X5Y12_EE4BEG[1] ,
    \Tile_X5Y12_EE4BEG[0] }),
    .FrameData({\Tile_X5Y12_FrameData_O[31] ,
    \Tile_X5Y12_FrameData_O[30] ,
    \Tile_X5Y12_FrameData_O[29] ,
    \Tile_X5Y12_FrameData_O[28] ,
    \Tile_X5Y12_FrameData_O[27] ,
    \Tile_X5Y12_FrameData_O[26] ,
    \Tile_X5Y12_FrameData_O[25] ,
    \Tile_X5Y12_FrameData_O[24] ,
    \Tile_X5Y12_FrameData_O[23] ,
    \Tile_X5Y12_FrameData_O[22] ,
    \Tile_X5Y12_FrameData_O[21] ,
    \Tile_X5Y12_FrameData_O[20] ,
    \Tile_X5Y12_FrameData_O[19] ,
    \Tile_X5Y12_FrameData_O[18] ,
    \Tile_X5Y12_FrameData_O[17] ,
    \Tile_X5Y12_FrameData_O[16] ,
    \Tile_X5Y12_FrameData_O[15] ,
    \Tile_X5Y12_FrameData_O[14] ,
    \Tile_X5Y12_FrameData_O[13] ,
    \Tile_X5Y12_FrameData_O[12] ,
    \Tile_X5Y12_FrameData_O[11] ,
    \Tile_X5Y12_FrameData_O[10] ,
    \Tile_X5Y12_FrameData_O[9] ,
    \Tile_X5Y12_FrameData_O[8] ,
    \Tile_X5Y12_FrameData_O[7] ,
    \Tile_X5Y12_FrameData_O[6] ,
    \Tile_X5Y12_FrameData_O[5] ,
    \Tile_X5Y12_FrameData_O[4] ,
    \Tile_X5Y12_FrameData_O[3] ,
    \Tile_X5Y12_FrameData_O[2] ,
    \Tile_X5Y12_FrameData_O[1] ,
    \Tile_X5Y12_FrameData_O[0] }),
    .FrameData_O({\Tile_X6Y12_FrameData_O[31] ,
    \Tile_X6Y12_FrameData_O[30] ,
    \Tile_X6Y12_FrameData_O[29] ,
    \Tile_X6Y12_FrameData_O[28] ,
    \Tile_X6Y12_FrameData_O[27] ,
    \Tile_X6Y12_FrameData_O[26] ,
    \Tile_X6Y12_FrameData_O[25] ,
    \Tile_X6Y12_FrameData_O[24] ,
    \Tile_X6Y12_FrameData_O[23] ,
    \Tile_X6Y12_FrameData_O[22] ,
    \Tile_X6Y12_FrameData_O[21] ,
    \Tile_X6Y12_FrameData_O[20] ,
    \Tile_X6Y12_FrameData_O[19] ,
    \Tile_X6Y12_FrameData_O[18] ,
    \Tile_X6Y12_FrameData_O[17] ,
    \Tile_X6Y12_FrameData_O[16] ,
    \Tile_X6Y12_FrameData_O[15] ,
    \Tile_X6Y12_FrameData_O[14] ,
    \Tile_X6Y12_FrameData_O[13] ,
    \Tile_X6Y12_FrameData_O[12] ,
    \Tile_X6Y12_FrameData_O[11] ,
    \Tile_X6Y12_FrameData_O[10] ,
    \Tile_X6Y12_FrameData_O[9] ,
    \Tile_X6Y12_FrameData_O[8] ,
    \Tile_X6Y12_FrameData_O[7] ,
    \Tile_X6Y12_FrameData_O[6] ,
    \Tile_X6Y12_FrameData_O[5] ,
    \Tile_X6Y12_FrameData_O[4] ,
    \Tile_X6Y12_FrameData_O[3] ,
    \Tile_X6Y12_FrameData_O[2] ,
    \Tile_X6Y12_FrameData_O[1] ,
    \Tile_X6Y12_FrameData_O[0] }),
    .FrameStrobe({\Tile_X6Y13_FrameStrobe_O[19] ,
    \Tile_X6Y13_FrameStrobe_O[18] ,
    \Tile_X6Y13_FrameStrobe_O[17] ,
    \Tile_X6Y13_FrameStrobe_O[16] ,
    \Tile_X6Y13_FrameStrobe_O[15] ,
    \Tile_X6Y13_FrameStrobe_O[14] ,
    \Tile_X6Y13_FrameStrobe_O[13] ,
    \Tile_X6Y13_FrameStrobe_O[12] ,
    \Tile_X6Y13_FrameStrobe_O[11] ,
    \Tile_X6Y13_FrameStrobe_O[10] ,
    \Tile_X6Y13_FrameStrobe_O[9] ,
    \Tile_X6Y13_FrameStrobe_O[8] ,
    \Tile_X6Y13_FrameStrobe_O[7] ,
    \Tile_X6Y13_FrameStrobe_O[6] ,
    \Tile_X6Y13_FrameStrobe_O[5] ,
    \Tile_X6Y13_FrameStrobe_O[4] ,
    \Tile_X6Y13_FrameStrobe_O[3] ,
    \Tile_X6Y13_FrameStrobe_O[2] ,
    \Tile_X6Y13_FrameStrobe_O[1] ,
    \Tile_X6Y13_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X6Y12_FrameStrobe_O[19] ,
    \Tile_X6Y12_FrameStrobe_O[18] ,
    \Tile_X6Y12_FrameStrobe_O[17] ,
    \Tile_X6Y12_FrameStrobe_O[16] ,
    \Tile_X6Y12_FrameStrobe_O[15] ,
    \Tile_X6Y12_FrameStrobe_O[14] ,
    \Tile_X6Y12_FrameStrobe_O[13] ,
    \Tile_X6Y12_FrameStrobe_O[12] ,
    \Tile_X6Y12_FrameStrobe_O[11] ,
    \Tile_X6Y12_FrameStrobe_O[10] ,
    \Tile_X6Y12_FrameStrobe_O[9] ,
    \Tile_X6Y12_FrameStrobe_O[8] ,
    \Tile_X6Y12_FrameStrobe_O[7] ,
    \Tile_X6Y12_FrameStrobe_O[6] ,
    \Tile_X6Y12_FrameStrobe_O[5] ,
    \Tile_X6Y12_FrameStrobe_O[4] ,
    \Tile_X6Y12_FrameStrobe_O[3] ,
    \Tile_X6Y12_FrameStrobe_O[2] ,
    \Tile_X6Y12_FrameStrobe_O[1] ,
    \Tile_X6Y12_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X6Y12_N1BEG[3] ,
    \Tile_X6Y12_N1BEG[2] ,
    \Tile_X6Y12_N1BEG[1] ,
    \Tile_X6Y12_N1BEG[0] }),
    .N1END({\Tile_X6Y13_N1BEG[3] ,
    \Tile_X6Y13_N1BEG[2] ,
    \Tile_X6Y13_N1BEG[1] ,
    \Tile_X6Y13_N1BEG[0] }),
    .N2BEG({\Tile_X6Y12_N2BEG[7] ,
    \Tile_X6Y12_N2BEG[6] ,
    \Tile_X6Y12_N2BEG[5] ,
    \Tile_X6Y12_N2BEG[4] ,
    \Tile_X6Y12_N2BEG[3] ,
    \Tile_X6Y12_N2BEG[2] ,
    \Tile_X6Y12_N2BEG[1] ,
    \Tile_X6Y12_N2BEG[0] }),
    .N2BEGb({\Tile_X6Y12_N2BEGb[7] ,
    \Tile_X6Y12_N2BEGb[6] ,
    \Tile_X6Y12_N2BEGb[5] ,
    \Tile_X6Y12_N2BEGb[4] ,
    \Tile_X6Y12_N2BEGb[3] ,
    \Tile_X6Y12_N2BEGb[2] ,
    \Tile_X6Y12_N2BEGb[1] ,
    \Tile_X6Y12_N2BEGb[0] }),
    .N2END({\Tile_X6Y13_N2BEGb[7] ,
    \Tile_X6Y13_N2BEGb[6] ,
    \Tile_X6Y13_N2BEGb[5] ,
    \Tile_X6Y13_N2BEGb[4] ,
    \Tile_X6Y13_N2BEGb[3] ,
    \Tile_X6Y13_N2BEGb[2] ,
    \Tile_X6Y13_N2BEGb[1] ,
    \Tile_X6Y13_N2BEGb[0] }),
    .N2MID({\Tile_X6Y13_N2BEG[7] ,
    \Tile_X6Y13_N2BEG[6] ,
    \Tile_X6Y13_N2BEG[5] ,
    \Tile_X6Y13_N2BEG[4] ,
    \Tile_X6Y13_N2BEG[3] ,
    \Tile_X6Y13_N2BEG[2] ,
    \Tile_X6Y13_N2BEG[1] ,
    \Tile_X6Y13_N2BEG[0] }),
    .N4BEG({\Tile_X6Y12_N4BEG[15] ,
    \Tile_X6Y12_N4BEG[14] ,
    \Tile_X6Y12_N4BEG[13] ,
    \Tile_X6Y12_N4BEG[12] ,
    \Tile_X6Y12_N4BEG[11] ,
    \Tile_X6Y12_N4BEG[10] ,
    \Tile_X6Y12_N4BEG[9] ,
    \Tile_X6Y12_N4BEG[8] ,
    \Tile_X6Y12_N4BEG[7] ,
    \Tile_X6Y12_N4BEG[6] ,
    \Tile_X6Y12_N4BEG[5] ,
    \Tile_X6Y12_N4BEG[4] ,
    \Tile_X6Y12_N4BEG[3] ,
    \Tile_X6Y12_N4BEG[2] ,
    \Tile_X6Y12_N4BEG[1] ,
    \Tile_X6Y12_N4BEG[0] }),
    .N4END({\Tile_X6Y13_N4BEG[15] ,
    \Tile_X6Y13_N4BEG[14] ,
    \Tile_X6Y13_N4BEG[13] ,
    \Tile_X6Y13_N4BEG[12] ,
    \Tile_X6Y13_N4BEG[11] ,
    \Tile_X6Y13_N4BEG[10] ,
    \Tile_X6Y13_N4BEG[9] ,
    \Tile_X6Y13_N4BEG[8] ,
    \Tile_X6Y13_N4BEG[7] ,
    \Tile_X6Y13_N4BEG[6] ,
    \Tile_X6Y13_N4BEG[5] ,
    \Tile_X6Y13_N4BEG[4] ,
    \Tile_X6Y13_N4BEG[3] ,
    \Tile_X6Y13_N4BEG[2] ,
    \Tile_X6Y13_N4BEG[1] ,
    \Tile_X6Y13_N4BEG[0] }),
    .NN4BEG({\Tile_X6Y12_NN4BEG[15] ,
    \Tile_X6Y12_NN4BEG[14] ,
    \Tile_X6Y12_NN4BEG[13] ,
    \Tile_X6Y12_NN4BEG[12] ,
    \Tile_X6Y12_NN4BEG[11] ,
    \Tile_X6Y12_NN4BEG[10] ,
    \Tile_X6Y12_NN4BEG[9] ,
    \Tile_X6Y12_NN4BEG[8] ,
    \Tile_X6Y12_NN4BEG[7] ,
    \Tile_X6Y12_NN4BEG[6] ,
    \Tile_X6Y12_NN4BEG[5] ,
    \Tile_X6Y12_NN4BEG[4] ,
    \Tile_X6Y12_NN4BEG[3] ,
    \Tile_X6Y12_NN4BEG[2] ,
    \Tile_X6Y12_NN4BEG[1] ,
    \Tile_X6Y12_NN4BEG[0] }),
    .NN4END({\Tile_X6Y13_NN4BEG[15] ,
    \Tile_X6Y13_NN4BEG[14] ,
    \Tile_X6Y13_NN4BEG[13] ,
    \Tile_X6Y13_NN4BEG[12] ,
    \Tile_X6Y13_NN4BEG[11] ,
    \Tile_X6Y13_NN4BEG[10] ,
    \Tile_X6Y13_NN4BEG[9] ,
    \Tile_X6Y13_NN4BEG[8] ,
    \Tile_X6Y13_NN4BEG[7] ,
    \Tile_X6Y13_NN4BEG[6] ,
    \Tile_X6Y13_NN4BEG[5] ,
    \Tile_X6Y13_NN4BEG[4] ,
    \Tile_X6Y13_NN4BEG[3] ,
    \Tile_X6Y13_NN4BEG[2] ,
    \Tile_X6Y13_NN4BEG[1] ,
    \Tile_X6Y13_NN4BEG[0] }),
    .S1BEG({\Tile_X6Y12_S1BEG[3] ,
    \Tile_X6Y12_S1BEG[2] ,
    \Tile_X6Y12_S1BEG[1] ,
    \Tile_X6Y12_S1BEG[0] }),
    .S1END({\Tile_X6Y11_S1BEG[3] ,
    \Tile_X6Y11_S1BEG[2] ,
    \Tile_X6Y11_S1BEG[1] ,
    \Tile_X6Y11_S1BEG[0] }),
    .S2BEG({\Tile_X6Y12_S2BEG[7] ,
    \Tile_X6Y12_S2BEG[6] ,
    \Tile_X6Y12_S2BEG[5] ,
    \Tile_X6Y12_S2BEG[4] ,
    \Tile_X6Y12_S2BEG[3] ,
    \Tile_X6Y12_S2BEG[2] ,
    \Tile_X6Y12_S2BEG[1] ,
    \Tile_X6Y12_S2BEG[0] }),
    .S2BEGb({\Tile_X6Y12_S2BEGb[7] ,
    \Tile_X6Y12_S2BEGb[6] ,
    \Tile_X6Y12_S2BEGb[5] ,
    \Tile_X6Y12_S2BEGb[4] ,
    \Tile_X6Y12_S2BEGb[3] ,
    \Tile_X6Y12_S2BEGb[2] ,
    \Tile_X6Y12_S2BEGb[1] ,
    \Tile_X6Y12_S2BEGb[0] }),
    .S2END({\Tile_X6Y11_S2BEGb[7] ,
    \Tile_X6Y11_S2BEGb[6] ,
    \Tile_X6Y11_S2BEGb[5] ,
    \Tile_X6Y11_S2BEGb[4] ,
    \Tile_X6Y11_S2BEGb[3] ,
    \Tile_X6Y11_S2BEGb[2] ,
    \Tile_X6Y11_S2BEGb[1] ,
    \Tile_X6Y11_S2BEGb[0] }),
    .S2MID({\Tile_X6Y11_S2BEG[7] ,
    \Tile_X6Y11_S2BEG[6] ,
    \Tile_X6Y11_S2BEG[5] ,
    \Tile_X6Y11_S2BEG[4] ,
    \Tile_X6Y11_S2BEG[3] ,
    \Tile_X6Y11_S2BEG[2] ,
    \Tile_X6Y11_S2BEG[1] ,
    \Tile_X6Y11_S2BEG[0] }),
    .S4BEG({\Tile_X6Y12_S4BEG[15] ,
    \Tile_X6Y12_S4BEG[14] ,
    \Tile_X6Y12_S4BEG[13] ,
    \Tile_X6Y12_S4BEG[12] ,
    \Tile_X6Y12_S4BEG[11] ,
    \Tile_X6Y12_S4BEG[10] ,
    \Tile_X6Y12_S4BEG[9] ,
    \Tile_X6Y12_S4BEG[8] ,
    \Tile_X6Y12_S4BEG[7] ,
    \Tile_X6Y12_S4BEG[6] ,
    \Tile_X6Y12_S4BEG[5] ,
    \Tile_X6Y12_S4BEG[4] ,
    \Tile_X6Y12_S4BEG[3] ,
    \Tile_X6Y12_S4BEG[2] ,
    \Tile_X6Y12_S4BEG[1] ,
    \Tile_X6Y12_S4BEG[0] }),
    .S4END({\Tile_X6Y11_S4BEG[15] ,
    \Tile_X6Y11_S4BEG[14] ,
    \Tile_X6Y11_S4BEG[13] ,
    \Tile_X6Y11_S4BEG[12] ,
    \Tile_X6Y11_S4BEG[11] ,
    \Tile_X6Y11_S4BEG[10] ,
    \Tile_X6Y11_S4BEG[9] ,
    \Tile_X6Y11_S4BEG[8] ,
    \Tile_X6Y11_S4BEG[7] ,
    \Tile_X6Y11_S4BEG[6] ,
    \Tile_X6Y11_S4BEG[5] ,
    \Tile_X6Y11_S4BEG[4] ,
    \Tile_X6Y11_S4BEG[3] ,
    \Tile_X6Y11_S4BEG[2] ,
    \Tile_X6Y11_S4BEG[1] ,
    \Tile_X6Y11_S4BEG[0] }),
    .SS4BEG({\Tile_X6Y12_SS4BEG[15] ,
    \Tile_X6Y12_SS4BEG[14] ,
    \Tile_X6Y12_SS4BEG[13] ,
    \Tile_X6Y12_SS4BEG[12] ,
    \Tile_X6Y12_SS4BEG[11] ,
    \Tile_X6Y12_SS4BEG[10] ,
    \Tile_X6Y12_SS4BEG[9] ,
    \Tile_X6Y12_SS4BEG[8] ,
    \Tile_X6Y12_SS4BEG[7] ,
    \Tile_X6Y12_SS4BEG[6] ,
    \Tile_X6Y12_SS4BEG[5] ,
    \Tile_X6Y12_SS4BEG[4] ,
    \Tile_X6Y12_SS4BEG[3] ,
    \Tile_X6Y12_SS4BEG[2] ,
    \Tile_X6Y12_SS4BEG[1] ,
    \Tile_X6Y12_SS4BEG[0] }),
    .SS4END({\Tile_X6Y11_SS4BEG[15] ,
    \Tile_X6Y11_SS4BEG[14] ,
    \Tile_X6Y11_SS4BEG[13] ,
    \Tile_X6Y11_SS4BEG[12] ,
    \Tile_X6Y11_SS4BEG[11] ,
    \Tile_X6Y11_SS4BEG[10] ,
    \Tile_X6Y11_SS4BEG[9] ,
    \Tile_X6Y11_SS4BEG[8] ,
    \Tile_X6Y11_SS4BEG[7] ,
    \Tile_X6Y11_SS4BEG[6] ,
    \Tile_X6Y11_SS4BEG[5] ,
    \Tile_X6Y11_SS4BEG[4] ,
    \Tile_X6Y11_SS4BEG[3] ,
    \Tile_X6Y11_SS4BEG[2] ,
    \Tile_X6Y11_SS4BEG[1] ,
    \Tile_X6Y11_SS4BEG[0] }),
    .W1BEG({\Tile_X6Y12_W1BEG[3] ,
    \Tile_X6Y12_W1BEG[2] ,
    \Tile_X6Y12_W1BEG[1] ,
    \Tile_X6Y12_W1BEG[0] }),
    .W1END({\Tile_X7Y12_W1BEG[3] ,
    \Tile_X7Y12_W1BEG[2] ,
    \Tile_X7Y12_W1BEG[1] ,
    \Tile_X7Y12_W1BEG[0] }),
    .W2BEG({\Tile_X6Y12_W2BEG[7] ,
    \Tile_X6Y12_W2BEG[6] ,
    \Tile_X6Y12_W2BEG[5] ,
    \Tile_X6Y12_W2BEG[4] ,
    \Tile_X6Y12_W2BEG[3] ,
    \Tile_X6Y12_W2BEG[2] ,
    \Tile_X6Y12_W2BEG[1] ,
    \Tile_X6Y12_W2BEG[0] }),
    .W2BEGb({\Tile_X6Y12_W2BEGb[7] ,
    \Tile_X6Y12_W2BEGb[6] ,
    \Tile_X6Y12_W2BEGb[5] ,
    \Tile_X6Y12_W2BEGb[4] ,
    \Tile_X6Y12_W2BEGb[3] ,
    \Tile_X6Y12_W2BEGb[2] ,
    \Tile_X6Y12_W2BEGb[1] ,
    \Tile_X6Y12_W2BEGb[0] }),
    .W2END({\Tile_X7Y12_W2BEGb[7] ,
    \Tile_X7Y12_W2BEGb[6] ,
    \Tile_X7Y12_W2BEGb[5] ,
    \Tile_X7Y12_W2BEGb[4] ,
    \Tile_X7Y12_W2BEGb[3] ,
    \Tile_X7Y12_W2BEGb[2] ,
    \Tile_X7Y12_W2BEGb[1] ,
    \Tile_X7Y12_W2BEGb[0] }),
    .W2MID({\Tile_X7Y12_W2BEG[7] ,
    \Tile_X7Y12_W2BEG[6] ,
    \Tile_X7Y12_W2BEG[5] ,
    \Tile_X7Y12_W2BEG[4] ,
    \Tile_X7Y12_W2BEG[3] ,
    \Tile_X7Y12_W2BEG[2] ,
    \Tile_X7Y12_W2BEG[1] ,
    \Tile_X7Y12_W2BEG[0] }),
    .W6BEG({\Tile_X6Y12_W6BEG[11] ,
    \Tile_X6Y12_W6BEG[10] ,
    \Tile_X6Y12_W6BEG[9] ,
    \Tile_X6Y12_W6BEG[8] ,
    \Tile_X6Y12_W6BEG[7] ,
    \Tile_X6Y12_W6BEG[6] ,
    \Tile_X6Y12_W6BEG[5] ,
    \Tile_X6Y12_W6BEG[4] ,
    \Tile_X6Y12_W6BEG[3] ,
    \Tile_X6Y12_W6BEG[2] ,
    \Tile_X6Y12_W6BEG[1] ,
    \Tile_X6Y12_W6BEG[0] }),
    .W6END({\Tile_X7Y12_W6BEG[11] ,
    \Tile_X7Y12_W6BEG[10] ,
    \Tile_X7Y12_W6BEG[9] ,
    \Tile_X7Y12_W6BEG[8] ,
    \Tile_X7Y12_W6BEG[7] ,
    \Tile_X7Y12_W6BEG[6] ,
    \Tile_X7Y12_W6BEG[5] ,
    \Tile_X7Y12_W6BEG[4] ,
    \Tile_X7Y12_W6BEG[3] ,
    \Tile_X7Y12_W6BEG[2] ,
    \Tile_X7Y12_W6BEG[1] ,
    \Tile_X7Y12_W6BEG[0] }),
    .WW4BEG({\Tile_X6Y12_WW4BEG[15] ,
    \Tile_X6Y12_WW4BEG[14] ,
    \Tile_X6Y12_WW4BEG[13] ,
    \Tile_X6Y12_WW4BEG[12] ,
    \Tile_X6Y12_WW4BEG[11] ,
    \Tile_X6Y12_WW4BEG[10] ,
    \Tile_X6Y12_WW4BEG[9] ,
    \Tile_X6Y12_WW4BEG[8] ,
    \Tile_X6Y12_WW4BEG[7] ,
    \Tile_X6Y12_WW4BEG[6] ,
    \Tile_X6Y12_WW4BEG[5] ,
    \Tile_X6Y12_WW4BEG[4] ,
    \Tile_X6Y12_WW4BEG[3] ,
    \Tile_X6Y12_WW4BEG[2] ,
    \Tile_X6Y12_WW4BEG[1] ,
    \Tile_X6Y12_WW4BEG[0] }),
    .WW4END({\Tile_X7Y12_WW4BEG[15] ,
    \Tile_X7Y12_WW4BEG[14] ,
    \Tile_X7Y12_WW4BEG[13] ,
    \Tile_X7Y12_WW4BEG[12] ,
    \Tile_X7Y12_WW4BEG[11] ,
    \Tile_X7Y12_WW4BEG[10] ,
    \Tile_X7Y12_WW4BEG[9] ,
    \Tile_X7Y12_WW4BEG[8] ,
    \Tile_X7Y12_WW4BEG[7] ,
    \Tile_X7Y12_WW4BEG[6] ,
    \Tile_X7Y12_WW4BEG[5] ,
    \Tile_X7Y12_WW4BEG[4] ,
    \Tile_X7Y12_WW4BEG[3] ,
    \Tile_X7Y12_WW4BEG[2] ,
    \Tile_X7Y12_WW4BEG[1] ,
    \Tile_X7Y12_WW4BEG[0] }));
 LUT4AB Tile_X6Y13_LUT4AB (.Ci(Tile_X6Y14_Co),
    .Co(Tile_X6Y13_Co),
    .UserCLK(Tile_X6Y14_UserCLKo),
    .UserCLKo(Tile_X6Y13_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X6Y13_E1BEG[3] ,
    \Tile_X6Y13_E1BEG[2] ,
    \Tile_X6Y13_E1BEG[1] ,
    \Tile_X6Y13_E1BEG[0] }),
    .E1END({\Tile_X5Y13_E1BEG[3] ,
    \Tile_X5Y13_E1BEG[2] ,
    \Tile_X5Y13_E1BEG[1] ,
    \Tile_X5Y13_E1BEG[0] }),
    .E2BEG({\Tile_X6Y13_E2BEG[7] ,
    \Tile_X6Y13_E2BEG[6] ,
    \Tile_X6Y13_E2BEG[5] ,
    \Tile_X6Y13_E2BEG[4] ,
    \Tile_X6Y13_E2BEG[3] ,
    \Tile_X6Y13_E2BEG[2] ,
    \Tile_X6Y13_E2BEG[1] ,
    \Tile_X6Y13_E2BEG[0] }),
    .E2BEGb({\Tile_X6Y13_E2BEGb[7] ,
    \Tile_X6Y13_E2BEGb[6] ,
    \Tile_X6Y13_E2BEGb[5] ,
    \Tile_X6Y13_E2BEGb[4] ,
    \Tile_X6Y13_E2BEGb[3] ,
    \Tile_X6Y13_E2BEGb[2] ,
    \Tile_X6Y13_E2BEGb[1] ,
    \Tile_X6Y13_E2BEGb[0] }),
    .E2END({\Tile_X5Y13_E2BEGb[7] ,
    \Tile_X5Y13_E2BEGb[6] ,
    \Tile_X5Y13_E2BEGb[5] ,
    \Tile_X5Y13_E2BEGb[4] ,
    \Tile_X5Y13_E2BEGb[3] ,
    \Tile_X5Y13_E2BEGb[2] ,
    \Tile_X5Y13_E2BEGb[1] ,
    \Tile_X5Y13_E2BEGb[0] }),
    .E2MID({\Tile_X5Y13_E2BEG[7] ,
    \Tile_X5Y13_E2BEG[6] ,
    \Tile_X5Y13_E2BEG[5] ,
    \Tile_X5Y13_E2BEG[4] ,
    \Tile_X5Y13_E2BEG[3] ,
    \Tile_X5Y13_E2BEG[2] ,
    \Tile_X5Y13_E2BEG[1] ,
    \Tile_X5Y13_E2BEG[0] }),
    .E6BEG({\Tile_X6Y13_E6BEG[11] ,
    \Tile_X6Y13_E6BEG[10] ,
    \Tile_X6Y13_E6BEG[9] ,
    \Tile_X6Y13_E6BEG[8] ,
    \Tile_X6Y13_E6BEG[7] ,
    \Tile_X6Y13_E6BEG[6] ,
    \Tile_X6Y13_E6BEG[5] ,
    \Tile_X6Y13_E6BEG[4] ,
    \Tile_X6Y13_E6BEG[3] ,
    \Tile_X6Y13_E6BEG[2] ,
    \Tile_X6Y13_E6BEG[1] ,
    \Tile_X6Y13_E6BEG[0] }),
    .E6END({\Tile_X5Y13_E6BEG[11] ,
    \Tile_X5Y13_E6BEG[10] ,
    \Tile_X5Y13_E6BEG[9] ,
    \Tile_X5Y13_E6BEG[8] ,
    \Tile_X5Y13_E6BEG[7] ,
    \Tile_X5Y13_E6BEG[6] ,
    \Tile_X5Y13_E6BEG[5] ,
    \Tile_X5Y13_E6BEG[4] ,
    \Tile_X5Y13_E6BEG[3] ,
    \Tile_X5Y13_E6BEG[2] ,
    \Tile_X5Y13_E6BEG[1] ,
    \Tile_X5Y13_E6BEG[0] }),
    .EE4BEG({\Tile_X6Y13_EE4BEG[15] ,
    \Tile_X6Y13_EE4BEG[14] ,
    \Tile_X6Y13_EE4BEG[13] ,
    \Tile_X6Y13_EE4BEG[12] ,
    \Tile_X6Y13_EE4BEG[11] ,
    \Tile_X6Y13_EE4BEG[10] ,
    \Tile_X6Y13_EE4BEG[9] ,
    \Tile_X6Y13_EE4BEG[8] ,
    \Tile_X6Y13_EE4BEG[7] ,
    \Tile_X6Y13_EE4BEG[6] ,
    \Tile_X6Y13_EE4BEG[5] ,
    \Tile_X6Y13_EE4BEG[4] ,
    \Tile_X6Y13_EE4BEG[3] ,
    \Tile_X6Y13_EE4BEG[2] ,
    \Tile_X6Y13_EE4BEG[1] ,
    \Tile_X6Y13_EE4BEG[0] }),
    .EE4END({\Tile_X5Y13_EE4BEG[15] ,
    \Tile_X5Y13_EE4BEG[14] ,
    \Tile_X5Y13_EE4BEG[13] ,
    \Tile_X5Y13_EE4BEG[12] ,
    \Tile_X5Y13_EE4BEG[11] ,
    \Tile_X5Y13_EE4BEG[10] ,
    \Tile_X5Y13_EE4BEG[9] ,
    \Tile_X5Y13_EE4BEG[8] ,
    \Tile_X5Y13_EE4BEG[7] ,
    \Tile_X5Y13_EE4BEG[6] ,
    \Tile_X5Y13_EE4BEG[5] ,
    \Tile_X5Y13_EE4BEG[4] ,
    \Tile_X5Y13_EE4BEG[3] ,
    \Tile_X5Y13_EE4BEG[2] ,
    \Tile_X5Y13_EE4BEG[1] ,
    \Tile_X5Y13_EE4BEG[0] }),
    .FrameData({\Tile_X5Y13_FrameData_O[31] ,
    \Tile_X5Y13_FrameData_O[30] ,
    \Tile_X5Y13_FrameData_O[29] ,
    \Tile_X5Y13_FrameData_O[28] ,
    \Tile_X5Y13_FrameData_O[27] ,
    \Tile_X5Y13_FrameData_O[26] ,
    \Tile_X5Y13_FrameData_O[25] ,
    \Tile_X5Y13_FrameData_O[24] ,
    \Tile_X5Y13_FrameData_O[23] ,
    \Tile_X5Y13_FrameData_O[22] ,
    \Tile_X5Y13_FrameData_O[21] ,
    \Tile_X5Y13_FrameData_O[20] ,
    \Tile_X5Y13_FrameData_O[19] ,
    \Tile_X5Y13_FrameData_O[18] ,
    \Tile_X5Y13_FrameData_O[17] ,
    \Tile_X5Y13_FrameData_O[16] ,
    \Tile_X5Y13_FrameData_O[15] ,
    \Tile_X5Y13_FrameData_O[14] ,
    \Tile_X5Y13_FrameData_O[13] ,
    \Tile_X5Y13_FrameData_O[12] ,
    \Tile_X5Y13_FrameData_O[11] ,
    \Tile_X5Y13_FrameData_O[10] ,
    \Tile_X5Y13_FrameData_O[9] ,
    \Tile_X5Y13_FrameData_O[8] ,
    \Tile_X5Y13_FrameData_O[7] ,
    \Tile_X5Y13_FrameData_O[6] ,
    \Tile_X5Y13_FrameData_O[5] ,
    \Tile_X5Y13_FrameData_O[4] ,
    \Tile_X5Y13_FrameData_O[3] ,
    \Tile_X5Y13_FrameData_O[2] ,
    \Tile_X5Y13_FrameData_O[1] ,
    \Tile_X5Y13_FrameData_O[0] }),
    .FrameData_O({\Tile_X6Y13_FrameData_O[31] ,
    \Tile_X6Y13_FrameData_O[30] ,
    \Tile_X6Y13_FrameData_O[29] ,
    \Tile_X6Y13_FrameData_O[28] ,
    \Tile_X6Y13_FrameData_O[27] ,
    \Tile_X6Y13_FrameData_O[26] ,
    \Tile_X6Y13_FrameData_O[25] ,
    \Tile_X6Y13_FrameData_O[24] ,
    \Tile_X6Y13_FrameData_O[23] ,
    \Tile_X6Y13_FrameData_O[22] ,
    \Tile_X6Y13_FrameData_O[21] ,
    \Tile_X6Y13_FrameData_O[20] ,
    \Tile_X6Y13_FrameData_O[19] ,
    \Tile_X6Y13_FrameData_O[18] ,
    \Tile_X6Y13_FrameData_O[17] ,
    \Tile_X6Y13_FrameData_O[16] ,
    \Tile_X6Y13_FrameData_O[15] ,
    \Tile_X6Y13_FrameData_O[14] ,
    \Tile_X6Y13_FrameData_O[13] ,
    \Tile_X6Y13_FrameData_O[12] ,
    \Tile_X6Y13_FrameData_O[11] ,
    \Tile_X6Y13_FrameData_O[10] ,
    \Tile_X6Y13_FrameData_O[9] ,
    \Tile_X6Y13_FrameData_O[8] ,
    \Tile_X6Y13_FrameData_O[7] ,
    \Tile_X6Y13_FrameData_O[6] ,
    \Tile_X6Y13_FrameData_O[5] ,
    \Tile_X6Y13_FrameData_O[4] ,
    \Tile_X6Y13_FrameData_O[3] ,
    \Tile_X6Y13_FrameData_O[2] ,
    \Tile_X6Y13_FrameData_O[1] ,
    \Tile_X6Y13_FrameData_O[0] }),
    .FrameStrobe({\Tile_X6Y14_FrameStrobe_O[19] ,
    \Tile_X6Y14_FrameStrobe_O[18] ,
    \Tile_X6Y14_FrameStrobe_O[17] ,
    \Tile_X6Y14_FrameStrobe_O[16] ,
    \Tile_X6Y14_FrameStrobe_O[15] ,
    \Tile_X6Y14_FrameStrobe_O[14] ,
    \Tile_X6Y14_FrameStrobe_O[13] ,
    \Tile_X6Y14_FrameStrobe_O[12] ,
    \Tile_X6Y14_FrameStrobe_O[11] ,
    \Tile_X6Y14_FrameStrobe_O[10] ,
    \Tile_X6Y14_FrameStrobe_O[9] ,
    \Tile_X6Y14_FrameStrobe_O[8] ,
    \Tile_X6Y14_FrameStrobe_O[7] ,
    \Tile_X6Y14_FrameStrobe_O[6] ,
    \Tile_X6Y14_FrameStrobe_O[5] ,
    \Tile_X6Y14_FrameStrobe_O[4] ,
    \Tile_X6Y14_FrameStrobe_O[3] ,
    \Tile_X6Y14_FrameStrobe_O[2] ,
    \Tile_X6Y14_FrameStrobe_O[1] ,
    \Tile_X6Y14_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X6Y13_FrameStrobe_O[19] ,
    \Tile_X6Y13_FrameStrobe_O[18] ,
    \Tile_X6Y13_FrameStrobe_O[17] ,
    \Tile_X6Y13_FrameStrobe_O[16] ,
    \Tile_X6Y13_FrameStrobe_O[15] ,
    \Tile_X6Y13_FrameStrobe_O[14] ,
    \Tile_X6Y13_FrameStrobe_O[13] ,
    \Tile_X6Y13_FrameStrobe_O[12] ,
    \Tile_X6Y13_FrameStrobe_O[11] ,
    \Tile_X6Y13_FrameStrobe_O[10] ,
    \Tile_X6Y13_FrameStrobe_O[9] ,
    \Tile_X6Y13_FrameStrobe_O[8] ,
    \Tile_X6Y13_FrameStrobe_O[7] ,
    \Tile_X6Y13_FrameStrobe_O[6] ,
    \Tile_X6Y13_FrameStrobe_O[5] ,
    \Tile_X6Y13_FrameStrobe_O[4] ,
    \Tile_X6Y13_FrameStrobe_O[3] ,
    \Tile_X6Y13_FrameStrobe_O[2] ,
    \Tile_X6Y13_FrameStrobe_O[1] ,
    \Tile_X6Y13_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X6Y13_N1BEG[3] ,
    \Tile_X6Y13_N1BEG[2] ,
    \Tile_X6Y13_N1BEG[1] ,
    \Tile_X6Y13_N1BEG[0] }),
    .N1END({\Tile_X6Y14_N1BEG[3] ,
    \Tile_X6Y14_N1BEG[2] ,
    \Tile_X6Y14_N1BEG[1] ,
    \Tile_X6Y14_N1BEG[0] }),
    .N2BEG({\Tile_X6Y13_N2BEG[7] ,
    \Tile_X6Y13_N2BEG[6] ,
    \Tile_X6Y13_N2BEG[5] ,
    \Tile_X6Y13_N2BEG[4] ,
    \Tile_X6Y13_N2BEG[3] ,
    \Tile_X6Y13_N2BEG[2] ,
    \Tile_X6Y13_N2BEG[1] ,
    \Tile_X6Y13_N2BEG[0] }),
    .N2BEGb({\Tile_X6Y13_N2BEGb[7] ,
    \Tile_X6Y13_N2BEGb[6] ,
    \Tile_X6Y13_N2BEGb[5] ,
    \Tile_X6Y13_N2BEGb[4] ,
    \Tile_X6Y13_N2BEGb[3] ,
    \Tile_X6Y13_N2BEGb[2] ,
    \Tile_X6Y13_N2BEGb[1] ,
    \Tile_X6Y13_N2BEGb[0] }),
    .N2END({\Tile_X6Y14_N2BEGb[7] ,
    \Tile_X6Y14_N2BEGb[6] ,
    \Tile_X6Y14_N2BEGb[5] ,
    \Tile_X6Y14_N2BEGb[4] ,
    \Tile_X6Y14_N2BEGb[3] ,
    \Tile_X6Y14_N2BEGb[2] ,
    \Tile_X6Y14_N2BEGb[1] ,
    \Tile_X6Y14_N2BEGb[0] }),
    .N2MID({\Tile_X6Y14_N2BEG[7] ,
    \Tile_X6Y14_N2BEG[6] ,
    \Tile_X6Y14_N2BEG[5] ,
    \Tile_X6Y14_N2BEG[4] ,
    \Tile_X6Y14_N2BEG[3] ,
    \Tile_X6Y14_N2BEG[2] ,
    \Tile_X6Y14_N2BEG[1] ,
    \Tile_X6Y14_N2BEG[0] }),
    .N4BEG({\Tile_X6Y13_N4BEG[15] ,
    \Tile_X6Y13_N4BEG[14] ,
    \Tile_X6Y13_N4BEG[13] ,
    \Tile_X6Y13_N4BEG[12] ,
    \Tile_X6Y13_N4BEG[11] ,
    \Tile_X6Y13_N4BEG[10] ,
    \Tile_X6Y13_N4BEG[9] ,
    \Tile_X6Y13_N4BEG[8] ,
    \Tile_X6Y13_N4BEG[7] ,
    \Tile_X6Y13_N4BEG[6] ,
    \Tile_X6Y13_N4BEG[5] ,
    \Tile_X6Y13_N4BEG[4] ,
    \Tile_X6Y13_N4BEG[3] ,
    \Tile_X6Y13_N4BEG[2] ,
    \Tile_X6Y13_N4BEG[1] ,
    \Tile_X6Y13_N4BEG[0] }),
    .N4END({\Tile_X6Y14_N4BEG[15] ,
    \Tile_X6Y14_N4BEG[14] ,
    \Tile_X6Y14_N4BEG[13] ,
    \Tile_X6Y14_N4BEG[12] ,
    \Tile_X6Y14_N4BEG[11] ,
    \Tile_X6Y14_N4BEG[10] ,
    \Tile_X6Y14_N4BEG[9] ,
    \Tile_X6Y14_N4BEG[8] ,
    \Tile_X6Y14_N4BEG[7] ,
    \Tile_X6Y14_N4BEG[6] ,
    \Tile_X6Y14_N4BEG[5] ,
    \Tile_X6Y14_N4BEG[4] ,
    \Tile_X6Y14_N4BEG[3] ,
    \Tile_X6Y14_N4BEG[2] ,
    \Tile_X6Y14_N4BEG[1] ,
    \Tile_X6Y14_N4BEG[0] }),
    .NN4BEG({\Tile_X6Y13_NN4BEG[15] ,
    \Tile_X6Y13_NN4BEG[14] ,
    \Tile_X6Y13_NN4BEG[13] ,
    \Tile_X6Y13_NN4BEG[12] ,
    \Tile_X6Y13_NN4BEG[11] ,
    \Tile_X6Y13_NN4BEG[10] ,
    \Tile_X6Y13_NN4BEG[9] ,
    \Tile_X6Y13_NN4BEG[8] ,
    \Tile_X6Y13_NN4BEG[7] ,
    \Tile_X6Y13_NN4BEG[6] ,
    \Tile_X6Y13_NN4BEG[5] ,
    \Tile_X6Y13_NN4BEG[4] ,
    \Tile_X6Y13_NN4BEG[3] ,
    \Tile_X6Y13_NN4BEG[2] ,
    \Tile_X6Y13_NN4BEG[1] ,
    \Tile_X6Y13_NN4BEG[0] }),
    .NN4END({\Tile_X6Y14_NN4BEG[15] ,
    \Tile_X6Y14_NN4BEG[14] ,
    \Tile_X6Y14_NN4BEG[13] ,
    \Tile_X6Y14_NN4BEG[12] ,
    \Tile_X6Y14_NN4BEG[11] ,
    \Tile_X6Y14_NN4BEG[10] ,
    \Tile_X6Y14_NN4BEG[9] ,
    \Tile_X6Y14_NN4BEG[8] ,
    \Tile_X6Y14_NN4BEG[7] ,
    \Tile_X6Y14_NN4BEG[6] ,
    \Tile_X6Y14_NN4BEG[5] ,
    \Tile_X6Y14_NN4BEG[4] ,
    \Tile_X6Y14_NN4BEG[3] ,
    \Tile_X6Y14_NN4BEG[2] ,
    \Tile_X6Y14_NN4BEG[1] ,
    \Tile_X6Y14_NN4BEG[0] }),
    .S1BEG({\Tile_X6Y13_S1BEG[3] ,
    \Tile_X6Y13_S1BEG[2] ,
    \Tile_X6Y13_S1BEG[1] ,
    \Tile_X6Y13_S1BEG[0] }),
    .S1END({\Tile_X6Y12_S1BEG[3] ,
    \Tile_X6Y12_S1BEG[2] ,
    \Tile_X6Y12_S1BEG[1] ,
    \Tile_X6Y12_S1BEG[0] }),
    .S2BEG({\Tile_X6Y13_S2BEG[7] ,
    \Tile_X6Y13_S2BEG[6] ,
    \Tile_X6Y13_S2BEG[5] ,
    \Tile_X6Y13_S2BEG[4] ,
    \Tile_X6Y13_S2BEG[3] ,
    \Tile_X6Y13_S2BEG[2] ,
    \Tile_X6Y13_S2BEG[1] ,
    \Tile_X6Y13_S2BEG[0] }),
    .S2BEGb({\Tile_X6Y13_S2BEGb[7] ,
    \Tile_X6Y13_S2BEGb[6] ,
    \Tile_X6Y13_S2BEGb[5] ,
    \Tile_X6Y13_S2BEGb[4] ,
    \Tile_X6Y13_S2BEGb[3] ,
    \Tile_X6Y13_S2BEGb[2] ,
    \Tile_X6Y13_S2BEGb[1] ,
    \Tile_X6Y13_S2BEGb[0] }),
    .S2END({\Tile_X6Y12_S2BEGb[7] ,
    \Tile_X6Y12_S2BEGb[6] ,
    \Tile_X6Y12_S2BEGb[5] ,
    \Tile_X6Y12_S2BEGb[4] ,
    \Tile_X6Y12_S2BEGb[3] ,
    \Tile_X6Y12_S2BEGb[2] ,
    \Tile_X6Y12_S2BEGb[1] ,
    \Tile_X6Y12_S2BEGb[0] }),
    .S2MID({\Tile_X6Y12_S2BEG[7] ,
    \Tile_X6Y12_S2BEG[6] ,
    \Tile_X6Y12_S2BEG[5] ,
    \Tile_X6Y12_S2BEG[4] ,
    \Tile_X6Y12_S2BEG[3] ,
    \Tile_X6Y12_S2BEG[2] ,
    \Tile_X6Y12_S2BEG[1] ,
    \Tile_X6Y12_S2BEG[0] }),
    .S4BEG({\Tile_X6Y13_S4BEG[15] ,
    \Tile_X6Y13_S4BEG[14] ,
    \Tile_X6Y13_S4BEG[13] ,
    \Tile_X6Y13_S4BEG[12] ,
    \Tile_X6Y13_S4BEG[11] ,
    \Tile_X6Y13_S4BEG[10] ,
    \Tile_X6Y13_S4BEG[9] ,
    \Tile_X6Y13_S4BEG[8] ,
    \Tile_X6Y13_S4BEG[7] ,
    \Tile_X6Y13_S4BEG[6] ,
    \Tile_X6Y13_S4BEG[5] ,
    \Tile_X6Y13_S4BEG[4] ,
    \Tile_X6Y13_S4BEG[3] ,
    \Tile_X6Y13_S4BEG[2] ,
    \Tile_X6Y13_S4BEG[1] ,
    \Tile_X6Y13_S4BEG[0] }),
    .S4END({\Tile_X6Y12_S4BEG[15] ,
    \Tile_X6Y12_S4BEG[14] ,
    \Tile_X6Y12_S4BEG[13] ,
    \Tile_X6Y12_S4BEG[12] ,
    \Tile_X6Y12_S4BEG[11] ,
    \Tile_X6Y12_S4BEG[10] ,
    \Tile_X6Y12_S4BEG[9] ,
    \Tile_X6Y12_S4BEG[8] ,
    \Tile_X6Y12_S4BEG[7] ,
    \Tile_X6Y12_S4BEG[6] ,
    \Tile_X6Y12_S4BEG[5] ,
    \Tile_X6Y12_S4BEG[4] ,
    \Tile_X6Y12_S4BEG[3] ,
    \Tile_X6Y12_S4BEG[2] ,
    \Tile_X6Y12_S4BEG[1] ,
    \Tile_X6Y12_S4BEG[0] }),
    .SS4BEG({\Tile_X6Y13_SS4BEG[15] ,
    \Tile_X6Y13_SS4BEG[14] ,
    \Tile_X6Y13_SS4BEG[13] ,
    \Tile_X6Y13_SS4BEG[12] ,
    \Tile_X6Y13_SS4BEG[11] ,
    \Tile_X6Y13_SS4BEG[10] ,
    \Tile_X6Y13_SS4BEG[9] ,
    \Tile_X6Y13_SS4BEG[8] ,
    \Tile_X6Y13_SS4BEG[7] ,
    \Tile_X6Y13_SS4BEG[6] ,
    \Tile_X6Y13_SS4BEG[5] ,
    \Tile_X6Y13_SS4BEG[4] ,
    \Tile_X6Y13_SS4BEG[3] ,
    \Tile_X6Y13_SS4BEG[2] ,
    \Tile_X6Y13_SS4BEG[1] ,
    \Tile_X6Y13_SS4BEG[0] }),
    .SS4END({\Tile_X6Y12_SS4BEG[15] ,
    \Tile_X6Y12_SS4BEG[14] ,
    \Tile_X6Y12_SS4BEG[13] ,
    \Tile_X6Y12_SS4BEG[12] ,
    \Tile_X6Y12_SS4BEG[11] ,
    \Tile_X6Y12_SS4BEG[10] ,
    \Tile_X6Y12_SS4BEG[9] ,
    \Tile_X6Y12_SS4BEG[8] ,
    \Tile_X6Y12_SS4BEG[7] ,
    \Tile_X6Y12_SS4BEG[6] ,
    \Tile_X6Y12_SS4BEG[5] ,
    \Tile_X6Y12_SS4BEG[4] ,
    \Tile_X6Y12_SS4BEG[3] ,
    \Tile_X6Y12_SS4BEG[2] ,
    \Tile_X6Y12_SS4BEG[1] ,
    \Tile_X6Y12_SS4BEG[0] }),
    .W1BEG({\Tile_X6Y13_W1BEG[3] ,
    \Tile_X6Y13_W1BEG[2] ,
    \Tile_X6Y13_W1BEG[1] ,
    \Tile_X6Y13_W1BEG[0] }),
    .W1END({\Tile_X7Y13_W1BEG[3] ,
    \Tile_X7Y13_W1BEG[2] ,
    \Tile_X7Y13_W1BEG[1] ,
    \Tile_X7Y13_W1BEG[0] }),
    .W2BEG({\Tile_X6Y13_W2BEG[7] ,
    \Tile_X6Y13_W2BEG[6] ,
    \Tile_X6Y13_W2BEG[5] ,
    \Tile_X6Y13_W2BEG[4] ,
    \Tile_X6Y13_W2BEG[3] ,
    \Tile_X6Y13_W2BEG[2] ,
    \Tile_X6Y13_W2BEG[1] ,
    \Tile_X6Y13_W2BEG[0] }),
    .W2BEGb({\Tile_X6Y13_W2BEGb[7] ,
    \Tile_X6Y13_W2BEGb[6] ,
    \Tile_X6Y13_W2BEGb[5] ,
    \Tile_X6Y13_W2BEGb[4] ,
    \Tile_X6Y13_W2BEGb[3] ,
    \Tile_X6Y13_W2BEGb[2] ,
    \Tile_X6Y13_W2BEGb[1] ,
    \Tile_X6Y13_W2BEGb[0] }),
    .W2END({\Tile_X7Y13_W2BEGb[7] ,
    \Tile_X7Y13_W2BEGb[6] ,
    \Tile_X7Y13_W2BEGb[5] ,
    \Tile_X7Y13_W2BEGb[4] ,
    \Tile_X7Y13_W2BEGb[3] ,
    \Tile_X7Y13_W2BEGb[2] ,
    \Tile_X7Y13_W2BEGb[1] ,
    \Tile_X7Y13_W2BEGb[0] }),
    .W2MID({\Tile_X7Y13_W2BEG[7] ,
    \Tile_X7Y13_W2BEG[6] ,
    \Tile_X7Y13_W2BEG[5] ,
    \Tile_X7Y13_W2BEG[4] ,
    \Tile_X7Y13_W2BEG[3] ,
    \Tile_X7Y13_W2BEG[2] ,
    \Tile_X7Y13_W2BEG[1] ,
    \Tile_X7Y13_W2BEG[0] }),
    .W6BEG({\Tile_X6Y13_W6BEG[11] ,
    \Tile_X6Y13_W6BEG[10] ,
    \Tile_X6Y13_W6BEG[9] ,
    \Tile_X6Y13_W6BEG[8] ,
    \Tile_X6Y13_W6BEG[7] ,
    \Tile_X6Y13_W6BEG[6] ,
    \Tile_X6Y13_W6BEG[5] ,
    \Tile_X6Y13_W6BEG[4] ,
    \Tile_X6Y13_W6BEG[3] ,
    \Tile_X6Y13_W6BEG[2] ,
    \Tile_X6Y13_W6BEG[1] ,
    \Tile_X6Y13_W6BEG[0] }),
    .W6END({\Tile_X7Y13_W6BEG[11] ,
    \Tile_X7Y13_W6BEG[10] ,
    \Tile_X7Y13_W6BEG[9] ,
    \Tile_X7Y13_W6BEG[8] ,
    \Tile_X7Y13_W6BEG[7] ,
    \Tile_X7Y13_W6BEG[6] ,
    \Tile_X7Y13_W6BEG[5] ,
    \Tile_X7Y13_W6BEG[4] ,
    \Tile_X7Y13_W6BEG[3] ,
    \Tile_X7Y13_W6BEG[2] ,
    \Tile_X7Y13_W6BEG[1] ,
    \Tile_X7Y13_W6BEG[0] }),
    .WW4BEG({\Tile_X6Y13_WW4BEG[15] ,
    \Tile_X6Y13_WW4BEG[14] ,
    \Tile_X6Y13_WW4BEG[13] ,
    \Tile_X6Y13_WW4BEG[12] ,
    \Tile_X6Y13_WW4BEG[11] ,
    \Tile_X6Y13_WW4BEG[10] ,
    \Tile_X6Y13_WW4BEG[9] ,
    \Tile_X6Y13_WW4BEG[8] ,
    \Tile_X6Y13_WW4BEG[7] ,
    \Tile_X6Y13_WW4BEG[6] ,
    \Tile_X6Y13_WW4BEG[5] ,
    \Tile_X6Y13_WW4BEG[4] ,
    \Tile_X6Y13_WW4BEG[3] ,
    \Tile_X6Y13_WW4BEG[2] ,
    \Tile_X6Y13_WW4BEG[1] ,
    \Tile_X6Y13_WW4BEG[0] }),
    .WW4END({\Tile_X7Y13_WW4BEG[15] ,
    \Tile_X7Y13_WW4BEG[14] ,
    \Tile_X7Y13_WW4BEG[13] ,
    \Tile_X7Y13_WW4BEG[12] ,
    \Tile_X7Y13_WW4BEG[11] ,
    \Tile_X7Y13_WW4BEG[10] ,
    \Tile_X7Y13_WW4BEG[9] ,
    \Tile_X7Y13_WW4BEG[8] ,
    \Tile_X7Y13_WW4BEG[7] ,
    \Tile_X7Y13_WW4BEG[6] ,
    \Tile_X7Y13_WW4BEG[5] ,
    \Tile_X7Y13_WW4BEG[4] ,
    \Tile_X7Y13_WW4BEG[3] ,
    \Tile_X7Y13_WW4BEG[2] ,
    \Tile_X7Y13_WW4BEG[1] ,
    \Tile_X7Y13_WW4BEG[0] }));
 LUT4AB Tile_X6Y14_LUT4AB (.Ci(Tile_X6Y15_Co),
    .Co(Tile_X6Y14_Co),
    .UserCLK(Tile_X6Y15_UserCLKo),
    .UserCLKo(Tile_X6Y14_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X6Y14_E1BEG[3] ,
    \Tile_X6Y14_E1BEG[2] ,
    \Tile_X6Y14_E1BEG[1] ,
    \Tile_X6Y14_E1BEG[0] }),
    .E1END({\Tile_X5Y14_E1BEG[3] ,
    \Tile_X5Y14_E1BEG[2] ,
    \Tile_X5Y14_E1BEG[1] ,
    \Tile_X5Y14_E1BEG[0] }),
    .E2BEG({\Tile_X6Y14_E2BEG[7] ,
    \Tile_X6Y14_E2BEG[6] ,
    \Tile_X6Y14_E2BEG[5] ,
    \Tile_X6Y14_E2BEG[4] ,
    \Tile_X6Y14_E2BEG[3] ,
    \Tile_X6Y14_E2BEG[2] ,
    \Tile_X6Y14_E2BEG[1] ,
    \Tile_X6Y14_E2BEG[0] }),
    .E2BEGb({\Tile_X6Y14_E2BEGb[7] ,
    \Tile_X6Y14_E2BEGb[6] ,
    \Tile_X6Y14_E2BEGb[5] ,
    \Tile_X6Y14_E2BEGb[4] ,
    \Tile_X6Y14_E2BEGb[3] ,
    \Tile_X6Y14_E2BEGb[2] ,
    \Tile_X6Y14_E2BEGb[1] ,
    \Tile_X6Y14_E2BEGb[0] }),
    .E2END({\Tile_X5Y14_E2BEGb[7] ,
    \Tile_X5Y14_E2BEGb[6] ,
    \Tile_X5Y14_E2BEGb[5] ,
    \Tile_X5Y14_E2BEGb[4] ,
    \Tile_X5Y14_E2BEGb[3] ,
    \Tile_X5Y14_E2BEGb[2] ,
    \Tile_X5Y14_E2BEGb[1] ,
    \Tile_X5Y14_E2BEGb[0] }),
    .E2MID({\Tile_X5Y14_E2BEG[7] ,
    \Tile_X5Y14_E2BEG[6] ,
    \Tile_X5Y14_E2BEG[5] ,
    \Tile_X5Y14_E2BEG[4] ,
    \Tile_X5Y14_E2BEG[3] ,
    \Tile_X5Y14_E2BEG[2] ,
    \Tile_X5Y14_E2BEG[1] ,
    \Tile_X5Y14_E2BEG[0] }),
    .E6BEG({\Tile_X6Y14_E6BEG[11] ,
    \Tile_X6Y14_E6BEG[10] ,
    \Tile_X6Y14_E6BEG[9] ,
    \Tile_X6Y14_E6BEG[8] ,
    \Tile_X6Y14_E6BEG[7] ,
    \Tile_X6Y14_E6BEG[6] ,
    \Tile_X6Y14_E6BEG[5] ,
    \Tile_X6Y14_E6BEG[4] ,
    \Tile_X6Y14_E6BEG[3] ,
    \Tile_X6Y14_E6BEG[2] ,
    \Tile_X6Y14_E6BEG[1] ,
    \Tile_X6Y14_E6BEG[0] }),
    .E6END({\Tile_X5Y14_E6BEG[11] ,
    \Tile_X5Y14_E6BEG[10] ,
    \Tile_X5Y14_E6BEG[9] ,
    \Tile_X5Y14_E6BEG[8] ,
    \Tile_X5Y14_E6BEG[7] ,
    \Tile_X5Y14_E6BEG[6] ,
    \Tile_X5Y14_E6BEG[5] ,
    \Tile_X5Y14_E6BEG[4] ,
    \Tile_X5Y14_E6BEG[3] ,
    \Tile_X5Y14_E6BEG[2] ,
    \Tile_X5Y14_E6BEG[1] ,
    \Tile_X5Y14_E6BEG[0] }),
    .EE4BEG({\Tile_X6Y14_EE4BEG[15] ,
    \Tile_X6Y14_EE4BEG[14] ,
    \Tile_X6Y14_EE4BEG[13] ,
    \Tile_X6Y14_EE4BEG[12] ,
    \Tile_X6Y14_EE4BEG[11] ,
    \Tile_X6Y14_EE4BEG[10] ,
    \Tile_X6Y14_EE4BEG[9] ,
    \Tile_X6Y14_EE4BEG[8] ,
    \Tile_X6Y14_EE4BEG[7] ,
    \Tile_X6Y14_EE4BEG[6] ,
    \Tile_X6Y14_EE4BEG[5] ,
    \Tile_X6Y14_EE4BEG[4] ,
    \Tile_X6Y14_EE4BEG[3] ,
    \Tile_X6Y14_EE4BEG[2] ,
    \Tile_X6Y14_EE4BEG[1] ,
    \Tile_X6Y14_EE4BEG[0] }),
    .EE4END({\Tile_X5Y14_EE4BEG[15] ,
    \Tile_X5Y14_EE4BEG[14] ,
    \Tile_X5Y14_EE4BEG[13] ,
    \Tile_X5Y14_EE4BEG[12] ,
    \Tile_X5Y14_EE4BEG[11] ,
    \Tile_X5Y14_EE4BEG[10] ,
    \Tile_X5Y14_EE4BEG[9] ,
    \Tile_X5Y14_EE4BEG[8] ,
    \Tile_X5Y14_EE4BEG[7] ,
    \Tile_X5Y14_EE4BEG[6] ,
    \Tile_X5Y14_EE4BEG[5] ,
    \Tile_X5Y14_EE4BEG[4] ,
    \Tile_X5Y14_EE4BEG[3] ,
    \Tile_X5Y14_EE4BEG[2] ,
    \Tile_X5Y14_EE4BEG[1] ,
    \Tile_X5Y14_EE4BEG[0] }),
    .FrameData({\Tile_X5Y14_FrameData_O[31] ,
    \Tile_X5Y14_FrameData_O[30] ,
    \Tile_X5Y14_FrameData_O[29] ,
    \Tile_X5Y14_FrameData_O[28] ,
    \Tile_X5Y14_FrameData_O[27] ,
    \Tile_X5Y14_FrameData_O[26] ,
    \Tile_X5Y14_FrameData_O[25] ,
    \Tile_X5Y14_FrameData_O[24] ,
    \Tile_X5Y14_FrameData_O[23] ,
    \Tile_X5Y14_FrameData_O[22] ,
    \Tile_X5Y14_FrameData_O[21] ,
    \Tile_X5Y14_FrameData_O[20] ,
    \Tile_X5Y14_FrameData_O[19] ,
    \Tile_X5Y14_FrameData_O[18] ,
    \Tile_X5Y14_FrameData_O[17] ,
    \Tile_X5Y14_FrameData_O[16] ,
    \Tile_X5Y14_FrameData_O[15] ,
    \Tile_X5Y14_FrameData_O[14] ,
    \Tile_X5Y14_FrameData_O[13] ,
    \Tile_X5Y14_FrameData_O[12] ,
    \Tile_X5Y14_FrameData_O[11] ,
    \Tile_X5Y14_FrameData_O[10] ,
    \Tile_X5Y14_FrameData_O[9] ,
    \Tile_X5Y14_FrameData_O[8] ,
    \Tile_X5Y14_FrameData_O[7] ,
    \Tile_X5Y14_FrameData_O[6] ,
    \Tile_X5Y14_FrameData_O[5] ,
    \Tile_X5Y14_FrameData_O[4] ,
    \Tile_X5Y14_FrameData_O[3] ,
    \Tile_X5Y14_FrameData_O[2] ,
    \Tile_X5Y14_FrameData_O[1] ,
    \Tile_X5Y14_FrameData_O[0] }),
    .FrameData_O({\Tile_X6Y14_FrameData_O[31] ,
    \Tile_X6Y14_FrameData_O[30] ,
    \Tile_X6Y14_FrameData_O[29] ,
    \Tile_X6Y14_FrameData_O[28] ,
    \Tile_X6Y14_FrameData_O[27] ,
    \Tile_X6Y14_FrameData_O[26] ,
    \Tile_X6Y14_FrameData_O[25] ,
    \Tile_X6Y14_FrameData_O[24] ,
    \Tile_X6Y14_FrameData_O[23] ,
    \Tile_X6Y14_FrameData_O[22] ,
    \Tile_X6Y14_FrameData_O[21] ,
    \Tile_X6Y14_FrameData_O[20] ,
    \Tile_X6Y14_FrameData_O[19] ,
    \Tile_X6Y14_FrameData_O[18] ,
    \Tile_X6Y14_FrameData_O[17] ,
    \Tile_X6Y14_FrameData_O[16] ,
    \Tile_X6Y14_FrameData_O[15] ,
    \Tile_X6Y14_FrameData_O[14] ,
    \Tile_X6Y14_FrameData_O[13] ,
    \Tile_X6Y14_FrameData_O[12] ,
    \Tile_X6Y14_FrameData_O[11] ,
    \Tile_X6Y14_FrameData_O[10] ,
    \Tile_X6Y14_FrameData_O[9] ,
    \Tile_X6Y14_FrameData_O[8] ,
    \Tile_X6Y14_FrameData_O[7] ,
    \Tile_X6Y14_FrameData_O[6] ,
    \Tile_X6Y14_FrameData_O[5] ,
    \Tile_X6Y14_FrameData_O[4] ,
    \Tile_X6Y14_FrameData_O[3] ,
    \Tile_X6Y14_FrameData_O[2] ,
    \Tile_X6Y14_FrameData_O[1] ,
    \Tile_X6Y14_FrameData_O[0] }),
    .FrameStrobe({\Tile_X6Y15_FrameStrobe_O[19] ,
    \Tile_X6Y15_FrameStrobe_O[18] ,
    \Tile_X6Y15_FrameStrobe_O[17] ,
    \Tile_X6Y15_FrameStrobe_O[16] ,
    \Tile_X6Y15_FrameStrobe_O[15] ,
    \Tile_X6Y15_FrameStrobe_O[14] ,
    \Tile_X6Y15_FrameStrobe_O[13] ,
    \Tile_X6Y15_FrameStrobe_O[12] ,
    \Tile_X6Y15_FrameStrobe_O[11] ,
    \Tile_X6Y15_FrameStrobe_O[10] ,
    \Tile_X6Y15_FrameStrobe_O[9] ,
    \Tile_X6Y15_FrameStrobe_O[8] ,
    \Tile_X6Y15_FrameStrobe_O[7] ,
    \Tile_X6Y15_FrameStrobe_O[6] ,
    \Tile_X6Y15_FrameStrobe_O[5] ,
    \Tile_X6Y15_FrameStrobe_O[4] ,
    \Tile_X6Y15_FrameStrobe_O[3] ,
    \Tile_X6Y15_FrameStrobe_O[2] ,
    \Tile_X6Y15_FrameStrobe_O[1] ,
    \Tile_X6Y15_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X6Y14_FrameStrobe_O[19] ,
    \Tile_X6Y14_FrameStrobe_O[18] ,
    \Tile_X6Y14_FrameStrobe_O[17] ,
    \Tile_X6Y14_FrameStrobe_O[16] ,
    \Tile_X6Y14_FrameStrobe_O[15] ,
    \Tile_X6Y14_FrameStrobe_O[14] ,
    \Tile_X6Y14_FrameStrobe_O[13] ,
    \Tile_X6Y14_FrameStrobe_O[12] ,
    \Tile_X6Y14_FrameStrobe_O[11] ,
    \Tile_X6Y14_FrameStrobe_O[10] ,
    \Tile_X6Y14_FrameStrobe_O[9] ,
    \Tile_X6Y14_FrameStrobe_O[8] ,
    \Tile_X6Y14_FrameStrobe_O[7] ,
    \Tile_X6Y14_FrameStrobe_O[6] ,
    \Tile_X6Y14_FrameStrobe_O[5] ,
    \Tile_X6Y14_FrameStrobe_O[4] ,
    \Tile_X6Y14_FrameStrobe_O[3] ,
    \Tile_X6Y14_FrameStrobe_O[2] ,
    \Tile_X6Y14_FrameStrobe_O[1] ,
    \Tile_X6Y14_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X6Y14_N1BEG[3] ,
    \Tile_X6Y14_N1BEG[2] ,
    \Tile_X6Y14_N1BEG[1] ,
    \Tile_X6Y14_N1BEG[0] }),
    .N1END({\Tile_X6Y15_N1BEG[3] ,
    \Tile_X6Y15_N1BEG[2] ,
    \Tile_X6Y15_N1BEG[1] ,
    \Tile_X6Y15_N1BEG[0] }),
    .N2BEG({\Tile_X6Y14_N2BEG[7] ,
    \Tile_X6Y14_N2BEG[6] ,
    \Tile_X6Y14_N2BEG[5] ,
    \Tile_X6Y14_N2BEG[4] ,
    \Tile_X6Y14_N2BEG[3] ,
    \Tile_X6Y14_N2BEG[2] ,
    \Tile_X6Y14_N2BEG[1] ,
    \Tile_X6Y14_N2BEG[0] }),
    .N2BEGb({\Tile_X6Y14_N2BEGb[7] ,
    \Tile_X6Y14_N2BEGb[6] ,
    \Tile_X6Y14_N2BEGb[5] ,
    \Tile_X6Y14_N2BEGb[4] ,
    \Tile_X6Y14_N2BEGb[3] ,
    \Tile_X6Y14_N2BEGb[2] ,
    \Tile_X6Y14_N2BEGb[1] ,
    \Tile_X6Y14_N2BEGb[0] }),
    .N2END({\Tile_X6Y15_N2BEGb[7] ,
    \Tile_X6Y15_N2BEGb[6] ,
    \Tile_X6Y15_N2BEGb[5] ,
    \Tile_X6Y15_N2BEGb[4] ,
    \Tile_X6Y15_N2BEGb[3] ,
    \Tile_X6Y15_N2BEGb[2] ,
    \Tile_X6Y15_N2BEGb[1] ,
    \Tile_X6Y15_N2BEGb[0] }),
    .N2MID({\Tile_X6Y15_N2BEG[7] ,
    \Tile_X6Y15_N2BEG[6] ,
    \Tile_X6Y15_N2BEG[5] ,
    \Tile_X6Y15_N2BEG[4] ,
    \Tile_X6Y15_N2BEG[3] ,
    \Tile_X6Y15_N2BEG[2] ,
    \Tile_X6Y15_N2BEG[1] ,
    \Tile_X6Y15_N2BEG[0] }),
    .N4BEG({\Tile_X6Y14_N4BEG[15] ,
    \Tile_X6Y14_N4BEG[14] ,
    \Tile_X6Y14_N4BEG[13] ,
    \Tile_X6Y14_N4BEG[12] ,
    \Tile_X6Y14_N4BEG[11] ,
    \Tile_X6Y14_N4BEG[10] ,
    \Tile_X6Y14_N4BEG[9] ,
    \Tile_X6Y14_N4BEG[8] ,
    \Tile_X6Y14_N4BEG[7] ,
    \Tile_X6Y14_N4BEG[6] ,
    \Tile_X6Y14_N4BEG[5] ,
    \Tile_X6Y14_N4BEG[4] ,
    \Tile_X6Y14_N4BEG[3] ,
    \Tile_X6Y14_N4BEG[2] ,
    \Tile_X6Y14_N4BEG[1] ,
    \Tile_X6Y14_N4BEG[0] }),
    .N4END({\Tile_X6Y15_N4BEG[15] ,
    \Tile_X6Y15_N4BEG[14] ,
    \Tile_X6Y15_N4BEG[13] ,
    \Tile_X6Y15_N4BEG[12] ,
    \Tile_X6Y15_N4BEG[11] ,
    \Tile_X6Y15_N4BEG[10] ,
    \Tile_X6Y15_N4BEG[9] ,
    \Tile_X6Y15_N4BEG[8] ,
    \Tile_X6Y15_N4BEG[7] ,
    \Tile_X6Y15_N4BEG[6] ,
    \Tile_X6Y15_N4BEG[5] ,
    \Tile_X6Y15_N4BEG[4] ,
    \Tile_X6Y15_N4BEG[3] ,
    \Tile_X6Y15_N4BEG[2] ,
    \Tile_X6Y15_N4BEG[1] ,
    \Tile_X6Y15_N4BEG[0] }),
    .NN4BEG({\Tile_X6Y14_NN4BEG[15] ,
    \Tile_X6Y14_NN4BEG[14] ,
    \Tile_X6Y14_NN4BEG[13] ,
    \Tile_X6Y14_NN4BEG[12] ,
    \Tile_X6Y14_NN4BEG[11] ,
    \Tile_X6Y14_NN4BEG[10] ,
    \Tile_X6Y14_NN4BEG[9] ,
    \Tile_X6Y14_NN4BEG[8] ,
    \Tile_X6Y14_NN4BEG[7] ,
    \Tile_X6Y14_NN4BEG[6] ,
    \Tile_X6Y14_NN4BEG[5] ,
    \Tile_X6Y14_NN4BEG[4] ,
    \Tile_X6Y14_NN4BEG[3] ,
    \Tile_X6Y14_NN4BEG[2] ,
    \Tile_X6Y14_NN4BEG[1] ,
    \Tile_X6Y14_NN4BEG[0] }),
    .NN4END({\Tile_X6Y15_NN4BEG[15] ,
    \Tile_X6Y15_NN4BEG[14] ,
    \Tile_X6Y15_NN4BEG[13] ,
    \Tile_X6Y15_NN4BEG[12] ,
    \Tile_X6Y15_NN4BEG[11] ,
    \Tile_X6Y15_NN4BEG[10] ,
    \Tile_X6Y15_NN4BEG[9] ,
    \Tile_X6Y15_NN4BEG[8] ,
    \Tile_X6Y15_NN4BEG[7] ,
    \Tile_X6Y15_NN4BEG[6] ,
    \Tile_X6Y15_NN4BEG[5] ,
    \Tile_X6Y15_NN4BEG[4] ,
    \Tile_X6Y15_NN4BEG[3] ,
    \Tile_X6Y15_NN4BEG[2] ,
    \Tile_X6Y15_NN4BEG[1] ,
    \Tile_X6Y15_NN4BEG[0] }),
    .S1BEG({\Tile_X6Y14_S1BEG[3] ,
    \Tile_X6Y14_S1BEG[2] ,
    \Tile_X6Y14_S1BEG[1] ,
    \Tile_X6Y14_S1BEG[0] }),
    .S1END({\Tile_X6Y13_S1BEG[3] ,
    \Tile_X6Y13_S1BEG[2] ,
    \Tile_X6Y13_S1BEG[1] ,
    \Tile_X6Y13_S1BEG[0] }),
    .S2BEG({\Tile_X6Y14_S2BEG[7] ,
    \Tile_X6Y14_S2BEG[6] ,
    \Tile_X6Y14_S2BEG[5] ,
    \Tile_X6Y14_S2BEG[4] ,
    \Tile_X6Y14_S2BEG[3] ,
    \Tile_X6Y14_S2BEG[2] ,
    \Tile_X6Y14_S2BEG[1] ,
    \Tile_X6Y14_S2BEG[0] }),
    .S2BEGb({\Tile_X6Y14_S2BEGb[7] ,
    \Tile_X6Y14_S2BEGb[6] ,
    \Tile_X6Y14_S2BEGb[5] ,
    \Tile_X6Y14_S2BEGb[4] ,
    \Tile_X6Y14_S2BEGb[3] ,
    \Tile_X6Y14_S2BEGb[2] ,
    \Tile_X6Y14_S2BEGb[1] ,
    \Tile_X6Y14_S2BEGb[0] }),
    .S2END({\Tile_X6Y13_S2BEGb[7] ,
    \Tile_X6Y13_S2BEGb[6] ,
    \Tile_X6Y13_S2BEGb[5] ,
    \Tile_X6Y13_S2BEGb[4] ,
    \Tile_X6Y13_S2BEGb[3] ,
    \Tile_X6Y13_S2BEGb[2] ,
    \Tile_X6Y13_S2BEGb[1] ,
    \Tile_X6Y13_S2BEGb[0] }),
    .S2MID({\Tile_X6Y13_S2BEG[7] ,
    \Tile_X6Y13_S2BEG[6] ,
    \Tile_X6Y13_S2BEG[5] ,
    \Tile_X6Y13_S2BEG[4] ,
    \Tile_X6Y13_S2BEG[3] ,
    \Tile_X6Y13_S2BEG[2] ,
    \Tile_X6Y13_S2BEG[1] ,
    \Tile_X6Y13_S2BEG[0] }),
    .S4BEG({\Tile_X6Y14_S4BEG[15] ,
    \Tile_X6Y14_S4BEG[14] ,
    \Tile_X6Y14_S4BEG[13] ,
    \Tile_X6Y14_S4BEG[12] ,
    \Tile_X6Y14_S4BEG[11] ,
    \Tile_X6Y14_S4BEG[10] ,
    \Tile_X6Y14_S4BEG[9] ,
    \Tile_X6Y14_S4BEG[8] ,
    \Tile_X6Y14_S4BEG[7] ,
    \Tile_X6Y14_S4BEG[6] ,
    \Tile_X6Y14_S4BEG[5] ,
    \Tile_X6Y14_S4BEG[4] ,
    \Tile_X6Y14_S4BEG[3] ,
    \Tile_X6Y14_S4BEG[2] ,
    \Tile_X6Y14_S4BEG[1] ,
    \Tile_X6Y14_S4BEG[0] }),
    .S4END({\Tile_X6Y13_S4BEG[15] ,
    \Tile_X6Y13_S4BEG[14] ,
    \Tile_X6Y13_S4BEG[13] ,
    \Tile_X6Y13_S4BEG[12] ,
    \Tile_X6Y13_S4BEG[11] ,
    \Tile_X6Y13_S4BEG[10] ,
    \Tile_X6Y13_S4BEG[9] ,
    \Tile_X6Y13_S4BEG[8] ,
    \Tile_X6Y13_S4BEG[7] ,
    \Tile_X6Y13_S4BEG[6] ,
    \Tile_X6Y13_S4BEG[5] ,
    \Tile_X6Y13_S4BEG[4] ,
    \Tile_X6Y13_S4BEG[3] ,
    \Tile_X6Y13_S4BEG[2] ,
    \Tile_X6Y13_S4BEG[1] ,
    \Tile_X6Y13_S4BEG[0] }),
    .SS4BEG({\Tile_X6Y14_SS4BEG[15] ,
    \Tile_X6Y14_SS4BEG[14] ,
    \Tile_X6Y14_SS4BEG[13] ,
    \Tile_X6Y14_SS4BEG[12] ,
    \Tile_X6Y14_SS4BEG[11] ,
    \Tile_X6Y14_SS4BEG[10] ,
    \Tile_X6Y14_SS4BEG[9] ,
    \Tile_X6Y14_SS4BEG[8] ,
    \Tile_X6Y14_SS4BEG[7] ,
    \Tile_X6Y14_SS4BEG[6] ,
    \Tile_X6Y14_SS4BEG[5] ,
    \Tile_X6Y14_SS4BEG[4] ,
    \Tile_X6Y14_SS4BEG[3] ,
    \Tile_X6Y14_SS4BEG[2] ,
    \Tile_X6Y14_SS4BEG[1] ,
    \Tile_X6Y14_SS4BEG[0] }),
    .SS4END({\Tile_X6Y13_SS4BEG[15] ,
    \Tile_X6Y13_SS4BEG[14] ,
    \Tile_X6Y13_SS4BEG[13] ,
    \Tile_X6Y13_SS4BEG[12] ,
    \Tile_X6Y13_SS4BEG[11] ,
    \Tile_X6Y13_SS4BEG[10] ,
    \Tile_X6Y13_SS4BEG[9] ,
    \Tile_X6Y13_SS4BEG[8] ,
    \Tile_X6Y13_SS4BEG[7] ,
    \Tile_X6Y13_SS4BEG[6] ,
    \Tile_X6Y13_SS4BEG[5] ,
    \Tile_X6Y13_SS4BEG[4] ,
    \Tile_X6Y13_SS4BEG[3] ,
    \Tile_X6Y13_SS4BEG[2] ,
    \Tile_X6Y13_SS4BEG[1] ,
    \Tile_X6Y13_SS4BEG[0] }),
    .W1BEG({\Tile_X6Y14_W1BEG[3] ,
    \Tile_X6Y14_W1BEG[2] ,
    \Tile_X6Y14_W1BEG[1] ,
    \Tile_X6Y14_W1BEG[0] }),
    .W1END({\Tile_X7Y14_W1BEG[3] ,
    \Tile_X7Y14_W1BEG[2] ,
    \Tile_X7Y14_W1BEG[1] ,
    \Tile_X7Y14_W1BEG[0] }),
    .W2BEG({\Tile_X6Y14_W2BEG[7] ,
    \Tile_X6Y14_W2BEG[6] ,
    \Tile_X6Y14_W2BEG[5] ,
    \Tile_X6Y14_W2BEG[4] ,
    \Tile_X6Y14_W2BEG[3] ,
    \Tile_X6Y14_W2BEG[2] ,
    \Tile_X6Y14_W2BEG[1] ,
    \Tile_X6Y14_W2BEG[0] }),
    .W2BEGb({\Tile_X6Y14_W2BEGb[7] ,
    \Tile_X6Y14_W2BEGb[6] ,
    \Tile_X6Y14_W2BEGb[5] ,
    \Tile_X6Y14_W2BEGb[4] ,
    \Tile_X6Y14_W2BEGb[3] ,
    \Tile_X6Y14_W2BEGb[2] ,
    \Tile_X6Y14_W2BEGb[1] ,
    \Tile_X6Y14_W2BEGb[0] }),
    .W2END({\Tile_X7Y14_W2BEGb[7] ,
    \Tile_X7Y14_W2BEGb[6] ,
    \Tile_X7Y14_W2BEGb[5] ,
    \Tile_X7Y14_W2BEGb[4] ,
    \Tile_X7Y14_W2BEGb[3] ,
    \Tile_X7Y14_W2BEGb[2] ,
    \Tile_X7Y14_W2BEGb[1] ,
    \Tile_X7Y14_W2BEGb[0] }),
    .W2MID({\Tile_X7Y14_W2BEG[7] ,
    \Tile_X7Y14_W2BEG[6] ,
    \Tile_X7Y14_W2BEG[5] ,
    \Tile_X7Y14_W2BEG[4] ,
    \Tile_X7Y14_W2BEG[3] ,
    \Tile_X7Y14_W2BEG[2] ,
    \Tile_X7Y14_W2BEG[1] ,
    \Tile_X7Y14_W2BEG[0] }),
    .W6BEG({\Tile_X6Y14_W6BEG[11] ,
    \Tile_X6Y14_W6BEG[10] ,
    \Tile_X6Y14_W6BEG[9] ,
    \Tile_X6Y14_W6BEG[8] ,
    \Tile_X6Y14_W6BEG[7] ,
    \Tile_X6Y14_W6BEG[6] ,
    \Tile_X6Y14_W6BEG[5] ,
    \Tile_X6Y14_W6BEG[4] ,
    \Tile_X6Y14_W6BEG[3] ,
    \Tile_X6Y14_W6BEG[2] ,
    \Tile_X6Y14_W6BEG[1] ,
    \Tile_X6Y14_W6BEG[0] }),
    .W6END({\Tile_X7Y14_W6BEG[11] ,
    \Tile_X7Y14_W6BEG[10] ,
    \Tile_X7Y14_W6BEG[9] ,
    \Tile_X7Y14_W6BEG[8] ,
    \Tile_X7Y14_W6BEG[7] ,
    \Tile_X7Y14_W6BEG[6] ,
    \Tile_X7Y14_W6BEG[5] ,
    \Tile_X7Y14_W6BEG[4] ,
    \Tile_X7Y14_W6BEG[3] ,
    \Tile_X7Y14_W6BEG[2] ,
    \Tile_X7Y14_W6BEG[1] ,
    \Tile_X7Y14_W6BEG[0] }),
    .WW4BEG({\Tile_X6Y14_WW4BEG[15] ,
    \Tile_X6Y14_WW4BEG[14] ,
    \Tile_X6Y14_WW4BEG[13] ,
    \Tile_X6Y14_WW4BEG[12] ,
    \Tile_X6Y14_WW4BEG[11] ,
    \Tile_X6Y14_WW4BEG[10] ,
    \Tile_X6Y14_WW4BEG[9] ,
    \Tile_X6Y14_WW4BEG[8] ,
    \Tile_X6Y14_WW4BEG[7] ,
    \Tile_X6Y14_WW4BEG[6] ,
    \Tile_X6Y14_WW4BEG[5] ,
    \Tile_X6Y14_WW4BEG[4] ,
    \Tile_X6Y14_WW4BEG[3] ,
    \Tile_X6Y14_WW4BEG[2] ,
    \Tile_X6Y14_WW4BEG[1] ,
    \Tile_X6Y14_WW4BEG[0] }),
    .WW4END({\Tile_X7Y14_WW4BEG[15] ,
    \Tile_X7Y14_WW4BEG[14] ,
    \Tile_X7Y14_WW4BEG[13] ,
    \Tile_X7Y14_WW4BEG[12] ,
    \Tile_X7Y14_WW4BEG[11] ,
    \Tile_X7Y14_WW4BEG[10] ,
    \Tile_X7Y14_WW4BEG[9] ,
    \Tile_X7Y14_WW4BEG[8] ,
    \Tile_X7Y14_WW4BEG[7] ,
    \Tile_X7Y14_WW4BEG[6] ,
    \Tile_X7Y14_WW4BEG[5] ,
    \Tile_X7Y14_WW4BEG[4] ,
    \Tile_X7Y14_WW4BEG[3] ,
    \Tile_X7Y14_WW4BEG[2] ,
    \Tile_X7Y14_WW4BEG[1] ,
    \Tile_X7Y14_WW4BEG[0] }));
 S_CPU_IF Tile_X6Y15_S_CPU_IF (.Co(Tile_X6Y15_Co),
    .I_top0(Tile_X6Y15_I_top0),
    .I_top1(Tile_X6Y15_I_top1),
    .I_top10(Tile_X6Y15_I_top10),
    .I_top11(Tile_X6Y15_I_top11),
    .I_top12(Tile_X6Y15_I_top12),
    .I_top13(Tile_X6Y15_I_top13),
    .I_top14(Tile_X6Y15_I_top14),
    .I_top15(Tile_X6Y15_I_top15),
    .I_top2(Tile_X6Y15_I_top2),
    .I_top3(Tile_X6Y15_I_top3),
    .I_top4(Tile_X6Y15_I_top4),
    .I_top5(Tile_X6Y15_I_top5),
    .I_top6(Tile_X6Y15_I_top6),
    .I_top7(Tile_X6Y15_I_top7),
    .I_top8(Tile_X6Y15_I_top8),
    .I_top9(Tile_X6Y15_I_top9),
    .O_top0(Tile_X6Y15_O_top0),
    .O_top1(Tile_X6Y15_O_top1),
    .O_top10(Tile_X6Y15_O_top10),
    .O_top11(Tile_X6Y15_O_top11),
    .O_top12(Tile_X6Y15_O_top12),
    .O_top13(Tile_X6Y15_O_top13),
    .O_top14(Tile_X6Y15_O_top14),
    .O_top15(Tile_X6Y15_O_top15),
    .O_top2(Tile_X6Y15_O_top2),
    .O_top3(Tile_X6Y15_O_top3),
    .O_top4(Tile_X6Y15_O_top4),
    .O_top5(Tile_X6Y15_O_top5),
    .O_top6(Tile_X6Y15_O_top6),
    .O_top7(Tile_X6Y15_O_top7),
    .O_top8(Tile_X6Y15_O_top8),
    .O_top9(Tile_X6Y15_O_top9),
    .UserCLK(UserCLK),
    .UserCLKo(Tile_X6Y15_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .FrameData({\Tile_X5Y15_FrameData_O[31] ,
    \Tile_X5Y15_FrameData_O[30] ,
    \Tile_X5Y15_FrameData_O[29] ,
    \Tile_X5Y15_FrameData_O[28] ,
    \Tile_X5Y15_FrameData_O[27] ,
    \Tile_X5Y15_FrameData_O[26] ,
    \Tile_X5Y15_FrameData_O[25] ,
    \Tile_X5Y15_FrameData_O[24] ,
    \Tile_X5Y15_FrameData_O[23] ,
    \Tile_X5Y15_FrameData_O[22] ,
    \Tile_X5Y15_FrameData_O[21] ,
    \Tile_X5Y15_FrameData_O[20] ,
    \Tile_X5Y15_FrameData_O[19] ,
    \Tile_X5Y15_FrameData_O[18] ,
    \Tile_X5Y15_FrameData_O[17] ,
    \Tile_X5Y15_FrameData_O[16] ,
    \Tile_X5Y15_FrameData_O[15] ,
    \Tile_X5Y15_FrameData_O[14] ,
    \Tile_X5Y15_FrameData_O[13] ,
    \Tile_X5Y15_FrameData_O[12] ,
    \Tile_X5Y15_FrameData_O[11] ,
    \Tile_X5Y15_FrameData_O[10] ,
    \Tile_X5Y15_FrameData_O[9] ,
    \Tile_X5Y15_FrameData_O[8] ,
    \Tile_X5Y15_FrameData_O[7] ,
    \Tile_X5Y15_FrameData_O[6] ,
    \Tile_X5Y15_FrameData_O[5] ,
    \Tile_X5Y15_FrameData_O[4] ,
    \Tile_X5Y15_FrameData_O[3] ,
    \Tile_X5Y15_FrameData_O[2] ,
    \Tile_X5Y15_FrameData_O[1] ,
    \Tile_X5Y15_FrameData_O[0] }),
    .FrameData_O({\Tile_X6Y15_FrameData_O[31] ,
    \Tile_X6Y15_FrameData_O[30] ,
    \Tile_X6Y15_FrameData_O[29] ,
    \Tile_X6Y15_FrameData_O[28] ,
    \Tile_X6Y15_FrameData_O[27] ,
    \Tile_X6Y15_FrameData_O[26] ,
    \Tile_X6Y15_FrameData_O[25] ,
    \Tile_X6Y15_FrameData_O[24] ,
    \Tile_X6Y15_FrameData_O[23] ,
    \Tile_X6Y15_FrameData_O[22] ,
    \Tile_X6Y15_FrameData_O[21] ,
    \Tile_X6Y15_FrameData_O[20] ,
    \Tile_X6Y15_FrameData_O[19] ,
    \Tile_X6Y15_FrameData_O[18] ,
    \Tile_X6Y15_FrameData_O[17] ,
    \Tile_X6Y15_FrameData_O[16] ,
    \Tile_X6Y15_FrameData_O[15] ,
    \Tile_X6Y15_FrameData_O[14] ,
    \Tile_X6Y15_FrameData_O[13] ,
    \Tile_X6Y15_FrameData_O[12] ,
    \Tile_X6Y15_FrameData_O[11] ,
    \Tile_X6Y15_FrameData_O[10] ,
    \Tile_X6Y15_FrameData_O[9] ,
    \Tile_X6Y15_FrameData_O[8] ,
    \Tile_X6Y15_FrameData_O[7] ,
    \Tile_X6Y15_FrameData_O[6] ,
    \Tile_X6Y15_FrameData_O[5] ,
    \Tile_X6Y15_FrameData_O[4] ,
    \Tile_X6Y15_FrameData_O[3] ,
    \Tile_X6Y15_FrameData_O[2] ,
    \Tile_X6Y15_FrameData_O[1] ,
    \Tile_X6Y15_FrameData_O[0] }),
    .FrameStrobe({FrameStrobe[139],
    FrameStrobe[138],
    FrameStrobe[137],
    FrameStrobe[136],
    FrameStrobe[135],
    FrameStrobe[134],
    FrameStrobe[133],
    FrameStrobe[132],
    FrameStrobe[131],
    FrameStrobe[130],
    FrameStrobe[129],
    FrameStrobe[128],
    FrameStrobe[127],
    FrameStrobe[126],
    FrameStrobe[125],
    FrameStrobe[124],
    FrameStrobe[123],
    FrameStrobe[122],
    FrameStrobe[121],
    FrameStrobe[120]}),
    .FrameStrobe_O({\Tile_X6Y15_FrameStrobe_O[19] ,
    \Tile_X6Y15_FrameStrobe_O[18] ,
    \Tile_X6Y15_FrameStrobe_O[17] ,
    \Tile_X6Y15_FrameStrobe_O[16] ,
    \Tile_X6Y15_FrameStrobe_O[15] ,
    \Tile_X6Y15_FrameStrobe_O[14] ,
    \Tile_X6Y15_FrameStrobe_O[13] ,
    \Tile_X6Y15_FrameStrobe_O[12] ,
    \Tile_X6Y15_FrameStrobe_O[11] ,
    \Tile_X6Y15_FrameStrobe_O[10] ,
    \Tile_X6Y15_FrameStrobe_O[9] ,
    \Tile_X6Y15_FrameStrobe_O[8] ,
    \Tile_X6Y15_FrameStrobe_O[7] ,
    \Tile_X6Y15_FrameStrobe_O[6] ,
    \Tile_X6Y15_FrameStrobe_O[5] ,
    \Tile_X6Y15_FrameStrobe_O[4] ,
    \Tile_X6Y15_FrameStrobe_O[3] ,
    \Tile_X6Y15_FrameStrobe_O[2] ,
    \Tile_X6Y15_FrameStrobe_O[1] ,
    \Tile_X6Y15_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X6Y15_N1BEG[3] ,
    \Tile_X6Y15_N1BEG[2] ,
    \Tile_X6Y15_N1BEG[1] ,
    \Tile_X6Y15_N1BEG[0] }),
    .N2BEG({\Tile_X6Y15_N2BEG[7] ,
    \Tile_X6Y15_N2BEG[6] ,
    \Tile_X6Y15_N2BEG[5] ,
    \Tile_X6Y15_N2BEG[4] ,
    \Tile_X6Y15_N2BEG[3] ,
    \Tile_X6Y15_N2BEG[2] ,
    \Tile_X6Y15_N2BEG[1] ,
    \Tile_X6Y15_N2BEG[0] }),
    .N2BEGb({\Tile_X6Y15_N2BEGb[7] ,
    \Tile_X6Y15_N2BEGb[6] ,
    \Tile_X6Y15_N2BEGb[5] ,
    \Tile_X6Y15_N2BEGb[4] ,
    \Tile_X6Y15_N2BEGb[3] ,
    \Tile_X6Y15_N2BEGb[2] ,
    \Tile_X6Y15_N2BEGb[1] ,
    \Tile_X6Y15_N2BEGb[0] }),
    .N4BEG({\Tile_X6Y15_N4BEG[15] ,
    \Tile_X6Y15_N4BEG[14] ,
    \Tile_X6Y15_N4BEG[13] ,
    \Tile_X6Y15_N4BEG[12] ,
    \Tile_X6Y15_N4BEG[11] ,
    \Tile_X6Y15_N4BEG[10] ,
    \Tile_X6Y15_N4BEG[9] ,
    \Tile_X6Y15_N4BEG[8] ,
    \Tile_X6Y15_N4BEG[7] ,
    \Tile_X6Y15_N4BEG[6] ,
    \Tile_X6Y15_N4BEG[5] ,
    \Tile_X6Y15_N4BEG[4] ,
    \Tile_X6Y15_N4BEG[3] ,
    \Tile_X6Y15_N4BEG[2] ,
    \Tile_X6Y15_N4BEG[1] ,
    \Tile_X6Y15_N4BEG[0] }),
    .NN4BEG({\Tile_X6Y15_NN4BEG[15] ,
    \Tile_X6Y15_NN4BEG[14] ,
    \Tile_X6Y15_NN4BEG[13] ,
    \Tile_X6Y15_NN4BEG[12] ,
    \Tile_X6Y15_NN4BEG[11] ,
    \Tile_X6Y15_NN4BEG[10] ,
    \Tile_X6Y15_NN4BEG[9] ,
    \Tile_X6Y15_NN4BEG[8] ,
    \Tile_X6Y15_NN4BEG[7] ,
    \Tile_X6Y15_NN4BEG[6] ,
    \Tile_X6Y15_NN4BEG[5] ,
    \Tile_X6Y15_NN4BEG[4] ,
    \Tile_X6Y15_NN4BEG[3] ,
    \Tile_X6Y15_NN4BEG[2] ,
    \Tile_X6Y15_NN4BEG[1] ,
    \Tile_X6Y15_NN4BEG[0] }),
    .S1END({\Tile_X6Y14_S1BEG[3] ,
    \Tile_X6Y14_S1BEG[2] ,
    \Tile_X6Y14_S1BEG[1] ,
    \Tile_X6Y14_S1BEG[0] }),
    .S2END({\Tile_X6Y14_S2BEGb[7] ,
    \Tile_X6Y14_S2BEGb[6] ,
    \Tile_X6Y14_S2BEGb[5] ,
    \Tile_X6Y14_S2BEGb[4] ,
    \Tile_X6Y14_S2BEGb[3] ,
    \Tile_X6Y14_S2BEGb[2] ,
    \Tile_X6Y14_S2BEGb[1] ,
    \Tile_X6Y14_S2BEGb[0] }),
    .S2MID({\Tile_X6Y14_S2BEG[7] ,
    \Tile_X6Y14_S2BEG[6] ,
    \Tile_X6Y14_S2BEG[5] ,
    \Tile_X6Y14_S2BEG[4] ,
    \Tile_X6Y14_S2BEG[3] ,
    \Tile_X6Y14_S2BEG[2] ,
    \Tile_X6Y14_S2BEG[1] ,
    \Tile_X6Y14_S2BEG[0] }),
    .S4END({\Tile_X6Y14_S4BEG[15] ,
    \Tile_X6Y14_S4BEG[14] ,
    \Tile_X6Y14_S4BEG[13] ,
    \Tile_X6Y14_S4BEG[12] ,
    \Tile_X6Y14_S4BEG[11] ,
    \Tile_X6Y14_S4BEG[10] ,
    \Tile_X6Y14_S4BEG[9] ,
    \Tile_X6Y14_S4BEG[8] ,
    \Tile_X6Y14_S4BEG[7] ,
    \Tile_X6Y14_S4BEG[6] ,
    \Tile_X6Y14_S4BEG[5] ,
    \Tile_X6Y14_S4BEG[4] ,
    \Tile_X6Y14_S4BEG[3] ,
    \Tile_X6Y14_S4BEG[2] ,
    \Tile_X6Y14_S4BEG[1] ,
    \Tile_X6Y14_S4BEG[0] }),
    .SS4END({\Tile_X6Y14_SS4BEG[15] ,
    \Tile_X6Y14_SS4BEG[14] ,
    \Tile_X6Y14_SS4BEG[13] ,
    \Tile_X6Y14_SS4BEG[12] ,
    \Tile_X6Y14_SS4BEG[11] ,
    \Tile_X6Y14_SS4BEG[10] ,
    \Tile_X6Y14_SS4BEG[9] ,
    \Tile_X6Y14_SS4BEG[8] ,
    \Tile_X6Y14_SS4BEG[7] ,
    \Tile_X6Y14_SS4BEG[6] ,
    \Tile_X6Y14_SS4BEG[5] ,
    \Tile_X6Y14_SS4BEG[4] ,
    \Tile_X6Y14_SS4BEG[3] ,
    \Tile_X6Y14_SS4BEG[2] ,
    \Tile_X6Y14_SS4BEG[1] ,
    \Tile_X6Y14_SS4BEG[0] }));
 LUT4AB Tile_X6Y1_LUT4AB (.Ci(Tile_X6Y2_Co),
    .Co(Tile_X6Y1_Co),
    .UserCLK(Tile_X6Y2_UserCLKo),
    .UserCLKo(Tile_X6Y1_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X6Y1_E1BEG[3] ,
    \Tile_X6Y1_E1BEG[2] ,
    \Tile_X6Y1_E1BEG[1] ,
    \Tile_X6Y1_E1BEG[0] }),
    .E1END({\Tile_X5Y1_E1BEG[3] ,
    \Tile_X5Y1_E1BEG[2] ,
    \Tile_X5Y1_E1BEG[1] ,
    \Tile_X5Y1_E1BEG[0] }),
    .E2BEG({\Tile_X6Y1_E2BEG[7] ,
    \Tile_X6Y1_E2BEG[6] ,
    \Tile_X6Y1_E2BEG[5] ,
    \Tile_X6Y1_E2BEG[4] ,
    \Tile_X6Y1_E2BEG[3] ,
    \Tile_X6Y1_E2BEG[2] ,
    \Tile_X6Y1_E2BEG[1] ,
    \Tile_X6Y1_E2BEG[0] }),
    .E2BEGb({\Tile_X6Y1_E2BEGb[7] ,
    \Tile_X6Y1_E2BEGb[6] ,
    \Tile_X6Y1_E2BEGb[5] ,
    \Tile_X6Y1_E2BEGb[4] ,
    \Tile_X6Y1_E2BEGb[3] ,
    \Tile_X6Y1_E2BEGb[2] ,
    \Tile_X6Y1_E2BEGb[1] ,
    \Tile_X6Y1_E2BEGb[0] }),
    .E2END({\Tile_X5Y1_E2BEGb[7] ,
    \Tile_X5Y1_E2BEGb[6] ,
    \Tile_X5Y1_E2BEGb[5] ,
    \Tile_X5Y1_E2BEGb[4] ,
    \Tile_X5Y1_E2BEGb[3] ,
    \Tile_X5Y1_E2BEGb[2] ,
    \Tile_X5Y1_E2BEGb[1] ,
    \Tile_X5Y1_E2BEGb[0] }),
    .E2MID({\Tile_X5Y1_E2BEG[7] ,
    \Tile_X5Y1_E2BEG[6] ,
    \Tile_X5Y1_E2BEG[5] ,
    \Tile_X5Y1_E2BEG[4] ,
    \Tile_X5Y1_E2BEG[3] ,
    \Tile_X5Y1_E2BEG[2] ,
    \Tile_X5Y1_E2BEG[1] ,
    \Tile_X5Y1_E2BEG[0] }),
    .E6BEG({\Tile_X6Y1_E6BEG[11] ,
    \Tile_X6Y1_E6BEG[10] ,
    \Tile_X6Y1_E6BEG[9] ,
    \Tile_X6Y1_E6BEG[8] ,
    \Tile_X6Y1_E6BEG[7] ,
    \Tile_X6Y1_E6BEG[6] ,
    \Tile_X6Y1_E6BEG[5] ,
    \Tile_X6Y1_E6BEG[4] ,
    \Tile_X6Y1_E6BEG[3] ,
    \Tile_X6Y1_E6BEG[2] ,
    \Tile_X6Y1_E6BEG[1] ,
    \Tile_X6Y1_E6BEG[0] }),
    .E6END({\Tile_X5Y1_E6BEG[11] ,
    \Tile_X5Y1_E6BEG[10] ,
    \Tile_X5Y1_E6BEG[9] ,
    \Tile_X5Y1_E6BEG[8] ,
    \Tile_X5Y1_E6BEG[7] ,
    \Tile_X5Y1_E6BEG[6] ,
    \Tile_X5Y1_E6BEG[5] ,
    \Tile_X5Y1_E6BEG[4] ,
    \Tile_X5Y1_E6BEG[3] ,
    \Tile_X5Y1_E6BEG[2] ,
    \Tile_X5Y1_E6BEG[1] ,
    \Tile_X5Y1_E6BEG[0] }),
    .EE4BEG({\Tile_X6Y1_EE4BEG[15] ,
    \Tile_X6Y1_EE4BEG[14] ,
    \Tile_X6Y1_EE4BEG[13] ,
    \Tile_X6Y1_EE4BEG[12] ,
    \Tile_X6Y1_EE4BEG[11] ,
    \Tile_X6Y1_EE4BEG[10] ,
    \Tile_X6Y1_EE4BEG[9] ,
    \Tile_X6Y1_EE4BEG[8] ,
    \Tile_X6Y1_EE4BEG[7] ,
    \Tile_X6Y1_EE4BEG[6] ,
    \Tile_X6Y1_EE4BEG[5] ,
    \Tile_X6Y1_EE4BEG[4] ,
    \Tile_X6Y1_EE4BEG[3] ,
    \Tile_X6Y1_EE4BEG[2] ,
    \Tile_X6Y1_EE4BEG[1] ,
    \Tile_X6Y1_EE4BEG[0] }),
    .EE4END({\Tile_X5Y1_EE4BEG[15] ,
    \Tile_X5Y1_EE4BEG[14] ,
    \Tile_X5Y1_EE4BEG[13] ,
    \Tile_X5Y1_EE4BEG[12] ,
    \Tile_X5Y1_EE4BEG[11] ,
    \Tile_X5Y1_EE4BEG[10] ,
    \Tile_X5Y1_EE4BEG[9] ,
    \Tile_X5Y1_EE4BEG[8] ,
    \Tile_X5Y1_EE4BEG[7] ,
    \Tile_X5Y1_EE4BEG[6] ,
    \Tile_X5Y1_EE4BEG[5] ,
    \Tile_X5Y1_EE4BEG[4] ,
    \Tile_X5Y1_EE4BEG[3] ,
    \Tile_X5Y1_EE4BEG[2] ,
    \Tile_X5Y1_EE4BEG[1] ,
    \Tile_X5Y1_EE4BEG[0] }),
    .FrameData({\Tile_X5Y1_FrameData_O[31] ,
    \Tile_X5Y1_FrameData_O[30] ,
    \Tile_X5Y1_FrameData_O[29] ,
    \Tile_X5Y1_FrameData_O[28] ,
    \Tile_X5Y1_FrameData_O[27] ,
    \Tile_X5Y1_FrameData_O[26] ,
    \Tile_X5Y1_FrameData_O[25] ,
    \Tile_X5Y1_FrameData_O[24] ,
    \Tile_X5Y1_FrameData_O[23] ,
    \Tile_X5Y1_FrameData_O[22] ,
    \Tile_X5Y1_FrameData_O[21] ,
    \Tile_X5Y1_FrameData_O[20] ,
    \Tile_X5Y1_FrameData_O[19] ,
    \Tile_X5Y1_FrameData_O[18] ,
    \Tile_X5Y1_FrameData_O[17] ,
    \Tile_X5Y1_FrameData_O[16] ,
    \Tile_X5Y1_FrameData_O[15] ,
    \Tile_X5Y1_FrameData_O[14] ,
    \Tile_X5Y1_FrameData_O[13] ,
    \Tile_X5Y1_FrameData_O[12] ,
    \Tile_X5Y1_FrameData_O[11] ,
    \Tile_X5Y1_FrameData_O[10] ,
    \Tile_X5Y1_FrameData_O[9] ,
    \Tile_X5Y1_FrameData_O[8] ,
    \Tile_X5Y1_FrameData_O[7] ,
    \Tile_X5Y1_FrameData_O[6] ,
    \Tile_X5Y1_FrameData_O[5] ,
    \Tile_X5Y1_FrameData_O[4] ,
    \Tile_X5Y1_FrameData_O[3] ,
    \Tile_X5Y1_FrameData_O[2] ,
    \Tile_X5Y1_FrameData_O[1] ,
    \Tile_X5Y1_FrameData_O[0] }),
    .FrameData_O({\Tile_X6Y1_FrameData_O[31] ,
    \Tile_X6Y1_FrameData_O[30] ,
    \Tile_X6Y1_FrameData_O[29] ,
    \Tile_X6Y1_FrameData_O[28] ,
    \Tile_X6Y1_FrameData_O[27] ,
    \Tile_X6Y1_FrameData_O[26] ,
    \Tile_X6Y1_FrameData_O[25] ,
    \Tile_X6Y1_FrameData_O[24] ,
    \Tile_X6Y1_FrameData_O[23] ,
    \Tile_X6Y1_FrameData_O[22] ,
    \Tile_X6Y1_FrameData_O[21] ,
    \Tile_X6Y1_FrameData_O[20] ,
    \Tile_X6Y1_FrameData_O[19] ,
    \Tile_X6Y1_FrameData_O[18] ,
    \Tile_X6Y1_FrameData_O[17] ,
    \Tile_X6Y1_FrameData_O[16] ,
    \Tile_X6Y1_FrameData_O[15] ,
    \Tile_X6Y1_FrameData_O[14] ,
    \Tile_X6Y1_FrameData_O[13] ,
    \Tile_X6Y1_FrameData_O[12] ,
    \Tile_X6Y1_FrameData_O[11] ,
    \Tile_X6Y1_FrameData_O[10] ,
    \Tile_X6Y1_FrameData_O[9] ,
    \Tile_X6Y1_FrameData_O[8] ,
    \Tile_X6Y1_FrameData_O[7] ,
    \Tile_X6Y1_FrameData_O[6] ,
    \Tile_X6Y1_FrameData_O[5] ,
    \Tile_X6Y1_FrameData_O[4] ,
    \Tile_X6Y1_FrameData_O[3] ,
    \Tile_X6Y1_FrameData_O[2] ,
    \Tile_X6Y1_FrameData_O[1] ,
    \Tile_X6Y1_FrameData_O[0] }),
    .FrameStrobe({\Tile_X6Y2_FrameStrobe_O[19] ,
    \Tile_X6Y2_FrameStrobe_O[18] ,
    \Tile_X6Y2_FrameStrobe_O[17] ,
    \Tile_X6Y2_FrameStrobe_O[16] ,
    \Tile_X6Y2_FrameStrobe_O[15] ,
    \Tile_X6Y2_FrameStrobe_O[14] ,
    \Tile_X6Y2_FrameStrobe_O[13] ,
    \Tile_X6Y2_FrameStrobe_O[12] ,
    \Tile_X6Y2_FrameStrobe_O[11] ,
    \Tile_X6Y2_FrameStrobe_O[10] ,
    \Tile_X6Y2_FrameStrobe_O[9] ,
    \Tile_X6Y2_FrameStrobe_O[8] ,
    \Tile_X6Y2_FrameStrobe_O[7] ,
    \Tile_X6Y2_FrameStrobe_O[6] ,
    \Tile_X6Y2_FrameStrobe_O[5] ,
    \Tile_X6Y2_FrameStrobe_O[4] ,
    \Tile_X6Y2_FrameStrobe_O[3] ,
    \Tile_X6Y2_FrameStrobe_O[2] ,
    \Tile_X6Y2_FrameStrobe_O[1] ,
    \Tile_X6Y2_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X6Y1_FrameStrobe_O[19] ,
    \Tile_X6Y1_FrameStrobe_O[18] ,
    \Tile_X6Y1_FrameStrobe_O[17] ,
    \Tile_X6Y1_FrameStrobe_O[16] ,
    \Tile_X6Y1_FrameStrobe_O[15] ,
    \Tile_X6Y1_FrameStrobe_O[14] ,
    \Tile_X6Y1_FrameStrobe_O[13] ,
    \Tile_X6Y1_FrameStrobe_O[12] ,
    \Tile_X6Y1_FrameStrobe_O[11] ,
    \Tile_X6Y1_FrameStrobe_O[10] ,
    \Tile_X6Y1_FrameStrobe_O[9] ,
    \Tile_X6Y1_FrameStrobe_O[8] ,
    \Tile_X6Y1_FrameStrobe_O[7] ,
    \Tile_X6Y1_FrameStrobe_O[6] ,
    \Tile_X6Y1_FrameStrobe_O[5] ,
    \Tile_X6Y1_FrameStrobe_O[4] ,
    \Tile_X6Y1_FrameStrobe_O[3] ,
    \Tile_X6Y1_FrameStrobe_O[2] ,
    \Tile_X6Y1_FrameStrobe_O[1] ,
    \Tile_X6Y1_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X6Y1_N1BEG[3] ,
    \Tile_X6Y1_N1BEG[2] ,
    \Tile_X6Y1_N1BEG[1] ,
    \Tile_X6Y1_N1BEG[0] }),
    .N1END({\Tile_X6Y2_N1BEG[3] ,
    \Tile_X6Y2_N1BEG[2] ,
    \Tile_X6Y2_N1BEG[1] ,
    \Tile_X6Y2_N1BEG[0] }),
    .N2BEG({\Tile_X6Y1_N2BEG[7] ,
    \Tile_X6Y1_N2BEG[6] ,
    \Tile_X6Y1_N2BEG[5] ,
    \Tile_X6Y1_N2BEG[4] ,
    \Tile_X6Y1_N2BEG[3] ,
    \Tile_X6Y1_N2BEG[2] ,
    \Tile_X6Y1_N2BEG[1] ,
    \Tile_X6Y1_N2BEG[0] }),
    .N2BEGb({\Tile_X6Y1_N2BEGb[7] ,
    \Tile_X6Y1_N2BEGb[6] ,
    \Tile_X6Y1_N2BEGb[5] ,
    \Tile_X6Y1_N2BEGb[4] ,
    \Tile_X6Y1_N2BEGb[3] ,
    \Tile_X6Y1_N2BEGb[2] ,
    \Tile_X6Y1_N2BEGb[1] ,
    \Tile_X6Y1_N2BEGb[0] }),
    .N2END({\Tile_X6Y2_N2BEGb[7] ,
    \Tile_X6Y2_N2BEGb[6] ,
    \Tile_X6Y2_N2BEGb[5] ,
    \Tile_X6Y2_N2BEGb[4] ,
    \Tile_X6Y2_N2BEGb[3] ,
    \Tile_X6Y2_N2BEGb[2] ,
    \Tile_X6Y2_N2BEGb[1] ,
    \Tile_X6Y2_N2BEGb[0] }),
    .N2MID({\Tile_X6Y2_N2BEG[7] ,
    \Tile_X6Y2_N2BEG[6] ,
    \Tile_X6Y2_N2BEG[5] ,
    \Tile_X6Y2_N2BEG[4] ,
    \Tile_X6Y2_N2BEG[3] ,
    \Tile_X6Y2_N2BEG[2] ,
    \Tile_X6Y2_N2BEG[1] ,
    \Tile_X6Y2_N2BEG[0] }),
    .N4BEG({\Tile_X6Y1_N4BEG[15] ,
    \Tile_X6Y1_N4BEG[14] ,
    \Tile_X6Y1_N4BEG[13] ,
    \Tile_X6Y1_N4BEG[12] ,
    \Tile_X6Y1_N4BEG[11] ,
    \Tile_X6Y1_N4BEG[10] ,
    \Tile_X6Y1_N4BEG[9] ,
    \Tile_X6Y1_N4BEG[8] ,
    \Tile_X6Y1_N4BEG[7] ,
    \Tile_X6Y1_N4BEG[6] ,
    \Tile_X6Y1_N4BEG[5] ,
    \Tile_X6Y1_N4BEG[4] ,
    \Tile_X6Y1_N4BEG[3] ,
    \Tile_X6Y1_N4BEG[2] ,
    \Tile_X6Y1_N4BEG[1] ,
    \Tile_X6Y1_N4BEG[0] }),
    .N4END({\Tile_X6Y2_N4BEG[15] ,
    \Tile_X6Y2_N4BEG[14] ,
    \Tile_X6Y2_N4BEG[13] ,
    \Tile_X6Y2_N4BEG[12] ,
    \Tile_X6Y2_N4BEG[11] ,
    \Tile_X6Y2_N4BEG[10] ,
    \Tile_X6Y2_N4BEG[9] ,
    \Tile_X6Y2_N4BEG[8] ,
    \Tile_X6Y2_N4BEG[7] ,
    \Tile_X6Y2_N4BEG[6] ,
    \Tile_X6Y2_N4BEG[5] ,
    \Tile_X6Y2_N4BEG[4] ,
    \Tile_X6Y2_N4BEG[3] ,
    \Tile_X6Y2_N4BEG[2] ,
    \Tile_X6Y2_N4BEG[1] ,
    \Tile_X6Y2_N4BEG[0] }),
    .NN4BEG({\Tile_X6Y1_NN4BEG[15] ,
    \Tile_X6Y1_NN4BEG[14] ,
    \Tile_X6Y1_NN4BEG[13] ,
    \Tile_X6Y1_NN4BEG[12] ,
    \Tile_X6Y1_NN4BEG[11] ,
    \Tile_X6Y1_NN4BEG[10] ,
    \Tile_X6Y1_NN4BEG[9] ,
    \Tile_X6Y1_NN4BEG[8] ,
    \Tile_X6Y1_NN4BEG[7] ,
    \Tile_X6Y1_NN4BEG[6] ,
    \Tile_X6Y1_NN4BEG[5] ,
    \Tile_X6Y1_NN4BEG[4] ,
    \Tile_X6Y1_NN4BEG[3] ,
    \Tile_X6Y1_NN4BEG[2] ,
    \Tile_X6Y1_NN4BEG[1] ,
    \Tile_X6Y1_NN4BEG[0] }),
    .NN4END({\Tile_X6Y2_NN4BEG[15] ,
    \Tile_X6Y2_NN4BEG[14] ,
    \Tile_X6Y2_NN4BEG[13] ,
    \Tile_X6Y2_NN4BEG[12] ,
    \Tile_X6Y2_NN4BEG[11] ,
    \Tile_X6Y2_NN4BEG[10] ,
    \Tile_X6Y2_NN4BEG[9] ,
    \Tile_X6Y2_NN4BEG[8] ,
    \Tile_X6Y2_NN4BEG[7] ,
    \Tile_X6Y2_NN4BEG[6] ,
    \Tile_X6Y2_NN4BEG[5] ,
    \Tile_X6Y2_NN4BEG[4] ,
    \Tile_X6Y2_NN4BEG[3] ,
    \Tile_X6Y2_NN4BEG[2] ,
    \Tile_X6Y2_NN4BEG[1] ,
    \Tile_X6Y2_NN4BEG[0] }),
    .S1BEG({\Tile_X6Y1_S1BEG[3] ,
    \Tile_X6Y1_S1BEG[2] ,
    \Tile_X6Y1_S1BEG[1] ,
    \Tile_X6Y1_S1BEG[0] }),
    .S1END({\Tile_X6Y0_S1BEG[3] ,
    \Tile_X6Y0_S1BEG[2] ,
    \Tile_X6Y0_S1BEG[1] ,
    \Tile_X6Y0_S1BEG[0] }),
    .S2BEG({\Tile_X6Y1_S2BEG[7] ,
    \Tile_X6Y1_S2BEG[6] ,
    \Tile_X6Y1_S2BEG[5] ,
    \Tile_X6Y1_S2BEG[4] ,
    \Tile_X6Y1_S2BEG[3] ,
    \Tile_X6Y1_S2BEG[2] ,
    \Tile_X6Y1_S2BEG[1] ,
    \Tile_X6Y1_S2BEG[0] }),
    .S2BEGb({\Tile_X6Y1_S2BEGb[7] ,
    \Tile_X6Y1_S2BEGb[6] ,
    \Tile_X6Y1_S2BEGb[5] ,
    \Tile_X6Y1_S2BEGb[4] ,
    \Tile_X6Y1_S2BEGb[3] ,
    \Tile_X6Y1_S2BEGb[2] ,
    \Tile_X6Y1_S2BEGb[1] ,
    \Tile_X6Y1_S2BEGb[0] }),
    .S2END({\Tile_X6Y0_S2BEGb[7] ,
    \Tile_X6Y0_S2BEGb[6] ,
    \Tile_X6Y0_S2BEGb[5] ,
    \Tile_X6Y0_S2BEGb[4] ,
    \Tile_X6Y0_S2BEGb[3] ,
    \Tile_X6Y0_S2BEGb[2] ,
    \Tile_X6Y0_S2BEGb[1] ,
    \Tile_X6Y0_S2BEGb[0] }),
    .S2MID({\Tile_X6Y0_S2BEG[7] ,
    \Tile_X6Y0_S2BEG[6] ,
    \Tile_X6Y0_S2BEG[5] ,
    \Tile_X6Y0_S2BEG[4] ,
    \Tile_X6Y0_S2BEG[3] ,
    \Tile_X6Y0_S2BEG[2] ,
    \Tile_X6Y0_S2BEG[1] ,
    \Tile_X6Y0_S2BEG[0] }),
    .S4BEG({\Tile_X6Y1_S4BEG[15] ,
    \Tile_X6Y1_S4BEG[14] ,
    \Tile_X6Y1_S4BEG[13] ,
    \Tile_X6Y1_S4BEG[12] ,
    \Tile_X6Y1_S4BEG[11] ,
    \Tile_X6Y1_S4BEG[10] ,
    \Tile_X6Y1_S4BEG[9] ,
    \Tile_X6Y1_S4BEG[8] ,
    \Tile_X6Y1_S4BEG[7] ,
    \Tile_X6Y1_S4BEG[6] ,
    \Tile_X6Y1_S4BEG[5] ,
    \Tile_X6Y1_S4BEG[4] ,
    \Tile_X6Y1_S4BEG[3] ,
    \Tile_X6Y1_S4BEG[2] ,
    \Tile_X6Y1_S4BEG[1] ,
    \Tile_X6Y1_S4BEG[0] }),
    .S4END({\Tile_X6Y0_S4BEG[15] ,
    \Tile_X6Y0_S4BEG[14] ,
    \Tile_X6Y0_S4BEG[13] ,
    \Tile_X6Y0_S4BEG[12] ,
    \Tile_X6Y0_S4BEG[11] ,
    \Tile_X6Y0_S4BEG[10] ,
    \Tile_X6Y0_S4BEG[9] ,
    \Tile_X6Y0_S4BEG[8] ,
    \Tile_X6Y0_S4BEG[7] ,
    \Tile_X6Y0_S4BEG[6] ,
    \Tile_X6Y0_S4BEG[5] ,
    \Tile_X6Y0_S4BEG[4] ,
    \Tile_X6Y0_S4BEG[3] ,
    \Tile_X6Y0_S4BEG[2] ,
    \Tile_X6Y0_S4BEG[1] ,
    \Tile_X6Y0_S4BEG[0] }),
    .SS4BEG({\Tile_X6Y1_SS4BEG[15] ,
    \Tile_X6Y1_SS4BEG[14] ,
    \Tile_X6Y1_SS4BEG[13] ,
    \Tile_X6Y1_SS4BEG[12] ,
    \Tile_X6Y1_SS4BEG[11] ,
    \Tile_X6Y1_SS4BEG[10] ,
    \Tile_X6Y1_SS4BEG[9] ,
    \Tile_X6Y1_SS4BEG[8] ,
    \Tile_X6Y1_SS4BEG[7] ,
    \Tile_X6Y1_SS4BEG[6] ,
    \Tile_X6Y1_SS4BEG[5] ,
    \Tile_X6Y1_SS4BEG[4] ,
    \Tile_X6Y1_SS4BEG[3] ,
    \Tile_X6Y1_SS4BEG[2] ,
    \Tile_X6Y1_SS4BEG[1] ,
    \Tile_X6Y1_SS4BEG[0] }),
    .SS4END({\Tile_X6Y0_SS4BEG[15] ,
    \Tile_X6Y0_SS4BEG[14] ,
    \Tile_X6Y0_SS4BEG[13] ,
    \Tile_X6Y0_SS4BEG[12] ,
    \Tile_X6Y0_SS4BEG[11] ,
    \Tile_X6Y0_SS4BEG[10] ,
    \Tile_X6Y0_SS4BEG[9] ,
    \Tile_X6Y0_SS4BEG[8] ,
    \Tile_X6Y0_SS4BEG[7] ,
    \Tile_X6Y0_SS4BEG[6] ,
    \Tile_X6Y0_SS4BEG[5] ,
    \Tile_X6Y0_SS4BEG[4] ,
    \Tile_X6Y0_SS4BEG[3] ,
    \Tile_X6Y0_SS4BEG[2] ,
    \Tile_X6Y0_SS4BEG[1] ,
    \Tile_X6Y0_SS4BEG[0] }),
    .W1BEG({\Tile_X6Y1_W1BEG[3] ,
    \Tile_X6Y1_W1BEG[2] ,
    \Tile_X6Y1_W1BEG[1] ,
    \Tile_X6Y1_W1BEG[0] }),
    .W1END({\Tile_X7Y1_W1BEG[3] ,
    \Tile_X7Y1_W1BEG[2] ,
    \Tile_X7Y1_W1BEG[1] ,
    \Tile_X7Y1_W1BEG[0] }),
    .W2BEG({\Tile_X6Y1_W2BEG[7] ,
    \Tile_X6Y1_W2BEG[6] ,
    \Tile_X6Y1_W2BEG[5] ,
    \Tile_X6Y1_W2BEG[4] ,
    \Tile_X6Y1_W2BEG[3] ,
    \Tile_X6Y1_W2BEG[2] ,
    \Tile_X6Y1_W2BEG[1] ,
    \Tile_X6Y1_W2BEG[0] }),
    .W2BEGb({\Tile_X6Y1_W2BEGb[7] ,
    \Tile_X6Y1_W2BEGb[6] ,
    \Tile_X6Y1_W2BEGb[5] ,
    \Tile_X6Y1_W2BEGb[4] ,
    \Tile_X6Y1_W2BEGb[3] ,
    \Tile_X6Y1_W2BEGb[2] ,
    \Tile_X6Y1_W2BEGb[1] ,
    \Tile_X6Y1_W2BEGb[0] }),
    .W2END({\Tile_X7Y1_W2BEGb[7] ,
    \Tile_X7Y1_W2BEGb[6] ,
    \Tile_X7Y1_W2BEGb[5] ,
    \Tile_X7Y1_W2BEGb[4] ,
    \Tile_X7Y1_W2BEGb[3] ,
    \Tile_X7Y1_W2BEGb[2] ,
    \Tile_X7Y1_W2BEGb[1] ,
    \Tile_X7Y1_W2BEGb[0] }),
    .W2MID({\Tile_X7Y1_W2BEG[7] ,
    \Tile_X7Y1_W2BEG[6] ,
    \Tile_X7Y1_W2BEG[5] ,
    \Tile_X7Y1_W2BEG[4] ,
    \Tile_X7Y1_W2BEG[3] ,
    \Tile_X7Y1_W2BEG[2] ,
    \Tile_X7Y1_W2BEG[1] ,
    \Tile_X7Y1_W2BEG[0] }),
    .W6BEG({\Tile_X6Y1_W6BEG[11] ,
    \Tile_X6Y1_W6BEG[10] ,
    \Tile_X6Y1_W6BEG[9] ,
    \Tile_X6Y1_W6BEG[8] ,
    \Tile_X6Y1_W6BEG[7] ,
    \Tile_X6Y1_W6BEG[6] ,
    \Tile_X6Y1_W6BEG[5] ,
    \Tile_X6Y1_W6BEG[4] ,
    \Tile_X6Y1_W6BEG[3] ,
    \Tile_X6Y1_W6BEG[2] ,
    \Tile_X6Y1_W6BEG[1] ,
    \Tile_X6Y1_W6BEG[0] }),
    .W6END({\Tile_X7Y1_W6BEG[11] ,
    \Tile_X7Y1_W6BEG[10] ,
    \Tile_X7Y1_W6BEG[9] ,
    \Tile_X7Y1_W6BEG[8] ,
    \Tile_X7Y1_W6BEG[7] ,
    \Tile_X7Y1_W6BEG[6] ,
    \Tile_X7Y1_W6BEG[5] ,
    \Tile_X7Y1_W6BEG[4] ,
    \Tile_X7Y1_W6BEG[3] ,
    \Tile_X7Y1_W6BEG[2] ,
    \Tile_X7Y1_W6BEG[1] ,
    \Tile_X7Y1_W6BEG[0] }),
    .WW4BEG({\Tile_X6Y1_WW4BEG[15] ,
    \Tile_X6Y1_WW4BEG[14] ,
    \Tile_X6Y1_WW4BEG[13] ,
    \Tile_X6Y1_WW4BEG[12] ,
    \Tile_X6Y1_WW4BEG[11] ,
    \Tile_X6Y1_WW4BEG[10] ,
    \Tile_X6Y1_WW4BEG[9] ,
    \Tile_X6Y1_WW4BEG[8] ,
    \Tile_X6Y1_WW4BEG[7] ,
    \Tile_X6Y1_WW4BEG[6] ,
    \Tile_X6Y1_WW4BEG[5] ,
    \Tile_X6Y1_WW4BEG[4] ,
    \Tile_X6Y1_WW4BEG[3] ,
    \Tile_X6Y1_WW4BEG[2] ,
    \Tile_X6Y1_WW4BEG[1] ,
    \Tile_X6Y1_WW4BEG[0] }),
    .WW4END({\Tile_X7Y1_WW4BEG[15] ,
    \Tile_X7Y1_WW4BEG[14] ,
    \Tile_X7Y1_WW4BEG[13] ,
    \Tile_X7Y1_WW4BEG[12] ,
    \Tile_X7Y1_WW4BEG[11] ,
    \Tile_X7Y1_WW4BEG[10] ,
    \Tile_X7Y1_WW4BEG[9] ,
    \Tile_X7Y1_WW4BEG[8] ,
    \Tile_X7Y1_WW4BEG[7] ,
    \Tile_X7Y1_WW4BEG[6] ,
    \Tile_X7Y1_WW4BEG[5] ,
    \Tile_X7Y1_WW4BEG[4] ,
    \Tile_X7Y1_WW4BEG[3] ,
    \Tile_X7Y1_WW4BEG[2] ,
    \Tile_X7Y1_WW4BEG[1] ,
    \Tile_X7Y1_WW4BEG[0] }));
 LUT4AB Tile_X6Y2_LUT4AB (.Ci(Tile_X6Y3_Co),
    .Co(Tile_X6Y2_Co),
    .UserCLK(Tile_X6Y3_UserCLKo),
    .UserCLKo(Tile_X6Y2_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X6Y2_E1BEG[3] ,
    \Tile_X6Y2_E1BEG[2] ,
    \Tile_X6Y2_E1BEG[1] ,
    \Tile_X6Y2_E1BEG[0] }),
    .E1END({\Tile_X5Y2_E1BEG[3] ,
    \Tile_X5Y2_E1BEG[2] ,
    \Tile_X5Y2_E1BEG[1] ,
    \Tile_X5Y2_E1BEG[0] }),
    .E2BEG({\Tile_X6Y2_E2BEG[7] ,
    \Tile_X6Y2_E2BEG[6] ,
    \Tile_X6Y2_E2BEG[5] ,
    \Tile_X6Y2_E2BEG[4] ,
    \Tile_X6Y2_E2BEG[3] ,
    \Tile_X6Y2_E2BEG[2] ,
    \Tile_X6Y2_E2BEG[1] ,
    \Tile_X6Y2_E2BEG[0] }),
    .E2BEGb({\Tile_X6Y2_E2BEGb[7] ,
    \Tile_X6Y2_E2BEGb[6] ,
    \Tile_X6Y2_E2BEGb[5] ,
    \Tile_X6Y2_E2BEGb[4] ,
    \Tile_X6Y2_E2BEGb[3] ,
    \Tile_X6Y2_E2BEGb[2] ,
    \Tile_X6Y2_E2BEGb[1] ,
    \Tile_X6Y2_E2BEGb[0] }),
    .E2END({\Tile_X5Y2_E2BEGb[7] ,
    \Tile_X5Y2_E2BEGb[6] ,
    \Tile_X5Y2_E2BEGb[5] ,
    \Tile_X5Y2_E2BEGb[4] ,
    \Tile_X5Y2_E2BEGb[3] ,
    \Tile_X5Y2_E2BEGb[2] ,
    \Tile_X5Y2_E2BEGb[1] ,
    \Tile_X5Y2_E2BEGb[0] }),
    .E2MID({\Tile_X5Y2_E2BEG[7] ,
    \Tile_X5Y2_E2BEG[6] ,
    \Tile_X5Y2_E2BEG[5] ,
    \Tile_X5Y2_E2BEG[4] ,
    \Tile_X5Y2_E2BEG[3] ,
    \Tile_X5Y2_E2BEG[2] ,
    \Tile_X5Y2_E2BEG[1] ,
    \Tile_X5Y2_E2BEG[0] }),
    .E6BEG({\Tile_X6Y2_E6BEG[11] ,
    \Tile_X6Y2_E6BEG[10] ,
    \Tile_X6Y2_E6BEG[9] ,
    \Tile_X6Y2_E6BEG[8] ,
    \Tile_X6Y2_E6BEG[7] ,
    \Tile_X6Y2_E6BEG[6] ,
    \Tile_X6Y2_E6BEG[5] ,
    \Tile_X6Y2_E6BEG[4] ,
    \Tile_X6Y2_E6BEG[3] ,
    \Tile_X6Y2_E6BEG[2] ,
    \Tile_X6Y2_E6BEG[1] ,
    \Tile_X6Y2_E6BEG[0] }),
    .E6END({\Tile_X5Y2_E6BEG[11] ,
    \Tile_X5Y2_E6BEG[10] ,
    \Tile_X5Y2_E6BEG[9] ,
    \Tile_X5Y2_E6BEG[8] ,
    \Tile_X5Y2_E6BEG[7] ,
    \Tile_X5Y2_E6BEG[6] ,
    \Tile_X5Y2_E6BEG[5] ,
    \Tile_X5Y2_E6BEG[4] ,
    \Tile_X5Y2_E6BEG[3] ,
    \Tile_X5Y2_E6BEG[2] ,
    \Tile_X5Y2_E6BEG[1] ,
    \Tile_X5Y2_E6BEG[0] }),
    .EE4BEG({\Tile_X6Y2_EE4BEG[15] ,
    \Tile_X6Y2_EE4BEG[14] ,
    \Tile_X6Y2_EE4BEG[13] ,
    \Tile_X6Y2_EE4BEG[12] ,
    \Tile_X6Y2_EE4BEG[11] ,
    \Tile_X6Y2_EE4BEG[10] ,
    \Tile_X6Y2_EE4BEG[9] ,
    \Tile_X6Y2_EE4BEG[8] ,
    \Tile_X6Y2_EE4BEG[7] ,
    \Tile_X6Y2_EE4BEG[6] ,
    \Tile_X6Y2_EE4BEG[5] ,
    \Tile_X6Y2_EE4BEG[4] ,
    \Tile_X6Y2_EE4BEG[3] ,
    \Tile_X6Y2_EE4BEG[2] ,
    \Tile_X6Y2_EE4BEG[1] ,
    \Tile_X6Y2_EE4BEG[0] }),
    .EE4END({\Tile_X5Y2_EE4BEG[15] ,
    \Tile_X5Y2_EE4BEG[14] ,
    \Tile_X5Y2_EE4BEG[13] ,
    \Tile_X5Y2_EE4BEG[12] ,
    \Tile_X5Y2_EE4BEG[11] ,
    \Tile_X5Y2_EE4BEG[10] ,
    \Tile_X5Y2_EE4BEG[9] ,
    \Tile_X5Y2_EE4BEG[8] ,
    \Tile_X5Y2_EE4BEG[7] ,
    \Tile_X5Y2_EE4BEG[6] ,
    \Tile_X5Y2_EE4BEG[5] ,
    \Tile_X5Y2_EE4BEG[4] ,
    \Tile_X5Y2_EE4BEG[3] ,
    \Tile_X5Y2_EE4BEG[2] ,
    \Tile_X5Y2_EE4BEG[1] ,
    \Tile_X5Y2_EE4BEG[0] }),
    .FrameData({\Tile_X5Y2_FrameData_O[31] ,
    \Tile_X5Y2_FrameData_O[30] ,
    \Tile_X5Y2_FrameData_O[29] ,
    \Tile_X5Y2_FrameData_O[28] ,
    \Tile_X5Y2_FrameData_O[27] ,
    \Tile_X5Y2_FrameData_O[26] ,
    \Tile_X5Y2_FrameData_O[25] ,
    \Tile_X5Y2_FrameData_O[24] ,
    \Tile_X5Y2_FrameData_O[23] ,
    \Tile_X5Y2_FrameData_O[22] ,
    \Tile_X5Y2_FrameData_O[21] ,
    \Tile_X5Y2_FrameData_O[20] ,
    \Tile_X5Y2_FrameData_O[19] ,
    \Tile_X5Y2_FrameData_O[18] ,
    \Tile_X5Y2_FrameData_O[17] ,
    \Tile_X5Y2_FrameData_O[16] ,
    \Tile_X5Y2_FrameData_O[15] ,
    \Tile_X5Y2_FrameData_O[14] ,
    \Tile_X5Y2_FrameData_O[13] ,
    \Tile_X5Y2_FrameData_O[12] ,
    \Tile_X5Y2_FrameData_O[11] ,
    \Tile_X5Y2_FrameData_O[10] ,
    \Tile_X5Y2_FrameData_O[9] ,
    \Tile_X5Y2_FrameData_O[8] ,
    \Tile_X5Y2_FrameData_O[7] ,
    \Tile_X5Y2_FrameData_O[6] ,
    \Tile_X5Y2_FrameData_O[5] ,
    \Tile_X5Y2_FrameData_O[4] ,
    \Tile_X5Y2_FrameData_O[3] ,
    \Tile_X5Y2_FrameData_O[2] ,
    \Tile_X5Y2_FrameData_O[1] ,
    \Tile_X5Y2_FrameData_O[0] }),
    .FrameData_O({\Tile_X6Y2_FrameData_O[31] ,
    \Tile_X6Y2_FrameData_O[30] ,
    \Tile_X6Y2_FrameData_O[29] ,
    \Tile_X6Y2_FrameData_O[28] ,
    \Tile_X6Y2_FrameData_O[27] ,
    \Tile_X6Y2_FrameData_O[26] ,
    \Tile_X6Y2_FrameData_O[25] ,
    \Tile_X6Y2_FrameData_O[24] ,
    \Tile_X6Y2_FrameData_O[23] ,
    \Tile_X6Y2_FrameData_O[22] ,
    \Tile_X6Y2_FrameData_O[21] ,
    \Tile_X6Y2_FrameData_O[20] ,
    \Tile_X6Y2_FrameData_O[19] ,
    \Tile_X6Y2_FrameData_O[18] ,
    \Tile_X6Y2_FrameData_O[17] ,
    \Tile_X6Y2_FrameData_O[16] ,
    \Tile_X6Y2_FrameData_O[15] ,
    \Tile_X6Y2_FrameData_O[14] ,
    \Tile_X6Y2_FrameData_O[13] ,
    \Tile_X6Y2_FrameData_O[12] ,
    \Tile_X6Y2_FrameData_O[11] ,
    \Tile_X6Y2_FrameData_O[10] ,
    \Tile_X6Y2_FrameData_O[9] ,
    \Tile_X6Y2_FrameData_O[8] ,
    \Tile_X6Y2_FrameData_O[7] ,
    \Tile_X6Y2_FrameData_O[6] ,
    \Tile_X6Y2_FrameData_O[5] ,
    \Tile_X6Y2_FrameData_O[4] ,
    \Tile_X6Y2_FrameData_O[3] ,
    \Tile_X6Y2_FrameData_O[2] ,
    \Tile_X6Y2_FrameData_O[1] ,
    \Tile_X6Y2_FrameData_O[0] }),
    .FrameStrobe({\Tile_X6Y3_FrameStrobe_O[19] ,
    \Tile_X6Y3_FrameStrobe_O[18] ,
    \Tile_X6Y3_FrameStrobe_O[17] ,
    \Tile_X6Y3_FrameStrobe_O[16] ,
    \Tile_X6Y3_FrameStrobe_O[15] ,
    \Tile_X6Y3_FrameStrobe_O[14] ,
    \Tile_X6Y3_FrameStrobe_O[13] ,
    \Tile_X6Y3_FrameStrobe_O[12] ,
    \Tile_X6Y3_FrameStrobe_O[11] ,
    \Tile_X6Y3_FrameStrobe_O[10] ,
    \Tile_X6Y3_FrameStrobe_O[9] ,
    \Tile_X6Y3_FrameStrobe_O[8] ,
    \Tile_X6Y3_FrameStrobe_O[7] ,
    \Tile_X6Y3_FrameStrobe_O[6] ,
    \Tile_X6Y3_FrameStrobe_O[5] ,
    \Tile_X6Y3_FrameStrobe_O[4] ,
    \Tile_X6Y3_FrameStrobe_O[3] ,
    \Tile_X6Y3_FrameStrobe_O[2] ,
    \Tile_X6Y3_FrameStrobe_O[1] ,
    \Tile_X6Y3_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X6Y2_FrameStrobe_O[19] ,
    \Tile_X6Y2_FrameStrobe_O[18] ,
    \Tile_X6Y2_FrameStrobe_O[17] ,
    \Tile_X6Y2_FrameStrobe_O[16] ,
    \Tile_X6Y2_FrameStrobe_O[15] ,
    \Tile_X6Y2_FrameStrobe_O[14] ,
    \Tile_X6Y2_FrameStrobe_O[13] ,
    \Tile_X6Y2_FrameStrobe_O[12] ,
    \Tile_X6Y2_FrameStrobe_O[11] ,
    \Tile_X6Y2_FrameStrobe_O[10] ,
    \Tile_X6Y2_FrameStrobe_O[9] ,
    \Tile_X6Y2_FrameStrobe_O[8] ,
    \Tile_X6Y2_FrameStrobe_O[7] ,
    \Tile_X6Y2_FrameStrobe_O[6] ,
    \Tile_X6Y2_FrameStrobe_O[5] ,
    \Tile_X6Y2_FrameStrobe_O[4] ,
    \Tile_X6Y2_FrameStrobe_O[3] ,
    \Tile_X6Y2_FrameStrobe_O[2] ,
    \Tile_X6Y2_FrameStrobe_O[1] ,
    \Tile_X6Y2_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X6Y2_N1BEG[3] ,
    \Tile_X6Y2_N1BEG[2] ,
    \Tile_X6Y2_N1BEG[1] ,
    \Tile_X6Y2_N1BEG[0] }),
    .N1END({\Tile_X6Y3_N1BEG[3] ,
    \Tile_X6Y3_N1BEG[2] ,
    \Tile_X6Y3_N1BEG[1] ,
    \Tile_X6Y3_N1BEG[0] }),
    .N2BEG({\Tile_X6Y2_N2BEG[7] ,
    \Tile_X6Y2_N2BEG[6] ,
    \Tile_X6Y2_N2BEG[5] ,
    \Tile_X6Y2_N2BEG[4] ,
    \Tile_X6Y2_N2BEG[3] ,
    \Tile_X6Y2_N2BEG[2] ,
    \Tile_X6Y2_N2BEG[1] ,
    \Tile_X6Y2_N2BEG[0] }),
    .N2BEGb({\Tile_X6Y2_N2BEGb[7] ,
    \Tile_X6Y2_N2BEGb[6] ,
    \Tile_X6Y2_N2BEGb[5] ,
    \Tile_X6Y2_N2BEGb[4] ,
    \Tile_X6Y2_N2BEGb[3] ,
    \Tile_X6Y2_N2BEGb[2] ,
    \Tile_X6Y2_N2BEGb[1] ,
    \Tile_X6Y2_N2BEGb[0] }),
    .N2END({\Tile_X6Y3_N2BEGb[7] ,
    \Tile_X6Y3_N2BEGb[6] ,
    \Tile_X6Y3_N2BEGb[5] ,
    \Tile_X6Y3_N2BEGb[4] ,
    \Tile_X6Y3_N2BEGb[3] ,
    \Tile_X6Y3_N2BEGb[2] ,
    \Tile_X6Y3_N2BEGb[1] ,
    \Tile_X6Y3_N2BEGb[0] }),
    .N2MID({\Tile_X6Y3_N2BEG[7] ,
    \Tile_X6Y3_N2BEG[6] ,
    \Tile_X6Y3_N2BEG[5] ,
    \Tile_X6Y3_N2BEG[4] ,
    \Tile_X6Y3_N2BEG[3] ,
    \Tile_X6Y3_N2BEG[2] ,
    \Tile_X6Y3_N2BEG[1] ,
    \Tile_X6Y3_N2BEG[0] }),
    .N4BEG({\Tile_X6Y2_N4BEG[15] ,
    \Tile_X6Y2_N4BEG[14] ,
    \Tile_X6Y2_N4BEG[13] ,
    \Tile_X6Y2_N4BEG[12] ,
    \Tile_X6Y2_N4BEG[11] ,
    \Tile_X6Y2_N4BEG[10] ,
    \Tile_X6Y2_N4BEG[9] ,
    \Tile_X6Y2_N4BEG[8] ,
    \Tile_X6Y2_N4BEG[7] ,
    \Tile_X6Y2_N4BEG[6] ,
    \Tile_X6Y2_N4BEG[5] ,
    \Tile_X6Y2_N4BEG[4] ,
    \Tile_X6Y2_N4BEG[3] ,
    \Tile_X6Y2_N4BEG[2] ,
    \Tile_X6Y2_N4BEG[1] ,
    \Tile_X6Y2_N4BEG[0] }),
    .N4END({\Tile_X6Y3_N4BEG[15] ,
    \Tile_X6Y3_N4BEG[14] ,
    \Tile_X6Y3_N4BEG[13] ,
    \Tile_X6Y3_N4BEG[12] ,
    \Tile_X6Y3_N4BEG[11] ,
    \Tile_X6Y3_N4BEG[10] ,
    \Tile_X6Y3_N4BEG[9] ,
    \Tile_X6Y3_N4BEG[8] ,
    \Tile_X6Y3_N4BEG[7] ,
    \Tile_X6Y3_N4BEG[6] ,
    \Tile_X6Y3_N4BEG[5] ,
    \Tile_X6Y3_N4BEG[4] ,
    \Tile_X6Y3_N4BEG[3] ,
    \Tile_X6Y3_N4BEG[2] ,
    \Tile_X6Y3_N4BEG[1] ,
    \Tile_X6Y3_N4BEG[0] }),
    .NN4BEG({\Tile_X6Y2_NN4BEG[15] ,
    \Tile_X6Y2_NN4BEG[14] ,
    \Tile_X6Y2_NN4BEG[13] ,
    \Tile_X6Y2_NN4BEG[12] ,
    \Tile_X6Y2_NN4BEG[11] ,
    \Tile_X6Y2_NN4BEG[10] ,
    \Tile_X6Y2_NN4BEG[9] ,
    \Tile_X6Y2_NN4BEG[8] ,
    \Tile_X6Y2_NN4BEG[7] ,
    \Tile_X6Y2_NN4BEG[6] ,
    \Tile_X6Y2_NN4BEG[5] ,
    \Tile_X6Y2_NN4BEG[4] ,
    \Tile_X6Y2_NN4BEG[3] ,
    \Tile_X6Y2_NN4BEG[2] ,
    \Tile_X6Y2_NN4BEG[1] ,
    \Tile_X6Y2_NN4BEG[0] }),
    .NN4END({\Tile_X6Y3_NN4BEG[15] ,
    \Tile_X6Y3_NN4BEG[14] ,
    \Tile_X6Y3_NN4BEG[13] ,
    \Tile_X6Y3_NN4BEG[12] ,
    \Tile_X6Y3_NN4BEG[11] ,
    \Tile_X6Y3_NN4BEG[10] ,
    \Tile_X6Y3_NN4BEG[9] ,
    \Tile_X6Y3_NN4BEG[8] ,
    \Tile_X6Y3_NN4BEG[7] ,
    \Tile_X6Y3_NN4BEG[6] ,
    \Tile_X6Y3_NN4BEG[5] ,
    \Tile_X6Y3_NN4BEG[4] ,
    \Tile_X6Y3_NN4BEG[3] ,
    \Tile_X6Y3_NN4BEG[2] ,
    \Tile_X6Y3_NN4BEG[1] ,
    \Tile_X6Y3_NN4BEG[0] }),
    .S1BEG({\Tile_X6Y2_S1BEG[3] ,
    \Tile_X6Y2_S1BEG[2] ,
    \Tile_X6Y2_S1BEG[1] ,
    \Tile_X6Y2_S1BEG[0] }),
    .S1END({\Tile_X6Y1_S1BEG[3] ,
    \Tile_X6Y1_S1BEG[2] ,
    \Tile_X6Y1_S1BEG[1] ,
    \Tile_X6Y1_S1BEG[0] }),
    .S2BEG({\Tile_X6Y2_S2BEG[7] ,
    \Tile_X6Y2_S2BEG[6] ,
    \Tile_X6Y2_S2BEG[5] ,
    \Tile_X6Y2_S2BEG[4] ,
    \Tile_X6Y2_S2BEG[3] ,
    \Tile_X6Y2_S2BEG[2] ,
    \Tile_X6Y2_S2BEG[1] ,
    \Tile_X6Y2_S2BEG[0] }),
    .S2BEGb({\Tile_X6Y2_S2BEGb[7] ,
    \Tile_X6Y2_S2BEGb[6] ,
    \Tile_X6Y2_S2BEGb[5] ,
    \Tile_X6Y2_S2BEGb[4] ,
    \Tile_X6Y2_S2BEGb[3] ,
    \Tile_X6Y2_S2BEGb[2] ,
    \Tile_X6Y2_S2BEGb[1] ,
    \Tile_X6Y2_S2BEGb[0] }),
    .S2END({\Tile_X6Y1_S2BEGb[7] ,
    \Tile_X6Y1_S2BEGb[6] ,
    \Tile_X6Y1_S2BEGb[5] ,
    \Tile_X6Y1_S2BEGb[4] ,
    \Tile_X6Y1_S2BEGb[3] ,
    \Tile_X6Y1_S2BEGb[2] ,
    \Tile_X6Y1_S2BEGb[1] ,
    \Tile_X6Y1_S2BEGb[0] }),
    .S2MID({\Tile_X6Y1_S2BEG[7] ,
    \Tile_X6Y1_S2BEG[6] ,
    \Tile_X6Y1_S2BEG[5] ,
    \Tile_X6Y1_S2BEG[4] ,
    \Tile_X6Y1_S2BEG[3] ,
    \Tile_X6Y1_S2BEG[2] ,
    \Tile_X6Y1_S2BEG[1] ,
    \Tile_X6Y1_S2BEG[0] }),
    .S4BEG({\Tile_X6Y2_S4BEG[15] ,
    \Tile_X6Y2_S4BEG[14] ,
    \Tile_X6Y2_S4BEG[13] ,
    \Tile_X6Y2_S4BEG[12] ,
    \Tile_X6Y2_S4BEG[11] ,
    \Tile_X6Y2_S4BEG[10] ,
    \Tile_X6Y2_S4BEG[9] ,
    \Tile_X6Y2_S4BEG[8] ,
    \Tile_X6Y2_S4BEG[7] ,
    \Tile_X6Y2_S4BEG[6] ,
    \Tile_X6Y2_S4BEG[5] ,
    \Tile_X6Y2_S4BEG[4] ,
    \Tile_X6Y2_S4BEG[3] ,
    \Tile_X6Y2_S4BEG[2] ,
    \Tile_X6Y2_S4BEG[1] ,
    \Tile_X6Y2_S4BEG[0] }),
    .S4END({\Tile_X6Y1_S4BEG[15] ,
    \Tile_X6Y1_S4BEG[14] ,
    \Tile_X6Y1_S4BEG[13] ,
    \Tile_X6Y1_S4BEG[12] ,
    \Tile_X6Y1_S4BEG[11] ,
    \Tile_X6Y1_S4BEG[10] ,
    \Tile_X6Y1_S4BEG[9] ,
    \Tile_X6Y1_S4BEG[8] ,
    \Tile_X6Y1_S4BEG[7] ,
    \Tile_X6Y1_S4BEG[6] ,
    \Tile_X6Y1_S4BEG[5] ,
    \Tile_X6Y1_S4BEG[4] ,
    \Tile_X6Y1_S4BEG[3] ,
    \Tile_X6Y1_S4BEG[2] ,
    \Tile_X6Y1_S4BEG[1] ,
    \Tile_X6Y1_S4BEG[0] }),
    .SS4BEG({\Tile_X6Y2_SS4BEG[15] ,
    \Tile_X6Y2_SS4BEG[14] ,
    \Tile_X6Y2_SS4BEG[13] ,
    \Tile_X6Y2_SS4BEG[12] ,
    \Tile_X6Y2_SS4BEG[11] ,
    \Tile_X6Y2_SS4BEG[10] ,
    \Tile_X6Y2_SS4BEG[9] ,
    \Tile_X6Y2_SS4BEG[8] ,
    \Tile_X6Y2_SS4BEG[7] ,
    \Tile_X6Y2_SS4BEG[6] ,
    \Tile_X6Y2_SS4BEG[5] ,
    \Tile_X6Y2_SS4BEG[4] ,
    \Tile_X6Y2_SS4BEG[3] ,
    \Tile_X6Y2_SS4BEG[2] ,
    \Tile_X6Y2_SS4BEG[1] ,
    \Tile_X6Y2_SS4BEG[0] }),
    .SS4END({\Tile_X6Y1_SS4BEG[15] ,
    \Tile_X6Y1_SS4BEG[14] ,
    \Tile_X6Y1_SS4BEG[13] ,
    \Tile_X6Y1_SS4BEG[12] ,
    \Tile_X6Y1_SS4BEG[11] ,
    \Tile_X6Y1_SS4BEG[10] ,
    \Tile_X6Y1_SS4BEG[9] ,
    \Tile_X6Y1_SS4BEG[8] ,
    \Tile_X6Y1_SS4BEG[7] ,
    \Tile_X6Y1_SS4BEG[6] ,
    \Tile_X6Y1_SS4BEG[5] ,
    \Tile_X6Y1_SS4BEG[4] ,
    \Tile_X6Y1_SS4BEG[3] ,
    \Tile_X6Y1_SS4BEG[2] ,
    \Tile_X6Y1_SS4BEG[1] ,
    \Tile_X6Y1_SS4BEG[0] }),
    .W1BEG({\Tile_X6Y2_W1BEG[3] ,
    \Tile_X6Y2_W1BEG[2] ,
    \Tile_X6Y2_W1BEG[1] ,
    \Tile_X6Y2_W1BEG[0] }),
    .W1END({\Tile_X7Y2_W1BEG[3] ,
    \Tile_X7Y2_W1BEG[2] ,
    \Tile_X7Y2_W1BEG[1] ,
    \Tile_X7Y2_W1BEG[0] }),
    .W2BEG({\Tile_X6Y2_W2BEG[7] ,
    \Tile_X6Y2_W2BEG[6] ,
    \Tile_X6Y2_W2BEG[5] ,
    \Tile_X6Y2_W2BEG[4] ,
    \Tile_X6Y2_W2BEG[3] ,
    \Tile_X6Y2_W2BEG[2] ,
    \Tile_X6Y2_W2BEG[1] ,
    \Tile_X6Y2_W2BEG[0] }),
    .W2BEGb({\Tile_X6Y2_W2BEGb[7] ,
    \Tile_X6Y2_W2BEGb[6] ,
    \Tile_X6Y2_W2BEGb[5] ,
    \Tile_X6Y2_W2BEGb[4] ,
    \Tile_X6Y2_W2BEGb[3] ,
    \Tile_X6Y2_W2BEGb[2] ,
    \Tile_X6Y2_W2BEGb[1] ,
    \Tile_X6Y2_W2BEGb[0] }),
    .W2END({\Tile_X7Y2_W2BEGb[7] ,
    \Tile_X7Y2_W2BEGb[6] ,
    \Tile_X7Y2_W2BEGb[5] ,
    \Tile_X7Y2_W2BEGb[4] ,
    \Tile_X7Y2_W2BEGb[3] ,
    \Tile_X7Y2_W2BEGb[2] ,
    \Tile_X7Y2_W2BEGb[1] ,
    \Tile_X7Y2_W2BEGb[0] }),
    .W2MID({\Tile_X7Y2_W2BEG[7] ,
    \Tile_X7Y2_W2BEG[6] ,
    \Tile_X7Y2_W2BEG[5] ,
    \Tile_X7Y2_W2BEG[4] ,
    \Tile_X7Y2_W2BEG[3] ,
    \Tile_X7Y2_W2BEG[2] ,
    \Tile_X7Y2_W2BEG[1] ,
    \Tile_X7Y2_W2BEG[0] }),
    .W6BEG({\Tile_X6Y2_W6BEG[11] ,
    \Tile_X6Y2_W6BEG[10] ,
    \Tile_X6Y2_W6BEG[9] ,
    \Tile_X6Y2_W6BEG[8] ,
    \Tile_X6Y2_W6BEG[7] ,
    \Tile_X6Y2_W6BEG[6] ,
    \Tile_X6Y2_W6BEG[5] ,
    \Tile_X6Y2_W6BEG[4] ,
    \Tile_X6Y2_W6BEG[3] ,
    \Tile_X6Y2_W6BEG[2] ,
    \Tile_X6Y2_W6BEG[1] ,
    \Tile_X6Y2_W6BEG[0] }),
    .W6END({\Tile_X7Y2_W6BEG[11] ,
    \Tile_X7Y2_W6BEG[10] ,
    \Tile_X7Y2_W6BEG[9] ,
    \Tile_X7Y2_W6BEG[8] ,
    \Tile_X7Y2_W6BEG[7] ,
    \Tile_X7Y2_W6BEG[6] ,
    \Tile_X7Y2_W6BEG[5] ,
    \Tile_X7Y2_W6BEG[4] ,
    \Tile_X7Y2_W6BEG[3] ,
    \Tile_X7Y2_W6BEG[2] ,
    \Tile_X7Y2_W6BEG[1] ,
    \Tile_X7Y2_W6BEG[0] }),
    .WW4BEG({\Tile_X6Y2_WW4BEG[15] ,
    \Tile_X6Y2_WW4BEG[14] ,
    \Tile_X6Y2_WW4BEG[13] ,
    \Tile_X6Y2_WW4BEG[12] ,
    \Tile_X6Y2_WW4BEG[11] ,
    \Tile_X6Y2_WW4BEG[10] ,
    \Tile_X6Y2_WW4BEG[9] ,
    \Tile_X6Y2_WW4BEG[8] ,
    \Tile_X6Y2_WW4BEG[7] ,
    \Tile_X6Y2_WW4BEG[6] ,
    \Tile_X6Y2_WW4BEG[5] ,
    \Tile_X6Y2_WW4BEG[4] ,
    \Tile_X6Y2_WW4BEG[3] ,
    \Tile_X6Y2_WW4BEG[2] ,
    \Tile_X6Y2_WW4BEG[1] ,
    \Tile_X6Y2_WW4BEG[0] }),
    .WW4END({\Tile_X7Y2_WW4BEG[15] ,
    \Tile_X7Y2_WW4BEG[14] ,
    \Tile_X7Y2_WW4BEG[13] ,
    \Tile_X7Y2_WW4BEG[12] ,
    \Tile_X7Y2_WW4BEG[11] ,
    \Tile_X7Y2_WW4BEG[10] ,
    \Tile_X7Y2_WW4BEG[9] ,
    \Tile_X7Y2_WW4BEG[8] ,
    \Tile_X7Y2_WW4BEG[7] ,
    \Tile_X7Y2_WW4BEG[6] ,
    \Tile_X7Y2_WW4BEG[5] ,
    \Tile_X7Y2_WW4BEG[4] ,
    \Tile_X7Y2_WW4BEG[3] ,
    \Tile_X7Y2_WW4BEG[2] ,
    \Tile_X7Y2_WW4BEG[1] ,
    \Tile_X7Y2_WW4BEG[0] }));
 LUT4AB Tile_X6Y3_LUT4AB (.Ci(Tile_X6Y4_Co),
    .Co(Tile_X6Y3_Co),
    .UserCLK(Tile_X6Y4_UserCLKo),
    .UserCLKo(Tile_X6Y3_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X6Y3_E1BEG[3] ,
    \Tile_X6Y3_E1BEG[2] ,
    \Tile_X6Y3_E1BEG[1] ,
    \Tile_X6Y3_E1BEG[0] }),
    .E1END({\Tile_X5Y3_E1BEG[3] ,
    \Tile_X5Y3_E1BEG[2] ,
    \Tile_X5Y3_E1BEG[1] ,
    \Tile_X5Y3_E1BEG[0] }),
    .E2BEG({\Tile_X6Y3_E2BEG[7] ,
    \Tile_X6Y3_E2BEG[6] ,
    \Tile_X6Y3_E2BEG[5] ,
    \Tile_X6Y3_E2BEG[4] ,
    \Tile_X6Y3_E2BEG[3] ,
    \Tile_X6Y3_E2BEG[2] ,
    \Tile_X6Y3_E2BEG[1] ,
    \Tile_X6Y3_E2BEG[0] }),
    .E2BEGb({\Tile_X6Y3_E2BEGb[7] ,
    \Tile_X6Y3_E2BEGb[6] ,
    \Tile_X6Y3_E2BEGb[5] ,
    \Tile_X6Y3_E2BEGb[4] ,
    \Tile_X6Y3_E2BEGb[3] ,
    \Tile_X6Y3_E2BEGb[2] ,
    \Tile_X6Y3_E2BEGb[1] ,
    \Tile_X6Y3_E2BEGb[0] }),
    .E2END({\Tile_X5Y3_E2BEGb[7] ,
    \Tile_X5Y3_E2BEGb[6] ,
    \Tile_X5Y3_E2BEGb[5] ,
    \Tile_X5Y3_E2BEGb[4] ,
    \Tile_X5Y3_E2BEGb[3] ,
    \Tile_X5Y3_E2BEGb[2] ,
    \Tile_X5Y3_E2BEGb[1] ,
    \Tile_X5Y3_E2BEGb[0] }),
    .E2MID({\Tile_X5Y3_E2BEG[7] ,
    \Tile_X5Y3_E2BEG[6] ,
    \Tile_X5Y3_E2BEG[5] ,
    \Tile_X5Y3_E2BEG[4] ,
    \Tile_X5Y3_E2BEG[3] ,
    \Tile_X5Y3_E2BEG[2] ,
    \Tile_X5Y3_E2BEG[1] ,
    \Tile_X5Y3_E2BEG[0] }),
    .E6BEG({\Tile_X6Y3_E6BEG[11] ,
    \Tile_X6Y3_E6BEG[10] ,
    \Tile_X6Y3_E6BEG[9] ,
    \Tile_X6Y3_E6BEG[8] ,
    \Tile_X6Y3_E6BEG[7] ,
    \Tile_X6Y3_E6BEG[6] ,
    \Tile_X6Y3_E6BEG[5] ,
    \Tile_X6Y3_E6BEG[4] ,
    \Tile_X6Y3_E6BEG[3] ,
    \Tile_X6Y3_E6BEG[2] ,
    \Tile_X6Y3_E6BEG[1] ,
    \Tile_X6Y3_E6BEG[0] }),
    .E6END({\Tile_X5Y3_E6BEG[11] ,
    \Tile_X5Y3_E6BEG[10] ,
    \Tile_X5Y3_E6BEG[9] ,
    \Tile_X5Y3_E6BEG[8] ,
    \Tile_X5Y3_E6BEG[7] ,
    \Tile_X5Y3_E6BEG[6] ,
    \Tile_X5Y3_E6BEG[5] ,
    \Tile_X5Y3_E6BEG[4] ,
    \Tile_X5Y3_E6BEG[3] ,
    \Tile_X5Y3_E6BEG[2] ,
    \Tile_X5Y3_E6BEG[1] ,
    \Tile_X5Y3_E6BEG[0] }),
    .EE4BEG({\Tile_X6Y3_EE4BEG[15] ,
    \Tile_X6Y3_EE4BEG[14] ,
    \Tile_X6Y3_EE4BEG[13] ,
    \Tile_X6Y3_EE4BEG[12] ,
    \Tile_X6Y3_EE4BEG[11] ,
    \Tile_X6Y3_EE4BEG[10] ,
    \Tile_X6Y3_EE4BEG[9] ,
    \Tile_X6Y3_EE4BEG[8] ,
    \Tile_X6Y3_EE4BEG[7] ,
    \Tile_X6Y3_EE4BEG[6] ,
    \Tile_X6Y3_EE4BEG[5] ,
    \Tile_X6Y3_EE4BEG[4] ,
    \Tile_X6Y3_EE4BEG[3] ,
    \Tile_X6Y3_EE4BEG[2] ,
    \Tile_X6Y3_EE4BEG[1] ,
    \Tile_X6Y3_EE4BEG[0] }),
    .EE4END({\Tile_X5Y3_EE4BEG[15] ,
    \Tile_X5Y3_EE4BEG[14] ,
    \Tile_X5Y3_EE4BEG[13] ,
    \Tile_X5Y3_EE4BEG[12] ,
    \Tile_X5Y3_EE4BEG[11] ,
    \Tile_X5Y3_EE4BEG[10] ,
    \Tile_X5Y3_EE4BEG[9] ,
    \Tile_X5Y3_EE4BEG[8] ,
    \Tile_X5Y3_EE4BEG[7] ,
    \Tile_X5Y3_EE4BEG[6] ,
    \Tile_X5Y3_EE4BEG[5] ,
    \Tile_X5Y3_EE4BEG[4] ,
    \Tile_X5Y3_EE4BEG[3] ,
    \Tile_X5Y3_EE4BEG[2] ,
    \Tile_X5Y3_EE4BEG[1] ,
    \Tile_X5Y3_EE4BEG[0] }),
    .FrameData({\Tile_X5Y3_FrameData_O[31] ,
    \Tile_X5Y3_FrameData_O[30] ,
    \Tile_X5Y3_FrameData_O[29] ,
    \Tile_X5Y3_FrameData_O[28] ,
    \Tile_X5Y3_FrameData_O[27] ,
    \Tile_X5Y3_FrameData_O[26] ,
    \Tile_X5Y3_FrameData_O[25] ,
    \Tile_X5Y3_FrameData_O[24] ,
    \Tile_X5Y3_FrameData_O[23] ,
    \Tile_X5Y3_FrameData_O[22] ,
    \Tile_X5Y3_FrameData_O[21] ,
    \Tile_X5Y3_FrameData_O[20] ,
    \Tile_X5Y3_FrameData_O[19] ,
    \Tile_X5Y3_FrameData_O[18] ,
    \Tile_X5Y3_FrameData_O[17] ,
    \Tile_X5Y3_FrameData_O[16] ,
    \Tile_X5Y3_FrameData_O[15] ,
    \Tile_X5Y3_FrameData_O[14] ,
    \Tile_X5Y3_FrameData_O[13] ,
    \Tile_X5Y3_FrameData_O[12] ,
    \Tile_X5Y3_FrameData_O[11] ,
    \Tile_X5Y3_FrameData_O[10] ,
    \Tile_X5Y3_FrameData_O[9] ,
    \Tile_X5Y3_FrameData_O[8] ,
    \Tile_X5Y3_FrameData_O[7] ,
    \Tile_X5Y3_FrameData_O[6] ,
    \Tile_X5Y3_FrameData_O[5] ,
    \Tile_X5Y3_FrameData_O[4] ,
    \Tile_X5Y3_FrameData_O[3] ,
    \Tile_X5Y3_FrameData_O[2] ,
    \Tile_X5Y3_FrameData_O[1] ,
    \Tile_X5Y3_FrameData_O[0] }),
    .FrameData_O({\Tile_X6Y3_FrameData_O[31] ,
    \Tile_X6Y3_FrameData_O[30] ,
    \Tile_X6Y3_FrameData_O[29] ,
    \Tile_X6Y3_FrameData_O[28] ,
    \Tile_X6Y3_FrameData_O[27] ,
    \Tile_X6Y3_FrameData_O[26] ,
    \Tile_X6Y3_FrameData_O[25] ,
    \Tile_X6Y3_FrameData_O[24] ,
    \Tile_X6Y3_FrameData_O[23] ,
    \Tile_X6Y3_FrameData_O[22] ,
    \Tile_X6Y3_FrameData_O[21] ,
    \Tile_X6Y3_FrameData_O[20] ,
    \Tile_X6Y3_FrameData_O[19] ,
    \Tile_X6Y3_FrameData_O[18] ,
    \Tile_X6Y3_FrameData_O[17] ,
    \Tile_X6Y3_FrameData_O[16] ,
    \Tile_X6Y3_FrameData_O[15] ,
    \Tile_X6Y3_FrameData_O[14] ,
    \Tile_X6Y3_FrameData_O[13] ,
    \Tile_X6Y3_FrameData_O[12] ,
    \Tile_X6Y3_FrameData_O[11] ,
    \Tile_X6Y3_FrameData_O[10] ,
    \Tile_X6Y3_FrameData_O[9] ,
    \Tile_X6Y3_FrameData_O[8] ,
    \Tile_X6Y3_FrameData_O[7] ,
    \Tile_X6Y3_FrameData_O[6] ,
    \Tile_X6Y3_FrameData_O[5] ,
    \Tile_X6Y3_FrameData_O[4] ,
    \Tile_X6Y3_FrameData_O[3] ,
    \Tile_X6Y3_FrameData_O[2] ,
    \Tile_X6Y3_FrameData_O[1] ,
    \Tile_X6Y3_FrameData_O[0] }),
    .FrameStrobe({\Tile_X6Y4_FrameStrobe_O[19] ,
    \Tile_X6Y4_FrameStrobe_O[18] ,
    \Tile_X6Y4_FrameStrobe_O[17] ,
    \Tile_X6Y4_FrameStrobe_O[16] ,
    \Tile_X6Y4_FrameStrobe_O[15] ,
    \Tile_X6Y4_FrameStrobe_O[14] ,
    \Tile_X6Y4_FrameStrobe_O[13] ,
    \Tile_X6Y4_FrameStrobe_O[12] ,
    \Tile_X6Y4_FrameStrobe_O[11] ,
    \Tile_X6Y4_FrameStrobe_O[10] ,
    \Tile_X6Y4_FrameStrobe_O[9] ,
    \Tile_X6Y4_FrameStrobe_O[8] ,
    \Tile_X6Y4_FrameStrobe_O[7] ,
    \Tile_X6Y4_FrameStrobe_O[6] ,
    \Tile_X6Y4_FrameStrobe_O[5] ,
    \Tile_X6Y4_FrameStrobe_O[4] ,
    \Tile_X6Y4_FrameStrobe_O[3] ,
    \Tile_X6Y4_FrameStrobe_O[2] ,
    \Tile_X6Y4_FrameStrobe_O[1] ,
    \Tile_X6Y4_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X6Y3_FrameStrobe_O[19] ,
    \Tile_X6Y3_FrameStrobe_O[18] ,
    \Tile_X6Y3_FrameStrobe_O[17] ,
    \Tile_X6Y3_FrameStrobe_O[16] ,
    \Tile_X6Y3_FrameStrobe_O[15] ,
    \Tile_X6Y3_FrameStrobe_O[14] ,
    \Tile_X6Y3_FrameStrobe_O[13] ,
    \Tile_X6Y3_FrameStrobe_O[12] ,
    \Tile_X6Y3_FrameStrobe_O[11] ,
    \Tile_X6Y3_FrameStrobe_O[10] ,
    \Tile_X6Y3_FrameStrobe_O[9] ,
    \Tile_X6Y3_FrameStrobe_O[8] ,
    \Tile_X6Y3_FrameStrobe_O[7] ,
    \Tile_X6Y3_FrameStrobe_O[6] ,
    \Tile_X6Y3_FrameStrobe_O[5] ,
    \Tile_X6Y3_FrameStrobe_O[4] ,
    \Tile_X6Y3_FrameStrobe_O[3] ,
    \Tile_X6Y3_FrameStrobe_O[2] ,
    \Tile_X6Y3_FrameStrobe_O[1] ,
    \Tile_X6Y3_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X6Y3_N1BEG[3] ,
    \Tile_X6Y3_N1BEG[2] ,
    \Tile_X6Y3_N1BEG[1] ,
    \Tile_X6Y3_N1BEG[0] }),
    .N1END({\Tile_X6Y4_N1BEG[3] ,
    \Tile_X6Y4_N1BEG[2] ,
    \Tile_X6Y4_N1BEG[1] ,
    \Tile_X6Y4_N1BEG[0] }),
    .N2BEG({\Tile_X6Y3_N2BEG[7] ,
    \Tile_X6Y3_N2BEG[6] ,
    \Tile_X6Y3_N2BEG[5] ,
    \Tile_X6Y3_N2BEG[4] ,
    \Tile_X6Y3_N2BEG[3] ,
    \Tile_X6Y3_N2BEG[2] ,
    \Tile_X6Y3_N2BEG[1] ,
    \Tile_X6Y3_N2BEG[0] }),
    .N2BEGb({\Tile_X6Y3_N2BEGb[7] ,
    \Tile_X6Y3_N2BEGb[6] ,
    \Tile_X6Y3_N2BEGb[5] ,
    \Tile_X6Y3_N2BEGb[4] ,
    \Tile_X6Y3_N2BEGb[3] ,
    \Tile_X6Y3_N2BEGb[2] ,
    \Tile_X6Y3_N2BEGb[1] ,
    \Tile_X6Y3_N2BEGb[0] }),
    .N2END({\Tile_X6Y4_N2BEGb[7] ,
    \Tile_X6Y4_N2BEGb[6] ,
    \Tile_X6Y4_N2BEGb[5] ,
    \Tile_X6Y4_N2BEGb[4] ,
    \Tile_X6Y4_N2BEGb[3] ,
    \Tile_X6Y4_N2BEGb[2] ,
    \Tile_X6Y4_N2BEGb[1] ,
    \Tile_X6Y4_N2BEGb[0] }),
    .N2MID({\Tile_X6Y4_N2BEG[7] ,
    \Tile_X6Y4_N2BEG[6] ,
    \Tile_X6Y4_N2BEG[5] ,
    \Tile_X6Y4_N2BEG[4] ,
    \Tile_X6Y4_N2BEG[3] ,
    \Tile_X6Y4_N2BEG[2] ,
    \Tile_X6Y4_N2BEG[1] ,
    \Tile_X6Y4_N2BEG[0] }),
    .N4BEG({\Tile_X6Y3_N4BEG[15] ,
    \Tile_X6Y3_N4BEG[14] ,
    \Tile_X6Y3_N4BEG[13] ,
    \Tile_X6Y3_N4BEG[12] ,
    \Tile_X6Y3_N4BEG[11] ,
    \Tile_X6Y3_N4BEG[10] ,
    \Tile_X6Y3_N4BEG[9] ,
    \Tile_X6Y3_N4BEG[8] ,
    \Tile_X6Y3_N4BEG[7] ,
    \Tile_X6Y3_N4BEG[6] ,
    \Tile_X6Y3_N4BEG[5] ,
    \Tile_X6Y3_N4BEG[4] ,
    \Tile_X6Y3_N4BEG[3] ,
    \Tile_X6Y3_N4BEG[2] ,
    \Tile_X6Y3_N4BEG[1] ,
    \Tile_X6Y3_N4BEG[0] }),
    .N4END({\Tile_X6Y4_N4BEG[15] ,
    \Tile_X6Y4_N4BEG[14] ,
    \Tile_X6Y4_N4BEG[13] ,
    \Tile_X6Y4_N4BEG[12] ,
    \Tile_X6Y4_N4BEG[11] ,
    \Tile_X6Y4_N4BEG[10] ,
    \Tile_X6Y4_N4BEG[9] ,
    \Tile_X6Y4_N4BEG[8] ,
    \Tile_X6Y4_N4BEG[7] ,
    \Tile_X6Y4_N4BEG[6] ,
    \Tile_X6Y4_N4BEG[5] ,
    \Tile_X6Y4_N4BEG[4] ,
    \Tile_X6Y4_N4BEG[3] ,
    \Tile_X6Y4_N4BEG[2] ,
    \Tile_X6Y4_N4BEG[1] ,
    \Tile_X6Y4_N4BEG[0] }),
    .NN4BEG({\Tile_X6Y3_NN4BEG[15] ,
    \Tile_X6Y3_NN4BEG[14] ,
    \Tile_X6Y3_NN4BEG[13] ,
    \Tile_X6Y3_NN4BEG[12] ,
    \Tile_X6Y3_NN4BEG[11] ,
    \Tile_X6Y3_NN4BEG[10] ,
    \Tile_X6Y3_NN4BEG[9] ,
    \Tile_X6Y3_NN4BEG[8] ,
    \Tile_X6Y3_NN4BEG[7] ,
    \Tile_X6Y3_NN4BEG[6] ,
    \Tile_X6Y3_NN4BEG[5] ,
    \Tile_X6Y3_NN4BEG[4] ,
    \Tile_X6Y3_NN4BEG[3] ,
    \Tile_X6Y3_NN4BEG[2] ,
    \Tile_X6Y3_NN4BEG[1] ,
    \Tile_X6Y3_NN4BEG[0] }),
    .NN4END({\Tile_X6Y4_NN4BEG[15] ,
    \Tile_X6Y4_NN4BEG[14] ,
    \Tile_X6Y4_NN4BEG[13] ,
    \Tile_X6Y4_NN4BEG[12] ,
    \Tile_X6Y4_NN4BEG[11] ,
    \Tile_X6Y4_NN4BEG[10] ,
    \Tile_X6Y4_NN4BEG[9] ,
    \Tile_X6Y4_NN4BEG[8] ,
    \Tile_X6Y4_NN4BEG[7] ,
    \Tile_X6Y4_NN4BEG[6] ,
    \Tile_X6Y4_NN4BEG[5] ,
    \Tile_X6Y4_NN4BEG[4] ,
    \Tile_X6Y4_NN4BEG[3] ,
    \Tile_X6Y4_NN4BEG[2] ,
    \Tile_X6Y4_NN4BEG[1] ,
    \Tile_X6Y4_NN4BEG[0] }),
    .S1BEG({\Tile_X6Y3_S1BEG[3] ,
    \Tile_X6Y3_S1BEG[2] ,
    \Tile_X6Y3_S1BEG[1] ,
    \Tile_X6Y3_S1BEG[0] }),
    .S1END({\Tile_X6Y2_S1BEG[3] ,
    \Tile_X6Y2_S1BEG[2] ,
    \Tile_X6Y2_S1BEG[1] ,
    \Tile_X6Y2_S1BEG[0] }),
    .S2BEG({\Tile_X6Y3_S2BEG[7] ,
    \Tile_X6Y3_S2BEG[6] ,
    \Tile_X6Y3_S2BEG[5] ,
    \Tile_X6Y3_S2BEG[4] ,
    \Tile_X6Y3_S2BEG[3] ,
    \Tile_X6Y3_S2BEG[2] ,
    \Tile_X6Y3_S2BEG[1] ,
    \Tile_X6Y3_S2BEG[0] }),
    .S2BEGb({\Tile_X6Y3_S2BEGb[7] ,
    \Tile_X6Y3_S2BEGb[6] ,
    \Tile_X6Y3_S2BEGb[5] ,
    \Tile_X6Y3_S2BEGb[4] ,
    \Tile_X6Y3_S2BEGb[3] ,
    \Tile_X6Y3_S2BEGb[2] ,
    \Tile_X6Y3_S2BEGb[1] ,
    \Tile_X6Y3_S2BEGb[0] }),
    .S2END({\Tile_X6Y2_S2BEGb[7] ,
    \Tile_X6Y2_S2BEGb[6] ,
    \Tile_X6Y2_S2BEGb[5] ,
    \Tile_X6Y2_S2BEGb[4] ,
    \Tile_X6Y2_S2BEGb[3] ,
    \Tile_X6Y2_S2BEGb[2] ,
    \Tile_X6Y2_S2BEGb[1] ,
    \Tile_X6Y2_S2BEGb[0] }),
    .S2MID({\Tile_X6Y2_S2BEG[7] ,
    \Tile_X6Y2_S2BEG[6] ,
    \Tile_X6Y2_S2BEG[5] ,
    \Tile_X6Y2_S2BEG[4] ,
    \Tile_X6Y2_S2BEG[3] ,
    \Tile_X6Y2_S2BEG[2] ,
    \Tile_X6Y2_S2BEG[1] ,
    \Tile_X6Y2_S2BEG[0] }),
    .S4BEG({\Tile_X6Y3_S4BEG[15] ,
    \Tile_X6Y3_S4BEG[14] ,
    \Tile_X6Y3_S4BEG[13] ,
    \Tile_X6Y3_S4BEG[12] ,
    \Tile_X6Y3_S4BEG[11] ,
    \Tile_X6Y3_S4BEG[10] ,
    \Tile_X6Y3_S4BEG[9] ,
    \Tile_X6Y3_S4BEG[8] ,
    \Tile_X6Y3_S4BEG[7] ,
    \Tile_X6Y3_S4BEG[6] ,
    \Tile_X6Y3_S4BEG[5] ,
    \Tile_X6Y3_S4BEG[4] ,
    \Tile_X6Y3_S4BEG[3] ,
    \Tile_X6Y3_S4BEG[2] ,
    \Tile_X6Y3_S4BEG[1] ,
    \Tile_X6Y3_S4BEG[0] }),
    .S4END({\Tile_X6Y2_S4BEG[15] ,
    \Tile_X6Y2_S4BEG[14] ,
    \Tile_X6Y2_S4BEG[13] ,
    \Tile_X6Y2_S4BEG[12] ,
    \Tile_X6Y2_S4BEG[11] ,
    \Tile_X6Y2_S4BEG[10] ,
    \Tile_X6Y2_S4BEG[9] ,
    \Tile_X6Y2_S4BEG[8] ,
    \Tile_X6Y2_S4BEG[7] ,
    \Tile_X6Y2_S4BEG[6] ,
    \Tile_X6Y2_S4BEG[5] ,
    \Tile_X6Y2_S4BEG[4] ,
    \Tile_X6Y2_S4BEG[3] ,
    \Tile_X6Y2_S4BEG[2] ,
    \Tile_X6Y2_S4BEG[1] ,
    \Tile_X6Y2_S4BEG[0] }),
    .SS4BEG({\Tile_X6Y3_SS4BEG[15] ,
    \Tile_X6Y3_SS4BEG[14] ,
    \Tile_X6Y3_SS4BEG[13] ,
    \Tile_X6Y3_SS4BEG[12] ,
    \Tile_X6Y3_SS4BEG[11] ,
    \Tile_X6Y3_SS4BEG[10] ,
    \Tile_X6Y3_SS4BEG[9] ,
    \Tile_X6Y3_SS4BEG[8] ,
    \Tile_X6Y3_SS4BEG[7] ,
    \Tile_X6Y3_SS4BEG[6] ,
    \Tile_X6Y3_SS4BEG[5] ,
    \Tile_X6Y3_SS4BEG[4] ,
    \Tile_X6Y3_SS4BEG[3] ,
    \Tile_X6Y3_SS4BEG[2] ,
    \Tile_X6Y3_SS4BEG[1] ,
    \Tile_X6Y3_SS4BEG[0] }),
    .SS4END({\Tile_X6Y2_SS4BEG[15] ,
    \Tile_X6Y2_SS4BEG[14] ,
    \Tile_X6Y2_SS4BEG[13] ,
    \Tile_X6Y2_SS4BEG[12] ,
    \Tile_X6Y2_SS4BEG[11] ,
    \Tile_X6Y2_SS4BEG[10] ,
    \Tile_X6Y2_SS4BEG[9] ,
    \Tile_X6Y2_SS4BEG[8] ,
    \Tile_X6Y2_SS4BEG[7] ,
    \Tile_X6Y2_SS4BEG[6] ,
    \Tile_X6Y2_SS4BEG[5] ,
    \Tile_X6Y2_SS4BEG[4] ,
    \Tile_X6Y2_SS4BEG[3] ,
    \Tile_X6Y2_SS4BEG[2] ,
    \Tile_X6Y2_SS4BEG[1] ,
    \Tile_X6Y2_SS4BEG[0] }),
    .W1BEG({\Tile_X6Y3_W1BEG[3] ,
    \Tile_X6Y3_W1BEG[2] ,
    \Tile_X6Y3_W1BEG[1] ,
    \Tile_X6Y3_W1BEG[0] }),
    .W1END({\Tile_X7Y3_W1BEG[3] ,
    \Tile_X7Y3_W1BEG[2] ,
    \Tile_X7Y3_W1BEG[1] ,
    \Tile_X7Y3_W1BEG[0] }),
    .W2BEG({\Tile_X6Y3_W2BEG[7] ,
    \Tile_X6Y3_W2BEG[6] ,
    \Tile_X6Y3_W2BEG[5] ,
    \Tile_X6Y3_W2BEG[4] ,
    \Tile_X6Y3_W2BEG[3] ,
    \Tile_X6Y3_W2BEG[2] ,
    \Tile_X6Y3_W2BEG[1] ,
    \Tile_X6Y3_W2BEG[0] }),
    .W2BEGb({\Tile_X6Y3_W2BEGb[7] ,
    \Tile_X6Y3_W2BEGb[6] ,
    \Tile_X6Y3_W2BEGb[5] ,
    \Tile_X6Y3_W2BEGb[4] ,
    \Tile_X6Y3_W2BEGb[3] ,
    \Tile_X6Y3_W2BEGb[2] ,
    \Tile_X6Y3_W2BEGb[1] ,
    \Tile_X6Y3_W2BEGb[0] }),
    .W2END({\Tile_X7Y3_W2BEGb[7] ,
    \Tile_X7Y3_W2BEGb[6] ,
    \Tile_X7Y3_W2BEGb[5] ,
    \Tile_X7Y3_W2BEGb[4] ,
    \Tile_X7Y3_W2BEGb[3] ,
    \Tile_X7Y3_W2BEGb[2] ,
    \Tile_X7Y3_W2BEGb[1] ,
    \Tile_X7Y3_W2BEGb[0] }),
    .W2MID({\Tile_X7Y3_W2BEG[7] ,
    \Tile_X7Y3_W2BEG[6] ,
    \Tile_X7Y3_W2BEG[5] ,
    \Tile_X7Y3_W2BEG[4] ,
    \Tile_X7Y3_W2BEG[3] ,
    \Tile_X7Y3_W2BEG[2] ,
    \Tile_X7Y3_W2BEG[1] ,
    \Tile_X7Y3_W2BEG[0] }),
    .W6BEG({\Tile_X6Y3_W6BEG[11] ,
    \Tile_X6Y3_W6BEG[10] ,
    \Tile_X6Y3_W6BEG[9] ,
    \Tile_X6Y3_W6BEG[8] ,
    \Tile_X6Y3_W6BEG[7] ,
    \Tile_X6Y3_W6BEG[6] ,
    \Tile_X6Y3_W6BEG[5] ,
    \Tile_X6Y3_W6BEG[4] ,
    \Tile_X6Y3_W6BEG[3] ,
    \Tile_X6Y3_W6BEG[2] ,
    \Tile_X6Y3_W6BEG[1] ,
    \Tile_X6Y3_W6BEG[0] }),
    .W6END({\Tile_X7Y3_W6BEG[11] ,
    \Tile_X7Y3_W6BEG[10] ,
    \Tile_X7Y3_W6BEG[9] ,
    \Tile_X7Y3_W6BEG[8] ,
    \Tile_X7Y3_W6BEG[7] ,
    \Tile_X7Y3_W6BEG[6] ,
    \Tile_X7Y3_W6BEG[5] ,
    \Tile_X7Y3_W6BEG[4] ,
    \Tile_X7Y3_W6BEG[3] ,
    \Tile_X7Y3_W6BEG[2] ,
    \Tile_X7Y3_W6BEG[1] ,
    \Tile_X7Y3_W6BEG[0] }),
    .WW4BEG({\Tile_X6Y3_WW4BEG[15] ,
    \Tile_X6Y3_WW4BEG[14] ,
    \Tile_X6Y3_WW4BEG[13] ,
    \Tile_X6Y3_WW4BEG[12] ,
    \Tile_X6Y3_WW4BEG[11] ,
    \Tile_X6Y3_WW4BEG[10] ,
    \Tile_X6Y3_WW4BEG[9] ,
    \Tile_X6Y3_WW4BEG[8] ,
    \Tile_X6Y3_WW4BEG[7] ,
    \Tile_X6Y3_WW4BEG[6] ,
    \Tile_X6Y3_WW4BEG[5] ,
    \Tile_X6Y3_WW4BEG[4] ,
    \Tile_X6Y3_WW4BEG[3] ,
    \Tile_X6Y3_WW4BEG[2] ,
    \Tile_X6Y3_WW4BEG[1] ,
    \Tile_X6Y3_WW4BEG[0] }),
    .WW4END({\Tile_X7Y3_WW4BEG[15] ,
    \Tile_X7Y3_WW4BEG[14] ,
    \Tile_X7Y3_WW4BEG[13] ,
    \Tile_X7Y3_WW4BEG[12] ,
    \Tile_X7Y3_WW4BEG[11] ,
    \Tile_X7Y3_WW4BEG[10] ,
    \Tile_X7Y3_WW4BEG[9] ,
    \Tile_X7Y3_WW4BEG[8] ,
    \Tile_X7Y3_WW4BEG[7] ,
    \Tile_X7Y3_WW4BEG[6] ,
    \Tile_X7Y3_WW4BEG[5] ,
    \Tile_X7Y3_WW4BEG[4] ,
    \Tile_X7Y3_WW4BEG[3] ,
    \Tile_X7Y3_WW4BEG[2] ,
    \Tile_X7Y3_WW4BEG[1] ,
    \Tile_X7Y3_WW4BEG[0] }));
 LUT4AB Tile_X6Y4_LUT4AB (.Ci(Tile_X6Y5_Co),
    .Co(Tile_X6Y4_Co),
    .UserCLK(Tile_X6Y5_UserCLKo),
    .UserCLKo(Tile_X6Y4_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X6Y4_E1BEG[3] ,
    \Tile_X6Y4_E1BEG[2] ,
    \Tile_X6Y4_E1BEG[1] ,
    \Tile_X6Y4_E1BEG[0] }),
    .E1END({\Tile_X5Y4_E1BEG[3] ,
    \Tile_X5Y4_E1BEG[2] ,
    \Tile_X5Y4_E1BEG[1] ,
    \Tile_X5Y4_E1BEG[0] }),
    .E2BEG({\Tile_X6Y4_E2BEG[7] ,
    \Tile_X6Y4_E2BEG[6] ,
    \Tile_X6Y4_E2BEG[5] ,
    \Tile_X6Y4_E2BEG[4] ,
    \Tile_X6Y4_E2BEG[3] ,
    \Tile_X6Y4_E2BEG[2] ,
    \Tile_X6Y4_E2BEG[1] ,
    \Tile_X6Y4_E2BEG[0] }),
    .E2BEGb({\Tile_X6Y4_E2BEGb[7] ,
    \Tile_X6Y4_E2BEGb[6] ,
    \Tile_X6Y4_E2BEGb[5] ,
    \Tile_X6Y4_E2BEGb[4] ,
    \Tile_X6Y4_E2BEGb[3] ,
    \Tile_X6Y4_E2BEGb[2] ,
    \Tile_X6Y4_E2BEGb[1] ,
    \Tile_X6Y4_E2BEGb[0] }),
    .E2END({\Tile_X5Y4_E2BEGb[7] ,
    \Tile_X5Y4_E2BEGb[6] ,
    \Tile_X5Y4_E2BEGb[5] ,
    \Tile_X5Y4_E2BEGb[4] ,
    \Tile_X5Y4_E2BEGb[3] ,
    \Tile_X5Y4_E2BEGb[2] ,
    \Tile_X5Y4_E2BEGb[1] ,
    \Tile_X5Y4_E2BEGb[0] }),
    .E2MID({\Tile_X5Y4_E2BEG[7] ,
    \Tile_X5Y4_E2BEG[6] ,
    \Tile_X5Y4_E2BEG[5] ,
    \Tile_X5Y4_E2BEG[4] ,
    \Tile_X5Y4_E2BEG[3] ,
    \Tile_X5Y4_E2BEG[2] ,
    \Tile_X5Y4_E2BEG[1] ,
    \Tile_X5Y4_E2BEG[0] }),
    .E6BEG({\Tile_X6Y4_E6BEG[11] ,
    \Tile_X6Y4_E6BEG[10] ,
    \Tile_X6Y4_E6BEG[9] ,
    \Tile_X6Y4_E6BEG[8] ,
    \Tile_X6Y4_E6BEG[7] ,
    \Tile_X6Y4_E6BEG[6] ,
    \Tile_X6Y4_E6BEG[5] ,
    \Tile_X6Y4_E6BEG[4] ,
    \Tile_X6Y4_E6BEG[3] ,
    \Tile_X6Y4_E6BEG[2] ,
    \Tile_X6Y4_E6BEG[1] ,
    \Tile_X6Y4_E6BEG[0] }),
    .E6END({\Tile_X5Y4_E6BEG[11] ,
    \Tile_X5Y4_E6BEG[10] ,
    \Tile_X5Y4_E6BEG[9] ,
    \Tile_X5Y4_E6BEG[8] ,
    \Tile_X5Y4_E6BEG[7] ,
    \Tile_X5Y4_E6BEG[6] ,
    \Tile_X5Y4_E6BEG[5] ,
    \Tile_X5Y4_E6BEG[4] ,
    \Tile_X5Y4_E6BEG[3] ,
    \Tile_X5Y4_E6BEG[2] ,
    \Tile_X5Y4_E6BEG[1] ,
    \Tile_X5Y4_E6BEG[0] }),
    .EE4BEG({\Tile_X6Y4_EE4BEG[15] ,
    \Tile_X6Y4_EE4BEG[14] ,
    \Tile_X6Y4_EE4BEG[13] ,
    \Tile_X6Y4_EE4BEG[12] ,
    \Tile_X6Y4_EE4BEG[11] ,
    \Tile_X6Y4_EE4BEG[10] ,
    \Tile_X6Y4_EE4BEG[9] ,
    \Tile_X6Y4_EE4BEG[8] ,
    \Tile_X6Y4_EE4BEG[7] ,
    \Tile_X6Y4_EE4BEG[6] ,
    \Tile_X6Y4_EE4BEG[5] ,
    \Tile_X6Y4_EE4BEG[4] ,
    \Tile_X6Y4_EE4BEG[3] ,
    \Tile_X6Y4_EE4BEG[2] ,
    \Tile_X6Y4_EE4BEG[1] ,
    \Tile_X6Y4_EE4BEG[0] }),
    .EE4END({\Tile_X5Y4_EE4BEG[15] ,
    \Tile_X5Y4_EE4BEG[14] ,
    \Tile_X5Y4_EE4BEG[13] ,
    \Tile_X5Y4_EE4BEG[12] ,
    \Tile_X5Y4_EE4BEG[11] ,
    \Tile_X5Y4_EE4BEG[10] ,
    \Tile_X5Y4_EE4BEG[9] ,
    \Tile_X5Y4_EE4BEG[8] ,
    \Tile_X5Y4_EE4BEG[7] ,
    \Tile_X5Y4_EE4BEG[6] ,
    \Tile_X5Y4_EE4BEG[5] ,
    \Tile_X5Y4_EE4BEG[4] ,
    \Tile_X5Y4_EE4BEG[3] ,
    \Tile_X5Y4_EE4BEG[2] ,
    \Tile_X5Y4_EE4BEG[1] ,
    \Tile_X5Y4_EE4BEG[0] }),
    .FrameData({\Tile_X5Y4_FrameData_O[31] ,
    \Tile_X5Y4_FrameData_O[30] ,
    \Tile_X5Y4_FrameData_O[29] ,
    \Tile_X5Y4_FrameData_O[28] ,
    \Tile_X5Y4_FrameData_O[27] ,
    \Tile_X5Y4_FrameData_O[26] ,
    \Tile_X5Y4_FrameData_O[25] ,
    \Tile_X5Y4_FrameData_O[24] ,
    \Tile_X5Y4_FrameData_O[23] ,
    \Tile_X5Y4_FrameData_O[22] ,
    \Tile_X5Y4_FrameData_O[21] ,
    \Tile_X5Y4_FrameData_O[20] ,
    \Tile_X5Y4_FrameData_O[19] ,
    \Tile_X5Y4_FrameData_O[18] ,
    \Tile_X5Y4_FrameData_O[17] ,
    \Tile_X5Y4_FrameData_O[16] ,
    \Tile_X5Y4_FrameData_O[15] ,
    \Tile_X5Y4_FrameData_O[14] ,
    \Tile_X5Y4_FrameData_O[13] ,
    \Tile_X5Y4_FrameData_O[12] ,
    \Tile_X5Y4_FrameData_O[11] ,
    \Tile_X5Y4_FrameData_O[10] ,
    \Tile_X5Y4_FrameData_O[9] ,
    \Tile_X5Y4_FrameData_O[8] ,
    \Tile_X5Y4_FrameData_O[7] ,
    \Tile_X5Y4_FrameData_O[6] ,
    \Tile_X5Y4_FrameData_O[5] ,
    \Tile_X5Y4_FrameData_O[4] ,
    \Tile_X5Y4_FrameData_O[3] ,
    \Tile_X5Y4_FrameData_O[2] ,
    \Tile_X5Y4_FrameData_O[1] ,
    \Tile_X5Y4_FrameData_O[0] }),
    .FrameData_O({\Tile_X6Y4_FrameData_O[31] ,
    \Tile_X6Y4_FrameData_O[30] ,
    \Tile_X6Y4_FrameData_O[29] ,
    \Tile_X6Y4_FrameData_O[28] ,
    \Tile_X6Y4_FrameData_O[27] ,
    \Tile_X6Y4_FrameData_O[26] ,
    \Tile_X6Y4_FrameData_O[25] ,
    \Tile_X6Y4_FrameData_O[24] ,
    \Tile_X6Y4_FrameData_O[23] ,
    \Tile_X6Y4_FrameData_O[22] ,
    \Tile_X6Y4_FrameData_O[21] ,
    \Tile_X6Y4_FrameData_O[20] ,
    \Tile_X6Y4_FrameData_O[19] ,
    \Tile_X6Y4_FrameData_O[18] ,
    \Tile_X6Y4_FrameData_O[17] ,
    \Tile_X6Y4_FrameData_O[16] ,
    \Tile_X6Y4_FrameData_O[15] ,
    \Tile_X6Y4_FrameData_O[14] ,
    \Tile_X6Y4_FrameData_O[13] ,
    \Tile_X6Y4_FrameData_O[12] ,
    \Tile_X6Y4_FrameData_O[11] ,
    \Tile_X6Y4_FrameData_O[10] ,
    \Tile_X6Y4_FrameData_O[9] ,
    \Tile_X6Y4_FrameData_O[8] ,
    \Tile_X6Y4_FrameData_O[7] ,
    \Tile_X6Y4_FrameData_O[6] ,
    \Tile_X6Y4_FrameData_O[5] ,
    \Tile_X6Y4_FrameData_O[4] ,
    \Tile_X6Y4_FrameData_O[3] ,
    \Tile_X6Y4_FrameData_O[2] ,
    \Tile_X6Y4_FrameData_O[1] ,
    \Tile_X6Y4_FrameData_O[0] }),
    .FrameStrobe({\Tile_X6Y5_FrameStrobe_O[19] ,
    \Tile_X6Y5_FrameStrobe_O[18] ,
    \Tile_X6Y5_FrameStrobe_O[17] ,
    \Tile_X6Y5_FrameStrobe_O[16] ,
    \Tile_X6Y5_FrameStrobe_O[15] ,
    \Tile_X6Y5_FrameStrobe_O[14] ,
    \Tile_X6Y5_FrameStrobe_O[13] ,
    \Tile_X6Y5_FrameStrobe_O[12] ,
    \Tile_X6Y5_FrameStrobe_O[11] ,
    \Tile_X6Y5_FrameStrobe_O[10] ,
    \Tile_X6Y5_FrameStrobe_O[9] ,
    \Tile_X6Y5_FrameStrobe_O[8] ,
    \Tile_X6Y5_FrameStrobe_O[7] ,
    \Tile_X6Y5_FrameStrobe_O[6] ,
    \Tile_X6Y5_FrameStrobe_O[5] ,
    \Tile_X6Y5_FrameStrobe_O[4] ,
    \Tile_X6Y5_FrameStrobe_O[3] ,
    \Tile_X6Y5_FrameStrobe_O[2] ,
    \Tile_X6Y5_FrameStrobe_O[1] ,
    \Tile_X6Y5_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X6Y4_FrameStrobe_O[19] ,
    \Tile_X6Y4_FrameStrobe_O[18] ,
    \Tile_X6Y4_FrameStrobe_O[17] ,
    \Tile_X6Y4_FrameStrobe_O[16] ,
    \Tile_X6Y4_FrameStrobe_O[15] ,
    \Tile_X6Y4_FrameStrobe_O[14] ,
    \Tile_X6Y4_FrameStrobe_O[13] ,
    \Tile_X6Y4_FrameStrobe_O[12] ,
    \Tile_X6Y4_FrameStrobe_O[11] ,
    \Tile_X6Y4_FrameStrobe_O[10] ,
    \Tile_X6Y4_FrameStrobe_O[9] ,
    \Tile_X6Y4_FrameStrobe_O[8] ,
    \Tile_X6Y4_FrameStrobe_O[7] ,
    \Tile_X6Y4_FrameStrobe_O[6] ,
    \Tile_X6Y4_FrameStrobe_O[5] ,
    \Tile_X6Y4_FrameStrobe_O[4] ,
    \Tile_X6Y4_FrameStrobe_O[3] ,
    \Tile_X6Y4_FrameStrobe_O[2] ,
    \Tile_X6Y4_FrameStrobe_O[1] ,
    \Tile_X6Y4_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X6Y4_N1BEG[3] ,
    \Tile_X6Y4_N1BEG[2] ,
    \Tile_X6Y4_N1BEG[1] ,
    \Tile_X6Y4_N1BEG[0] }),
    .N1END({\Tile_X6Y5_N1BEG[3] ,
    \Tile_X6Y5_N1BEG[2] ,
    \Tile_X6Y5_N1BEG[1] ,
    \Tile_X6Y5_N1BEG[0] }),
    .N2BEG({\Tile_X6Y4_N2BEG[7] ,
    \Tile_X6Y4_N2BEG[6] ,
    \Tile_X6Y4_N2BEG[5] ,
    \Tile_X6Y4_N2BEG[4] ,
    \Tile_X6Y4_N2BEG[3] ,
    \Tile_X6Y4_N2BEG[2] ,
    \Tile_X6Y4_N2BEG[1] ,
    \Tile_X6Y4_N2BEG[0] }),
    .N2BEGb({\Tile_X6Y4_N2BEGb[7] ,
    \Tile_X6Y4_N2BEGb[6] ,
    \Tile_X6Y4_N2BEGb[5] ,
    \Tile_X6Y4_N2BEGb[4] ,
    \Tile_X6Y4_N2BEGb[3] ,
    \Tile_X6Y4_N2BEGb[2] ,
    \Tile_X6Y4_N2BEGb[1] ,
    \Tile_X6Y4_N2BEGb[0] }),
    .N2END({\Tile_X6Y5_N2BEGb[7] ,
    \Tile_X6Y5_N2BEGb[6] ,
    \Tile_X6Y5_N2BEGb[5] ,
    \Tile_X6Y5_N2BEGb[4] ,
    \Tile_X6Y5_N2BEGb[3] ,
    \Tile_X6Y5_N2BEGb[2] ,
    \Tile_X6Y5_N2BEGb[1] ,
    \Tile_X6Y5_N2BEGb[0] }),
    .N2MID({\Tile_X6Y5_N2BEG[7] ,
    \Tile_X6Y5_N2BEG[6] ,
    \Tile_X6Y5_N2BEG[5] ,
    \Tile_X6Y5_N2BEG[4] ,
    \Tile_X6Y5_N2BEG[3] ,
    \Tile_X6Y5_N2BEG[2] ,
    \Tile_X6Y5_N2BEG[1] ,
    \Tile_X6Y5_N2BEG[0] }),
    .N4BEG({\Tile_X6Y4_N4BEG[15] ,
    \Tile_X6Y4_N4BEG[14] ,
    \Tile_X6Y4_N4BEG[13] ,
    \Tile_X6Y4_N4BEG[12] ,
    \Tile_X6Y4_N4BEG[11] ,
    \Tile_X6Y4_N4BEG[10] ,
    \Tile_X6Y4_N4BEG[9] ,
    \Tile_X6Y4_N4BEG[8] ,
    \Tile_X6Y4_N4BEG[7] ,
    \Tile_X6Y4_N4BEG[6] ,
    \Tile_X6Y4_N4BEG[5] ,
    \Tile_X6Y4_N4BEG[4] ,
    \Tile_X6Y4_N4BEG[3] ,
    \Tile_X6Y4_N4BEG[2] ,
    \Tile_X6Y4_N4BEG[1] ,
    \Tile_X6Y4_N4BEG[0] }),
    .N4END({\Tile_X6Y5_N4BEG[15] ,
    \Tile_X6Y5_N4BEG[14] ,
    \Tile_X6Y5_N4BEG[13] ,
    \Tile_X6Y5_N4BEG[12] ,
    \Tile_X6Y5_N4BEG[11] ,
    \Tile_X6Y5_N4BEG[10] ,
    \Tile_X6Y5_N4BEG[9] ,
    \Tile_X6Y5_N4BEG[8] ,
    \Tile_X6Y5_N4BEG[7] ,
    \Tile_X6Y5_N4BEG[6] ,
    \Tile_X6Y5_N4BEG[5] ,
    \Tile_X6Y5_N4BEG[4] ,
    \Tile_X6Y5_N4BEG[3] ,
    \Tile_X6Y5_N4BEG[2] ,
    \Tile_X6Y5_N4BEG[1] ,
    \Tile_X6Y5_N4BEG[0] }),
    .NN4BEG({\Tile_X6Y4_NN4BEG[15] ,
    \Tile_X6Y4_NN4BEG[14] ,
    \Tile_X6Y4_NN4BEG[13] ,
    \Tile_X6Y4_NN4BEG[12] ,
    \Tile_X6Y4_NN4BEG[11] ,
    \Tile_X6Y4_NN4BEG[10] ,
    \Tile_X6Y4_NN4BEG[9] ,
    \Tile_X6Y4_NN4BEG[8] ,
    \Tile_X6Y4_NN4BEG[7] ,
    \Tile_X6Y4_NN4BEG[6] ,
    \Tile_X6Y4_NN4BEG[5] ,
    \Tile_X6Y4_NN4BEG[4] ,
    \Tile_X6Y4_NN4BEG[3] ,
    \Tile_X6Y4_NN4BEG[2] ,
    \Tile_X6Y4_NN4BEG[1] ,
    \Tile_X6Y4_NN4BEG[0] }),
    .NN4END({\Tile_X6Y5_NN4BEG[15] ,
    \Tile_X6Y5_NN4BEG[14] ,
    \Tile_X6Y5_NN4BEG[13] ,
    \Tile_X6Y5_NN4BEG[12] ,
    \Tile_X6Y5_NN4BEG[11] ,
    \Tile_X6Y5_NN4BEG[10] ,
    \Tile_X6Y5_NN4BEG[9] ,
    \Tile_X6Y5_NN4BEG[8] ,
    \Tile_X6Y5_NN4BEG[7] ,
    \Tile_X6Y5_NN4BEG[6] ,
    \Tile_X6Y5_NN4BEG[5] ,
    \Tile_X6Y5_NN4BEG[4] ,
    \Tile_X6Y5_NN4BEG[3] ,
    \Tile_X6Y5_NN4BEG[2] ,
    \Tile_X6Y5_NN4BEG[1] ,
    \Tile_X6Y5_NN4BEG[0] }),
    .S1BEG({\Tile_X6Y4_S1BEG[3] ,
    \Tile_X6Y4_S1BEG[2] ,
    \Tile_X6Y4_S1BEG[1] ,
    \Tile_X6Y4_S1BEG[0] }),
    .S1END({\Tile_X6Y3_S1BEG[3] ,
    \Tile_X6Y3_S1BEG[2] ,
    \Tile_X6Y3_S1BEG[1] ,
    \Tile_X6Y3_S1BEG[0] }),
    .S2BEG({\Tile_X6Y4_S2BEG[7] ,
    \Tile_X6Y4_S2BEG[6] ,
    \Tile_X6Y4_S2BEG[5] ,
    \Tile_X6Y4_S2BEG[4] ,
    \Tile_X6Y4_S2BEG[3] ,
    \Tile_X6Y4_S2BEG[2] ,
    \Tile_X6Y4_S2BEG[1] ,
    \Tile_X6Y4_S2BEG[0] }),
    .S2BEGb({\Tile_X6Y4_S2BEGb[7] ,
    \Tile_X6Y4_S2BEGb[6] ,
    \Tile_X6Y4_S2BEGb[5] ,
    \Tile_X6Y4_S2BEGb[4] ,
    \Tile_X6Y4_S2BEGb[3] ,
    \Tile_X6Y4_S2BEGb[2] ,
    \Tile_X6Y4_S2BEGb[1] ,
    \Tile_X6Y4_S2BEGb[0] }),
    .S2END({\Tile_X6Y3_S2BEGb[7] ,
    \Tile_X6Y3_S2BEGb[6] ,
    \Tile_X6Y3_S2BEGb[5] ,
    \Tile_X6Y3_S2BEGb[4] ,
    \Tile_X6Y3_S2BEGb[3] ,
    \Tile_X6Y3_S2BEGb[2] ,
    \Tile_X6Y3_S2BEGb[1] ,
    \Tile_X6Y3_S2BEGb[0] }),
    .S2MID({\Tile_X6Y3_S2BEG[7] ,
    \Tile_X6Y3_S2BEG[6] ,
    \Tile_X6Y3_S2BEG[5] ,
    \Tile_X6Y3_S2BEG[4] ,
    \Tile_X6Y3_S2BEG[3] ,
    \Tile_X6Y3_S2BEG[2] ,
    \Tile_X6Y3_S2BEG[1] ,
    \Tile_X6Y3_S2BEG[0] }),
    .S4BEG({\Tile_X6Y4_S4BEG[15] ,
    \Tile_X6Y4_S4BEG[14] ,
    \Tile_X6Y4_S4BEG[13] ,
    \Tile_X6Y4_S4BEG[12] ,
    \Tile_X6Y4_S4BEG[11] ,
    \Tile_X6Y4_S4BEG[10] ,
    \Tile_X6Y4_S4BEG[9] ,
    \Tile_X6Y4_S4BEG[8] ,
    \Tile_X6Y4_S4BEG[7] ,
    \Tile_X6Y4_S4BEG[6] ,
    \Tile_X6Y4_S4BEG[5] ,
    \Tile_X6Y4_S4BEG[4] ,
    \Tile_X6Y4_S4BEG[3] ,
    \Tile_X6Y4_S4BEG[2] ,
    \Tile_X6Y4_S4BEG[1] ,
    \Tile_X6Y4_S4BEG[0] }),
    .S4END({\Tile_X6Y3_S4BEG[15] ,
    \Tile_X6Y3_S4BEG[14] ,
    \Tile_X6Y3_S4BEG[13] ,
    \Tile_X6Y3_S4BEG[12] ,
    \Tile_X6Y3_S4BEG[11] ,
    \Tile_X6Y3_S4BEG[10] ,
    \Tile_X6Y3_S4BEG[9] ,
    \Tile_X6Y3_S4BEG[8] ,
    \Tile_X6Y3_S4BEG[7] ,
    \Tile_X6Y3_S4BEG[6] ,
    \Tile_X6Y3_S4BEG[5] ,
    \Tile_X6Y3_S4BEG[4] ,
    \Tile_X6Y3_S4BEG[3] ,
    \Tile_X6Y3_S4BEG[2] ,
    \Tile_X6Y3_S4BEG[1] ,
    \Tile_X6Y3_S4BEG[0] }),
    .SS4BEG({\Tile_X6Y4_SS4BEG[15] ,
    \Tile_X6Y4_SS4BEG[14] ,
    \Tile_X6Y4_SS4BEG[13] ,
    \Tile_X6Y4_SS4BEG[12] ,
    \Tile_X6Y4_SS4BEG[11] ,
    \Tile_X6Y4_SS4BEG[10] ,
    \Tile_X6Y4_SS4BEG[9] ,
    \Tile_X6Y4_SS4BEG[8] ,
    \Tile_X6Y4_SS4BEG[7] ,
    \Tile_X6Y4_SS4BEG[6] ,
    \Tile_X6Y4_SS4BEG[5] ,
    \Tile_X6Y4_SS4BEG[4] ,
    \Tile_X6Y4_SS4BEG[3] ,
    \Tile_X6Y4_SS4BEG[2] ,
    \Tile_X6Y4_SS4BEG[1] ,
    \Tile_X6Y4_SS4BEG[0] }),
    .SS4END({\Tile_X6Y3_SS4BEG[15] ,
    \Tile_X6Y3_SS4BEG[14] ,
    \Tile_X6Y3_SS4BEG[13] ,
    \Tile_X6Y3_SS4BEG[12] ,
    \Tile_X6Y3_SS4BEG[11] ,
    \Tile_X6Y3_SS4BEG[10] ,
    \Tile_X6Y3_SS4BEG[9] ,
    \Tile_X6Y3_SS4BEG[8] ,
    \Tile_X6Y3_SS4BEG[7] ,
    \Tile_X6Y3_SS4BEG[6] ,
    \Tile_X6Y3_SS4BEG[5] ,
    \Tile_X6Y3_SS4BEG[4] ,
    \Tile_X6Y3_SS4BEG[3] ,
    \Tile_X6Y3_SS4BEG[2] ,
    \Tile_X6Y3_SS4BEG[1] ,
    \Tile_X6Y3_SS4BEG[0] }),
    .W1BEG({\Tile_X6Y4_W1BEG[3] ,
    \Tile_X6Y4_W1BEG[2] ,
    \Tile_X6Y4_W1BEG[1] ,
    \Tile_X6Y4_W1BEG[0] }),
    .W1END({\Tile_X7Y4_W1BEG[3] ,
    \Tile_X7Y4_W1BEG[2] ,
    \Tile_X7Y4_W1BEG[1] ,
    \Tile_X7Y4_W1BEG[0] }),
    .W2BEG({\Tile_X6Y4_W2BEG[7] ,
    \Tile_X6Y4_W2BEG[6] ,
    \Tile_X6Y4_W2BEG[5] ,
    \Tile_X6Y4_W2BEG[4] ,
    \Tile_X6Y4_W2BEG[3] ,
    \Tile_X6Y4_W2BEG[2] ,
    \Tile_X6Y4_W2BEG[1] ,
    \Tile_X6Y4_W2BEG[0] }),
    .W2BEGb({\Tile_X6Y4_W2BEGb[7] ,
    \Tile_X6Y4_W2BEGb[6] ,
    \Tile_X6Y4_W2BEGb[5] ,
    \Tile_X6Y4_W2BEGb[4] ,
    \Tile_X6Y4_W2BEGb[3] ,
    \Tile_X6Y4_W2BEGb[2] ,
    \Tile_X6Y4_W2BEGb[1] ,
    \Tile_X6Y4_W2BEGb[0] }),
    .W2END({\Tile_X7Y4_W2BEGb[7] ,
    \Tile_X7Y4_W2BEGb[6] ,
    \Tile_X7Y4_W2BEGb[5] ,
    \Tile_X7Y4_W2BEGb[4] ,
    \Tile_X7Y4_W2BEGb[3] ,
    \Tile_X7Y4_W2BEGb[2] ,
    \Tile_X7Y4_W2BEGb[1] ,
    \Tile_X7Y4_W2BEGb[0] }),
    .W2MID({\Tile_X7Y4_W2BEG[7] ,
    \Tile_X7Y4_W2BEG[6] ,
    \Tile_X7Y4_W2BEG[5] ,
    \Tile_X7Y4_W2BEG[4] ,
    \Tile_X7Y4_W2BEG[3] ,
    \Tile_X7Y4_W2BEG[2] ,
    \Tile_X7Y4_W2BEG[1] ,
    \Tile_X7Y4_W2BEG[0] }),
    .W6BEG({\Tile_X6Y4_W6BEG[11] ,
    \Tile_X6Y4_W6BEG[10] ,
    \Tile_X6Y4_W6BEG[9] ,
    \Tile_X6Y4_W6BEG[8] ,
    \Tile_X6Y4_W6BEG[7] ,
    \Tile_X6Y4_W6BEG[6] ,
    \Tile_X6Y4_W6BEG[5] ,
    \Tile_X6Y4_W6BEG[4] ,
    \Tile_X6Y4_W6BEG[3] ,
    \Tile_X6Y4_W6BEG[2] ,
    \Tile_X6Y4_W6BEG[1] ,
    \Tile_X6Y4_W6BEG[0] }),
    .W6END({\Tile_X7Y4_W6BEG[11] ,
    \Tile_X7Y4_W6BEG[10] ,
    \Tile_X7Y4_W6BEG[9] ,
    \Tile_X7Y4_W6BEG[8] ,
    \Tile_X7Y4_W6BEG[7] ,
    \Tile_X7Y4_W6BEG[6] ,
    \Tile_X7Y4_W6BEG[5] ,
    \Tile_X7Y4_W6BEG[4] ,
    \Tile_X7Y4_W6BEG[3] ,
    \Tile_X7Y4_W6BEG[2] ,
    \Tile_X7Y4_W6BEG[1] ,
    \Tile_X7Y4_W6BEG[0] }),
    .WW4BEG({\Tile_X6Y4_WW4BEG[15] ,
    \Tile_X6Y4_WW4BEG[14] ,
    \Tile_X6Y4_WW4BEG[13] ,
    \Tile_X6Y4_WW4BEG[12] ,
    \Tile_X6Y4_WW4BEG[11] ,
    \Tile_X6Y4_WW4BEG[10] ,
    \Tile_X6Y4_WW4BEG[9] ,
    \Tile_X6Y4_WW4BEG[8] ,
    \Tile_X6Y4_WW4BEG[7] ,
    \Tile_X6Y4_WW4BEG[6] ,
    \Tile_X6Y4_WW4BEG[5] ,
    \Tile_X6Y4_WW4BEG[4] ,
    \Tile_X6Y4_WW4BEG[3] ,
    \Tile_X6Y4_WW4BEG[2] ,
    \Tile_X6Y4_WW4BEG[1] ,
    \Tile_X6Y4_WW4BEG[0] }),
    .WW4END({\Tile_X7Y4_WW4BEG[15] ,
    \Tile_X7Y4_WW4BEG[14] ,
    \Tile_X7Y4_WW4BEG[13] ,
    \Tile_X7Y4_WW4BEG[12] ,
    \Tile_X7Y4_WW4BEG[11] ,
    \Tile_X7Y4_WW4BEG[10] ,
    \Tile_X7Y4_WW4BEG[9] ,
    \Tile_X7Y4_WW4BEG[8] ,
    \Tile_X7Y4_WW4BEG[7] ,
    \Tile_X7Y4_WW4BEG[6] ,
    \Tile_X7Y4_WW4BEG[5] ,
    \Tile_X7Y4_WW4BEG[4] ,
    \Tile_X7Y4_WW4BEG[3] ,
    \Tile_X7Y4_WW4BEG[2] ,
    \Tile_X7Y4_WW4BEG[1] ,
    \Tile_X7Y4_WW4BEG[0] }));
 LUT4AB Tile_X6Y5_LUT4AB (.Ci(Tile_X6Y6_Co),
    .Co(Tile_X6Y5_Co),
    .UserCLK(Tile_X6Y6_UserCLKo),
    .UserCLKo(Tile_X6Y5_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X6Y5_E1BEG[3] ,
    \Tile_X6Y5_E1BEG[2] ,
    \Tile_X6Y5_E1BEG[1] ,
    \Tile_X6Y5_E1BEG[0] }),
    .E1END({\Tile_X5Y5_E1BEG[3] ,
    \Tile_X5Y5_E1BEG[2] ,
    \Tile_X5Y5_E1BEG[1] ,
    \Tile_X5Y5_E1BEG[0] }),
    .E2BEG({\Tile_X6Y5_E2BEG[7] ,
    \Tile_X6Y5_E2BEG[6] ,
    \Tile_X6Y5_E2BEG[5] ,
    \Tile_X6Y5_E2BEG[4] ,
    \Tile_X6Y5_E2BEG[3] ,
    \Tile_X6Y5_E2BEG[2] ,
    \Tile_X6Y5_E2BEG[1] ,
    \Tile_X6Y5_E2BEG[0] }),
    .E2BEGb({\Tile_X6Y5_E2BEGb[7] ,
    \Tile_X6Y5_E2BEGb[6] ,
    \Tile_X6Y5_E2BEGb[5] ,
    \Tile_X6Y5_E2BEGb[4] ,
    \Tile_X6Y5_E2BEGb[3] ,
    \Tile_X6Y5_E2BEGb[2] ,
    \Tile_X6Y5_E2BEGb[1] ,
    \Tile_X6Y5_E2BEGb[0] }),
    .E2END({\Tile_X5Y5_E2BEGb[7] ,
    \Tile_X5Y5_E2BEGb[6] ,
    \Tile_X5Y5_E2BEGb[5] ,
    \Tile_X5Y5_E2BEGb[4] ,
    \Tile_X5Y5_E2BEGb[3] ,
    \Tile_X5Y5_E2BEGb[2] ,
    \Tile_X5Y5_E2BEGb[1] ,
    \Tile_X5Y5_E2BEGb[0] }),
    .E2MID({\Tile_X5Y5_E2BEG[7] ,
    \Tile_X5Y5_E2BEG[6] ,
    \Tile_X5Y5_E2BEG[5] ,
    \Tile_X5Y5_E2BEG[4] ,
    \Tile_X5Y5_E2BEG[3] ,
    \Tile_X5Y5_E2BEG[2] ,
    \Tile_X5Y5_E2BEG[1] ,
    \Tile_X5Y5_E2BEG[0] }),
    .E6BEG({\Tile_X6Y5_E6BEG[11] ,
    \Tile_X6Y5_E6BEG[10] ,
    \Tile_X6Y5_E6BEG[9] ,
    \Tile_X6Y5_E6BEG[8] ,
    \Tile_X6Y5_E6BEG[7] ,
    \Tile_X6Y5_E6BEG[6] ,
    \Tile_X6Y5_E6BEG[5] ,
    \Tile_X6Y5_E6BEG[4] ,
    \Tile_X6Y5_E6BEG[3] ,
    \Tile_X6Y5_E6BEG[2] ,
    \Tile_X6Y5_E6BEG[1] ,
    \Tile_X6Y5_E6BEG[0] }),
    .E6END({\Tile_X5Y5_E6BEG[11] ,
    \Tile_X5Y5_E6BEG[10] ,
    \Tile_X5Y5_E6BEG[9] ,
    \Tile_X5Y5_E6BEG[8] ,
    \Tile_X5Y5_E6BEG[7] ,
    \Tile_X5Y5_E6BEG[6] ,
    \Tile_X5Y5_E6BEG[5] ,
    \Tile_X5Y5_E6BEG[4] ,
    \Tile_X5Y5_E6BEG[3] ,
    \Tile_X5Y5_E6BEG[2] ,
    \Tile_X5Y5_E6BEG[1] ,
    \Tile_X5Y5_E6BEG[0] }),
    .EE4BEG({\Tile_X6Y5_EE4BEG[15] ,
    \Tile_X6Y5_EE4BEG[14] ,
    \Tile_X6Y5_EE4BEG[13] ,
    \Tile_X6Y5_EE4BEG[12] ,
    \Tile_X6Y5_EE4BEG[11] ,
    \Tile_X6Y5_EE4BEG[10] ,
    \Tile_X6Y5_EE4BEG[9] ,
    \Tile_X6Y5_EE4BEG[8] ,
    \Tile_X6Y5_EE4BEG[7] ,
    \Tile_X6Y5_EE4BEG[6] ,
    \Tile_X6Y5_EE4BEG[5] ,
    \Tile_X6Y5_EE4BEG[4] ,
    \Tile_X6Y5_EE4BEG[3] ,
    \Tile_X6Y5_EE4BEG[2] ,
    \Tile_X6Y5_EE4BEG[1] ,
    \Tile_X6Y5_EE4BEG[0] }),
    .EE4END({\Tile_X5Y5_EE4BEG[15] ,
    \Tile_X5Y5_EE4BEG[14] ,
    \Tile_X5Y5_EE4BEG[13] ,
    \Tile_X5Y5_EE4BEG[12] ,
    \Tile_X5Y5_EE4BEG[11] ,
    \Tile_X5Y5_EE4BEG[10] ,
    \Tile_X5Y5_EE4BEG[9] ,
    \Tile_X5Y5_EE4BEG[8] ,
    \Tile_X5Y5_EE4BEG[7] ,
    \Tile_X5Y5_EE4BEG[6] ,
    \Tile_X5Y5_EE4BEG[5] ,
    \Tile_X5Y5_EE4BEG[4] ,
    \Tile_X5Y5_EE4BEG[3] ,
    \Tile_X5Y5_EE4BEG[2] ,
    \Tile_X5Y5_EE4BEG[1] ,
    \Tile_X5Y5_EE4BEG[0] }),
    .FrameData({\Tile_X5Y5_FrameData_O[31] ,
    \Tile_X5Y5_FrameData_O[30] ,
    \Tile_X5Y5_FrameData_O[29] ,
    \Tile_X5Y5_FrameData_O[28] ,
    \Tile_X5Y5_FrameData_O[27] ,
    \Tile_X5Y5_FrameData_O[26] ,
    \Tile_X5Y5_FrameData_O[25] ,
    \Tile_X5Y5_FrameData_O[24] ,
    \Tile_X5Y5_FrameData_O[23] ,
    \Tile_X5Y5_FrameData_O[22] ,
    \Tile_X5Y5_FrameData_O[21] ,
    \Tile_X5Y5_FrameData_O[20] ,
    \Tile_X5Y5_FrameData_O[19] ,
    \Tile_X5Y5_FrameData_O[18] ,
    \Tile_X5Y5_FrameData_O[17] ,
    \Tile_X5Y5_FrameData_O[16] ,
    \Tile_X5Y5_FrameData_O[15] ,
    \Tile_X5Y5_FrameData_O[14] ,
    \Tile_X5Y5_FrameData_O[13] ,
    \Tile_X5Y5_FrameData_O[12] ,
    \Tile_X5Y5_FrameData_O[11] ,
    \Tile_X5Y5_FrameData_O[10] ,
    \Tile_X5Y5_FrameData_O[9] ,
    \Tile_X5Y5_FrameData_O[8] ,
    \Tile_X5Y5_FrameData_O[7] ,
    \Tile_X5Y5_FrameData_O[6] ,
    \Tile_X5Y5_FrameData_O[5] ,
    \Tile_X5Y5_FrameData_O[4] ,
    \Tile_X5Y5_FrameData_O[3] ,
    \Tile_X5Y5_FrameData_O[2] ,
    \Tile_X5Y5_FrameData_O[1] ,
    \Tile_X5Y5_FrameData_O[0] }),
    .FrameData_O({\Tile_X6Y5_FrameData_O[31] ,
    \Tile_X6Y5_FrameData_O[30] ,
    \Tile_X6Y5_FrameData_O[29] ,
    \Tile_X6Y5_FrameData_O[28] ,
    \Tile_X6Y5_FrameData_O[27] ,
    \Tile_X6Y5_FrameData_O[26] ,
    \Tile_X6Y5_FrameData_O[25] ,
    \Tile_X6Y5_FrameData_O[24] ,
    \Tile_X6Y5_FrameData_O[23] ,
    \Tile_X6Y5_FrameData_O[22] ,
    \Tile_X6Y5_FrameData_O[21] ,
    \Tile_X6Y5_FrameData_O[20] ,
    \Tile_X6Y5_FrameData_O[19] ,
    \Tile_X6Y5_FrameData_O[18] ,
    \Tile_X6Y5_FrameData_O[17] ,
    \Tile_X6Y5_FrameData_O[16] ,
    \Tile_X6Y5_FrameData_O[15] ,
    \Tile_X6Y5_FrameData_O[14] ,
    \Tile_X6Y5_FrameData_O[13] ,
    \Tile_X6Y5_FrameData_O[12] ,
    \Tile_X6Y5_FrameData_O[11] ,
    \Tile_X6Y5_FrameData_O[10] ,
    \Tile_X6Y5_FrameData_O[9] ,
    \Tile_X6Y5_FrameData_O[8] ,
    \Tile_X6Y5_FrameData_O[7] ,
    \Tile_X6Y5_FrameData_O[6] ,
    \Tile_X6Y5_FrameData_O[5] ,
    \Tile_X6Y5_FrameData_O[4] ,
    \Tile_X6Y5_FrameData_O[3] ,
    \Tile_X6Y5_FrameData_O[2] ,
    \Tile_X6Y5_FrameData_O[1] ,
    \Tile_X6Y5_FrameData_O[0] }),
    .FrameStrobe({\Tile_X6Y6_FrameStrobe_O[19] ,
    \Tile_X6Y6_FrameStrobe_O[18] ,
    \Tile_X6Y6_FrameStrobe_O[17] ,
    \Tile_X6Y6_FrameStrobe_O[16] ,
    \Tile_X6Y6_FrameStrobe_O[15] ,
    \Tile_X6Y6_FrameStrobe_O[14] ,
    \Tile_X6Y6_FrameStrobe_O[13] ,
    \Tile_X6Y6_FrameStrobe_O[12] ,
    \Tile_X6Y6_FrameStrobe_O[11] ,
    \Tile_X6Y6_FrameStrobe_O[10] ,
    \Tile_X6Y6_FrameStrobe_O[9] ,
    \Tile_X6Y6_FrameStrobe_O[8] ,
    \Tile_X6Y6_FrameStrobe_O[7] ,
    \Tile_X6Y6_FrameStrobe_O[6] ,
    \Tile_X6Y6_FrameStrobe_O[5] ,
    \Tile_X6Y6_FrameStrobe_O[4] ,
    \Tile_X6Y6_FrameStrobe_O[3] ,
    \Tile_X6Y6_FrameStrobe_O[2] ,
    \Tile_X6Y6_FrameStrobe_O[1] ,
    \Tile_X6Y6_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X6Y5_FrameStrobe_O[19] ,
    \Tile_X6Y5_FrameStrobe_O[18] ,
    \Tile_X6Y5_FrameStrobe_O[17] ,
    \Tile_X6Y5_FrameStrobe_O[16] ,
    \Tile_X6Y5_FrameStrobe_O[15] ,
    \Tile_X6Y5_FrameStrobe_O[14] ,
    \Tile_X6Y5_FrameStrobe_O[13] ,
    \Tile_X6Y5_FrameStrobe_O[12] ,
    \Tile_X6Y5_FrameStrobe_O[11] ,
    \Tile_X6Y5_FrameStrobe_O[10] ,
    \Tile_X6Y5_FrameStrobe_O[9] ,
    \Tile_X6Y5_FrameStrobe_O[8] ,
    \Tile_X6Y5_FrameStrobe_O[7] ,
    \Tile_X6Y5_FrameStrobe_O[6] ,
    \Tile_X6Y5_FrameStrobe_O[5] ,
    \Tile_X6Y5_FrameStrobe_O[4] ,
    \Tile_X6Y5_FrameStrobe_O[3] ,
    \Tile_X6Y5_FrameStrobe_O[2] ,
    \Tile_X6Y5_FrameStrobe_O[1] ,
    \Tile_X6Y5_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X6Y5_N1BEG[3] ,
    \Tile_X6Y5_N1BEG[2] ,
    \Tile_X6Y5_N1BEG[1] ,
    \Tile_X6Y5_N1BEG[0] }),
    .N1END({\Tile_X6Y6_N1BEG[3] ,
    \Tile_X6Y6_N1BEG[2] ,
    \Tile_X6Y6_N1BEG[1] ,
    \Tile_X6Y6_N1BEG[0] }),
    .N2BEG({\Tile_X6Y5_N2BEG[7] ,
    \Tile_X6Y5_N2BEG[6] ,
    \Tile_X6Y5_N2BEG[5] ,
    \Tile_X6Y5_N2BEG[4] ,
    \Tile_X6Y5_N2BEG[3] ,
    \Tile_X6Y5_N2BEG[2] ,
    \Tile_X6Y5_N2BEG[1] ,
    \Tile_X6Y5_N2BEG[0] }),
    .N2BEGb({\Tile_X6Y5_N2BEGb[7] ,
    \Tile_X6Y5_N2BEGb[6] ,
    \Tile_X6Y5_N2BEGb[5] ,
    \Tile_X6Y5_N2BEGb[4] ,
    \Tile_X6Y5_N2BEGb[3] ,
    \Tile_X6Y5_N2BEGb[2] ,
    \Tile_X6Y5_N2BEGb[1] ,
    \Tile_X6Y5_N2BEGb[0] }),
    .N2END({\Tile_X6Y6_N2BEGb[7] ,
    \Tile_X6Y6_N2BEGb[6] ,
    \Tile_X6Y6_N2BEGb[5] ,
    \Tile_X6Y6_N2BEGb[4] ,
    \Tile_X6Y6_N2BEGb[3] ,
    \Tile_X6Y6_N2BEGb[2] ,
    \Tile_X6Y6_N2BEGb[1] ,
    \Tile_X6Y6_N2BEGb[0] }),
    .N2MID({\Tile_X6Y6_N2BEG[7] ,
    \Tile_X6Y6_N2BEG[6] ,
    \Tile_X6Y6_N2BEG[5] ,
    \Tile_X6Y6_N2BEG[4] ,
    \Tile_X6Y6_N2BEG[3] ,
    \Tile_X6Y6_N2BEG[2] ,
    \Tile_X6Y6_N2BEG[1] ,
    \Tile_X6Y6_N2BEG[0] }),
    .N4BEG({\Tile_X6Y5_N4BEG[15] ,
    \Tile_X6Y5_N4BEG[14] ,
    \Tile_X6Y5_N4BEG[13] ,
    \Tile_X6Y5_N4BEG[12] ,
    \Tile_X6Y5_N4BEG[11] ,
    \Tile_X6Y5_N4BEG[10] ,
    \Tile_X6Y5_N4BEG[9] ,
    \Tile_X6Y5_N4BEG[8] ,
    \Tile_X6Y5_N4BEG[7] ,
    \Tile_X6Y5_N4BEG[6] ,
    \Tile_X6Y5_N4BEG[5] ,
    \Tile_X6Y5_N4BEG[4] ,
    \Tile_X6Y5_N4BEG[3] ,
    \Tile_X6Y5_N4BEG[2] ,
    \Tile_X6Y5_N4BEG[1] ,
    \Tile_X6Y5_N4BEG[0] }),
    .N4END({\Tile_X6Y6_N4BEG[15] ,
    \Tile_X6Y6_N4BEG[14] ,
    \Tile_X6Y6_N4BEG[13] ,
    \Tile_X6Y6_N4BEG[12] ,
    \Tile_X6Y6_N4BEG[11] ,
    \Tile_X6Y6_N4BEG[10] ,
    \Tile_X6Y6_N4BEG[9] ,
    \Tile_X6Y6_N4BEG[8] ,
    \Tile_X6Y6_N4BEG[7] ,
    \Tile_X6Y6_N4BEG[6] ,
    \Tile_X6Y6_N4BEG[5] ,
    \Tile_X6Y6_N4BEG[4] ,
    \Tile_X6Y6_N4BEG[3] ,
    \Tile_X6Y6_N4BEG[2] ,
    \Tile_X6Y6_N4BEG[1] ,
    \Tile_X6Y6_N4BEG[0] }),
    .NN4BEG({\Tile_X6Y5_NN4BEG[15] ,
    \Tile_X6Y5_NN4BEG[14] ,
    \Tile_X6Y5_NN4BEG[13] ,
    \Tile_X6Y5_NN4BEG[12] ,
    \Tile_X6Y5_NN4BEG[11] ,
    \Tile_X6Y5_NN4BEG[10] ,
    \Tile_X6Y5_NN4BEG[9] ,
    \Tile_X6Y5_NN4BEG[8] ,
    \Tile_X6Y5_NN4BEG[7] ,
    \Tile_X6Y5_NN4BEG[6] ,
    \Tile_X6Y5_NN4BEG[5] ,
    \Tile_X6Y5_NN4BEG[4] ,
    \Tile_X6Y5_NN4BEG[3] ,
    \Tile_X6Y5_NN4BEG[2] ,
    \Tile_X6Y5_NN4BEG[1] ,
    \Tile_X6Y5_NN4BEG[0] }),
    .NN4END({\Tile_X6Y6_NN4BEG[15] ,
    \Tile_X6Y6_NN4BEG[14] ,
    \Tile_X6Y6_NN4BEG[13] ,
    \Tile_X6Y6_NN4BEG[12] ,
    \Tile_X6Y6_NN4BEG[11] ,
    \Tile_X6Y6_NN4BEG[10] ,
    \Tile_X6Y6_NN4BEG[9] ,
    \Tile_X6Y6_NN4BEG[8] ,
    \Tile_X6Y6_NN4BEG[7] ,
    \Tile_X6Y6_NN4BEG[6] ,
    \Tile_X6Y6_NN4BEG[5] ,
    \Tile_X6Y6_NN4BEG[4] ,
    \Tile_X6Y6_NN4BEG[3] ,
    \Tile_X6Y6_NN4BEG[2] ,
    \Tile_X6Y6_NN4BEG[1] ,
    \Tile_X6Y6_NN4BEG[0] }),
    .S1BEG({\Tile_X6Y5_S1BEG[3] ,
    \Tile_X6Y5_S1BEG[2] ,
    \Tile_X6Y5_S1BEG[1] ,
    \Tile_X6Y5_S1BEG[0] }),
    .S1END({\Tile_X6Y4_S1BEG[3] ,
    \Tile_X6Y4_S1BEG[2] ,
    \Tile_X6Y4_S1BEG[1] ,
    \Tile_X6Y4_S1BEG[0] }),
    .S2BEG({\Tile_X6Y5_S2BEG[7] ,
    \Tile_X6Y5_S2BEG[6] ,
    \Tile_X6Y5_S2BEG[5] ,
    \Tile_X6Y5_S2BEG[4] ,
    \Tile_X6Y5_S2BEG[3] ,
    \Tile_X6Y5_S2BEG[2] ,
    \Tile_X6Y5_S2BEG[1] ,
    \Tile_X6Y5_S2BEG[0] }),
    .S2BEGb({\Tile_X6Y5_S2BEGb[7] ,
    \Tile_X6Y5_S2BEGb[6] ,
    \Tile_X6Y5_S2BEGb[5] ,
    \Tile_X6Y5_S2BEGb[4] ,
    \Tile_X6Y5_S2BEGb[3] ,
    \Tile_X6Y5_S2BEGb[2] ,
    \Tile_X6Y5_S2BEGb[1] ,
    \Tile_X6Y5_S2BEGb[0] }),
    .S2END({\Tile_X6Y4_S2BEGb[7] ,
    \Tile_X6Y4_S2BEGb[6] ,
    \Tile_X6Y4_S2BEGb[5] ,
    \Tile_X6Y4_S2BEGb[4] ,
    \Tile_X6Y4_S2BEGb[3] ,
    \Tile_X6Y4_S2BEGb[2] ,
    \Tile_X6Y4_S2BEGb[1] ,
    \Tile_X6Y4_S2BEGb[0] }),
    .S2MID({\Tile_X6Y4_S2BEG[7] ,
    \Tile_X6Y4_S2BEG[6] ,
    \Tile_X6Y4_S2BEG[5] ,
    \Tile_X6Y4_S2BEG[4] ,
    \Tile_X6Y4_S2BEG[3] ,
    \Tile_X6Y4_S2BEG[2] ,
    \Tile_X6Y4_S2BEG[1] ,
    \Tile_X6Y4_S2BEG[0] }),
    .S4BEG({\Tile_X6Y5_S4BEG[15] ,
    \Tile_X6Y5_S4BEG[14] ,
    \Tile_X6Y5_S4BEG[13] ,
    \Tile_X6Y5_S4BEG[12] ,
    \Tile_X6Y5_S4BEG[11] ,
    \Tile_X6Y5_S4BEG[10] ,
    \Tile_X6Y5_S4BEG[9] ,
    \Tile_X6Y5_S4BEG[8] ,
    \Tile_X6Y5_S4BEG[7] ,
    \Tile_X6Y5_S4BEG[6] ,
    \Tile_X6Y5_S4BEG[5] ,
    \Tile_X6Y5_S4BEG[4] ,
    \Tile_X6Y5_S4BEG[3] ,
    \Tile_X6Y5_S4BEG[2] ,
    \Tile_X6Y5_S4BEG[1] ,
    \Tile_X6Y5_S4BEG[0] }),
    .S4END({\Tile_X6Y4_S4BEG[15] ,
    \Tile_X6Y4_S4BEG[14] ,
    \Tile_X6Y4_S4BEG[13] ,
    \Tile_X6Y4_S4BEG[12] ,
    \Tile_X6Y4_S4BEG[11] ,
    \Tile_X6Y4_S4BEG[10] ,
    \Tile_X6Y4_S4BEG[9] ,
    \Tile_X6Y4_S4BEG[8] ,
    \Tile_X6Y4_S4BEG[7] ,
    \Tile_X6Y4_S4BEG[6] ,
    \Tile_X6Y4_S4BEG[5] ,
    \Tile_X6Y4_S4BEG[4] ,
    \Tile_X6Y4_S4BEG[3] ,
    \Tile_X6Y4_S4BEG[2] ,
    \Tile_X6Y4_S4BEG[1] ,
    \Tile_X6Y4_S4BEG[0] }),
    .SS4BEG({\Tile_X6Y5_SS4BEG[15] ,
    \Tile_X6Y5_SS4BEG[14] ,
    \Tile_X6Y5_SS4BEG[13] ,
    \Tile_X6Y5_SS4BEG[12] ,
    \Tile_X6Y5_SS4BEG[11] ,
    \Tile_X6Y5_SS4BEG[10] ,
    \Tile_X6Y5_SS4BEG[9] ,
    \Tile_X6Y5_SS4BEG[8] ,
    \Tile_X6Y5_SS4BEG[7] ,
    \Tile_X6Y5_SS4BEG[6] ,
    \Tile_X6Y5_SS4BEG[5] ,
    \Tile_X6Y5_SS4BEG[4] ,
    \Tile_X6Y5_SS4BEG[3] ,
    \Tile_X6Y5_SS4BEG[2] ,
    \Tile_X6Y5_SS4BEG[1] ,
    \Tile_X6Y5_SS4BEG[0] }),
    .SS4END({\Tile_X6Y4_SS4BEG[15] ,
    \Tile_X6Y4_SS4BEG[14] ,
    \Tile_X6Y4_SS4BEG[13] ,
    \Tile_X6Y4_SS4BEG[12] ,
    \Tile_X6Y4_SS4BEG[11] ,
    \Tile_X6Y4_SS4BEG[10] ,
    \Tile_X6Y4_SS4BEG[9] ,
    \Tile_X6Y4_SS4BEG[8] ,
    \Tile_X6Y4_SS4BEG[7] ,
    \Tile_X6Y4_SS4BEG[6] ,
    \Tile_X6Y4_SS4BEG[5] ,
    \Tile_X6Y4_SS4BEG[4] ,
    \Tile_X6Y4_SS4BEG[3] ,
    \Tile_X6Y4_SS4BEG[2] ,
    \Tile_X6Y4_SS4BEG[1] ,
    \Tile_X6Y4_SS4BEG[0] }),
    .W1BEG({\Tile_X6Y5_W1BEG[3] ,
    \Tile_X6Y5_W1BEG[2] ,
    \Tile_X6Y5_W1BEG[1] ,
    \Tile_X6Y5_W1BEG[0] }),
    .W1END({\Tile_X7Y5_W1BEG[3] ,
    \Tile_X7Y5_W1BEG[2] ,
    \Tile_X7Y5_W1BEG[1] ,
    \Tile_X7Y5_W1BEG[0] }),
    .W2BEG({\Tile_X6Y5_W2BEG[7] ,
    \Tile_X6Y5_W2BEG[6] ,
    \Tile_X6Y5_W2BEG[5] ,
    \Tile_X6Y5_W2BEG[4] ,
    \Tile_X6Y5_W2BEG[3] ,
    \Tile_X6Y5_W2BEG[2] ,
    \Tile_X6Y5_W2BEG[1] ,
    \Tile_X6Y5_W2BEG[0] }),
    .W2BEGb({\Tile_X6Y5_W2BEGb[7] ,
    \Tile_X6Y5_W2BEGb[6] ,
    \Tile_X6Y5_W2BEGb[5] ,
    \Tile_X6Y5_W2BEGb[4] ,
    \Tile_X6Y5_W2BEGb[3] ,
    \Tile_X6Y5_W2BEGb[2] ,
    \Tile_X6Y5_W2BEGb[1] ,
    \Tile_X6Y5_W2BEGb[0] }),
    .W2END({\Tile_X7Y5_W2BEGb[7] ,
    \Tile_X7Y5_W2BEGb[6] ,
    \Tile_X7Y5_W2BEGb[5] ,
    \Tile_X7Y5_W2BEGb[4] ,
    \Tile_X7Y5_W2BEGb[3] ,
    \Tile_X7Y5_W2BEGb[2] ,
    \Tile_X7Y5_W2BEGb[1] ,
    \Tile_X7Y5_W2BEGb[0] }),
    .W2MID({\Tile_X7Y5_W2BEG[7] ,
    \Tile_X7Y5_W2BEG[6] ,
    \Tile_X7Y5_W2BEG[5] ,
    \Tile_X7Y5_W2BEG[4] ,
    \Tile_X7Y5_W2BEG[3] ,
    \Tile_X7Y5_W2BEG[2] ,
    \Tile_X7Y5_W2BEG[1] ,
    \Tile_X7Y5_W2BEG[0] }),
    .W6BEG({\Tile_X6Y5_W6BEG[11] ,
    \Tile_X6Y5_W6BEG[10] ,
    \Tile_X6Y5_W6BEG[9] ,
    \Tile_X6Y5_W6BEG[8] ,
    \Tile_X6Y5_W6BEG[7] ,
    \Tile_X6Y5_W6BEG[6] ,
    \Tile_X6Y5_W6BEG[5] ,
    \Tile_X6Y5_W6BEG[4] ,
    \Tile_X6Y5_W6BEG[3] ,
    \Tile_X6Y5_W6BEG[2] ,
    \Tile_X6Y5_W6BEG[1] ,
    \Tile_X6Y5_W6BEG[0] }),
    .W6END({\Tile_X7Y5_W6BEG[11] ,
    \Tile_X7Y5_W6BEG[10] ,
    \Tile_X7Y5_W6BEG[9] ,
    \Tile_X7Y5_W6BEG[8] ,
    \Tile_X7Y5_W6BEG[7] ,
    \Tile_X7Y5_W6BEG[6] ,
    \Tile_X7Y5_W6BEG[5] ,
    \Tile_X7Y5_W6BEG[4] ,
    \Tile_X7Y5_W6BEG[3] ,
    \Tile_X7Y5_W6BEG[2] ,
    \Tile_X7Y5_W6BEG[1] ,
    \Tile_X7Y5_W6BEG[0] }),
    .WW4BEG({\Tile_X6Y5_WW4BEG[15] ,
    \Tile_X6Y5_WW4BEG[14] ,
    \Tile_X6Y5_WW4BEG[13] ,
    \Tile_X6Y5_WW4BEG[12] ,
    \Tile_X6Y5_WW4BEG[11] ,
    \Tile_X6Y5_WW4BEG[10] ,
    \Tile_X6Y5_WW4BEG[9] ,
    \Tile_X6Y5_WW4BEG[8] ,
    \Tile_X6Y5_WW4BEG[7] ,
    \Tile_X6Y5_WW4BEG[6] ,
    \Tile_X6Y5_WW4BEG[5] ,
    \Tile_X6Y5_WW4BEG[4] ,
    \Tile_X6Y5_WW4BEG[3] ,
    \Tile_X6Y5_WW4BEG[2] ,
    \Tile_X6Y5_WW4BEG[1] ,
    \Tile_X6Y5_WW4BEG[0] }),
    .WW4END({\Tile_X7Y5_WW4BEG[15] ,
    \Tile_X7Y5_WW4BEG[14] ,
    \Tile_X7Y5_WW4BEG[13] ,
    \Tile_X7Y5_WW4BEG[12] ,
    \Tile_X7Y5_WW4BEG[11] ,
    \Tile_X7Y5_WW4BEG[10] ,
    \Tile_X7Y5_WW4BEG[9] ,
    \Tile_X7Y5_WW4BEG[8] ,
    \Tile_X7Y5_WW4BEG[7] ,
    \Tile_X7Y5_WW4BEG[6] ,
    \Tile_X7Y5_WW4BEG[5] ,
    \Tile_X7Y5_WW4BEG[4] ,
    \Tile_X7Y5_WW4BEG[3] ,
    \Tile_X7Y5_WW4BEG[2] ,
    \Tile_X7Y5_WW4BEG[1] ,
    \Tile_X7Y5_WW4BEG[0] }));
 LUT4AB Tile_X6Y6_LUT4AB (.Ci(Tile_X6Y7_Co),
    .Co(Tile_X6Y6_Co),
    .UserCLK(Tile_X6Y7_UserCLKo),
    .UserCLKo(Tile_X6Y6_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X6Y6_E1BEG[3] ,
    \Tile_X6Y6_E1BEG[2] ,
    \Tile_X6Y6_E1BEG[1] ,
    \Tile_X6Y6_E1BEG[0] }),
    .E1END({\Tile_X5Y6_E1BEG[3] ,
    \Tile_X5Y6_E1BEG[2] ,
    \Tile_X5Y6_E1BEG[1] ,
    \Tile_X5Y6_E1BEG[0] }),
    .E2BEG({\Tile_X6Y6_E2BEG[7] ,
    \Tile_X6Y6_E2BEG[6] ,
    \Tile_X6Y6_E2BEG[5] ,
    \Tile_X6Y6_E2BEG[4] ,
    \Tile_X6Y6_E2BEG[3] ,
    \Tile_X6Y6_E2BEG[2] ,
    \Tile_X6Y6_E2BEG[1] ,
    \Tile_X6Y6_E2BEG[0] }),
    .E2BEGb({\Tile_X6Y6_E2BEGb[7] ,
    \Tile_X6Y6_E2BEGb[6] ,
    \Tile_X6Y6_E2BEGb[5] ,
    \Tile_X6Y6_E2BEGb[4] ,
    \Tile_X6Y6_E2BEGb[3] ,
    \Tile_X6Y6_E2BEGb[2] ,
    \Tile_X6Y6_E2BEGb[1] ,
    \Tile_X6Y6_E2BEGb[0] }),
    .E2END({\Tile_X5Y6_E2BEGb[7] ,
    \Tile_X5Y6_E2BEGb[6] ,
    \Tile_X5Y6_E2BEGb[5] ,
    \Tile_X5Y6_E2BEGb[4] ,
    \Tile_X5Y6_E2BEGb[3] ,
    \Tile_X5Y6_E2BEGb[2] ,
    \Tile_X5Y6_E2BEGb[1] ,
    \Tile_X5Y6_E2BEGb[0] }),
    .E2MID({\Tile_X5Y6_E2BEG[7] ,
    \Tile_X5Y6_E2BEG[6] ,
    \Tile_X5Y6_E2BEG[5] ,
    \Tile_X5Y6_E2BEG[4] ,
    \Tile_X5Y6_E2BEG[3] ,
    \Tile_X5Y6_E2BEG[2] ,
    \Tile_X5Y6_E2BEG[1] ,
    \Tile_X5Y6_E2BEG[0] }),
    .E6BEG({\Tile_X6Y6_E6BEG[11] ,
    \Tile_X6Y6_E6BEG[10] ,
    \Tile_X6Y6_E6BEG[9] ,
    \Tile_X6Y6_E6BEG[8] ,
    \Tile_X6Y6_E6BEG[7] ,
    \Tile_X6Y6_E6BEG[6] ,
    \Tile_X6Y6_E6BEG[5] ,
    \Tile_X6Y6_E6BEG[4] ,
    \Tile_X6Y6_E6BEG[3] ,
    \Tile_X6Y6_E6BEG[2] ,
    \Tile_X6Y6_E6BEG[1] ,
    \Tile_X6Y6_E6BEG[0] }),
    .E6END({\Tile_X5Y6_E6BEG[11] ,
    \Tile_X5Y6_E6BEG[10] ,
    \Tile_X5Y6_E6BEG[9] ,
    \Tile_X5Y6_E6BEG[8] ,
    \Tile_X5Y6_E6BEG[7] ,
    \Tile_X5Y6_E6BEG[6] ,
    \Tile_X5Y6_E6BEG[5] ,
    \Tile_X5Y6_E6BEG[4] ,
    \Tile_X5Y6_E6BEG[3] ,
    \Tile_X5Y6_E6BEG[2] ,
    \Tile_X5Y6_E6BEG[1] ,
    \Tile_X5Y6_E6BEG[0] }),
    .EE4BEG({\Tile_X6Y6_EE4BEG[15] ,
    \Tile_X6Y6_EE4BEG[14] ,
    \Tile_X6Y6_EE4BEG[13] ,
    \Tile_X6Y6_EE4BEG[12] ,
    \Tile_X6Y6_EE4BEG[11] ,
    \Tile_X6Y6_EE4BEG[10] ,
    \Tile_X6Y6_EE4BEG[9] ,
    \Tile_X6Y6_EE4BEG[8] ,
    \Tile_X6Y6_EE4BEG[7] ,
    \Tile_X6Y6_EE4BEG[6] ,
    \Tile_X6Y6_EE4BEG[5] ,
    \Tile_X6Y6_EE4BEG[4] ,
    \Tile_X6Y6_EE4BEG[3] ,
    \Tile_X6Y6_EE4BEG[2] ,
    \Tile_X6Y6_EE4BEG[1] ,
    \Tile_X6Y6_EE4BEG[0] }),
    .EE4END({\Tile_X5Y6_EE4BEG[15] ,
    \Tile_X5Y6_EE4BEG[14] ,
    \Tile_X5Y6_EE4BEG[13] ,
    \Tile_X5Y6_EE4BEG[12] ,
    \Tile_X5Y6_EE4BEG[11] ,
    \Tile_X5Y6_EE4BEG[10] ,
    \Tile_X5Y6_EE4BEG[9] ,
    \Tile_X5Y6_EE4BEG[8] ,
    \Tile_X5Y6_EE4BEG[7] ,
    \Tile_X5Y6_EE4BEG[6] ,
    \Tile_X5Y6_EE4BEG[5] ,
    \Tile_X5Y6_EE4BEG[4] ,
    \Tile_X5Y6_EE4BEG[3] ,
    \Tile_X5Y6_EE4BEG[2] ,
    \Tile_X5Y6_EE4BEG[1] ,
    \Tile_X5Y6_EE4BEG[0] }),
    .FrameData({\Tile_X5Y6_FrameData_O[31] ,
    \Tile_X5Y6_FrameData_O[30] ,
    \Tile_X5Y6_FrameData_O[29] ,
    \Tile_X5Y6_FrameData_O[28] ,
    \Tile_X5Y6_FrameData_O[27] ,
    \Tile_X5Y6_FrameData_O[26] ,
    \Tile_X5Y6_FrameData_O[25] ,
    \Tile_X5Y6_FrameData_O[24] ,
    \Tile_X5Y6_FrameData_O[23] ,
    \Tile_X5Y6_FrameData_O[22] ,
    \Tile_X5Y6_FrameData_O[21] ,
    \Tile_X5Y6_FrameData_O[20] ,
    \Tile_X5Y6_FrameData_O[19] ,
    \Tile_X5Y6_FrameData_O[18] ,
    \Tile_X5Y6_FrameData_O[17] ,
    \Tile_X5Y6_FrameData_O[16] ,
    \Tile_X5Y6_FrameData_O[15] ,
    \Tile_X5Y6_FrameData_O[14] ,
    \Tile_X5Y6_FrameData_O[13] ,
    \Tile_X5Y6_FrameData_O[12] ,
    \Tile_X5Y6_FrameData_O[11] ,
    \Tile_X5Y6_FrameData_O[10] ,
    \Tile_X5Y6_FrameData_O[9] ,
    \Tile_X5Y6_FrameData_O[8] ,
    \Tile_X5Y6_FrameData_O[7] ,
    \Tile_X5Y6_FrameData_O[6] ,
    \Tile_X5Y6_FrameData_O[5] ,
    \Tile_X5Y6_FrameData_O[4] ,
    \Tile_X5Y6_FrameData_O[3] ,
    \Tile_X5Y6_FrameData_O[2] ,
    \Tile_X5Y6_FrameData_O[1] ,
    \Tile_X5Y6_FrameData_O[0] }),
    .FrameData_O({\Tile_X6Y6_FrameData_O[31] ,
    \Tile_X6Y6_FrameData_O[30] ,
    \Tile_X6Y6_FrameData_O[29] ,
    \Tile_X6Y6_FrameData_O[28] ,
    \Tile_X6Y6_FrameData_O[27] ,
    \Tile_X6Y6_FrameData_O[26] ,
    \Tile_X6Y6_FrameData_O[25] ,
    \Tile_X6Y6_FrameData_O[24] ,
    \Tile_X6Y6_FrameData_O[23] ,
    \Tile_X6Y6_FrameData_O[22] ,
    \Tile_X6Y6_FrameData_O[21] ,
    \Tile_X6Y6_FrameData_O[20] ,
    \Tile_X6Y6_FrameData_O[19] ,
    \Tile_X6Y6_FrameData_O[18] ,
    \Tile_X6Y6_FrameData_O[17] ,
    \Tile_X6Y6_FrameData_O[16] ,
    \Tile_X6Y6_FrameData_O[15] ,
    \Tile_X6Y6_FrameData_O[14] ,
    \Tile_X6Y6_FrameData_O[13] ,
    \Tile_X6Y6_FrameData_O[12] ,
    \Tile_X6Y6_FrameData_O[11] ,
    \Tile_X6Y6_FrameData_O[10] ,
    \Tile_X6Y6_FrameData_O[9] ,
    \Tile_X6Y6_FrameData_O[8] ,
    \Tile_X6Y6_FrameData_O[7] ,
    \Tile_X6Y6_FrameData_O[6] ,
    \Tile_X6Y6_FrameData_O[5] ,
    \Tile_X6Y6_FrameData_O[4] ,
    \Tile_X6Y6_FrameData_O[3] ,
    \Tile_X6Y6_FrameData_O[2] ,
    \Tile_X6Y6_FrameData_O[1] ,
    \Tile_X6Y6_FrameData_O[0] }),
    .FrameStrobe({\Tile_X6Y7_FrameStrobe_O[19] ,
    \Tile_X6Y7_FrameStrobe_O[18] ,
    \Tile_X6Y7_FrameStrobe_O[17] ,
    \Tile_X6Y7_FrameStrobe_O[16] ,
    \Tile_X6Y7_FrameStrobe_O[15] ,
    \Tile_X6Y7_FrameStrobe_O[14] ,
    \Tile_X6Y7_FrameStrobe_O[13] ,
    \Tile_X6Y7_FrameStrobe_O[12] ,
    \Tile_X6Y7_FrameStrobe_O[11] ,
    \Tile_X6Y7_FrameStrobe_O[10] ,
    \Tile_X6Y7_FrameStrobe_O[9] ,
    \Tile_X6Y7_FrameStrobe_O[8] ,
    \Tile_X6Y7_FrameStrobe_O[7] ,
    \Tile_X6Y7_FrameStrobe_O[6] ,
    \Tile_X6Y7_FrameStrobe_O[5] ,
    \Tile_X6Y7_FrameStrobe_O[4] ,
    \Tile_X6Y7_FrameStrobe_O[3] ,
    \Tile_X6Y7_FrameStrobe_O[2] ,
    \Tile_X6Y7_FrameStrobe_O[1] ,
    \Tile_X6Y7_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X6Y6_FrameStrobe_O[19] ,
    \Tile_X6Y6_FrameStrobe_O[18] ,
    \Tile_X6Y6_FrameStrobe_O[17] ,
    \Tile_X6Y6_FrameStrobe_O[16] ,
    \Tile_X6Y6_FrameStrobe_O[15] ,
    \Tile_X6Y6_FrameStrobe_O[14] ,
    \Tile_X6Y6_FrameStrobe_O[13] ,
    \Tile_X6Y6_FrameStrobe_O[12] ,
    \Tile_X6Y6_FrameStrobe_O[11] ,
    \Tile_X6Y6_FrameStrobe_O[10] ,
    \Tile_X6Y6_FrameStrobe_O[9] ,
    \Tile_X6Y6_FrameStrobe_O[8] ,
    \Tile_X6Y6_FrameStrobe_O[7] ,
    \Tile_X6Y6_FrameStrobe_O[6] ,
    \Tile_X6Y6_FrameStrobe_O[5] ,
    \Tile_X6Y6_FrameStrobe_O[4] ,
    \Tile_X6Y6_FrameStrobe_O[3] ,
    \Tile_X6Y6_FrameStrobe_O[2] ,
    \Tile_X6Y6_FrameStrobe_O[1] ,
    \Tile_X6Y6_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X6Y6_N1BEG[3] ,
    \Tile_X6Y6_N1BEG[2] ,
    \Tile_X6Y6_N1BEG[1] ,
    \Tile_X6Y6_N1BEG[0] }),
    .N1END({\Tile_X6Y7_N1BEG[3] ,
    \Tile_X6Y7_N1BEG[2] ,
    \Tile_X6Y7_N1BEG[1] ,
    \Tile_X6Y7_N1BEG[0] }),
    .N2BEG({\Tile_X6Y6_N2BEG[7] ,
    \Tile_X6Y6_N2BEG[6] ,
    \Tile_X6Y6_N2BEG[5] ,
    \Tile_X6Y6_N2BEG[4] ,
    \Tile_X6Y6_N2BEG[3] ,
    \Tile_X6Y6_N2BEG[2] ,
    \Tile_X6Y6_N2BEG[1] ,
    \Tile_X6Y6_N2BEG[0] }),
    .N2BEGb({\Tile_X6Y6_N2BEGb[7] ,
    \Tile_X6Y6_N2BEGb[6] ,
    \Tile_X6Y6_N2BEGb[5] ,
    \Tile_X6Y6_N2BEGb[4] ,
    \Tile_X6Y6_N2BEGb[3] ,
    \Tile_X6Y6_N2BEGb[2] ,
    \Tile_X6Y6_N2BEGb[1] ,
    \Tile_X6Y6_N2BEGb[0] }),
    .N2END({\Tile_X6Y7_N2BEGb[7] ,
    \Tile_X6Y7_N2BEGb[6] ,
    \Tile_X6Y7_N2BEGb[5] ,
    \Tile_X6Y7_N2BEGb[4] ,
    \Tile_X6Y7_N2BEGb[3] ,
    \Tile_X6Y7_N2BEGb[2] ,
    \Tile_X6Y7_N2BEGb[1] ,
    \Tile_X6Y7_N2BEGb[0] }),
    .N2MID({\Tile_X6Y7_N2BEG[7] ,
    \Tile_X6Y7_N2BEG[6] ,
    \Tile_X6Y7_N2BEG[5] ,
    \Tile_X6Y7_N2BEG[4] ,
    \Tile_X6Y7_N2BEG[3] ,
    \Tile_X6Y7_N2BEG[2] ,
    \Tile_X6Y7_N2BEG[1] ,
    \Tile_X6Y7_N2BEG[0] }),
    .N4BEG({\Tile_X6Y6_N4BEG[15] ,
    \Tile_X6Y6_N4BEG[14] ,
    \Tile_X6Y6_N4BEG[13] ,
    \Tile_X6Y6_N4BEG[12] ,
    \Tile_X6Y6_N4BEG[11] ,
    \Tile_X6Y6_N4BEG[10] ,
    \Tile_X6Y6_N4BEG[9] ,
    \Tile_X6Y6_N4BEG[8] ,
    \Tile_X6Y6_N4BEG[7] ,
    \Tile_X6Y6_N4BEG[6] ,
    \Tile_X6Y6_N4BEG[5] ,
    \Tile_X6Y6_N4BEG[4] ,
    \Tile_X6Y6_N4BEG[3] ,
    \Tile_X6Y6_N4BEG[2] ,
    \Tile_X6Y6_N4BEG[1] ,
    \Tile_X6Y6_N4BEG[0] }),
    .N4END({\Tile_X6Y7_N4BEG[15] ,
    \Tile_X6Y7_N4BEG[14] ,
    \Tile_X6Y7_N4BEG[13] ,
    \Tile_X6Y7_N4BEG[12] ,
    \Tile_X6Y7_N4BEG[11] ,
    \Tile_X6Y7_N4BEG[10] ,
    \Tile_X6Y7_N4BEG[9] ,
    \Tile_X6Y7_N4BEG[8] ,
    \Tile_X6Y7_N4BEG[7] ,
    \Tile_X6Y7_N4BEG[6] ,
    \Tile_X6Y7_N4BEG[5] ,
    \Tile_X6Y7_N4BEG[4] ,
    \Tile_X6Y7_N4BEG[3] ,
    \Tile_X6Y7_N4BEG[2] ,
    \Tile_X6Y7_N4BEG[1] ,
    \Tile_X6Y7_N4BEG[0] }),
    .NN4BEG({\Tile_X6Y6_NN4BEG[15] ,
    \Tile_X6Y6_NN4BEG[14] ,
    \Tile_X6Y6_NN4BEG[13] ,
    \Tile_X6Y6_NN4BEG[12] ,
    \Tile_X6Y6_NN4BEG[11] ,
    \Tile_X6Y6_NN4BEG[10] ,
    \Tile_X6Y6_NN4BEG[9] ,
    \Tile_X6Y6_NN4BEG[8] ,
    \Tile_X6Y6_NN4BEG[7] ,
    \Tile_X6Y6_NN4BEG[6] ,
    \Tile_X6Y6_NN4BEG[5] ,
    \Tile_X6Y6_NN4BEG[4] ,
    \Tile_X6Y6_NN4BEG[3] ,
    \Tile_X6Y6_NN4BEG[2] ,
    \Tile_X6Y6_NN4BEG[1] ,
    \Tile_X6Y6_NN4BEG[0] }),
    .NN4END({\Tile_X6Y7_NN4BEG[15] ,
    \Tile_X6Y7_NN4BEG[14] ,
    \Tile_X6Y7_NN4BEG[13] ,
    \Tile_X6Y7_NN4BEG[12] ,
    \Tile_X6Y7_NN4BEG[11] ,
    \Tile_X6Y7_NN4BEG[10] ,
    \Tile_X6Y7_NN4BEG[9] ,
    \Tile_X6Y7_NN4BEG[8] ,
    \Tile_X6Y7_NN4BEG[7] ,
    \Tile_X6Y7_NN4BEG[6] ,
    \Tile_X6Y7_NN4BEG[5] ,
    \Tile_X6Y7_NN4BEG[4] ,
    \Tile_X6Y7_NN4BEG[3] ,
    \Tile_X6Y7_NN4BEG[2] ,
    \Tile_X6Y7_NN4BEG[1] ,
    \Tile_X6Y7_NN4BEG[0] }),
    .S1BEG({\Tile_X6Y6_S1BEG[3] ,
    \Tile_X6Y6_S1BEG[2] ,
    \Tile_X6Y6_S1BEG[1] ,
    \Tile_X6Y6_S1BEG[0] }),
    .S1END({\Tile_X6Y5_S1BEG[3] ,
    \Tile_X6Y5_S1BEG[2] ,
    \Tile_X6Y5_S1BEG[1] ,
    \Tile_X6Y5_S1BEG[0] }),
    .S2BEG({\Tile_X6Y6_S2BEG[7] ,
    \Tile_X6Y6_S2BEG[6] ,
    \Tile_X6Y6_S2BEG[5] ,
    \Tile_X6Y6_S2BEG[4] ,
    \Tile_X6Y6_S2BEG[3] ,
    \Tile_X6Y6_S2BEG[2] ,
    \Tile_X6Y6_S2BEG[1] ,
    \Tile_X6Y6_S2BEG[0] }),
    .S2BEGb({\Tile_X6Y6_S2BEGb[7] ,
    \Tile_X6Y6_S2BEGb[6] ,
    \Tile_X6Y6_S2BEGb[5] ,
    \Tile_X6Y6_S2BEGb[4] ,
    \Tile_X6Y6_S2BEGb[3] ,
    \Tile_X6Y6_S2BEGb[2] ,
    \Tile_X6Y6_S2BEGb[1] ,
    \Tile_X6Y6_S2BEGb[0] }),
    .S2END({\Tile_X6Y5_S2BEGb[7] ,
    \Tile_X6Y5_S2BEGb[6] ,
    \Tile_X6Y5_S2BEGb[5] ,
    \Tile_X6Y5_S2BEGb[4] ,
    \Tile_X6Y5_S2BEGb[3] ,
    \Tile_X6Y5_S2BEGb[2] ,
    \Tile_X6Y5_S2BEGb[1] ,
    \Tile_X6Y5_S2BEGb[0] }),
    .S2MID({\Tile_X6Y5_S2BEG[7] ,
    \Tile_X6Y5_S2BEG[6] ,
    \Tile_X6Y5_S2BEG[5] ,
    \Tile_X6Y5_S2BEG[4] ,
    \Tile_X6Y5_S2BEG[3] ,
    \Tile_X6Y5_S2BEG[2] ,
    \Tile_X6Y5_S2BEG[1] ,
    \Tile_X6Y5_S2BEG[0] }),
    .S4BEG({\Tile_X6Y6_S4BEG[15] ,
    \Tile_X6Y6_S4BEG[14] ,
    \Tile_X6Y6_S4BEG[13] ,
    \Tile_X6Y6_S4BEG[12] ,
    \Tile_X6Y6_S4BEG[11] ,
    \Tile_X6Y6_S4BEG[10] ,
    \Tile_X6Y6_S4BEG[9] ,
    \Tile_X6Y6_S4BEG[8] ,
    \Tile_X6Y6_S4BEG[7] ,
    \Tile_X6Y6_S4BEG[6] ,
    \Tile_X6Y6_S4BEG[5] ,
    \Tile_X6Y6_S4BEG[4] ,
    \Tile_X6Y6_S4BEG[3] ,
    \Tile_X6Y6_S4BEG[2] ,
    \Tile_X6Y6_S4BEG[1] ,
    \Tile_X6Y6_S4BEG[0] }),
    .S4END({\Tile_X6Y5_S4BEG[15] ,
    \Tile_X6Y5_S4BEG[14] ,
    \Tile_X6Y5_S4BEG[13] ,
    \Tile_X6Y5_S4BEG[12] ,
    \Tile_X6Y5_S4BEG[11] ,
    \Tile_X6Y5_S4BEG[10] ,
    \Tile_X6Y5_S4BEG[9] ,
    \Tile_X6Y5_S4BEG[8] ,
    \Tile_X6Y5_S4BEG[7] ,
    \Tile_X6Y5_S4BEG[6] ,
    \Tile_X6Y5_S4BEG[5] ,
    \Tile_X6Y5_S4BEG[4] ,
    \Tile_X6Y5_S4BEG[3] ,
    \Tile_X6Y5_S4BEG[2] ,
    \Tile_X6Y5_S4BEG[1] ,
    \Tile_X6Y5_S4BEG[0] }),
    .SS4BEG({\Tile_X6Y6_SS4BEG[15] ,
    \Tile_X6Y6_SS4BEG[14] ,
    \Tile_X6Y6_SS4BEG[13] ,
    \Tile_X6Y6_SS4BEG[12] ,
    \Tile_X6Y6_SS4BEG[11] ,
    \Tile_X6Y6_SS4BEG[10] ,
    \Tile_X6Y6_SS4BEG[9] ,
    \Tile_X6Y6_SS4BEG[8] ,
    \Tile_X6Y6_SS4BEG[7] ,
    \Tile_X6Y6_SS4BEG[6] ,
    \Tile_X6Y6_SS4BEG[5] ,
    \Tile_X6Y6_SS4BEG[4] ,
    \Tile_X6Y6_SS4BEG[3] ,
    \Tile_X6Y6_SS4BEG[2] ,
    \Tile_X6Y6_SS4BEG[1] ,
    \Tile_X6Y6_SS4BEG[0] }),
    .SS4END({\Tile_X6Y5_SS4BEG[15] ,
    \Tile_X6Y5_SS4BEG[14] ,
    \Tile_X6Y5_SS4BEG[13] ,
    \Tile_X6Y5_SS4BEG[12] ,
    \Tile_X6Y5_SS4BEG[11] ,
    \Tile_X6Y5_SS4BEG[10] ,
    \Tile_X6Y5_SS4BEG[9] ,
    \Tile_X6Y5_SS4BEG[8] ,
    \Tile_X6Y5_SS4BEG[7] ,
    \Tile_X6Y5_SS4BEG[6] ,
    \Tile_X6Y5_SS4BEG[5] ,
    \Tile_X6Y5_SS4BEG[4] ,
    \Tile_X6Y5_SS4BEG[3] ,
    \Tile_X6Y5_SS4BEG[2] ,
    \Tile_X6Y5_SS4BEG[1] ,
    \Tile_X6Y5_SS4BEG[0] }),
    .W1BEG({\Tile_X6Y6_W1BEG[3] ,
    \Tile_X6Y6_W1BEG[2] ,
    \Tile_X6Y6_W1BEG[1] ,
    \Tile_X6Y6_W1BEG[0] }),
    .W1END({\Tile_X7Y6_W1BEG[3] ,
    \Tile_X7Y6_W1BEG[2] ,
    \Tile_X7Y6_W1BEG[1] ,
    \Tile_X7Y6_W1BEG[0] }),
    .W2BEG({\Tile_X6Y6_W2BEG[7] ,
    \Tile_X6Y6_W2BEG[6] ,
    \Tile_X6Y6_W2BEG[5] ,
    \Tile_X6Y6_W2BEG[4] ,
    \Tile_X6Y6_W2BEG[3] ,
    \Tile_X6Y6_W2BEG[2] ,
    \Tile_X6Y6_W2BEG[1] ,
    \Tile_X6Y6_W2BEG[0] }),
    .W2BEGb({\Tile_X6Y6_W2BEGb[7] ,
    \Tile_X6Y6_W2BEGb[6] ,
    \Tile_X6Y6_W2BEGb[5] ,
    \Tile_X6Y6_W2BEGb[4] ,
    \Tile_X6Y6_W2BEGb[3] ,
    \Tile_X6Y6_W2BEGb[2] ,
    \Tile_X6Y6_W2BEGb[1] ,
    \Tile_X6Y6_W2BEGb[0] }),
    .W2END({\Tile_X7Y6_W2BEGb[7] ,
    \Tile_X7Y6_W2BEGb[6] ,
    \Tile_X7Y6_W2BEGb[5] ,
    \Tile_X7Y6_W2BEGb[4] ,
    \Tile_X7Y6_W2BEGb[3] ,
    \Tile_X7Y6_W2BEGb[2] ,
    \Tile_X7Y6_W2BEGb[1] ,
    \Tile_X7Y6_W2BEGb[0] }),
    .W2MID({\Tile_X7Y6_W2BEG[7] ,
    \Tile_X7Y6_W2BEG[6] ,
    \Tile_X7Y6_W2BEG[5] ,
    \Tile_X7Y6_W2BEG[4] ,
    \Tile_X7Y6_W2BEG[3] ,
    \Tile_X7Y6_W2BEG[2] ,
    \Tile_X7Y6_W2BEG[1] ,
    \Tile_X7Y6_W2BEG[0] }),
    .W6BEG({\Tile_X6Y6_W6BEG[11] ,
    \Tile_X6Y6_W6BEG[10] ,
    \Tile_X6Y6_W6BEG[9] ,
    \Tile_X6Y6_W6BEG[8] ,
    \Tile_X6Y6_W6BEG[7] ,
    \Tile_X6Y6_W6BEG[6] ,
    \Tile_X6Y6_W6BEG[5] ,
    \Tile_X6Y6_W6BEG[4] ,
    \Tile_X6Y6_W6BEG[3] ,
    \Tile_X6Y6_W6BEG[2] ,
    \Tile_X6Y6_W6BEG[1] ,
    \Tile_X6Y6_W6BEG[0] }),
    .W6END({\Tile_X7Y6_W6BEG[11] ,
    \Tile_X7Y6_W6BEG[10] ,
    \Tile_X7Y6_W6BEG[9] ,
    \Tile_X7Y6_W6BEG[8] ,
    \Tile_X7Y6_W6BEG[7] ,
    \Tile_X7Y6_W6BEG[6] ,
    \Tile_X7Y6_W6BEG[5] ,
    \Tile_X7Y6_W6BEG[4] ,
    \Tile_X7Y6_W6BEG[3] ,
    \Tile_X7Y6_W6BEG[2] ,
    \Tile_X7Y6_W6BEG[1] ,
    \Tile_X7Y6_W6BEG[0] }),
    .WW4BEG({\Tile_X6Y6_WW4BEG[15] ,
    \Tile_X6Y6_WW4BEG[14] ,
    \Tile_X6Y6_WW4BEG[13] ,
    \Tile_X6Y6_WW4BEG[12] ,
    \Tile_X6Y6_WW4BEG[11] ,
    \Tile_X6Y6_WW4BEG[10] ,
    \Tile_X6Y6_WW4BEG[9] ,
    \Tile_X6Y6_WW4BEG[8] ,
    \Tile_X6Y6_WW4BEG[7] ,
    \Tile_X6Y6_WW4BEG[6] ,
    \Tile_X6Y6_WW4BEG[5] ,
    \Tile_X6Y6_WW4BEG[4] ,
    \Tile_X6Y6_WW4BEG[3] ,
    \Tile_X6Y6_WW4BEG[2] ,
    \Tile_X6Y6_WW4BEG[1] ,
    \Tile_X6Y6_WW4BEG[0] }),
    .WW4END({\Tile_X7Y6_WW4BEG[15] ,
    \Tile_X7Y6_WW4BEG[14] ,
    \Tile_X7Y6_WW4BEG[13] ,
    \Tile_X7Y6_WW4BEG[12] ,
    \Tile_X7Y6_WW4BEG[11] ,
    \Tile_X7Y6_WW4BEG[10] ,
    \Tile_X7Y6_WW4BEG[9] ,
    \Tile_X7Y6_WW4BEG[8] ,
    \Tile_X7Y6_WW4BEG[7] ,
    \Tile_X7Y6_WW4BEG[6] ,
    \Tile_X7Y6_WW4BEG[5] ,
    \Tile_X7Y6_WW4BEG[4] ,
    \Tile_X7Y6_WW4BEG[3] ,
    \Tile_X7Y6_WW4BEG[2] ,
    \Tile_X7Y6_WW4BEG[1] ,
    \Tile_X7Y6_WW4BEG[0] }));
 LUT4AB Tile_X6Y7_LUT4AB (.Ci(Tile_X6Y8_Co),
    .Co(Tile_X6Y7_Co),
    .UserCLK(Tile_X6Y8_UserCLKo),
    .UserCLKo(Tile_X6Y7_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X6Y7_E1BEG[3] ,
    \Tile_X6Y7_E1BEG[2] ,
    \Tile_X6Y7_E1BEG[1] ,
    \Tile_X6Y7_E1BEG[0] }),
    .E1END({\Tile_X5Y7_E1BEG[3] ,
    \Tile_X5Y7_E1BEG[2] ,
    \Tile_X5Y7_E1BEG[1] ,
    \Tile_X5Y7_E1BEG[0] }),
    .E2BEG({\Tile_X6Y7_E2BEG[7] ,
    \Tile_X6Y7_E2BEG[6] ,
    \Tile_X6Y7_E2BEG[5] ,
    \Tile_X6Y7_E2BEG[4] ,
    \Tile_X6Y7_E2BEG[3] ,
    \Tile_X6Y7_E2BEG[2] ,
    \Tile_X6Y7_E2BEG[1] ,
    \Tile_X6Y7_E2BEG[0] }),
    .E2BEGb({\Tile_X6Y7_E2BEGb[7] ,
    \Tile_X6Y7_E2BEGb[6] ,
    \Tile_X6Y7_E2BEGb[5] ,
    \Tile_X6Y7_E2BEGb[4] ,
    \Tile_X6Y7_E2BEGb[3] ,
    \Tile_X6Y7_E2BEGb[2] ,
    \Tile_X6Y7_E2BEGb[1] ,
    \Tile_X6Y7_E2BEGb[0] }),
    .E2END({\Tile_X5Y7_E2BEGb[7] ,
    \Tile_X5Y7_E2BEGb[6] ,
    \Tile_X5Y7_E2BEGb[5] ,
    \Tile_X5Y7_E2BEGb[4] ,
    \Tile_X5Y7_E2BEGb[3] ,
    \Tile_X5Y7_E2BEGb[2] ,
    \Tile_X5Y7_E2BEGb[1] ,
    \Tile_X5Y7_E2BEGb[0] }),
    .E2MID({\Tile_X5Y7_E2BEG[7] ,
    \Tile_X5Y7_E2BEG[6] ,
    \Tile_X5Y7_E2BEG[5] ,
    \Tile_X5Y7_E2BEG[4] ,
    \Tile_X5Y7_E2BEG[3] ,
    \Tile_X5Y7_E2BEG[2] ,
    \Tile_X5Y7_E2BEG[1] ,
    \Tile_X5Y7_E2BEG[0] }),
    .E6BEG({\Tile_X6Y7_E6BEG[11] ,
    \Tile_X6Y7_E6BEG[10] ,
    \Tile_X6Y7_E6BEG[9] ,
    \Tile_X6Y7_E6BEG[8] ,
    \Tile_X6Y7_E6BEG[7] ,
    \Tile_X6Y7_E6BEG[6] ,
    \Tile_X6Y7_E6BEG[5] ,
    \Tile_X6Y7_E6BEG[4] ,
    \Tile_X6Y7_E6BEG[3] ,
    \Tile_X6Y7_E6BEG[2] ,
    \Tile_X6Y7_E6BEG[1] ,
    \Tile_X6Y7_E6BEG[0] }),
    .E6END({\Tile_X5Y7_E6BEG[11] ,
    \Tile_X5Y7_E6BEG[10] ,
    \Tile_X5Y7_E6BEG[9] ,
    \Tile_X5Y7_E6BEG[8] ,
    \Tile_X5Y7_E6BEG[7] ,
    \Tile_X5Y7_E6BEG[6] ,
    \Tile_X5Y7_E6BEG[5] ,
    \Tile_X5Y7_E6BEG[4] ,
    \Tile_X5Y7_E6BEG[3] ,
    \Tile_X5Y7_E6BEG[2] ,
    \Tile_X5Y7_E6BEG[1] ,
    \Tile_X5Y7_E6BEG[0] }),
    .EE4BEG({\Tile_X6Y7_EE4BEG[15] ,
    \Tile_X6Y7_EE4BEG[14] ,
    \Tile_X6Y7_EE4BEG[13] ,
    \Tile_X6Y7_EE4BEG[12] ,
    \Tile_X6Y7_EE4BEG[11] ,
    \Tile_X6Y7_EE4BEG[10] ,
    \Tile_X6Y7_EE4BEG[9] ,
    \Tile_X6Y7_EE4BEG[8] ,
    \Tile_X6Y7_EE4BEG[7] ,
    \Tile_X6Y7_EE4BEG[6] ,
    \Tile_X6Y7_EE4BEG[5] ,
    \Tile_X6Y7_EE4BEG[4] ,
    \Tile_X6Y7_EE4BEG[3] ,
    \Tile_X6Y7_EE4BEG[2] ,
    \Tile_X6Y7_EE4BEG[1] ,
    \Tile_X6Y7_EE4BEG[0] }),
    .EE4END({\Tile_X5Y7_EE4BEG[15] ,
    \Tile_X5Y7_EE4BEG[14] ,
    \Tile_X5Y7_EE4BEG[13] ,
    \Tile_X5Y7_EE4BEG[12] ,
    \Tile_X5Y7_EE4BEG[11] ,
    \Tile_X5Y7_EE4BEG[10] ,
    \Tile_X5Y7_EE4BEG[9] ,
    \Tile_X5Y7_EE4BEG[8] ,
    \Tile_X5Y7_EE4BEG[7] ,
    \Tile_X5Y7_EE4BEG[6] ,
    \Tile_X5Y7_EE4BEG[5] ,
    \Tile_X5Y7_EE4BEG[4] ,
    \Tile_X5Y7_EE4BEG[3] ,
    \Tile_X5Y7_EE4BEG[2] ,
    \Tile_X5Y7_EE4BEG[1] ,
    \Tile_X5Y7_EE4BEG[0] }),
    .FrameData({\Tile_X5Y7_FrameData_O[31] ,
    \Tile_X5Y7_FrameData_O[30] ,
    \Tile_X5Y7_FrameData_O[29] ,
    \Tile_X5Y7_FrameData_O[28] ,
    \Tile_X5Y7_FrameData_O[27] ,
    \Tile_X5Y7_FrameData_O[26] ,
    \Tile_X5Y7_FrameData_O[25] ,
    \Tile_X5Y7_FrameData_O[24] ,
    \Tile_X5Y7_FrameData_O[23] ,
    \Tile_X5Y7_FrameData_O[22] ,
    \Tile_X5Y7_FrameData_O[21] ,
    \Tile_X5Y7_FrameData_O[20] ,
    \Tile_X5Y7_FrameData_O[19] ,
    \Tile_X5Y7_FrameData_O[18] ,
    \Tile_X5Y7_FrameData_O[17] ,
    \Tile_X5Y7_FrameData_O[16] ,
    \Tile_X5Y7_FrameData_O[15] ,
    \Tile_X5Y7_FrameData_O[14] ,
    \Tile_X5Y7_FrameData_O[13] ,
    \Tile_X5Y7_FrameData_O[12] ,
    \Tile_X5Y7_FrameData_O[11] ,
    \Tile_X5Y7_FrameData_O[10] ,
    \Tile_X5Y7_FrameData_O[9] ,
    \Tile_X5Y7_FrameData_O[8] ,
    \Tile_X5Y7_FrameData_O[7] ,
    \Tile_X5Y7_FrameData_O[6] ,
    \Tile_X5Y7_FrameData_O[5] ,
    \Tile_X5Y7_FrameData_O[4] ,
    \Tile_X5Y7_FrameData_O[3] ,
    \Tile_X5Y7_FrameData_O[2] ,
    \Tile_X5Y7_FrameData_O[1] ,
    \Tile_X5Y7_FrameData_O[0] }),
    .FrameData_O({\Tile_X6Y7_FrameData_O[31] ,
    \Tile_X6Y7_FrameData_O[30] ,
    \Tile_X6Y7_FrameData_O[29] ,
    \Tile_X6Y7_FrameData_O[28] ,
    \Tile_X6Y7_FrameData_O[27] ,
    \Tile_X6Y7_FrameData_O[26] ,
    \Tile_X6Y7_FrameData_O[25] ,
    \Tile_X6Y7_FrameData_O[24] ,
    \Tile_X6Y7_FrameData_O[23] ,
    \Tile_X6Y7_FrameData_O[22] ,
    \Tile_X6Y7_FrameData_O[21] ,
    \Tile_X6Y7_FrameData_O[20] ,
    \Tile_X6Y7_FrameData_O[19] ,
    \Tile_X6Y7_FrameData_O[18] ,
    \Tile_X6Y7_FrameData_O[17] ,
    \Tile_X6Y7_FrameData_O[16] ,
    \Tile_X6Y7_FrameData_O[15] ,
    \Tile_X6Y7_FrameData_O[14] ,
    \Tile_X6Y7_FrameData_O[13] ,
    \Tile_X6Y7_FrameData_O[12] ,
    \Tile_X6Y7_FrameData_O[11] ,
    \Tile_X6Y7_FrameData_O[10] ,
    \Tile_X6Y7_FrameData_O[9] ,
    \Tile_X6Y7_FrameData_O[8] ,
    \Tile_X6Y7_FrameData_O[7] ,
    \Tile_X6Y7_FrameData_O[6] ,
    \Tile_X6Y7_FrameData_O[5] ,
    \Tile_X6Y7_FrameData_O[4] ,
    \Tile_X6Y7_FrameData_O[3] ,
    \Tile_X6Y7_FrameData_O[2] ,
    \Tile_X6Y7_FrameData_O[1] ,
    \Tile_X6Y7_FrameData_O[0] }),
    .FrameStrobe({\Tile_X6Y8_FrameStrobe_O[19] ,
    \Tile_X6Y8_FrameStrobe_O[18] ,
    \Tile_X6Y8_FrameStrobe_O[17] ,
    \Tile_X6Y8_FrameStrobe_O[16] ,
    \Tile_X6Y8_FrameStrobe_O[15] ,
    \Tile_X6Y8_FrameStrobe_O[14] ,
    \Tile_X6Y8_FrameStrobe_O[13] ,
    \Tile_X6Y8_FrameStrobe_O[12] ,
    \Tile_X6Y8_FrameStrobe_O[11] ,
    \Tile_X6Y8_FrameStrobe_O[10] ,
    \Tile_X6Y8_FrameStrobe_O[9] ,
    \Tile_X6Y8_FrameStrobe_O[8] ,
    \Tile_X6Y8_FrameStrobe_O[7] ,
    \Tile_X6Y8_FrameStrobe_O[6] ,
    \Tile_X6Y8_FrameStrobe_O[5] ,
    \Tile_X6Y8_FrameStrobe_O[4] ,
    \Tile_X6Y8_FrameStrobe_O[3] ,
    \Tile_X6Y8_FrameStrobe_O[2] ,
    \Tile_X6Y8_FrameStrobe_O[1] ,
    \Tile_X6Y8_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X6Y7_FrameStrobe_O[19] ,
    \Tile_X6Y7_FrameStrobe_O[18] ,
    \Tile_X6Y7_FrameStrobe_O[17] ,
    \Tile_X6Y7_FrameStrobe_O[16] ,
    \Tile_X6Y7_FrameStrobe_O[15] ,
    \Tile_X6Y7_FrameStrobe_O[14] ,
    \Tile_X6Y7_FrameStrobe_O[13] ,
    \Tile_X6Y7_FrameStrobe_O[12] ,
    \Tile_X6Y7_FrameStrobe_O[11] ,
    \Tile_X6Y7_FrameStrobe_O[10] ,
    \Tile_X6Y7_FrameStrobe_O[9] ,
    \Tile_X6Y7_FrameStrobe_O[8] ,
    \Tile_X6Y7_FrameStrobe_O[7] ,
    \Tile_X6Y7_FrameStrobe_O[6] ,
    \Tile_X6Y7_FrameStrobe_O[5] ,
    \Tile_X6Y7_FrameStrobe_O[4] ,
    \Tile_X6Y7_FrameStrobe_O[3] ,
    \Tile_X6Y7_FrameStrobe_O[2] ,
    \Tile_X6Y7_FrameStrobe_O[1] ,
    \Tile_X6Y7_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X6Y7_N1BEG[3] ,
    \Tile_X6Y7_N1BEG[2] ,
    \Tile_X6Y7_N1BEG[1] ,
    \Tile_X6Y7_N1BEG[0] }),
    .N1END({\Tile_X6Y8_N1BEG[3] ,
    \Tile_X6Y8_N1BEG[2] ,
    \Tile_X6Y8_N1BEG[1] ,
    \Tile_X6Y8_N1BEG[0] }),
    .N2BEG({\Tile_X6Y7_N2BEG[7] ,
    \Tile_X6Y7_N2BEG[6] ,
    \Tile_X6Y7_N2BEG[5] ,
    \Tile_X6Y7_N2BEG[4] ,
    \Tile_X6Y7_N2BEG[3] ,
    \Tile_X6Y7_N2BEG[2] ,
    \Tile_X6Y7_N2BEG[1] ,
    \Tile_X6Y7_N2BEG[0] }),
    .N2BEGb({\Tile_X6Y7_N2BEGb[7] ,
    \Tile_X6Y7_N2BEGb[6] ,
    \Tile_X6Y7_N2BEGb[5] ,
    \Tile_X6Y7_N2BEGb[4] ,
    \Tile_X6Y7_N2BEGb[3] ,
    \Tile_X6Y7_N2BEGb[2] ,
    \Tile_X6Y7_N2BEGb[1] ,
    \Tile_X6Y7_N2BEGb[0] }),
    .N2END({\Tile_X6Y8_N2BEGb[7] ,
    \Tile_X6Y8_N2BEGb[6] ,
    \Tile_X6Y8_N2BEGb[5] ,
    \Tile_X6Y8_N2BEGb[4] ,
    \Tile_X6Y8_N2BEGb[3] ,
    \Tile_X6Y8_N2BEGb[2] ,
    \Tile_X6Y8_N2BEGb[1] ,
    \Tile_X6Y8_N2BEGb[0] }),
    .N2MID({\Tile_X6Y8_N2BEG[7] ,
    \Tile_X6Y8_N2BEG[6] ,
    \Tile_X6Y8_N2BEG[5] ,
    \Tile_X6Y8_N2BEG[4] ,
    \Tile_X6Y8_N2BEG[3] ,
    \Tile_X6Y8_N2BEG[2] ,
    \Tile_X6Y8_N2BEG[1] ,
    \Tile_X6Y8_N2BEG[0] }),
    .N4BEG({\Tile_X6Y7_N4BEG[15] ,
    \Tile_X6Y7_N4BEG[14] ,
    \Tile_X6Y7_N4BEG[13] ,
    \Tile_X6Y7_N4BEG[12] ,
    \Tile_X6Y7_N4BEG[11] ,
    \Tile_X6Y7_N4BEG[10] ,
    \Tile_X6Y7_N4BEG[9] ,
    \Tile_X6Y7_N4BEG[8] ,
    \Tile_X6Y7_N4BEG[7] ,
    \Tile_X6Y7_N4BEG[6] ,
    \Tile_X6Y7_N4BEG[5] ,
    \Tile_X6Y7_N4BEG[4] ,
    \Tile_X6Y7_N4BEG[3] ,
    \Tile_X6Y7_N4BEG[2] ,
    \Tile_X6Y7_N4BEG[1] ,
    \Tile_X6Y7_N4BEG[0] }),
    .N4END({\Tile_X6Y8_N4BEG[15] ,
    \Tile_X6Y8_N4BEG[14] ,
    \Tile_X6Y8_N4BEG[13] ,
    \Tile_X6Y8_N4BEG[12] ,
    \Tile_X6Y8_N4BEG[11] ,
    \Tile_X6Y8_N4BEG[10] ,
    \Tile_X6Y8_N4BEG[9] ,
    \Tile_X6Y8_N4BEG[8] ,
    \Tile_X6Y8_N4BEG[7] ,
    \Tile_X6Y8_N4BEG[6] ,
    \Tile_X6Y8_N4BEG[5] ,
    \Tile_X6Y8_N4BEG[4] ,
    \Tile_X6Y8_N4BEG[3] ,
    \Tile_X6Y8_N4BEG[2] ,
    \Tile_X6Y8_N4BEG[1] ,
    \Tile_X6Y8_N4BEG[0] }),
    .NN4BEG({\Tile_X6Y7_NN4BEG[15] ,
    \Tile_X6Y7_NN4BEG[14] ,
    \Tile_X6Y7_NN4BEG[13] ,
    \Tile_X6Y7_NN4BEG[12] ,
    \Tile_X6Y7_NN4BEG[11] ,
    \Tile_X6Y7_NN4BEG[10] ,
    \Tile_X6Y7_NN4BEG[9] ,
    \Tile_X6Y7_NN4BEG[8] ,
    \Tile_X6Y7_NN4BEG[7] ,
    \Tile_X6Y7_NN4BEG[6] ,
    \Tile_X6Y7_NN4BEG[5] ,
    \Tile_X6Y7_NN4BEG[4] ,
    \Tile_X6Y7_NN4BEG[3] ,
    \Tile_X6Y7_NN4BEG[2] ,
    \Tile_X6Y7_NN4BEG[1] ,
    \Tile_X6Y7_NN4BEG[0] }),
    .NN4END({\Tile_X6Y8_NN4BEG[15] ,
    \Tile_X6Y8_NN4BEG[14] ,
    \Tile_X6Y8_NN4BEG[13] ,
    \Tile_X6Y8_NN4BEG[12] ,
    \Tile_X6Y8_NN4BEG[11] ,
    \Tile_X6Y8_NN4BEG[10] ,
    \Tile_X6Y8_NN4BEG[9] ,
    \Tile_X6Y8_NN4BEG[8] ,
    \Tile_X6Y8_NN4BEG[7] ,
    \Tile_X6Y8_NN4BEG[6] ,
    \Tile_X6Y8_NN4BEG[5] ,
    \Tile_X6Y8_NN4BEG[4] ,
    \Tile_X6Y8_NN4BEG[3] ,
    \Tile_X6Y8_NN4BEG[2] ,
    \Tile_X6Y8_NN4BEG[1] ,
    \Tile_X6Y8_NN4BEG[0] }),
    .S1BEG({\Tile_X6Y7_S1BEG[3] ,
    \Tile_X6Y7_S1BEG[2] ,
    \Tile_X6Y7_S1BEG[1] ,
    \Tile_X6Y7_S1BEG[0] }),
    .S1END({\Tile_X6Y6_S1BEG[3] ,
    \Tile_X6Y6_S1BEG[2] ,
    \Tile_X6Y6_S1BEG[1] ,
    \Tile_X6Y6_S1BEG[0] }),
    .S2BEG({\Tile_X6Y7_S2BEG[7] ,
    \Tile_X6Y7_S2BEG[6] ,
    \Tile_X6Y7_S2BEG[5] ,
    \Tile_X6Y7_S2BEG[4] ,
    \Tile_X6Y7_S2BEG[3] ,
    \Tile_X6Y7_S2BEG[2] ,
    \Tile_X6Y7_S2BEG[1] ,
    \Tile_X6Y7_S2BEG[0] }),
    .S2BEGb({\Tile_X6Y7_S2BEGb[7] ,
    \Tile_X6Y7_S2BEGb[6] ,
    \Tile_X6Y7_S2BEGb[5] ,
    \Tile_X6Y7_S2BEGb[4] ,
    \Tile_X6Y7_S2BEGb[3] ,
    \Tile_X6Y7_S2BEGb[2] ,
    \Tile_X6Y7_S2BEGb[1] ,
    \Tile_X6Y7_S2BEGb[0] }),
    .S2END({\Tile_X6Y6_S2BEGb[7] ,
    \Tile_X6Y6_S2BEGb[6] ,
    \Tile_X6Y6_S2BEGb[5] ,
    \Tile_X6Y6_S2BEGb[4] ,
    \Tile_X6Y6_S2BEGb[3] ,
    \Tile_X6Y6_S2BEGb[2] ,
    \Tile_X6Y6_S2BEGb[1] ,
    \Tile_X6Y6_S2BEGb[0] }),
    .S2MID({\Tile_X6Y6_S2BEG[7] ,
    \Tile_X6Y6_S2BEG[6] ,
    \Tile_X6Y6_S2BEG[5] ,
    \Tile_X6Y6_S2BEG[4] ,
    \Tile_X6Y6_S2BEG[3] ,
    \Tile_X6Y6_S2BEG[2] ,
    \Tile_X6Y6_S2BEG[1] ,
    \Tile_X6Y6_S2BEG[0] }),
    .S4BEG({\Tile_X6Y7_S4BEG[15] ,
    \Tile_X6Y7_S4BEG[14] ,
    \Tile_X6Y7_S4BEG[13] ,
    \Tile_X6Y7_S4BEG[12] ,
    \Tile_X6Y7_S4BEG[11] ,
    \Tile_X6Y7_S4BEG[10] ,
    \Tile_X6Y7_S4BEG[9] ,
    \Tile_X6Y7_S4BEG[8] ,
    \Tile_X6Y7_S4BEG[7] ,
    \Tile_X6Y7_S4BEG[6] ,
    \Tile_X6Y7_S4BEG[5] ,
    \Tile_X6Y7_S4BEG[4] ,
    \Tile_X6Y7_S4BEG[3] ,
    \Tile_X6Y7_S4BEG[2] ,
    \Tile_X6Y7_S4BEG[1] ,
    \Tile_X6Y7_S4BEG[0] }),
    .S4END({\Tile_X6Y6_S4BEG[15] ,
    \Tile_X6Y6_S4BEG[14] ,
    \Tile_X6Y6_S4BEG[13] ,
    \Tile_X6Y6_S4BEG[12] ,
    \Tile_X6Y6_S4BEG[11] ,
    \Tile_X6Y6_S4BEG[10] ,
    \Tile_X6Y6_S4BEG[9] ,
    \Tile_X6Y6_S4BEG[8] ,
    \Tile_X6Y6_S4BEG[7] ,
    \Tile_X6Y6_S4BEG[6] ,
    \Tile_X6Y6_S4BEG[5] ,
    \Tile_X6Y6_S4BEG[4] ,
    \Tile_X6Y6_S4BEG[3] ,
    \Tile_X6Y6_S4BEG[2] ,
    \Tile_X6Y6_S4BEG[1] ,
    \Tile_X6Y6_S4BEG[0] }),
    .SS4BEG({\Tile_X6Y7_SS4BEG[15] ,
    \Tile_X6Y7_SS4BEG[14] ,
    \Tile_X6Y7_SS4BEG[13] ,
    \Tile_X6Y7_SS4BEG[12] ,
    \Tile_X6Y7_SS4BEG[11] ,
    \Tile_X6Y7_SS4BEG[10] ,
    \Tile_X6Y7_SS4BEG[9] ,
    \Tile_X6Y7_SS4BEG[8] ,
    \Tile_X6Y7_SS4BEG[7] ,
    \Tile_X6Y7_SS4BEG[6] ,
    \Tile_X6Y7_SS4BEG[5] ,
    \Tile_X6Y7_SS4BEG[4] ,
    \Tile_X6Y7_SS4BEG[3] ,
    \Tile_X6Y7_SS4BEG[2] ,
    \Tile_X6Y7_SS4BEG[1] ,
    \Tile_X6Y7_SS4BEG[0] }),
    .SS4END({\Tile_X6Y6_SS4BEG[15] ,
    \Tile_X6Y6_SS4BEG[14] ,
    \Tile_X6Y6_SS4BEG[13] ,
    \Tile_X6Y6_SS4BEG[12] ,
    \Tile_X6Y6_SS4BEG[11] ,
    \Tile_X6Y6_SS4BEG[10] ,
    \Tile_X6Y6_SS4BEG[9] ,
    \Tile_X6Y6_SS4BEG[8] ,
    \Tile_X6Y6_SS4BEG[7] ,
    \Tile_X6Y6_SS4BEG[6] ,
    \Tile_X6Y6_SS4BEG[5] ,
    \Tile_X6Y6_SS4BEG[4] ,
    \Tile_X6Y6_SS4BEG[3] ,
    \Tile_X6Y6_SS4BEG[2] ,
    \Tile_X6Y6_SS4BEG[1] ,
    \Tile_X6Y6_SS4BEG[0] }),
    .W1BEG({\Tile_X6Y7_W1BEG[3] ,
    \Tile_X6Y7_W1BEG[2] ,
    \Tile_X6Y7_W1BEG[1] ,
    \Tile_X6Y7_W1BEG[0] }),
    .W1END({\Tile_X7Y7_W1BEG[3] ,
    \Tile_X7Y7_W1BEG[2] ,
    \Tile_X7Y7_W1BEG[1] ,
    \Tile_X7Y7_W1BEG[0] }),
    .W2BEG({\Tile_X6Y7_W2BEG[7] ,
    \Tile_X6Y7_W2BEG[6] ,
    \Tile_X6Y7_W2BEG[5] ,
    \Tile_X6Y7_W2BEG[4] ,
    \Tile_X6Y7_W2BEG[3] ,
    \Tile_X6Y7_W2BEG[2] ,
    \Tile_X6Y7_W2BEG[1] ,
    \Tile_X6Y7_W2BEG[0] }),
    .W2BEGb({\Tile_X6Y7_W2BEGb[7] ,
    \Tile_X6Y7_W2BEGb[6] ,
    \Tile_X6Y7_W2BEGb[5] ,
    \Tile_X6Y7_W2BEGb[4] ,
    \Tile_X6Y7_W2BEGb[3] ,
    \Tile_X6Y7_W2BEGb[2] ,
    \Tile_X6Y7_W2BEGb[1] ,
    \Tile_X6Y7_W2BEGb[0] }),
    .W2END({\Tile_X7Y7_W2BEGb[7] ,
    \Tile_X7Y7_W2BEGb[6] ,
    \Tile_X7Y7_W2BEGb[5] ,
    \Tile_X7Y7_W2BEGb[4] ,
    \Tile_X7Y7_W2BEGb[3] ,
    \Tile_X7Y7_W2BEGb[2] ,
    \Tile_X7Y7_W2BEGb[1] ,
    \Tile_X7Y7_W2BEGb[0] }),
    .W2MID({\Tile_X7Y7_W2BEG[7] ,
    \Tile_X7Y7_W2BEG[6] ,
    \Tile_X7Y7_W2BEG[5] ,
    \Tile_X7Y7_W2BEG[4] ,
    \Tile_X7Y7_W2BEG[3] ,
    \Tile_X7Y7_W2BEG[2] ,
    \Tile_X7Y7_W2BEG[1] ,
    \Tile_X7Y7_W2BEG[0] }),
    .W6BEG({\Tile_X6Y7_W6BEG[11] ,
    \Tile_X6Y7_W6BEG[10] ,
    \Tile_X6Y7_W6BEG[9] ,
    \Tile_X6Y7_W6BEG[8] ,
    \Tile_X6Y7_W6BEG[7] ,
    \Tile_X6Y7_W6BEG[6] ,
    \Tile_X6Y7_W6BEG[5] ,
    \Tile_X6Y7_W6BEG[4] ,
    \Tile_X6Y7_W6BEG[3] ,
    \Tile_X6Y7_W6BEG[2] ,
    \Tile_X6Y7_W6BEG[1] ,
    \Tile_X6Y7_W6BEG[0] }),
    .W6END({\Tile_X7Y7_W6BEG[11] ,
    \Tile_X7Y7_W6BEG[10] ,
    \Tile_X7Y7_W6BEG[9] ,
    \Tile_X7Y7_W6BEG[8] ,
    \Tile_X7Y7_W6BEG[7] ,
    \Tile_X7Y7_W6BEG[6] ,
    \Tile_X7Y7_W6BEG[5] ,
    \Tile_X7Y7_W6BEG[4] ,
    \Tile_X7Y7_W6BEG[3] ,
    \Tile_X7Y7_W6BEG[2] ,
    \Tile_X7Y7_W6BEG[1] ,
    \Tile_X7Y7_W6BEG[0] }),
    .WW4BEG({\Tile_X6Y7_WW4BEG[15] ,
    \Tile_X6Y7_WW4BEG[14] ,
    \Tile_X6Y7_WW4BEG[13] ,
    \Tile_X6Y7_WW4BEG[12] ,
    \Tile_X6Y7_WW4BEG[11] ,
    \Tile_X6Y7_WW4BEG[10] ,
    \Tile_X6Y7_WW4BEG[9] ,
    \Tile_X6Y7_WW4BEG[8] ,
    \Tile_X6Y7_WW4BEG[7] ,
    \Tile_X6Y7_WW4BEG[6] ,
    \Tile_X6Y7_WW4BEG[5] ,
    \Tile_X6Y7_WW4BEG[4] ,
    \Tile_X6Y7_WW4BEG[3] ,
    \Tile_X6Y7_WW4BEG[2] ,
    \Tile_X6Y7_WW4BEG[1] ,
    \Tile_X6Y7_WW4BEG[0] }),
    .WW4END({\Tile_X7Y7_WW4BEG[15] ,
    \Tile_X7Y7_WW4BEG[14] ,
    \Tile_X7Y7_WW4BEG[13] ,
    \Tile_X7Y7_WW4BEG[12] ,
    \Tile_X7Y7_WW4BEG[11] ,
    \Tile_X7Y7_WW4BEG[10] ,
    \Tile_X7Y7_WW4BEG[9] ,
    \Tile_X7Y7_WW4BEG[8] ,
    \Tile_X7Y7_WW4BEG[7] ,
    \Tile_X7Y7_WW4BEG[6] ,
    \Tile_X7Y7_WW4BEG[5] ,
    \Tile_X7Y7_WW4BEG[4] ,
    \Tile_X7Y7_WW4BEG[3] ,
    \Tile_X7Y7_WW4BEG[2] ,
    \Tile_X7Y7_WW4BEG[1] ,
    \Tile_X7Y7_WW4BEG[0] }));
 LUT4AB Tile_X6Y8_LUT4AB (.Ci(Tile_X6Y9_Co),
    .Co(Tile_X6Y8_Co),
    .UserCLK(Tile_X6Y9_UserCLKo),
    .UserCLKo(Tile_X6Y8_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X6Y8_E1BEG[3] ,
    \Tile_X6Y8_E1BEG[2] ,
    \Tile_X6Y8_E1BEG[1] ,
    \Tile_X6Y8_E1BEG[0] }),
    .E1END({\Tile_X5Y8_E1BEG[3] ,
    \Tile_X5Y8_E1BEG[2] ,
    \Tile_X5Y8_E1BEG[1] ,
    \Tile_X5Y8_E1BEG[0] }),
    .E2BEG({\Tile_X6Y8_E2BEG[7] ,
    \Tile_X6Y8_E2BEG[6] ,
    \Tile_X6Y8_E2BEG[5] ,
    \Tile_X6Y8_E2BEG[4] ,
    \Tile_X6Y8_E2BEG[3] ,
    \Tile_X6Y8_E2BEG[2] ,
    \Tile_X6Y8_E2BEG[1] ,
    \Tile_X6Y8_E2BEG[0] }),
    .E2BEGb({\Tile_X6Y8_E2BEGb[7] ,
    \Tile_X6Y8_E2BEGb[6] ,
    \Tile_X6Y8_E2BEGb[5] ,
    \Tile_X6Y8_E2BEGb[4] ,
    \Tile_X6Y8_E2BEGb[3] ,
    \Tile_X6Y8_E2BEGb[2] ,
    \Tile_X6Y8_E2BEGb[1] ,
    \Tile_X6Y8_E2BEGb[0] }),
    .E2END({\Tile_X5Y8_E2BEGb[7] ,
    \Tile_X5Y8_E2BEGb[6] ,
    \Tile_X5Y8_E2BEGb[5] ,
    \Tile_X5Y8_E2BEGb[4] ,
    \Tile_X5Y8_E2BEGb[3] ,
    \Tile_X5Y8_E2BEGb[2] ,
    \Tile_X5Y8_E2BEGb[1] ,
    \Tile_X5Y8_E2BEGb[0] }),
    .E2MID({\Tile_X5Y8_E2BEG[7] ,
    \Tile_X5Y8_E2BEG[6] ,
    \Tile_X5Y8_E2BEG[5] ,
    \Tile_X5Y8_E2BEG[4] ,
    \Tile_X5Y8_E2BEG[3] ,
    \Tile_X5Y8_E2BEG[2] ,
    \Tile_X5Y8_E2BEG[1] ,
    \Tile_X5Y8_E2BEG[0] }),
    .E6BEG({\Tile_X6Y8_E6BEG[11] ,
    \Tile_X6Y8_E6BEG[10] ,
    \Tile_X6Y8_E6BEG[9] ,
    \Tile_X6Y8_E6BEG[8] ,
    \Tile_X6Y8_E6BEG[7] ,
    \Tile_X6Y8_E6BEG[6] ,
    \Tile_X6Y8_E6BEG[5] ,
    \Tile_X6Y8_E6BEG[4] ,
    \Tile_X6Y8_E6BEG[3] ,
    \Tile_X6Y8_E6BEG[2] ,
    \Tile_X6Y8_E6BEG[1] ,
    \Tile_X6Y8_E6BEG[0] }),
    .E6END({\Tile_X5Y8_E6BEG[11] ,
    \Tile_X5Y8_E6BEG[10] ,
    \Tile_X5Y8_E6BEG[9] ,
    \Tile_X5Y8_E6BEG[8] ,
    \Tile_X5Y8_E6BEG[7] ,
    \Tile_X5Y8_E6BEG[6] ,
    \Tile_X5Y8_E6BEG[5] ,
    \Tile_X5Y8_E6BEG[4] ,
    \Tile_X5Y8_E6BEG[3] ,
    \Tile_X5Y8_E6BEG[2] ,
    \Tile_X5Y8_E6BEG[1] ,
    \Tile_X5Y8_E6BEG[0] }),
    .EE4BEG({\Tile_X6Y8_EE4BEG[15] ,
    \Tile_X6Y8_EE4BEG[14] ,
    \Tile_X6Y8_EE4BEG[13] ,
    \Tile_X6Y8_EE4BEG[12] ,
    \Tile_X6Y8_EE4BEG[11] ,
    \Tile_X6Y8_EE4BEG[10] ,
    \Tile_X6Y8_EE4BEG[9] ,
    \Tile_X6Y8_EE4BEG[8] ,
    \Tile_X6Y8_EE4BEG[7] ,
    \Tile_X6Y8_EE4BEG[6] ,
    \Tile_X6Y8_EE4BEG[5] ,
    \Tile_X6Y8_EE4BEG[4] ,
    \Tile_X6Y8_EE4BEG[3] ,
    \Tile_X6Y8_EE4BEG[2] ,
    \Tile_X6Y8_EE4BEG[1] ,
    \Tile_X6Y8_EE4BEG[0] }),
    .EE4END({\Tile_X5Y8_EE4BEG[15] ,
    \Tile_X5Y8_EE4BEG[14] ,
    \Tile_X5Y8_EE4BEG[13] ,
    \Tile_X5Y8_EE4BEG[12] ,
    \Tile_X5Y8_EE4BEG[11] ,
    \Tile_X5Y8_EE4BEG[10] ,
    \Tile_X5Y8_EE4BEG[9] ,
    \Tile_X5Y8_EE4BEG[8] ,
    \Tile_X5Y8_EE4BEG[7] ,
    \Tile_X5Y8_EE4BEG[6] ,
    \Tile_X5Y8_EE4BEG[5] ,
    \Tile_X5Y8_EE4BEG[4] ,
    \Tile_X5Y8_EE4BEG[3] ,
    \Tile_X5Y8_EE4BEG[2] ,
    \Tile_X5Y8_EE4BEG[1] ,
    \Tile_X5Y8_EE4BEG[0] }),
    .FrameData({\Tile_X5Y8_FrameData_O[31] ,
    \Tile_X5Y8_FrameData_O[30] ,
    \Tile_X5Y8_FrameData_O[29] ,
    \Tile_X5Y8_FrameData_O[28] ,
    \Tile_X5Y8_FrameData_O[27] ,
    \Tile_X5Y8_FrameData_O[26] ,
    \Tile_X5Y8_FrameData_O[25] ,
    \Tile_X5Y8_FrameData_O[24] ,
    \Tile_X5Y8_FrameData_O[23] ,
    \Tile_X5Y8_FrameData_O[22] ,
    \Tile_X5Y8_FrameData_O[21] ,
    \Tile_X5Y8_FrameData_O[20] ,
    \Tile_X5Y8_FrameData_O[19] ,
    \Tile_X5Y8_FrameData_O[18] ,
    \Tile_X5Y8_FrameData_O[17] ,
    \Tile_X5Y8_FrameData_O[16] ,
    \Tile_X5Y8_FrameData_O[15] ,
    \Tile_X5Y8_FrameData_O[14] ,
    \Tile_X5Y8_FrameData_O[13] ,
    \Tile_X5Y8_FrameData_O[12] ,
    \Tile_X5Y8_FrameData_O[11] ,
    \Tile_X5Y8_FrameData_O[10] ,
    \Tile_X5Y8_FrameData_O[9] ,
    \Tile_X5Y8_FrameData_O[8] ,
    \Tile_X5Y8_FrameData_O[7] ,
    \Tile_X5Y8_FrameData_O[6] ,
    \Tile_X5Y8_FrameData_O[5] ,
    \Tile_X5Y8_FrameData_O[4] ,
    \Tile_X5Y8_FrameData_O[3] ,
    \Tile_X5Y8_FrameData_O[2] ,
    \Tile_X5Y8_FrameData_O[1] ,
    \Tile_X5Y8_FrameData_O[0] }),
    .FrameData_O({\Tile_X6Y8_FrameData_O[31] ,
    \Tile_X6Y8_FrameData_O[30] ,
    \Tile_X6Y8_FrameData_O[29] ,
    \Tile_X6Y8_FrameData_O[28] ,
    \Tile_X6Y8_FrameData_O[27] ,
    \Tile_X6Y8_FrameData_O[26] ,
    \Tile_X6Y8_FrameData_O[25] ,
    \Tile_X6Y8_FrameData_O[24] ,
    \Tile_X6Y8_FrameData_O[23] ,
    \Tile_X6Y8_FrameData_O[22] ,
    \Tile_X6Y8_FrameData_O[21] ,
    \Tile_X6Y8_FrameData_O[20] ,
    \Tile_X6Y8_FrameData_O[19] ,
    \Tile_X6Y8_FrameData_O[18] ,
    \Tile_X6Y8_FrameData_O[17] ,
    \Tile_X6Y8_FrameData_O[16] ,
    \Tile_X6Y8_FrameData_O[15] ,
    \Tile_X6Y8_FrameData_O[14] ,
    \Tile_X6Y8_FrameData_O[13] ,
    \Tile_X6Y8_FrameData_O[12] ,
    \Tile_X6Y8_FrameData_O[11] ,
    \Tile_X6Y8_FrameData_O[10] ,
    \Tile_X6Y8_FrameData_O[9] ,
    \Tile_X6Y8_FrameData_O[8] ,
    \Tile_X6Y8_FrameData_O[7] ,
    \Tile_X6Y8_FrameData_O[6] ,
    \Tile_X6Y8_FrameData_O[5] ,
    \Tile_X6Y8_FrameData_O[4] ,
    \Tile_X6Y8_FrameData_O[3] ,
    \Tile_X6Y8_FrameData_O[2] ,
    \Tile_X6Y8_FrameData_O[1] ,
    \Tile_X6Y8_FrameData_O[0] }),
    .FrameStrobe({\Tile_X6Y9_FrameStrobe_O[19] ,
    \Tile_X6Y9_FrameStrobe_O[18] ,
    \Tile_X6Y9_FrameStrobe_O[17] ,
    \Tile_X6Y9_FrameStrobe_O[16] ,
    \Tile_X6Y9_FrameStrobe_O[15] ,
    \Tile_X6Y9_FrameStrobe_O[14] ,
    \Tile_X6Y9_FrameStrobe_O[13] ,
    \Tile_X6Y9_FrameStrobe_O[12] ,
    \Tile_X6Y9_FrameStrobe_O[11] ,
    \Tile_X6Y9_FrameStrobe_O[10] ,
    \Tile_X6Y9_FrameStrobe_O[9] ,
    \Tile_X6Y9_FrameStrobe_O[8] ,
    \Tile_X6Y9_FrameStrobe_O[7] ,
    \Tile_X6Y9_FrameStrobe_O[6] ,
    \Tile_X6Y9_FrameStrobe_O[5] ,
    \Tile_X6Y9_FrameStrobe_O[4] ,
    \Tile_X6Y9_FrameStrobe_O[3] ,
    \Tile_X6Y9_FrameStrobe_O[2] ,
    \Tile_X6Y9_FrameStrobe_O[1] ,
    \Tile_X6Y9_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X6Y8_FrameStrobe_O[19] ,
    \Tile_X6Y8_FrameStrobe_O[18] ,
    \Tile_X6Y8_FrameStrobe_O[17] ,
    \Tile_X6Y8_FrameStrobe_O[16] ,
    \Tile_X6Y8_FrameStrobe_O[15] ,
    \Tile_X6Y8_FrameStrobe_O[14] ,
    \Tile_X6Y8_FrameStrobe_O[13] ,
    \Tile_X6Y8_FrameStrobe_O[12] ,
    \Tile_X6Y8_FrameStrobe_O[11] ,
    \Tile_X6Y8_FrameStrobe_O[10] ,
    \Tile_X6Y8_FrameStrobe_O[9] ,
    \Tile_X6Y8_FrameStrobe_O[8] ,
    \Tile_X6Y8_FrameStrobe_O[7] ,
    \Tile_X6Y8_FrameStrobe_O[6] ,
    \Tile_X6Y8_FrameStrobe_O[5] ,
    \Tile_X6Y8_FrameStrobe_O[4] ,
    \Tile_X6Y8_FrameStrobe_O[3] ,
    \Tile_X6Y8_FrameStrobe_O[2] ,
    \Tile_X6Y8_FrameStrobe_O[1] ,
    \Tile_X6Y8_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X6Y8_N1BEG[3] ,
    \Tile_X6Y8_N1BEG[2] ,
    \Tile_X6Y8_N1BEG[1] ,
    \Tile_X6Y8_N1BEG[0] }),
    .N1END({\Tile_X6Y9_N1BEG[3] ,
    \Tile_X6Y9_N1BEG[2] ,
    \Tile_X6Y9_N1BEG[1] ,
    \Tile_X6Y9_N1BEG[0] }),
    .N2BEG({\Tile_X6Y8_N2BEG[7] ,
    \Tile_X6Y8_N2BEG[6] ,
    \Tile_X6Y8_N2BEG[5] ,
    \Tile_X6Y8_N2BEG[4] ,
    \Tile_X6Y8_N2BEG[3] ,
    \Tile_X6Y8_N2BEG[2] ,
    \Tile_X6Y8_N2BEG[1] ,
    \Tile_X6Y8_N2BEG[0] }),
    .N2BEGb({\Tile_X6Y8_N2BEGb[7] ,
    \Tile_X6Y8_N2BEGb[6] ,
    \Tile_X6Y8_N2BEGb[5] ,
    \Tile_X6Y8_N2BEGb[4] ,
    \Tile_X6Y8_N2BEGb[3] ,
    \Tile_X6Y8_N2BEGb[2] ,
    \Tile_X6Y8_N2BEGb[1] ,
    \Tile_X6Y8_N2BEGb[0] }),
    .N2END({\Tile_X6Y9_N2BEGb[7] ,
    \Tile_X6Y9_N2BEGb[6] ,
    \Tile_X6Y9_N2BEGb[5] ,
    \Tile_X6Y9_N2BEGb[4] ,
    \Tile_X6Y9_N2BEGb[3] ,
    \Tile_X6Y9_N2BEGb[2] ,
    \Tile_X6Y9_N2BEGb[1] ,
    \Tile_X6Y9_N2BEGb[0] }),
    .N2MID({\Tile_X6Y9_N2BEG[7] ,
    \Tile_X6Y9_N2BEG[6] ,
    \Tile_X6Y9_N2BEG[5] ,
    \Tile_X6Y9_N2BEG[4] ,
    \Tile_X6Y9_N2BEG[3] ,
    \Tile_X6Y9_N2BEG[2] ,
    \Tile_X6Y9_N2BEG[1] ,
    \Tile_X6Y9_N2BEG[0] }),
    .N4BEG({\Tile_X6Y8_N4BEG[15] ,
    \Tile_X6Y8_N4BEG[14] ,
    \Tile_X6Y8_N4BEG[13] ,
    \Tile_X6Y8_N4BEG[12] ,
    \Tile_X6Y8_N4BEG[11] ,
    \Tile_X6Y8_N4BEG[10] ,
    \Tile_X6Y8_N4BEG[9] ,
    \Tile_X6Y8_N4BEG[8] ,
    \Tile_X6Y8_N4BEG[7] ,
    \Tile_X6Y8_N4BEG[6] ,
    \Tile_X6Y8_N4BEG[5] ,
    \Tile_X6Y8_N4BEG[4] ,
    \Tile_X6Y8_N4BEG[3] ,
    \Tile_X6Y8_N4BEG[2] ,
    \Tile_X6Y8_N4BEG[1] ,
    \Tile_X6Y8_N4BEG[0] }),
    .N4END({\Tile_X6Y9_N4BEG[15] ,
    \Tile_X6Y9_N4BEG[14] ,
    \Tile_X6Y9_N4BEG[13] ,
    \Tile_X6Y9_N4BEG[12] ,
    \Tile_X6Y9_N4BEG[11] ,
    \Tile_X6Y9_N4BEG[10] ,
    \Tile_X6Y9_N4BEG[9] ,
    \Tile_X6Y9_N4BEG[8] ,
    \Tile_X6Y9_N4BEG[7] ,
    \Tile_X6Y9_N4BEG[6] ,
    \Tile_X6Y9_N4BEG[5] ,
    \Tile_X6Y9_N4BEG[4] ,
    \Tile_X6Y9_N4BEG[3] ,
    \Tile_X6Y9_N4BEG[2] ,
    \Tile_X6Y9_N4BEG[1] ,
    \Tile_X6Y9_N4BEG[0] }),
    .NN4BEG({\Tile_X6Y8_NN4BEG[15] ,
    \Tile_X6Y8_NN4BEG[14] ,
    \Tile_X6Y8_NN4BEG[13] ,
    \Tile_X6Y8_NN4BEG[12] ,
    \Tile_X6Y8_NN4BEG[11] ,
    \Tile_X6Y8_NN4BEG[10] ,
    \Tile_X6Y8_NN4BEG[9] ,
    \Tile_X6Y8_NN4BEG[8] ,
    \Tile_X6Y8_NN4BEG[7] ,
    \Tile_X6Y8_NN4BEG[6] ,
    \Tile_X6Y8_NN4BEG[5] ,
    \Tile_X6Y8_NN4BEG[4] ,
    \Tile_X6Y8_NN4BEG[3] ,
    \Tile_X6Y8_NN4BEG[2] ,
    \Tile_X6Y8_NN4BEG[1] ,
    \Tile_X6Y8_NN4BEG[0] }),
    .NN4END({\Tile_X6Y9_NN4BEG[15] ,
    \Tile_X6Y9_NN4BEG[14] ,
    \Tile_X6Y9_NN4BEG[13] ,
    \Tile_X6Y9_NN4BEG[12] ,
    \Tile_X6Y9_NN4BEG[11] ,
    \Tile_X6Y9_NN4BEG[10] ,
    \Tile_X6Y9_NN4BEG[9] ,
    \Tile_X6Y9_NN4BEG[8] ,
    \Tile_X6Y9_NN4BEG[7] ,
    \Tile_X6Y9_NN4BEG[6] ,
    \Tile_X6Y9_NN4BEG[5] ,
    \Tile_X6Y9_NN4BEG[4] ,
    \Tile_X6Y9_NN4BEG[3] ,
    \Tile_X6Y9_NN4BEG[2] ,
    \Tile_X6Y9_NN4BEG[1] ,
    \Tile_X6Y9_NN4BEG[0] }),
    .S1BEG({\Tile_X6Y8_S1BEG[3] ,
    \Tile_X6Y8_S1BEG[2] ,
    \Tile_X6Y8_S1BEG[1] ,
    \Tile_X6Y8_S1BEG[0] }),
    .S1END({\Tile_X6Y7_S1BEG[3] ,
    \Tile_X6Y7_S1BEG[2] ,
    \Tile_X6Y7_S1BEG[1] ,
    \Tile_X6Y7_S1BEG[0] }),
    .S2BEG({\Tile_X6Y8_S2BEG[7] ,
    \Tile_X6Y8_S2BEG[6] ,
    \Tile_X6Y8_S2BEG[5] ,
    \Tile_X6Y8_S2BEG[4] ,
    \Tile_X6Y8_S2BEG[3] ,
    \Tile_X6Y8_S2BEG[2] ,
    \Tile_X6Y8_S2BEG[1] ,
    \Tile_X6Y8_S2BEG[0] }),
    .S2BEGb({\Tile_X6Y8_S2BEGb[7] ,
    \Tile_X6Y8_S2BEGb[6] ,
    \Tile_X6Y8_S2BEGb[5] ,
    \Tile_X6Y8_S2BEGb[4] ,
    \Tile_X6Y8_S2BEGb[3] ,
    \Tile_X6Y8_S2BEGb[2] ,
    \Tile_X6Y8_S2BEGb[1] ,
    \Tile_X6Y8_S2BEGb[0] }),
    .S2END({\Tile_X6Y7_S2BEGb[7] ,
    \Tile_X6Y7_S2BEGb[6] ,
    \Tile_X6Y7_S2BEGb[5] ,
    \Tile_X6Y7_S2BEGb[4] ,
    \Tile_X6Y7_S2BEGb[3] ,
    \Tile_X6Y7_S2BEGb[2] ,
    \Tile_X6Y7_S2BEGb[1] ,
    \Tile_X6Y7_S2BEGb[0] }),
    .S2MID({\Tile_X6Y7_S2BEG[7] ,
    \Tile_X6Y7_S2BEG[6] ,
    \Tile_X6Y7_S2BEG[5] ,
    \Tile_X6Y7_S2BEG[4] ,
    \Tile_X6Y7_S2BEG[3] ,
    \Tile_X6Y7_S2BEG[2] ,
    \Tile_X6Y7_S2BEG[1] ,
    \Tile_X6Y7_S2BEG[0] }),
    .S4BEG({\Tile_X6Y8_S4BEG[15] ,
    \Tile_X6Y8_S4BEG[14] ,
    \Tile_X6Y8_S4BEG[13] ,
    \Tile_X6Y8_S4BEG[12] ,
    \Tile_X6Y8_S4BEG[11] ,
    \Tile_X6Y8_S4BEG[10] ,
    \Tile_X6Y8_S4BEG[9] ,
    \Tile_X6Y8_S4BEG[8] ,
    \Tile_X6Y8_S4BEG[7] ,
    \Tile_X6Y8_S4BEG[6] ,
    \Tile_X6Y8_S4BEG[5] ,
    \Tile_X6Y8_S4BEG[4] ,
    \Tile_X6Y8_S4BEG[3] ,
    \Tile_X6Y8_S4BEG[2] ,
    \Tile_X6Y8_S4BEG[1] ,
    \Tile_X6Y8_S4BEG[0] }),
    .S4END({\Tile_X6Y7_S4BEG[15] ,
    \Tile_X6Y7_S4BEG[14] ,
    \Tile_X6Y7_S4BEG[13] ,
    \Tile_X6Y7_S4BEG[12] ,
    \Tile_X6Y7_S4BEG[11] ,
    \Tile_X6Y7_S4BEG[10] ,
    \Tile_X6Y7_S4BEG[9] ,
    \Tile_X6Y7_S4BEG[8] ,
    \Tile_X6Y7_S4BEG[7] ,
    \Tile_X6Y7_S4BEG[6] ,
    \Tile_X6Y7_S4BEG[5] ,
    \Tile_X6Y7_S4BEG[4] ,
    \Tile_X6Y7_S4BEG[3] ,
    \Tile_X6Y7_S4BEG[2] ,
    \Tile_X6Y7_S4BEG[1] ,
    \Tile_X6Y7_S4BEG[0] }),
    .SS4BEG({\Tile_X6Y8_SS4BEG[15] ,
    \Tile_X6Y8_SS4BEG[14] ,
    \Tile_X6Y8_SS4BEG[13] ,
    \Tile_X6Y8_SS4BEG[12] ,
    \Tile_X6Y8_SS4BEG[11] ,
    \Tile_X6Y8_SS4BEG[10] ,
    \Tile_X6Y8_SS4BEG[9] ,
    \Tile_X6Y8_SS4BEG[8] ,
    \Tile_X6Y8_SS4BEG[7] ,
    \Tile_X6Y8_SS4BEG[6] ,
    \Tile_X6Y8_SS4BEG[5] ,
    \Tile_X6Y8_SS4BEG[4] ,
    \Tile_X6Y8_SS4BEG[3] ,
    \Tile_X6Y8_SS4BEG[2] ,
    \Tile_X6Y8_SS4BEG[1] ,
    \Tile_X6Y8_SS4BEG[0] }),
    .SS4END({\Tile_X6Y7_SS4BEG[15] ,
    \Tile_X6Y7_SS4BEG[14] ,
    \Tile_X6Y7_SS4BEG[13] ,
    \Tile_X6Y7_SS4BEG[12] ,
    \Tile_X6Y7_SS4BEG[11] ,
    \Tile_X6Y7_SS4BEG[10] ,
    \Tile_X6Y7_SS4BEG[9] ,
    \Tile_X6Y7_SS4BEG[8] ,
    \Tile_X6Y7_SS4BEG[7] ,
    \Tile_X6Y7_SS4BEG[6] ,
    \Tile_X6Y7_SS4BEG[5] ,
    \Tile_X6Y7_SS4BEG[4] ,
    \Tile_X6Y7_SS4BEG[3] ,
    \Tile_X6Y7_SS4BEG[2] ,
    \Tile_X6Y7_SS4BEG[1] ,
    \Tile_X6Y7_SS4BEG[0] }),
    .W1BEG({\Tile_X6Y8_W1BEG[3] ,
    \Tile_X6Y8_W1BEG[2] ,
    \Tile_X6Y8_W1BEG[1] ,
    \Tile_X6Y8_W1BEG[0] }),
    .W1END({\Tile_X7Y8_W1BEG[3] ,
    \Tile_X7Y8_W1BEG[2] ,
    \Tile_X7Y8_W1BEG[1] ,
    \Tile_X7Y8_W1BEG[0] }),
    .W2BEG({\Tile_X6Y8_W2BEG[7] ,
    \Tile_X6Y8_W2BEG[6] ,
    \Tile_X6Y8_W2BEG[5] ,
    \Tile_X6Y8_W2BEG[4] ,
    \Tile_X6Y8_W2BEG[3] ,
    \Tile_X6Y8_W2BEG[2] ,
    \Tile_X6Y8_W2BEG[1] ,
    \Tile_X6Y8_W2BEG[0] }),
    .W2BEGb({\Tile_X6Y8_W2BEGb[7] ,
    \Tile_X6Y8_W2BEGb[6] ,
    \Tile_X6Y8_W2BEGb[5] ,
    \Tile_X6Y8_W2BEGb[4] ,
    \Tile_X6Y8_W2BEGb[3] ,
    \Tile_X6Y8_W2BEGb[2] ,
    \Tile_X6Y8_W2BEGb[1] ,
    \Tile_X6Y8_W2BEGb[0] }),
    .W2END({\Tile_X7Y8_W2BEGb[7] ,
    \Tile_X7Y8_W2BEGb[6] ,
    \Tile_X7Y8_W2BEGb[5] ,
    \Tile_X7Y8_W2BEGb[4] ,
    \Tile_X7Y8_W2BEGb[3] ,
    \Tile_X7Y8_W2BEGb[2] ,
    \Tile_X7Y8_W2BEGb[1] ,
    \Tile_X7Y8_W2BEGb[0] }),
    .W2MID({\Tile_X7Y8_W2BEG[7] ,
    \Tile_X7Y8_W2BEG[6] ,
    \Tile_X7Y8_W2BEG[5] ,
    \Tile_X7Y8_W2BEG[4] ,
    \Tile_X7Y8_W2BEG[3] ,
    \Tile_X7Y8_W2BEG[2] ,
    \Tile_X7Y8_W2BEG[1] ,
    \Tile_X7Y8_W2BEG[0] }),
    .W6BEG({\Tile_X6Y8_W6BEG[11] ,
    \Tile_X6Y8_W6BEG[10] ,
    \Tile_X6Y8_W6BEG[9] ,
    \Tile_X6Y8_W6BEG[8] ,
    \Tile_X6Y8_W6BEG[7] ,
    \Tile_X6Y8_W6BEG[6] ,
    \Tile_X6Y8_W6BEG[5] ,
    \Tile_X6Y8_W6BEG[4] ,
    \Tile_X6Y8_W6BEG[3] ,
    \Tile_X6Y8_W6BEG[2] ,
    \Tile_X6Y8_W6BEG[1] ,
    \Tile_X6Y8_W6BEG[0] }),
    .W6END({\Tile_X7Y8_W6BEG[11] ,
    \Tile_X7Y8_W6BEG[10] ,
    \Tile_X7Y8_W6BEG[9] ,
    \Tile_X7Y8_W6BEG[8] ,
    \Tile_X7Y8_W6BEG[7] ,
    \Tile_X7Y8_W6BEG[6] ,
    \Tile_X7Y8_W6BEG[5] ,
    \Tile_X7Y8_W6BEG[4] ,
    \Tile_X7Y8_W6BEG[3] ,
    \Tile_X7Y8_W6BEG[2] ,
    \Tile_X7Y8_W6BEG[1] ,
    \Tile_X7Y8_W6BEG[0] }),
    .WW4BEG({\Tile_X6Y8_WW4BEG[15] ,
    \Tile_X6Y8_WW4BEG[14] ,
    \Tile_X6Y8_WW4BEG[13] ,
    \Tile_X6Y8_WW4BEG[12] ,
    \Tile_X6Y8_WW4BEG[11] ,
    \Tile_X6Y8_WW4BEG[10] ,
    \Tile_X6Y8_WW4BEG[9] ,
    \Tile_X6Y8_WW4BEG[8] ,
    \Tile_X6Y8_WW4BEG[7] ,
    \Tile_X6Y8_WW4BEG[6] ,
    \Tile_X6Y8_WW4BEG[5] ,
    \Tile_X6Y8_WW4BEG[4] ,
    \Tile_X6Y8_WW4BEG[3] ,
    \Tile_X6Y8_WW4BEG[2] ,
    \Tile_X6Y8_WW4BEG[1] ,
    \Tile_X6Y8_WW4BEG[0] }),
    .WW4END({\Tile_X7Y8_WW4BEG[15] ,
    \Tile_X7Y8_WW4BEG[14] ,
    \Tile_X7Y8_WW4BEG[13] ,
    \Tile_X7Y8_WW4BEG[12] ,
    \Tile_X7Y8_WW4BEG[11] ,
    \Tile_X7Y8_WW4BEG[10] ,
    \Tile_X7Y8_WW4BEG[9] ,
    \Tile_X7Y8_WW4BEG[8] ,
    \Tile_X7Y8_WW4BEG[7] ,
    \Tile_X7Y8_WW4BEG[6] ,
    \Tile_X7Y8_WW4BEG[5] ,
    \Tile_X7Y8_WW4BEG[4] ,
    \Tile_X7Y8_WW4BEG[3] ,
    \Tile_X7Y8_WW4BEG[2] ,
    \Tile_X7Y8_WW4BEG[1] ,
    \Tile_X7Y8_WW4BEG[0] }));
 LUT4AB Tile_X6Y9_LUT4AB (.Ci(Tile_X6Y10_Co),
    .Co(Tile_X6Y9_Co),
    .UserCLK(Tile_X6Y10_UserCLKo),
    .UserCLKo(Tile_X6Y9_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X6Y9_E1BEG[3] ,
    \Tile_X6Y9_E1BEG[2] ,
    \Tile_X6Y9_E1BEG[1] ,
    \Tile_X6Y9_E1BEG[0] }),
    .E1END({\Tile_X5Y9_E1BEG[3] ,
    \Tile_X5Y9_E1BEG[2] ,
    \Tile_X5Y9_E1BEG[1] ,
    \Tile_X5Y9_E1BEG[0] }),
    .E2BEG({\Tile_X6Y9_E2BEG[7] ,
    \Tile_X6Y9_E2BEG[6] ,
    \Tile_X6Y9_E2BEG[5] ,
    \Tile_X6Y9_E2BEG[4] ,
    \Tile_X6Y9_E2BEG[3] ,
    \Tile_X6Y9_E2BEG[2] ,
    \Tile_X6Y9_E2BEG[1] ,
    \Tile_X6Y9_E2BEG[0] }),
    .E2BEGb({\Tile_X6Y9_E2BEGb[7] ,
    \Tile_X6Y9_E2BEGb[6] ,
    \Tile_X6Y9_E2BEGb[5] ,
    \Tile_X6Y9_E2BEGb[4] ,
    \Tile_X6Y9_E2BEGb[3] ,
    \Tile_X6Y9_E2BEGb[2] ,
    \Tile_X6Y9_E2BEGb[1] ,
    \Tile_X6Y9_E2BEGb[0] }),
    .E2END({\Tile_X5Y9_E2BEGb[7] ,
    \Tile_X5Y9_E2BEGb[6] ,
    \Tile_X5Y9_E2BEGb[5] ,
    \Tile_X5Y9_E2BEGb[4] ,
    \Tile_X5Y9_E2BEGb[3] ,
    \Tile_X5Y9_E2BEGb[2] ,
    \Tile_X5Y9_E2BEGb[1] ,
    \Tile_X5Y9_E2BEGb[0] }),
    .E2MID({\Tile_X5Y9_E2BEG[7] ,
    \Tile_X5Y9_E2BEG[6] ,
    \Tile_X5Y9_E2BEG[5] ,
    \Tile_X5Y9_E2BEG[4] ,
    \Tile_X5Y9_E2BEG[3] ,
    \Tile_X5Y9_E2BEG[2] ,
    \Tile_X5Y9_E2BEG[1] ,
    \Tile_X5Y9_E2BEG[0] }),
    .E6BEG({\Tile_X6Y9_E6BEG[11] ,
    \Tile_X6Y9_E6BEG[10] ,
    \Tile_X6Y9_E6BEG[9] ,
    \Tile_X6Y9_E6BEG[8] ,
    \Tile_X6Y9_E6BEG[7] ,
    \Tile_X6Y9_E6BEG[6] ,
    \Tile_X6Y9_E6BEG[5] ,
    \Tile_X6Y9_E6BEG[4] ,
    \Tile_X6Y9_E6BEG[3] ,
    \Tile_X6Y9_E6BEG[2] ,
    \Tile_X6Y9_E6BEG[1] ,
    \Tile_X6Y9_E6BEG[0] }),
    .E6END({\Tile_X5Y9_E6BEG[11] ,
    \Tile_X5Y9_E6BEG[10] ,
    \Tile_X5Y9_E6BEG[9] ,
    \Tile_X5Y9_E6BEG[8] ,
    \Tile_X5Y9_E6BEG[7] ,
    \Tile_X5Y9_E6BEG[6] ,
    \Tile_X5Y9_E6BEG[5] ,
    \Tile_X5Y9_E6BEG[4] ,
    \Tile_X5Y9_E6BEG[3] ,
    \Tile_X5Y9_E6BEG[2] ,
    \Tile_X5Y9_E6BEG[1] ,
    \Tile_X5Y9_E6BEG[0] }),
    .EE4BEG({\Tile_X6Y9_EE4BEG[15] ,
    \Tile_X6Y9_EE4BEG[14] ,
    \Tile_X6Y9_EE4BEG[13] ,
    \Tile_X6Y9_EE4BEG[12] ,
    \Tile_X6Y9_EE4BEG[11] ,
    \Tile_X6Y9_EE4BEG[10] ,
    \Tile_X6Y9_EE4BEG[9] ,
    \Tile_X6Y9_EE4BEG[8] ,
    \Tile_X6Y9_EE4BEG[7] ,
    \Tile_X6Y9_EE4BEG[6] ,
    \Tile_X6Y9_EE4BEG[5] ,
    \Tile_X6Y9_EE4BEG[4] ,
    \Tile_X6Y9_EE4BEG[3] ,
    \Tile_X6Y9_EE4BEG[2] ,
    \Tile_X6Y9_EE4BEG[1] ,
    \Tile_X6Y9_EE4BEG[0] }),
    .EE4END({\Tile_X5Y9_EE4BEG[15] ,
    \Tile_X5Y9_EE4BEG[14] ,
    \Tile_X5Y9_EE4BEG[13] ,
    \Tile_X5Y9_EE4BEG[12] ,
    \Tile_X5Y9_EE4BEG[11] ,
    \Tile_X5Y9_EE4BEG[10] ,
    \Tile_X5Y9_EE4BEG[9] ,
    \Tile_X5Y9_EE4BEG[8] ,
    \Tile_X5Y9_EE4BEG[7] ,
    \Tile_X5Y9_EE4BEG[6] ,
    \Tile_X5Y9_EE4BEG[5] ,
    \Tile_X5Y9_EE4BEG[4] ,
    \Tile_X5Y9_EE4BEG[3] ,
    \Tile_X5Y9_EE4BEG[2] ,
    \Tile_X5Y9_EE4BEG[1] ,
    \Tile_X5Y9_EE4BEG[0] }),
    .FrameData({\Tile_X5Y9_FrameData_O[31] ,
    \Tile_X5Y9_FrameData_O[30] ,
    \Tile_X5Y9_FrameData_O[29] ,
    \Tile_X5Y9_FrameData_O[28] ,
    \Tile_X5Y9_FrameData_O[27] ,
    \Tile_X5Y9_FrameData_O[26] ,
    \Tile_X5Y9_FrameData_O[25] ,
    \Tile_X5Y9_FrameData_O[24] ,
    \Tile_X5Y9_FrameData_O[23] ,
    \Tile_X5Y9_FrameData_O[22] ,
    \Tile_X5Y9_FrameData_O[21] ,
    \Tile_X5Y9_FrameData_O[20] ,
    \Tile_X5Y9_FrameData_O[19] ,
    \Tile_X5Y9_FrameData_O[18] ,
    \Tile_X5Y9_FrameData_O[17] ,
    \Tile_X5Y9_FrameData_O[16] ,
    \Tile_X5Y9_FrameData_O[15] ,
    \Tile_X5Y9_FrameData_O[14] ,
    \Tile_X5Y9_FrameData_O[13] ,
    \Tile_X5Y9_FrameData_O[12] ,
    \Tile_X5Y9_FrameData_O[11] ,
    \Tile_X5Y9_FrameData_O[10] ,
    \Tile_X5Y9_FrameData_O[9] ,
    \Tile_X5Y9_FrameData_O[8] ,
    \Tile_X5Y9_FrameData_O[7] ,
    \Tile_X5Y9_FrameData_O[6] ,
    \Tile_X5Y9_FrameData_O[5] ,
    \Tile_X5Y9_FrameData_O[4] ,
    \Tile_X5Y9_FrameData_O[3] ,
    \Tile_X5Y9_FrameData_O[2] ,
    \Tile_X5Y9_FrameData_O[1] ,
    \Tile_X5Y9_FrameData_O[0] }),
    .FrameData_O({\Tile_X6Y9_FrameData_O[31] ,
    \Tile_X6Y9_FrameData_O[30] ,
    \Tile_X6Y9_FrameData_O[29] ,
    \Tile_X6Y9_FrameData_O[28] ,
    \Tile_X6Y9_FrameData_O[27] ,
    \Tile_X6Y9_FrameData_O[26] ,
    \Tile_X6Y9_FrameData_O[25] ,
    \Tile_X6Y9_FrameData_O[24] ,
    \Tile_X6Y9_FrameData_O[23] ,
    \Tile_X6Y9_FrameData_O[22] ,
    \Tile_X6Y9_FrameData_O[21] ,
    \Tile_X6Y9_FrameData_O[20] ,
    \Tile_X6Y9_FrameData_O[19] ,
    \Tile_X6Y9_FrameData_O[18] ,
    \Tile_X6Y9_FrameData_O[17] ,
    \Tile_X6Y9_FrameData_O[16] ,
    \Tile_X6Y9_FrameData_O[15] ,
    \Tile_X6Y9_FrameData_O[14] ,
    \Tile_X6Y9_FrameData_O[13] ,
    \Tile_X6Y9_FrameData_O[12] ,
    \Tile_X6Y9_FrameData_O[11] ,
    \Tile_X6Y9_FrameData_O[10] ,
    \Tile_X6Y9_FrameData_O[9] ,
    \Tile_X6Y9_FrameData_O[8] ,
    \Tile_X6Y9_FrameData_O[7] ,
    \Tile_X6Y9_FrameData_O[6] ,
    \Tile_X6Y9_FrameData_O[5] ,
    \Tile_X6Y9_FrameData_O[4] ,
    \Tile_X6Y9_FrameData_O[3] ,
    \Tile_X6Y9_FrameData_O[2] ,
    \Tile_X6Y9_FrameData_O[1] ,
    \Tile_X6Y9_FrameData_O[0] }),
    .FrameStrobe({\Tile_X6Y10_FrameStrobe_O[19] ,
    \Tile_X6Y10_FrameStrobe_O[18] ,
    \Tile_X6Y10_FrameStrobe_O[17] ,
    \Tile_X6Y10_FrameStrobe_O[16] ,
    \Tile_X6Y10_FrameStrobe_O[15] ,
    \Tile_X6Y10_FrameStrobe_O[14] ,
    \Tile_X6Y10_FrameStrobe_O[13] ,
    \Tile_X6Y10_FrameStrobe_O[12] ,
    \Tile_X6Y10_FrameStrobe_O[11] ,
    \Tile_X6Y10_FrameStrobe_O[10] ,
    \Tile_X6Y10_FrameStrobe_O[9] ,
    \Tile_X6Y10_FrameStrobe_O[8] ,
    \Tile_X6Y10_FrameStrobe_O[7] ,
    \Tile_X6Y10_FrameStrobe_O[6] ,
    \Tile_X6Y10_FrameStrobe_O[5] ,
    \Tile_X6Y10_FrameStrobe_O[4] ,
    \Tile_X6Y10_FrameStrobe_O[3] ,
    \Tile_X6Y10_FrameStrobe_O[2] ,
    \Tile_X6Y10_FrameStrobe_O[1] ,
    \Tile_X6Y10_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X6Y9_FrameStrobe_O[19] ,
    \Tile_X6Y9_FrameStrobe_O[18] ,
    \Tile_X6Y9_FrameStrobe_O[17] ,
    \Tile_X6Y9_FrameStrobe_O[16] ,
    \Tile_X6Y9_FrameStrobe_O[15] ,
    \Tile_X6Y9_FrameStrobe_O[14] ,
    \Tile_X6Y9_FrameStrobe_O[13] ,
    \Tile_X6Y9_FrameStrobe_O[12] ,
    \Tile_X6Y9_FrameStrobe_O[11] ,
    \Tile_X6Y9_FrameStrobe_O[10] ,
    \Tile_X6Y9_FrameStrobe_O[9] ,
    \Tile_X6Y9_FrameStrobe_O[8] ,
    \Tile_X6Y9_FrameStrobe_O[7] ,
    \Tile_X6Y9_FrameStrobe_O[6] ,
    \Tile_X6Y9_FrameStrobe_O[5] ,
    \Tile_X6Y9_FrameStrobe_O[4] ,
    \Tile_X6Y9_FrameStrobe_O[3] ,
    \Tile_X6Y9_FrameStrobe_O[2] ,
    \Tile_X6Y9_FrameStrobe_O[1] ,
    \Tile_X6Y9_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X6Y9_N1BEG[3] ,
    \Tile_X6Y9_N1BEG[2] ,
    \Tile_X6Y9_N1BEG[1] ,
    \Tile_X6Y9_N1BEG[0] }),
    .N1END({\Tile_X6Y10_N1BEG[3] ,
    \Tile_X6Y10_N1BEG[2] ,
    \Tile_X6Y10_N1BEG[1] ,
    \Tile_X6Y10_N1BEG[0] }),
    .N2BEG({\Tile_X6Y9_N2BEG[7] ,
    \Tile_X6Y9_N2BEG[6] ,
    \Tile_X6Y9_N2BEG[5] ,
    \Tile_X6Y9_N2BEG[4] ,
    \Tile_X6Y9_N2BEG[3] ,
    \Tile_X6Y9_N2BEG[2] ,
    \Tile_X6Y9_N2BEG[1] ,
    \Tile_X6Y9_N2BEG[0] }),
    .N2BEGb({\Tile_X6Y9_N2BEGb[7] ,
    \Tile_X6Y9_N2BEGb[6] ,
    \Tile_X6Y9_N2BEGb[5] ,
    \Tile_X6Y9_N2BEGb[4] ,
    \Tile_X6Y9_N2BEGb[3] ,
    \Tile_X6Y9_N2BEGb[2] ,
    \Tile_X6Y9_N2BEGb[1] ,
    \Tile_X6Y9_N2BEGb[0] }),
    .N2END({\Tile_X6Y10_N2BEGb[7] ,
    \Tile_X6Y10_N2BEGb[6] ,
    \Tile_X6Y10_N2BEGb[5] ,
    \Tile_X6Y10_N2BEGb[4] ,
    \Tile_X6Y10_N2BEGb[3] ,
    \Tile_X6Y10_N2BEGb[2] ,
    \Tile_X6Y10_N2BEGb[1] ,
    \Tile_X6Y10_N2BEGb[0] }),
    .N2MID({\Tile_X6Y10_N2BEG[7] ,
    \Tile_X6Y10_N2BEG[6] ,
    \Tile_X6Y10_N2BEG[5] ,
    \Tile_X6Y10_N2BEG[4] ,
    \Tile_X6Y10_N2BEG[3] ,
    \Tile_X6Y10_N2BEG[2] ,
    \Tile_X6Y10_N2BEG[1] ,
    \Tile_X6Y10_N2BEG[0] }),
    .N4BEG({\Tile_X6Y9_N4BEG[15] ,
    \Tile_X6Y9_N4BEG[14] ,
    \Tile_X6Y9_N4BEG[13] ,
    \Tile_X6Y9_N4BEG[12] ,
    \Tile_X6Y9_N4BEG[11] ,
    \Tile_X6Y9_N4BEG[10] ,
    \Tile_X6Y9_N4BEG[9] ,
    \Tile_X6Y9_N4BEG[8] ,
    \Tile_X6Y9_N4BEG[7] ,
    \Tile_X6Y9_N4BEG[6] ,
    \Tile_X6Y9_N4BEG[5] ,
    \Tile_X6Y9_N4BEG[4] ,
    \Tile_X6Y9_N4BEG[3] ,
    \Tile_X6Y9_N4BEG[2] ,
    \Tile_X6Y9_N4BEG[1] ,
    \Tile_X6Y9_N4BEG[0] }),
    .N4END({\Tile_X6Y10_N4BEG[15] ,
    \Tile_X6Y10_N4BEG[14] ,
    \Tile_X6Y10_N4BEG[13] ,
    \Tile_X6Y10_N4BEG[12] ,
    \Tile_X6Y10_N4BEG[11] ,
    \Tile_X6Y10_N4BEG[10] ,
    \Tile_X6Y10_N4BEG[9] ,
    \Tile_X6Y10_N4BEG[8] ,
    \Tile_X6Y10_N4BEG[7] ,
    \Tile_X6Y10_N4BEG[6] ,
    \Tile_X6Y10_N4BEG[5] ,
    \Tile_X6Y10_N4BEG[4] ,
    \Tile_X6Y10_N4BEG[3] ,
    \Tile_X6Y10_N4BEG[2] ,
    \Tile_X6Y10_N4BEG[1] ,
    \Tile_X6Y10_N4BEG[0] }),
    .NN4BEG({\Tile_X6Y9_NN4BEG[15] ,
    \Tile_X6Y9_NN4BEG[14] ,
    \Tile_X6Y9_NN4BEG[13] ,
    \Tile_X6Y9_NN4BEG[12] ,
    \Tile_X6Y9_NN4BEG[11] ,
    \Tile_X6Y9_NN4BEG[10] ,
    \Tile_X6Y9_NN4BEG[9] ,
    \Tile_X6Y9_NN4BEG[8] ,
    \Tile_X6Y9_NN4BEG[7] ,
    \Tile_X6Y9_NN4BEG[6] ,
    \Tile_X6Y9_NN4BEG[5] ,
    \Tile_X6Y9_NN4BEG[4] ,
    \Tile_X6Y9_NN4BEG[3] ,
    \Tile_X6Y9_NN4BEG[2] ,
    \Tile_X6Y9_NN4BEG[1] ,
    \Tile_X6Y9_NN4BEG[0] }),
    .NN4END({\Tile_X6Y10_NN4BEG[15] ,
    \Tile_X6Y10_NN4BEG[14] ,
    \Tile_X6Y10_NN4BEG[13] ,
    \Tile_X6Y10_NN4BEG[12] ,
    \Tile_X6Y10_NN4BEG[11] ,
    \Tile_X6Y10_NN4BEG[10] ,
    \Tile_X6Y10_NN4BEG[9] ,
    \Tile_X6Y10_NN4BEG[8] ,
    \Tile_X6Y10_NN4BEG[7] ,
    \Tile_X6Y10_NN4BEG[6] ,
    \Tile_X6Y10_NN4BEG[5] ,
    \Tile_X6Y10_NN4BEG[4] ,
    \Tile_X6Y10_NN4BEG[3] ,
    \Tile_X6Y10_NN4BEG[2] ,
    \Tile_X6Y10_NN4BEG[1] ,
    \Tile_X6Y10_NN4BEG[0] }),
    .S1BEG({\Tile_X6Y9_S1BEG[3] ,
    \Tile_X6Y9_S1BEG[2] ,
    \Tile_X6Y9_S1BEG[1] ,
    \Tile_X6Y9_S1BEG[0] }),
    .S1END({\Tile_X6Y8_S1BEG[3] ,
    \Tile_X6Y8_S1BEG[2] ,
    \Tile_X6Y8_S1BEG[1] ,
    \Tile_X6Y8_S1BEG[0] }),
    .S2BEG({\Tile_X6Y9_S2BEG[7] ,
    \Tile_X6Y9_S2BEG[6] ,
    \Tile_X6Y9_S2BEG[5] ,
    \Tile_X6Y9_S2BEG[4] ,
    \Tile_X6Y9_S2BEG[3] ,
    \Tile_X6Y9_S2BEG[2] ,
    \Tile_X6Y9_S2BEG[1] ,
    \Tile_X6Y9_S2BEG[0] }),
    .S2BEGb({\Tile_X6Y9_S2BEGb[7] ,
    \Tile_X6Y9_S2BEGb[6] ,
    \Tile_X6Y9_S2BEGb[5] ,
    \Tile_X6Y9_S2BEGb[4] ,
    \Tile_X6Y9_S2BEGb[3] ,
    \Tile_X6Y9_S2BEGb[2] ,
    \Tile_X6Y9_S2BEGb[1] ,
    \Tile_X6Y9_S2BEGb[0] }),
    .S2END({\Tile_X6Y8_S2BEGb[7] ,
    \Tile_X6Y8_S2BEGb[6] ,
    \Tile_X6Y8_S2BEGb[5] ,
    \Tile_X6Y8_S2BEGb[4] ,
    \Tile_X6Y8_S2BEGb[3] ,
    \Tile_X6Y8_S2BEGb[2] ,
    \Tile_X6Y8_S2BEGb[1] ,
    \Tile_X6Y8_S2BEGb[0] }),
    .S2MID({\Tile_X6Y8_S2BEG[7] ,
    \Tile_X6Y8_S2BEG[6] ,
    \Tile_X6Y8_S2BEG[5] ,
    \Tile_X6Y8_S2BEG[4] ,
    \Tile_X6Y8_S2BEG[3] ,
    \Tile_X6Y8_S2BEG[2] ,
    \Tile_X6Y8_S2BEG[1] ,
    \Tile_X6Y8_S2BEG[0] }),
    .S4BEG({\Tile_X6Y9_S4BEG[15] ,
    \Tile_X6Y9_S4BEG[14] ,
    \Tile_X6Y9_S4BEG[13] ,
    \Tile_X6Y9_S4BEG[12] ,
    \Tile_X6Y9_S4BEG[11] ,
    \Tile_X6Y9_S4BEG[10] ,
    \Tile_X6Y9_S4BEG[9] ,
    \Tile_X6Y9_S4BEG[8] ,
    \Tile_X6Y9_S4BEG[7] ,
    \Tile_X6Y9_S4BEG[6] ,
    \Tile_X6Y9_S4BEG[5] ,
    \Tile_X6Y9_S4BEG[4] ,
    \Tile_X6Y9_S4BEG[3] ,
    \Tile_X6Y9_S4BEG[2] ,
    \Tile_X6Y9_S4BEG[1] ,
    \Tile_X6Y9_S4BEG[0] }),
    .S4END({\Tile_X6Y8_S4BEG[15] ,
    \Tile_X6Y8_S4BEG[14] ,
    \Tile_X6Y8_S4BEG[13] ,
    \Tile_X6Y8_S4BEG[12] ,
    \Tile_X6Y8_S4BEG[11] ,
    \Tile_X6Y8_S4BEG[10] ,
    \Tile_X6Y8_S4BEG[9] ,
    \Tile_X6Y8_S4BEG[8] ,
    \Tile_X6Y8_S4BEG[7] ,
    \Tile_X6Y8_S4BEG[6] ,
    \Tile_X6Y8_S4BEG[5] ,
    \Tile_X6Y8_S4BEG[4] ,
    \Tile_X6Y8_S4BEG[3] ,
    \Tile_X6Y8_S4BEG[2] ,
    \Tile_X6Y8_S4BEG[1] ,
    \Tile_X6Y8_S4BEG[0] }),
    .SS4BEG({\Tile_X6Y9_SS4BEG[15] ,
    \Tile_X6Y9_SS4BEG[14] ,
    \Tile_X6Y9_SS4BEG[13] ,
    \Tile_X6Y9_SS4BEG[12] ,
    \Tile_X6Y9_SS4BEG[11] ,
    \Tile_X6Y9_SS4BEG[10] ,
    \Tile_X6Y9_SS4BEG[9] ,
    \Tile_X6Y9_SS4BEG[8] ,
    \Tile_X6Y9_SS4BEG[7] ,
    \Tile_X6Y9_SS4BEG[6] ,
    \Tile_X6Y9_SS4BEG[5] ,
    \Tile_X6Y9_SS4BEG[4] ,
    \Tile_X6Y9_SS4BEG[3] ,
    \Tile_X6Y9_SS4BEG[2] ,
    \Tile_X6Y9_SS4BEG[1] ,
    \Tile_X6Y9_SS4BEG[0] }),
    .SS4END({\Tile_X6Y8_SS4BEG[15] ,
    \Tile_X6Y8_SS4BEG[14] ,
    \Tile_X6Y8_SS4BEG[13] ,
    \Tile_X6Y8_SS4BEG[12] ,
    \Tile_X6Y8_SS4BEG[11] ,
    \Tile_X6Y8_SS4BEG[10] ,
    \Tile_X6Y8_SS4BEG[9] ,
    \Tile_X6Y8_SS4BEG[8] ,
    \Tile_X6Y8_SS4BEG[7] ,
    \Tile_X6Y8_SS4BEG[6] ,
    \Tile_X6Y8_SS4BEG[5] ,
    \Tile_X6Y8_SS4BEG[4] ,
    \Tile_X6Y8_SS4BEG[3] ,
    \Tile_X6Y8_SS4BEG[2] ,
    \Tile_X6Y8_SS4BEG[1] ,
    \Tile_X6Y8_SS4BEG[0] }),
    .W1BEG({\Tile_X6Y9_W1BEG[3] ,
    \Tile_X6Y9_W1BEG[2] ,
    \Tile_X6Y9_W1BEG[1] ,
    \Tile_X6Y9_W1BEG[0] }),
    .W1END({\Tile_X7Y9_W1BEG[3] ,
    \Tile_X7Y9_W1BEG[2] ,
    \Tile_X7Y9_W1BEG[1] ,
    \Tile_X7Y9_W1BEG[0] }),
    .W2BEG({\Tile_X6Y9_W2BEG[7] ,
    \Tile_X6Y9_W2BEG[6] ,
    \Tile_X6Y9_W2BEG[5] ,
    \Tile_X6Y9_W2BEG[4] ,
    \Tile_X6Y9_W2BEG[3] ,
    \Tile_X6Y9_W2BEG[2] ,
    \Tile_X6Y9_W2BEG[1] ,
    \Tile_X6Y9_W2BEG[0] }),
    .W2BEGb({\Tile_X6Y9_W2BEGb[7] ,
    \Tile_X6Y9_W2BEGb[6] ,
    \Tile_X6Y9_W2BEGb[5] ,
    \Tile_X6Y9_W2BEGb[4] ,
    \Tile_X6Y9_W2BEGb[3] ,
    \Tile_X6Y9_W2BEGb[2] ,
    \Tile_X6Y9_W2BEGb[1] ,
    \Tile_X6Y9_W2BEGb[0] }),
    .W2END({\Tile_X7Y9_W2BEGb[7] ,
    \Tile_X7Y9_W2BEGb[6] ,
    \Tile_X7Y9_W2BEGb[5] ,
    \Tile_X7Y9_W2BEGb[4] ,
    \Tile_X7Y9_W2BEGb[3] ,
    \Tile_X7Y9_W2BEGb[2] ,
    \Tile_X7Y9_W2BEGb[1] ,
    \Tile_X7Y9_W2BEGb[0] }),
    .W2MID({\Tile_X7Y9_W2BEG[7] ,
    \Tile_X7Y9_W2BEG[6] ,
    \Tile_X7Y9_W2BEG[5] ,
    \Tile_X7Y9_W2BEG[4] ,
    \Tile_X7Y9_W2BEG[3] ,
    \Tile_X7Y9_W2BEG[2] ,
    \Tile_X7Y9_W2BEG[1] ,
    \Tile_X7Y9_W2BEG[0] }),
    .W6BEG({\Tile_X6Y9_W6BEG[11] ,
    \Tile_X6Y9_W6BEG[10] ,
    \Tile_X6Y9_W6BEG[9] ,
    \Tile_X6Y9_W6BEG[8] ,
    \Tile_X6Y9_W6BEG[7] ,
    \Tile_X6Y9_W6BEG[6] ,
    \Tile_X6Y9_W6BEG[5] ,
    \Tile_X6Y9_W6BEG[4] ,
    \Tile_X6Y9_W6BEG[3] ,
    \Tile_X6Y9_W6BEG[2] ,
    \Tile_X6Y9_W6BEG[1] ,
    \Tile_X6Y9_W6BEG[0] }),
    .W6END({\Tile_X7Y9_W6BEG[11] ,
    \Tile_X7Y9_W6BEG[10] ,
    \Tile_X7Y9_W6BEG[9] ,
    \Tile_X7Y9_W6BEG[8] ,
    \Tile_X7Y9_W6BEG[7] ,
    \Tile_X7Y9_W6BEG[6] ,
    \Tile_X7Y9_W6BEG[5] ,
    \Tile_X7Y9_W6BEG[4] ,
    \Tile_X7Y9_W6BEG[3] ,
    \Tile_X7Y9_W6BEG[2] ,
    \Tile_X7Y9_W6BEG[1] ,
    \Tile_X7Y9_W6BEG[0] }),
    .WW4BEG({\Tile_X6Y9_WW4BEG[15] ,
    \Tile_X6Y9_WW4BEG[14] ,
    \Tile_X6Y9_WW4BEG[13] ,
    \Tile_X6Y9_WW4BEG[12] ,
    \Tile_X6Y9_WW4BEG[11] ,
    \Tile_X6Y9_WW4BEG[10] ,
    \Tile_X6Y9_WW4BEG[9] ,
    \Tile_X6Y9_WW4BEG[8] ,
    \Tile_X6Y9_WW4BEG[7] ,
    \Tile_X6Y9_WW4BEG[6] ,
    \Tile_X6Y9_WW4BEG[5] ,
    \Tile_X6Y9_WW4BEG[4] ,
    \Tile_X6Y9_WW4BEG[3] ,
    \Tile_X6Y9_WW4BEG[2] ,
    \Tile_X6Y9_WW4BEG[1] ,
    \Tile_X6Y9_WW4BEG[0] }),
    .WW4END({\Tile_X7Y9_WW4BEG[15] ,
    \Tile_X7Y9_WW4BEG[14] ,
    \Tile_X7Y9_WW4BEG[13] ,
    \Tile_X7Y9_WW4BEG[12] ,
    \Tile_X7Y9_WW4BEG[11] ,
    \Tile_X7Y9_WW4BEG[10] ,
    \Tile_X7Y9_WW4BEG[9] ,
    \Tile_X7Y9_WW4BEG[8] ,
    \Tile_X7Y9_WW4BEG[7] ,
    \Tile_X7Y9_WW4BEG[6] ,
    \Tile_X7Y9_WW4BEG[5] ,
    \Tile_X7Y9_WW4BEG[4] ,
    \Tile_X7Y9_WW4BEG[3] ,
    \Tile_X7Y9_WW4BEG[2] ,
    \Tile_X7Y9_WW4BEG[1] ,
    \Tile_X7Y9_WW4BEG[0] }));
 N_term_DSP Tile_X7Y0_N_term_DSP (.UserCLK(Tile_X7Y1_UserCLKo),
    .UserCLKo(Tile_X7Y0_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .FrameData({\Tile_X6Y0_FrameData_O[31] ,
    \Tile_X6Y0_FrameData_O[30] ,
    \Tile_X6Y0_FrameData_O[29] ,
    \Tile_X6Y0_FrameData_O[28] ,
    \Tile_X6Y0_FrameData_O[27] ,
    \Tile_X6Y0_FrameData_O[26] ,
    \Tile_X6Y0_FrameData_O[25] ,
    \Tile_X6Y0_FrameData_O[24] ,
    \Tile_X6Y0_FrameData_O[23] ,
    \Tile_X6Y0_FrameData_O[22] ,
    \Tile_X6Y0_FrameData_O[21] ,
    \Tile_X6Y0_FrameData_O[20] ,
    \Tile_X6Y0_FrameData_O[19] ,
    \Tile_X6Y0_FrameData_O[18] ,
    \Tile_X6Y0_FrameData_O[17] ,
    \Tile_X6Y0_FrameData_O[16] ,
    \Tile_X6Y0_FrameData_O[15] ,
    \Tile_X6Y0_FrameData_O[14] ,
    \Tile_X6Y0_FrameData_O[13] ,
    \Tile_X6Y0_FrameData_O[12] ,
    \Tile_X6Y0_FrameData_O[11] ,
    \Tile_X6Y0_FrameData_O[10] ,
    \Tile_X6Y0_FrameData_O[9] ,
    \Tile_X6Y0_FrameData_O[8] ,
    \Tile_X6Y0_FrameData_O[7] ,
    \Tile_X6Y0_FrameData_O[6] ,
    \Tile_X6Y0_FrameData_O[5] ,
    \Tile_X6Y0_FrameData_O[4] ,
    \Tile_X6Y0_FrameData_O[3] ,
    \Tile_X6Y0_FrameData_O[2] ,
    \Tile_X6Y0_FrameData_O[1] ,
    \Tile_X6Y0_FrameData_O[0] }),
    .FrameData_O({\Tile_X7Y0_FrameData_O[31] ,
    \Tile_X7Y0_FrameData_O[30] ,
    \Tile_X7Y0_FrameData_O[29] ,
    \Tile_X7Y0_FrameData_O[28] ,
    \Tile_X7Y0_FrameData_O[27] ,
    \Tile_X7Y0_FrameData_O[26] ,
    \Tile_X7Y0_FrameData_O[25] ,
    \Tile_X7Y0_FrameData_O[24] ,
    \Tile_X7Y0_FrameData_O[23] ,
    \Tile_X7Y0_FrameData_O[22] ,
    \Tile_X7Y0_FrameData_O[21] ,
    \Tile_X7Y0_FrameData_O[20] ,
    \Tile_X7Y0_FrameData_O[19] ,
    \Tile_X7Y0_FrameData_O[18] ,
    \Tile_X7Y0_FrameData_O[17] ,
    \Tile_X7Y0_FrameData_O[16] ,
    \Tile_X7Y0_FrameData_O[15] ,
    \Tile_X7Y0_FrameData_O[14] ,
    \Tile_X7Y0_FrameData_O[13] ,
    \Tile_X7Y0_FrameData_O[12] ,
    \Tile_X7Y0_FrameData_O[11] ,
    \Tile_X7Y0_FrameData_O[10] ,
    \Tile_X7Y0_FrameData_O[9] ,
    \Tile_X7Y0_FrameData_O[8] ,
    \Tile_X7Y0_FrameData_O[7] ,
    \Tile_X7Y0_FrameData_O[6] ,
    \Tile_X7Y0_FrameData_O[5] ,
    \Tile_X7Y0_FrameData_O[4] ,
    \Tile_X7Y0_FrameData_O[3] ,
    \Tile_X7Y0_FrameData_O[2] ,
    \Tile_X7Y0_FrameData_O[1] ,
    \Tile_X7Y0_FrameData_O[0] }),
    .FrameStrobe({\Tile_X7Y1_FrameStrobe_O[19] ,
    \Tile_X7Y1_FrameStrobe_O[18] ,
    \Tile_X7Y1_FrameStrobe_O[17] ,
    \Tile_X7Y1_FrameStrobe_O[16] ,
    \Tile_X7Y1_FrameStrobe_O[15] ,
    \Tile_X7Y1_FrameStrobe_O[14] ,
    \Tile_X7Y1_FrameStrobe_O[13] ,
    \Tile_X7Y1_FrameStrobe_O[12] ,
    \Tile_X7Y1_FrameStrobe_O[11] ,
    \Tile_X7Y1_FrameStrobe_O[10] ,
    \Tile_X7Y1_FrameStrobe_O[9] ,
    \Tile_X7Y1_FrameStrobe_O[8] ,
    \Tile_X7Y1_FrameStrobe_O[7] ,
    \Tile_X7Y1_FrameStrobe_O[6] ,
    \Tile_X7Y1_FrameStrobe_O[5] ,
    \Tile_X7Y1_FrameStrobe_O[4] ,
    \Tile_X7Y1_FrameStrobe_O[3] ,
    \Tile_X7Y1_FrameStrobe_O[2] ,
    \Tile_X7Y1_FrameStrobe_O[1] ,
    \Tile_X7Y1_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X7Y0_FrameStrobe_O[19] ,
    \Tile_X7Y0_FrameStrobe_O[18] ,
    \Tile_X7Y0_FrameStrobe_O[17] ,
    \Tile_X7Y0_FrameStrobe_O[16] ,
    \Tile_X7Y0_FrameStrobe_O[15] ,
    \Tile_X7Y0_FrameStrobe_O[14] ,
    \Tile_X7Y0_FrameStrobe_O[13] ,
    \Tile_X7Y0_FrameStrobe_O[12] ,
    \Tile_X7Y0_FrameStrobe_O[11] ,
    \Tile_X7Y0_FrameStrobe_O[10] ,
    \Tile_X7Y0_FrameStrobe_O[9] ,
    \Tile_X7Y0_FrameStrobe_O[8] ,
    \Tile_X7Y0_FrameStrobe_O[7] ,
    \Tile_X7Y0_FrameStrobe_O[6] ,
    \Tile_X7Y0_FrameStrobe_O[5] ,
    \Tile_X7Y0_FrameStrobe_O[4] ,
    \Tile_X7Y0_FrameStrobe_O[3] ,
    \Tile_X7Y0_FrameStrobe_O[2] ,
    \Tile_X7Y0_FrameStrobe_O[1] ,
    \Tile_X7Y0_FrameStrobe_O[0] }),
    .N1END({\Tile_X7Y1_N1BEG[3] ,
    \Tile_X7Y1_N1BEG[2] ,
    \Tile_X7Y1_N1BEG[1] ,
    \Tile_X7Y1_N1BEG[0] }),
    .N2END({\Tile_X7Y1_N2BEGb[7] ,
    \Tile_X7Y1_N2BEGb[6] ,
    \Tile_X7Y1_N2BEGb[5] ,
    \Tile_X7Y1_N2BEGb[4] ,
    \Tile_X7Y1_N2BEGb[3] ,
    \Tile_X7Y1_N2BEGb[2] ,
    \Tile_X7Y1_N2BEGb[1] ,
    \Tile_X7Y1_N2BEGb[0] }),
    .N2MID({\Tile_X7Y1_N2BEG[7] ,
    \Tile_X7Y1_N2BEG[6] ,
    \Tile_X7Y1_N2BEG[5] ,
    \Tile_X7Y1_N2BEG[4] ,
    \Tile_X7Y1_N2BEG[3] ,
    \Tile_X7Y1_N2BEG[2] ,
    \Tile_X7Y1_N2BEG[1] ,
    \Tile_X7Y1_N2BEG[0] }),
    .N4END({\Tile_X7Y1_N4BEG[15] ,
    \Tile_X7Y1_N4BEG[14] ,
    \Tile_X7Y1_N4BEG[13] ,
    \Tile_X7Y1_N4BEG[12] ,
    \Tile_X7Y1_N4BEG[11] ,
    \Tile_X7Y1_N4BEG[10] ,
    \Tile_X7Y1_N4BEG[9] ,
    \Tile_X7Y1_N4BEG[8] ,
    \Tile_X7Y1_N4BEG[7] ,
    \Tile_X7Y1_N4BEG[6] ,
    \Tile_X7Y1_N4BEG[5] ,
    \Tile_X7Y1_N4BEG[4] ,
    \Tile_X7Y1_N4BEG[3] ,
    \Tile_X7Y1_N4BEG[2] ,
    \Tile_X7Y1_N4BEG[1] ,
    \Tile_X7Y1_N4BEG[0] }),
    .NN4END({\Tile_X7Y1_NN4BEG[15] ,
    \Tile_X7Y1_NN4BEG[14] ,
    \Tile_X7Y1_NN4BEG[13] ,
    \Tile_X7Y1_NN4BEG[12] ,
    \Tile_X7Y1_NN4BEG[11] ,
    \Tile_X7Y1_NN4BEG[10] ,
    \Tile_X7Y1_NN4BEG[9] ,
    \Tile_X7Y1_NN4BEG[8] ,
    \Tile_X7Y1_NN4BEG[7] ,
    \Tile_X7Y1_NN4BEG[6] ,
    \Tile_X7Y1_NN4BEG[5] ,
    \Tile_X7Y1_NN4BEG[4] ,
    \Tile_X7Y1_NN4BEG[3] ,
    \Tile_X7Y1_NN4BEG[2] ,
    \Tile_X7Y1_NN4BEG[1] ,
    \Tile_X7Y1_NN4BEG[0] }),
    .S1BEG({\Tile_X7Y0_S1BEG[3] ,
    \Tile_X7Y0_S1BEG[2] ,
    \Tile_X7Y0_S1BEG[1] ,
    \Tile_X7Y0_S1BEG[0] }),
    .S2BEG({\Tile_X7Y0_S2BEG[7] ,
    \Tile_X7Y0_S2BEG[6] ,
    \Tile_X7Y0_S2BEG[5] ,
    \Tile_X7Y0_S2BEG[4] ,
    \Tile_X7Y0_S2BEG[3] ,
    \Tile_X7Y0_S2BEG[2] ,
    \Tile_X7Y0_S2BEG[1] ,
    \Tile_X7Y0_S2BEG[0] }),
    .S2BEGb({\Tile_X7Y0_S2BEGb[7] ,
    \Tile_X7Y0_S2BEGb[6] ,
    \Tile_X7Y0_S2BEGb[5] ,
    \Tile_X7Y0_S2BEGb[4] ,
    \Tile_X7Y0_S2BEGb[3] ,
    \Tile_X7Y0_S2BEGb[2] ,
    \Tile_X7Y0_S2BEGb[1] ,
    \Tile_X7Y0_S2BEGb[0] }),
    .S4BEG({\Tile_X7Y0_S4BEG[15] ,
    \Tile_X7Y0_S4BEG[14] ,
    \Tile_X7Y0_S4BEG[13] ,
    \Tile_X7Y0_S4BEG[12] ,
    \Tile_X7Y0_S4BEG[11] ,
    \Tile_X7Y0_S4BEG[10] ,
    \Tile_X7Y0_S4BEG[9] ,
    \Tile_X7Y0_S4BEG[8] ,
    \Tile_X7Y0_S4BEG[7] ,
    \Tile_X7Y0_S4BEG[6] ,
    \Tile_X7Y0_S4BEG[5] ,
    \Tile_X7Y0_S4BEG[4] ,
    \Tile_X7Y0_S4BEG[3] ,
    \Tile_X7Y0_S4BEG[2] ,
    \Tile_X7Y0_S4BEG[1] ,
    \Tile_X7Y0_S4BEG[0] }),
    .SS4BEG({\Tile_X7Y0_SS4BEG[15] ,
    \Tile_X7Y0_SS4BEG[14] ,
    \Tile_X7Y0_SS4BEG[13] ,
    \Tile_X7Y0_SS4BEG[12] ,
    \Tile_X7Y0_SS4BEG[11] ,
    \Tile_X7Y0_SS4BEG[10] ,
    \Tile_X7Y0_SS4BEG[9] ,
    \Tile_X7Y0_SS4BEG[8] ,
    \Tile_X7Y0_SS4BEG[7] ,
    \Tile_X7Y0_SS4BEG[6] ,
    \Tile_X7Y0_SS4BEG[5] ,
    \Tile_X7Y0_SS4BEG[4] ,
    \Tile_X7Y0_SS4BEG[3] ,
    \Tile_X7Y0_SS4BEG[2] ,
    \Tile_X7Y0_SS4BEG[1] ,
    \Tile_X7Y0_SS4BEG[0] }));
 DSP Tile_X7Y11_DSP (.Tile_X0Y0_UserCLKo(Tile_X7Y11_UserCLKo),
    .Tile_X0Y1_UserCLK(Tile_X7Y13_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .Tile_X0Y0_E1BEG({\Tile_X7Y11_E1BEG[3] ,
    \Tile_X7Y11_E1BEG[2] ,
    \Tile_X7Y11_E1BEG[1] ,
    \Tile_X7Y11_E1BEG[0] }),
    .Tile_X0Y0_E1END({\Tile_X6Y11_E1BEG[3] ,
    \Tile_X6Y11_E1BEG[2] ,
    \Tile_X6Y11_E1BEG[1] ,
    \Tile_X6Y11_E1BEG[0] }),
    .Tile_X0Y0_E2BEG({\Tile_X7Y11_E2BEG[7] ,
    \Tile_X7Y11_E2BEG[6] ,
    \Tile_X7Y11_E2BEG[5] ,
    \Tile_X7Y11_E2BEG[4] ,
    \Tile_X7Y11_E2BEG[3] ,
    \Tile_X7Y11_E2BEG[2] ,
    \Tile_X7Y11_E2BEG[1] ,
    \Tile_X7Y11_E2BEG[0] }),
    .Tile_X0Y0_E2BEGb({\Tile_X7Y11_E2BEGb[7] ,
    \Tile_X7Y11_E2BEGb[6] ,
    \Tile_X7Y11_E2BEGb[5] ,
    \Tile_X7Y11_E2BEGb[4] ,
    \Tile_X7Y11_E2BEGb[3] ,
    \Tile_X7Y11_E2BEGb[2] ,
    \Tile_X7Y11_E2BEGb[1] ,
    \Tile_X7Y11_E2BEGb[0] }),
    .Tile_X0Y0_E2END({\Tile_X6Y11_E2BEGb[7] ,
    \Tile_X6Y11_E2BEGb[6] ,
    \Tile_X6Y11_E2BEGb[5] ,
    \Tile_X6Y11_E2BEGb[4] ,
    \Tile_X6Y11_E2BEGb[3] ,
    \Tile_X6Y11_E2BEGb[2] ,
    \Tile_X6Y11_E2BEGb[1] ,
    \Tile_X6Y11_E2BEGb[0] }),
    .Tile_X0Y0_E2MID({\Tile_X6Y11_E2BEG[7] ,
    \Tile_X6Y11_E2BEG[6] ,
    \Tile_X6Y11_E2BEG[5] ,
    \Tile_X6Y11_E2BEG[4] ,
    \Tile_X6Y11_E2BEG[3] ,
    \Tile_X6Y11_E2BEG[2] ,
    \Tile_X6Y11_E2BEG[1] ,
    \Tile_X6Y11_E2BEG[0] }),
    .Tile_X0Y0_E6BEG({\Tile_X7Y11_E6BEG[11] ,
    \Tile_X7Y11_E6BEG[10] ,
    \Tile_X7Y11_E6BEG[9] ,
    \Tile_X7Y11_E6BEG[8] ,
    \Tile_X7Y11_E6BEG[7] ,
    \Tile_X7Y11_E6BEG[6] ,
    \Tile_X7Y11_E6BEG[5] ,
    \Tile_X7Y11_E6BEG[4] ,
    \Tile_X7Y11_E6BEG[3] ,
    \Tile_X7Y11_E6BEG[2] ,
    \Tile_X7Y11_E6BEG[1] ,
    \Tile_X7Y11_E6BEG[0] }),
    .Tile_X0Y0_E6END({\Tile_X6Y11_E6BEG[11] ,
    \Tile_X6Y11_E6BEG[10] ,
    \Tile_X6Y11_E6BEG[9] ,
    \Tile_X6Y11_E6BEG[8] ,
    \Tile_X6Y11_E6BEG[7] ,
    \Tile_X6Y11_E6BEG[6] ,
    \Tile_X6Y11_E6BEG[5] ,
    \Tile_X6Y11_E6BEG[4] ,
    \Tile_X6Y11_E6BEG[3] ,
    \Tile_X6Y11_E6BEG[2] ,
    \Tile_X6Y11_E6BEG[1] ,
    \Tile_X6Y11_E6BEG[0] }),
    .Tile_X0Y0_EE4BEG({\Tile_X7Y11_EE4BEG[15] ,
    \Tile_X7Y11_EE4BEG[14] ,
    \Tile_X7Y11_EE4BEG[13] ,
    \Tile_X7Y11_EE4BEG[12] ,
    \Tile_X7Y11_EE4BEG[11] ,
    \Tile_X7Y11_EE4BEG[10] ,
    \Tile_X7Y11_EE4BEG[9] ,
    \Tile_X7Y11_EE4BEG[8] ,
    \Tile_X7Y11_EE4BEG[7] ,
    \Tile_X7Y11_EE4BEG[6] ,
    \Tile_X7Y11_EE4BEG[5] ,
    \Tile_X7Y11_EE4BEG[4] ,
    \Tile_X7Y11_EE4BEG[3] ,
    \Tile_X7Y11_EE4BEG[2] ,
    \Tile_X7Y11_EE4BEG[1] ,
    \Tile_X7Y11_EE4BEG[0] }),
    .Tile_X0Y0_EE4END({\Tile_X6Y11_EE4BEG[15] ,
    \Tile_X6Y11_EE4BEG[14] ,
    \Tile_X6Y11_EE4BEG[13] ,
    \Tile_X6Y11_EE4BEG[12] ,
    \Tile_X6Y11_EE4BEG[11] ,
    \Tile_X6Y11_EE4BEG[10] ,
    \Tile_X6Y11_EE4BEG[9] ,
    \Tile_X6Y11_EE4BEG[8] ,
    \Tile_X6Y11_EE4BEG[7] ,
    \Tile_X6Y11_EE4BEG[6] ,
    \Tile_X6Y11_EE4BEG[5] ,
    \Tile_X6Y11_EE4BEG[4] ,
    \Tile_X6Y11_EE4BEG[3] ,
    \Tile_X6Y11_EE4BEG[2] ,
    \Tile_X6Y11_EE4BEG[1] ,
    \Tile_X6Y11_EE4BEG[0] }),
    .Tile_X0Y0_FrameData({\Tile_X6Y11_FrameData_O[31] ,
    \Tile_X6Y11_FrameData_O[30] ,
    \Tile_X6Y11_FrameData_O[29] ,
    \Tile_X6Y11_FrameData_O[28] ,
    \Tile_X6Y11_FrameData_O[27] ,
    \Tile_X6Y11_FrameData_O[26] ,
    \Tile_X6Y11_FrameData_O[25] ,
    \Tile_X6Y11_FrameData_O[24] ,
    \Tile_X6Y11_FrameData_O[23] ,
    \Tile_X6Y11_FrameData_O[22] ,
    \Tile_X6Y11_FrameData_O[21] ,
    \Tile_X6Y11_FrameData_O[20] ,
    \Tile_X6Y11_FrameData_O[19] ,
    \Tile_X6Y11_FrameData_O[18] ,
    \Tile_X6Y11_FrameData_O[17] ,
    \Tile_X6Y11_FrameData_O[16] ,
    \Tile_X6Y11_FrameData_O[15] ,
    \Tile_X6Y11_FrameData_O[14] ,
    \Tile_X6Y11_FrameData_O[13] ,
    \Tile_X6Y11_FrameData_O[12] ,
    \Tile_X6Y11_FrameData_O[11] ,
    \Tile_X6Y11_FrameData_O[10] ,
    \Tile_X6Y11_FrameData_O[9] ,
    \Tile_X6Y11_FrameData_O[8] ,
    \Tile_X6Y11_FrameData_O[7] ,
    \Tile_X6Y11_FrameData_O[6] ,
    \Tile_X6Y11_FrameData_O[5] ,
    \Tile_X6Y11_FrameData_O[4] ,
    \Tile_X6Y11_FrameData_O[3] ,
    \Tile_X6Y11_FrameData_O[2] ,
    \Tile_X6Y11_FrameData_O[1] ,
    \Tile_X6Y11_FrameData_O[0] }),
    .Tile_X0Y0_FrameData_O({\Tile_X7Y11_FrameData_O[31] ,
    \Tile_X7Y11_FrameData_O[30] ,
    \Tile_X7Y11_FrameData_O[29] ,
    \Tile_X7Y11_FrameData_O[28] ,
    \Tile_X7Y11_FrameData_O[27] ,
    \Tile_X7Y11_FrameData_O[26] ,
    \Tile_X7Y11_FrameData_O[25] ,
    \Tile_X7Y11_FrameData_O[24] ,
    \Tile_X7Y11_FrameData_O[23] ,
    \Tile_X7Y11_FrameData_O[22] ,
    \Tile_X7Y11_FrameData_O[21] ,
    \Tile_X7Y11_FrameData_O[20] ,
    \Tile_X7Y11_FrameData_O[19] ,
    \Tile_X7Y11_FrameData_O[18] ,
    \Tile_X7Y11_FrameData_O[17] ,
    \Tile_X7Y11_FrameData_O[16] ,
    \Tile_X7Y11_FrameData_O[15] ,
    \Tile_X7Y11_FrameData_O[14] ,
    \Tile_X7Y11_FrameData_O[13] ,
    \Tile_X7Y11_FrameData_O[12] ,
    \Tile_X7Y11_FrameData_O[11] ,
    \Tile_X7Y11_FrameData_O[10] ,
    \Tile_X7Y11_FrameData_O[9] ,
    \Tile_X7Y11_FrameData_O[8] ,
    \Tile_X7Y11_FrameData_O[7] ,
    \Tile_X7Y11_FrameData_O[6] ,
    \Tile_X7Y11_FrameData_O[5] ,
    \Tile_X7Y11_FrameData_O[4] ,
    \Tile_X7Y11_FrameData_O[3] ,
    \Tile_X7Y11_FrameData_O[2] ,
    \Tile_X7Y11_FrameData_O[1] ,
    \Tile_X7Y11_FrameData_O[0] }),
    .Tile_X0Y0_FrameStrobe_O({\Tile_X7Y11_FrameStrobe_O[19] ,
    \Tile_X7Y11_FrameStrobe_O[18] ,
    \Tile_X7Y11_FrameStrobe_O[17] ,
    \Tile_X7Y11_FrameStrobe_O[16] ,
    \Tile_X7Y11_FrameStrobe_O[15] ,
    \Tile_X7Y11_FrameStrobe_O[14] ,
    \Tile_X7Y11_FrameStrobe_O[13] ,
    \Tile_X7Y11_FrameStrobe_O[12] ,
    \Tile_X7Y11_FrameStrobe_O[11] ,
    \Tile_X7Y11_FrameStrobe_O[10] ,
    \Tile_X7Y11_FrameStrobe_O[9] ,
    \Tile_X7Y11_FrameStrobe_O[8] ,
    \Tile_X7Y11_FrameStrobe_O[7] ,
    \Tile_X7Y11_FrameStrobe_O[6] ,
    \Tile_X7Y11_FrameStrobe_O[5] ,
    \Tile_X7Y11_FrameStrobe_O[4] ,
    \Tile_X7Y11_FrameStrobe_O[3] ,
    \Tile_X7Y11_FrameStrobe_O[2] ,
    \Tile_X7Y11_FrameStrobe_O[1] ,
    \Tile_X7Y11_FrameStrobe_O[0] }),
    .Tile_X0Y0_N1BEG({\Tile_X7Y11_N1BEG[3] ,
    \Tile_X7Y11_N1BEG[2] ,
    \Tile_X7Y11_N1BEG[1] ,
    \Tile_X7Y11_N1BEG[0] }),
    .Tile_X0Y0_N2BEG({\Tile_X7Y11_N2BEG[7] ,
    \Tile_X7Y11_N2BEG[6] ,
    \Tile_X7Y11_N2BEG[5] ,
    \Tile_X7Y11_N2BEG[4] ,
    \Tile_X7Y11_N2BEG[3] ,
    \Tile_X7Y11_N2BEG[2] ,
    \Tile_X7Y11_N2BEG[1] ,
    \Tile_X7Y11_N2BEG[0] }),
    .Tile_X0Y0_N2BEGb({\Tile_X7Y11_N2BEGb[7] ,
    \Tile_X7Y11_N2BEGb[6] ,
    \Tile_X7Y11_N2BEGb[5] ,
    \Tile_X7Y11_N2BEGb[4] ,
    \Tile_X7Y11_N2BEGb[3] ,
    \Tile_X7Y11_N2BEGb[2] ,
    \Tile_X7Y11_N2BEGb[1] ,
    \Tile_X7Y11_N2BEGb[0] }),
    .Tile_X0Y0_N4BEG({\Tile_X7Y11_N4BEG[15] ,
    \Tile_X7Y11_N4BEG[14] ,
    \Tile_X7Y11_N4BEG[13] ,
    \Tile_X7Y11_N4BEG[12] ,
    \Tile_X7Y11_N4BEG[11] ,
    \Tile_X7Y11_N4BEG[10] ,
    \Tile_X7Y11_N4BEG[9] ,
    \Tile_X7Y11_N4BEG[8] ,
    \Tile_X7Y11_N4BEG[7] ,
    \Tile_X7Y11_N4BEG[6] ,
    \Tile_X7Y11_N4BEG[5] ,
    \Tile_X7Y11_N4BEG[4] ,
    \Tile_X7Y11_N4BEG[3] ,
    \Tile_X7Y11_N4BEG[2] ,
    \Tile_X7Y11_N4BEG[1] ,
    \Tile_X7Y11_N4BEG[0] }),
    .Tile_X0Y0_NN4BEG({\Tile_X7Y11_NN4BEG[15] ,
    \Tile_X7Y11_NN4BEG[14] ,
    \Tile_X7Y11_NN4BEG[13] ,
    \Tile_X7Y11_NN4BEG[12] ,
    \Tile_X7Y11_NN4BEG[11] ,
    \Tile_X7Y11_NN4BEG[10] ,
    \Tile_X7Y11_NN4BEG[9] ,
    \Tile_X7Y11_NN4BEG[8] ,
    \Tile_X7Y11_NN4BEG[7] ,
    \Tile_X7Y11_NN4BEG[6] ,
    \Tile_X7Y11_NN4BEG[5] ,
    \Tile_X7Y11_NN4BEG[4] ,
    \Tile_X7Y11_NN4BEG[3] ,
    \Tile_X7Y11_NN4BEG[2] ,
    \Tile_X7Y11_NN4BEG[1] ,
    \Tile_X7Y11_NN4BEG[0] }),
    .Tile_X0Y0_S1END({\Tile_X7Y10_S1BEG[3] ,
    \Tile_X7Y10_S1BEG[2] ,
    \Tile_X7Y10_S1BEG[1] ,
    \Tile_X7Y10_S1BEG[0] }),
    .Tile_X0Y0_S2END({\Tile_X7Y10_S2BEGb[7] ,
    \Tile_X7Y10_S2BEGb[6] ,
    \Tile_X7Y10_S2BEGb[5] ,
    \Tile_X7Y10_S2BEGb[4] ,
    \Tile_X7Y10_S2BEGb[3] ,
    \Tile_X7Y10_S2BEGb[2] ,
    \Tile_X7Y10_S2BEGb[1] ,
    \Tile_X7Y10_S2BEGb[0] }),
    .Tile_X0Y0_S2MID({\Tile_X7Y10_S2BEG[7] ,
    \Tile_X7Y10_S2BEG[6] ,
    \Tile_X7Y10_S2BEG[5] ,
    \Tile_X7Y10_S2BEG[4] ,
    \Tile_X7Y10_S2BEG[3] ,
    \Tile_X7Y10_S2BEG[2] ,
    \Tile_X7Y10_S2BEG[1] ,
    \Tile_X7Y10_S2BEG[0] }),
    .Tile_X0Y0_S4END({\Tile_X7Y10_S4BEG[15] ,
    \Tile_X7Y10_S4BEG[14] ,
    \Tile_X7Y10_S4BEG[13] ,
    \Tile_X7Y10_S4BEG[12] ,
    \Tile_X7Y10_S4BEG[11] ,
    \Tile_X7Y10_S4BEG[10] ,
    \Tile_X7Y10_S4BEG[9] ,
    \Tile_X7Y10_S4BEG[8] ,
    \Tile_X7Y10_S4BEG[7] ,
    \Tile_X7Y10_S4BEG[6] ,
    \Tile_X7Y10_S4BEG[5] ,
    \Tile_X7Y10_S4BEG[4] ,
    \Tile_X7Y10_S4BEG[3] ,
    \Tile_X7Y10_S4BEG[2] ,
    \Tile_X7Y10_S4BEG[1] ,
    \Tile_X7Y10_S4BEG[0] }),
    .Tile_X0Y0_SS4END({\Tile_X7Y10_SS4BEG[15] ,
    \Tile_X7Y10_SS4BEG[14] ,
    \Tile_X7Y10_SS4BEG[13] ,
    \Tile_X7Y10_SS4BEG[12] ,
    \Tile_X7Y10_SS4BEG[11] ,
    \Tile_X7Y10_SS4BEG[10] ,
    \Tile_X7Y10_SS4BEG[9] ,
    \Tile_X7Y10_SS4BEG[8] ,
    \Tile_X7Y10_SS4BEG[7] ,
    \Tile_X7Y10_SS4BEG[6] ,
    \Tile_X7Y10_SS4BEG[5] ,
    \Tile_X7Y10_SS4BEG[4] ,
    \Tile_X7Y10_SS4BEG[3] ,
    \Tile_X7Y10_SS4BEG[2] ,
    \Tile_X7Y10_SS4BEG[1] ,
    \Tile_X7Y10_SS4BEG[0] }),
    .Tile_X0Y0_W1BEG({\Tile_X7Y11_W1BEG[3] ,
    \Tile_X7Y11_W1BEG[2] ,
    \Tile_X7Y11_W1BEG[1] ,
    \Tile_X7Y11_W1BEG[0] }),
    .Tile_X0Y0_W1END({\Tile_X8Y11_W1BEG[3] ,
    \Tile_X8Y11_W1BEG[2] ,
    \Tile_X8Y11_W1BEG[1] ,
    \Tile_X8Y11_W1BEG[0] }),
    .Tile_X0Y0_W2BEG({\Tile_X7Y11_W2BEG[7] ,
    \Tile_X7Y11_W2BEG[6] ,
    \Tile_X7Y11_W2BEG[5] ,
    \Tile_X7Y11_W2BEG[4] ,
    \Tile_X7Y11_W2BEG[3] ,
    \Tile_X7Y11_W2BEG[2] ,
    \Tile_X7Y11_W2BEG[1] ,
    \Tile_X7Y11_W2BEG[0] }),
    .Tile_X0Y0_W2BEGb({\Tile_X7Y11_W2BEGb[7] ,
    \Tile_X7Y11_W2BEGb[6] ,
    \Tile_X7Y11_W2BEGb[5] ,
    \Tile_X7Y11_W2BEGb[4] ,
    \Tile_X7Y11_W2BEGb[3] ,
    \Tile_X7Y11_W2BEGb[2] ,
    \Tile_X7Y11_W2BEGb[1] ,
    \Tile_X7Y11_W2BEGb[0] }),
    .Tile_X0Y0_W2END({\Tile_X8Y11_W2BEGb[7] ,
    \Tile_X8Y11_W2BEGb[6] ,
    \Tile_X8Y11_W2BEGb[5] ,
    \Tile_X8Y11_W2BEGb[4] ,
    \Tile_X8Y11_W2BEGb[3] ,
    \Tile_X8Y11_W2BEGb[2] ,
    \Tile_X8Y11_W2BEGb[1] ,
    \Tile_X8Y11_W2BEGb[0] }),
    .Tile_X0Y0_W2MID({\Tile_X8Y11_W2BEG[7] ,
    \Tile_X8Y11_W2BEG[6] ,
    \Tile_X8Y11_W2BEG[5] ,
    \Tile_X8Y11_W2BEG[4] ,
    \Tile_X8Y11_W2BEG[3] ,
    \Tile_X8Y11_W2BEG[2] ,
    \Tile_X8Y11_W2BEG[1] ,
    \Tile_X8Y11_W2BEG[0] }),
    .Tile_X0Y0_W6BEG({\Tile_X7Y11_W6BEG[11] ,
    \Tile_X7Y11_W6BEG[10] ,
    \Tile_X7Y11_W6BEG[9] ,
    \Tile_X7Y11_W6BEG[8] ,
    \Tile_X7Y11_W6BEG[7] ,
    \Tile_X7Y11_W6BEG[6] ,
    \Tile_X7Y11_W6BEG[5] ,
    \Tile_X7Y11_W6BEG[4] ,
    \Tile_X7Y11_W6BEG[3] ,
    \Tile_X7Y11_W6BEG[2] ,
    \Tile_X7Y11_W6BEG[1] ,
    \Tile_X7Y11_W6BEG[0] }),
    .Tile_X0Y0_W6END({\Tile_X8Y11_W6BEG[11] ,
    \Tile_X8Y11_W6BEG[10] ,
    \Tile_X8Y11_W6BEG[9] ,
    \Tile_X8Y11_W6BEG[8] ,
    \Tile_X8Y11_W6BEG[7] ,
    \Tile_X8Y11_W6BEG[6] ,
    \Tile_X8Y11_W6BEG[5] ,
    \Tile_X8Y11_W6BEG[4] ,
    \Tile_X8Y11_W6BEG[3] ,
    \Tile_X8Y11_W6BEG[2] ,
    \Tile_X8Y11_W6BEG[1] ,
    \Tile_X8Y11_W6BEG[0] }),
    .Tile_X0Y0_WW4BEG({\Tile_X7Y11_WW4BEG[15] ,
    \Tile_X7Y11_WW4BEG[14] ,
    \Tile_X7Y11_WW4BEG[13] ,
    \Tile_X7Y11_WW4BEG[12] ,
    \Tile_X7Y11_WW4BEG[11] ,
    \Tile_X7Y11_WW4BEG[10] ,
    \Tile_X7Y11_WW4BEG[9] ,
    \Tile_X7Y11_WW4BEG[8] ,
    \Tile_X7Y11_WW4BEG[7] ,
    \Tile_X7Y11_WW4BEG[6] ,
    \Tile_X7Y11_WW4BEG[5] ,
    \Tile_X7Y11_WW4BEG[4] ,
    \Tile_X7Y11_WW4BEG[3] ,
    \Tile_X7Y11_WW4BEG[2] ,
    \Tile_X7Y11_WW4BEG[1] ,
    \Tile_X7Y11_WW4BEG[0] }),
    .Tile_X0Y0_WW4END({\Tile_X8Y11_WW4BEG[15] ,
    \Tile_X8Y11_WW4BEG[14] ,
    \Tile_X8Y11_WW4BEG[13] ,
    \Tile_X8Y11_WW4BEG[12] ,
    \Tile_X8Y11_WW4BEG[11] ,
    \Tile_X8Y11_WW4BEG[10] ,
    \Tile_X8Y11_WW4BEG[9] ,
    \Tile_X8Y11_WW4BEG[8] ,
    \Tile_X8Y11_WW4BEG[7] ,
    \Tile_X8Y11_WW4BEG[6] ,
    \Tile_X8Y11_WW4BEG[5] ,
    \Tile_X8Y11_WW4BEG[4] ,
    \Tile_X8Y11_WW4BEG[3] ,
    \Tile_X8Y11_WW4BEG[2] ,
    \Tile_X8Y11_WW4BEG[1] ,
    \Tile_X8Y11_WW4BEG[0] }),
    .Tile_X0Y1_E1BEG({\Tile_X7Y12_E1BEG[3] ,
    \Tile_X7Y12_E1BEG[2] ,
    \Tile_X7Y12_E1BEG[1] ,
    \Tile_X7Y12_E1BEG[0] }),
    .Tile_X0Y1_E1END({\Tile_X6Y12_E1BEG[3] ,
    \Tile_X6Y12_E1BEG[2] ,
    \Tile_X6Y12_E1BEG[1] ,
    \Tile_X6Y12_E1BEG[0] }),
    .Tile_X0Y1_E2BEG({\Tile_X7Y12_E2BEG[7] ,
    \Tile_X7Y12_E2BEG[6] ,
    \Tile_X7Y12_E2BEG[5] ,
    \Tile_X7Y12_E2BEG[4] ,
    \Tile_X7Y12_E2BEG[3] ,
    \Tile_X7Y12_E2BEG[2] ,
    \Tile_X7Y12_E2BEG[1] ,
    \Tile_X7Y12_E2BEG[0] }),
    .Tile_X0Y1_E2BEGb({\Tile_X7Y12_E2BEGb[7] ,
    \Tile_X7Y12_E2BEGb[6] ,
    \Tile_X7Y12_E2BEGb[5] ,
    \Tile_X7Y12_E2BEGb[4] ,
    \Tile_X7Y12_E2BEGb[3] ,
    \Tile_X7Y12_E2BEGb[2] ,
    \Tile_X7Y12_E2BEGb[1] ,
    \Tile_X7Y12_E2BEGb[0] }),
    .Tile_X0Y1_E2END({\Tile_X6Y12_E2BEGb[7] ,
    \Tile_X6Y12_E2BEGb[6] ,
    \Tile_X6Y12_E2BEGb[5] ,
    \Tile_X6Y12_E2BEGb[4] ,
    \Tile_X6Y12_E2BEGb[3] ,
    \Tile_X6Y12_E2BEGb[2] ,
    \Tile_X6Y12_E2BEGb[1] ,
    \Tile_X6Y12_E2BEGb[0] }),
    .Tile_X0Y1_E2MID({\Tile_X6Y12_E2BEG[7] ,
    \Tile_X6Y12_E2BEG[6] ,
    \Tile_X6Y12_E2BEG[5] ,
    \Tile_X6Y12_E2BEG[4] ,
    \Tile_X6Y12_E2BEG[3] ,
    \Tile_X6Y12_E2BEG[2] ,
    \Tile_X6Y12_E2BEG[1] ,
    \Tile_X6Y12_E2BEG[0] }),
    .Tile_X0Y1_E6BEG({\Tile_X7Y12_E6BEG[11] ,
    \Tile_X7Y12_E6BEG[10] ,
    \Tile_X7Y12_E6BEG[9] ,
    \Tile_X7Y12_E6BEG[8] ,
    \Tile_X7Y12_E6BEG[7] ,
    \Tile_X7Y12_E6BEG[6] ,
    \Tile_X7Y12_E6BEG[5] ,
    \Tile_X7Y12_E6BEG[4] ,
    \Tile_X7Y12_E6BEG[3] ,
    \Tile_X7Y12_E6BEG[2] ,
    \Tile_X7Y12_E6BEG[1] ,
    \Tile_X7Y12_E6BEG[0] }),
    .Tile_X0Y1_E6END({\Tile_X6Y12_E6BEG[11] ,
    \Tile_X6Y12_E6BEG[10] ,
    \Tile_X6Y12_E6BEG[9] ,
    \Tile_X6Y12_E6BEG[8] ,
    \Tile_X6Y12_E6BEG[7] ,
    \Tile_X6Y12_E6BEG[6] ,
    \Tile_X6Y12_E6BEG[5] ,
    \Tile_X6Y12_E6BEG[4] ,
    \Tile_X6Y12_E6BEG[3] ,
    \Tile_X6Y12_E6BEG[2] ,
    \Tile_X6Y12_E6BEG[1] ,
    \Tile_X6Y12_E6BEG[0] }),
    .Tile_X0Y1_EE4BEG({\Tile_X7Y12_EE4BEG[15] ,
    \Tile_X7Y12_EE4BEG[14] ,
    \Tile_X7Y12_EE4BEG[13] ,
    \Tile_X7Y12_EE4BEG[12] ,
    \Tile_X7Y12_EE4BEG[11] ,
    \Tile_X7Y12_EE4BEG[10] ,
    \Tile_X7Y12_EE4BEG[9] ,
    \Tile_X7Y12_EE4BEG[8] ,
    \Tile_X7Y12_EE4BEG[7] ,
    \Tile_X7Y12_EE4BEG[6] ,
    \Tile_X7Y12_EE4BEG[5] ,
    \Tile_X7Y12_EE4BEG[4] ,
    \Tile_X7Y12_EE4BEG[3] ,
    \Tile_X7Y12_EE4BEG[2] ,
    \Tile_X7Y12_EE4BEG[1] ,
    \Tile_X7Y12_EE4BEG[0] }),
    .Tile_X0Y1_EE4END({\Tile_X6Y12_EE4BEG[15] ,
    \Tile_X6Y12_EE4BEG[14] ,
    \Tile_X6Y12_EE4BEG[13] ,
    \Tile_X6Y12_EE4BEG[12] ,
    \Tile_X6Y12_EE4BEG[11] ,
    \Tile_X6Y12_EE4BEG[10] ,
    \Tile_X6Y12_EE4BEG[9] ,
    \Tile_X6Y12_EE4BEG[8] ,
    \Tile_X6Y12_EE4BEG[7] ,
    \Tile_X6Y12_EE4BEG[6] ,
    \Tile_X6Y12_EE4BEG[5] ,
    \Tile_X6Y12_EE4BEG[4] ,
    \Tile_X6Y12_EE4BEG[3] ,
    \Tile_X6Y12_EE4BEG[2] ,
    \Tile_X6Y12_EE4BEG[1] ,
    \Tile_X6Y12_EE4BEG[0] }),
    .Tile_X0Y1_FrameData({\Tile_X6Y12_FrameData_O[31] ,
    \Tile_X6Y12_FrameData_O[30] ,
    \Tile_X6Y12_FrameData_O[29] ,
    \Tile_X6Y12_FrameData_O[28] ,
    \Tile_X6Y12_FrameData_O[27] ,
    \Tile_X6Y12_FrameData_O[26] ,
    \Tile_X6Y12_FrameData_O[25] ,
    \Tile_X6Y12_FrameData_O[24] ,
    \Tile_X6Y12_FrameData_O[23] ,
    \Tile_X6Y12_FrameData_O[22] ,
    \Tile_X6Y12_FrameData_O[21] ,
    \Tile_X6Y12_FrameData_O[20] ,
    \Tile_X6Y12_FrameData_O[19] ,
    \Tile_X6Y12_FrameData_O[18] ,
    \Tile_X6Y12_FrameData_O[17] ,
    \Tile_X6Y12_FrameData_O[16] ,
    \Tile_X6Y12_FrameData_O[15] ,
    \Tile_X6Y12_FrameData_O[14] ,
    \Tile_X6Y12_FrameData_O[13] ,
    \Tile_X6Y12_FrameData_O[12] ,
    \Tile_X6Y12_FrameData_O[11] ,
    \Tile_X6Y12_FrameData_O[10] ,
    \Tile_X6Y12_FrameData_O[9] ,
    \Tile_X6Y12_FrameData_O[8] ,
    \Tile_X6Y12_FrameData_O[7] ,
    \Tile_X6Y12_FrameData_O[6] ,
    \Tile_X6Y12_FrameData_O[5] ,
    \Tile_X6Y12_FrameData_O[4] ,
    \Tile_X6Y12_FrameData_O[3] ,
    \Tile_X6Y12_FrameData_O[2] ,
    \Tile_X6Y12_FrameData_O[1] ,
    \Tile_X6Y12_FrameData_O[0] }),
    .Tile_X0Y1_FrameData_O({\Tile_X7Y12_FrameData_O[31] ,
    \Tile_X7Y12_FrameData_O[30] ,
    \Tile_X7Y12_FrameData_O[29] ,
    \Tile_X7Y12_FrameData_O[28] ,
    \Tile_X7Y12_FrameData_O[27] ,
    \Tile_X7Y12_FrameData_O[26] ,
    \Tile_X7Y12_FrameData_O[25] ,
    \Tile_X7Y12_FrameData_O[24] ,
    \Tile_X7Y12_FrameData_O[23] ,
    \Tile_X7Y12_FrameData_O[22] ,
    \Tile_X7Y12_FrameData_O[21] ,
    \Tile_X7Y12_FrameData_O[20] ,
    \Tile_X7Y12_FrameData_O[19] ,
    \Tile_X7Y12_FrameData_O[18] ,
    \Tile_X7Y12_FrameData_O[17] ,
    \Tile_X7Y12_FrameData_O[16] ,
    \Tile_X7Y12_FrameData_O[15] ,
    \Tile_X7Y12_FrameData_O[14] ,
    \Tile_X7Y12_FrameData_O[13] ,
    \Tile_X7Y12_FrameData_O[12] ,
    \Tile_X7Y12_FrameData_O[11] ,
    \Tile_X7Y12_FrameData_O[10] ,
    \Tile_X7Y12_FrameData_O[9] ,
    \Tile_X7Y12_FrameData_O[8] ,
    \Tile_X7Y12_FrameData_O[7] ,
    \Tile_X7Y12_FrameData_O[6] ,
    \Tile_X7Y12_FrameData_O[5] ,
    \Tile_X7Y12_FrameData_O[4] ,
    \Tile_X7Y12_FrameData_O[3] ,
    \Tile_X7Y12_FrameData_O[2] ,
    \Tile_X7Y12_FrameData_O[1] ,
    \Tile_X7Y12_FrameData_O[0] }),
    .Tile_X0Y1_FrameStrobe({\Tile_X7Y13_FrameStrobe_O[19] ,
    \Tile_X7Y13_FrameStrobe_O[18] ,
    \Tile_X7Y13_FrameStrobe_O[17] ,
    \Tile_X7Y13_FrameStrobe_O[16] ,
    \Tile_X7Y13_FrameStrobe_O[15] ,
    \Tile_X7Y13_FrameStrobe_O[14] ,
    \Tile_X7Y13_FrameStrobe_O[13] ,
    \Tile_X7Y13_FrameStrobe_O[12] ,
    \Tile_X7Y13_FrameStrobe_O[11] ,
    \Tile_X7Y13_FrameStrobe_O[10] ,
    \Tile_X7Y13_FrameStrobe_O[9] ,
    \Tile_X7Y13_FrameStrobe_O[8] ,
    \Tile_X7Y13_FrameStrobe_O[7] ,
    \Tile_X7Y13_FrameStrobe_O[6] ,
    \Tile_X7Y13_FrameStrobe_O[5] ,
    \Tile_X7Y13_FrameStrobe_O[4] ,
    \Tile_X7Y13_FrameStrobe_O[3] ,
    \Tile_X7Y13_FrameStrobe_O[2] ,
    \Tile_X7Y13_FrameStrobe_O[1] ,
    \Tile_X7Y13_FrameStrobe_O[0] }),
    .Tile_X0Y1_N1END({\Tile_X7Y13_N1BEG[3] ,
    \Tile_X7Y13_N1BEG[2] ,
    \Tile_X7Y13_N1BEG[1] ,
    \Tile_X7Y13_N1BEG[0] }),
    .Tile_X0Y1_N2END({\Tile_X7Y13_N2BEGb[7] ,
    \Tile_X7Y13_N2BEGb[6] ,
    \Tile_X7Y13_N2BEGb[5] ,
    \Tile_X7Y13_N2BEGb[4] ,
    \Tile_X7Y13_N2BEGb[3] ,
    \Tile_X7Y13_N2BEGb[2] ,
    \Tile_X7Y13_N2BEGb[1] ,
    \Tile_X7Y13_N2BEGb[0] }),
    .Tile_X0Y1_N2MID({\Tile_X7Y13_N2BEG[7] ,
    \Tile_X7Y13_N2BEG[6] ,
    \Tile_X7Y13_N2BEG[5] ,
    \Tile_X7Y13_N2BEG[4] ,
    \Tile_X7Y13_N2BEG[3] ,
    \Tile_X7Y13_N2BEG[2] ,
    \Tile_X7Y13_N2BEG[1] ,
    \Tile_X7Y13_N2BEG[0] }),
    .Tile_X0Y1_N4END({\Tile_X7Y13_N4BEG[15] ,
    \Tile_X7Y13_N4BEG[14] ,
    \Tile_X7Y13_N4BEG[13] ,
    \Tile_X7Y13_N4BEG[12] ,
    \Tile_X7Y13_N4BEG[11] ,
    \Tile_X7Y13_N4BEG[10] ,
    \Tile_X7Y13_N4BEG[9] ,
    \Tile_X7Y13_N4BEG[8] ,
    \Tile_X7Y13_N4BEG[7] ,
    \Tile_X7Y13_N4BEG[6] ,
    \Tile_X7Y13_N4BEG[5] ,
    \Tile_X7Y13_N4BEG[4] ,
    \Tile_X7Y13_N4BEG[3] ,
    \Tile_X7Y13_N4BEG[2] ,
    \Tile_X7Y13_N4BEG[1] ,
    \Tile_X7Y13_N4BEG[0] }),
    .Tile_X0Y1_NN4END({\Tile_X7Y13_NN4BEG[15] ,
    \Tile_X7Y13_NN4BEG[14] ,
    \Tile_X7Y13_NN4BEG[13] ,
    \Tile_X7Y13_NN4BEG[12] ,
    \Tile_X7Y13_NN4BEG[11] ,
    \Tile_X7Y13_NN4BEG[10] ,
    \Tile_X7Y13_NN4BEG[9] ,
    \Tile_X7Y13_NN4BEG[8] ,
    \Tile_X7Y13_NN4BEG[7] ,
    \Tile_X7Y13_NN4BEG[6] ,
    \Tile_X7Y13_NN4BEG[5] ,
    \Tile_X7Y13_NN4BEG[4] ,
    \Tile_X7Y13_NN4BEG[3] ,
    \Tile_X7Y13_NN4BEG[2] ,
    \Tile_X7Y13_NN4BEG[1] ,
    \Tile_X7Y13_NN4BEG[0] }),
    .Tile_X0Y1_S1BEG({\Tile_X7Y12_S1BEG[3] ,
    \Tile_X7Y12_S1BEG[2] ,
    \Tile_X7Y12_S1BEG[1] ,
    \Tile_X7Y12_S1BEG[0] }),
    .Tile_X0Y1_S2BEG({\Tile_X7Y12_S2BEG[7] ,
    \Tile_X7Y12_S2BEG[6] ,
    \Tile_X7Y12_S2BEG[5] ,
    \Tile_X7Y12_S2BEG[4] ,
    \Tile_X7Y12_S2BEG[3] ,
    \Tile_X7Y12_S2BEG[2] ,
    \Tile_X7Y12_S2BEG[1] ,
    \Tile_X7Y12_S2BEG[0] }),
    .Tile_X0Y1_S2BEGb({\Tile_X7Y12_S2BEGb[7] ,
    \Tile_X7Y12_S2BEGb[6] ,
    \Tile_X7Y12_S2BEGb[5] ,
    \Tile_X7Y12_S2BEGb[4] ,
    \Tile_X7Y12_S2BEGb[3] ,
    \Tile_X7Y12_S2BEGb[2] ,
    \Tile_X7Y12_S2BEGb[1] ,
    \Tile_X7Y12_S2BEGb[0] }),
    .Tile_X0Y1_S4BEG({\Tile_X7Y12_S4BEG[15] ,
    \Tile_X7Y12_S4BEG[14] ,
    \Tile_X7Y12_S4BEG[13] ,
    \Tile_X7Y12_S4BEG[12] ,
    \Tile_X7Y12_S4BEG[11] ,
    \Tile_X7Y12_S4BEG[10] ,
    \Tile_X7Y12_S4BEG[9] ,
    \Tile_X7Y12_S4BEG[8] ,
    \Tile_X7Y12_S4BEG[7] ,
    \Tile_X7Y12_S4BEG[6] ,
    \Tile_X7Y12_S4BEG[5] ,
    \Tile_X7Y12_S4BEG[4] ,
    \Tile_X7Y12_S4BEG[3] ,
    \Tile_X7Y12_S4BEG[2] ,
    \Tile_X7Y12_S4BEG[1] ,
    \Tile_X7Y12_S4BEG[0] }),
    .Tile_X0Y1_SS4BEG({\Tile_X7Y12_SS4BEG[15] ,
    \Tile_X7Y12_SS4BEG[14] ,
    \Tile_X7Y12_SS4BEG[13] ,
    \Tile_X7Y12_SS4BEG[12] ,
    \Tile_X7Y12_SS4BEG[11] ,
    \Tile_X7Y12_SS4BEG[10] ,
    \Tile_X7Y12_SS4BEG[9] ,
    \Tile_X7Y12_SS4BEG[8] ,
    \Tile_X7Y12_SS4BEG[7] ,
    \Tile_X7Y12_SS4BEG[6] ,
    \Tile_X7Y12_SS4BEG[5] ,
    \Tile_X7Y12_SS4BEG[4] ,
    \Tile_X7Y12_SS4BEG[3] ,
    \Tile_X7Y12_SS4BEG[2] ,
    \Tile_X7Y12_SS4BEG[1] ,
    \Tile_X7Y12_SS4BEG[0] }),
    .Tile_X0Y1_W1BEG({\Tile_X7Y12_W1BEG[3] ,
    \Tile_X7Y12_W1BEG[2] ,
    \Tile_X7Y12_W1BEG[1] ,
    \Tile_X7Y12_W1BEG[0] }),
    .Tile_X0Y1_W1END({\Tile_X8Y12_W1BEG[3] ,
    \Tile_X8Y12_W1BEG[2] ,
    \Tile_X8Y12_W1BEG[1] ,
    \Tile_X8Y12_W1BEG[0] }),
    .Tile_X0Y1_W2BEG({\Tile_X7Y12_W2BEG[7] ,
    \Tile_X7Y12_W2BEG[6] ,
    \Tile_X7Y12_W2BEG[5] ,
    \Tile_X7Y12_W2BEG[4] ,
    \Tile_X7Y12_W2BEG[3] ,
    \Tile_X7Y12_W2BEG[2] ,
    \Tile_X7Y12_W2BEG[1] ,
    \Tile_X7Y12_W2BEG[0] }),
    .Tile_X0Y1_W2BEGb({\Tile_X7Y12_W2BEGb[7] ,
    \Tile_X7Y12_W2BEGb[6] ,
    \Tile_X7Y12_W2BEGb[5] ,
    \Tile_X7Y12_W2BEGb[4] ,
    \Tile_X7Y12_W2BEGb[3] ,
    \Tile_X7Y12_W2BEGb[2] ,
    \Tile_X7Y12_W2BEGb[1] ,
    \Tile_X7Y12_W2BEGb[0] }),
    .Tile_X0Y1_W2END({\Tile_X8Y12_W2BEGb[7] ,
    \Tile_X8Y12_W2BEGb[6] ,
    \Tile_X8Y12_W2BEGb[5] ,
    \Tile_X8Y12_W2BEGb[4] ,
    \Tile_X8Y12_W2BEGb[3] ,
    \Tile_X8Y12_W2BEGb[2] ,
    \Tile_X8Y12_W2BEGb[1] ,
    \Tile_X8Y12_W2BEGb[0] }),
    .Tile_X0Y1_W2MID({\Tile_X8Y12_W2BEG[7] ,
    \Tile_X8Y12_W2BEG[6] ,
    \Tile_X8Y12_W2BEG[5] ,
    \Tile_X8Y12_W2BEG[4] ,
    \Tile_X8Y12_W2BEG[3] ,
    \Tile_X8Y12_W2BEG[2] ,
    \Tile_X8Y12_W2BEG[1] ,
    \Tile_X8Y12_W2BEG[0] }),
    .Tile_X0Y1_W6BEG({\Tile_X7Y12_W6BEG[11] ,
    \Tile_X7Y12_W6BEG[10] ,
    \Tile_X7Y12_W6BEG[9] ,
    \Tile_X7Y12_W6BEG[8] ,
    \Tile_X7Y12_W6BEG[7] ,
    \Tile_X7Y12_W6BEG[6] ,
    \Tile_X7Y12_W6BEG[5] ,
    \Tile_X7Y12_W6BEG[4] ,
    \Tile_X7Y12_W6BEG[3] ,
    \Tile_X7Y12_W6BEG[2] ,
    \Tile_X7Y12_W6BEG[1] ,
    \Tile_X7Y12_W6BEG[0] }),
    .Tile_X0Y1_W6END({\Tile_X8Y12_W6BEG[11] ,
    \Tile_X8Y12_W6BEG[10] ,
    \Tile_X8Y12_W6BEG[9] ,
    \Tile_X8Y12_W6BEG[8] ,
    \Tile_X8Y12_W6BEG[7] ,
    \Tile_X8Y12_W6BEG[6] ,
    \Tile_X8Y12_W6BEG[5] ,
    \Tile_X8Y12_W6BEG[4] ,
    \Tile_X8Y12_W6BEG[3] ,
    \Tile_X8Y12_W6BEG[2] ,
    \Tile_X8Y12_W6BEG[1] ,
    \Tile_X8Y12_W6BEG[0] }),
    .Tile_X0Y1_WW4BEG({\Tile_X7Y12_WW4BEG[15] ,
    \Tile_X7Y12_WW4BEG[14] ,
    \Tile_X7Y12_WW4BEG[13] ,
    \Tile_X7Y12_WW4BEG[12] ,
    \Tile_X7Y12_WW4BEG[11] ,
    \Tile_X7Y12_WW4BEG[10] ,
    \Tile_X7Y12_WW4BEG[9] ,
    \Tile_X7Y12_WW4BEG[8] ,
    \Tile_X7Y12_WW4BEG[7] ,
    \Tile_X7Y12_WW4BEG[6] ,
    \Tile_X7Y12_WW4BEG[5] ,
    \Tile_X7Y12_WW4BEG[4] ,
    \Tile_X7Y12_WW4BEG[3] ,
    \Tile_X7Y12_WW4BEG[2] ,
    \Tile_X7Y12_WW4BEG[1] ,
    \Tile_X7Y12_WW4BEG[0] }),
    .Tile_X0Y1_WW4END({\Tile_X8Y12_WW4BEG[15] ,
    \Tile_X8Y12_WW4BEG[14] ,
    \Tile_X8Y12_WW4BEG[13] ,
    \Tile_X8Y12_WW4BEG[12] ,
    \Tile_X8Y12_WW4BEG[11] ,
    \Tile_X8Y12_WW4BEG[10] ,
    \Tile_X8Y12_WW4BEG[9] ,
    \Tile_X8Y12_WW4BEG[8] ,
    \Tile_X8Y12_WW4BEG[7] ,
    \Tile_X8Y12_WW4BEG[6] ,
    \Tile_X8Y12_WW4BEG[5] ,
    \Tile_X8Y12_WW4BEG[4] ,
    \Tile_X8Y12_WW4BEG[3] ,
    \Tile_X8Y12_WW4BEG[2] ,
    \Tile_X8Y12_WW4BEG[1] ,
    \Tile_X8Y12_WW4BEG[0] }));
 DSP Tile_X7Y13_DSP (.Tile_X0Y0_UserCLKo(Tile_X7Y13_UserCLKo),
    .Tile_X0Y1_UserCLK(Tile_X7Y15_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .Tile_X0Y0_E1BEG({\Tile_X7Y13_E1BEG[3] ,
    \Tile_X7Y13_E1BEG[2] ,
    \Tile_X7Y13_E1BEG[1] ,
    \Tile_X7Y13_E1BEG[0] }),
    .Tile_X0Y0_E1END({\Tile_X6Y13_E1BEG[3] ,
    \Tile_X6Y13_E1BEG[2] ,
    \Tile_X6Y13_E1BEG[1] ,
    \Tile_X6Y13_E1BEG[0] }),
    .Tile_X0Y0_E2BEG({\Tile_X7Y13_E2BEG[7] ,
    \Tile_X7Y13_E2BEG[6] ,
    \Tile_X7Y13_E2BEG[5] ,
    \Tile_X7Y13_E2BEG[4] ,
    \Tile_X7Y13_E2BEG[3] ,
    \Tile_X7Y13_E2BEG[2] ,
    \Tile_X7Y13_E2BEG[1] ,
    \Tile_X7Y13_E2BEG[0] }),
    .Tile_X0Y0_E2BEGb({\Tile_X7Y13_E2BEGb[7] ,
    \Tile_X7Y13_E2BEGb[6] ,
    \Tile_X7Y13_E2BEGb[5] ,
    \Tile_X7Y13_E2BEGb[4] ,
    \Tile_X7Y13_E2BEGb[3] ,
    \Tile_X7Y13_E2BEGb[2] ,
    \Tile_X7Y13_E2BEGb[1] ,
    \Tile_X7Y13_E2BEGb[0] }),
    .Tile_X0Y0_E2END({\Tile_X6Y13_E2BEGb[7] ,
    \Tile_X6Y13_E2BEGb[6] ,
    \Tile_X6Y13_E2BEGb[5] ,
    \Tile_X6Y13_E2BEGb[4] ,
    \Tile_X6Y13_E2BEGb[3] ,
    \Tile_X6Y13_E2BEGb[2] ,
    \Tile_X6Y13_E2BEGb[1] ,
    \Tile_X6Y13_E2BEGb[0] }),
    .Tile_X0Y0_E2MID({\Tile_X6Y13_E2BEG[7] ,
    \Tile_X6Y13_E2BEG[6] ,
    \Tile_X6Y13_E2BEG[5] ,
    \Tile_X6Y13_E2BEG[4] ,
    \Tile_X6Y13_E2BEG[3] ,
    \Tile_X6Y13_E2BEG[2] ,
    \Tile_X6Y13_E2BEG[1] ,
    \Tile_X6Y13_E2BEG[0] }),
    .Tile_X0Y0_E6BEG({\Tile_X7Y13_E6BEG[11] ,
    \Tile_X7Y13_E6BEG[10] ,
    \Tile_X7Y13_E6BEG[9] ,
    \Tile_X7Y13_E6BEG[8] ,
    \Tile_X7Y13_E6BEG[7] ,
    \Tile_X7Y13_E6BEG[6] ,
    \Tile_X7Y13_E6BEG[5] ,
    \Tile_X7Y13_E6BEG[4] ,
    \Tile_X7Y13_E6BEG[3] ,
    \Tile_X7Y13_E6BEG[2] ,
    \Tile_X7Y13_E6BEG[1] ,
    \Tile_X7Y13_E6BEG[0] }),
    .Tile_X0Y0_E6END({\Tile_X6Y13_E6BEG[11] ,
    \Tile_X6Y13_E6BEG[10] ,
    \Tile_X6Y13_E6BEG[9] ,
    \Tile_X6Y13_E6BEG[8] ,
    \Tile_X6Y13_E6BEG[7] ,
    \Tile_X6Y13_E6BEG[6] ,
    \Tile_X6Y13_E6BEG[5] ,
    \Tile_X6Y13_E6BEG[4] ,
    \Tile_X6Y13_E6BEG[3] ,
    \Tile_X6Y13_E6BEG[2] ,
    \Tile_X6Y13_E6BEG[1] ,
    \Tile_X6Y13_E6BEG[0] }),
    .Tile_X0Y0_EE4BEG({\Tile_X7Y13_EE4BEG[15] ,
    \Tile_X7Y13_EE4BEG[14] ,
    \Tile_X7Y13_EE4BEG[13] ,
    \Tile_X7Y13_EE4BEG[12] ,
    \Tile_X7Y13_EE4BEG[11] ,
    \Tile_X7Y13_EE4BEG[10] ,
    \Tile_X7Y13_EE4BEG[9] ,
    \Tile_X7Y13_EE4BEG[8] ,
    \Tile_X7Y13_EE4BEG[7] ,
    \Tile_X7Y13_EE4BEG[6] ,
    \Tile_X7Y13_EE4BEG[5] ,
    \Tile_X7Y13_EE4BEG[4] ,
    \Tile_X7Y13_EE4BEG[3] ,
    \Tile_X7Y13_EE4BEG[2] ,
    \Tile_X7Y13_EE4BEG[1] ,
    \Tile_X7Y13_EE4BEG[0] }),
    .Tile_X0Y0_EE4END({\Tile_X6Y13_EE4BEG[15] ,
    \Tile_X6Y13_EE4BEG[14] ,
    \Tile_X6Y13_EE4BEG[13] ,
    \Tile_X6Y13_EE4BEG[12] ,
    \Tile_X6Y13_EE4BEG[11] ,
    \Tile_X6Y13_EE4BEG[10] ,
    \Tile_X6Y13_EE4BEG[9] ,
    \Tile_X6Y13_EE4BEG[8] ,
    \Tile_X6Y13_EE4BEG[7] ,
    \Tile_X6Y13_EE4BEG[6] ,
    \Tile_X6Y13_EE4BEG[5] ,
    \Tile_X6Y13_EE4BEG[4] ,
    \Tile_X6Y13_EE4BEG[3] ,
    \Tile_X6Y13_EE4BEG[2] ,
    \Tile_X6Y13_EE4BEG[1] ,
    \Tile_X6Y13_EE4BEG[0] }),
    .Tile_X0Y0_FrameData({\Tile_X6Y13_FrameData_O[31] ,
    \Tile_X6Y13_FrameData_O[30] ,
    \Tile_X6Y13_FrameData_O[29] ,
    \Tile_X6Y13_FrameData_O[28] ,
    \Tile_X6Y13_FrameData_O[27] ,
    \Tile_X6Y13_FrameData_O[26] ,
    \Tile_X6Y13_FrameData_O[25] ,
    \Tile_X6Y13_FrameData_O[24] ,
    \Tile_X6Y13_FrameData_O[23] ,
    \Tile_X6Y13_FrameData_O[22] ,
    \Tile_X6Y13_FrameData_O[21] ,
    \Tile_X6Y13_FrameData_O[20] ,
    \Tile_X6Y13_FrameData_O[19] ,
    \Tile_X6Y13_FrameData_O[18] ,
    \Tile_X6Y13_FrameData_O[17] ,
    \Tile_X6Y13_FrameData_O[16] ,
    \Tile_X6Y13_FrameData_O[15] ,
    \Tile_X6Y13_FrameData_O[14] ,
    \Tile_X6Y13_FrameData_O[13] ,
    \Tile_X6Y13_FrameData_O[12] ,
    \Tile_X6Y13_FrameData_O[11] ,
    \Tile_X6Y13_FrameData_O[10] ,
    \Tile_X6Y13_FrameData_O[9] ,
    \Tile_X6Y13_FrameData_O[8] ,
    \Tile_X6Y13_FrameData_O[7] ,
    \Tile_X6Y13_FrameData_O[6] ,
    \Tile_X6Y13_FrameData_O[5] ,
    \Tile_X6Y13_FrameData_O[4] ,
    \Tile_X6Y13_FrameData_O[3] ,
    \Tile_X6Y13_FrameData_O[2] ,
    \Tile_X6Y13_FrameData_O[1] ,
    \Tile_X6Y13_FrameData_O[0] }),
    .Tile_X0Y0_FrameData_O({\Tile_X7Y13_FrameData_O[31] ,
    \Tile_X7Y13_FrameData_O[30] ,
    \Tile_X7Y13_FrameData_O[29] ,
    \Tile_X7Y13_FrameData_O[28] ,
    \Tile_X7Y13_FrameData_O[27] ,
    \Tile_X7Y13_FrameData_O[26] ,
    \Tile_X7Y13_FrameData_O[25] ,
    \Tile_X7Y13_FrameData_O[24] ,
    \Tile_X7Y13_FrameData_O[23] ,
    \Tile_X7Y13_FrameData_O[22] ,
    \Tile_X7Y13_FrameData_O[21] ,
    \Tile_X7Y13_FrameData_O[20] ,
    \Tile_X7Y13_FrameData_O[19] ,
    \Tile_X7Y13_FrameData_O[18] ,
    \Tile_X7Y13_FrameData_O[17] ,
    \Tile_X7Y13_FrameData_O[16] ,
    \Tile_X7Y13_FrameData_O[15] ,
    \Tile_X7Y13_FrameData_O[14] ,
    \Tile_X7Y13_FrameData_O[13] ,
    \Tile_X7Y13_FrameData_O[12] ,
    \Tile_X7Y13_FrameData_O[11] ,
    \Tile_X7Y13_FrameData_O[10] ,
    \Tile_X7Y13_FrameData_O[9] ,
    \Tile_X7Y13_FrameData_O[8] ,
    \Tile_X7Y13_FrameData_O[7] ,
    \Tile_X7Y13_FrameData_O[6] ,
    \Tile_X7Y13_FrameData_O[5] ,
    \Tile_X7Y13_FrameData_O[4] ,
    \Tile_X7Y13_FrameData_O[3] ,
    \Tile_X7Y13_FrameData_O[2] ,
    \Tile_X7Y13_FrameData_O[1] ,
    \Tile_X7Y13_FrameData_O[0] }),
    .Tile_X0Y0_FrameStrobe_O({\Tile_X7Y13_FrameStrobe_O[19] ,
    \Tile_X7Y13_FrameStrobe_O[18] ,
    \Tile_X7Y13_FrameStrobe_O[17] ,
    \Tile_X7Y13_FrameStrobe_O[16] ,
    \Tile_X7Y13_FrameStrobe_O[15] ,
    \Tile_X7Y13_FrameStrobe_O[14] ,
    \Tile_X7Y13_FrameStrobe_O[13] ,
    \Tile_X7Y13_FrameStrobe_O[12] ,
    \Tile_X7Y13_FrameStrobe_O[11] ,
    \Tile_X7Y13_FrameStrobe_O[10] ,
    \Tile_X7Y13_FrameStrobe_O[9] ,
    \Tile_X7Y13_FrameStrobe_O[8] ,
    \Tile_X7Y13_FrameStrobe_O[7] ,
    \Tile_X7Y13_FrameStrobe_O[6] ,
    \Tile_X7Y13_FrameStrobe_O[5] ,
    \Tile_X7Y13_FrameStrobe_O[4] ,
    \Tile_X7Y13_FrameStrobe_O[3] ,
    \Tile_X7Y13_FrameStrobe_O[2] ,
    \Tile_X7Y13_FrameStrobe_O[1] ,
    \Tile_X7Y13_FrameStrobe_O[0] }),
    .Tile_X0Y0_N1BEG({\Tile_X7Y13_N1BEG[3] ,
    \Tile_X7Y13_N1BEG[2] ,
    \Tile_X7Y13_N1BEG[1] ,
    \Tile_X7Y13_N1BEG[0] }),
    .Tile_X0Y0_N2BEG({\Tile_X7Y13_N2BEG[7] ,
    \Tile_X7Y13_N2BEG[6] ,
    \Tile_X7Y13_N2BEG[5] ,
    \Tile_X7Y13_N2BEG[4] ,
    \Tile_X7Y13_N2BEG[3] ,
    \Tile_X7Y13_N2BEG[2] ,
    \Tile_X7Y13_N2BEG[1] ,
    \Tile_X7Y13_N2BEG[0] }),
    .Tile_X0Y0_N2BEGb({\Tile_X7Y13_N2BEGb[7] ,
    \Tile_X7Y13_N2BEGb[6] ,
    \Tile_X7Y13_N2BEGb[5] ,
    \Tile_X7Y13_N2BEGb[4] ,
    \Tile_X7Y13_N2BEGb[3] ,
    \Tile_X7Y13_N2BEGb[2] ,
    \Tile_X7Y13_N2BEGb[1] ,
    \Tile_X7Y13_N2BEGb[0] }),
    .Tile_X0Y0_N4BEG({\Tile_X7Y13_N4BEG[15] ,
    \Tile_X7Y13_N4BEG[14] ,
    \Tile_X7Y13_N4BEG[13] ,
    \Tile_X7Y13_N4BEG[12] ,
    \Tile_X7Y13_N4BEG[11] ,
    \Tile_X7Y13_N4BEG[10] ,
    \Tile_X7Y13_N4BEG[9] ,
    \Tile_X7Y13_N4BEG[8] ,
    \Tile_X7Y13_N4BEG[7] ,
    \Tile_X7Y13_N4BEG[6] ,
    \Tile_X7Y13_N4BEG[5] ,
    \Tile_X7Y13_N4BEG[4] ,
    \Tile_X7Y13_N4BEG[3] ,
    \Tile_X7Y13_N4BEG[2] ,
    \Tile_X7Y13_N4BEG[1] ,
    \Tile_X7Y13_N4BEG[0] }),
    .Tile_X0Y0_NN4BEG({\Tile_X7Y13_NN4BEG[15] ,
    \Tile_X7Y13_NN4BEG[14] ,
    \Tile_X7Y13_NN4BEG[13] ,
    \Tile_X7Y13_NN4BEG[12] ,
    \Tile_X7Y13_NN4BEG[11] ,
    \Tile_X7Y13_NN4BEG[10] ,
    \Tile_X7Y13_NN4BEG[9] ,
    \Tile_X7Y13_NN4BEG[8] ,
    \Tile_X7Y13_NN4BEG[7] ,
    \Tile_X7Y13_NN4BEG[6] ,
    \Tile_X7Y13_NN4BEG[5] ,
    \Tile_X7Y13_NN4BEG[4] ,
    \Tile_X7Y13_NN4BEG[3] ,
    \Tile_X7Y13_NN4BEG[2] ,
    \Tile_X7Y13_NN4BEG[1] ,
    \Tile_X7Y13_NN4BEG[0] }),
    .Tile_X0Y0_S1END({\Tile_X7Y12_S1BEG[3] ,
    \Tile_X7Y12_S1BEG[2] ,
    \Tile_X7Y12_S1BEG[1] ,
    \Tile_X7Y12_S1BEG[0] }),
    .Tile_X0Y0_S2END({\Tile_X7Y12_S2BEGb[7] ,
    \Tile_X7Y12_S2BEGb[6] ,
    \Tile_X7Y12_S2BEGb[5] ,
    \Tile_X7Y12_S2BEGb[4] ,
    \Tile_X7Y12_S2BEGb[3] ,
    \Tile_X7Y12_S2BEGb[2] ,
    \Tile_X7Y12_S2BEGb[1] ,
    \Tile_X7Y12_S2BEGb[0] }),
    .Tile_X0Y0_S2MID({\Tile_X7Y12_S2BEG[7] ,
    \Tile_X7Y12_S2BEG[6] ,
    \Tile_X7Y12_S2BEG[5] ,
    \Tile_X7Y12_S2BEG[4] ,
    \Tile_X7Y12_S2BEG[3] ,
    \Tile_X7Y12_S2BEG[2] ,
    \Tile_X7Y12_S2BEG[1] ,
    \Tile_X7Y12_S2BEG[0] }),
    .Tile_X0Y0_S4END({\Tile_X7Y12_S4BEG[15] ,
    \Tile_X7Y12_S4BEG[14] ,
    \Tile_X7Y12_S4BEG[13] ,
    \Tile_X7Y12_S4BEG[12] ,
    \Tile_X7Y12_S4BEG[11] ,
    \Tile_X7Y12_S4BEG[10] ,
    \Tile_X7Y12_S4BEG[9] ,
    \Tile_X7Y12_S4BEG[8] ,
    \Tile_X7Y12_S4BEG[7] ,
    \Tile_X7Y12_S4BEG[6] ,
    \Tile_X7Y12_S4BEG[5] ,
    \Tile_X7Y12_S4BEG[4] ,
    \Tile_X7Y12_S4BEG[3] ,
    \Tile_X7Y12_S4BEG[2] ,
    \Tile_X7Y12_S4BEG[1] ,
    \Tile_X7Y12_S4BEG[0] }),
    .Tile_X0Y0_SS4END({\Tile_X7Y12_SS4BEG[15] ,
    \Tile_X7Y12_SS4BEG[14] ,
    \Tile_X7Y12_SS4BEG[13] ,
    \Tile_X7Y12_SS4BEG[12] ,
    \Tile_X7Y12_SS4BEG[11] ,
    \Tile_X7Y12_SS4BEG[10] ,
    \Tile_X7Y12_SS4BEG[9] ,
    \Tile_X7Y12_SS4BEG[8] ,
    \Tile_X7Y12_SS4BEG[7] ,
    \Tile_X7Y12_SS4BEG[6] ,
    \Tile_X7Y12_SS4BEG[5] ,
    \Tile_X7Y12_SS4BEG[4] ,
    \Tile_X7Y12_SS4BEG[3] ,
    \Tile_X7Y12_SS4BEG[2] ,
    \Tile_X7Y12_SS4BEG[1] ,
    \Tile_X7Y12_SS4BEG[0] }),
    .Tile_X0Y0_W1BEG({\Tile_X7Y13_W1BEG[3] ,
    \Tile_X7Y13_W1BEG[2] ,
    \Tile_X7Y13_W1BEG[1] ,
    \Tile_X7Y13_W1BEG[0] }),
    .Tile_X0Y0_W1END({\Tile_X8Y13_W1BEG[3] ,
    \Tile_X8Y13_W1BEG[2] ,
    \Tile_X8Y13_W1BEG[1] ,
    \Tile_X8Y13_W1BEG[0] }),
    .Tile_X0Y0_W2BEG({\Tile_X7Y13_W2BEG[7] ,
    \Tile_X7Y13_W2BEG[6] ,
    \Tile_X7Y13_W2BEG[5] ,
    \Tile_X7Y13_W2BEG[4] ,
    \Tile_X7Y13_W2BEG[3] ,
    \Tile_X7Y13_W2BEG[2] ,
    \Tile_X7Y13_W2BEG[1] ,
    \Tile_X7Y13_W2BEG[0] }),
    .Tile_X0Y0_W2BEGb({\Tile_X7Y13_W2BEGb[7] ,
    \Tile_X7Y13_W2BEGb[6] ,
    \Tile_X7Y13_W2BEGb[5] ,
    \Tile_X7Y13_W2BEGb[4] ,
    \Tile_X7Y13_W2BEGb[3] ,
    \Tile_X7Y13_W2BEGb[2] ,
    \Tile_X7Y13_W2BEGb[1] ,
    \Tile_X7Y13_W2BEGb[0] }),
    .Tile_X0Y0_W2END({\Tile_X8Y13_W2BEGb[7] ,
    \Tile_X8Y13_W2BEGb[6] ,
    \Tile_X8Y13_W2BEGb[5] ,
    \Tile_X8Y13_W2BEGb[4] ,
    \Tile_X8Y13_W2BEGb[3] ,
    \Tile_X8Y13_W2BEGb[2] ,
    \Tile_X8Y13_W2BEGb[1] ,
    \Tile_X8Y13_W2BEGb[0] }),
    .Tile_X0Y0_W2MID({\Tile_X8Y13_W2BEG[7] ,
    \Tile_X8Y13_W2BEG[6] ,
    \Tile_X8Y13_W2BEG[5] ,
    \Tile_X8Y13_W2BEG[4] ,
    \Tile_X8Y13_W2BEG[3] ,
    \Tile_X8Y13_W2BEG[2] ,
    \Tile_X8Y13_W2BEG[1] ,
    \Tile_X8Y13_W2BEG[0] }),
    .Tile_X0Y0_W6BEG({\Tile_X7Y13_W6BEG[11] ,
    \Tile_X7Y13_W6BEG[10] ,
    \Tile_X7Y13_W6BEG[9] ,
    \Tile_X7Y13_W6BEG[8] ,
    \Tile_X7Y13_W6BEG[7] ,
    \Tile_X7Y13_W6BEG[6] ,
    \Tile_X7Y13_W6BEG[5] ,
    \Tile_X7Y13_W6BEG[4] ,
    \Tile_X7Y13_W6BEG[3] ,
    \Tile_X7Y13_W6BEG[2] ,
    \Tile_X7Y13_W6BEG[1] ,
    \Tile_X7Y13_W6BEG[0] }),
    .Tile_X0Y0_W6END({\Tile_X8Y13_W6BEG[11] ,
    \Tile_X8Y13_W6BEG[10] ,
    \Tile_X8Y13_W6BEG[9] ,
    \Tile_X8Y13_W6BEG[8] ,
    \Tile_X8Y13_W6BEG[7] ,
    \Tile_X8Y13_W6BEG[6] ,
    \Tile_X8Y13_W6BEG[5] ,
    \Tile_X8Y13_W6BEG[4] ,
    \Tile_X8Y13_W6BEG[3] ,
    \Tile_X8Y13_W6BEG[2] ,
    \Tile_X8Y13_W6BEG[1] ,
    \Tile_X8Y13_W6BEG[0] }),
    .Tile_X0Y0_WW4BEG({\Tile_X7Y13_WW4BEG[15] ,
    \Tile_X7Y13_WW4BEG[14] ,
    \Tile_X7Y13_WW4BEG[13] ,
    \Tile_X7Y13_WW4BEG[12] ,
    \Tile_X7Y13_WW4BEG[11] ,
    \Tile_X7Y13_WW4BEG[10] ,
    \Tile_X7Y13_WW4BEG[9] ,
    \Tile_X7Y13_WW4BEG[8] ,
    \Tile_X7Y13_WW4BEG[7] ,
    \Tile_X7Y13_WW4BEG[6] ,
    \Tile_X7Y13_WW4BEG[5] ,
    \Tile_X7Y13_WW4BEG[4] ,
    \Tile_X7Y13_WW4BEG[3] ,
    \Tile_X7Y13_WW4BEG[2] ,
    \Tile_X7Y13_WW4BEG[1] ,
    \Tile_X7Y13_WW4BEG[0] }),
    .Tile_X0Y0_WW4END({\Tile_X8Y13_WW4BEG[15] ,
    \Tile_X8Y13_WW4BEG[14] ,
    \Tile_X8Y13_WW4BEG[13] ,
    \Tile_X8Y13_WW4BEG[12] ,
    \Tile_X8Y13_WW4BEG[11] ,
    \Tile_X8Y13_WW4BEG[10] ,
    \Tile_X8Y13_WW4BEG[9] ,
    \Tile_X8Y13_WW4BEG[8] ,
    \Tile_X8Y13_WW4BEG[7] ,
    \Tile_X8Y13_WW4BEG[6] ,
    \Tile_X8Y13_WW4BEG[5] ,
    \Tile_X8Y13_WW4BEG[4] ,
    \Tile_X8Y13_WW4BEG[3] ,
    \Tile_X8Y13_WW4BEG[2] ,
    \Tile_X8Y13_WW4BEG[1] ,
    \Tile_X8Y13_WW4BEG[0] }),
    .Tile_X0Y1_E1BEG({\Tile_X7Y14_E1BEG[3] ,
    \Tile_X7Y14_E1BEG[2] ,
    \Tile_X7Y14_E1BEG[1] ,
    \Tile_X7Y14_E1BEG[0] }),
    .Tile_X0Y1_E1END({\Tile_X6Y14_E1BEG[3] ,
    \Tile_X6Y14_E1BEG[2] ,
    \Tile_X6Y14_E1BEG[1] ,
    \Tile_X6Y14_E1BEG[0] }),
    .Tile_X0Y1_E2BEG({\Tile_X7Y14_E2BEG[7] ,
    \Tile_X7Y14_E2BEG[6] ,
    \Tile_X7Y14_E2BEG[5] ,
    \Tile_X7Y14_E2BEG[4] ,
    \Tile_X7Y14_E2BEG[3] ,
    \Tile_X7Y14_E2BEG[2] ,
    \Tile_X7Y14_E2BEG[1] ,
    \Tile_X7Y14_E2BEG[0] }),
    .Tile_X0Y1_E2BEGb({\Tile_X7Y14_E2BEGb[7] ,
    \Tile_X7Y14_E2BEGb[6] ,
    \Tile_X7Y14_E2BEGb[5] ,
    \Tile_X7Y14_E2BEGb[4] ,
    \Tile_X7Y14_E2BEGb[3] ,
    \Tile_X7Y14_E2BEGb[2] ,
    \Tile_X7Y14_E2BEGb[1] ,
    \Tile_X7Y14_E2BEGb[0] }),
    .Tile_X0Y1_E2END({\Tile_X6Y14_E2BEGb[7] ,
    \Tile_X6Y14_E2BEGb[6] ,
    \Tile_X6Y14_E2BEGb[5] ,
    \Tile_X6Y14_E2BEGb[4] ,
    \Tile_X6Y14_E2BEGb[3] ,
    \Tile_X6Y14_E2BEGb[2] ,
    \Tile_X6Y14_E2BEGb[1] ,
    \Tile_X6Y14_E2BEGb[0] }),
    .Tile_X0Y1_E2MID({\Tile_X6Y14_E2BEG[7] ,
    \Tile_X6Y14_E2BEG[6] ,
    \Tile_X6Y14_E2BEG[5] ,
    \Tile_X6Y14_E2BEG[4] ,
    \Tile_X6Y14_E2BEG[3] ,
    \Tile_X6Y14_E2BEG[2] ,
    \Tile_X6Y14_E2BEG[1] ,
    \Tile_X6Y14_E2BEG[0] }),
    .Tile_X0Y1_E6BEG({\Tile_X7Y14_E6BEG[11] ,
    \Tile_X7Y14_E6BEG[10] ,
    \Tile_X7Y14_E6BEG[9] ,
    \Tile_X7Y14_E6BEG[8] ,
    \Tile_X7Y14_E6BEG[7] ,
    \Tile_X7Y14_E6BEG[6] ,
    \Tile_X7Y14_E6BEG[5] ,
    \Tile_X7Y14_E6BEG[4] ,
    \Tile_X7Y14_E6BEG[3] ,
    \Tile_X7Y14_E6BEG[2] ,
    \Tile_X7Y14_E6BEG[1] ,
    \Tile_X7Y14_E6BEG[0] }),
    .Tile_X0Y1_E6END({\Tile_X6Y14_E6BEG[11] ,
    \Tile_X6Y14_E6BEG[10] ,
    \Tile_X6Y14_E6BEG[9] ,
    \Tile_X6Y14_E6BEG[8] ,
    \Tile_X6Y14_E6BEG[7] ,
    \Tile_X6Y14_E6BEG[6] ,
    \Tile_X6Y14_E6BEG[5] ,
    \Tile_X6Y14_E6BEG[4] ,
    \Tile_X6Y14_E6BEG[3] ,
    \Tile_X6Y14_E6BEG[2] ,
    \Tile_X6Y14_E6BEG[1] ,
    \Tile_X6Y14_E6BEG[0] }),
    .Tile_X0Y1_EE4BEG({\Tile_X7Y14_EE4BEG[15] ,
    \Tile_X7Y14_EE4BEG[14] ,
    \Tile_X7Y14_EE4BEG[13] ,
    \Tile_X7Y14_EE4BEG[12] ,
    \Tile_X7Y14_EE4BEG[11] ,
    \Tile_X7Y14_EE4BEG[10] ,
    \Tile_X7Y14_EE4BEG[9] ,
    \Tile_X7Y14_EE4BEG[8] ,
    \Tile_X7Y14_EE4BEG[7] ,
    \Tile_X7Y14_EE4BEG[6] ,
    \Tile_X7Y14_EE4BEG[5] ,
    \Tile_X7Y14_EE4BEG[4] ,
    \Tile_X7Y14_EE4BEG[3] ,
    \Tile_X7Y14_EE4BEG[2] ,
    \Tile_X7Y14_EE4BEG[1] ,
    \Tile_X7Y14_EE4BEG[0] }),
    .Tile_X0Y1_EE4END({\Tile_X6Y14_EE4BEG[15] ,
    \Tile_X6Y14_EE4BEG[14] ,
    \Tile_X6Y14_EE4BEG[13] ,
    \Tile_X6Y14_EE4BEG[12] ,
    \Tile_X6Y14_EE4BEG[11] ,
    \Tile_X6Y14_EE4BEG[10] ,
    \Tile_X6Y14_EE4BEG[9] ,
    \Tile_X6Y14_EE4BEG[8] ,
    \Tile_X6Y14_EE4BEG[7] ,
    \Tile_X6Y14_EE4BEG[6] ,
    \Tile_X6Y14_EE4BEG[5] ,
    \Tile_X6Y14_EE4BEG[4] ,
    \Tile_X6Y14_EE4BEG[3] ,
    \Tile_X6Y14_EE4BEG[2] ,
    \Tile_X6Y14_EE4BEG[1] ,
    \Tile_X6Y14_EE4BEG[0] }),
    .Tile_X0Y1_FrameData({\Tile_X6Y14_FrameData_O[31] ,
    \Tile_X6Y14_FrameData_O[30] ,
    \Tile_X6Y14_FrameData_O[29] ,
    \Tile_X6Y14_FrameData_O[28] ,
    \Tile_X6Y14_FrameData_O[27] ,
    \Tile_X6Y14_FrameData_O[26] ,
    \Tile_X6Y14_FrameData_O[25] ,
    \Tile_X6Y14_FrameData_O[24] ,
    \Tile_X6Y14_FrameData_O[23] ,
    \Tile_X6Y14_FrameData_O[22] ,
    \Tile_X6Y14_FrameData_O[21] ,
    \Tile_X6Y14_FrameData_O[20] ,
    \Tile_X6Y14_FrameData_O[19] ,
    \Tile_X6Y14_FrameData_O[18] ,
    \Tile_X6Y14_FrameData_O[17] ,
    \Tile_X6Y14_FrameData_O[16] ,
    \Tile_X6Y14_FrameData_O[15] ,
    \Tile_X6Y14_FrameData_O[14] ,
    \Tile_X6Y14_FrameData_O[13] ,
    \Tile_X6Y14_FrameData_O[12] ,
    \Tile_X6Y14_FrameData_O[11] ,
    \Tile_X6Y14_FrameData_O[10] ,
    \Tile_X6Y14_FrameData_O[9] ,
    \Tile_X6Y14_FrameData_O[8] ,
    \Tile_X6Y14_FrameData_O[7] ,
    \Tile_X6Y14_FrameData_O[6] ,
    \Tile_X6Y14_FrameData_O[5] ,
    \Tile_X6Y14_FrameData_O[4] ,
    \Tile_X6Y14_FrameData_O[3] ,
    \Tile_X6Y14_FrameData_O[2] ,
    \Tile_X6Y14_FrameData_O[1] ,
    \Tile_X6Y14_FrameData_O[0] }),
    .Tile_X0Y1_FrameData_O({\Tile_X7Y14_FrameData_O[31] ,
    \Tile_X7Y14_FrameData_O[30] ,
    \Tile_X7Y14_FrameData_O[29] ,
    \Tile_X7Y14_FrameData_O[28] ,
    \Tile_X7Y14_FrameData_O[27] ,
    \Tile_X7Y14_FrameData_O[26] ,
    \Tile_X7Y14_FrameData_O[25] ,
    \Tile_X7Y14_FrameData_O[24] ,
    \Tile_X7Y14_FrameData_O[23] ,
    \Tile_X7Y14_FrameData_O[22] ,
    \Tile_X7Y14_FrameData_O[21] ,
    \Tile_X7Y14_FrameData_O[20] ,
    \Tile_X7Y14_FrameData_O[19] ,
    \Tile_X7Y14_FrameData_O[18] ,
    \Tile_X7Y14_FrameData_O[17] ,
    \Tile_X7Y14_FrameData_O[16] ,
    \Tile_X7Y14_FrameData_O[15] ,
    \Tile_X7Y14_FrameData_O[14] ,
    \Tile_X7Y14_FrameData_O[13] ,
    \Tile_X7Y14_FrameData_O[12] ,
    \Tile_X7Y14_FrameData_O[11] ,
    \Tile_X7Y14_FrameData_O[10] ,
    \Tile_X7Y14_FrameData_O[9] ,
    \Tile_X7Y14_FrameData_O[8] ,
    \Tile_X7Y14_FrameData_O[7] ,
    \Tile_X7Y14_FrameData_O[6] ,
    \Tile_X7Y14_FrameData_O[5] ,
    \Tile_X7Y14_FrameData_O[4] ,
    \Tile_X7Y14_FrameData_O[3] ,
    \Tile_X7Y14_FrameData_O[2] ,
    \Tile_X7Y14_FrameData_O[1] ,
    \Tile_X7Y14_FrameData_O[0] }),
    .Tile_X0Y1_FrameStrobe({\Tile_X7Y15_FrameStrobe_O[19] ,
    \Tile_X7Y15_FrameStrobe_O[18] ,
    \Tile_X7Y15_FrameStrobe_O[17] ,
    \Tile_X7Y15_FrameStrobe_O[16] ,
    \Tile_X7Y15_FrameStrobe_O[15] ,
    \Tile_X7Y15_FrameStrobe_O[14] ,
    \Tile_X7Y15_FrameStrobe_O[13] ,
    \Tile_X7Y15_FrameStrobe_O[12] ,
    \Tile_X7Y15_FrameStrobe_O[11] ,
    \Tile_X7Y15_FrameStrobe_O[10] ,
    \Tile_X7Y15_FrameStrobe_O[9] ,
    \Tile_X7Y15_FrameStrobe_O[8] ,
    \Tile_X7Y15_FrameStrobe_O[7] ,
    \Tile_X7Y15_FrameStrobe_O[6] ,
    \Tile_X7Y15_FrameStrobe_O[5] ,
    \Tile_X7Y15_FrameStrobe_O[4] ,
    \Tile_X7Y15_FrameStrobe_O[3] ,
    \Tile_X7Y15_FrameStrobe_O[2] ,
    \Tile_X7Y15_FrameStrobe_O[1] ,
    \Tile_X7Y15_FrameStrobe_O[0] }),
    .Tile_X0Y1_N1END({\Tile_X7Y15_N1BEG[3] ,
    \Tile_X7Y15_N1BEG[2] ,
    \Tile_X7Y15_N1BEG[1] ,
    \Tile_X7Y15_N1BEG[0] }),
    .Tile_X0Y1_N2END({\Tile_X7Y15_N2BEGb[7] ,
    \Tile_X7Y15_N2BEGb[6] ,
    \Tile_X7Y15_N2BEGb[5] ,
    \Tile_X7Y15_N2BEGb[4] ,
    \Tile_X7Y15_N2BEGb[3] ,
    \Tile_X7Y15_N2BEGb[2] ,
    \Tile_X7Y15_N2BEGb[1] ,
    \Tile_X7Y15_N2BEGb[0] }),
    .Tile_X0Y1_N2MID({\Tile_X7Y15_N2BEG[7] ,
    \Tile_X7Y15_N2BEG[6] ,
    \Tile_X7Y15_N2BEG[5] ,
    \Tile_X7Y15_N2BEG[4] ,
    \Tile_X7Y15_N2BEG[3] ,
    \Tile_X7Y15_N2BEG[2] ,
    \Tile_X7Y15_N2BEG[1] ,
    \Tile_X7Y15_N2BEG[0] }),
    .Tile_X0Y1_N4END({\Tile_X7Y15_N4BEG[15] ,
    \Tile_X7Y15_N4BEG[14] ,
    \Tile_X7Y15_N4BEG[13] ,
    \Tile_X7Y15_N4BEG[12] ,
    \Tile_X7Y15_N4BEG[11] ,
    \Tile_X7Y15_N4BEG[10] ,
    \Tile_X7Y15_N4BEG[9] ,
    \Tile_X7Y15_N4BEG[8] ,
    \Tile_X7Y15_N4BEG[7] ,
    \Tile_X7Y15_N4BEG[6] ,
    \Tile_X7Y15_N4BEG[5] ,
    \Tile_X7Y15_N4BEG[4] ,
    \Tile_X7Y15_N4BEG[3] ,
    \Tile_X7Y15_N4BEG[2] ,
    \Tile_X7Y15_N4BEG[1] ,
    \Tile_X7Y15_N4BEG[0] }),
    .Tile_X0Y1_NN4END({\Tile_X7Y15_NN4BEG[15] ,
    \Tile_X7Y15_NN4BEG[14] ,
    \Tile_X7Y15_NN4BEG[13] ,
    \Tile_X7Y15_NN4BEG[12] ,
    \Tile_X7Y15_NN4BEG[11] ,
    \Tile_X7Y15_NN4BEG[10] ,
    \Tile_X7Y15_NN4BEG[9] ,
    \Tile_X7Y15_NN4BEG[8] ,
    \Tile_X7Y15_NN4BEG[7] ,
    \Tile_X7Y15_NN4BEG[6] ,
    \Tile_X7Y15_NN4BEG[5] ,
    \Tile_X7Y15_NN4BEG[4] ,
    \Tile_X7Y15_NN4BEG[3] ,
    \Tile_X7Y15_NN4BEG[2] ,
    \Tile_X7Y15_NN4BEG[1] ,
    \Tile_X7Y15_NN4BEG[0] }),
    .Tile_X0Y1_S1BEG({\Tile_X7Y14_S1BEG[3] ,
    \Tile_X7Y14_S1BEG[2] ,
    \Tile_X7Y14_S1BEG[1] ,
    \Tile_X7Y14_S1BEG[0] }),
    .Tile_X0Y1_S2BEG({\Tile_X7Y14_S2BEG[7] ,
    \Tile_X7Y14_S2BEG[6] ,
    \Tile_X7Y14_S2BEG[5] ,
    \Tile_X7Y14_S2BEG[4] ,
    \Tile_X7Y14_S2BEG[3] ,
    \Tile_X7Y14_S2BEG[2] ,
    \Tile_X7Y14_S2BEG[1] ,
    \Tile_X7Y14_S2BEG[0] }),
    .Tile_X0Y1_S2BEGb({\Tile_X7Y14_S2BEGb[7] ,
    \Tile_X7Y14_S2BEGb[6] ,
    \Tile_X7Y14_S2BEGb[5] ,
    \Tile_X7Y14_S2BEGb[4] ,
    \Tile_X7Y14_S2BEGb[3] ,
    \Tile_X7Y14_S2BEGb[2] ,
    \Tile_X7Y14_S2BEGb[1] ,
    \Tile_X7Y14_S2BEGb[0] }),
    .Tile_X0Y1_S4BEG({\Tile_X7Y14_S4BEG[15] ,
    \Tile_X7Y14_S4BEG[14] ,
    \Tile_X7Y14_S4BEG[13] ,
    \Tile_X7Y14_S4BEG[12] ,
    \Tile_X7Y14_S4BEG[11] ,
    \Tile_X7Y14_S4BEG[10] ,
    \Tile_X7Y14_S4BEG[9] ,
    \Tile_X7Y14_S4BEG[8] ,
    \Tile_X7Y14_S4BEG[7] ,
    \Tile_X7Y14_S4BEG[6] ,
    \Tile_X7Y14_S4BEG[5] ,
    \Tile_X7Y14_S4BEG[4] ,
    \Tile_X7Y14_S4BEG[3] ,
    \Tile_X7Y14_S4BEG[2] ,
    \Tile_X7Y14_S4BEG[1] ,
    \Tile_X7Y14_S4BEG[0] }),
    .Tile_X0Y1_SS4BEG({\Tile_X7Y14_SS4BEG[15] ,
    \Tile_X7Y14_SS4BEG[14] ,
    \Tile_X7Y14_SS4BEG[13] ,
    \Tile_X7Y14_SS4BEG[12] ,
    \Tile_X7Y14_SS4BEG[11] ,
    \Tile_X7Y14_SS4BEG[10] ,
    \Tile_X7Y14_SS4BEG[9] ,
    \Tile_X7Y14_SS4BEG[8] ,
    \Tile_X7Y14_SS4BEG[7] ,
    \Tile_X7Y14_SS4BEG[6] ,
    \Tile_X7Y14_SS4BEG[5] ,
    \Tile_X7Y14_SS4BEG[4] ,
    \Tile_X7Y14_SS4BEG[3] ,
    \Tile_X7Y14_SS4BEG[2] ,
    \Tile_X7Y14_SS4BEG[1] ,
    \Tile_X7Y14_SS4BEG[0] }),
    .Tile_X0Y1_W1BEG({\Tile_X7Y14_W1BEG[3] ,
    \Tile_X7Y14_W1BEG[2] ,
    \Tile_X7Y14_W1BEG[1] ,
    \Tile_X7Y14_W1BEG[0] }),
    .Tile_X0Y1_W1END({\Tile_X8Y14_W1BEG[3] ,
    \Tile_X8Y14_W1BEG[2] ,
    \Tile_X8Y14_W1BEG[1] ,
    \Tile_X8Y14_W1BEG[0] }),
    .Tile_X0Y1_W2BEG({\Tile_X7Y14_W2BEG[7] ,
    \Tile_X7Y14_W2BEG[6] ,
    \Tile_X7Y14_W2BEG[5] ,
    \Tile_X7Y14_W2BEG[4] ,
    \Tile_X7Y14_W2BEG[3] ,
    \Tile_X7Y14_W2BEG[2] ,
    \Tile_X7Y14_W2BEG[1] ,
    \Tile_X7Y14_W2BEG[0] }),
    .Tile_X0Y1_W2BEGb({\Tile_X7Y14_W2BEGb[7] ,
    \Tile_X7Y14_W2BEGb[6] ,
    \Tile_X7Y14_W2BEGb[5] ,
    \Tile_X7Y14_W2BEGb[4] ,
    \Tile_X7Y14_W2BEGb[3] ,
    \Tile_X7Y14_W2BEGb[2] ,
    \Tile_X7Y14_W2BEGb[1] ,
    \Tile_X7Y14_W2BEGb[0] }),
    .Tile_X0Y1_W2END({\Tile_X8Y14_W2BEGb[7] ,
    \Tile_X8Y14_W2BEGb[6] ,
    \Tile_X8Y14_W2BEGb[5] ,
    \Tile_X8Y14_W2BEGb[4] ,
    \Tile_X8Y14_W2BEGb[3] ,
    \Tile_X8Y14_W2BEGb[2] ,
    \Tile_X8Y14_W2BEGb[1] ,
    \Tile_X8Y14_W2BEGb[0] }),
    .Tile_X0Y1_W2MID({\Tile_X8Y14_W2BEG[7] ,
    \Tile_X8Y14_W2BEG[6] ,
    \Tile_X8Y14_W2BEG[5] ,
    \Tile_X8Y14_W2BEG[4] ,
    \Tile_X8Y14_W2BEG[3] ,
    \Tile_X8Y14_W2BEG[2] ,
    \Tile_X8Y14_W2BEG[1] ,
    \Tile_X8Y14_W2BEG[0] }),
    .Tile_X0Y1_W6BEG({\Tile_X7Y14_W6BEG[11] ,
    \Tile_X7Y14_W6BEG[10] ,
    \Tile_X7Y14_W6BEG[9] ,
    \Tile_X7Y14_W6BEG[8] ,
    \Tile_X7Y14_W6BEG[7] ,
    \Tile_X7Y14_W6BEG[6] ,
    \Tile_X7Y14_W6BEG[5] ,
    \Tile_X7Y14_W6BEG[4] ,
    \Tile_X7Y14_W6BEG[3] ,
    \Tile_X7Y14_W6BEG[2] ,
    \Tile_X7Y14_W6BEG[1] ,
    \Tile_X7Y14_W6BEG[0] }),
    .Tile_X0Y1_W6END({\Tile_X8Y14_W6BEG[11] ,
    \Tile_X8Y14_W6BEG[10] ,
    \Tile_X8Y14_W6BEG[9] ,
    \Tile_X8Y14_W6BEG[8] ,
    \Tile_X8Y14_W6BEG[7] ,
    \Tile_X8Y14_W6BEG[6] ,
    \Tile_X8Y14_W6BEG[5] ,
    \Tile_X8Y14_W6BEG[4] ,
    \Tile_X8Y14_W6BEG[3] ,
    \Tile_X8Y14_W6BEG[2] ,
    \Tile_X8Y14_W6BEG[1] ,
    \Tile_X8Y14_W6BEG[0] }),
    .Tile_X0Y1_WW4BEG({\Tile_X7Y14_WW4BEG[15] ,
    \Tile_X7Y14_WW4BEG[14] ,
    \Tile_X7Y14_WW4BEG[13] ,
    \Tile_X7Y14_WW4BEG[12] ,
    \Tile_X7Y14_WW4BEG[11] ,
    \Tile_X7Y14_WW4BEG[10] ,
    \Tile_X7Y14_WW4BEG[9] ,
    \Tile_X7Y14_WW4BEG[8] ,
    \Tile_X7Y14_WW4BEG[7] ,
    \Tile_X7Y14_WW4BEG[6] ,
    \Tile_X7Y14_WW4BEG[5] ,
    \Tile_X7Y14_WW4BEG[4] ,
    \Tile_X7Y14_WW4BEG[3] ,
    \Tile_X7Y14_WW4BEG[2] ,
    \Tile_X7Y14_WW4BEG[1] ,
    \Tile_X7Y14_WW4BEG[0] }),
    .Tile_X0Y1_WW4END({\Tile_X8Y14_WW4BEG[15] ,
    \Tile_X8Y14_WW4BEG[14] ,
    \Tile_X8Y14_WW4BEG[13] ,
    \Tile_X8Y14_WW4BEG[12] ,
    \Tile_X8Y14_WW4BEG[11] ,
    \Tile_X8Y14_WW4BEG[10] ,
    \Tile_X8Y14_WW4BEG[9] ,
    \Tile_X8Y14_WW4BEG[8] ,
    \Tile_X8Y14_WW4BEG[7] ,
    \Tile_X8Y14_WW4BEG[6] ,
    \Tile_X8Y14_WW4BEG[5] ,
    \Tile_X8Y14_WW4BEG[4] ,
    \Tile_X8Y14_WW4BEG[3] ,
    \Tile_X8Y14_WW4BEG[2] ,
    \Tile_X8Y14_WW4BEG[1] ,
    \Tile_X8Y14_WW4BEG[0] }));
 S_term_DSP Tile_X7Y15_S_term_DSP (.UserCLK(UserCLK),
    .UserCLKo(Tile_X7Y15_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .FrameData({\Tile_X6Y15_FrameData_O[31] ,
    \Tile_X6Y15_FrameData_O[30] ,
    \Tile_X6Y15_FrameData_O[29] ,
    \Tile_X6Y15_FrameData_O[28] ,
    \Tile_X6Y15_FrameData_O[27] ,
    \Tile_X6Y15_FrameData_O[26] ,
    \Tile_X6Y15_FrameData_O[25] ,
    \Tile_X6Y15_FrameData_O[24] ,
    \Tile_X6Y15_FrameData_O[23] ,
    \Tile_X6Y15_FrameData_O[22] ,
    \Tile_X6Y15_FrameData_O[21] ,
    \Tile_X6Y15_FrameData_O[20] ,
    \Tile_X6Y15_FrameData_O[19] ,
    \Tile_X6Y15_FrameData_O[18] ,
    \Tile_X6Y15_FrameData_O[17] ,
    \Tile_X6Y15_FrameData_O[16] ,
    \Tile_X6Y15_FrameData_O[15] ,
    \Tile_X6Y15_FrameData_O[14] ,
    \Tile_X6Y15_FrameData_O[13] ,
    \Tile_X6Y15_FrameData_O[12] ,
    \Tile_X6Y15_FrameData_O[11] ,
    \Tile_X6Y15_FrameData_O[10] ,
    \Tile_X6Y15_FrameData_O[9] ,
    \Tile_X6Y15_FrameData_O[8] ,
    \Tile_X6Y15_FrameData_O[7] ,
    \Tile_X6Y15_FrameData_O[6] ,
    \Tile_X6Y15_FrameData_O[5] ,
    \Tile_X6Y15_FrameData_O[4] ,
    \Tile_X6Y15_FrameData_O[3] ,
    \Tile_X6Y15_FrameData_O[2] ,
    \Tile_X6Y15_FrameData_O[1] ,
    \Tile_X6Y15_FrameData_O[0] }),
    .FrameData_O({\Tile_X7Y15_FrameData_O[31] ,
    \Tile_X7Y15_FrameData_O[30] ,
    \Tile_X7Y15_FrameData_O[29] ,
    \Tile_X7Y15_FrameData_O[28] ,
    \Tile_X7Y15_FrameData_O[27] ,
    \Tile_X7Y15_FrameData_O[26] ,
    \Tile_X7Y15_FrameData_O[25] ,
    \Tile_X7Y15_FrameData_O[24] ,
    \Tile_X7Y15_FrameData_O[23] ,
    \Tile_X7Y15_FrameData_O[22] ,
    \Tile_X7Y15_FrameData_O[21] ,
    \Tile_X7Y15_FrameData_O[20] ,
    \Tile_X7Y15_FrameData_O[19] ,
    \Tile_X7Y15_FrameData_O[18] ,
    \Tile_X7Y15_FrameData_O[17] ,
    \Tile_X7Y15_FrameData_O[16] ,
    \Tile_X7Y15_FrameData_O[15] ,
    \Tile_X7Y15_FrameData_O[14] ,
    \Tile_X7Y15_FrameData_O[13] ,
    \Tile_X7Y15_FrameData_O[12] ,
    \Tile_X7Y15_FrameData_O[11] ,
    \Tile_X7Y15_FrameData_O[10] ,
    \Tile_X7Y15_FrameData_O[9] ,
    \Tile_X7Y15_FrameData_O[8] ,
    \Tile_X7Y15_FrameData_O[7] ,
    \Tile_X7Y15_FrameData_O[6] ,
    \Tile_X7Y15_FrameData_O[5] ,
    \Tile_X7Y15_FrameData_O[4] ,
    \Tile_X7Y15_FrameData_O[3] ,
    \Tile_X7Y15_FrameData_O[2] ,
    \Tile_X7Y15_FrameData_O[1] ,
    \Tile_X7Y15_FrameData_O[0] }),
    .FrameStrobe({FrameStrobe[159],
    FrameStrobe[158],
    FrameStrobe[157],
    FrameStrobe[156],
    FrameStrobe[155],
    FrameStrobe[154],
    FrameStrobe[153],
    FrameStrobe[152],
    FrameStrobe[151],
    FrameStrobe[150],
    FrameStrobe[149],
    FrameStrobe[148],
    FrameStrobe[147],
    FrameStrobe[146],
    FrameStrobe[145],
    FrameStrobe[144],
    FrameStrobe[143],
    FrameStrobe[142],
    FrameStrobe[141],
    FrameStrobe[140]}),
    .FrameStrobe_O({\Tile_X7Y15_FrameStrobe_O[19] ,
    \Tile_X7Y15_FrameStrobe_O[18] ,
    \Tile_X7Y15_FrameStrobe_O[17] ,
    \Tile_X7Y15_FrameStrobe_O[16] ,
    \Tile_X7Y15_FrameStrobe_O[15] ,
    \Tile_X7Y15_FrameStrobe_O[14] ,
    \Tile_X7Y15_FrameStrobe_O[13] ,
    \Tile_X7Y15_FrameStrobe_O[12] ,
    \Tile_X7Y15_FrameStrobe_O[11] ,
    \Tile_X7Y15_FrameStrobe_O[10] ,
    \Tile_X7Y15_FrameStrobe_O[9] ,
    \Tile_X7Y15_FrameStrobe_O[8] ,
    \Tile_X7Y15_FrameStrobe_O[7] ,
    \Tile_X7Y15_FrameStrobe_O[6] ,
    \Tile_X7Y15_FrameStrobe_O[5] ,
    \Tile_X7Y15_FrameStrobe_O[4] ,
    \Tile_X7Y15_FrameStrobe_O[3] ,
    \Tile_X7Y15_FrameStrobe_O[2] ,
    \Tile_X7Y15_FrameStrobe_O[1] ,
    \Tile_X7Y15_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X7Y15_N1BEG[3] ,
    \Tile_X7Y15_N1BEG[2] ,
    \Tile_X7Y15_N1BEG[1] ,
    \Tile_X7Y15_N1BEG[0] }),
    .N2BEG({\Tile_X7Y15_N2BEG[7] ,
    \Tile_X7Y15_N2BEG[6] ,
    \Tile_X7Y15_N2BEG[5] ,
    \Tile_X7Y15_N2BEG[4] ,
    \Tile_X7Y15_N2BEG[3] ,
    \Tile_X7Y15_N2BEG[2] ,
    \Tile_X7Y15_N2BEG[1] ,
    \Tile_X7Y15_N2BEG[0] }),
    .N2BEGb({\Tile_X7Y15_N2BEGb[7] ,
    \Tile_X7Y15_N2BEGb[6] ,
    \Tile_X7Y15_N2BEGb[5] ,
    \Tile_X7Y15_N2BEGb[4] ,
    \Tile_X7Y15_N2BEGb[3] ,
    \Tile_X7Y15_N2BEGb[2] ,
    \Tile_X7Y15_N2BEGb[1] ,
    \Tile_X7Y15_N2BEGb[0] }),
    .N4BEG({\Tile_X7Y15_N4BEG[15] ,
    \Tile_X7Y15_N4BEG[14] ,
    \Tile_X7Y15_N4BEG[13] ,
    \Tile_X7Y15_N4BEG[12] ,
    \Tile_X7Y15_N4BEG[11] ,
    \Tile_X7Y15_N4BEG[10] ,
    \Tile_X7Y15_N4BEG[9] ,
    \Tile_X7Y15_N4BEG[8] ,
    \Tile_X7Y15_N4BEG[7] ,
    \Tile_X7Y15_N4BEG[6] ,
    \Tile_X7Y15_N4BEG[5] ,
    \Tile_X7Y15_N4BEG[4] ,
    \Tile_X7Y15_N4BEG[3] ,
    \Tile_X7Y15_N4BEG[2] ,
    \Tile_X7Y15_N4BEG[1] ,
    \Tile_X7Y15_N4BEG[0] }),
    .NN4BEG({\Tile_X7Y15_NN4BEG[15] ,
    \Tile_X7Y15_NN4BEG[14] ,
    \Tile_X7Y15_NN4BEG[13] ,
    \Tile_X7Y15_NN4BEG[12] ,
    \Tile_X7Y15_NN4BEG[11] ,
    \Tile_X7Y15_NN4BEG[10] ,
    \Tile_X7Y15_NN4BEG[9] ,
    \Tile_X7Y15_NN4BEG[8] ,
    \Tile_X7Y15_NN4BEG[7] ,
    \Tile_X7Y15_NN4BEG[6] ,
    \Tile_X7Y15_NN4BEG[5] ,
    \Tile_X7Y15_NN4BEG[4] ,
    \Tile_X7Y15_NN4BEG[3] ,
    \Tile_X7Y15_NN4BEG[2] ,
    \Tile_X7Y15_NN4BEG[1] ,
    \Tile_X7Y15_NN4BEG[0] }),
    .S1END({\Tile_X7Y14_S1BEG[3] ,
    \Tile_X7Y14_S1BEG[2] ,
    \Tile_X7Y14_S1BEG[1] ,
    \Tile_X7Y14_S1BEG[0] }),
    .S2END({\Tile_X7Y14_S2BEGb[7] ,
    \Tile_X7Y14_S2BEGb[6] ,
    \Tile_X7Y14_S2BEGb[5] ,
    \Tile_X7Y14_S2BEGb[4] ,
    \Tile_X7Y14_S2BEGb[3] ,
    \Tile_X7Y14_S2BEGb[2] ,
    \Tile_X7Y14_S2BEGb[1] ,
    \Tile_X7Y14_S2BEGb[0] }),
    .S2MID({\Tile_X7Y14_S2BEG[7] ,
    \Tile_X7Y14_S2BEG[6] ,
    \Tile_X7Y14_S2BEG[5] ,
    \Tile_X7Y14_S2BEG[4] ,
    \Tile_X7Y14_S2BEG[3] ,
    \Tile_X7Y14_S2BEG[2] ,
    \Tile_X7Y14_S2BEG[1] ,
    \Tile_X7Y14_S2BEG[0] }),
    .S4END({\Tile_X7Y14_S4BEG[15] ,
    \Tile_X7Y14_S4BEG[14] ,
    \Tile_X7Y14_S4BEG[13] ,
    \Tile_X7Y14_S4BEG[12] ,
    \Tile_X7Y14_S4BEG[11] ,
    \Tile_X7Y14_S4BEG[10] ,
    \Tile_X7Y14_S4BEG[9] ,
    \Tile_X7Y14_S4BEG[8] ,
    \Tile_X7Y14_S4BEG[7] ,
    \Tile_X7Y14_S4BEG[6] ,
    \Tile_X7Y14_S4BEG[5] ,
    \Tile_X7Y14_S4BEG[4] ,
    \Tile_X7Y14_S4BEG[3] ,
    \Tile_X7Y14_S4BEG[2] ,
    \Tile_X7Y14_S4BEG[1] ,
    \Tile_X7Y14_S4BEG[0] }),
    .SS4END({\Tile_X7Y14_SS4BEG[15] ,
    \Tile_X7Y14_SS4BEG[14] ,
    \Tile_X7Y14_SS4BEG[13] ,
    \Tile_X7Y14_SS4BEG[12] ,
    \Tile_X7Y14_SS4BEG[11] ,
    \Tile_X7Y14_SS4BEG[10] ,
    \Tile_X7Y14_SS4BEG[9] ,
    \Tile_X7Y14_SS4BEG[8] ,
    \Tile_X7Y14_SS4BEG[7] ,
    \Tile_X7Y14_SS4BEG[6] ,
    \Tile_X7Y14_SS4BEG[5] ,
    \Tile_X7Y14_SS4BEG[4] ,
    \Tile_X7Y14_SS4BEG[3] ,
    \Tile_X7Y14_SS4BEG[2] ,
    \Tile_X7Y14_SS4BEG[1] ,
    \Tile_X7Y14_SS4BEG[0] }));
 DSP Tile_X7Y1_DSP (.Tile_X0Y0_UserCLKo(Tile_X7Y1_UserCLKo),
    .Tile_X0Y1_UserCLK(Tile_X7Y3_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .Tile_X0Y0_E1BEG({\Tile_X7Y1_E1BEG[3] ,
    \Tile_X7Y1_E1BEG[2] ,
    \Tile_X7Y1_E1BEG[1] ,
    \Tile_X7Y1_E1BEG[0] }),
    .Tile_X0Y0_E1END({\Tile_X6Y1_E1BEG[3] ,
    \Tile_X6Y1_E1BEG[2] ,
    \Tile_X6Y1_E1BEG[1] ,
    \Tile_X6Y1_E1BEG[0] }),
    .Tile_X0Y0_E2BEG({\Tile_X7Y1_E2BEG[7] ,
    \Tile_X7Y1_E2BEG[6] ,
    \Tile_X7Y1_E2BEG[5] ,
    \Tile_X7Y1_E2BEG[4] ,
    \Tile_X7Y1_E2BEG[3] ,
    \Tile_X7Y1_E2BEG[2] ,
    \Tile_X7Y1_E2BEG[1] ,
    \Tile_X7Y1_E2BEG[0] }),
    .Tile_X0Y0_E2BEGb({\Tile_X7Y1_E2BEGb[7] ,
    \Tile_X7Y1_E2BEGb[6] ,
    \Tile_X7Y1_E2BEGb[5] ,
    \Tile_X7Y1_E2BEGb[4] ,
    \Tile_X7Y1_E2BEGb[3] ,
    \Tile_X7Y1_E2BEGb[2] ,
    \Tile_X7Y1_E2BEGb[1] ,
    \Tile_X7Y1_E2BEGb[0] }),
    .Tile_X0Y0_E2END({\Tile_X6Y1_E2BEGb[7] ,
    \Tile_X6Y1_E2BEGb[6] ,
    \Tile_X6Y1_E2BEGb[5] ,
    \Tile_X6Y1_E2BEGb[4] ,
    \Tile_X6Y1_E2BEGb[3] ,
    \Tile_X6Y1_E2BEGb[2] ,
    \Tile_X6Y1_E2BEGb[1] ,
    \Tile_X6Y1_E2BEGb[0] }),
    .Tile_X0Y0_E2MID({\Tile_X6Y1_E2BEG[7] ,
    \Tile_X6Y1_E2BEG[6] ,
    \Tile_X6Y1_E2BEG[5] ,
    \Tile_X6Y1_E2BEG[4] ,
    \Tile_X6Y1_E2BEG[3] ,
    \Tile_X6Y1_E2BEG[2] ,
    \Tile_X6Y1_E2BEG[1] ,
    \Tile_X6Y1_E2BEG[0] }),
    .Tile_X0Y0_E6BEG({\Tile_X7Y1_E6BEG[11] ,
    \Tile_X7Y1_E6BEG[10] ,
    \Tile_X7Y1_E6BEG[9] ,
    \Tile_X7Y1_E6BEG[8] ,
    \Tile_X7Y1_E6BEG[7] ,
    \Tile_X7Y1_E6BEG[6] ,
    \Tile_X7Y1_E6BEG[5] ,
    \Tile_X7Y1_E6BEG[4] ,
    \Tile_X7Y1_E6BEG[3] ,
    \Tile_X7Y1_E6BEG[2] ,
    \Tile_X7Y1_E6BEG[1] ,
    \Tile_X7Y1_E6BEG[0] }),
    .Tile_X0Y0_E6END({\Tile_X6Y1_E6BEG[11] ,
    \Tile_X6Y1_E6BEG[10] ,
    \Tile_X6Y1_E6BEG[9] ,
    \Tile_X6Y1_E6BEG[8] ,
    \Tile_X6Y1_E6BEG[7] ,
    \Tile_X6Y1_E6BEG[6] ,
    \Tile_X6Y1_E6BEG[5] ,
    \Tile_X6Y1_E6BEG[4] ,
    \Tile_X6Y1_E6BEG[3] ,
    \Tile_X6Y1_E6BEG[2] ,
    \Tile_X6Y1_E6BEG[1] ,
    \Tile_X6Y1_E6BEG[0] }),
    .Tile_X0Y0_EE4BEG({\Tile_X7Y1_EE4BEG[15] ,
    \Tile_X7Y1_EE4BEG[14] ,
    \Tile_X7Y1_EE4BEG[13] ,
    \Tile_X7Y1_EE4BEG[12] ,
    \Tile_X7Y1_EE4BEG[11] ,
    \Tile_X7Y1_EE4BEG[10] ,
    \Tile_X7Y1_EE4BEG[9] ,
    \Tile_X7Y1_EE4BEG[8] ,
    \Tile_X7Y1_EE4BEG[7] ,
    \Tile_X7Y1_EE4BEG[6] ,
    \Tile_X7Y1_EE4BEG[5] ,
    \Tile_X7Y1_EE4BEG[4] ,
    \Tile_X7Y1_EE4BEG[3] ,
    \Tile_X7Y1_EE4BEG[2] ,
    \Tile_X7Y1_EE4BEG[1] ,
    \Tile_X7Y1_EE4BEG[0] }),
    .Tile_X0Y0_EE4END({\Tile_X6Y1_EE4BEG[15] ,
    \Tile_X6Y1_EE4BEG[14] ,
    \Tile_X6Y1_EE4BEG[13] ,
    \Tile_X6Y1_EE4BEG[12] ,
    \Tile_X6Y1_EE4BEG[11] ,
    \Tile_X6Y1_EE4BEG[10] ,
    \Tile_X6Y1_EE4BEG[9] ,
    \Tile_X6Y1_EE4BEG[8] ,
    \Tile_X6Y1_EE4BEG[7] ,
    \Tile_X6Y1_EE4BEG[6] ,
    \Tile_X6Y1_EE4BEG[5] ,
    \Tile_X6Y1_EE4BEG[4] ,
    \Tile_X6Y1_EE4BEG[3] ,
    \Tile_X6Y1_EE4BEG[2] ,
    \Tile_X6Y1_EE4BEG[1] ,
    \Tile_X6Y1_EE4BEG[0] }),
    .Tile_X0Y0_FrameData({\Tile_X6Y1_FrameData_O[31] ,
    \Tile_X6Y1_FrameData_O[30] ,
    \Tile_X6Y1_FrameData_O[29] ,
    \Tile_X6Y1_FrameData_O[28] ,
    \Tile_X6Y1_FrameData_O[27] ,
    \Tile_X6Y1_FrameData_O[26] ,
    \Tile_X6Y1_FrameData_O[25] ,
    \Tile_X6Y1_FrameData_O[24] ,
    \Tile_X6Y1_FrameData_O[23] ,
    \Tile_X6Y1_FrameData_O[22] ,
    \Tile_X6Y1_FrameData_O[21] ,
    \Tile_X6Y1_FrameData_O[20] ,
    \Tile_X6Y1_FrameData_O[19] ,
    \Tile_X6Y1_FrameData_O[18] ,
    \Tile_X6Y1_FrameData_O[17] ,
    \Tile_X6Y1_FrameData_O[16] ,
    \Tile_X6Y1_FrameData_O[15] ,
    \Tile_X6Y1_FrameData_O[14] ,
    \Tile_X6Y1_FrameData_O[13] ,
    \Tile_X6Y1_FrameData_O[12] ,
    \Tile_X6Y1_FrameData_O[11] ,
    \Tile_X6Y1_FrameData_O[10] ,
    \Tile_X6Y1_FrameData_O[9] ,
    \Tile_X6Y1_FrameData_O[8] ,
    \Tile_X6Y1_FrameData_O[7] ,
    \Tile_X6Y1_FrameData_O[6] ,
    \Tile_X6Y1_FrameData_O[5] ,
    \Tile_X6Y1_FrameData_O[4] ,
    \Tile_X6Y1_FrameData_O[3] ,
    \Tile_X6Y1_FrameData_O[2] ,
    \Tile_X6Y1_FrameData_O[1] ,
    \Tile_X6Y1_FrameData_O[0] }),
    .Tile_X0Y0_FrameData_O({\Tile_X7Y1_FrameData_O[31] ,
    \Tile_X7Y1_FrameData_O[30] ,
    \Tile_X7Y1_FrameData_O[29] ,
    \Tile_X7Y1_FrameData_O[28] ,
    \Tile_X7Y1_FrameData_O[27] ,
    \Tile_X7Y1_FrameData_O[26] ,
    \Tile_X7Y1_FrameData_O[25] ,
    \Tile_X7Y1_FrameData_O[24] ,
    \Tile_X7Y1_FrameData_O[23] ,
    \Tile_X7Y1_FrameData_O[22] ,
    \Tile_X7Y1_FrameData_O[21] ,
    \Tile_X7Y1_FrameData_O[20] ,
    \Tile_X7Y1_FrameData_O[19] ,
    \Tile_X7Y1_FrameData_O[18] ,
    \Tile_X7Y1_FrameData_O[17] ,
    \Tile_X7Y1_FrameData_O[16] ,
    \Tile_X7Y1_FrameData_O[15] ,
    \Tile_X7Y1_FrameData_O[14] ,
    \Tile_X7Y1_FrameData_O[13] ,
    \Tile_X7Y1_FrameData_O[12] ,
    \Tile_X7Y1_FrameData_O[11] ,
    \Tile_X7Y1_FrameData_O[10] ,
    \Tile_X7Y1_FrameData_O[9] ,
    \Tile_X7Y1_FrameData_O[8] ,
    \Tile_X7Y1_FrameData_O[7] ,
    \Tile_X7Y1_FrameData_O[6] ,
    \Tile_X7Y1_FrameData_O[5] ,
    \Tile_X7Y1_FrameData_O[4] ,
    \Tile_X7Y1_FrameData_O[3] ,
    \Tile_X7Y1_FrameData_O[2] ,
    \Tile_X7Y1_FrameData_O[1] ,
    \Tile_X7Y1_FrameData_O[0] }),
    .Tile_X0Y0_FrameStrobe_O({\Tile_X7Y1_FrameStrobe_O[19] ,
    \Tile_X7Y1_FrameStrobe_O[18] ,
    \Tile_X7Y1_FrameStrobe_O[17] ,
    \Tile_X7Y1_FrameStrobe_O[16] ,
    \Tile_X7Y1_FrameStrobe_O[15] ,
    \Tile_X7Y1_FrameStrobe_O[14] ,
    \Tile_X7Y1_FrameStrobe_O[13] ,
    \Tile_X7Y1_FrameStrobe_O[12] ,
    \Tile_X7Y1_FrameStrobe_O[11] ,
    \Tile_X7Y1_FrameStrobe_O[10] ,
    \Tile_X7Y1_FrameStrobe_O[9] ,
    \Tile_X7Y1_FrameStrobe_O[8] ,
    \Tile_X7Y1_FrameStrobe_O[7] ,
    \Tile_X7Y1_FrameStrobe_O[6] ,
    \Tile_X7Y1_FrameStrobe_O[5] ,
    \Tile_X7Y1_FrameStrobe_O[4] ,
    \Tile_X7Y1_FrameStrobe_O[3] ,
    \Tile_X7Y1_FrameStrobe_O[2] ,
    \Tile_X7Y1_FrameStrobe_O[1] ,
    \Tile_X7Y1_FrameStrobe_O[0] }),
    .Tile_X0Y0_N1BEG({\Tile_X7Y1_N1BEG[3] ,
    \Tile_X7Y1_N1BEG[2] ,
    \Tile_X7Y1_N1BEG[1] ,
    \Tile_X7Y1_N1BEG[0] }),
    .Tile_X0Y0_N2BEG({\Tile_X7Y1_N2BEG[7] ,
    \Tile_X7Y1_N2BEG[6] ,
    \Tile_X7Y1_N2BEG[5] ,
    \Tile_X7Y1_N2BEG[4] ,
    \Tile_X7Y1_N2BEG[3] ,
    \Tile_X7Y1_N2BEG[2] ,
    \Tile_X7Y1_N2BEG[1] ,
    \Tile_X7Y1_N2BEG[0] }),
    .Tile_X0Y0_N2BEGb({\Tile_X7Y1_N2BEGb[7] ,
    \Tile_X7Y1_N2BEGb[6] ,
    \Tile_X7Y1_N2BEGb[5] ,
    \Tile_X7Y1_N2BEGb[4] ,
    \Tile_X7Y1_N2BEGb[3] ,
    \Tile_X7Y1_N2BEGb[2] ,
    \Tile_X7Y1_N2BEGb[1] ,
    \Tile_X7Y1_N2BEGb[0] }),
    .Tile_X0Y0_N4BEG({\Tile_X7Y1_N4BEG[15] ,
    \Tile_X7Y1_N4BEG[14] ,
    \Tile_X7Y1_N4BEG[13] ,
    \Tile_X7Y1_N4BEG[12] ,
    \Tile_X7Y1_N4BEG[11] ,
    \Tile_X7Y1_N4BEG[10] ,
    \Tile_X7Y1_N4BEG[9] ,
    \Tile_X7Y1_N4BEG[8] ,
    \Tile_X7Y1_N4BEG[7] ,
    \Tile_X7Y1_N4BEG[6] ,
    \Tile_X7Y1_N4BEG[5] ,
    \Tile_X7Y1_N4BEG[4] ,
    \Tile_X7Y1_N4BEG[3] ,
    \Tile_X7Y1_N4BEG[2] ,
    \Tile_X7Y1_N4BEG[1] ,
    \Tile_X7Y1_N4BEG[0] }),
    .Tile_X0Y0_NN4BEG({\Tile_X7Y1_NN4BEG[15] ,
    \Tile_X7Y1_NN4BEG[14] ,
    \Tile_X7Y1_NN4BEG[13] ,
    \Tile_X7Y1_NN4BEG[12] ,
    \Tile_X7Y1_NN4BEG[11] ,
    \Tile_X7Y1_NN4BEG[10] ,
    \Tile_X7Y1_NN4BEG[9] ,
    \Tile_X7Y1_NN4BEG[8] ,
    \Tile_X7Y1_NN4BEG[7] ,
    \Tile_X7Y1_NN4BEG[6] ,
    \Tile_X7Y1_NN4BEG[5] ,
    \Tile_X7Y1_NN4BEG[4] ,
    \Tile_X7Y1_NN4BEG[3] ,
    \Tile_X7Y1_NN4BEG[2] ,
    \Tile_X7Y1_NN4BEG[1] ,
    \Tile_X7Y1_NN4BEG[0] }),
    .Tile_X0Y0_S1END({\Tile_X7Y0_S1BEG[3] ,
    \Tile_X7Y0_S1BEG[2] ,
    \Tile_X7Y0_S1BEG[1] ,
    \Tile_X7Y0_S1BEG[0] }),
    .Tile_X0Y0_S2END({\Tile_X7Y0_S2BEGb[7] ,
    \Tile_X7Y0_S2BEGb[6] ,
    \Tile_X7Y0_S2BEGb[5] ,
    \Tile_X7Y0_S2BEGb[4] ,
    \Tile_X7Y0_S2BEGb[3] ,
    \Tile_X7Y0_S2BEGb[2] ,
    \Tile_X7Y0_S2BEGb[1] ,
    \Tile_X7Y0_S2BEGb[0] }),
    .Tile_X0Y0_S2MID({\Tile_X7Y0_S2BEG[7] ,
    \Tile_X7Y0_S2BEG[6] ,
    \Tile_X7Y0_S2BEG[5] ,
    \Tile_X7Y0_S2BEG[4] ,
    \Tile_X7Y0_S2BEG[3] ,
    \Tile_X7Y0_S2BEG[2] ,
    \Tile_X7Y0_S2BEG[1] ,
    \Tile_X7Y0_S2BEG[0] }),
    .Tile_X0Y0_S4END({\Tile_X7Y0_S4BEG[15] ,
    \Tile_X7Y0_S4BEG[14] ,
    \Tile_X7Y0_S4BEG[13] ,
    \Tile_X7Y0_S4BEG[12] ,
    \Tile_X7Y0_S4BEG[11] ,
    \Tile_X7Y0_S4BEG[10] ,
    \Tile_X7Y0_S4BEG[9] ,
    \Tile_X7Y0_S4BEG[8] ,
    \Tile_X7Y0_S4BEG[7] ,
    \Tile_X7Y0_S4BEG[6] ,
    \Tile_X7Y0_S4BEG[5] ,
    \Tile_X7Y0_S4BEG[4] ,
    \Tile_X7Y0_S4BEG[3] ,
    \Tile_X7Y0_S4BEG[2] ,
    \Tile_X7Y0_S4BEG[1] ,
    \Tile_X7Y0_S4BEG[0] }),
    .Tile_X0Y0_SS4END({\Tile_X7Y0_SS4BEG[15] ,
    \Tile_X7Y0_SS4BEG[14] ,
    \Tile_X7Y0_SS4BEG[13] ,
    \Tile_X7Y0_SS4BEG[12] ,
    \Tile_X7Y0_SS4BEG[11] ,
    \Tile_X7Y0_SS4BEG[10] ,
    \Tile_X7Y0_SS4BEG[9] ,
    \Tile_X7Y0_SS4BEG[8] ,
    \Tile_X7Y0_SS4BEG[7] ,
    \Tile_X7Y0_SS4BEG[6] ,
    \Tile_X7Y0_SS4BEG[5] ,
    \Tile_X7Y0_SS4BEG[4] ,
    \Tile_X7Y0_SS4BEG[3] ,
    \Tile_X7Y0_SS4BEG[2] ,
    \Tile_X7Y0_SS4BEG[1] ,
    \Tile_X7Y0_SS4BEG[0] }),
    .Tile_X0Y0_W1BEG({\Tile_X7Y1_W1BEG[3] ,
    \Tile_X7Y1_W1BEG[2] ,
    \Tile_X7Y1_W1BEG[1] ,
    \Tile_X7Y1_W1BEG[0] }),
    .Tile_X0Y0_W1END({\Tile_X8Y1_W1BEG[3] ,
    \Tile_X8Y1_W1BEG[2] ,
    \Tile_X8Y1_W1BEG[1] ,
    \Tile_X8Y1_W1BEG[0] }),
    .Tile_X0Y0_W2BEG({\Tile_X7Y1_W2BEG[7] ,
    \Tile_X7Y1_W2BEG[6] ,
    \Tile_X7Y1_W2BEG[5] ,
    \Tile_X7Y1_W2BEG[4] ,
    \Tile_X7Y1_W2BEG[3] ,
    \Tile_X7Y1_W2BEG[2] ,
    \Tile_X7Y1_W2BEG[1] ,
    \Tile_X7Y1_W2BEG[0] }),
    .Tile_X0Y0_W2BEGb({\Tile_X7Y1_W2BEGb[7] ,
    \Tile_X7Y1_W2BEGb[6] ,
    \Tile_X7Y1_W2BEGb[5] ,
    \Tile_X7Y1_W2BEGb[4] ,
    \Tile_X7Y1_W2BEGb[3] ,
    \Tile_X7Y1_W2BEGb[2] ,
    \Tile_X7Y1_W2BEGb[1] ,
    \Tile_X7Y1_W2BEGb[0] }),
    .Tile_X0Y0_W2END({\Tile_X8Y1_W2BEGb[7] ,
    \Tile_X8Y1_W2BEGb[6] ,
    \Tile_X8Y1_W2BEGb[5] ,
    \Tile_X8Y1_W2BEGb[4] ,
    \Tile_X8Y1_W2BEGb[3] ,
    \Tile_X8Y1_W2BEGb[2] ,
    \Tile_X8Y1_W2BEGb[1] ,
    \Tile_X8Y1_W2BEGb[0] }),
    .Tile_X0Y0_W2MID({\Tile_X8Y1_W2BEG[7] ,
    \Tile_X8Y1_W2BEG[6] ,
    \Tile_X8Y1_W2BEG[5] ,
    \Tile_X8Y1_W2BEG[4] ,
    \Tile_X8Y1_W2BEG[3] ,
    \Tile_X8Y1_W2BEG[2] ,
    \Tile_X8Y1_W2BEG[1] ,
    \Tile_X8Y1_W2BEG[0] }),
    .Tile_X0Y0_W6BEG({\Tile_X7Y1_W6BEG[11] ,
    \Tile_X7Y1_W6BEG[10] ,
    \Tile_X7Y1_W6BEG[9] ,
    \Tile_X7Y1_W6BEG[8] ,
    \Tile_X7Y1_W6BEG[7] ,
    \Tile_X7Y1_W6BEG[6] ,
    \Tile_X7Y1_W6BEG[5] ,
    \Tile_X7Y1_W6BEG[4] ,
    \Tile_X7Y1_W6BEG[3] ,
    \Tile_X7Y1_W6BEG[2] ,
    \Tile_X7Y1_W6BEG[1] ,
    \Tile_X7Y1_W6BEG[0] }),
    .Tile_X0Y0_W6END({\Tile_X8Y1_W6BEG[11] ,
    \Tile_X8Y1_W6BEG[10] ,
    \Tile_X8Y1_W6BEG[9] ,
    \Tile_X8Y1_W6BEG[8] ,
    \Tile_X8Y1_W6BEG[7] ,
    \Tile_X8Y1_W6BEG[6] ,
    \Tile_X8Y1_W6BEG[5] ,
    \Tile_X8Y1_W6BEG[4] ,
    \Tile_X8Y1_W6BEG[3] ,
    \Tile_X8Y1_W6BEG[2] ,
    \Tile_X8Y1_W6BEG[1] ,
    \Tile_X8Y1_W6BEG[0] }),
    .Tile_X0Y0_WW4BEG({\Tile_X7Y1_WW4BEG[15] ,
    \Tile_X7Y1_WW4BEG[14] ,
    \Tile_X7Y1_WW4BEG[13] ,
    \Tile_X7Y1_WW4BEG[12] ,
    \Tile_X7Y1_WW4BEG[11] ,
    \Tile_X7Y1_WW4BEG[10] ,
    \Tile_X7Y1_WW4BEG[9] ,
    \Tile_X7Y1_WW4BEG[8] ,
    \Tile_X7Y1_WW4BEG[7] ,
    \Tile_X7Y1_WW4BEG[6] ,
    \Tile_X7Y1_WW4BEG[5] ,
    \Tile_X7Y1_WW4BEG[4] ,
    \Tile_X7Y1_WW4BEG[3] ,
    \Tile_X7Y1_WW4BEG[2] ,
    \Tile_X7Y1_WW4BEG[1] ,
    \Tile_X7Y1_WW4BEG[0] }),
    .Tile_X0Y0_WW4END({\Tile_X8Y1_WW4BEG[15] ,
    \Tile_X8Y1_WW4BEG[14] ,
    \Tile_X8Y1_WW4BEG[13] ,
    \Tile_X8Y1_WW4BEG[12] ,
    \Tile_X8Y1_WW4BEG[11] ,
    \Tile_X8Y1_WW4BEG[10] ,
    \Tile_X8Y1_WW4BEG[9] ,
    \Tile_X8Y1_WW4BEG[8] ,
    \Tile_X8Y1_WW4BEG[7] ,
    \Tile_X8Y1_WW4BEG[6] ,
    \Tile_X8Y1_WW4BEG[5] ,
    \Tile_X8Y1_WW4BEG[4] ,
    \Tile_X8Y1_WW4BEG[3] ,
    \Tile_X8Y1_WW4BEG[2] ,
    \Tile_X8Y1_WW4BEG[1] ,
    \Tile_X8Y1_WW4BEG[0] }),
    .Tile_X0Y1_E1BEG({\Tile_X7Y2_E1BEG[3] ,
    \Tile_X7Y2_E1BEG[2] ,
    \Tile_X7Y2_E1BEG[1] ,
    \Tile_X7Y2_E1BEG[0] }),
    .Tile_X0Y1_E1END({\Tile_X6Y2_E1BEG[3] ,
    \Tile_X6Y2_E1BEG[2] ,
    \Tile_X6Y2_E1BEG[1] ,
    \Tile_X6Y2_E1BEG[0] }),
    .Tile_X0Y1_E2BEG({\Tile_X7Y2_E2BEG[7] ,
    \Tile_X7Y2_E2BEG[6] ,
    \Tile_X7Y2_E2BEG[5] ,
    \Tile_X7Y2_E2BEG[4] ,
    \Tile_X7Y2_E2BEG[3] ,
    \Tile_X7Y2_E2BEG[2] ,
    \Tile_X7Y2_E2BEG[1] ,
    \Tile_X7Y2_E2BEG[0] }),
    .Tile_X0Y1_E2BEGb({\Tile_X7Y2_E2BEGb[7] ,
    \Tile_X7Y2_E2BEGb[6] ,
    \Tile_X7Y2_E2BEGb[5] ,
    \Tile_X7Y2_E2BEGb[4] ,
    \Tile_X7Y2_E2BEGb[3] ,
    \Tile_X7Y2_E2BEGb[2] ,
    \Tile_X7Y2_E2BEGb[1] ,
    \Tile_X7Y2_E2BEGb[0] }),
    .Tile_X0Y1_E2END({\Tile_X6Y2_E2BEGb[7] ,
    \Tile_X6Y2_E2BEGb[6] ,
    \Tile_X6Y2_E2BEGb[5] ,
    \Tile_X6Y2_E2BEGb[4] ,
    \Tile_X6Y2_E2BEGb[3] ,
    \Tile_X6Y2_E2BEGb[2] ,
    \Tile_X6Y2_E2BEGb[1] ,
    \Tile_X6Y2_E2BEGb[0] }),
    .Tile_X0Y1_E2MID({\Tile_X6Y2_E2BEG[7] ,
    \Tile_X6Y2_E2BEG[6] ,
    \Tile_X6Y2_E2BEG[5] ,
    \Tile_X6Y2_E2BEG[4] ,
    \Tile_X6Y2_E2BEG[3] ,
    \Tile_X6Y2_E2BEG[2] ,
    \Tile_X6Y2_E2BEG[1] ,
    \Tile_X6Y2_E2BEG[0] }),
    .Tile_X0Y1_E6BEG({\Tile_X7Y2_E6BEG[11] ,
    \Tile_X7Y2_E6BEG[10] ,
    \Tile_X7Y2_E6BEG[9] ,
    \Tile_X7Y2_E6BEG[8] ,
    \Tile_X7Y2_E6BEG[7] ,
    \Tile_X7Y2_E6BEG[6] ,
    \Tile_X7Y2_E6BEG[5] ,
    \Tile_X7Y2_E6BEG[4] ,
    \Tile_X7Y2_E6BEG[3] ,
    \Tile_X7Y2_E6BEG[2] ,
    \Tile_X7Y2_E6BEG[1] ,
    \Tile_X7Y2_E6BEG[0] }),
    .Tile_X0Y1_E6END({\Tile_X6Y2_E6BEG[11] ,
    \Tile_X6Y2_E6BEG[10] ,
    \Tile_X6Y2_E6BEG[9] ,
    \Tile_X6Y2_E6BEG[8] ,
    \Tile_X6Y2_E6BEG[7] ,
    \Tile_X6Y2_E6BEG[6] ,
    \Tile_X6Y2_E6BEG[5] ,
    \Tile_X6Y2_E6BEG[4] ,
    \Tile_X6Y2_E6BEG[3] ,
    \Tile_X6Y2_E6BEG[2] ,
    \Tile_X6Y2_E6BEG[1] ,
    \Tile_X6Y2_E6BEG[0] }),
    .Tile_X0Y1_EE4BEG({\Tile_X7Y2_EE4BEG[15] ,
    \Tile_X7Y2_EE4BEG[14] ,
    \Tile_X7Y2_EE4BEG[13] ,
    \Tile_X7Y2_EE4BEG[12] ,
    \Tile_X7Y2_EE4BEG[11] ,
    \Tile_X7Y2_EE4BEG[10] ,
    \Tile_X7Y2_EE4BEG[9] ,
    \Tile_X7Y2_EE4BEG[8] ,
    \Tile_X7Y2_EE4BEG[7] ,
    \Tile_X7Y2_EE4BEG[6] ,
    \Tile_X7Y2_EE4BEG[5] ,
    \Tile_X7Y2_EE4BEG[4] ,
    \Tile_X7Y2_EE4BEG[3] ,
    \Tile_X7Y2_EE4BEG[2] ,
    \Tile_X7Y2_EE4BEG[1] ,
    \Tile_X7Y2_EE4BEG[0] }),
    .Tile_X0Y1_EE4END({\Tile_X6Y2_EE4BEG[15] ,
    \Tile_X6Y2_EE4BEG[14] ,
    \Tile_X6Y2_EE4BEG[13] ,
    \Tile_X6Y2_EE4BEG[12] ,
    \Tile_X6Y2_EE4BEG[11] ,
    \Tile_X6Y2_EE4BEG[10] ,
    \Tile_X6Y2_EE4BEG[9] ,
    \Tile_X6Y2_EE4BEG[8] ,
    \Tile_X6Y2_EE4BEG[7] ,
    \Tile_X6Y2_EE4BEG[6] ,
    \Tile_X6Y2_EE4BEG[5] ,
    \Tile_X6Y2_EE4BEG[4] ,
    \Tile_X6Y2_EE4BEG[3] ,
    \Tile_X6Y2_EE4BEG[2] ,
    \Tile_X6Y2_EE4BEG[1] ,
    \Tile_X6Y2_EE4BEG[0] }),
    .Tile_X0Y1_FrameData({\Tile_X6Y2_FrameData_O[31] ,
    \Tile_X6Y2_FrameData_O[30] ,
    \Tile_X6Y2_FrameData_O[29] ,
    \Tile_X6Y2_FrameData_O[28] ,
    \Tile_X6Y2_FrameData_O[27] ,
    \Tile_X6Y2_FrameData_O[26] ,
    \Tile_X6Y2_FrameData_O[25] ,
    \Tile_X6Y2_FrameData_O[24] ,
    \Tile_X6Y2_FrameData_O[23] ,
    \Tile_X6Y2_FrameData_O[22] ,
    \Tile_X6Y2_FrameData_O[21] ,
    \Tile_X6Y2_FrameData_O[20] ,
    \Tile_X6Y2_FrameData_O[19] ,
    \Tile_X6Y2_FrameData_O[18] ,
    \Tile_X6Y2_FrameData_O[17] ,
    \Tile_X6Y2_FrameData_O[16] ,
    \Tile_X6Y2_FrameData_O[15] ,
    \Tile_X6Y2_FrameData_O[14] ,
    \Tile_X6Y2_FrameData_O[13] ,
    \Tile_X6Y2_FrameData_O[12] ,
    \Tile_X6Y2_FrameData_O[11] ,
    \Tile_X6Y2_FrameData_O[10] ,
    \Tile_X6Y2_FrameData_O[9] ,
    \Tile_X6Y2_FrameData_O[8] ,
    \Tile_X6Y2_FrameData_O[7] ,
    \Tile_X6Y2_FrameData_O[6] ,
    \Tile_X6Y2_FrameData_O[5] ,
    \Tile_X6Y2_FrameData_O[4] ,
    \Tile_X6Y2_FrameData_O[3] ,
    \Tile_X6Y2_FrameData_O[2] ,
    \Tile_X6Y2_FrameData_O[1] ,
    \Tile_X6Y2_FrameData_O[0] }),
    .Tile_X0Y1_FrameData_O({\Tile_X7Y2_FrameData_O[31] ,
    \Tile_X7Y2_FrameData_O[30] ,
    \Tile_X7Y2_FrameData_O[29] ,
    \Tile_X7Y2_FrameData_O[28] ,
    \Tile_X7Y2_FrameData_O[27] ,
    \Tile_X7Y2_FrameData_O[26] ,
    \Tile_X7Y2_FrameData_O[25] ,
    \Tile_X7Y2_FrameData_O[24] ,
    \Tile_X7Y2_FrameData_O[23] ,
    \Tile_X7Y2_FrameData_O[22] ,
    \Tile_X7Y2_FrameData_O[21] ,
    \Tile_X7Y2_FrameData_O[20] ,
    \Tile_X7Y2_FrameData_O[19] ,
    \Tile_X7Y2_FrameData_O[18] ,
    \Tile_X7Y2_FrameData_O[17] ,
    \Tile_X7Y2_FrameData_O[16] ,
    \Tile_X7Y2_FrameData_O[15] ,
    \Tile_X7Y2_FrameData_O[14] ,
    \Tile_X7Y2_FrameData_O[13] ,
    \Tile_X7Y2_FrameData_O[12] ,
    \Tile_X7Y2_FrameData_O[11] ,
    \Tile_X7Y2_FrameData_O[10] ,
    \Tile_X7Y2_FrameData_O[9] ,
    \Tile_X7Y2_FrameData_O[8] ,
    \Tile_X7Y2_FrameData_O[7] ,
    \Tile_X7Y2_FrameData_O[6] ,
    \Tile_X7Y2_FrameData_O[5] ,
    \Tile_X7Y2_FrameData_O[4] ,
    \Tile_X7Y2_FrameData_O[3] ,
    \Tile_X7Y2_FrameData_O[2] ,
    \Tile_X7Y2_FrameData_O[1] ,
    \Tile_X7Y2_FrameData_O[0] }),
    .Tile_X0Y1_FrameStrobe({\Tile_X7Y3_FrameStrobe_O[19] ,
    \Tile_X7Y3_FrameStrobe_O[18] ,
    \Tile_X7Y3_FrameStrobe_O[17] ,
    \Tile_X7Y3_FrameStrobe_O[16] ,
    \Tile_X7Y3_FrameStrobe_O[15] ,
    \Tile_X7Y3_FrameStrobe_O[14] ,
    \Tile_X7Y3_FrameStrobe_O[13] ,
    \Tile_X7Y3_FrameStrobe_O[12] ,
    \Tile_X7Y3_FrameStrobe_O[11] ,
    \Tile_X7Y3_FrameStrobe_O[10] ,
    \Tile_X7Y3_FrameStrobe_O[9] ,
    \Tile_X7Y3_FrameStrobe_O[8] ,
    \Tile_X7Y3_FrameStrobe_O[7] ,
    \Tile_X7Y3_FrameStrobe_O[6] ,
    \Tile_X7Y3_FrameStrobe_O[5] ,
    \Tile_X7Y3_FrameStrobe_O[4] ,
    \Tile_X7Y3_FrameStrobe_O[3] ,
    \Tile_X7Y3_FrameStrobe_O[2] ,
    \Tile_X7Y3_FrameStrobe_O[1] ,
    \Tile_X7Y3_FrameStrobe_O[0] }),
    .Tile_X0Y1_N1END({\Tile_X7Y3_N1BEG[3] ,
    \Tile_X7Y3_N1BEG[2] ,
    \Tile_X7Y3_N1BEG[1] ,
    \Tile_X7Y3_N1BEG[0] }),
    .Tile_X0Y1_N2END({\Tile_X7Y3_N2BEGb[7] ,
    \Tile_X7Y3_N2BEGb[6] ,
    \Tile_X7Y3_N2BEGb[5] ,
    \Tile_X7Y3_N2BEGb[4] ,
    \Tile_X7Y3_N2BEGb[3] ,
    \Tile_X7Y3_N2BEGb[2] ,
    \Tile_X7Y3_N2BEGb[1] ,
    \Tile_X7Y3_N2BEGb[0] }),
    .Tile_X0Y1_N2MID({\Tile_X7Y3_N2BEG[7] ,
    \Tile_X7Y3_N2BEG[6] ,
    \Tile_X7Y3_N2BEG[5] ,
    \Tile_X7Y3_N2BEG[4] ,
    \Tile_X7Y3_N2BEG[3] ,
    \Tile_X7Y3_N2BEG[2] ,
    \Tile_X7Y3_N2BEG[1] ,
    \Tile_X7Y3_N2BEG[0] }),
    .Tile_X0Y1_N4END({\Tile_X7Y3_N4BEG[15] ,
    \Tile_X7Y3_N4BEG[14] ,
    \Tile_X7Y3_N4BEG[13] ,
    \Tile_X7Y3_N4BEG[12] ,
    \Tile_X7Y3_N4BEG[11] ,
    \Tile_X7Y3_N4BEG[10] ,
    \Tile_X7Y3_N4BEG[9] ,
    \Tile_X7Y3_N4BEG[8] ,
    \Tile_X7Y3_N4BEG[7] ,
    \Tile_X7Y3_N4BEG[6] ,
    \Tile_X7Y3_N4BEG[5] ,
    \Tile_X7Y3_N4BEG[4] ,
    \Tile_X7Y3_N4BEG[3] ,
    \Tile_X7Y3_N4BEG[2] ,
    \Tile_X7Y3_N4BEG[1] ,
    \Tile_X7Y3_N4BEG[0] }),
    .Tile_X0Y1_NN4END({\Tile_X7Y3_NN4BEG[15] ,
    \Tile_X7Y3_NN4BEG[14] ,
    \Tile_X7Y3_NN4BEG[13] ,
    \Tile_X7Y3_NN4BEG[12] ,
    \Tile_X7Y3_NN4BEG[11] ,
    \Tile_X7Y3_NN4BEG[10] ,
    \Tile_X7Y3_NN4BEG[9] ,
    \Tile_X7Y3_NN4BEG[8] ,
    \Tile_X7Y3_NN4BEG[7] ,
    \Tile_X7Y3_NN4BEG[6] ,
    \Tile_X7Y3_NN4BEG[5] ,
    \Tile_X7Y3_NN4BEG[4] ,
    \Tile_X7Y3_NN4BEG[3] ,
    \Tile_X7Y3_NN4BEG[2] ,
    \Tile_X7Y3_NN4BEG[1] ,
    \Tile_X7Y3_NN4BEG[0] }),
    .Tile_X0Y1_S1BEG({\Tile_X7Y2_S1BEG[3] ,
    \Tile_X7Y2_S1BEG[2] ,
    \Tile_X7Y2_S1BEG[1] ,
    \Tile_X7Y2_S1BEG[0] }),
    .Tile_X0Y1_S2BEG({\Tile_X7Y2_S2BEG[7] ,
    \Tile_X7Y2_S2BEG[6] ,
    \Tile_X7Y2_S2BEG[5] ,
    \Tile_X7Y2_S2BEG[4] ,
    \Tile_X7Y2_S2BEG[3] ,
    \Tile_X7Y2_S2BEG[2] ,
    \Tile_X7Y2_S2BEG[1] ,
    \Tile_X7Y2_S2BEG[0] }),
    .Tile_X0Y1_S2BEGb({\Tile_X7Y2_S2BEGb[7] ,
    \Tile_X7Y2_S2BEGb[6] ,
    \Tile_X7Y2_S2BEGb[5] ,
    \Tile_X7Y2_S2BEGb[4] ,
    \Tile_X7Y2_S2BEGb[3] ,
    \Tile_X7Y2_S2BEGb[2] ,
    \Tile_X7Y2_S2BEGb[1] ,
    \Tile_X7Y2_S2BEGb[0] }),
    .Tile_X0Y1_S4BEG({\Tile_X7Y2_S4BEG[15] ,
    \Tile_X7Y2_S4BEG[14] ,
    \Tile_X7Y2_S4BEG[13] ,
    \Tile_X7Y2_S4BEG[12] ,
    \Tile_X7Y2_S4BEG[11] ,
    \Tile_X7Y2_S4BEG[10] ,
    \Tile_X7Y2_S4BEG[9] ,
    \Tile_X7Y2_S4BEG[8] ,
    \Tile_X7Y2_S4BEG[7] ,
    \Tile_X7Y2_S4BEG[6] ,
    \Tile_X7Y2_S4BEG[5] ,
    \Tile_X7Y2_S4BEG[4] ,
    \Tile_X7Y2_S4BEG[3] ,
    \Tile_X7Y2_S4BEG[2] ,
    \Tile_X7Y2_S4BEG[1] ,
    \Tile_X7Y2_S4BEG[0] }),
    .Tile_X0Y1_SS4BEG({\Tile_X7Y2_SS4BEG[15] ,
    \Tile_X7Y2_SS4BEG[14] ,
    \Tile_X7Y2_SS4BEG[13] ,
    \Tile_X7Y2_SS4BEG[12] ,
    \Tile_X7Y2_SS4BEG[11] ,
    \Tile_X7Y2_SS4BEG[10] ,
    \Tile_X7Y2_SS4BEG[9] ,
    \Tile_X7Y2_SS4BEG[8] ,
    \Tile_X7Y2_SS4BEG[7] ,
    \Tile_X7Y2_SS4BEG[6] ,
    \Tile_X7Y2_SS4BEG[5] ,
    \Tile_X7Y2_SS4BEG[4] ,
    \Tile_X7Y2_SS4BEG[3] ,
    \Tile_X7Y2_SS4BEG[2] ,
    \Tile_X7Y2_SS4BEG[1] ,
    \Tile_X7Y2_SS4BEG[0] }),
    .Tile_X0Y1_W1BEG({\Tile_X7Y2_W1BEG[3] ,
    \Tile_X7Y2_W1BEG[2] ,
    \Tile_X7Y2_W1BEG[1] ,
    \Tile_X7Y2_W1BEG[0] }),
    .Tile_X0Y1_W1END({\Tile_X8Y2_W1BEG[3] ,
    \Tile_X8Y2_W1BEG[2] ,
    \Tile_X8Y2_W1BEG[1] ,
    \Tile_X8Y2_W1BEG[0] }),
    .Tile_X0Y1_W2BEG({\Tile_X7Y2_W2BEG[7] ,
    \Tile_X7Y2_W2BEG[6] ,
    \Tile_X7Y2_W2BEG[5] ,
    \Tile_X7Y2_W2BEG[4] ,
    \Tile_X7Y2_W2BEG[3] ,
    \Tile_X7Y2_W2BEG[2] ,
    \Tile_X7Y2_W2BEG[1] ,
    \Tile_X7Y2_W2BEG[0] }),
    .Tile_X0Y1_W2BEGb({\Tile_X7Y2_W2BEGb[7] ,
    \Tile_X7Y2_W2BEGb[6] ,
    \Tile_X7Y2_W2BEGb[5] ,
    \Tile_X7Y2_W2BEGb[4] ,
    \Tile_X7Y2_W2BEGb[3] ,
    \Tile_X7Y2_W2BEGb[2] ,
    \Tile_X7Y2_W2BEGb[1] ,
    \Tile_X7Y2_W2BEGb[0] }),
    .Tile_X0Y1_W2END({\Tile_X8Y2_W2BEGb[7] ,
    \Tile_X8Y2_W2BEGb[6] ,
    \Tile_X8Y2_W2BEGb[5] ,
    \Tile_X8Y2_W2BEGb[4] ,
    \Tile_X8Y2_W2BEGb[3] ,
    \Tile_X8Y2_W2BEGb[2] ,
    \Tile_X8Y2_W2BEGb[1] ,
    \Tile_X8Y2_W2BEGb[0] }),
    .Tile_X0Y1_W2MID({\Tile_X8Y2_W2BEG[7] ,
    \Tile_X8Y2_W2BEG[6] ,
    \Tile_X8Y2_W2BEG[5] ,
    \Tile_X8Y2_W2BEG[4] ,
    \Tile_X8Y2_W2BEG[3] ,
    \Tile_X8Y2_W2BEG[2] ,
    \Tile_X8Y2_W2BEG[1] ,
    \Tile_X8Y2_W2BEG[0] }),
    .Tile_X0Y1_W6BEG({\Tile_X7Y2_W6BEG[11] ,
    \Tile_X7Y2_W6BEG[10] ,
    \Tile_X7Y2_W6BEG[9] ,
    \Tile_X7Y2_W6BEG[8] ,
    \Tile_X7Y2_W6BEG[7] ,
    \Tile_X7Y2_W6BEG[6] ,
    \Tile_X7Y2_W6BEG[5] ,
    \Tile_X7Y2_W6BEG[4] ,
    \Tile_X7Y2_W6BEG[3] ,
    \Tile_X7Y2_W6BEG[2] ,
    \Tile_X7Y2_W6BEG[1] ,
    \Tile_X7Y2_W6BEG[0] }),
    .Tile_X0Y1_W6END({\Tile_X8Y2_W6BEG[11] ,
    \Tile_X8Y2_W6BEG[10] ,
    \Tile_X8Y2_W6BEG[9] ,
    \Tile_X8Y2_W6BEG[8] ,
    \Tile_X8Y2_W6BEG[7] ,
    \Tile_X8Y2_W6BEG[6] ,
    \Tile_X8Y2_W6BEG[5] ,
    \Tile_X8Y2_W6BEG[4] ,
    \Tile_X8Y2_W6BEG[3] ,
    \Tile_X8Y2_W6BEG[2] ,
    \Tile_X8Y2_W6BEG[1] ,
    \Tile_X8Y2_W6BEG[0] }),
    .Tile_X0Y1_WW4BEG({\Tile_X7Y2_WW4BEG[15] ,
    \Tile_X7Y2_WW4BEG[14] ,
    \Tile_X7Y2_WW4BEG[13] ,
    \Tile_X7Y2_WW4BEG[12] ,
    \Tile_X7Y2_WW4BEG[11] ,
    \Tile_X7Y2_WW4BEG[10] ,
    \Tile_X7Y2_WW4BEG[9] ,
    \Tile_X7Y2_WW4BEG[8] ,
    \Tile_X7Y2_WW4BEG[7] ,
    \Tile_X7Y2_WW4BEG[6] ,
    \Tile_X7Y2_WW4BEG[5] ,
    \Tile_X7Y2_WW4BEG[4] ,
    \Tile_X7Y2_WW4BEG[3] ,
    \Tile_X7Y2_WW4BEG[2] ,
    \Tile_X7Y2_WW4BEG[1] ,
    \Tile_X7Y2_WW4BEG[0] }),
    .Tile_X0Y1_WW4END({\Tile_X8Y2_WW4BEG[15] ,
    \Tile_X8Y2_WW4BEG[14] ,
    \Tile_X8Y2_WW4BEG[13] ,
    \Tile_X8Y2_WW4BEG[12] ,
    \Tile_X8Y2_WW4BEG[11] ,
    \Tile_X8Y2_WW4BEG[10] ,
    \Tile_X8Y2_WW4BEG[9] ,
    \Tile_X8Y2_WW4BEG[8] ,
    \Tile_X8Y2_WW4BEG[7] ,
    \Tile_X8Y2_WW4BEG[6] ,
    \Tile_X8Y2_WW4BEG[5] ,
    \Tile_X8Y2_WW4BEG[4] ,
    \Tile_X8Y2_WW4BEG[3] ,
    \Tile_X8Y2_WW4BEG[2] ,
    \Tile_X8Y2_WW4BEG[1] ,
    \Tile_X8Y2_WW4BEG[0] }));
 DSP Tile_X7Y3_DSP (.Tile_X0Y0_UserCLKo(Tile_X7Y3_UserCLKo),
    .Tile_X0Y1_UserCLK(Tile_X7Y5_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .Tile_X0Y0_E1BEG({\Tile_X7Y3_E1BEG[3] ,
    \Tile_X7Y3_E1BEG[2] ,
    \Tile_X7Y3_E1BEG[1] ,
    \Tile_X7Y3_E1BEG[0] }),
    .Tile_X0Y0_E1END({\Tile_X6Y3_E1BEG[3] ,
    \Tile_X6Y3_E1BEG[2] ,
    \Tile_X6Y3_E1BEG[1] ,
    \Tile_X6Y3_E1BEG[0] }),
    .Tile_X0Y0_E2BEG({\Tile_X7Y3_E2BEG[7] ,
    \Tile_X7Y3_E2BEG[6] ,
    \Tile_X7Y3_E2BEG[5] ,
    \Tile_X7Y3_E2BEG[4] ,
    \Tile_X7Y3_E2BEG[3] ,
    \Tile_X7Y3_E2BEG[2] ,
    \Tile_X7Y3_E2BEG[1] ,
    \Tile_X7Y3_E2BEG[0] }),
    .Tile_X0Y0_E2BEGb({\Tile_X7Y3_E2BEGb[7] ,
    \Tile_X7Y3_E2BEGb[6] ,
    \Tile_X7Y3_E2BEGb[5] ,
    \Tile_X7Y3_E2BEGb[4] ,
    \Tile_X7Y3_E2BEGb[3] ,
    \Tile_X7Y3_E2BEGb[2] ,
    \Tile_X7Y3_E2BEGb[1] ,
    \Tile_X7Y3_E2BEGb[0] }),
    .Tile_X0Y0_E2END({\Tile_X6Y3_E2BEGb[7] ,
    \Tile_X6Y3_E2BEGb[6] ,
    \Tile_X6Y3_E2BEGb[5] ,
    \Tile_X6Y3_E2BEGb[4] ,
    \Tile_X6Y3_E2BEGb[3] ,
    \Tile_X6Y3_E2BEGb[2] ,
    \Tile_X6Y3_E2BEGb[1] ,
    \Tile_X6Y3_E2BEGb[0] }),
    .Tile_X0Y0_E2MID({\Tile_X6Y3_E2BEG[7] ,
    \Tile_X6Y3_E2BEG[6] ,
    \Tile_X6Y3_E2BEG[5] ,
    \Tile_X6Y3_E2BEG[4] ,
    \Tile_X6Y3_E2BEG[3] ,
    \Tile_X6Y3_E2BEG[2] ,
    \Tile_X6Y3_E2BEG[1] ,
    \Tile_X6Y3_E2BEG[0] }),
    .Tile_X0Y0_E6BEG({\Tile_X7Y3_E6BEG[11] ,
    \Tile_X7Y3_E6BEG[10] ,
    \Tile_X7Y3_E6BEG[9] ,
    \Tile_X7Y3_E6BEG[8] ,
    \Tile_X7Y3_E6BEG[7] ,
    \Tile_X7Y3_E6BEG[6] ,
    \Tile_X7Y3_E6BEG[5] ,
    \Tile_X7Y3_E6BEG[4] ,
    \Tile_X7Y3_E6BEG[3] ,
    \Tile_X7Y3_E6BEG[2] ,
    \Tile_X7Y3_E6BEG[1] ,
    \Tile_X7Y3_E6BEG[0] }),
    .Tile_X0Y0_E6END({\Tile_X6Y3_E6BEG[11] ,
    \Tile_X6Y3_E6BEG[10] ,
    \Tile_X6Y3_E6BEG[9] ,
    \Tile_X6Y3_E6BEG[8] ,
    \Tile_X6Y3_E6BEG[7] ,
    \Tile_X6Y3_E6BEG[6] ,
    \Tile_X6Y3_E6BEG[5] ,
    \Tile_X6Y3_E6BEG[4] ,
    \Tile_X6Y3_E6BEG[3] ,
    \Tile_X6Y3_E6BEG[2] ,
    \Tile_X6Y3_E6BEG[1] ,
    \Tile_X6Y3_E6BEG[0] }),
    .Tile_X0Y0_EE4BEG({\Tile_X7Y3_EE4BEG[15] ,
    \Tile_X7Y3_EE4BEG[14] ,
    \Tile_X7Y3_EE4BEG[13] ,
    \Tile_X7Y3_EE4BEG[12] ,
    \Tile_X7Y3_EE4BEG[11] ,
    \Tile_X7Y3_EE4BEG[10] ,
    \Tile_X7Y3_EE4BEG[9] ,
    \Tile_X7Y3_EE4BEG[8] ,
    \Tile_X7Y3_EE4BEG[7] ,
    \Tile_X7Y3_EE4BEG[6] ,
    \Tile_X7Y3_EE4BEG[5] ,
    \Tile_X7Y3_EE4BEG[4] ,
    \Tile_X7Y3_EE4BEG[3] ,
    \Tile_X7Y3_EE4BEG[2] ,
    \Tile_X7Y3_EE4BEG[1] ,
    \Tile_X7Y3_EE4BEG[0] }),
    .Tile_X0Y0_EE4END({\Tile_X6Y3_EE4BEG[15] ,
    \Tile_X6Y3_EE4BEG[14] ,
    \Tile_X6Y3_EE4BEG[13] ,
    \Tile_X6Y3_EE4BEG[12] ,
    \Tile_X6Y3_EE4BEG[11] ,
    \Tile_X6Y3_EE4BEG[10] ,
    \Tile_X6Y3_EE4BEG[9] ,
    \Tile_X6Y3_EE4BEG[8] ,
    \Tile_X6Y3_EE4BEG[7] ,
    \Tile_X6Y3_EE4BEG[6] ,
    \Tile_X6Y3_EE4BEG[5] ,
    \Tile_X6Y3_EE4BEG[4] ,
    \Tile_X6Y3_EE4BEG[3] ,
    \Tile_X6Y3_EE4BEG[2] ,
    \Tile_X6Y3_EE4BEG[1] ,
    \Tile_X6Y3_EE4BEG[0] }),
    .Tile_X0Y0_FrameData({\Tile_X6Y3_FrameData_O[31] ,
    \Tile_X6Y3_FrameData_O[30] ,
    \Tile_X6Y3_FrameData_O[29] ,
    \Tile_X6Y3_FrameData_O[28] ,
    \Tile_X6Y3_FrameData_O[27] ,
    \Tile_X6Y3_FrameData_O[26] ,
    \Tile_X6Y3_FrameData_O[25] ,
    \Tile_X6Y3_FrameData_O[24] ,
    \Tile_X6Y3_FrameData_O[23] ,
    \Tile_X6Y3_FrameData_O[22] ,
    \Tile_X6Y3_FrameData_O[21] ,
    \Tile_X6Y3_FrameData_O[20] ,
    \Tile_X6Y3_FrameData_O[19] ,
    \Tile_X6Y3_FrameData_O[18] ,
    \Tile_X6Y3_FrameData_O[17] ,
    \Tile_X6Y3_FrameData_O[16] ,
    \Tile_X6Y3_FrameData_O[15] ,
    \Tile_X6Y3_FrameData_O[14] ,
    \Tile_X6Y3_FrameData_O[13] ,
    \Tile_X6Y3_FrameData_O[12] ,
    \Tile_X6Y3_FrameData_O[11] ,
    \Tile_X6Y3_FrameData_O[10] ,
    \Tile_X6Y3_FrameData_O[9] ,
    \Tile_X6Y3_FrameData_O[8] ,
    \Tile_X6Y3_FrameData_O[7] ,
    \Tile_X6Y3_FrameData_O[6] ,
    \Tile_X6Y3_FrameData_O[5] ,
    \Tile_X6Y3_FrameData_O[4] ,
    \Tile_X6Y3_FrameData_O[3] ,
    \Tile_X6Y3_FrameData_O[2] ,
    \Tile_X6Y3_FrameData_O[1] ,
    \Tile_X6Y3_FrameData_O[0] }),
    .Tile_X0Y0_FrameData_O({\Tile_X7Y3_FrameData_O[31] ,
    \Tile_X7Y3_FrameData_O[30] ,
    \Tile_X7Y3_FrameData_O[29] ,
    \Tile_X7Y3_FrameData_O[28] ,
    \Tile_X7Y3_FrameData_O[27] ,
    \Tile_X7Y3_FrameData_O[26] ,
    \Tile_X7Y3_FrameData_O[25] ,
    \Tile_X7Y3_FrameData_O[24] ,
    \Tile_X7Y3_FrameData_O[23] ,
    \Tile_X7Y3_FrameData_O[22] ,
    \Tile_X7Y3_FrameData_O[21] ,
    \Tile_X7Y3_FrameData_O[20] ,
    \Tile_X7Y3_FrameData_O[19] ,
    \Tile_X7Y3_FrameData_O[18] ,
    \Tile_X7Y3_FrameData_O[17] ,
    \Tile_X7Y3_FrameData_O[16] ,
    \Tile_X7Y3_FrameData_O[15] ,
    \Tile_X7Y3_FrameData_O[14] ,
    \Tile_X7Y3_FrameData_O[13] ,
    \Tile_X7Y3_FrameData_O[12] ,
    \Tile_X7Y3_FrameData_O[11] ,
    \Tile_X7Y3_FrameData_O[10] ,
    \Tile_X7Y3_FrameData_O[9] ,
    \Tile_X7Y3_FrameData_O[8] ,
    \Tile_X7Y3_FrameData_O[7] ,
    \Tile_X7Y3_FrameData_O[6] ,
    \Tile_X7Y3_FrameData_O[5] ,
    \Tile_X7Y3_FrameData_O[4] ,
    \Tile_X7Y3_FrameData_O[3] ,
    \Tile_X7Y3_FrameData_O[2] ,
    \Tile_X7Y3_FrameData_O[1] ,
    \Tile_X7Y3_FrameData_O[0] }),
    .Tile_X0Y0_FrameStrobe_O({\Tile_X7Y3_FrameStrobe_O[19] ,
    \Tile_X7Y3_FrameStrobe_O[18] ,
    \Tile_X7Y3_FrameStrobe_O[17] ,
    \Tile_X7Y3_FrameStrobe_O[16] ,
    \Tile_X7Y3_FrameStrobe_O[15] ,
    \Tile_X7Y3_FrameStrobe_O[14] ,
    \Tile_X7Y3_FrameStrobe_O[13] ,
    \Tile_X7Y3_FrameStrobe_O[12] ,
    \Tile_X7Y3_FrameStrobe_O[11] ,
    \Tile_X7Y3_FrameStrobe_O[10] ,
    \Tile_X7Y3_FrameStrobe_O[9] ,
    \Tile_X7Y3_FrameStrobe_O[8] ,
    \Tile_X7Y3_FrameStrobe_O[7] ,
    \Tile_X7Y3_FrameStrobe_O[6] ,
    \Tile_X7Y3_FrameStrobe_O[5] ,
    \Tile_X7Y3_FrameStrobe_O[4] ,
    \Tile_X7Y3_FrameStrobe_O[3] ,
    \Tile_X7Y3_FrameStrobe_O[2] ,
    \Tile_X7Y3_FrameStrobe_O[1] ,
    \Tile_X7Y3_FrameStrobe_O[0] }),
    .Tile_X0Y0_N1BEG({\Tile_X7Y3_N1BEG[3] ,
    \Tile_X7Y3_N1BEG[2] ,
    \Tile_X7Y3_N1BEG[1] ,
    \Tile_X7Y3_N1BEG[0] }),
    .Tile_X0Y0_N2BEG({\Tile_X7Y3_N2BEG[7] ,
    \Tile_X7Y3_N2BEG[6] ,
    \Tile_X7Y3_N2BEG[5] ,
    \Tile_X7Y3_N2BEG[4] ,
    \Tile_X7Y3_N2BEG[3] ,
    \Tile_X7Y3_N2BEG[2] ,
    \Tile_X7Y3_N2BEG[1] ,
    \Tile_X7Y3_N2BEG[0] }),
    .Tile_X0Y0_N2BEGb({\Tile_X7Y3_N2BEGb[7] ,
    \Tile_X7Y3_N2BEGb[6] ,
    \Tile_X7Y3_N2BEGb[5] ,
    \Tile_X7Y3_N2BEGb[4] ,
    \Tile_X7Y3_N2BEGb[3] ,
    \Tile_X7Y3_N2BEGb[2] ,
    \Tile_X7Y3_N2BEGb[1] ,
    \Tile_X7Y3_N2BEGb[0] }),
    .Tile_X0Y0_N4BEG({\Tile_X7Y3_N4BEG[15] ,
    \Tile_X7Y3_N4BEG[14] ,
    \Tile_X7Y3_N4BEG[13] ,
    \Tile_X7Y3_N4BEG[12] ,
    \Tile_X7Y3_N4BEG[11] ,
    \Tile_X7Y3_N4BEG[10] ,
    \Tile_X7Y3_N4BEG[9] ,
    \Tile_X7Y3_N4BEG[8] ,
    \Tile_X7Y3_N4BEG[7] ,
    \Tile_X7Y3_N4BEG[6] ,
    \Tile_X7Y3_N4BEG[5] ,
    \Tile_X7Y3_N4BEG[4] ,
    \Tile_X7Y3_N4BEG[3] ,
    \Tile_X7Y3_N4BEG[2] ,
    \Tile_X7Y3_N4BEG[1] ,
    \Tile_X7Y3_N4BEG[0] }),
    .Tile_X0Y0_NN4BEG({\Tile_X7Y3_NN4BEG[15] ,
    \Tile_X7Y3_NN4BEG[14] ,
    \Tile_X7Y3_NN4BEG[13] ,
    \Tile_X7Y3_NN4BEG[12] ,
    \Tile_X7Y3_NN4BEG[11] ,
    \Tile_X7Y3_NN4BEG[10] ,
    \Tile_X7Y3_NN4BEG[9] ,
    \Tile_X7Y3_NN4BEG[8] ,
    \Tile_X7Y3_NN4BEG[7] ,
    \Tile_X7Y3_NN4BEG[6] ,
    \Tile_X7Y3_NN4BEG[5] ,
    \Tile_X7Y3_NN4BEG[4] ,
    \Tile_X7Y3_NN4BEG[3] ,
    \Tile_X7Y3_NN4BEG[2] ,
    \Tile_X7Y3_NN4BEG[1] ,
    \Tile_X7Y3_NN4BEG[0] }),
    .Tile_X0Y0_S1END({\Tile_X7Y2_S1BEG[3] ,
    \Tile_X7Y2_S1BEG[2] ,
    \Tile_X7Y2_S1BEG[1] ,
    \Tile_X7Y2_S1BEG[0] }),
    .Tile_X0Y0_S2END({\Tile_X7Y2_S2BEGb[7] ,
    \Tile_X7Y2_S2BEGb[6] ,
    \Tile_X7Y2_S2BEGb[5] ,
    \Tile_X7Y2_S2BEGb[4] ,
    \Tile_X7Y2_S2BEGb[3] ,
    \Tile_X7Y2_S2BEGb[2] ,
    \Tile_X7Y2_S2BEGb[1] ,
    \Tile_X7Y2_S2BEGb[0] }),
    .Tile_X0Y0_S2MID({\Tile_X7Y2_S2BEG[7] ,
    \Tile_X7Y2_S2BEG[6] ,
    \Tile_X7Y2_S2BEG[5] ,
    \Tile_X7Y2_S2BEG[4] ,
    \Tile_X7Y2_S2BEG[3] ,
    \Tile_X7Y2_S2BEG[2] ,
    \Tile_X7Y2_S2BEG[1] ,
    \Tile_X7Y2_S2BEG[0] }),
    .Tile_X0Y0_S4END({\Tile_X7Y2_S4BEG[15] ,
    \Tile_X7Y2_S4BEG[14] ,
    \Tile_X7Y2_S4BEG[13] ,
    \Tile_X7Y2_S4BEG[12] ,
    \Tile_X7Y2_S4BEG[11] ,
    \Tile_X7Y2_S4BEG[10] ,
    \Tile_X7Y2_S4BEG[9] ,
    \Tile_X7Y2_S4BEG[8] ,
    \Tile_X7Y2_S4BEG[7] ,
    \Tile_X7Y2_S4BEG[6] ,
    \Tile_X7Y2_S4BEG[5] ,
    \Tile_X7Y2_S4BEG[4] ,
    \Tile_X7Y2_S4BEG[3] ,
    \Tile_X7Y2_S4BEG[2] ,
    \Tile_X7Y2_S4BEG[1] ,
    \Tile_X7Y2_S4BEG[0] }),
    .Tile_X0Y0_SS4END({\Tile_X7Y2_SS4BEG[15] ,
    \Tile_X7Y2_SS4BEG[14] ,
    \Tile_X7Y2_SS4BEG[13] ,
    \Tile_X7Y2_SS4BEG[12] ,
    \Tile_X7Y2_SS4BEG[11] ,
    \Tile_X7Y2_SS4BEG[10] ,
    \Tile_X7Y2_SS4BEG[9] ,
    \Tile_X7Y2_SS4BEG[8] ,
    \Tile_X7Y2_SS4BEG[7] ,
    \Tile_X7Y2_SS4BEG[6] ,
    \Tile_X7Y2_SS4BEG[5] ,
    \Tile_X7Y2_SS4BEG[4] ,
    \Tile_X7Y2_SS4BEG[3] ,
    \Tile_X7Y2_SS4BEG[2] ,
    \Tile_X7Y2_SS4BEG[1] ,
    \Tile_X7Y2_SS4BEG[0] }),
    .Tile_X0Y0_W1BEG({\Tile_X7Y3_W1BEG[3] ,
    \Tile_X7Y3_W1BEG[2] ,
    \Tile_X7Y3_W1BEG[1] ,
    \Tile_X7Y3_W1BEG[0] }),
    .Tile_X0Y0_W1END({\Tile_X8Y3_W1BEG[3] ,
    \Tile_X8Y3_W1BEG[2] ,
    \Tile_X8Y3_W1BEG[1] ,
    \Tile_X8Y3_W1BEG[0] }),
    .Tile_X0Y0_W2BEG({\Tile_X7Y3_W2BEG[7] ,
    \Tile_X7Y3_W2BEG[6] ,
    \Tile_X7Y3_W2BEG[5] ,
    \Tile_X7Y3_W2BEG[4] ,
    \Tile_X7Y3_W2BEG[3] ,
    \Tile_X7Y3_W2BEG[2] ,
    \Tile_X7Y3_W2BEG[1] ,
    \Tile_X7Y3_W2BEG[0] }),
    .Tile_X0Y0_W2BEGb({\Tile_X7Y3_W2BEGb[7] ,
    \Tile_X7Y3_W2BEGb[6] ,
    \Tile_X7Y3_W2BEGb[5] ,
    \Tile_X7Y3_W2BEGb[4] ,
    \Tile_X7Y3_W2BEGb[3] ,
    \Tile_X7Y3_W2BEGb[2] ,
    \Tile_X7Y3_W2BEGb[1] ,
    \Tile_X7Y3_W2BEGb[0] }),
    .Tile_X0Y0_W2END({\Tile_X8Y3_W2BEGb[7] ,
    \Tile_X8Y3_W2BEGb[6] ,
    \Tile_X8Y3_W2BEGb[5] ,
    \Tile_X8Y3_W2BEGb[4] ,
    \Tile_X8Y3_W2BEGb[3] ,
    \Tile_X8Y3_W2BEGb[2] ,
    \Tile_X8Y3_W2BEGb[1] ,
    \Tile_X8Y3_W2BEGb[0] }),
    .Tile_X0Y0_W2MID({\Tile_X8Y3_W2BEG[7] ,
    \Tile_X8Y3_W2BEG[6] ,
    \Tile_X8Y3_W2BEG[5] ,
    \Tile_X8Y3_W2BEG[4] ,
    \Tile_X8Y3_W2BEG[3] ,
    \Tile_X8Y3_W2BEG[2] ,
    \Tile_X8Y3_W2BEG[1] ,
    \Tile_X8Y3_W2BEG[0] }),
    .Tile_X0Y0_W6BEG({\Tile_X7Y3_W6BEG[11] ,
    \Tile_X7Y3_W6BEG[10] ,
    \Tile_X7Y3_W6BEG[9] ,
    \Tile_X7Y3_W6BEG[8] ,
    \Tile_X7Y3_W6BEG[7] ,
    \Tile_X7Y3_W6BEG[6] ,
    \Tile_X7Y3_W6BEG[5] ,
    \Tile_X7Y3_W6BEG[4] ,
    \Tile_X7Y3_W6BEG[3] ,
    \Tile_X7Y3_W6BEG[2] ,
    \Tile_X7Y3_W6BEG[1] ,
    \Tile_X7Y3_W6BEG[0] }),
    .Tile_X0Y0_W6END({\Tile_X8Y3_W6BEG[11] ,
    \Tile_X8Y3_W6BEG[10] ,
    \Tile_X8Y3_W6BEG[9] ,
    \Tile_X8Y3_W6BEG[8] ,
    \Tile_X8Y3_W6BEG[7] ,
    \Tile_X8Y3_W6BEG[6] ,
    \Tile_X8Y3_W6BEG[5] ,
    \Tile_X8Y3_W6BEG[4] ,
    \Tile_X8Y3_W6BEG[3] ,
    \Tile_X8Y3_W6BEG[2] ,
    \Tile_X8Y3_W6BEG[1] ,
    \Tile_X8Y3_W6BEG[0] }),
    .Tile_X0Y0_WW4BEG({\Tile_X7Y3_WW4BEG[15] ,
    \Tile_X7Y3_WW4BEG[14] ,
    \Tile_X7Y3_WW4BEG[13] ,
    \Tile_X7Y3_WW4BEG[12] ,
    \Tile_X7Y3_WW4BEG[11] ,
    \Tile_X7Y3_WW4BEG[10] ,
    \Tile_X7Y3_WW4BEG[9] ,
    \Tile_X7Y3_WW4BEG[8] ,
    \Tile_X7Y3_WW4BEG[7] ,
    \Tile_X7Y3_WW4BEG[6] ,
    \Tile_X7Y3_WW4BEG[5] ,
    \Tile_X7Y3_WW4BEG[4] ,
    \Tile_X7Y3_WW4BEG[3] ,
    \Tile_X7Y3_WW4BEG[2] ,
    \Tile_X7Y3_WW4BEG[1] ,
    \Tile_X7Y3_WW4BEG[0] }),
    .Tile_X0Y0_WW4END({\Tile_X8Y3_WW4BEG[15] ,
    \Tile_X8Y3_WW4BEG[14] ,
    \Tile_X8Y3_WW4BEG[13] ,
    \Tile_X8Y3_WW4BEG[12] ,
    \Tile_X8Y3_WW4BEG[11] ,
    \Tile_X8Y3_WW4BEG[10] ,
    \Tile_X8Y3_WW4BEG[9] ,
    \Tile_X8Y3_WW4BEG[8] ,
    \Tile_X8Y3_WW4BEG[7] ,
    \Tile_X8Y3_WW4BEG[6] ,
    \Tile_X8Y3_WW4BEG[5] ,
    \Tile_X8Y3_WW4BEG[4] ,
    \Tile_X8Y3_WW4BEG[3] ,
    \Tile_X8Y3_WW4BEG[2] ,
    \Tile_X8Y3_WW4BEG[1] ,
    \Tile_X8Y3_WW4BEG[0] }),
    .Tile_X0Y1_E1BEG({\Tile_X7Y4_E1BEG[3] ,
    \Tile_X7Y4_E1BEG[2] ,
    \Tile_X7Y4_E1BEG[1] ,
    \Tile_X7Y4_E1BEG[0] }),
    .Tile_X0Y1_E1END({\Tile_X6Y4_E1BEG[3] ,
    \Tile_X6Y4_E1BEG[2] ,
    \Tile_X6Y4_E1BEG[1] ,
    \Tile_X6Y4_E1BEG[0] }),
    .Tile_X0Y1_E2BEG({\Tile_X7Y4_E2BEG[7] ,
    \Tile_X7Y4_E2BEG[6] ,
    \Tile_X7Y4_E2BEG[5] ,
    \Tile_X7Y4_E2BEG[4] ,
    \Tile_X7Y4_E2BEG[3] ,
    \Tile_X7Y4_E2BEG[2] ,
    \Tile_X7Y4_E2BEG[1] ,
    \Tile_X7Y4_E2BEG[0] }),
    .Tile_X0Y1_E2BEGb({\Tile_X7Y4_E2BEGb[7] ,
    \Tile_X7Y4_E2BEGb[6] ,
    \Tile_X7Y4_E2BEGb[5] ,
    \Tile_X7Y4_E2BEGb[4] ,
    \Tile_X7Y4_E2BEGb[3] ,
    \Tile_X7Y4_E2BEGb[2] ,
    \Tile_X7Y4_E2BEGb[1] ,
    \Tile_X7Y4_E2BEGb[0] }),
    .Tile_X0Y1_E2END({\Tile_X6Y4_E2BEGb[7] ,
    \Tile_X6Y4_E2BEGb[6] ,
    \Tile_X6Y4_E2BEGb[5] ,
    \Tile_X6Y4_E2BEGb[4] ,
    \Tile_X6Y4_E2BEGb[3] ,
    \Tile_X6Y4_E2BEGb[2] ,
    \Tile_X6Y4_E2BEGb[1] ,
    \Tile_X6Y4_E2BEGb[0] }),
    .Tile_X0Y1_E2MID({\Tile_X6Y4_E2BEG[7] ,
    \Tile_X6Y4_E2BEG[6] ,
    \Tile_X6Y4_E2BEG[5] ,
    \Tile_X6Y4_E2BEG[4] ,
    \Tile_X6Y4_E2BEG[3] ,
    \Tile_X6Y4_E2BEG[2] ,
    \Tile_X6Y4_E2BEG[1] ,
    \Tile_X6Y4_E2BEG[0] }),
    .Tile_X0Y1_E6BEG({\Tile_X7Y4_E6BEG[11] ,
    \Tile_X7Y4_E6BEG[10] ,
    \Tile_X7Y4_E6BEG[9] ,
    \Tile_X7Y4_E6BEG[8] ,
    \Tile_X7Y4_E6BEG[7] ,
    \Tile_X7Y4_E6BEG[6] ,
    \Tile_X7Y4_E6BEG[5] ,
    \Tile_X7Y4_E6BEG[4] ,
    \Tile_X7Y4_E6BEG[3] ,
    \Tile_X7Y4_E6BEG[2] ,
    \Tile_X7Y4_E6BEG[1] ,
    \Tile_X7Y4_E6BEG[0] }),
    .Tile_X0Y1_E6END({\Tile_X6Y4_E6BEG[11] ,
    \Tile_X6Y4_E6BEG[10] ,
    \Tile_X6Y4_E6BEG[9] ,
    \Tile_X6Y4_E6BEG[8] ,
    \Tile_X6Y4_E6BEG[7] ,
    \Tile_X6Y4_E6BEG[6] ,
    \Tile_X6Y4_E6BEG[5] ,
    \Tile_X6Y4_E6BEG[4] ,
    \Tile_X6Y4_E6BEG[3] ,
    \Tile_X6Y4_E6BEG[2] ,
    \Tile_X6Y4_E6BEG[1] ,
    \Tile_X6Y4_E6BEG[0] }),
    .Tile_X0Y1_EE4BEG({\Tile_X7Y4_EE4BEG[15] ,
    \Tile_X7Y4_EE4BEG[14] ,
    \Tile_X7Y4_EE4BEG[13] ,
    \Tile_X7Y4_EE4BEG[12] ,
    \Tile_X7Y4_EE4BEG[11] ,
    \Tile_X7Y4_EE4BEG[10] ,
    \Tile_X7Y4_EE4BEG[9] ,
    \Tile_X7Y4_EE4BEG[8] ,
    \Tile_X7Y4_EE4BEG[7] ,
    \Tile_X7Y4_EE4BEG[6] ,
    \Tile_X7Y4_EE4BEG[5] ,
    \Tile_X7Y4_EE4BEG[4] ,
    \Tile_X7Y4_EE4BEG[3] ,
    \Tile_X7Y4_EE4BEG[2] ,
    \Tile_X7Y4_EE4BEG[1] ,
    \Tile_X7Y4_EE4BEG[0] }),
    .Tile_X0Y1_EE4END({\Tile_X6Y4_EE4BEG[15] ,
    \Tile_X6Y4_EE4BEG[14] ,
    \Tile_X6Y4_EE4BEG[13] ,
    \Tile_X6Y4_EE4BEG[12] ,
    \Tile_X6Y4_EE4BEG[11] ,
    \Tile_X6Y4_EE4BEG[10] ,
    \Tile_X6Y4_EE4BEG[9] ,
    \Tile_X6Y4_EE4BEG[8] ,
    \Tile_X6Y4_EE4BEG[7] ,
    \Tile_X6Y4_EE4BEG[6] ,
    \Tile_X6Y4_EE4BEG[5] ,
    \Tile_X6Y4_EE4BEG[4] ,
    \Tile_X6Y4_EE4BEG[3] ,
    \Tile_X6Y4_EE4BEG[2] ,
    \Tile_X6Y4_EE4BEG[1] ,
    \Tile_X6Y4_EE4BEG[0] }),
    .Tile_X0Y1_FrameData({\Tile_X6Y4_FrameData_O[31] ,
    \Tile_X6Y4_FrameData_O[30] ,
    \Tile_X6Y4_FrameData_O[29] ,
    \Tile_X6Y4_FrameData_O[28] ,
    \Tile_X6Y4_FrameData_O[27] ,
    \Tile_X6Y4_FrameData_O[26] ,
    \Tile_X6Y4_FrameData_O[25] ,
    \Tile_X6Y4_FrameData_O[24] ,
    \Tile_X6Y4_FrameData_O[23] ,
    \Tile_X6Y4_FrameData_O[22] ,
    \Tile_X6Y4_FrameData_O[21] ,
    \Tile_X6Y4_FrameData_O[20] ,
    \Tile_X6Y4_FrameData_O[19] ,
    \Tile_X6Y4_FrameData_O[18] ,
    \Tile_X6Y4_FrameData_O[17] ,
    \Tile_X6Y4_FrameData_O[16] ,
    \Tile_X6Y4_FrameData_O[15] ,
    \Tile_X6Y4_FrameData_O[14] ,
    \Tile_X6Y4_FrameData_O[13] ,
    \Tile_X6Y4_FrameData_O[12] ,
    \Tile_X6Y4_FrameData_O[11] ,
    \Tile_X6Y4_FrameData_O[10] ,
    \Tile_X6Y4_FrameData_O[9] ,
    \Tile_X6Y4_FrameData_O[8] ,
    \Tile_X6Y4_FrameData_O[7] ,
    \Tile_X6Y4_FrameData_O[6] ,
    \Tile_X6Y4_FrameData_O[5] ,
    \Tile_X6Y4_FrameData_O[4] ,
    \Tile_X6Y4_FrameData_O[3] ,
    \Tile_X6Y4_FrameData_O[2] ,
    \Tile_X6Y4_FrameData_O[1] ,
    \Tile_X6Y4_FrameData_O[0] }),
    .Tile_X0Y1_FrameData_O({\Tile_X7Y4_FrameData_O[31] ,
    \Tile_X7Y4_FrameData_O[30] ,
    \Tile_X7Y4_FrameData_O[29] ,
    \Tile_X7Y4_FrameData_O[28] ,
    \Tile_X7Y4_FrameData_O[27] ,
    \Tile_X7Y4_FrameData_O[26] ,
    \Tile_X7Y4_FrameData_O[25] ,
    \Tile_X7Y4_FrameData_O[24] ,
    \Tile_X7Y4_FrameData_O[23] ,
    \Tile_X7Y4_FrameData_O[22] ,
    \Tile_X7Y4_FrameData_O[21] ,
    \Tile_X7Y4_FrameData_O[20] ,
    \Tile_X7Y4_FrameData_O[19] ,
    \Tile_X7Y4_FrameData_O[18] ,
    \Tile_X7Y4_FrameData_O[17] ,
    \Tile_X7Y4_FrameData_O[16] ,
    \Tile_X7Y4_FrameData_O[15] ,
    \Tile_X7Y4_FrameData_O[14] ,
    \Tile_X7Y4_FrameData_O[13] ,
    \Tile_X7Y4_FrameData_O[12] ,
    \Tile_X7Y4_FrameData_O[11] ,
    \Tile_X7Y4_FrameData_O[10] ,
    \Tile_X7Y4_FrameData_O[9] ,
    \Tile_X7Y4_FrameData_O[8] ,
    \Tile_X7Y4_FrameData_O[7] ,
    \Tile_X7Y4_FrameData_O[6] ,
    \Tile_X7Y4_FrameData_O[5] ,
    \Tile_X7Y4_FrameData_O[4] ,
    \Tile_X7Y4_FrameData_O[3] ,
    \Tile_X7Y4_FrameData_O[2] ,
    \Tile_X7Y4_FrameData_O[1] ,
    \Tile_X7Y4_FrameData_O[0] }),
    .Tile_X0Y1_FrameStrobe({\Tile_X7Y5_FrameStrobe_O[19] ,
    \Tile_X7Y5_FrameStrobe_O[18] ,
    \Tile_X7Y5_FrameStrobe_O[17] ,
    \Tile_X7Y5_FrameStrobe_O[16] ,
    \Tile_X7Y5_FrameStrobe_O[15] ,
    \Tile_X7Y5_FrameStrobe_O[14] ,
    \Tile_X7Y5_FrameStrobe_O[13] ,
    \Tile_X7Y5_FrameStrobe_O[12] ,
    \Tile_X7Y5_FrameStrobe_O[11] ,
    \Tile_X7Y5_FrameStrobe_O[10] ,
    \Tile_X7Y5_FrameStrobe_O[9] ,
    \Tile_X7Y5_FrameStrobe_O[8] ,
    \Tile_X7Y5_FrameStrobe_O[7] ,
    \Tile_X7Y5_FrameStrobe_O[6] ,
    \Tile_X7Y5_FrameStrobe_O[5] ,
    \Tile_X7Y5_FrameStrobe_O[4] ,
    \Tile_X7Y5_FrameStrobe_O[3] ,
    \Tile_X7Y5_FrameStrobe_O[2] ,
    \Tile_X7Y5_FrameStrobe_O[1] ,
    \Tile_X7Y5_FrameStrobe_O[0] }),
    .Tile_X0Y1_N1END({\Tile_X7Y5_N1BEG[3] ,
    \Tile_X7Y5_N1BEG[2] ,
    \Tile_X7Y5_N1BEG[1] ,
    \Tile_X7Y5_N1BEG[0] }),
    .Tile_X0Y1_N2END({\Tile_X7Y5_N2BEGb[7] ,
    \Tile_X7Y5_N2BEGb[6] ,
    \Tile_X7Y5_N2BEGb[5] ,
    \Tile_X7Y5_N2BEGb[4] ,
    \Tile_X7Y5_N2BEGb[3] ,
    \Tile_X7Y5_N2BEGb[2] ,
    \Tile_X7Y5_N2BEGb[1] ,
    \Tile_X7Y5_N2BEGb[0] }),
    .Tile_X0Y1_N2MID({\Tile_X7Y5_N2BEG[7] ,
    \Tile_X7Y5_N2BEG[6] ,
    \Tile_X7Y5_N2BEG[5] ,
    \Tile_X7Y5_N2BEG[4] ,
    \Tile_X7Y5_N2BEG[3] ,
    \Tile_X7Y5_N2BEG[2] ,
    \Tile_X7Y5_N2BEG[1] ,
    \Tile_X7Y5_N2BEG[0] }),
    .Tile_X0Y1_N4END({\Tile_X7Y5_N4BEG[15] ,
    \Tile_X7Y5_N4BEG[14] ,
    \Tile_X7Y5_N4BEG[13] ,
    \Tile_X7Y5_N4BEG[12] ,
    \Tile_X7Y5_N4BEG[11] ,
    \Tile_X7Y5_N4BEG[10] ,
    \Tile_X7Y5_N4BEG[9] ,
    \Tile_X7Y5_N4BEG[8] ,
    \Tile_X7Y5_N4BEG[7] ,
    \Tile_X7Y5_N4BEG[6] ,
    \Tile_X7Y5_N4BEG[5] ,
    \Tile_X7Y5_N4BEG[4] ,
    \Tile_X7Y5_N4BEG[3] ,
    \Tile_X7Y5_N4BEG[2] ,
    \Tile_X7Y5_N4BEG[1] ,
    \Tile_X7Y5_N4BEG[0] }),
    .Tile_X0Y1_NN4END({\Tile_X7Y5_NN4BEG[15] ,
    \Tile_X7Y5_NN4BEG[14] ,
    \Tile_X7Y5_NN4BEG[13] ,
    \Tile_X7Y5_NN4BEG[12] ,
    \Tile_X7Y5_NN4BEG[11] ,
    \Tile_X7Y5_NN4BEG[10] ,
    \Tile_X7Y5_NN4BEG[9] ,
    \Tile_X7Y5_NN4BEG[8] ,
    \Tile_X7Y5_NN4BEG[7] ,
    \Tile_X7Y5_NN4BEG[6] ,
    \Tile_X7Y5_NN4BEG[5] ,
    \Tile_X7Y5_NN4BEG[4] ,
    \Tile_X7Y5_NN4BEG[3] ,
    \Tile_X7Y5_NN4BEG[2] ,
    \Tile_X7Y5_NN4BEG[1] ,
    \Tile_X7Y5_NN4BEG[0] }),
    .Tile_X0Y1_S1BEG({\Tile_X7Y4_S1BEG[3] ,
    \Tile_X7Y4_S1BEG[2] ,
    \Tile_X7Y4_S1BEG[1] ,
    \Tile_X7Y4_S1BEG[0] }),
    .Tile_X0Y1_S2BEG({\Tile_X7Y4_S2BEG[7] ,
    \Tile_X7Y4_S2BEG[6] ,
    \Tile_X7Y4_S2BEG[5] ,
    \Tile_X7Y4_S2BEG[4] ,
    \Tile_X7Y4_S2BEG[3] ,
    \Tile_X7Y4_S2BEG[2] ,
    \Tile_X7Y4_S2BEG[1] ,
    \Tile_X7Y4_S2BEG[0] }),
    .Tile_X0Y1_S2BEGb({\Tile_X7Y4_S2BEGb[7] ,
    \Tile_X7Y4_S2BEGb[6] ,
    \Tile_X7Y4_S2BEGb[5] ,
    \Tile_X7Y4_S2BEGb[4] ,
    \Tile_X7Y4_S2BEGb[3] ,
    \Tile_X7Y4_S2BEGb[2] ,
    \Tile_X7Y4_S2BEGb[1] ,
    \Tile_X7Y4_S2BEGb[0] }),
    .Tile_X0Y1_S4BEG({\Tile_X7Y4_S4BEG[15] ,
    \Tile_X7Y4_S4BEG[14] ,
    \Tile_X7Y4_S4BEG[13] ,
    \Tile_X7Y4_S4BEG[12] ,
    \Tile_X7Y4_S4BEG[11] ,
    \Tile_X7Y4_S4BEG[10] ,
    \Tile_X7Y4_S4BEG[9] ,
    \Tile_X7Y4_S4BEG[8] ,
    \Tile_X7Y4_S4BEG[7] ,
    \Tile_X7Y4_S4BEG[6] ,
    \Tile_X7Y4_S4BEG[5] ,
    \Tile_X7Y4_S4BEG[4] ,
    \Tile_X7Y4_S4BEG[3] ,
    \Tile_X7Y4_S4BEG[2] ,
    \Tile_X7Y4_S4BEG[1] ,
    \Tile_X7Y4_S4BEG[0] }),
    .Tile_X0Y1_SS4BEG({\Tile_X7Y4_SS4BEG[15] ,
    \Tile_X7Y4_SS4BEG[14] ,
    \Tile_X7Y4_SS4BEG[13] ,
    \Tile_X7Y4_SS4BEG[12] ,
    \Tile_X7Y4_SS4BEG[11] ,
    \Tile_X7Y4_SS4BEG[10] ,
    \Tile_X7Y4_SS4BEG[9] ,
    \Tile_X7Y4_SS4BEG[8] ,
    \Tile_X7Y4_SS4BEG[7] ,
    \Tile_X7Y4_SS4BEG[6] ,
    \Tile_X7Y4_SS4BEG[5] ,
    \Tile_X7Y4_SS4BEG[4] ,
    \Tile_X7Y4_SS4BEG[3] ,
    \Tile_X7Y4_SS4BEG[2] ,
    \Tile_X7Y4_SS4BEG[1] ,
    \Tile_X7Y4_SS4BEG[0] }),
    .Tile_X0Y1_W1BEG({\Tile_X7Y4_W1BEG[3] ,
    \Tile_X7Y4_W1BEG[2] ,
    \Tile_X7Y4_W1BEG[1] ,
    \Tile_X7Y4_W1BEG[0] }),
    .Tile_X0Y1_W1END({\Tile_X8Y4_W1BEG[3] ,
    \Tile_X8Y4_W1BEG[2] ,
    \Tile_X8Y4_W1BEG[1] ,
    \Tile_X8Y4_W1BEG[0] }),
    .Tile_X0Y1_W2BEG({\Tile_X7Y4_W2BEG[7] ,
    \Tile_X7Y4_W2BEG[6] ,
    \Tile_X7Y4_W2BEG[5] ,
    \Tile_X7Y4_W2BEG[4] ,
    \Tile_X7Y4_W2BEG[3] ,
    \Tile_X7Y4_W2BEG[2] ,
    \Tile_X7Y4_W2BEG[1] ,
    \Tile_X7Y4_W2BEG[0] }),
    .Tile_X0Y1_W2BEGb({\Tile_X7Y4_W2BEGb[7] ,
    \Tile_X7Y4_W2BEGb[6] ,
    \Tile_X7Y4_W2BEGb[5] ,
    \Tile_X7Y4_W2BEGb[4] ,
    \Tile_X7Y4_W2BEGb[3] ,
    \Tile_X7Y4_W2BEGb[2] ,
    \Tile_X7Y4_W2BEGb[1] ,
    \Tile_X7Y4_W2BEGb[0] }),
    .Tile_X0Y1_W2END({\Tile_X8Y4_W2BEGb[7] ,
    \Tile_X8Y4_W2BEGb[6] ,
    \Tile_X8Y4_W2BEGb[5] ,
    \Tile_X8Y4_W2BEGb[4] ,
    \Tile_X8Y4_W2BEGb[3] ,
    \Tile_X8Y4_W2BEGb[2] ,
    \Tile_X8Y4_W2BEGb[1] ,
    \Tile_X8Y4_W2BEGb[0] }),
    .Tile_X0Y1_W2MID({\Tile_X8Y4_W2BEG[7] ,
    \Tile_X8Y4_W2BEG[6] ,
    \Tile_X8Y4_W2BEG[5] ,
    \Tile_X8Y4_W2BEG[4] ,
    \Tile_X8Y4_W2BEG[3] ,
    \Tile_X8Y4_W2BEG[2] ,
    \Tile_X8Y4_W2BEG[1] ,
    \Tile_X8Y4_W2BEG[0] }),
    .Tile_X0Y1_W6BEG({\Tile_X7Y4_W6BEG[11] ,
    \Tile_X7Y4_W6BEG[10] ,
    \Tile_X7Y4_W6BEG[9] ,
    \Tile_X7Y4_W6BEG[8] ,
    \Tile_X7Y4_W6BEG[7] ,
    \Tile_X7Y4_W6BEG[6] ,
    \Tile_X7Y4_W6BEG[5] ,
    \Tile_X7Y4_W6BEG[4] ,
    \Tile_X7Y4_W6BEG[3] ,
    \Tile_X7Y4_W6BEG[2] ,
    \Tile_X7Y4_W6BEG[1] ,
    \Tile_X7Y4_W6BEG[0] }),
    .Tile_X0Y1_W6END({\Tile_X8Y4_W6BEG[11] ,
    \Tile_X8Y4_W6BEG[10] ,
    \Tile_X8Y4_W6BEG[9] ,
    \Tile_X8Y4_W6BEG[8] ,
    \Tile_X8Y4_W6BEG[7] ,
    \Tile_X8Y4_W6BEG[6] ,
    \Tile_X8Y4_W6BEG[5] ,
    \Tile_X8Y4_W6BEG[4] ,
    \Tile_X8Y4_W6BEG[3] ,
    \Tile_X8Y4_W6BEG[2] ,
    \Tile_X8Y4_W6BEG[1] ,
    \Tile_X8Y4_W6BEG[0] }),
    .Tile_X0Y1_WW4BEG({\Tile_X7Y4_WW4BEG[15] ,
    \Tile_X7Y4_WW4BEG[14] ,
    \Tile_X7Y4_WW4BEG[13] ,
    \Tile_X7Y4_WW4BEG[12] ,
    \Tile_X7Y4_WW4BEG[11] ,
    \Tile_X7Y4_WW4BEG[10] ,
    \Tile_X7Y4_WW4BEG[9] ,
    \Tile_X7Y4_WW4BEG[8] ,
    \Tile_X7Y4_WW4BEG[7] ,
    \Tile_X7Y4_WW4BEG[6] ,
    \Tile_X7Y4_WW4BEG[5] ,
    \Tile_X7Y4_WW4BEG[4] ,
    \Tile_X7Y4_WW4BEG[3] ,
    \Tile_X7Y4_WW4BEG[2] ,
    \Tile_X7Y4_WW4BEG[1] ,
    \Tile_X7Y4_WW4BEG[0] }),
    .Tile_X0Y1_WW4END({\Tile_X8Y4_WW4BEG[15] ,
    \Tile_X8Y4_WW4BEG[14] ,
    \Tile_X8Y4_WW4BEG[13] ,
    \Tile_X8Y4_WW4BEG[12] ,
    \Tile_X8Y4_WW4BEG[11] ,
    \Tile_X8Y4_WW4BEG[10] ,
    \Tile_X8Y4_WW4BEG[9] ,
    \Tile_X8Y4_WW4BEG[8] ,
    \Tile_X8Y4_WW4BEG[7] ,
    \Tile_X8Y4_WW4BEG[6] ,
    \Tile_X8Y4_WW4BEG[5] ,
    \Tile_X8Y4_WW4BEG[4] ,
    \Tile_X8Y4_WW4BEG[3] ,
    \Tile_X8Y4_WW4BEG[2] ,
    \Tile_X8Y4_WW4BEG[1] ,
    \Tile_X8Y4_WW4BEG[0] }));
 DSP Tile_X7Y5_DSP (.Tile_X0Y0_UserCLKo(Tile_X7Y5_UserCLKo),
    .Tile_X0Y1_UserCLK(Tile_X7Y7_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .Tile_X0Y0_E1BEG({\Tile_X7Y5_E1BEG[3] ,
    \Tile_X7Y5_E1BEG[2] ,
    \Tile_X7Y5_E1BEG[1] ,
    \Tile_X7Y5_E1BEG[0] }),
    .Tile_X0Y0_E1END({\Tile_X6Y5_E1BEG[3] ,
    \Tile_X6Y5_E1BEG[2] ,
    \Tile_X6Y5_E1BEG[1] ,
    \Tile_X6Y5_E1BEG[0] }),
    .Tile_X0Y0_E2BEG({\Tile_X7Y5_E2BEG[7] ,
    \Tile_X7Y5_E2BEG[6] ,
    \Tile_X7Y5_E2BEG[5] ,
    \Tile_X7Y5_E2BEG[4] ,
    \Tile_X7Y5_E2BEG[3] ,
    \Tile_X7Y5_E2BEG[2] ,
    \Tile_X7Y5_E2BEG[1] ,
    \Tile_X7Y5_E2BEG[0] }),
    .Tile_X0Y0_E2BEGb({\Tile_X7Y5_E2BEGb[7] ,
    \Tile_X7Y5_E2BEGb[6] ,
    \Tile_X7Y5_E2BEGb[5] ,
    \Tile_X7Y5_E2BEGb[4] ,
    \Tile_X7Y5_E2BEGb[3] ,
    \Tile_X7Y5_E2BEGb[2] ,
    \Tile_X7Y5_E2BEGb[1] ,
    \Tile_X7Y5_E2BEGb[0] }),
    .Tile_X0Y0_E2END({\Tile_X6Y5_E2BEGb[7] ,
    \Tile_X6Y5_E2BEGb[6] ,
    \Tile_X6Y5_E2BEGb[5] ,
    \Tile_X6Y5_E2BEGb[4] ,
    \Tile_X6Y5_E2BEGb[3] ,
    \Tile_X6Y5_E2BEGb[2] ,
    \Tile_X6Y5_E2BEGb[1] ,
    \Tile_X6Y5_E2BEGb[0] }),
    .Tile_X0Y0_E2MID({\Tile_X6Y5_E2BEG[7] ,
    \Tile_X6Y5_E2BEG[6] ,
    \Tile_X6Y5_E2BEG[5] ,
    \Tile_X6Y5_E2BEG[4] ,
    \Tile_X6Y5_E2BEG[3] ,
    \Tile_X6Y5_E2BEG[2] ,
    \Tile_X6Y5_E2BEG[1] ,
    \Tile_X6Y5_E2BEG[0] }),
    .Tile_X0Y0_E6BEG({\Tile_X7Y5_E6BEG[11] ,
    \Tile_X7Y5_E6BEG[10] ,
    \Tile_X7Y5_E6BEG[9] ,
    \Tile_X7Y5_E6BEG[8] ,
    \Tile_X7Y5_E6BEG[7] ,
    \Tile_X7Y5_E6BEG[6] ,
    \Tile_X7Y5_E6BEG[5] ,
    \Tile_X7Y5_E6BEG[4] ,
    \Tile_X7Y5_E6BEG[3] ,
    \Tile_X7Y5_E6BEG[2] ,
    \Tile_X7Y5_E6BEG[1] ,
    \Tile_X7Y5_E6BEG[0] }),
    .Tile_X0Y0_E6END({\Tile_X6Y5_E6BEG[11] ,
    \Tile_X6Y5_E6BEG[10] ,
    \Tile_X6Y5_E6BEG[9] ,
    \Tile_X6Y5_E6BEG[8] ,
    \Tile_X6Y5_E6BEG[7] ,
    \Tile_X6Y5_E6BEG[6] ,
    \Tile_X6Y5_E6BEG[5] ,
    \Tile_X6Y5_E6BEG[4] ,
    \Tile_X6Y5_E6BEG[3] ,
    \Tile_X6Y5_E6BEG[2] ,
    \Tile_X6Y5_E6BEG[1] ,
    \Tile_X6Y5_E6BEG[0] }),
    .Tile_X0Y0_EE4BEG({\Tile_X7Y5_EE4BEG[15] ,
    \Tile_X7Y5_EE4BEG[14] ,
    \Tile_X7Y5_EE4BEG[13] ,
    \Tile_X7Y5_EE4BEG[12] ,
    \Tile_X7Y5_EE4BEG[11] ,
    \Tile_X7Y5_EE4BEG[10] ,
    \Tile_X7Y5_EE4BEG[9] ,
    \Tile_X7Y5_EE4BEG[8] ,
    \Tile_X7Y5_EE4BEG[7] ,
    \Tile_X7Y5_EE4BEG[6] ,
    \Tile_X7Y5_EE4BEG[5] ,
    \Tile_X7Y5_EE4BEG[4] ,
    \Tile_X7Y5_EE4BEG[3] ,
    \Tile_X7Y5_EE4BEG[2] ,
    \Tile_X7Y5_EE4BEG[1] ,
    \Tile_X7Y5_EE4BEG[0] }),
    .Tile_X0Y0_EE4END({\Tile_X6Y5_EE4BEG[15] ,
    \Tile_X6Y5_EE4BEG[14] ,
    \Tile_X6Y5_EE4BEG[13] ,
    \Tile_X6Y5_EE4BEG[12] ,
    \Tile_X6Y5_EE4BEG[11] ,
    \Tile_X6Y5_EE4BEG[10] ,
    \Tile_X6Y5_EE4BEG[9] ,
    \Tile_X6Y5_EE4BEG[8] ,
    \Tile_X6Y5_EE4BEG[7] ,
    \Tile_X6Y5_EE4BEG[6] ,
    \Tile_X6Y5_EE4BEG[5] ,
    \Tile_X6Y5_EE4BEG[4] ,
    \Tile_X6Y5_EE4BEG[3] ,
    \Tile_X6Y5_EE4BEG[2] ,
    \Tile_X6Y5_EE4BEG[1] ,
    \Tile_X6Y5_EE4BEG[0] }),
    .Tile_X0Y0_FrameData({\Tile_X6Y5_FrameData_O[31] ,
    \Tile_X6Y5_FrameData_O[30] ,
    \Tile_X6Y5_FrameData_O[29] ,
    \Tile_X6Y5_FrameData_O[28] ,
    \Tile_X6Y5_FrameData_O[27] ,
    \Tile_X6Y5_FrameData_O[26] ,
    \Tile_X6Y5_FrameData_O[25] ,
    \Tile_X6Y5_FrameData_O[24] ,
    \Tile_X6Y5_FrameData_O[23] ,
    \Tile_X6Y5_FrameData_O[22] ,
    \Tile_X6Y5_FrameData_O[21] ,
    \Tile_X6Y5_FrameData_O[20] ,
    \Tile_X6Y5_FrameData_O[19] ,
    \Tile_X6Y5_FrameData_O[18] ,
    \Tile_X6Y5_FrameData_O[17] ,
    \Tile_X6Y5_FrameData_O[16] ,
    \Tile_X6Y5_FrameData_O[15] ,
    \Tile_X6Y5_FrameData_O[14] ,
    \Tile_X6Y5_FrameData_O[13] ,
    \Tile_X6Y5_FrameData_O[12] ,
    \Tile_X6Y5_FrameData_O[11] ,
    \Tile_X6Y5_FrameData_O[10] ,
    \Tile_X6Y5_FrameData_O[9] ,
    \Tile_X6Y5_FrameData_O[8] ,
    \Tile_X6Y5_FrameData_O[7] ,
    \Tile_X6Y5_FrameData_O[6] ,
    \Tile_X6Y5_FrameData_O[5] ,
    \Tile_X6Y5_FrameData_O[4] ,
    \Tile_X6Y5_FrameData_O[3] ,
    \Tile_X6Y5_FrameData_O[2] ,
    \Tile_X6Y5_FrameData_O[1] ,
    \Tile_X6Y5_FrameData_O[0] }),
    .Tile_X0Y0_FrameData_O({\Tile_X7Y5_FrameData_O[31] ,
    \Tile_X7Y5_FrameData_O[30] ,
    \Tile_X7Y5_FrameData_O[29] ,
    \Tile_X7Y5_FrameData_O[28] ,
    \Tile_X7Y5_FrameData_O[27] ,
    \Tile_X7Y5_FrameData_O[26] ,
    \Tile_X7Y5_FrameData_O[25] ,
    \Tile_X7Y5_FrameData_O[24] ,
    \Tile_X7Y5_FrameData_O[23] ,
    \Tile_X7Y5_FrameData_O[22] ,
    \Tile_X7Y5_FrameData_O[21] ,
    \Tile_X7Y5_FrameData_O[20] ,
    \Tile_X7Y5_FrameData_O[19] ,
    \Tile_X7Y5_FrameData_O[18] ,
    \Tile_X7Y5_FrameData_O[17] ,
    \Tile_X7Y5_FrameData_O[16] ,
    \Tile_X7Y5_FrameData_O[15] ,
    \Tile_X7Y5_FrameData_O[14] ,
    \Tile_X7Y5_FrameData_O[13] ,
    \Tile_X7Y5_FrameData_O[12] ,
    \Tile_X7Y5_FrameData_O[11] ,
    \Tile_X7Y5_FrameData_O[10] ,
    \Tile_X7Y5_FrameData_O[9] ,
    \Tile_X7Y5_FrameData_O[8] ,
    \Tile_X7Y5_FrameData_O[7] ,
    \Tile_X7Y5_FrameData_O[6] ,
    \Tile_X7Y5_FrameData_O[5] ,
    \Tile_X7Y5_FrameData_O[4] ,
    \Tile_X7Y5_FrameData_O[3] ,
    \Tile_X7Y5_FrameData_O[2] ,
    \Tile_X7Y5_FrameData_O[1] ,
    \Tile_X7Y5_FrameData_O[0] }),
    .Tile_X0Y0_FrameStrobe_O({\Tile_X7Y5_FrameStrobe_O[19] ,
    \Tile_X7Y5_FrameStrobe_O[18] ,
    \Tile_X7Y5_FrameStrobe_O[17] ,
    \Tile_X7Y5_FrameStrobe_O[16] ,
    \Tile_X7Y5_FrameStrobe_O[15] ,
    \Tile_X7Y5_FrameStrobe_O[14] ,
    \Tile_X7Y5_FrameStrobe_O[13] ,
    \Tile_X7Y5_FrameStrobe_O[12] ,
    \Tile_X7Y5_FrameStrobe_O[11] ,
    \Tile_X7Y5_FrameStrobe_O[10] ,
    \Tile_X7Y5_FrameStrobe_O[9] ,
    \Tile_X7Y5_FrameStrobe_O[8] ,
    \Tile_X7Y5_FrameStrobe_O[7] ,
    \Tile_X7Y5_FrameStrobe_O[6] ,
    \Tile_X7Y5_FrameStrobe_O[5] ,
    \Tile_X7Y5_FrameStrobe_O[4] ,
    \Tile_X7Y5_FrameStrobe_O[3] ,
    \Tile_X7Y5_FrameStrobe_O[2] ,
    \Tile_X7Y5_FrameStrobe_O[1] ,
    \Tile_X7Y5_FrameStrobe_O[0] }),
    .Tile_X0Y0_N1BEG({\Tile_X7Y5_N1BEG[3] ,
    \Tile_X7Y5_N1BEG[2] ,
    \Tile_X7Y5_N1BEG[1] ,
    \Tile_X7Y5_N1BEG[0] }),
    .Tile_X0Y0_N2BEG({\Tile_X7Y5_N2BEG[7] ,
    \Tile_X7Y5_N2BEG[6] ,
    \Tile_X7Y5_N2BEG[5] ,
    \Tile_X7Y5_N2BEG[4] ,
    \Tile_X7Y5_N2BEG[3] ,
    \Tile_X7Y5_N2BEG[2] ,
    \Tile_X7Y5_N2BEG[1] ,
    \Tile_X7Y5_N2BEG[0] }),
    .Tile_X0Y0_N2BEGb({\Tile_X7Y5_N2BEGb[7] ,
    \Tile_X7Y5_N2BEGb[6] ,
    \Tile_X7Y5_N2BEGb[5] ,
    \Tile_X7Y5_N2BEGb[4] ,
    \Tile_X7Y5_N2BEGb[3] ,
    \Tile_X7Y5_N2BEGb[2] ,
    \Tile_X7Y5_N2BEGb[1] ,
    \Tile_X7Y5_N2BEGb[0] }),
    .Tile_X0Y0_N4BEG({\Tile_X7Y5_N4BEG[15] ,
    \Tile_X7Y5_N4BEG[14] ,
    \Tile_X7Y5_N4BEG[13] ,
    \Tile_X7Y5_N4BEG[12] ,
    \Tile_X7Y5_N4BEG[11] ,
    \Tile_X7Y5_N4BEG[10] ,
    \Tile_X7Y5_N4BEG[9] ,
    \Tile_X7Y5_N4BEG[8] ,
    \Tile_X7Y5_N4BEG[7] ,
    \Tile_X7Y5_N4BEG[6] ,
    \Tile_X7Y5_N4BEG[5] ,
    \Tile_X7Y5_N4BEG[4] ,
    \Tile_X7Y5_N4BEG[3] ,
    \Tile_X7Y5_N4BEG[2] ,
    \Tile_X7Y5_N4BEG[1] ,
    \Tile_X7Y5_N4BEG[0] }),
    .Tile_X0Y0_NN4BEG({\Tile_X7Y5_NN4BEG[15] ,
    \Tile_X7Y5_NN4BEG[14] ,
    \Tile_X7Y5_NN4BEG[13] ,
    \Tile_X7Y5_NN4BEG[12] ,
    \Tile_X7Y5_NN4BEG[11] ,
    \Tile_X7Y5_NN4BEG[10] ,
    \Tile_X7Y5_NN4BEG[9] ,
    \Tile_X7Y5_NN4BEG[8] ,
    \Tile_X7Y5_NN4BEG[7] ,
    \Tile_X7Y5_NN4BEG[6] ,
    \Tile_X7Y5_NN4BEG[5] ,
    \Tile_X7Y5_NN4BEG[4] ,
    \Tile_X7Y5_NN4BEG[3] ,
    \Tile_X7Y5_NN4BEG[2] ,
    \Tile_X7Y5_NN4BEG[1] ,
    \Tile_X7Y5_NN4BEG[0] }),
    .Tile_X0Y0_S1END({\Tile_X7Y4_S1BEG[3] ,
    \Tile_X7Y4_S1BEG[2] ,
    \Tile_X7Y4_S1BEG[1] ,
    \Tile_X7Y4_S1BEG[0] }),
    .Tile_X0Y0_S2END({\Tile_X7Y4_S2BEGb[7] ,
    \Tile_X7Y4_S2BEGb[6] ,
    \Tile_X7Y4_S2BEGb[5] ,
    \Tile_X7Y4_S2BEGb[4] ,
    \Tile_X7Y4_S2BEGb[3] ,
    \Tile_X7Y4_S2BEGb[2] ,
    \Tile_X7Y4_S2BEGb[1] ,
    \Tile_X7Y4_S2BEGb[0] }),
    .Tile_X0Y0_S2MID({\Tile_X7Y4_S2BEG[7] ,
    \Tile_X7Y4_S2BEG[6] ,
    \Tile_X7Y4_S2BEG[5] ,
    \Tile_X7Y4_S2BEG[4] ,
    \Tile_X7Y4_S2BEG[3] ,
    \Tile_X7Y4_S2BEG[2] ,
    \Tile_X7Y4_S2BEG[1] ,
    \Tile_X7Y4_S2BEG[0] }),
    .Tile_X0Y0_S4END({\Tile_X7Y4_S4BEG[15] ,
    \Tile_X7Y4_S4BEG[14] ,
    \Tile_X7Y4_S4BEG[13] ,
    \Tile_X7Y4_S4BEG[12] ,
    \Tile_X7Y4_S4BEG[11] ,
    \Tile_X7Y4_S4BEG[10] ,
    \Tile_X7Y4_S4BEG[9] ,
    \Tile_X7Y4_S4BEG[8] ,
    \Tile_X7Y4_S4BEG[7] ,
    \Tile_X7Y4_S4BEG[6] ,
    \Tile_X7Y4_S4BEG[5] ,
    \Tile_X7Y4_S4BEG[4] ,
    \Tile_X7Y4_S4BEG[3] ,
    \Tile_X7Y4_S4BEG[2] ,
    \Tile_X7Y4_S4BEG[1] ,
    \Tile_X7Y4_S4BEG[0] }),
    .Tile_X0Y0_SS4END({\Tile_X7Y4_SS4BEG[15] ,
    \Tile_X7Y4_SS4BEG[14] ,
    \Tile_X7Y4_SS4BEG[13] ,
    \Tile_X7Y4_SS4BEG[12] ,
    \Tile_X7Y4_SS4BEG[11] ,
    \Tile_X7Y4_SS4BEG[10] ,
    \Tile_X7Y4_SS4BEG[9] ,
    \Tile_X7Y4_SS4BEG[8] ,
    \Tile_X7Y4_SS4BEG[7] ,
    \Tile_X7Y4_SS4BEG[6] ,
    \Tile_X7Y4_SS4BEG[5] ,
    \Tile_X7Y4_SS4BEG[4] ,
    \Tile_X7Y4_SS4BEG[3] ,
    \Tile_X7Y4_SS4BEG[2] ,
    \Tile_X7Y4_SS4BEG[1] ,
    \Tile_X7Y4_SS4BEG[0] }),
    .Tile_X0Y0_W1BEG({\Tile_X7Y5_W1BEG[3] ,
    \Tile_X7Y5_W1BEG[2] ,
    \Tile_X7Y5_W1BEG[1] ,
    \Tile_X7Y5_W1BEG[0] }),
    .Tile_X0Y0_W1END({\Tile_X8Y5_W1BEG[3] ,
    \Tile_X8Y5_W1BEG[2] ,
    \Tile_X8Y5_W1BEG[1] ,
    \Tile_X8Y5_W1BEG[0] }),
    .Tile_X0Y0_W2BEG({\Tile_X7Y5_W2BEG[7] ,
    \Tile_X7Y5_W2BEG[6] ,
    \Tile_X7Y5_W2BEG[5] ,
    \Tile_X7Y5_W2BEG[4] ,
    \Tile_X7Y5_W2BEG[3] ,
    \Tile_X7Y5_W2BEG[2] ,
    \Tile_X7Y5_W2BEG[1] ,
    \Tile_X7Y5_W2BEG[0] }),
    .Tile_X0Y0_W2BEGb({\Tile_X7Y5_W2BEGb[7] ,
    \Tile_X7Y5_W2BEGb[6] ,
    \Tile_X7Y5_W2BEGb[5] ,
    \Tile_X7Y5_W2BEGb[4] ,
    \Tile_X7Y5_W2BEGb[3] ,
    \Tile_X7Y5_W2BEGb[2] ,
    \Tile_X7Y5_W2BEGb[1] ,
    \Tile_X7Y5_W2BEGb[0] }),
    .Tile_X0Y0_W2END({\Tile_X8Y5_W2BEGb[7] ,
    \Tile_X8Y5_W2BEGb[6] ,
    \Tile_X8Y5_W2BEGb[5] ,
    \Tile_X8Y5_W2BEGb[4] ,
    \Tile_X8Y5_W2BEGb[3] ,
    \Tile_X8Y5_W2BEGb[2] ,
    \Tile_X8Y5_W2BEGb[1] ,
    \Tile_X8Y5_W2BEGb[0] }),
    .Tile_X0Y0_W2MID({\Tile_X8Y5_W2BEG[7] ,
    \Tile_X8Y5_W2BEG[6] ,
    \Tile_X8Y5_W2BEG[5] ,
    \Tile_X8Y5_W2BEG[4] ,
    \Tile_X8Y5_W2BEG[3] ,
    \Tile_X8Y5_W2BEG[2] ,
    \Tile_X8Y5_W2BEG[1] ,
    \Tile_X8Y5_W2BEG[0] }),
    .Tile_X0Y0_W6BEG({\Tile_X7Y5_W6BEG[11] ,
    \Tile_X7Y5_W6BEG[10] ,
    \Tile_X7Y5_W6BEG[9] ,
    \Tile_X7Y5_W6BEG[8] ,
    \Tile_X7Y5_W6BEG[7] ,
    \Tile_X7Y5_W6BEG[6] ,
    \Tile_X7Y5_W6BEG[5] ,
    \Tile_X7Y5_W6BEG[4] ,
    \Tile_X7Y5_W6BEG[3] ,
    \Tile_X7Y5_W6BEG[2] ,
    \Tile_X7Y5_W6BEG[1] ,
    \Tile_X7Y5_W6BEG[0] }),
    .Tile_X0Y0_W6END({\Tile_X8Y5_W6BEG[11] ,
    \Tile_X8Y5_W6BEG[10] ,
    \Tile_X8Y5_W6BEG[9] ,
    \Tile_X8Y5_W6BEG[8] ,
    \Tile_X8Y5_W6BEG[7] ,
    \Tile_X8Y5_W6BEG[6] ,
    \Tile_X8Y5_W6BEG[5] ,
    \Tile_X8Y5_W6BEG[4] ,
    \Tile_X8Y5_W6BEG[3] ,
    \Tile_X8Y5_W6BEG[2] ,
    \Tile_X8Y5_W6BEG[1] ,
    \Tile_X8Y5_W6BEG[0] }),
    .Tile_X0Y0_WW4BEG({\Tile_X7Y5_WW4BEG[15] ,
    \Tile_X7Y5_WW4BEG[14] ,
    \Tile_X7Y5_WW4BEG[13] ,
    \Tile_X7Y5_WW4BEG[12] ,
    \Tile_X7Y5_WW4BEG[11] ,
    \Tile_X7Y5_WW4BEG[10] ,
    \Tile_X7Y5_WW4BEG[9] ,
    \Tile_X7Y5_WW4BEG[8] ,
    \Tile_X7Y5_WW4BEG[7] ,
    \Tile_X7Y5_WW4BEG[6] ,
    \Tile_X7Y5_WW4BEG[5] ,
    \Tile_X7Y5_WW4BEG[4] ,
    \Tile_X7Y5_WW4BEG[3] ,
    \Tile_X7Y5_WW4BEG[2] ,
    \Tile_X7Y5_WW4BEG[1] ,
    \Tile_X7Y5_WW4BEG[0] }),
    .Tile_X0Y0_WW4END({\Tile_X8Y5_WW4BEG[15] ,
    \Tile_X8Y5_WW4BEG[14] ,
    \Tile_X8Y5_WW4BEG[13] ,
    \Tile_X8Y5_WW4BEG[12] ,
    \Tile_X8Y5_WW4BEG[11] ,
    \Tile_X8Y5_WW4BEG[10] ,
    \Tile_X8Y5_WW4BEG[9] ,
    \Tile_X8Y5_WW4BEG[8] ,
    \Tile_X8Y5_WW4BEG[7] ,
    \Tile_X8Y5_WW4BEG[6] ,
    \Tile_X8Y5_WW4BEG[5] ,
    \Tile_X8Y5_WW4BEG[4] ,
    \Tile_X8Y5_WW4BEG[3] ,
    \Tile_X8Y5_WW4BEG[2] ,
    \Tile_X8Y5_WW4BEG[1] ,
    \Tile_X8Y5_WW4BEG[0] }),
    .Tile_X0Y1_E1BEG({\Tile_X7Y6_E1BEG[3] ,
    \Tile_X7Y6_E1BEG[2] ,
    \Tile_X7Y6_E1BEG[1] ,
    \Tile_X7Y6_E1BEG[0] }),
    .Tile_X0Y1_E1END({\Tile_X6Y6_E1BEG[3] ,
    \Tile_X6Y6_E1BEG[2] ,
    \Tile_X6Y6_E1BEG[1] ,
    \Tile_X6Y6_E1BEG[0] }),
    .Tile_X0Y1_E2BEG({\Tile_X7Y6_E2BEG[7] ,
    \Tile_X7Y6_E2BEG[6] ,
    \Tile_X7Y6_E2BEG[5] ,
    \Tile_X7Y6_E2BEG[4] ,
    \Tile_X7Y6_E2BEG[3] ,
    \Tile_X7Y6_E2BEG[2] ,
    \Tile_X7Y6_E2BEG[1] ,
    \Tile_X7Y6_E2BEG[0] }),
    .Tile_X0Y1_E2BEGb({\Tile_X7Y6_E2BEGb[7] ,
    \Tile_X7Y6_E2BEGb[6] ,
    \Tile_X7Y6_E2BEGb[5] ,
    \Tile_X7Y6_E2BEGb[4] ,
    \Tile_X7Y6_E2BEGb[3] ,
    \Tile_X7Y6_E2BEGb[2] ,
    \Tile_X7Y6_E2BEGb[1] ,
    \Tile_X7Y6_E2BEGb[0] }),
    .Tile_X0Y1_E2END({\Tile_X6Y6_E2BEGb[7] ,
    \Tile_X6Y6_E2BEGb[6] ,
    \Tile_X6Y6_E2BEGb[5] ,
    \Tile_X6Y6_E2BEGb[4] ,
    \Tile_X6Y6_E2BEGb[3] ,
    \Tile_X6Y6_E2BEGb[2] ,
    \Tile_X6Y6_E2BEGb[1] ,
    \Tile_X6Y6_E2BEGb[0] }),
    .Tile_X0Y1_E2MID({\Tile_X6Y6_E2BEG[7] ,
    \Tile_X6Y6_E2BEG[6] ,
    \Tile_X6Y6_E2BEG[5] ,
    \Tile_X6Y6_E2BEG[4] ,
    \Tile_X6Y6_E2BEG[3] ,
    \Tile_X6Y6_E2BEG[2] ,
    \Tile_X6Y6_E2BEG[1] ,
    \Tile_X6Y6_E2BEG[0] }),
    .Tile_X0Y1_E6BEG({\Tile_X7Y6_E6BEG[11] ,
    \Tile_X7Y6_E6BEG[10] ,
    \Tile_X7Y6_E6BEG[9] ,
    \Tile_X7Y6_E6BEG[8] ,
    \Tile_X7Y6_E6BEG[7] ,
    \Tile_X7Y6_E6BEG[6] ,
    \Tile_X7Y6_E6BEG[5] ,
    \Tile_X7Y6_E6BEG[4] ,
    \Tile_X7Y6_E6BEG[3] ,
    \Tile_X7Y6_E6BEG[2] ,
    \Tile_X7Y6_E6BEG[1] ,
    \Tile_X7Y6_E6BEG[0] }),
    .Tile_X0Y1_E6END({\Tile_X6Y6_E6BEG[11] ,
    \Tile_X6Y6_E6BEG[10] ,
    \Tile_X6Y6_E6BEG[9] ,
    \Tile_X6Y6_E6BEG[8] ,
    \Tile_X6Y6_E6BEG[7] ,
    \Tile_X6Y6_E6BEG[6] ,
    \Tile_X6Y6_E6BEG[5] ,
    \Tile_X6Y6_E6BEG[4] ,
    \Tile_X6Y6_E6BEG[3] ,
    \Tile_X6Y6_E6BEG[2] ,
    \Tile_X6Y6_E6BEG[1] ,
    \Tile_X6Y6_E6BEG[0] }),
    .Tile_X0Y1_EE4BEG({\Tile_X7Y6_EE4BEG[15] ,
    \Tile_X7Y6_EE4BEG[14] ,
    \Tile_X7Y6_EE4BEG[13] ,
    \Tile_X7Y6_EE4BEG[12] ,
    \Tile_X7Y6_EE4BEG[11] ,
    \Tile_X7Y6_EE4BEG[10] ,
    \Tile_X7Y6_EE4BEG[9] ,
    \Tile_X7Y6_EE4BEG[8] ,
    \Tile_X7Y6_EE4BEG[7] ,
    \Tile_X7Y6_EE4BEG[6] ,
    \Tile_X7Y6_EE4BEG[5] ,
    \Tile_X7Y6_EE4BEG[4] ,
    \Tile_X7Y6_EE4BEG[3] ,
    \Tile_X7Y6_EE4BEG[2] ,
    \Tile_X7Y6_EE4BEG[1] ,
    \Tile_X7Y6_EE4BEG[0] }),
    .Tile_X0Y1_EE4END({\Tile_X6Y6_EE4BEG[15] ,
    \Tile_X6Y6_EE4BEG[14] ,
    \Tile_X6Y6_EE4BEG[13] ,
    \Tile_X6Y6_EE4BEG[12] ,
    \Tile_X6Y6_EE4BEG[11] ,
    \Tile_X6Y6_EE4BEG[10] ,
    \Tile_X6Y6_EE4BEG[9] ,
    \Tile_X6Y6_EE4BEG[8] ,
    \Tile_X6Y6_EE4BEG[7] ,
    \Tile_X6Y6_EE4BEG[6] ,
    \Tile_X6Y6_EE4BEG[5] ,
    \Tile_X6Y6_EE4BEG[4] ,
    \Tile_X6Y6_EE4BEG[3] ,
    \Tile_X6Y6_EE4BEG[2] ,
    \Tile_X6Y6_EE4BEG[1] ,
    \Tile_X6Y6_EE4BEG[0] }),
    .Tile_X0Y1_FrameData({\Tile_X6Y6_FrameData_O[31] ,
    \Tile_X6Y6_FrameData_O[30] ,
    \Tile_X6Y6_FrameData_O[29] ,
    \Tile_X6Y6_FrameData_O[28] ,
    \Tile_X6Y6_FrameData_O[27] ,
    \Tile_X6Y6_FrameData_O[26] ,
    \Tile_X6Y6_FrameData_O[25] ,
    \Tile_X6Y6_FrameData_O[24] ,
    \Tile_X6Y6_FrameData_O[23] ,
    \Tile_X6Y6_FrameData_O[22] ,
    \Tile_X6Y6_FrameData_O[21] ,
    \Tile_X6Y6_FrameData_O[20] ,
    \Tile_X6Y6_FrameData_O[19] ,
    \Tile_X6Y6_FrameData_O[18] ,
    \Tile_X6Y6_FrameData_O[17] ,
    \Tile_X6Y6_FrameData_O[16] ,
    \Tile_X6Y6_FrameData_O[15] ,
    \Tile_X6Y6_FrameData_O[14] ,
    \Tile_X6Y6_FrameData_O[13] ,
    \Tile_X6Y6_FrameData_O[12] ,
    \Tile_X6Y6_FrameData_O[11] ,
    \Tile_X6Y6_FrameData_O[10] ,
    \Tile_X6Y6_FrameData_O[9] ,
    \Tile_X6Y6_FrameData_O[8] ,
    \Tile_X6Y6_FrameData_O[7] ,
    \Tile_X6Y6_FrameData_O[6] ,
    \Tile_X6Y6_FrameData_O[5] ,
    \Tile_X6Y6_FrameData_O[4] ,
    \Tile_X6Y6_FrameData_O[3] ,
    \Tile_X6Y6_FrameData_O[2] ,
    \Tile_X6Y6_FrameData_O[1] ,
    \Tile_X6Y6_FrameData_O[0] }),
    .Tile_X0Y1_FrameData_O({\Tile_X7Y6_FrameData_O[31] ,
    \Tile_X7Y6_FrameData_O[30] ,
    \Tile_X7Y6_FrameData_O[29] ,
    \Tile_X7Y6_FrameData_O[28] ,
    \Tile_X7Y6_FrameData_O[27] ,
    \Tile_X7Y6_FrameData_O[26] ,
    \Tile_X7Y6_FrameData_O[25] ,
    \Tile_X7Y6_FrameData_O[24] ,
    \Tile_X7Y6_FrameData_O[23] ,
    \Tile_X7Y6_FrameData_O[22] ,
    \Tile_X7Y6_FrameData_O[21] ,
    \Tile_X7Y6_FrameData_O[20] ,
    \Tile_X7Y6_FrameData_O[19] ,
    \Tile_X7Y6_FrameData_O[18] ,
    \Tile_X7Y6_FrameData_O[17] ,
    \Tile_X7Y6_FrameData_O[16] ,
    \Tile_X7Y6_FrameData_O[15] ,
    \Tile_X7Y6_FrameData_O[14] ,
    \Tile_X7Y6_FrameData_O[13] ,
    \Tile_X7Y6_FrameData_O[12] ,
    \Tile_X7Y6_FrameData_O[11] ,
    \Tile_X7Y6_FrameData_O[10] ,
    \Tile_X7Y6_FrameData_O[9] ,
    \Tile_X7Y6_FrameData_O[8] ,
    \Tile_X7Y6_FrameData_O[7] ,
    \Tile_X7Y6_FrameData_O[6] ,
    \Tile_X7Y6_FrameData_O[5] ,
    \Tile_X7Y6_FrameData_O[4] ,
    \Tile_X7Y6_FrameData_O[3] ,
    \Tile_X7Y6_FrameData_O[2] ,
    \Tile_X7Y6_FrameData_O[1] ,
    \Tile_X7Y6_FrameData_O[0] }),
    .Tile_X0Y1_FrameStrobe({\Tile_X7Y7_FrameStrobe_O[19] ,
    \Tile_X7Y7_FrameStrobe_O[18] ,
    \Tile_X7Y7_FrameStrobe_O[17] ,
    \Tile_X7Y7_FrameStrobe_O[16] ,
    \Tile_X7Y7_FrameStrobe_O[15] ,
    \Tile_X7Y7_FrameStrobe_O[14] ,
    \Tile_X7Y7_FrameStrobe_O[13] ,
    \Tile_X7Y7_FrameStrobe_O[12] ,
    \Tile_X7Y7_FrameStrobe_O[11] ,
    \Tile_X7Y7_FrameStrobe_O[10] ,
    \Tile_X7Y7_FrameStrobe_O[9] ,
    \Tile_X7Y7_FrameStrobe_O[8] ,
    \Tile_X7Y7_FrameStrobe_O[7] ,
    \Tile_X7Y7_FrameStrobe_O[6] ,
    \Tile_X7Y7_FrameStrobe_O[5] ,
    \Tile_X7Y7_FrameStrobe_O[4] ,
    \Tile_X7Y7_FrameStrobe_O[3] ,
    \Tile_X7Y7_FrameStrobe_O[2] ,
    \Tile_X7Y7_FrameStrobe_O[1] ,
    \Tile_X7Y7_FrameStrobe_O[0] }),
    .Tile_X0Y1_N1END({\Tile_X7Y7_N1BEG[3] ,
    \Tile_X7Y7_N1BEG[2] ,
    \Tile_X7Y7_N1BEG[1] ,
    \Tile_X7Y7_N1BEG[0] }),
    .Tile_X0Y1_N2END({\Tile_X7Y7_N2BEGb[7] ,
    \Tile_X7Y7_N2BEGb[6] ,
    \Tile_X7Y7_N2BEGb[5] ,
    \Tile_X7Y7_N2BEGb[4] ,
    \Tile_X7Y7_N2BEGb[3] ,
    \Tile_X7Y7_N2BEGb[2] ,
    \Tile_X7Y7_N2BEGb[1] ,
    \Tile_X7Y7_N2BEGb[0] }),
    .Tile_X0Y1_N2MID({\Tile_X7Y7_N2BEG[7] ,
    \Tile_X7Y7_N2BEG[6] ,
    \Tile_X7Y7_N2BEG[5] ,
    \Tile_X7Y7_N2BEG[4] ,
    \Tile_X7Y7_N2BEG[3] ,
    \Tile_X7Y7_N2BEG[2] ,
    \Tile_X7Y7_N2BEG[1] ,
    \Tile_X7Y7_N2BEG[0] }),
    .Tile_X0Y1_N4END({\Tile_X7Y7_N4BEG[15] ,
    \Tile_X7Y7_N4BEG[14] ,
    \Tile_X7Y7_N4BEG[13] ,
    \Tile_X7Y7_N4BEG[12] ,
    \Tile_X7Y7_N4BEG[11] ,
    \Tile_X7Y7_N4BEG[10] ,
    \Tile_X7Y7_N4BEG[9] ,
    \Tile_X7Y7_N4BEG[8] ,
    \Tile_X7Y7_N4BEG[7] ,
    \Tile_X7Y7_N4BEG[6] ,
    \Tile_X7Y7_N4BEG[5] ,
    \Tile_X7Y7_N4BEG[4] ,
    \Tile_X7Y7_N4BEG[3] ,
    \Tile_X7Y7_N4BEG[2] ,
    \Tile_X7Y7_N4BEG[1] ,
    \Tile_X7Y7_N4BEG[0] }),
    .Tile_X0Y1_NN4END({\Tile_X7Y7_NN4BEG[15] ,
    \Tile_X7Y7_NN4BEG[14] ,
    \Tile_X7Y7_NN4BEG[13] ,
    \Tile_X7Y7_NN4BEG[12] ,
    \Tile_X7Y7_NN4BEG[11] ,
    \Tile_X7Y7_NN4BEG[10] ,
    \Tile_X7Y7_NN4BEG[9] ,
    \Tile_X7Y7_NN4BEG[8] ,
    \Tile_X7Y7_NN4BEG[7] ,
    \Tile_X7Y7_NN4BEG[6] ,
    \Tile_X7Y7_NN4BEG[5] ,
    \Tile_X7Y7_NN4BEG[4] ,
    \Tile_X7Y7_NN4BEG[3] ,
    \Tile_X7Y7_NN4BEG[2] ,
    \Tile_X7Y7_NN4BEG[1] ,
    \Tile_X7Y7_NN4BEG[0] }),
    .Tile_X0Y1_S1BEG({\Tile_X7Y6_S1BEG[3] ,
    \Tile_X7Y6_S1BEG[2] ,
    \Tile_X7Y6_S1BEG[1] ,
    \Tile_X7Y6_S1BEG[0] }),
    .Tile_X0Y1_S2BEG({\Tile_X7Y6_S2BEG[7] ,
    \Tile_X7Y6_S2BEG[6] ,
    \Tile_X7Y6_S2BEG[5] ,
    \Tile_X7Y6_S2BEG[4] ,
    \Tile_X7Y6_S2BEG[3] ,
    \Tile_X7Y6_S2BEG[2] ,
    \Tile_X7Y6_S2BEG[1] ,
    \Tile_X7Y6_S2BEG[0] }),
    .Tile_X0Y1_S2BEGb({\Tile_X7Y6_S2BEGb[7] ,
    \Tile_X7Y6_S2BEGb[6] ,
    \Tile_X7Y6_S2BEGb[5] ,
    \Tile_X7Y6_S2BEGb[4] ,
    \Tile_X7Y6_S2BEGb[3] ,
    \Tile_X7Y6_S2BEGb[2] ,
    \Tile_X7Y6_S2BEGb[1] ,
    \Tile_X7Y6_S2BEGb[0] }),
    .Tile_X0Y1_S4BEG({\Tile_X7Y6_S4BEG[15] ,
    \Tile_X7Y6_S4BEG[14] ,
    \Tile_X7Y6_S4BEG[13] ,
    \Tile_X7Y6_S4BEG[12] ,
    \Tile_X7Y6_S4BEG[11] ,
    \Tile_X7Y6_S4BEG[10] ,
    \Tile_X7Y6_S4BEG[9] ,
    \Tile_X7Y6_S4BEG[8] ,
    \Tile_X7Y6_S4BEG[7] ,
    \Tile_X7Y6_S4BEG[6] ,
    \Tile_X7Y6_S4BEG[5] ,
    \Tile_X7Y6_S4BEG[4] ,
    \Tile_X7Y6_S4BEG[3] ,
    \Tile_X7Y6_S4BEG[2] ,
    \Tile_X7Y6_S4BEG[1] ,
    \Tile_X7Y6_S4BEG[0] }),
    .Tile_X0Y1_SS4BEG({\Tile_X7Y6_SS4BEG[15] ,
    \Tile_X7Y6_SS4BEG[14] ,
    \Tile_X7Y6_SS4BEG[13] ,
    \Tile_X7Y6_SS4BEG[12] ,
    \Tile_X7Y6_SS4BEG[11] ,
    \Tile_X7Y6_SS4BEG[10] ,
    \Tile_X7Y6_SS4BEG[9] ,
    \Tile_X7Y6_SS4BEG[8] ,
    \Tile_X7Y6_SS4BEG[7] ,
    \Tile_X7Y6_SS4BEG[6] ,
    \Tile_X7Y6_SS4BEG[5] ,
    \Tile_X7Y6_SS4BEG[4] ,
    \Tile_X7Y6_SS4BEG[3] ,
    \Tile_X7Y6_SS4BEG[2] ,
    \Tile_X7Y6_SS4BEG[1] ,
    \Tile_X7Y6_SS4BEG[0] }),
    .Tile_X0Y1_W1BEG({\Tile_X7Y6_W1BEG[3] ,
    \Tile_X7Y6_W1BEG[2] ,
    \Tile_X7Y6_W1BEG[1] ,
    \Tile_X7Y6_W1BEG[0] }),
    .Tile_X0Y1_W1END({\Tile_X8Y6_W1BEG[3] ,
    \Tile_X8Y6_W1BEG[2] ,
    \Tile_X8Y6_W1BEG[1] ,
    \Tile_X8Y6_W1BEG[0] }),
    .Tile_X0Y1_W2BEG({\Tile_X7Y6_W2BEG[7] ,
    \Tile_X7Y6_W2BEG[6] ,
    \Tile_X7Y6_W2BEG[5] ,
    \Tile_X7Y6_W2BEG[4] ,
    \Tile_X7Y6_W2BEG[3] ,
    \Tile_X7Y6_W2BEG[2] ,
    \Tile_X7Y6_W2BEG[1] ,
    \Tile_X7Y6_W2BEG[0] }),
    .Tile_X0Y1_W2BEGb({\Tile_X7Y6_W2BEGb[7] ,
    \Tile_X7Y6_W2BEGb[6] ,
    \Tile_X7Y6_W2BEGb[5] ,
    \Tile_X7Y6_W2BEGb[4] ,
    \Tile_X7Y6_W2BEGb[3] ,
    \Tile_X7Y6_W2BEGb[2] ,
    \Tile_X7Y6_W2BEGb[1] ,
    \Tile_X7Y6_W2BEGb[0] }),
    .Tile_X0Y1_W2END({\Tile_X8Y6_W2BEGb[7] ,
    \Tile_X8Y6_W2BEGb[6] ,
    \Tile_X8Y6_W2BEGb[5] ,
    \Tile_X8Y6_W2BEGb[4] ,
    \Tile_X8Y6_W2BEGb[3] ,
    \Tile_X8Y6_W2BEGb[2] ,
    \Tile_X8Y6_W2BEGb[1] ,
    \Tile_X8Y6_W2BEGb[0] }),
    .Tile_X0Y1_W2MID({\Tile_X8Y6_W2BEG[7] ,
    \Tile_X8Y6_W2BEG[6] ,
    \Tile_X8Y6_W2BEG[5] ,
    \Tile_X8Y6_W2BEG[4] ,
    \Tile_X8Y6_W2BEG[3] ,
    \Tile_X8Y6_W2BEG[2] ,
    \Tile_X8Y6_W2BEG[1] ,
    \Tile_X8Y6_W2BEG[0] }),
    .Tile_X0Y1_W6BEG({\Tile_X7Y6_W6BEG[11] ,
    \Tile_X7Y6_W6BEG[10] ,
    \Tile_X7Y6_W6BEG[9] ,
    \Tile_X7Y6_W6BEG[8] ,
    \Tile_X7Y6_W6BEG[7] ,
    \Tile_X7Y6_W6BEG[6] ,
    \Tile_X7Y6_W6BEG[5] ,
    \Tile_X7Y6_W6BEG[4] ,
    \Tile_X7Y6_W6BEG[3] ,
    \Tile_X7Y6_W6BEG[2] ,
    \Tile_X7Y6_W6BEG[1] ,
    \Tile_X7Y6_W6BEG[0] }),
    .Tile_X0Y1_W6END({\Tile_X8Y6_W6BEG[11] ,
    \Tile_X8Y6_W6BEG[10] ,
    \Tile_X8Y6_W6BEG[9] ,
    \Tile_X8Y6_W6BEG[8] ,
    \Tile_X8Y6_W6BEG[7] ,
    \Tile_X8Y6_W6BEG[6] ,
    \Tile_X8Y6_W6BEG[5] ,
    \Tile_X8Y6_W6BEG[4] ,
    \Tile_X8Y6_W6BEG[3] ,
    \Tile_X8Y6_W6BEG[2] ,
    \Tile_X8Y6_W6BEG[1] ,
    \Tile_X8Y6_W6BEG[0] }),
    .Tile_X0Y1_WW4BEG({\Tile_X7Y6_WW4BEG[15] ,
    \Tile_X7Y6_WW4BEG[14] ,
    \Tile_X7Y6_WW4BEG[13] ,
    \Tile_X7Y6_WW4BEG[12] ,
    \Tile_X7Y6_WW4BEG[11] ,
    \Tile_X7Y6_WW4BEG[10] ,
    \Tile_X7Y6_WW4BEG[9] ,
    \Tile_X7Y6_WW4BEG[8] ,
    \Tile_X7Y6_WW4BEG[7] ,
    \Tile_X7Y6_WW4BEG[6] ,
    \Tile_X7Y6_WW4BEG[5] ,
    \Tile_X7Y6_WW4BEG[4] ,
    \Tile_X7Y6_WW4BEG[3] ,
    \Tile_X7Y6_WW4BEG[2] ,
    \Tile_X7Y6_WW4BEG[1] ,
    \Tile_X7Y6_WW4BEG[0] }),
    .Tile_X0Y1_WW4END({\Tile_X8Y6_WW4BEG[15] ,
    \Tile_X8Y6_WW4BEG[14] ,
    \Tile_X8Y6_WW4BEG[13] ,
    \Tile_X8Y6_WW4BEG[12] ,
    \Tile_X8Y6_WW4BEG[11] ,
    \Tile_X8Y6_WW4BEG[10] ,
    \Tile_X8Y6_WW4BEG[9] ,
    \Tile_X8Y6_WW4BEG[8] ,
    \Tile_X8Y6_WW4BEG[7] ,
    \Tile_X8Y6_WW4BEG[6] ,
    \Tile_X8Y6_WW4BEG[5] ,
    \Tile_X8Y6_WW4BEG[4] ,
    \Tile_X8Y6_WW4BEG[3] ,
    \Tile_X8Y6_WW4BEG[2] ,
    \Tile_X8Y6_WW4BEG[1] ,
    \Tile_X8Y6_WW4BEG[0] }));
 DSP Tile_X7Y7_DSP (.Tile_X0Y0_UserCLKo(Tile_X7Y7_UserCLKo),
    .Tile_X0Y1_UserCLK(Tile_X7Y9_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .Tile_X0Y0_E1BEG({\Tile_X7Y7_E1BEG[3] ,
    \Tile_X7Y7_E1BEG[2] ,
    \Tile_X7Y7_E1BEG[1] ,
    \Tile_X7Y7_E1BEG[0] }),
    .Tile_X0Y0_E1END({\Tile_X6Y7_E1BEG[3] ,
    \Tile_X6Y7_E1BEG[2] ,
    \Tile_X6Y7_E1BEG[1] ,
    \Tile_X6Y7_E1BEG[0] }),
    .Tile_X0Y0_E2BEG({\Tile_X7Y7_E2BEG[7] ,
    \Tile_X7Y7_E2BEG[6] ,
    \Tile_X7Y7_E2BEG[5] ,
    \Tile_X7Y7_E2BEG[4] ,
    \Tile_X7Y7_E2BEG[3] ,
    \Tile_X7Y7_E2BEG[2] ,
    \Tile_X7Y7_E2BEG[1] ,
    \Tile_X7Y7_E2BEG[0] }),
    .Tile_X0Y0_E2BEGb({\Tile_X7Y7_E2BEGb[7] ,
    \Tile_X7Y7_E2BEGb[6] ,
    \Tile_X7Y7_E2BEGb[5] ,
    \Tile_X7Y7_E2BEGb[4] ,
    \Tile_X7Y7_E2BEGb[3] ,
    \Tile_X7Y7_E2BEGb[2] ,
    \Tile_X7Y7_E2BEGb[1] ,
    \Tile_X7Y7_E2BEGb[0] }),
    .Tile_X0Y0_E2END({\Tile_X6Y7_E2BEGb[7] ,
    \Tile_X6Y7_E2BEGb[6] ,
    \Tile_X6Y7_E2BEGb[5] ,
    \Tile_X6Y7_E2BEGb[4] ,
    \Tile_X6Y7_E2BEGb[3] ,
    \Tile_X6Y7_E2BEGb[2] ,
    \Tile_X6Y7_E2BEGb[1] ,
    \Tile_X6Y7_E2BEGb[0] }),
    .Tile_X0Y0_E2MID({\Tile_X6Y7_E2BEG[7] ,
    \Tile_X6Y7_E2BEG[6] ,
    \Tile_X6Y7_E2BEG[5] ,
    \Tile_X6Y7_E2BEG[4] ,
    \Tile_X6Y7_E2BEG[3] ,
    \Tile_X6Y7_E2BEG[2] ,
    \Tile_X6Y7_E2BEG[1] ,
    \Tile_X6Y7_E2BEG[0] }),
    .Tile_X0Y0_E6BEG({\Tile_X7Y7_E6BEG[11] ,
    \Tile_X7Y7_E6BEG[10] ,
    \Tile_X7Y7_E6BEG[9] ,
    \Tile_X7Y7_E6BEG[8] ,
    \Tile_X7Y7_E6BEG[7] ,
    \Tile_X7Y7_E6BEG[6] ,
    \Tile_X7Y7_E6BEG[5] ,
    \Tile_X7Y7_E6BEG[4] ,
    \Tile_X7Y7_E6BEG[3] ,
    \Tile_X7Y7_E6BEG[2] ,
    \Tile_X7Y7_E6BEG[1] ,
    \Tile_X7Y7_E6BEG[0] }),
    .Tile_X0Y0_E6END({\Tile_X6Y7_E6BEG[11] ,
    \Tile_X6Y7_E6BEG[10] ,
    \Tile_X6Y7_E6BEG[9] ,
    \Tile_X6Y7_E6BEG[8] ,
    \Tile_X6Y7_E6BEG[7] ,
    \Tile_X6Y7_E6BEG[6] ,
    \Tile_X6Y7_E6BEG[5] ,
    \Tile_X6Y7_E6BEG[4] ,
    \Tile_X6Y7_E6BEG[3] ,
    \Tile_X6Y7_E6BEG[2] ,
    \Tile_X6Y7_E6BEG[1] ,
    \Tile_X6Y7_E6BEG[0] }),
    .Tile_X0Y0_EE4BEG({\Tile_X7Y7_EE4BEG[15] ,
    \Tile_X7Y7_EE4BEG[14] ,
    \Tile_X7Y7_EE4BEG[13] ,
    \Tile_X7Y7_EE4BEG[12] ,
    \Tile_X7Y7_EE4BEG[11] ,
    \Tile_X7Y7_EE4BEG[10] ,
    \Tile_X7Y7_EE4BEG[9] ,
    \Tile_X7Y7_EE4BEG[8] ,
    \Tile_X7Y7_EE4BEG[7] ,
    \Tile_X7Y7_EE4BEG[6] ,
    \Tile_X7Y7_EE4BEG[5] ,
    \Tile_X7Y7_EE4BEG[4] ,
    \Tile_X7Y7_EE4BEG[3] ,
    \Tile_X7Y7_EE4BEG[2] ,
    \Tile_X7Y7_EE4BEG[1] ,
    \Tile_X7Y7_EE4BEG[0] }),
    .Tile_X0Y0_EE4END({\Tile_X6Y7_EE4BEG[15] ,
    \Tile_X6Y7_EE4BEG[14] ,
    \Tile_X6Y7_EE4BEG[13] ,
    \Tile_X6Y7_EE4BEG[12] ,
    \Tile_X6Y7_EE4BEG[11] ,
    \Tile_X6Y7_EE4BEG[10] ,
    \Tile_X6Y7_EE4BEG[9] ,
    \Tile_X6Y7_EE4BEG[8] ,
    \Tile_X6Y7_EE4BEG[7] ,
    \Tile_X6Y7_EE4BEG[6] ,
    \Tile_X6Y7_EE4BEG[5] ,
    \Tile_X6Y7_EE4BEG[4] ,
    \Tile_X6Y7_EE4BEG[3] ,
    \Tile_X6Y7_EE4BEG[2] ,
    \Tile_X6Y7_EE4BEG[1] ,
    \Tile_X6Y7_EE4BEG[0] }),
    .Tile_X0Y0_FrameData({\Tile_X6Y7_FrameData_O[31] ,
    \Tile_X6Y7_FrameData_O[30] ,
    \Tile_X6Y7_FrameData_O[29] ,
    \Tile_X6Y7_FrameData_O[28] ,
    \Tile_X6Y7_FrameData_O[27] ,
    \Tile_X6Y7_FrameData_O[26] ,
    \Tile_X6Y7_FrameData_O[25] ,
    \Tile_X6Y7_FrameData_O[24] ,
    \Tile_X6Y7_FrameData_O[23] ,
    \Tile_X6Y7_FrameData_O[22] ,
    \Tile_X6Y7_FrameData_O[21] ,
    \Tile_X6Y7_FrameData_O[20] ,
    \Tile_X6Y7_FrameData_O[19] ,
    \Tile_X6Y7_FrameData_O[18] ,
    \Tile_X6Y7_FrameData_O[17] ,
    \Tile_X6Y7_FrameData_O[16] ,
    \Tile_X6Y7_FrameData_O[15] ,
    \Tile_X6Y7_FrameData_O[14] ,
    \Tile_X6Y7_FrameData_O[13] ,
    \Tile_X6Y7_FrameData_O[12] ,
    \Tile_X6Y7_FrameData_O[11] ,
    \Tile_X6Y7_FrameData_O[10] ,
    \Tile_X6Y7_FrameData_O[9] ,
    \Tile_X6Y7_FrameData_O[8] ,
    \Tile_X6Y7_FrameData_O[7] ,
    \Tile_X6Y7_FrameData_O[6] ,
    \Tile_X6Y7_FrameData_O[5] ,
    \Tile_X6Y7_FrameData_O[4] ,
    \Tile_X6Y7_FrameData_O[3] ,
    \Tile_X6Y7_FrameData_O[2] ,
    \Tile_X6Y7_FrameData_O[1] ,
    \Tile_X6Y7_FrameData_O[0] }),
    .Tile_X0Y0_FrameData_O({\Tile_X7Y7_FrameData_O[31] ,
    \Tile_X7Y7_FrameData_O[30] ,
    \Tile_X7Y7_FrameData_O[29] ,
    \Tile_X7Y7_FrameData_O[28] ,
    \Tile_X7Y7_FrameData_O[27] ,
    \Tile_X7Y7_FrameData_O[26] ,
    \Tile_X7Y7_FrameData_O[25] ,
    \Tile_X7Y7_FrameData_O[24] ,
    \Tile_X7Y7_FrameData_O[23] ,
    \Tile_X7Y7_FrameData_O[22] ,
    \Tile_X7Y7_FrameData_O[21] ,
    \Tile_X7Y7_FrameData_O[20] ,
    \Tile_X7Y7_FrameData_O[19] ,
    \Tile_X7Y7_FrameData_O[18] ,
    \Tile_X7Y7_FrameData_O[17] ,
    \Tile_X7Y7_FrameData_O[16] ,
    \Tile_X7Y7_FrameData_O[15] ,
    \Tile_X7Y7_FrameData_O[14] ,
    \Tile_X7Y7_FrameData_O[13] ,
    \Tile_X7Y7_FrameData_O[12] ,
    \Tile_X7Y7_FrameData_O[11] ,
    \Tile_X7Y7_FrameData_O[10] ,
    \Tile_X7Y7_FrameData_O[9] ,
    \Tile_X7Y7_FrameData_O[8] ,
    \Tile_X7Y7_FrameData_O[7] ,
    \Tile_X7Y7_FrameData_O[6] ,
    \Tile_X7Y7_FrameData_O[5] ,
    \Tile_X7Y7_FrameData_O[4] ,
    \Tile_X7Y7_FrameData_O[3] ,
    \Tile_X7Y7_FrameData_O[2] ,
    \Tile_X7Y7_FrameData_O[1] ,
    \Tile_X7Y7_FrameData_O[0] }),
    .Tile_X0Y0_FrameStrobe_O({\Tile_X7Y7_FrameStrobe_O[19] ,
    \Tile_X7Y7_FrameStrobe_O[18] ,
    \Tile_X7Y7_FrameStrobe_O[17] ,
    \Tile_X7Y7_FrameStrobe_O[16] ,
    \Tile_X7Y7_FrameStrobe_O[15] ,
    \Tile_X7Y7_FrameStrobe_O[14] ,
    \Tile_X7Y7_FrameStrobe_O[13] ,
    \Tile_X7Y7_FrameStrobe_O[12] ,
    \Tile_X7Y7_FrameStrobe_O[11] ,
    \Tile_X7Y7_FrameStrobe_O[10] ,
    \Tile_X7Y7_FrameStrobe_O[9] ,
    \Tile_X7Y7_FrameStrobe_O[8] ,
    \Tile_X7Y7_FrameStrobe_O[7] ,
    \Tile_X7Y7_FrameStrobe_O[6] ,
    \Tile_X7Y7_FrameStrobe_O[5] ,
    \Tile_X7Y7_FrameStrobe_O[4] ,
    \Tile_X7Y7_FrameStrobe_O[3] ,
    \Tile_X7Y7_FrameStrobe_O[2] ,
    \Tile_X7Y7_FrameStrobe_O[1] ,
    \Tile_X7Y7_FrameStrobe_O[0] }),
    .Tile_X0Y0_N1BEG({\Tile_X7Y7_N1BEG[3] ,
    \Tile_X7Y7_N1BEG[2] ,
    \Tile_X7Y7_N1BEG[1] ,
    \Tile_X7Y7_N1BEG[0] }),
    .Tile_X0Y0_N2BEG({\Tile_X7Y7_N2BEG[7] ,
    \Tile_X7Y7_N2BEG[6] ,
    \Tile_X7Y7_N2BEG[5] ,
    \Tile_X7Y7_N2BEG[4] ,
    \Tile_X7Y7_N2BEG[3] ,
    \Tile_X7Y7_N2BEG[2] ,
    \Tile_X7Y7_N2BEG[1] ,
    \Tile_X7Y7_N2BEG[0] }),
    .Tile_X0Y0_N2BEGb({\Tile_X7Y7_N2BEGb[7] ,
    \Tile_X7Y7_N2BEGb[6] ,
    \Tile_X7Y7_N2BEGb[5] ,
    \Tile_X7Y7_N2BEGb[4] ,
    \Tile_X7Y7_N2BEGb[3] ,
    \Tile_X7Y7_N2BEGb[2] ,
    \Tile_X7Y7_N2BEGb[1] ,
    \Tile_X7Y7_N2BEGb[0] }),
    .Tile_X0Y0_N4BEG({\Tile_X7Y7_N4BEG[15] ,
    \Tile_X7Y7_N4BEG[14] ,
    \Tile_X7Y7_N4BEG[13] ,
    \Tile_X7Y7_N4BEG[12] ,
    \Tile_X7Y7_N4BEG[11] ,
    \Tile_X7Y7_N4BEG[10] ,
    \Tile_X7Y7_N4BEG[9] ,
    \Tile_X7Y7_N4BEG[8] ,
    \Tile_X7Y7_N4BEG[7] ,
    \Tile_X7Y7_N4BEG[6] ,
    \Tile_X7Y7_N4BEG[5] ,
    \Tile_X7Y7_N4BEG[4] ,
    \Tile_X7Y7_N4BEG[3] ,
    \Tile_X7Y7_N4BEG[2] ,
    \Tile_X7Y7_N4BEG[1] ,
    \Tile_X7Y7_N4BEG[0] }),
    .Tile_X0Y0_NN4BEG({\Tile_X7Y7_NN4BEG[15] ,
    \Tile_X7Y7_NN4BEG[14] ,
    \Tile_X7Y7_NN4BEG[13] ,
    \Tile_X7Y7_NN4BEG[12] ,
    \Tile_X7Y7_NN4BEG[11] ,
    \Tile_X7Y7_NN4BEG[10] ,
    \Tile_X7Y7_NN4BEG[9] ,
    \Tile_X7Y7_NN4BEG[8] ,
    \Tile_X7Y7_NN4BEG[7] ,
    \Tile_X7Y7_NN4BEG[6] ,
    \Tile_X7Y7_NN4BEG[5] ,
    \Tile_X7Y7_NN4BEG[4] ,
    \Tile_X7Y7_NN4BEG[3] ,
    \Tile_X7Y7_NN4BEG[2] ,
    \Tile_X7Y7_NN4BEG[1] ,
    \Tile_X7Y7_NN4BEG[0] }),
    .Tile_X0Y0_S1END({\Tile_X7Y6_S1BEG[3] ,
    \Tile_X7Y6_S1BEG[2] ,
    \Tile_X7Y6_S1BEG[1] ,
    \Tile_X7Y6_S1BEG[0] }),
    .Tile_X0Y0_S2END({\Tile_X7Y6_S2BEGb[7] ,
    \Tile_X7Y6_S2BEGb[6] ,
    \Tile_X7Y6_S2BEGb[5] ,
    \Tile_X7Y6_S2BEGb[4] ,
    \Tile_X7Y6_S2BEGb[3] ,
    \Tile_X7Y6_S2BEGb[2] ,
    \Tile_X7Y6_S2BEGb[1] ,
    \Tile_X7Y6_S2BEGb[0] }),
    .Tile_X0Y0_S2MID({\Tile_X7Y6_S2BEG[7] ,
    \Tile_X7Y6_S2BEG[6] ,
    \Tile_X7Y6_S2BEG[5] ,
    \Tile_X7Y6_S2BEG[4] ,
    \Tile_X7Y6_S2BEG[3] ,
    \Tile_X7Y6_S2BEG[2] ,
    \Tile_X7Y6_S2BEG[1] ,
    \Tile_X7Y6_S2BEG[0] }),
    .Tile_X0Y0_S4END({\Tile_X7Y6_S4BEG[15] ,
    \Tile_X7Y6_S4BEG[14] ,
    \Tile_X7Y6_S4BEG[13] ,
    \Tile_X7Y6_S4BEG[12] ,
    \Tile_X7Y6_S4BEG[11] ,
    \Tile_X7Y6_S4BEG[10] ,
    \Tile_X7Y6_S4BEG[9] ,
    \Tile_X7Y6_S4BEG[8] ,
    \Tile_X7Y6_S4BEG[7] ,
    \Tile_X7Y6_S4BEG[6] ,
    \Tile_X7Y6_S4BEG[5] ,
    \Tile_X7Y6_S4BEG[4] ,
    \Tile_X7Y6_S4BEG[3] ,
    \Tile_X7Y6_S4BEG[2] ,
    \Tile_X7Y6_S4BEG[1] ,
    \Tile_X7Y6_S4BEG[0] }),
    .Tile_X0Y0_SS4END({\Tile_X7Y6_SS4BEG[15] ,
    \Tile_X7Y6_SS4BEG[14] ,
    \Tile_X7Y6_SS4BEG[13] ,
    \Tile_X7Y6_SS4BEG[12] ,
    \Tile_X7Y6_SS4BEG[11] ,
    \Tile_X7Y6_SS4BEG[10] ,
    \Tile_X7Y6_SS4BEG[9] ,
    \Tile_X7Y6_SS4BEG[8] ,
    \Tile_X7Y6_SS4BEG[7] ,
    \Tile_X7Y6_SS4BEG[6] ,
    \Tile_X7Y6_SS4BEG[5] ,
    \Tile_X7Y6_SS4BEG[4] ,
    \Tile_X7Y6_SS4BEG[3] ,
    \Tile_X7Y6_SS4BEG[2] ,
    \Tile_X7Y6_SS4BEG[1] ,
    \Tile_X7Y6_SS4BEG[0] }),
    .Tile_X0Y0_W1BEG({\Tile_X7Y7_W1BEG[3] ,
    \Tile_X7Y7_W1BEG[2] ,
    \Tile_X7Y7_W1BEG[1] ,
    \Tile_X7Y7_W1BEG[0] }),
    .Tile_X0Y0_W1END({\Tile_X8Y7_W1BEG[3] ,
    \Tile_X8Y7_W1BEG[2] ,
    \Tile_X8Y7_W1BEG[1] ,
    \Tile_X8Y7_W1BEG[0] }),
    .Tile_X0Y0_W2BEG({\Tile_X7Y7_W2BEG[7] ,
    \Tile_X7Y7_W2BEG[6] ,
    \Tile_X7Y7_W2BEG[5] ,
    \Tile_X7Y7_W2BEG[4] ,
    \Tile_X7Y7_W2BEG[3] ,
    \Tile_X7Y7_W2BEG[2] ,
    \Tile_X7Y7_W2BEG[1] ,
    \Tile_X7Y7_W2BEG[0] }),
    .Tile_X0Y0_W2BEGb({\Tile_X7Y7_W2BEGb[7] ,
    \Tile_X7Y7_W2BEGb[6] ,
    \Tile_X7Y7_W2BEGb[5] ,
    \Tile_X7Y7_W2BEGb[4] ,
    \Tile_X7Y7_W2BEGb[3] ,
    \Tile_X7Y7_W2BEGb[2] ,
    \Tile_X7Y7_W2BEGb[1] ,
    \Tile_X7Y7_W2BEGb[0] }),
    .Tile_X0Y0_W2END({\Tile_X8Y7_W2BEGb[7] ,
    \Tile_X8Y7_W2BEGb[6] ,
    \Tile_X8Y7_W2BEGb[5] ,
    \Tile_X8Y7_W2BEGb[4] ,
    \Tile_X8Y7_W2BEGb[3] ,
    \Tile_X8Y7_W2BEGb[2] ,
    \Tile_X8Y7_W2BEGb[1] ,
    \Tile_X8Y7_W2BEGb[0] }),
    .Tile_X0Y0_W2MID({\Tile_X8Y7_W2BEG[7] ,
    \Tile_X8Y7_W2BEG[6] ,
    \Tile_X8Y7_W2BEG[5] ,
    \Tile_X8Y7_W2BEG[4] ,
    \Tile_X8Y7_W2BEG[3] ,
    \Tile_X8Y7_W2BEG[2] ,
    \Tile_X8Y7_W2BEG[1] ,
    \Tile_X8Y7_W2BEG[0] }),
    .Tile_X0Y0_W6BEG({\Tile_X7Y7_W6BEG[11] ,
    \Tile_X7Y7_W6BEG[10] ,
    \Tile_X7Y7_W6BEG[9] ,
    \Tile_X7Y7_W6BEG[8] ,
    \Tile_X7Y7_W6BEG[7] ,
    \Tile_X7Y7_W6BEG[6] ,
    \Tile_X7Y7_W6BEG[5] ,
    \Tile_X7Y7_W6BEG[4] ,
    \Tile_X7Y7_W6BEG[3] ,
    \Tile_X7Y7_W6BEG[2] ,
    \Tile_X7Y7_W6BEG[1] ,
    \Tile_X7Y7_W6BEG[0] }),
    .Tile_X0Y0_W6END({\Tile_X8Y7_W6BEG[11] ,
    \Tile_X8Y7_W6BEG[10] ,
    \Tile_X8Y7_W6BEG[9] ,
    \Tile_X8Y7_W6BEG[8] ,
    \Tile_X8Y7_W6BEG[7] ,
    \Tile_X8Y7_W6BEG[6] ,
    \Tile_X8Y7_W6BEG[5] ,
    \Tile_X8Y7_W6BEG[4] ,
    \Tile_X8Y7_W6BEG[3] ,
    \Tile_X8Y7_W6BEG[2] ,
    \Tile_X8Y7_W6BEG[1] ,
    \Tile_X8Y7_W6BEG[0] }),
    .Tile_X0Y0_WW4BEG({\Tile_X7Y7_WW4BEG[15] ,
    \Tile_X7Y7_WW4BEG[14] ,
    \Tile_X7Y7_WW4BEG[13] ,
    \Tile_X7Y7_WW4BEG[12] ,
    \Tile_X7Y7_WW4BEG[11] ,
    \Tile_X7Y7_WW4BEG[10] ,
    \Tile_X7Y7_WW4BEG[9] ,
    \Tile_X7Y7_WW4BEG[8] ,
    \Tile_X7Y7_WW4BEG[7] ,
    \Tile_X7Y7_WW4BEG[6] ,
    \Tile_X7Y7_WW4BEG[5] ,
    \Tile_X7Y7_WW4BEG[4] ,
    \Tile_X7Y7_WW4BEG[3] ,
    \Tile_X7Y7_WW4BEG[2] ,
    \Tile_X7Y7_WW4BEG[1] ,
    \Tile_X7Y7_WW4BEG[0] }),
    .Tile_X0Y0_WW4END({\Tile_X8Y7_WW4BEG[15] ,
    \Tile_X8Y7_WW4BEG[14] ,
    \Tile_X8Y7_WW4BEG[13] ,
    \Tile_X8Y7_WW4BEG[12] ,
    \Tile_X8Y7_WW4BEG[11] ,
    \Tile_X8Y7_WW4BEG[10] ,
    \Tile_X8Y7_WW4BEG[9] ,
    \Tile_X8Y7_WW4BEG[8] ,
    \Tile_X8Y7_WW4BEG[7] ,
    \Tile_X8Y7_WW4BEG[6] ,
    \Tile_X8Y7_WW4BEG[5] ,
    \Tile_X8Y7_WW4BEG[4] ,
    \Tile_X8Y7_WW4BEG[3] ,
    \Tile_X8Y7_WW4BEG[2] ,
    \Tile_X8Y7_WW4BEG[1] ,
    \Tile_X8Y7_WW4BEG[0] }),
    .Tile_X0Y1_E1BEG({\Tile_X7Y8_E1BEG[3] ,
    \Tile_X7Y8_E1BEG[2] ,
    \Tile_X7Y8_E1BEG[1] ,
    \Tile_X7Y8_E1BEG[0] }),
    .Tile_X0Y1_E1END({\Tile_X6Y8_E1BEG[3] ,
    \Tile_X6Y8_E1BEG[2] ,
    \Tile_X6Y8_E1BEG[1] ,
    \Tile_X6Y8_E1BEG[0] }),
    .Tile_X0Y1_E2BEG({\Tile_X7Y8_E2BEG[7] ,
    \Tile_X7Y8_E2BEG[6] ,
    \Tile_X7Y8_E2BEG[5] ,
    \Tile_X7Y8_E2BEG[4] ,
    \Tile_X7Y8_E2BEG[3] ,
    \Tile_X7Y8_E2BEG[2] ,
    \Tile_X7Y8_E2BEG[1] ,
    \Tile_X7Y8_E2BEG[0] }),
    .Tile_X0Y1_E2BEGb({\Tile_X7Y8_E2BEGb[7] ,
    \Tile_X7Y8_E2BEGb[6] ,
    \Tile_X7Y8_E2BEGb[5] ,
    \Tile_X7Y8_E2BEGb[4] ,
    \Tile_X7Y8_E2BEGb[3] ,
    \Tile_X7Y8_E2BEGb[2] ,
    \Tile_X7Y8_E2BEGb[1] ,
    \Tile_X7Y8_E2BEGb[0] }),
    .Tile_X0Y1_E2END({\Tile_X6Y8_E2BEGb[7] ,
    \Tile_X6Y8_E2BEGb[6] ,
    \Tile_X6Y8_E2BEGb[5] ,
    \Tile_X6Y8_E2BEGb[4] ,
    \Tile_X6Y8_E2BEGb[3] ,
    \Tile_X6Y8_E2BEGb[2] ,
    \Tile_X6Y8_E2BEGb[1] ,
    \Tile_X6Y8_E2BEGb[0] }),
    .Tile_X0Y1_E2MID({\Tile_X6Y8_E2BEG[7] ,
    \Tile_X6Y8_E2BEG[6] ,
    \Tile_X6Y8_E2BEG[5] ,
    \Tile_X6Y8_E2BEG[4] ,
    \Tile_X6Y8_E2BEG[3] ,
    \Tile_X6Y8_E2BEG[2] ,
    \Tile_X6Y8_E2BEG[1] ,
    \Tile_X6Y8_E2BEG[0] }),
    .Tile_X0Y1_E6BEG({\Tile_X7Y8_E6BEG[11] ,
    \Tile_X7Y8_E6BEG[10] ,
    \Tile_X7Y8_E6BEG[9] ,
    \Tile_X7Y8_E6BEG[8] ,
    \Tile_X7Y8_E6BEG[7] ,
    \Tile_X7Y8_E6BEG[6] ,
    \Tile_X7Y8_E6BEG[5] ,
    \Tile_X7Y8_E6BEG[4] ,
    \Tile_X7Y8_E6BEG[3] ,
    \Tile_X7Y8_E6BEG[2] ,
    \Tile_X7Y8_E6BEG[1] ,
    \Tile_X7Y8_E6BEG[0] }),
    .Tile_X0Y1_E6END({\Tile_X6Y8_E6BEG[11] ,
    \Tile_X6Y8_E6BEG[10] ,
    \Tile_X6Y8_E6BEG[9] ,
    \Tile_X6Y8_E6BEG[8] ,
    \Tile_X6Y8_E6BEG[7] ,
    \Tile_X6Y8_E6BEG[6] ,
    \Tile_X6Y8_E6BEG[5] ,
    \Tile_X6Y8_E6BEG[4] ,
    \Tile_X6Y8_E6BEG[3] ,
    \Tile_X6Y8_E6BEG[2] ,
    \Tile_X6Y8_E6BEG[1] ,
    \Tile_X6Y8_E6BEG[0] }),
    .Tile_X0Y1_EE4BEG({\Tile_X7Y8_EE4BEG[15] ,
    \Tile_X7Y8_EE4BEG[14] ,
    \Tile_X7Y8_EE4BEG[13] ,
    \Tile_X7Y8_EE4BEG[12] ,
    \Tile_X7Y8_EE4BEG[11] ,
    \Tile_X7Y8_EE4BEG[10] ,
    \Tile_X7Y8_EE4BEG[9] ,
    \Tile_X7Y8_EE4BEG[8] ,
    \Tile_X7Y8_EE4BEG[7] ,
    \Tile_X7Y8_EE4BEG[6] ,
    \Tile_X7Y8_EE4BEG[5] ,
    \Tile_X7Y8_EE4BEG[4] ,
    \Tile_X7Y8_EE4BEG[3] ,
    \Tile_X7Y8_EE4BEG[2] ,
    \Tile_X7Y8_EE4BEG[1] ,
    \Tile_X7Y8_EE4BEG[0] }),
    .Tile_X0Y1_EE4END({\Tile_X6Y8_EE4BEG[15] ,
    \Tile_X6Y8_EE4BEG[14] ,
    \Tile_X6Y8_EE4BEG[13] ,
    \Tile_X6Y8_EE4BEG[12] ,
    \Tile_X6Y8_EE4BEG[11] ,
    \Tile_X6Y8_EE4BEG[10] ,
    \Tile_X6Y8_EE4BEG[9] ,
    \Tile_X6Y8_EE4BEG[8] ,
    \Tile_X6Y8_EE4BEG[7] ,
    \Tile_X6Y8_EE4BEG[6] ,
    \Tile_X6Y8_EE4BEG[5] ,
    \Tile_X6Y8_EE4BEG[4] ,
    \Tile_X6Y8_EE4BEG[3] ,
    \Tile_X6Y8_EE4BEG[2] ,
    \Tile_X6Y8_EE4BEG[1] ,
    \Tile_X6Y8_EE4BEG[0] }),
    .Tile_X0Y1_FrameData({\Tile_X6Y8_FrameData_O[31] ,
    \Tile_X6Y8_FrameData_O[30] ,
    \Tile_X6Y8_FrameData_O[29] ,
    \Tile_X6Y8_FrameData_O[28] ,
    \Tile_X6Y8_FrameData_O[27] ,
    \Tile_X6Y8_FrameData_O[26] ,
    \Tile_X6Y8_FrameData_O[25] ,
    \Tile_X6Y8_FrameData_O[24] ,
    \Tile_X6Y8_FrameData_O[23] ,
    \Tile_X6Y8_FrameData_O[22] ,
    \Tile_X6Y8_FrameData_O[21] ,
    \Tile_X6Y8_FrameData_O[20] ,
    \Tile_X6Y8_FrameData_O[19] ,
    \Tile_X6Y8_FrameData_O[18] ,
    \Tile_X6Y8_FrameData_O[17] ,
    \Tile_X6Y8_FrameData_O[16] ,
    \Tile_X6Y8_FrameData_O[15] ,
    \Tile_X6Y8_FrameData_O[14] ,
    \Tile_X6Y8_FrameData_O[13] ,
    \Tile_X6Y8_FrameData_O[12] ,
    \Tile_X6Y8_FrameData_O[11] ,
    \Tile_X6Y8_FrameData_O[10] ,
    \Tile_X6Y8_FrameData_O[9] ,
    \Tile_X6Y8_FrameData_O[8] ,
    \Tile_X6Y8_FrameData_O[7] ,
    \Tile_X6Y8_FrameData_O[6] ,
    \Tile_X6Y8_FrameData_O[5] ,
    \Tile_X6Y8_FrameData_O[4] ,
    \Tile_X6Y8_FrameData_O[3] ,
    \Tile_X6Y8_FrameData_O[2] ,
    \Tile_X6Y8_FrameData_O[1] ,
    \Tile_X6Y8_FrameData_O[0] }),
    .Tile_X0Y1_FrameData_O({\Tile_X7Y8_FrameData_O[31] ,
    \Tile_X7Y8_FrameData_O[30] ,
    \Tile_X7Y8_FrameData_O[29] ,
    \Tile_X7Y8_FrameData_O[28] ,
    \Tile_X7Y8_FrameData_O[27] ,
    \Tile_X7Y8_FrameData_O[26] ,
    \Tile_X7Y8_FrameData_O[25] ,
    \Tile_X7Y8_FrameData_O[24] ,
    \Tile_X7Y8_FrameData_O[23] ,
    \Tile_X7Y8_FrameData_O[22] ,
    \Tile_X7Y8_FrameData_O[21] ,
    \Tile_X7Y8_FrameData_O[20] ,
    \Tile_X7Y8_FrameData_O[19] ,
    \Tile_X7Y8_FrameData_O[18] ,
    \Tile_X7Y8_FrameData_O[17] ,
    \Tile_X7Y8_FrameData_O[16] ,
    \Tile_X7Y8_FrameData_O[15] ,
    \Tile_X7Y8_FrameData_O[14] ,
    \Tile_X7Y8_FrameData_O[13] ,
    \Tile_X7Y8_FrameData_O[12] ,
    \Tile_X7Y8_FrameData_O[11] ,
    \Tile_X7Y8_FrameData_O[10] ,
    \Tile_X7Y8_FrameData_O[9] ,
    \Tile_X7Y8_FrameData_O[8] ,
    \Tile_X7Y8_FrameData_O[7] ,
    \Tile_X7Y8_FrameData_O[6] ,
    \Tile_X7Y8_FrameData_O[5] ,
    \Tile_X7Y8_FrameData_O[4] ,
    \Tile_X7Y8_FrameData_O[3] ,
    \Tile_X7Y8_FrameData_O[2] ,
    \Tile_X7Y8_FrameData_O[1] ,
    \Tile_X7Y8_FrameData_O[0] }),
    .Tile_X0Y1_FrameStrobe({\Tile_X7Y9_FrameStrobe_O[19] ,
    \Tile_X7Y9_FrameStrobe_O[18] ,
    \Tile_X7Y9_FrameStrobe_O[17] ,
    \Tile_X7Y9_FrameStrobe_O[16] ,
    \Tile_X7Y9_FrameStrobe_O[15] ,
    \Tile_X7Y9_FrameStrobe_O[14] ,
    \Tile_X7Y9_FrameStrobe_O[13] ,
    \Tile_X7Y9_FrameStrobe_O[12] ,
    \Tile_X7Y9_FrameStrobe_O[11] ,
    \Tile_X7Y9_FrameStrobe_O[10] ,
    \Tile_X7Y9_FrameStrobe_O[9] ,
    \Tile_X7Y9_FrameStrobe_O[8] ,
    \Tile_X7Y9_FrameStrobe_O[7] ,
    \Tile_X7Y9_FrameStrobe_O[6] ,
    \Tile_X7Y9_FrameStrobe_O[5] ,
    \Tile_X7Y9_FrameStrobe_O[4] ,
    \Tile_X7Y9_FrameStrobe_O[3] ,
    \Tile_X7Y9_FrameStrobe_O[2] ,
    \Tile_X7Y9_FrameStrobe_O[1] ,
    \Tile_X7Y9_FrameStrobe_O[0] }),
    .Tile_X0Y1_N1END({\Tile_X7Y9_N1BEG[3] ,
    \Tile_X7Y9_N1BEG[2] ,
    \Tile_X7Y9_N1BEG[1] ,
    \Tile_X7Y9_N1BEG[0] }),
    .Tile_X0Y1_N2END({\Tile_X7Y9_N2BEGb[7] ,
    \Tile_X7Y9_N2BEGb[6] ,
    \Tile_X7Y9_N2BEGb[5] ,
    \Tile_X7Y9_N2BEGb[4] ,
    \Tile_X7Y9_N2BEGb[3] ,
    \Tile_X7Y9_N2BEGb[2] ,
    \Tile_X7Y9_N2BEGb[1] ,
    \Tile_X7Y9_N2BEGb[0] }),
    .Tile_X0Y1_N2MID({\Tile_X7Y9_N2BEG[7] ,
    \Tile_X7Y9_N2BEG[6] ,
    \Tile_X7Y9_N2BEG[5] ,
    \Tile_X7Y9_N2BEG[4] ,
    \Tile_X7Y9_N2BEG[3] ,
    \Tile_X7Y9_N2BEG[2] ,
    \Tile_X7Y9_N2BEG[1] ,
    \Tile_X7Y9_N2BEG[0] }),
    .Tile_X0Y1_N4END({\Tile_X7Y9_N4BEG[15] ,
    \Tile_X7Y9_N4BEG[14] ,
    \Tile_X7Y9_N4BEG[13] ,
    \Tile_X7Y9_N4BEG[12] ,
    \Tile_X7Y9_N4BEG[11] ,
    \Tile_X7Y9_N4BEG[10] ,
    \Tile_X7Y9_N4BEG[9] ,
    \Tile_X7Y9_N4BEG[8] ,
    \Tile_X7Y9_N4BEG[7] ,
    \Tile_X7Y9_N4BEG[6] ,
    \Tile_X7Y9_N4BEG[5] ,
    \Tile_X7Y9_N4BEG[4] ,
    \Tile_X7Y9_N4BEG[3] ,
    \Tile_X7Y9_N4BEG[2] ,
    \Tile_X7Y9_N4BEG[1] ,
    \Tile_X7Y9_N4BEG[0] }),
    .Tile_X0Y1_NN4END({\Tile_X7Y9_NN4BEG[15] ,
    \Tile_X7Y9_NN4BEG[14] ,
    \Tile_X7Y9_NN4BEG[13] ,
    \Tile_X7Y9_NN4BEG[12] ,
    \Tile_X7Y9_NN4BEG[11] ,
    \Tile_X7Y9_NN4BEG[10] ,
    \Tile_X7Y9_NN4BEG[9] ,
    \Tile_X7Y9_NN4BEG[8] ,
    \Tile_X7Y9_NN4BEG[7] ,
    \Tile_X7Y9_NN4BEG[6] ,
    \Tile_X7Y9_NN4BEG[5] ,
    \Tile_X7Y9_NN4BEG[4] ,
    \Tile_X7Y9_NN4BEG[3] ,
    \Tile_X7Y9_NN4BEG[2] ,
    \Tile_X7Y9_NN4BEG[1] ,
    \Tile_X7Y9_NN4BEG[0] }),
    .Tile_X0Y1_S1BEG({\Tile_X7Y8_S1BEG[3] ,
    \Tile_X7Y8_S1BEG[2] ,
    \Tile_X7Y8_S1BEG[1] ,
    \Tile_X7Y8_S1BEG[0] }),
    .Tile_X0Y1_S2BEG({\Tile_X7Y8_S2BEG[7] ,
    \Tile_X7Y8_S2BEG[6] ,
    \Tile_X7Y8_S2BEG[5] ,
    \Tile_X7Y8_S2BEG[4] ,
    \Tile_X7Y8_S2BEG[3] ,
    \Tile_X7Y8_S2BEG[2] ,
    \Tile_X7Y8_S2BEG[1] ,
    \Tile_X7Y8_S2BEG[0] }),
    .Tile_X0Y1_S2BEGb({\Tile_X7Y8_S2BEGb[7] ,
    \Tile_X7Y8_S2BEGb[6] ,
    \Tile_X7Y8_S2BEGb[5] ,
    \Tile_X7Y8_S2BEGb[4] ,
    \Tile_X7Y8_S2BEGb[3] ,
    \Tile_X7Y8_S2BEGb[2] ,
    \Tile_X7Y8_S2BEGb[1] ,
    \Tile_X7Y8_S2BEGb[0] }),
    .Tile_X0Y1_S4BEG({\Tile_X7Y8_S4BEG[15] ,
    \Tile_X7Y8_S4BEG[14] ,
    \Tile_X7Y8_S4BEG[13] ,
    \Tile_X7Y8_S4BEG[12] ,
    \Tile_X7Y8_S4BEG[11] ,
    \Tile_X7Y8_S4BEG[10] ,
    \Tile_X7Y8_S4BEG[9] ,
    \Tile_X7Y8_S4BEG[8] ,
    \Tile_X7Y8_S4BEG[7] ,
    \Tile_X7Y8_S4BEG[6] ,
    \Tile_X7Y8_S4BEG[5] ,
    \Tile_X7Y8_S4BEG[4] ,
    \Tile_X7Y8_S4BEG[3] ,
    \Tile_X7Y8_S4BEG[2] ,
    \Tile_X7Y8_S4BEG[1] ,
    \Tile_X7Y8_S4BEG[0] }),
    .Tile_X0Y1_SS4BEG({\Tile_X7Y8_SS4BEG[15] ,
    \Tile_X7Y8_SS4BEG[14] ,
    \Tile_X7Y8_SS4BEG[13] ,
    \Tile_X7Y8_SS4BEG[12] ,
    \Tile_X7Y8_SS4BEG[11] ,
    \Tile_X7Y8_SS4BEG[10] ,
    \Tile_X7Y8_SS4BEG[9] ,
    \Tile_X7Y8_SS4BEG[8] ,
    \Tile_X7Y8_SS4BEG[7] ,
    \Tile_X7Y8_SS4BEG[6] ,
    \Tile_X7Y8_SS4BEG[5] ,
    \Tile_X7Y8_SS4BEG[4] ,
    \Tile_X7Y8_SS4BEG[3] ,
    \Tile_X7Y8_SS4BEG[2] ,
    \Tile_X7Y8_SS4BEG[1] ,
    \Tile_X7Y8_SS4BEG[0] }),
    .Tile_X0Y1_W1BEG({\Tile_X7Y8_W1BEG[3] ,
    \Tile_X7Y8_W1BEG[2] ,
    \Tile_X7Y8_W1BEG[1] ,
    \Tile_X7Y8_W1BEG[0] }),
    .Tile_X0Y1_W1END({\Tile_X8Y8_W1BEG[3] ,
    \Tile_X8Y8_W1BEG[2] ,
    \Tile_X8Y8_W1BEG[1] ,
    \Tile_X8Y8_W1BEG[0] }),
    .Tile_X0Y1_W2BEG({\Tile_X7Y8_W2BEG[7] ,
    \Tile_X7Y8_W2BEG[6] ,
    \Tile_X7Y8_W2BEG[5] ,
    \Tile_X7Y8_W2BEG[4] ,
    \Tile_X7Y8_W2BEG[3] ,
    \Tile_X7Y8_W2BEG[2] ,
    \Tile_X7Y8_W2BEG[1] ,
    \Tile_X7Y8_W2BEG[0] }),
    .Tile_X0Y1_W2BEGb({\Tile_X7Y8_W2BEGb[7] ,
    \Tile_X7Y8_W2BEGb[6] ,
    \Tile_X7Y8_W2BEGb[5] ,
    \Tile_X7Y8_W2BEGb[4] ,
    \Tile_X7Y8_W2BEGb[3] ,
    \Tile_X7Y8_W2BEGb[2] ,
    \Tile_X7Y8_W2BEGb[1] ,
    \Tile_X7Y8_W2BEGb[0] }),
    .Tile_X0Y1_W2END({\Tile_X8Y8_W2BEGb[7] ,
    \Tile_X8Y8_W2BEGb[6] ,
    \Tile_X8Y8_W2BEGb[5] ,
    \Tile_X8Y8_W2BEGb[4] ,
    \Tile_X8Y8_W2BEGb[3] ,
    \Tile_X8Y8_W2BEGb[2] ,
    \Tile_X8Y8_W2BEGb[1] ,
    \Tile_X8Y8_W2BEGb[0] }),
    .Tile_X0Y1_W2MID({\Tile_X8Y8_W2BEG[7] ,
    \Tile_X8Y8_W2BEG[6] ,
    \Tile_X8Y8_W2BEG[5] ,
    \Tile_X8Y8_W2BEG[4] ,
    \Tile_X8Y8_W2BEG[3] ,
    \Tile_X8Y8_W2BEG[2] ,
    \Tile_X8Y8_W2BEG[1] ,
    \Tile_X8Y8_W2BEG[0] }),
    .Tile_X0Y1_W6BEG({\Tile_X7Y8_W6BEG[11] ,
    \Tile_X7Y8_W6BEG[10] ,
    \Tile_X7Y8_W6BEG[9] ,
    \Tile_X7Y8_W6BEG[8] ,
    \Tile_X7Y8_W6BEG[7] ,
    \Tile_X7Y8_W6BEG[6] ,
    \Tile_X7Y8_W6BEG[5] ,
    \Tile_X7Y8_W6BEG[4] ,
    \Tile_X7Y8_W6BEG[3] ,
    \Tile_X7Y8_W6BEG[2] ,
    \Tile_X7Y8_W6BEG[1] ,
    \Tile_X7Y8_W6BEG[0] }),
    .Tile_X0Y1_W6END({\Tile_X8Y8_W6BEG[11] ,
    \Tile_X8Y8_W6BEG[10] ,
    \Tile_X8Y8_W6BEG[9] ,
    \Tile_X8Y8_W6BEG[8] ,
    \Tile_X8Y8_W6BEG[7] ,
    \Tile_X8Y8_W6BEG[6] ,
    \Tile_X8Y8_W6BEG[5] ,
    \Tile_X8Y8_W6BEG[4] ,
    \Tile_X8Y8_W6BEG[3] ,
    \Tile_X8Y8_W6BEG[2] ,
    \Tile_X8Y8_W6BEG[1] ,
    \Tile_X8Y8_W6BEG[0] }),
    .Tile_X0Y1_WW4BEG({\Tile_X7Y8_WW4BEG[15] ,
    \Tile_X7Y8_WW4BEG[14] ,
    \Tile_X7Y8_WW4BEG[13] ,
    \Tile_X7Y8_WW4BEG[12] ,
    \Tile_X7Y8_WW4BEG[11] ,
    \Tile_X7Y8_WW4BEG[10] ,
    \Tile_X7Y8_WW4BEG[9] ,
    \Tile_X7Y8_WW4BEG[8] ,
    \Tile_X7Y8_WW4BEG[7] ,
    \Tile_X7Y8_WW4BEG[6] ,
    \Tile_X7Y8_WW4BEG[5] ,
    \Tile_X7Y8_WW4BEG[4] ,
    \Tile_X7Y8_WW4BEG[3] ,
    \Tile_X7Y8_WW4BEG[2] ,
    \Tile_X7Y8_WW4BEG[1] ,
    \Tile_X7Y8_WW4BEG[0] }),
    .Tile_X0Y1_WW4END({\Tile_X8Y8_WW4BEG[15] ,
    \Tile_X8Y8_WW4BEG[14] ,
    \Tile_X8Y8_WW4BEG[13] ,
    \Tile_X8Y8_WW4BEG[12] ,
    \Tile_X8Y8_WW4BEG[11] ,
    \Tile_X8Y8_WW4BEG[10] ,
    \Tile_X8Y8_WW4BEG[9] ,
    \Tile_X8Y8_WW4BEG[8] ,
    \Tile_X8Y8_WW4BEG[7] ,
    \Tile_X8Y8_WW4BEG[6] ,
    \Tile_X8Y8_WW4BEG[5] ,
    \Tile_X8Y8_WW4BEG[4] ,
    \Tile_X8Y8_WW4BEG[3] ,
    \Tile_X8Y8_WW4BEG[2] ,
    \Tile_X8Y8_WW4BEG[1] ,
    \Tile_X8Y8_WW4BEG[0] }));
 DSP Tile_X7Y9_DSP (.Tile_X0Y0_UserCLKo(Tile_X7Y9_UserCLKo),
    .Tile_X0Y1_UserCLK(Tile_X7Y11_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .Tile_X0Y0_E1BEG({\Tile_X7Y9_E1BEG[3] ,
    \Tile_X7Y9_E1BEG[2] ,
    \Tile_X7Y9_E1BEG[1] ,
    \Tile_X7Y9_E1BEG[0] }),
    .Tile_X0Y0_E1END({\Tile_X6Y9_E1BEG[3] ,
    \Tile_X6Y9_E1BEG[2] ,
    \Tile_X6Y9_E1BEG[1] ,
    \Tile_X6Y9_E1BEG[0] }),
    .Tile_X0Y0_E2BEG({\Tile_X7Y9_E2BEG[7] ,
    \Tile_X7Y9_E2BEG[6] ,
    \Tile_X7Y9_E2BEG[5] ,
    \Tile_X7Y9_E2BEG[4] ,
    \Tile_X7Y9_E2BEG[3] ,
    \Tile_X7Y9_E2BEG[2] ,
    \Tile_X7Y9_E2BEG[1] ,
    \Tile_X7Y9_E2BEG[0] }),
    .Tile_X0Y0_E2BEGb({\Tile_X7Y9_E2BEGb[7] ,
    \Tile_X7Y9_E2BEGb[6] ,
    \Tile_X7Y9_E2BEGb[5] ,
    \Tile_X7Y9_E2BEGb[4] ,
    \Tile_X7Y9_E2BEGb[3] ,
    \Tile_X7Y9_E2BEGb[2] ,
    \Tile_X7Y9_E2BEGb[1] ,
    \Tile_X7Y9_E2BEGb[0] }),
    .Tile_X0Y0_E2END({\Tile_X6Y9_E2BEGb[7] ,
    \Tile_X6Y9_E2BEGb[6] ,
    \Tile_X6Y9_E2BEGb[5] ,
    \Tile_X6Y9_E2BEGb[4] ,
    \Tile_X6Y9_E2BEGb[3] ,
    \Tile_X6Y9_E2BEGb[2] ,
    \Tile_X6Y9_E2BEGb[1] ,
    \Tile_X6Y9_E2BEGb[0] }),
    .Tile_X0Y0_E2MID({\Tile_X6Y9_E2BEG[7] ,
    \Tile_X6Y9_E2BEG[6] ,
    \Tile_X6Y9_E2BEG[5] ,
    \Tile_X6Y9_E2BEG[4] ,
    \Tile_X6Y9_E2BEG[3] ,
    \Tile_X6Y9_E2BEG[2] ,
    \Tile_X6Y9_E2BEG[1] ,
    \Tile_X6Y9_E2BEG[0] }),
    .Tile_X0Y0_E6BEG({\Tile_X7Y9_E6BEG[11] ,
    \Tile_X7Y9_E6BEG[10] ,
    \Tile_X7Y9_E6BEG[9] ,
    \Tile_X7Y9_E6BEG[8] ,
    \Tile_X7Y9_E6BEG[7] ,
    \Tile_X7Y9_E6BEG[6] ,
    \Tile_X7Y9_E6BEG[5] ,
    \Tile_X7Y9_E6BEG[4] ,
    \Tile_X7Y9_E6BEG[3] ,
    \Tile_X7Y9_E6BEG[2] ,
    \Tile_X7Y9_E6BEG[1] ,
    \Tile_X7Y9_E6BEG[0] }),
    .Tile_X0Y0_E6END({\Tile_X6Y9_E6BEG[11] ,
    \Tile_X6Y9_E6BEG[10] ,
    \Tile_X6Y9_E6BEG[9] ,
    \Tile_X6Y9_E6BEG[8] ,
    \Tile_X6Y9_E6BEG[7] ,
    \Tile_X6Y9_E6BEG[6] ,
    \Tile_X6Y9_E6BEG[5] ,
    \Tile_X6Y9_E6BEG[4] ,
    \Tile_X6Y9_E6BEG[3] ,
    \Tile_X6Y9_E6BEG[2] ,
    \Tile_X6Y9_E6BEG[1] ,
    \Tile_X6Y9_E6BEG[0] }),
    .Tile_X0Y0_EE4BEG({\Tile_X7Y9_EE4BEG[15] ,
    \Tile_X7Y9_EE4BEG[14] ,
    \Tile_X7Y9_EE4BEG[13] ,
    \Tile_X7Y9_EE4BEG[12] ,
    \Tile_X7Y9_EE4BEG[11] ,
    \Tile_X7Y9_EE4BEG[10] ,
    \Tile_X7Y9_EE4BEG[9] ,
    \Tile_X7Y9_EE4BEG[8] ,
    \Tile_X7Y9_EE4BEG[7] ,
    \Tile_X7Y9_EE4BEG[6] ,
    \Tile_X7Y9_EE4BEG[5] ,
    \Tile_X7Y9_EE4BEG[4] ,
    \Tile_X7Y9_EE4BEG[3] ,
    \Tile_X7Y9_EE4BEG[2] ,
    \Tile_X7Y9_EE4BEG[1] ,
    \Tile_X7Y9_EE4BEG[0] }),
    .Tile_X0Y0_EE4END({\Tile_X6Y9_EE4BEG[15] ,
    \Tile_X6Y9_EE4BEG[14] ,
    \Tile_X6Y9_EE4BEG[13] ,
    \Tile_X6Y9_EE4BEG[12] ,
    \Tile_X6Y9_EE4BEG[11] ,
    \Tile_X6Y9_EE4BEG[10] ,
    \Tile_X6Y9_EE4BEG[9] ,
    \Tile_X6Y9_EE4BEG[8] ,
    \Tile_X6Y9_EE4BEG[7] ,
    \Tile_X6Y9_EE4BEG[6] ,
    \Tile_X6Y9_EE4BEG[5] ,
    \Tile_X6Y9_EE4BEG[4] ,
    \Tile_X6Y9_EE4BEG[3] ,
    \Tile_X6Y9_EE4BEG[2] ,
    \Tile_X6Y9_EE4BEG[1] ,
    \Tile_X6Y9_EE4BEG[0] }),
    .Tile_X0Y0_FrameData({\Tile_X6Y9_FrameData_O[31] ,
    \Tile_X6Y9_FrameData_O[30] ,
    \Tile_X6Y9_FrameData_O[29] ,
    \Tile_X6Y9_FrameData_O[28] ,
    \Tile_X6Y9_FrameData_O[27] ,
    \Tile_X6Y9_FrameData_O[26] ,
    \Tile_X6Y9_FrameData_O[25] ,
    \Tile_X6Y9_FrameData_O[24] ,
    \Tile_X6Y9_FrameData_O[23] ,
    \Tile_X6Y9_FrameData_O[22] ,
    \Tile_X6Y9_FrameData_O[21] ,
    \Tile_X6Y9_FrameData_O[20] ,
    \Tile_X6Y9_FrameData_O[19] ,
    \Tile_X6Y9_FrameData_O[18] ,
    \Tile_X6Y9_FrameData_O[17] ,
    \Tile_X6Y9_FrameData_O[16] ,
    \Tile_X6Y9_FrameData_O[15] ,
    \Tile_X6Y9_FrameData_O[14] ,
    \Tile_X6Y9_FrameData_O[13] ,
    \Tile_X6Y9_FrameData_O[12] ,
    \Tile_X6Y9_FrameData_O[11] ,
    \Tile_X6Y9_FrameData_O[10] ,
    \Tile_X6Y9_FrameData_O[9] ,
    \Tile_X6Y9_FrameData_O[8] ,
    \Tile_X6Y9_FrameData_O[7] ,
    \Tile_X6Y9_FrameData_O[6] ,
    \Tile_X6Y9_FrameData_O[5] ,
    \Tile_X6Y9_FrameData_O[4] ,
    \Tile_X6Y9_FrameData_O[3] ,
    \Tile_X6Y9_FrameData_O[2] ,
    \Tile_X6Y9_FrameData_O[1] ,
    \Tile_X6Y9_FrameData_O[0] }),
    .Tile_X0Y0_FrameData_O({\Tile_X7Y9_FrameData_O[31] ,
    \Tile_X7Y9_FrameData_O[30] ,
    \Tile_X7Y9_FrameData_O[29] ,
    \Tile_X7Y9_FrameData_O[28] ,
    \Tile_X7Y9_FrameData_O[27] ,
    \Tile_X7Y9_FrameData_O[26] ,
    \Tile_X7Y9_FrameData_O[25] ,
    \Tile_X7Y9_FrameData_O[24] ,
    \Tile_X7Y9_FrameData_O[23] ,
    \Tile_X7Y9_FrameData_O[22] ,
    \Tile_X7Y9_FrameData_O[21] ,
    \Tile_X7Y9_FrameData_O[20] ,
    \Tile_X7Y9_FrameData_O[19] ,
    \Tile_X7Y9_FrameData_O[18] ,
    \Tile_X7Y9_FrameData_O[17] ,
    \Tile_X7Y9_FrameData_O[16] ,
    \Tile_X7Y9_FrameData_O[15] ,
    \Tile_X7Y9_FrameData_O[14] ,
    \Tile_X7Y9_FrameData_O[13] ,
    \Tile_X7Y9_FrameData_O[12] ,
    \Tile_X7Y9_FrameData_O[11] ,
    \Tile_X7Y9_FrameData_O[10] ,
    \Tile_X7Y9_FrameData_O[9] ,
    \Tile_X7Y9_FrameData_O[8] ,
    \Tile_X7Y9_FrameData_O[7] ,
    \Tile_X7Y9_FrameData_O[6] ,
    \Tile_X7Y9_FrameData_O[5] ,
    \Tile_X7Y9_FrameData_O[4] ,
    \Tile_X7Y9_FrameData_O[3] ,
    \Tile_X7Y9_FrameData_O[2] ,
    \Tile_X7Y9_FrameData_O[1] ,
    \Tile_X7Y9_FrameData_O[0] }),
    .Tile_X0Y0_FrameStrobe_O({\Tile_X7Y9_FrameStrobe_O[19] ,
    \Tile_X7Y9_FrameStrobe_O[18] ,
    \Tile_X7Y9_FrameStrobe_O[17] ,
    \Tile_X7Y9_FrameStrobe_O[16] ,
    \Tile_X7Y9_FrameStrobe_O[15] ,
    \Tile_X7Y9_FrameStrobe_O[14] ,
    \Tile_X7Y9_FrameStrobe_O[13] ,
    \Tile_X7Y9_FrameStrobe_O[12] ,
    \Tile_X7Y9_FrameStrobe_O[11] ,
    \Tile_X7Y9_FrameStrobe_O[10] ,
    \Tile_X7Y9_FrameStrobe_O[9] ,
    \Tile_X7Y9_FrameStrobe_O[8] ,
    \Tile_X7Y9_FrameStrobe_O[7] ,
    \Tile_X7Y9_FrameStrobe_O[6] ,
    \Tile_X7Y9_FrameStrobe_O[5] ,
    \Tile_X7Y9_FrameStrobe_O[4] ,
    \Tile_X7Y9_FrameStrobe_O[3] ,
    \Tile_X7Y9_FrameStrobe_O[2] ,
    \Tile_X7Y9_FrameStrobe_O[1] ,
    \Tile_X7Y9_FrameStrobe_O[0] }),
    .Tile_X0Y0_N1BEG({\Tile_X7Y9_N1BEG[3] ,
    \Tile_X7Y9_N1BEG[2] ,
    \Tile_X7Y9_N1BEG[1] ,
    \Tile_X7Y9_N1BEG[0] }),
    .Tile_X0Y0_N2BEG({\Tile_X7Y9_N2BEG[7] ,
    \Tile_X7Y9_N2BEG[6] ,
    \Tile_X7Y9_N2BEG[5] ,
    \Tile_X7Y9_N2BEG[4] ,
    \Tile_X7Y9_N2BEG[3] ,
    \Tile_X7Y9_N2BEG[2] ,
    \Tile_X7Y9_N2BEG[1] ,
    \Tile_X7Y9_N2BEG[0] }),
    .Tile_X0Y0_N2BEGb({\Tile_X7Y9_N2BEGb[7] ,
    \Tile_X7Y9_N2BEGb[6] ,
    \Tile_X7Y9_N2BEGb[5] ,
    \Tile_X7Y9_N2BEGb[4] ,
    \Tile_X7Y9_N2BEGb[3] ,
    \Tile_X7Y9_N2BEGb[2] ,
    \Tile_X7Y9_N2BEGb[1] ,
    \Tile_X7Y9_N2BEGb[0] }),
    .Tile_X0Y0_N4BEG({\Tile_X7Y9_N4BEG[15] ,
    \Tile_X7Y9_N4BEG[14] ,
    \Tile_X7Y9_N4BEG[13] ,
    \Tile_X7Y9_N4BEG[12] ,
    \Tile_X7Y9_N4BEG[11] ,
    \Tile_X7Y9_N4BEG[10] ,
    \Tile_X7Y9_N4BEG[9] ,
    \Tile_X7Y9_N4BEG[8] ,
    \Tile_X7Y9_N4BEG[7] ,
    \Tile_X7Y9_N4BEG[6] ,
    \Tile_X7Y9_N4BEG[5] ,
    \Tile_X7Y9_N4BEG[4] ,
    \Tile_X7Y9_N4BEG[3] ,
    \Tile_X7Y9_N4BEG[2] ,
    \Tile_X7Y9_N4BEG[1] ,
    \Tile_X7Y9_N4BEG[0] }),
    .Tile_X0Y0_NN4BEG({\Tile_X7Y9_NN4BEG[15] ,
    \Tile_X7Y9_NN4BEG[14] ,
    \Tile_X7Y9_NN4BEG[13] ,
    \Tile_X7Y9_NN4BEG[12] ,
    \Tile_X7Y9_NN4BEG[11] ,
    \Tile_X7Y9_NN4BEG[10] ,
    \Tile_X7Y9_NN4BEG[9] ,
    \Tile_X7Y9_NN4BEG[8] ,
    \Tile_X7Y9_NN4BEG[7] ,
    \Tile_X7Y9_NN4BEG[6] ,
    \Tile_X7Y9_NN4BEG[5] ,
    \Tile_X7Y9_NN4BEG[4] ,
    \Tile_X7Y9_NN4BEG[3] ,
    \Tile_X7Y9_NN4BEG[2] ,
    \Tile_X7Y9_NN4BEG[1] ,
    \Tile_X7Y9_NN4BEG[0] }),
    .Tile_X0Y0_S1END({\Tile_X7Y8_S1BEG[3] ,
    \Tile_X7Y8_S1BEG[2] ,
    \Tile_X7Y8_S1BEG[1] ,
    \Tile_X7Y8_S1BEG[0] }),
    .Tile_X0Y0_S2END({\Tile_X7Y8_S2BEGb[7] ,
    \Tile_X7Y8_S2BEGb[6] ,
    \Tile_X7Y8_S2BEGb[5] ,
    \Tile_X7Y8_S2BEGb[4] ,
    \Tile_X7Y8_S2BEGb[3] ,
    \Tile_X7Y8_S2BEGb[2] ,
    \Tile_X7Y8_S2BEGb[1] ,
    \Tile_X7Y8_S2BEGb[0] }),
    .Tile_X0Y0_S2MID({\Tile_X7Y8_S2BEG[7] ,
    \Tile_X7Y8_S2BEG[6] ,
    \Tile_X7Y8_S2BEG[5] ,
    \Tile_X7Y8_S2BEG[4] ,
    \Tile_X7Y8_S2BEG[3] ,
    \Tile_X7Y8_S2BEG[2] ,
    \Tile_X7Y8_S2BEG[1] ,
    \Tile_X7Y8_S2BEG[0] }),
    .Tile_X0Y0_S4END({\Tile_X7Y8_S4BEG[15] ,
    \Tile_X7Y8_S4BEG[14] ,
    \Tile_X7Y8_S4BEG[13] ,
    \Tile_X7Y8_S4BEG[12] ,
    \Tile_X7Y8_S4BEG[11] ,
    \Tile_X7Y8_S4BEG[10] ,
    \Tile_X7Y8_S4BEG[9] ,
    \Tile_X7Y8_S4BEG[8] ,
    \Tile_X7Y8_S4BEG[7] ,
    \Tile_X7Y8_S4BEG[6] ,
    \Tile_X7Y8_S4BEG[5] ,
    \Tile_X7Y8_S4BEG[4] ,
    \Tile_X7Y8_S4BEG[3] ,
    \Tile_X7Y8_S4BEG[2] ,
    \Tile_X7Y8_S4BEG[1] ,
    \Tile_X7Y8_S4BEG[0] }),
    .Tile_X0Y0_SS4END({\Tile_X7Y8_SS4BEG[15] ,
    \Tile_X7Y8_SS4BEG[14] ,
    \Tile_X7Y8_SS4BEG[13] ,
    \Tile_X7Y8_SS4BEG[12] ,
    \Tile_X7Y8_SS4BEG[11] ,
    \Tile_X7Y8_SS4BEG[10] ,
    \Tile_X7Y8_SS4BEG[9] ,
    \Tile_X7Y8_SS4BEG[8] ,
    \Tile_X7Y8_SS4BEG[7] ,
    \Tile_X7Y8_SS4BEG[6] ,
    \Tile_X7Y8_SS4BEG[5] ,
    \Tile_X7Y8_SS4BEG[4] ,
    \Tile_X7Y8_SS4BEG[3] ,
    \Tile_X7Y8_SS4BEG[2] ,
    \Tile_X7Y8_SS4BEG[1] ,
    \Tile_X7Y8_SS4BEG[0] }),
    .Tile_X0Y0_W1BEG({\Tile_X7Y9_W1BEG[3] ,
    \Tile_X7Y9_W1BEG[2] ,
    \Tile_X7Y9_W1BEG[1] ,
    \Tile_X7Y9_W1BEG[0] }),
    .Tile_X0Y0_W1END({\Tile_X8Y9_W1BEG[3] ,
    \Tile_X8Y9_W1BEG[2] ,
    \Tile_X8Y9_W1BEG[1] ,
    \Tile_X8Y9_W1BEG[0] }),
    .Tile_X0Y0_W2BEG({\Tile_X7Y9_W2BEG[7] ,
    \Tile_X7Y9_W2BEG[6] ,
    \Tile_X7Y9_W2BEG[5] ,
    \Tile_X7Y9_W2BEG[4] ,
    \Tile_X7Y9_W2BEG[3] ,
    \Tile_X7Y9_W2BEG[2] ,
    \Tile_X7Y9_W2BEG[1] ,
    \Tile_X7Y9_W2BEG[0] }),
    .Tile_X0Y0_W2BEGb({\Tile_X7Y9_W2BEGb[7] ,
    \Tile_X7Y9_W2BEGb[6] ,
    \Tile_X7Y9_W2BEGb[5] ,
    \Tile_X7Y9_W2BEGb[4] ,
    \Tile_X7Y9_W2BEGb[3] ,
    \Tile_X7Y9_W2BEGb[2] ,
    \Tile_X7Y9_W2BEGb[1] ,
    \Tile_X7Y9_W2BEGb[0] }),
    .Tile_X0Y0_W2END({\Tile_X8Y9_W2BEGb[7] ,
    \Tile_X8Y9_W2BEGb[6] ,
    \Tile_X8Y9_W2BEGb[5] ,
    \Tile_X8Y9_W2BEGb[4] ,
    \Tile_X8Y9_W2BEGb[3] ,
    \Tile_X8Y9_W2BEGb[2] ,
    \Tile_X8Y9_W2BEGb[1] ,
    \Tile_X8Y9_W2BEGb[0] }),
    .Tile_X0Y0_W2MID({\Tile_X8Y9_W2BEG[7] ,
    \Tile_X8Y9_W2BEG[6] ,
    \Tile_X8Y9_W2BEG[5] ,
    \Tile_X8Y9_W2BEG[4] ,
    \Tile_X8Y9_W2BEG[3] ,
    \Tile_X8Y9_W2BEG[2] ,
    \Tile_X8Y9_W2BEG[1] ,
    \Tile_X8Y9_W2BEG[0] }),
    .Tile_X0Y0_W6BEG({\Tile_X7Y9_W6BEG[11] ,
    \Tile_X7Y9_W6BEG[10] ,
    \Tile_X7Y9_W6BEG[9] ,
    \Tile_X7Y9_W6BEG[8] ,
    \Tile_X7Y9_W6BEG[7] ,
    \Tile_X7Y9_W6BEG[6] ,
    \Tile_X7Y9_W6BEG[5] ,
    \Tile_X7Y9_W6BEG[4] ,
    \Tile_X7Y9_W6BEG[3] ,
    \Tile_X7Y9_W6BEG[2] ,
    \Tile_X7Y9_W6BEG[1] ,
    \Tile_X7Y9_W6BEG[0] }),
    .Tile_X0Y0_W6END({\Tile_X8Y9_W6BEG[11] ,
    \Tile_X8Y9_W6BEG[10] ,
    \Tile_X8Y9_W6BEG[9] ,
    \Tile_X8Y9_W6BEG[8] ,
    \Tile_X8Y9_W6BEG[7] ,
    \Tile_X8Y9_W6BEG[6] ,
    \Tile_X8Y9_W6BEG[5] ,
    \Tile_X8Y9_W6BEG[4] ,
    \Tile_X8Y9_W6BEG[3] ,
    \Tile_X8Y9_W6BEG[2] ,
    \Tile_X8Y9_W6BEG[1] ,
    \Tile_X8Y9_W6BEG[0] }),
    .Tile_X0Y0_WW4BEG({\Tile_X7Y9_WW4BEG[15] ,
    \Tile_X7Y9_WW4BEG[14] ,
    \Tile_X7Y9_WW4BEG[13] ,
    \Tile_X7Y9_WW4BEG[12] ,
    \Tile_X7Y9_WW4BEG[11] ,
    \Tile_X7Y9_WW4BEG[10] ,
    \Tile_X7Y9_WW4BEG[9] ,
    \Tile_X7Y9_WW4BEG[8] ,
    \Tile_X7Y9_WW4BEG[7] ,
    \Tile_X7Y9_WW4BEG[6] ,
    \Tile_X7Y9_WW4BEG[5] ,
    \Tile_X7Y9_WW4BEG[4] ,
    \Tile_X7Y9_WW4BEG[3] ,
    \Tile_X7Y9_WW4BEG[2] ,
    \Tile_X7Y9_WW4BEG[1] ,
    \Tile_X7Y9_WW4BEG[0] }),
    .Tile_X0Y0_WW4END({\Tile_X8Y9_WW4BEG[15] ,
    \Tile_X8Y9_WW4BEG[14] ,
    \Tile_X8Y9_WW4BEG[13] ,
    \Tile_X8Y9_WW4BEG[12] ,
    \Tile_X8Y9_WW4BEG[11] ,
    \Tile_X8Y9_WW4BEG[10] ,
    \Tile_X8Y9_WW4BEG[9] ,
    \Tile_X8Y9_WW4BEG[8] ,
    \Tile_X8Y9_WW4BEG[7] ,
    \Tile_X8Y9_WW4BEG[6] ,
    \Tile_X8Y9_WW4BEG[5] ,
    \Tile_X8Y9_WW4BEG[4] ,
    \Tile_X8Y9_WW4BEG[3] ,
    \Tile_X8Y9_WW4BEG[2] ,
    \Tile_X8Y9_WW4BEG[1] ,
    \Tile_X8Y9_WW4BEG[0] }),
    .Tile_X0Y1_E1BEG({\Tile_X7Y10_E1BEG[3] ,
    \Tile_X7Y10_E1BEG[2] ,
    \Tile_X7Y10_E1BEG[1] ,
    \Tile_X7Y10_E1BEG[0] }),
    .Tile_X0Y1_E1END({\Tile_X6Y10_E1BEG[3] ,
    \Tile_X6Y10_E1BEG[2] ,
    \Tile_X6Y10_E1BEG[1] ,
    \Tile_X6Y10_E1BEG[0] }),
    .Tile_X0Y1_E2BEG({\Tile_X7Y10_E2BEG[7] ,
    \Tile_X7Y10_E2BEG[6] ,
    \Tile_X7Y10_E2BEG[5] ,
    \Tile_X7Y10_E2BEG[4] ,
    \Tile_X7Y10_E2BEG[3] ,
    \Tile_X7Y10_E2BEG[2] ,
    \Tile_X7Y10_E2BEG[1] ,
    \Tile_X7Y10_E2BEG[0] }),
    .Tile_X0Y1_E2BEGb({\Tile_X7Y10_E2BEGb[7] ,
    \Tile_X7Y10_E2BEGb[6] ,
    \Tile_X7Y10_E2BEGb[5] ,
    \Tile_X7Y10_E2BEGb[4] ,
    \Tile_X7Y10_E2BEGb[3] ,
    \Tile_X7Y10_E2BEGb[2] ,
    \Tile_X7Y10_E2BEGb[1] ,
    \Tile_X7Y10_E2BEGb[0] }),
    .Tile_X0Y1_E2END({\Tile_X6Y10_E2BEGb[7] ,
    \Tile_X6Y10_E2BEGb[6] ,
    \Tile_X6Y10_E2BEGb[5] ,
    \Tile_X6Y10_E2BEGb[4] ,
    \Tile_X6Y10_E2BEGb[3] ,
    \Tile_X6Y10_E2BEGb[2] ,
    \Tile_X6Y10_E2BEGb[1] ,
    \Tile_X6Y10_E2BEGb[0] }),
    .Tile_X0Y1_E2MID({\Tile_X6Y10_E2BEG[7] ,
    \Tile_X6Y10_E2BEG[6] ,
    \Tile_X6Y10_E2BEG[5] ,
    \Tile_X6Y10_E2BEG[4] ,
    \Tile_X6Y10_E2BEG[3] ,
    \Tile_X6Y10_E2BEG[2] ,
    \Tile_X6Y10_E2BEG[1] ,
    \Tile_X6Y10_E2BEG[0] }),
    .Tile_X0Y1_E6BEG({\Tile_X7Y10_E6BEG[11] ,
    \Tile_X7Y10_E6BEG[10] ,
    \Tile_X7Y10_E6BEG[9] ,
    \Tile_X7Y10_E6BEG[8] ,
    \Tile_X7Y10_E6BEG[7] ,
    \Tile_X7Y10_E6BEG[6] ,
    \Tile_X7Y10_E6BEG[5] ,
    \Tile_X7Y10_E6BEG[4] ,
    \Tile_X7Y10_E6BEG[3] ,
    \Tile_X7Y10_E6BEG[2] ,
    \Tile_X7Y10_E6BEG[1] ,
    \Tile_X7Y10_E6BEG[0] }),
    .Tile_X0Y1_E6END({\Tile_X6Y10_E6BEG[11] ,
    \Tile_X6Y10_E6BEG[10] ,
    \Tile_X6Y10_E6BEG[9] ,
    \Tile_X6Y10_E6BEG[8] ,
    \Tile_X6Y10_E6BEG[7] ,
    \Tile_X6Y10_E6BEG[6] ,
    \Tile_X6Y10_E6BEG[5] ,
    \Tile_X6Y10_E6BEG[4] ,
    \Tile_X6Y10_E6BEG[3] ,
    \Tile_X6Y10_E6BEG[2] ,
    \Tile_X6Y10_E6BEG[1] ,
    \Tile_X6Y10_E6BEG[0] }),
    .Tile_X0Y1_EE4BEG({\Tile_X7Y10_EE4BEG[15] ,
    \Tile_X7Y10_EE4BEG[14] ,
    \Tile_X7Y10_EE4BEG[13] ,
    \Tile_X7Y10_EE4BEG[12] ,
    \Tile_X7Y10_EE4BEG[11] ,
    \Tile_X7Y10_EE4BEG[10] ,
    \Tile_X7Y10_EE4BEG[9] ,
    \Tile_X7Y10_EE4BEG[8] ,
    \Tile_X7Y10_EE4BEG[7] ,
    \Tile_X7Y10_EE4BEG[6] ,
    \Tile_X7Y10_EE4BEG[5] ,
    \Tile_X7Y10_EE4BEG[4] ,
    \Tile_X7Y10_EE4BEG[3] ,
    \Tile_X7Y10_EE4BEG[2] ,
    \Tile_X7Y10_EE4BEG[1] ,
    \Tile_X7Y10_EE4BEG[0] }),
    .Tile_X0Y1_EE4END({\Tile_X6Y10_EE4BEG[15] ,
    \Tile_X6Y10_EE4BEG[14] ,
    \Tile_X6Y10_EE4BEG[13] ,
    \Tile_X6Y10_EE4BEG[12] ,
    \Tile_X6Y10_EE4BEG[11] ,
    \Tile_X6Y10_EE4BEG[10] ,
    \Tile_X6Y10_EE4BEG[9] ,
    \Tile_X6Y10_EE4BEG[8] ,
    \Tile_X6Y10_EE4BEG[7] ,
    \Tile_X6Y10_EE4BEG[6] ,
    \Tile_X6Y10_EE4BEG[5] ,
    \Tile_X6Y10_EE4BEG[4] ,
    \Tile_X6Y10_EE4BEG[3] ,
    \Tile_X6Y10_EE4BEG[2] ,
    \Tile_X6Y10_EE4BEG[1] ,
    \Tile_X6Y10_EE4BEG[0] }),
    .Tile_X0Y1_FrameData({\Tile_X6Y10_FrameData_O[31] ,
    \Tile_X6Y10_FrameData_O[30] ,
    \Tile_X6Y10_FrameData_O[29] ,
    \Tile_X6Y10_FrameData_O[28] ,
    \Tile_X6Y10_FrameData_O[27] ,
    \Tile_X6Y10_FrameData_O[26] ,
    \Tile_X6Y10_FrameData_O[25] ,
    \Tile_X6Y10_FrameData_O[24] ,
    \Tile_X6Y10_FrameData_O[23] ,
    \Tile_X6Y10_FrameData_O[22] ,
    \Tile_X6Y10_FrameData_O[21] ,
    \Tile_X6Y10_FrameData_O[20] ,
    \Tile_X6Y10_FrameData_O[19] ,
    \Tile_X6Y10_FrameData_O[18] ,
    \Tile_X6Y10_FrameData_O[17] ,
    \Tile_X6Y10_FrameData_O[16] ,
    \Tile_X6Y10_FrameData_O[15] ,
    \Tile_X6Y10_FrameData_O[14] ,
    \Tile_X6Y10_FrameData_O[13] ,
    \Tile_X6Y10_FrameData_O[12] ,
    \Tile_X6Y10_FrameData_O[11] ,
    \Tile_X6Y10_FrameData_O[10] ,
    \Tile_X6Y10_FrameData_O[9] ,
    \Tile_X6Y10_FrameData_O[8] ,
    \Tile_X6Y10_FrameData_O[7] ,
    \Tile_X6Y10_FrameData_O[6] ,
    \Tile_X6Y10_FrameData_O[5] ,
    \Tile_X6Y10_FrameData_O[4] ,
    \Tile_X6Y10_FrameData_O[3] ,
    \Tile_X6Y10_FrameData_O[2] ,
    \Tile_X6Y10_FrameData_O[1] ,
    \Tile_X6Y10_FrameData_O[0] }),
    .Tile_X0Y1_FrameData_O({\Tile_X7Y10_FrameData_O[31] ,
    \Tile_X7Y10_FrameData_O[30] ,
    \Tile_X7Y10_FrameData_O[29] ,
    \Tile_X7Y10_FrameData_O[28] ,
    \Tile_X7Y10_FrameData_O[27] ,
    \Tile_X7Y10_FrameData_O[26] ,
    \Tile_X7Y10_FrameData_O[25] ,
    \Tile_X7Y10_FrameData_O[24] ,
    \Tile_X7Y10_FrameData_O[23] ,
    \Tile_X7Y10_FrameData_O[22] ,
    \Tile_X7Y10_FrameData_O[21] ,
    \Tile_X7Y10_FrameData_O[20] ,
    \Tile_X7Y10_FrameData_O[19] ,
    \Tile_X7Y10_FrameData_O[18] ,
    \Tile_X7Y10_FrameData_O[17] ,
    \Tile_X7Y10_FrameData_O[16] ,
    \Tile_X7Y10_FrameData_O[15] ,
    \Tile_X7Y10_FrameData_O[14] ,
    \Tile_X7Y10_FrameData_O[13] ,
    \Tile_X7Y10_FrameData_O[12] ,
    \Tile_X7Y10_FrameData_O[11] ,
    \Tile_X7Y10_FrameData_O[10] ,
    \Tile_X7Y10_FrameData_O[9] ,
    \Tile_X7Y10_FrameData_O[8] ,
    \Tile_X7Y10_FrameData_O[7] ,
    \Tile_X7Y10_FrameData_O[6] ,
    \Tile_X7Y10_FrameData_O[5] ,
    \Tile_X7Y10_FrameData_O[4] ,
    \Tile_X7Y10_FrameData_O[3] ,
    \Tile_X7Y10_FrameData_O[2] ,
    \Tile_X7Y10_FrameData_O[1] ,
    \Tile_X7Y10_FrameData_O[0] }),
    .Tile_X0Y1_FrameStrobe({\Tile_X7Y11_FrameStrobe_O[19] ,
    \Tile_X7Y11_FrameStrobe_O[18] ,
    \Tile_X7Y11_FrameStrobe_O[17] ,
    \Tile_X7Y11_FrameStrobe_O[16] ,
    \Tile_X7Y11_FrameStrobe_O[15] ,
    \Tile_X7Y11_FrameStrobe_O[14] ,
    \Tile_X7Y11_FrameStrobe_O[13] ,
    \Tile_X7Y11_FrameStrobe_O[12] ,
    \Tile_X7Y11_FrameStrobe_O[11] ,
    \Tile_X7Y11_FrameStrobe_O[10] ,
    \Tile_X7Y11_FrameStrobe_O[9] ,
    \Tile_X7Y11_FrameStrobe_O[8] ,
    \Tile_X7Y11_FrameStrobe_O[7] ,
    \Tile_X7Y11_FrameStrobe_O[6] ,
    \Tile_X7Y11_FrameStrobe_O[5] ,
    \Tile_X7Y11_FrameStrobe_O[4] ,
    \Tile_X7Y11_FrameStrobe_O[3] ,
    \Tile_X7Y11_FrameStrobe_O[2] ,
    \Tile_X7Y11_FrameStrobe_O[1] ,
    \Tile_X7Y11_FrameStrobe_O[0] }),
    .Tile_X0Y1_N1END({\Tile_X7Y11_N1BEG[3] ,
    \Tile_X7Y11_N1BEG[2] ,
    \Tile_X7Y11_N1BEG[1] ,
    \Tile_X7Y11_N1BEG[0] }),
    .Tile_X0Y1_N2END({\Tile_X7Y11_N2BEGb[7] ,
    \Tile_X7Y11_N2BEGb[6] ,
    \Tile_X7Y11_N2BEGb[5] ,
    \Tile_X7Y11_N2BEGb[4] ,
    \Tile_X7Y11_N2BEGb[3] ,
    \Tile_X7Y11_N2BEGb[2] ,
    \Tile_X7Y11_N2BEGb[1] ,
    \Tile_X7Y11_N2BEGb[0] }),
    .Tile_X0Y1_N2MID({\Tile_X7Y11_N2BEG[7] ,
    \Tile_X7Y11_N2BEG[6] ,
    \Tile_X7Y11_N2BEG[5] ,
    \Tile_X7Y11_N2BEG[4] ,
    \Tile_X7Y11_N2BEG[3] ,
    \Tile_X7Y11_N2BEG[2] ,
    \Tile_X7Y11_N2BEG[1] ,
    \Tile_X7Y11_N2BEG[0] }),
    .Tile_X0Y1_N4END({\Tile_X7Y11_N4BEG[15] ,
    \Tile_X7Y11_N4BEG[14] ,
    \Tile_X7Y11_N4BEG[13] ,
    \Tile_X7Y11_N4BEG[12] ,
    \Tile_X7Y11_N4BEG[11] ,
    \Tile_X7Y11_N4BEG[10] ,
    \Tile_X7Y11_N4BEG[9] ,
    \Tile_X7Y11_N4BEG[8] ,
    \Tile_X7Y11_N4BEG[7] ,
    \Tile_X7Y11_N4BEG[6] ,
    \Tile_X7Y11_N4BEG[5] ,
    \Tile_X7Y11_N4BEG[4] ,
    \Tile_X7Y11_N4BEG[3] ,
    \Tile_X7Y11_N4BEG[2] ,
    \Tile_X7Y11_N4BEG[1] ,
    \Tile_X7Y11_N4BEG[0] }),
    .Tile_X0Y1_NN4END({\Tile_X7Y11_NN4BEG[15] ,
    \Tile_X7Y11_NN4BEG[14] ,
    \Tile_X7Y11_NN4BEG[13] ,
    \Tile_X7Y11_NN4BEG[12] ,
    \Tile_X7Y11_NN4BEG[11] ,
    \Tile_X7Y11_NN4BEG[10] ,
    \Tile_X7Y11_NN4BEG[9] ,
    \Tile_X7Y11_NN4BEG[8] ,
    \Tile_X7Y11_NN4BEG[7] ,
    \Tile_X7Y11_NN4BEG[6] ,
    \Tile_X7Y11_NN4BEG[5] ,
    \Tile_X7Y11_NN4BEG[4] ,
    \Tile_X7Y11_NN4BEG[3] ,
    \Tile_X7Y11_NN4BEG[2] ,
    \Tile_X7Y11_NN4BEG[1] ,
    \Tile_X7Y11_NN4BEG[0] }),
    .Tile_X0Y1_S1BEG({\Tile_X7Y10_S1BEG[3] ,
    \Tile_X7Y10_S1BEG[2] ,
    \Tile_X7Y10_S1BEG[1] ,
    \Tile_X7Y10_S1BEG[0] }),
    .Tile_X0Y1_S2BEG({\Tile_X7Y10_S2BEG[7] ,
    \Tile_X7Y10_S2BEG[6] ,
    \Tile_X7Y10_S2BEG[5] ,
    \Tile_X7Y10_S2BEG[4] ,
    \Tile_X7Y10_S2BEG[3] ,
    \Tile_X7Y10_S2BEG[2] ,
    \Tile_X7Y10_S2BEG[1] ,
    \Tile_X7Y10_S2BEG[0] }),
    .Tile_X0Y1_S2BEGb({\Tile_X7Y10_S2BEGb[7] ,
    \Tile_X7Y10_S2BEGb[6] ,
    \Tile_X7Y10_S2BEGb[5] ,
    \Tile_X7Y10_S2BEGb[4] ,
    \Tile_X7Y10_S2BEGb[3] ,
    \Tile_X7Y10_S2BEGb[2] ,
    \Tile_X7Y10_S2BEGb[1] ,
    \Tile_X7Y10_S2BEGb[0] }),
    .Tile_X0Y1_S4BEG({\Tile_X7Y10_S4BEG[15] ,
    \Tile_X7Y10_S4BEG[14] ,
    \Tile_X7Y10_S4BEG[13] ,
    \Tile_X7Y10_S4BEG[12] ,
    \Tile_X7Y10_S4BEG[11] ,
    \Tile_X7Y10_S4BEG[10] ,
    \Tile_X7Y10_S4BEG[9] ,
    \Tile_X7Y10_S4BEG[8] ,
    \Tile_X7Y10_S4BEG[7] ,
    \Tile_X7Y10_S4BEG[6] ,
    \Tile_X7Y10_S4BEG[5] ,
    \Tile_X7Y10_S4BEG[4] ,
    \Tile_X7Y10_S4BEG[3] ,
    \Tile_X7Y10_S4BEG[2] ,
    \Tile_X7Y10_S4BEG[1] ,
    \Tile_X7Y10_S4BEG[0] }),
    .Tile_X0Y1_SS4BEG({\Tile_X7Y10_SS4BEG[15] ,
    \Tile_X7Y10_SS4BEG[14] ,
    \Tile_X7Y10_SS4BEG[13] ,
    \Tile_X7Y10_SS4BEG[12] ,
    \Tile_X7Y10_SS4BEG[11] ,
    \Tile_X7Y10_SS4BEG[10] ,
    \Tile_X7Y10_SS4BEG[9] ,
    \Tile_X7Y10_SS4BEG[8] ,
    \Tile_X7Y10_SS4BEG[7] ,
    \Tile_X7Y10_SS4BEG[6] ,
    \Tile_X7Y10_SS4BEG[5] ,
    \Tile_X7Y10_SS4BEG[4] ,
    \Tile_X7Y10_SS4BEG[3] ,
    \Tile_X7Y10_SS4BEG[2] ,
    \Tile_X7Y10_SS4BEG[1] ,
    \Tile_X7Y10_SS4BEG[0] }),
    .Tile_X0Y1_W1BEG({\Tile_X7Y10_W1BEG[3] ,
    \Tile_X7Y10_W1BEG[2] ,
    \Tile_X7Y10_W1BEG[1] ,
    \Tile_X7Y10_W1BEG[0] }),
    .Tile_X0Y1_W1END({\Tile_X8Y10_W1BEG[3] ,
    \Tile_X8Y10_W1BEG[2] ,
    \Tile_X8Y10_W1BEG[1] ,
    \Tile_X8Y10_W1BEG[0] }),
    .Tile_X0Y1_W2BEG({\Tile_X7Y10_W2BEG[7] ,
    \Tile_X7Y10_W2BEG[6] ,
    \Tile_X7Y10_W2BEG[5] ,
    \Tile_X7Y10_W2BEG[4] ,
    \Tile_X7Y10_W2BEG[3] ,
    \Tile_X7Y10_W2BEG[2] ,
    \Tile_X7Y10_W2BEG[1] ,
    \Tile_X7Y10_W2BEG[0] }),
    .Tile_X0Y1_W2BEGb({\Tile_X7Y10_W2BEGb[7] ,
    \Tile_X7Y10_W2BEGb[6] ,
    \Tile_X7Y10_W2BEGb[5] ,
    \Tile_X7Y10_W2BEGb[4] ,
    \Tile_X7Y10_W2BEGb[3] ,
    \Tile_X7Y10_W2BEGb[2] ,
    \Tile_X7Y10_W2BEGb[1] ,
    \Tile_X7Y10_W2BEGb[0] }),
    .Tile_X0Y1_W2END({\Tile_X8Y10_W2BEGb[7] ,
    \Tile_X8Y10_W2BEGb[6] ,
    \Tile_X8Y10_W2BEGb[5] ,
    \Tile_X8Y10_W2BEGb[4] ,
    \Tile_X8Y10_W2BEGb[3] ,
    \Tile_X8Y10_W2BEGb[2] ,
    \Tile_X8Y10_W2BEGb[1] ,
    \Tile_X8Y10_W2BEGb[0] }),
    .Tile_X0Y1_W2MID({\Tile_X8Y10_W2BEG[7] ,
    \Tile_X8Y10_W2BEG[6] ,
    \Tile_X8Y10_W2BEG[5] ,
    \Tile_X8Y10_W2BEG[4] ,
    \Tile_X8Y10_W2BEG[3] ,
    \Tile_X8Y10_W2BEG[2] ,
    \Tile_X8Y10_W2BEG[1] ,
    \Tile_X8Y10_W2BEG[0] }),
    .Tile_X0Y1_W6BEG({\Tile_X7Y10_W6BEG[11] ,
    \Tile_X7Y10_W6BEG[10] ,
    \Tile_X7Y10_W6BEG[9] ,
    \Tile_X7Y10_W6BEG[8] ,
    \Tile_X7Y10_W6BEG[7] ,
    \Tile_X7Y10_W6BEG[6] ,
    \Tile_X7Y10_W6BEG[5] ,
    \Tile_X7Y10_W6BEG[4] ,
    \Tile_X7Y10_W6BEG[3] ,
    \Tile_X7Y10_W6BEG[2] ,
    \Tile_X7Y10_W6BEG[1] ,
    \Tile_X7Y10_W6BEG[0] }),
    .Tile_X0Y1_W6END({\Tile_X8Y10_W6BEG[11] ,
    \Tile_X8Y10_W6BEG[10] ,
    \Tile_X8Y10_W6BEG[9] ,
    \Tile_X8Y10_W6BEG[8] ,
    \Tile_X8Y10_W6BEG[7] ,
    \Tile_X8Y10_W6BEG[6] ,
    \Tile_X8Y10_W6BEG[5] ,
    \Tile_X8Y10_W6BEG[4] ,
    \Tile_X8Y10_W6BEG[3] ,
    \Tile_X8Y10_W6BEG[2] ,
    \Tile_X8Y10_W6BEG[1] ,
    \Tile_X8Y10_W6BEG[0] }),
    .Tile_X0Y1_WW4BEG({\Tile_X7Y10_WW4BEG[15] ,
    \Tile_X7Y10_WW4BEG[14] ,
    \Tile_X7Y10_WW4BEG[13] ,
    \Tile_X7Y10_WW4BEG[12] ,
    \Tile_X7Y10_WW4BEG[11] ,
    \Tile_X7Y10_WW4BEG[10] ,
    \Tile_X7Y10_WW4BEG[9] ,
    \Tile_X7Y10_WW4BEG[8] ,
    \Tile_X7Y10_WW4BEG[7] ,
    \Tile_X7Y10_WW4BEG[6] ,
    \Tile_X7Y10_WW4BEG[5] ,
    \Tile_X7Y10_WW4BEG[4] ,
    \Tile_X7Y10_WW4BEG[3] ,
    \Tile_X7Y10_WW4BEG[2] ,
    \Tile_X7Y10_WW4BEG[1] ,
    \Tile_X7Y10_WW4BEG[0] }),
    .Tile_X0Y1_WW4END({\Tile_X8Y10_WW4BEG[15] ,
    \Tile_X8Y10_WW4BEG[14] ,
    \Tile_X8Y10_WW4BEG[13] ,
    \Tile_X8Y10_WW4BEG[12] ,
    \Tile_X8Y10_WW4BEG[11] ,
    \Tile_X8Y10_WW4BEG[10] ,
    \Tile_X8Y10_WW4BEG[9] ,
    \Tile_X8Y10_WW4BEG[8] ,
    \Tile_X8Y10_WW4BEG[7] ,
    \Tile_X8Y10_WW4BEG[6] ,
    \Tile_X8Y10_WW4BEG[5] ,
    \Tile_X8Y10_WW4BEG[4] ,
    \Tile_X8Y10_WW4BEG[3] ,
    \Tile_X8Y10_WW4BEG[2] ,
    \Tile_X8Y10_WW4BEG[1] ,
    \Tile_X8Y10_WW4BEG[0] }));
 N_term_single Tile_X8Y0_N_term_single (.Ci(Tile_X8Y1_Co),
    .UserCLK(Tile_X8Y1_UserCLKo),
    .UserCLKo(Tile_X8Y0_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .FrameData({\Tile_X7Y0_FrameData_O[31] ,
    \Tile_X7Y0_FrameData_O[30] ,
    \Tile_X7Y0_FrameData_O[29] ,
    \Tile_X7Y0_FrameData_O[28] ,
    \Tile_X7Y0_FrameData_O[27] ,
    \Tile_X7Y0_FrameData_O[26] ,
    \Tile_X7Y0_FrameData_O[25] ,
    \Tile_X7Y0_FrameData_O[24] ,
    \Tile_X7Y0_FrameData_O[23] ,
    \Tile_X7Y0_FrameData_O[22] ,
    \Tile_X7Y0_FrameData_O[21] ,
    \Tile_X7Y0_FrameData_O[20] ,
    \Tile_X7Y0_FrameData_O[19] ,
    \Tile_X7Y0_FrameData_O[18] ,
    \Tile_X7Y0_FrameData_O[17] ,
    \Tile_X7Y0_FrameData_O[16] ,
    \Tile_X7Y0_FrameData_O[15] ,
    \Tile_X7Y0_FrameData_O[14] ,
    \Tile_X7Y0_FrameData_O[13] ,
    \Tile_X7Y0_FrameData_O[12] ,
    \Tile_X7Y0_FrameData_O[11] ,
    \Tile_X7Y0_FrameData_O[10] ,
    \Tile_X7Y0_FrameData_O[9] ,
    \Tile_X7Y0_FrameData_O[8] ,
    \Tile_X7Y0_FrameData_O[7] ,
    \Tile_X7Y0_FrameData_O[6] ,
    \Tile_X7Y0_FrameData_O[5] ,
    \Tile_X7Y0_FrameData_O[4] ,
    \Tile_X7Y0_FrameData_O[3] ,
    \Tile_X7Y0_FrameData_O[2] ,
    \Tile_X7Y0_FrameData_O[1] ,
    \Tile_X7Y0_FrameData_O[0] }),
    .FrameData_O({\Tile_X8Y0_FrameData_O[31] ,
    \Tile_X8Y0_FrameData_O[30] ,
    \Tile_X8Y0_FrameData_O[29] ,
    \Tile_X8Y0_FrameData_O[28] ,
    \Tile_X8Y0_FrameData_O[27] ,
    \Tile_X8Y0_FrameData_O[26] ,
    \Tile_X8Y0_FrameData_O[25] ,
    \Tile_X8Y0_FrameData_O[24] ,
    \Tile_X8Y0_FrameData_O[23] ,
    \Tile_X8Y0_FrameData_O[22] ,
    \Tile_X8Y0_FrameData_O[21] ,
    \Tile_X8Y0_FrameData_O[20] ,
    \Tile_X8Y0_FrameData_O[19] ,
    \Tile_X8Y0_FrameData_O[18] ,
    \Tile_X8Y0_FrameData_O[17] ,
    \Tile_X8Y0_FrameData_O[16] ,
    \Tile_X8Y0_FrameData_O[15] ,
    \Tile_X8Y0_FrameData_O[14] ,
    \Tile_X8Y0_FrameData_O[13] ,
    \Tile_X8Y0_FrameData_O[12] ,
    \Tile_X8Y0_FrameData_O[11] ,
    \Tile_X8Y0_FrameData_O[10] ,
    \Tile_X8Y0_FrameData_O[9] ,
    \Tile_X8Y0_FrameData_O[8] ,
    \Tile_X8Y0_FrameData_O[7] ,
    \Tile_X8Y0_FrameData_O[6] ,
    \Tile_X8Y0_FrameData_O[5] ,
    \Tile_X8Y0_FrameData_O[4] ,
    \Tile_X8Y0_FrameData_O[3] ,
    \Tile_X8Y0_FrameData_O[2] ,
    \Tile_X8Y0_FrameData_O[1] ,
    \Tile_X8Y0_FrameData_O[0] }),
    .FrameStrobe({\Tile_X8Y1_FrameStrobe_O[19] ,
    \Tile_X8Y1_FrameStrobe_O[18] ,
    \Tile_X8Y1_FrameStrobe_O[17] ,
    \Tile_X8Y1_FrameStrobe_O[16] ,
    \Tile_X8Y1_FrameStrobe_O[15] ,
    \Tile_X8Y1_FrameStrobe_O[14] ,
    \Tile_X8Y1_FrameStrobe_O[13] ,
    \Tile_X8Y1_FrameStrobe_O[12] ,
    \Tile_X8Y1_FrameStrobe_O[11] ,
    \Tile_X8Y1_FrameStrobe_O[10] ,
    \Tile_X8Y1_FrameStrobe_O[9] ,
    \Tile_X8Y1_FrameStrobe_O[8] ,
    \Tile_X8Y1_FrameStrobe_O[7] ,
    \Tile_X8Y1_FrameStrobe_O[6] ,
    \Tile_X8Y1_FrameStrobe_O[5] ,
    \Tile_X8Y1_FrameStrobe_O[4] ,
    \Tile_X8Y1_FrameStrobe_O[3] ,
    \Tile_X8Y1_FrameStrobe_O[2] ,
    \Tile_X8Y1_FrameStrobe_O[1] ,
    \Tile_X8Y1_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X8Y0_FrameStrobe_O[19] ,
    \Tile_X8Y0_FrameStrobe_O[18] ,
    \Tile_X8Y0_FrameStrobe_O[17] ,
    \Tile_X8Y0_FrameStrobe_O[16] ,
    \Tile_X8Y0_FrameStrobe_O[15] ,
    \Tile_X8Y0_FrameStrobe_O[14] ,
    \Tile_X8Y0_FrameStrobe_O[13] ,
    \Tile_X8Y0_FrameStrobe_O[12] ,
    \Tile_X8Y0_FrameStrobe_O[11] ,
    \Tile_X8Y0_FrameStrobe_O[10] ,
    \Tile_X8Y0_FrameStrobe_O[9] ,
    \Tile_X8Y0_FrameStrobe_O[8] ,
    \Tile_X8Y0_FrameStrobe_O[7] ,
    \Tile_X8Y0_FrameStrobe_O[6] ,
    \Tile_X8Y0_FrameStrobe_O[5] ,
    \Tile_X8Y0_FrameStrobe_O[4] ,
    \Tile_X8Y0_FrameStrobe_O[3] ,
    \Tile_X8Y0_FrameStrobe_O[2] ,
    \Tile_X8Y0_FrameStrobe_O[1] ,
    \Tile_X8Y0_FrameStrobe_O[0] }),
    .N1END({\Tile_X8Y1_N1BEG[3] ,
    \Tile_X8Y1_N1BEG[2] ,
    \Tile_X8Y1_N1BEG[1] ,
    \Tile_X8Y1_N1BEG[0] }),
    .N2END({\Tile_X8Y1_N2BEGb[7] ,
    \Tile_X8Y1_N2BEGb[6] ,
    \Tile_X8Y1_N2BEGb[5] ,
    \Tile_X8Y1_N2BEGb[4] ,
    \Tile_X8Y1_N2BEGb[3] ,
    \Tile_X8Y1_N2BEGb[2] ,
    \Tile_X8Y1_N2BEGb[1] ,
    \Tile_X8Y1_N2BEGb[0] }),
    .N2MID({\Tile_X8Y1_N2BEG[7] ,
    \Tile_X8Y1_N2BEG[6] ,
    \Tile_X8Y1_N2BEG[5] ,
    \Tile_X8Y1_N2BEG[4] ,
    \Tile_X8Y1_N2BEG[3] ,
    \Tile_X8Y1_N2BEG[2] ,
    \Tile_X8Y1_N2BEG[1] ,
    \Tile_X8Y1_N2BEG[0] }),
    .N4END({\Tile_X8Y1_N4BEG[15] ,
    \Tile_X8Y1_N4BEG[14] ,
    \Tile_X8Y1_N4BEG[13] ,
    \Tile_X8Y1_N4BEG[12] ,
    \Tile_X8Y1_N4BEG[11] ,
    \Tile_X8Y1_N4BEG[10] ,
    \Tile_X8Y1_N4BEG[9] ,
    \Tile_X8Y1_N4BEG[8] ,
    \Tile_X8Y1_N4BEG[7] ,
    \Tile_X8Y1_N4BEG[6] ,
    \Tile_X8Y1_N4BEG[5] ,
    \Tile_X8Y1_N4BEG[4] ,
    \Tile_X8Y1_N4BEG[3] ,
    \Tile_X8Y1_N4BEG[2] ,
    \Tile_X8Y1_N4BEG[1] ,
    \Tile_X8Y1_N4BEG[0] }),
    .NN4END({\Tile_X8Y1_NN4BEG[15] ,
    \Tile_X8Y1_NN4BEG[14] ,
    \Tile_X8Y1_NN4BEG[13] ,
    \Tile_X8Y1_NN4BEG[12] ,
    \Tile_X8Y1_NN4BEG[11] ,
    \Tile_X8Y1_NN4BEG[10] ,
    \Tile_X8Y1_NN4BEG[9] ,
    \Tile_X8Y1_NN4BEG[8] ,
    \Tile_X8Y1_NN4BEG[7] ,
    \Tile_X8Y1_NN4BEG[6] ,
    \Tile_X8Y1_NN4BEG[5] ,
    \Tile_X8Y1_NN4BEG[4] ,
    \Tile_X8Y1_NN4BEG[3] ,
    \Tile_X8Y1_NN4BEG[2] ,
    \Tile_X8Y1_NN4BEG[1] ,
    \Tile_X8Y1_NN4BEG[0] }),
    .S1BEG({\Tile_X8Y0_S1BEG[3] ,
    \Tile_X8Y0_S1BEG[2] ,
    \Tile_X8Y0_S1BEG[1] ,
    \Tile_X8Y0_S1BEG[0] }),
    .S2BEG({\Tile_X8Y0_S2BEG[7] ,
    \Tile_X8Y0_S2BEG[6] ,
    \Tile_X8Y0_S2BEG[5] ,
    \Tile_X8Y0_S2BEG[4] ,
    \Tile_X8Y0_S2BEG[3] ,
    \Tile_X8Y0_S2BEG[2] ,
    \Tile_X8Y0_S2BEG[1] ,
    \Tile_X8Y0_S2BEG[0] }),
    .S2BEGb({\Tile_X8Y0_S2BEGb[7] ,
    \Tile_X8Y0_S2BEGb[6] ,
    \Tile_X8Y0_S2BEGb[5] ,
    \Tile_X8Y0_S2BEGb[4] ,
    \Tile_X8Y0_S2BEGb[3] ,
    \Tile_X8Y0_S2BEGb[2] ,
    \Tile_X8Y0_S2BEGb[1] ,
    \Tile_X8Y0_S2BEGb[0] }),
    .S4BEG({\Tile_X8Y0_S4BEG[15] ,
    \Tile_X8Y0_S4BEG[14] ,
    \Tile_X8Y0_S4BEG[13] ,
    \Tile_X8Y0_S4BEG[12] ,
    \Tile_X8Y0_S4BEG[11] ,
    \Tile_X8Y0_S4BEG[10] ,
    \Tile_X8Y0_S4BEG[9] ,
    \Tile_X8Y0_S4BEG[8] ,
    \Tile_X8Y0_S4BEG[7] ,
    \Tile_X8Y0_S4BEG[6] ,
    \Tile_X8Y0_S4BEG[5] ,
    \Tile_X8Y0_S4BEG[4] ,
    \Tile_X8Y0_S4BEG[3] ,
    \Tile_X8Y0_S4BEG[2] ,
    \Tile_X8Y0_S4BEG[1] ,
    \Tile_X8Y0_S4BEG[0] }),
    .SS4BEG({\Tile_X8Y0_SS4BEG[15] ,
    \Tile_X8Y0_SS4BEG[14] ,
    \Tile_X8Y0_SS4BEG[13] ,
    \Tile_X8Y0_SS4BEG[12] ,
    \Tile_X8Y0_SS4BEG[11] ,
    \Tile_X8Y0_SS4BEG[10] ,
    \Tile_X8Y0_SS4BEG[9] ,
    \Tile_X8Y0_SS4BEG[8] ,
    \Tile_X8Y0_SS4BEG[7] ,
    \Tile_X8Y0_SS4BEG[6] ,
    \Tile_X8Y0_SS4BEG[5] ,
    \Tile_X8Y0_SS4BEG[4] ,
    \Tile_X8Y0_SS4BEG[3] ,
    \Tile_X8Y0_SS4BEG[2] ,
    \Tile_X8Y0_SS4BEG[1] ,
    \Tile_X8Y0_SS4BEG[0] }));
 LUT4AB Tile_X8Y10_LUT4AB (.Ci(Tile_X8Y11_Co),
    .Co(Tile_X8Y10_Co),
    .UserCLK(Tile_X8Y11_UserCLKo),
    .UserCLKo(Tile_X8Y10_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X8Y10_E1BEG[3] ,
    \Tile_X8Y10_E1BEG[2] ,
    \Tile_X8Y10_E1BEG[1] ,
    \Tile_X8Y10_E1BEG[0] }),
    .E1END({\Tile_X7Y10_E1BEG[3] ,
    \Tile_X7Y10_E1BEG[2] ,
    \Tile_X7Y10_E1BEG[1] ,
    \Tile_X7Y10_E1BEG[0] }),
    .E2BEG({\Tile_X8Y10_E2BEG[7] ,
    \Tile_X8Y10_E2BEG[6] ,
    \Tile_X8Y10_E2BEG[5] ,
    \Tile_X8Y10_E2BEG[4] ,
    \Tile_X8Y10_E2BEG[3] ,
    \Tile_X8Y10_E2BEG[2] ,
    \Tile_X8Y10_E2BEG[1] ,
    \Tile_X8Y10_E2BEG[0] }),
    .E2BEGb({\Tile_X8Y10_E2BEGb[7] ,
    \Tile_X8Y10_E2BEGb[6] ,
    \Tile_X8Y10_E2BEGb[5] ,
    \Tile_X8Y10_E2BEGb[4] ,
    \Tile_X8Y10_E2BEGb[3] ,
    \Tile_X8Y10_E2BEGb[2] ,
    \Tile_X8Y10_E2BEGb[1] ,
    \Tile_X8Y10_E2BEGb[0] }),
    .E2END({\Tile_X7Y10_E2BEGb[7] ,
    \Tile_X7Y10_E2BEGb[6] ,
    \Tile_X7Y10_E2BEGb[5] ,
    \Tile_X7Y10_E2BEGb[4] ,
    \Tile_X7Y10_E2BEGb[3] ,
    \Tile_X7Y10_E2BEGb[2] ,
    \Tile_X7Y10_E2BEGb[1] ,
    \Tile_X7Y10_E2BEGb[0] }),
    .E2MID({\Tile_X7Y10_E2BEG[7] ,
    \Tile_X7Y10_E2BEG[6] ,
    \Tile_X7Y10_E2BEG[5] ,
    \Tile_X7Y10_E2BEG[4] ,
    \Tile_X7Y10_E2BEG[3] ,
    \Tile_X7Y10_E2BEG[2] ,
    \Tile_X7Y10_E2BEG[1] ,
    \Tile_X7Y10_E2BEG[0] }),
    .E6BEG({\Tile_X8Y10_E6BEG[11] ,
    \Tile_X8Y10_E6BEG[10] ,
    \Tile_X8Y10_E6BEG[9] ,
    \Tile_X8Y10_E6BEG[8] ,
    \Tile_X8Y10_E6BEG[7] ,
    \Tile_X8Y10_E6BEG[6] ,
    \Tile_X8Y10_E6BEG[5] ,
    \Tile_X8Y10_E6BEG[4] ,
    \Tile_X8Y10_E6BEG[3] ,
    \Tile_X8Y10_E6BEG[2] ,
    \Tile_X8Y10_E6BEG[1] ,
    \Tile_X8Y10_E6BEG[0] }),
    .E6END({\Tile_X7Y10_E6BEG[11] ,
    \Tile_X7Y10_E6BEG[10] ,
    \Tile_X7Y10_E6BEG[9] ,
    \Tile_X7Y10_E6BEG[8] ,
    \Tile_X7Y10_E6BEG[7] ,
    \Tile_X7Y10_E6BEG[6] ,
    \Tile_X7Y10_E6BEG[5] ,
    \Tile_X7Y10_E6BEG[4] ,
    \Tile_X7Y10_E6BEG[3] ,
    \Tile_X7Y10_E6BEG[2] ,
    \Tile_X7Y10_E6BEG[1] ,
    \Tile_X7Y10_E6BEG[0] }),
    .EE4BEG({\Tile_X8Y10_EE4BEG[15] ,
    \Tile_X8Y10_EE4BEG[14] ,
    \Tile_X8Y10_EE4BEG[13] ,
    \Tile_X8Y10_EE4BEG[12] ,
    \Tile_X8Y10_EE4BEG[11] ,
    \Tile_X8Y10_EE4BEG[10] ,
    \Tile_X8Y10_EE4BEG[9] ,
    \Tile_X8Y10_EE4BEG[8] ,
    \Tile_X8Y10_EE4BEG[7] ,
    \Tile_X8Y10_EE4BEG[6] ,
    \Tile_X8Y10_EE4BEG[5] ,
    \Tile_X8Y10_EE4BEG[4] ,
    \Tile_X8Y10_EE4BEG[3] ,
    \Tile_X8Y10_EE4BEG[2] ,
    \Tile_X8Y10_EE4BEG[1] ,
    \Tile_X8Y10_EE4BEG[0] }),
    .EE4END({\Tile_X7Y10_EE4BEG[15] ,
    \Tile_X7Y10_EE4BEG[14] ,
    \Tile_X7Y10_EE4BEG[13] ,
    \Tile_X7Y10_EE4BEG[12] ,
    \Tile_X7Y10_EE4BEG[11] ,
    \Tile_X7Y10_EE4BEG[10] ,
    \Tile_X7Y10_EE4BEG[9] ,
    \Tile_X7Y10_EE4BEG[8] ,
    \Tile_X7Y10_EE4BEG[7] ,
    \Tile_X7Y10_EE4BEG[6] ,
    \Tile_X7Y10_EE4BEG[5] ,
    \Tile_X7Y10_EE4BEG[4] ,
    \Tile_X7Y10_EE4BEG[3] ,
    \Tile_X7Y10_EE4BEG[2] ,
    \Tile_X7Y10_EE4BEG[1] ,
    \Tile_X7Y10_EE4BEG[0] }),
    .FrameData({\Tile_X7Y10_FrameData_O[31] ,
    \Tile_X7Y10_FrameData_O[30] ,
    \Tile_X7Y10_FrameData_O[29] ,
    \Tile_X7Y10_FrameData_O[28] ,
    \Tile_X7Y10_FrameData_O[27] ,
    \Tile_X7Y10_FrameData_O[26] ,
    \Tile_X7Y10_FrameData_O[25] ,
    \Tile_X7Y10_FrameData_O[24] ,
    \Tile_X7Y10_FrameData_O[23] ,
    \Tile_X7Y10_FrameData_O[22] ,
    \Tile_X7Y10_FrameData_O[21] ,
    \Tile_X7Y10_FrameData_O[20] ,
    \Tile_X7Y10_FrameData_O[19] ,
    \Tile_X7Y10_FrameData_O[18] ,
    \Tile_X7Y10_FrameData_O[17] ,
    \Tile_X7Y10_FrameData_O[16] ,
    \Tile_X7Y10_FrameData_O[15] ,
    \Tile_X7Y10_FrameData_O[14] ,
    \Tile_X7Y10_FrameData_O[13] ,
    \Tile_X7Y10_FrameData_O[12] ,
    \Tile_X7Y10_FrameData_O[11] ,
    \Tile_X7Y10_FrameData_O[10] ,
    \Tile_X7Y10_FrameData_O[9] ,
    \Tile_X7Y10_FrameData_O[8] ,
    \Tile_X7Y10_FrameData_O[7] ,
    \Tile_X7Y10_FrameData_O[6] ,
    \Tile_X7Y10_FrameData_O[5] ,
    \Tile_X7Y10_FrameData_O[4] ,
    \Tile_X7Y10_FrameData_O[3] ,
    \Tile_X7Y10_FrameData_O[2] ,
    \Tile_X7Y10_FrameData_O[1] ,
    \Tile_X7Y10_FrameData_O[0] }),
    .FrameData_O({\Tile_X8Y10_FrameData_O[31] ,
    \Tile_X8Y10_FrameData_O[30] ,
    \Tile_X8Y10_FrameData_O[29] ,
    \Tile_X8Y10_FrameData_O[28] ,
    \Tile_X8Y10_FrameData_O[27] ,
    \Tile_X8Y10_FrameData_O[26] ,
    \Tile_X8Y10_FrameData_O[25] ,
    \Tile_X8Y10_FrameData_O[24] ,
    \Tile_X8Y10_FrameData_O[23] ,
    \Tile_X8Y10_FrameData_O[22] ,
    \Tile_X8Y10_FrameData_O[21] ,
    \Tile_X8Y10_FrameData_O[20] ,
    \Tile_X8Y10_FrameData_O[19] ,
    \Tile_X8Y10_FrameData_O[18] ,
    \Tile_X8Y10_FrameData_O[17] ,
    \Tile_X8Y10_FrameData_O[16] ,
    \Tile_X8Y10_FrameData_O[15] ,
    \Tile_X8Y10_FrameData_O[14] ,
    \Tile_X8Y10_FrameData_O[13] ,
    \Tile_X8Y10_FrameData_O[12] ,
    \Tile_X8Y10_FrameData_O[11] ,
    \Tile_X8Y10_FrameData_O[10] ,
    \Tile_X8Y10_FrameData_O[9] ,
    \Tile_X8Y10_FrameData_O[8] ,
    \Tile_X8Y10_FrameData_O[7] ,
    \Tile_X8Y10_FrameData_O[6] ,
    \Tile_X8Y10_FrameData_O[5] ,
    \Tile_X8Y10_FrameData_O[4] ,
    \Tile_X8Y10_FrameData_O[3] ,
    \Tile_X8Y10_FrameData_O[2] ,
    \Tile_X8Y10_FrameData_O[1] ,
    \Tile_X8Y10_FrameData_O[0] }),
    .FrameStrobe({\Tile_X8Y11_FrameStrobe_O[19] ,
    \Tile_X8Y11_FrameStrobe_O[18] ,
    \Tile_X8Y11_FrameStrobe_O[17] ,
    \Tile_X8Y11_FrameStrobe_O[16] ,
    \Tile_X8Y11_FrameStrobe_O[15] ,
    \Tile_X8Y11_FrameStrobe_O[14] ,
    \Tile_X8Y11_FrameStrobe_O[13] ,
    \Tile_X8Y11_FrameStrobe_O[12] ,
    \Tile_X8Y11_FrameStrobe_O[11] ,
    \Tile_X8Y11_FrameStrobe_O[10] ,
    \Tile_X8Y11_FrameStrobe_O[9] ,
    \Tile_X8Y11_FrameStrobe_O[8] ,
    \Tile_X8Y11_FrameStrobe_O[7] ,
    \Tile_X8Y11_FrameStrobe_O[6] ,
    \Tile_X8Y11_FrameStrobe_O[5] ,
    \Tile_X8Y11_FrameStrobe_O[4] ,
    \Tile_X8Y11_FrameStrobe_O[3] ,
    \Tile_X8Y11_FrameStrobe_O[2] ,
    \Tile_X8Y11_FrameStrobe_O[1] ,
    \Tile_X8Y11_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X8Y10_FrameStrobe_O[19] ,
    \Tile_X8Y10_FrameStrobe_O[18] ,
    \Tile_X8Y10_FrameStrobe_O[17] ,
    \Tile_X8Y10_FrameStrobe_O[16] ,
    \Tile_X8Y10_FrameStrobe_O[15] ,
    \Tile_X8Y10_FrameStrobe_O[14] ,
    \Tile_X8Y10_FrameStrobe_O[13] ,
    \Tile_X8Y10_FrameStrobe_O[12] ,
    \Tile_X8Y10_FrameStrobe_O[11] ,
    \Tile_X8Y10_FrameStrobe_O[10] ,
    \Tile_X8Y10_FrameStrobe_O[9] ,
    \Tile_X8Y10_FrameStrobe_O[8] ,
    \Tile_X8Y10_FrameStrobe_O[7] ,
    \Tile_X8Y10_FrameStrobe_O[6] ,
    \Tile_X8Y10_FrameStrobe_O[5] ,
    \Tile_X8Y10_FrameStrobe_O[4] ,
    \Tile_X8Y10_FrameStrobe_O[3] ,
    \Tile_X8Y10_FrameStrobe_O[2] ,
    \Tile_X8Y10_FrameStrobe_O[1] ,
    \Tile_X8Y10_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X8Y10_N1BEG[3] ,
    \Tile_X8Y10_N1BEG[2] ,
    \Tile_X8Y10_N1BEG[1] ,
    \Tile_X8Y10_N1BEG[0] }),
    .N1END({\Tile_X8Y11_N1BEG[3] ,
    \Tile_X8Y11_N1BEG[2] ,
    \Tile_X8Y11_N1BEG[1] ,
    \Tile_X8Y11_N1BEG[0] }),
    .N2BEG({\Tile_X8Y10_N2BEG[7] ,
    \Tile_X8Y10_N2BEG[6] ,
    \Tile_X8Y10_N2BEG[5] ,
    \Tile_X8Y10_N2BEG[4] ,
    \Tile_X8Y10_N2BEG[3] ,
    \Tile_X8Y10_N2BEG[2] ,
    \Tile_X8Y10_N2BEG[1] ,
    \Tile_X8Y10_N2BEG[0] }),
    .N2BEGb({\Tile_X8Y10_N2BEGb[7] ,
    \Tile_X8Y10_N2BEGb[6] ,
    \Tile_X8Y10_N2BEGb[5] ,
    \Tile_X8Y10_N2BEGb[4] ,
    \Tile_X8Y10_N2BEGb[3] ,
    \Tile_X8Y10_N2BEGb[2] ,
    \Tile_X8Y10_N2BEGb[1] ,
    \Tile_X8Y10_N2BEGb[0] }),
    .N2END({\Tile_X8Y11_N2BEGb[7] ,
    \Tile_X8Y11_N2BEGb[6] ,
    \Tile_X8Y11_N2BEGb[5] ,
    \Tile_X8Y11_N2BEGb[4] ,
    \Tile_X8Y11_N2BEGb[3] ,
    \Tile_X8Y11_N2BEGb[2] ,
    \Tile_X8Y11_N2BEGb[1] ,
    \Tile_X8Y11_N2BEGb[0] }),
    .N2MID({\Tile_X8Y11_N2BEG[7] ,
    \Tile_X8Y11_N2BEG[6] ,
    \Tile_X8Y11_N2BEG[5] ,
    \Tile_X8Y11_N2BEG[4] ,
    \Tile_X8Y11_N2BEG[3] ,
    \Tile_X8Y11_N2BEG[2] ,
    \Tile_X8Y11_N2BEG[1] ,
    \Tile_X8Y11_N2BEG[0] }),
    .N4BEG({\Tile_X8Y10_N4BEG[15] ,
    \Tile_X8Y10_N4BEG[14] ,
    \Tile_X8Y10_N4BEG[13] ,
    \Tile_X8Y10_N4BEG[12] ,
    \Tile_X8Y10_N4BEG[11] ,
    \Tile_X8Y10_N4BEG[10] ,
    \Tile_X8Y10_N4BEG[9] ,
    \Tile_X8Y10_N4BEG[8] ,
    \Tile_X8Y10_N4BEG[7] ,
    \Tile_X8Y10_N4BEG[6] ,
    \Tile_X8Y10_N4BEG[5] ,
    \Tile_X8Y10_N4BEG[4] ,
    \Tile_X8Y10_N4BEG[3] ,
    \Tile_X8Y10_N4BEG[2] ,
    \Tile_X8Y10_N4BEG[1] ,
    \Tile_X8Y10_N4BEG[0] }),
    .N4END({\Tile_X8Y11_N4BEG[15] ,
    \Tile_X8Y11_N4BEG[14] ,
    \Tile_X8Y11_N4BEG[13] ,
    \Tile_X8Y11_N4BEG[12] ,
    \Tile_X8Y11_N4BEG[11] ,
    \Tile_X8Y11_N4BEG[10] ,
    \Tile_X8Y11_N4BEG[9] ,
    \Tile_X8Y11_N4BEG[8] ,
    \Tile_X8Y11_N4BEG[7] ,
    \Tile_X8Y11_N4BEG[6] ,
    \Tile_X8Y11_N4BEG[5] ,
    \Tile_X8Y11_N4BEG[4] ,
    \Tile_X8Y11_N4BEG[3] ,
    \Tile_X8Y11_N4BEG[2] ,
    \Tile_X8Y11_N4BEG[1] ,
    \Tile_X8Y11_N4BEG[0] }),
    .NN4BEG({\Tile_X8Y10_NN4BEG[15] ,
    \Tile_X8Y10_NN4BEG[14] ,
    \Tile_X8Y10_NN4BEG[13] ,
    \Tile_X8Y10_NN4BEG[12] ,
    \Tile_X8Y10_NN4BEG[11] ,
    \Tile_X8Y10_NN4BEG[10] ,
    \Tile_X8Y10_NN4BEG[9] ,
    \Tile_X8Y10_NN4BEG[8] ,
    \Tile_X8Y10_NN4BEG[7] ,
    \Tile_X8Y10_NN4BEG[6] ,
    \Tile_X8Y10_NN4BEG[5] ,
    \Tile_X8Y10_NN4BEG[4] ,
    \Tile_X8Y10_NN4BEG[3] ,
    \Tile_X8Y10_NN4BEG[2] ,
    \Tile_X8Y10_NN4BEG[1] ,
    \Tile_X8Y10_NN4BEG[0] }),
    .NN4END({\Tile_X8Y11_NN4BEG[15] ,
    \Tile_X8Y11_NN4BEG[14] ,
    \Tile_X8Y11_NN4BEG[13] ,
    \Tile_X8Y11_NN4BEG[12] ,
    \Tile_X8Y11_NN4BEG[11] ,
    \Tile_X8Y11_NN4BEG[10] ,
    \Tile_X8Y11_NN4BEG[9] ,
    \Tile_X8Y11_NN4BEG[8] ,
    \Tile_X8Y11_NN4BEG[7] ,
    \Tile_X8Y11_NN4BEG[6] ,
    \Tile_X8Y11_NN4BEG[5] ,
    \Tile_X8Y11_NN4BEG[4] ,
    \Tile_X8Y11_NN4BEG[3] ,
    \Tile_X8Y11_NN4BEG[2] ,
    \Tile_X8Y11_NN4BEG[1] ,
    \Tile_X8Y11_NN4BEG[0] }),
    .S1BEG({\Tile_X8Y10_S1BEG[3] ,
    \Tile_X8Y10_S1BEG[2] ,
    \Tile_X8Y10_S1BEG[1] ,
    \Tile_X8Y10_S1BEG[0] }),
    .S1END({\Tile_X8Y9_S1BEG[3] ,
    \Tile_X8Y9_S1BEG[2] ,
    \Tile_X8Y9_S1BEG[1] ,
    \Tile_X8Y9_S1BEG[0] }),
    .S2BEG({\Tile_X8Y10_S2BEG[7] ,
    \Tile_X8Y10_S2BEG[6] ,
    \Tile_X8Y10_S2BEG[5] ,
    \Tile_X8Y10_S2BEG[4] ,
    \Tile_X8Y10_S2BEG[3] ,
    \Tile_X8Y10_S2BEG[2] ,
    \Tile_X8Y10_S2BEG[1] ,
    \Tile_X8Y10_S2BEG[0] }),
    .S2BEGb({\Tile_X8Y10_S2BEGb[7] ,
    \Tile_X8Y10_S2BEGb[6] ,
    \Tile_X8Y10_S2BEGb[5] ,
    \Tile_X8Y10_S2BEGb[4] ,
    \Tile_X8Y10_S2BEGb[3] ,
    \Tile_X8Y10_S2BEGb[2] ,
    \Tile_X8Y10_S2BEGb[1] ,
    \Tile_X8Y10_S2BEGb[0] }),
    .S2END({\Tile_X8Y9_S2BEGb[7] ,
    \Tile_X8Y9_S2BEGb[6] ,
    \Tile_X8Y9_S2BEGb[5] ,
    \Tile_X8Y9_S2BEGb[4] ,
    \Tile_X8Y9_S2BEGb[3] ,
    \Tile_X8Y9_S2BEGb[2] ,
    \Tile_X8Y9_S2BEGb[1] ,
    \Tile_X8Y9_S2BEGb[0] }),
    .S2MID({\Tile_X8Y9_S2BEG[7] ,
    \Tile_X8Y9_S2BEG[6] ,
    \Tile_X8Y9_S2BEG[5] ,
    \Tile_X8Y9_S2BEG[4] ,
    \Tile_X8Y9_S2BEG[3] ,
    \Tile_X8Y9_S2BEG[2] ,
    \Tile_X8Y9_S2BEG[1] ,
    \Tile_X8Y9_S2BEG[0] }),
    .S4BEG({\Tile_X8Y10_S4BEG[15] ,
    \Tile_X8Y10_S4BEG[14] ,
    \Tile_X8Y10_S4BEG[13] ,
    \Tile_X8Y10_S4BEG[12] ,
    \Tile_X8Y10_S4BEG[11] ,
    \Tile_X8Y10_S4BEG[10] ,
    \Tile_X8Y10_S4BEG[9] ,
    \Tile_X8Y10_S4BEG[8] ,
    \Tile_X8Y10_S4BEG[7] ,
    \Tile_X8Y10_S4BEG[6] ,
    \Tile_X8Y10_S4BEG[5] ,
    \Tile_X8Y10_S4BEG[4] ,
    \Tile_X8Y10_S4BEG[3] ,
    \Tile_X8Y10_S4BEG[2] ,
    \Tile_X8Y10_S4BEG[1] ,
    \Tile_X8Y10_S4BEG[0] }),
    .S4END({\Tile_X8Y9_S4BEG[15] ,
    \Tile_X8Y9_S4BEG[14] ,
    \Tile_X8Y9_S4BEG[13] ,
    \Tile_X8Y9_S4BEG[12] ,
    \Tile_X8Y9_S4BEG[11] ,
    \Tile_X8Y9_S4BEG[10] ,
    \Tile_X8Y9_S4BEG[9] ,
    \Tile_X8Y9_S4BEG[8] ,
    \Tile_X8Y9_S4BEG[7] ,
    \Tile_X8Y9_S4BEG[6] ,
    \Tile_X8Y9_S4BEG[5] ,
    \Tile_X8Y9_S4BEG[4] ,
    \Tile_X8Y9_S4BEG[3] ,
    \Tile_X8Y9_S4BEG[2] ,
    \Tile_X8Y9_S4BEG[1] ,
    \Tile_X8Y9_S4BEG[0] }),
    .SS4BEG({\Tile_X8Y10_SS4BEG[15] ,
    \Tile_X8Y10_SS4BEG[14] ,
    \Tile_X8Y10_SS4BEG[13] ,
    \Tile_X8Y10_SS4BEG[12] ,
    \Tile_X8Y10_SS4BEG[11] ,
    \Tile_X8Y10_SS4BEG[10] ,
    \Tile_X8Y10_SS4BEG[9] ,
    \Tile_X8Y10_SS4BEG[8] ,
    \Tile_X8Y10_SS4BEG[7] ,
    \Tile_X8Y10_SS4BEG[6] ,
    \Tile_X8Y10_SS4BEG[5] ,
    \Tile_X8Y10_SS4BEG[4] ,
    \Tile_X8Y10_SS4BEG[3] ,
    \Tile_X8Y10_SS4BEG[2] ,
    \Tile_X8Y10_SS4BEG[1] ,
    \Tile_X8Y10_SS4BEG[0] }),
    .SS4END({\Tile_X8Y9_SS4BEG[15] ,
    \Tile_X8Y9_SS4BEG[14] ,
    \Tile_X8Y9_SS4BEG[13] ,
    \Tile_X8Y9_SS4BEG[12] ,
    \Tile_X8Y9_SS4BEG[11] ,
    \Tile_X8Y9_SS4BEG[10] ,
    \Tile_X8Y9_SS4BEG[9] ,
    \Tile_X8Y9_SS4BEG[8] ,
    \Tile_X8Y9_SS4BEG[7] ,
    \Tile_X8Y9_SS4BEG[6] ,
    \Tile_X8Y9_SS4BEG[5] ,
    \Tile_X8Y9_SS4BEG[4] ,
    \Tile_X8Y9_SS4BEG[3] ,
    \Tile_X8Y9_SS4BEG[2] ,
    \Tile_X8Y9_SS4BEG[1] ,
    \Tile_X8Y9_SS4BEG[0] }),
    .W1BEG({\Tile_X8Y10_W1BEG[3] ,
    \Tile_X8Y10_W1BEG[2] ,
    \Tile_X8Y10_W1BEG[1] ,
    \Tile_X8Y10_W1BEG[0] }),
    .W1END({\Tile_X9Y10_W1BEG[3] ,
    \Tile_X9Y10_W1BEG[2] ,
    \Tile_X9Y10_W1BEG[1] ,
    \Tile_X9Y10_W1BEG[0] }),
    .W2BEG({\Tile_X8Y10_W2BEG[7] ,
    \Tile_X8Y10_W2BEG[6] ,
    \Tile_X8Y10_W2BEG[5] ,
    \Tile_X8Y10_W2BEG[4] ,
    \Tile_X8Y10_W2BEG[3] ,
    \Tile_X8Y10_W2BEG[2] ,
    \Tile_X8Y10_W2BEG[1] ,
    \Tile_X8Y10_W2BEG[0] }),
    .W2BEGb({\Tile_X8Y10_W2BEGb[7] ,
    \Tile_X8Y10_W2BEGb[6] ,
    \Tile_X8Y10_W2BEGb[5] ,
    \Tile_X8Y10_W2BEGb[4] ,
    \Tile_X8Y10_W2BEGb[3] ,
    \Tile_X8Y10_W2BEGb[2] ,
    \Tile_X8Y10_W2BEGb[1] ,
    \Tile_X8Y10_W2BEGb[0] }),
    .W2END({\Tile_X9Y10_W2BEGb[7] ,
    \Tile_X9Y10_W2BEGb[6] ,
    \Tile_X9Y10_W2BEGb[5] ,
    \Tile_X9Y10_W2BEGb[4] ,
    \Tile_X9Y10_W2BEGb[3] ,
    \Tile_X9Y10_W2BEGb[2] ,
    \Tile_X9Y10_W2BEGb[1] ,
    \Tile_X9Y10_W2BEGb[0] }),
    .W2MID({\Tile_X9Y10_W2BEG[7] ,
    \Tile_X9Y10_W2BEG[6] ,
    \Tile_X9Y10_W2BEG[5] ,
    \Tile_X9Y10_W2BEG[4] ,
    \Tile_X9Y10_W2BEG[3] ,
    \Tile_X9Y10_W2BEG[2] ,
    \Tile_X9Y10_W2BEG[1] ,
    \Tile_X9Y10_W2BEG[0] }),
    .W6BEG({\Tile_X8Y10_W6BEG[11] ,
    \Tile_X8Y10_W6BEG[10] ,
    \Tile_X8Y10_W6BEG[9] ,
    \Tile_X8Y10_W6BEG[8] ,
    \Tile_X8Y10_W6BEG[7] ,
    \Tile_X8Y10_W6BEG[6] ,
    \Tile_X8Y10_W6BEG[5] ,
    \Tile_X8Y10_W6BEG[4] ,
    \Tile_X8Y10_W6BEG[3] ,
    \Tile_X8Y10_W6BEG[2] ,
    \Tile_X8Y10_W6BEG[1] ,
    \Tile_X8Y10_W6BEG[0] }),
    .W6END({\Tile_X9Y10_W6BEG[11] ,
    \Tile_X9Y10_W6BEG[10] ,
    \Tile_X9Y10_W6BEG[9] ,
    \Tile_X9Y10_W6BEG[8] ,
    \Tile_X9Y10_W6BEG[7] ,
    \Tile_X9Y10_W6BEG[6] ,
    \Tile_X9Y10_W6BEG[5] ,
    \Tile_X9Y10_W6BEG[4] ,
    \Tile_X9Y10_W6BEG[3] ,
    \Tile_X9Y10_W6BEG[2] ,
    \Tile_X9Y10_W6BEG[1] ,
    \Tile_X9Y10_W6BEG[0] }),
    .WW4BEG({\Tile_X8Y10_WW4BEG[15] ,
    \Tile_X8Y10_WW4BEG[14] ,
    \Tile_X8Y10_WW4BEG[13] ,
    \Tile_X8Y10_WW4BEG[12] ,
    \Tile_X8Y10_WW4BEG[11] ,
    \Tile_X8Y10_WW4BEG[10] ,
    \Tile_X8Y10_WW4BEG[9] ,
    \Tile_X8Y10_WW4BEG[8] ,
    \Tile_X8Y10_WW4BEG[7] ,
    \Tile_X8Y10_WW4BEG[6] ,
    \Tile_X8Y10_WW4BEG[5] ,
    \Tile_X8Y10_WW4BEG[4] ,
    \Tile_X8Y10_WW4BEG[3] ,
    \Tile_X8Y10_WW4BEG[2] ,
    \Tile_X8Y10_WW4BEG[1] ,
    \Tile_X8Y10_WW4BEG[0] }),
    .WW4END({\Tile_X9Y10_WW4BEG[15] ,
    \Tile_X9Y10_WW4BEG[14] ,
    \Tile_X9Y10_WW4BEG[13] ,
    \Tile_X9Y10_WW4BEG[12] ,
    \Tile_X9Y10_WW4BEG[11] ,
    \Tile_X9Y10_WW4BEG[10] ,
    \Tile_X9Y10_WW4BEG[9] ,
    \Tile_X9Y10_WW4BEG[8] ,
    \Tile_X9Y10_WW4BEG[7] ,
    \Tile_X9Y10_WW4BEG[6] ,
    \Tile_X9Y10_WW4BEG[5] ,
    \Tile_X9Y10_WW4BEG[4] ,
    \Tile_X9Y10_WW4BEG[3] ,
    \Tile_X9Y10_WW4BEG[2] ,
    \Tile_X9Y10_WW4BEG[1] ,
    \Tile_X9Y10_WW4BEG[0] }));
 LUT4AB Tile_X8Y11_LUT4AB (.Ci(Tile_X8Y12_Co),
    .Co(Tile_X8Y11_Co),
    .UserCLK(Tile_X8Y12_UserCLKo),
    .UserCLKo(Tile_X8Y11_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X8Y11_E1BEG[3] ,
    \Tile_X8Y11_E1BEG[2] ,
    \Tile_X8Y11_E1BEG[1] ,
    \Tile_X8Y11_E1BEG[0] }),
    .E1END({\Tile_X7Y11_E1BEG[3] ,
    \Tile_X7Y11_E1BEG[2] ,
    \Tile_X7Y11_E1BEG[1] ,
    \Tile_X7Y11_E1BEG[0] }),
    .E2BEG({\Tile_X8Y11_E2BEG[7] ,
    \Tile_X8Y11_E2BEG[6] ,
    \Tile_X8Y11_E2BEG[5] ,
    \Tile_X8Y11_E2BEG[4] ,
    \Tile_X8Y11_E2BEG[3] ,
    \Tile_X8Y11_E2BEG[2] ,
    \Tile_X8Y11_E2BEG[1] ,
    \Tile_X8Y11_E2BEG[0] }),
    .E2BEGb({\Tile_X8Y11_E2BEGb[7] ,
    \Tile_X8Y11_E2BEGb[6] ,
    \Tile_X8Y11_E2BEGb[5] ,
    \Tile_X8Y11_E2BEGb[4] ,
    \Tile_X8Y11_E2BEGb[3] ,
    \Tile_X8Y11_E2BEGb[2] ,
    \Tile_X8Y11_E2BEGb[1] ,
    \Tile_X8Y11_E2BEGb[0] }),
    .E2END({\Tile_X7Y11_E2BEGb[7] ,
    \Tile_X7Y11_E2BEGb[6] ,
    \Tile_X7Y11_E2BEGb[5] ,
    \Tile_X7Y11_E2BEGb[4] ,
    \Tile_X7Y11_E2BEGb[3] ,
    \Tile_X7Y11_E2BEGb[2] ,
    \Tile_X7Y11_E2BEGb[1] ,
    \Tile_X7Y11_E2BEGb[0] }),
    .E2MID({\Tile_X7Y11_E2BEG[7] ,
    \Tile_X7Y11_E2BEG[6] ,
    \Tile_X7Y11_E2BEG[5] ,
    \Tile_X7Y11_E2BEG[4] ,
    \Tile_X7Y11_E2BEG[3] ,
    \Tile_X7Y11_E2BEG[2] ,
    \Tile_X7Y11_E2BEG[1] ,
    \Tile_X7Y11_E2BEG[0] }),
    .E6BEG({\Tile_X8Y11_E6BEG[11] ,
    \Tile_X8Y11_E6BEG[10] ,
    \Tile_X8Y11_E6BEG[9] ,
    \Tile_X8Y11_E6BEG[8] ,
    \Tile_X8Y11_E6BEG[7] ,
    \Tile_X8Y11_E6BEG[6] ,
    \Tile_X8Y11_E6BEG[5] ,
    \Tile_X8Y11_E6BEG[4] ,
    \Tile_X8Y11_E6BEG[3] ,
    \Tile_X8Y11_E6BEG[2] ,
    \Tile_X8Y11_E6BEG[1] ,
    \Tile_X8Y11_E6BEG[0] }),
    .E6END({\Tile_X7Y11_E6BEG[11] ,
    \Tile_X7Y11_E6BEG[10] ,
    \Tile_X7Y11_E6BEG[9] ,
    \Tile_X7Y11_E6BEG[8] ,
    \Tile_X7Y11_E6BEG[7] ,
    \Tile_X7Y11_E6BEG[6] ,
    \Tile_X7Y11_E6BEG[5] ,
    \Tile_X7Y11_E6BEG[4] ,
    \Tile_X7Y11_E6BEG[3] ,
    \Tile_X7Y11_E6BEG[2] ,
    \Tile_X7Y11_E6BEG[1] ,
    \Tile_X7Y11_E6BEG[0] }),
    .EE4BEG({\Tile_X8Y11_EE4BEG[15] ,
    \Tile_X8Y11_EE4BEG[14] ,
    \Tile_X8Y11_EE4BEG[13] ,
    \Tile_X8Y11_EE4BEG[12] ,
    \Tile_X8Y11_EE4BEG[11] ,
    \Tile_X8Y11_EE4BEG[10] ,
    \Tile_X8Y11_EE4BEG[9] ,
    \Tile_X8Y11_EE4BEG[8] ,
    \Tile_X8Y11_EE4BEG[7] ,
    \Tile_X8Y11_EE4BEG[6] ,
    \Tile_X8Y11_EE4BEG[5] ,
    \Tile_X8Y11_EE4BEG[4] ,
    \Tile_X8Y11_EE4BEG[3] ,
    \Tile_X8Y11_EE4BEG[2] ,
    \Tile_X8Y11_EE4BEG[1] ,
    \Tile_X8Y11_EE4BEG[0] }),
    .EE4END({\Tile_X7Y11_EE4BEG[15] ,
    \Tile_X7Y11_EE4BEG[14] ,
    \Tile_X7Y11_EE4BEG[13] ,
    \Tile_X7Y11_EE4BEG[12] ,
    \Tile_X7Y11_EE4BEG[11] ,
    \Tile_X7Y11_EE4BEG[10] ,
    \Tile_X7Y11_EE4BEG[9] ,
    \Tile_X7Y11_EE4BEG[8] ,
    \Tile_X7Y11_EE4BEG[7] ,
    \Tile_X7Y11_EE4BEG[6] ,
    \Tile_X7Y11_EE4BEG[5] ,
    \Tile_X7Y11_EE4BEG[4] ,
    \Tile_X7Y11_EE4BEG[3] ,
    \Tile_X7Y11_EE4BEG[2] ,
    \Tile_X7Y11_EE4BEG[1] ,
    \Tile_X7Y11_EE4BEG[0] }),
    .FrameData({\Tile_X7Y11_FrameData_O[31] ,
    \Tile_X7Y11_FrameData_O[30] ,
    \Tile_X7Y11_FrameData_O[29] ,
    \Tile_X7Y11_FrameData_O[28] ,
    \Tile_X7Y11_FrameData_O[27] ,
    \Tile_X7Y11_FrameData_O[26] ,
    \Tile_X7Y11_FrameData_O[25] ,
    \Tile_X7Y11_FrameData_O[24] ,
    \Tile_X7Y11_FrameData_O[23] ,
    \Tile_X7Y11_FrameData_O[22] ,
    \Tile_X7Y11_FrameData_O[21] ,
    \Tile_X7Y11_FrameData_O[20] ,
    \Tile_X7Y11_FrameData_O[19] ,
    \Tile_X7Y11_FrameData_O[18] ,
    \Tile_X7Y11_FrameData_O[17] ,
    \Tile_X7Y11_FrameData_O[16] ,
    \Tile_X7Y11_FrameData_O[15] ,
    \Tile_X7Y11_FrameData_O[14] ,
    \Tile_X7Y11_FrameData_O[13] ,
    \Tile_X7Y11_FrameData_O[12] ,
    \Tile_X7Y11_FrameData_O[11] ,
    \Tile_X7Y11_FrameData_O[10] ,
    \Tile_X7Y11_FrameData_O[9] ,
    \Tile_X7Y11_FrameData_O[8] ,
    \Tile_X7Y11_FrameData_O[7] ,
    \Tile_X7Y11_FrameData_O[6] ,
    \Tile_X7Y11_FrameData_O[5] ,
    \Tile_X7Y11_FrameData_O[4] ,
    \Tile_X7Y11_FrameData_O[3] ,
    \Tile_X7Y11_FrameData_O[2] ,
    \Tile_X7Y11_FrameData_O[1] ,
    \Tile_X7Y11_FrameData_O[0] }),
    .FrameData_O({\Tile_X8Y11_FrameData_O[31] ,
    \Tile_X8Y11_FrameData_O[30] ,
    \Tile_X8Y11_FrameData_O[29] ,
    \Tile_X8Y11_FrameData_O[28] ,
    \Tile_X8Y11_FrameData_O[27] ,
    \Tile_X8Y11_FrameData_O[26] ,
    \Tile_X8Y11_FrameData_O[25] ,
    \Tile_X8Y11_FrameData_O[24] ,
    \Tile_X8Y11_FrameData_O[23] ,
    \Tile_X8Y11_FrameData_O[22] ,
    \Tile_X8Y11_FrameData_O[21] ,
    \Tile_X8Y11_FrameData_O[20] ,
    \Tile_X8Y11_FrameData_O[19] ,
    \Tile_X8Y11_FrameData_O[18] ,
    \Tile_X8Y11_FrameData_O[17] ,
    \Tile_X8Y11_FrameData_O[16] ,
    \Tile_X8Y11_FrameData_O[15] ,
    \Tile_X8Y11_FrameData_O[14] ,
    \Tile_X8Y11_FrameData_O[13] ,
    \Tile_X8Y11_FrameData_O[12] ,
    \Tile_X8Y11_FrameData_O[11] ,
    \Tile_X8Y11_FrameData_O[10] ,
    \Tile_X8Y11_FrameData_O[9] ,
    \Tile_X8Y11_FrameData_O[8] ,
    \Tile_X8Y11_FrameData_O[7] ,
    \Tile_X8Y11_FrameData_O[6] ,
    \Tile_X8Y11_FrameData_O[5] ,
    \Tile_X8Y11_FrameData_O[4] ,
    \Tile_X8Y11_FrameData_O[3] ,
    \Tile_X8Y11_FrameData_O[2] ,
    \Tile_X8Y11_FrameData_O[1] ,
    \Tile_X8Y11_FrameData_O[0] }),
    .FrameStrobe({\Tile_X8Y12_FrameStrobe_O[19] ,
    \Tile_X8Y12_FrameStrobe_O[18] ,
    \Tile_X8Y12_FrameStrobe_O[17] ,
    \Tile_X8Y12_FrameStrobe_O[16] ,
    \Tile_X8Y12_FrameStrobe_O[15] ,
    \Tile_X8Y12_FrameStrobe_O[14] ,
    \Tile_X8Y12_FrameStrobe_O[13] ,
    \Tile_X8Y12_FrameStrobe_O[12] ,
    \Tile_X8Y12_FrameStrobe_O[11] ,
    \Tile_X8Y12_FrameStrobe_O[10] ,
    \Tile_X8Y12_FrameStrobe_O[9] ,
    \Tile_X8Y12_FrameStrobe_O[8] ,
    \Tile_X8Y12_FrameStrobe_O[7] ,
    \Tile_X8Y12_FrameStrobe_O[6] ,
    \Tile_X8Y12_FrameStrobe_O[5] ,
    \Tile_X8Y12_FrameStrobe_O[4] ,
    \Tile_X8Y12_FrameStrobe_O[3] ,
    \Tile_X8Y12_FrameStrobe_O[2] ,
    \Tile_X8Y12_FrameStrobe_O[1] ,
    \Tile_X8Y12_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X8Y11_FrameStrobe_O[19] ,
    \Tile_X8Y11_FrameStrobe_O[18] ,
    \Tile_X8Y11_FrameStrobe_O[17] ,
    \Tile_X8Y11_FrameStrobe_O[16] ,
    \Tile_X8Y11_FrameStrobe_O[15] ,
    \Tile_X8Y11_FrameStrobe_O[14] ,
    \Tile_X8Y11_FrameStrobe_O[13] ,
    \Tile_X8Y11_FrameStrobe_O[12] ,
    \Tile_X8Y11_FrameStrobe_O[11] ,
    \Tile_X8Y11_FrameStrobe_O[10] ,
    \Tile_X8Y11_FrameStrobe_O[9] ,
    \Tile_X8Y11_FrameStrobe_O[8] ,
    \Tile_X8Y11_FrameStrobe_O[7] ,
    \Tile_X8Y11_FrameStrobe_O[6] ,
    \Tile_X8Y11_FrameStrobe_O[5] ,
    \Tile_X8Y11_FrameStrobe_O[4] ,
    \Tile_X8Y11_FrameStrobe_O[3] ,
    \Tile_X8Y11_FrameStrobe_O[2] ,
    \Tile_X8Y11_FrameStrobe_O[1] ,
    \Tile_X8Y11_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X8Y11_N1BEG[3] ,
    \Tile_X8Y11_N1BEG[2] ,
    \Tile_X8Y11_N1BEG[1] ,
    \Tile_X8Y11_N1BEG[0] }),
    .N1END({\Tile_X8Y12_N1BEG[3] ,
    \Tile_X8Y12_N1BEG[2] ,
    \Tile_X8Y12_N1BEG[1] ,
    \Tile_X8Y12_N1BEG[0] }),
    .N2BEG({\Tile_X8Y11_N2BEG[7] ,
    \Tile_X8Y11_N2BEG[6] ,
    \Tile_X8Y11_N2BEG[5] ,
    \Tile_X8Y11_N2BEG[4] ,
    \Tile_X8Y11_N2BEG[3] ,
    \Tile_X8Y11_N2BEG[2] ,
    \Tile_X8Y11_N2BEG[1] ,
    \Tile_X8Y11_N2BEG[0] }),
    .N2BEGb({\Tile_X8Y11_N2BEGb[7] ,
    \Tile_X8Y11_N2BEGb[6] ,
    \Tile_X8Y11_N2BEGb[5] ,
    \Tile_X8Y11_N2BEGb[4] ,
    \Tile_X8Y11_N2BEGb[3] ,
    \Tile_X8Y11_N2BEGb[2] ,
    \Tile_X8Y11_N2BEGb[1] ,
    \Tile_X8Y11_N2BEGb[0] }),
    .N2END({\Tile_X8Y12_N2BEGb[7] ,
    \Tile_X8Y12_N2BEGb[6] ,
    \Tile_X8Y12_N2BEGb[5] ,
    \Tile_X8Y12_N2BEGb[4] ,
    \Tile_X8Y12_N2BEGb[3] ,
    \Tile_X8Y12_N2BEGb[2] ,
    \Tile_X8Y12_N2BEGb[1] ,
    \Tile_X8Y12_N2BEGb[0] }),
    .N2MID({\Tile_X8Y12_N2BEG[7] ,
    \Tile_X8Y12_N2BEG[6] ,
    \Tile_X8Y12_N2BEG[5] ,
    \Tile_X8Y12_N2BEG[4] ,
    \Tile_X8Y12_N2BEG[3] ,
    \Tile_X8Y12_N2BEG[2] ,
    \Tile_X8Y12_N2BEG[1] ,
    \Tile_X8Y12_N2BEG[0] }),
    .N4BEG({\Tile_X8Y11_N4BEG[15] ,
    \Tile_X8Y11_N4BEG[14] ,
    \Tile_X8Y11_N4BEG[13] ,
    \Tile_X8Y11_N4BEG[12] ,
    \Tile_X8Y11_N4BEG[11] ,
    \Tile_X8Y11_N4BEG[10] ,
    \Tile_X8Y11_N4BEG[9] ,
    \Tile_X8Y11_N4BEG[8] ,
    \Tile_X8Y11_N4BEG[7] ,
    \Tile_X8Y11_N4BEG[6] ,
    \Tile_X8Y11_N4BEG[5] ,
    \Tile_X8Y11_N4BEG[4] ,
    \Tile_X8Y11_N4BEG[3] ,
    \Tile_X8Y11_N4BEG[2] ,
    \Tile_X8Y11_N4BEG[1] ,
    \Tile_X8Y11_N4BEG[0] }),
    .N4END({\Tile_X8Y12_N4BEG[15] ,
    \Tile_X8Y12_N4BEG[14] ,
    \Tile_X8Y12_N4BEG[13] ,
    \Tile_X8Y12_N4BEG[12] ,
    \Tile_X8Y12_N4BEG[11] ,
    \Tile_X8Y12_N4BEG[10] ,
    \Tile_X8Y12_N4BEG[9] ,
    \Tile_X8Y12_N4BEG[8] ,
    \Tile_X8Y12_N4BEG[7] ,
    \Tile_X8Y12_N4BEG[6] ,
    \Tile_X8Y12_N4BEG[5] ,
    \Tile_X8Y12_N4BEG[4] ,
    \Tile_X8Y12_N4BEG[3] ,
    \Tile_X8Y12_N4BEG[2] ,
    \Tile_X8Y12_N4BEG[1] ,
    \Tile_X8Y12_N4BEG[0] }),
    .NN4BEG({\Tile_X8Y11_NN4BEG[15] ,
    \Tile_X8Y11_NN4BEG[14] ,
    \Tile_X8Y11_NN4BEG[13] ,
    \Tile_X8Y11_NN4BEG[12] ,
    \Tile_X8Y11_NN4BEG[11] ,
    \Tile_X8Y11_NN4BEG[10] ,
    \Tile_X8Y11_NN4BEG[9] ,
    \Tile_X8Y11_NN4BEG[8] ,
    \Tile_X8Y11_NN4BEG[7] ,
    \Tile_X8Y11_NN4BEG[6] ,
    \Tile_X8Y11_NN4BEG[5] ,
    \Tile_X8Y11_NN4BEG[4] ,
    \Tile_X8Y11_NN4BEG[3] ,
    \Tile_X8Y11_NN4BEG[2] ,
    \Tile_X8Y11_NN4BEG[1] ,
    \Tile_X8Y11_NN4BEG[0] }),
    .NN4END({\Tile_X8Y12_NN4BEG[15] ,
    \Tile_X8Y12_NN4BEG[14] ,
    \Tile_X8Y12_NN4BEG[13] ,
    \Tile_X8Y12_NN4BEG[12] ,
    \Tile_X8Y12_NN4BEG[11] ,
    \Tile_X8Y12_NN4BEG[10] ,
    \Tile_X8Y12_NN4BEG[9] ,
    \Tile_X8Y12_NN4BEG[8] ,
    \Tile_X8Y12_NN4BEG[7] ,
    \Tile_X8Y12_NN4BEG[6] ,
    \Tile_X8Y12_NN4BEG[5] ,
    \Tile_X8Y12_NN4BEG[4] ,
    \Tile_X8Y12_NN4BEG[3] ,
    \Tile_X8Y12_NN4BEG[2] ,
    \Tile_X8Y12_NN4BEG[1] ,
    \Tile_X8Y12_NN4BEG[0] }),
    .S1BEG({\Tile_X8Y11_S1BEG[3] ,
    \Tile_X8Y11_S1BEG[2] ,
    \Tile_X8Y11_S1BEG[1] ,
    \Tile_X8Y11_S1BEG[0] }),
    .S1END({\Tile_X8Y10_S1BEG[3] ,
    \Tile_X8Y10_S1BEG[2] ,
    \Tile_X8Y10_S1BEG[1] ,
    \Tile_X8Y10_S1BEG[0] }),
    .S2BEG({\Tile_X8Y11_S2BEG[7] ,
    \Tile_X8Y11_S2BEG[6] ,
    \Tile_X8Y11_S2BEG[5] ,
    \Tile_X8Y11_S2BEG[4] ,
    \Tile_X8Y11_S2BEG[3] ,
    \Tile_X8Y11_S2BEG[2] ,
    \Tile_X8Y11_S2BEG[1] ,
    \Tile_X8Y11_S2BEG[0] }),
    .S2BEGb({\Tile_X8Y11_S2BEGb[7] ,
    \Tile_X8Y11_S2BEGb[6] ,
    \Tile_X8Y11_S2BEGb[5] ,
    \Tile_X8Y11_S2BEGb[4] ,
    \Tile_X8Y11_S2BEGb[3] ,
    \Tile_X8Y11_S2BEGb[2] ,
    \Tile_X8Y11_S2BEGb[1] ,
    \Tile_X8Y11_S2BEGb[0] }),
    .S2END({\Tile_X8Y10_S2BEGb[7] ,
    \Tile_X8Y10_S2BEGb[6] ,
    \Tile_X8Y10_S2BEGb[5] ,
    \Tile_X8Y10_S2BEGb[4] ,
    \Tile_X8Y10_S2BEGb[3] ,
    \Tile_X8Y10_S2BEGb[2] ,
    \Tile_X8Y10_S2BEGb[1] ,
    \Tile_X8Y10_S2BEGb[0] }),
    .S2MID({\Tile_X8Y10_S2BEG[7] ,
    \Tile_X8Y10_S2BEG[6] ,
    \Tile_X8Y10_S2BEG[5] ,
    \Tile_X8Y10_S2BEG[4] ,
    \Tile_X8Y10_S2BEG[3] ,
    \Tile_X8Y10_S2BEG[2] ,
    \Tile_X8Y10_S2BEG[1] ,
    \Tile_X8Y10_S2BEG[0] }),
    .S4BEG({\Tile_X8Y11_S4BEG[15] ,
    \Tile_X8Y11_S4BEG[14] ,
    \Tile_X8Y11_S4BEG[13] ,
    \Tile_X8Y11_S4BEG[12] ,
    \Tile_X8Y11_S4BEG[11] ,
    \Tile_X8Y11_S4BEG[10] ,
    \Tile_X8Y11_S4BEG[9] ,
    \Tile_X8Y11_S4BEG[8] ,
    \Tile_X8Y11_S4BEG[7] ,
    \Tile_X8Y11_S4BEG[6] ,
    \Tile_X8Y11_S4BEG[5] ,
    \Tile_X8Y11_S4BEG[4] ,
    \Tile_X8Y11_S4BEG[3] ,
    \Tile_X8Y11_S4BEG[2] ,
    \Tile_X8Y11_S4BEG[1] ,
    \Tile_X8Y11_S4BEG[0] }),
    .S4END({\Tile_X8Y10_S4BEG[15] ,
    \Tile_X8Y10_S4BEG[14] ,
    \Tile_X8Y10_S4BEG[13] ,
    \Tile_X8Y10_S4BEG[12] ,
    \Tile_X8Y10_S4BEG[11] ,
    \Tile_X8Y10_S4BEG[10] ,
    \Tile_X8Y10_S4BEG[9] ,
    \Tile_X8Y10_S4BEG[8] ,
    \Tile_X8Y10_S4BEG[7] ,
    \Tile_X8Y10_S4BEG[6] ,
    \Tile_X8Y10_S4BEG[5] ,
    \Tile_X8Y10_S4BEG[4] ,
    \Tile_X8Y10_S4BEG[3] ,
    \Tile_X8Y10_S4BEG[2] ,
    \Tile_X8Y10_S4BEG[1] ,
    \Tile_X8Y10_S4BEG[0] }),
    .SS4BEG({\Tile_X8Y11_SS4BEG[15] ,
    \Tile_X8Y11_SS4BEG[14] ,
    \Tile_X8Y11_SS4BEG[13] ,
    \Tile_X8Y11_SS4BEG[12] ,
    \Tile_X8Y11_SS4BEG[11] ,
    \Tile_X8Y11_SS4BEG[10] ,
    \Tile_X8Y11_SS4BEG[9] ,
    \Tile_X8Y11_SS4BEG[8] ,
    \Tile_X8Y11_SS4BEG[7] ,
    \Tile_X8Y11_SS4BEG[6] ,
    \Tile_X8Y11_SS4BEG[5] ,
    \Tile_X8Y11_SS4BEG[4] ,
    \Tile_X8Y11_SS4BEG[3] ,
    \Tile_X8Y11_SS4BEG[2] ,
    \Tile_X8Y11_SS4BEG[1] ,
    \Tile_X8Y11_SS4BEG[0] }),
    .SS4END({\Tile_X8Y10_SS4BEG[15] ,
    \Tile_X8Y10_SS4BEG[14] ,
    \Tile_X8Y10_SS4BEG[13] ,
    \Tile_X8Y10_SS4BEG[12] ,
    \Tile_X8Y10_SS4BEG[11] ,
    \Tile_X8Y10_SS4BEG[10] ,
    \Tile_X8Y10_SS4BEG[9] ,
    \Tile_X8Y10_SS4BEG[8] ,
    \Tile_X8Y10_SS4BEG[7] ,
    \Tile_X8Y10_SS4BEG[6] ,
    \Tile_X8Y10_SS4BEG[5] ,
    \Tile_X8Y10_SS4BEG[4] ,
    \Tile_X8Y10_SS4BEG[3] ,
    \Tile_X8Y10_SS4BEG[2] ,
    \Tile_X8Y10_SS4BEG[1] ,
    \Tile_X8Y10_SS4BEG[0] }),
    .W1BEG({\Tile_X8Y11_W1BEG[3] ,
    \Tile_X8Y11_W1BEG[2] ,
    \Tile_X8Y11_W1BEG[1] ,
    \Tile_X8Y11_W1BEG[0] }),
    .W1END({\Tile_X9Y11_W1BEG[3] ,
    \Tile_X9Y11_W1BEG[2] ,
    \Tile_X9Y11_W1BEG[1] ,
    \Tile_X9Y11_W1BEG[0] }),
    .W2BEG({\Tile_X8Y11_W2BEG[7] ,
    \Tile_X8Y11_W2BEG[6] ,
    \Tile_X8Y11_W2BEG[5] ,
    \Tile_X8Y11_W2BEG[4] ,
    \Tile_X8Y11_W2BEG[3] ,
    \Tile_X8Y11_W2BEG[2] ,
    \Tile_X8Y11_W2BEG[1] ,
    \Tile_X8Y11_W2BEG[0] }),
    .W2BEGb({\Tile_X8Y11_W2BEGb[7] ,
    \Tile_X8Y11_W2BEGb[6] ,
    \Tile_X8Y11_W2BEGb[5] ,
    \Tile_X8Y11_W2BEGb[4] ,
    \Tile_X8Y11_W2BEGb[3] ,
    \Tile_X8Y11_W2BEGb[2] ,
    \Tile_X8Y11_W2BEGb[1] ,
    \Tile_X8Y11_W2BEGb[0] }),
    .W2END({\Tile_X9Y11_W2BEGb[7] ,
    \Tile_X9Y11_W2BEGb[6] ,
    \Tile_X9Y11_W2BEGb[5] ,
    \Tile_X9Y11_W2BEGb[4] ,
    \Tile_X9Y11_W2BEGb[3] ,
    \Tile_X9Y11_W2BEGb[2] ,
    \Tile_X9Y11_W2BEGb[1] ,
    \Tile_X9Y11_W2BEGb[0] }),
    .W2MID({\Tile_X9Y11_W2BEG[7] ,
    \Tile_X9Y11_W2BEG[6] ,
    \Tile_X9Y11_W2BEG[5] ,
    \Tile_X9Y11_W2BEG[4] ,
    \Tile_X9Y11_W2BEG[3] ,
    \Tile_X9Y11_W2BEG[2] ,
    \Tile_X9Y11_W2BEG[1] ,
    \Tile_X9Y11_W2BEG[0] }),
    .W6BEG({\Tile_X8Y11_W6BEG[11] ,
    \Tile_X8Y11_W6BEG[10] ,
    \Tile_X8Y11_W6BEG[9] ,
    \Tile_X8Y11_W6BEG[8] ,
    \Tile_X8Y11_W6BEG[7] ,
    \Tile_X8Y11_W6BEG[6] ,
    \Tile_X8Y11_W6BEG[5] ,
    \Tile_X8Y11_W6BEG[4] ,
    \Tile_X8Y11_W6BEG[3] ,
    \Tile_X8Y11_W6BEG[2] ,
    \Tile_X8Y11_W6BEG[1] ,
    \Tile_X8Y11_W6BEG[0] }),
    .W6END({\Tile_X9Y11_W6BEG[11] ,
    \Tile_X9Y11_W6BEG[10] ,
    \Tile_X9Y11_W6BEG[9] ,
    \Tile_X9Y11_W6BEG[8] ,
    \Tile_X9Y11_W6BEG[7] ,
    \Tile_X9Y11_W6BEG[6] ,
    \Tile_X9Y11_W6BEG[5] ,
    \Tile_X9Y11_W6BEG[4] ,
    \Tile_X9Y11_W6BEG[3] ,
    \Tile_X9Y11_W6BEG[2] ,
    \Tile_X9Y11_W6BEG[1] ,
    \Tile_X9Y11_W6BEG[0] }),
    .WW4BEG({\Tile_X8Y11_WW4BEG[15] ,
    \Tile_X8Y11_WW4BEG[14] ,
    \Tile_X8Y11_WW4BEG[13] ,
    \Tile_X8Y11_WW4BEG[12] ,
    \Tile_X8Y11_WW4BEG[11] ,
    \Tile_X8Y11_WW4BEG[10] ,
    \Tile_X8Y11_WW4BEG[9] ,
    \Tile_X8Y11_WW4BEG[8] ,
    \Tile_X8Y11_WW4BEG[7] ,
    \Tile_X8Y11_WW4BEG[6] ,
    \Tile_X8Y11_WW4BEG[5] ,
    \Tile_X8Y11_WW4BEG[4] ,
    \Tile_X8Y11_WW4BEG[3] ,
    \Tile_X8Y11_WW4BEG[2] ,
    \Tile_X8Y11_WW4BEG[1] ,
    \Tile_X8Y11_WW4BEG[0] }),
    .WW4END({\Tile_X9Y11_WW4BEG[15] ,
    \Tile_X9Y11_WW4BEG[14] ,
    \Tile_X9Y11_WW4BEG[13] ,
    \Tile_X9Y11_WW4BEG[12] ,
    \Tile_X9Y11_WW4BEG[11] ,
    \Tile_X9Y11_WW4BEG[10] ,
    \Tile_X9Y11_WW4BEG[9] ,
    \Tile_X9Y11_WW4BEG[8] ,
    \Tile_X9Y11_WW4BEG[7] ,
    \Tile_X9Y11_WW4BEG[6] ,
    \Tile_X9Y11_WW4BEG[5] ,
    \Tile_X9Y11_WW4BEG[4] ,
    \Tile_X9Y11_WW4BEG[3] ,
    \Tile_X9Y11_WW4BEG[2] ,
    \Tile_X9Y11_WW4BEG[1] ,
    \Tile_X9Y11_WW4BEG[0] }));
 LUT4AB Tile_X8Y12_LUT4AB (.Ci(Tile_X8Y13_Co),
    .Co(Tile_X8Y12_Co),
    .UserCLK(Tile_X8Y13_UserCLKo),
    .UserCLKo(Tile_X8Y12_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X8Y12_E1BEG[3] ,
    \Tile_X8Y12_E1BEG[2] ,
    \Tile_X8Y12_E1BEG[1] ,
    \Tile_X8Y12_E1BEG[0] }),
    .E1END({\Tile_X7Y12_E1BEG[3] ,
    \Tile_X7Y12_E1BEG[2] ,
    \Tile_X7Y12_E1BEG[1] ,
    \Tile_X7Y12_E1BEG[0] }),
    .E2BEG({\Tile_X8Y12_E2BEG[7] ,
    \Tile_X8Y12_E2BEG[6] ,
    \Tile_X8Y12_E2BEG[5] ,
    \Tile_X8Y12_E2BEG[4] ,
    \Tile_X8Y12_E2BEG[3] ,
    \Tile_X8Y12_E2BEG[2] ,
    \Tile_X8Y12_E2BEG[1] ,
    \Tile_X8Y12_E2BEG[0] }),
    .E2BEGb({\Tile_X8Y12_E2BEGb[7] ,
    \Tile_X8Y12_E2BEGb[6] ,
    \Tile_X8Y12_E2BEGb[5] ,
    \Tile_X8Y12_E2BEGb[4] ,
    \Tile_X8Y12_E2BEGb[3] ,
    \Tile_X8Y12_E2BEGb[2] ,
    \Tile_X8Y12_E2BEGb[1] ,
    \Tile_X8Y12_E2BEGb[0] }),
    .E2END({\Tile_X7Y12_E2BEGb[7] ,
    \Tile_X7Y12_E2BEGb[6] ,
    \Tile_X7Y12_E2BEGb[5] ,
    \Tile_X7Y12_E2BEGb[4] ,
    \Tile_X7Y12_E2BEGb[3] ,
    \Tile_X7Y12_E2BEGb[2] ,
    \Tile_X7Y12_E2BEGb[1] ,
    \Tile_X7Y12_E2BEGb[0] }),
    .E2MID({\Tile_X7Y12_E2BEG[7] ,
    \Tile_X7Y12_E2BEG[6] ,
    \Tile_X7Y12_E2BEG[5] ,
    \Tile_X7Y12_E2BEG[4] ,
    \Tile_X7Y12_E2BEG[3] ,
    \Tile_X7Y12_E2BEG[2] ,
    \Tile_X7Y12_E2BEG[1] ,
    \Tile_X7Y12_E2BEG[0] }),
    .E6BEG({\Tile_X8Y12_E6BEG[11] ,
    \Tile_X8Y12_E6BEG[10] ,
    \Tile_X8Y12_E6BEG[9] ,
    \Tile_X8Y12_E6BEG[8] ,
    \Tile_X8Y12_E6BEG[7] ,
    \Tile_X8Y12_E6BEG[6] ,
    \Tile_X8Y12_E6BEG[5] ,
    \Tile_X8Y12_E6BEG[4] ,
    \Tile_X8Y12_E6BEG[3] ,
    \Tile_X8Y12_E6BEG[2] ,
    \Tile_X8Y12_E6BEG[1] ,
    \Tile_X8Y12_E6BEG[0] }),
    .E6END({\Tile_X7Y12_E6BEG[11] ,
    \Tile_X7Y12_E6BEG[10] ,
    \Tile_X7Y12_E6BEG[9] ,
    \Tile_X7Y12_E6BEG[8] ,
    \Tile_X7Y12_E6BEG[7] ,
    \Tile_X7Y12_E6BEG[6] ,
    \Tile_X7Y12_E6BEG[5] ,
    \Tile_X7Y12_E6BEG[4] ,
    \Tile_X7Y12_E6BEG[3] ,
    \Tile_X7Y12_E6BEG[2] ,
    \Tile_X7Y12_E6BEG[1] ,
    \Tile_X7Y12_E6BEG[0] }),
    .EE4BEG({\Tile_X8Y12_EE4BEG[15] ,
    \Tile_X8Y12_EE4BEG[14] ,
    \Tile_X8Y12_EE4BEG[13] ,
    \Tile_X8Y12_EE4BEG[12] ,
    \Tile_X8Y12_EE4BEG[11] ,
    \Tile_X8Y12_EE4BEG[10] ,
    \Tile_X8Y12_EE4BEG[9] ,
    \Tile_X8Y12_EE4BEG[8] ,
    \Tile_X8Y12_EE4BEG[7] ,
    \Tile_X8Y12_EE4BEG[6] ,
    \Tile_X8Y12_EE4BEG[5] ,
    \Tile_X8Y12_EE4BEG[4] ,
    \Tile_X8Y12_EE4BEG[3] ,
    \Tile_X8Y12_EE4BEG[2] ,
    \Tile_X8Y12_EE4BEG[1] ,
    \Tile_X8Y12_EE4BEG[0] }),
    .EE4END({\Tile_X7Y12_EE4BEG[15] ,
    \Tile_X7Y12_EE4BEG[14] ,
    \Tile_X7Y12_EE4BEG[13] ,
    \Tile_X7Y12_EE4BEG[12] ,
    \Tile_X7Y12_EE4BEG[11] ,
    \Tile_X7Y12_EE4BEG[10] ,
    \Tile_X7Y12_EE4BEG[9] ,
    \Tile_X7Y12_EE4BEG[8] ,
    \Tile_X7Y12_EE4BEG[7] ,
    \Tile_X7Y12_EE4BEG[6] ,
    \Tile_X7Y12_EE4BEG[5] ,
    \Tile_X7Y12_EE4BEG[4] ,
    \Tile_X7Y12_EE4BEG[3] ,
    \Tile_X7Y12_EE4BEG[2] ,
    \Tile_X7Y12_EE4BEG[1] ,
    \Tile_X7Y12_EE4BEG[0] }),
    .FrameData({\Tile_X7Y12_FrameData_O[31] ,
    \Tile_X7Y12_FrameData_O[30] ,
    \Tile_X7Y12_FrameData_O[29] ,
    \Tile_X7Y12_FrameData_O[28] ,
    \Tile_X7Y12_FrameData_O[27] ,
    \Tile_X7Y12_FrameData_O[26] ,
    \Tile_X7Y12_FrameData_O[25] ,
    \Tile_X7Y12_FrameData_O[24] ,
    \Tile_X7Y12_FrameData_O[23] ,
    \Tile_X7Y12_FrameData_O[22] ,
    \Tile_X7Y12_FrameData_O[21] ,
    \Tile_X7Y12_FrameData_O[20] ,
    \Tile_X7Y12_FrameData_O[19] ,
    \Tile_X7Y12_FrameData_O[18] ,
    \Tile_X7Y12_FrameData_O[17] ,
    \Tile_X7Y12_FrameData_O[16] ,
    \Tile_X7Y12_FrameData_O[15] ,
    \Tile_X7Y12_FrameData_O[14] ,
    \Tile_X7Y12_FrameData_O[13] ,
    \Tile_X7Y12_FrameData_O[12] ,
    \Tile_X7Y12_FrameData_O[11] ,
    \Tile_X7Y12_FrameData_O[10] ,
    \Tile_X7Y12_FrameData_O[9] ,
    \Tile_X7Y12_FrameData_O[8] ,
    \Tile_X7Y12_FrameData_O[7] ,
    \Tile_X7Y12_FrameData_O[6] ,
    \Tile_X7Y12_FrameData_O[5] ,
    \Tile_X7Y12_FrameData_O[4] ,
    \Tile_X7Y12_FrameData_O[3] ,
    \Tile_X7Y12_FrameData_O[2] ,
    \Tile_X7Y12_FrameData_O[1] ,
    \Tile_X7Y12_FrameData_O[0] }),
    .FrameData_O({\Tile_X8Y12_FrameData_O[31] ,
    \Tile_X8Y12_FrameData_O[30] ,
    \Tile_X8Y12_FrameData_O[29] ,
    \Tile_X8Y12_FrameData_O[28] ,
    \Tile_X8Y12_FrameData_O[27] ,
    \Tile_X8Y12_FrameData_O[26] ,
    \Tile_X8Y12_FrameData_O[25] ,
    \Tile_X8Y12_FrameData_O[24] ,
    \Tile_X8Y12_FrameData_O[23] ,
    \Tile_X8Y12_FrameData_O[22] ,
    \Tile_X8Y12_FrameData_O[21] ,
    \Tile_X8Y12_FrameData_O[20] ,
    \Tile_X8Y12_FrameData_O[19] ,
    \Tile_X8Y12_FrameData_O[18] ,
    \Tile_X8Y12_FrameData_O[17] ,
    \Tile_X8Y12_FrameData_O[16] ,
    \Tile_X8Y12_FrameData_O[15] ,
    \Tile_X8Y12_FrameData_O[14] ,
    \Tile_X8Y12_FrameData_O[13] ,
    \Tile_X8Y12_FrameData_O[12] ,
    \Tile_X8Y12_FrameData_O[11] ,
    \Tile_X8Y12_FrameData_O[10] ,
    \Tile_X8Y12_FrameData_O[9] ,
    \Tile_X8Y12_FrameData_O[8] ,
    \Tile_X8Y12_FrameData_O[7] ,
    \Tile_X8Y12_FrameData_O[6] ,
    \Tile_X8Y12_FrameData_O[5] ,
    \Tile_X8Y12_FrameData_O[4] ,
    \Tile_X8Y12_FrameData_O[3] ,
    \Tile_X8Y12_FrameData_O[2] ,
    \Tile_X8Y12_FrameData_O[1] ,
    \Tile_X8Y12_FrameData_O[0] }),
    .FrameStrobe({\Tile_X8Y13_FrameStrobe_O[19] ,
    \Tile_X8Y13_FrameStrobe_O[18] ,
    \Tile_X8Y13_FrameStrobe_O[17] ,
    \Tile_X8Y13_FrameStrobe_O[16] ,
    \Tile_X8Y13_FrameStrobe_O[15] ,
    \Tile_X8Y13_FrameStrobe_O[14] ,
    \Tile_X8Y13_FrameStrobe_O[13] ,
    \Tile_X8Y13_FrameStrobe_O[12] ,
    \Tile_X8Y13_FrameStrobe_O[11] ,
    \Tile_X8Y13_FrameStrobe_O[10] ,
    \Tile_X8Y13_FrameStrobe_O[9] ,
    \Tile_X8Y13_FrameStrobe_O[8] ,
    \Tile_X8Y13_FrameStrobe_O[7] ,
    \Tile_X8Y13_FrameStrobe_O[6] ,
    \Tile_X8Y13_FrameStrobe_O[5] ,
    \Tile_X8Y13_FrameStrobe_O[4] ,
    \Tile_X8Y13_FrameStrobe_O[3] ,
    \Tile_X8Y13_FrameStrobe_O[2] ,
    \Tile_X8Y13_FrameStrobe_O[1] ,
    \Tile_X8Y13_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X8Y12_FrameStrobe_O[19] ,
    \Tile_X8Y12_FrameStrobe_O[18] ,
    \Tile_X8Y12_FrameStrobe_O[17] ,
    \Tile_X8Y12_FrameStrobe_O[16] ,
    \Tile_X8Y12_FrameStrobe_O[15] ,
    \Tile_X8Y12_FrameStrobe_O[14] ,
    \Tile_X8Y12_FrameStrobe_O[13] ,
    \Tile_X8Y12_FrameStrobe_O[12] ,
    \Tile_X8Y12_FrameStrobe_O[11] ,
    \Tile_X8Y12_FrameStrobe_O[10] ,
    \Tile_X8Y12_FrameStrobe_O[9] ,
    \Tile_X8Y12_FrameStrobe_O[8] ,
    \Tile_X8Y12_FrameStrobe_O[7] ,
    \Tile_X8Y12_FrameStrobe_O[6] ,
    \Tile_X8Y12_FrameStrobe_O[5] ,
    \Tile_X8Y12_FrameStrobe_O[4] ,
    \Tile_X8Y12_FrameStrobe_O[3] ,
    \Tile_X8Y12_FrameStrobe_O[2] ,
    \Tile_X8Y12_FrameStrobe_O[1] ,
    \Tile_X8Y12_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X8Y12_N1BEG[3] ,
    \Tile_X8Y12_N1BEG[2] ,
    \Tile_X8Y12_N1BEG[1] ,
    \Tile_X8Y12_N1BEG[0] }),
    .N1END({\Tile_X8Y13_N1BEG[3] ,
    \Tile_X8Y13_N1BEG[2] ,
    \Tile_X8Y13_N1BEG[1] ,
    \Tile_X8Y13_N1BEG[0] }),
    .N2BEG({\Tile_X8Y12_N2BEG[7] ,
    \Tile_X8Y12_N2BEG[6] ,
    \Tile_X8Y12_N2BEG[5] ,
    \Tile_X8Y12_N2BEG[4] ,
    \Tile_X8Y12_N2BEG[3] ,
    \Tile_X8Y12_N2BEG[2] ,
    \Tile_X8Y12_N2BEG[1] ,
    \Tile_X8Y12_N2BEG[0] }),
    .N2BEGb({\Tile_X8Y12_N2BEGb[7] ,
    \Tile_X8Y12_N2BEGb[6] ,
    \Tile_X8Y12_N2BEGb[5] ,
    \Tile_X8Y12_N2BEGb[4] ,
    \Tile_X8Y12_N2BEGb[3] ,
    \Tile_X8Y12_N2BEGb[2] ,
    \Tile_X8Y12_N2BEGb[1] ,
    \Tile_X8Y12_N2BEGb[0] }),
    .N2END({\Tile_X8Y13_N2BEGb[7] ,
    \Tile_X8Y13_N2BEGb[6] ,
    \Tile_X8Y13_N2BEGb[5] ,
    \Tile_X8Y13_N2BEGb[4] ,
    \Tile_X8Y13_N2BEGb[3] ,
    \Tile_X8Y13_N2BEGb[2] ,
    \Tile_X8Y13_N2BEGb[1] ,
    \Tile_X8Y13_N2BEGb[0] }),
    .N2MID({\Tile_X8Y13_N2BEG[7] ,
    \Tile_X8Y13_N2BEG[6] ,
    \Tile_X8Y13_N2BEG[5] ,
    \Tile_X8Y13_N2BEG[4] ,
    \Tile_X8Y13_N2BEG[3] ,
    \Tile_X8Y13_N2BEG[2] ,
    \Tile_X8Y13_N2BEG[1] ,
    \Tile_X8Y13_N2BEG[0] }),
    .N4BEG({\Tile_X8Y12_N4BEG[15] ,
    \Tile_X8Y12_N4BEG[14] ,
    \Tile_X8Y12_N4BEG[13] ,
    \Tile_X8Y12_N4BEG[12] ,
    \Tile_X8Y12_N4BEG[11] ,
    \Tile_X8Y12_N4BEG[10] ,
    \Tile_X8Y12_N4BEG[9] ,
    \Tile_X8Y12_N4BEG[8] ,
    \Tile_X8Y12_N4BEG[7] ,
    \Tile_X8Y12_N4BEG[6] ,
    \Tile_X8Y12_N4BEG[5] ,
    \Tile_X8Y12_N4BEG[4] ,
    \Tile_X8Y12_N4BEG[3] ,
    \Tile_X8Y12_N4BEG[2] ,
    \Tile_X8Y12_N4BEG[1] ,
    \Tile_X8Y12_N4BEG[0] }),
    .N4END({\Tile_X8Y13_N4BEG[15] ,
    \Tile_X8Y13_N4BEG[14] ,
    \Tile_X8Y13_N4BEG[13] ,
    \Tile_X8Y13_N4BEG[12] ,
    \Tile_X8Y13_N4BEG[11] ,
    \Tile_X8Y13_N4BEG[10] ,
    \Tile_X8Y13_N4BEG[9] ,
    \Tile_X8Y13_N4BEG[8] ,
    \Tile_X8Y13_N4BEG[7] ,
    \Tile_X8Y13_N4BEG[6] ,
    \Tile_X8Y13_N4BEG[5] ,
    \Tile_X8Y13_N4BEG[4] ,
    \Tile_X8Y13_N4BEG[3] ,
    \Tile_X8Y13_N4BEG[2] ,
    \Tile_X8Y13_N4BEG[1] ,
    \Tile_X8Y13_N4BEG[0] }),
    .NN4BEG({\Tile_X8Y12_NN4BEG[15] ,
    \Tile_X8Y12_NN4BEG[14] ,
    \Tile_X8Y12_NN4BEG[13] ,
    \Tile_X8Y12_NN4BEG[12] ,
    \Tile_X8Y12_NN4BEG[11] ,
    \Tile_X8Y12_NN4BEG[10] ,
    \Tile_X8Y12_NN4BEG[9] ,
    \Tile_X8Y12_NN4BEG[8] ,
    \Tile_X8Y12_NN4BEG[7] ,
    \Tile_X8Y12_NN4BEG[6] ,
    \Tile_X8Y12_NN4BEG[5] ,
    \Tile_X8Y12_NN4BEG[4] ,
    \Tile_X8Y12_NN4BEG[3] ,
    \Tile_X8Y12_NN4BEG[2] ,
    \Tile_X8Y12_NN4BEG[1] ,
    \Tile_X8Y12_NN4BEG[0] }),
    .NN4END({\Tile_X8Y13_NN4BEG[15] ,
    \Tile_X8Y13_NN4BEG[14] ,
    \Tile_X8Y13_NN4BEG[13] ,
    \Tile_X8Y13_NN4BEG[12] ,
    \Tile_X8Y13_NN4BEG[11] ,
    \Tile_X8Y13_NN4BEG[10] ,
    \Tile_X8Y13_NN4BEG[9] ,
    \Tile_X8Y13_NN4BEG[8] ,
    \Tile_X8Y13_NN4BEG[7] ,
    \Tile_X8Y13_NN4BEG[6] ,
    \Tile_X8Y13_NN4BEG[5] ,
    \Tile_X8Y13_NN4BEG[4] ,
    \Tile_X8Y13_NN4BEG[3] ,
    \Tile_X8Y13_NN4BEG[2] ,
    \Tile_X8Y13_NN4BEG[1] ,
    \Tile_X8Y13_NN4BEG[0] }),
    .S1BEG({\Tile_X8Y12_S1BEG[3] ,
    \Tile_X8Y12_S1BEG[2] ,
    \Tile_X8Y12_S1BEG[1] ,
    \Tile_X8Y12_S1BEG[0] }),
    .S1END({\Tile_X8Y11_S1BEG[3] ,
    \Tile_X8Y11_S1BEG[2] ,
    \Tile_X8Y11_S1BEG[1] ,
    \Tile_X8Y11_S1BEG[0] }),
    .S2BEG({\Tile_X8Y12_S2BEG[7] ,
    \Tile_X8Y12_S2BEG[6] ,
    \Tile_X8Y12_S2BEG[5] ,
    \Tile_X8Y12_S2BEG[4] ,
    \Tile_X8Y12_S2BEG[3] ,
    \Tile_X8Y12_S2BEG[2] ,
    \Tile_X8Y12_S2BEG[1] ,
    \Tile_X8Y12_S2BEG[0] }),
    .S2BEGb({\Tile_X8Y12_S2BEGb[7] ,
    \Tile_X8Y12_S2BEGb[6] ,
    \Tile_X8Y12_S2BEGb[5] ,
    \Tile_X8Y12_S2BEGb[4] ,
    \Tile_X8Y12_S2BEGb[3] ,
    \Tile_X8Y12_S2BEGb[2] ,
    \Tile_X8Y12_S2BEGb[1] ,
    \Tile_X8Y12_S2BEGb[0] }),
    .S2END({\Tile_X8Y11_S2BEGb[7] ,
    \Tile_X8Y11_S2BEGb[6] ,
    \Tile_X8Y11_S2BEGb[5] ,
    \Tile_X8Y11_S2BEGb[4] ,
    \Tile_X8Y11_S2BEGb[3] ,
    \Tile_X8Y11_S2BEGb[2] ,
    \Tile_X8Y11_S2BEGb[1] ,
    \Tile_X8Y11_S2BEGb[0] }),
    .S2MID({\Tile_X8Y11_S2BEG[7] ,
    \Tile_X8Y11_S2BEG[6] ,
    \Tile_X8Y11_S2BEG[5] ,
    \Tile_X8Y11_S2BEG[4] ,
    \Tile_X8Y11_S2BEG[3] ,
    \Tile_X8Y11_S2BEG[2] ,
    \Tile_X8Y11_S2BEG[1] ,
    \Tile_X8Y11_S2BEG[0] }),
    .S4BEG({\Tile_X8Y12_S4BEG[15] ,
    \Tile_X8Y12_S4BEG[14] ,
    \Tile_X8Y12_S4BEG[13] ,
    \Tile_X8Y12_S4BEG[12] ,
    \Tile_X8Y12_S4BEG[11] ,
    \Tile_X8Y12_S4BEG[10] ,
    \Tile_X8Y12_S4BEG[9] ,
    \Tile_X8Y12_S4BEG[8] ,
    \Tile_X8Y12_S4BEG[7] ,
    \Tile_X8Y12_S4BEG[6] ,
    \Tile_X8Y12_S4BEG[5] ,
    \Tile_X8Y12_S4BEG[4] ,
    \Tile_X8Y12_S4BEG[3] ,
    \Tile_X8Y12_S4BEG[2] ,
    \Tile_X8Y12_S4BEG[1] ,
    \Tile_X8Y12_S4BEG[0] }),
    .S4END({\Tile_X8Y11_S4BEG[15] ,
    \Tile_X8Y11_S4BEG[14] ,
    \Tile_X8Y11_S4BEG[13] ,
    \Tile_X8Y11_S4BEG[12] ,
    \Tile_X8Y11_S4BEG[11] ,
    \Tile_X8Y11_S4BEG[10] ,
    \Tile_X8Y11_S4BEG[9] ,
    \Tile_X8Y11_S4BEG[8] ,
    \Tile_X8Y11_S4BEG[7] ,
    \Tile_X8Y11_S4BEG[6] ,
    \Tile_X8Y11_S4BEG[5] ,
    \Tile_X8Y11_S4BEG[4] ,
    \Tile_X8Y11_S4BEG[3] ,
    \Tile_X8Y11_S4BEG[2] ,
    \Tile_X8Y11_S4BEG[1] ,
    \Tile_X8Y11_S4BEG[0] }),
    .SS4BEG({\Tile_X8Y12_SS4BEG[15] ,
    \Tile_X8Y12_SS4BEG[14] ,
    \Tile_X8Y12_SS4BEG[13] ,
    \Tile_X8Y12_SS4BEG[12] ,
    \Tile_X8Y12_SS4BEG[11] ,
    \Tile_X8Y12_SS4BEG[10] ,
    \Tile_X8Y12_SS4BEG[9] ,
    \Tile_X8Y12_SS4BEG[8] ,
    \Tile_X8Y12_SS4BEG[7] ,
    \Tile_X8Y12_SS4BEG[6] ,
    \Tile_X8Y12_SS4BEG[5] ,
    \Tile_X8Y12_SS4BEG[4] ,
    \Tile_X8Y12_SS4BEG[3] ,
    \Tile_X8Y12_SS4BEG[2] ,
    \Tile_X8Y12_SS4BEG[1] ,
    \Tile_X8Y12_SS4BEG[0] }),
    .SS4END({\Tile_X8Y11_SS4BEG[15] ,
    \Tile_X8Y11_SS4BEG[14] ,
    \Tile_X8Y11_SS4BEG[13] ,
    \Tile_X8Y11_SS4BEG[12] ,
    \Tile_X8Y11_SS4BEG[11] ,
    \Tile_X8Y11_SS4BEG[10] ,
    \Tile_X8Y11_SS4BEG[9] ,
    \Tile_X8Y11_SS4BEG[8] ,
    \Tile_X8Y11_SS4BEG[7] ,
    \Tile_X8Y11_SS4BEG[6] ,
    \Tile_X8Y11_SS4BEG[5] ,
    \Tile_X8Y11_SS4BEG[4] ,
    \Tile_X8Y11_SS4BEG[3] ,
    \Tile_X8Y11_SS4BEG[2] ,
    \Tile_X8Y11_SS4BEG[1] ,
    \Tile_X8Y11_SS4BEG[0] }),
    .W1BEG({\Tile_X8Y12_W1BEG[3] ,
    \Tile_X8Y12_W1BEG[2] ,
    \Tile_X8Y12_W1BEG[1] ,
    \Tile_X8Y12_W1BEG[0] }),
    .W1END({\Tile_X9Y12_W1BEG[3] ,
    \Tile_X9Y12_W1BEG[2] ,
    \Tile_X9Y12_W1BEG[1] ,
    \Tile_X9Y12_W1BEG[0] }),
    .W2BEG({\Tile_X8Y12_W2BEG[7] ,
    \Tile_X8Y12_W2BEG[6] ,
    \Tile_X8Y12_W2BEG[5] ,
    \Tile_X8Y12_W2BEG[4] ,
    \Tile_X8Y12_W2BEG[3] ,
    \Tile_X8Y12_W2BEG[2] ,
    \Tile_X8Y12_W2BEG[1] ,
    \Tile_X8Y12_W2BEG[0] }),
    .W2BEGb({\Tile_X8Y12_W2BEGb[7] ,
    \Tile_X8Y12_W2BEGb[6] ,
    \Tile_X8Y12_W2BEGb[5] ,
    \Tile_X8Y12_W2BEGb[4] ,
    \Tile_X8Y12_W2BEGb[3] ,
    \Tile_X8Y12_W2BEGb[2] ,
    \Tile_X8Y12_W2BEGb[1] ,
    \Tile_X8Y12_W2BEGb[0] }),
    .W2END({\Tile_X9Y12_W2BEGb[7] ,
    \Tile_X9Y12_W2BEGb[6] ,
    \Tile_X9Y12_W2BEGb[5] ,
    \Tile_X9Y12_W2BEGb[4] ,
    \Tile_X9Y12_W2BEGb[3] ,
    \Tile_X9Y12_W2BEGb[2] ,
    \Tile_X9Y12_W2BEGb[1] ,
    \Tile_X9Y12_W2BEGb[0] }),
    .W2MID({\Tile_X9Y12_W2BEG[7] ,
    \Tile_X9Y12_W2BEG[6] ,
    \Tile_X9Y12_W2BEG[5] ,
    \Tile_X9Y12_W2BEG[4] ,
    \Tile_X9Y12_W2BEG[3] ,
    \Tile_X9Y12_W2BEG[2] ,
    \Tile_X9Y12_W2BEG[1] ,
    \Tile_X9Y12_W2BEG[0] }),
    .W6BEG({\Tile_X8Y12_W6BEG[11] ,
    \Tile_X8Y12_W6BEG[10] ,
    \Tile_X8Y12_W6BEG[9] ,
    \Tile_X8Y12_W6BEG[8] ,
    \Tile_X8Y12_W6BEG[7] ,
    \Tile_X8Y12_W6BEG[6] ,
    \Tile_X8Y12_W6BEG[5] ,
    \Tile_X8Y12_W6BEG[4] ,
    \Tile_X8Y12_W6BEG[3] ,
    \Tile_X8Y12_W6BEG[2] ,
    \Tile_X8Y12_W6BEG[1] ,
    \Tile_X8Y12_W6BEG[0] }),
    .W6END({\Tile_X9Y12_W6BEG[11] ,
    \Tile_X9Y12_W6BEG[10] ,
    \Tile_X9Y12_W6BEG[9] ,
    \Tile_X9Y12_W6BEG[8] ,
    \Tile_X9Y12_W6BEG[7] ,
    \Tile_X9Y12_W6BEG[6] ,
    \Tile_X9Y12_W6BEG[5] ,
    \Tile_X9Y12_W6BEG[4] ,
    \Tile_X9Y12_W6BEG[3] ,
    \Tile_X9Y12_W6BEG[2] ,
    \Tile_X9Y12_W6BEG[1] ,
    \Tile_X9Y12_W6BEG[0] }),
    .WW4BEG({\Tile_X8Y12_WW4BEG[15] ,
    \Tile_X8Y12_WW4BEG[14] ,
    \Tile_X8Y12_WW4BEG[13] ,
    \Tile_X8Y12_WW4BEG[12] ,
    \Tile_X8Y12_WW4BEG[11] ,
    \Tile_X8Y12_WW4BEG[10] ,
    \Tile_X8Y12_WW4BEG[9] ,
    \Tile_X8Y12_WW4BEG[8] ,
    \Tile_X8Y12_WW4BEG[7] ,
    \Tile_X8Y12_WW4BEG[6] ,
    \Tile_X8Y12_WW4BEG[5] ,
    \Tile_X8Y12_WW4BEG[4] ,
    \Tile_X8Y12_WW4BEG[3] ,
    \Tile_X8Y12_WW4BEG[2] ,
    \Tile_X8Y12_WW4BEG[1] ,
    \Tile_X8Y12_WW4BEG[0] }),
    .WW4END({\Tile_X9Y12_WW4BEG[15] ,
    \Tile_X9Y12_WW4BEG[14] ,
    \Tile_X9Y12_WW4BEG[13] ,
    \Tile_X9Y12_WW4BEG[12] ,
    \Tile_X9Y12_WW4BEG[11] ,
    \Tile_X9Y12_WW4BEG[10] ,
    \Tile_X9Y12_WW4BEG[9] ,
    \Tile_X9Y12_WW4BEG[8] ,
    \Tile_X9Y12_WW4BEG[7] ,
    \Tile_X9Y12_WW4BEG[6] ,
    \Tile_X9Y12_WW4BEG[5] ,
    \Tile_X9Y12_WW4BEG[4] ,
    \Tile_X9Y12_WW4BEG[3] ,
    \Tile_X9Y12_WW4BEG[2] ,
    \Tile_X9Y12_WW4BEG[1] ,
    \Tile_X9Y12_WW4BEG[0] }));
 LUT4AB Tile_X8Y13_LUT4AB (.Ci(Tile_X8Y14_Co),
    .Co(Tile_X8Y13_Co),
    .UserCLK(Tile_X8Y14_UserCLKo),
    .UserCLKo(Tile_X8Y13_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X8Y13_E1BEG[3] ,
    \Tile_X8Y13_E1BEG[2] ,
    \Tile_X8Y13_E1BEG[1] ,
    \Tile_X8Y13_E1BEG[0] }),
    .E1END({\Tile_X7Y13_E1BEG[3] ,
    \Tile_X7Y13_E1BEG[2] ,
    \Tile_X7Y13_E1BEG[1] ,
    \Tile_X7Y13_E1BEG[0] }),
    .E2BEG({\Tile_X8Y13_E2BEG[7] ,
    \Tile_X8Y13_E2BEG[6] ,
    \Tile_X8Y13_E2BEG[5] ,
    \Tile_X8Y13_E2BEG[4] ,
    \Tile_X8Y13_E2BEG[3] ,
    \Tile_X8Y13_E2BEG[2] ,
    \Tile_X8Y13_E2BEG[1] ,
    \Tile_X8Y13_E2BEG[0] }),
    .E2BEGb({\Tile_X8Y13_E2BEGb[7] ,
    \Tile_X8Y13_E2BEGb[6] ,
    \Tile_X8Y13_E2BEGb[5] ,
    \Tile_X8Y13_E2BEGb[4] ,
    \Tile_X8Y13_E2BEGb[3] ,
    \Tile_X8Y13_E2BEGb[2] ,
    \Tile_X8Y13_E2BEGb[1] ,
    \Tile_X8Y13_E2BEGb[0] }),
    .E2END({\Tile_X7Y13_E2BEGb[7] ,
    \Tile_X7Y13_E2BEGb[6] ,
    \Tile_X7Y13_E2BEGb[5] ,
    \Tile_X7Y13_E2BEGb[4] ,
    \Tile_X7Y13_E2BEGb[3] ,
    \Tile_X7Y13_E2BEGb[2] ,
    \Tile_X7Y13_E2BEGb[1] ,
    \Tile_X7Y13_E2BEGb[0] }),
    .E2MID({\Tile_X7Y13_E2BEG[7] ,
    \Tile_X7Y13_E2BEG[6] ,
    \Tile_X7Y13_E2BEG[5] ,
    \Tile_X7Y13_E2BEG[4] ,
    \Tile_X7Y13_E2BEG[3] ,
    \Tile_X7Y13_E2BEG[2] ,
    \Tile_X7Y13_E2BEG[1] ,
    \Tile_X7Y13_E2BEG[0] }),
    .E6BEG({\Tile_X8Y13_E6BEG[11] ,
    \Tile_X8Y13_E6BEG[10] ,
    \Tile_X8Y13_E6BEG[9] ,
    \Tile_X8Y13_E6BEG[8] ,
    \Tile_X8Y13_E6BEG[7] ,
    \Tile_X8Y13_E6BEG[6] ,
    \Tile_X8Y13_E6BEG[5] ,
    \Tile_X8Y13_E6BEG[4] ,
    \Tile_X8Y13_E6BEG[3] ,
    \Tile_X8Y13_E6BEG[2] ,
    \Tile_X8Y13_E6BEG[1] ,
    \Tile_X8Y13_E6BEG[0] }),
    .E6END({\Tile_X7Y13_E6BEG[11] ,
    \Tile_X7Y13_E6BEG[10] ,
    \Tile_X7Y13_E6BEG[9] ,
    \Tile_X7Y13_E6BEG[8] ,
    \Tile_X7Y13_E6BEG[7] ,
    \Tile_X7Y13_E6BEG[6] ,
    \Tile_X7Y13_E6BEG[5] ,
    \Tile_X7Y13_E6BEG[4] ,
    \Tile_X7Y13_E6BEG[3] ,
    \Tile_X7Y13_E6BEG[2] ,
    \Tile_X7Y13_E6BEG[1] ,
    \Tile_X7Y13_E6BEG[0] }),
    .EE4BEG({\Tile_X8Y13_EE4BEG[15] ,
    \Tile_X8Y13_EE4BEG[14] ,
    \Tile_X8Y13_EE4BEG[13] ,
    \Tile_X8Y13_EE4BEG[12] ,
    \Tile_X8Y13_EE4BEG[11] ,
    \Tile_X8Y13_EE4BEG[10] ,
    \Tile_X8Y13_EE4BEG[9] ,
    \Tile_X8Y13_EE4BEG[8] ,
    \Tile_X8Y13_EE4BEG[7] ,
    \Tile_X8Y13_EE4BEG[6] ,
    \Tile_X8Y13_EE4BEG[5] ,
    \Tile_X8Y13_EE4BEG[4] ,
    \Tile_X8Y13_EE4BEG[3] ,
    \Tile_X8Y13_EE4BEG[2] ,
    \Tile_X8Y13_EE4BEG[1] ,
    \Tile_X8Y13_EE4BEG[0] }),
    .EE4END({\Tile_X7Y13_EE4BEG[15] ,
    \Tile_X7Y13_EE4BEG[14] ,
    \Tile_X7Y13_EE4BEG[13] ,
    \Tile_X7Y13_EE4BEG[12] ,
    \Tile_X7Y13_EE4BEG[11] ,
    \Tile_X7Y13_EE4BEG[10] ,
    \Tile_X7Y13_EE4BEG[9] ,
    \Tile_X7Y13_EE4BEG[8] ,
    \Tile_X7Y13_EE4BEG[7] ,
    \Tile_X7Y13_EE4BEG[6] ,
    \Tile_X7Y13_EE4BEG[5] ,
    \Tile_X7Y13_EE4BEG[4] ,
    \Tile_X7Y13_EE4BEG[3] ,
    \Tile_X7Y13_EE4BEG[2] ,
    \Tile_X7Y13_EE4BEG[1] ,
    \Tile_X7Y13_EE4BEG[0] }),
    .FrameData({\Tile_X7Y13_FrameData_O[31] ,
    \Tile_X7Y13_FrameData_O[30] ,
    \Tile_X7Y13_FrameData_O[29] ,
    \Tile_X7Y13_FrameData_O[28] ,
    \Tile_X7Y13_FrameData_O[27] ,
    \Tile_X7Y13_FrameData_O[26] ,
    \Tile_X7Y13_FrameData_O[25] ,
    \Tile_X7Y13_FrameData_O[24] ,
    \Tile_X7Y13_FrameData_O[23] ,
    \Tile_X7Y13_FrameData_O[22] ,
    \Tile_X7Y13_FrameData_O[21] ,
    \Tile_X7Y13_FrameData_O[20] ,
    \Tile_X7Y13_FrameData_O[19] ,
    \Tile_X7Y13_FrameData_O[18] ,
    \Tile_X7Y13_FrameData_O[17] ,
    \Tile_X7Y13_FrameData_O[16] ,
    \Tile_X7Y13_FrameData_O[15] ,
    \Tile_X7Y13_FrameData_O[14] ,
    \Tile_X7Y13_FrameData_O[13] ,
    \Tile_X7Y13_FrameData_O[12] ,
    \Tile_X7Y13_FrameData_O[11] ,
    \Tile_X7Y13_FrameData_O[10] ,
    \Tile_X7Y13_FrameData_O[9] ,
    \Tile_X7Y13_FrameData_O[8] ,
    \Tile_X7Y13_FrameData_O[7] ,
    \Tile_X7Y13_FrameData_O[6] ,
    \Tile_X7Y13_FrameData_O[5] ,
    \Tile_X7Y13_FrameData_O[4] ,
    \Tile_X7Y13_FrameData_O[3] ,
    \Tile_X7Y13_FrameData_O[2] ,
    \Tile_X7Y13_FrameData_O[1] ,
    \Tile_X7Y13_FrameData_O[0] }),
    .FrameData_O({\Tile_X8Y13_FrameData_O[31] ,
    \Tile_X8Y13_FrameData_O[30] ,
    \Tile_X8Y13_FrameData_O[29] ,
    \Tile_X8Y13_FrameData_O[28] ,
    \Tile_X8Y13_FrameData_O[27] ,
    \Tile_X8Y13_FrameData_O[26] ,
    \Tile_X8Y13_FrameData_O[25] ,
    \Tile_X8Y13_FrameData_O[24] ,
    \Tile_X8Y13_FrameData_O[23] ,
    \Tile_X8Y13_FrameData_O[22] ,
    \Tile_X8Y13_FrameData_O[21] ,
    \Tile_X8Y13_FrameData_O[20] ,
    \Tile_X8Y13_FrameData_O[19] ,
    \Tile_X8Y13_FrameData_O[18] ,
    \Tile_X8Y13_FrameData_O[17] ,
    \Tile_X8Y13_FrameData_O[16] ,
    \Tile_X8Y13_FrameData_O[15] ,
    \Tile_X8Y13_FrameData_O[14] ,
    \Tile_X8Y13_FrameData_O[13] ,
    \Tile_X8Y13_FrameData_O[12] ,
    \Tile_X8Y13_FrameData_O[11] ,
    \Tile_X8Y13_FrameData_O[10] ,
    \Tile_X8Y13_FrameData_O[9] ,
    \Tile_X8Y13_FrameData_O[8] ,
    \Tile_X8Y13_FrameData_O[7] ,
    \Tile_X8Y13_FrameData_O[6] ,
    \Tile_X8Y13_FrameData_O[5] ,
    \Tile_X8Y13_FrameData_O[4] ,
    \Tile_X8Y13_FrameData_O[3] ,
    \Tile_X8Y13_FrameData_O[2] ,
    \Tile_X8Y13_FrameData_O[1] ,
    \Tile_X8Y13_FrameData_O[0] }),
    .FrameStrobe({\Tile_X8Y14_FrameStrobe_O[19] ,
    \Tile_X8Y14_FrameStrobe_O[18] ,
    \Tile_X8Y14_FrameStrobe_O[17] ,
    \Tile_X8Y14_FrameStrobe_O[16] ,
    \Tile_X8Y14_FrameStrobe_O[15] ,
    \Tile_X8Y14_FrameStrobe_O[14] ,
    \Tile_X8Y14_FrameStrobe_O[13] ,
    \Tile_X8Y14_FrameStrobe_O[12] ,
    \Tile_X8Y14_FrameStrobe_O[11] ,
    \Tile_X8Y14_FrameStrobe_O[10] ,
    \Tile_X8Y14_FrameStrobe_O[9] ,
    \Tile_X8Y14_FrameStrobe_O[8] ,
    \Tile_X8Y14_FrameStrobe_O[7] ,
    \Tile_X8Y14_FrameStrobe_O[6] ,
    \Tile_X8Y14_FrameStrobe_O[5] ,
    \Tile_X8Y14_FrameStrobe_O[4] ,
    \Tile_X8Y14_FrameStrobe_O[3] ,
    \Tile_X8Y14_FrameStrobe_O[2] ,
    \Tile_X8Y14_FrameStrobe_O[1] ,
    \Tile_X8Y14_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X8Y13_FrameStrobe_O[19] ,
    \Tile_X8Y13_FrameStrobe_O[18] ,
    \Tile_X8Y13_FrameStrobe_O[17] ,
    \Tile_X8Y13_FrameStrobe_O[16] ,
    \Tile_X8Y13_FrameStrobe_O[15] ,
    \Tile_X8Y13_FrameStrobe_O[14] ,
    \Tile_X8Y13_FrameStrobe_O[13] ,
    \Tile_X8Y13_FrameStrobe_O[12] ,
    \Tile_X8Y13_FrameStrobe_O[11] ,
    \Tile_X8Y13_FrameStrobe_O[10] ,
    \Tile_X8Y13_FrameStrobe_O[9] ,
    \Tile_X8Y13_FrameStrobe_O[8] ,
    \Tile_X8Y13_FrameStrobe_O[7] ,
    \Tile_X8Y13_FrameStrobe_O[6] ,
    \Tile_X8Y13_FrameStrobe_O[5] ,
    \Tile_X8Y13_FrameStrobe_O[4] ,
    \Tile_X8Y13_FrameStrobe_O[3] ,
    \Tile_X8Y13_FrameStrobe_O[2] ,
    \Tile_X8Y13_FrameStrobe_O[1] ,
    \Tile_X8Y13_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X8Y13_N1BEG[3] ,
    \Tile_X8Y13_N1BEG[2] ,
    \Tile_X8Y13_N1BEG[1] ,
    \Tile_X8Y13_N1BEG[0] }),
    .N1END({\Tile_X8Y14_N1BEG[3] ,
    \Tile_X8Y14_N1BEG[2] ,
    \Tile_X8Y14_N1BEG[1] ,
    \Tile_X8Y14_N1BEG[0] }),
    .N2BEG({\Tile_X8Y13_N2BEG[7] ,
    \Tile_X8Y13_N2BEG[6] ,
    \Tile_X8Y13_N2BEG[5] ,
    \Tile_X8Y13_N2BEG[4] ,
    \Tile_X8Y13_N2BEG[3] ,
    \Tile_X8Y13_N2BEG[2] ,
    \Tile_X8Y13_N2BEG[1] ,
    \Tile_X8Y13_N2BEG[0] }),
    .N2BEGb({\Tile_X8Y13_N2BEGb[7] ,
    \Tile_X8Y13_N2BEGb[6] ,
    \Tile_X8Y13_N2BEGb[5] ,
    \Tile_X8Y13_N2BEGb[4] ,
    \Tile_X8Y13_N2BEGb[3] ,
    \Tile_X8Y13_N2BEGb[2] ,
    \Tile_X8Y13_N2BEGb[1] ,
    \Tile_X8Y13_N2BEGb[0] }),
    .N2END({\Tile_X8Y14_N2BEGb[7] ,
    \Tile_X8Y14_N2BEGb[6] ,
    \Tile_X8Y14_N2BEGb[5] ,
    \Tile_X8Y14_N2BEGb[4] ,
    \Tile_X8Y14_N2BEGb[3] ,
    \Tile_X8Y14_N2BEGb[2] ,
    \Tile_X8Y14_N2BEGb[1] ,
    \Tile_X8Y14_N2BEGb[0] }),
    .N2MID({\Tile_X8Y14_N2BEG[7] ,
    \Tile_X8Y14_N2BEG[6] ,
    \Tile_X8Y14_N2BEG[5] ,
    \Tile_X8Y14_N2BEG[4] ,
    \Tile_X8Y14_N2BEG[3] ,
    \Tile_X8Y14_N2BEG[2] ,
    \Tile_X8Y14_N2BEG[1] ,
    \Tile_X8Y14_N2BEG[0] }),
    .N4BEG({\Tile_X8Y13_N4BEG[15] ,
    \Tile_X8Y13_N4BEG[14] ,
    \Tile_X8Y13_N4BEG[13] ,
    \Tile_X8Y13_N4BEG[12] ,
    \Tile_X8Y13_N4BEG[11] ,
    \Tile_X8Y13_N4BEG[10] ,
    \Tile_X8Y13_N4BEG[9] ,
    \Tile_X8Y13_N4BEG[8] ,
    \Tile_X8Y13_N4BEG[7] ,
    \Tile_X8Y13_N4BEG[6] ,
    \Tile_X8Y13_N4BEG[5] ,
    \Tile_X8Y13_N4BEG[4] ,
    \Tile_X8Y13_N4BEG[3] ,
    \Tile_X8Y13_N4BEG[2] ,
    \Tile_X8Y13_N4BEG[1] ,
    \Tile_X8Y13_N4BEG[0] }),
    .N4END({\Tile_X8Y14_N4BEG[15] ,
    \Tile_X8Y14_N4BEG[14] ,
    \Tile_X8Y14_N4BEG[13] ,
    \Tile_X8Y14_N4BEG[12] ,
    \Tile_X8Y14_N4BEG[11] ,
    \Tile_X8Y14_N4BEG[10] ,
    \Tile_X8Y14_N4BEG[9] ,
    \Tile_X8Y14_N4BEG[8] ,
    \Tile_X8Y14_N4BEG[7] ,
    \Tile_X8Y14_N4BEG[6] ,
    \Tile_X8Y14_N4BEG[5] ,
    \Tile_X8Y14_N4BEG[4] ,
    \Tile_X8Y14_N4BEG[3] ,
    \Tile_X8Y14_N4BEG[2] ,
    \Tile_X8Y14_N4BEG[1] ,
    \Tile_X8Y14_N4BEG[0] }),
    .NN4BEG({\Tile_X8Y13_NN4BEG[15] ,
    \Tile_X8Y13_NN4BEG[14] ,
    \Tile_X8Y13_NN4BEG[13] ,
    \Tile_X8Y13_NN4BEG[12] ,
    \Tile_X8Y13_NN4BEG[11] ,
    \Tile_X8Y13_NN4BEG[10] ,
    \Tile_X8Y13_NN4BEG[9] ,
    \Tile_X8Y13_NN4BEG[8] ,
    \Tile_X8Y13_NN4BEG[7] ,
    \Tile_X8Y13_NN4BEG[6] ,
    \Tile_X8Y13_NN4BEG[5] ,
    \Tile_X8Y13_NN4BEG[4] ,
    \Tile_X8Y13_NN4BEG[3] ,
    \Tile_X8Y13_NN4BEG[2] ,
    \Tile_X8Y13_NN4BEG[1] ,
    \Tile_X8Y13_NN4BEG[0] }),
    .NN4END({\Tile_X8Y14_NN4BEG[15] ,
    \Tile_X8Y14_NN4BEG[14] ,
    \Tile_X8Y14_NN4BEG[13] ,
    \Tile_X8Y14_NN4BEG[12] ,
    \Tile_X8Y14_NN4BEG[11] ,
    \Tile_X8Y14_NN4BEG[10] ,
    \Tile_X8Y14_NN4BEG[9] ,
    \Tile_X8Y14_NN4BEG[8] ,
    \Tile_X8Y14_NN4BEG[7] ,
    \Tile_X8Y14_NN4BEG[6] ,
    \Tile_X8Y14_NN4BEG[5] ,
    \Tile_X8Y14_NN4BEG[4] ,
    \Tile_X8Y14_NN4BEG[3] ,
    \Tile_X8Y14_NN4BEG[2] ,
    \Tile_X8Y14_NN4BEG[1] ,
    \Tile_X8Y14_NN4BEG[0] }),
    .S1BEG({\Tile_X8Y13_S1BEG[3] ,
    \Tile_X8Y13_S1BEG[2] ,
    \Tile_X8Y13_S1BEG[1] ,
    \Tile_X8Y13_S1BEG[0] }),
    .S1END({\Tile_X8Y12_S1BEG[3] ,
    \Tile_X8Y12_S1BEG[2] ,
    \Tile_X8Y12_S1BEG[1] ,
    \Tile_X8Y12_S1BEG[0] }),
    .S2BEG({\Tile_X8Y13_S2BEG[7] ,
    \Tile_X8Y13_S2BEG[6] ,
    \Tile_X8Y13_S2BEG[5] ,
    \Tile_X8Y13_S2BEG[4] ,
    \Tile_X8Y13_S2BEG[3] ,
    \Tile_X8Y13_S2BEG[2] ,
    \Tile_X8Y13_S2BEG[1] ,
    \Tile_X8Y13_S2BEG[0] }),
    .S2BEGb({\Tile_X8Y13_S2BEGb[7] ,
    \Tile_X8Y13_S2BEGb[6] ,
    \Tile_X8Y13_S2BEGb[5] ,
    \Tile_X8Y13_S2BEGb[4] ,
    \Tile_X8Y13_S2BEGb[3] ,
    \Tile_X8Y13_S2BEGb[2] ,
    \Tile_X8Y13_S2BEGb[1] ,
    \Tile_X8Y13_S2BEGb[0] }),
    .S2END({\Tile_X8Y12_S2BEGb[7] ,
    \Tile_X8Y12_S2BEGb[6] ,
    \Tile_X8Y12_S2BEGb[5] ,
    \Tile_X8Y12_S2BEGb[4] ,
    \Tile_X8Y12_S2BEGb[3] ,
    \Tile_X8Y12_S2BEGb[2] ,
    \Tile_X8Y12_S2BEGb[1] ,
    \Tile_X8Y12_S2BEGb[0] }),
    .S2MID({\Tile_X8Y12_S2BEG[7] ,
    \Tile_X8Y12_S2BEG[6] ,
    \Tile_X8Y12_S2BEG[5] ,
    \Tile_X8Y12_S2BEG[4] ,
    \Tile_X8Y12_S2BEG[3] ,
    \Tile_X8Y12_S2BEG[2] ,
    \Tile_X8Y12_S2BEG[1] ,
    \Tile_X8Y12_S2BEG[0] }),
    .S4BEG({\Tile_X8Y13_S4BEG[15] ,
    \Tile_X8Y13_S4BEG[14] ,
    \Tile_X8Y13_S4BEG[13] ,
    \Tile_X8Y13_S4BEG[12] ,
    \Tile_X8Y13_S4BEG[11] ,
    \Tile_X8Y13_S4BEG[10] ,
    \Tile_X8Y13_S4BEG[9] ,
    \Tile_X8Y13_S4BEG[8] ,
    \Tile_X8Y13_S4BEG[7] ,
    \Tile_X8Y13_S4BEG[6] ,
    \Tile_X8Y13_S4BEG[5] ,
    \Tile_X8Y13_S4BEG[4] ,
    \Tile_X8Y13_S4BEG[3] ,
    \Tile_X8Y13_S4BEG[2] ,
    \Tile_X8Y13_S4BEG[1] ,
    \Tile_X8Y13_S4BEG[0] }),
    .S4END({\Tile_X8Y12_S4BEG[15] ,
    \Tile_X8Y12_S4BEG[14] ,
    \Tile_X8Y12_S4BEG[13] ,
    \Tile_X8Y12_S4BEG[12] ,
    \Tile_X8Y12_S4BEG[11] ,
    \Tile_X8Y12_S4BEG[10] ,
    \Tile_X8Y12_S4BEG[9] ,
    \Tile_X8Y12_S4BEG[8] ,
    \Tile_X8Y12_S4BEG[7] ,
    \Tile_X8Y12_S4BEG[6] ,
    \Tile_X8Y12_S4BEG[5] ,
    \Tile_X8Y12_S4BEG[4] ,
    \Tile_X8Y12_S4BEG[3] ,
    \Tile_X8Y12_S4BEG[2] ,
    \Tile_X8Y12_S4BEG[1] ,
    \Tile_X8Y12_S4BEG[0] }),
    .SS4BEG({\Tile_X8Y13_SS4BEG[15] ,
    \Tile_X8Y13_SS4BEG[14] ,
    \Tile_X8Y13_SS4BEG[13] ,
    \Tile_X8Y13_SS4BEG[12] ,
    \Tile_X8Y13_SS4BEG[11] ,
    \Tile_X8Y13_SS4BEG[10] ,
    \Tile_X8Y13_SS4BEG[9] ,
    \Tile_X8Y13_SS4BEG[8] ,
    \Tile_X8Y13_SS4BEG[7] ,
    \Tile_X8Y13_SS4BEG[6] ,
    \Tile_X8Y13_SS4BEG[5] ,
    \Tile_X8Y13_SS4BEG[4] ,
    \Tile_X8Y13_SS4BEG[3] ,
    \Tile_X8Y13_SS4BEG[2] ,
    \Tile_X8Y13_SS4BEG[1] ,
    \Tile_X8Y13_SS4BEG[0] }),
    .SS4END({\Tile_X8Y12_SS4BEG[15] ,
    \Tile_X8Y12_SS4BEG[14] ,
    \Tile_X8Y12_SS4BEG[13] ,
    \Tile_X8Y12_SS4BEG[12] ,
    \Tile_X8Y12_SS4BEG[11] ,
    \Tile_X8Y12_SS4BEG[10] ,
    \Tile_X8Y12_SS4BEG[9] ,
    \Tile_X8Y12_SS4BEG[8] ,
    \Tile_X8Y12_SS4BEG[7] ,
    \Tile_X8Y12_SS4BEG[6] ,
    \Tile_X8Y12_SS4BEG[5] ,
    \Tile_X8Y12_SS4BEG[4] ,
    \Tile_X8Y12_SS4BEG[3] ,
    \Tile_X8Y12_SS4BEG[2] ,
    \Tile_X8Y12_SS4BEG[1] ,
    \Tile_X8Y12_SS4BEG[0] }),
    .W1BEG({\Tile_X8Y13_W1BEG[3] ,
    \Tile_X8Y13_W1BEG[2] ,
    \Tile_X8Y13_W1BEG[1] ,
    \Tile_X8Y13_W1BEG[0] }),
    .W1END({\Tile_X9Y13_W1BEG[3] ,
    \Tile_X9Y13_W1BEG[2] ,
    \Tile_X9Y13_W1BEG[1] ,
    \Tile_X9Y13_W1BEG[0] }),
    .W2BEG({\Tile_X8Y13_W2BEG[7] ,
    \Tile_X8Y13_W2BEG[6] ,
    \Tile_X8Y13_W2BEG[5] ,
    \Tile_X8Y13_W2BEG[4] ,
    \Tile_X8Y13_W2BEG[3] ,
    \Tile_X8Y13_W2BEG[2] ,
    \Tile_X8Y13_W2BEG[1] ,
    \Tile_X8Y13_W2BEG[0] }),
    .W2BEGb({\Tile_X8Y13_W2BEGb[7] ,
    \Tile_X8Y13_W2BEGb[6] ,
    \Tile_X8Y13_W2BEGb[5] ,
    \Tile_X8Y13_W2BEGb[4] ,
    \Tile_X8Y13_W2BEGb[3] ,
    \Tile_X8Y13_W2BEGb[2] ,
    \Tile_X8Y13_W2BEGb[1] ,
    \Tile_X8Y13_W2BEGb[0] }),
    .W2END({\Tile_X9Y13_W2BEGb[7] ,
    \Tile_X9Y13_W2BEGb[6] ,
    \Tile_X9Y13_W2BEGb[5] ,
    \Tile_X9Y13_W2BEGb[4] ,
    \Tile_X9Y13_W2BEGb[3] ,
    \Tile_X9Y13_W2BEGb[2] ,
    \Tile_X9Y13_W2BEGb[1] ,
    \Tile_X9Y13_W2BEGb[0] }),
    .W2MID({\Tile_X9Y13_W2BEG[7] ,
    \Tile_X9Y13_W2BEG[6] ,
    \Tile_X9Y13_W2BEG[5] ,
    \Tile_X9Y13_W2BEG[4] ,
    \Tile_X9Y13_W2BEG[3] ,
    \Tile_X9Y13_W2BEG[2] ,
    \Tile_X9Y13_W2BEG[1] ,
    \Tile_X9Y13_W2BEG[0] }),
    .W6BEG({\Tile_X8Y13_W6BEG[11] ,
    \Tile_X8Y13_W6BEG[10] ,
    \Tile_X8Y13_W6BEG[9] ,
    \Tile_X8Y13_W6BEG[8] ,
    \Tile_X8Y13_W6BEG[7] ,
    \Tile_X8Y13_W6BEG[6] ,
    \Tile_X8Y13_W6BEG[5] ,
    \Tile_X8Y13_W6BEG[4] ,
    \Tile_X8Y13_W6BEG[3] ,
    \Tile_X8Y13_W6BEG[2] ,
    \Tile_X8Y13_W6BEG[1] ,
    \Tile_X8Y13_W6BEG[0] }),
    .W6END({\Tile_X9Y13_W6BEG[11] ,
    \Tile_X9Y13_W6BEG[10] ,
    \Tile_X9Y13_W6BEG[9] ,
    \Tile_X9Y13_W6BEG[8] ,
    \Tile_X9Y13_W6BEG[7] ,
    \Tile_X9Y13_W6BEG[6] ,
    \Tile_X9Y13_W6BEG[5] ,
    \Tile_X9Y13_W6BEG[4] ,
    \Tile_X9Y13_W6BEG[3] ,
    \Tile_X9Y13_W6BEG[2] ,
    \Tile_X9Y13_W6BEG[1] ,
    \Tile_X9Y13_W6BEG[0] }),
    .WW4BEG({\Tile_X8Y13_WW4BEG[15] ,
    \Tile_X8Y13_WW4BEG[14] ,
    \Tile_X8Y13_WW4BEG[13] ,
    \Tile_X8Y13_WW4BEG[12] ,
    \Tile_X8Y13_WW4BEG[11] ,
    \Tile_X8Y13_WW4BEG[10] ,
    \Tile_X8Y13_WW4BEG[9] ,
    \Tile_X8Y13_WW4BEG[8] ,
    \Tile_X8Y13_WW4BEG[7] ,
    \Tile_X8Y13_WW4BEG[6] ,
    \Tile_X8Y13_WW4BEG[5] ,
    \Tile_X8Y13_WW4BEG[4] ,
    \Tile_X8Y13_WW4BEG[3] ,
    \Tile_X8Y13_WW4BEG[2] ,
    \Tile_X8Y13_WW4BEG[1] ,
    \Tile_X8Y13_WW4BEG[0] }),
    .WW4END({\Tile_X9Y13_WW4BEG[15] ,
    \Tile_X9Y13_WW4BEG[14] ,
    \Tile_X9Y13_WW4BEG[13] ,
    \Tile_X9Y13_WW4BEG[12] ,
    \Tile_X9Y13_WW4BEG[11] ,
    \Tile_X9Y13_WW4BEG[10] ,
    \Tile_X9Y13_WW4BEG[9] ,
    \Tile_X9Y13_WW4BEG[8] ,
    \Tile_X9Y13_WW4BEG[7] ,
    \Tile_X9Y13_WW4BEG[6] ,
    \Tile_X9Y13_WW4BEG[5] ,
    \Tile_X9Y13_WW4BEG[4] ,
    \Tile_X9Y13_WW4BEG[3] ,
    \Tile_X9Y13_WW4BEG[2] ,
    \Tile_X9Y13_WW4BEG[1] ,
    \Tile_X9Y13_WW4BEG[0] }));
 LUT4AB Tile_X8Y14_LUT4AB (.Ci(Tile_X8Y15_Co),
    .Co(Tile_X8Y14_Co),
    .UserCLK(Tile_X8Y15_UserCLKo),
    .UserCLKo(Tile_X8Y14_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X8Y14_E1BEG[3] ,
    \Tile_X8Y14_E1BEG[2] ,
    \Tile_X8Y14_E1BEG[1] ,
    \Tile_X8Y14_E1BEG[0] }),
    .E1END({\Tile_X7Y14_E1BEG[3] ,
    \Tile_X7Y14_E1BEG[2] ,
    \Tile_X7Y14_E1BEG[1] ,
    \Tile_X7Y14_E1BEG[0] }),
    .E2BEG({\Tile_X8Y14_E2BEG[7] ,
    \Tile_X8Y14_E2BEG[6] ,
    \Tile_X8Y14_E2BEG[5] ,
    \Tile_X8Y14_E2BEG[4] ,
    \Tile_X8Y14_E2BEG[3] ,
    \Tile_X8Y14_E2BEG[2] ,
    \Tile_X8Y14_E2BEG[1] ,
    \Tile_X8Y14_E2BEG[0] }),
    .E2BEGb({\Tile_X8Y14_E2BEGb[7] ,
    \Tile_X8Y14_E2BEGb[6] ,
    \Tile_X8Y14_E2BEGb[5] ,
    \Tile_X8Y14_E2BEGb[4] ,
    \Tile_X8Y14_E2BEGb[3] ,
    \Tile_X8Y14_E2BEGb[2] ,
    \Tile_X8Y14_E2BEGb[1] ,
    \Tile_X8Y14_E2BEGb[0] }),
    .E2END({\Tile_X7Y14_E2BEGb[7] ,
    \Tile_X7Y14_E2BEGb[6] ,
    \Tile_X7Y14_E2BEGb[5] ,
    \Tile_X7Y14_E2BEGb[4] ,
    \Tile_X7Y14_E2BEGb[3] ,
    \Tile_X7Y14_E2BEGb[2] ,
    \Tile_X7Y14_E2BEGb[1] ,
    \Tile_X7Y14_E2BEGb[0] }),
    .E2MID({\Tile_X7Y14_E2BEG[7] ,
    \Tile_X7Y14_E2BEG[6] ,
    \Tile_X7Y14_E2BEG[5] ,
    \Tile_X7Y14_E2BEG[4] ,
    \Tile_X7Y14_E2BEG[3] ,
    \Tile_X7Y14_E2BEG[2] ,
    \Tile_X7Y14_E2BEG[1] ,
    \Tile_X7Y14_E2BEG[0] }),
    .E6BEG({\Tile_X8Y14_E6BEG[11] ,
    \Tile_X8Y14_E6BEG[10] ,
    \Tile_X8Y14_E6BEG[9] ,
    \Tile_X8Y14_E6BEG[8] ,
    \Tile_X8Y14_E6BEG[7] ,
    \Tile_X8Y14_E6BEG[6] ,
    \Tile_X8Y14_E6BEG[5] ,
    \Tile_X8Y14_E6BEG[4] ,
    \Tile_X8Y14_E6BEG[3] ,
    \Tile_X8Y14_E6BEG[2] ,
    \Tile_X8Y14_E6BEG[1] ,
    \Tile_X8Y14_E6BEG[0] }),
    .E6END({\Tile_X7Y14_E6BEG[11] ,
    \Tile_X7Y14_E6BEG[10] ,
    \Tile_X7Y14_E6BEG[9] ,
    \Tile_X7Y14_E6BEG[8] ,
    \Tile_X7Y14_E6BEG[7] ,
    \Tile_X7Y14_E6BEG[6] ,
    \Tile_X7Y14_E6BEG[5] ,
    \Tile_X7Y14_E6BEG[4] ,
    \Tile_X7Y14_E6BEG[3] ,
    \Tile_X7Y14_E6BEG[2] ,
    \Tile_X7Y14_E6BEG[1] ,
    \Tile_X7Y14_E6BEG[0] }),
    .EE4BEG({\Tile_X8Y14_EE4BEG[15] ,
    \Tile_X8Y14_EE4BEG[14] ,
    \Tile_X8Y14_EE4BEG[13] ,
    \Tile_X8Y14_EE4BEG[12] ,
    \Tile_X8Y14_EE4BEG[11] ,
    \Tile_X8Y14_EE4BEG[10] ,
    \Tile_X8Y14_EE4BEG[9] ,
    \Tile_X8Y14_EE4BEG[8] ,
    \Tile_X8Y14_EE4BEG[7] ,
    \Tile_X8Y14_EE4BEG[6] ,
    \Tile_X8Y14_EE4BEG[5] ,
    \Tile_X8Y14_EE4BEG[4] ,
    \Tile_X8Y14_EE4BEG[3] ,
    \Tile_X8Y14_EE4BEG[2] ,
    \Tile_X8Y14_EE4BEG[1] ,
    \Tile_X8Y14_EE4BEG[0] }),
    .EE4END({\Tile_X7Y14_EE4BEG[15] ,
    \Tile_X7Y14_EE4BEG[14] ,
    \Tile_X7Y14_EE4BEG[13] ,
    \Tile_X7Y14_EE4BEG[12] ,
    \Tile_X7Y14_EE4BEG[11] ,
    \Tile_X7Y14_EE4BEG[10] ,
    \Tile_X7Y14_EE4BEG[9] ,
    \Tile_X7Y14_EE4BEG[8] ,
    \Tile_X7Y14_EE4BEG[7] ,
    \Tile_X7Y14_EE4BEG[6] ,
    \Tile_X7Y14_EE4BEG[5] ,
    \Tile_X7Y14_EE4BEG[4] ,
    \Tile_X7Y14_EE4BEG[3] ,
    \Tile_X7Y14_EE4BEG[2] ,
    \Tile_X7Y14_EE4BEG[1] ,
    \Tile_X7Y14_EE4BEG[0] }),
    .FrameData({\Tile_X7Y14_FrameData_O[31] ,
    \Tile_X7Y14_FrameData_O[30] ,
    \Tile_X7Y14_FrameData_O[29] ,
    \Tile_X7Y14_FrameData_O[28] ,
    \Tile_X7Y14_FrameData_O[27] ,
    \Tile_X7Y14_FrameData_O[26] ,
    \Tile_X7Y14_FrameData_O[25] ,
    \Tile_X7Y14_FrameData_O[24] ,
    \Tile_X7Y14_FrameData_O[23] ,
    \Tile_X7Y14_FrameData_O[22] ,
    \Tile_X7Y14_FrameData_O[21] ,
    \Tile_X7Y14_FrameData_O[20] ,
    \Tile_X7Y14_FrameData_O[19] ,
    \Tile_X7Y14_FrameData_O[18] ,
    \Tile_X7Y14_FrameData_O[17] ,
    \Tile_X7Y14_FrameData_O[16] ,
    \Tile_X7Y14_FrameData_O[15] ,
    \Tile_X7Y14_FrameData_O[14] ,
    \Tile_X7Y14_FrameData_O[13] ,
    \Tile_X7Y14_FrameData_O[12] ,
    \Tile_X7Y14_FrameData_O[11] ,
    \Tile_X7Y14_FrameData_O[10] ,
    \Tile_X7Y14_FrameData_O[9] ,
    \Tile_X7Y14_FrameData_O[8] ,
    \Tile_X7Y14_FrameData_O[7] ,
    \Tile_X7Y14_FrameData_O[6] ,
    \Tile_X7Y14_FrameData_O[5] ,
    \Tile_X7Y14_FrameData_O[4] ,
    \Tile_X7Y14_FrameData_O[3] ,
    \Tile_X7Y14_FrameData_O[2] ,
    \Tile_X7Y14_FrameData_O[1] ,
    \Tile_X7Y14_FrameData_O[0] }),
    .FrameData_O({\Tile_X8Y14_FrameData_O[31] ,
    \Tile_X8Y14_FrameData_O[30] ,
    \Tile_X8Y14_FrameData_O[29] ,
    \Tile_X8Y14_FrameData_O[28] ,
    \Tile_X8Y14_FrameData_O[27] ,
    \Tile_X8Y14_FrameData_O[26] ,
    \Tile_X8Y14_FrameData_O[25] ,
    \Tile_X8Y14_FrameData_O[24] ,
    \Tile_X8Y14_FrameData_O[23] ,
    \Tile_X8Y14_FrameData_O[22] ,
    \Tile_X8Y14_FrameData_O[21] ,
    \Tile_X8Y14_FrameData_O[20] ,
    \Tile_X8Y14_FrameData_O[19] ,
    \Tile_X8Y14_FrameData_O[18] ,
    \Tile_X8Y14_FrameData_O[17] ,
    \Tile_X8Y14_FrameData_O[16] ,
    \Tile_X8Y14_FrameData_O[15] ,
    \Tile_X8Y14_FrameData_O[14] ,
    \Tile_X8Y14_FrameData_O[13] ,
    \Tile_X8Y14_FrameData_O[12] ,
    \Tile_X8Y14_FrameData_O[11] ,
    \Tile_X8Y14_FrameData_O[10] ,
    \Tile_X8Y14_FrameData_O[9] ,
    \Tile_X8Y14_FrameData_O[8] ,
    \Tile_X8Y14_FrameData_O[7] ,
    \Tile_X8Y14_FrameData_O[6] ,
    \Tile_X8Y14_FrameData_O[5] ,
    \Tile_X8Y14_FrameData_O[4] ,
    \Tile_X8Y14_FrameData_O[3] ,
    \Tile_X8Y14_FrameData_O[2] ,
    \Tile_X8Y14_FrameData_O[1] ,
    \Tile_X8Y14_FrameData_O[0] }),
    .FrameStrobe({\Tile_X8Y15_FrameStrobe_O[19] ,
    \Tile_X8Y15_FrameStrobe_O[18] ,
    \Tile_X8Y15_FrameStrobe_O[17] ,
    \Tile_X8Y15_FrameStrobe_O[16] ,
    \Tile_X8Y15_FrameStrobe_O[15] ,
    \Tile_X8Y15_FrameStrobe_O[14] ,
    \Tile_X8Y15_FrameStrobe_O[13] ,
    \Tile_X8Y15_FrameStrobe_O[12] ,
    \Tile_X8Y15_FrameStrobe_O[11] ,
    \Tile_X8Y15_FrameStrobe_O[10] ,
    \Tile_X8Y15_FrameStrobe_O[9] ,
    \Tile_X8Y15_FrameStrobe_O[8] ,
    \Tile_X8Y15_FrameStrobe_O[7] ,
    \Tile_X8Y15_FrameStrobe_O[6] ,
    \Tile_X8Y15_FrameStrobe_O[5] ,
    \Tile_X8Y15_FrameStrobe_O[4] ,
    \Tile_X8Y15_FrameStrobe_O[3] ,
    \Tile_X8Y15_FrameStrobe_O[2] ,
    \Tile_X8Y15_FrameStrobe_O[1] ,
    \Tile_X8Y15_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X8Y14_FrameStrobe_O[19] ,
    \Tile_X8Y14_FrameStrobe_O[18] ,
    \Tile_X8Y14_FrameStrobe_O[17] ,
    \Tile_X8Y14_FrameStrobe_O[16] ,
    \Tile_X8Y14_FrameStrobe_O[15] ,
    \Tile_X8Y14_FrameStrobe_O[14] ,
    \Tile_X8Y14_FrameStrobe_O[13] ,
    \Tile_X8Y14_FrameStrobe_O[12] ,
    \Tile_X8Y14_FrameStrobe_O[11] ,
    \Tile_X8Y14_FrameStrobe_O[10] ,
    \Tile_X8Y14_FrameStrobe_O[9] ,
    \Tile_X8Y14_FrameStrobe_O[8] ,
    \Tile_X8Y14_FrameStrobe_O[7] ,
    \Tile_X8Y14_FrameStrobe_O[6] ,
    \Tile_X8Y14_FrameStrobe_O[5] ,
    \Tile_X8Y14_FrameStrobe_O[4] ,
    \Tile_X8Y14_FrameStrobe_O[3] ,
    \Tile_X8Y14_FrameStrobe_O[2] ,
    \Tile_X8Y14_FrameStrobe_O[1] ,
    \Tile_X8Y14_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X8Y14_N1BEG[3] ,
    \Tile_X8Y14_N1BEG[2] ,
    \Tile_X8Y14_N1BEG[1] ,
    \Tile_X8Y14_N1BEG[0] }),
    .N1END({\Tile_X8Y15_N1BEG[3] ,
    \Tile_X8Y15_N1BEG[2] ,
    \Tile_X8Y15_N1BEG[1] ,
    \Tile_X8Y15_N1BEG[0] }),
    .N2BEG({\Tile_X8Y14_N2BEG[7] ,
    \Tile_X8Y14_N2BEG[6] ,
    \Tile_X8Y14_N2BEG[5] ,
    \Tile_X8Y14_N2BEG[4] ,
    \Tile_X8Y14_N2BEG[3] ,
    \Tile_X8Y14_N2BEG[2] ,
    \Tile_X8Y14_N2BEG[1] ,
    \Tile_X8Y14_N2BEG[0] }),
    .N2BEGb({\Tile_X8Y14_N2BEGb[7] ,
    \Tile_X8Y14_N2BEGb[6] ,
    \Tile_X8Y14_N2BEGb[5] ,
    \Tile_X8Y14_N2BEGb[4] ,
    \Tile_X8Y14_N2BEGb[3] ,
    \Tile_X8Y14_N2BEGb[2] ,
    \Tile_X8Y14_N2BEGb[1] ,
    \Tile_X8Y14_N2BEGb[0] }),
    .N2END({\Tile_X8Y15_N2BEGb[7] ,
    \Tile_X8Y15_N2BEGb[6] ,
    \Tile_X8Y15_N2BEGb[5] ,
    \Tile_X8Y15_N2BEGb[4] ,
    \Tile_X8Y15_N2BEGb[3] ,
    \Tile_X8Y15_N2BEGb[2] ,
    \Tile_X8Y15_N2BEGb[1] ,
    \Tile_X8Y15_N2BEGb[0] }),
    .N2MID({\Tile_X8Y15_N2BEG[7] ,
    \Tile_X8Y15_N2BEG[6] ,
    \Tile_X8Y15_N2BEG[5] ,
    \Tile_X8Y15_N2BEG[4] ,
    \Tile_X8Y15_N2BEG[3] ,
    \Tile_X8Y15_N2BEG[2] ,
    \Tile_X8Y15_N2BEG[1] ,
    \Tile_X8Y15_N2BEG[0] }),
    .N4BEG({\Tile_X8Y14_N4BEG[15] ,
    \Tile_X8Y14_N4BEG[14] ,
    \Tile_X8Y14_N4BEG[13] ,
    \Tile_X8Y14_N4BEG[12] ,
    \Tile_X8Y14_N4BEG[11] ,
    \Tile_X8Y14_N4BEG[10] ,
    \Tile_X8Y14_N4BEG[9] ,
    \Tile_X8Y14_N4BEG[8] ,
    \Tile_X8Y14_N4BEG[7] ,
    \Tile_X8Y14_N4BEG[6] ,
    \Tile_X8Y14_N4BEG[5] ,
    \Tile_X8Y14_N4BEG[4] ,
    \Tile_X8Y14_N4BEG[3] ,
    \Tile_X8Y14_N4BEG[2] ,
    \Tile_X8Y14_N4BEG[1] ,
    \Tile_X8Y14_N4BEG[0] }),
    .N4END({\Tile_X8Y15_N4BEG[15] ,
    \Tile_X8Y15_N4BEG[14] ,
    \Tile_X8Y15_N4BEG[13] ,
    \Tile_X8Y15_N4BEG[12] ,
    \Tile_X8Y15_N4BEG[11] ,
    \Tile_X8Y15_N4BEG[10] ,
    \Tile_X8Y15_N4BEG[9] ,
    \Tile_X8Y15_N4BEG[8] ,
    \Tile_X8Y15_N4BEG[7] ,
    \Tile_X8Y15_N4BEG[6] ,
    \Tile_X8Y15_N4BEG[5] ,
    \Tile_X8Y15_N4BEG[4] ,
    \Tile_X8Y15_N4BEG[3] ,
    \Tile_X8Y15_N4BEG[2] ,
    \Tile_X8Y15_N4BEG[1] ,
    \Tile_X8Y15_N4BEG[0] }),
    .NN4BEG({\Tile_X8Y14_NN4BEG[15] ,
    \Tile_X8Y14_NN4BEG[14] ,
    \Tile_X8Y14_NN4BEG[13] ,
    \Tile_X8Y14_NN4BEG[12] ,
    \Tile_X8Y14_NN4BEG[11] ,
    \Tile_X8Y14_NN4BEG[10] ,
    \Tile_X8Y14_NN4BEG[9] ,
    \Tile_X8Y14_NN4BEG[8] ,
    \Tile_X8Y14_NN4BEG[7] ,
    \Tile_X8Y14_NN4BEG[6] ,
    \Tile_X8Y14_NN4BEG[5] ,
    \Tile_X8Y14_NN4BEG[4] ,
    \Tile_X8Y14_NN4BEG[3] ,
    \Tile_X8Y14_NN4BEG[2] ,
    \Tile_X8Y14_NN4BEG[1] ,
    \Tile_X8Y14_NN4BEG[0] }),
    .NN4END({\Tile_X8Y15_NN4BEG[15] ,
    \Tile_X8Y15_NN4BEG[14] ,
    \Tile_X8Y15_NN4BEG[13] ,
    \Tile_X8Y15_NN4BEG[12] ,
    \Tile_X8Y15_NN4BEG[11] ,
    \Tile_X8Y15_NN4BEG[10] ,
    \Tile_X8Y15_NN4BEG[9] ,
    \Tile_X8Y15_NN4BEG[8] ,
    \Tile_X8Y15_NN4BEG[7] ,
    \Tile_X8Y15_NN4BEG[6] ,
    \Tile_X8Y15_NN4BEG[5] ,
    \Tile_X8Y15_NN4BEG[4] ,
    \Tile_X8Y15_NN4BEG[3] ,
    \Tile_X8Y15_NN4BEG[2] ,
    \Tile_X8Y15_NN4BEG[1] ,
    \Tile_X8Y15_NN4BEG[0] }),
    .S1BEG({\Tile_X8Y14_S1BEG[3] ,
    \Tile_X8Y14_S1BEG[2] ,
    \Tile_X8Y14_S1BEG[1] ,
    \Tile_X8Y14_S1BEG[0] }),
    .S1END({\Tile_X8Y13_S1BEG[3] ,
    \Tile_X8Y13_S1BEG[2] ,
    \Tile_X8Y13_S1BEG[1] ,
    \Tile_X8Y13_S1BEG[0] }),
    .S2BEG({\Tile_X8Y14_S2BEG[7] ,
    \Tile_X8Y14_S2BEG[6] ,
    \Tile_X8Y14_S2BEG[5] ,
    \Tile_X8Y14_S2BEG[4] ,
    \Tile_X8Y14_S2BEG[3] ,
    \Tile_X8Y14_S2BEG[2] ,
    \Tile_X8Y14_S2BEG[1] ,
    \Tile_X8Y14_S2BEG[0] }),
    .S2BEGb({\Tile_X8Y14_S2BEGb[7] ,
    \Tile_X8Y14_S2BEGb[6] ,
    \Tile_X8Y14_S2BEGb[5] ,
    \Tile_X8Y14_S2BEGb[4] ,
    \Tile_X8Y14_S2BEGb[3] ,
    \Tile_X8Y14_S2BEGb[2] ,
    \Tile_X8Y14_S2BEGb[1] ,
    \Tile_X8Y14_S2BEGb[0] }),
    .S2END({\Tile_X8Y13_S2BEGb[7] ,
    \Tile_X8Y13_S2BEGb[6] ,
    \Tile_X8Y13_S2BEGb[5] ,
    \Tile_X8Y13_S2BEGb[4] ,
    \Tile_X8Y13_S2BEGb[3] ,
    \Tile_X8Y13_S2BEGb[2] ,
    \Tile_X8Y13_S2BEGb[1] ,
    \Tile_X8Y13_S2BEGb[0] }),
    .S2MID({\Tile_X8Y13_S2BEG[7] ,
    \Tile_X8Y13_S2BEG[6] ,
    \Tile_X8Y13_S2BEG[5] ,
    \Tile_X8Y13_S2BEG[4] ,
    \Tile_X8Y13_S2BEG[3] ,
    \Tile_X8Y13_S2BEG[2] ,
    \Tile_X8Y13_S2BEG[1] ,
    \Tile_X8Y13_S2BEG[0] }),
    .S4BEG({\Tile_X8Y14_S4BEG[15] ,
    \Tile_X8Y14_S4BEG[14] ,
    \Tile_X8Y14_S4BEG[13] ,
    \Tile_X8Y14_S4BEG[12] ,
    \Tile_X8Y14_S4BEG[11] ,
    \Tile_X8Y14_S4BEG[10] ,
    \Tile_X8Y14_S4BEG[9] ,
    \Tile_X8Y14_S4BEG[8] ,
    \Tile_X8Y14_S4BEG[7] ,
    \Tile_X8Y14_S4BEG[6] ,
    \Tile_X8Y14_S4BEG[5] ,
    \Tile_X8Y14_S4BEG[4] ,
    \Tile_X8Y14_S4BEG[3] ,
    \Tile_X8Y14_S4BEG[2] ,
    \Tile_X8Y14_S4BEG[1] ,
    \Tile_X8Y14_S4BEG[0] }),
    .S4END({\Tile_X8Y13_S4BEG[15] ,
    \Tile_X8Y13_S4BEG[14] ,
    \Tile_X8Y13_S4BEG[13] ,
    \Tile_X8Y13_S4BEG[12] ,
    \Tile_X8Y13_S4BEG[11] ,
    \Tile_X8Y13_S4BEG[10] ,
    \Tile_X8Y13_S4BEG[9] ,
    \Tile_X8Y13_S4BEG[8] ,
    \Tile_X8Y13_S4BEG[7] ,
    \Tile_X8Y13_S4BEG[6] ,
    \Tile_X8Y13_S4BEG[5] ,
    \Tile_X8Y13_S4BEG[4] ,
    \Tile_X8Y13_S4BEG[3] ,
    \Tile_X8Y13_S4BEG[2] ,
    \Tile_X8Y13_S4BEG[1] ,
    \Tile_X8Y13_S4BEG[0] }),
    .SS4BEG({\Tile_X8Y14_SS4BEG[15] ,
    \Tile_X8Y14_SS4BEG[14] ,
    \Tile_X8Y14_SS4BEG[13] ,
    \Tile_X8Y14_SS4BEG[12] ,
    \Tile_X8Y14_SS4BEG[11] ,
    \Tile_X8Y14_SS4BEG[10] ,
    \Tile_X8Y14_SS4BEG[9] ,
    \Tile_X8Y14_SS4BEG[8] ,
    \Tile_X8Y14_SS4BEG[7] ,
    \Tile_X8Y14_SS4BEG[6] ,
    \Tile_X8Y14_SS4BEG[5] ,
    \Tile_X8Y14_SS4BEG[4] ,
    \Tile_X8Y14_SS4BEG[3] ,
    \Tile_X8Y14_SS4BEG[2] ,
    \Tile_X8Y14_SS4BEG[1] ,
    \Tile_X8Y14_SS4BEG[0] }),
    .SS4END({\Tile_X8Y13_SS4BEG[15] ,
    \Tile_X8Y13_SS4BEG[14] ,
    \Tile_X8Y13_SS4BEG[13] ,
    \Tile_X8Y13_SS4BEG[12] ,
    \Tile_X8Y13_SS4BEG[11] ,
    \Tile_X8Y13_SS4BEG[10] ,
    \Tile_X8Y13_SS4BEG[9] ,
    \Tile_X8Y13_SS4BEG[8] ,
    \Tile_X8Y13_SS4BEG[7] ,
    \Tile_X8Y13_SS4BEG[6] ,
    \Tile_X8Y13_SS4BEG[5] ,
    \Tile_X8Y13_SS4BEG[4] ,
    \Tile_X8Y13_SS4BEG[3] ,
    \Tile_X8Y13_SS4BEG[2] ,
    \Tile_X8Y13_SS4BEG[1] ,
    \Tile_X8Y13_SS4BEG[0] }),
    .W1BEG({\Tile_X8Y14_W1BEG[3] ,
    \Tile_X8Y14_W1BEG[2] ,
    \Tile_X8Y14_W1BEG[1] ,
    \Tile_X8Y14_W1BEG[0] }),
    .W1END({\Tile_X9Y14_W1BEG[3] ,
    \Tile_X9Y14_W1BEG[2] ,
    \Tile_X9Y14_W1BEG[1] ,
    \Tile_X9Y14_W1BEG[0] }),
    .W2BEG({\Tile_X8Y14_W2BEG[7] ,
    \Tile_X8Y14_W2BEG[6] ,
    \Tile_X8Y14_W2BEG[5] ,
    \Tile_X8Y14_W2BEG[4] ,
    \Tile_X8Y14_W2BEG[3] ,
    \Tile_X8Y14_W2BEG[2] ,
    \Tile_X8Y14_W2BEG[1] ,
    \Tile_X8Y14_W2BEG[0] }),
    .W2BEGb({\Tile_X8Y14_W2BEGb[7] ,
    \Tile_X8Y14_W2BEGb[6] ,
    \Tile_X8Y14_W2BEGb[5] ,
    \Tile_X8Y14_W2BEGb[4] ,
    \Tile_X8Y14_W2BEGb[3] ,
    \Tile_X8Y14_W2BEGb[2] ,
    \Tile_X8Y14_W2BEGb[1] ,
    \Tile_X8Y14_W2BEGb[0] }),
    .W2END({\Tile_X9Y14_W2BEGb[7] ,
    \Tile_X9Y14_W2BEGb[6] ,
    \Tile_X9Y14_W2BEGb[5] ,
    \Tile_X9Y14_W2BEGb[4] ,
    \Tile_X9Y14_W2BEGb[3] ,
    \Tile_X9Y14_W2BEGb[2] ,
    \Tile_X9Y14_W2BEGb[1] ,
    \Tile_X9Y14_W2BEGb[0] }),
    .W2MID({\Tile_X9Y14_W2BEG[7] ,
    \Tile_X9Y14_W2BEG[6] ,
    \Tile_X9Y14_W2BEG[5] ,
    \Tile_X9Y14_W2BEG[4] ,
    \Tile_X9Y14_W2BEG[3] ,
    \Tile_X9Y14_W2BEG[2] ,
    \Tile_X9Y14_W2BEG[1] ,
    \Tile_X9Y14_W2BEG[0] }),
    .W6BEG({\Tile_X8Y14_W6BEG[11] ,
    \Tile_X8Y14_W6BEG[10] ,
    \Tile_X8Y14_W6BEG[9] ,
    \Tile_X8Y14_W6BEG[8] ,
    \Tile_X8Y14_W6BEG[7] ,
    \Tile_X8Y14_W6BEG[6] ,
    \Tile_X8Y14_W6BEG[5] ,
    \Tile_X8Y14_W6BEG[4] ,
    \Tile_X8Y14_W6BEG[3] ,
    \Tile_X8Y14_W6BEG[2] ,
    \Tile_X8Y14_W6BEG[1] ,
    \Tile_X8Y14_W6BEG[0] }),
    .W6END({\Tile_X9Y14_W6BEG[11] ,
    \Tile_X9Y14_W6BEG[10] ,
    \Tile_X9Y14_W6BEG[9] ,
    \Tile_X9Y14_W6BEG[8] ,
    \Tile_X9Y14_W6BEG[7] ,
    \Tile_X9Y14_W6BEG[6] ,
    \Tile_X9Y14_W6BEG[5] ,
    \Tile_X9Y14_W6BEG[4] ,
    \Tile_X9Y14_W6BEG[3] ,
    \Tile_X9Y14_W6BEG[2] ,
    \Tile_X9Y14_W6BEG[1] ,
    \Tile_X9Y14_W6BEG[0] }),
    .WW4BEG({\Tile_X8Y14_WW4BEG[15] ,
    \Tile_X8Y14_WW4BEG[14] ,
    \Tile_X8Y14_WW4BEG[13] ,
    \Tile_X8Y14_WW4BEG[12] ,
    \Tile_X8Y14_WW4BEG[11] ,
    \Tile_X8Y14_WW4BEG[10] ,
    \Tile_X8Y14_WW4BEG[9] ,
    \Tile_X8Y14_WW4BEG[8] ,
    \Tile_X8Y14_WW4BEG[7] ,
    \Tile_X8Y14_WW4BEG[6] ,
    \Tile_X8Y14_WW4BEG[5] ,
    \Tile_X8Y14_WW4BEG[4] ,
    \Tile_X8Y14_WW4BEG[3] ,
    \Tile_X8Y14_WW4BEG[2] ,
    \Tile_X8Y14_WW4BEG[1] ,
    \Tile_X8Y14_WW4BEG[0] }),
    .WW4END({\Tile_X9Y14_WW4BEG[15] ,
    \Tile_X9Y14_WW4BEG[14] ,
    \Tile_X9Y14_WW4BEG[13] ,
    \Tile_X9Y14_WW4BEG[12] ,
    \Tile_X9Y14_WW4BEG[11] ,
    \Tile_X9Y14_WW4BEG[10] ,
    \Tile_X9Y14_WW4BEG[9] ,
    \Tile_X9Y14_WW4BEG[8] ,
    \Tile_X9Y14_WW4BEG[7] ,
    \Tile_X9Y14_WW4BEG[6] ,
    \Tile_X9Y14_WW4BEG[5] ,
    \Tile_X9Y14_WW4BEG[4] ,
    \Tile_X9Y14_WW4BEG[3] ,
    \Tile_X9Y14_WW4BEG[2] ,
    \Tile_X9Y14_WW4BEG[1] ,
    \Tile_X9Y14_WW4BEG[0] }));
 S_CPU_IF Tile_X8Y15_S_CPU_IF (.Co(Tile_X8Y15_Co),
    .I_top0(Tile_X8Y15_I_top0),
    .I_top1(Tile_X8Y15_I_top1),
    .I_top10(Tile_X8Y15_I_top10),
    .I_top11(Tile_X8Y15_I_top11),
    .I_top12(Tile_X8Y15_I_top12),
    .I_top13(Tile_X8Y15_I_top13),
    .I_top14(Tile_X8Y15_I_top14),
    .I_top15(Tile_X8Y15_I_top15),
    .I_top2(Tile_X8Y15_I_top2),
    .I_top3(Tile_X8Y15_I_top3),
    .I_top4(Tile_X8Y15_I_top4),
    .I_top5(Tile_X8Y15_I_top5),
    .I_top6(Tile_X8Y15_I_top6),
    .I_top7(Tile_X8Y15_I_top7),
    .I_top8(Tile_X8Y15_I_top8),
    .I_top9(Tile_X8Y15_I_top9),
    .O_top0(Tile_X8Y15_O_top0),
    .O_top1(Tile_X8Y15_O_top1),
    .O_top10(Tile_X8Y15_O_top10),
    .O_top11(Tile_X8Y15_O_top11),
    .O_top12(Tile_X8Y15_O_top12),
    .O_top13(Tile_X8Y15_O_top13),
    .O_top14(Tile_X8Y15_O_top14),
    .O_top15(Tile_X8Y15_O_top15),
    .O_top2(Tile_X8Y15_O_top2),
    .O_top3(Tile_X8Y15_O_top3),
    .O_top4(Tile_X8Y15_O_top4),
    .O_top5(Tile_X8Y15_O_top5),
    .O_top6(Tile_X8Y15_O_top6),
    .O_top7(Tile_X8Y15_O_top7),
    .O_top8(Tile_X8Y15_O_top8),
    .O_top9(Tile_X8Y15_O_top9),
    .UserCLK(UserCLK),
    .UserCLKo(Tile_X8Y15_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .FrameData({\Tile_X7Y15_FrameData_O[31] ,
    \Tile_X7Y15_FrameData_O[30] ,
    \Tile_X7Y15_FrameData_O[29] ,
    \Tile_X7Y15_FrameData_O[28] ,
    \Tile_X7Y15_FrameData_O[27] ,
    \Tile_X7Y15_FrameData_O[26] ,
    \Tile_X7Y15_FrameData_O[25] ,
    \Tile_X7Y15_FrameData_O[24] ,
    \Tile_X7Y15_FrameData_O[23] ,
    \Tile_X7Y15_FrameData_O[22] ,
    \Tile_X7Y15_FrameData_O[21] ,
    \Tile_X7Y15_FrameData_O[20] ,
    \Tile_X7Y15_FrameData_O[19] ,
    \Tile_X7Y15_FrameData_O[18] ,
    \Tile_X7Y15_FrameData_O[17] ,
    \Tile_X7Y15_FrameData_O[16] ,
    \Tile_X7Y15_FrameData_O[15] ,
    \Tile_X7Y15_FrameData_O[14] ,
    \Tile_X7Y15_FrameData_O[13] ,
    \Tile_X7Y15_FrameData_O[12] ,
    \Tile_X7Y15_FrameData_O[11] ,
    \Tile_X7Y15_FrameData_O[10] ,
    \Tile_X7Y15_FrameData_O[9] ,
    \Tile_X7Y15_FrameData_O[8] ,
    \Tile_X7Y15_FrameData_O[7] ,
    \Tile_X7Y15_FrameData_O[6] ,
    \Tile_X7Y15_FrameData_O[5] ,
    \Tile_X7Y15_FrameData_O[4] ,
    \Tile_X7Y15_FrameData_O[3] ,
    \Tile_X7Y15_FrameData_O[2] ,
    \Tile_X7Y15_FrameData_O[1] ,
    \Tile_X7Y15_FrameData_O[0] }),
    .FrameData_O({\Tile_X8Y15_FrameData_O[31] ,
    \Tile_X8Y15_FrameData_O[30] ,
    \Tile_X8Y15_FrameData_O[29] ,
    \Tile_X8Y15_FrameData_O[28] ,
    \Tile_X8Y15_FrameData_O[27] ,
    \Tile_X8Y15_FrameData_O[26] ,
    \Tile_X8Y15_FrameData_O[25] ,
    \Tile_X8Y15_FrameData_O[24] ,
    \Tile_X8Y15_FrameData_O[23] ,
    \Tile_X8Y15_FrameData_O[22] ,
    \Tile_X8Y15_FrameData_O[21] ,
    \Tile_X8Y15_FrameData_O[20] ,
    \Tile_X8Y15_FrameData_O[19] ,
    \Tile_X8Y15_FrameData_O[18] ,
    \Tile_X8Y15_FrameData_O[17] ,
    \Tile_X8Y15_FrameData_O[16] ,
    \Tile_X8Y15_FrameData_O[15] ,
    \Tile_X8Y15_FrameData_O[14] ,
    \Tile_X8Y15_FrameData_O[13] ,
    \Tile_X8Y15_FrameData_O[12] ,
    \Tile_X8Y15_FrameData_O[11] ,
    \Tile_X8Y15_FrameData_O[10] ,
    \Tile_X8Y15_FrameData_O[9] ,
    \Tile_X8Y15_FrameData_O[8] ,
    \Tile_X8Y15_FrameData_O[7] ,
    \Tile_X8Y15_FrameData_O[6] ,
    \Tile_X8Y15_FrameData_O[5] ,
    \Tile_X8Y15_FrameData_O[4] ,
    \Tile_X8Y15_FrameData_O[3] ,
    \Tile_X8Y15_FrameData_O[2] ,
    \Tile_X8Y15_FrameData_O[1] ,
    \Tile_X8Y15_FrameData_O[0] }),
    .FrameStrobe({FrameStrobe[179],
    FrameStrobe[178],
    FrameStrobe[177],
    FrameStrobe[176],
    FrameStrobe[175],
    FrameStrobe[174],
    FrameStrobe[173],
    FrameStrobe[172],
    FrameStrobe[171],
    FrameStrobe[170],
    FrameStrobe[169],
    FrameStrobe[168],
    FrameStrobe[167],
    FrameStrobe[166],
    FrameStrobe[165],
    FrameStrobe[164],
    FrameStrobe[163],
    FrameStrobe[162],
    FrameStrobe[161],
    FrameStrobe[160]}),
    .FrameStrobe_O({\Tile_X8Y15_FrameStrobe_O[19] ,
    \Tile_X8Y15_FrameStrobe_O[18] ,
    \Tile_X8Y15_FrameStrobe_O[17] ,
    \Tile_X8Y15_FrameStrobe_O[16] ,
    \Tile_X8Y15_FrameStrobe_O[15] ,
    \Tile_X8Y15_FrameStrobe_O[14] ,
    \Tile_X8Y15_FrameStrobe_O[13] ,
    \Tile_X8Y15_FrameStrobe_O[12] ,
    \Tile_X8Y15_FrameStrobe_O[11] ,
    \Tile_X8Y15_FrameStrobe_O[10] ,
    \Tile_X8Y15_FrameStrobe_O[9] ,
    \Tile_X8Y15_FrameStrobe_O[8] ,
    \Tile_X8Y15_FrameStrobe_O[7] ,
    \Tile_X8Y15_FrameStrobe_O[6] ,
    \Tile_X8Y15_FrameStrobe_O[5] ,
    \Tile_X8Y15_FrameStrobe_O[4] ,
    \Tile_X8Y15_FrameStrobe_O[3] ,
    \Tile_X8Y15_FrameStrobe_O[2] ,
    \Tile_X8Y15_FrameStrobe_O[1] ,
    \Tile_X8Y15_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X8Y15_N1BEG[3] ,
    \Tile_X8Y15_N1BEG[2] ,
    \Tile_X8Y15_N1BEG[1] ,
    \Tile_X8Y15_N1BEG[0] }),
    .N2BEG({\Tile_X8Y15_N2BEG[7] ,
    \Tile_X8Y15_N2BEG[6] ,
    \Tile_X8Y15_N2BEG[5] ,
    \Tile_X8Y15_N2BEG[4] ,
    \Tile_X8Y15_N2BEG[3] ,
    \Tile_X8Y15_N2BEG[2] ,
    \Tile_X8Y15_N2BEG[1] ,
    \Tile_X8Y15_N2BEG[0] }),
    .N2BEGb({\Tile_X8Y15_N2BEGb[7] ,
    \Tile_X8Y15_N2BEGb[6] ,
    \Tile_X8Y15_N2BEGb[5] ,
    \Tile_X8Y15_N2BEGb[4] ,
    \Tile_X8Y15_N2BEGb[3] ,
    \Tile_X8Y15_N2BEGb[2] ,
    \Tile_X8Y15_N2BEGb[1] ,
    \Tile_X8Y15_N2BEGb[0] }),
    .N4BEG({\Tile_X8Y15_N4BEG[15] ,
    \Tile_X8Y15_N4BEG[14] ,
    \Tile_X8Y15_N4BEG[13] ,
    \Tile_X8Y15_N4BEG[12] ,
    \Tile_X8Y15_N4BEG[11] ,
    \Tile_X8Y15_N4BEG[10] ,
    \Tile_X8Y15_N4BEG[9] ,
    \Tile_X8Y15_N4BEG[8] ,
    \Tile_X8Y15_N4BEG[7] ,
    \Tile_X8Y15_N4BEG[6] ,
    \Tile_X8Y15_N4BEG[5] ,
    \Tile_X8Y15_N4BEG[4] ,
    \Tile_X8Y15_N4BEG[3] ,
    \Tile_X8Y15_N4BEG[2] ,
    \Tile_X8Y15_N4BEG[1] ,
    \Tile_X8Y15_N4BEG[0] }),
    .NN4BEG({\Tile_X8Y15_NN4BEG[15] ,
    \Tile_X8Y15_NN4BEG[14] ,
    \Tile_X8Y15_NN4BEG[13] ,
    \Tile_X8Y15_NN4BEG[12] ,
    \Tile_X8Y15_NN4BEG[11] ,
    \Tile_X8Y15_NN4BEG[10] ,
    \Tile_X8Y15_NN4BEG[9] ,
    \Tile_X8Y15_NN4BEG[8] ,
    \Tile_X8Y15_NN4BEG[7] ,
    \Tile_X8Y15_NN4BEG[6] ,
    \Tile_X8Y15_NN4BEG[5] ,
    \Tile_X8Y15_NN4BEG[4] ,
    \Tile_X8Y15_NN4BEG[3] ,
    \Tile_X8Y15_NN4BEG[2] ,
    \Tile_X8Y15_NN4BEG[1] ,
    \Tile_X8Y15_NN4BEG[0] }),
    .S1END({\Tile_X8Y14_S1BEG[3] ,
    \Tile_X8Y14_S1BEG[2] ,
    \Tile_X8Y14_S1BEG[1] ,
    \Tile_X8Y14_S1BEG[0] }),
    .S2END({\Tile_X8Y14_S2BEGb[7] ,
    \Tile_X8Y14_S2BEGb[6] ,
    \Tile_X8Y14_S2BEGb[5] ,
    \Tile_X8Y14_S2BEGb[4] ,
    \Tile_X8Y14_S2BEGb[3] ,
    \Tile_X8Y14_S2BEGb[2] ,
    \Tile_X8Y14_S2BEGb[1] ,
    \Tile_X8Y14_S2BEGb[0] }),
    .S2MID({\Tile_X8Y14_S2BEG[7] ,
    \Tile_X8Y14_S2BEG[6] ,
    \Tile_X8Y14_S2BEG[5] ,
    \Tile_X8Y14_S2BEG[4] ,
    \Tile_X8Y14_S2BEG[3] ,
    \Tile_X8Y14_S2BEG[2] ,
    \Tile_X8Y14_S2BEG[1] ,
    \Tile_X8Y14_S2BEG[0] }),
    .S4END({\Tile_X8Y14_S4BEG[15] ,
    \Tile_X8Y14_S4BEG[14] ,
    \Tile_X8Y14_S4BEG[13] ,
    \Tile_X8Y14_S4BEG[12] ,
    \Tile_X8Y14_S4BEG[11] ,
    \Tile_X8Y14_S4BEG[10] ,
    \Tile_X8Y14_S4BEG[9] ,
    \Tile_X8Y14_S4BEG[8] ,
    \Tile_X8Y14_S4BEG[7] ,
    \Tile_X8Y14_S4BEG[6] ,
    \Tile_X8Y14_S4BEG[5] ,
    \Tile_X8Y14_S4BEG[4] ,
    \Tile_X8Y14_S4BEG[3] ,
    \Tile_X8Y14_S4BEG[2] ,
    \Tile_X8Y14_S4BEG[1] ,
    \Tile_X8Y14_S4BEG[0] }),
    .SS4END({\Tile_X8Y14_SS4BEG[15] ,
    \Tile_X8Y14_SS4BEG[14] ,
    \Tile_X8Y14_SS4BEG[13] ,
    \Tile_X8Y14_SS4BEG[12] ,
    \Tile_X8Y14_SS4BEG[11] ,
    \Tile_X8Y14_SS4BEG[10] ,
    \Tile_X8Y14_SS4BEG[9] ,
    \Tile_X8Y14_SS4BEG[8] ,
    \Tile_X8Y14_SS4BEG[7] ,
    \Tile_X8Y14_SS4BEG[6] ,
    \Tile_X8Y14_SS4BEG[5] ,
    \Tile_X8Y14_SS4BEG[4] ,
    \Tile_X8Y14_SS4BEG[3] ,
    \Tile_X8Y14_SS4BEG[2] ,
    \Tile_X8Y14_SS4BEG[1] ,
    \Tile_X8Y14_SS4BEG[0] }));
 LUT4AB Tile_X8Y1_LUT4AB (.Ci(Tile_X8Y2_Co),
    .Co(Tile_X8Y1_Co),
    .UserCLK(Tile_X8Y2_UserCLKo),
    .UserCLKo(Tile_X8Y1_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X8Y1_E1BEG[3] ,
    \Tile_X8Y1_E1BEG[2] ,
    \Tile_X8Y1_E1BEG[1] ,
    \Tile_X8Y1_E1BEG[0] }),
    .E1END({\Tile_X7Y1_E1BEG[3] ,
    \Tile_X7Y1_E1BEG[2] ,
    \Tile_X7Y1_E1BEG[1] ,
    \Tile_X7Y1_E1BEG[0] }),
    .E2BEG({\Tile_X8Y1_E2BEG[7] ,
    \Tile_X8Y1_E2BEG[6] ,
    \Tile_X8Y1_E2BEG[5] ,
    \Tile_X8Y1_E2BEG[4] ,
    \Tile_X8Y1_E2BEG[3] ,
    \Tile_X8Y1_E2BEG[2] ,
    \Tile_X8Y1_E2BEG[1] ,
    \Tile_X8Y1_E2BEG[0] }),
    .E2BEGb({\Tile_X8Y1_E2BEGb[7] ,
    \Tile_X8Y1_E2BEGb[6] ,
    \Tile_X8Y1_E2BEGb[5] ,
    \Tile_X8Y1_E2BEGb[4] ,
    \Tile_X8Y1_E2BEGb[3] ,
    \Tile_X8Y1_E2BEGb[2] ,
    \Tile_X8Y1_E2BEGb[1] ,
    \Tile_X8Y1_E2BEGb[0] }),
    .E2END({\Tile_X7Y1_E2BEGb[7] ,
    \Tile_X7Y1_E2BEGb[6] ,
    \Tile_X7Y1_E2BEGb[5] ,
    \Tile_X7Y1_E2BEGb[4] ,
    \Tile_X7Y1_E2BEGb[3] ,
    \Tile_X7Y1_E2BEGb[2] ,
    \Tile_X7Y1_E2BEGb[1] ,
    \Tile_X7Y1_E2BEGb[0] }),
    .E2MID({\Tile_X7Y1_E2BEG[7] ,
    \Tile_X7Y1_E2BEG[6] ,
    \Tile_X7Y1_E2BEG[5] ,
    \Tile_X7Y1_E2BEG[4] ,
    \Tile_X7Y1_E2BEG[3] ,
    \Tile_X7Y1_E2BEG[2] ,
    \Tile_X7Y1_E2BEG[1] ,
    \Tile_X7Y1_E2BEG[0] }),
    .E6BEG({\Tile_X8Y1_E6BEG[11] ,
    \Tile_X8Y1_E6BEG[10] ,
    \Tile_X8Y1_E6BEG[9] ,
    \Tile_X8Y1_E6BEG[8] ,
    \Tile_X8Y1_E6BEG[7] ,
    \Tile_X8Y1_E6BEG[6] ,
    \Tile_X8Y1_E6BEG[5] ,
    \Tile_X8Y1_E6BEG[4] ,
    \Tile_X8Y1_E6BEG[3] ,
    \Tile_X8Y1_E6BEG[2] ,
    \Tile_X8Y1_E6BEG[1] ,
    \Tile_X8Y1_E6BEG[0] }),
    .E6END({\Tile_X7Y1_E6BEG[11] ,
    \Tile_X7Y1_E6BEG[10] ,
    \Tile_X7Y1_E6BEG[9] ,
    \Tile_X7Y1_E6BEG[8] ,
    \Tile_X7Y1_E6BEG[7] ,
    \Tile_X7Y1_E6BEG[6] ,
    \Tile_X7Y1_E6BEG[5] ,
    \Tile_X7Y1_E6BEG[4] ,
    \Tile_X7Y1_E6BEG[3] ,
    \Tile_X7Y1_E6BEG[2] ,
    \Tile_X7Y1_E6BEG[1] ,
    \Tile_X7Y1_E6BEG[0] }),
    .EE4BEG({\Tile_X8Y1_EE4BEG[15] ,
    \Tile_X8Y1_EE4BEG[14] ,
    \Tile_X8Y1_EE4BEG[13] ,
    \Tile_X8Y1_EE4BEG[12] ,
    \Tile_X8Y1_EE4BEG[11] ,
    \Tile_X8Y1_EE4BEG[10] ,
    \Tile_X8Y1_EE4BEG[9] ,
    \Tile_X8Y1_EE4BEG[8] ,
    \Tile_X8Y1_EE4BEG[7] ,
    \Tile_X8Y1_EE4BEG[6] ,
    \Tile_X8Y1_EE4BEG[5] ,
    \Tile_X8Y1_EE4BEG[4] ,
    \Tile_X8Y1_EE4BEG[3] ,
    \Tile_X8Y1_EE4BEG[2] ,
    \Tile_X8Y1_EE4BEG[1] ,
    \Tile_X8Y1_EE4BEG[0] }),
    .EE4END({\Tile_X7Y1_EE4BEG[15] ,
    \Tile_X7Y1_EE4BEG[14] ,
    \Tile_X7Y1_EE4BEG[13] ,
    \Tile_X7Y1_EE4BEG[12] ,
    \Tile_X7Y1_EE4BEG[11] ,
    \Tile_X7Y1_EE4BEG[10] ,
    \Tile_X7Y1_EE4BEG[9] ,
    \Tile_X7Y1_EE4BEG[8] ,
    \Tile_X7Y1_EE4BEG[7] ,
    \Tile_X7Y1_EE4BEG[6] ,
    \Tile_X7Y1_EE4BEG[5] ,
    \Tile_X7Y1_EE4BEG[4] ,
    \Tile_X7Y1_EE4BEG[3] ,
    \Tile_X7Y1_EE4BEG[2] ,
    \Tile_X7Y1_EE4BEG[1] ,
    \Tile_X7Y1_EE4BEG[0] }),
    .FrameData({\Tile_X7Y1_FrameData_O[31] ,
    \Tile_X7Y1_FrameData_O[30] ,
    \Tile_X7Y1_FrameData_O[29] ,
    \Tile_X7Y1_FrameData_O[28] ,
    \Tile_X7Y1_FrameData_O[27] ,
    \Tile_X7Y1_FrameData_O[26] ,
    \Tile_X7Y1_FrameData_O[25] ,
    \Tile_X7Y1_FrameData_O[24] ,
    \Tile_X7Y1_FrameData_O[23] ,
    \Tile_X7Y1_FrameData_O[22] ,
    \Tile_X7Y1_FrameData_O[21] ,
    \Tile_X7Y1_FrameData_O[20] ,
    \Tile_X7Y1_FrameData_O[19] ,
    \Tile_X7Y1_FrameData_O[18] ,
    \Tile_X7Y1_FrameData_O[17] ,
    \Tile_X7Y1_FrameData_O[16] ,
    \Tile_X7Y1_FrameData_O[15] ,
    \Tile_X7Y1_FrameData_O[14] ,
    \Tile_X7Y1_FrameData_O[13] ,
    \Tile_X7Y1_FrameData_O[12] ,
    \Tile_X7Y1_FrameData_O[11] ,
    \Tile_X7Y1_FrameData_O[10] ,
    \Tile_X7Y1_FrameData_O[9] ,
    \Tile_X7Y1_FrameData_O[8] ,
    \Tile_X7Y1_FrameData_O[7] ,
    \Tile_X7Y1_FrameData_O[6] ,
    \Tile_X7Y1_FrameData_O[5] ,
    \Tile_X7Y1_FrameData_O[4] ,
    \Tile_X7Y1_FrameData_O[3] ,
    \Tile_X7Y1_FrameData_O[2] ,
    \Tile_X7Y1_FrameData_O[1] ,
    \Tile_X7Y1_FrameData_O[0] }),
    .FrameData_O({\Tile_X8Y1_FrameData_O[31] ,
    \Tile_X8Y1_FrameData_O[30] ,
    \Tile_X8Y1_FrameData_O[29] ,
    \Tile_X8Y1_FrameData_O[28] ,
    \Tile_X8Y1_FrameData_O[27] ,
    \Tile_X8Y1_FrameData_O[26] ,
    \Tile_X8Y1_FrameData_O[25] ,
    \Tile_X8Y1_FrameData_O[24] ,
    \Tile_X8Y1_FrameData_O[23] ,
    \Tile_X8Y1_FrameData_O[22] ,
    \Tile_X8Y1_FrameData_O[21] ,
    \Tile_X8Y1_FrameData_O[20] ,
    \Tile_X8Y1_FrameData_O[19] ,
    \Tile_X8Y1_FrameData_O[18] ,
    \Tile_X8Y1_FrameData_O[17] ,
    \Tile_X8Y1_FrameData_O[16] ,
    \Tile_X8Y1_FrameData_O[15] ,
    \Tile_X8Y1_FrameData_O[14] ,
    \Tile_X8Y1_FrameData_O[13] ,
    \Tile_X8Y1_FrameData_O[12] ,
    \Tile_X8Y1_FrameData_O[11] ,
    \Tile_X8Y1_FrameData_O[10] ,
    \Tile_X8Y1_FrameData_O[9] ,
    \Tile_X8Y1_FrameData_O[8] ,
    \Tile_X8Y1_FrameData_O[7] ,
    \Tile_X8Y1_FrameData_O[6] ,
    \Tile_X8Y1_FrameData_O[5] ,
    \Tile_X8Y1_FrameData_O[4] ,
    \Tile_X8Y1_FrameData_O[3] ,
    \Tile_X8Y1_FrameData_O[2] ,
    \Tile_X8Y1_FrameData_O[1] ,
    \Tile_X8Y1_FrameData_O[0] }),
    .FrameStrobe({\Tile_X8Y2_FrameStrobe_O[19] ,
    \Tile_X8Y2_FrameStrobe_O[18] ,
    \Tile_X8Y2_FrameStrobe_O[17] ,
    \Tile_X8Y2_FrameStrobe_O[16] ,
    \Tile_X8Y2_FrameStrobe_O[15] ,
    \Tile_X8Y2_FrameStrobe_O[14] ,
    \Tile_X8Y2_FrameStrobe_O[13] ,
    \Tile_X8Y2_FrameStrobe_O[12] ,
    \Tile_X8Y2_FrameStrobe_O[11] ,
    \Tile_X8Y2_FrameStrobe_O[10] ,
    \Tile_X8Y2_FrameStrobe_O[9] ,
    \Tile_X8Y2_FrameStrobe_O[8] ,
    \Tile_X8Y2_FrameStrobe_O[7] ,
    \Tile_X8Y2_FrameStrobe_O[6] ,
    \Tile_X8Y2_FrameStrobe_O[5] ,
    \Tile_X8Y2_FrameStrobe_O[4] ,
    \Tile_X8Y2_FrameStrobe_O[3] ,
    \Tile_X8Y2_FrameStrobe_O[2] ,
    \Tile_X8Y2_FrameStrobe_O[1] ,
    \Tile_X8Y2_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X8Y1_FrameStrobe_O[19] ,
    \Tile_X8Y1_FrameStrobe_O[18] ,
    \Tile_X8Y1_FrameStrobe_O[17] ,
    \Tile_X8Y1_FrameStrobe_O[16] ,
    \Tile_X8Y1_FrameStrobe_O[15] ,
    \Tile_X8Y1_FrameStrobe_O[14] ,
    \Tile_X8Y1_FrameStrobe_O[13] ,
    \Tile_X8Y1_FrameStrobe_O[12] ,
    \Tile_X8Y1_FrameStrobe_O[11] ,
    \Tile_X8Y1_FrameStrobe_O[10] ,
    \Tile_X8Y1_FrameStrobe_O[9] ,
    \Tile_X8Y1_FrameStrobe_O[8] ,
    \Tile_X8Y1_FrameStrobe_O[7] ,
    \Tile_X8Y1_FrameStrobe_O[6] ,
    \Tile_X8Y1_FrameStrobe_O[5] ,
    \Tile_X8Y1_FrameStrobe_O[4] ,
    \Tile_X8Y1_FrameStrobe_O[3] ,
    \Tile_X8Y1_FrameStrobe_O[2] ,
    \Tile_X8Y1_FrameStrobe_O[1] ,
    \Tile_X8Y1_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X8Y1_N1BEG[3] ,
    \Tile_X8Y1_N1BEG[2] ,
    \Tile_X8Y1_N1BEG[1] ,
    \Tile_X8Y1_N1BEG[0] }),
    .N1END({\Tile_X8Y2_N1BEG[3] ,
    \Tile_X8Y2_N1BEG[2] ,
    \Tile_X8Y2_N1BEG[1] ,
    \Tile_X8Y2_N1BEG[0] }),
    .N2BEG({\Tile_X8Y1_N2BEG[7] ,
    \Tile_X8Y1_N2BEG[6] ,
    \Tile_X8Y1_N2BEG[5] ,
    \Tile_X8Y1_N2BEG[4] ,
    \Tile_X8Y1_N2BEG[3] ,
    \Tile_X8Y1_N2BEG[2] ,
    \Tile_X8Y1_N2BEG[1] ,
    \Tile_X8Y1_N2BEG[0] }),
    .N2BEGb({\Tile_X8Y1_N2BEGb[7] ,
    \Tile_X8Y1_N2BEGb[6] ,
    \Tile_X8Y1_N2BEGb[5] ,
    \Tile_X8Y1_N2BEGb[4] ,
    \Tile_X8Y1_N2BEGb[3] ,
    \Tile_X8Y1_N2BEGb[2] ,
    \Tile_X8Y1_N2BEGb[1] ,
    \Tile_X8Y1_N2BEGb[0] }),
    .N2END({\Tile_X8Y2_N2BEGb[7] ,
    \Tile_X8Y2_N2BEGb[6] ,
    \Tile_X8Y2_N2BEGb[5] ,
    \Tile_X8Y2_N2BEGb[4] ,
    \Tile_X8Y2_N2BEGb[3] ,
    \Tile_X8Y2_N2BEGb[2] ,
    \Tile_X8Y2_N2BEGb[1] ,
    \Tile_X8Y2_N2BEGb[0] }),
    .N2MID({\Tile_X8Y2_N2BEG[7] ,
    \Tile_X8Y2_N2BEG[6] ,
    \Tile_X8Y2_N2BEG[5] ,
    \Tile_X8Y2_N2BEG[4] ,
    \Tile_X8Y2_N2BEG[3] ,
    \Tile_X8Y2_N2BEG[2] ,
    \Tile_X8Y2_N2BEG[1] ,
    \Tile_X8Y2_N2BEG[0] }),
    .N4BEG({\Tile_X8Y1_N4BEG[15] ,
    \Tile_X8Y1_N4BEG[14] ,
    \Tile_X8Y1_N4BEG[13] ,
    \Tile_X8Y1_N4BEG[12] ,
    \Tile_X8Y1_N4BEG[11] ,
    \Tile_X8Y1_N4BEG[10] ,
    \Tile_X8Y1_N4BEG[9] ,
    \Tile_X8Y1_N4BEG[8] ,
    \Tile_X8Y1_N4BEG[7] ,
    \Tile_X8Y1_N4BEG[6] ,
    \Tile_X8Y1_N4BEG[5] ,
    \Tile_X8Y1_N4BEG[4] ,
    \Tile_X8Y1_N4BEG[3] ,
    \Tile_X8Y1_N4BEG[2] ,
    \Tile_X8Y1_N4BEG[1] ,
    \Tile_X8Y1_N4BEG[0] }),
    .N4END({\Tile_X8Y2_N4BEG[15] ,
    \Tile_X8Y2_N4BEG[14] ,
    \Tile_X8Y2_N4BEG[13] ,
    \Tile_X8Y2_N4BEG[12] ,
    \Tile_X8Y2_N4BEG[11] ,
    \Tile_X8Y2_N4BEG[10] ,
    \Tile_X8Y2_N4BEG[9] ,
    \Tile_X8Y2_N4BEG[8] ,
    \Tile_X8Y2_N4BEG[7] ,
    \Tile_X8Y2_N4BEG[6] ,
    \Tile_X8Y2_N4BEG[5] ,
    \Tile_X8Y2_N4BEG[4] ,
    \Tile_X8Y2_N4BEG[3] ,
    \Tile_X8Y2_N4BEG[2] ,
    \Tile_X8Y2_N4BEG[1] ,
    \Tile_X8Y2_N4BEG[0] }),
    .NN4BEG({\Tile_X8Y1_NN4BEG[15] ,
    \Tile_X8Y1_NN4BEG[14] ,
    \Tile_X8Y1_NN4BEG[13] ,
    \Tile_X8Y1_NN4BEG[12] ,
    \Tile_X8Y1_NN4BEG[11] ,
    \Tile_X8Y1_NN4BEG[10] ,
    \Tile_X8Y1_NN4BEG[9] ,
    \Tile_X8Y1_NN4BEG[8] ,
    \Tile_X8Y1_NN4BEG[7] ,
    \Tile_X8Y1_NN4BEG[6] ,
    \Tile_X8Y1_NN4BEG[5] ,
    \Tile_X8Y1_NN4BEG[4] ,
    \Tile_X8Y1_NN4BEG[3] ,
    \Tile_X8Y1_NN4BEG[2] ,
    \Tile_X8Y1_NN4BEG[1] ,
    \Tile_X8Y1_NN4BEG[0] }),
    .NN4END({\Tile_X8Y2_NN4BEG[15] ,
    \Tile_X8Y2_NN4BEG[14] ,
    \Tile_X8Y2_NN4BEG[13] ,
    \Tile_X8Y2_NN4BEG[12] ,
    \Tile_X8Y2_NN4BEG[11] ,
    \Tile_X8Y2_NN4BEG[10] ,
    \Tile_X8Y2_NN4BEG[9] ,
    \Tile_X8Y2_NN4BEG[8] ,
    \Tile_X8Y2_NN4BEG[7] ,
    \Tile_X8Y2_NN4BEG[6] ,
    \Tile_X8Y2_NN4BEG[5] ,
    \Tile_X8Y2_NN4BEG[4] ,
    \Tile_X8Y2_NN4BEG[3] ,
    \Tile_X8Y2_NN4BEG[2] ,
    \Tile_X8Y2_NN4BEG[1] ,
    \Tile_X8Y2_NN4BEG[0] }),
    .S1BEG({\Tile_X8Y1_S1BEG[3] ,
    \Tile_X8Y1_S1BEG[2] ,
    \Tile_X8Y1_S1BEG[1] ,
    \Tile_X8Y1_S1BEG[0] }),
    .S1END({\Tile_X8Y0_S1BEG[3] ,
    \Tile_X8Y0_S1BEG[2] ,
    \Tile_X8Y0_S1BEG[1] ,
    \Tile_X8Y0_S1BEG[0] }),
    .S2BEG({\Tile_X8Y1_S2BEG[7] ,
    \Tile_X8Y1_S2BEG[6] ,
    \Tile_X8Y1_S2BEG[5] ,
    \Tile_X8Y1_S2BEG[4] ,
    \Tile_X8Y1_S2BEG[3] ,
    \Tile_X8Y1_S2BEG[2] ,
    \Tile_X8Y1_S2BEG[1] ,
    \Tile_X8Y1_S2BEG[0] }),
    .S2BEGb({\Tile_X8Y1_S2BEGb[7] ,
    \Tile_X8Y1_S2BEGb[6] ,
    \Tile_X8Y1_S2BEGb[5] ,
    \Tile_X8Y1_S2BEGb[4] ,
    \Tile_X8Y1_S2BEGb[3] ,
    \Tile_X8Y1_S2BEGb[2] ,
    \Tile_X8Y1_S2BEGb[1] ,
    \Tile_X8Y1_S2BEGb[0] }),
    .S2END({\Tile_X8Y0_S2BEGb[7] ,
    \Tile_X8Y0_S2BEGb[6] ,
    \Tile_X8Y0_S2BEGb[5] ,
    \Tile_X8Y0_S2BEGb[4] ,
    \Tile_X8Y0_S2BEGb[3] ,
    \Tile_X8Y0_S2BEGb[2] ,
    \Tile_X8Y0_S2BEGb[1] ,
    \Tile_X8Y0_S2BEGb[0] }),
    .S2MID({\Tile_X8Y0_S2BEG[7] ,
    \Tile_X8Y0_S2BEG[6] ,
    \Tile_X8Y0_S2BEG[5] ,
    \Tile_X8Y0_S2BEG[4] ,
    \Tile_X8Y0_S2BEG[3] ,
    \Tile_X8Y0_S2BEG[2] ,
    \Tile_X8Y0_S2BEG[1] ,
    \Tile_X8Y0_S2BEG[0] }),
    .S4BEG({\Tile_X8Y1_S4BEG[15] ,
    \Tile_X8Y1_S4BEG[14] ,
    \Tile_X8Y1_S4BEG[13] ,
    \Tile_X8Y1_S4BEG[12] ,
    \Tile_X8Y1_S4BEG[11] ,
    \Tile_X8Y1_S4BEG[10] ,
    \Tile_X8Y1_S4BEG[9] ,
    \Tile_X8Y1_S4BEG[8] ,
    \Tile_X8Y1_S4BEG[7] ,
    \Tile_X8Y1_S4BEG[6] ,
    \Tile_X8Y1_S4BEG[5] ,
    \Tile_X8Y1_S4BEG[4] ,
    \Tile_X8Y1_S4BEG[3] ,
    \Tile_X8Y1_S4BEG[2] ,
    \Tile_X8Y1_S4BEG[1] ,
    \Tile_X8Y1_S4BEG[0] }),
    .S4END({\Tile_X8Y0_S4BEG[15] ,
    \Tile_X8Y0_S4BEG[14] ,
    \Tile_X8Y0_S4BEG[13] ,
    \Tile_X8Y0_S4BEG[12] ,
    \Tile_X8Y0_S4BEG[11] ,
    \Tile_X8Y0_S4BEG[10] ,
    \Tile_X8Y0_S4BEG[9] ,
    \Tile_X8Y0_S4BEG[8] ,
    \Tile_X8Y0_S4BEG[7] ,
    \Tile_X8Y0_S4BEG[6] ,
    \Tile_X8Y0_S4BEG[5] ,
    \Tile_X8Y0_S4BEG[4] ,
    \Tile_X8Y0_S4BEG[3] ,
    \Tile_X8Y0_S4BEG[2] ,
    \Tile_X8Y0_S4BEG[1] ,
    \Tile_X8Y0_S4BEG[0] }),
    .SS4BEG({\Tile_X8Y1_SS4BEG[15] ,
    \Tile_X8Y1_SS4BEG[14] ,
    \Tile_X8Y1_SS4BEG[13] ,
    \Tile_X8Y1_SS4BEG[12] ,
    \Tile_X8Y1_SS4BEG[11] ,
    \Tile_X8Y1_SS4BEG[10] ,
    \Tile_X8Y1_SS4BEG[9] ,
    \Tile_X8Y1_SS4BEG[8] ,
    \Tile_X8Y1_SS4BEG[7] ,
    \Tile_X8Y1_SS4BEG[6] ,
    \Tile_X8Y1_SS4BEG[5] ,
    \Tile_X8Y1_SS4BEG[4] ,
    \Tile_X8Y1_SS4BEG[3] ,
    \Tile_X8Y1_SS4BEG[2] ,
    \Tile_X8Y1_SS4BEG[1] ,
    \Tile_X8Y1_SS4BEG[0] }),
    .SS4END({\Tile_X8Y0_SS4BEG[15] ,
    \Tile_X8Y0_SS4BEG[14] ,
    \Tile_X8Y0_SS4BEG[13] ,
    \Tile_X8Y0_SS4BEG[12] ,
    \Tile_X8Y0_SS4BEG[11] ,
    \Tile_X8Y0_SS4BEG[10] ,
    \Tile_X8Y0_SS4BEG[9] ,
    \Tile_X8Y0_SS4BEG[8] ,
    \Tile_X8Y0_SS4BEG[7] ,
    \Tile_X8Y0_SS4BEG[6] ,
    \Tile_X8Y0_SS4BEG[5] ,
    \Tile_X8Y0_SS4BEG[4] ,
    \Tile_X8Y0_SS4BEG[3] ,
    \Tile_X8Y0_SS4BEG[2] ,
    \Tile_X8Y0_SS4BEG[1] ,
    \Tile_X8Y0_SS4BEG[0] }),
    .W1BEG({\Tile_X8Y1_W1BEG[3] ,
    \Tile_X8Y1_W1BEG[2] ,
    \Tile_X8Y1_W1BEG[1] ,
    \Tile_X8Y1_W1BEG[0] }),
    .W1END({\Tile_X9Y1_W1BEG[3] ,
    \Tile_X9Y1_W1BEG[2] ,
    \Tile_X9Y1_W1BEG[1] ,
    \Tile_X9Y1_W1BEG[0] }),
    .W2BEG({\Tile_X8Y1_W2BEG[7] ,
    \Tile_X8Y1_W2BEG[6] ,
    \Tile_X8Y1_W2BEG[5] ,
    \Tile_X8Y1_W2BEG[4] ,
    \Tile_X8Y1_W2BEG[3] ,
    \Tile_X8Y1_W2BEG[2] ,
    \Tile_X8Y1_W2BEG[1] ,
    \Tile_X8Y1_W2BEG[0] }),
    .W2BEGb({\Tile_X8Y1_W2BEGb[7] ,
    \Tile_X8Y1_W2BEGb[6] ,
    \Tile_X8Y1_W2BEGb[5] ,
    \Tile_X8Y1_W2BEGb[4] ,
    \Tile_X8Y1_W2BEGb[3] ,
    \Tile_X8Y1_W2BEGb[2] ,
    \Tile_X8Y1_W2BEGb[1] ,
    \Tile_X8Y1_W2BEGb[0] }),
    .W2END({\Tile_X9Y1_W2BEGb[7] ,
    \Tile_X9Y1_W2BEGb[6] ,
    \Tile_X9Y1_W2BEGb[5] ,
    \Tile_X9Y1_W2BEGb[4] ,
    \Tile_X9Y1_W2BEGb[3] ,
    \Tile_X9Y1_W2BEGb[2] ,
    \Tile_X9Y1_W2BEGb[1] ,
    \Tile_X9Y1_W2BEGb[0] }),
    .W2MID({\Tile_X9Y1_W2BEG[7] ,
    \Tile_X9Y1_W2BEG[6] ,
    \Tile_X9Y1_W2BEG[5] ,
    \Tile_X9Y1_W2BEG[4] ,
    \Tile_X9Y1_W2BEG[3] ,
    \Tile_X9Y1_W2BEG[2] ,
    \Tile_X9Y1_W2BEG[1] ,
    \Tile_X9Y1_W2BEG[0] }),
    .W6BEG({\Tile_X8Y1_W6BEG[11] ,
    \Tile_X8Y1_W6BEG[10] ,
    \Tile_X8Y1_W6BEG[9] ,
    \Tile_X8Y1_W6BEG[8] ,
    \Tile_X8Y1_W6BEG[7] ,
    \Tile_X8Y1_W6BEG[6] ,
    \Tile_X8Y1_W6BEG[5] ,
    \Tile_X8Y1_W6BEG[4] ,
    \Tile_X8Y1_W6BEG[3] ,
    \Tile_X8Y1_W6BEG[2] ,
    \Tile_X8Y1_W6BEG[1] ,
    \Tile_X8Y1_W6BEG[0] }),
    .W6END({\Tile_X9Y1_W6BEG[11] ,
    \Tile_X9Y1_W6BEG[10] ,
    \Tile_X9Y1_W6BEG[9] ,
    \Tile_X9Y1_W6BEG[8] ,
    \Tile_X9Y1_W6BEG[7] ,
    \Tile_X9Y1_W6BEG[6] ,
    \Tile_X9Y1_W6BEG[5] ,
    \Tile_X9Y1_W6BEG[4] ,
    \Tile_X9Y1_W6BEG[3] ,
    \Tile_X9Y1_W6BEG[2] ,
    \Tile_X9Y1_W6BEG[1] ,
    \Tile_X9Y1_W6BEG[0] }),
    .WW4BEG({\Tile_X8Y1_WW4BEG[15] ,
    \Tile_X8Y1_WW4BEG[14] ,
    \Tile_X8Y1_WW4BEG[13] ,
    \Tile_X8Y1_WW4BEG[12] ,
    \Tile_X8Y1_WW4BEG[11] ,
    \Tile_X8Y1_WW4BEG[10] ,
    \Tile_X8Y1_WW4BEG[9] ,
    \Tile_X8Y1_WW4BEG[8] ,
    \Tile_X8Y1_WW4BEG[7] ,
    \Tile_X8Y1_WW4BEG[6] ,
    \Tile_X8Y1_WW4BEG[5] ,
    \Tile_X8Y1_WW4BEG[4] ,
    \Tile_X8Y1_WW4BEG[3] ,
    \Tile_X8Y1_WW4BEG[2] ,
    \Tile_X8Y1_WW4BEG[1] ,
    \Tile_X8Y1_WW4BEG[0] }),
    .WW4END({\Tile_X9Y1_WW4BEG[15] ,
    \Tile_X9Y1_WW4BEG[14] ,
    \Tile_X9Y1_WW4BEG[13] ,
    \Tile_X9Y1_WW4BEG[12] ,
    \Tile_X9Y1_WW4BEG[11] ,
    \Tile_X9Y1_WW4BEG[10] ,
    \Tile_X9Y1_WW4BEG[9] ,
    \Tile_X9Y1_WW4BEG[8] ,
    \Tile_X9Y1_WW4BEG[7] ,
    \Tile_X9Y1_WW4BEG[6] ,
    \Tile_X9Y1_WW4BEG[5] ,
    \Tile_X9Y1_WW4BEG[4] ,
    \Tile_X9Y1_WW4BEG[3] ,
    \Tile_X9Y1_WW4BEG[2] ,
    \Tile_X9Y1_WW4BEG[1] ,
    \Tile_X9Y1_WW4BEG[0] }));
 LUT4AB Tile_X8Y2_LUT4AB (.Ci(Tile_X8Y3_Co),
    .Co(Tile_X8Y2_Co),
    .UserCLK(Tile_X8Y3_UserCLKo),
    .UserCLKo(Tile_X8Y2_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X8Y2_E1BEG[3] ,
    \Tile_X8Y2_E1BEG[2] ,
    \Tile_X8Y2_E1BEG[1] ,
    \Tile_X8Y2_E1BEG[0] }),
    .E1END({\Tile_X7Y2_E1BEG[3] ,
    \Tile_X7Y2_E1BEG[2] ,
    \Tile_X7Y2_E1BEG[1] ,
    \Tile_X7Y2_E1BEG[0] }),
    .E2BEG({\Tile_X8Y2_E2BEG[7] ,
    \Tile_X8Y2_E2BEG[6] ,
    \Tile_X8Y2_E2BEG[5] ,
    \Tile_X8Y2_E2BEG[4] ,
    \Tile_X8Y2_E2BEG[3] ,
    \Tile_X8Y2_E2BEG[2] ,
    \Tile_X8Y2_E2BEG[1] ,
    \Tile_X8Y2_E2BEG[0] }),
    .E2BEGb({\Tile_X8Y2_E2BEGb[7] ,
    \Tile_X8Y2_E2BEGb[6] ,
    \Tile_X8Y2_E2BEGb[5] ,
    \Tile_X8Y2_E2BEGb[4] ,
    \Tile_X8Y2_E2BEGb[3] ,
    \Tile_X8Y2_E2BEGb[2] ,
    \Tile_X8Y2_E2BEGb[1] ,
    \Tile_X8Y2_E2BEGb[0] }),
    .E2END({\Tile_X7Y2_E2BEGb[7] ,
    \Tile_X7Y2_E2BEGb[6] ,
    \Tile_X7Y2_E2BEGb[5] ,
    \Tile_X7Y2_E2BEGb[4] ,
    \Tile_X7Y2_E2BEGb[3] ,
    \Tile_X7Y2_E2BEGb[2] ,
    \Tile_X7Y2_E2BEGb[1] ,
    \Tile_X7Y2_E2BEGb[0] }),
    .E2MID({\Tile_X7Y2_E2BEG[7] ,
    \Tile_X7Y2_E2BEG[6] ,
    \Tile_X7Y2_E2BEG[5] ,
    \Tile_X7Y2_E2BEG[4] ,
    \Tile_X7Y2_E2BEG[3] ,
    \Tile_X7Y2_E2BEG[2] ,
    \Tile_X7Y2_E2BEG[1] ,
    \Tile_X7Y2_E2BEG[0] }),
    .E6BEG({\Tile_X8Y2_E6BEG[11] ,
    \Tile_X8Y2_E6BEG[10] ,
    \Tile_X8Y2_E6BEG[9] ,
    \Tile_X8Y2_E6BEG[8] ,
    \Tile_X8Y2_E6BEG[7] ,
    \Tile_X8Y2_E6BEG[6] ,
    \Tile_X8Y2_E6BEG[5] ,
    \Tile_X8Y2_E6BEG[4] ,
    \Tile_X8Y2_E6BEG[3] ,
    \Tile_X8Y2_E6BEG[2] ,
    \Tile_X8Y2_E6BEG[1] ,
    \Tile_X8Y2_E6BEG[0] }),
    .E6END({\Tile_X7Y2_E6BEG[11] ,
    \Tile_X7Y2_E6BEG[10] ,
    \Tile_X7Y2_E6BEG[9] ,
    \Tile_X7Y2_E6BEG[8] ,
    \Tile_X7Y2_E6BEG[7] ,
    \Tile_X7Y2_E6BEG[6] ,
    \Tile_X7Y2_E6BEG[5] ,
    \Tile_X7Y2_E6BEG[4] ,
    \Tile_X7Y2_E6BEG[3] ,
    \Tile_X7Y2_E6BEG[2] ,
    \Tile_X7Y2_E6BEG[1] ,
    \Tile_X7Y2_E6BEG[0] }),
    .EE4BEG({\Tile_X8Y2_EE4BEG[15] ,
    \Tile_X8Y2_EE4BEG[14] ,
    \Tile_X8Y2_EE4BEG[13] ,
    \Tile_X8Y2_EE4BEG[12] ,
    \Tile_X8Y2_EE4BEG[11] ,
    \Tile_X8Y2_EE4BEG[10] ,
    \Tile_X8Y2_EE4BEG[9] ,
    \Tile_X8Y2_EE4BEG[8] ,
    \Tile_X8Y2_EE4BEG[7] ,
    \Tile_X8Y2_EE4BEG[6] ,
    \Tile_X8Y2_EE4BEG[5] ,
    \Tile_X8Y2_EE4BEG[4] ,
    \Tile_X8Y2_EE4BEG[3] ,
    \Tile_X8Y2_EE4BEG[2] ,
    \Tile_X8Y2_EE4BEG[1] ,
    \Tile_X8Y2_EE4BEG[0] }),
    .EE4END({\Tile_X7Y2_EE4BEG[15] ,
    \Tile_X7Y2_EE4BEG[14] ,
    \Tile_X7Y2_EE4BEG[13] ,
    \Tile_X7Y2_EE4BEG[12] ,
    \Tile_X7Y2_EE4BEG[11] ,
    \Tile_X7Y2_EE4BEG[10] ,
    \Tile_X7Y2_EE4BEG[9] ,
    \Tile_X7Y2_EE4BEG[8] ,
    \Tile_X7Y2_EE4BEG[7] ,
    \Tile_X7Y2_EE4BEG[6] ,
    \Tile_X7Y2_EE4BEG[5] ,
    \Tile_X7Y2_EE4BEG[4] ,
    \Tile_X7Y2_EE4BEG[3] ,
    \Tile_X7Y2_EE4BEG[2] ,
    \Tile_X7Y2_EE4BEG[1] ,
    \Tile_X7Y2_EE4BEG[0] }),
    .FrameData({\Tile_X7Y2_FrameData_O[31] ,
    \Tile_X7Y2_FrameData_O[30] ,
    \Tile_X7Y2_FrameData_O[29] ,
    \Tile_X7Y2_FrameData_O[28] ,
    \Tile_X7Y2_FrameData_O[27] ,
    \Tile_X7Y2_FrameData_O[26] ,
    \Tile_X7Y2_FrameData_O[25] ,
    \Tile_X7Y2_FrameData_O[24] ,
    \Tile_X7Y2_FrameData_O[23] ,
    \Tile_X7Y2_FrameData_O[22] ,
    \Tile_X7Y2_FrameData_O[21] ,
    \Tile_X7Y2_FrameData_O[20] ,
    \Tile_X7Y2_FrameData_O[19] ,
    \Tile_X7Y2_FrameData_O[18] ,
    \Tile_X7Y2_FrameData_O[17] ,
    \Tile_X7Y2_FrameData_O[16] ,
    \Tile_X7Y2_FrameData_O[15] ,
    \Tile_X7Y2_FrameData_O[14] ,
    \Tile_X7Y2_FrameData_O[13] ,
    \Tile_X7Y2_FrameData_O[12] ,
    \Tile_X7Y2_FrameData_O[11] ,
    \Tile_X7Y2_FrameData_O[10] ,
    \Tile_X7Y2_FrameData_O[9] ,
    \Tile_X7Y2_FrameData_O[8] ,
    \Tile_X7Y2_FrameData_O[7] ,
    \Tile_X7Y2_FrameData_O[6] ,
    \Tile_X7Y2_FrameData_O[5] ,
    \Tile_X7Y2_FrameData_O[4] ,
    \Tile_X7Y2_FrameData_O[3] ,
    \Tile_X7Y2_FrameData_O[2] ,
    \Tile_X7Y2_FrameData_O[1] ,
    \Tile_X7Y2_FrameData_O[0] }),
    .FrameData_O({\Tile_X8Y2_FrameData_O[31] ,
    \Tile_X8Y2_FrameData_O[30] ,
    \Tile_X8Y2_FrameData_O[29] ,
    \Tile_X8Y2_FrameData_O[28] ,
    \Tile_X8Y2_FrameData_O[27] ,
    \Tile_X8Y2_FrameData_O[26] ,
    \Tile_X8Y2_FrameData_O[25] ,
    \Tile_X8Y2_FrameData_O[24] ,
    \Tile_X8Y2_FrameData_O[23] ,
    \Tile_X8Y2_FrameData_O[22] ,
    \Tile_X8Y2_FrameData_O[21] ,
    \Tile_X8Y2_FrameData_O[20] ,
    \Tile_X8Y2_FrameData_O[19] ,
    \Tile_X8Y2_FrameData_O[18] ,
    \Tile_X8Y2_FrameData_O[17] ,
    \Tile_X8Y2_FrameData_O[16] ,
    \Tile_X8Y2_FrameData_O[15] ,
    \Tile_X8Y2_FrameData_O[14] ,
    \Tile_X8Y2_FrameData_O[13] ,
    \Tile_X8Y2_FrameData_O[12] ,
    \Tile_X8Y2_FrameData_O[11] ,
    \Tile_X8Y2_FrameData_O[10] ,
    \Tile_X8Y2_FrameData_O[9] ,
    \Tile_X8Y2_FrameData_O[8] ,
    \Tile_X8Y2_FrameData_O[7] ,
    \Tile_X8Y2_FrameData_O[6] ,
    \Tile_X8Y2_FrameData_O[5] ,
    \Tile_X8Y2_FrameData_O[4] ,
    \Tile_X8Y2_FrameData_O[3] ,
    \Tile_X8Y2_FrameData_O[2] ,
    \Tile_X8Y2_FrameData_O[1] ,
    \Tile_X8Y2_FrameData_O[0] }),
    .FrameStrobe({\Tile_X8Y3_FrameStrobe_O[19] ,
    \Tile_X8Y3_FrameStrobe_O[18] ,
    \Tile_X8Y3_FrameStrobe_O[17] ,
    \Tile_X8Y3_FrameStrobe_O[16] ,
    \Tile_X8Y3_FrameStrobe_O[15] ,
    \Tile_X8Y3_FrameStrobe_O[14] ,
    \Tile_X8Y3_FrameStrobe_O[13] ,
    \Tile_X8Y3_FrameStrobe_O[12] ,
    \Tile_X8Y3_FrameStrobe_O[11] ,
    \Tile_X8Y3_FrameStrobe_O[10] ,
    \Tile_X8Y3_FrameStrobe_O[9] ,
    \Tile_X8Y3_FrameStrobe_O[8] ,
    \Tile_X8Y3_FrameStrobe_O[7] ,
    \Tile_X8Y3_FrameStrobe_O[6] ,
    \Tile_X8Y3_FrameStrobe_O[5] ,
    \Tile_X8Y3_FrameStrobe_O[4] ,
    \Tile_X8Y3_FrameStrobe_O[3] ,
    \Tile_X8Y3_FrameStrobe_O[2] ,
    \Tile_X8Y3_FrameStrobe_O[1] ,
    \Tile_X8Y3_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X8Y2_FrameStrobe_O[19] ,
    \Tile_X8Y2_FrameStrobe_O[18] ,
    \Tile_X8Y2_FrameStrobe_O[17] ,
    \Tile_X8Y2_FrameStrobe_O[16] ,
    \Tile_X8Y2_FrameStrobe_O[15] ,
    \Tile_X8Y2_FrameStrobe_O[14] ,
    \Tile_X8Y2_FrameStrobe_O[13] ,
    \Tile_X8Y2_FrameStrobe_O[12] ,
    \Tile_X8Y2_FrameStrobe_O[11] ,
    \Tile_X8Y2_FrameStrobe_O[10] ,
    \Tile_X8Y2_FrameStrobe_O[9] ,
    \Tile_X8Y2_FrameStrobe_O[8] ,
    \Tile_X8Y2_FrameStrobe_O[7] ,
    \Tile_X8Y2_FrameStrobe_O[6] ,
    \Tile_X8Y2_FrameStrobe_O[5] ,
    \Tile_X8Y2_FrameStrobe_O[4] ,
    \Tile_X8Y2_FrameStrobe_O[3] ,
    \Tile_X8Y2_FrameStrobe_O[2] ,
    \Tile_X8Y2_FrameStrobe_O[1] ,
    \Tile_X8Y2_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X8Y2_N1BEG[3] ,
    \Tile_X8Y2_N1BEG[2] ,
    \Tile_X8Y2_N1BEG[1] ,
    \Tile_X8Y2_N1BEG[0] }),
    .N1END({\Tile_X8Y3_N1BEG[3] ,
    \Tile_X8Y3_N1BEG[2] ,
    \Tile_X8Y3_N1BEG[1] ,
    \Tile_X8Y3_N1BEG[0] }),
    .N2BEG({\Tile_X8Y2_N2BEG[7] ,
    \Tile_X8Y2_N2BEG[6] ,
    \Tile_X8Y2_N2BEG[5] ,
    \Tile_X8Y2_N2BEG[4] ,
    \Tile_X8Y2_N2BEG[3] ,
    \Tile_X8Y2_N2BEG[2] ,
    \Tile_X8Y2_N2BEG[1] ,
    \Tile_X8Y2_N2BEG[0] }),
    .N2BEGb({\Tile_X8Y2_N2BEGb[7] ,
    \Tile_X8Y2_N2BEGb[6] ,
    \Tile_X8Y2_N2BEGb[5] ,
    \Tile_X8Y2_N2BEGb[4] ,
    \Tile_X8Y2_N2BEGb[3] ,
    \Tile_X8Y2_N2BEGb[2] ,
    \Tile_X8Y2_N2BEGb[1] ,
    \Tile_X8Y2_N2BEGb[0] }),
    .N2END({\Tile_X8Y3_N2BEGb[7] ,
    \Tile_X8Y3_N2BEGb[6] ,
    \Tile_X8Y3_N2BEGb[5] ,
    \Tile_X8Y3_N2BEGb[4] ,
    \Tile_X8Y3_N2BEGb[3] ,
    \Tile_X8Y3_N2BEGb[2] ,
    \Tile_X8Y3_N2BEGb[1] ,
    \Tile_X8Y3_N2BEGb[0] }),
    .N2MID({\Tile_X8Y3_N2BEG[7] ,
    \Tile_X8Y3_N2BEG[6] ,
    \Tile_X8Y3_N2BEG[5] ,
    \Tile_X8Y3_N2BEG[4] ,
    \Tile_X8Y3_N2BEG[3] ,
    \Tile_X8Y3_N2BEG[2] ,
    \Tile_X8Y3_N2BEG[1] ,
    \Tile_X8Y3_N2BEG[0] }),
    .N4BEG({\Tile_X8Y2_N4BEG[15] ,
    \Tile_X8Y2_N4BEG[14] ,
    \Tile_X8Y2_N4BEG[13] ,
    \Tile_X8Y2_N4BEG[12] ,
    \Tile_X8Y2_N4BEG[11] ,
    \Tile_X8Y2_N4BEG[10] ,
    \Tile_X8Y2_N4BEG[9] ,
    \Tile_X8Y2_N4BEG[8] ,
    \Tile_X8Y2_N4BEG[7] ,
    \Tile_X8Y2_N4BEG[6] ,
    \Tile_X8Y2_N4BEG[5] ,
    \Tile_X8Y2_N4BEG[4] ,
    \Tile_X8Y2_N4BEG[3] ,
    \Tile_X8Y2_N4BEG[2] ,
    \Tile_X8Y2_N4BEG[1] ,
    \Tile_X8Y2_N4BEG[0] }),
    .N4END({\Tile_X8Y3_N4BEG[15] ,
    \Tile_X8Y3_N4BEG[14] ,
    \Tile_X8Y3_N4BEG[13] ,
    \Tile_X8Y3_N4BEG[12] ,
    \Tile_X8Y3_N4BEG[11] ,
    \Tile_X8Y3_N4BEG[10] ,
    \Tile_X8Y3_N4BEG[9] ,
    \Tile_X8Y3_N4BEG[8] ,
    \Tile_X8Y3_N4BEG[7] ,
    \Tile_X8Y3_N4BEG[6] ,
    \Tile_X8Y3_N4BEG[5] ,
    \Tile_X8Y3_N4BEG[4] ,
    \Tile_X8Y3_N4BEG[3] ,
    \Tile_X8Y3_N4BEG[2] ,
    \Tile_X8Y3_N4BEG[1] ,
    \Tile_X8Y3_N4BEG[0] }),
    .NN4BEG({\Tile_X8Y2_NN4BEG[15] ,
    \Tile_X8Y2_NN4BEG[14] ,
    \Tile_X8Y2_NN4BEG[13] ,
    \Tile_X8Y2_NN4BEG[12] ,
    \Tile_X8Y2_NN4BEG[11] ,
    \Tile_X8Y2_NN4BEG[10] ,
    \Tile_X8Y2_NN4BEG[9] ,
    \Tile_X8Y2_NN4BEG[8] ,
    \Tile_X8Y2_NN4BEG[7] ,
    \Tile_X8Y2_NN4BEG[6] ,
    \Tile_X8Y2_NN4BEG[5] ,
    \Tile_X8Y2_NN4BEG[4] ,
    \Tile_X8Y2_NN4BEG[3] ,
    \Tile_X8Y2_NN4BEG[2] ,
    \Tile_X8Y2_NN4BEG[1] ,
    \Tile_X8Y2_NN4BEG[0] }),
    .NN4END({\Tile_X8Y3_NN4BEG[15] ,
    \Tile_X8Y3_NN4BEG[14] ,
    \Tile_X8Y3_NN4BEG[13] ,
    \Tile_X8Y3_NN4BEG[12] ,
    \Tile_X8Y3_NN4BEG[11] ,
    \Tile_X8Y3_NN4BEG[10] ,
    \Tile_X8Y3_NN4BEG[9] ,
    \Tile_X8Y3_NN4BEG[8] ,
    \Tile_X8Y3_NN4BEG[7] ,
    \Tile_X8Y3_NN4BEG[6] ,
    \Tile_X8Y3_NN4BEG[5] ,
    \Tile_X8Y3_NN4BEG[4] ,
    \Tile_X8Y3_NN4BEG[3] ,
    \Tile_X8Y3_NN4BEG[2] ,
    \Tile_X8Y3_NN4BEG[1] ,
    \Tile_X8Y3_NN4BEG[0] }),
    .S1BEG({\Tile_X8Y2_S1BEG[3] ,
    \Tile_X8Y2_S1BEG[2] ,
    \Tile_X8Y2_S1BEG[1] ,
    \Tile_X8Y2_S1BEG[0] }),
    .S1END({\Tile_X8Y1_S1BEG[3] ,
    \Tile_X8Y1_S1BEG[2] ,
    \Tile_X8Y1_S1BEG[1] ,
    \Tile_X8Y1_S1BEG[0] }),
    .S2BEG({\Tile_X8Y2_S2BEG[7] ,
    \Tile_X8Y2_S2BEG[6] ,
    \Tile_X8Y2_S2BEG[5] ,
    \Tile_X8Y2_S2BEG[4] ,
    \Tile_X8Y2_S2BEG[3] ,
    \Tile_X8Y2_S2BEG[2] ,
    \Tile_X8Y2_S2BEG[1] ,
    \Tile_X8Y2_S2BEG[0] }),
    .S2BEGb({\Tile_X8Y2_S2BEGb[7] ,
    \Tile_X8Y2_S2BEGb[6] ,
    \Tile_X8Y2_S2BEGb[5] ,
    \Tile_X8Y2_S2BEGb[4] ,
    \Tile_X8Y2_S2BEGb[3] ,
    \Tile_X8Y2_S2BEGb[2] ,
    \Tile_X8Y2_S2BEGb[1] ,
    \Tile_X8Y2_S2BEGb[0] }),
    .S2END({\Tile_X8Y1_S2BEGb[7] ,
    \Tile_X8Y1_S2BEGb[6] ,
    \Tile_X8Y1_S2BEGb[5] ,
    \Tile_X8Y1_S2BEGb[4] ,
    \Tile_X8Y1_S2BEGb[3] ,
    \Tile_X8Y1_S2BEGb[2] ,
    \Tile_X8Y1_S2BEGb[1] ,
    \Tile_X8Y1_S2BEGb[0] }),
    .S2MID({\Tile_X8Y1_S2BEG[7] ,
    \Tile_X8Y1_S2BEG[6] ,
    \Tile_X8Y1_S2BEG[5] ,
    \Tile_X8Y1_S2BEG[4] ,
    \Tile_X8Y1_S2BEG[3] ,
    \Tile_X8Y1_S2BEG[2] ,
    \Tile_X8Y1_S2BEG[1] ,
    \Tile_X8Y1_S2BEG[0] }),
    .S4BEG({\Tile_X8Y2_S4BEG[15] ,
    \Tile_X8Y2_S4BEG[14] ,
    \Tile_X8Y2_S4BEG[13] ,
    \Tile_X8Y2_S4BEG[12] ,
    \Tile_X8Y2_S4BEG[11] ,
    \Tile_X8Y2_S4BEG[10] ,
    \Tile_X8Y2_S4BEG[9] ,
    \Tile_X8Y2_S4BEG[8] ,
    \Tile_X8Y2_S4BEG[7] ,
    \Tile_X8Y2_S4BEG[6] ,
    \Tile_X8Y2_S4BEG[5] ,
    \Tile_X8Y2_S4BEG[4] ,
    \Tile_X8Y2_S4BEG[3] ,
    \Tile_X8Y2_S4BEG[2] ,
    \Tile_X8Y2_S4BEG[1] ,
    \Tile_X8Y2_S4BEG[0] }),
    .S4END({\Tile_X8Y1_S4BEG[15] ,
    \Tile_X8Y1_S4BEG[14] ,
    \Tile_X8Y1_S4BEG[13] ,
    \Tile_X8Y1_S4BEG[12] ,
    \Tile_X8Y1_S4BEG[11] ,
    \Tile_X8Y1_S4BEG[10] ,
    \Tile_X8Y1_S4BEG[9] ,
    \Tile_X8Y1_S4BEG[8] ,
    \Tile_X8Y1_S4BEG[7] ,
    \Tile_X8Y1_S4BEG[6] ,
    \Tile_X8Y1_S4BEG[5] ,
    \Tile_X8Y1_S4BEG[4] ,
    \Tile_X8Y1_S4BEG[3] ,
    \Tile_X8Y1_S4BEG[2] ,
    \Tile_X8Y1_S4BEG[1] ,
    \Tile_X8Y1_S4BEG[0] }),
    .SS4BEG({\Tile_X8Y2_SS4BEG[15] ,
    \Tile_X8Y2_SS4BEG[14] ,
    \Tile_X8Y2_SS4BEG[13] ,
    \Tile_X8Y2_SS4BEG[12] ,
    \Tile_X8Y2_SS4BEG[11] ,
    \Tile_X8Y2_SS4BEG[10] ,
    \Tile_X8Y2_SS4BEG[9] ,
    \Tile_X8Y2_SS4BEG[8] ,
    \Tile_X8Y2_SS4BEG[7] ,
    \Tile_X8Y2_SS4BEG[6] ,
    \Tile_X8Y2_SS4BEG[5] ,
    \Tile_X8Y2_SS4BEG[4] ,
    \Tile_X8Y2_SS4BEG[3] ,
    \Tile_X8Y2_SS4BEG[2] ,
    \Tile_X8Y2_SS4BEG[1] ,
    \Tile_X8Y2_SS4BEG[0] }),
    .SS4END({\Tile_X8Y1_SS4BEG[15] ,
    \Tile_X8Y1_SS4BEG[14] ,
    \Tile_X8Y1_SS4BEG[13] ,
    \Tile_X8Y1_SS4BEG[12] ,
    \Tile_X8Y1_SS4BEG[11] ,
    \Tile_X8Y1_SS4BEG[10] ,
    \Tile_X8Y1_SS4BEG[9] ,
    \Tile_X8Y1_SS4BEG[8] ,
    \Tile_X8Y1_SS4BEG[7] ,
    \Tile_X8Y1_SS4BEG[6] ,
    \Tile_X8Y1_SS4BEG[5] ,
    \Tile_X8Y1_SS4BEG[4] ,
    \Tile_X8Y1_SS4BEG[3] ,
    \Tile_X8Y1_SS4BEG[2] ,
    \Tile_X8Y1_SS4BEG[1] ,
    \Tile_X8Y1_SS4BEG[0] }),
    .W1BEG({\Tile_X8Y2_W1BEG[3] ,
    \Tile_X8Y2_W1BEG[2] ,
    \Tile_X8Y2_W1BEG[1] ,
    \Tile_X8Y2_W1BEG[0] }),
    .W1END({\Tile_X9Y2_W1BEG[3] ,
    \Tile_X9Y2_W1BEG[2] ,
    \Tile_X9Y2_W1BEG[1] ,
    \Tile_X9Y2_W1BEG[0] }),
    .W2BEG({\Tile_X8Y2_W2BEG[7] ,
    \Tile_X8Y2_W2BEG[6] ,
    \Tile_X8Y2_W2BEG[5] ,
    \Tile_X8Y2_W2BEG[4] ,
    \Tile_X8Y2_W2BEG[3] ,
    \Tile_X8Y2_W2BEG[2] ,
    \Tile_X8Y2_W2BEG[1] ,
    \Tile_X8Y2_W2BEG[0] }),
    .W2BEGb({\Tile_X8Y2_W2BEGb[7] ,
    \Tile_X8Y2_W2BEGb[6] ,
    \Tile_X8Y2_W2BEGb[5] ,
    \Tile_X8Y2_W2BEGb[4] ,
    \Tile_X8Y2_W2BEGb[3] ,
    \Tile_X8Y2_W2BEGb[2] ,
    \Tile_X8Y2_W2BEGb[1] ,
    \Tile_X8Y2_W2BEGb[0] }),
    .W2END({\Tile_X9Y2_W2BEGb[7] ,
    \Tile_X9Y2_W2BEGb[6] ,
    \Tile_X9Y2_W2BEGb[5] ,
    \Tile_X9Y2_W2BEGb[4] ,
    \Tile_X9Y2_W2BEGb[3] ,
    \Tile_X9Y2_W2BEGb[2] ,
    \Tile_X9Y2_W2BEGb[1] ,
    \Tile_X9Y2_W2BEGb[0] }),
    .W2MID({\Tile_X9Y2_W2BEG[7] ,
    \Tile_X9Y2_W2BEG[6] ,
    \Tile_X9Y2_W2BEG[5] ,
    \Tile_X9Y2_W2BEG[4] ,
    \Tile_X9Y2_W2BEG[3] ,
    \Tile_X9Y2_W2BEG[2] ,
    \Tile_X9Y2_W2BEG[1] ,
    \Tile_X9Y2_W2BEG[0] }),
    .W6BEG({\Tile_X8Y2_W6BEG[11] ,
    \Tile_X8Y2_W6BEG[10] ,
    \Tile_X8Y2_W6BEG[9] ,
    \Tile_X8Y2_W6BEG[8] ,
    \Tile_X8Y2_W6BEG[7] ,
    \Tile_X8Y2_W6BEG[6] ,
    \Tile_X8Y2_W6BEG[5] ,
    \Tile_X8Y2_W6BEG[4] ,
    \Tile_X8Y2_W6BEG[3] ,
    \Tile_X8Y2_W6BEG[2] ,
    \Tile_X8Y2_W6BEG[1] ,
    \Tile_X8Y2_W6BEG[0] }),
    .W6END({\Tile_X9Y2_W6BEG[11] ,
    \Tile_X9Y2_W6BEG[10] ,
    \Tile_X9Y2_W6BEG[9] ,
    \Tile_X9Y2_W6BEG[8] ,
    \Tile_X9Y2_W6BEG[7] ,
    \Tile_X9Y2_W6BEG[6] ,
    \Tile_X9Y2_W6BEG[5] ,
    \Tile_X9Y2_W6BEG[4] ,
    \Tile_X9Y2_W6BEG[3] ,
    \Tile_X9Y2_W6BEG[2] ,
    \Tile_X9Y2_W6BEG[1] ,
    \Tile_X9Y2_W6BEG[0] }),
    .WW4BEG({\Tile_X8Y2_WW4BEG[15] ,
    \Tile_X8Y2_WW4BEG[14] ,
    \Tile_X8Y2_WW4BEG[13] ,
    \Tile_X8Y2_WW4BEG[12] ,
    \Tile_X8Y2_WW4BEG[11] ,
    \Tile_X8Y2_WW4BEG[10] ,
    \Tile_X8Y2_WW4BEG[9] ,
    \Tile_X8Y2_WW4BEG[8] ,
    \Tile_X8Y2_WW4BEG[7] ,
    \Tile_X8Y2_WW4BEG[6] ,
    \Tile_X8Y2_WW4BEG[5] ,
    \Tile_X8Y2_WW4BEG[4] ,
    \Tile_X8Y2_WW4BEG[3] ,
    \Tile_X8Y2_WW4BEG[2] ,
    \Tile_X8Y2_WW4BEG[1] ,
    \Tile_X8Y2_WW4BEG[0] }),
    .WW4END({\Tile_X9Y2_WW4BEG[15] ,
    \Tile_X9Y2_WW4BEG[14] ,
    \Tile_X9Y2_WW4BEG[13] ,
    \Tile_X9Y2_WW4BEG[12] ,
    \Tile_X9Y2_WW4BEG[11] ,
    \Tile_X9Y2_WW4BEG[10] ,
    \Tile_X9Y2_WW4BEG[9] ,
    \Tile_X9Y2_WW4BEG[8] ,
    \Tile_X9Y2_WW4BEG[7] ,
    \Tile_X9Y2_WW4BEG[6] ,
    \Tile_X9Y2_WW4BEG[5] ,
    \Tile_X9Y2_WW4BEG[4] ,
    \Tile_X9Y2_WW4BEG[3] ,
    \Tile_X9Y2_WW4BEG[2] ,
    \Tile_X9Y2_WW4BEG[1] ,
    \Tile_X9Y2_WW4BEG[0] }));
 LUT4AB Tile_X8Y3_LUT4AB (.Ci(Tile_X8Y4_Co),
    .Co(Tile_X8Y3_Co),
    .UserCLK(Tile_X8Y4_UserCLKo),
    .UserCLKo(Tile_X8Y3_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X8Y3_E1BEG[3] ,
    \Tile_X8Y3_E1BEG[2] ,
    \Tile_X8Y3_E1BEG[1] ,
    \Tile_X8Y3_E1BEG[0] }),
    .E1END({\Tile_X7Y3_E1BEG[3] ,
    \Tile_X7Y3_E1BEG[2] ,
    \Tile_X7Y3_E1BEG[1] ,
    \Tile_X7Y3_E1BEG[0] }),
    .E2BEG({\Tile_X8Y3_E2BEG[7] ,
    \Tile_X8Y3_E2BEG[6] ,
    \Tile_X8Y3_E2BEG[5] ,
    \Tile_X8Y3_E2BEG[4] ,
    \Tile_X8Y3_E2BEG[3] ,
    \Tile_X8Y3_E2BEG[2] ,
    \Tile_X8Y3_E2BEG[1] ,
    \Tile_X8Y3_E2BEG[0] }),
    .E2BEGb({\Tile_X8Y3_E2BEGb[7] ,
    \Tile_X8Y3_E2BEGb[6] ,
    \Tile_X8Y3_E2BEGb[5] ,
    \Tile_X8Y3_E2BEGb[4] ,
    \Tile_X8Y3_E2BEGb[3] ,
    \Tile_X8Y3_E2BEGb[2] ,
    \Tile_X8Y3_E2BEGb[1] ,
    \Tile_X8Y3_E2BEGb[0] }),
    .E2END({\Tile_X7Y3_E2BEGb[7] ,
    \Tile_X7Y3_E2BEGb[6] ,
    \Tile_X7Y3_E2BEGb[5] ,
    \Tile_X7Y3_E2BEGb[4] ,
    \Tile_X7Y3_E2BEGb[3] ,
    \Tile_X7Y3_E2BEGb[2] ,
    \Tile_X7Y3_E2BEGb[1] ,
    \Tile_X7Y3_E2BEGb[0] }),
    .E2MID({\Tile_X7Y3_E2BEG[7] ,
    \Tile_X7Y3_E2BEG[6] ,
    \Tile_X7Y3_E2BEG[5] ,
    \Tile_X7Y3_E2BEG[4] ,
    \Tile_X7Y3_E2BEG[3] ,
    \Tile_X7Y3_E2BEG[2] ,
    \Tile_X7Y3_E2BEG[1] ,
    \Tile_X7Y3_E2BEG[0] }),
    .E6BEG({\Tile_X8Y3_E6BEG[11] ,
    \Tile_X8Y3_E6BEG[10] ,
    \Tile_X8Y3_E6BEG[9] ,
    \Tile_X8Y3_E6BEG[8] ,
    \Tile_X8Y3_E6BEG[7] ,
    \Tile_X8Y3_E6BEG[6] ,
    \Tile_X8Y3_E6BEG[5] ,
    \Tile_X8Y3_E6BEG[4] ,
    \Tile_X8Y3_E6BEG[3] ,
    \Tile_X8Y3_E6BEG[2] ,
    \Tile_X8Y3_E6BEG[1] ,
    \Tile_X8Y3_E6BEG[0] }),
    .E6END({\Tile_X7Y3_E6BEG[11] ,
    \Tile_X7Y3_E6BEG[10] ,
    \Tile_X7Y3_E6BEG[9] ,
    \Tile_X7Y3_E6BEG[8] ,
    \Tile_X7Y3_E6BEG[7] ,
    \Tile_X7Y3_E6BEG[6] ,
    \Tile_X7Y3_E6BEG[5] ,
    \Tile_X7Y3_E6BEG[4] ,
    \Tile_X7Y3_E6BEG[3] ,
    \Tile_X7Y3_E6BEG[2] ,
    \Tile_X7Y3_E6BEG[1] ,
    \Tile_X7Y3_E6BEG[0] }),
    .EE4BEG({\Tile_X8Y3_EE4BEG[15] ,
    \Tile_X8Y3_EE4BEG[14] ,
    \Tile_X8Y3_EE4BEG[13] ,
    \Tile_X8Y3_EE4BEG[12] ,
    \Tile_X8Y3_EE4BEG[11] ,
    \Tile_X8Y3_EE4BEG[10] ,
    \Tile_X8Y3_EE4BEG[9] ,
    \Tile_X8Y3_EE4BEG[8] ,
    \Tile_X8Y3_EE4BEG[7] ,
    \Tile_X8Y3_EE4BEG[6] ,
    \Tile_X8Y3_EE4BEG[5] ,
    \Tile_X8Y3_EE4BEG[4] ,
    \Tile_X8Y3_EE4BEG[3] ,
    \Tile_X8Y3_EE4BEG[2] ,
    \Tile_X8Y3_EE4BEG[1] ,
    \Tile_X8Y3_EE4BEG[0] }),
    .EE4END({\Tile_X7Y3_EE4BEG[15] ,
    \Tile_X7Y3_EE4BEG[14] ,
    \Tile_X7Y3_EE4BEG[13] ,
    \Tile_X7Y3_EE4BEG[12] ,
    \Tile_X7Y3_EE4BEG[11] ,
    \Tile_X7Y3_EE4BEG[10] ,
    \Tile_X7Y3_EE4BEG[9] ,
    \Tile_X7Y3_EE4BEG[8] ,
    \Tile_X7Y3_EE4BEG[7] ,
    \Tile_X7Y3_EE4BEG[6] ,
    \Tile_X7Y3_EE4BEG[5] ,
    \Tile_X7Y3_EE4BEG[4] ,
    \Tile_X7Y3_EE4BEG[3] ,
    \Tile_X7Y3_EE4BEG[2] ,
    \Tile_X7Y3_EE4BEG[1] ,
    \Tile_X7Y3_EE4BEG[0] }),
    .FrameData({\Tile_X7Y3_FrameData_O[31] ,
    \Tile_X7Y3_FrameData_O[30] ,
    \Tile_X7Y3_FrameData_O[29] ,
    \Tile_X7Y3_FrameData_O[28] ,
    \Tile_X7Y3_FrameData_O[27] ,
    \Tile_X7Y3_FrameData_O[26] ,
    \Tile_X7Y3_FrameData_O[25] ,
    \Tile_X7Y3_FrameData_O[24] ,
    \Tile_X7Y3_FrameData_O[23] ,
    \Tile_X7Y3_FrameData_O[22] ,
    \Tile_X7Y3_FrameData_O[21] ,
    \Tile_X7Y3_FrameData_O[20] ,
    \Tile_X7Y3_FrameData_O[19] ,
    \Tile_X7Y3_FrameData_O[18] ,
    \Tile_X7Y3_FrameData_O[17] ,
    \Tile_X7Y3_FrameData_O[16] ,
    \Tile_X7Y3_FrameData_O[15] ,
    \Tile_X7Y3_FrameData_O[14] ,
    \Tile_X7Y3_FrameData_O[13] ,
    \Tile_X7Y3_FrameData_O[12] ,
    \Tile_X7Y3_FrameData_O[11] ,
    \Tile_X7Y3_FrameData_O[10] ,
    \Tile_X7Y3_FrameData_O[9] ,
    \Tile_X7Y3_FrameData_O[8] ,
    \Tile_X7Y3_FrameData_O[7] ,
    \Tile_X7Y3_FrameData_O[6] ,
    \Tile_X7Y3_FrameData_O[5] ,
    \Tile_X7Y3_FrameData_O[4] ,
    \Tile_X7Y3_FrameData_O[3] ,
    \Tile_X7Y3_FrameData_O[2] ,
    \Tile_X7Y3_FrameData_O[1] ,
    \Tile_X7Y3_FrameData_O[0] }),
    .FrameData_O({\Tile_X8Y3_FrameData_O[31] ,
    \Tile_X8Y3_FrameData_O[30] ,
    \Tile_X8Y3_FrameData_O[29] ,
    \Tile_X8Y3_FrameData_O[28] ,
    \Tile_X8Y3_FrameData_O[27] ,
    \Tile_X8Y3_FrameData_O[26] ,
    \Tile_X8Y3_FrameData_O[25] ,
    \Tile_X8Y3_FrameData_O[24] ,
    \Tile_X8Y3_FrameData_O[23] ,
    \Tile_X8Y3_FrameData_O[22] ,
    \Tile_X8Y3_FrameData_O[21] ,
    \Tile_X8Y3_FrameData_O[20] ,
    \Tile_X8Y3_FrameData_O[19] ,
    \Tile_X8Y3_FrameData_O[18] ,
    \Tile_X8Y3_FrameData_O[17] ,
    \Tile_X8Y3_FrameData_O[16] ,
    \Tile_X8Y3_FrameData_O[15] ,
    \Tile_X8Y3_FrameData_O[14] ,
    \Tile_X8Y3_FrameData_O[13] ,
    \Tile_X8Y3_FrameData_O[12] ,
    \Tile_X8Y3_FrameData_O[11] ,
    \Tile_X8Y3_FrameData_O[10] ,
    \Tile_X8Y3_FrameData_O[9] ,
    \Tile_X8Y3_FrameData_O[8] ,
    \Tile_X8Y3_FrameData_O[7] ,
    \Tile_X8Y3_FrameData_O[6] ,
    \Tile_X8Y3_FrameData_O[5] ,
    \Tile_X8Y3_FrameData_O[4] ,
    \Tile_X8Y3_FrameData_O[3] ,
    \Tile_X8Y3_FrameData_O[2] ,
    \Tile_X8Y3_FrameData_O[1] ,
    \Tile_X8Y3_FrameData_O[0] }),
    .FrameStrobe({\Tile_X8Y4_FrameStrobe_O[19] ,
    \Tile_X8Y4_FrameStrobe_O[18] ,
    \Tile_X8Y4_FrameStrobe_O[17] ,
    \Tile_X8Y4_FrameStrobe_O[16] ,
    \Tile_X8Y4_FrameStrobe_O[15] ,
    \Tile_X8Y4_FrameStrobe_O[14] ,
    \Tile_X8Y4_FrameStrobe_O[13] ,
    \Tile_X8Y4_FrameStrobe_O[12] ,
    \Tile_X8Y4_FrameStrobe_O[11] ,
    \Tile_X8Y4_FrameStrobe_O[10] ,
    \Tile_X8Y4_FrameStrobe_O[9] ,
    \Tile_X8Y4_FrameStrobe_O[8] ,
    \Tile_X8Y4_FrameStrobe_O[7] ,
    \Tile_X8Y4_FrameStrobe_O[6] ,
    \Tile_X8Y4_FrameStrobe_O[5] ,
    \Tile_X8Y4_FrameStrobe_O[4] ,
    \Tile_X8Y4_FrameStrobe_O[3] ,
    \Tile_X8Y4_FrameStrobe_O[2] ,
    \Tile_X8Y4_FrameStrobe_O[1] ,
    \Tile_X8Y4_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X8Y3_FrameStrobe_O[19] ,
    \Tile_X8Y3_FrameStrobe_O[18] ,
    \Tile_X8Y3_FrameStrobe_O[17] ,
    \Tile_X8Y3_FrameStrobe_O[16] ,
    \Tile_X8Y3_FrameStrobe_O[15] ,
    \Tile_X8Y3_FrameStrobe_O[14] ,
    \Tile_X8Y3_FrameStrobe_O[13] ,
    \Tile_X8Y3_FrameStrobe_O[12] ,
    \Tile_X8Y3_FrameStrobe_O[11] ,
    \Tile_X8Y3_FrameStrobe_O[10] ,
    \Tile_X8Y3_FrameStrobe_O[9] ,
    \Tile_X8Y3_FrameStrobe_O[8] ,
    \Tile_X8Y3_FrameStrobe_O[7] ,
    \Tile_X8Y3_FrameStrobe_O[6] ,
    \Tile_X8Y3_FrameStrobe_O[5] ,
    \Tile_X8Y3_FrameStrobe_O[4] ,
    \Tile_X8Y3_FrameStrobe_O[3] ,
    \Tile_X8Y3_FrameStrobe_O[2] ,
    \Tile_X8Y3_FrameStrobe_O[1] ,
    \Tile_X8Y3_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X8Y3_N1BEG[3] ,
    \Tile_X8Y3_N1BEG[2] ,
    \Tile_X8Y3_N1BEG[1] ,
    \Tile_X8Y3_N1BEG[0] }),
    .N1END({\Tile_X8Y4_N1BEG[3] ,
    \Tile_X8Y4_N1BEG[2] ,
    \Tile_X8Y4_N1BEG[1] ,
    \Tile_X8Y4_N1BEG[0] }),
    .N2BEG({\Tile_X8Y3_N2BEG[7] ,
    \Tile_X8Y3_N2BEG[6] ,
    \Tile_X8Y3_N2BEG[5] ,
    \Tile_X8Y3_N2BEG[4] ,
    \Tile_X8Y3_N2BEG[3] ,
    \Tile_X8Y3_N2BEG[2] ,
    \Tile_X8Y3_N2BEG[1] ,
    \Tile_X8Y3_N2BEG[0] }),
    .N2BEGb({\Tile_X8Y3_N2BEGb[7] ,
    \Tile_X8Y3_N2BEGb[6] ,
    \Tile_X8Y3_N2BEGb[5] ,
    \Tile_X8Y3_N2BEGb[4] ,
    \Tile_X8Y3_N2BEGb[3] ,
    \Tile_X8Y3_N2BEGb[2] ,
    \Tile_X8Y3_N2BEGb[1] ,
    \Tile_X8Y3_N2BEGb[0] }),
    .N2END({\Tile_X8Y4_N2BEGb[7] ,
    \Tile_X8Y4_N2BEGb[6] ,
    \Tile_X8Y4_N2BEGb[5] ,
    \Tile_X8Y4_N2BEGb[4] ,
    \Tile_X8Y4_N2BEGb[3] ,
    \Tile_X8Y4_N2BEGb[2] ,
    \Tile_X8Y4_N2BEGb[1] ,
    \Tile_X8Y4_N2BEGb[0] }),
    .N2MID({\Tile_X8Y4_N2BEG[7] ,
    \Tile_X8Y4_N2BEG[6] ,
    \Tile_X8Y4_N2BEG[5] ,
    \Tile_X8Y4_N2BEG[4] ,
    \Tile_X8Y4_N2BEG[3] ,
    \Tile_X8Y4_N2BEG[2] ,
    \Tile_X8Y4_N2BEG[1] ,
    \Tile_X8Y4_N2BEG[0] }),
    .N4BEG({\Tile_X8Y3_N4BEG[15] ,
    \Tile_X8Y3_N4BEG[14] ,
    \Tile_X8Y3_N4BEG[13] ,
    \Tile_X8Y3_N4BEG[12] ,
    \Tile_X8Y3_N4BEG[11] ,
    \Tile_X8Y3_N4BEG[10] ,
    \Tile_X8Y3_N4BEG[9] ,
    \Tile_X8Y3_N4BEG[8] ,
    \Tile_X8Y3_N4BEG[7] ,
    \Tile_X8Y3_N4BEG[6] ,
    \Tile_X8Y3_N4BEG[5] ,
    \Tile_X8Y3_N4BEG[4] ,
    \Tile_X8Y3_N4BEG[3] ,
    \Tile_X8Y3_N4BEG[2] ,
    \Tile_X8Y3_N4BEG[1] ,
    \Tile_X8Y3_N4BEG[0] }),
    .N4END({\Tile_X8Y4_N4BEG[15] ,
    \Tile_X8Y4_N4BEG[14] ,
    \Tile_X8Y4_N4BEG[13] ,
    \Tile_X8Y4_N4BEG[12] ,
    \Tile_X8Y4_N4BEG[11] ,
    \Tile_X8Y4_N4BEG[10] ,
    \Tile_X8Y4_N4BEG[9] ,
    \Tile_X8Y4_N4BEG[8] ,
    \Tile_X8Y4_N4BEG[7] ,
    \Tile_X8Y4_N4BEG[6] ,
    \Tile_X8Y4_N4BEG[5] ,
    \Tile_X8Y4_N4BEG[4] ,
    \Tile_X8Y4_N4BEG[3] ,
    \Tile_X8Y4_N4BEG[2] ,
    \Tile_X8Y4_N4BEG[1] ,
    \Tile_X8Y4_N4BEG[0] }),
    .NN4BEG({\Tile_X8Y3_NN4BEG[15] ,
    \Tile_X8Y3_NN4BEG[14] ,
    \Tile_X8Y3_NN4BEG[13] ,
    \Tile_X8Y3_NN4BEG[12] ,
    \Tile_X8Y3_NN4BEG[11] ,
    \Tile_X8Y3_NN4BEG[10] ,
    \Tile_X8Y3_NN4BEG[9] ,
    \Tile_X8Y3_NN4BEG[8] ,
    \Tile_X8Y3_NN4BEG[7] ,
    \Tile_X8Y3_NN4BEG[6] ,
    \Tile_X8Y3_NN4BEG[5] ,
    \Tile_X8Y3_NN4BEG[4] ,
    \Tile_X8Y3_NN4BEG[3] ,
    \Tile_X8Y3_NN4BEG[2] ,
    \Tile_X8Y3_NN4BEG[1] ,
    \Tile_X8Y3_NN4BEG[0] }),
    .NN4END({\Tile_X8Y4_NN4BEG[15] ,
    \Tile_X8Y4_NN4BEG[14] ,
    \Tile_X8Y4_NN4BEG[13] ,
    \Tile_X8Y4_NN4BEG[12] ,
    \Tile_X8Y4_NN4BEG[11] ,
    \Tile_X8Y4_NN4BEG[10] ,
    \Tile_X8Y4_NN4BEG[9] ,
    \Tile_X8Y4_NN4BEG[8] ,
    \Tile_X8Y4_NN4BEG[7] ,
    \Tile_X8Y4_NN4BEG[6] ,
    \Tile_X8Y4_NN4BEG[5] ,
    \Tile_X8Y4_NN4BEG[4] ,
    \Tile_X8Y4_NN4BEG[3] ,
    \Tile_X8Y4_NN4BEG[2] ,
    \Tile_X8Y4_NN4BEG[1] ,
    \Tile_X8Y4_NN4BEG[0] }),
    .S1BEG({\Tile_X8Y3_S1BEG[3] ,
    \Tile_X8Y3_S1BEG[2] ,
    \Tile_X8Y3_S1BEG[1] ,
    \Tile_X8Y3_S1BEG[0] }),
    .S1END({\Tile_X8Y2_S1BEG[3] ,
    \Tile_X8Y2_S1BEG[2] ,
    \Tile_X8Y2_S1BEG[1] ,
    \Tile_X8Y2_S1BEG[0] }),
    .S2BEG({\Tile_X8Y3_S2BEG[7] ,
    \Tile_X8Y3_S2BEG[6] ,
    \Tile_X8Y3_S2BEG[5] ,
    \Tile_X8Y3_S2BEG[4] ,
    \Tile_X8Y3_S2BEG[3] ,
    \Tile_X8Y3_S2BEG[2] ,
    \Tile_X8Y3_S2BEG[1] ,
    \Tile_X8Y3_S2BEG[0] }),
    .S2BEGb({\Tile_X8Y3_S2BEGb[7] ,
    \Tile_X8Y3_S2BEGb[6] ,
    \Tile_X8Y3_S2BEGb[5] ,
    \Tile_X8Y3_S2BEGb[4] ,
    \Tile_X8Y3_S2BEGb[3] ,
    \Tile_X8Y3_S2BEGb[2] ,
    \Tile_X8Y3_S2BEGb[1] ,
    \Tile_X8Y3_S2BEGb[0] }),
    .S2END({\Tile_X8Y2_S2BEGb[7] ,
    \Tile_X8Y2_S2BEGb[6] ,
    \Tile_X8Y2_S2BEGb[5] ,
    \Tile_X8Y2_S2BEGb[4] ,
    \Tile_X8Y2_S2BEGb[3] ,
    \Tile_X8Y2_S2BEGb[2] ,
    \Tile_X8Y2_S2BEGb[1] ,
    \Tile_X8Y2_S2BEGb[0] }),
    .S2MID({\Tile_X8Y2_S2BEG[7] ,
    \Tile_X8Y2_S2BEG[6] ,
    \Tile_X8Y2_S2BEG[5] ,
    \Tile_X8Y2_S2BEG[4] ,
    \Tile_X8Y2_S2BEG[3] ,
    \Tile_X8Y2_S2BEG[2] ,
    \Tile_X8Y2_S2BEG[1] ,
    \Tile_X8Y2_S2BEG[0] }),
    .S4BEG({\Tile_X8Y3_S4BEG[15] ,
    \Tile_X8Y3_S4BEG[14] ,
    \Tile_X8Y3_S4BEG[13] ,
    \Tile_X8Y3_S4BEG[12] ,
    \Tile_X8Y3_S4BEG[11] ,
    \Tile_X8Y3_S4BEG[10] ,
    \Tile_X8Y3_S4BEG[9] ,
    \Tile_X8Y3_S4BEG[8] ,
    \Tile_X8Y3_S4BEG[7] ,
    \Tile_X8Y3_S4BEG[6] ,
    \Tile_X8Y3_S4BEG[5] ,
    \Tile_X8Y3_S4BEG[4] ,
    \Tile_X8Y3_S4BEG[3] ,
    \Tile_X8Y3_S4BEG[2] ,
    \Tile_X8Y3_S4BEG[1] ,
    \Tile_X8Y3_S4BEG[0] }),
    .S4END({\Tile_X8Y2_S4BEG[15] ,
    \Tile_X8Y2_S4BEG[14] ,
    \Tile_X8Y2_S4BEG[13] ,
    \Tile_X8Y2_S4BEG[12] ,
    \Tile_X8Y2_S4BEG[11] ,
    \Tile_X8Y2_S4BEG[10] ,
    \Tile_X8Y2_S4BEG[9] ,
    \Tile_X8Y2_S4BEG[8] ,
    \Tile_X8Y2_S4BEG[7] ,
    \Tile_X8Y2_S4BEG[6] ,
    \Tile_X8Y2_S4BEG[5] ,
    \Tile_X8Y2_S4BEG[4] ,
    \Tile_X8Y2_S4BEG[3] ,
    \Tile_X8Y2_S4BEG[2] ,
    \Tile_X8Y2_S4BEG[1] ,
    \Tile_X8Y2_S4BEG[0] }),
    .SS4BEG({\Tile_X8Y3_SS4BEG[15] ,
    \Tile_X8Y3_SS4BEG[14] ,
    \Tile_X8Y3_SS4BEG[13] ,
    \Tile_X8Y3_SS4BEG[12] ,
    \Tile_X8Y3_SS4BEG[11] ,
    \Tile_X8Y3_SS4BEG[10] ,
    \Tile_X8Y3_SS4BEG[9] ,
    \Tile_X8Y3_SS4BEG[8] ,
    \Tile_X8Y3_SS4BEG[7] ,
    \Tile_X8Y3_SS4BEG[6] ,
    \Tile_X8Y3_SS4BEG[5] ,
    \Tile_X8Y3_SS4BEG[4] ,
    \Tile_X8Y3_SS4BEG[3] ,
    \Tile_X8Y3_SS4BEG[2] ,
    \Tile_X8Y3_SS4BEG[1] ,
    \Tile_X8Y3_SS4BEG[0] }),
    .SS4END({\Tile_X8Y2_SS4BEG[15] ,
    \Tile_X8Y2_SS4BEG[14] ,
    \Tile_X8Y2_SS4BEG[13] ,
    \Tile_X8Y2_SS4BEG[12] ,
    \Tile_X8Y2_SS4BEG[11] ,
    \Tile_X8Y2_SS4BEG[10] ,
    \Tile_X8Y2_SS4BEG[9] ,
    \Tile_X8Y2_SS4BEG[8] ,
    \Tile_X8Y2_SS4BEG[7] ,
    \Tile_X8Y2_SS4BEG[6] ,
    \Tile_X8Y2_SS4BEG[5] ,
    \Tile_X8Y2_SS4BEG[4] ,
    \Tile_X8Y2_SS4BEG[3] ,
    \Tile_X8Y2_SS4BEG[2] ,
    \Tile_X8Y2_SS4BEG[1] ,
    \Tile_X8Y2_SS4BEG[0] }),
    .W1BEG({\Tile_X8Y3_W1BEG[3] ,
    \Tile_X8Y3_W1BEG[2] ,
    \Tile_X8Y3_W1BEG[1] ,
    \Tile_X8Y3_W1BEG[0] }),
    .W1END({\Tile_X9Y3_W1BEG[3] ,
    \Tile_X9Y3_W1BEG[2] ,
    \Tile_X9Y3_W1BEG[1] ,
    \Tile_X9Y3_W1BEG[0] }),
    .W2BEG({\Tile_X8Y3_W2BEG[7] ,
    \Tile_X8Y3_W2BEG[6] ,
    \Tile_X8Y3_W2BEG[5] ,
    \Tile_X8Y3_W2BEG[4] ,
    \Tile_X8Y3_W2BEG[3] ,
    \Tile_X8Y3_W2BEG[2] ,
    \Tile_X8Y3_W2BEG[1] ,
    \Tile_X8Y3_W2BEG[0] }),
    .W2BEGb({\Tile_X8Y3_W2BEGb[7] ,
    \Tile_X8Y3_W2BEGb[6] ,
    \Tile_X8Y3_W2BEGb[5] ,
    \Tile_X8Y3_W2BEGb[4] ,
    \Tile_X8Y3_W2BEGb[3] ,
    \Tile_X8Y3_W2BEGb[2] ,
    \Tile_X8Y3_W2BEGb[1] ,
    \Tile_X8Y3_W2BEGb[0] }),
    .W2END({\Tile_X9Y3_W2BEGb[7] ,
    \Tile_X9Y3_W2BEGb[6] ,
    \Tile_X9Y3_W2BEGb[5] ,
    \Tile_X9Y3_W2BEGb[4] ,
    \Tile_X9Y3_W2BEGb[3] ,
    \Tile_X9Y3_W2BEGb[2] ,
    \Tile_X9Y3_W2BEGb[1] ,
    \Tile_X9Y3_W2BEGb[0] }),
    .W2MID({\Tile_X9Y3_W2BEG[7] ,
    \Tile_X9Y3_W2BEG[6] ,
    \Tile_X9Y3_W2BEG[5] ,
    \Tile_X9Y3_W2BEG[4] ,
    \Tile_X9Y3_W2BEG[3] ,
    \Tile_X9Y3_W2BEG[2] ,
    \Tile_X9Y3_W2BEG[1] ,
    \Tile_X9Y3_W2BEG[0] }),
    .W6BEG({\Tile_X8Y3_W6BEG[11] ,
    \Tile_X8Y3_W6BEG[10] ,
    \Tile_X8Y3_W6BEG[9] ,
    \Tile_X8Y3_W6BEG[8] ,
    \Tile_X8Y3_W6BEG[7] ,
    \Tile_X8Y3_W6BEG[6] ,
    \Tile_X8Y3_W6BEG[5] ,
    \Tile_X8Y3_W6BEG[4] ,
    \Tile_X8Y3_W6BEG[3] ,
    \Tile_X8Y3_W6BEG[2] ,
    \Tile_X8Y3_W6BEG[1] ,
    \Tile_X8Y3_W6BEG[0] }),
    .W6END({\Tile_X9Y3_W6BEG[11] ,
    \Tile_X9Y3_W6BEG[10] ,
    \Tile_X9Y3_W6BEG[9] ,
    \Tile_X9Y3_W6BEG[8] ,
    \Tile_X9Y3_W6BEG[7] ,
    \Tile_X9Y3_W6BEG[6] ,
    \Tile_X9Y3_W6BEG[5] ,
    \Tile_X9Y3_W6BEG[4] ,
    \Tile_X9Y3_W6BEG[3] ,
    \Tile_X9Y3_W6BEG[2] ,
    \Tile_X9Y3_W6BEG[1] ,
    \Tile_X9Y3_W6BEG[0] }),
    .WW4BEG({\Tile_X8Y3_WW4BEG[15] ,
    \Tile_X8Y3_WW4BEG[14] ,
    \Tile_X8Y3_WW4BEG[13] ,
    \Tile_X8Y3_WW4BEG[12] ,
    \Tile_X8Y3_WW4BEG[11] ,
    \Tile_X8Y3_WW4BEG[10] ,
    \Tile_X8Y3_WW4BEG[9] ,
    \Tile_X8Y3_WW4BEG[8] ,
    \Tile_X8Y3_WW4BEG[7] ,
    \Tile_X8Y3_WW4BEG[6] ,
    \Tile_X8Y3_WW4BEG[5] ,
    \Tile_X8Y3_WW4BEG[4] ,
    \Tile_X8Y3_WW4BEG[3] ,
    \Tile_X8Y3_WW4BEG[2] ,
    \Tile_X8Y3_WW4BEG[1] ,
    \Tile_X8Y3_WW4BEG[0] }),
    .WW4END({\Tile_X9Y3_WW4BEG[15] ,
    \Tile_X9Y3_WW4BEG[14] ,
    \Tile_X9Y3_WW4BEG[13] ,
    \Tile_X9Y3_WW4BEG[12] ,
    \Tile_X9Y3_WW4BEG[11] ,
    \Tile_X9Y3_WW4BEG[10] ,
    \Tile_X9Y3_WW4BEG[9] ,
    \Tile_X9Y3_WW4BEG[8] ,
    \Tile_X9Y3_WW4BEG[7] ,
    \Tile_X9Y3_WW4BEG[6] ,
    \Tile_X9Y3_WW4BEG[5] ,
    \Tile_X9Y3_WW4BEG[4] ,
    \Tile_X9Y3_WW4BEG[3] ,
    \Tile_X9Y3_WW4BEG[2] ,
    \Tile_X9Y3_WW4BEG[1] ,
    \Tile_X9Y3_WW4BEG[0] }));
 LUT4AB Tile_X8Y4_LUT4AB (.Ci(Tile_X8Y5_Co),
    .Co(Tile_X8Y4_Co),
    .UserCLK(Tile_X8Y5_UserCLKo),
    .UserCLKo(Tile_X8Y4_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X8Y4_E1BEG[3] ,
    \Tile_X8Y4_E1BEG[2] ,
    \Tile_X8Y4_E1BEG[1] ,
    \Tile_X8Y4_E1BEG[0] }),
    .E1END({\Tile_X7Y4_E1BEG[3] ,
    \Tile_X7Y4_E1BEG[2] ,
    \Tile_X7Y4_E1BEG[1] ,
    \Tile_X7Y4_E1BEG[0] }),
    .E2BEG({\Tile_X8Y4_E2BEG[7] ,
    \Tile_X8Y4_E2BEG[6] ,
    \Tile_X8Y4_E2BEG[5] ,
    \Tile_X8Y4_E2BEG[4] ,
    \Tile_X8Y4_E2BEG[3] ,
    \Tile_X8Y4_E2BEG[2] ,
    \Tile_X8Y4_E2BEG[1] ,
    \Tile_X8Y4_E2BEG[0] }),
    .E2BEGb({\Tile_X8Y4_E2BEGb[7] ,
    \Tile_X8Y4_E2BEGb[6] ,
    \Tile_X8Y4_E2BEGb[5] ,
    \Tile_X8Y4_E2BEGb[4] ,
    \Tile_X8Y4_E2BEGb[3] ,
    \Tile_X8Y4_E2BEGb[2] ,
    \Tile_X8Y4_E2BEGb[1] ,
    \Tile_X8Y4_E2BEGb[0] }),
    .E2END({\Tile_X7Y4_E2BEGb[7] ,
    \Tile_X7Y4_E2BEGb[6] ,
    \Tile_X7Y4_E2BEGb[5] ,
    \Tile_X7Y4_E2BEGb[4] ,
    \Tile_X7Y4_E2BEGb[3] ,
    \Tile_X7Y4_E2BEGb[2] ,
    \Tile_X7Y4_E2BEGb[1] ,
    \Tile_X7Y4_E2BEGb[0] }),
    .E2MID({\Tile_X7Y4_E2BEG[7] ,
    \Tile_X7Y4_E2BEG[6] ,
    \Tile_X7Y4_E2BEG[5] ,
    \Tile_X7Y4_E2BEG[4] ,
    \Tile_X7Y4_E2BEG[3] ,
    \Tile_X7Y4_E2BEG[2] ,
    \Tile_X7Y4_E2BEG[1] ,
    \Tile_X7Y4_E2BEG[0] }),
    .E6BEG({\Tile_X8Y4_E6BEG[11] ,
    \Tile_X8Y4_E6BEG[10] ,
    \Tile_X8Y4_E6BEG[9] ,
    \Tile_X8Y4_E6BEG[8] ,
    \Tile_X8Y4_E6BEG[7] ,
    \Tile_X8Y4_E6BEG[6] ,
    \Tile_X8Y4_E6BEG[5] ,
    \Tile_X8Y4_E6BEG[4] ,
    \Tile_X8Y4_E6BEG[3] ,
    \Tile_X8Y4_E6BEG[2] ,
    \Tile_X8Y4_E6BEG[1] ,
    \Tile_X8Y4_E6BEG[0] }),
    .E6END({\Tile_X7Y4_E6BEG[11] ,
    \Tile_X7Y4_E6BEG[10] ,
    \Tile_X7Y4_E6BEG[9] ,
    \Tile_X7Y4_E6BEG[8] ,
    \Tile_X7Y4_E6BEG[7] ,
    \Tile_X7Y4_E6BEG[6] ,
    \Tile_X7Y4_E6BEG[5] ,
    \Tile_X7Y4_E6BEG[4] ,
    \Tile_X7Y4_E6BEG[3] ,
    \Tile_X7Y4_E6BEG[2] ,
    \Tile_X7Y4_E6BEG[1] ,
    \Tile_X7Y4_E6BEG[0] }),
    .EE4BEG({\Tile_X8Y4_EE4BEG[15] ,
    \Tile_X8Y4_EE4BEG[14] ,
    \Tile_X8Y4_EE4BEG[13] ,
    \Tile_X8Y4_EE4BEG[12] ,
    \Tile_X8Y4_EE4BEG[11] ,
    \Tile_X8Y4_EE4BEG[10] ,
    \Tile_X8Y4_EE4BEG[9] ,
    \Tile_X8Y4_EE4BEG[8] ,
    \Tile_X8Y4_EE4BEG[7] ,
    \Tile_X8Y4_EE4BEG[6] ,
    \Tile_X8Y4_EE4BEG[5] ,
    \Tile_X8Y4_EE4BEG[4] ,
    \Tile_X8Y4_EE4BEG[3] ,
    \Tile_X8Y4_EE4BEG[2] ,
    \Tile_X8Y4_EE4BEG[1] ,
    \Tile_X8Y4_EE4BEG[0] }),
    .EE4END({\Tile_X7Y4_EE4BEG[15] ,
    \Tile_X7Y4_EE4BEG[14] ,
    \Tile_X7Y4_EE4BEG[13] ,
    \Tile_X7Y4_EE4BEG[12] ,
    \Tile_X7Y4_EE4BEG[11] ,
    \Tile_X7Y4_EE4BEG[10] ,
    \Tile_X7Y4_EE4BEG[9] ,
    \Tile_X7Y4_EE4BEG[8] ,
    \Tile_X7Y4_EE4BEG[7] ,
    \Tile_X7Y4_EE4BEG[6] ,
    \Tile_X7Y4_EE4BEG[5] ,
    \Tile_X7Y4_EE4BEG[4] ,
    \Tile_X7Y4_EE4BEG[3] ,
    \Tile_X7Y4_EE4BEG[2] ,
    \Tile_X7Y4_EE4BEG[1] ,
    \Tile_X7Y4_EE4BEG[0] }),
    .FrameData({\Tile_X7Y4_FrameData_O[31] ,
    \Tile_X7Y4_FrameData_O[30] ,
    \Tile_X7Y4_FrameData_O[29] ,
    \Tile_X7Y4_FrameData_O[28] ,
    \Tile_X7Y4_FrameData_O[27] ,
    \Tile_X7Y4_FrameData_O[26] ,
    \Tile_X7Y4_FrameData_O[25] ,
    \Tile_X7Y4_FrameData_O[24] ,
    \Tile_X7Y4_FrameData_O[23] ,
    \Tile_X7Y4_FrameData_O[22] ,
    \Tile_X7Y4_FrameData_O[21] ,
    \Tile_X7Y4_FrameData_O[20] ,
    \Tile_X7Y4_FrameData_O[19] ,
    \Tile_X7Y4_FrameData_O[18] ,
    \Tile_X7Y4_FrameData_O[17] ,
    \Tile_X7Y4_FrameData_O[16] ,
    \Tile_X7Y4_FrameData_O[15] ,
    \Tile_X7Y4_FrameData_O[14] ,
    \Tile_X7Y4_FrameData_O[13] ,
    \Tile_X7Y4_FrameData_O[12] ,
    \Tile_X7Y4_FrameData_O[11] ,
    \Tile_X7Y4_FrameData_O[10] ,
    \Tile_X7Y4_FrameData_O[9] ,
    \Tile_X7Y4_FrameData_O[8] ,
    \Tile_X7Y4_FrameData_O[7] ,
    \Tile_X7Y4_FrameData_O[6] ,
    \Tile_X7Y4_FrameData_O[5] ,
    \Tile_X7Y4_FrameData_O[4] ,
    \Tile_X7Y4_FrameData_O[3] ,
    \Tile_X7Y4_FrameData_O[2] ,
    \Tile_X7Y4_FrameData_O[1] ,
    \Tile_X7Y4_FrameData_O[0] }),
    .FrameData_O({\Tile_X8Y4_FrameData_O[31] ,
    \Tile_X8Y4_FrameData_O[30] ,
    \Tile_X8Y4_FrameData_O[29] ,
    \Tile_X8Y4_FrameData_O[28] ,
    \Tile_X8Y4_FrameData_O[27] ,
    \Tile_X8Y4_FrameData_O[26] ,
    \Tile_X8Y4_FrameData_O[25] ,
    \Tile_X8Y4_FrameData_O[24] ,
    \Tile_X8Y4_FrameData_O[23] ,
    \Tile_X8Y4_FrameData_O[22] ,
    \Tile_X8Y4_FrameData_O[21] ,
    \Tile_X8Y4_FrameData_O[20] ,
    \Tile_X8Y4_FrameData_O[19] ,
    \Tile_X8Y4_FrameData_O[18] ,
    \Tile_X8Y4_FrameData_O[17] ,
    \Tile_X8Y4_FrameData_O[16] ,
    \Tile_X8Y4_FrameData_O[15] ,
    \Tile_X8Y4_FrameData_O[14] ,
    \Tile_X8Y4_FrameData_O[13] ,
    \Tile_X8Y4_FrameData_O[12] ,
    \Tile_X8Y4_FrameData_O[11] ,
    \Tile_X8Y4_FrameData_O[10] ,
    \Tile_X8Y4_FrameData_O[9] ,
    \Tile_X8Y4_FrameData_O[8] ,
    \Tile_X8Y4_FrameData_O[7] ,
    \Tile_X8Y4_FrameData_O[6] ,
    \Tile_X8Y4_FrameData_O[5] ,
    \Tile_X8Y4_FrameData_O[4] ,
    \Tile_X8Y4_FrameData_O[3] ,
    \Tile_X8Y4_FrameData_O[2] ,
    \Tile_X8Y4_FrameData_O[1] ,
    \Tile_X8Y4_FrameData_O[0] }),
    .FrameStrobe({\Tile_X8Y5_FrameStrobe_O[19] ,
    \Tile_X8Y5_FrameStrobe_O[18] ,
    \Tile_X8Y5_FrameStrobe_O[17] ,
    \Tile_X8Y5_FrameStrobe_O[16] ,
    \Tile_X8Y5_FrameStrobe_O[15] ,
    \Tile_X8Y5_FrameStrobe_O[14] ,
    \Tile_X8Y5_FrameStrobe_O[13] ,
    \Tile_X8Y5_FrameStrobe_O[12] ,
    \Tile_X8Y5_FrameStrobe_O[11] ,
    \Tile_X8Y5_FrameStrobe_O[10] ,
    \Tile_X8Y5_FrameStrobe_O[9] ,
    \Tile_X8Y5_FrameStrobe_O[8] ,
    \Tile_X8Y5_FrameStrobe_O[7] ,
    \Tile_X8Y5_FrameStrobe_O[6] ,
    \Tile_X8Y5_FrameStrobe_O[5] ,
    \Tile_X8Y5_FrameStrobe_O[4] ,
    \Tile_X8Y5_FrameStrobe_O[3] ,
    \Tile_X8Y5_FrameStrobe_O[2] ,
    \Tile_X8Y5_FrameStrobe_O[1] ,
    \Tile_X8Y5_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X8Y4_FrameStrobe_O[19] ,
    \Tile_X8Y4_FrameStrobe_O[18] ,
    \Tile_X8Y4_FrameStrobe_O[17] ,
    \Tile_X8Y4_FrameStrobe_O[16] ,
    \Tile_X8Y4_FrameStrobe_O[15] ,
    \Tile_X8Y4_FrameStrobe_O[14] ,
    \Tile_X8Y4_FrameStrobe_O[13] ,
    \Tile_X8Y4_FrameStrobe_O[12] ,
    \Tile_X8Y4_FrameStrobe_O[11] ,
    \Tile_X8Y4_FrameStrobe_O[10] ,
    \Tile_X8Y4_FrameStrobe_O[9] ,
    \Tile_X8Y4_FrameStrobe_O[8] ,
    \Tile_X8Y4_FrameStrobe_O[7] ,
    \Tile_X8Y4_FrameStrobe_O[6] ,
    \Tile_X8Y4_FrameStrobe_O[5] ,
    \Tile_X8Y4_FrameStrobe_O[4] ,
    \Tile_X8Y4_FrameStrobe_O[3] ,
    \Tile_X8Y4_FrameStrobe_O[2] ,
    \Tile_X8Y4_FrameStrobe_O[1] ,
    \Tile_X8Y4_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X8Y4_N1BEG[3] ,
    \Tile_X8Y4_N1BEG[2] ,
    \Tile_X8Y4_N1BEG[1] ,
    \Tile_X8Y4_N1BEG[0] }),
    .N1END({\Tile_X8Y5_N1BEG[3] ,
    \Tile_X8Y5_N1BEG[2] ,
    \Tile_X8Y5_N1BEG[1] ,
    \Tile_X8Y5_N1BEG[0] }),
    .N2BEG({\Tile_X8Y4_N2BEG[7] ,
    \Tile_X8Y4_N2BEG[6] ,
    \Tile_X8Y4_N2BEG[5] ,
    \Tile_X8Y4_N2BEG[4] ,
    \Tile_X8Y4_N2BEG[3] ,
    \Tile_X8Y4_N2BEG[2] ,
    \Tile_X8Y4_N2BEG[1] ,
    \Tile_X8Y4_N2BEG[0] }),
    .N2BEGb({\Tile_X8Y4_N2BEGb[7] ,
    \Tile_X8Y4_N2BEGb[6] ,
    \Tile_X8Y4_N2BEGb[5] ,
    \Tile_X8Y4_N2BEGb[4] ,
    \Tile_X8Y4_N2BEGb[3] ,
    \Tile_X8Y4_N2BEGb[2] ,
    \Tile_X8Y4_N2BEGb[1] ,
    \Tile_X8Y4_N2BEGb[0] }),
    .N2END({\Tile_X8Y5_N2BEGb[7] ,
    \Tile_X8Y5_N2BEGb[6] ,
    \Tile_X8Y5_N2BEGb[5] ,
    \Tile_X8Y5_N2BEGb[4] ,
    \Tile_X8Y5_N2BEGb[3] ,
    \Tile_X8Y5_N2BEGb[2] ,
    \Tile_X8Y5_N2BEGb[1] ,
    \Tile_X8Y5_N2BEGb[0] }),
    .N2MID({\Tile_X8Y5_N2BEG[7] ,
    \Tile_X8Y5_N2BEG[6] ,
    \Tile_X8Y5_N2BEG[5] ,
    \Tile_X8Y5_N2BEG[4] ,
    \Tile_X8Y5_N2BEG[3] ,
    \Tile_X8Y5_N2BEG[2] ,
    \Tile_X8Y5_N2BEG[1] ,
    \Tile_X8Y5_N2BEG[0] }),
    .N4BEG({\Tile_X8Y4_N4BEG[15] ,
    \Tile_X8Y4_N4BEG[14] ,
    \Tile_X8Y4_N4BEG[13] ,
    \Tile_X8Y4_N4BEG[12] ,
    \Tile_X8Y4_N4BEG[11] ,
    \Tile_X8Y4_N4BEG[10] ,
    \Tile_X8Y4_N4BEG[9] ,
    \Tile_X8Y4_N4BEG[8] ,
    \Tile_X8Y4_N4BEG[7] ,
    \Tile_X8Y4_N4BEG[6] ,
    \Tile_X8Y4_N4BEG[5] ,
    \Tile_X8Y4_N4BEG[4] ,
    \Tile_X8Y4_N4BEG[3] ,
    \Tile_X8Y4_N4BEG[2] ,
    \Tile_X8Y4_N4BEG[1] ,
    \Tile_X8Y4_N4BEG[0] }),
    .N4END({\Tile_X8Y5_N4BEG[15] ,
    \Tile_X8Y5_N4BEG[14] ,
    \Tile_X8Y5_N4BEG[13] ,
    \Tile_X8Y5_N4BEG[12] ,
    \Tile_X8Y5_N4BEG[11] ,
    \Tile_X8Y5_N4BEG[10] ,
    \Tile_X8Y5_N4BEG[9] ,
    \Tile_X8Y5_N4BEG[8] ,
    \Tile_X8Y5_N4BEG[7] ,
    \Tile_X8Y5_N4BEG[6] ,
    \Tile_X8Y5_N4BEG[5] ,
    \Tile_X8Y5_N4BEG[4] ,
    \Tile_X8Y5_N4BEG[3] ,
    \Tile_X8Y5_N4BEG[2] ,
    \Tile_X8Y5_N4BEG[1] ,
    \Tile_X8Y5_N4BEG[0] }),
    .NN4BEG({\Tile_X8Y4_NN4BEG[15] ,
    \Tile_X8Y4_NN4BEG[14] ,
    \Tile_X8Y4_NN4BEG[13] ,
    \Tile_X8Y4_NN4BEG[12] ,
    \Tile_X8Y4_NN4BEG[11] ,
    \Tile_X8Y4_NN4BEG[10] ,
    \Tile_X8Y4_NN4BEG[9] ,
    \Tile_X8Y4_NN4BEG[8] ,
    \Tile_X8Y4_NN4BEG[7] ,
    \Tile_X8Y4_NN4BEG[6] ,
    \Tile_X8Y4_NN4BEG[5] ,
    \Tile_X8Y4_NN4BEG[4] ,
    \Tile_X8Y4_NN4BEG[3] ,
    \Tile_X8Y4_NN4BEG[2] ,
    \Tile_X8Y4_NN4BEG[1] ,
    \Tile_X8Y4_NN4BEG[0] }),
    .NN4END({\Tile_X8Y5_NN4BEG[15] ,
    \Tile_X8Y5_NN4BEG[14] ,
    \Tile_X8Y5_NN4BEG[13] ,
    \Tile_X8Y5_NN4BEG[12] ,
    \Tile_X8Y5_NN4BEG[11] ,
    \Tile_X8Y5_NN4BEG[10] ,
    \Tile_X8Y5_NN4BEG[9] ,
    \Tile_X8Y5_NN4BEG[8] ,
    \Tile_X8Y5_NN4BEG[7] ,
    \Tile_X8Y5_NN4BEG[6] ,
    \Tile_X8Y5_NN4BEG[5] ,
    \Tile_X8Y5_NN4BEG[4] ,
    \Tile_X8Y5_NN4BEG[3] ,
    \Tile_X8Y5_NN4BEG[2] ,
    \Tile_X8Y5_NN4BEG[1] ,
    \Tile_X8Y5_NN4BEG[0] }),
    .S1BEG({\Tile_X8Y4_S1BEG[3] ,
    \Tile_X8Y4_S1BEG[2] ,
    \Tile_X8Y4_S1BEG[1] ,
    \Tile_X8Y4_S1BEG[0] }),
    .S1END({\Tile_X8Y3_S1BEG[3] ,
    \Tile_X8Y3_S1BEG[2] ,
    \Tile_X8Y3_S1BEG[1] ,
    \Tile_X8Y3_S1BEG[0] }),
    .S2BEG({\Tile_X8Y4_S2BEG[7] ,
    \Tile_X8Y4_S2BEG[6] ,
    \Tile_X8Y4_S2BEG[5] ,
    \Tile_X8Y4_S2BEG[4] ,
    \Tile_X8Y4_S2BEG[3] ,
    \Tile_X8Y4_S2BEG[2] ,
    \Tile_X8Y4_S2BEG[1] ,
    \Tile_X8Y4_S2BEG[0] }),
    .S2BEGb({\Tile_X8Y4_S2BEGb[7] ,
    \Tile_X8Y4_S2BEGb[6] ,
    \Tile_X8Y4_S2BEGb[5] ,
    \Tile_X8Y4_S2BEGb[4] ,
    \Tile_X8Y4_S2BEGb[3] ,
    \Tile_X8Y4_S2BEGb[2] ,
    \Tile_X8Y4_S2BEGb[1] ,
    \Tile_X8Y4_S2BEGb[0] }),
    .S2END({\Tile_X8Y3_S2BEGb[7] ,
    \Tile_X8Y3_S2BEGb[6] ,
    \Tile_X8Y3_S2BEGb[5] ,
    \Tile_X8Y3_S2BEGb[4] ,
    \Tile_X8Y3_S2BEGb[3] ,
    \Tile_X8Y3_S2BEGb[2] ,
    \Tile_X8Y3_S2BEGb[1] ,
    \Tile_X8Y3_S2BEGb[0] }),
    .S2MID({\Tile_X8Y3_S2BEG[7] ,
    \Tile_X8Y3_S2BEG[6] ,
    \Tile_X8Y3_S2BEG[5] ,
    \Tile_X8Y3_S2BEG[4] ,
    \Tile_X8Y3_S2BEG[3] ,
    \Tile_X8Y3_S2BEG[2] ,
    \Tile_X8Y3_S2BEG[1] ,
    \Tile_X8Y3_S2BEG[0] }),
    .S4BEG({\Tile_X8Y4_S4BEG[15] ,
    \Tile_X8Y4_S4BEG[14] ,
    \Tile_X8Y4_S4BEG[13] ,
    \Tile_X8Y4_S4BEG[12] ,
    \Tile_X8Y4_S4BEG[11] ,
    \Tile_X8Y4_S4BEG[10] ,
    \Tile_X8Y4_S4BEG[9] ,
    \Tile_X8Y4_S4BEG[8] ,
    \Tile_X8Y4_S4BEG[7] ,
    \Tile_X8Y4_S4BEG[6] ,
    \Tile_X8Y4_S4BEG[5] ,
    \Tile_X8Y4_S4BEG[4] ,
    \Tile_X8Y4_S4BEG[3] ,
    \Tile_X8Y4_S4BEG[2] ,
    \Tile_X8Y4_S4BEG[1] ,
    \Tile_X8Y4_S4BEG[0] }),
    .S4END({\Tile_X8Y3_S4BEG[15] ,
    \Tile_X8Y3_S4BEG[14] ,
    \Tile_X8Y3_S4BEG[13] ,
    \Tile_X8Y3_S4BEG[12] ,
    \Tile_X8Y3_S4BEG[11] ,
    \Tile_X8Y3_S4BEG[10] ,
    \Tile_X8Y3_S4BEG[9] ,
    \Tile_X8Y3_S4BEG[8] ,
    \Tile_X8Y3_S4BEG[7] ,
    \Tile_X8Y3_S4BEG[6] ,
    \Tile_X8Y3_S4BEG[5] ,
    \Tile_X8Y3_S4BEG[4] ,
    \Tile_X8Y3_S4BEG[3] ,
    \Tile_X8Y3_S4BEG[2] ,
    \Tile_X8Y3_S4BEG[1] ,
    \Tile_X8Y3_S4BEG[0] }),
    .SS4BEG({\Tile_X8Y4_SS4BEG[15] ,
    \Tile_X8Y4_SS4BEG[14] ,
    \Tile_X8Y4_SS4BEG[13] ,
    \Tile_X8Y4_SS4BEG[12] ,
    \Tile_X8Y4_SS4BEG[11] ,
    \Tile_X8Y4_SS4BEG[10] ,
    \Tile_X8Y4_SS4BEG[9] ,
    \Tile_X8Y4_SS4BEG[8] ,
    \Tile_X8Y4_SS4BEG[7] ,
    \Tile_X8Y4_SS4BEG[6] ,
    \Tile_X8Y4_SS4BEG[5] ,
    \Tile_X8Y4_SS4BEG[4] ,
    \Tile_X8Y4_SS4BEG[3] ,
    \Tile_X8Y4_SS4BEG[2] ,
    \Tile_X8Y4_SS4BEG[1] ,
    \Tile_X8Y4_SS4BEG[0] }),
    .SS4END({\Tile_X8Y3_SS4BEG[15] ,
    \Tile_X8Y3_SS4BEG[14] ,
    \Tile_X8Y3_SS4BEG[13] ,
    \Tile_X8Y3_SS4BEG[12] ,
    \Tile_X8Y3_SS4BEG[11] ,
    \Tile_X8Y3_SS4BEG[10] ,
    \Tile_X8Y3_SS4BEG[9] ,
    \Tile_X8Y3_SS4BEG[8] ,
    \Tile_X8Y3_SS4BEG[7] ,
    \Tile_X8Y3_SS4BEG[6] ,
    \Tile_X8Y3_SS4BEG[5] ,
    \Tile_X8Y3_SS4BEG[4] ,
    \Tile_X8Y3_SS4BEG[3] ,
    \Tile_X8Y3_SS4BEG[2] ,
    \Tile_X8Y3_SS4BEG[1] ,
    \Tile_X8Y3_SS4BEG[0] }),
    .W1BEG({\Tile_X8Y4_W1BEG[3] ,
    \Tile_X8Y4_W1BEG[2] ,
    \Tile_X8Y4_W1BEG[1] ,
    \Tile_X8Y4_W1BEG[0] }),
    .W1END({\Tile_X9Y4_W1BEG[3] ,
    \Tile_X9Y4_W1BEG[2] ,
    \Tile_X9Y4_W1BEG[1] ,
    \Tile_X9Y4_W1BEG[0] }),
    .W2BEG({\Tile_X8Y4_W2BEG[7] ,
    \Tile_X8Y4_W2BEG[6] ,
    \Tile_X8Y4_W2BEG[5] ,
    \Tile_X8Y4_W2BEG[4] ,
    \Tile_X8Y4_W2BEG[3] ,
    \Tile_X8Y4_W2BEG[2] ,
    \Tile_X8Y4_W2BEG[1] ,
    \Tile_X8Y4_W2BEG[0] }),
    .W2BEGb({\Tile_X8Y4_W2BEGb[7] ,
    \Tile_X8Y4_W2BEGb[6] ,
    \Tile_X8Y4_W2BEGb[5] ,
    \Tile_X8Y4_W2BEGb[4] ,
    \Tile_X8Y4_W2BEGb[3] ,
    \Tile_X8Y4_W2BEGb[2] ,
    \Tile_X8Y4_W2BEGb[1] ,
    \Tile_X8Y4_W2BEGb[0] }),
    .W2END({\Tile_X9Y4_W2BEGb[7] ,
    \Tile_X9Y4_W2BEGb[6] ,
    \Tile_X9Y4_W2BEGb[5] ,
    \Tile_X9Y4_W2BEGb[4] ,
    \Tile_X9Y4_W2BEGb[3] ,
    \Tile_X9Y4_W2BEGb[2] ,
    \Tile_X9Y4_W2BEGb[1] ,
    \Tile_X9Y4_W2BEGb[0] }),
    .W2MID({\Tile_X9Y4_W2BEG[7] ,
    \Tile_X9Y4_W2BEG[6] ,
    \Tile_X9Y4_W2BEG[5] ,
    \Tile_X9Y4_W2BEG[4] ,
    \Tile_X9Y4_W2BEG[3] ,
    \Tile_X9Y4_W2BEG[2] ,
    \Tile_X9Y4_W2BEG[1] ,
    \Tile_X9Y4_W2BEG[0] }),
    .W6BEG({\Tile_X8Y4_W6BEG[11] ,
    \Tile_X8Y4_W6BEG[10] ,
    \Tile_X8Y4_W6BEG[9] ,
    \Tile_X8Y4_W6BEG[8] ,
    \Tile_X8Y4_W6BEG[7] ,
    \Tile_X8Y4_W6BEG[6] ,
    \Tile_X8Y4_W6BEG[5] ,
    \Tile_X8Y4_W6BEG[4] ,
    \Tile_X8Y4_W6BEG[3] ,
    \Tile_X8Y4_W6BEG[2] ,
    \Tile_X8Y4_W6BEG[1] ,
    \Tile_X8Y4_W6BEG[0] }),
    .W6END({\Tile_X9Y4_W6BEG[11] ,
    \Tile_X9Y4_W6BEG[10] ,
    \Tile_X9Y4_W6BEG[9] ,
    \Tile_X9Y4_W6BEG[8] ,
    \Tile_X9Y4_W6BEG[7] ,
    \Tile_X9Y4_W6BEG[6] ,
    \Tile_X9Y4_W6BEG[5] ,
    \Tile_X9Y4_W6BEG[4] ,
    \Tile_X9Y4_W6BEG[3] ,
    \Tile_X9Y4_W6BEG[2] ,
    \Tile_X9Y4_W6BEG[1] ,
    \Tile_X9Y4_W6BEG[0] }),
    .WW4BEG({\Tile_X8Y4_WW4BEG[15] ,
    \Tile_X8Y4_WW4BEG[14] ,
    \Tile_X8Y4_WW4BEG[13] ,
    \Tile_X8Y4_WW4BEG[12] ,
    \Tile_X8Y4_WW4BEG[11] ,
    \Tile_X8Y4_WW4BEG[10] ,
    \Tile_X8Y4_WW4BEG[9] ,
    \Tile_X8Y4_WW4BEG[8] ,
    \Tile_X8Y4_WW4BEG[7] ,
    \Tile_X8Y4_WW4BEG[6] ,
    \Tile_X8Y4_WW4BEG[5] ,
    \Tile_X8Y4_WW4BEG[4] ,
    \Tile_X8Y4_WW4BEG[3] ,
    \Tile_X8Y4_WW4BEG[2] ,
    \Tile_X8Y4_WW4BEG[1] ,
    \Tile_X8Y4_WW4BEG[0] }),
    .WW4END({\Tile_X9Y4_WW4BEG[15] ,
    \Tile_X9Y4_WW4BEG[14] ,
    \Tile_X9Y4_WW4BEG[13] ,
    \Tile_X9Y4_WW4BEG[12] ,
    \Tile_X9Y4_WW4BEG[11] ,
    \Tile_X9Y4_WW4BEG[10] ,
    \Tile_X9Y4_WW4BEG[9] ,
    \Tile_X9Y4_WW4BEG[8] ,
    \Tile_X9Y4_WW4BEG[7] ,
    \Tile_X9Y4_WW4BEG[6] ,
    \Tile_X9Y4_WW4BEG[5] ,
    \Tile_X9Y4_WW4BEG[4] ,
    \Tile_X9Y4_WW4BEG[3] ,
    \Tile_X9Y4_WW4BEG[2] ,
    \Tile_X9Y4_WW4BEG[1] ,
    \Tile_X9Y4_WW4BEG[0] }));
 LUT4AB Tile_X8Y5_LUT4AB (.Ci(Tile_X8Y6_Co),
    .Co(Tile_X8Y5_Co),
    .UserCLK(Tile_X8Y6_UserCLKo),
    .UserCLKo(Tile_X8Y5_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X8Y5_E1BEG[3] ,
    \Tile_X8Y5_E1BEG[2] ,
    \Tile_X8Y5_E1BEG[1] ,
    \Tile_X8Y5_E1BEG[0] }),
    .E1END({\Tile_X7Y5_E1BEG[3] ,
    \Tile_X7Y5_E1BEG[2] ,
    \Tile_X7Y5_E1BEG[1] ,
    \Tile_X7Y5_E1BEG[0] }),
    .E2BEG({\Tile_X8Y5_E2BEG[7] ,
    \Tile_X8Y5_E2BEG[6] ,
    \Tile_X8Y5_E2BEG[5] ,
    \Tile_X8Y5_E2BEG[4] ,
    \Tile_X8Y5_E2BEG[3] ,
    \Tile_X8Y5_E2BEG[2] ,
    \Tile_X8Y5_E2BEG[1] ,
    \Tile_X8Y5_E2BEG[0] }),
    .E2BEGb({\Tile_X8Y5_E2BEGb[7] ,
    \Tile_X8Y5_E2BEGb[6] ,
    \Tile_X8Y5_E2BEGb[5] ,
    \Tile_X8Y5_E2BEGb[4] ,
    \Tile_X8Y5_E2BEGb[3] ,
    \Tile_X8Y5_E2BEGb[2] ,
    \Tile_X8Y5_E2BEGb[1] ,
    \Tile_X8Y5_E2BEGb[0] }),
    .E2END({\Tile_X7Y5_E2BEGb[7] ,
    \Tile_X7Y5_E2BEGb[6] ,
    \Tile_X7Y5_E2BEGb[5] ,
    \Tile_X7Y5_E2BEGb[4] ,
    \Tile_X7Y5_E2BEGb[3] ,
    \Tile_X7Y5_E2BEGb[2] ,
    \Tile_X7Y5_E2BEGb[1] ,
    \Tile_X7Y5_E2BEGb[0] }),
    .E2MID({\Tile_X7Y5_E2BEG[7] ,
    \Tile_X7Y5_E2BEG[6] ,
    \Tile_X7Y5_E2BEG[5] ,
    \Tile_X7Y5_E2BEG[4] ,
    \Tile_X7Y5_E2BEG[3] ,
    \Tile_X7Y5_E2BEG[2] ,
    \Tile_X7Y5_E2BEG[1] ,
    \Tile_X7Y5_E2BEG[0] }),
    .E6BEG({\Tile_X8Y5_E6BEG[11] ,
    \Tile_X8Y5_E6BEG[10] ,
    \Tile_X8Y5_E6BEG[9] ,
    \Tile_X8Y5_E6BEG[8] ,
    \Tile_X8Y5_E6BEG[7] ,
    \Tile_X8Y5_E6BEG[6] ,
    \Tile_X8Y5_E6BEG[5] ,
    \Tile_X8Y5_E6BEG[4] ,
    \Tile_X8Y5_E6BEG[3] ,
    \Tile_X8Y5_E6BEG[2] ,
    \Tile_X8Y5_E6BEG[1] ,
    \Tile_X8Y5_E6BEG[0] }),
    .E6END({\Tile_X7Y5_E6BEG[11] ,
    \Tile_X7Y5_E6BEG[10] ,
    \Tile_X7Y5_E6BEG[9] ,
    \Tile_X7Y5_E6BEG[8] ,
    \Tile_X7Y5_E6BEG[7] ,
    \Tile_X7Y5_E6BEG[6] ,
    \Tile_X7Y5_E6BEG[5] ,
    \Tile_X7Y5_E6BEG[4] ,
    \Tile_X7Y5_E6BEG[3] ,
    \Tile_X7Y5_E6BEG[2] ,
    \Tile_X7Y5_E6BEG[1] ,
    \Tile_X7Y5_E6BEG[0] }),
    .EE4BEG({\Tile_X8Y5_EE4BEG[15] ,
    \Tile_X8Y5_EE4BEG[14] ,
    \Tile_X8Y5_EE4BEG[13] ,
    \Tile_X8Y5_EE4BEG[12] ,
    \Tile_X8Y5_EE4BEG[11] ,
    \Tile_X8Y5_EE4BEG[10] ,
    \Tile_X8Y5_EE4BEG[9] ,
    \Tile_X8Y5_EE4BEG[8] ,
    \Tile_X8Y5_EE4BEG[7] ,
    \Tile_X8Y5_EE4BEG[6] ,
    \Tile_X8Y5_EE4BEG[5] ,
    \Tile_X8Y5_EE4BEG[4] ,
    \Tile_X8Y5_EE4BEG[3] ,
    \Tile_X8Y5_EE4BEG[2] ,
    \Tile_X8Y5_EE4BEG[1] ,
    \Tile_X8Y5_EE4BEG[0] }),
    .EE4END({\Tile_X7Y5_EE4BEG[15] ,
    \Tile_X7Y5_EE4BEG[14] ,
    \Tile_X7Y5_EE4BEG[13] ,
    \Tile_X7Y5_EE4BEG[12] ,
    \Tile_X7Y5_EE4BEG[11] ,
    \Tile_X7Y5_EE4BEG[10] ,
    \Tile_X7Y5_EE4BEG[9] ,
    \Tile_X7Y5_EE4BEG[8] ,
    \Tile_X7Y5_EE4BEG[7] ,
    \Tile_X7Y5_EE4BEG[6] ,
    \Tile_X7Y5_EE4BEG[5] ,
    \Tile_X7Y5_EE4BEG[4] ,
    \Tile_X7Y5_EE4BEG[3] ,
    \Tile_X7Y5_EE4BEG[2] ,
    \Tile_X7Y5_EE4BEG[1] ,
    \Tile_X7Y5_EE4BEG[0] }),
    .FrameData({\Tile_X7Y5_FrameData_O[31] ,
    \Tile_X7Y5_FrameData_O[30] ,
    \Tile_X7Y5_FrameData_O[29] ,
    \Tile_X7Y5_FrameData_O[28] ,
    \Tile_X7Y5_FrameData_O[27] ,
    \Tile_X7Y5_FrameData_O[26] ,
    \Tile_X7Y5_FrameData_O[25] ,
    \Tile_X7Y5_FrameData_O[24] ,
    \Tile_X7Y5_FrameData_O[23] ,
    \Tile_X7Y5_FrameData_O[22] ,
    \Tile_X7Y5_FrameData_O[21] ,
    \Tile_X7Y5_FrameData_O[20] ,
    \Tile_X7Y5_FrameData_O[19] ,
    \Tile_X7Y5_FrameData_O[18] ,
    \Tile_X7Y5_FrameData_O[17] ,
    \Tile_X7Y5_FrameData_O[16] ,
    \Tile_X7Y5_FrameData_O[15] ,
    \Tile_X7Y5_FrameData_O[14] ,
    \Tile_X7Y5_FrameData_O[13] ,
    \Tile_X7Y5_FrameData_O[12] ,
    \Tile_X7Y5_FrameData_O[11] ,
    \Tile_X7Y5_FrameData_O[10] ,
    \Tile_X7Y5_FrameData_O[9] ,
    \Tile_X7Y5_FrameData_O[8] ,
    \Tile_X7Y5_FrameData_O[7] ,
    \Tile_X7Y5_FrameData_O[6] ,
    \Tile_X7Y5_FrameData_O[5] ,
    \Tile_X7Y5_FrameData_O[4] ,
    \Tile_X7Y5_FrameData_O[3] ,
    \Tile_X7Y5_FrameData_O[2] ,
    \Tile_X7Y5_FrameData_O[1] ,
    \Tile_X7Y5_FrameData_O[0] }),
    .FrameData_O({\Tile_X8Y5_FrameData_O[31] ,
    \Tile_X8Y5_FrameData_O[30] ,
    \Tile_X8Y5_FrameData_O[29] ,
    \Tile_X8Y5_FrameData_O[28] ,
    \Tile_X8Y5_FrameData_O[27] ,
    \Tile_X8Y5_FrameData_O[26] ,
    \Tile_X8Y5_FrameData_O[25] ,
    \Tile_X8Y5_FrameData_O[24] ,
    \Tile_X8Y5_FrameData_O[23] ,
    \Tile_X8Y5_FrameData_O[22] ,
    \Tile_X8Y5_FrameData_O[21] ,
    \Tile_X8Y5_FrameData_O[20] ,
    \Tile_X8Y5_FrameData_O[19] ,
    \Tile_X8Y5_FrameData_O[18] ,
    \Tile_X8Y5_FrameData_O[17] ,
    \Tile_X8Y5_FrameData_O[16] ,
    \Tile_X8Y5_FrameData_O[15] ,
    \Tile_X8Y5_FrameData_O[14] ,
    \Tile_X8Y5_FrameData_O[13] ,
    \Tile_X8Y5_FrameData_O[12] ,
    \Tile_X8Y5_FrameData_O[11] ,
    \Tile_X8Y5_FrameData_O[10] ,
    \Tile_X8Y5_FrameData_O[9] ,
    \Tile_X8Y5_FrameData_O[8] ,
    \Tile_X8Y5_FrameData_O[7] ,
    \Tile_X8Y5_FrameData_O[6] ,
    \Tile_X8Y5_FrameData_O[5] ,
    \Tile_X8Y5_FrameData_O[4] ,
    \Tile_X8Y5_FrameData_O[3] ,
    \Tile_X8Y5_FrameData_O[2] ,
    \Tile_X8Y5_FrameData_O[1] ,
    \Tile_X8Y5_FrameData_O[0] }),
    .FrameStrobe({\Tile_X8Y6_FrameStrobe_O[19] ,
    \Tile_X8Y6_FrameStrobe_O[18] ,
    \Tile_X8Y6_FrameStrobe_O[17] ,
    \Tile_X8Y6_FrameStrobe_O[16] ,
    \Tile_X8Y6_FrameStrobe_O[15] ,
    \Tile_X8Y6_FrameStrobe_O[14] ,
    \Tile_X8Y6_FrameStrobe_O[13] ,
    \Tile_X8Y6_FrameStrobe_O[12] ,
    \Tile_X8Y6_FrameStrobe_O[11] ,
    \Tile_X8Y6_FrameStrobe_O[10] ,
    \Tile_X8Y6_FrameStrobe_O[9] ,
    \Tile_X8Y6_FrameStrobe_O[8] ,
    \Tile_X8Y6_FrameStrobe_O[7] ,
    \Tile_X8Y6_FrameStrobe_O[6] ,
    \Tile_X8Y6_FrameStrobe_O[5] ,
    \Tile_X8Y6_FrameStrobe_O[4] ,
    \Tile_X8Y6_FrameStrobe_O[3] ,
    \Tile_X8Y6_FrameStrobe_O[2] ,
    \Tile_X8Y6_FrameStrobe_O[1] ,
    \Tile_X8Y6_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X8Y5_FrameStrobe_O[19] ,
    \Tile_X8Y5_FrameStrobe_O[18] ,
    \Tile_X8Y5_FrameStrobe_O[17] ,
    \Tile_X8Y5_FrameStrobe_O[16] ,
    \Tile_X8Y5_FrameStrobe_O[15] ,
    \Tile_X8Y5_FrameStrobe_O[14] ,
    \Tile_X8Y5_FrameStrobe_O[13] ,
    \Tile_X8Y5_FrameStrobe_O[12] ,
    \Tile_X8Y5_FrameStrobe_O[11] ,
    \Tile_X8Y5_FrameStrobe_O[10] ,
    \Tile_X8Y5_FrameStrobe_O[9] ,
    \Tile_X8Y5_FrameStrobe_O[8] ,
    \Tile_X8Y5_FrameStrobe_O[7] ,
    \Tile_X8Y5_FrameStrobe_O[6] ,
    \Tile_X8Y5_FrameStrobe_O[5] ,
    \Tile_X8Y5_FrameStrobe_O[4] ,
    \Tile_X8Y5_FrameStrobe_O[3] ,
    \Tile_X8Y5_FrameStrobe_O[2] ,
    \Tile_X8Y5_FrameStrobe_O[1] ,
    \Tile_X8Y5_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X8Y5_N1BEG[3] ,
    \Tile_X8Y5_N1BEG[2] ,
    \Tile_X8Y5_N1BEG[1] ,
    \Tile_X8Y5_N1BEG[0] }),
    .N1END({\Tile_X8Y6_N1BEG[3] ,
    \Tile_X8Y6_N1BEG[2] ,
    \Tile_X8Y6_N1BEG[1] ,
    \Tile_X8Y6_N1BEG[0] }),
    .N2BEG({\Tile_X8Y5_N2BEG[7] ,
    \Tile_X8Y5_N2BEG[6] ,
    \Tile_X8Y5_N2BEG[5] ,
    \Tile_X8Y5_N2BEG[4] ,
    \Tile_X8Y5_N2BEG[3] ,
    \Tile_X8Y5_N2BEG[2] ,
    \Tile_X8Y5_N2BEG[1] ,
    \Tile_X8Y5_N2BEG[0] }),
    .N2BEGb({\Tile_X8Y5_N2BEGb[7] ,
    \Tile_X8Y5_N2BEGb[6] ,
    \Tile_X8Y5_N2BEGb[5] ,
    \Tile_X8Y5_N2BEGb[4] ,
    \Tile_X8Y5_N2BEGb[3] ,
    \Tile_X8Y5_N2BEGb[2] ,
    \Tile_X8Y5_N2BEGb[1] ,
    \Tile_X8Y5_N2BEGb[0] }),
    .N2END({\Tile_X8Y6_N2BEGb[7] ,
    \Tile_X8Y6_N2BEGb[6] ,
    \Tile_X8Y6_N2BEGb[5] ,
    \Tile_X8Y6_N2BEGb[4] ,
    \Tile_X8Y6_N2BEGb[3] ,
    \Tile_X8Y6_N2BEGb[2] ,
    \Tile_X8Y6_N2BEGb[1] ,
    \Tile_X8Y6_N2BEGb[0] }),
    .N2MID({\Tile_X8Y6_N2BEG[7] ,
    \Tile_X8Y6_N2BEG[6] ,
    \Tile_X8Y6_N2BEG[5] ,
    \Tile_X8Y6_N2BEG[4] ,
    \Tile_X8Y6_N2BEG[3] ,
    \Tile_X8Y6_N2BEG[2] ,
    \Tile_X8Y6_N2BEG[1] ,
    \Tile_X8Y6_N2BEG[0] }),
    .N4BEG({\Tile_X8Y5_N4BEG[15] ,
    \Tile_X8Y5_N4BEG[14] ,
    \Tile_X8Y5_N4BEG[13] ,
    \Tile_X8Y5_N4BEG[12] ,
    \Tile_X8Y5_N4BEG[11] ,
    \Tile_X8Y5_N4BEG[10] ,
    \Tile_X8Y5_N4BEG[9] ,
    \Tile_X8Y5_N4BEG[8] ,
    \Tile_X8Y5_N4BEG[7] ,
    \Tile_X8Y5_N4BEG[6] ,
    \Tile_X8Y5_N4BEG[5] ,
    \Tile_X8Y5_N4BEG[4] ,
    \Tile_X8Y5_N4BEG[3] ,
    \Tile_X8Y5_N4BEG[2] ,
    \Tile_X8Y5_N4BEG[1] ,
    \Tile_X8Y5_N4BEG[0] }),
    .N4END({\Tile_X8Y6_N4BEG[15] ,
    \Tile_X8Y6_N4BEG[14] ,
    \Tile_X8Y6_N4BEG[13] ,
    \Tile_X8Y6_N4BEG[12] ,
    \Tile_X8Y6_N4BEG[11] ,
    \Tile_X8Y6_N4BEG[10] ,
    \Tile_X8Y6_N4BEG[9] ,
    \Tile_X8Y6_N4BEG[8] ,
    \Tile_X8Y6_N4BEG[7] ,
    \Tile_X8Y6_N4BEG[6] ,
    \Tile_X8Y6_N4BEG[5] ,
    \Tile_X8Y6_N4BEG[4] ,
    \Tile_X8Y6_N4BEG[3] ,
    \Tile_X8Y6_N4BEG[2] ,
    \Tile_X8Y6_N4BEG[1] ,
    \Tile_X8Y6_N4BEG[0] }),
    .NN4BEG({\Tile_X8Y5_NN4BEG[15] ,
    \Tile_X8Y5_NN4BEG[14] ,
    \Tile_X8Y5_NN4BEG[13] ,
    \Tile_X8Y5_NN4BEG[12] ,
    \Tile_X8Y5_NN4BEG[11] ,
    \Tile_X8Y5_NN4BEG[10] ,
    \Tile_X8Y5_NN4BEG[9] ,
    \Tile_X8Y5_NN4BEG[8] ,
    \Tile_X8Y5_NN4BEG[7] ,
    \Tile_X8Y5_NN4BEG[6] ,
    \Tile_X8Y5_NN4BEG[5] ,
    \Tile_X8Y5_NN4BEG[4] ,
    \Tile_X8Y5_NN4BEG[3] ,
    \Tile_X8Y5_NN4BEG[2] ,
    \Tile_X8Y5_NN4BEG[1] ,
    \Tile_X8Y5_NN4BEG[0] }),
    .NN4END({\Tile_X8Y6_NN4BEG[15] ,
    \Tile_X8Y6_NN4BEG[14] ,
    \Tile_X8Y6_NN4BEG[13] ,
    \Tile_X8Y6_NN4BEG[12] ,
    \Tile_X8Y6_NN4BEG[11] ,
    \Tile_X8Y6_NN4BEG[10] ,
    \Tile_X8Y6_NN4BEG[9] ,
    \Tile_X8Y6_NN4BEG[8] ,
    \Tile_X8Y6_NN4BEG[7] ,
    \Tile_X8Y6_NN4BEG[6] ,
    \Tile_X8Y6_NN4BEG[5] ,
    \Tile_X8Y6_NN4BEG[4] ,
    \Tile_X8Y6_NN4BEG[3] ,
    \Tile_X8Y6_NN4BEG[2] ,
    \Tile_X8Y6_NN4BEG[1] ,
    \Tile_X8Y6_NN4BEG[0] }),
    .S1BEG({\Tile_X8Y5_S1BEG[3] ,
    \Tile_X8Y5_S1BEG[2] ,
    \Tile_X8Y5_S1BEG[1] ,
    \Tile_X8Y5_S1BEG[0] }),
    .S1END({\Tile_X8Y4_S1BEG[3] ,
    \Tile_X8Y4_S1BEG[2] ,
    \Tile_X8Y4_S1BEG[1] ,
    \Tile_X8Y4_S1BEG[0] }),
    .S2BEG({\Tile_X8Y5_S2BEG[7] ,
    \Tile_X8Y5_S2BEG[6] ,
    \Tile_X8Y5_S2BEG[5] ,
    \Tile_X8Y5_S2BEG[4] ,
    \Tile_X8Y5_S2BEG[3] ,
    \Tile_X8Y5_S2BEG[2] ,
    \Tile_X8Y5_S2BEG[1] ,
    \Tile_X8Y5_S2BEG[0] }),
    .S2BEGb({\Tile_X8Y5_S2BEGb[7] ,
    \Tile_X8Y5_S2BEGb[6] ,
    \Tile_X8Y5_S2BEGb[5] ,
    \Tile_X8Y5_S2BEGb[4] ,
    \Tile_X8Y5_S2BEGb[3] ,
    \Tile_X8Y5_S2BEGb[2] ,
    \Tile_X8Y5_S2BEGb[1] ,
    \Tile_X8Y5_S2BEGb[0] }),
    .S2END({\Tile_X8Y4_S2BEGb[7] ,
    \Tile_X8Y4_S2BEGb[6] ,
    \Tile_X8Y4_S2BEGb[5] ,
    \Tile_X8Y4_S2BEGb[4] ,
    \Tile_X8Y4_S2BEGb[3] ,
    \Tile_X8Y4_S2BEGb[2] ,
    \Tile_X8Y4_S2BEGb[1] ,
    \Tile_X8Y4_S2BEGb[0] }),
    .S2MID({\Tile_X8Y4_S2BEG[7] ,
    \Tile_X8Y4_S2BEG[6] ,
    \Tile_X8Y4_S2BEG[5] ,
    \Tile_X8Y4_S2BEG[4] ,
    \Tile_X8Y4_S2BEG[3] ,
    \Tile_X8Y4_S2BEG[2] ,
    \Tile_X8Y4_S2BEG[1] ,
    \Tile_X8Y4_S2BEG[0] }),
    .S4BEG({\Tile_X8Y5_S4BEG[15] ,
    \Tile_X8Y5_S4BEG[14] ,
    \Tile_X8Y5_S4BEG[13] ,
    \Tile_X8Y5_S4BEG[12] ,
    \Tile_X8Y5_S4BEG[11] ,
    \Tile_X8Y5_S4BEG[10] ,
    \Tile_X8Y5_S4BEG[9] ,
    \Tile_X8Y5_S4BEG[8] ,
    \Tile_X8Y5_S4BEG[7] ,
    \Tile_X8Y5_S4BEG[6] ,
    \Tile_X8Y5_S4BEG[5] ,
    \Tile_X8Y5_S4BEG[4] ,
    \Tile_X8Y5_S4BEG[3] ,
    \Tile_X8Y5_S4BEG[2] ,
    \Tile_X8Y5_S4BEG[1] ,
    \Tile_X8Y5_S4BEG[0] }),
    .S4END({\Tile_X8Y4_S4BEG[15] ,
    \Tile_X8Y4_S4BEG[14] ,
    \Tile_X8Y4_S4BEG[13] ,
    \Tile_X8Y4_S4BEG[12] ,
    \Tile_X8Y4_S4BEG[11] ,
    \Tile_X8Y4_S4BEG[10] ,
    \Tile_X8Y4_S4BEG[9] ,
    \Tile_X8Y4_S4BEG[8] ,
    \Tile_X8Y4_S4BEG[7] ,
    \Tile_X8Y4_S4BEG[6] ,
    \Tile_X8Y4_S4BEG[5] ,
    \Tile_X8Y4_S4BEG[4] ,
    \Tile_X8Y4_S4BEG[3] ,
    \Tile_X8Y4_S4BEG[2] ,
    \Tile_X8Y4_S4BEG[1] ,
    \Tile_X8Y4_S4BEG[0] }),
    .SS4BEG({\Tile_X8Y5_SS4BEG[15] ,
    \Tile_X8Y5_SS4BEG[14] ,
    \Tile_X8Y5_SS4BEG[13] ,
    \Tile_X8Y5_SS4BEG[12] ,
    \Tile_X8Y5_SS4BEG[11] ,
    \Tile_X8Y5_SS4BEG[10] ,
    \Tile_X8Y5_SS4BEG[9] ,
    \Tile_X8Y5_SS4BEG[8] ,
    \Tile_X8Y5_SS4BEG[7] ,
    \Tile_X8Y5_SS4BEG[6] ,
    \Tile_X8Y5_SS4BEG[5] ,
    \Tile_X8Y5_SS4BEG[4] ,
    \Tile_X8Y5_SS4BEG[3] ,
    \Tile_X8Y5_SS4BEG[2] ,
    \Tile_X8Y5_SS4BEG[1] ,
    \Tile_X8Y5_SS4BEG[0] }),
    .SS4END({\Tile_X8Y4_SS4BEG[15] ,
    \Tile_X8Y4_SS4BEG[14] ,
    \Tile_X8Y4_SS4BEG[13] ,
    \Tile_X8Y4_SS4BEG[12] ,
    \Tile_X8Y4_SS4BEG[11] ,
    \Tile_X8Y4_SS4BEG[10] ,
    \Tile_X8Y4_SS4BEG[9] ,
    \Tile_X8Y4_SS4BEG[8] ,
    \Tile_X8Y4_SS4BEG[7] ,
    \Tile_X8Y4_SS4BEG[6] ,
    \Tile_X8Y4_SS4BEG[5] ,
    \Tile_X8Y4_SS4BEG[4] ,
    \Tile_X8Y4_SS4BEG[3] ,
    \Tile_X8Y4_SS4BEG[2] ,
    \Tile_X8Y4_SS4BEG[1] ,
    \Tile_X8Y4_SS4BEG[0] }),
    .W1BEG({\Tile_X8Y5_W1BEG[3] ,
    \Tile_X8Y5_W1BEG[2] ,
    \Tile_X8Y5_W1BEG[1] ,
    \Tile_X8Y5_W1BEG[0] }),
    .W1END({\Tile_X9Y5_W1BEG[3] ,
    \Tile_X9Y5_W1BEG[2] ,
    \Tile_X9Y5_W1BEG[1] ,
    \Tile_X9Y5_W1BEG[0] }),
    .W2BEG({\Tile_X8Y5_W2BEG[7] ,
    \Tile_X8Y5_W2BEG[6] ,
    \Tile_X8Y5_W2BEG[5] ,
    \Tile_X8Y5_W2BEG[4] ,
    \Tile_X8Y5_W2BEG[3] ,
    \Tile_X8Y5_W2BEG[2] ,
    \Tile_X8Y5_W2BEG[1] ,
    \Tile_X8Y5_W2BEG[0] }),
    .W2BEGb({\Tile_X8Y5_W2BEGb[7] ,
    \Tile_X8Y5_W2BEGb[6] ,
    \Tile_X8Y5_W2BEGb[5] ,
    \Tile_X8Y5_W2BEGb[4] ,
    \Tile_X8Y5_W2BEGb[3] ,
    \Tile_X8Y5_W2BEGb[2] ,
    \Tile_X8Y5_W2BEGb[1] ,
    \Tile_X8Y5_W2BEGb[0] }),
    .W2END({\Tile_X9Y5_W2BEGb[7] ,
    \Tile_X9Y5_W2BEGb[6] ,
    \Tile_X9Y5_W2BEGb[5] ,
    \Tile_X9Y5_W2BEGb[4] ,
    \Tile_X9Y5_W2BEGb[3] ,
    \Tile_X9Y5_W2BEGb[2] ,
    \Tile_X9Y5_W2BEGb[1] ,
    \Tile_X9Y5_W2BEGb[0] }),
    .W2MID({\Tile_X9Y5_W2BEG[7] ,
    \Tile_X9Y5_W2BEG[6] ,
    \Tile_X9Y5_W2BEG[5] ,
    \Tile_X9Y5_W2BEG[4] ,
    \Tile_X9Y5_W2BEG[3] ,
    \Tile_X9Y5_W2BEG[2] ,
    \Tile_X9Y5_W2BEG[1] ,
    \Tile_X9Y5_W2BEG[0] }),
    .W6BEG({\Tile_X8Y5_W6BEG[11] ,
    \Tile_X8Y5_W6BEG[10] ,
    \Tile_X8Y5_W6BEG[9] ,
    \Tile_X8Y5_W6BEG[8] ,
    \Tile_X8Y5_W6BEG[7] ,
    \Tile_X8Y5_W6BEG[6] ,
    \Tile_X8Y5_W6BEG[5] ,
    \Tile_X8Y5_W6BEG[4] ,
    \Tile_X8Y5_W6BEG[3] ,
    \Tile_X8Y5_W6BEG[2] ,
    \Tile_X8Y5_W6BEG[1] ,
    \Tile_X8Y5_W6BEG[0] }),
    .W6END({\Tile_X9Y5_W6BEG[11] ,
    \Tile_X9Y5_W6BEG[10] ,
    \Tile_X9Y5_W6BEG[9] ,
    \Tile_X9Y5_W6BEG[8] ,
    \Tile_X9Y5_W6BEG[7] ,
    \Tile_X9Y5_W6BEG[6] ,
    \Tile_X9Y5_W6BEG[5] ,
    \Tile_X9Y5_W6BEG[4] ,
    \Tile_X9Y5_W6BEG[3] ,
    \Tile_X9Y5_W6BEG[2] ,
    \Tile_X9Y5_W6BEG[1] ,
    \Tile_X9Y5_W6BEG[0] }),
    .WW4BEG({\Tile_X8Y5_WW4BEG[15] ,
    \Tile_X8Y5_WW4BEG[14] ,
    \Tile_X8Y5_WW4BEG[13] ,
    \Tile_X8Y5_WW4BEG[12] ,
    \Tile_X8Y5_WW4BEG[11] ,
    \Tile_X8Y5_WW4BEG[10] ,
    \Tile_X8Y5_WW4BEG[9] ,
    \Tile_X8Y5_WW4BEG[8] ,
    \Tile_X8Y5_WW4BEG[7] ,
    \Tile_X8Y5_WW4BEG[6] ,
    \Tile_X8Y5_WW4BEG[5] ,
    \Tile_X8Y5_WW4BEG[4] ,
    \Tile_X8Y5_WW4BEG[3] ,
    \Tile_X8Y5_WW4BEG[2] ,
    \Tile_X8Y5_WW4BEG[1] ,
    \Tile_X8Y5_WW4BEG[0] }),
    .WW4END({\Tile_X9Y5_WW4BEG[15] ,
    \Tile_X9Y5_WW4BEG[14] ,
    \Tile_X9Y5_WW4BEG[13] ,
    \Tile_X9Y5_WW4BEG[12] ,
    \Tile_X9Y5_WW4BEG[11] ,
    \Tile_X9Y5_WW4BEG[10] ,
    \Tile_X9Y5_WW4BEG[9] ,
    \Tile_X9Y5_WW4BEG[8] ,
    \Tile_X9Y5_WW4BEG[7] ,
    \Tile_X9Y5_WW4BEG[6] ,
    \Tile_X9Y5_WW4BEG[5] ,
    \Tile_X9Y5_WW4BEG[4] ,
    \Tile_X9Y5_WW4BEG[3] ,
    \Tile_X9Y5_WW4BEG[2] ,
    \Tile_X9Y5_WW4BEG[1] ,
    \Tile_X9Y5_WW4BEG[0] }));
 LUT4AB Tile_X8Y6_LUT4AB (.Ci(Tile_X8Y7_Co),
    .Co(Tile_X8Y6_Co),
    .UserCLK(Tile_X8Y7_UserCLKo),
    .UserCLKo(Tile_X8Y6_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X8Y6_E1BEG[3] ,
    \Tile_X8Y6_E1BEG[2] ,
    \Tile_X8Y6_E1BEG[1] ,
    \Tile_X8Y6_E1BEG[0] }),
    .E1END({\Tile_X7Y6_E1BEG[3] ,
    \Tile_X7Y6_E1BEG[2] ,
    \Tile_X7Y6_E1BEG[1] ,
    \Tile_X7Y6_E1BEG[0] }),
    .E2BEG({\Tile_X8Y6_E2BEG[7] ,
    \Tile_X8Y6_E2BEG[6] ,
    \Tile_X8Y6_E2BEG[5] ,
    \Tile_X8Y6_E2BEG[4] ,
    \Tile_X8Y6_E2BEG[3] ,
    \Tile_X8Y6_E2BEG[2] ,
    \Tile_X8Y6_E2BEG[1] ,
    \Tile_X8Y6_E2BEG[0] }),
    .E2BEGb({\Tile_X8Y6_E2BEGb[7] ,
    \Tile_X8Y6_E2BEGb[6] ,
    \Tile_X8Y6_E2BEGb[5] ,
    \Tile_X8Y6_E2BEGb[4] ,
    \Tile_X8Y6_E2BEGb[3] ,
    \Tile_X8Y6_E2BEGb[2] ,
    \Tile_X8Y6_E2BEGb[1] ,
    \Tile_X8Y6_E2BEGb[0] }),
    .E2END({\Tile_X7Y6_E2BEGb[7] ,
    \Tile_X7Y6_E2BEGb[6] ,
    \Tile_X7Y6_E2BEGb[5] ,
    \Tile_X7Y6_E2BEGb[4] ,
    \Tile_X7Y6_E2BEGb[3] ,
    \Tile_X7Y6_E2BEGb[2] ,
    \Tile_X7Y6_E2BEGb[1] ,
    \Tile_X7Y6_E2BEGb[0] }),
    .E2MID({\Tile_X7Y6_E2BEG[7] ,
    \Tile_X7Y6_E2BEG[6] ,
    \Tile_X7Y6_E2BEG[5] ,
    \Tile_X7Y6_E2BEG[4] ,
    \Tile_X7Y6_E2BEG[3] ,
    \Tile_X7Y6_E2BEG[2] ,
    \Tile_X7Y6_E2BEG[1] ,
    \Tile_X7Y6_E2BEG[0] }),
    .E6BEG({\Tile_X8Y6_E6BEG[11] ,
    \Tile_X8Y6_E6BEG[10] ,
    \Tile_X8Y6_E6BEG[9] ,
    \Tile_X8Y6_E6BEG[8] ,
    \Tile_X8Y6_E6BEG[7] ,
    \Tile_X8Y6_E6BEG[6] ,
    \Tile_X8Y6_E6BEG[5] ,
    \Tile_X8Y6_E6BEG[4] ,
    \Tile_X8Y6_E6BEG[3] ,
    \Tile_X8Y6_E6BEG[2] ,
    \Tile_X8Y6_E6BEG[1] ,
    \Tile_X8Y6_E6BEG[0] }),
    .E6END({\Tile_X7Y6_E6BEG[11] ,
    \Tile_X7Y6_E6BEG[10] ,
    \Tile_X7Y6_E6BEG[9] ,
    \Tile_X7Y6_E6BEG[8] ,
    \Tile_X7Y6_E6BEG[7] ,
    \Tile_X7Y6_E6BEG[6] ,
    \Tile_X7Y6_E6BEG[5] ,
    \Tile_X7Y6_E6BEG[4] ,
    \Tile_X7Y6_E6BEG[3] ,
    \Tile_X7Y6_E6BEG[2] ,
    \Tile_X7Y6_E6BEG[1] ,
    \Tile_X7Y6_E6BEG[0] }),
    .EE4BEG({\Tile_X8Y6_EE4BEG[15] ,
    \Tile_X8Y6_EE4BEG[14] ,
    \Tile_X8Y6_EE4BEG[13] ,
    \Tile_X8Y6_EE4BEG[12] ,
    \Tile_X8Y6_EE4BEG[11] ,
    \Tile_X8Y6_EE4BEG[10] ,
    \Tile_X8Y6_EE4BEG[9] ,
    \Tile_X8Y6_EE4BEG[8] ,
    \Tile_X8Y6_EE4BEG[7] ,
    \Tile_X8Y6_EE4BEG[6] ,
    \Tile_X8Y6_EE4BEG[5] ,
    \Tile_X8Y6_EE4BEG[4] ,
    \Tile_X8Y6_EE4BEG[3] ,
    \Tile_X8Y6_EE4BEG[2] ,
    \Tile_X8Y6_EE4BEG[1] ,
    \Tile_X8Y6_EE4BEG[0] }),
    .EE4END({\Tile_X7Y6_EE4BEG[15] ,
    \Tile_X7Y6_EE4BEG[14] ,
    \Tile_X7Y6_EE4BEG[13] ,
    \Tile_X7Y6_EE4BEG[12] ,
    \Tile_X7Y6_EE4BEG[11] ,
    \Tile_X7Y6_EE4BEG[10] ,
    \Tile_X7Y6_EE4BEG[9] ,
    \Tile_X7Y6_EE4BEG[8] ,
    \Tile_X7Y6_EE4BEG[7] ,
    \Tile_X7Y6_EE4BEG[6] ,
    \Tile_X7Y6_EE4BEG[5] ,
    \Tile_X7Y6_EE4BEG[4] ,
    \Tile_X7Y6_EE4BEG[3] ,
    \Tile_X7Y6_EE4BEG[2] ,
    \Tile_X7Y6_EE4BEG[1] ,
    \Tile_X7Y6_EE4BEG[0] }),
    .FrameData({\Tile_X7Y6_FrameData_O[31] ,
    \Tile_X7Y6_FrameData_O[30] ,
    \Tile_X7Y6_FrameData_O[29] ,
    \Tile_X7Y6_FrameData_O[28] ,
    \Tile_X7Y6_FrameData_O[27] ,
    \Tile_X7Y6_FrameData_O[26] ,
    \Tile_X7Y6_FrameData_O[25] ,
    \Tile_X7Y6_FrameData_O[24] ,
    \Tile_X7Y6_FrameData_O[23] ,
    \Tile_X7Y6_FrameData_O[22] ,
    \Tile_X7Y6_FrameData_O[21] ,
    \Tile_X7Y6_FrameData_O[20] ,
    \Tile_X7Y6_FrameData_O[19] ,
    \Tile_X7Y6_FrameData_O[18] ,
    \Tile_X7Y6_FrameData_O[17] ,
    \Tile_X7Y6_FrameData_O[16] ,
    \Tile_X7Y6_FrameData_O[15] ,
    \Tile_X7Y6_FrameData_O[14] ,
    \Tile_X7Y6_FrameData_O[13] ,
    \Tile_X7Y6_FrameData_O[12] ,
    \Tile_X7Y6_FrameData_O[11] ,
    \Tile_X7Y6_FrameData_O[10] ,
    \Tile_X7Y6_FrameData_O[9] ,
    \Tile_X7Y6_FrameData_O[8] ,
    \Tile_X7Y6_FrameData_O[7] ,
    \Tile_X7Y6_FrameData_O[6] ,
    \Tile_X7Y6_FrameData_O[5] ,
    \Tile_X7Y6_FrameData_O[4] ,
    \Tile_X7Y6_FrameData_O[3] ,
    \Tile_X7Y6_FrameData_O[2] ,
    \Tile_X7Y6_FrameData_O[1] ,
    \Tile_X7Y6_FrameData_O[0] }),
    .FrameData_O({\Tile_X8Y6_FrameData_O[31] ,
    \Tile_X8Y6_FrameData_O[30] ,
    \Tile_X8Y6_FrameData_O[29] ,
    \Tile_X8Y6_FrameData_O[28] ,
    \Tile_X8Y6_FrameData_O[27] ,
    \Tile_X8Y6_FrameData_O[26] ,
    \Tile_X8Y6_FrameData_O[25] ,
    \Tile_X8Y6_FrameData_O[24] ,
    \Tile_X8Y6_FrameData_O[23] ,
    \Tile_X8Y6_FrameData_O[22] ,
    \Tile_X8Y6_FrameData_O[21] ,
    \Tile_X8Y6_FrameData_O[20] ,
    \Tile_X8Y6_FrameData_O[19] ,
    \Tile_X8Y6_FrameData_O[18] ,
    \Tile_X8Y6_FrameData_O[17] ,
    \Tile_X8Y6_FrameData_O[16] ,
    \Tile_X8Y6_FrameData_O[15] ,
    \Tile_X8Y6_FrameData_O[14] ,
    \Tile_X8Y6_FrameData_O[13] ,
    \Tile_X8Y6_FrameData_O[12] ,
    \Tile_X8Y6_FrameData_O[11] ,
    \Tile_X8Y6_FrameData_O[10] ,
    \Tile_X8Y6_FrameData_O[9] ,
    \Tile_X8Y6_FrameData_O[8] ,
    \Tile_X8Y6_FrameData_O[7] ,
    \Tile_X8Y6_FrameData_O[6] ,
    \Tile_X8Y6_FrameData_O[5] ,
    \Tile_X8Y6_FrameData_O[4] ,
    \Tile_X8Y6_FrameData_O[3] ,
    \Tile_X8Y6_FrameData_O[2] ,
    \Tile_X8Y6_FrameData_O[1] ,
    \Tile_X8Y6_FrameData_O[0] }),
    .FrameStrobe({\Tile_X8Y7_FrameStrobe_O[19] ,
    \Tile_X8Y7_FrameStrobe_O[18] ,
    \Tile_X8Y7_FrameStrobe_O[17] ,
    \Tile_X8Y7_FrameStrobe_O[16] ,
    \Tile_X8Y7_FrameStrobe_O[15] ,
    \Tile_X8Y7_FrameStrobe_O[14] ,
    \Tile_X8Y7_FrameStrobe_O[13] ,
    \Tile_X8Y7_FrameStrobe_O[12] ,
    \Tile_X8Y7_FrameStrobe_O[11] ,
    \Tile_X8Y7_FrameStrobe_O[10] ,
    \Tile_X8Y7_FrameStrobe_O[9] ,
    \Tile_X8Y7_FrameStrobe_O[8] ,
    \Tile_X8Y7_FrameStrobe_O[7] ,
    \Tile_X8Y7_FrameStrobe_O[6] ,
    \Tile_X8Y7_FrameStrobe_O[5] ,
    \Tile_X8Y7_FrameStrobe_O[4] ,
    \Tile_X8Y7_FrameStrobe_O[3] ,
    \Tile_X8Y7_FrameStrobe_O[2] ,
    \Tile_X8Y7_FrameStrobe_O[1] ,
    \Tile_X8Y7_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X8Y6_FrameStrobe_O[19] ,
    \Tile_X8Y6_FrameStrobe_O[18] ,
    \Tile_X8Y6_FrameStrobe_O[17] ,
    \Tile_X8Y6_FrameStrobe_O[16] ,
    \Tile_X8Y6_FrameStrobe_O[15] ,
    \Tile_X8Y6_FrameStrobe_O[14] ,
    \Tile_X8Y6_FrameStrobe_O[13] ,
    \Tile_X8Y6_FrameStrobe_O[12] ,
    \Tile_X8Y6_FrameStrobe_O[11] ,
    \Tile_X8Y6_FrameStrobe_O[10] ,
    \Tile_X8Y6_FrameStrobe_O[9] ,
    \Tile_X8Y6_FrameStrobe_O[8] ,
    \Tile_X8Y6_FrameStrobe_O[7] ,
    \Tile_X8Y6_FrameStrobe_O[6] ,
    \Tile_X8Y6_FrameStrobe_O[5] ,
    \Tile_X8Y6_FrameStrobe_O[4] ,
    \Tile_X8Y6_FrameStrobe_O[3] ,
    \Tile_X8Y6_FrameStrobe_O[2] ,
    \Tile_X8Y6_FrameStrobe_O[1] ,
    \Tile_X8Y6_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X8Y6_N1BEG[3] ,
    \Tile_X8Y6_N1BEG[2] ,
    \Tile_X8Y6_N1BEG[1] ,
    \Tile_X8Y6_N1BEG[0] }),
    .N1END({\Tile_X8Y7_N1BEG[3] ,
    \Tile_X8Y7_N1BEG[2] ,
    \Tile_X8Y7_N1BEG[1] ,
    \Tile_X8Y7_N1BEG[0] }),
    .N2BEG({\Tile_X8Y6_N2BEG[7] ,
    \Tile_X8Y6_N2BEG[6] ,
    \Tile_X8Y6_N2BEG[5] ,
    \Tile_X8Y6_N2BEG[4] ,
    \Tile_X8Y6_N2BEG[3] ,
    \Tile_X8Y6_N2BEG[2] ,
    \Tile_X8Y6_N2BEG[1] ,
    \Tile_X8Y6_N2BEG[0] }),
    .N2BEGb({\Tile_X8Y6_N2BEGb[7] ,
    \Tile_X8Y6_N2BEGb[6] ,
    \Tile_X8Y6_N2BEGb[5] ,
    \Tile_X8Y6_N2BEGb[4] ,
    \Tile_X8Y6_N2BEGb[3] ,
    \Tile_X8Y6_N2BEGb[2] ,
    \Tile_X8Y6_N2BEGb[1] ,
    \Tile_X8Y6_N2BEGb[0] }),
    .N2END({\Tile_X8Y7_N2BEGb[7] ,
    \Tile_X8Y7_N2BEGb[6] ,
    \Tile_X8Y7_N2BEGb[5] ,
    \Tile_X8Y7_N2BEGb[4] ,
    \Tile_X8Y7_N2BEGb[3] ,
    \Tile_X8Y7_N2BEGb[2] ,
    \Tile_X8Y7_N2BEGb[1] ,
    \Tile_X8Y7_N2BEGb[0] }),
    .N2MID({\Tile_X8Y7_N2BEG[7] ,
    \Tile_X8Y7_N2BEG[6] ,
    \Tile_X8Y7_N2BEG[5] ,
    \Tile_X8Y7_N2BEG[4] ,
    \Tile_X8Y7_N2BEG[3] ,
    \Tile_X8Y7_N2BEG[2] ,
    \Tile_X8Y7_N2BEG[1] ,
    \Tile_X8Y7_N2BEG[0] }),
    .N4BEG({\Tile_X8Y6_N4BEG[15] ,
    \Tile_X8Y6_N4BEG[14] ,
    \Tile_X8Y6_N4BEG[13] ,
    \Tile_X8Y6_N4BEG[12] ,
    \Tile_X8Y6_N4BEG[11] ,
    \Tile_X8Y6_N4BEG[10] ,
    \Tile_X8Y6_N4BEG[9] ,
    \Tile_X8Y6_N4BEG[8] ,
    \Tile_X8Y6_N4BEG[7] ,
    \Tile_X8Y6_N4BEG[6] ,
    \Tile_X8Y6_N4BEG[5] ,
    \Tile_X8Y6_N4BEG[4] ,
    \Tile_X8Y6_N4BEG[3] ,
    \Tile_X8Y6_N4BEG[2] ,
    \Tile_X8Y6_N4BEG[1] ,
    \Tile_X8Y6_N4BEG[0] }),
    .N4END({\Tile_X8Y7_N4BEG[15] ,
    \Tile_X8Y7_N4BEG[14] ,
    \Tile_X8Y7_N4BEG[13] ,
    \Tile_X8Y7_N4BEG[12] ,
    \Tile_X8Y7_N4BEG[11] ,
    \Tile_X8Y7_N4BEG[10] ,
    \Tile_X8Y7_N4BEG[9] ,
    \Tile_X8Y7_N4BEG[8] ,
    \Tile_X8Y7_N4BEG[7] ,
    \Tile_X8Y7_N4BEG[6] ,
    \Tile_X8Y7_N4BEG[5] ,
    \Tile_X8Y7_N4BEG[4] ,
    \Tile_X8Y7_N4BEG[3] ,
    \Tile_X8Y7_N4BEG[2] ,
    \Tile_X8Y7_N4BEG[1] ,
    \Tile_X8Y7_N4BEG[0] }),
    .NN4BEG({\Tile_X8Y6_NN4BEG[15] ,
    \Tile_X8Y6_NN4BEG[14] ,
    \Tile_X8Y6_NN4BEG[13] ,
    \Tile_X8Y6_NN4BEG[12] ,
    \Tile_X8Y6_NN4BEG[11] ,
    \Tile_X8Y6_NN4BEG[10] ,
    \Tile_X8Y6_NN4BEG[9] ,
    \Tile_X8Y6_NN4BEG[8] ,
    \Tile_X8Y6_NN4BEG[7] ,
    \Tile_X8Y6_NN4BEG[6] ,
    \Tile_X8Y6_NN4BEG[5] ,
    \Tile_X8Y6_NN4BEG[4] ,
    \Tile_X8Y6_NN4BEG[3] ,
    \Tile_X8Y6_NN4BEG[2] ,
    \Tile_X8Y6_NN4BEG[1] ,
    \Tile_X8Y6_NN4BEG[0] }),
    .NN4END({\Tile_X8Y7_NN4BEG[15] ,
    \Tile_X8Y7_NN4BEG[14] ,
    \Tile_X8Y7_NN4BEG[13] ,
    \Tile_X8Y7_NN4BEG[12] ,
    \Tile_X8Y7_NN4BEG[11] ,
    \Tile_X8Y7_NN4BEG[10] ,
    \Tile_X8Y7_NN4BEG[9] ,
    \Tile_X8Y7_NN4BEG[8] ,
    \Tile_X8Y7_NN4BEG[7] ,
    \Tile_X8Y7_NN4BEG[6] ,
    \Tile_X8Y7_NN4BEG[5] ,
    \Tile_X8Y7_NN4BEG[4] ,
    \Tile_X8Y7_NN4BEG[3] ,
    \Tile_X8Y7_NN4BEG[2] ,
    \Tile_X8Y7_NN4BEG[1] ,
    \Tile_X8Y7_NN4BEG[0] }),
    .S1BEG({\Tile_X8Y6_S1BEG[3] ,
    \Tile_X8Y6_S1BEG[2] ,
    \Tile_X8Y6_S1BEG[1] ,
    \Tile_X8Y6_S1BEG[0] }),
    .S1END({\Tile_X8Y5_S1BEG[3] ,
    \Tile_X8Y5_S1BEG[2] ,
    \Tile_X8Y5_S1BEG[1] ,
    \Tile_X8Y5_S1BEG[0] }),
    .S2BEG({\Tile_X8Y6_S2BEG[7] ,
    \Tile_X8Y6_S2BEG[6] ,
    \Tile_X8Y6_S2BEG[5] ,
    \Tile_X8Y6_S2BEG[4] ,
    \Tile_X8Y6_S2BEG[3] ,
    \Tile_X8Y6_S2BEG[2] ,
    \Tile_X8Y6_S2BEG[1] ,
    \Tile_X8Y6_S2BEG[0] }),
    .S2BEGb({\Tile_X8Y6_S2BEGb[7] ,
    \Tile_X8Y6_S2BEGb[6] ,
    \Tile_X8Y6_S2BEGb[5] ,
    \Tile_X8Y6_S2BEGb[4] ,
    \Tile_X8Y6_S2BEGb[3] ,
    \Tile_X8Y6_S2BEGb[2] ,
    \Tile_X8Y6_S2BEGb[1] ,
    \Tile_X8Y6_S2BEGb[0] }),
    .S2END({\Tile_X8Y5_S2BEGb[7] ,
    \Tile_X8Y5_S2BEGb[6] ,
    \Tile_X8Y5_S2BEGb[5] ,
    \Tile_X8Y5_S2BEGb[4] ,
    \Tile_X8Y5_S2BEGb[3] ,
    \Tile_X8Y5_S2BEGb[2] ,
    \Tile_X8Y5_S2BEGb[1] ,
    \Tile_X8Y5_S2BEGb[0] }),
    .S2MID({\Tile_X8Y5_S2BEG[7] ,
    \Tile_X8Y5_S2BEG[6] ,
    \Tile_X8Y5_S2BEG[5] ,
    \Tile_X8Y5_S2BEG[4] ,
    \Tile_X8Y5_S2BEG[3] ,
    \Tile_X8Y5_S2BEG[2] ,
    \Tile_X8Y5_S2BEG[1] ,
    \Tile_X8Y5_S2BEG[0] }),
    .S4BEG({\Tile_X8Y6_S4BEG[15] ,
    \Tile_X8Y6_S4BEG[14] ,
    \Tile_X8Y6_S4BEG[13] ,
    \Tile_X8Y6_S4BEG[12] ,
    \Tile_X8Y6_S4BEG[11] ,
    \Tile_X8Y6_S4BEG[10] ,
    \Tile_X8Y6_S4BEG[9] ,
    \Tile_X8Y6_S4BEG[8] ,
    \Tile_X8Y6_S4BEG[7] ,
    \Tile_X8Y6_S4BEG[6] ,
    \Tile_X8Y6_S4BEG[5] ,
    \Tile_X8Y6_S4BEG[4] ,
    \Tile_X8Y6_S4BEG[3] ,
    \Tile_X8Y6_S4BEG[2] ,
    \Tile_X8Y6_S4BEG[1] ,
    \Tile_X8Y6_S4BEG[0] }),
    .S4END({\Tile_X8Y5_S4BEG[15] ,
    \Tile_X8Y5_S4BEG[14] ,
    \Tile_X8Y5_S4BEG[13] ,
    \Tile_X8Y5_S4BEG[12] ,
    \Tile_X8Y5_S4BEG[11] ,
    \Tile_X8Y5_S4BEG[10] ,
    \Tile_X8Y5_S4BEG[9] ,
    \Tile_X8Y5_S4BEG[8] ,
    \Tile_X8Y5_S4BEG[7] ,
    \Tile_X8Y5_S4BEG[6] ,
    \Tile_X8Y5_S4BEG[5] ,
    \Tile_X8Y5_S4BEG[4] ,
    \Tile_X8Y5_S4BEG[3] ,
    \Tile_X8Y5_S4BEG[2] ,
    \Tile_X8Y5_S4BEG[1] ,
    \Tile_X8Y5_S4BEG[0] }),
    .SS4BEG({\Tile_X8Y6_SS4BEG[15] ,
    \Tile_X8Y6_SS4BEG[14] ,
    \Tile_X8Y6_SS4BEG[13] ,
    \Tile_X8Y6_SS4BEG[12] ,
    \Tile_X8Y6_SS4BEG[11] ,
    \Tile_X8Y6_SS4BEG[10] ,
    \Tile_X8Y6_SS4BEG[9] ,
    \Tile_X8Y6_SS4BEG[8] ,
    \Tile_X8Y6_SS4BEG[7] ,
    \Tile_X8Y6_SS4BEG[6] ,
    \Tile_X8Y6_SS4BEG[5] ,
    \Tile_X8Y6_SS4BEG[4] ,
    \Tile_X8Y6_SS4BEG[3] ,
    \Tile_X8Y6_SS4BEG[2] ,
    \Tile_X8Y6_SS4BEG[1] ,
    \Tile_X8Y6_SS4BEG[0] }),
    .SS4END({\Tile_X8Y5_SS4BEG[15] ,
    \Tile_X8Y5_SS4BEG[14] ,
    \Tile_X8Y5_SS4BEG[13] ,
    \Tile_X8Y5_SS4BEG[12] ,
    \Tile_X8Y5_SS4BEG[11] ,
    \Tile_X8Y5_SS4BEG[10] ,
    \Tile_X8Y5_SS4BEG[9] ,
    \Tile_X8Y5_SS4BEG[8] ,
    \Tile_X8Y5_SS4BEG[7] ,
    \Tile_X8Y5_SS4BEG[6] ,
    \Tile_X8Y5_SS4BEG[5] ,
    \Tile_X8Y5_SS4BEG[4] ,
    \Tile_X8Y5_SS4BEG[3] ,
    \Tile_X8Y5_SS4BEG[2] ,
    \Tile_X8Y5_SS4BEG[1] ,
    \Tile_X8Y5_SS4BEG[0] }),
    .W1BEG({\Tile_X8Y6_W1BEG[3] ,
    \Tile_X8Y6_W1BEG[2] ,
    \Tile_X8Y6_W1BEG[1] ,
    \Tile_X8Y6_W1BEG[0] }),
    .W1END({\Tile_X9Y6_W1BEG[3] ,
    \Tile_X9Y6_W1BEG[2] ,
    \Tile_X9Y6_W1BEG[1] ,
    \Tile_X9Y6_W1BEG[0] }),
    .W2BEG({\Tile_X8Y6_W2BEG[7] ,
    \Tile_X8Y6_W2BEG[6] ,
    \Tile_X8Y6_W2BEG[5] ,
    \Tile_X8Y6_W2BEG[4] ,
    \Tile_X8Y6_W2BEG[3] ,
    \Tile_X8Y6_W2BEG[2] ,
    \Tile_X8Y6_W2BEG[1] ,
    \Tile_X8Y6_W2BEG[0] }),
    .W2BEGb({\Tile_X8Y6_W2BEGb[7] ,
    \Tile_X8Y6_W2BEGb[6] ,
    \Tile_X8Y6_W2BEGb[5] ,
    \Tile_X8Y6_W2BEGb[4] ,
    \Tile_X8Y6_W2BEGb[3] ,
    \Tile_X8Y6_W2BEGb[2] ,
    \Tile_X8Y6_W2BEGb[1] ,
    \Tile_X8Y6_W2BEGb[0] }),
    .W2END({\Tile_X9Y6_W2BEGb[7] ,
    \Tile_X9Y6_W2BEGb[6] ,
    \Tile_X9Y6_W2BEGb[5] ,
    \Tile_X9Y6_W2BEGb[4] ,
    \Tile_X9Y6_W2BEGb[3] ,
    \Tile_X9Y6_W2BEGb[2] ,
    \Tile_X9Y6_W2BEGb[1] ,
    \Tile_X9Y6_W2BEGb[0] }),
    .W2MID({\Tile_X9Y6_W2BEG[7] ,
    \Tile_X9Y6_W2BEG[6] ,
    \Tile_X9Y6_W2BEG[5] ,
    \Tile_X9Y6_W2BEG[4] ,
    \Tile_X9Y6_W2BEG[3] ,
    \Tile_X9Y6_W2BEG[2] ,
    \Tile_X9Y6_W2BEG[1] ,
    \Tile_X9Y6_W2BEG[0] }),
    .W6BEG({\Tile_X8Y6_W6BEG[11] ,
    \Tile_X8Y6_W6BEG[10] ,
    \Tile_X8Y6_W6BEG[9] ,
    \Tile_X8Y6_W6BEG[8] ,
    \Tile_X8Y6_W6BEG[7] ,
    \Tile_X8Y6_W6BEG[6] ,
    \Tile_X8Y6_W6BEG[5] ,
    \Tile_X8Y6_W6BEG[4] ,
    \Tile_X8Y6_W6BEG[3] ,
    \Tile_X8Y6_W6BEG[2] ,
    \Tile_X8Y6_W6BEG[1] ,
    \Tile_X8Y6_W6BEG[0] }),
    .W6END({\Tile_X9Y6_W6BEG[11] ,
    \Tile_X9Y6_W6BEG[10] ,
    \Tile_X9Y6_W6BEG[9] ,
    \Tile_X9Y6_W6BEG[8] ,
    \Tile_X9Y6_W6BEG[7] ,
    \Tile_X9Y6_W6BEG[6] ,
    \Tile_X9Y6_W6BEG[5] ,
    \Tile_X9Y6_W6BEG[4] ,
    \Tile_X9Y6_W6BEG[3] ,
    \Tile_X9Y6_W6BEG[2] ,
    \Tile_X9Y6_W6BEG[1] ,
    \Tile_X9Y6_W6BEG[0] }),
    .WW4BEG({\Tile_X8Y6_WW4BEG[15] ,
    \Tile_X8Y6_WW4BEG[14] ,
    \Tile_X8Y6_WW4BEG[13] ,
    \Tile_X8Y6_WW4BEG[12] ,
    \Tile_X8Y6_WW4BEG[11] ,
    \Tile_X8Y6_WW4BEG[10] ,
    \Tile_X8Y6_WW4BEG[9] ,
    \Tile_X8Y6_WW4BEG[8] ,
    \Tile_X8Y6_WW4BEG[7] ,
    \Tile_X8Y6_WW4BEG[6] ,
    \Tile_X8Y6_WW4BEG[5] ,
    \Tile_X8Y6_WW4BEG[4] ,
    \Tile_X8Y6_WW4BEG[3] ,
    \Tile_X8Y6_WW4BEG[2] ,
    \Tile_X8Y6_WW4BEG[1] ,
    \Tile_X8Y6_WW4BEG[0] }),
    .WW4END({\Tile_X9Y6_WW4BEG[15] ,
    \Tile_X9Y6_WW4BEG[14] ,
    \Tile_X9Y6_WW4BEG[13] ,
    \Tile_X9Y6_WW4BEG[12] ,
    \Tile_X9Y6_WW4BEG[11] ,
    \Tile_X9Y6_WW4BEG[10] ,
    \Tile_X9Y6_WW4BEG[9] ,
    \Tile_X9Y6_WW4BEG[8] ,
    \Tile_X9Y6_WW4BEG[7] ,
    \Tile_X9Y6_WW4BEG[6] ,
    \Tile_X9Y6_WW4BEG[5] ,
    \Tile_X9Y6_WW4BEG[4] ,
    \Tile_X9Y6_WW4BEG[3] ,
    \Tile_X9Y6_WW4BEG[2] ,
    \Tile_X9Y6_WW4BEG[1] ,
    \Tile_X9Y6_WW4BEG[0] }));
 LUT4AB Tile_X8Y7_LUT4AB (.Ci(Tile_X8Y8_Co),
    .Co(Tile_X8Y7_Co),
    .UserCLK(Tile_X8Y8_UserCLKo),
    .UserCLKo(Tile_X8Y7_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X8Y7_E1BEG[3] ,
    \Tile_X8Y7_E1BEG[2] ,
    \Tile_X8Y7_E1BEG[1] ,
    \Tile_X8Y7_E1BEG[0] }),
    .E1END({\Tile_X7Y7_E1BEG[3] ,
    \Tile_X7Y7_E1BEG[2] ,
    \Tile_X7Y7_E1BEG[1] ,
    \Tile_X7Y7_E1BEG[0] }),
    .E2BEG({\Tile_X8Y7_E2BEG[7] ,
    \Tile_X8Y7_E2BEG[6] ,
    \Tile_X8Y7_E2BEG[5] ,
    \Tile_X8Y7_E2BEG[4] ,
    \Tile_X8Y7_E2BEG[3] ,
    \Tile_X8Y7_E2BEG[2] ,
    \Tile_X8Y7_E2BEG[1] ,
    \Tile_X8Y7_E2BEG[0] }),
    .E2BEGb({\Tile_X8Y7_E2BEGb[7] ,
    \Tile_X8Y7_E2BEGb[6] ,
    \Tile_X8Y7_E2BEGb[5] ,
    \Tile_X8Y7_E2BEGb[4] ,
    \Tile_X8Y7_E2BEGb[3] ,
    \Tile_X8Y7_E2BEGb[2] ,
    \Tile_X8Y7_E2BEGb[1] ,
    \Tile_X8Y7_E2BEGb[0] }),
    .E2END({\Tile_X7Y7_E2BEGb[7] ,
    \Tile_X7Y7_E2BEGb[6] ,
    \Tile_X7Y7_E2BEGb[5] ,
    \Tile_X7Y7_E2BEGb[4] ,
    \Tile_X7Y7_E2BEGb[3] ,
    \Tile_X7Y7_E2BEGb[2] ,
    \Tile_X7Y7_E2BEGb[1] ,
    \Tile_X7Y7_E2BEGb[0] }),
    .E2MID({\Tile_X7Y7_E2BEG[7] ,
    \Tile_X7Y7_E2BEG[6] ,
    \Tile_X7Y7_E2BEG[5] ,
    \Tile_X7Y7_E2BEG[4] ,
    \Tile_X7Y7_E2BEG[3] ,
    \Tile_X7Y7_E2BEG[2] ,
    \Tile_X7Y7_E2BEG[1] ,
    \Tile_X7Y7_E2BEG[0] }),
    .E6BEG({\Tile_X8Y7_E6BEG[11] ,
    \Tile_X8Y7_E6BEG[10] ,
    \Tile_X8Y7_E6BEG[9] ,
    \Tile_X8Y7_E6BEG[8] ,
    \Tile_X8Y7_E6BEG[7] ,
    \Tile_X8Y7_E6BEG[6] ,
    \Tile_X8Y7_E6BEG[5] ,
    \Tile_X8Y7_E6BEG[4] ,
    \Tile_X8Y7_E6BEG[3] ,
    \Tile_X8Y7_E6BEG[2] ,
    \Tile_X8Y7_E6BEG[1] ,
    \Tile_X8Y7_E6BEG[0] }),
    .E6END({\Tile_X7Y7_E6BEG[11] ,
    \Tile_X7Y7_E6BEG[10] ,
    \Tile_X7Y7_E6BEG[9] ,
    \Tile_X7Y7_E6BEG[8] ,
    \Tile_X7Y7_E6BEG[7] ,
    \Tile_X7Y7_E6BEG[6] ,
    \Tile_X7Y7_E6BEG[5] ,
    \Tile_X7Y7_E6BEG[4] ,
    \Tile_X7Y7_E6BEG[3] ,
    \Tile_X7Y7_E6BEG[2] ,
    \Tile_X7Y7_E6BEG[1] ,
    \Tile_X7Y7_E6BEG[0] }),
    .EE4BEG({\Tile_X8Y7_EE4BEG[15] ,
    \Tile_X8Y7_EE4BEG[14] ,
    \Tile_X8Y7_EE4BEG[13] ,
    \Tile_X8Y7_EE4BEG[12] ,
    \Tile_X8Y7_EE4BEG[11] ,
    \Tile_X8Y7_EE4BEG[10] ,
    \Tile_X8Y7_EE4BEG[9] ,
    \Tile_X8Y7_EE4BEG[8] ,
    \Tile_X8Y7_EE4BEG[7] ,
    \Tile_X8Y7_EE4BEG[6] ,
    \Tile_X8Y7_EE4BEG[5] ,
    \Tile_X8Y7_EE4BEG[4] ,
    \Tile_X8Y7_EE4BEG[3] ,
    \Tile_X8Y7_EE4BEG[2] ,
    \Tile_X8Y7_EE4BEG[1] ,
    \Tile_X8Y7_EE4BEG[0] }),
    .EE4END({\Tile_X7Y7_EE4BEG[15] ,
    \Tile_X7Y7_EE4BEG[14] ,
    \Tile_X7Y7_EE4BEG[13] ,
    \Tile_X7Y7_EE4BEG[12] ,
    \Tile_X7Y7_EE4BEG[11] ,
    \Tile_X7Y7_EE4BEG[10] ,
    \Tile_X7Y7_EE4BEG[9] ,
    \Tile_X7Y7_EE4BEG[8] ,
    \Tile_X7Y7_EE4BEG[7] ,
    \Tile_X7Y7_EE4BEG[6] ,
    \Tile_X7Y7_EE4BEG[5] ,
    \Tile_X7Y7_EE4BEG[4] ,
    \Tile_X7Y7_EE4BEG[3] ,
    \Tile_X7Y7_EE4BEG[2] ,
    \Tile_X7Y7_EE4BEG[1] ,
    \Tile_X7Y7_EE4BEG[0] }),
    .FrameData({\Tile_X7Y7_FrameData_O[31] ,
    \Tile_X7Y7_FrameData_O[30] ,
    \Tile_X7Y7_FrameData_O[29] ,
    \Tile_X7Y7_FrameData_O[28] ,
    \Tile_X7Y7_FrameData_O[27] ,
    \Tile_X7Y7_FrameData_O[26] ,
    \Tile_X7Y7_FrameData_O[25] ,
    \Tile_X7Y7_FrameData_O[24] ,
    \Tile_X7Y7_FrameData_O[23] ,
    \Tile_X7Y7_FrameData_O[22] ,
    \Tile_X7Y7_FrameData_O[21] ,
    \Tile_X7Y7_FrameData_O[20] ,
    \Tile_X7Y7_FrameData_O[19] ,
    \Tile_X7Y7_FrameData_O[18] ,
    \Tile_X7Y7_FrameData_O[17] ,
    \Tile_X7Y7_FrameData_O[16] ,
    \Tile_X7Y7_FrameData_O[15] ,
    \Tile_X7Y7_FrameData_O[14] ,
    \Tile_X7Y7_FrameData_O[13] ,
    \Tile_X7Y7_FrameData_O[12] ,
    \Tile_X7Y7_FrameData_O[11] ,
    \Tile_X7Y7_FrameData_O[10] ,
    \Tile_X7Y7_FrameData_O[9] ,
    \Tile_X7Y7_FrameData_O[8] ,
    \Tile_X7Y7_FrameData_O[7] ,
    \Tile_X7Y7_FrameData_O[6] ,
    \Tile_X7Y7_FrameData_O[5] ,
    \Tile_X7Y7_FrameData_O[4] ,
    \Tile_X7Y7_FrameData_O[3] ,
    \Tile_X7Y7_FrameData_O[2] ,
    \Tile_X7Y7_FrameData_O[1] ,
    \Tile_X7Y7_FrameData_O[0] }),
    .FrameData_O({\Tile_X8Y7_FrameData_O[31] ,
    \Tile_X8Y7_FrameData_O[30] ,
    \Tile_X8Y7_FrameData_O[29] ,
    \Tile_X8Y7_FrameData_O[28] ,
    \Tile_X8Y7_FrameData_O[27] ,
    \Tile_X8Y7_FrameData_O[26] ,
    \Tile_X8Y7_FrameData_O[25] ,
    \Tile_X8Y7_FrameData_O[24] ,
    \Tile_X8Y7_FrameData_O[23] ,
    \Tile_X8Y7_FrameData_O[22] ,
    \Tile_X8Y7_FrameData_O[21] ,
    \Tile_X8Y7_FrameData_O[20] ,
    \Tile_X8Y7_FrameData_O[19] ,
    \Tile_X8Y7_FrameData_O[18] ,
    \Tile_X8Y7_FrameData_O[17] ,
    \Tile_X8Y7_FrameData_O[16] ,
    \Tile_X8Y7_FrameData_O[15] ,
    \Tile_X8Y7_FrameData_O[14] ,
    \Tile_X8Y7_FrameData_O[13] ,
    \Tile_X8Y7_FrameData_O[12] ,
    \Tile_X8Y7_FrameData_O[11] ,
    \Tile_X8Y7_FrameData_O[10] ,
    \Tile_X8Y7_FrameData_O[9] ,
    \Tile_X8Y7_FrameData_O[8] ,
    \Tile_X8Y7_FrameData_O[7] ,
    \Tile_X8Y7_FrameData_O[6] ,
    \Tile_X8Y7_FrameData_O[5] ,
    \Tile_X8Y7_FrameData_O[4] ,
    \Tile_X8Y7_FrameData_O[3] ,
    \Tile_X8Y7_FrameData_O[2] ,
    \Tile_X8Y7_FrameData_O[1] ,
    \Tile_X8Y7_FrameData_O[0] }),
    .FrameStrobe({\Tile_X8Y8_FrameStrobe_O[19] ,
    \Tile_X8Y8_FrameStrobe_O[18] ,
    \Tile_X8Y8_FrameStrobe_O[17] ,
    \Tile_X8Y8_FrameStrobe_O[16] ,
    \Tile_X8Y8_FrameStrobe_O[15] ,
    \Tile_X8Y8_FrameStrobe_O[14] ,
    \Tile_X8Y8_FrameStrobe_O[13] ,
    \Tile_X8Y8_FrameStrobe_O[12] ,
    \Tile_X8Y8_FrameStrobe_O[11] ,
    \Tile_X8Y8_FrameStrobe_O[10] ,
    \Tile_X8Y8_FrameStrobe_O[9] ,
    \Tile_X8Y8_FrameStrobe_O[8] ,
    \Tile_X8Y8_FrameStrobe_O[7] ,
    \Tile_X8Y8_FrameStrobe_O[6] ,
    \Tile_X8Y8_FrameStrobe_O[5] ,
    \Tile_X8Y8_FrameStrobe_O[4] ,
    \Tile_X8Y8_FrameStrobe_O[3] ,
    \Tile_X8Y8_FrameStrobe_O[2] ,
    \Tile_X8Y8_FrameStrobe_O[1] ,
    \Tile_X8Y8_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X8Y7_FrameStrobe_O[19] ,
    \Tile_X8Y7_FrameStrobe_O[18] ,
    \Tile_X8Y7_FrameStrobe_O[17] ,
    \Tile_X8Y7_FrameStrobe_O[16] ,
    \Tile_X8Y7_FrameStrobe_O[15] ,
    \Tile_X8Y7_FrameStrobe_O[14] ,
    \Tile_X8Y7_FrameStrobe_O[13] ,
    \Tile_X8Y7_FrameStrobe_O[12] ,
    \Tile_X8Y7_FrameStrobe_O[11] ,
    \Tile_X8Y7_FrameStrobe_O[10] ,
    \Tile_X8Y7_FrameStrobe_O[9] ,
    \Tile_X8Y7_FrameStrobe_O[8] ,
    \Tile_X8Y7_FrameStrobe_O[7] ,
    \Tile_X8Y7_FrameStrobe_O[6] ,
    \Tile_X8Y7_FrameStrobe_O[5] ,
    \Tile_X8Y7_FrameStrobe_O[4] ,
    \Tile_X8Y7_FrameStrobe_O[3] ,
    \Tile_X8Y7_FrameStrobe_O[2] ,
    \Tile_X8Y7_FrameStrobe_O[1] ,
    \Tile_X8Y7_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X8Y7_N1BEG[3] ,
    \Tile_X8Y7_N1BEG[2] ,
    \Tile_X8Y7_N1BEG[1] ,
    \Tile_X8Y7_N1BEG[0] }),
    .N1END({\Tile_X8Y8_N1BEG[3] ,
    \Tile_X8Y8_N1BEG[2] ,
    \Tile_X8Y8_N1BEG[1] ,
    \Tile_X8Y8_N1BEG[0] }),
    .N2BEG({\Tile_X8Y7_N2BEG[7] ,
    \Tile_X8Y7_N2BEG[6] ,
    \Tile_X8Y7_N2BEG[5] ,
    \Tile_X8Y7_N2BEG[4] ,
    \Tile_X8Y7_N2BEG[3] ,
    \Tile_X8Y7_N2BEG[2] ,
    \Tile_X8Y7_N2BEG[1] ,
    \Tile_X8Y7_N2BEG[0] }),
    .N2BEGb({\Tile_X8Y7_N2BEGb[7] ,
    \Tile_X8Y7_N2BEGb[6] ,
    \Tile_X8Y7_N2BEGb[5] ,
    \Tile_X8Y7_N2BEGb[4] ,
    \Tile_X8Y7_N2BEGb[3] ,
    \Tile_X8Y7_N2BEGb[2] ,
    \Tile_X8Y7_N2BEGb[1] ,
    \Tile_X8Y7_N2BEGb[0] }),
    .N2END({\Tile_X8Y8_N2BEGb[7] ,
    \Tile_X8Y8_N2BEGb[6] ,
    \Tile_X8Y8_N2BEGb[5] ,
    \Tile_X8Y8_N2BEGb[4] ,
    \Tile_X8Y8_N2BEGb[3] ,
    \Tile_X8Y8_N2BEGb[2] ,
    \Tile_X8Y8_N2BEGb[1] ,
    \Tile_X8Y8_N2BEGb[0] }),
    .N2MID({\Tile_X8Y8_N2BEG[7] ,
    \Tile_X8Y8_N2BEG[6] ,
    \Tile_X8Y8_N2BEG[5] ,
    \Tile_X8Y8_N2BEG[4] ,
    \Tile_X8Y8_N2BEG[3] ,
    \Tile_X8Y8_N2BEG[2] ,
    \Tile_X8Y8_N2BEG[1] ,
    \Tile_X8Y8_N2BEG[0] }),
    .N4BEG({\Tile_X8Y7_N4BEG[15] ,
    \Tile_X8Y7_N4BEG[14] ,
    \Tile_X8Y7_N4BEG[13] ,
    \Tile_X8Y7_N4BEG[12] ,
    \Tile_X8Y7_N4BEG[11] ,
    \Tile_X8Y7_N4BEG[10] ,
    \Tile_X8Y7_N4BEG[9] ,
    \Tile_X8Y7_N4BEG[8] ,
    \Tile_X8Y7_N4BEG[7] ,
    \Tile_X8Y7_N4BEG[6] ,
    \Tile_X8Y7_N4BEG[5] ,
    \Tile_X8Y7_N4BEG[4] ,
    \Tile_X8Y7_N4BEG[3] ,
    \Tile_X8Y7_N4BEG[2] ,
    \Tile_X8Y7_N4BEG[1] ,
    \Tile_X8Y7_N4BEG[0] }),
    .N4END({\Tile_X8Y8_N4BEG[15] ,
    \Tile_X8Y8_N4BEG[14] ,
    \Tile_X8Y8_N4BEG[13] ,
    \Tile_X8Y8_N4BEG[12] ,
    \Tile_X8Y8_N4BEG[11] ,
    \Tile_X8Y8_N4BEG[10] ,
    \Tile_X8Y8_N4BEG[9] ,
    \Tile_X8Y8_N4BEG[8] ,
    \Tile_X8Y8_N4BEG[7] ,
    \Tile_X8Y8_N4BEG[6] ,
    \Tile_X8Y8_N4BEG[5] ,
    \Tile_X8Y8_N4BEG[4] ,
    \Tile_X8Y8_N4BEG[3] ,
    \Tile_X8Y8_N4BEG[2] ,
    \Tile_X8Y8_N4BEG[1] ,
    \Tile_X8Y8_N4BEG[0] }),
    .NN4BEG({\Tile_X8Y7_NN4BEG[15] ,
    \Tile_X8Y7_NN4BEG[14] ,
    \Tile_X8Y7_NN4BEG[13] ,
    \Tile_X8Y7_NN4BEG[12] ,
    \Tile_X8Y7_NN4BEG[11] ,
    \Tile_X8Y7_NN4BEG[10] ,
    \Tile_X8Y7_NN4BEG[9] ,
    \Tile_X8Y7_NN4BEG[8] ,
    \Tile_X8Y7_NN4BEG[7] ,
    \Tile_X8Y7_NN4BEG[6] ,
    \Tile_X8Y7_NN4BEG[5] ,
    \Tile_X8Y7_NN4BEG[4] ,
    \Tile_X8Y7_NN4BEG[3] ,
    \Tile_X8Y7_NN4BEG[2] ,
    \Tile_X8Y7_NN4BEG[1] ,
    \Tile_X8Y7_NN4BEG[0] }),
    .NN4END({\Tile_X8Y8_NN4BEG[15] ,
    \Tile_X8Y8_NN4BEG[14] ,
    \Tile_X8Y8_NN4BEG[13] ,
    \Tile_X8Y8_NN4BEG[12] ,
    \Tile_X8Y8_NN4BEG[11] ,
    \Tile_X8Y8_NN4BEG[10] ,
    \Tile_X8Y8_NN4BEG[9] ,
    \Tile_X8Y8_NN4BEG[8] ,
    \Tile_X8Y8_NN4BEG[7] ,
    \Tile_X8Y8_NN4BEG[6] ,
    \Tile_X8Y8_NN4BEG[5] ,
    \Tile_X8Y8_NN4BEG[4] ,
    \Tile_X8Y8_NN4BEG[3] ,
    \Tile_X8Y8_NN4BEG[2] ,
    \Tile_X8Y8_NN4BEG[1] ,
    \Tile_X8Y8_NN4BEG[0] }),
    .S1BEG({\Tile_X8Y7_S1BEG[3] ,
    \Tile_X8Y7_S1BEG[2] ,
    \Tile_X8Y7_S1BEG[1] ,
    \Tile_X8Y7_S1BEG[0] }),
    .S1END({\Tile_X8Y6_S1BEG[3] ,
    \Tile_X8Y6_S1BEG[2] ,
    \Tile_X8Y6_S1BEG[1] ,
    \Tile_X8Y6_S1BEG[0] }),
    .S2BEG({\Tile_X8Y7_S2BEG[7] ,
    \Tile_X8Y7_S2BEG[6] ,
    \Tile_X8Y7_S2BEG[5] ,
    \Tile_X8Y7_S2BEG[4] ,
    \Tile_X8Y7_S2BEG[3] ,
    \Tile_X8Y7_S2BEG[2] ,
    \Tile_X8Y7_S2BEG[1] ,
    \Tile_X8Y7_S2BEG[0] }),
    .S2BEGb({\Tile_X8Y7_S2BEGb[7] ,
    \Tile_X8Y7_S2BEGb[6] ,
    \Tile_X8Y7_S2BEGb[5] ,
    \Tile_X8Y7_S2BEGb[4] ,
    \Tile_X8Y7_S2BEGb[3] ,
    \Tile_X8Y7_S2BEGb[2] ,
    \Tile_X8Y7_S2BEGb[1] ,
    \Tile_X8Y7_S2BEGb[0] }),
    .S2END({\Tile_X8Y6_S2BEGb[7] ,
    \Tile_X8Y6_S2BEGb[6] ,
    \Tile_X8Y6_S2BEGb[5] ,
    \Tile_X8Y6_S2BEGb[4] ,
    \Tile_X8Y6_S2BEGb[3] ,
    \Tile_X8Y6_S2BEGb[2] ,
    \Tile_X8Y6_S2BEGb[1] ,
    \Tile_X8Y6_S2BEGb[0] }),
    .S2MID({\Tile_X8Y6_S2BEG[7] ,
    \Tile_X8Y6_S2BEG[6] ,
    \Tile_X8Y6_S2BEG[5] ,
    \Tile_X8Y6_S2BEG[4] ,
    \Tile_X8Y6_S2BEG[3] ,
    \Tile_X8Y6_S2BEG[2] ,
    \Tile_X8Y6_S2BEG[1] ,
    \Tile_X8Y6_S2BEG[0] }),
    .S4BEG({\Tile_X8Y7_S4BEG[15] ,
    \Tile_X8Y7_S4BEG[14] ,
    \Tile_X8Y7_S4BEG[13] ,
    \Tile_X8Y7_S4BEG[12] ,
    \Tile_X8Y7_S4BEG[11] ,
    \Tile_X8Y7_S4BEG[10] ,
    \Tile_X8Y7_S4BEG[9] ,
    \Tile_X8Y7_S4BEG[8] ,
    \Tile_X8Y7_S4BEG[7] ,
    \Tile_X8Y7_S4BEG[6] ,
    \Tile_X8Y7_S4BEG[5] ,
    \Tile_X8Y7_S4BEG[4] ,
    \Tile_X8Y7_S4BEG[3] ,
    \Tile_X8Y7_S4BEG[2] ,
    \Tile_X8Y7_S4BEG[1] ,
    \Tile_X8Y7_S4BEG[0] }),
    .S4END({\Tile_X8Y6_S4BEG[15] ,
    \Tile_X8Y6_S4BEG[14] ,
    \Tile_X8Y6_S4BEG[13] ,
    \Tile_X8Y6_S4BEG[12] ,
    \Tile_X8Y6_S4BEG[11] ,
    \Tile_X8Y6_S4BEG[10] ,
    \Tile_X8Y6_S4BEG[9] ,
    \Tile_X8Y6_S4BEG[8] ,
    \Tile_X8Y6_S4BEG[7] ,
    \Tile_X8Y6_S4BEG[6] ,
    \Tile_X8Y6_S4BEG[5] ,
    \Tile_X8Y6_S4BEG[4] ,
    \Tile_X8Y6_S4BEG[3] ,
    \Tile_X8Y6_S4BEG[2] ,
    \Tile_X8Y6_S4BEG[1] ,
    \Tile_X8Y6_S4BEG[0] }),
    .SS4BEG({\Tile_X8Y7_SS4BEG[15] ,
    \Tile_X8Y7_SS4BEG[14] ,
    \Tile_X8Y7_SS4BEG[13] ,
    \Tile_X8Y7_SS4BEG[12] ,
    \Tile_X8Y7_SS4BEG[11] ,
    \Tile_X8Y7_SS4BEG[10] ,
    \Tile_X8Y7_SS4BEG[9] ,
    \Tile_X8Y7_SS4BEG[8] ,
    \Tile_X8Y7_SS4BEG[7] ,
    \Tile_X8Y7_SS4BEG[6] ,
    \Tile_X8Y7_SS4BEG[5] ,
    \Tile_X8Y7_SS4BEG[4] ,
    \Tile_X8Y7_SS4BEG[3] ,
    \Tile_X8Y7_SS4BEG[2] ,
    \Tile_X8Y7_SS4BEG[1] ,
    \Tile_X8Y7_SS4BEG[0] }),
    .SS4END({\Tile_X8Y6_SS4BEG[15] ,
    \Tile_X8Y6_SS4BEG[14] ,
    \Tile_X8Y6_SS4BEG[13] ,
    \Tile_X8Y6_SS4BEG[12] ,
    \Tile_X8Y6_SS4BEG[11] ,
    \Tile_X8Y6_SS4BEG[10] ,
    \Tile_X8Y6_SS4BEG[9] ,
    \Tile_X8Y6_SS4BEG[8] ,
    \Tile_X8Y6_SS4BEG[7] ,
    \Tile_X8Y6_SS4BEG[6] ,
    \Tile_X8Y6_SS4BEG[5] ,
    \Tile_X8Y6_SS4BEG[4] ,
    \Tile_X8Y6_SS4BEG[3] ,
    \Tile_X8Y6_SS4BEG[2] ,
    \Tile_X8Y6_SS4BEG[1] ,
    \Tile_X8Y6_SS4BEG[0] }),
    .W1BEG({\Tile_X8Y7_W1BEG[3] ,
    \Tile_X8Y7_W1BEG[2] ,
    \Tile_X8Y7_W1BEG[1] ,
    \Tile_X8Y7_W1BEG[0] }),
    .W1END({\Tile_X9Y7_W1BEG[3] ,
    \Tile_X9Y7_W1BEG[2] ,
    \Tile_X9Y7_W1BEG[1] ,
    \Tile_X9Y7_W1BEG[0] }),
    .W2BEG({\Tile_X8Y7_W2BEG[7] ,
    \Tile_X8Y7_W2BEG[6] ,
    \Tile_X8Y7_W2BEG[5] ,
    \Tile_X8Y7_W2BEG[4] ,
    \Tile_X8Y7_W2BEG[3] ,
    \Tile_X8Y7_W2BEG[2] ,
    \Tile_X8Y7_W2BEG[1] ,
    \Tile_X8Y7_W2BEG[0] }),
    .W2BEGb({\Tile_X8Y7_W2BEGb[7] ,
    \Tile_X8Y7_W2BEGb[6] ,
    \Tile_X8Y7_W2BEGb[5] ,
    \Tile_X8Y7_W2BEGb[4] ,
    \Tile_X8Y7_W2BEGb[3] ,
    \Tile_X8Y7_W2BEGb[2] ,
    \Tile_X8Y7_W2BEGb[1] ,
    \Tile_X8Y7_W2BEGb[0] }),
    .W2END({\Tile_X9Y7_W2BEGb[7] ,
    \Tile_X9Y7_W2BEGb[6] ,
    \Tile_X9Y7_W2BEGb[5] ,
    \Tile_X9Y7_W2BEGb[4] ,
    \Tile_X9Y7_W2BEGb[3] ,
    \Tile_X9Y7_W2BEGb[2] ,
    \Tile_X9Y7_W2BEGb[1] ,
    \Tile_X9Y7_W2BEGb[0] }),
    .W2MID({\Tile_X9Y7_W2BEG[7] ,
    \Tile_X9Y7_W2BEG[6] ,
    \Tile_X9Y7_W2BEG[5] ,
    \Tile_X9Y7_W2BEG[4] ,
    \Tile_X9Y7_W2BEG[3] ,
    \Tile_X9Y7_W2BEG[2] ,
    \Tile_X9Y7_W2BEG[1] ,
    \Tile_X9Y7_W2BEG[0] }),
    .W6BEG({\Tile_X8Y7_W6BEG[11] ,
    \Tile_X8Y7_W6BEG[10] ,
    \Tile_X8Y7_W6BEG[9] ,
    \Tile_X8Y7_W6BEG[8] ,
    \Tile_X8Y7_W6BEG[7] ,
    \Tile_X8Y7_W6BEG[6] ,
    \Tile_X8Y7_W6BEG[5] ,
    \Tile_X8Y7_W6BEG[4] ,
    \Tile_X8Y7_W6BEG[3] ,
    \Tile_X8Y7_W6BEG[2] ,
    \Tile_X8Y7_W6BEG[1] ,
    \Tile_X8Y7_W6BEG[0] }),
    .W6END({\Tile_X9Y7_W6BEG[11] ,
    \Tile_X9Y7_W6BEG[10] ,
    \Tile_X9Y7_W6BEG[9] ,
    \Tile_X9Y7_W6BEG[8] ,
    \Tile_X9Y7_W6BEG[7] ,
    \Tile_X9Y7_W6BEG[6] ,
    \Tile_X9Y7_W6BEG[5] ,
    \Tile_X9Y7_W6BEG[4] ,
    \Tile_X9Y7_W6BEG[3] ,
    \Tile_X9Y7_W6BEG[2] ,
    \Tile_X9Y7_W6BEG[1] ,
    \Tile_X9Y7_W6BEG[0] }),
    .WW4BEG({\Tile_X8Y7_WW4BEG[15] ,
    \Tile_X8Y7_WW4BEG[14] ,
    \Tile_X8Y7_WW4BEG[13] ,
    \Tile_X8Y7_WW4BEG[12] ,
    \Tile_X8Y7_WW4BEG[11] ,
    \Tile_X8Y7_WW4BEG[10] ,
    \Tile_X8Y7_WW4BEG[9] ,
    \Tile_X8Y7_WW4BEG[8] ,
    \Tile_X8Y7_WW4BEG[7] ,
    \Tile_X8Y7_WW4BEG[6] ,
    \Tile_X8Y7_WW4BEG[5] ,
    \Tile_X8Y7_WW4BEG[4] ,
    \Tile_X8Y7_WW4BEG[3] ,
    \Tile_X8Y7_WW4BEG[2] ,
    \Tile_X8Y7_WW4BEG[1] ,
    \Tile_X8Y7_WW4BEG[0] }),
    .WW4END({\Tile_X9Y7_WW4BEG[15] ,
    \Tile_X9Y7_WW4BEG[14] ,
    \Tile_X9Y7_WW4BEG[13] ,
    \Tile_X9Y7_WW4BEG[12] ,
    \Tile_X9Y7_WW4BEG[11] ,
    \Tile_X9Y7_WW4BEG[10] ,
    \Tile_X9Y7_WW4BEG[9] ,
    \Tile_X9Y7_WW4BEG[8] ,
    \Tile_X9Y7_WW4BEG[7] ,
    \Tile_X9Y7_WW4BEG[6] ,
    \Tile_X9Y7_WW4BEG[5] ,
    \Tile_X9Y7_WW4BEG[4] ,
    \Tile_X9Y7_WW4BEG[3] ,
    \Tile_X9Y7_WW4BEG[2] ,
    \Tile_X9Y7_WW4BEG[1] ,
    \Tile_X9Y7_WW4BEG[0] }));
 LUT4AB Tile_X8Y8_LUT4AB (.Ci(Tile_X8Y9_Co),
    .Co(Tile_X8Y8_Co),
    .UserCLK(Tile_X8Y9_UserCLKo),
    .UserCLKo(Tile_X8Y8_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X8Y8_E1BEG[3] ,
    \Tile_X8Y8_E1BEG[2] ,
    \Tile_X8Y8_E1BEG[1] ,
    \Tile_X8Y8_E1BEG[0] }),
    .E1END({\Tile_X7Y8_E1BEG[3] ,
    \Tile_X7Y8_E1BEG[2] ,
    \Tile_X7Y8_E1BEG[1] ,
    \Tile_X7Y8_E1BEG[0] }),
    .E2BEG({\Tile_X8Y8_E2BEG[7] ,
    \Tile_X8Y8_E2BEG[6] ,
    \Tile_X8Y8_E2BEG[5] ,
    \Tile_X8Y8_E2BEG[4] ,
    \Tile_X8Y8_E2BEG[3] ,
    \Tile_X8Y8_E2BEG[2] ,
    \Tile_X8Y8_E2BEG[1] ,
    \Tile_X8Y8_E2BEG[0] }),
    .E2BEGb({\Tile_X8Y8_E2BEGb[7] ,
    \Tile_X8Y8_E2BEGb[6] ,
    \Tile_X8Y8_E2BEGb[5] ,
    \Tile_X8Y8_E2BEGb[4] ,
    \Tile_X8Y8_E2BEGb[3] ,
    \Tile_X8Y8_E2BEGb[2] ,
    \Tile_X8Y8_E2BEGb[1] ,
    \Tile_X8Y8_E2BEGb[0] }),
    .E2END({\Tile_X7Y8_E2BEGb[7] ,
    \Tile_X7Y8_E2BEGb[6] ,
    \Tile_X7Y8_E2BEGb[5] ,
    \Tile_X7Y8_E2BEGb[4] ,
    \Tile_X7Y8_E2BEGb[3] ,
    \Tile_X7Y8_E2BEGb[2] ,
    \Tile_X7Y8_E2BEGb[1] ,
    \Tile_X7Y8_E2BEGb[0] }),
    .E2MID({\Tile_X7Y8_E2BEG[7] ,
    \Tile_X7Y8_E2BEG[6] ,
    \Tile_X7Y8_E2BEG[5] ,
    \Tile_X7Y8_E2BEG[4] ,
    \Tile_X7Y8_E2BEG[3] ,
    \Tile_X7Y8_E2BEG[2] ,
    \Tile_X7Y8_E2BEG[1] ,
    \Tile_X7Y8_E2BEG[0] }),
    .E6BEG({\Tile_X8Y8_E6BEG[11] ,
    \Tile_X8Y8_E6BEG[10] ,
    \Tile_X8Y8_E6BEG[9] ,
    \Tile_X8Y8_E6BEG[8] ,
    \Tile_X8Y8_E6BEG[7] ,
    \Tile_X8Y8_E6BEG[6] ,
    \Tile_X8Y8_E6BEG[5] ,
    \Tile_X8Y8_E6BEG[4] ,
    \Tile_X8Y8_E6BEG[3] ,
    \Tile_X8Y8_E6BEG[2] ,
    \Tile_X8Y8_E6BEG[1] ,
    \Tile_X8Y8_E6BEG[0] }),
    .E6END({\Tile_X7Y8_E6BEG[11] ,
    \Tile_X7Y8_E6BEG[10] ,
    \Tile_X7Y8_E6BEG[9] ,
    \Tile_X7Y8_E6BEG[8] ,
    \Tile_X7Y8_E6BEG[7] ,
    \Tile_X7Y8_E6BEG[6] ,
    \Tile_X7Y8_E6BEG[5] ,
    \Tile_X7Y8_E6BEG[4] ,
    \Tile_X7Y8_E6BEG[3] ,
    \Tile_X7Y8_E6BEG[2] ,
    \Tile_X7Y8_E6BEG[1] ,
    \Tile_X7Y8_E6BEG[0] }),
    .EE4BEG({\Tile_X8Y8_EE4BEG[15] ,
    \Tile_X8Y8_EE4BEG[14] ,
    \Tile_X8Y8_EE4BEG[13] ,
    \Tile_X8Y8_EE4BEG[12] ,
    \Tile_X8Y8_EE4BEG[11] ,
    \Tile_X8Y8_EE4BEG[10] ,
    \Tile_X8Y8_EE4BEG[9] ,
    \Tile_X8Y8_EE4BEG[8] ,
    \Tile_X8Y8_EE4BEG[7] ,
    \Tile_X8Y8_EE4BEG[6] ,
    \Tile_X8Y8_EE4BEG[5] ,
    \Tile_X8Y8_EE4BEG[4] ,
    \Tile_X8Y8_EE4BEG[3] ,
    \Tile_X8Y8_EE4BEG[2] ,
    \Tile_X8Y8_EE4BEG[1] ,
    \Tile_X8Y8_EE4BEG[0] }),
    .EE4END({\Tile_X7Y8_EE4BEG[15] ,
    \Tile_X7Y8_EE4BEG[14] ,
    \Tile_X7Y8_EE4BEG[13] ,
    \Tile_X7Y8_EE4BEG[12] ,
    \Tile_X7Y8_EE4BEG[11] ,
    \Tile_X7Y8_EE4BEG[10] ,
    \Tile_X7Y8_EE4BEG[9] ,
    \Tile_X7Y8_EE4BEG[8] ,
    \Tile_X7Y8_EE4BEG[7] ,
    \Tile_X7Y8_EE4BEG[6] ,
    \Tile_X7Y8_EE4BEG[5] ,
    \Tile_X7Y8_EE4BEG[4] ,
    \Tile_X7Y8_EE4BEG[3] ,
    \Tile_X7Y8_EE4BEG[2] ,
    \Tile_X7Y8_EE4BEG[1] ,
    \Tile_X7Y8_EE4BEG[0] }),
    .FrameData({\Tile_X7Y8_FrameData_O[31] ,
    \Tile_X7Y8_FrameData_O[30] ,
    \Tile_X7Y8_FrameData_O[29] ,
    \Tile_X7Y8_FrameData_O[28] ,
    \Tile_X7Y8_FrameData_O[27] ,
    \Tile_X7Y8_FrameData_O[26] ,
    \Tile_X7Y8_FrameData_O[25] ,
    \Tile_X7Y8_FrameData_O[24] ,
    \Tile_X7Y8_FrameData_O[23] ,
    \Tile_X7Y8_FrameData_O[22] ,
    \Tile_X7Y8_FrameData_O[21] ,
    \Tile_X7Y8_FrameData_O[20] ,
    \Tile_X7Y8_FrameData_O[19] ,
    \Tile_X7Y8_FrameData_O[18] ,
    \Tile_X7Y8_FrameData_O[17] ,
    \Tile_X7Y8_FrameData_O[16] ,
    \Tile_X7Y8_FrameData_O[15] ,
    \Tile_X7Y8_FrameData_O[14] ,
    \Tile_X7Y8_FrameData_O[13] ,
    \Tile_X7Y8_FrameData_O[12] ,
    \Tile_X7Y8_FrameData_O[11] ,
    \Tile_X7Y8_FrameData_O[10] ,
    \Tile_X7Y8_FrameData_O[9] ,
    \Tile_X7Y8_FrameData_O[8] ,
    \Tile_X7Y8_FrameData_O[7] ,
    \Tile_X7Y8_FrameData_O[6] ,
    \Tile_X7Y8_FrameData_O[5] ,
    \Tile_X7Y8_FrameData_O[4] ,
    \Tile_X7Y8_FrameData_O[3] ,
    \Tile_X7Y8_FrameData_O[2] ,
    \Tile_X7Y8_FrameData_O[1] ,
    \Tile_X7Y8_FrameData_O[0] }),
    .FrameData_O({\Tile_X8Y8_FrameData_O[31] ,
    \Tile_X8Y8_FrameData_O[30] ,
    \Tile_X8Y8_FrameData_O[29] ,
    \Tile_X8Y8_FrameData_O[28] ,
    \Tile_X8Y8_FrameData_O[27] ,
    \Tile_X8Y8_FrameData_O[26] ,
    \Tile_X8Y8_FrameData_O[25] ,
    \Tile_X8Y8_FrameData_O[24] ,
    \Tile_X8Y8_FrameData_O[23] ,
    \Tile_X8Y8_FrameData_O[22] ,
    \Tile_X8Y8_FrameData_O[21] ,
    \Tile_X8Y8_FrameData_O[20] ,
    \Tile_X8Y8_FrameData_O[19] ,
    \Tile_X8Y8_FrameData_O[18] ,
    \Tile_X8Y8_FrameData_O[17] ,
    \Tile_X8Y8_FrameData_O[16] ,
    \Tile_X8Y8_FrameData_O[15] ,
    \Tile_X8Y8_FrameData_O[14] ,
    \Tile_X8Y8_FrameData_O[13] ,
    \Tile_X8Y8_FrameData_O[12] ,
    \Tile_X8Y8_FrameData_O[11] ,
    \Tile_X8Y8_FrameData_O[10] ,
    \Tile_X8Y8_FrameData_O[9] ,
    \Tile_X8Y8_FrameData_O[8] ,
    \Tile_X8Y8_FrameData_O[7] ,
    \Tile_X8Y8_FrameData_O[6] ,
    \Tile_X8Y8_FrameData_O[5] ,
    \Tile_X8Y8_FrameData_O[4] ,
    \Tile_X8Y8_FrameData_O[3] ,
    \Tile_X8Y8_FrameData_O[2] ,
    \Tile_X8Y8_FrameData_O[1] ,
    \Tile_X8Y8_FrameData_O[0] }),
    .FrameStrobe({\Tile_X8Y9_FrameStrobe_O[19] ,
    \Tile_X8Y9_FrameStrobe_O[18] ,
    \Tile_X8Y9_FrameStrobe_O[17] ,
    \Tile_X8Y9_FrameStrobe_O[16] ,
    \Tile_X8Y9_FrameStrobe_O[15] ,
    \Tile_X8Y9_FrameStrobe_O[14] ,
    \Tile_X8Y9_FrameStrobe_O[13] ,
    \Tile_X8Y9_FrameStrobe_O[12] ,
    \Tile_X8Y9_FrameStrobe_O[11] ,
    \Tile_X8Y9_FrameStrobe_O[10] ,
    \Tile_X8Y9_FrameStrobe_O[9] ,
    \Tile_X8Y9_FrameStrobe_O[8] ,
    \Tile_X8Y9_FrameStrobe_O[7] ,
    \Tile_X8Y9_FrameStrobe_O[6] ,
    \Tile_X8Y9_FrameStrobe_O[5] ,
    \Tile_X8Y9_FrameStrobe_O[4] ,
    \Tile_X8Y9_FrameStrobe_O[3] ,
    \Tile_X8Y9_FrameStrobe_O[2] ,
    \Tile_X8Y9_FrameStrobe_O[1] ,
    \Tile_X8Y9_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X8Y8_FrameStrobe_O[19] ,
    \Tile_X8Y8_FrameStrobe_O[18] ,
    \Tile_X8Y8_FrameStrobe_O[17] ,
    \Tile_X8Y8_FrameStrobe_O[16] ,
    \Tile_X8Y8_FrameStrobe_O[15] ,
    \Tile_X8Y8_FrameStrobe_O[14] ,
    \Tile_X8Y8_FrameStrobe_O[13] ,
    \Tile_X8Y8_FrameStrobe_O[12] ,
    \Tile_X8Y8_FrameStrobe_O[11] ,
    \Tile_X8Y8_FrameStrobe_O[10] ,
    \Tile_X8Y8_FrameStrobe_O[9] ,
    \Tile_X8Y8_FrameStrobe_O[8] ,
    \Tile_X8Y8_FrameStrobe_O[7] ,
    \Tile_X8Y8_FrameStrobe_O[6] ,
    \Tile_X8Y8_FrameStrobe_O[5] ,
    \Tile_X8Y8_FrameStrobe_O[4] ,
    \Tile_X8Y8_FrameStrobe_O[3] ,
    \Tile_X8Y8_FrameStrobe_O[2] ,
    \Tile_X8Y8_FrameStrobe_O[1] ,
    \Tile_X8Y8_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X8Y8_N1BEG[3] ,
    \Tile_X8Y8_N1BEG[2] ,
    \Tile_X8Y8_N1BEG[1] ,
    \Tile_X8Y8_N1BEG[0] }),
    .N1END({\Tile_X8Y9_N1BEG[3] ,
    \Tile_X8Y9_N1BEG[2] ,
    \Tile_X8Y9_N1BEG[1] ,
    \Tile_X8Y9_N1BEG[0] }),
    .N2BEG({\Tile_X8Y8_N2BEG[7] ,
    \Tile_X8Y8_N2BEG[6] ,
    \Tile_X8Y8_N2BEG[5] ,
    \Tile_X8Y8_N2BEG[4] ,
    \Tile_X8Y8_N2BEG[3] ,
    \Tile_X8Y8_N2BEG[2] ,
    \Tile_X8Y8_N2BEG[1] ,
    \Tile_X8Y8_N2BEG[0] }),
    .N2BEGb({\Tile_X8Y8_N2BEGb[7] ,
    \Tile_X8Y8_N2BEGb[6] ,
    \Tile_X8Y8_N2BEGb[5] ,
    \Tile_X8Y8_N2BEGb[4] ,
    \Tile_X8Y8_N2BEGb[3] ,
    \Tile_X8Y8_N2BEGb[2] ,
    \Tile_X8Y8_N2BEGb[1] ,
    \Tile_X8Y8_N2BEGb[0] }),
    .N2END({\Tile_X8Y9_N2BEGb[7] ,
    \Tile_X8Y9_N2BEGb[6] ,
    \Tile_X8Y9_N2BEGb[5] ,
    \Tile_X8Y9_N2BEGb[4] ,
    \Tile_X8Y9_N2BEGb[3] ,
    \Tile_X8Y9_N2BEGb[2] ,
    \Tile_X8Y9_N2BEGb[1] ,
    \Tile_X8Y9_N2BEGb[0] }),
    .N2MID({\Tile_X8Y9_N2BEG[7] ,
    \Tile_X8Y9_N2BEG[6] ,
    \Tile_X8Y9_N2BEG[5] ,
    \Tile_X8Y9_N2BEG[4] ,
    \Tile_X8Y9_N2BEG[3] ,
    \Tile_X8Y9_N2BEG[2] ,
    \Tile_X8Y9_N2BEG[1] ,
    \Tile_X8Y9_N2BEG[0] }),
    .N4BEG({\Tile_X8Y8_N4BEG[15] ,
    \Tile_X8Y8_N4BEG[14] ,
    \Tile_X8Y8_N4BEG[13] ,
    \Tile_X8Y8_N4BEG[12] ,
    \Tile_X8Y8_N4BEG[11] ,
    \Tile_X8Y8_N4BEG[10] ,
    \Tile_X8Y8_N4BEG[9] ,
    \Tile_X8Y8_N4BEG[8] ,
    \Tile_X8Y8_N4BEG[7] ,
    \Tile_X8Y8_N4BEG[6] ,
    \Tile_X8Y8_N4BEG[5] ,
    \Tile_X8Y8_N4BEG[4] ,
    \Tile_X8Y8_N4BEG[3] ,
    \Tile_X8Y8_N4BEG[2] ,
    \Tile_X8Y8_N4BEG[1] ,
    \Tile_X8Y8_N4BEG[0] }),
    .N4END({\Tile_X8Y9_N4BEG[15] ,
    \Tile_X8Y9_N4BEG[14] ,
    \Tile_X8Y9_N4BEG[13] ,
    \Tile_X8Y9_N4BEG[12] ,
    \Tile_X8Y9_N4BEG[11] ,
    \Tile_X8Y9_N4BEG[10] ,
    \Tile_X8Y9_N4BEG[9] ,
    \Tile_X8Y9_N4BEG[8] ,
    \Tile_X8Y9_N4BEG[7] ,
    \Tile_X8Y9_N4BEG[6] ,
    \Tile_X8Y9_N4BEG[5] ,
    \Tile_X8Y9_N4BEG[4] ,
    \Tile_X8Y9_N4BEG[3] ,
    \Tile_X8Y9_N4BEG[2] ,
    \Tile_X8Y9_N4BEG[1] ,
    \Tile_X8Y9_N4BEG[0] }),
    .NN4BEG({\Tile_X8Y8_NN4BEG[15] ,
    \Tile_X8Y8_NN4BEG[14] ,
    \Tile_X8Y8_NN4BEG[13] ,
    \Tile_X8Y8_NN4BEG[12] ,
    \Tile_X8Y8_NN4BEG[11] ,
    \Tile_X8Y8_NN4BEG[10] ,
    \Tile_X8Y8_NN4BEG[9] ,
    \Tile_X8Y8_NN4BEG[8] ,
    \Tile_X8Y8_NN4BEG[7] ,
    \Tile_X8Y8_NN4BEG[6] ,
    \Tile_X8Y8_NN4BEG[5] ,
    \Tile_X8Y8_NN4BEG[4] ,
    \Tile_X8Y8_NN4BEG[3] ,
    \Tile_X8Y8_NN4BEG[2] ,
    \Tile_X8Y8_NN4BEG[1] ,
    \Tile_X8Y8_NN4BEG[0] }),
    .NN4END({\Tile_X8Y9_NN4BEG[15] ,
    \Tile_X8Y9_NN4BEG[14] ,
    \Tile_X8Y9_NN4BEG[13] ,
    \Tile_X8Y9_NN4BEG[12] ,
    \Tile_X8Y9_NN4BEG[11] ,
    \Tile_X8Y9_NN4BEG[10] ,
    \Tile_X8Y9_NN4BEG[9] ,
    \Tile_X8Y9_NN4BEG[8] ,
    \Tile_X8Y9_NN4BEG[7] ,
    \Tile_X8Y9_NN4BEG[6] ,
    \Tile_X8Y9_NN4BEG[5] ,
    \Tile_X8Y9_NN4BEG[4] ,
    \Tile_X8Y9_NN4BEG[3] ,
    \Tile_X8Y9_NN4BEG[2] ,
    \Tile_X8Y9_NN4BEG[1] ,
    \Tile_X8Y9_NN4BEG[0] }),
    .S1BEG({\Tile_X8Y8_S1BEG[3] ,
    \Tile_X8Y8_S1BEG[2] ,
    \Tile_X8Y8_S1BEG[1] ,
    \Tile_X8Y8_S1BEG[0] }),
    .S1END({\Tile_X8Y7_S1BEG[3] ,
    \Tile_X8Y7_S1BEG[2] ,
    \Tile_X8Y7_S1BEG[1] ,
    \Tile_X8Y7_S1BEG[0] }),
    .S2BEG({\Tile_X8Y8_S2BEG[7] ,
    \Tile_X8Y8_S2BEG[6] ,
    \Tile_X8Y8_S2BEG[5] ,
    \Tile_X8Y8_S2BEG[4] ,
    \Tile_X8Y8_S2BEG[3] ,
    \Tile_X8Y8_S2BEG[2] ,
    \Tile_X8Y8_S2BEG[1] ,
    \Tile_X8Y8_S2BEG[0] }),
    .S2BEGb({\Tile_X8Y8_S2BEGb[7] ,
    \Tile_X8Y8_S2BEGb[6] ,
    \Tile_X8Y8_S2BEGb[5] ,
    \Tile_X8Y8_S2BEGb[4] ,
    \Tile_X8Y8_S2BEGb[3] ,
    \Tile_X8Y8_S2BEGb[2] ,
    \Tile_X8Y8_S2BEGb[1] ,
    \Tile_X8Y8_S2BEGb[0] }),
    .S2END({\Tile_X8Y7_S2BEGb[7] ,
    \Tile_X8Y7_S2BEGb[6] ,
    \Tile_X8Y7_S2BEGb[5] ,
    \Tile_X8Y7_S2BEGb[4] ,
    \Tile_X8Y7_S2BEGb[3] ,
    \Tile_X8Y7_S2BEGb[2] ,
    \Tile_X8Y7_S2BEGb[1] ,
    \Tile_X8Y7_S2BEGb[0] }),
    .S2MID({\Tile_X8Y7_S2BEG[7] ,
    \Tile_X8Y7_S2BEG[6] ,
    \Tile_X8Y7_S2BEG[5] ,
    \Tile_X8Y7_S2BEG[4] ,
    \Tile_X8Y7_S2BEG[3] ,
    \Tile_X8Y7_S2BEG[2] ,
    \Tile_X8Y7_S2BEG[1] ,
    \Tile_X8Y7_S2BEG[0] }),
    .S4BEG({\Tile_X8Y8_S4BEG[15] ,
    \Tile_X8Y8_S4BEG[14] ,
    \Tile_X8Y8_S4BEG[13] ,
    \Tile_X8Y8_S4BEG[12] ,
    \Tile_X8Y8_S4BEG[11] ,
    \Tile_X8Y8_S4BEG[10] ,
    \Tile_X8Y8_S4BEG[9] ,
    \Tile_X8Y8_S4BEG[8] ,
    \Tile_X8Y8_S4BEG[7] ,
    \Tile_X8Y8_S4BEG[6] ,
    \Tile_X8Y8_S4BEG[5] ,
    \Tile_X8Y8_S4BEG[4] ,
    \Tile_X8Y8_S4BEG[3] ,
    \Tile_X8Y8_S4BEG[2] ,
    \Tile_X8Y8_S4BEG[1] ,
    \Tile_X8Y8_S4BEG[0] }),
    .S4END({\Tile_X8Y7_S4BEG[15] ,
    \Tile_X8Y7_S4BEG[14] ,
    \Tile_X8Y7_S4BEG[13] ,
    \Tile_X8Y7_S4BEG[12] ,
    \Tile_X8Y7_S4BEG[11] ,
    \Tile_X8Y7_S4BEG[10] ,
    \Tile_X8Y7_S4BEG[9] ,
    \Tile_X8Y7_S4BEG[8] ,
    \Tile_X8Y7_S4BEG[7] ,
    \Tile_X8Y7_S4BEG[6] ,
    \Tile_X8Y7_S4BEG[5] ,
    \Tile_X8Y7_S4BEG[4] ,
    \Tile_X8Y7_S4BEG[3] ,
    \Tile_X8Y7_S4BEG[2] ,
    \Tile_X8Y7_S4BEG[1] ,
    \Tile_X8Y7_S4BEG[0] }),
    .SS4BEG({\Tile_X8Y8_SS4BEG[15] ,
    \Tile_X8Y8_SS4BEG[14] ,
    \Tile_X8Y8_SS4BEG[13] ,
    \Tile_X8Y8_SS4BEG[12] ,
    \Tile_X8Y8_SS4BEG[11] ,
    \Tile_X8Y8_SS4BEG[10] ,
    \Tile_X8Y8_SS4BEG[9] ,
    \Tile_X8Y8_SS4BEG[8] ,
    \Tile_X8Y8_SS4BEG[7] ,
    \Tile_X8Y8_SS4BEG[6] ,
    \Tile_X8Y8_SS4BEG[5] ,
    \Tile_X8Y8_SS4BEG[4] ,
    \Tile_X8Y8_SS4BEG[3] ,
    \Tile_X8Y8_SS4BEG[2] ,
    \Tile_X8Y8_SS4BEG[1] ,
    \Tile_X8Y8_SS4BEG[0] }),
    .SS4END({\Tile_X8Y7_SS4BEG[15] ,
    \Tile_X8Y7_SS4BEG[14] ,
    \Tile_X8Y7_SS4BEG[13] ,
    \Tile_X8Y7_SS4BEG[12] ,
    \Tile_X8Y7_SS4BEG[11] ,
    \Tile_X8Y7_SS4BEG[10] ,
    \Tile_X8Y7_SS4BEG[9] ,
    \Tile_X8Y7_SS4BEG[8] ,
    \Tile_X8Y7_SS4BEG[7] ,
    \Tile_X8Y7_SS4BEG[6] ,
    \Tile_X8Y7_SS4BEG[5] ,
    \Tile_X8Y7_SS4BEG[4] ,
    \Tile_X8Y7_SS4BEG[3] ,
    \Tile_X8Y7_SS4BEG[2] ,
    \Tile_X8Y7_SS4BEG[1] ,
    \Tile_X8Y7_SS4BEG[0] }),
    .W1BEG({\Tile_X8Y8_W1BEG[3] ,
    \Tile_X8Y8_W1BEG[2] ,
    \Tile_X8Y8_W1BEG[1] ,
    \Tile_X8Y8_W1BEG[0] }),
    .W1END({\Tile_X9Y8_W1BEG[3] ,
    \Tile_X9Y8_W1BEG[2] ,
    \Tile_X9Y8_W1BEG[1] ,
    \Tile_X9Y8_W1BEG[0] }),
    .W2BEG({\Tile_X8Y8_W2BEG[7] ,
    \Tile_X8Y8_W2BEG[6] ,
    \Tile_X8Y8_W2BEG[5] ,
    \Tile_X8Y8_W2BEG[4] ,
    \Tile_X8Y8_W2BEG[3] ,
    \Tile_X8Y8_W2BEG[2] ,
    \Tile_X8Y8_W2BEG[1] ,
    \Tile_X8Y8_W2BEG[0] }),
    .W2BEGb({\Tile_X8Y8_W2BEGb[7] ,
    \Tile_X8Y8_W2BEGb[6] ,
    \Tile_X8Y8_W2BEGb[5] ,
    \Tile_X8Y8_W2BEGb[4] ,
    \Tile_X8Y8_W2BEGb[3] ,
    \Tile_X8Y8_W2BEGb[2] ,
    \Tile_X8Y8_W2BEGb[1] ,
    \Tile_X8Y8_W2BEGb[0] }),
    .W2END({\Tile_X9Y8_W2BEGb[7] ,
    \Tile_X9Y8_W2BEGb[6] ,
    \Tile_X9Y8_W2BEGb[5] ,
    \Tile_X9Y8_W2BEGb[4] ,
    \Tile_X9Y8_W2BEGb[3] ,
    \Tile_X9Y8_W2BEGb[2] ,
    \Tile_X9Y8_W2BEGb[1] ,
    \Tile_X9Y8_W2BEGb[0] }),
    .W2MID({\Tile_X9Y8_W2BEG[7] ,
    \Tile_X9Y8_W2BEG[6] ,
    \Tile_X9Y8_W2BEG[5] ,
    \Tile_X9Y8_W2BEG[4] ,
    \Tile_X9Y8_W2BEG[3] ,
    \Tile_X9Y8_W2BEG[2] ,
    \Tile_X9Y8_W2BEG[1] ,
    \Tile_X9Y8_W2BEG[0] }),
    .W6BEG({\Tile_X8Y8_W6BEG[11] ,
    \Tile_X8Y8_W6BEG[10] ,
    \Tile_X8Y8_W6BEG[9] ,
    \Tile_X8Y8_W6BEG[8] ,
    \Tile_X8Y8_W6BEG[7] ,
    \Tile_X8Y8_W6BEG[6] ,
    \Tile_X8Y8_W6BEG[5] ,
    \Tile_X8Y8_W6BEG[4] ,
    \Tile_X8Y8_W6BEG[3] ,
    \Tile_X8Y8_W6BEG[2] ,
    \Tile_X8Y8_W6BEG[1] ,
    \Tile_X8Y8_W6BEG[0] }),
    .W6END({\Tile_X9Y8_W6BEG[11] ,
    \Tile_X9Y8_W6BEG[10] ,
    \Tile_X9Y8_W6BEG[9] ,
    \Tile_X9Y8_W6BEG[8] ,
    \Tile_X9Y8_W6BEG[7] ,
    \Tile_X9Y8_W6BEG[6] ,
    \Tile_X9Y8_W6BEG[5] ,
    \Tile_X9Y8_W6BEG[4] ,
    \Tile_X9Y8_W6BEG[3] ,
    \Tile_X9Y8_W6BEG[2] ,
    \Tile_X9Y8_W6BEG[1] ,
    \Tile_X9Y8_W6BEG[0] }),
    .WW4BEG({\Tile_X8Y8_WW4BEG[15] ,
    \Tile_X8Y8_WW4BEG[14] ,
    \Tile_X8Y8_WW4BEG[13] ,
    \Tile_X8Y8_WW4BEG[12] ,
    \Tile_X8Y8_WW4BEG[11] ,
    \Tile_X8Y8_WW4BEG[10] ,
    \Tile_X8Y8_WW4BEG[9] ,
    \Tile_X8Y8_WW4BEG[8] ,
    \Tile_X8Y8_WW4BEG[7] ,
    \Tile_X8Y8_WW4BEG[6] ,
    \Tile_X8Y8_WW4BEG[5] ,
    \Tile_X8Y8_WW4BEG[4] ,
    \Tile_X8Y8_WW4BEG[3] ,
    \Tile_X8Y8_WW4BEG[2] ,
    \Tile_X8Y8_WW4BEG[1] ,
    \Tile_X8Y8_WW4BEG[0] }),
    .WW4END({\Tile_X9Y8_WW4BEG[15] ,
    \Tile_X9Y8_WW4BEG[14] ,
    \Tile_X9Y8_WW4BEG[13] ,
    \Tile_X9Y8_WW4BEG[12] ,
    \Tile_X9Y8_WW4BEG[11] ,
    \Tile_X9Y8_WW4BEG[10] ,
    \Tile_X9Y8_WW4BEG[9] ,
    \Tile_X9Y8_WW4BEG[8] ,
    \Tile_X9Y8_WW4BEG[7] ,
    \Tile_X9Y8_WW4BEG[6] ,
    \Tile_X9Y8_WW4BEG[5] ,
    \Tile_X9Y8_WW4BEG[4] ,
    \Tile_X9Y8_WW4BEG[3] ,
    \Tile_X9Y8_WW4BEG[2] ,
    \Tile_X9Y8_WW4BEG[1] ,
    \Tile_X9Y8_WW4BEG[0] }));
 LUT4AB Tile_X8Y9_LUT4AB (.Ci(Tile_X8Y10_Co),
    .Co(Tile_X8Y9_Co),
    .UserCLK(Tile_X8Y10_UserCLKo),
    .UserCLKo(Tile_X8Y9_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X8Y9_E1BEG[3] ,
    \Tile_X8Y9_E1BEG[2] ,
    \Tile_X8Y9_E1BEG[1] ,
    \Tile_X8Y9_E1BEG[0] }),
    .E1END({\Tile_X7Y9_E1BEG[3] ,
    \Tile_X7Y9_E1BEG[2] ,
    \Tile_X7Y9_E1BEG[1] ,
    \Tile_X7Y9_E1BEG[0] }),
    .E2BEG({\Tile_X8Y9_E2BEG[7] ,
    \Tile_X8Y9_E2BEG[6] ,
    \Tile_X8Y9_E2BEG[5] ,
    \Tile_X8Y9_E2BEG[4] ,
    \Tile_X8Y9_E2BEG[3] ,
    \Tile_X8Y9_E2BEG[2] ,
    \Tile_X8Y9_E2BEG[1] ,
    \Tile_X8Y9_E2BEG[0] }),
    .E2BEGb({\Tile_X8Y9_E2BEGb[7] ,
    \Tile_X8Y9_E2BEGb[6] ,
    \Tile_X8Y9_E2BEGb[5] ,
    \Tile_X8Y9_E2BEGb[4] ,
    \Tile_X8Y9_E2BEGb[3] ,
    \Tile_X8Y9_E2BEGb[2] ,
    \Tile_X8Y9_E2BEGb[1] ,
    \Tile_X8Y9_E2BEGb[0] }),
    .E2END({\Tile_X7Y9_E2BEGb[7] ,
    \Tile_X7Y9_E2BEGb[6] ,
    \Tile_X7Y9_E2BEGb[5] ,
    \Tile_X7Y9_E2BEGb[4] ,
    \Tile_X7Y9_E2BEGb[3] ,
    \Tile_X7Y9_E2BEGb[2] ,
    \Tile_X7Y9_E2BEGb[1] ,
    \Tile_X7Y9_E2BEGb[0] }),
    .E2MID({\Tile_X7Y9_E2BEG[7] ,
    \Tile_X7Y9_E2BEG[6] ,
    \Tile_X7Y9_E2BEG[5] ,
    \Tile_X7Y9_E2BEG[4] ,
    \Tile_X7Y9_E2BEG[3] ,
    \Tile_X7Y9_E2BEG[2] ,
    \Tile_X7Y9_E2BEG[1] ,
    \Tile_X7Y9_E2BEG[0] }),
    .E6BEG({\Tile_X8Y9_E6BEG[11] ,
    \Tile_X8Y9_E6BEG[10] ,
    \Tile_X8Y9_E6BEG[9] ,
    \Tile_X8Y9_E6BEG[8] ,
    \Tile_X8Y9_E6BEG[7] ,
    \Tile_X8Y9_E6BEG[6] ,
    \Tile_X8Y9_E6BEG[5] ,
    \Tile_X8Y9_E6BEG[4] ,
    \Tile_X8Y9_E6BEG[3] ,
    \Tile_X8Y9_E6BEG[2] ,
    \Tile_X8Y9_E6BEG[1] ,
    \Tile_X8Y9_E6BEG[0] }),
    .E6END({\Tile_X7Y9_E6BEG[11] ,
    \Tile_X7Y9_E6BEG[10] ,
    \Tile_X7Y9_E6BEG[9] ,
    \Tile_X7Y9_E6BEG[8] ,
    \Tile_X7Y9_E6BEG[7] ,
    \Tile_X7Y9_E6BEG[6] ,
    \Tile_X7Y9_E6BEG[5] ,
    \Tile_X7Y9_E6BEG[4] ,
    \Tile_X7Y9_E6BEG[3] ,
    \Tile_X7Y9_E6BEG[2] ,
    \Tile_X7Y9_E6BEG[1] ,
    \Tile_X7Y9_E6BEG[0] }),
    .EE4BEG({\Tile_X8Y9_EE4BEG[15] ,
    \Tile_X8Y9_EE4BEG[14] ,
    \Tile_X8Y9_EE4BEG[13] ,
    \Tile_X8Y9_EE4BEG[12] ,
    \Tile_X8Y9_EE4BEG[11] ,
    \Tile_X8Y9_EE4BEG[10] ,
    \Tile_X8Y9_EE4BEG[9] ,
    \Tile_X8Y9_EE4BEG[8] ,
    \Tile_X8Y9_EE4BEG[7] ,
    \Tile_X8Y9_EE4BEG[6] ,
    \Tile_X8Y9_EE4BEG[5] ,
    \Tile_X8Y9_EE4BEG[4] ,
    \Tile_X8Y9_EE4BEG[3] ,
    \Tile_X8Y9_EE4BEG[2] ,
    \Tile_X8Y9_EE4BEG[1] ,
    \Tile_X8Y9_EE4BEG[0] }),
    .EE4END({\Tile_X7Y9_EE4BEG[15] ,
    \Tile_X7Y9_EE4BEG[14] ,
    \Tile_X7Y9_EE4BEG[13] ,
    \Tile_X7Y9_EE4BEG[12] ,
    \Tile_X7Y9_EE4BEG[11] ,
    \Tile_X7Y9_EE4BEG[10] ,
    \Tile_X7Y9_EE4BEG[9] ,
    \Tile_X7Y9_EE4BEG[8] ,
    \Tile_X7Y9_EE4BEG[7] ,
    \Tile_X7Y9_EE4BEG[6] ,
    \Tile_X7Y9_EE4BEG[5] ,
    \Tile_X7Y9_EE4BEG[4] ,
    \Tile_X7Y9_EE4BEG[3] ,
    \Tile_X7Y9_EE4BEG[2] ,
    \Tile_X7Y9_EE4BEG[1] ,
    \Tile_X7Y9_EE4BEG[0] }),
    .FrameData({\Tile_X7Y9_FrameData_O[31] ,
    \Tile_X7Y9_FrameData_O[30] ,
    \Tile_X7Y9_FrameData_O[29] ,
    \Tile_X7Y9_FrameData_O[28] ,
    \Tile_X7Y9_FrameData_O[27] ,
    \Tile_X7Y9_FrameData_O[26] ,
    \Tile_X7Y9_FrameData_O[25] ,
    \Tile_X7Y9_FrameData_O[24] ,
    \Tile_X7Y9_FrameData_O[23] ,
    \Tile_X7Y9_FrameData_O[22] ,
    \Tile_X7Y9_FrameData_O[21] ,
    \Tile_X7Y9_FrameData_O[20] ,
    \Tile_X7Y9_FrameData_O[19] ,
    \Tile_X7Y9_FrameData_O[18] ,
    \Tile_X7Y9_FrameData_O[17] ,
    \Tile_X7Y9_FrameData_O[16] ,
    \Tile_X7Y9_FrameData_O[15] ,
    \Tile_X7Y9_FrameData_O[14] ,
    \Tile_X7Y9_FrameData_O[13] ,
    \Tile_X7Y9_FrameData_O[12] ,
    \Tile_X7Y9_FrameData_O[11] ,
    \Tile_X7Y9_FrameData_O[10] ,
    \Tile_X7Y9_FrameData_O[9] ,
    \Tile_X7Y9_FrameData_O[8] ,
    \Tile_X7Y9_FrameData_O[7] ,
    \Tile_X7Y9_FrameData_O[6] ,
    \Tile_X7Y9_FrameData_O[5] ,
    \Tile_X7Y9_FrameData_O[4] ,
    \Tile_X7Y9_FrameData_O[3] ,
    \Tile_X7Y9_FrameData_O[2] ,
    \Tile_X7Y9_FrameData_O[1] ,
    \Tile_X7Y9_FrameData_O[0] }),
    .FrameData_O({\Tile_X8Y9_FrameData_O[31] ,
    \Tile_X8Y9_FrameData_O[30] ,
    \Tile_X8Y9_FrameData_O[29] ,
    \Tile_X8Y9_FrameData_O[28] ,
    \Tile_X8Y9_FrameData_O[27] ,
    \Tile_X8Y9_FrameData_O[26] ,
    \Tile_X8Y9_FrameData_O[25] ,
    \Tile_X8Y9_FrameData_O[24] ,
    \Tile_X8Y9_FrameData_O[23] ,
    \Tile_X8Y9_FrameData_O[22] ,
    \Tile_X8Y9_FrameData_O[21] ,
    \Tile_X8Y9_FrameData_O[20] ,
    \Tile_X8Y9_FrameData_O[19] ,
    \Tile_X8Y9_FrameData_O[18] ,
    \Tile_X8Y9_FrameData_O[17] ,
    \Tile_X8Y9_FrameData_O[16] ,
    \Tile_X8Y9_FrameData_O[15] ,
    \Tile_X8Y9_FrameData_O[14] ,
    \Tile_X8Y9_FrameData_O[13] ,
    \Tile_X8Y9_FrameData_O[12] ,
    \Tile_X8Y9_FrameData_O[11] ,
    \Tile_X8Y9_FrameData_O[10] ,
    \Tile_X8Y9_FrameData_O[9] ,
    \Tile_X8Y9_FrameData_O[8] ,
    \Tile_X8Y9_FrameData_O[7] ,
    \Tile_X8Y9_FrameData_O[6] ,
    \Tile_X8Y9_FrameData_O[5] ,
    \Tile_X8Y9_FrameData_O[4] ,
    \Tile_X8Y9_FrameData_O[3] ,
    \Tile_X8Y9_FrameData_O[2] ,
    \Tile_X8Y9_FrameData_O[1] ,
    \Tile_X8Y9_FrameData_O[0] }),
    .FrameStrobe({\Tile_X8Y10_FrameStrobe_O[19] ,
    \Tile_X8Y10_FrameStrobe_O[18] ,
    \Tile_X8Y10_FrameStrobe_O[17] ,
    \Tile_X8Y10_FrameStrobe_O[16] ,
    \Tile_X8Y10_FrameStrobe_O[15] ,
    \Tile_X8Y10_FrameStrobe_O[14] ,
    \Tile_X8Y10_FrameStrobe_O[13] ,
    \Tile_X8Y10_FrameStrobe_O[12] ,
    \Tile_X8Y10_FrameStrobe_O[11] ,
    \Tile_X8Y10_FrameStrobe_O[10] ,
    \Tile_X8Y10_FrameStrobe_O[9] ,
    \Tile_X8Y10_FrameStrobe_O[8] ,
    \Tile_X8Y10_FrameStrobe_O[7] ,
    \Tile_X8Y10_FrameStrobe_O[6] ,
    \Tile_X8Y10_FrameStrobe_O[5] ,
    \Tile_X8Y10_FrameStrobe_O[4] ,
    \Tile_X8Y10_FrameStrobe_O[3] ,
    \Tile_X8Y10_FrameStrobe_O[2] ,
    \Tile_X8Y10_FrameStrobe_O[1] ,
    \Tile_X8Y10_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X8Y9_FrameStrobe_O[19] ,
    \Tile_X8Y9_FrameStrobe_O[18] ,
    \Tile_X8Y9_FrameStrobe_O[17] ,
    \Tile_X8Y9_FrameStrobe_O[16] ,
    \Tile_X8Y9_FrameStrobe_O[15] ,
    \Tile_X8Y9_FrameStrobe_O[14] ,
    \Tile_X8Y9_FrameStrobe_O[13] ,
    \Tile_X8Y9_FrameStrobe_O[12] ,
    \Tile_X8Y9_FrameStrobe_O[11] ,
    \Tile_X8Y9_FrameStrobe_O[10] ,
    \Tile_X8Y9_FrameStrobe_O[9] ,
    \Tile_X8Y9_FrameStrobe_O[8] ,
    \Tile_X8Y9_FrameStrobe_O[7] ,
    \Tile_X8Y9_FrameStrobe_O[6] ,
    \Tile_X8Y9_FrameStrobe_O[5] ,
    \Tile_X8Y9_FrameStrobe_O[4] ,
    \Tile_X8Y9_FrameStrobe_O[3] ,
    \Tile_X8Y9_FrameStrobe_O[2] ,
    \Tile_X8Y9_FrameStrobe_O[1] ,
    \Tile_X8Y9_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X8Y9_N1BEG[3] ,
    \Tile_X8Y9_N1BEG[2] ,
    \Tile_X8Y9_N1BEG[1] ,
    \Tile_X8Y9_N1BEG[0] }),
    .N1END({\Tile_X8Y10_N1BEG[3] ,
    \Tile_X8Y10_N1BEG[2] ,
    \Tile_X8Y10_N1BEG[1] ,
    \Tile_X8Y10_N1BEG[0] }),
    .N2BEG({\Tile_X8Y9_N2BEG[7] ,
    \Tile_X8Y9_N2BEG[6] ,
    \Tile_X8Y9_N2BEG[5] ,
    \Tile_X8Y9_N2BEG[4] ,
    \Tile_X8Y9_N2BEG[3] ,
    \Tile_X8Y9_N2BEG[2] ,
    \Tile_X8Y9_N2BEG[1] ,
    \Tile_X8Y9_N2BEG[0] }),
    .N2BEGb({\Tile_X8Y9_N2BEGb[7] ,
    \Tile_X8Y9_N2BEGb[6] ,
    \Tile_X8Y9_N2BEGb[5] ,
    \Tile_X8Y9_N2BEGb[4] ,
    \Tile_X8Y9_N2BEGb[3] ,
    \Tile_X8Y9_N2BEGb[2] ,
    \Tile_X8Y9_N2BEGb[1] ,
    \Tile_X8Y9_N2BEGb[0] }),
    .N2END({\Tile_X8Y10_N2BEGb[7] ,
    \Tile_X8Y10_N2BEGb[6] ,
    \Tile_X8Y10_N2BEGb[5] ,
    \Tile_X8Y10_N2BEGb[4] ,
    \Tile_X8Y10_N2BEGb[3] ,
    \Tile_X8Y10_N2BEGb[2] ,
    \Tile_X8Y10_N2BEGb[1] ,
    \Tile_X8Y10_N2BEGb[0] }),
    .N2MID({\Tile_X8Y10_N2BEG[7] ,
    \Tile_X8Y10_N2BEG[6] ,
    \Tile_X8Y10_N2BEG[5] ,
    \Tile_X8Y10_N2BEG[4] ,
    \Tile_X8Y10_N2BEG[3] ,
    \Tile_X8Y10_N2BEG[2] ,
    \Tile_X8Y10_N2BEG[1] ,
    \Tile_X8Y10_N2BEG[0] }),
    .N4BEG({\Tile_X8Y9_N4BEG[15] ,
    \Tile_X8Y9_N4BEG[14] ,
    \Tile_X8Y9_N4BEG[13] ,
    \Tile_X8Y9_N4BEG[12] ,
    \Tile_X8Y9_N4BEG[11] ,
    \Tile_X8Y9_N4BEG[10] ,
    \Tile_X8Y9_N4BEG[9] ,
    \Tile_X8Y9_N4BEG[8] ,
    \Tile_X8Y9_N4BEG[7] ,
    \Tile_X8Y9_N4BEG[6] ,
    \Tile_X8Y9_N4BEG[5] ,
    \Tile_X8Y9_N4BEG[4] ,
    \Tile_X8Y9_N4BEG[3] ,
    \Tile_X8Y9_N4BEG[2] ,
    \Tile_X8Y9_N4BEG[1] ,
    \Tile_X8Y9_N4BEG[0] }),
    .N4END({\Tile_X8Y10_N4BEG[15] ,
    \Tile_X8Y10_N4BEG[14] ,
    \Tile_X8Y10_N4BEG[13] ,
    \Tile_X8Y10_N4BEG[12] ,
    \Tile_X8Y10_N4BEG[11] ,
    \Tile_X8Y10_N4BEG[10] ,
    \Tile_X8Y10_N4BEG[9] ,
    \Tile_X8Y10_N4BEG[8] ,
    \Tile_X8Y10_N4BEG[7] ,
    \Tile_X8Y10_N4BEG[6] ,
    \Tile_X8Y10_N4BEG[5] ,
    \Tile_X8Y10_N4BEG[4] ,
    \Tile_X8Y10_N4BEG[3] ,
    \Tile_X8Y10_N4BEG[2] ,
    \Tile_X8Y10_N4BEG[1] ,
    \Tile_X8Y10_N4BEG[0] }),
    .NN4BEG({\Tile_X8Y9_NN4BEG[15] ,
    \Tile_X8Y9_NN4BEG[14] ,
    \Tile_X8Y9_NN4BEG[13] ,
    \Tile_X8Y9_NN4BEG[12] ,
    \Tile_X8Y9_NN4BEG[11] ,
    \Tile_X8Y9_NN4BEG[10] ,
    \Tile_X8Y9_NN4BEG[9] ,
    \Tile_X8Y9_NN4BEG[8] ,
    \Tile_X8Y9_NN4BEG[7] ,
    \Tile_X8Y9_NN4BEG[6] ,
    \Tile_X8Y9_NN4BEG[5] ,
    \Tile_X8Y9_NN4BEG[4] ,
    \Tile_X8Y9_NN4BEG[3] ,
    \Tile_X8Y9_NN4BEG[2] ,
    \Tile_X8Y9_NN4BEG[1] ,
    \Tile_X8Y9_NN4BEG[0] }),
    .NN4END({\Tile_X8Y10_NN4BEG[15] ,
    \Tile_X8Y10_NN4BEG[14] ,
    \Tile_X8Y10_NN4BEG[13] ,
    \Tile_X8Y10_NN4BEG[12] ,
    \Tile_X8Y10_NN4BEG[11] ,
    \Tile_X8Y10_NN4BEG[10] ,
    \Tile_X8Y10_NN4BEG[9] ,
    \Tile_X8Y10_NN4BEG[8] ,
    \Tile_X8Y10_NN4BEG[7] ,
    \Tile_X8Y10_NN4BEG[6] ,
    \Tile_X8Y10_NN4BEG[5] ,
    \Tile_X8Y10_NN4BEG[4] ,
    \Tile_X8Y10_NN4BEG[3] ,
    \Tile_X8Y10_NN4BEG[2] ,
    \Tile_X8Y10_NN4BEG[1] ,
    \Tile_X8Y10_NN4BEG[0] }),
    .S1BEG({\Tile_X8Y9_S1BEG[3] ,
    \Tile_X8Y9_S1BEG[2] ,
    \Tile_X8Y9_S1BEG[1] ,
    \Tile_X8Y9_S1BEG[0] }),
    .S1END({\Tile_X8Y8_S1BEG[3] ,
    \Tile_X8Y8_S1BEG[2] ,
    \Tile_X8Y8_S1BEG[1] ,
    \Tile_X8Y8_S1BEG[0] }),
    .S2BEG({\Tile_X8Y9_S2BEG[7] ,
    \Tile_X8Y9_S2BEG[6] ,
    \Tile_X8Y9_S2BEG[5] ,
    \Tile_X8Y9_S2BEG[4] ,
    \Tile_X8Y9_S2BEG[3] ,
    \Tile_X8Y9_S2BEG[2] ,
    \Tile_X8Y9_S2BEG[1] ,
    \Tile_X8Y9_S2BEG[0] }),
    .S2BEGb({\Tile_X8Y9_S2BEGb[7] ,
    \Tile_X8Y9_S2BEGb[6] ,
    \Tile_X8Y9_S2BEGb[5] ,
    \Tile_X8Y9_S2BEGb[4] ,
    \Tile_X8Y9_S2BEGb[3] ,
    \Tile_X8Y9_S2BEGb[2] ,
    \Tile_X8Y9_S2BEGb[1] ,
    \Tile_X8Y9_S2BEGb[0] }),
    .S2END({\Tile_X8Y8_S2BEGb[7] ,
    \Tile_X8Y8_S2BEGb[6] ,
    \Tile_X8Y8_S2BEGb[5] ,
    \Tile_X8Y8_S2BEGb[4] ,
    \Tile_X8Y8_S2BEGb[3] ,
    \Tile_X8Y8_S2BEGb[2] ,
    \Tile_X8Y8_S2BEGb[1] ,
    \Tile_X8Y8_S2BEGb[0] }),
    .S2MID({\Tile_X8Y8_S2BEG[7] ,
    \Tile_X8Y8_S2BEG[6] ,
    \Tile_X8Y8_S2BEG[5] ,
    \Tile_X8Y8_S2BEG[4] ,
    \Tile_X8Y8_S2BEG[3] ,
    \Tile_X8Y8_S2BEG[2] ,
    \Tile_X8Y8_S2BEG[1] ,
    \Tile_X8Y8_S2BEG[0] }),
    .S4BEG({\Tile_X8Y9_S4BEG[15] ,
    \Tile_X8Y9_S4BEG[14] ,
    \Tile_X8Y9_S4BEG[13] ,
    \Tile_X8Y9_S4BEG[12] ,
    \Tile_X8Y9_S4BEG[11] ,
    \Tile_X8Y9_S4BEG[10] ,
    \Tile_X8Y9_S4BEG[9] ,
    \Tile_X8Y9_S4BEG[8] ,
    \Tile_X8Y9_S4BEG[7] ,
    \Tile_X8Y9_S4BEG[6] ,
    \Tile_X8Y9_S4BEG[5] ,
    \Tile_X8Y9_S4BEG[4] ,
    \Tile_X8Y9_S4BEG[3] ,
    \Tile_X8Y9_S4BEG[2] ,
    \Tile_X8Y9_S4BEG[1] ,
    \Tile_X8Y9_S4BEG[0] }),
    .S4END({\Tile_X8Y8_S4BEG[15] ,
    \Tile_X8Y8_S4BEG[14] ,
    \Tile_X8Y8_S4BEG[13] ,
    \Tile_X8Y8_S4BEG[12] ,
    \Tile_X8Y8_S4BEG[11] ,
    \Tile_X8Y8_S4BEG[10] ,
    \Tile_X8Y8_S4BEG[9] ,
    \Tile_X8Y8_S4BEG[8] ,
    \Tile_X8Y8_S4BEG[7] ,
    \Tile_X8Y8_S4BEG[6] ,
    \Tile_X8Y8_S4BEG[5] ,
    \Tile_X8Y8_S4BEG[4] ,
    \Tile_X8Y8_S4BEG[3] ,
    \Tile_X8Y8_S4BEG[2] ,
    \Tile_X8Y8_S4BEG[1] ,
    \Tile_X8Y8_S4BEG[0] }),
    .SS4BEG({\Tile_X8Y9_SS4BEG[15] ,
    \Tile_X8Y9_SS4BEG[14] ,
    \Tile_X8Y9_SS4BEG[13] ,
    \Tile_X8Y9_SS4BEG[12] ,
    \Tile_X8Y9_SS4BEG[11] ,
    \Tile_X8Y9_SS4BEG[10] ,
    \Tile_X8Y9_SS4BEG[9] ,
    \Tile_X8Y9_SS4BEG[8] ,
    \Tile_X8Y9_SS4BEG[7] ,
    \Tile_X8Y9_SS4BEG[6] ,
    \Tile_X8Y9_SS4BEG[5] ,
    \Tile_X8Y9_SS4BEG[4] ,
    \Tile_X8Y9_SS4BEG[3] ,
    \Tile_X8Y9_SS4BEG[2] ,
    \Tile_X8Y9_SS4BEG[1] ,
    \Tile_X8Y9_SS4BEG[0] }),
    .SS4END({\Tile_X8Y8_SS4BEG[15] ,
    \Tile_X8Y8_SS4BEG[14] ,
    \Tile_X8Y8_SS4BEG[13] ,
    \Tile_X8Y8_SS4BEG[12] ,
    \Tile_X8Y8_SS4BEG[11] ,
    \Tile_X8Y8_SS4BEG[10] ,
    \Tile_X8Y8_SS4BEG[9] ,
    \Tile_X8Y8_SS4BEG[8] ,
    \Tile_X8Y8_SS4BEG[7] ,
    \Tile_X8Y8_SS4BEG[6] ,
    \Tile_X8Y8_SS4BEG[5] ,
    \Tile_X8Y8_SS4BEG[4] ,
    \Tile_X8Y8_SS4BEG[3] ,
    \Tile_X8Y8_SS4BEG[2] ,
    \Tile_X8Y8_SS4BEG[1] ,
    \Tile_X8Y8_SS4BEG[0] }),
    .W1BEG({\Tile_X8Y9_W1BEG[3] ,
    \Tile_X8Y9_W1BEG[2] ,
    \Tile_X8Y9_W1BEG[1] ,
    \Tile_X8Y9_W1BEG[0] }),
    .W1END({\Tile_X9Y9_W1BEG[3] ,
    \Tile_X9Y9_W1BEG[2] ,
    \Tile_X9Y9_W1BEG[1] ,
    \Tile_X9Y9_W1BEG[0] }),
    .W2BEG({\Tile_X8Y9_W2BEG[7] ,
    \Tile_X8Y9_W2BEG[6] ,
    \Tile_X8Y9_W2BEG[5] ,
    \Tile_X8Y9_W2BEG[4] ,
    \Tile_X8Y9_W2BEG[3] ,
    \Tile_X8Y9_W2BEG[2] ,
    \Tile_X8Y9_W2BEG[1] ,
    \Tile_X8Y9_W2BEG[0] }),
    .W2BEGb({\Tile_X8Y9_W2BEGb[7] ,
    \Tile_X8Y9_W2BEGb[6] ,
    \Tile_X8Y9_W2BEGb[5] ,
    \Tile_X8Y9_W2BEGb[4] ,
    \Tile_X8Y9_W2BEGb[3] ,
    \Tile_X8Y9_W2BEGb[2] ,
    \Tile_X8Y9_W2BEGb[1] ,
    \Tile_X8Y9_W2BEGb[0] }),
    .W2END({\Tile_X9Y9_W2BEGb[7] ,
    \Tile_X9Y9_W2BEGb[6] ,
    \Tile_X9Y9_W2BEGb[5] ,
    \Tile_X9Y9_W2BEGb[4] ,
    \Tile_X9Y9_W2BEGb[3] ,
    \Tile_X9Y9_W2BEGb[2] ,
    \Tile_X9Y9_W2BEGb[1] ,
    \Tile_X9Y9_W2BEGb[0] }),
    .W2MID({\Tile_X9Y9_W2BEG[7] ,
    \Tile_X9Y9_W2BEG[6] ,
    \Tile_X9Y9_W2BEG[5] ,
    \Tile_X9Y9_W2BEG[4] ,
    \Tile_X9Y9_W2BEG[3] ,
    \Tile_X9Y9_W2BEG[2] ,
    \Tile_X9Y9_W2BEG[1] ,
    \Tile_X9Y9_W2BEG[0] }),
    .W6BEG({\Tile_X8Y9_W6BEG[11] ,
    \Tile_X8Y9_W6BEG[10] ,
    \Tile_X8Y9_W6BEG[9] ,
    \Tile_X8Y9_W6BEG[8] ,
    \Tile_X8Y9_W6BEG[7] ,
    \Tile_X8Y9_W6BEG[6] ,
    \Tile_X8Y9_W6BEG[5] ,
    \Tile_X8Y9_W6BEG[4] ,
    \Tile_X8Y9_W6BEG[3] ,
    \Tile_X8Y9_W6BEG[2] ,
    \Tile_X8Y9_W6BEG[1] ,
    \Tile_X8Y9_W6BEG[0] }),
    .W6END({\Tile_X9Y9_W6BEG[11] ,
    \Tile_X9Y9_W6BEG[10] ,
    \Tile_X9Y9_W6BEG[9] ,
    \Tile_X9Y9_W6BEG[8] ,
    \Tile_X9Y9_W6BEG[7] ,
    \Tile_X9Y9_W6BEG[6] ,
    \Tile_X9Y9_W6BEG[5] ,
    \Tile_X9Y9_W6BEG[4] ,
    \Tile_X9Y9_W6BEG[3] ,
    \Tile_X9Y9_W6BEG[2] ,
    \Tile_X9Y9_W6BEG[1] ,
    \Tile_X9Y9_W6BEG[0] }),
    .WW4BEG({\Tile_X8Y9_WW4BEG[15] ,
    \Tile_X8Y9_WW4BEG[14] ,
    \Tile_X8Y9_WW4BEG[13] ,
    \Tile_X8Y9_WW4BEG[12] ,
    \Tile_X8Y9_WW4BEG[11] ,
    \Tile_X8Y9_WW4BEG[10] ,
    \Tile_X8Y9_WW4BEG[9] ,
    \Tile_X8Y9_WW4BEG[8] ,
    \Tile_X8Y9_WW4BEG[7] ,
    \Tile_X8Y9_WW4BEG[6] ,
    \Tile_X8Y9_WW4BEG[5] ,
    \Tile_X8Y9_WW4BEG[4] ,
    \Tile_X8Y9_WW4BEG[3] ,
    \Tile_X8Y9_WW4BEG[2] ,
    \Tile_X8Y9_WW4BEG[1] ,
    \Tile_X8Y9_WW4BEG[0] }),
    .WW4END({\Tile_X9Y9_WW4BEG[15] ,
    \Tile_X9Y9_WW4BEG[14] ,
    \Tile_X9Y9_WW4BEG[13] ,
    \Tile_X9Y9_WW4BEG[12] ,
    \Tile_X9Y9_WW4BEG[11] ,
    \Tile_X9Y9_WW4BEG[10] ,
    \Tile_X9Y9_WW4BEG[9] ,
    \Tile_X9Y9_WW4BEG[8] ,
    \Tile_X9Y9_WW4BEG[7] ,
    \Tile_X9Y9_WW4BEG[6] ,
    \Tile_X9Y9_WW4BEG[5] ,
    \Tile_X9Y9_WW4BEG[4] ,
    \Tile_X9Y9_WW4BEG[3] ,
    \Tile_X9Y9_WW4BEG[2] ,
    \Tile_X9Y9_WW4BEG[1] ,
    \Tile_X9Y9_WW4BEG[0] }));
 N_term_single Tile_X9Y0_N_term_single (.Ci(Tile_X9Y1_Co),
    .UserCLK(Tile_X9Y1_UserCLKo),
    .UserCLKo(Tile_X9Y0_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .FrameData({\Tile_X8Y0_FrameData_O[31] ,
    \Tile_X8Y0_FrameData_O[30] ,
    \Tile_X8Y0_FrameData_O[29] ,
    \Tile_X8Y0_FrameData_O[28] ,
    \Tile_X8Y0_FrameData_O[27] ,
    \Tile_X8Y0_FrameData_O[26] ,
    \Tile_X8Y0_FrameData_O[25] ,
    \Tile_X8Y0_FrameData_O[24] ,
    \Tile_X8Y0_FrameData_O[23] ,
    \Tile_X8Y0_FrameData_O[22] ,
    \Tile_X8Y0_FrameData_O[21] ,
    \Tile_X8Y0_FrameData_O[20] ,
    \Tile_X8Y0_FrameData_O[19] ,
    \Tile_X8Y0_FrameData_O[18] ,
    \Tile_X8Y0_FrameData_O[17] ,
    \Tile_X8Y0_FrameData_O[16] ,
    \Tile_X8Y0_FrameData_O[15] ,
    \Tile_X8Y0_FrameData_O[14] ,
    \Tile_X8Y0_FrameData_O[13] ,
    \Tile_X8Y0_FrameData_O[12] ,
    \Tile_X8Y0_FrameData_O[11] ,
    \Tile_X8Y0_FrameData_O[10] ,
    \Tile_X8Y0_FrameData_O[9] ,
    \Tile_X8Y0_FrameData_O[8] ,
    \Tile_X8Y0_FrameData_O[7] ,
    \Tile_X8Y0_FrameData_O[6] ,
    \Tile_X8Y0_FrameData_O[5] ,
    \Tile_X8Y0_FrameData_O[4] ,
    \Tile_X8Y0_FrameData_O[3] ,
    \Tile_X8Y0_FrameData_O[2] ,
    \Tile_X8Y0_FrameData_O[1] ,
    \Tile_X8Y0_FrameData_O[0] }),
    .FrameData_O({\Tile_X9Y0_FrameData_O[31] ,
    \Tile_X9Y0_FrameData_O[30] ,
    \Tile_X9Y0_FrameData_O[29] ,
    \Tile_X9Y0_FrameData_O[28] ,
    \Tile_X9Y0_FrameData_O[27] ,
    \Tile_X9Y0_FrameData_O[26] ,
    \Tile_X9Y0_FrameData_O[25] ,
    \Tile_X9Y0_FrameData_O[24] ,
    \Tile_X9Y0_FrameData_O[23] ,
    \Tile_X9Y0_FrameData_O[22] ,
    \Tile_X9Y0_FrameData_O[21] ,
    \Tile_X9Y0_FrameData_O[20] ,
    \Tile_X9Y0_FrameData_O[19] ,
    \Tile_X9Y0_FrameData_O[18] ,
    \Tile_X9Y0_FrameData_O[17] ,
    \Tile_X9Y0_FrameData_O[16] ,
    \Tile_X9Y0_FrameData_O[15] ,
    \Tile_X9Y0_FrameData_O[14] ,
    \Tile_X9Y0_FrameData_O[13] ,
    \Tile_X9Y0_FrameData_O[12] ,
    \Tile_X9Y0_FrameData_O[11] ,
    \Tile_X9Y0_FrameData_O[10] ,
    \Tile_X9Y0_FrameData_O[9] ,
    \Tile_X9Y0_FrameData_O[8] ,
    \Tile_X9Y0_FrameData_O[7] ,
    \Tile_X9Y0_FrameData_O[6] ,
    \Tile_X9Y0_FrameData_O[5] ,
    \Tile_X9Y0_FrameData_O[4] ,
    \Tile_X9Y0_FrameData_O[3] ,
    \Tile_X9Y0_FrameData_O[2] ,
    \Tile_X9Y0_FrameData_O[1] ,
    \Tile_X9Y0_FrameData_O[0] }),
    .FrameStrobe({\Tile_X9Y1_FrameStrobe_O[19] ,
    \Tile_X9Y1_FrameStrobe_O[18] ,
    \Tile_X9Y1_FrameStrobe_O[17] ,
    \Tile_X9Y1_FrameStrobe_O[16] ,
    \Tile_X9Y1_FrameStrobe_O[15] ,
    \Tile_X9Y1_FrameStrobe_O[14] ,
    \Tile_X9Y1_FrameStrobe_O[13] ,
    \Tile_X9Y1_FrameStrobe_O[12] ,
    \Tile_X9Y1_FrameStrobe_O[11] ,
    \Tile_X9Y1_FrameStrobe_O[10] ,
    \Tile_X9Y1_FrameStrobe_O[9] ,
    \Tile_X9Y1_FrameStrobe_O[8] ,
    \Tile_X9Y1_FrameStrobe_O[7] ,
    \Tile_X9Y1_FrameStrobe_O[6] ,
    \Tile_X9Y1_FrameStrobe_O[5] ,
    \Tile_X9Y1_FrameStrobe_O[4] ,
    \Tile_X9Y1_FrameStrobe_O[3] ,
    \Tile_X9Y1_FrameStrobe_O[2] ,
    \Tile_X9Y1_FrameStrobe_O[1] ,
    \Tile_X9Y1_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X9Y0_FrameStrobe_O[19] ,
    \Tile_X9Y0_FrameStrobe_O[18] ,
    \Tile_X9Y0_FrameStrobe_O[17] ,
    \Tile_X9Y0_FrameStrobe_O[16] ,
    \Tile_X9Y0_FrameStrobe_O[15] ,
    \Tile_X9Y0_FrameStrobe_O[14] ,
    \Tile_X9Y0_FrameStrobe_O[13] ,
    \Tile_X9Y0_FrameStrobe_O[12] ,
    \Tile_X9Y0_FrameStrobe_O[11] ,
    \Tile_X9Y0_FrameStrobe_O[10] ,
    \Tile_X9Y0_FrameStrobe_O[9] ,
    \Tile_X9Y0_FrameStrobe_O[8] ,
    \Tile_X9Y0_FrameStrobe_O[7] ,
    \Tile_X9Y0_FrameStrobe_O[6] ,
    \Tile_X9Y0_FrameStrobe_O[5] ,
    \Tile_X9Y0_FrameStrobe_O[4] ,
    \Tile_X9Y0_FrameStrobe_O[3] ,
    \Tile_X9Y0_FrameStrobe_O[2] ,
    \Tile_X9Y0_FrameStrobe_O[1] ,
    \Tile_X9Y0_FrameStrobe_O[0] }),
    .N1END({\Tile_X9Y1_N1BEG[3] ,
    \Tile_X9Y1_N1BEG[2] ,
    \Tile_X9Y1_N1BEG[1] ,
    \Tile_X9Y1_N1BEG[0] }),
    .N2END({\Tile_X9Y1_N2BEGb[7] ,
    \Tile_X9Y1_N2BEGb[6] ,
    \Tile_X9Y1_N2BEGb[5] ,
    \Tile_X9Y1_N2BEGb[4] ,
    \Tile_X9Y1_N2BEGb[3] ,
    \Tile_X9Y1_N2BEGb[2] ,
    \Tile_X9Y1_N2BEGb[1] ,
    \Tile_X9Y1_N2BEGb[0] }),
    .N2MID({\Tile_X9Y1_N2BEG[7] ,
    \Tile_X9Y1_N2BEG[6] ,
    \Tile_X9Y1_N2BEG[5] ,
    \Tile_X9Y1_N2BEG[4] ,
    \Tile_X9Y1_N2BEG[3] ,
    \Tile_X9Y1_N2BEG[2] ,
    \Tile_X9Y1_N2BEG[1] ,
    \Tile_X9Y1_N2BEG[0] }),
    .N4END({\Tile_X9Y1_N4BEG[15] ,
    \Tile_X9Y1_N4BEG[14] ,
    \Tile_X9Y1_N4BEG[13] ,
    \Tile_X9Y1_N4BEG[12] ,
    \Tile_X9Y1_N4BEG[11] ,
    \Tile_X9Y1_N4BEG[10] ,
    \Tile_X9Y1_N4BEG[9] ,
    \Tile_X9Y1_N4BEG[8] ,
    \Tile_X9Y1_N4BEG[7] ,
    \Tile_X9Y1_N4BEG[6] ,
    \Tile_X9Y1_N4BEG[5] ,
    \Tile_X9Y1_N4BEG[4] ,
    \Tile_X9Y1_N4BEG[3] ,
    \Tile_X9Y1_N4BEG[2] ,
    \Tile_X9Y1_N4BEG[1] ,
    \Tile_X9Y1_N4BEG[0] }),
    .NN4END({\Tile_X9Y1_NN4BEG[15] ,
    \Tile_X9Y1_NN4BEG[14] ,
    \Tile_X9Y1_NN4BEG[13] ,
    \Tile_X9Y1_NN4BEG[12] ,
    \Tile_X9Y1_NN4BEG[11] ,
    \Tile_X9Y1_NN4BEG[10] ,
    \Tile_X9Y1_NN4BEG[9] ,
    \Tile_X9Y1_NN4BEG[8] ,
    \Tile_X9Y1_NN4BEG[7] ,
    \Tile_X9Y1_NN4BEG[6] ,
    \Tile_X9Y1_NN4BEG[5] ,
    \Tile_X9Y1_NN4BEG[4] ,
    \Tile_X9Y1_NN4BEG[3] ,
    \Tile_X9Y1_NN4BEG[2] ,
    \Tile_X9Y1_NN4BEG[1] ,
    \Tile_X9Y1_NN4BEG[0] }),
    .S1BEG({\Tile_X9Y0_S1BEG[3] ,
    \Tile_X9Y0_S1BEG[2] ,
    \Tile_X9Y0_S1BEG[1] ,
    \Tile_X9Y0_S1BEG[0] }),
    .S2BEG({\Tile_X9Y0_S2BEG[7] ,
    \Tile_X9Y0_S2BEG[6] ,
    \Tile_X9Y0_S2BEG[5] ,
    \Tile_X9Y0_S2BEG[4] ,
    \Tile_X9Y0_S2BEG[3] ,
    \Tile_X9Y0_S2BEG[2] ,
    \Tile_X9Y0_S2BEG[1] ,
    \Tile_X9Y0_S2BEG[0] }),
    .S2BEGb({\Tile_X9Y0_S2BEGb[7] ,
    \Tile_X9Y0_S2BEGb[6] ,
    \Tile_X9Y0_S2BEGb[5] ,
    \Tile_X9Y0_S2BEGb[4] ,
    \Tile_X9Y0_S2BEGb[3] ,
    \Tile_X9Y0_S2BEGb[2] ,
    \Tile_X9Y0_S2BEGb[1] ,
    \Tile_X9Y0_S2BEGb[0] }),
    .S4BEG({\Tile_X9Y0_S4BEG[15] ,
    \Tile_X9Y0_S4BEG[14] ,
    \Tile_X9Y0_S4BEG[13] ,
    \Tile_X9Y0_S4BEG[12] ,
    \Tile_X9Y0_S4BEG[11] ,
    \Tile_X9Y0_S4BEG[10] ,
    \Tile_X9Y0_S4BEG[9] ,
    \Tile_X9Y0_S4BEG[8] ,
    \Tile_X9Y0_S4BEG[7] ,
    \Tile_X9Y0_S4BEG[6] ,
    \Tile_X9Y0_S4BEG[5] ,
    \Tile_X9Y0_S4BEG[4] ,
    \Tile_X9Y0_S4BEG[3] ,
    \Tile_X9Y0_S4BEG[2] ,
    \Tile_X9Y0_S4BEG[1] ,
    \Tile_X9Y0_S4BEG[0] }),
    .SS4BEG({\Tile_X9Y0_SS4BEG[15] ,
    \Tile_X9Y0_SS4BEG[14] ,
    \Tile_X9Y0_SS4BEG[13] ,
    \Tile_X9Y0_SS4BEG[12] ,
    \Tile_X9Y0_SS4BEG[11] ,
    \Tile_X9Y0_SS4BEG[10] ,
    \Tile_X9Y0_SS4BEG[9] ,
    \Tile_X9Y0_SS4BEG[8] ,
    \Tile_X9Y0_SS4BEG[7] ,
    \Tile_X9Y0_SS4BEG[6] ,
    \Tile_X9Y0_SS4BEG[5] ,
    \Tile_X9Y0_SS4BEG[4] ,
    \Tile_X9Y0_SS4BEG[3] ,
    \Tile_X9Y0_SS4BEG[2] ,
    \Tile_X9Y0_SS4BEG[1] ,
    \Tile_X9Y0_SS4BEG[0] }));
 LUT4AB Tile_X9Y10_LUT4AB (.Ci(Tile_X9Y11_Co),
    .Co(Tile_X9Y10_Co),
    .UserCLK(Tile_X9Y11_UserCLKo),
    .UserCLKo(Tile_X9Y10_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X9Y10_E1BEG[3] ,
    \Tile_X9Y10_E1BEG[2] ,
    \Tile_X9Y10_E1BEG[1] ,
    \Tile_X9Y10_E1BEG[0] }),
    .E1END({\Tile_X8Y10_E1BEG[3] ,
    \Tile_X8Y10_E1BEG[2] ,
    \Tile_X8Y10_E1BEG[1] ,
    \Tile_X8Y10_E1BEG[0] }),
    .E2BEG({\Tile_X9Y10_E2BEG[7] ,
    \Tile_X9Y10_E2BEG[6] ,
    \Tile_X9Y10_E2BEG[5] ,
    \Tile_X9Y10_E2BEG[4] ,
    \Tile_X9Y10_E2BEG[3] ,
    \Tile_X9Y10_E2BEG[2] ,
    \Tile_X9Y10_E2BEG[1] ,
    \Tile_X9Y10_E2BEG[0] }),
    .E2BEGb({\Tile_X9Y10_E2BEGb[7] ,
    \Tile_X9Y10_E2BEGb[6] ,
    \Tile_X9Y10_E2BEGb[5] ,
    \Tile_X9Y10_E2BEGb[4] ,
    \Tile_X9Y10_E2BEGb[3] ,
    \Tile_X9Y10_E2BEGb[2] ,
    \Tile_X9Y10_E2BEGb[1] ,
    \Tile_X9Y10_E2BEGb[0] }),
    .E2END({\Tile_X8Y10_E2BEGb[7] ,
    \Tile_X8Y10_E2BEGb[6] ,
    \Tile_X8Y10_E2BEGb[5] ,
    \Tile_X8Y10_E2BEGb[4] ,
    \Tile_X8Y10_E2BEGb[3] ,
    \Tile_X8Y10_E2BEGb[2] ,
    \Tile_X8Y10_E2BEGb[1] ,
    \Tile_X8Y10_E2BEGb[0] }),
    .E2MID({\Tile_X8Y10_E2BEG[7] ,
    \Tile_X8Y10_E2BEG[6] ,
    \Tile_X8Y10_E2BEG[5] ,
    \Tile_X8Y10_E2BEG[4] ,
    \Tile_X8Y10_E2BEG[3] ,
    \Tile_X8Y10_E2BEG[2] ,
    \Tile_X8Y10_E2BEG[1] ,
    \Tile_X8Y10_E2BEG[0] }),
    .E6BEG({\Tile_X9Y10_E6BEG[11] ,
    \Tile_X9Y10_E6BEG[10] ,
    \Tile_X9Y10_E6BEG[9] ,
    \Tile_X9Y10_E6BEG[8] ,
    \Tile_X9Y10_E6BEG[7] ,
    \Tile_X9Y10_E6BEG[6] ,
    \Tile_X9Y10_E6BEG[5] ,
    \Tile_X9Y10_E6BEG[4] ,
    \Tile_X9Y10_E6BEG[3] ,
    \Tile_X9Y10_E6BEG[2] ,
    \Tile_X9Y10_E6BEG[1] ,
    \Tile_X9Y10_E6BEG[0] }),
    .E6END({\Tile_X8Y10_E6BEG[11] ,
    \Tile_X8Y10_E6BEG[10] ,
    \Tile_X8Y10_E6BEG[9] ,
    \Tile_X8Y10_E6BEG[8] ,
    \Tile_X8Y10_E6BEG[7] ,
    \Tile_X8Y10_E6BEG[6] ,
    \Tile_X8Y10_E6BEG[5] ,
    \Tile_X8Y10_E6BEG[4] ,
    \Tile_X8Y10_E6BEG[3] ,
    \Tile_X8Y10_E6BEG[2] ,
    \Tile_X8Y10_E6BEG[1] ,
    \Tile_X8Y10_E6BEG[0] }),
    .EE4BEG({\Tile_X9Y10_EE4BEG[15] ,
    \Tile_X9Y10_EE4BEG[14] ,
    \Tile_X9Y10_EE4BEG[13] ,
    \Tile_X9Y10_EE4BEG[12] ,
    \Tile_X9Y10_EE4BEG[11] ,
    \Tile_X9Y10_EE4BEG[10] ,
    \Tile_X9Y10_EE4BEG[9] ,
    \Tile_X9Y10_EE4BEG[8] ,
    \Tile_X9Y10_EE4BEG[7] ,
    \Tile_X9Y10_EE4BEG[6] ,
    \Tile_X9Y10_EE4BEG[5] ,
    \Tile_X9Y10_EE4BEG[4] ,
    \Tile_X9Y10_EE4BEG[3] ,
    \Tile_X9Y10_EE4BEG[2] ,
    \Tile_X9Y10_EE4BEG[1] ,
    \Tile_X9Y10_EE4BEG[0] }),
    .EE4END({\Tile_X8Y10_EE4BEG[15] ,
    \Tile_X8Y10_EE4BEG[14] ,
    \Tile_X8Y10_EE4BEG[13] ,
    \Tile_X8Y10_EE4BEG[12] ,
    \Tile_X8Y10_EE4BEG[11] ,
    \Tile_X8Y10_EE4BEG[10] ,
    \Tile_X8Y10_EE4BEG[9] ,
    \Tile_X8Y10_EE4BEG[8] ,
    \Tile_X8Y10_EE4BEG[7] ,
    \Tile_X8Y10_EE4BEG[6] ,
    \Tile_X8Y10_EE4BEG[5] ,
    \Tile_X8Y10_EE4BEG[4] ,
    \Tile_X8Y10_EE4BEG[3] ,
    \Tile_X8Y10_EE4BEG[2] ,
    \Tile_X8Y10_EE4BEG[1] ,
    \Tile_X8Y10_EE4BEG[0] }),
    .FrameData({\Tile_X8Y10_FrameData_O[31] ,
    \Tile_X8Y10_FrameData_O[30] ,
    \Tile_X8Y10_FrameData_O[29] ,
    \Tile_X8Y10_FrameData_O[28] ,
    \Tile_X8Y10_FrameData_O[27] ,
    \Tile_X8Y10_FrameData_O[26] ,
    \Tile_X8Y10_FrameData_O[25] ,
    \Tile_X8Y10_FrameData_O[24] ,
    \Tile_X8Y10_FrameData_O[23] ,
    \Tile_X8Y10_FrameData_O[22] ,
    \Tile_X8Y10_FrameData_O[21] ,
    \Tile_X8Y10_FrameData_O[20] ,
    \Tile_X8Y10_FrameData_O[19] ,
    \Tile_X8Y10_FrameData_O[18] ,
    \Tile_X8Y10_FrameData_O[17] ,
    \Tile_X8Y10_FrameData_O[16] ,
    \Tile_X8Y10_FrameData_O[15] ,
    \Tile_X8Y10_FrameData_O[14] ,
    \Tile_X8Y10_FrameData_O[13] ,
    \Tile_X8Y10_FrameData_O[12] ,
    \Tile_X8Y10_FrameData_O[11] ,
    \Tile_X8Y10_FrameData_O[10] ,
    \Tile_X8Y10_FrameData_O[9] ,
    \Tile_X8Y10_FrameData_O[8] ,
    \Tile_X8Y10_FrameData_O[7] ,
    \Tile_X8Y10_FrameData_O[6] ,
    \Tile_X8Y10_FrameData_O[5] ,
    \Tile_X8Y10_FrameData_O[4] ,
    \Tile_X8Y10_FrameData_O[3] ,
    \Tile_X8Y10_FrameData_O[2] ,
    \Tile_X8Y10_FrameData_O[1] ,
    \Tile_X8Y10_FrameData_O[0] }),
    .FrameData_O({\Tile_X9Y10_FrameData_O[31] ,
    \Tile_X9Y10_FrameData_O[30] ,
    \Tile_X9Y10_FrameData_O[29] ,
    \Tile_X9Y10_FrameData_O[28] ,
    \Tile_X9Y10_FrameData_O[27] ,
    \Tile_X9Y10_FrameData_O[26] ,
    \Tile_X9Y10_FrameData_O[25] ,
    \Tile_X9Y10_FrameData_O[24] ,
    \Tile_X9Y10_FrameData_O[23] ,
    \Tile_X9Y10_FrameData_O[22] ,
    \Tile_X9Y10_FrameData_O[21] ,
    \Tile_X9Y10_FrameData_O[20] ,
    \Tile_X9Y10_FrameData_O[19] ,
    \Tile_X9Y10_FrameData_O[18] ,
    \Tile_X9Y10_FrameData_O[17] ,
    \Tile_X9Y10_FrameData_O[16] ,
    \Tile_X9Y10_FrameData_O[15] ,
    \Tile_X9Y10_FrameData_O[14] ,
    \Tile_X9Y10_FrameData_O[13] ,
    \Tile_X9Y10_FrameData_O[12] ,
    \Tile_X9Y10_FrameData_O[11] ,
    \Tile_X9Y10_FrameData_O[10] ,
    \Tile_X9Y10_FrameData_O[9] ,
    \Tile_X9Y10_FrameData_O[8] ,
    \Tile_X9Y10_FrameData_O[7] ,
    \Tile_X9Y10_FrameData_O[6] ,
    \Tile_X9Y10_FrameData_O[5] ,
    \Tile_X9Y10_FrameData_O[4] ,
    \Tile_X9Y10_FrameData_O[3] ,
    \Tile_X9Y10_FrameData_O[2] ,
    \Tile_X9Y10_FrameData_O[1] ,
    \Tile_X9Y10_FrameData_O[0] }),
    .FrameStrobe({\Tile_X9Y11_FrameStrobe_O[19] ,
    \Tile_X9Y11_FrameStrobe_O[18] ,
    \Tile_X9Y11_FrameStrobe_O[17] ,
    \Tile_X9Y11_FrameStrobe_O[16] ,
    \Tile_X9Y11_FrameStrobe_O[15] ,
    \Tile_X9Y11_FrameStrobe_O[14] ,
    \Tile_X9Y11_FrameStrobe_O[13] ,
    \Tile_X9Y11_FrameStrobe_O[12] ,
    \Tile_X9Y11_FrameStrobe_O[11] ,
    \Tile_X9Y11_FrameStrobe_O[10] ,
    \Tile_X9Y11_FrameStrobe_O[9] ,
    \Tile_X9Y11_FrameStrobe_O[8] ,
    \Tile_X9Y11_FrameStrobe_O[7] ,
    \Tile_X9Y11_FrameStrobe_O[6] ,
    \Tile_X9Y11_FrameStrobe_O[5] ,
    \Tile_X9Y11_FrameStrobe_O[4] ,
    \Tile_X9Y11_FrameStrobe_O[3] ,
    \Tile_X9Y11_FrameStrobe_O[2] ,
    \Tile_X9Y11_FrameStrobe_O[1] ,
    \Tile_X9Y11_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X9Y10_FrameStrobe_O[19] ,
    \Tile_X9Y10_FrameStrobe_O[18] ,
    \Tile_X9Y10_FrameStrobe_O[17] ,
    \Tile_X9Y10_FrameStrobe_O[16] ,
    \Tile_X9Y10_FrameStrobe_O[15] ,
    \Tile_X9Y10_FrameStrobe_O[14] ,
    \Tile_X9Y10_FrameStrobe_O[13] ,
    \Tile_X9Y10_FrameStrobe_O[12] ,
    \Tile_X9Y10_FrameStrobe_O[11] ,
    \Tile_X9Y10_FrameStrobe_O[10] ,
    \Tile_X9Y10_FrameStrobe_O[9] ,
    \Tile_X9Y10_FrameStrobe_O[8] ,
    \Tile_X9Y10_FrameStrobe_O[7] ,
    \Tile_X9Y10_FrameStrobe_O[6] ,
    \Tile_X9Y10_FrameStrobe_O[5] ,
    \Tile_X9Y10_FrameStrobe_O[4] ,
    \Tile_X9Y10_FrameStrobe_O[3] ,
    \Tile_X9Y10_FrameStrobe_O[2] ,
    \Tile_X9Y10_FrameStrobe_O[1] ,
    \Tile_X9Y10_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X9Y10_N1BEG[3] ,
    \Tile_X9Y10_N1BEG[2] ,
    \Tile_X9Y10_N1BEG[1] ,
    \Tile_X9Y10_N1BEG[0] }),
    .N1END({\Tile_X9Y11_N1BEG[3] ,
    \Tile_X9Y11_N1BEG[2] ,
    \Tile_X9Y11_N1BEG[1] ,
    \Tile_X9Y11_N1BEG[0] }),
    .N2BEG({\Tile_X9Y10_N2BEG[7] ,
    \Tile_X9Y10_N2BEG[6] ,
    \Tile_X9Y10_N2BEG[5] ,
    \Tile_X9Y10_N2BEG[4] ,
    \Tile_X9Y10_N2BEG[3] ,
    \Tile_X9Y10_N2BEG[2] ,
    \Tile_X9Y10_N2BEG[1] ,
    \Tile_X9Y10_N2BEG[0] }),
    .N2BEGb({\Tile_X9Y10_N2BEGb[7] ,
    \Tile_X9Y10_N2BEGb[6] ,
    \Tile_X9Y10_N2BEGb[5] ,
    \Tile_X9Y10_N2BEGb[4] ,
    \Tile_X9Y10_N2BEGb[3] ,
    \Tile_X9Y10_N2BEGb[2] ,
    \Tile_X9Y10_N2BEGb[1] ,
    \Tile_X9Y10_N2BEGb[0] }),
    .N2END({\Tile_X9Y11_N2BEGb[7] ,
    \Tile_X9Y11_N2BEGb[6] ,
    \Tile_X9Y11_N2BEGb[5] ,
    \Tile_X9Y11_N2BEGb[4] ,
    \Tile_X9Y11_N2BEGb[3] ,
    \Tile_X9Y11_N2BEGb[2] ,
    \Tile_X9Y11_N2BEGb[1] ,
    \Tile_X9Y11_N2BEGb[0] }),
    .N2MID({\Tile_X9Y11_N2BEG[7] ,
    \Tile_X9Y11_N2BEG[6] ,
    \Tile_X9Y11_N2BEG[5] ,
    \Tile_X9Y11_N2BEG[4] ,
    \Tile_X9Y11_N2BEG[3] ,
    \Tile_X9Y11_N2BEG[2] ,
    \Tile_X9Y11_N2BEG[1] ,
    \Tile_X9Y11_N2BEG[0] }),
    .N4BEG({\Tile_X9Y10_N4BEG[15] ,
    \Tile_X9Y10_N4BEG[14] ,
    \Tile_X9Y10_N4BEG[13] ,
    \Tile_X9Y10_N4BEG[12] ,
    \Tile_X9Y10_N4BEG[11] ,
    \Tile_X9Y10_N4BEG[10] ,
    \Tile_X9Y10_N4BEG[9] ,
    \Tile_X9Y10_N4BEG[8] ,
    \Tile_X9Y10_N4BEG[7] ,
    \Tile_X9Y10_N4BEG[6] ,
    \Tile_X9Y10_N4BEG[5] ,
    \Tile_X9Y10_N4BEG[4] ,
    \Tile_X9Y10_N4BEG[3] ,
    \Tile_X9Y10_N4BEG[2] ,
    \Tile_X9Y10_N4BEG[1] ,
    \Tile_X9Y10_N4BEG[0] }),
    .N4END({\Tile_X9Y11_N4BEG[15] ,
    \Tile_X9Y11_N4BEG[14] ,
    \Tile_X9Y11_N4BEG[13] ,
    \Tile_X9Y11_N4BEG[12] ,
    \Tile_X9Y11_N4BEG[11] ,
    \Tile_X9Y11_N4BEG[10] ,
    \Tile_X9Y11_N4BEG[9] ,
    \Tile_X9Y11_N4BEG[8] ,
    \Tile_X9Y11_N4BEG[7] ,
    \Tile_X9Y11_N4BEG[6] ,
    \Tile_X9Y11_N4BEG[5] ,
    \Tile_X9Y11_N4BEG[4] ,
    \Tile_X9Y11_N4BEG[3] ,
    \Tile_X9Y11_N4BEG[2] ,
    \Tile_X9Y11_N4BEG[1] ,
    \Tile_X9Y11_N4BEG[0] }),
    .NN4BEG({\Tile_X9Y10_NN4BEG[15] ,
    \Tile_X9Y10_NN4BEG[14] ,
    \Tile_X9Y10_NN4BEG[13] ,
    \Tile_X9Y10_NN4BEG[12] ,
    \Tile_X9Y10_NN4BEG[11] ,
    \Tile_X9Y10_NN4BEG[10] ,
    \Tile_X9Y10_NN4BEG[9] ,
    \Tile_X9Y10_NN4BEG[8] ,
    \Tile_X9Y10_NN4BEG[7] ,
    \Tile_X9Y10_NN4BEG[6] ,
    \Tile_X9Y10_NN4BEG[5] ,
    \Tile_X9Y10_NN4BEG[4] ,
    \Tile_X9Y10_NN4BEG[3] ,
    \Tile_X9Y10_NN4BEG[2] ,
    \Tile_X9Y10_NN4BEG[1] ,
    \Tile_X9Y10_NN4BEG[0] }),
    .NN4END({\Tile_X9Y11_NN4BEG[15] ,
    \Tile_X9Y11_NN4BEG[14] ,
    \Tile_X9Y11_NN4BEG[13] ,
    \Tile_X9Y11_NN4BEG[12] ,
    \Tile_X9Y11_NN4BEG[11] ,
    \Tile_X9Y11_NN4BEG[10] ,
    \Tile_X9Y11_NN4BEG[9] ,
    \Tile_X9Y11_NN4BEG[8] ,
    \Tile_X9Y11_NN4BEG[7] ,
    \Tile_X9Y11_NN4BEG[6] ,
    \Tile_X9Y11_NN4BEG[5] ,
    \Tile_X9Y11_NN4BEG[4] ,
    \Tile_X9Y11_NN4BEG[3] ,
    \Tile_X9Y11_NN4BEG[2] ,
    \Tile_X9Y11_NN4BEG[1] ,
    \Tile_X9Y11_NN4BEG[0] }),
    .S1BEG({\Tile_X9Y10_S1BEG[3] ,
    \Tile_X9Y10_S1BEG[2] ,
    \Tile_X9Y10_S1BEG[1] ,
    \Tile_X9Y10_S1BEG[0] }),
    .S1END({\Tile_X9Y9_S1BEG[3] ,
    \Tile_X9Y9_S1BEG[2] ,
    \Tile_X9Y9_S1BEG[1] ,
    \Tile_X9Y9_S1BEG[0] }),
    .S2BEG({\Tile_X9Y10_S2BEG[7] ,
    \Tile_X9Y10_S2BEG[6] ,
    \Tile_X9Y10_S2BEG[5] ,
    \Tile_X9Y10_S2BEG[4] ,
    \Tile_X9Y10_S2BEG[3] ,
    \Tile_X9Y10_S2BEG[2] ,
    \Tile_X9Y10_S2BEG[1] ,
    \Tile_X9Y10_S2BEG[0] }),
    .S2BEGb({\Tile_X9Y10_S2BEGb[7] ,
    \Tile_X9Y10_S2BEGb[6] ,
    \Tile_X9Y10_S2BEGb[5] ,
    \Tile_X9Y10_S2BEGb[4] ,
    \Tile_X9Y10_S2BEGb[3] ,
    \Tile_X9Y10_S2BEGb[2] ,
    \Tile_X9Y10_S2BEGb[1] ,
    \Tile_X9Y10_S2BEGb[0] }),
    .S2END({\Tile_X9Y9_S2BEGb[7] ,
    \Tile_X9Y9_S2BEGb[6] ,
    \Tile_X9Y9_S2BEGb[5] ,
    \Tile_X9Y9_S2BEGb[4] ,
    \Tile_X9Y9_S2BEGb[3] ,
    \Tile_X9Y9_S2BEGb[2] ,
    \Tile_X9Y9_S2BEGb[1] ,
    \Tile_X9Y9_S2BEGb[0] }),
    .S2MID({\Tile_X9Y9_S2BEG[7] ,
    \Tile_X9Y9_S2BEG[6] ,
    \Tile_X9Y9_S2BEG[5] ,
    \Tile_X9Y9_S2BEG[4] ,
    \Tile_X9Y9_S2BEG[3] ,
    \Tile_X9Y9_S2BEG[2] ,
    \Tile_X9Y9_S2BEG[1] ,
    \Tile_X9Y9_S2BEG[0] }),
    .S4BEG({\Tile_X9Y10_S4BEG[15] ,
    \Tile_X9Y10_S4BEG[14] ,
    \Tile_X9Y10_S4BEG[13] ,
    \Tile_X9Y10_S4BEG[12] ,
    \Tile_X9Y10_S4BEG[11] ,
    \Tile_X9Y10_S4BEG[10] ,
    \Tile_X9Y10_S4BEG[9] ,
    \Tile_X9Y10_S4BEG[8] ,
    \Tile_X9Y10_S4BEG[7] ,
    \Tile_X9Y10_S4BEG[6] ,
    \Tile_X9Y10_S4BEG[5] ,
    \Tile_X9Y10_S4BEG[4] ,
    \Tile_X9Y10_S4BEG[3] ,
    \Tile_X9Y10_S4BEG[2] ,
    \Tile_X9Y10_S4BEG[1] ,
    \Tile_X9Y10_S4BEG[0] }),
    .S4END({\Tile_X9Y9_S4BEG[15] ,
    \Tile_X9Y9_S4BEG[14] ,
    \Tile_X9Y9_S4BEG[13] ,
    \Tile_X9Y9_S4BEG[12] ,
    \Tile_X9Y9_S4BEG[11] ,
    \Tile_X9Y9_S4BEG[10] ,
    \Tile_X9Y9_S4BEG[9] ,
    \Tile_X9Y9_S4BEG[8] ,
    \Tile_X9Y9_S4BEG[7] ,
    \Tile_X9Y9_S4BEG[6] ,
    \Tile_X9Y9_S4BEG[5] ,
    \Tile_X9Y9_S4BEG[4] ,
    \Tile_X9Y9_S4BEG[3] ,
    \Tile_X9Y9_S4BEG[2] ,
    \Tile_X9Y9_S4BEG[1] ,
    \Tile_X9Y9_S4BEG[0] }),
    .SS4BEG({\Tile_X9Y10_SS4BEG[15] ,
    \Tile_X9Y10_SS4BEG[14] ,
    \Tile_X9Y10_SS4BEG[13] ,
    \Tile_X9Y10_SS4BEG[12] ,
    \Tile_X9Y10_SS4BEG[11] ,
    \Tile_X9Y10_SS4BEG[10] ,
    \Tile_X9Y10_SS4BEG[9] ,
    \Tile_X9Y10_SS4BEG[8] ,
    \Tile_X9Y10_SS4BEG[7] ,
    \Tile_X9Y10_SS4BEG[6] ,
    \Tile_X9Y10_SS4BEG[5] ,
    \Tile_X9Y10_SS4BEG[4] ,
    \Tile_X9Y10_SS4BEG[3] ,
    \Tile_X9Y10_SS4BEG[2] ,
    \Tile_X9Y10_SS4BEG[1] ,
    \Tile_X9Y10_SS4BEG[0] }),
    .SS4END({\Tile_X9Y9_SS4BEG[15] ,
    \Tile_X9Y9_SS4BEG[14] ,
    \Tile_X9Y9_SS4BEG[13] ,
    \Tile_X9Y9_SS4BEG[12] ,
    \Tile_X9Y9_SS4BEG[11] ,
    \Tile_X9Y9_SS4BEG[10] ,
    \Tile_X9Y9_SS4BEG[9] ,
    \Tile_X9Y9_SS4BEG[8] ,
    \Tile_X9Y9_SS4BEG[7] ,
    \Tile_X9Y9_SS4BEG[6] ,
    \Tile_X9Y9_SS4BEG[5] ,
    \Tile_X9Y9_SS4BEG[4] ,
    \Tile_X9Y9_SS4BEG[3] ,
    \Tile_X9Y9_SS4BEG[2] ,
    \Tile_X9Y9_SS4BEG[1] ,
    \Tile_X9Y9_SS4BEG[0] }),
    .W1BEG({\Tile_X9Y10_W1BEG[3] ,
    \Tile_X9Y10_W1BEG[2] ,
    \Tile_X9Y10_W1BEG[1] ,
    \Tile_X9Y10_W1BEG[0] }),
    .W1END({\Tile_X10Y10_W1BEG[3] ,
    \Tile_X10Y10_W1BEG[2] ,
    \Tile_X10Y10_W1BEG[1] ,
    \Tile_X10Y10_W1BEG[0] }),
    .W2BEG({\Tile_X9Y10_W2BEG[7] ,
    \Tile_X9Y10_W2BEG[6] ,
    \Tile_X9Y10_W2BEG[5] ,
    \Tile_X9Y10_W2BEG[4] ,
    \Tile_X9Y10_W2BEG[3] ,
    \Tile_X9Y10_W2BEG[2] ,
    \Tile_X9Y10_W2BEG[1] ,
    \Tile_X9Y10_W2BEG[0] }),
    .W2BEGb({\Tile_X9Y10_W2BEGb[7] ,
    \Tile_X9Y10_W2BEGb[6] ,
    \Tile_X9Y10_W2BEGb[5] ,
    \Tile_X9Y10_W2BEGb[4] ,
    \Tile_X9Y10_W2BEGb[3] ,
    \Tile_X9Y10_W2BEGb[2] ,
    \Tile_X9Y10_W2BEGb[1] ,
    \Tile_X9Y10_W2BEGb[0] }),
    .W2END({\Tile_X10Y10_W2BEGb[7] ,
    \Tile_X10Y10_W2BEGb[6] ,
    \Tile_X10Y10_W2BEGb[5] ,
    \Tile_X10Y10_W2BEGb[4] ,
    \Tile_X10Y10_W2BEGb[3] ,
    \Tile_X10Y10_W2BEGb[2] ,
    \Tile_X10Y10_W2BEGb[1] ,
    \Tile_X10Y10_W2BEGb[0] }),
    .W2MID({\Tile_X10Y10_W2BEG[7] ,
    \Tile_X10Y10_W2BEG[6] ,
    \Tile_X10Y10_W2BEG[5] ,
    \Tile_X10Y10_W2BEG[4] ,
    \Tile_X10Y10_W2BEG[3] ,
    \Tile_X10Y10_W2BEG[2] ,
    \Tile_X10Y10_W2BEG[1] ,
    \Tile_X10Y10_W2BEG[0] }),
    .W6BEG({\Tile_X9Y10_W6BEG[11] ,
    \Tile_X9Y10_W6BEG[10] ,
    \Tile_X9Y10_W6BEG[9] ,
    \Tile_X9Y10_W6BEG[8] ,
    \Tile_X9Y10_W6BEG[7] ,
    \Tile_X9Y10_W6BEG[6] ,
    \Tile_X9Y10_W6BEG[5] ,
    \Tile_X9Y10_W6BEG[4] ,
    \Tile_X9Y10_W6BEG[3] ,
    \Tile_X9Y10_W6BEG[2] ,
    \Tile_X9Y10_W6BEG[1] ,
    \Tile_X9Y10_W6BEG[0] }),
    .W6END({\Tile_X10Y10_W6BEG[11] ,
    \Tile_X10Y10_W6BEG[10] ,
    \Tile_X10Y10_W6BEG[9] ,
    \Tile_X10Y10_W6BEG[8] ,
    \Tile_X10Y10_W6BEG[7] ,
    \Tile_X10Y10_W6BEG[6] ,
    \Tile_X10Y10_W6BEG[5] ,
    \Tile_X10Y10_W6BEG[4] ,
    \Tile_X10Y10_W6BEG[3] ,
    \Tile_X10Y10_W6BEG[2] ,
    \Tile_X10Y10_W6BEG[1] ,
    \Tile_X10Y10_W6BEG[0] }),
    .WW4BEG({\Tile_X9Y10_WW4BEG[15] ,
    \Tile_X9Y10_WW4BEG[14] ,
    \Tile_X9Y10_WW4BEG[13] ,
    \Tile_X9Y10_WW4BEG[12] ,
    \Tile_X9Y10_WW4BEG[11] ,
    \Tile_X9Y10_WW4BEG[10] ,
    \Tile_X9Y10_WW4BEG[9] ,
    \Tile_X9Y10_WW4BEG[8] ,
    \Tile_X9Y10_WW4BEG[7] ,
    \Tile_X9Y10_WW4BEG[6] ,
    \Tile_X9Y10_WW4BEG[5] ,
    \Tile_X9Y10_WW4BEG[4] ,
    \Tile_X9Y10_WW4BEG[3] ,
    \Tile_X9Y10_WW4BEG[2] ,
    \Tile_X9Y10_WW4BEG[1] ,
    \Tile_X9Y10_WW4BEG[0] }),
    .WW4END({\Tile_X10Y10_WW4BEG[15] ,
    \Tile_X10Y10_WW4BEG[14] ,
    \Tile_X10Y10_WW4BEG[13] ,
    \Tile_X10Y10_WW4BEG[12] ,
    \Tile_X10Y10_WW4BEG[11] ,
    \Tile_X10Y10_WW4BEG[10] ,
    \Tile_X10Y10_WW4BEG[9] ,
    \Tile_X10Y10_WW4BEG[8] ,
    \Tile_X10Y10_WW4BEG[7] ,
    \Tile_X10Y10_WW4BEG[6] ,
    \Tile_X10Y10_WW4BEG[5] ,
    \Tile_X10Y10_WW4BEG[4] ,
    \Tile_X10Y10_WW4BEG[3] ,
    \Tile_X10Y10_WW4BEG[2] ,
    \Tile_X10Y10_WW4BEG[1] ,
    \Tile_X10Y10_WW4BEG[0] }));
 LUT4AB Tile_X9Y11_LUT4AB (.Ci(Tile_X9Y12_Co),
    .Co(Tile_X9Y11_Co),
    .UserCLK(Tile_X9Y12_UserCLKo),
    .UserCLKo(Tile_X9Y11_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X9Y11_E1BEG[3] ,
    \Tile_X9Y11_E1BEG[2] ,
    \Tile_X9Y11_E1BEG[1] ,
    \Tile_X9Y11_E1BEG[0] }),
    .E1END({\Tile_X8Y11_E1BEG[3] ,
    \Tile_X8Y11_E1BEG[2] ,
    \Tile_X8Y11_E1BEG[1] ,
    \Tile_X8Y11_E1BEG[0] }),
    .E2BEG({\Tile_X9Y11_E2BEG[7] ,
    \Tile_X9Y11_E2BEG[6] ,
    \Tile_X9Y11_E2BEG[5] ,
    \Tile_X9Y11_E2BEG[4] ,
    \Tile_X9Y11_E2BEG[3] ,
    \Tile_X9Y11_E2BEG[2] ,
    \Tile_X9Y11_E2BEG[1] ,
    \Tile_X9Y11_E2BEG[0] }),
    .E2BEGb({\Tile_X9Y11_E2BEGb[7] ,
    \Tile_X9Y11_E2BEGb[6] ,
    \Tile_X9Y11_E2BEGb[5] ,
    \Tile_X9Y11_E2BEGb[4] ,
    \Tile_X9Y11_E2BEGb[3] ,
    \Tile_X9Y11_E2BEGb[2] ,
    \Tile_X9Y11_E2BEGb[1] ,
    \Tile_X9Y11_E2BEGb[0] }),
    .E2END({\Tile_X8Y11_E2BEGb[7] ,
    \Tile_X8Y11_E2BEGb[6] ,
    \Tile_X8Y11_E2BEGb[5] ,
    \Tile_X8Y11_E2BEGb[4] ,
    \Tile_X8Y11_E2BEGb[3] ,
    \Tile_X8Y11_E2BEGb[2] ,
    \Tile_X8Y11_E2BEGb[1] ,
    \Tile_X8Y11_E2BEGb[0] }),
    .E2MID({\Tile_X8Y11_E2BEG[7] ,
    \Tile_X8Y11_E2BEG[6] ,
    \Tile_X8Y11_E2BEG[5] ,
    \Tile_X8Y11_E2BEG[4] ,
    \Tile_X8Y11_E2BEG[3] ,
    \Tile_X8Y11_E2BEG[2] ,
    \Tile_X8Y11_E2BEG[1] ,
    \Tile_X8Y11_E2BEG[0] }),
    .E6BEG({\Tile_X9Y11_E6BEG[11] ,
    \Tile_X9Y11_E6BEG[10] ,
    \Tile_X9Y11_E6BEG[9] ,
    \Tile_X9Y11_E6BEG[8] ,
    \Tile_X9Y11_E6BEG[7] ,
    \Tile_X9Y11_E6BEG[6] ,
    \Tile_X9Y11_E6BEG[5] ,
    \Tile_X9Y11_E6BEG[4] ,
    \Tile_X9Y11_E6BEG[3] ,
    \Tile_X9Y11_E6BEG[2] ,
    \Tile_X9Y11_E6BEG[1] ,
    \Tile_X9Y11_E6BEG[0] }),
    .E6END({\Tile_X8Y11_E6BEG[11] ,
    \Tile_X8Y11_E6BEG[10] ,
    \Tile_X8Y11_E6BEG[9] ,
    \Tile_X8Y11_E6BEG[8] ,
    \Tile_X8Y11_E6BEG[7] ,
    \Tile_X8Y11_E6BEG[6] ,
    \Tile_X8Y11_E6BEG[5] ,
    \Tile_X8Y11_E6BEG[4] ,
    \Tile_X8Y11_E6BEG[3] ,
    \Tile_X8Y11_E6BEG[2] ,
    \Tile_X8Y11_E6BEG[1] ,
    \Tile_X8Y11_E6BEG[0] }),
    .EE4BEG({\Tile_X9Y11_EE4BEG[15] ,
    \Tile_X9Y11_EE4BEG[14] ,
    \Tile_X9Y11_EE4BEG[13] ,
    \Tile_X9Y11_EE4BEG[12] ,
    \Tile_X9Y11_EE4BEG[11] ,
    \Tile_X9Y11_EE4BEG[10] ,
    \Tile_X9Y11_EE4BEG[9] ,
    \Tile_X9Y11_EE4BEG[8] ,
    \Tile_X9Y11_EE4BEG[7] ,
    \Tile_X9Y11_EE4BEG[6] ,
    \Tile_X9Y11_EE4BEG[5] ,
    \Tile_X9Y11_EE4BEG[4] ,
    \Tile_X9Y11_EE4BEG[3] ,
    \Tile_X9Y11_EE4BEG[2] ,
    \Tile_X9Y11_EE4BEG[1] ,
    \Tile_X9Y11_EE4BEG[0] }),
    .EE4END({\Tile_X8Y11_EE4BEG[15] ,
    \Tile_X8Y11_EE4BEG[14] ,
    \Tile_X8Y11_EE4BEG[13] ,
    \Tile_X8Y11_EE4BEG[12] ,
    \Tile_X8Y11_EE4BEG[11] ,
    \Tile_X8Y11_EE4BEG[10] ,
    \Tile_X8Y11_EE4BEG[9] ,
    \Tile_X8Y11_EE4BEG[8] ,
    \Tile_X8Y11_EE4BEG[7] ,
    \Tile_X8Y11_EE4BEG[6] ,
    \Tile_X8Y11_EE4BEG[5] ,
    \Tile_X8Y11_EE4BEG[4] ,
    \Tile_X8Y11_EE4BEG[3] ,
    \Tile_X8Y11_EE4BEG[2] ,
    \Tile_X8Y11_EE4BEG[1] ,
    \Tile_X8Y11_EE4BEG[0] }),
    .FrameData({\Tile_X8Y11_FrameData_O[31] ,
    \Tile_X8Y11_FrameData_O[30] ,
    \Tile_X8Y11_FrameData_O[29] ,
    \Tile_X8Y11_FrameData_O[28] ,
    \Tile_X8Y11_FrameData_O[27] ,
    \Tile_X8Y11_FrameData_O[26] ,
    \Tile_X8Y11_FrameData_O[25] ,
    \Tile_X8Y11_FrameData_O[24] ,
    \Tile_X8Y11_FrameData_O[23] ,
    \Tile_X8Y11_FrameData_O[22] ,
    \Tile_X8Y11_FrameData_O[21] ,
    \Tile_X8Y11_FrameData_O[20] ,
    \Tile_X8Y11_FrameData_O[19] ,
    \Tile_X8Y11_FrameData_O[18] ,
    \Tile_X8Y11_FrameData_O[17] ,
    \Tile_X8Y11_FrameData_O[16] ,
    \Tile_X8Y11_FrameData_O[15] ,
    \Tile_X8Y11_FrameData_O[14] ,
    \Tile_X8Y11_FrameData_O[13] ,
    \Tile_X8Y11_FrameData_O[12] ,
    \Tile_X8Y11_FrameData_O[11] ,
    \Tile_X8Y11_FrameData_O[10] ,
    \Tile_X8Y11_FrameData_O[9] ,
    \Tile_X8Y11_FrameData_O[8] ,
    \Tile_X8Y11_FrameData_O[7] ,
    \Tile_X8Y11_FrameData_O[6] ,
    \Tile_X8Y11_FrameData_O[5] ,
    \Tile_X8Y11_FrameData_O[4] ,
    \Tile_X8Y11_FrameData_O[3] ,
    \Tile_X8Y11_FrameData_O[2] ,
    \Tile_X8Y11_FrameData_O[1] ,
    \Tile_X8Y11_FrameData_O[0] }),
    .FrameData_O({\Tile_X9Y11_FrameData_O[31] ,
    \Tile_X9Y11_FrameData_O[30] ,
    \Tile_X9Y11_FrameData_O[29] ,
    \Tile_X9Y11_FrameData_O[28] ,
    \Tile_X9Y11_FrameData_O[27] ,
    \Tile_X9Y11_FrameData_O[26] ,
    \Tile_X9Y11_FrameData_O[25] ,
    \Tile_X9Y11_FrameData_O[24] ,
    \Tile_X9Y11_FrameData_O[23] ,
    \Tile_X9Y11_FrameData_O[22] ,
    \Tile_X9Y11_FrameData_O[21] ,
    \Tile_X9Y11_FrameData_O[20] ,
    \Tile_X9Y11_FrameData_O[19] ,
    \Tile_X9Y11_FrameData_O[18] ,
    \Tile_X9Y11_FrameData_O[17] ,
    \Tile_X9Y11_FrameData_O[16] ,
    \Tile_X9Y11_FrameData_O[15] ,
    \Tile_X9Y11_FrameData_O[14] ,
    \Tile_X9Y11_FrameData_O[13] ,
    \Tile_X9Y11_FrameData_O[12] ,
    \Tile_X9Y11_FrameData_O[11] ,
    \Tile_X9Y11_FrameData_O[10] ,
    \Tile_X9Y11_FrameData_O[9] ,
    \Tile_X9Y11_FrameData_O[8] ,
    \Tile_X9Y11_FrameData_O[7] ,
    \Tile_X9Y11_FrameData_O[6] ,
    \Tile_X9Y11_FrameData_O[5] ,
    \Tile_X9Y11_FrameData_O[4] ,
    \Tile_X9Y11_FrameData_O[3] ,
    \Tile_X9Y11_FrameData_O[2] ,
    \Tile_X9Y11_FrameData_O[1] ,
    \Tile_X9Y11_FrameData_O[0] }),
    .FrameStrobe({\Tile_X9Y12_FrameStrobe_O[19] ,
    \Tile_X9Y12_FrameStrobe_O[18] ,
    \Tile_X9Y12_FrameStrobe_O[17] ,
    \Tile_X9Y12_FrameStrobe_O[16] ,
    \Tile_X9Y12_FrameStrobe_O[15] ,
    \Tile_X9Y12_FrameStrobe_O[14] ,
    \Tile_X9Y12_FrameStrobe_O[13] ,
    \Tile_X9Y12_FrameStrobe_O[12] ,
    \Tile_X9Y12_FrameStrobe_O[11] ,
    \Tile_X9Y12_FrameStrobe_O[10] ,
    \Tile_X9Y12_FrameStrobe_O[9] ,
    \Tile_X9Y12_FrameStrobe_O[8] ,
    \Tile_X9Y12_FrameStrobe_O[7] ,
    \Tile_X9Y12_FrameStrobe_O[6] ,
    \Tile_X9Y12_FrameStrobe_O[5] ,
    \Tile_X9Y12_FrameStrobe_O[4] ,
    \Tile_X9Y12_FrameStrobe_O[3] ,
    \Tile_X9Y12_FrameStrobe_O[2] ,
    \Tile_X9Y12_FrameStrobe_O[1] ,
    \Tile_X9Y12_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X9Y11_FrameStrobe_O[19] ,
    \Tile_X9Y11_FrameStrobe_O[18] ,
    \Tile_X9Y11_FrameStrobe_O[17] ,
    \Tile_X9Y11_FrameStrobe_O[16] ,
    \Tile_X9Y11_FrameStrobe_O[15] ,
    \Tile_X9Y11_FrameStrobe_O[14] ,
    \Tile_X9Y11_FrameStrobe_O[13] ,
    \Tile_X9Y11_FrameStrobe_O[12] ,
    \Tile_X9Y11_FrameStrobe_O[11] ,
    \Tile_X9Y11_FrameStrobe_O[10] ,
    \Tile_X9Y11_FrameStrobe_O[9] ,
    \Tile_X9Y11_FrameStrobe_O[8] ,
    \Tile_X9Y11_FrameStrobe_O[7] ,
    \Tile_X9Y11_FrameStrobe_O[6] ,
    \Tile_X9Y11_FrameStrobe_O[5] ,
    \Tile_X9Y11_FrameStrobe_O[4] ,
    \Tile_X9Y11_FrameStrobe_O[3] ,
    \Tile_X9Y11_FrameStrobe_O[2] ,
    \Tile_X9Y11_FrameStrobe_O[1] ,
    \Tile_X9Y11_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X9Y11_N1BEG[3] ,
    \Tile_X9Y11_N1BEG[2] ,
    \Tile_X9Y11_N1BEG[1] ,
    \Tile_X9Y11_N1BEG[0] }),
    .N1END({\Tile_X9Y12_N1BEG[3] ,
    \Tile_X9Y12_N1BEG[2] ,
    \Tile_X9Y12_N1BEG[1] ,
    \Tile_X9Y12_N1BEG[0] }),
    .N2BEG({\Tile_X9Y11_N2BEG[7] ,
    \Tile_X9Y11_N2BEG[6] ,
    \Tile_X9Y11_N2BEG[5] ,
    \Tile_X9Y11_N2BEG[4] ,
    \Tile_X9Y11_N2BEG[3] ,
    \Tile_X9Y11_N2BEG[2] ,
    \Tile_X9Y11_N2BEG[1] ,
    \Tile_X9Y11_N2BEG[0] }),
    .N2BEGb({\Tile_X9Y11_N2BEGb[7] ,
    \Tile_X9Y11_N2BEGb[6] ,
    \Tile_X9Y11_N2BEGb[5] ,
    \Tile_X9Y11_N2BEGb[4] ,
    \Tile_X9Y11_N2BEGb[3] ,
    \Tile_X9Y11_N2BEGb[2] ,
    \Tile_X9Y11_N2BEGb[1] ,
    \Tile_X9Y11_N2BEGb[0] }),
    .N2END({\Tile_X9Y12_N2BEGb[7] ,
    \Tile_X9Y12_N2BEGb[6] ,
    \Tile_X9Y12_N2BEGb[5] ,
    \Tile_X9Y12_N2BEGb[4] ,
    \Tile_X9Y12_N2BEGb[3] ,
    \Tile_X9Y12_N2BEGb[2] ,
    \Tile_X9Y12_N2BEGb[1] ,
    \Tile_X9Y12_N2BEGb[0] }),
    .N2MID({\Tile_X9Y12_N2BEG[7] ,
    \Tile_X9Y12_N2BEG[6] ,
    \Tile_X9Y12_N2BEG[5] ,
    \Tile_X9Y12_N2BEG[4] ,
    \Tile_X9Y12_N2BEG[3] ,
    \Tile_X9Y12_N2BEG[2] ,
    \Tile_X9Y12_N2BEG[1] ,
    \Tile_X9Y12_N2BEG[0] }),
    .N4BEG({\Tile_X9Y11_N4BEG[15] ,
    \Tile_X9Y11_N4BEG[14] ,
    \Tile_X9Y11_N4BEG[13] ,
    \Tile_X9Y11_N4BEG[12] ,
    \Tile_X9Y11_N4BEG[11] ,
    \Tile_X9Y11_N4BEG[10] ,
    \Tile_X9Y11_N4BEG[9] ,
    \Tile_X9Y11_N4BEG[8] ,
    \Tile_X9Y11_N4BEG[7] ,
    \Tile_X9Y11_N4BEG[6] ,
    \Tile_X9Y11_N4BEG[5] ,
    \Tile_X9Y11_N4BEG[4] ,
    \Tile_X9Y11_N4BEG[3] ,
    \Tile_X9Y11_N4BEG[2] ,
    \Tile_X9Y11_N4BEG[1] ,
    \Tile_X9Y11_N4BEG[0] }),
    .N4END({\Tile_X9Y12_N4BEG[15] ,
    \Tile_X9Y12_N4BEG[14] ,
    \Tile_X9Y12_N4BEG[13] ,
    \Tile_X9Y12_N4BEG[12] ,
    \Tile_X9Y12_N4BEG[11] ,
    \Tile_X9Y12_N4BEG[10] ,
    \Tile_X9Y12_N4BEG[9] ,
    \Tile_X9Y12_N4BEG[8] ,
    \Tile_X9Y12_N4BEG[7] ,
    \Tile_X9Y12_N4BEG[6] ,
    \Tile_X9Y12_N4BEG[5] ,
    \Tile_X9Y12_N4BEG[4] ,
    \Tile_X9Y12_N4BEG[3] ,
    \Tile_X9Y12_N4BEG[2] ,
    \Tile_X9Y12_N4BEG[1] ,
    \Tile_X9Y12_N4BEG[0] }),
    .NN4BEG({\Tile_X9Y11_NN4BEG[15] ,
    \Tile_X9Y11_NN4BEG[14] ,
    \Tile_X9Y11_NN4BEG[13] ,
    \Tile_X9Y11_NN4BEG[12] ,
    \Tile_X9Y11_NN4BEG[11] ,
    \Tile_X9Y11_NN4BEG[10] ,
    \Tile_X9Y11_NN4BEG[9] ,
    \Tile_X9Y11_NN4BEG[8] ,
    \Tile_X9Y11_NN4BEG[7] ,
    \Tile_X9Y11_NN4BEG[6] ,
    \Tile_X9Y11_NN4BEG[5] ,
    \Tile_X9Y11_NN4BEG[4] ,
    \Tile_X9Y11_NN4BEG[3] ,
    \Tile_X9Y11_NN4BEG[2] ,
    \Tile_X9Y11_NN4BEG[1] ,
    \Tile_X9Y11_NN4BEG[0] }),
    .NN4END({\Tile_X9Y12_NN4BEG[15] ,
    \Tile_X9Y12_NN4BEG[14] ,
    \Tile_X9Y12_NN4BEG[13] ,
    \Tile_X9Y12_NN4BEG[12] ,
    \Tile_X9Y12_NN4BEG[11] ,
    \Tile_X9Y12_NN4BEG[10] ,
    \Tile_X9Y12_NN4BEG[9] ,
    \Tile_X9Y12_NN4BEG[8] ,
    \Tile_X9Y12_NN4BEG[7] ,
    \Tile_X9Y12_NN4BEG[6] ,
    \Tile_X9Y12_NN4BEG[5] ,
    \Tile_X9Y12_NN4BEG[4] ,
    \Tile_X9Y12_NN4BEG[3] ,
    \Tile_X9Y12_NN4BEG[2] ,
    \Tile_X9Y12_NN4BEG[1] ,
    \Tile_X9Y12_NN4BEG[0] }),
    .S1BEG({\Tile_X9Y11_S1BEG[3] ,
    \Tile_X9Y11_S1BEG[2] ,
    \Tile_X9Y11_S1BEG[1] ,
    \Tile_X9Y11_S1BEG[0] }),
    .S1END({\Tile_X9Y10_S1BEG[3] ,
    \Tile_X9Y10_S1BEG[2] ,
    \Tile_X9Y10_S1BEG[1] ,
    \Tile_X9Y10_S1BEG[0] }),
    .S2BEG({\Tile_X9Y11_S2BEG[7] ,
    \Tile_X9Y11_S2BEG[6] ,
    \Tile_X9Y11_S2BEG[5] ,
    \Tile_X9Y11_S2BEG[4] ,
    \Tile_X9Y11_S2BEG[3] ,
    \Tile_X9Y11_S2BEG[2] ,
    \Tile_X9Y11_S2BEG[1] ,
    \Tile_X9Y11_S2BEG[0] }),
    .S2BEGb({\Tile_X9Y11_S2BEGb[7] ,
    \Tile_X9Y11_S2BEGb[6] ,
    \Tile_X9Y11_S2BEGb[5] ,
    \Tile_X9Y11_S2BEGb[4] ,
    \Tile_X9Y11_S2BEGb[3] ,
    \Tile_X9Y11_S2BEGb[2] ,
    \Tile_X9Y11_S2BEGb[1] ,
    \Tile_X9Y11_S2BEGb[0] }),
    .S2END({\Tile_X9Y10_S2BEGb[7] ,
    \Tile_X9Y10_S2BEGb[6] ,
    \Tile_X9Y10_S2BEGb[5] ,
    \Tile_X9Y10_S2BEGb[4] ,
    \Tile_X9Y10_S2BEGb[3] ,
    \Tile_X9Y10_S2BEGb[2] ,
    \Tile_X9Y10_S2BEGb[1] ,
    \Tile_X9Y10_S2BEGb[0] }),
    .S2MID({\Tile_X9Y10_S2BEG[7] ,
    \Tile_X9Y10_S2BEG[6] ,
    \Tile_X9Y10_S2BEG[5] ,
    \Tile_X9Y10_S2BEG[4] ,
    \Tile_X9Y10_S2BEG[3] ,
    \Tile_X9Y10_S2BEG[2] ,
    \Tile_X9Y10_S2BEG[1] ,
    \Tile_X9Y10_S2BEG[0] }),
    .S4BEG({\Tile_X9Y11_S4BEG[15] ,
    \Tile_X9Y11_S4BEG[14] ,
    \Tile_X9Y11_S4BEG[13] ,
    \Tile_X9Y11_S4BEG[12] ,
    \Tile_X9Y11_S4BEG[11] ,
    \Tile_X9Y11_S4BEG[10] ,
    \Tile_X9Y11_S4BEG[9] ,
    \Tile_X9Y11_S4BEG[8] ,
    \Tile_X9Y11_S4BEG[7] ,
    \Tile_X9Y11_S4BEG[6] ,
    \Tile_X9Y11_S4BEG[5] ,
    \Tile_X9Y11_S4BEG[4] ,
    \Tile_X9Y11_S4BEG[3] ,
    \Tile_X9Y11_S4BEG[2] ,
    \Tile_X9Y11_S4BEG[1] ,
    \Tile_X9Y11_S4BEG[0] }),
    .S4END({\Tile_X9Y10_S4BEG[15] ,
    \Tile_X9Y10_S4BEG[14] ,
    \Tile_X9Y10_S4BEG[13] ,
    \Tile_X9Y10_S4BEG[12] ,
    \Tile_X9Y10_S4BEG[11] ,
    \Tile_X9Y10_S4BEG[10] ,
    \Tile_X9Y10_S4BEG[9] ,
    \Tile_X9Y10_S4BEG[8] ,
    \Tile_X9Y10_S4BEG[7] ,
    \Tile_X9Y10_S4BEG[6] ,
    \Tile_X9Y10_S4BEG[5] ,
    \Tile_X9Y10_S4BEG[4] ,
    \Tile_X9Y10_S4BEG[3] ,
    \Tile_X9Y10_S4BEG[2] ,
    \Tile_X9Y10_S4BEG[1] ,
    \Tile_X9Y10_S4BEG[0] }),
    .SS4BEG({\Tile_X9Y11_SS4BEG[15] ,
    \Tile_X9Y11_SS4BEG[14] ,
    \Tile_X9Y11_SS4BEG[13] ,
    \Tile_X9Y11_SS4BEG[12] ,
    \Tile_X9Y11_SS4BEG[11] ,
    \Tile_X9Y11_SS4BEG[10] ,
    \Tile_X9Y11_SS4BEG[9] ,
    \Tile_X9Y11_SS4BEG[8] ,
    \Tile_X9Y11_SS4BEG[7] ,
    \Tile_X9Y11_SS4BEG[6] ,
    \Tile_X9Y11_SS4BEG[5] ,
    \Tile_X9Y11_SS4BEG[4] ,
    \Tile_X9Y11_SS4BEG[3] ,
    \Tile_X9Y11_SS4BEG[2] ,
    \Tile_X9Y11_SS4BEG[1] ,
    \Tile_X9Y11_SS4BEG[0] }),
    .SS4END({\Tile_X9Y10_SS4BEG[15] ,
    \Tile_X9Y10_SS4BEG[14] ,
    \Tile_X9Y10_SS4BEG[13] ,
    \Tile_X9Y10_SS4BEG[12] ,
    \Tile_X9Y10_SS4BEG[11] ,
    \Tile_X9Y10_SS4BEG[10] ,
    \Tile_X9Y10_SS4BEG[9] ,
    \Tile_X9Y10_SS4BEG[8] ,
    \Tile_X9Y10_SS4BEG[7] ,
    \Tile_X9Y10_SS4BEG[6] ,
    \Tile_X9Y10_SS4BEG[5] ,
    \Tile_X9Y10_SS4BEG[4] ,
    \Tile_X9Y10_SS4BEG[3] ,
    \Tile_X9Y10_SS4BEG[2] ,
    \Tile_X9Y10_SS4BEG[1] ,
    \Tile_X9Y10_SS4BEG[0] }),
    .W1BEG({\Tile_X9Y11_W1BEG[3] ,
    \Tile_X9Y11_W1BEG[2] ,
    \Tile_X9Y11_W1BEG[1] ,
    \Tile_X9Y11_W1BEG[0] }),
    .W1END({\Tile_X10Y11_W1BEG[3] ,
    \Tile_X10Y11_W1BEG[2] ,
    \Tile_X10Y11_W1BEG[1] ,
    \Tile_X10Y11_W1BEG[0] }),
    .W2BEG({\Tile_X9Y11_W2BEG[7] ,
    \Tile_X9Y11_W2BEG[6] ,
    \Tile_X9Y11_W2BEG[5] ,
    \Tile_X9Y11_W2BEG[4] ,
    \Tile_X9Y11_W2BEG[3] ,
    \Tile_X9Y11_W2BEG[2] ,
    \Tile_X9Y11_W2BEG[1] ,
    \Tile_X9Y11_W2BEG[0] }),
    .W2BEGb({\Tile_X9Y11_W2BEGb[7] ,
    \Tile_X9Y11_W2BEGb[6] ,
    \Tile_X9Y11_W2BEGb[5] ,
    \Tile_X9Y11_W2BEGb[4] ,
    \Tile_X9Y11_W2BEGb[3] ,
    \Tile_X9Y11_W2BEGb[2] ,
    \Tile_X9Y11_W2BEGb[1] ,
    \Tile_X9Y11_W2BEGb[0] }),
    .W2END({\Tile_X10Y11_W2BEGb[7] ,
    \Tile_X10Y11_W2BEGb[6] ,
    \Tile_X10Y11_W2BEGb[5] ,
    \Tile_X10Y11_W2BEGb[4] ,
    \Tile_X10Y11_W2BEGb[3] ,
    \Tile_X10Y11_W2BEGb[2] ,
    \Tile_X10Y11_W2BEGb[1] ,
    \Tile_X10Y11_W2BEGb[0] }),
    .W2MID({\Tile_X10Y11_W2BEG[7] ,
    \Tile_X10Y11_W2BEG[6] ,
    \Tile_X10Y11_W2BEG[5] ,
    \Tile_X10Y11_W2BEG[4] ,
    \Tile_X10Y11_W2BEG[3] ,
    \Tile_X10Y11_W2BEG[2] ,
    \Tile_X10Y11_W2BEG[1] ,
    \Tile_X10Y11_W2BEG[0] }),
    .W6BEG({\Tile_X9Y11_W6BEG[11] ,
    \Tile_X9Y11_W6BEG[10] ,
    \Tile_X9Y11_W6BEG[9] ,
    \Tile_X9Y11_W6BEG[8] ,
    \Tile_X9Y11_W6BEG[7] ,
    \Tile_X9Y11_W6BEG[6] ,
    \Tile_X9Y11_W6BEG[5] ,
    \Tile_X9Y11_W6BEG[4] ,
    \Tile_X9Y11_W6BEG[3] ,
    \Tile_X9Y11_W6BEG[2] ,
    \Tile_X9Y11_W6BEG[1] ,
    \Tile_X9Y11_W6BEG[0] }),
    .W6END({\Tile_X10Y11_W6BEG[11] ,
    \Tile_X10Y11_W6BEG[10] ,
    \Tile_X10Y11_W6BEG[9] ,
    \Tile_X10Y11_W6BEG[8] ,
    \Tile_X10Y11_W6BEG[7] ,
    \Tile_X10Y11_W6BEG[6] ,
    \Tile_X10Y11_W6BEG[5] ,
    \Tile_X10Y11_W6BEG[4] ,
    \Tile_X10Y11_W6BEG[3] ,
    \Tile_X10Y11_W6BEG[2] ,
    \Tile_X10Y11_W6BEG[1] ,
    \Tile_X10Y11_W6BEG[0] }),
    .WW4BEG({\Tile_X9Y11_WW4BEG[15] ,
    \Tile_X9Y11_WW4BEG[14] ,
    \Tile_X9Y11_WW4BEG[13] ,
    \Tile_X9Y11_WW4BEG[12] ,
    \Tile_X9Y11_WW4BEG[11] ,
    \Tile_X9Y11_WW4BEG[10] ,
    \Tile_X9Y11_WW4BEG[9] ,
    \Tile_X9Y11_WW4BEG[8] ,
    \Tile_X9Y11_WW4BEG[7] ,
    \Tile_X9Y11_WW4BEG[6] ,
    \Tile_X9Y11_WW4BEG[5] ,
    \Tile_X9Y11_WW4BEG[4] ,
    \Tile_X9Y11_WW4BEG[3] ,
    \Tile_X9Y11_WW4BEG[2] ,
    \Tile_X9Y11_WW4BEG[1] ,
    \Tile_X9Y11_WW4BEG[0] }),
    .WW4END({\Tile_X10Y11_WW4BEG[15] ,
    \Tile_X10Y11_WW4BEG[14] ,
    \Tile_X10Y11_WW4BEG[13] ,
    \Tile_X10Y11_WW4BEG[12] ,
    \Tile_X10Y11_WW4BEG[11] ,
    \Tile_X10Y11_WW4BEG[10] ,
    \Tile_X10Y11_WW4BEG[9] ,
    \Tile_X10Y11_WW4BEG[8] ,
    \Tile_X10Y11_WW4BEG[7] ,
    \Tile_X10Y11_WW4BEG[6] ,
    \Tile_X10Y11_WW4BEG[5] ,
    \Tile_X10Y11_WW4BEG[4] ,
    \Tile_X10Y11_WW4BEG[3] ,
    \Tile_X10Y11_WW4BEG[2] ,
    \Tile_X10Y11_WW4BEG[1] ,
    \Tile_X10Y11_WW4BEG[0] }));
 LUT4AB Tile_X9Y12_LUT4AB (.Ci(Tile_X9Y13_Co),
    .Co(Tile_X9Y12_Co),
    .UserCLK(Tile_X9Y13_UserCLKo),
    .UserCLKo(Tile_X9Y12_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X9Y12_E1BEG[3] ,
    \Tile_X9Y12_E1BEG[2] ,
    \Tile_X9Y12_E1BEG[1] ,
    \Tile_X9Y12_E1BEG[0] }),
    .E1END({\Tile_X8Y12_E1BEG[3] ,
    \Tile_X8Y12_E1BEG[2] ,
    \Tile_X8Y12_E1BEG[1] ,
    \Tile_X8Y12_E1BEG[0] }),
    .E2BEG({\Tile_X9Y12_E2BEG[7] ,
    \Tile_X9Y12_E2BEG[6] ,
    \Tile_X9Y12_E2BEG[5] ,
    \Tile_X9Y12_E2BEG[4] ,
    \Tile_X9Y12_E2BEG[3] ,
    \Tile_X9Y12_E2BEG[2] ,
    \Tile_X9Y12_E2BEG[1] ,
    \Tile_X9Y12_E2BEG[0] }),
    .E2BEGb({\Tile_X9Y12_E2BEGb[7] ,
    \Tile_X9Y12_E2BEGb[6] ,
    \Tile_X9Y12_E2BEGb[5] ,
    \Tile_X9Y12_E2BEGb[4] ,
    \Tile_X9Y12_E2BEGb[3] ,
    \Tile_X9Y12_E2BEGb[2] ,
    \Tile_X9Y12_E2BEGb[1] ,
    \Tile_X9Y12_E2BEGb[0] }),
    .E2END({\Tile_X8Y12_E2BEGb[7] ,
    \Tile_X8Y12_E2BEGb[6] ,
    \Tile_X8Y12_E2BEGb[5] ,
    \Tile_X8Y12_E2BEGb[4] ,
    \Tile_X8Y12_E2BEGb[3] ,
    \Tile_X8Y12_E2BEGb[2] ,
    \Tile_X8Y12_E2BEGb[1] ,
    \Tile_X8Y12_E2BEGb[0] }),
    .E2MID({\Tile_X8Y12_E2BEG[7] ,
    \Tile_X8Y12_E2BEG[6] ,
    \Tile_X8Y12_E2BEG[5] ,
    \Tile_X8Y12_E2BEG[4] ,
    \Tile_X8Y12_E2BEG[3] ,
    \Tile_X8Y12_E2BEG[2] ,
    \Tile_X8Y12_E2BEG[1] ,
    \Tile_X8Y12_E2BEG[0] }),
    .E6BEG({\Tile_X9Y12_E6BEG[11] ,
    \Tile_X9Y12_E6BEG[10] ,
    \Tile_X9Y12_E6BEG[9] ,
    \Tile_X9Y12_E6BEG[8] ,
    \Tile_X9Y12_E6BEG[7] ,
    \Tile_X9Y12_E6BEG[6] ,
    \Tile_X9Y12_E6BEG[5] ,
    \Tile_X9Y12_E6BEG[4] ,
    \Tile_X9Y12_E6BEG[3] ,
    \Tile_X9Y12_E6BEG[2] ,
    \Tile_X9Y12_E6BEG[1] ,
    \Tile_X9Y12_E6BEG[0] }),
    .E6END({\Tile_X8Y12_E6BEG[11] ,
    \Tile_X8Y12_E6BEG[10] ,
    \Tile_X8Y12_E6BEG[9] ,
    \Tile_X8Y12_E6BEG[8] ,
    \Tile_X8Y12_E6BEG[7] ,
    \Tile_X8Y12_E6BEG[6] ,
    \Tile_X8Y12_E6BEG[5] ,
    \Tile_X8Y12_E6BEG[4] ,
    \Tile_X8Y12_E6BEG[3] ,
    \Tile_X8Y12_E6BEG[2] ,
    \Tile_X8Y12_E6BEG[1] ,
    \Tile_X8Y12_E6BEG[0] }),
    .EE4BEG({\Tile_X9Y12_EE4BEG[15] ,
    \Tile_X9Y12_EE4BEG[14] ,
    \Tile_X9Y12_EE4BEG[13] ,
    \Tile_X9Y12_EE4BEG[12] ,
    \Tile_X9Y12_EE4BEG[11] ,
    \Tile_X9Y12_EE4BEG[10] ,
    \Tile_X9Y12_EE4BEG[9] ,
    \Tile_X9Y12_EE4BEG[8] ,
    \Tile_X9Y12_EE4BEG[7] ,
    \Tile_X9Y12_EE4BEG[6] ,
    \Tile_X9Y12_EE4BEG[5] ,
    \Tile_X9Y12_EE4BEG[4] ,
    \Tile_X9Y12_EE4BEG[3] ,
    \Tile_X9Y12_EE4BEG[2] ,
    \Tile_X9Y12_EE4BEG[1] ,
    \Tile_X9Y12_EE4BEG[0] }),
    .EE4END({\Tile_X8Y12_EE4BEG[15] ,
    \Tile_X8Y12_EE4BEG[14] ,
    \Tile_X8Y12_EE4BEG[13] ,
    \Tile_X8Y12_EE4BEG[12] ,
    \Tile_X8Y12_EE4BEG[11] ,
    \Tile_X8Y12_EE4BEG[10] ,
    \Tile_X8Y12_EE4BEG[9] ,
    \Tile_X8Y12_EE4BEG[8] ,
    \Tile_X8Y12_EE4BEG[7] ,
    \Tile_X8Y12_EE4BEG[6] ,
    \Tile_X8Y12_EE4BEG[5] ,
    \Tile_X8Y12_EE4BEG[4] ,
    \Tile_X8Y12_EE4BEG[3] ,
    \Tile_X8Y12_EE4BEG[2] ,
    \Tile_X8Y12_EE4BEG[1] ,
    \Tile_X8Y12_EE4BEG[0] }),
    .FrameData({\Tile_X8Y12_FrameData_O[31] ,
    \Tile_X8Y12_FrameData_O[30] ,
    \Tile_X8Y12_FrameData_O[29] ,
    \Tile_X8Y12_FrameData_O[28] ,
    \Tile_X8Y12_FrameData_O[27] ,
    \Tile_X8Y12_FrameData_O[26] ,
    \Tile_X8Y12_FrameData_O[25] ,
    \Tile_X8Y12_FrameData_O[24] ,
    \Tile_X8Y12_FrameData_O[23] ,
    \Tile_X8Y12_FrameData_O[22] ,
    \Tile_X8Y12_FrameData_O[21] ,
    \Tile_X8Y12_FrameData_O[20] ,
    \Tile_X8Y12_FrameData_O[19] ,
    \Tile_X8Y12_FrameData_O[18] ,
    \Tile_X8Y12_FrameData_O[17] ,
    \Tile_X8Y12_FrameData_O[16] ,
    \Tile_X8Y12_FrameData_O[15] ,
    \Tile_X8Y12_FrameData_O[14] ,
    \Tile_X8Y12_FrameData_O[13] ,
    \Tile_X8Y12_FrameData_O[12] ,
    \Tile_X8Y12_FrameData_O[11] ,
    \Tile_X8Y12_FrameData_O[10] ,
    \Tile_X8Y12_FrameData_O[9] ,
    \Tile_X8Y12_FrameData_O[8] ,
    \Tile_X8Y12_FrameData_O[7] ,
    \Tile_X8Y12_FrameData_O[6] ,
    \Tile_X8Y12_FrameData_O[5] ,
    \Tile_X8Y12_FrameData_O[4] ,
    \Tile_X8Y12_FrameData_O[3] ,
    \Tile_X8Y12_FrameData_O[2] ,
    \Tile_X8Y12_FrameData_O[1] ,
    \Tile_X8Y12_FrameData_O[0] }),
    .FrameData_O({\Tile_X9Y12_FrameData_O[31] ,
    \Tile_X9Y12_FrameData_O[30] ,
    \Tile_X9Y12_FrameData_O[29] ,
    \Tile_X9Y12_FrameData_O[28] ,
    \Tile_X9Y12_FrameData_O[27] ,
    \Tile_X9Y12_FrameData_O[26] ,
    \Tile_X9Y12_FrameData_O[25] ,
    \Tile_X9Y12_FrameData_O[24] ,
    \Tile_X9Y12_FrameData_O[23] ,
    \Tile_X9Y12_FrameData_O[22] ,
    \Tile_X9Y12_FrameData_O[21] ,
    \Tile_X9Y12_FrameData_O[20] ,
    \Tile_X9Y12_FrameData_O[19] ,
    \Tile_X9Y12_FrameData_O[18] ,
    \Tile_X9Y12_FrameData_O[17] ,
    \Tile_X9Y12_FrameData_O[16] ,
    \Tile_X9Y12_FrameData_O[15] ,
    \Tile_X9Y12_FrameData_O[14] ,
    \Tile_X9Y12_FrameData_O[13] ,
    \Tile_X9Y12_FrameData_O[12] ,
    \Tile_X9Y12_FrameData_O[11] ,
    \Tile_X9Y12_FrameData_O[10] ,
    \Tile_X9Y12_FrameData_O[9] ,
    \Tile_X9Y12_FrameData_O[8] ,
    \Tile_X9Y12_FrameData_O[7] ,
    \Tile_X9Y12_FrameData_O[6] ,
    \Tile_X9Y12_FrameData_O[5] ,
    \Tile_X9Y12_FrameData_O[4] ,
    \Tile_X9Y12_FrameData_O[3] ,
    \Tile_X9Y12_FrameData_O[2] ,
    \Tile_X9Y12_FrameData_O[1] ,
    \Tile_X9Y12_FrameData_O[0] }),
    .FrameStrobe({\Tile_X9Y13_FrameStrobe_O[19] ,
    \Tile_X9Y13_FrameStrobe_O[18] ,
    \Tile_X9Y13_FrameStrobe_O[17] ,
    \Tile_X9Y13_FrameStrobe_O[16] ,
    \Tile_X9Y13_FrameStrobe_O[15] ,
    \Tile_X9Y13_FrameStrobe_O[14] ,
    \Tile_X9Y13_FrameStrobe_O[13] ,
    \Tile_X9Y13_FrameStrobe_O[12] ,
    \Tile_X9Y13_FrameStrobe_O[11] ,
    \Tile_X9Y13_FrameStrobe_O[10] ,
    \Tile_X9Y13_FrameStrobe_O[9] ,
    \Tile_X9Y13_FrameStrobe_O[8] ,
    \Tile_X9Y13_FrameStrobe_O[7] ,
    \Tile_X9Y13_FrameStrobe_O[6] ,
    \Tile_X9Y13_FrameStrobe_O[5] ,
    \Tile_X9Y13_FrameStrobe_O[4] ,
    \Tile_X9Y13_FrameStrobe_O[3] ,
    \Tile_X9Y13_FrameStrobe_O[2] ,
    \Tile_X9Y13_FrameStrobe_O[1] ,
    \Tile_X9Y13_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X9Y12_FrameStrobe_O[19] ,
    \Tile_X9Y12_FrameStrobe_O[18] ,
    \Tile_X9Y12_FrameStrobe_O[17] ,
    \Tile_X9Y12_FrameStrobe_O[16] ,
    \Tile_X9Y12_FrameStrobe_O[15] ,
    \Tile_X9Y12_FrameStrobe_O[14] ,
    \Tile_X9Y12_FrameStrobe_O[13] ,
    \Tile_X9Y12_FrameStrobe_O[12] ,
    \Tile_X9Y12_FrameStrobe_O[11] ,
    \Tile_X9Y12_FrameStrobe_O[10] ,
    \Tile_X9Y12_FrameStrobe_O[9] ,
    \Tile_X9Y12_FrameStrobe_O[8] ,
    \Tile_X9Y12_FrameStrobe_O[7] ,
    \Tile_X9Y12_FrameStrobe_O[6] ,
    \Tile_X9Y12_FrameStrobe_O[5] ,
    \Tile_X9Y12_FrameStrobe_O[4] ,
    \Tile_X9Y12_FrameStrobe_O[3] ,
    \Tile_X9Y12_FrameStrobe_O[2] ,
    \Tile_X9Y12_FrameStrobe_O[1] ,
    \Tile_X9Y12_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X9Y12_N1BEG[3] ,
    \Tile_X9Y12_N1BEG[2] ,
    \Tile_X9Y12_N1BEG[1] ,
    \Tile_X9Y12_N1BEG[0] }),
    .N1END({\Tile_X9Y13_N1BEG[3] ,
    \Tile_X9Y13_N1BEG[2] ,
    \Tile_X9Y13_N1BEG[1] ,
    \Tile_X9Y13_N1BEG[0] }),
    .N2BEG({\Tile_X9Y12_N2BEG[7] ,
    \Tile_X9Y12_N2BEG[6] ,
    \Tile_X9Y12_N2BEG[5] ,
    \Tile_X9Y12_N2BEG[4] ,
    \Tile_X9Y12_N2BEG[3] ,
    \Tile_X9Y12_N2BEG[2] ,
    \Tile_X9Y12_N2BEG[1] ,
    \Tile_X9Y12_N2BEG[0] }),
    .N2BEGb({\Tile_X9Y12_N2BEGb[7] ,
    \Tile_X9Y12_N2BEGb[6] ,
    \Tile_X9Y12_N2BEGb[5] ,
    \Tile_X9Y12_N2BEGb[4] ,
    \Tile_X9Y12_N2BEGb[3] ,
    \Tile_X9Y12_N2BEGb[2] ,
    \Tile_X9Y12_N2BEGb[1] ,
    \Tile_X9Y12_N2BEGb[0] }),
    .N2END({\Tile_X9Y13_N2BEGb[7] ,
    \Tile_X9Y13_N2BEGb[6] ,
    \Tile_X9Y13_N2BEGb[5] ,
    \Tile_X9Y13_N2BEGb[4] ,
    \Tile_X9Y13_N2BEGb[3] ,
    \Tile_X9Y13_N2BEGb[2] ,
    \Tile_X9Y13_N2BEGb[1] ,
    \Tile_X9Y13_N2BEGb[0] }),
    .N2MID({\Tile_X9Y13_N2BEG[7] ,
    \Tile_X9Y13_N2BEG[6] ,
    \Tile_X9Y13_N2BEG[5] ,
    \Tile_X9Y13_N2BEG[4] ,
    \Tile_X9Y13_N2BEG[3] ,
    \Tile_X9Y13_N2BEG[2] ,
    \Tile_X9Y13_N2BEG[1] ,
    \Tile_X9Y13_N2BEG[0] }),
    .N4BEG({\Tile_X9Y12_N4BEG[15] ,
    \Tile_X9Y12_N4BEG[14] ,
    \Tile_X9Y12_N4BEG[13] ,
    \Tile_X9Y12_N4BEG[12] ,
    \Tile_X9Y12_N4BEG[11] ,
    \Tile_X9Y12_N4BEG[10] ,
    \Tile_X9Y12_N4BEG[9] ,
    \Tile_X9Y12_N4BEG[8] ,
    \Tile_X9Y12_N4BEG[7] ,
    \Tile_X9Y12_N4BEG[6] ,
    \Tile_X9Y12_N4BEG[5] ,
    \Tile_X9Y12_N4BEG[4] ,
    \Tile_X9Y12_N4BEG[3] ,
    \Tile_X9Y12_N4BEG[2] ,
    \Tile_X9Y12_N4BEG[1] ,
    \Tile_X9Y12_N4BEG[0] }),
    .N4END({\Tile_X9Y13_N4BEG[15] ,
    \Tile_X9Y13_N4BEG[14] ,
    \Tile_X9Y13_N4BEG[13] ,
    \Tile_X9Y13_N4BEG[12] ,
    \Tile_X9Y13_N4BEG[11] ,
    \Tile_X9Y13_N4BEG[10] ,
    \Tile_X9Y13_N4BEG[9] ,
    \Tile_X9Y13_N4BEG[8] ,
    \Tile_X9Y13_N4BEG[7] ,
    \Tile_X9Y13_N4BEG[6] ,
    \Tile_X9Y13_N4BEG[5] ,
    \Tile_X9Y13_N4BEG[4] ,
    \Tile_X9Y13_N4BEG[3] ,
    \Tile_X9Y13_N4BEG[2] ,
    \Tile_X9Y13_N4BEG[1] ,
    \Tile_X9Y13_N4BEG[0] }),
    .NN4BEG({\Tile_X9Y12_NN4BEG[15] ,
    \Tile_X9Y12_NN4BEG[14] ,
    \Tile_X9Y12_NN4BEG[13] ,
    \Tile_X9Y12_NN4BEG[12] ,
    \Tile_X9Y12_NN4BEG[11] ,
    \Tile_X9Y12_NN4BEG[10] ,
    \Tile_X9Y12_NN4BEG[9] ,
    \Tile_X9Y12_NN4BEG[8] ,
    \Tile_X9Y12_NN4BEG[7] ,
    \Tile_X9Y12_NN4BEG[6] ,
    \Tile_X9Y12_NN4BEG[5] ,
    \Tile_X9Y12_NN4BEG[4] ,
    \Tile_X9Y12_NN4BEG[3] ,
    \Tile_X9Y12_NN4BEG[2] ,
    \Tile_X9Y12_NN4BEG[1] ,
    \Tile_X9Y12_NN4BEG[0] }),
    .NN4END({\Tile_X9Y13_NN4BEG[15] ,
    \Tile_X9Y13_NN4BEG[14] ,
    \Tile_X9Y13_NN4BEG[13] ,
    \Tile_X9Y13_NN4BEG[12] ,
    \Tile_X9Y13_NN4BEG[11] ,
    \Tile_X9Y13_NN4BEG[10] ,
    \Tile_X9Y13_NN4BEG[9] ,
    \Tile_X9Y13_NN4BEG[8] ,
    \Tile_X9Y13_NN4BEG[7] ,
    \Tile_X9Y13_NN4BEG[6] ,
    \Tile_X9Y13_NN4BEG[5] ,
    \Tile_X9Y13_NN4BEG[4] ,
    \Tile_X9Y13_NN4BEG[3] ,
    \Tile_X9Y13_NN4BEG[2] ,
    \Tile_X9Y13_NN4BEG[1] ,
    \Tile_X9Y13_NN4BEG[0] }),
    .S1BEG({\Tile_X9Y12_S1BEG[3] ,
    \Tile_X9Y12_S1BEG[2] ,
    \Tile_X9Y12_S1BEG[1] ,
    \Tile_X9Y12_S1BEG[0] }),
    .S1END({\Tile_X9Y11_S1BEG[3] ,
    \Tile_X9Y11_S1BEG[2] ,
    \Tile_X9Y11_S1BEG[1] ,
    \Tile_X9Y11_S1BEG[0] }),
    .S2BEG({\Tile_X9Y12_S2BEG[7] ,
    \Tile_X9Y12_S2BEG[6] ,
    \Tile_X9Y12_S2BEG[5] ,
    \Tile_X9Y12_S2BEG[4] ,
    \Tile_X9Y12_S2BEG[3] ,
    \Tile_X9Y12_S2BEG[2] ,
    \Tile_X9Y12_S2BEG[1] ,
    \Tile_X9Y12_S2BEG[0] }),
    .S2BEGb({\Tile_X9Y12_S2BEGb[7] ,
    \Tile_X9Y12_S2BEGb[6] ,
    \Tile_X9Y12_S2BEGb[5] ,
    \Tile_X9Y12_S2BEGb[4] ,
    \Tile_X9Y12_S2BEGb[3] ,
    \Tile_X9Y12_S2BEGb[2] ,
    \Tile_X9Y12_S2BEGb[1] ,
    \Tile_X9Y12_S2BEGb[0] }),
    .S2END({\Tile_X9Y11_S2BEGb[7] ,
    \Tile_X9Y11_S2BEGb[6] ,
    \Tile_X9Y11_S2BEGb[5] ,
    \Tile_X9Y11_S2BEGb[4] ,
    \Tile_X9Y11_S2BEGb[3] ,
    \Tile_X9Y11_S2BEGb[2] ,
    \Tile_X9Y11_S2BEGb[1] ,
    \Tile_X9Y11_S2BEGb[0] }),
    .S2MID({\Tile_X9Y11_S2BEG[7] ,
    \Tile_X9Y11_S2BEG[6] ,
    \Tile_X9Y11_S2BEG[5] ,
    \Tile_X9Y11_S2BEG[4] ,
    \Tile_X9Y11_S2BEG[3] ,
    \Tile_X9Y11_S2BEG[2] ,
    \Tile_X9Y11_S2BEG[1] ,
    \Tile_X9Y11_S2BEG[0] }),
    .S4BEG({\Tile_X9Y12_S4BEG[15] ,
    \Tile_X9Y12_S4BEG[14] ,
    \Tile_X9Y12_S4BEG[13] ,
    \Tile_X9Y12_S4BEG[12] ,
    \Tile_X9Y12_S4BEG[11] ,
    \Tile_X9Y12_S4BEG[10] ,
    \Tile_X9Y12_S4BEG[9] ,
    \Tile_X9Y12_S4BEG[8] ,
    \Tile_X9Y12_S4BEG[7] ,
    \Tile_X9Y12_S4BEG[6] ,
    \Tile_X9Y12_S4BEG[5] ,
    \Tile_X9Y12_S4BEG[4] ,
    \Tile_X9Y12_S4BEG[3] ,
    \Tile_X9Y12_S4BEG[2] ,
    \Tile_X9Y12_S4BEG[1] ,
    \Tile_X9Y12_S4BEG[0] }),
    .S4END({\Tile_X9Y11_S4BEG[15] ,
    \Tile_X9Y11_S4BEG[14] ,
    \Tile_X9Y11_S4BEG[13] ,
    \Tile_X9Y11_S4BEG[12] ,
    \Tile_X9Y11_S4BEG[11] ,
    \Tile_X9Y11_S4BEG[10] ,
    \Tile_X9Y11_S4BEG[9] ,
    \Tile_X9Y11_S4BEG[8] ,
    \Tile_X9Y11_S4BEG[7] ,
    \Tile_X9Y11_S4BEG[6] ,
    \Tile_X9Y11_S4BEG[5] ,
    \Tile_X9Y11_S4BEG[4] ,
    \Tile_X9Y11_S4BEG[3] ,
    \Tile_X9Y11_S4BEG[2] ,
    \Tile_X9Y11_S4BEG[1] ,
    \Tile_X9Y11_S4BEG[0] }),
    .SS4BEG({\Tile_X9Y12_SS4BEG[15] ,
    \Tile_X9Y12_SS4BEG[14] ,
    \Tile_X9Y12_SS4BEG[13] ,
    \Tile_X9Y12_SS4BEG[12] ,
    \Tile_X9Y12_SS4BEG[11] ,
    \Tile_X9Y12_SS4BEG[10] ,
    \Tile_X9Y12_SS4BEG[9] ,
    \Tile_X9Y12_SS4BEG[8] ,
    \Tile_X9Y12_SS4BEG[7] ,
    \Tile_X9Y12_SS4BEG[6] ,
    \Tile_X9Y12_SS4BEG[5] ,
    \Tile_X9Y12_SS4BEG[4] ,
    \Tile_X9Y12_SS4BEG[3] ,
    \Tile_X9Y12_SS4BEG[2] ,
    \Tile_X9Y12_SS4BEG[1] ,
    \Tile_X9Y12_SS4BEG[0] }),
    .SS4END({\Tile_X9Y11_SS4BEG[15] ,
    \Tile_X9Y11_SS4BEG[14] ,
    \Tile_X9Y11_SS4BEG[13] ,
    \Tile_X9Y11_SS4BEG[12] ,
    \Tile_X9Y11_SS4BEG[11] ,
    \Tile_X9Y11_SS4BEG[10] ,
    \Tile_X9Y11_SS4BEG[9] ,
    \Tile_X9Y11_SS4BEG[8] ,
    \Tile_X9Y11_SS4BEG[7] ,
    \Tile_X9Y11_SS4BEG[6] ,
    \Tile_X9Y11_SS4BEG[5] ,
    \Tile_X9Y11_SS4BEG[4] ,
    \Tile_X9Y11_SS4BEG[3] ,
    \Tile_X9Y11_SS4BEG[2] ,
    \Tile_X9Y11_SS4BEG[1] ,
    \Tile_X9Y11_SS4BEG[0] }),
    .W1BEG({\Tile_X9Y12_W1BEG[3] ,
    \Tile_X9Y12_W1BEG[2] ,
    \Tile_X9Y12_W1BEG[1] ,
    \Tile_X9Y12_W1BEG[0] }),
    .W1END({\Tile_X10Y12_W1BEG[3] ,
    \Tile_X10Y12_W1BEG[2] ,
    \Tile_X10Y12_W1BEG[1] ,
    \Tile_X10Y12_W1BEG[0] }),
    .W2BEG({\Tile_X9Y12_W2BEG[7] ,
    \Tile_X9Y12_W2BEG[6] ,
    \Tile_X9Y12_W2BEG[5] ,
    \Tile_X9Y12_W2BEG[4] ,
    \Tile_X9Y12_W2BEG[3] ,
    \Tile_X9Y12_W2BEG[2] ,
    \Tile_X9Y12_W2BEG[1] ,
    \Tile_X9Y12_W2BEG[0] }),
    .W2BEGb({\Tile_X9Y12_W2BEGb[7] ,
    \Tile_X9Y12_W2BEGb[6] ,
    \Tile_X9Y12_W2BEGb[5] ,
    \Tile_X9Y12_W2BEGb[4] ,
    \Tile_X9Y12_W2BEGb[3] ,
    \Tile_X9Y12_W2BEGb[2] ,
    \Tile_X9Y12_W2BEGb[1] ,
    \Tile_X9Y12_W2BEGb[0] }),
    .W2END({\Tile_X10Y12_W2BEGb[7] ,
    \Tile_X10Y12_W2BEGb[6] ,
    \Tile_X10Y12_W2BEGb[5] ,
    \Tile_X10Y12_W2BEGb[4] ,
    \Tile_X10Y12_W2BEGb[3] ,
    \Tile_X10Y12_W2BEGb[2] ,
    \Tile_X10Y12_W2BEGb[1] ,
    \Tile_X10Y12_W2BEGb[0] }),
    .W2MID({\Tile_X10Y12_W2BEG[7] ,
    \Tile_X10Y12_W2BEG[6] ,
    \Tile_X10Y12_W2BEG[5] ,
    \Tile_X10Y12_W2BEG[4] ,
    \Tile_X10Y12_W2BEG[3] ,
    \Tile_X10Y12_W2BEG[2] ,
    \Tile_X10Y12_W2BEG[1] ,
    \Tile_X10Y12_W2BEG[0] }),
    .W6BEG({\Tile_X9Y12_W6BEG[11] ,
    \Tile_X9Y12_W6BEG[10] ,
    \Tile_X9Y12_W6BEG[9] ,
    \Tile_X9Y12_W6BEG[8] ,
    \Tile_X9Y12_W6BEG[7] ,
    \Tile_X9Y12_W6BEG[6] ,
    \Tile_X9Y12_W6BEG[5] ,
    \Tile_X9Y12_W6BEG[4] ,
    \Tile_X9Y12_W6BEG[3] ,
    \Tile_X9Y12_W6BEG[2] ,
    \Tile_X9Y12_W6BEG[1] ,
    \Tile_X9Y12_W6BEG[0] }),
    .W6END({\Tile_X10Y12_W6BEG[11] ,
    \Tile_X10Y12_W6BEG[10] ,
    \Tile_X10Y12_W6BEG[9] ,
    \Tile_X10Y12_W6BEG[8] ,
    \Tile_X10Y12_W6BEG[7] ,
    \Tile_X10Y12_W6BEG[6] ,
    \Tile_X10Y12_W6BEG[5] ,
    \Tile_X10Y12_W6BEG[4] ,
    \Tile_X10Y12_W6BEG[3] ,
    \Tile_X10Y12_W6BEG[2] ,
    \Tile_X10Y12_W6BEG[1] ,
    \Tile_X10Y12_W6BEG[0] }),
    .WW4BEG({\Tile_X9Y12_WW4BEG[15] ,
    \Tile_X9Y12_WW4BEG[14] ,
    \Tile_X9Y12_WW4BEG[13] ,
    \Tile_X9Y12_WW4BEG[12] ,
    \Tile_X9Y12_WW4BEG[11] ,
    \Tile_X9Y12_WW4BEG[10] ,
    \Tile_X9Y12_WW4BEG[9] ,
    \Tile_X9Y12_WW4BEG[8] ,
    \Tile_X9Y12_WW4BEG[7] ,
    \Tile_X9Y12_WW4BEG[6] ,
    \Tile_X9Y12_WW4BEG[5] ,
    \Tile_X9Y12_WW4BEG[4] ,
    \Tile_X9Y12_WW4BEG[3] ,
    \Tile_X9Y12_WW4BEG[2] ,
    \Tile_X9Y12_WW4BEG[1] ,
    \Tile_X9Y12_WW4BEG[0] }),
    .WW4END({\Tile_X10Y12_WW4BEG[15] ,
    \Tile_X10Y12_WW4BEG[14] ,
    \Tile_X10Y12_WW4BEG[13] ,
    \Tile_X10Y12_WW4BEG[12] ,
    \Tile_X10Y12_WW4BEG[11] ,
    \Tile_X10Y12_WW4BEG[10] ,
    \Tile_X10Y12_WW4BEG[9] ,
    \Tile_X10Y12_WW4BEG[8] ,
    \Tile_X10Y12_WW4BEG[7] ,
    \Tile_X10Y12_WW4BEG[6] ,
    \Tile_X10Y12_WW4BEG[5] ,
    \Tile_X10Y12_WW4BEG[4] ,
    \Tile_X10Y12_WW4BEG[3] ,
    \Tile_X10Y12_WW4BEG[2] ,
    \Tile_X10Y12_WW4BEG[1] ,
    \Tile_X10Y12_WW4BEG[0] }));
 LUT4AB Tile_X9Y13_LUT4AB (.Ci(Tile_X9Y14_Co),
    .Co(Tile_X9Y13_Co),
    .UserCLK(Tile_X9Y14_UserCLKo),
    .UserCLKo(Tile_X9Y13_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X9Y13_E1BEG[3] ,
    \Tile_X9Y13_E1BEG[2] ,
    \Tile_X9Y13_E1BEG[1] ,
    \Tile_X9Y13_E1BEG[0] }),
    .E1END({\Tile_X8Y13_E1BEG[3] ,
    \Tile_X8Y13_E1BEG[2] ,
    \Tile_X8Y13_E1BEG[1] ,
    \Tile_X8Y13_E1BEG[0] }),
    .E2BEG({\Tile_X9Y13_E2BEG[7] ,
    \Tile_X9Y13_E2BEG[6] ,
    \Tile_X9Y13_E2BEG[5] ,
    \Tile_X9Y13_E2BEG[4] ,
    \Tile_X9Y13_E2BEG[3] ,
    \Tile_X9Y13_E2BEG[2] ,
    \Tile_X9Y13_E2BEG[1] ,
    \Tile_X9Y13_E2BEG[0] }),
    .E2BEGb({\Tile_X9Y13_E2BEGb[7] ,
    \Tile_X9Y13_E2BEGb[6] ,
    \Tile_X9Y13_E2BEGb[5] ,
    \Tile_X9Y13_E2BEGb[4] ,
    \Tile_X9Y13_E2BEGb[3] ,
    \Tile_X9Y13_E2BEGb[2] ,
    \Tile_X9Y13_E2BEGb[1] ,
    \Tile_X9Y13_E2BEGb[0] }),
    .E2END({\Tile_X8Y13_E2BEGb[7] ,
    \Tile_X8Y13_E2BEGb[6] ,
    \Tile_X8Y13_E2BEGb[5] ,
    \Tile_X8Y13_E2BEGb[4] ,
    \Tile_X8Y13_E2BEGb[3] ,
    \Tile_X8Y13_E2BEGb[2] ,
    \Tile_X8Y13_E2BEGb[1] ,
    \Tile_X8Y13_E2BEGb[0] }),
    .E2MID({\Tile_X8Y13_E2BEG[7] ,
    \Tile_X8Y13_E2BEG[6] ,
    \Tile_X8Y13_E2BEG[5] ,
    \Tile_X8Y13_E2BEG[4] ,
    \Tile_X8Y13_E2BEG[3] ,
    \Tile_X8Y13_E2BEG[2] ,
    \Tile_X8Y13_E2BEG[1] ,
    \Tile_X8Y13_E2BEG[0] }),
    .E6BEG({\Tile_X9Y13_E6BEG[11] ,
    \Tile_X9Y13_E6BEG[10] ,
    \Tile_X9Y13_E6BEG[9] ,
    \Tile_X9Y13_E6BEG[8] ,
    \Tile_X9Y13_E6BEG[7] ,
    \Tile_X9Y13_E6BEG[6] ,
    \Tile_X9Y13_E6BEG[5] ,
    \Tile_X9Y13_E6BEG[4] ,
    \Tile_X9Y13_E6BEG[3] ,
    \Tile_X9Y13_E6BEG[2] ,
    \Tile_X9Y13_E6BEG[1] ,
    \Tile_X9Y13_E6BEG[0] }),
    .E6END({\Tile_X8Y13_E6BEG[11] ,
    \Tile_X8Y13_E6BEG[10] ,
    \Tile_X8Y13_E6BEG[9] ,
    \Tile_X8Y13_E6BEG[8] ,
    \Tile_X8Y13_E6BEG[7] ,
    \Tile_X8Y13_E6BEG[6] ,
    \Tile_X8Y13_E6BEG[5] ,
    \Tile_X8Y13_E6BEG[4] ,
    \Tile_X8Y13_E6BEG[3] ,
    \Tile_X8Y13_E6BEG[2] ,
    \Tile_X8Y13_E6BEG[1] ,
    \Tile_X8Y13_E6BEG[0] }),
    .EE4BEG({\Tile_X9Y13_EE4BEG[15] ,
    \Tile_X9Y13_EE4BEG[14] ,
    \Tile_X9Y13_EE4BEG[13] ,
    \Tile_X9Y13_EE4BEG[12] ,
    \Tile_X9Y13_EE4BEG[11] ,
    \Tile_X9Y13_EE4BEG[10] ,
    \Tile_X9Y13_EE4BEG[9] ,
    \Tile_X9Y13_EE4BEG[8] ,
    \Tile_X9Y13_EE4BEG[7] ,
    \Tile_X9Y13_EE4BEG[6] ,
    \Tile_X9Y13_EE4BEG[5] ,
    \Tile_X9Y13_EE4BEG[4] ,
    \Tile_X9Y13_EE4BEG[3] ,
    \Tile_X9Y13_EE4BEG[2] ,
    \Tile_X9Y13_EE4BEG[1] ,
    \Tile_X9Y13_EE4BEG[0] }),
    .EE4END({\Tile_X8Y13_EE4BEG[15] ,
    \Tile_X8Y13_EE4BEG[14] ,
    \Tile_X8Y13_EE4BEG[13] ,
    \Tile_X8Y13_EE4BEG[12] ,
    \Tile_X8Y13_EE4BEG[11] ,
    \Tile_X8Y13_EE4BEG[10] ,
    \Tile_X8Y13_EE4BEG[9] ,
    \Tile_X8Y13_EE4BEG[8] ,
    \Tile_X8Y13_EE4BEG[7] ,
    \Tile_X8Y13_EE4BEG[6] ,
    \Tile_X8Y13_EE4BEG[5] ,
    \Tile_X8Y13_EE4BEG[4] ,
    \Tile_X8Y13_EE4BEG[3] ,
    \Tile_X8Y13_EE4BEG[2] ,
    \Tile_X8Y13_EE4BEG[1] ,
    \Tile_X8Y13_EE4BEG[0] }),
    .FrameData({\Tile_X8Y13_FrameData_O[31] ,
    \Tile_X8Y13_FrameData_O[30] ,
    \Tile_X8Y13_FrameData_O[29] ,
    \Tile_X8Y13_FrameData_O[28] ,
    \Tile_X8Y13_FrameData_O[27] ,
    \Tile_X8Y13_FrameData_O[26] ,
    \Tile_X8Y13_FrameData_O[25] ,
    \Tile_X8Y13_FrameData_O[24] ,
    \Tile_X8Y13_FrameData_O[23] ,
    \Tile_X8Y13_FrameData_O[22] ,
    \Tile_X8Y13_FrameData_O[21] ,
    \Tile_X8Y13_FrameData_O[20] ,
    \Tile_X8Y13_FrameData_O[19] ,
    \Tile_X8Y13_FrameData_O[18] ,
    \Tile_X8Y13_FrameData_O[17] ,
    \Tile_X8Y13_FrameData_O[16] ,
    \Tile_X8Y13_FrameData_O[15] ,
    \Tile_X8Y13_FrameData_O[14] ,
    \Tile_X8Y13_FrameData_O[13] ,
    \Tile_X8Y13_FrameData_O[12] ,
    \Tile_X8Y13_FrameData_O[11] ,
    \Tile_X8Y13_FrameData_O[10] ,
    \Tile_X8Y13_FrameData_O[9] ,
    \Tile_X8Y13_FrameData_O[8] ,
    \Tile_X8Y13_FrameData_O[7] ,
    \Tile_X8Y13_FrameData_O[6] ,
    \Tile_X8Y13_FrameData_O[5] ,
    \Tile_X8Y13_FrameData_O[4] ,
    \Tile_X8Y13_FrameData_O[3] ,
    \Tile_X8Y13_FrameData_O[2] ,
    \Tile_X8Y13_FrameData_O[1] ,
    \Tile_X8Y13_FrameData_O[0] }),
    .FrameData_O({\Tile_X9Y13_FrameData_O[31] ,
    \Tile_X9Y13_FrameData_O[30] ,
    \Tile_X9Y13_FrameData_O[29] ,
    \Tile_X9Y13_FrameData_O[28] ,
    \Tile_X9Y13_FrameData_O[27] ,
    \Tile_X9Y13_FrameData_O[26] ,
    \Tile_X9Y13_FrameData_O[25] ,
    \Tile_X9Y13_FrameData_O[24] ,
    \Tile_X9Y13_FrameData_O[23] ,
    \Tile_X9Y13_FrameData_O[22] ,
    \Tile_X9Y13_FrameData_O[21] ,
    \Tile_X9Y13_FrameData_O[20] ,
    \Tile_X9Y13_FrameData_O[19] ,
    \Tile_X9Y13_FrameData_O[18] ,
    \Tile_X9Y13_FrameData_O[17] ,
    \Tile_X9Y13_FrameData_O[16] ,
    \Tile_X9Y13_FrameData_O[15] ,
    \Tile_X9Y13_FrameData_O[14] ,
    \Tile_X9Y13_FrameData_O[13] ,
    \Tile_X9Y13_FrameData_O[12] ,
    \Tile_X9Y13_FrameData_O[11] ,
    \Tile_X9Y13_FrameData_O[10] ,
    \Tile_X9Y13_FrameData_O[9] ,
    \Tile_X9Y13_FrameData_O[8] ,
    \Tile_X9Y13_FrameData_O[7] ,
    \Tile_X9Y13_FrameData_O[6] ,
    \Tile_X9Y13_FrameData_O[5] ,
    \Tile_X9Y13_FrameData_O[4] ,
    \Tile_X9Y13_FrameData_O[3] ,
    \Tile_X9Y13_FrameData_O[2] ,
    \Tile_X9Y13_FrameData_O[1] ,
    \Tile_X9Y13_FrameData_O[0] }),
    .FrameStrobe({\Tile_X9Y14_FrameStrobe_O[19] ,
    \Tile_X9Y14_FrameStrobe_O[18] ,
    \Tile_X9Y14_FrameStrobe_O[17] ,
    \Tile_X9Y14_FrameStrobe_O[16] ,
    \Tile_X9Y14_FrameStrobe_O[15] ,
    \Tile_X9Y14_FrameStrobe_O[14] ,
    \Tile_X9Y14_FrameStrobe_O[13] ,
    \Tile_X9Y14_FrameStrobe_O[12] ,
    \Tile_X9Y14_FrameStrobe_O[11] ,
    \Tile_X9Y14_FrameStrobe_O[10] ,
    \Tile_X9Y14_FrameStrobe_O[9] ,
    \Tile_X9Y14_FrameStrobe_O[8] ,
    \Tile_X9Y14_FrameStrobe_O[7] ,
    \Tile_X9Y14_FrameStrobe_O[6] ,
    \Tile_X9Y14_FrameStrobe_O[5] ,
    \Tile_X9Y14_FrameStrobe_O[4] ,
    \Tile_X9Y14_FrameStrobe_O[3] ,
    \Tile_X9Y14_FrameStrobe_O[2] ,
    \Tile_X9Y14_FrameStrobe_O[1] ,
    \Tile_X9Y14_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X9Y13_FrameStrobe_O[19] ,
    \Tile_X9Y13_FrameStrobe_O[18] ,
    \Tile_X9Y13_FrameStrobe_O[17] ,
    \Tile_X9Y13_FrameStrobe_O[16] ,
    \Tile_X9Y13_FrameStrobe_O[15] ,
    \Tile_X9Y13_FrameStrobe_O[14] ,
    \Tile_X9Y13_FrameStrobe_O[13] ,
    \Tile_X9Y13_FrameStrobe_O[12] ,
    \Tile_X9Y13_FrameStrobe_O[11] ,
    \Tile_X9Y13_FrameStrobe_O[10] ,
    \Tile_X9Y13_FrameStrobe_O[9] ,
    \Tile_X9Y13_FrameStrobe_O[8] ,
    \Tile_X9Y13_FrameStrobe_O[7] ,
    \Tile_X9Y13_FrameStrobe_O[6] ,
    \Tile_X9Y13_FrameStrobe_O[5] ,
    \Tile_X9Y13_FrameStrobe_O[4] ,
    \Tile_X9Y13_FrameStrobe_O[3] ,
    \Tile_X9Y13_FrameStrobe_O[2] ,
    \Tile_X9Y13_FrameStrobe_O[1] ,
    \Tile_X9Y13_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X9Y13_N1BEG[3] ,
    \Tile_X9Y13_N1BEG[2] ,
    \Tile_X9Y13_N1BEG[1] ,
    \Tile_X9Y13_N1BEG[0] }),
    .N1END({\Tile_X9Y14_N1BEG[3] ,
    \Tile_X9Y14_N1BEG[2] ,
    \Tile_X9Y14_N1BEG[1] ,
    \Tile_X9Y14_N1BEG[0] }),
    .N2BEG({\Tile_X9Y13_N2BEG[7] ,
    \Tile_X9Y13_N2BEG[6] ,
    \Tile_X9Y13_N2BEG[5] ,
    \Tile_X9Y13_N2BEG[4] ,
    \Tile_X9Y13_N2BEG[3] ,
    \Tile_X9Y13_N2BEG[2] ,
    \Tile_X9Y13_N2BEG[1] ,
    \Tile_X9Y13_N2BEG[0] }),
    .N2BEGb({\Tile_X9Y13_N2BEGb[7] ,
    \Tile_X9Y13_N2BEGb[6] ,
    \Tile_X9Y13_N2BEGb[5] ,
    \Tile_X9Y13_N2BEGb[4] ,
    \Tile_X9Y13_N2BEGb[3] ,
    \Tile_X9Y13_N2BEGb[2] ,
    \Tile_X9Y13_N2BEGb[1] ,
    \Tile_X9Y13_N2BEGb[0] }),
    .N2END({\Tile_X9Y14_N2BEGb[7] ,
    \Tile_X9Y14_N2BEGb[6] ,
    \Tile_X9Y14_N2BEGb[5] ,
    \Tile_X9Y14_N2BEGb[4] ,
    \Tile_X9Y14_N2BEGb[3] ,
    \Tile_X9Y14_N2BEGb[2] ,
    \Tile_X9Y14_N2BEGb[1] ,
    \Tile_X9Y14_N2BEGb[0] }),
    .N2MID({\Tile_X9Y14_N2BEG[7] ,
    \Tile_X9Y14_N2BEG[6] ,
    \Tile_X9Y14_N2BEG[5] ,
    \Tile_X9Y14_N2BEG[4] ,
    \Tile_X9Y14_N2BEG[3] ,
    \Tile_X9Y14_N2BEG[2] ,
    \Tile_X9Y14_N2BEG[1] ,
    \Tile_X9Y14_N2BEG[0] }),
    .N4BEG({\Tile_X9Y13_N4BEG[15] ,
    \Tile_X9Y13_N4BEG[14] ,
    \Tile_X9Y13_N4BEG[13] ,
    \Tile_X9Y13_N4BEG[12] ,
    \Tile_X9Y13_N4BEG[11] ,
    \Tile_X9Y13_N4BEG[10] ,
    \Tile_X9Y13_N4BEG[9] ,
    \Tile_X9Y13_N4BEG[8] ,
    \Tile_X9Y13_N4BEG[7] ,
    \Tile_X9Y13_N4BEG[6] ,
    \Tile_X9Y13_N4BEG[5] ,
    \Tile_X9Y13_N4BEG[4] ,
    \Tile_X9Y13_N4BEG[3] ,
    \Tile_X9Y13_N4BEG[2] ,
    \Tile_X9Y13_N4BEG[1] ,
    \Tile_X9Y13_N4BEG[0] }),
    .N4END({\Tile_X9Y14_N4BEG[15] ,
    \Tile_X9Y14_N4BEG[14] ,
    \Tile_X9Y14_N4BEG[13] ,
    \Tile_X9Y14_N4BEG[12] ,
    \Tile_X9Y14_N4BEG[11] ,
    \Tile_X9Y14_N4BEG[10] ,
    \Tile_X9Y14_N4BEG[9] ,
    \Tile_X9Y14_N4BEG[8] ,
    \Tile_X9Y14_N4BEG[7] ,
    \Tile_X9Y14_N4BEG[6] ,
    \Tile_X9Y14_N4BEG[5] ,
    \Tile_X9Y14_N4BEG[4] ,
    \Tile_X9Y14_N4BEG[3] ,
    \Tile_X9Y14_N4BEG[2] ,
    \Tile_X9Y14_N4BEG[1] ,
    \Tile_X9Y14_N4BEG[0] }),
    .NN4BEG({\Tile_X9Y13_NN4BEG[15] ,
    \Tile_X9Y13_NN4BEG[14] ,
    \Tile_X9Y13_NN4BEG[13] ,
    \Tile_X9Y13_NN4BEG[12] ,
    \Tile_X9Y13_NN4BEG[11] ,
    \Tile_X9Y13_NN4BEG[10] ,
    \Tile_X9Y13_NN4BEG[9] ,
    \Tile_X9Y13_NN4BEG[8] ,
    \Tile_X9Y13_NN4BEG[7] ,
    \Tile_X9Y13_NN4BEG[6] ,
    \Tile_X9Y13_NN4BEG[5] ,
    \Tile_X9Y13_NN4BEG[4] ,
    \Tile_X9Y13_NN4BEG[3] ,
    \Tile_X9Y13_NN4BEG[2] ,
    \Tile_X9Y13_NN4BEG[1] ,
    \Tile_X9Y13_NN4BEG[0] }),
    .NN4END({\Tile_X9Y14_NN4BEG[15] ,
    \Tile_X9Y14_NN4BEG[14] ,
    \Tile_X9Y14_NN4BEG[13] ,
    \Tile_X9Y14_NN4BEG[12] ,
    \Tile_X9Y14_NN4BEG[11] ,
    \Tile_X9Y14_NN4BEG[10] ,
    \Tile_X9Y14_NN4BEG[9] ,
    \Tile_X9Y14_NN4BEG[8] ,
    \Tile_X9Y14_NN4BEG[7] ,
    \Tile_X9Y14_NN4BEG[6] ,
    \Tile_X9Y14_NN4BEG[5] ,
    \Tile_X9Y14_NN4BEG[4] ,
    \Tile_X9Y14_NN4BEG[3] ,
    \Tile_X9Y14_NN4BEG[2] ,
    \Tile_X9Y14_NN4BEG[1] ,
    \Tile_X9Y14_NN4BEG[0] }),
    .S1BEG({\Tile_X9Y13_S1BEG[3] ,
    \Tile_X9Y13_S1BEG[2] ,
    \Tile_X9Y13_S1BEG[1] ,
    \Tile_X9Y13_S1BEG[0] }),
    .S1END({\Tile_X9Y12_S1BEG[3] ,
    \Tile_X9Y12_S1BEG[2] ,
    \Tile_X9Y12_S1BEG[1] ,
    \Tile_X9Y12_S1BEG[0] }),
    .S2BEG({\Tile_X9Y13_S2BEG[7] ,
    \Tile_X9Y13_S2BEG[6] ,
    \Tile_X9Y13_S2BEG[5] ,
    \Tile_X9Y13_S2BEG[4] ,
    \Tile_X9Y13_S2BEG[3] ,
    \Tile_X9Y13_S2BEG[2] ,
    \Tile_X9Y13_S2BEG[1] ,
    \Tile_X9Y13_S2BEG[0] }),
    .S2BEGb({\Tile_X9Y13_S2BEGb[7] ,
    \Tile_X9Y13_S2BEGb[6] ,
    \Tile_X9Y13_S2BEGb[5] ,
    \Tile_X9Y13_S2BEGb[4] ,
    \Tile_X9Y13_S2BEGb[3] ,
    \Tile_X9Y13_S2BEGb[2] ,
    \Tile_X9Y13_S2BEGb[1] ,
    \Tile_X9Y13_S2BEGb[0] }),
    .S2END({\Tile_X9Y12_S2BEGb[7] ,
    \Tile_X9Y12_S2BEGb[6] ,
    \Tile_X9Y12_S2BEGb[5] ,
    \Tile_X9Y12_S2BEGb[4] ,
    \Tile_X9Y12_S2BEGb[3] ,
    \Tile_X9Y12_S2BEGb[2] ,
    \Tile_X9Y12_S2BEGb[1] ,
    \Tile_X9Y12_S2BEGb[0] }),
    .S2MID({\Tile_X9Y12_S2BEG[7] ,
    \Tile_X9Y12_S2BEG[6] ,
    \Tile_X9Y12_S2BEG[5] ,
    \Tile_X9Y12_S2BEG[4] ,
    \Tile_X9Y12_S2BEG[3] ,
    \Tile_X9Y12_S2BEG[2] ,
    \Tile_X9Y12_S2BEG[1] ,
    \Tile_X9Y12_S2BEG[0] }),
    .S4BEG({\Tile_X9Y13_S4BEG[15] ,
    \Tile_X9Y13_S4BEG[14] ,
    \Tile_X9Y13_S4BEG[13] ,
    \Tile_X9Y13_S4BEG[12] ,
    \Tile_X9Y13_S4BEG[11] ,
    \Tile_X9Y13_S4BEG[10] ,
    \Tile_X9Y13_S4BEG[9] ,
    \Tile_X9Y13_S4BEG[8] ,
    \Tile_X9Y13_S4BEG[7] ,
    \Tile_X9Y13_S4BEG[6] ,
    \Tile_X9Y13_S4BEG[5] ,
    \Tile_X9Y13_S4BEG[4] ,
    \Tile_X9Y13_S4BEG[3] ,
    \Tile_X9Y13_S4BEG[2] ,
    \Tile_X9Y13_S4BEG[1] ,
    \Tile_X9Y13_S4BEG[0] }),
    .S4END({\Tile_X9Y12_S4BEG[15] ,
    \Tile_X9Y12_S4BEG[14] ,
    \Tile_X9Y12_S4BEG[13] ,
    \Tile_X9Y12_S4BEG[12] ,
    \Tile_X9Y12_S4BEG[11] ,
    \Tile_X9Y12_S4BEG[10] ,
    \Tile_X9Y12_S4BEG[9] ,
    \Tile_X9Y12_S4BEG[8] ,
    \Tile_X9Y12_S4BEG[7] ,
    \Tile_X9Y12_S4BEG[6] ,
    \Tile_X9Y12_S4BEG[5] ,
    \Tile_X9Y12_S4BEG[4] ,
    \Tile_X9Y12_S4BEG[3] ,
    \Tile_X9Y12_S4BEG[2] ,
    \Tile_X9Y12_S4BEG[1] ,
    \Tile_X9Y12_S4BEG[0] }),
    .SS4BEG({\Tile_X9Y13_SS4BEG[15] ,
    \Tile_X9Y13_SS4BEG[14] ,
    \Tile_X9Y13_SS4BEG[13] ,
    \Tile_X9Y13_SS4BEG[12] ,
    \Tile_X9Y13_SS4BEG[11] ,
    \Tile_X9Y13_SS4BEG[10] ,
    \Tile_X9Y13_SS4BEG[9] ,
    \Tile_X9Y13_SS4BEG[8] ,
    \Tile_X9Y13_SS4BEG[7] ,
    \Tile_X9Y13_SS4BEG[6] ,
    \Tile_X9Y13_SS4BEG[5] ,
    \Tile_X9Y13_SS4BEG[4] ,
    \Tile_X9Y13_SS4BEG[3] ,
    \Tile_X9Y13_SS4BEG[2] ,
    \Tile_X9Y13_SS4BEG[1] ,
    \Tile_X9Y13_SS4BEG[0] }),
    .SS4END({\Tile_X9Y12_SS4BEG[15] ,
    \Tile_X9Y12_SS4BEG[14] ,
    \Tile_X9Y12_SS4BEG[13] ,
    \Tile_X9Y12_SS4BEG[12] ,
    \Tile_X9Y12_SS4BEG[11] ,
    \Tile_X9Y12_SS4BEG[10] ,
    \Tile_X9Y12_SS4BEG[9] ,
    \Tile_X9Y12_SS4BEG[8] ,
    \Tile_X9Y12_SS4BEG[7] ,
    \Tile_X9Y12_SS4BEG[6] ,
    \Tile_X9Y12_SS4BEG[5] ,
    \Tile_X9Y12_SS4BEG[4] ,
    \Tile_X9Y12_SS4BEG[3] ,
    \Tile_X9Y12_SS4BEG[2] ,
    \Tile_X9Y12_SS4BEG[1] ,
    \Tile_X9Y12_SS4BEG[0] }),
    .W1BEG({\Tile_X9Y13_W1BEG[3] ,
    \Tile_X9Y13_W1BEG[2] ,
    \Tile_X9Y13_W1BEG[1] ,
    \Tile_X9Y13_W1BEG[0] }),
    .W1END({\Tile_X10Y13_W1BEG[3] ,
    \Tile_X10Y13_W1BEG[2] ,
    \Tile_X10Y13_W1BEG[1] ,
    \Tile_X10Y13_W1BEG[0] }),
    .W2BEG({\Tile_X9Y13_W2BEG[7] ,
    \Tile_X9Y13_W2BEG[6] ,
    \Tile_X9Y13_W2BEG[5] ,
    \Tile_X9Y13_W2BEG[4] ,
    \Tile_X9Y13_W2BEG[3] ,
    \Tile_X9Y13_W2BEG[2] ,
    \Tile_X9Y13_W2BEG[1] ,
    \Tile_X9Y13_W2BEG[0] }),
    .W2BEGb({\Tile_X9Y13_W2BEGb[7] ,
    \Tile_X9Y13_W2BEGb[6] ,
    \Tile_X9Y13_W2BEGb[5] ,
    \Tile_X9Y13_W2BEGb[4] ,
    \Tile_X9Y13_W2BEGb[3] ,
    \Tile_X9Y13_W2BEGb[2] ,
    \Tile_X9Y13_W2BEGb[1] ,
    \Tile_X9Y13_W2BEGb[0] }),
    .W2END({\Tile_X10Y13_W2BEGb[7] ,
    \Tile_X10Y13_W2BEGb[6] ,
    \Tile_X10Y13_W2BEGb[5] ,
    \Tile_X10Y13_W2BEGb[4] ,
    \Tile_X10Y13_W2BEGb[3] ,
    \Tile_X10Y13_W2BEGb[2] ,
    \Tile_X10Y13_W2BEGb[1] ,
    \Tile_X10Y13_W2BEGb[0] }),
    .W2MID({\Tile_X10Y13_W2BEG[7] ,
    \Tile_X10Y13_W2BEG[6] ,
    \Tile_X10Y13_W2BEG[5] ,
    \Tile_X10Y13_W2BEG[4] ,
    \Tile_X10Y13_W2BEG[3] ,
    \Tile_X10Y13_W2BEG[2] ,
    \Tile_X10Y13_W2BEG[1] ,
    \Tile_X10Y13_W2BEG[0] }),
    .W6BEG({\Tile_X9Y13_W6BEG[11] ,
    \Tile_X9Y13_W6BEG[10] ,
    \Tile_X9Y13_W6BEG[9] ,
    \Tile_X9Y13_W6BEG[8] ,
    \Tile_X9Y13_W6BEG[7] ,
    \Tile_X9Y13_W6BEG[6] ,
    \Tile_X9Y13_W6BEG[5] ,
    \Tile_X9Y13_W6BEG[4] ,
    \Tile_X9Y13_W6BEG[3] ,
    \Tile_X9Y13_W6BEG[2] ,
    \Tile_X9Y13_W6BEG[1] ,
    \Tile_X9Y13_W6BEG[0] }),
    .W6END({\Tile_X10Y13_W6BEG[11] ,
    \Tile_X10Y13_W6BEG[10] ,
    \Tile_X10Y13_W6BEG[9] ,
    \Tile_X10Y13_W6BEG[8] ,
    \Tile_X10Y13_W6BEG[7] ,
    \Tile_X10Y13_W6BEG[6] ,
    \Tile_X10Y13_W6BEG[5] ,
    \Tile_X10Y13_W6BEG[4] ,
    \Tile_X10Y13_W6BEG[3] ,
    \Tile_X10Y13_W6BEG[2] ,
    \Tile_X10Y13_W6BEG[1] ,
    \Tile_X10Y13_W6BEG[0] }),
    .WW4BEG({\Tile_X9Y13_WW4BEG[15] ,
    \Tile_X9Y13_WW4BEG[14] ,
    \Tile_X9Y13_WW4BEG[13] ,
    \Tile_X9Y13_WW4BEG[12] ,
    \Tile_X9Y13_WW4BEG[11] ,
    \Tile_X9Y13_WW4BEG[10] ,
    \Tile_X9Y13_WW4BEG[9] ,
    \Tile_X9Y13_WW4BEG[8] ,
    \Tile_X9Y13_WW4BEG[7] ,
    \Tile_X9Y13_WW4BEG[6] ,
    \Tile_X9Y13_WW4BEG[5] ,
    \Tile_X9Y13_WW4BEG[4] ,
    \Tile_X9Y13_WW4BEG[3] ,
    \Tile_X9Y13_WW4BEG[2] ,
    \Tile_X9Y13_WW4BEG[1] ,
    \Tile_X9Y13_WW4BEG[0] }),
    .WW4END({\Tile_X10Y13_WW4BEG[15] ,
    \Tile_X10Y13_WW4BEG[14] ,
    \Tile_X10Y13_WW4BEG[13] ,
    \Tile_X10Y13_WW4BEG[12] ,
    \Tile_X10Y13_WW4BEG[11] ,
    \Tile_X10Y13_WW4BEG[10] ,
    \Tile_X10Y13_WW4BEG[9] ,
    \Tile_X10Y13_WW4BEG[8] ,
    \Tile_X10Y13_WW4BEG[7] ,
    \Tile_X10Y13_WW4BEG[6] ,
    \Tile_X10Y13_WW4BEG[5] ,
    \Tile_X10Y13_WW4BEG[4] ,
    \Tile_X10Y13_WW4BEG[3] ,
    \Tile_X10Y13_WW4BEG[2] ,
    \Tile_X10Y13_WW4BEG[1] ,
    \Tile_X10Y13_WW4BEG[0] }));
 LUT4AB Tile_X9Y14_LUT4AB (.Ci(Tile_X9Y15_Co),
    .Co(Tile_X9Y14_Co),
    .UserCLK(Tile_X9Y15_UserCLKo),
    .UserCLKo(Tile_X9Y14_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X9Y14_E1BEG[3] ,
    \Tile_X9Y14_E1BEG[2] ,
    \Tile_X9Y14_E1BEG[1] ,
    \Tile_X9Y14_E1BEG[0] }),
    .E1END({\Tile_X8Y14_E1BEG[3] ,
    \Tile_X8Y14_E1BEG[2] ,
    \Tile_X8Y14_E1BEG[1] ,
    \Tile_X8Y14_E1BEG[0] }),
    .E2BEG({\Tile_X9Y14_E2BEG[7] ,
    \Tile_X9Y14_E2BEG[6] ,
    \Tile_X9Y14_E2BEG[5] ,
    \Tile_X9Y14_E2BEG[4] ,
    \Tile_X9Y14_E2BEG[3] ,
    \Tile_X9Y14_E2BEG[2] ,
    \Tile_X9Y14_E2BEG[1] ,
    \Tile_X9Y14_E2BEG[0] }),
    .E2BEGb({\Tile_X9Y14_E2BEGb[7] ,
    \Tile_X9Y14_E2BEGb[6] ,
    \Tile_X9Y14_E2BEGb[5] ,
    \Tile_X9Y14_E2BEGb[4] ,
    \Tile_X9Y14_E2BEGb[3] ,
    \Tile_X9Y14_E2BEGb[2] ,
    \Tile_X9Y14_E2BEGb[1] ,
    \Tile_X9Y14_E2BEGb[0] }),
    .E2END({\Tile_X8Y14_E2BEGb[7] ,
    \Tile_X8Y14_E2BEGb[6] ,
    \Tile_X8Y14_E2BEGb[5] ,
    \Tile_X8Y14_E2BEGb[4] ,
    \Tile_X8Y14_E2BEGb[3] ,
    \Tile_X8Y14_E2BEGb[2] ,
    \Tile_X8Y14_E2BEGb[1] ,
    \Tile_X8Y14_E2BEGb[0] }),
    .E2MID({\Tile_X8Y14_E2BEG[7] ,
    \Tile_X8Y14_E2BEG[6] ,
    \Tile_X8Y14_E2BEG[5] ,
    \Tile_X8Y14_E2BEG[4] ,
    \Tile_X8Y14_E2BEG[3] ,
    \Tile_X8Y14_E2BEG[2] ,
    \Tile_X8Y14_E2BEG[1] ,
    \Tile_X8Y14_E2BEG[0] }),
    .E6BEG({\Tile_X9Y14_E6BEG[11] ,
    \Tile_X9Y14_E6BEG[10] ,
    \Tile_X9Y14_E6BEG[9] ,
    \Tile_X9Y14_E6BEG[8] ,
    \Tile_X9Y14_E6BEG[7] ,
    \Tile_X9Y14_E6BEG[6] ,
    \Tile_X9Y14_E6BEG[5] ,
    \Tile_X9Y14_E6BEG[4] ,
    \Tile_X9Y14_E6BEG[3] ,
    \Tile_X9Y14_E6BEG[2] ,
    \Tile_X9Y14_E6BEG[1] ,
    \Tile_X9Y14_E6BEG[0] }),
    .E6END({\Tile_X8Y14_E6BEG[11] ,
    \Tile_X8Y14_E6BEG[10] ,
    \Tile_X8Y14_E6BEG[9] ,
    \Tile_X8Y14_E6BEG[8] ,
    \Tile_X8Y14_E6BEG[7] ,
    \Tile_X8Y14_E6BEG[6] ,
    \Tile_X8Y14_E6BEG[5] ,
    \Tile_X8Y14_E6BEG[4] ,
    \Tile_X8Y14_E6BEG[3] ,
    \Tile_X8Y14_E6BEG[2] ,
    \Tile_X8Y14_E6BEG[1] ,
    \Tile_X8Y14_E6BEG[0] }),
    .EE4BEG({\Tile_X9Y14_EE4BEG[15] ,
    \Tile_X9Y14_EE4BEG[14] ,
    \Tile_X9Y14_EE4BEG[13] ,
    \Tile_X9Y14_EE4BEG[12] ,
    \Tile_X9Y14_EE4BEG[11] ,
    \Tile_X9Y14_EE4BEG[10] ,
    \Tile_X9Y14_EE4BEG[9] ,
    \Tile_X9Y14_EE4BEG[8] ,
    \Tile_X9Y14_EE4BEG[7] ,
    \Tile_X9Y14_EE4BEG[6] ,
    \Tile_X9Y14_EE4BEG[5] ,
    \Tile_X9Y14_EE4BEG[4] ,
    \Tile_X9Y14_EE4BEG[3] ,
    \Tile_X9Y14_EE4BEG[2] ,
    \Tile_X9Y14_EE4BEG[1] ,
    \Tile_X9Y14_EE4BEG[0] }),
    .EE4END({\Tile_X8Y14_EE4BEG[15] ,
    \Tile_X8Y14_EE4BEG[14] ,
    \Tile_X8Y14_EE4BEG[13] ,
    \Tile_X8Y14_EE4BEG[12] ,
    \Tile_X8Y14_EE4BEG[11] ,
    \Tile_X8Y14_EE4BEG[10] ,
    \Tile_X8Y14_EE4BEG[9] ,
    \Tile_X8Y14_EE4BEG[8] ,
    \Tile_X8Y14_EE4BEG[7] ,
    \Tile_X8Y14_EE4BEG[6] ,
    \Tile_X8Y14_EE4BEG[5] ,
    \Tile_X8Y14_EE4BEG[4] ,
    \Tile_X8Y14_EE4BEG[3] ,
    \Tile_X8Y14_EE4BEG[2] ,
    \Tile_X8Y14_EE4BEG[1] ,
    \Tile_X8Y14_EE4BEG[0] }),
    .FrameData({\Tile_X8Y14_FrameData_O[31] ,
    \Tile_X8Y14_FrameData_O[30] ,
    \Tile_X8Y14_FrameData_O[29] ,
    \Tile_X8Y14_FrameData_O[28] ,
    \Tile_X8Y14_FrameData_O[27] ,
    \Tile_X8Y14_FrameData_O[26] ,
    \Tile_X8Y14_FrameData_O[25] ,
    \Tile_X8Y14_FrameData_O[24] ,
    \Tile_X8Y14_FrameData_O[23] ,
    \Tile_X8Y14_FrameData_O[22] ,
    \Tile_X8Y14_FrameData_O[21] ,
    \Tile_X8Y14_FrameData_O[20] ,
    \Tile_X8Y14_FrameData_O[19] ,
    \Tile_X8Y14_FrameData_O[18] ,
    \Tile_X8Y14_FrameData_O[17] ,
    \Tile_X8Y14_FrameData_O[16] ,
    \Tile_X8Y14_FrameData_O[15] ,
    \Tile_X8Y14_FrameData_O[14] ,
    \Tile_X8Y14_FrameData_O[13] ,
    \Tile_X8Y14_FrameData_O[12] ,
    \Tile_X8Y14_FrameData_O[11] ,
    \Tile_X8Y14_FrameData_O[10] ,
    \Tile_X8Y14_FrameData_O[9] ,
    \Tile_X8Y14_FrameData_O[8] ,
    \Tile_X8Y14_FrameData_O[7] ,
    \Tile_X8Y14_FrameData_O[6] ,
    \Tile_X8Y14_FrameData_O[5] ,
    \Tile_X8Y14_FrameData_O[4] ,
    \Tile_X8Y14_FrameData_O[3] ,
    \Tile_X8Y14_FrameData_O[2] ,
    \Tile_X8Y14_FrameData_O[1] ,
    \Tile_X8Y14_FrameData_O[0] }),
    .FrameData_O({\Tile_X9Y14_FrameData_O[31] ,
    \Tile_X9Y14_FrameData_O[30] ,
    \Tile_X9Y14_FrameData_O[29] ,
    \Tile_X9Y14_FrameData_O[28] ,
    \Tile_X9Y14_FrameData_O[27] ,
    \Tile_X9Y14_FrameData_O[26] ,
    \Tile_X9Y14_FrameData_O[25] ,
    \Tile_X9Y14_FrameData_O[24] ,
    \Tile_X9Y14_FrameData_O[23] ,
    \Tile_X9Y14_FrameData_O[22] ,
    \Tile_X9Y14_FrameData_O[21] ,
    \Tile_X9Y14_FrameData_O[20] ,
    \Tile_X9Y14_FrameData_O[19] ,
    \Tile_X9Y14_FrameData_O[18] ,
    \Tile_X9Y14_FrameData_O[17] ,
    \Tile_X9Y14_FrameData_O[16] ,
    \Tile_X9Y14_FrameData_O[15] ,
    \Tile_X9Y14_FrameData_O[14] ,
    \Tile_X9Y14_FrameData_O[13] ,
    \Tile_X9Y14_FrameData_O[12] ,
    \Tile_X9Y14_FrameData_O[11] ,
    \Tile_X9Y14_FrameData_O[10] ,
    \Tile_X9Y14_FrameData_O[9] ,
    \Tile_X9Y14_FrameData_O[8] ,
    \Tile_X9Y14_FrameData_O[7] ,
    \Tile_X9Y14_FrameData_O[6] ,
    \Tile_X9Y14_FrameData_O[5] ,
    \Tile_X9Y14_FrameData_O[4] ,
    \Tile_X9Y14_FrameData_O[3] ,
    \Tile_X9Y14_FrameData_O[2] ,
    \Tile_X9Y14_FrameData_O[1] ,
    \Tile_X9Y14_FrameData_O[0] }),
    .FrameStrobe({\Tile_X9Y15_FrameStrobe_O[19] ,
    \Tile_X9Y15_FrameStrobe_O[18] ,
    \Tile_X9Y15_FrameStrobe_O[17] ,
    \Tile_X9Y15_FrameStrobe_O[16] ,
    \Tile_X9Y15_FrameStrobe_O[15] ,
    \Tile_X9Y15_FrameStrobe_O[14] ,
    \Tile_X9Y15_FrameStrobe_O[13] ,
    \Tile_X9Y15_FrameStrobe_O[12] ,
    \Tile_X9Y15_FrameStrobe_O[11] ,
    \Tile_X9Y15_FrameStrobe_O[10] ,
    \Tile_X9Y15_FrameStrobe_O[9] ,
    \Tile_X9Y15_FrameStrobe_O[8] ,
    \Tile_X9Y15_FrameStrobe_O[7] ,
    \Tile_X9Y15_FrameStrobe_O[6] ,
    \Tile_X9Y15_FrameStrobe_O[5] ,
    \Tile_X9Y15_FrameStrobe_O[4] ,
    \Tile_X9Y15_FrameStrobe_O[3] ,
    \Tile_X9Y15_FrameStrobe_O[2] ,
    \Tile_X9Y15_FrameStrobe_O[1] ,
    \Tile_X9Y15_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X9Y14_FrameStrobe_O[19] ,
    \Tile_X9Y14_FrameStrobe_O[18] ,
    \Tile_X9Y14_FrameStrobe_O[17] ,
    \Tile_X9Y14_FrameStrobe_O[16] ,
    \Tile_X9Y14_FrameStrobe_O[15] ,
    \Tile_X9Y14_FrameStrobe_O[14] ,
    \Tile_X9Y14_FrameStrobe_O[13] ,
    \Tile_X9Y14_FrameStrobe_O[12] ,
    \Tile_X9Y14_FrameStrobe_O[11] ,
    \Tile_X9Y14_FrameStrobe_O[10] ,
    \Tile_X9Y14_FrameStrobe_O[9] ,
    \Tile_X9Y14_FrameStrobe_O[8] ,
    \Tile_X9Y14_FrameStrobe_O[7] ,
    \Tile_X9Y14_FrameStrobe_O[6] ,
    \Tile_X9Y14_FrameStrobe_O[5] ,
    \Tile_X9Y14_FrameStrobe_O[4] ,
    \Tile_X9Y14_FrameStrobe_O[3] ,
    \Tile_X9Y14_FrameStrobe_O[2] ,
    \Tile_X9Y14_FrameStrobe_O[1] ,
    \Tile_X9Y14_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X9Y14_N1BEG[3] ,
    \Tile_X9Y14_N1BEG[2] ,
    \Tile_X9Y14_N1BEG[1] ,
    \Tile_X9Y14_N1BEG[0] }),
    .N1END({\Tile_X9Y15_N1BEG[3] ,
    \Tile_X9Y15_N1BEG[2] ,
    \Tile_X9Y15_N1BEG[1] ,
    \Tile_X9Y15_N1BEG[0] }),
    .N2BEG({\Tile_X9Y14_N2BEG[7] ,
    \Tile_X9Y14_N2BEG[6] ,
    \Tile_X9Y14_N2BEG[5] ,
    \Tile_X9Y14_N2BEG[4] ,
    \Tile_X9Y14_N2BEG[3] ,
    \Tile_X9Y14_N2BEG[2] ,
    \Tile_X9Y14_N2BEG[1] ,
    \Tile_X9Y14_N2BEG[0] }),
    .N2BEGb({\Tile_X9Y14_N2BEGb[7] ,
    \Tile_X9Y14_N2BEGb[6] ,
    \Tile_X9Y14_N2BEGb[5] ,
    \Tile_X9Y14_N2BEGb[4] ,
    \Tile_X9Y14_N2BEGb[3] ,
    \Tile_X9Y14_N2BEGb[2] ,
    \Tile_X9Y14_N2BEGb[1] ,
    \Tile_X9Y14_N2BEGb[0] }),
    .N2END({\Tile_X9Y15_N2BEGb[7] ,
    \Tile_X9Y15_N2BEGb[6] ,
    \Tile_X9Y15_N2BEGb[5] ,
    \Tile_X9Y15_N2BEGb[4] ,
    \Tile_X9Y15_N2BEGb[3] ,
    \Tile_X9Y15_N2BEGb[2] ,
    \Tile_X9Y15_N2BEGb[1] ,
    \Tile_X9Y15_N2BEGb[0] }),
    .N2MID({\Tile_X9Y15_N2BEG[7] ,
    \Tile_X9Y15_N2BEG[6] ,
    \Tile_X9Y15_N2BEG[5] ,
    \Tile_X9Y15_N2BEG[4] ,
    \Tile_X9Y15_N2BEG[3] ,
    \Tile_X9Y15_N2BEG[2] ,
    \Tile_X9Y15_N2BEG[1] ,
    \Tile_X9Y15_N2BEG[0] }),
    .N4BEG({\Tile_X9Y14_N4BEG[15] ,
    \Tile_X9Y14_N4BEG[14] ,
    \Tile_X9Y14_N4BEG[13] ,
    \Tile_X9Y14_N4BEG[12] ,
    \Tile_X9Y14_N4BEG[11] ,
    \Tile_X9Y14_N4BEG[10] ,
    \Tile_X9Y14_N4BEG[9] ,
    \Tile_X9Y14_N4BEG[8] ,
    \Tile_X9Y14_N4BEG[7] ,
    \Tile_X9Y14_N4BEG[6] ,
    \Tile_X9Y14_N4BEG[5] ,
    \Tile_X9Y14_N4BEG[4] ,
    \Tile_X9Y14_N4BEG[3] ,
    \Tile_X9Y14_N4BEG[2] ,
    \Tile_X9Y14_N4BEG[1] ,
    \Tile_X9Y14_N4BEG[0] }),
    .N4END({\Tile_X9Y15_N4BEG[15] ,
    \Tile_X9Y15_N4BEG[14] ,
    \Tile_X9Y15_N4BEG[13] ,
    \Tile_X9Y15_N4BEG[12] ,
    \Tile_X9Y15_N4BEG[11] ,
    \Tile_X9Y15_N4BEG[10] ,
    \Tile_X9Y15_N4BEG[9] ,
    \Tile_X9Y15_N4BEG[8] ,
    \Tile_X9Y15_N4BEG[7] ,
    \Tile_X9Y15_N4BEG[6] ,
    \Tile_X9Y15_N4BEG[5] ,
    \Tile_X9Y15_N4BEG[4] ,
    \Tile_X9Y15_N4BEG[3] ,
    \Tile_X9Y15_N4BEG[2] ,
    \Tile_X9Y15_N4BEG[1] ,
    \Tile_X9Y15_N4BEG[0] }),
    .NN4BEG({\Tile_X9Y14_NN4BEG[15] ,
    \Tile_X9Y14_NN4BEG[14] ,
    \Tile_X9Y14_NN4BEG[13] ,
    \Tile_X9Y14_NN4BEG[12] ,
    \Tile_X9Y14_NN4BEG[11] ,
    \Tile_X9Y14_NN4BEG[10] ,
    \Tile_X9Y14_NN4BEG[9] ,
    \Tile_X9Y14_NN4BEG[8] ,
    \Tile_X9Y14_NN4BEG[7] ,
    \Tile_X9Y14_NN4BEG[6] ,
    \Tile_X9Y14_NN4BEG[5] ,
    \Tile_X9Y14_NN4BEG[4] ,
    \Tile_X9Y14_NN4BEG[3] ,
    \Tile_X9Y14_NN4BEG[2] ,
    \Tile_X9Y14_NN4BEG[1] ,
    \Tile_X9Y14_NN4BEG[0] }),
    .NN4END({\Tile_X9Y15_NN4BEG[15] ,
    \Tile_X9Y15_NN4BEG[14] ,
    \Tile_X9Y15_NN4BEG[13] ,
    \Tile_X9Y15_NN4BEG[12] ,
    \Tile_X9Y15_NN4BEG[11] ,
    \Tile_X9Y15_NN4BEG[10] ,
    \Tile_X9Y15_NN4BEG[9] ,
    \Tile_X9Y15_NN4BEG[8] ,
    \Tile_X9Y15_NN4BEG[7] ,
    \Tile_X9Y15_NN4BEG[6] ,
    \Tile_X9Y15_NN4BEG[5] ,
    \Tile_X9Y15_NN4BEG[4] ,
    \Tile_X9Y15_NN4BEG[3] ,
    \Tile_X9Y15_NN4BEG[2] ,
    \Tile_X9Y15_NN4BEG[1] ,
    \Tile_X9Y15_NN4BEG[0] }),
    .S1BEG({\Tile_X9Y14_S1BEG[3] ,
    \Tile_X9Y14_S1BEG[2] ,
    \Tile_X9Y14_S1BEG[1] ,
    \Tile_X9Y14_S1BEG[0] }),
    .S1END({\Tile_X9Y13_S1BEG[3] ,
    \Tile_X9Y13_S1BEG[2] ,
    \Tile_X9Y13_S1BEG[1] ,
    \Tile_X9Y13_S1BEG[0] }),
    .S2BEG({\Tile_X9Y14_S2BEG[7] ,
    \Tile_X9Y14_S2BEG[6] ,
    \Tile_X9Y14_S2BEG[5] ,
    \Tile_X9Y14_S2BEG[4] ,
    \Tile_X9Y14_S2BEG[3] ,
    \Tile_X9Y14_S2BEG[2] ,
    \Tile_X9Y14_S2BEG[1] ,
    \Tile_X9Y14_S2BEG[0] }),
    .S2BEGb({\Tile_X9Y14_S2BEGb[7] ,
    \Tile_X9Y14_S2BEGb[6] ,
    \Tile_X9Y14_S2BEGb[5] ,
    \Tile_X9Y14_S2BEGb[4] ,
    \Tile_X9Y14_S2BEGb[3] ,
    \Tile_X9Y14_S2BEGb[2] ,
    \Tile_X9Y14_S2BEGb[1] ,
    \Tile_X9Y14_S2BEGb[0] }),
    .S2END({\Tile_X9Y13_S2BEGb[7] ,
    \Tile_X9Y13_S2BEGb[6] ,
    \Tile_X9Y13_S2BEGb[5] ,
    \Tile_X9Y13_S2BEGb[4] ,
    \Tile_X9Y13_S2BEGb[3] ,
    \Tile_X9Y13_S2BEGb[2] ,
    \Tile_X9Y13_S2BEGb[1] ,
    \Tile_X9Y13_S2BEGb[0] }),
    .S2MID({\Tile_X9Y13_S2BEG[7] ,
    \Tile_X9Y13_S2BEG[6] ,
    \Tile_X9Y13_S2BEG[5] ,
    \Tile_X9Y13_S2BEG[4] ,
    \Tile_X9Y13_S2BEG[3] ,
    \Tile_X9Y13_S2BEG[2] ,
    \Tile_X9Y13_S2BEG[1] ,
    \Tile_X9Y13_S2BEG[0] }),
    .S4BEG({\Tile_X9Y14_S4BEG[15] ,
    \Tile_X9Y14_S4BEG[14] ,
    \Tile_X9Y14_S4BEG[13] ,
    \Tile_X9Y14_S4BEG[12] ,
    \Tile_X9Y14_S4BEG[11] ,
    \Tile_X9Y14_S4BEG[10] ,
    \Tile_X9Y14_S4BEG[9] ,
    \Tile_X9Y14_S4BEG[8] ,
    \Tile_X9Y14_S4BEG[7] ,
    \Tile_X9Y14_S4BEG[6] ,
    \Tile_X9Y14_S4BEG[5] ,
    \Tile_X9Y14_S4BEG[4] ,
    \Tile_X9Y14_S4BEG[3] ,
    \Tile_X9Y14_S4BEG[2] ,
    \Tile_X9Y14_S4BEG[1] ,
    \Tile_X9Y14_S4BEG[0] }),
    .S4END({\Tile_X9Y13_S4BEG[15] ,
    \Tile_X9Y13_S4BEG[14] ,
    \Tile_X9Y13_S4BEG[13] ,
    \Tile_X9Y13_S4BEG[12] ,
    \Tile_X9Y13_S4BEG[11] ,
    \Tile_X9Y13_S4BEG[10] ,
    \Tile_X9Y13_S4BEG[9] ,
    \Tile_X9Y13_S4BEG[8] ,
    \Tile_X9Y13_S4BEG[7] ,
    \Tile_X9Y13_S4BEG[6] ,
    \Tile_X9Y13_S4BEG[5] ,
    \Tile_X9Y13_S4BEG[4] ,
    \Tile_X9Y13_S4BEG[3] ,
    \Tile_X9Y13_S4BEG[2] ,
    \Tile_X9Y13_S4BEG[1] ,
    \Tile_X9Y13_S4BEG[0] }),
    .SS4BEG({\Tile_X9Y14_SS4BEG[15] ,
    \Tile_X9Y14_SS4BEG[14] ,
    \Tile_X9Y14_SS4BEG[13] ,
    \Tile_X9Y14_SS4BEG[12] ,
    \Tile_X9Y14_SS4BEG[11] ,
    \Tile_X9Y14_SS4BEG[10] ,
    \Tile_X9Y14_SS4BEG[9] ,
    \Tile_X9Y14_SS4BEG[8] ,
    \Tile_X9Y14_SS4BEG[7] ,
    \Tile_X9Y14_SS4BEG[6] ,
    \Tile_X9Y14_SS4BEG[5] ,
    \Tile_X9Y14_SS4BEG[4] ,
    \Tile_X9Y14_SS4BEG[3] ,
    \Tile_X9Y14_SS4BEG[2] ,
    \Tile_X9Y14_SS4BEG[1] ,
    \Tile_X9Y14_SS4BEG[0] }),
    .SS4END({\Tile_X9Y13_SS4BEG[15] ,
    \Tile_X9Y13_SS4BEG[14] ,
    \Tile_X9Y13_SS4BEG[13] ,
    \Tile_X9Y13_SS4BEG[12] ,
    \Tile_X9Y13_SS4BEG[11] ,
    \Tile_X9Y13_SS4BEG[10] ,
    \Tile_X9Y13_SS4BEG[9] ,
    \Tile_X9Y13_SS4BEG[8] ,
    \Tile_X9Y13_SS4BEG[7] ,
    \Tile_X9Y13_SS4BEG[6] ,
    \Tile_X9Y13_SS4BEG[5] ,
    \Tile_X9Y13_SS4BEG[4] ,
    \Tile_X9Y13_SS4BEG[3] ,
    \Tile_X9Y13_SS4BEG[2] ,
    \Tile_X9Y13_SS4BEG[1] ,
    \Tile_X9Y13_SS4BEG[0] }),
    .W1BEG({\Tile_X9Y14_W1BEG[3] ,
    \Tile_X9Y14_W1BEG[2] ,
    \Tile_X9Y14_W1BEG[1] ,
    \Tile_X9Y14_W1BEG[0] }),
    .W1END({\Tile_X10Y14_W1BEG[3] ,
    \Tile_X10Y14_W1BEG[2] ,
    \Tile_X10Y14_W1BEG[1] ,
    \Tile_X10Y14_W1BEG[0] }),
    .W2BEG({\Tile_X9Y14_W2BEG[7] ,
    \Tile_X9Y14_W2BEG[6] ,
    \Tile_X9Y14_W2BEG[5] ,
    \Tile_X9Y14_W2BEG[4] ,
    \Tile_X9Y14_W2BEG[3] ,
    \Tile_X9Y14_W2BEG[2] ,
    \Tile_X9Y14_W2BEG[1] ,
    \Tile_X9Y14_W2BEG[0] }),
    .W2BEGb({\Tile_X9Y14_W2BEGb[7] ,
    \Tile_X9Y14_W2BEGb[6] ,
    \Tile_X9Y14_W2BEGb[5] ,
    \Tile_X9Y14_W2BEGb[4] ,
    \Tile_X9Y14_W2BEGb[3] ,
    \Tile_X9Y14_W2BEGb[2] ,
    \Tile_X9Y14_W2BEGb[1] ,
    \Tile_X9Y14_W2BEGb[0] }),
    .W2END({\Tile_X10Y14_W2BEGb[7] ,
    \Tile_X10Y14_W2BEGb[6] ,
    \Tile_X10Y14_W2BEGb[5] ,
    \Tile_X10Y14_W2BEGb[4] ,
    \Tile_X10Y14_W2BEGb[3] ,
    \Tile_X10Y14_W2BEGb[2] ,
    \Tile_X10Y14_W2BEGb[1] ,
    \Tile_X10Y14_W2BEGb[0] }),
    .W2MID({\Tile_X10Y14_W2BEG[7] ,
    \Tile_X10Y14_W2BEG[6] ,
    \Tile_X10Y14_W2BEG[5] ,
    \Tile_X10Y14_W2BEG[4] ,
    \Tile_X10Y14_W2BEG[3] ,
    \Tile_X10Y14_W2BEG[2] ,
    \Tile_X10Y14_W2BEG[1] ,
    \Tile_X10Y14_W2BEG[0] }),
    .W6BEG({\Tile_X9Y14_W6BEG[11] ,
    \Tile_X9Y14_W6BEG[10] ,
    \Tile_X9Y14_W6BEG[9] ,
    \Tile_X9Y14_W6BEG[8] ,
    \Tile_X9Y14_W6BEG[7] ,
    \Tile_X9Y14_W6BEG[6] ,
    \Tile_X9Y14_W6BEG[5] ,
    \Tile_X9Y14_W6BEG[4] ,
    \Tile_X9Y14_W6BEG[3] ,
    \Tile_X9Y14_W6BEG[2] ,
    \Tile_X9Y14_W6BEG[1] ,
    \Tile_X9Y14_W6BEG[0] }),
    .W6END({\Tile_X10Y14_W6BEG[11] ,
    \Tile_X10Y14_W6BEG[10] ,
    \Tile_X10Y14_W6BEG[9] ,
    \Tile_X10Y14_W6BEG[8] ,
    \Tile_X10Y14_W6BEG[7] ,
    \Tile_X10Y14_W6BEG[6] ,
    \Tile_X10Y14_W6BEG[5] ,
    \Tile_X10Y14_W6BEG[4] ,
    \Tile_X10Y14_W6BEG[3] ,
    \Tile_X10Y14_W6BEG[2] ,
    \Tile_X10Y14_W6BEG[1] ,
    \Tile_X10Y14_W6BEG[0] }),
    .WW4BEG({\Tile_X9Y14_WW4BEG[15] ,
    \Tile_X9Y14_WW4BEG[14] ,
    \Tile_X9Y14_WW4BEG[13] ,
    \Tile_X9Y14_WW4BEG[12] ,
    \Tile_X9Y14_WW4BEG[11] ,
    \Tile_X9Y14_WW4BEG[10] ,
    \Tile_X9Y14_WW4BEG[9] ,
    \Tile_X9Y14_WW4BEG[8] ,
    \Tile_X9Y14_WW4BEG[7] ,
    \Tile_X9Y14_WW4BEG[6] ,
    \Tile_X9Y14_WW4BEG[5] ,
    \Tile_X9Y14_WW4BEG[4] ,
    \Tile_X9Y14_WW4BEG[3] ,
    \Tile_X9Y14_WW4BEG[2] ,
    \Tile_X9Y14_WW4BEG[1] ,
    \Tile_X9Y14_WW4BEG[0] }),
    .WW4END({\Tile_X10Y14_WW4BEG[15] ,
    \Tile_X10Y14_WW4BEG[14] ,
    \Tile_X10Y14_WW4BEG[13] ,
    \Tile_X10Y14_WW4BEG[12] ,
    \Tile_X10Y14_WW4BEG[11] ,
    \Tile_X10Y14_WW4BEG[10] ,
    \Tile_X10Y14_WW4BEG[9] ,
    \Tile_X10Y14_WW4BEG[8] ,
    \Tile_X10Y14_WW4BEG[7] ,
    \Tile_X10Y14_WW4BEG[6] ,
    \Tile_X10Y14_WW4BEG[5] ,
    \Tile_X10Y14_WW4BEG[4] ,
    \Tile_X10Y14_WW4BEG[3] ,
    \Tile_X10Y14_WW4BEG[2] ,
    \Tile_X10Y14_WW4BEG[1] ,
    \Tile_X10Y14_WW4BEG[0] }));
 S_CPU_IF Tile_X9Y15_S_CPU_IF (.Co(Tile_X9Y15_Co),
    .I_top0(Tile_X9Y15_I_top0),
    .I_top1(Tile_X9Y15_I_top1),
    .I_top10(Tile_X9Y15_I_top10),
    .I_top11(Tile_X9Y15_I_top11),
    .I_top12(Tile_X9Y15_I_top12),
    .I_top13(Tile_X9Y15_I_top13),
    .I_top14(Tile_X9Y15_I_top14),
    .I_top15(Tile_X9Y15_I_top15),
    .I_top2(Tile_X9Y15_I_top2),
    .I_top3(Tile_X9Y15_I_top3),
    .I_top4(Tile_X9Y15_I_top4),
    .I_top5(Tile_X9Y15_I_top5),
    .I_top6(Tile_X9Y15_I_top6),
    .I_top7(Tile_X9Y15_I_top7),
    .I_top8(Tile_X9Y15_I_top8),
    .I_top9(Tile_X9Y15_I_top9),
    .O_top0(Tile_X9Y15_O_top0),
    .O_top1(Tile_X9Y15_O_top1),
    .O_top10(Tile_X9Y15_O_top10),
    .O_top11(Tile_X9Y15_O_top11),
    .O_top12(Tile_X9Y15_O_top12),
    .O_top13(Tile_X9Y15_O_top13),
    .O_top14(Tile_X9Y15_O_top14),
    .O_top15(Tile_X9Y15_O_top15),
    .O_top2(Tile_X9Y15_O_top2),
    .O_top3(Tile_X9Y15_O_top3),
    .O_top4(Tile_X9Y15_O_top4),
    .O_top5(Tile_X9Y15_O_top5),
    .O_top6(Tile_X9Y15_O_top6),
    .O_top7(Tile_X9Y15_O_top7),
    .O_top8(Tile_X9Y15_O_top8),
    .O_top9(Tile_X9Y15_O_top9),
    .UserCLK(UserCLK),
    .UserCLKo(Tile_X9Y15_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .FrameData({\Tile_X8Y15_FrameData_O[31] ,
    \Tile_X8Y15_FrameData_O[30] ,
    \Tile_X8Y15_FrameData_O[29] ,
    \Tile_X8Y15_FrameData_O[28] ,
    \Tile_X8Y15_FrameData_O[27] ,
    \Tile_X8Y15_FrameData_O[26] ,
    \Tile_X8Y15_FrameData_O[25] ,
    \Tile_X8Y15_FrameData_O[24] ,
    \Tile_X8Y15_FrameData_O[23] ,
    \Tile_X8Y15_FrameData_O[22] ,
    \Tile_X8Y15_FrameData_O[21] ,
    \Tile_X8Y15_FrameData_O[20] ,
    \Tile_X8Y15_FrameData_O[19] ,
    \Tile_X8Y15_FrameData_O[18] ,
    \Tile_X8Y15_FrameData_O[17] ,
    \Tile_X8Y15_FrameData_O[16] ,
    \Tile_X8Y15_FrameData_O[15] ,
    \Tile_X8Y15_FrameData_O[14] ,
    \Tile_X8Y15_FrameData_O[13] ,
    \Tile_X8Y15_FrameData_O[12] ,
    \Tile_X8Y15_FrameData_O[11] ,
    \Tile_X8Y15_FrameData_O[10] ,
    \Tile_X8Y15_FrameData_O[9] ,
    \Tile_X8Y15_FrameData_O[8] ,
    \Tile_X8Y15_FrameData_O[7] ,
    \Tile_X8Y15_FrameData_O[6] ,
    \Tile_X8Y15_FrameData_O[5] ,
    \Tile_X8Y15_FrameData_O[4] ,
    \Tile_X8Y15_FrameData_O[3] ,
    \Tile_X8Y15_FrameData_O[2] ,
    \Tile_X8Y15_FrameData_O[1] ,
    \Tile_X8Y15_FrameData_O[0] }),
    .FrameData_O({\Tile_X9Y15_FrameData_O[31] ,
    \Tile_X9Y15_FrameData_O[30] ,
    \Tile_X9Y15_FrameData_O[29] ,
    \Tile_X9Y15_FrameData_O[28] ,
    \Tile_X9Y15_FrameData_O[27] ,
    \Tile_X9Y15_FrameData_O[26] ,
    \Tile_X9Y15_FrameData_O[25] ,
    \Tile_X9Y15_FrameData_O[24] ,
    \Tile_X9Y15_FrameData_O[23] ,
    \Tile_X9Y15_FrameData_O[22] ,
    \Tile_X9Y15_FrameData_O[21] ,
    \Tile_X9Y15_FrameData_O[20] ,
    \Tile_X9Y15_FrameData_O[19] ,
    \Tile_X9Y15_FrameData_O[18] ,
    \Tile_X9Y15_FrameData_O[17] ,
    \Tile_X9Y15_FrameData_O[16] ,
    \Tile_X9Y15_FrameData_O[15] ,
    \Tile_X9Y15_FrameData_O[14] ,
    \Tile_X9Y15_FrameData_O[13] ,
    \Tile_X9Y15_FrameData_O[12] ,
    \Tile_X9Y15_FrameData_O[11] ,
    \Tile_X9Y15_FrameData_O[10] ,
    \Tile_X9Y15_FrameData_O[9] ,
    \Tile_X9Y15_FrameData_O[8] ,
    \Tile_X9Y15_FrameData_O[7] ,
    \Tile_X9Y15_FrameData_O[6] ,
    \Tile_X9Y15_FrameData_O[5] ,
    \Tile_X9Y15_FrameData_O[4] ,
    \Tile_X9Y15_FrameData_O[3] ,
    \Tile_X9Y15_FrameData_O[2] ,
    \Tile_X9Y15_FrameData_O[1] ,
    \Tile_X9Y15_FrameData_O[0] }),
    .FrameStrobe({FrameStrobe[199],
    FrameStrobe[198],
    FrameStrobe[197],
    FrameStrobe[196],
    FrameStrobe[195],
    FrameStrobe[194],
    FrameStrobe[193],
    FrameStrobe[192],
    FrameStrobe[191],
    FrameStrobe[190],
    FrameStrobe[189],
    FrameStrobe[188],
    FrameStrobe[187],
    FrameStrobe[186],
    FrameStrobe[185],
    FrameStrobe[184],
    FrameStrobe[183],
    FrameStrobe[182],
    FrameStrobe[181],
    FrameStrobe[180]}),
    .FrameStrobe_O({\Tile_X9Y15_FrameStrobe_O[19] ,
    \Tile_X9Y15_FrameStrobe_O[18] ,
    \Tile_X9Y15_FrameStrobe_O[17] ,
    \Tile_X9Y15_FrameStrobe_O[16] ,
    \Tile_X9Y15_FrameStrobe_O[15] ,
    \Tile_X9Y15_FrameStrobe_O[14] ,
    \Tile_X9Y15_FrameStrobe_O[13] ,
    \Tile_X9Y15_FrameStrobe_O[12] ,
    \Tile_X9Y15_FrameStrobe_O[11] ,
    \Tile_X9Y15_FrameStrobe_O[10] ,
    \Tile_X9Y15_FrameStrobe_O[9] ,
    \Tile_X9Y15_FrameStrobe_O[8] ,
    \Tile_X9Y15_FrameStrobe_O[7] ,
    \Tile_X9Y15_FrameStrobe_O[6] ,
    \Tile_X9Y15_FrameStrobe_O[5] ,
    \Tile_X9Y15_FrameStrobe_O[4] ,
    \Tile_X9Y15_FrameStrobe_O[3] ,
    \Tile_X9Y15_FrameStrobe_O[2] ,
    \Tile_X9Y15_FrameStrobe_O[1] ,
    \Tile_X9Y15_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X9Y15_N1BEG[3] ,
    \Tile_X9Y15_N1BEG[2] ,
    \Tile_X9Y15_N1BEG[1] ,
    \Tile_X9Y15_N1BEG[0] }),
    .N2BEG({\Tile_X9Y15_N2BEG[7] ,
    \Tile_X9Y15_N2BEG[6] ,
    \Tile_X9Y15_N2BEG[5] ,
    \Tile_X9Y15_N2BEG[4] ,
    \Tile_X9Y15_N2BEG[3] ,
    \Tile_X9Y15_N2BEG[2] ,
    \Tile_X9Y15_N2BEG[1] ,
    \Tile_X9Y15_N2BEG[0] }),
    .N2BEGb({\Tile_X9Y15_N2BEGb[7] ,
    \Tile_X9Y15_N2BEGb[6] ,
    \Tile_X9Y15_N2BEGb[5] ,
    \Tile_X9Y15_N2BEGb[4] ,
    \Tile_X9Y15_N2BEGb[3] ,
    \Tile_X9Y15_N2BEGb[2] ,
    \Tile_X9Y15_N2BEGb[1] ,
    \Tile_X9Y15_N2BEGb[0] }),
    .N4BEG({\Tile_X9Y15_N4BEG[15] ,
    \Tile_X9Y15_N4BEG[14] ,
    \Tile_X9Y15_N4BEG[13] ,
    \Tile_X9Y15_N4BEG[12] ,
    \Tile_X9Y15_N4BEG[11] ,
    \Tile_X9Y15_N4BEG[10] ,
    \Tile_X9Y15_N4BEG[9] ,
    \Tile_X9Y15_N4BEG[8] ,
    \Tile_X9Y15_N4BEG[7] ,
    \Tile_X9Y15_N4BEG[6] ,
    \Tile_X9Y15_N4BEG[5] ,
    \Tile_X9Y15_N4BEG[4] ,
    \Tile_X9Y15_N4BEG[3] ,
    \Tile_X9Y15_N4BEG[2] ,
    \Tile_X9Y15_N4BEG[1] ,
    \Tile_X9Y15_N4BEG[0] }),
    .NN4BEG({\Tile_X9Y15_NN4BEG[15] ,
    \Tile_X9Y15_NN4BEG[14] ,
    \Tile_X9Y15_NN4BEG[13] ,
    \Tile_X9Y15_NN4BEG[12] ,
    \Tile_X9Y15_NN4BEG[11] ,
    \Tile_X9Y15_NN4BEG[10] ,
    \Tile_X9Y15_NN4BEG[9] ,
    \Tile_X9Y15_NN4BEG[8] ,
    \Tile_X9Y15_NN4BEG[7] ,
    \Tile_X9Y15_NN4BEG[6] ,
    \Tile_X9Y15_NN4BEG[5] ,
    \Tile_X9Y15_NN4BEG[4] ,
    \Tile_X9Y15_NN4BEG[3] ,
    \Tile_X9Y15_NN4BEG[2] ,
    \Tile_X9Y15_NN4BEG[1] ,
    \Tile_X9Y15_NN4BEG[0] }),
    .S1END({\Tile_X9Y14_S1BEG[3] ,
    \Tile_X9Y14_S1BEG[2] ,
    \Tile_X9Y14_S1BEG[1] ,
    \Tile_X9Y14_S1BEG[0] }),
    .S2END({\Tile_X9Y14_S2BEGb[7] ,
    \Tile_X9Y14_S2BEGb[6] ,
    \Tile_X9Y14_S2BEGb[5] ,
    \Tile_X9Y14_S2BEGb[4] ,
    \Tile_X9Y14_S2BEGb[3] ,
    \Tile_X9Y14_S2BEGb[2] ,
    \Tile_X9Y14_S2BEGb[1] ,
    \Tile_X9Y14_S2BEGb[0] }),
    .S2MID({\Tile_X9Y14_S2BEG[7] ,
    \Tile_X9Y14_S2BEG[6] ,
    \Tile_X9Y14_S2BEG[5] ,
    \Tile_X9Y14_S2BEG[4] ,
    \Tile_X9Y14_S2BEG[3] ,
    \Tile_X9Y14_S2BEG[2] ,
    \Tile_X9Y14_S2BEG[1] ,
    \Tile_X9Y14_S2BEG[0] }),
    .S4END({\Tile_X9Y14_S4BEG[15] ,
    \Tile_X9Y14_S4BEG[14] ,
    \Tile_X9Y14_S4BEG[13] ,
    \Tile_X9Y14_S4BEG[12] ,
    \Tile_X9Y14_S4BEG[11] ,
    \Tile_X9Y14_S4BEG[10] ,
    \Tile_X9Y14_S4BEG[9] ,
    \Tile_X9Y14_S4BEG[8] ,
    \Tile_X9Y14_S4BEG[7] ,
    \Tile_X9Y14_S4BEG[6] ,
    \Tile_X9Y14_S4BEG[5] ,
    \Tile_X9Y14_S4BEG[4] ,
    \Tile_X9Y14_S4BEG[3] ,
    \Tile_X9Y14_S4BEG[2] ,
    \Tile_X9Y14_S4BEG[1] ,
    \Tile_X9Y14_S4BEG[0] }),
    .SS4END({\Tile_X9Y14_SS4BEG[15] ,
    \Tile_X9Y14_SS4BEG[14] ,
    \Tile_X9Y14_SS4BEG[13] ,
    \Tile_X9Y14_SS4BEG[12] ,
    \Tile_X9Y14_SS4BEG[11] ,
    \Tile_X9Y14_SS4BEG[10] ,
    \Tile_X9Y14_SS4BEG[9] ,
    \Tile_X9Y14_SS4BEG[8] ,
    \Tile_X9Y14_SS4BEG[7] ,
    \Tile_X9Y14_SS4BEG[6] ,
    \Tile_X9Y14_SS4BEG[5] ,
    \Tile_X9Y14_SS4BEG[4] ,
    \Tile_X9Y14_SS4BEG[3] ,
    \Tile_X9Y14_SS4BEG[2] ,
    \Tile_X9Y14_SS4BEG[1] ,
    \Tile_X9Y14_SS4BEG[0] }));
 LUT4AB Tile_X9Y1_LUT4AB (.Ci(Tile_X9Y2_Co),
    .Co(Tile_X9Y1_Co),
    .UserCLK(Tile_X9Y2_UserCLKo),
    .UserCLKo(Tile_X9Y1_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X9Y1_E1BEG[3] ,
    \Tile_X9Y1_E1BEG[2] ,
    \Tile_X9Y1_E1BEG[1] ,
    \Tile_X9Y1_E1BEG[0] }),
    .E1END({\Tile_X8Y1_E1BEG[3] ,
    \Tile_X8Y1_E1BEG[2] ,
    \Tile_X8Y1_E1BEG[1] ,
    \Tile_X8Y1_E1BEG[0] }),
    .E2BEG({\Tile_X9Y1_E2BEG[7] ,
    \Tile_X9Y1_E2BEG[6] ,
    \Tile_X9Y1_E2BEG[5] ,
    \Tile_X9Y1_E2BEG[4] ,
    \Tile_X9Y1_E2BEG[3] ,
    \Tile_X9Y1_E2BEG[2] ,
    \Tile_X9Y1_E2BEG[1] ,
    \Tile_X9Y1_E2BEG[0] }),
    .E2BEGb({\Tile_X9Y1_E2BEGb[7] ,
    \Tile_X9Y1_E2BEGb[6] ,
    \Tile_X9Y1_E2BEGb[5] ,
    \Tile_X9Y1_E2BEGb[4] ,
    \Tile_X9Y1_E2BEGb[3] ,
    \Tile_X9Y1_E2BEGb[2] ,
    \Tile_X9Y1_E2BEGb[1] ,
    \Tile_X9Y1_E2BEGb[0] }),
    .E2END({\Tile_X8Y1_E2BEGb[7] ,
    \Tile_X8Y1_E2BEGb[6] ,
    \Tile_X8Y1_E2BEGb[5] ,
    \Tile_X8Y1_E2BEGb[4] ,
    \Tile_X8Y1_E2BEGb[3] ,
    \Tile_X8Y1_E2BEGb[2] ,
    \Tile_X8Y1_E2BEGb[1] ,
    \Tile_X8Y1_E2BEGb[0] }),
    .E2MID({\Tile_X8Y1_E2BEG[7] ,
    \Tile_X8Y1_E2BEG[6] ,
    \Tile_X8Y1_E2BEG[5] ,
    \Tile_X8Y1_E2BEG[4] ,
    \Tile_X8Y1_E2BEG[3] ,
    \Tile_X8Y1_E2BEG[2] ,
    \Tile_X8Y1_E2BEG[1] ,
    \Tile_X8Y1_E2BEG[0] }),
    .E6BEG({\Tile_X9Y1_E6BEG[11] ,
    \Tile_X9Y1_E6BEG[10] ,
    \Tile_X9Y1_E6BEG[9] ,
    \Tile_X9Y1_E6BEG[8] ,
    \Tile_X9Y1_E6BEG[7] ,
    \Tile_X9Y1_E6BEG[6] ,
    \Tile_X9Y1_E6BEG[5] ,
    \Tile_X9Y1_E6BEG[4] ,
    \Tile_X9Y1_E6BEG[3] ,
    \Tile_X9Y1_E6BEG[2] ,
    \Tile_X9Y1_E6BEG[1] ,
    \Tile_X9Y1_E6BEG[0] }),
    .E6END({\Tile_X8Y1_E6BEG[11] ,
    \Tile_X8Y1_E6BEG[10] ,
    \Tile_X8Y1_E6BEG[9] ,
    \Tile_X8Y1_E6BEG[8] ,
    \Tile_X8Y1_E6BEG[7] ,
    \Tile_X8Y1_E6BEG[6] ,
    \Tile_X8Y1_E6BEG[5] ,
    \Tile_X8Y1_E6BEG[4] ,
    \Tile_X8Y1_E6BEG[3] ,
    \Tile_X8Y1_E6BEG[2] ,
    \Tile_X8Y1_E6BEG[1] ,
    \Tile_X8Y1_E6BEG[0] }),
    .EE4BEG({\Tile_X9Y1_EE4BEG[15] ,
    \Tile_X9Y1_EE4BEG[14] ,
    \Tile_X9Y1_EE4BEG[13] ,
    \Tile_X9Y1_EE4BEG[12] ,
    \Tile_X9Y1_EE4BEG[11] ,
    \Tile_X9Y1_EE4BEG[10] ,
    \Tile_X9Y1_EE4BEG[9] ,
    \Tile_X9Y1_EE4BEG[8] ,
    \Tile_X9Y1_EE4BEG[7] ,
    \Tile_X9Y1_EE4BEG[6] ,
    \Tile_X9Y1_EE4BEG[5] ,
    \Tile_X9Y1_EE4BEG[4] ,
    \Tile_X9Y1_EE4BEG[3] ,
    \Tile_X9Y1_EE4BEG[2] ,
    \Tile_X9Y1_EE4BEG[1] ,
    \Tile_X9Y1_EE4BEG[0] }),
    .EE4END({\Tile_X8Y1_EE4BEG[15] ,
    \Tile_X8Y1_EE4BEG[14] ,
    \Tile_X8Y1_EE4BEG[13] ,
    \Tile_X8Y1_EE4BEG[12] ,
    \Tile_X8Y1_EE4BEG[11] ,
    \Tile_X8Y1_EE4BEG[10] ,
    \Tile_X8Y1_EE4BEG[9] ,
    \Tile_X8Y1_EE4BEG[8] ,
    \Tile_X8Y1_EE4BEG[7] ,
    \Tile_X8Y1_EE4BEG[6] ,
    \Tile_X8Y1_EE4BEG[5] ,
    \Tile_X8Y1_EE4BEG[4] ,
    \Tile_X8Y1_EE4BEG[3] ,
    \Tile_X8Y1_EE4BEG[2] ,
    \Tile_X8Y1_EE4BEG[1] ,
    \Tile_X8Y1_EE4BEG[0] }),
    .FrameData({\Tile_X8Y1_FrameData_O[31] ,
    \Tile_X8Y1_FrameData_O[30] ,
    \Tile_X8Y1_FrameData_O[29] ,
    \Tile_X8Y1_FrameData_O[28] ,
    \Tile_X8Y1_FrameData_O[27] ,
    \Tile_X8Y1_FrameData_O[26] ,
    \Tile_X8Y1_FrameData_O[25] ,
    \Tile_X8Y1_FrameData_O[24] ,
    \Tile_X8Y1_FrameData_O[23] ,
    \Tile_X8Y1_FrameData_O[22] ,
    \Tile_X8Y1_FrameData_O[21] ,
    \Tile_X8Y1_FrameData_O[20] ,
    \Tile_X8Y1_FrameData_O[19] ,
    \Tile_X8Y1_FrameData_O[18] ,
    \Tile_X8Y1_FrameData_O[17] ,
    \Tile_X8Y1_FrameData_O[16] ,
    \Tile_X8Y1_FrameData_O[15] ,
    \Tile_X8Y1_FrameData_O[14] ,
    \Tile_X8Y1_FrameData_O[13] ,
    \Tile_X8Y1_FrameData_O[12] ,
    \Tile_X8Y1_FrameData_O[11] ,
    \Tile_X8Y1_FrameData_O[10] ,
    \Tile_X8Y1_FrameData_O[9] ,
    \Tile_X8Y1_FrameData_O[8] ,
    \Tile_X8Y1_FrameData_O[7] ,
    \Tile_X8Y1_FrameData_O[6] ,
    \Tile_X8Y1_FrameData_O[5] ,
    \Tile_X8Y1_FrameData_O[4] ,
    \Tile_X8Y1_FrameData_O[3] ,
    \Tile_X8Y1_FrameData_O[2] ,
    \Tile_X8Y1_FrameData_O[1] ,
    \Tile_X8Y1_FrameData_O[0] }),
    .FrameData_O({\Tile_X9Y1_FrameData_O[31] ,
    \Tile_X9Y1_FrameData_O[30] ,
    \Tile_X9Y1_FrameData_O[29] ,
    \Tile_X9Y1_FrameData_O[28] ,
    \Tile_X9Y1_FrameData_O[27] ,
    \Tile_X9Y1_FrameData_O[26] ,
    \Tile_X9Y1_FrameData_O[25] ,
    \Tile_X9Y1_FrameData_O[24] ,
    \Tile_X9Y1_FrameData_O[23] ,
    \Tile_X9Y1_FrameData_O[22] ,
    \Tile_X9Y1_FrameData_O[21] ,
    \Tile_X9Y1_FrameData_O[20] ,
    \Tile_X9Y1_FrameData_O[19] ,
    \Tile_X9Y1_FrameData_O[18] ,
    \Tile_X9Y1_FrameData_O[17] ,
    \Tile_X9Y1_FrameData_O[16] ,
    \Tile_X9Y1_FrameData_O[15] ,
    \Tile_X9Y1_FrameData_O[14] ,
    \Tile_X9Y1_FrameData_O[13] ,
    \Tile_X9Y1_FrameData_O[12] ,
    \Tile_X9Y1_FrameData_O[11] ,
    \Tile_X9Y1_FrameData_O[10] ,
    \Tile_X9Y1_FrameData_O[9] ,
    \Tile_X9Y1_FrameData_O[8] ,
    \Tile_X9Y1_FrameData_O[7] ,
    \Tile_X9Y1_FrameData_O[6] ,
    \Tile_X9Y1_FrameData_O[5] ,
    \Tile_X9Y1_FrameData_O[4] ,
    \Tile_X9Y1_FrameData_O[3] ,
    \Tile_X9Y1_FrameData_O[2] ,
    \Tile_X9Y1_FrameData_O[1] ,
    \Tile_X9Y1_FrameData_O[0] }),
    .FrameStrobe({\Tile_X9Y2_FrameStrobe_O[19] ,
    \Tile_X9Y2_FrameStrobe_O[18] ,
    \Tile_X9Y2_FrameStrobe_O[17] ,
    \Tile_X9Y2_FrameStrobe_O[16] ,
    \Tile_X9Y2_FrameStrobe_O[15] ,
    \Tile_X9Y2_FrameStrobe_O[14] ,
    \Tile_X9Y2_FrameStrobe_O[13] ,
    \Tile_X9Y2_FrameStrobe_O[12] ,
    \Tile_X9Y2_FrameStrobe_O[11] ,
    \Tile_X9Y2_FrameStrobe_O[10] ,
    \Tile_X9Y2_FrameStrobe_O[9] ,
    \Tile_X9Y2_FrameStrobe_O[8] ,
    \Tile_X9Y2_FrameStrobe_O[7] ,
    \Tile_X9Y2_FrameStrobe_O[6] ,
    \Tile_X9Y2_FrameStrobe_O[5] ,
    \Tile_X9Y2_FrameStrobe_O[4] ,
    \Tile_X9Y2_FrameStrobe_O[3] ,
    \Tile_X9Y2_FrameStrobe_O[2] ,
    \Tile_X9Y2_FrameStrobe_O[1] ,
    \Tile_X9Y2_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X9Y1_FrameStrobe_O[19] ,
    \Tile_X9Y1_FrameStrobe_O[18] ,
    \Tile_X9Y1_FrameStrobe_O[17] ,
    \Tile_X9Y1_FrameStrobe_O[16] ,
    \Tile_X9Y1_FrameStrobe_O[15] ,
    \Tile_X9Y1_FrameStrobe_O[14] ,
    \Tile_X9Y1_FrameStrobe_O[13] ,
    \Tile_X9Y1_FrameStrobe_O[12] ,
    \Tile_X9Y1_FrameStrobe_O[11] ,
    \Tile_X9Y1_FrameStrobe_O[10] ,
    \Tile_X9Y1_FrameStrobe_O[9] ,
    \Tile_X9Y1_FrameStrobe_O[8] ,
    \Tile_X9Y1_FrameStrobe_O[7] ,
    \Tile_X9Y1_FrameStrobe_O[6] ,
    \Tile_X9Y1_FrameStrobe_O[5] ,
    \Tile_X9Y1_FrameStrobe_O[4] ,
    \Tile_X9Y1_FrameStrobe_O[3] ,
    \Tile_X9Y1_FrameStrobe_O[2] ,
    \Tile_X9Y1_FrameStrobe_O[1] ,
    \Tile_X9Y1_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X9Y1_N1BEG[3] ,
    \Tile_X9Y1_N1BEG[2] ,
    \Tile_X9Y1_N1BEG[1] ,
    \Tile_X9Y1_N1BEG[0] }),
    .N1END({\Tile_X9Y2_N1BEG[3] ,
    \Tile_X9Y2_N1BEG[2] ,
    \Tile_X9Y2_N1BEG[1] ,
    \Tile_X9Y2_N1BEG[0] }),
    .N2BEG({\Tile_X9Y1_N2BEG[7] ,
    \Tile_X9Y1_N2BEG[6] ,
    \Tile_X9Y1_N2BEG[5] ,
    \Tile_X9Y1_N2BEG[4] ,
    \Tile_X9Y1_N2BEG[3] ,
    \Tile_X9Y1_N2BEG[2] ,
    \Tile_X9Y1_N2BEG[1] ,
    \Tile_X9Y1_N2BEG[0] }),
    .N2BEGb({\Tile_X9Y1_N2BEGb[7] ,
    \Tile_X9Y1_N2BEGb[6] ,
    \Tile_X9Y1_N2BEGb[5] ,
    \Tile_X9Y1_N2BEGb[4] ,
    \Tile_X9Y1_N2BEGb[3] ,
    \Tile_X9Y1_N2BEGb[2] ,
    \Tile_X9Y1_N2BEGb[1] ,
    \Tile_X9Y1_N2BEGb[0] }),
    .N2END({\Tile_X9Y2_N2BEGb[7] ,
    \Tile_X9Y2_N2BEGb[6] ,
    \Tile_X9Y2_N2BEGb[5] ,
    \Tile_X9Y2_N2BEGb[4] ,
    \Tile_X9Y2_N2BEGb[3] ,
    \Tile_X9Y2_N2BEGb[2] ,
    \Tile_X9Y2_N2BEGb[1] ,
    \Tile_X9Y2_N2BEGb[0] }),
    .N2MID({\Tile_X9Y2_N2BEG[7] ,
    \Tile_X9Y2_N2BEG[6] ,
    \Tile_X9Y2_N2BEG[5] ,
    \Tile_X9Y2_N2BEG[4] ,
    \Tile_X9Y2_N2BEG[3] ,
    \Tile_X9Y2_N2BEG[2] ,
    \Tile_X9Y2_N2BEG[1] ,
    \Tile_X9Y2_N2BEG[0] }),
    .N4BEG({\Tile_X9Y1_N4BEG[15] ,
    \Tile_X9Y1_N4BEG[14] ,
    \Tile_X9Y1_N4BEG[13] ,
    \Tile_X9Y1_N4BEG[12] ,
    \Tile_X9Y1_N4BEG[11] ,
    \Tile_X9Y1_N4BEG[10] ,
    \Tile_X9Y1_N4BEG[9] ,
    \Tile_X9Y1_N4BEG[8] ,
    \Tile_X9Y1_N4BEG[7] ,
    \Tile_X9Y1_N4BEG[6] ,
    \Tile_X9Y1_N4BEG[5] ,
    \Tile_X9Y1_N4BEG[4] ,
    \Tile_X9Y1_N4BEG[3] ,
    \Tile_X9Y1_N4BEG[2] ,
    \Tile_X9Y1_N4BEG[1] ,
    \Tile_X9Y1_N4BEG[0] }),
    .N4END({\Tile_X9Y2_N4BEG[15] ,
    \Tile_X9Y2_N4BEG[14] ,
    \Tile_X9Y2_N4BEG[13] ,
    \Tile_X9Y2_N4BEG[12] ,
    \Tile_X9Y2_N4BEG[11] ,
    \Tile_X9Y2_N4BEG[10] ,
    \Tile_X9Y2_N4BEG[9] ,
    \Tile_X9Y2_N4BEG[8] ,
    \Tile_X9Y2_N4BEG[7] ,
    \Tile_X9Y2_N4BEG[6] ,
    \Tile_X9Y2_N4BEG[5] ,
    \Tile_X9Y2_N4BEG[4] ,
    \Tile_X9Y2_N4BEG[3] ,
    \Tile_X9Y2_N4BEG[2] ,
    \Tile_X9Y2_N4BEG[1] ,
    \Tile_X9Y2_N4BEG[0] }),
    .NN4BEG({\Tile_X9Y1_NN4BEG[15] ,
    \Tile_X9Y1_NN4BEG[14] ,
    \Tile_X9Y1_NN4BEG[13] ,
    \Tile_X9Y1_NN4BEG[12] ,
    \Tile_X9Y1_NN4BEG[11] ,
    \Tile_X9Y1_NN4BEG[10] ,
    \Tile_X9Y1_NN4BEG[9] ,
    \Tile_X9Y1_NN4BEG[8] ,
    \Tile_X9Y1_NN4BEG[7] ,
    \Tile_X9Y1_NN4BEG[6] ,
    \Tile_X9Y1_NN4BEG[5] ,
    \Tile_X9Y1_NN4BEG[4] ,
    \Tile_X9Y1_NN4BEG[3] ,
    \Tile_X9Y1_NN4BEG[2] ,
    \Tile_X9Y1_NN4BEG[1] ,
    \Tile_X9Y1_NN4BEG[0] }),
    .NN4END({\Tile_X9Y2_NN4BEG[15] ,
    \Tile_X9Y2_NN4BEG[14] ,
    \Tile_X9Y2_NN4BEG[13] ,
    \Tile_X9Y2_NN4BEG[12] ,
    \Tile_X9Y2_NN4BEG[11] ,
    \Tile_X9Y2_NN4BEG[10] ,
    \Tile_X9Y2_NN4BEG[9] ,
    \Tile_X9Y2_NN4BEG[8] ,
    \Tile_X9Y2_NN4BEG[7] ,
    \Tile_X9Y2_NN4BEG[6] ,
    \Tile_X9Y2_NN4BEG[5] ,
    \Tile_X9Y2_NN4BEG[4] ,
    \Tile_X9Y2_NN4BEG[3] ,
    \Tile_X9Y2_NN4BEG[2] ,
    \Tile_X9Y2_NN4BEG[1] ,
    \Tile_X9Y2_NN4BEG[0] }),
    .S1BEG({\Tile_X9Y1_S1BEG[3] ,
    \Tile_X9Y1_S1BEG[2] ,
    \Tile_X9Y1_S1BEG[1] ,
    \Tile_X9Y1_S1BEG[0] }),
    .S1END({\Tile_X9Y0_S1BEG[3] ,
    \Tile_X9Y0_S1BEG[2] ,
    \Tile_X9Y0_S1BEG[1] ,
    \Tile_X9Y0_S1BEG[0] }),
    .S2BEG({\Tile_X9Y1_S2BEG[7] ,
    \Tile_X9Y1_S2BEG[6] ,
    \Tile_X9Y1_S2BEG[5] ,
    \Tile_X9Y1_S2BEG[4] ,
    \Tile_X9Y1_S2BEG[3] ,
    \Tile_X9Y1_S2BEG[2] ,
    \Tile_X9Y1_S2BEG[1] ,
    \Tile_X9Y1_S2BEG[0] }),
    .S2BEGb({\Tile_X9Y1_S2BEGb[7] ,
    \Tile_X9Y1_S2BEGb[6] ,
    \Tile_X9Y1_S2BEGb[5] ,
    \Tile_X9Y1_S2BEGb[4] ,
    \Tile_X9Y1_S2BEGb[3] ,
    \Tile_X9Y1_S2BEGb[2] ,
    \Tile_X9Y1_S2BEGb[1] ,
    \Tile_X9Y1_S2BEGb[0] }),
    .S2END({\Tile_X9Y0_S2BEGb[7] ,
    \Tile_X9Y0_S2BEGb[6] ,
    \Tile_X9Y0_S2BEGb[5] ,
    \Tile_X9Y0_S2BEGb[4] ,
    \Tile_X9Y0_S2BEGb[3] ,
    \Tile_X9Y0_S2BEGb[2] ,
    \Tile_X9Y0_S2BEGb[1] ,
    \Tile_X9Y0_S2BEGb[0] }),
    .S2MID({\Tile_X9Y0_S2BEG[7] ,
    \Tile_X9Y0_S2BEG[6] ,
    \Tile_X9Y0_S2BEG[5] ,
    \Tile_X9Y0_S2BEG[4] ,
    \Tile_X9Y0_S2BEG[3] ,
    \Tile_X9Y0_S2BEG[2] ,
    \Tile_X9Y0_S2BEG[1] ,
    \Tile_X9Y0_S2BEG[0] }),
    .S4BEG({\Tile_X9Y1_S4BEG[15] ,
    \Tile_X9Y1_S4BEG[14] ,
    \Tile_X9Y1_S4BEG[13] ,
    \Tile_X9Y1_S4BEG[12] ,
    \Tile_X9Y1_S4BEG[11] ,
    \Tile_X9Y1_S4BEG[10] ,
    \Tile_X9Y1_S4BEG[9] ,
    \Tile_X9Y1_S4BEG[8] ,
    \Tile_X9Y1_S4BEG[7] ,
    \Tile_X9Y1_S4BEG[6] ,
    \Tile_X9Y1_S4BEG[5] ,
    \Tile_X9Y1_S4BEG[4] ,
    \Tile_X9Y1_S4BEG[3] ,
    \Tile_X9Y1_S4BEG[2] ,
    \Tile_X9Y1_S4BEG[1] ,
    \Tile_X9Y1_S4BEG[0] }),
    .S4END({\Tile_X9Y0_S4BEG[15] ,
    \Tile_X9Y0_S4BEG[14] ,
    \Tile_X9Y0_S4BEG[13] ,
    \Tile_X9Y0_S4BEG[12] ,
    \Tile_X9Y0_S4BEG[11] ,
    \Tile_X9Y0_S4BEG[10] ,
    \Tile_X9Y0_S4BEG[9] ,
    \Tile_X9Y0_S4BEG[8] ,
    \Tile_X9Y0_S4BEG[7] ,
    \Tile_X9Y0_S4BEG[6] ,
    \Tile_X9Y0_S4BEG[5] ,
    \Tile_X9Y0_S4BEG[4] ,
    \Tile_X9Y0_S4BEG[3] ,
    \Tile_X9Y0_S4BEG[2] ,
    \Tile_X9Y0_S4BEG[1] ,
    \Tile_X9Y0_S4BEG[0] }),
    .SS4BEG({\Tile_X9Y1_SS4BEG[15] ,
    \Tile_X9Y1_SS4BEG[14] ,
    \Tile_X9Y1_SS4BEG[13] ,
    \Tile_X9Y1_SS4BEG[12] ,
    \Tile_X9Y1_SS4BEG[11] ,
    \Tile_X9Y1_SS4BEG[10] ,
    \Tile_X9Y1_SS4BEG[9] ,
    \Tile_X9Y1_SS4BEG[8] ,
    \Tile_X9Y1_SS4BEG[7] ,
    \Tile_X9Y1_SS4BEG[6] ,
    \Tile_X9Y1_SS4BEG[5] ,
    \Tile_X9Y1_SS4BEG[4] ,
    \Tile_X9Y1_SS4BEG[3] ,
    \Tile_X9Y1_SS4BEG[2] ,
    \Tile_X9Y1_SS4BEG[1] ,
    \Tile_X9Y1_SS4BEG[0] }),
    .SS4END({\Tile_X9Y0_SS4BEG[15] ,
    \Tile_X9Y0_SS4BEG[14] ,
    \Tile_X9Y0_SS4BEG[13] ,
    \Tile_X9Y0_SS4BEG[12] ,
    \Tile_X9Y0_SS4BEG[11] ,
    \Tile_X9Y0_SS4BEG[10] ,
    \Tile_X9Y0_SS4BEG[9] ,
    \Tile_X9Y0_SS4BEG[8] ,
    \Tile_X9Y0_SS4BEG[7] ,
    \Tile_X9Y0_SS4BEG[6] ,
    \Tile_X9Y0_SS4BEG[5] ,
    \Tile_X9Y0_SS4BEG[4] ,
    \Tile_X9Y0_SS4BEG[3] ,
    \Tile_X9Y0_SS4BEG[2] ,
    \Tile_X9Y0_SS4BEG[1] ,
    \Tile_X9Y0_SS4BEG[0] }),
    .W1BEG({\Tile_X9Y1_W1BEG[3] ,
    \Tile_X9Y1_W1BEG[2] ,
    \Tile_X9Y1_W1BEG[1] ,
    \Tile_X9Y1_W1BEG[0] }),
    .W1END({\Tile_X10Y1_W1BEG[3] ,
    \Tile_X10Y1_W1BEG[2] ,
    \Tile_X10Y1_W1BEG[1] ,
    \Tile_X10Y1_W1BEG[0] }),
    .W2BEG({\Tile_X9Y1_W2BEG[7] ,
    \Tile_X9Y1_W2BEG[6] ,
    \Tile_X9Y1_W2BEG[5] ,
    \Tile_X9Y1_W2BEG[4] ,
    \Tile_X9Y1_W2BEG[3] ,
    \Tile_X9Y1_W2BEG[2] ,
    \Tile_X9Y1_W2BEG[1] ,
    \Tile_X9Y1_W2BEG[0] }),
    .W2BEGb({\Tile_X9Y1_W2BEGb[7] ,
    \Tile_X9Y1_W2BEGb[6] ,
    \Tile_X9Y1_W2BEGb[5] ,
    \Tile_X9Y1_W2BEGb[4] ,
    \Tile_X9Y1_W2BEGb[3] ,
    \Tile_X9Y1_W2BEGb[2] ,
    \Tile_X9Y1_W2BEGb[1] ,
    \Tile_X9Y1_W2BEGb[0] }),
    .W2END({\Tile_X10Y1_W2BEGb[7] ,
    \Tile_X10Y1_W2BEGb[6] ,
    \Tile_X10Y1_W2BEGb[5] ,
    \Tile_X10Y1_W2BEGb[4] ,
    \Tile_X10Y1_W2BEGb[3] ,
    \Tile_X10Y1_W2BEGb[2] ,
    \Tile_X10Y1_W2BEGb[1] ,
    \Tile_X10Y1_W2BEGb[0] }),
    .W2MID({\Tile_X10Y1_W2BEG[7] ,
    \Tile_X10Y1_W2BEG[6] ,
    \Tile_X10Y1_W2BEG[5] ,
    \Tile_X10Y1_W2BEG[4] ,
    \Tile_X10Y1_W2BEG[3] ,
    \Tile_X10Y1_W2BEG[2] ,
    \Tile_X10Y1_W2BEG[1] ,
    \Tile_X10Y1_W2BEG[0] }),
    .W6BEG({\Tile_X9Y1_W6BEG[11] ,
    \Tile_X9Y1_W6BEG[10] ,
    \Tile_X9Y1_W6BEG[9] ,
    \Tile_X9Y1_W6BEG[8] ,
    \Tile_X9Y1_W6BEG[7] ,
    \Tile_X9Y1_W6BEG[6] ,
    \Tile_X9Y1_W6BEG[5] ,
    \Tile_X9Y1_W6BEG[4] ,
    \Tile_X9Y1_W6BEG[3] ,
    \Tile_X9Y1_W6BEG[2] ,
    \Tile_X9Y1_W6BEG[1] ,
    \Tile_X9Y1_W6BEG[0] }),
    .W6END({\Tile_X10Y1_W6BEG[11] ,
    \Tile_X10Y1_W6BEG[10] ,
    \Tile_X10Y1_W6BEG[9] ,
    \Tile_X10Y1_W6BEG[8] ,
    \Tile_X10Y1_W6BEG[7] ,
    \Tile_X10Y1_W6BEG[6] ,
    \Tile_X10Y1_W6BEG[5] ,
    \Tile_X10Y1_W6BEG[4] ,
    \Tile_X10Y1_W6BEG[3] ,
    \Tile_X10Y1_W6BEG[2] ,
    \Tile_X10Y1_W6BEG[1] ,
    \Tile_X10Y1_W6BEG[0] }),
    .WW4BEG({\Tile_X9Y1_WW4BEG[15] ,
    \Tile_X9Y1_WW4BEG[14] ,
    \Tile_X9Y1_WW4BEG[13] ,
    \Tile_X9Y1_WW4BEG[12] ,
    \Tile_X9Y1_WW4BEG[11] ,
    \Tile_X9Y1_WW4BEG[10] ,
    \Tile_X9Y1_WW4BEG[9] ,
    \Tile_X9Y1_WW4BEG[8] ,
    \Tile_X9Y1_WW4BEG[7] ,
    \Tile_X9Y1_WW4BEG[6] ,
    \Tile_X9Y1_WW4BEG[5] ,
    \Tile_X9Y1_WW4BEG[4] ,
    \Tile_X9Y1_WW4BEG[3] ,
    \Tile_X9Y1_WW4BEG[2] ,
    \Tile_X9Y1_WW4BEG[1] ,
    \Tile_X9Y1_WW4BEG[0] }),
    .WW4END({\Tile_X10Y1_WW4BEG[15] ,
    \Tile_X10Y1_WW4BEG[14] ,
    \Tile_X10Y1_WW4BEG[13] ,
    \Tile_X10Y1_WW4BEG[12] ,
    \Tile_X10Y1_WW4BEG[11] ,
    \Tile_X10Y1_WW4BEG[10] ,
    \Tile_X10Y1_WW4BEG[9] ,
    \Tile_X10Y1_WW4BEG[8] ,
    \Tile_X10Y1_WW4BEG[7] ,
    \Tile_X10Y1_WW4BEG[6] ,
    \Tile_X10Y1_WW4BEG[5] ,
    \Tile_X10Y1_WW4BEG[4] ,
    \Tile_X10Y1_WW4BEG[3] ,
    \Tile_X10Y1_WW4BEG[2] ,
    \Tile_X10Y1_WW4BEG[1] ,
    \Tile_X10Y1_WW4BEG[0] }));
 LUT4AB Tile_X9Y2_LUT4AB (.Ci(Tile_X9Y3_Co),
    .Co(Tile_X9Y2_Co),
    .UserCLK(Tile_X9Y3_UserCLKo),
    .UserCLKo(Tile_X9Y2_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X9Y2_E1BEG[3] ,
    \Tile_X9Y2_E1BEG[2] ,
    \Tile_X9Y2_E1BEG[1] ,
    \Tile_X9Y2_E1BEG[0] }),
    .E1END({\Tile_X8Y2_E1BEG[3] ,
    \Tile_X8Y2_E1BEG[2] ,
    \Tile_X8Y2_E1BEG[1] ,
    \Tile_X8Y2_E1BEG[0] }),
    .E2BEG({\Tile_X9Y2_E2BEG[7] ,
    \Tile_X9Y2_E2BEG[6] ,
    \Tile_X9Y2_E2BEG[5] ,
    \Tile_X9Y2_E2BEG[4] ,
    \Tile_X9Y2_E2BEG[3] ,
    \Tile_X9Y2_E2BEG[2] ,
    \Tile_X9Y2_E2BEG[1] ,
    \Tile_X9Y2_E2BEG[0] }),
    .E2BEGb({\Tile_X9Y2_E2BEGb[7] ,
    \Tile_X9Y2_E2BEGb[6] ,
    \Tile_X9Y2_E2BEGb[5] ,
    \Tile_X9Y2_E2BEGb[4] ,
    \Tile_X9Y2_E2BEGb[3] ,
    \Tile_X9Y2_E2BEGb[2] ,
    \Tile_X9Y2_E2BEGb[1] ,
    \Tile_X9Y2_E2BEGb[0] }),
    .E2END({\Tile_X8Y2_E2BEGb[7] ,
    \Tile_X8Y2_E2BEGb[6] ,
    \Tile_X8Y2_E2BEGb[5] ,
    \Tile_X8Y2_E2BEGb[4] ,
    \Tile_X8Y2_E2BEGb[3] ,
    \Tile_X8Y2_E2BEGb[2] ,
    \Tile_X8Y2_E2BEGb[1] ,
    \Tile_X8Y2_E2BEGb[0] }),
    .E2MID({\Tile_X8Y2_E2BEG[7] ,
    \Tile_X8Y2_E2BEG[6] ,
    \Tile_X8Y2_E2BEG[5] ,
    \Tile_X8Y2_E2BEG[4] ,
    \Tile_X8Y2_E2BEG[3] ,
    \Tile_X8Y2_E2BEG[2] ,
    \Tile_X8Y2_E2BEG[1] ,
    \Tile_X8Y2_E2BEG[0] }),
    .E6BEG({\Tile_X9Y2_E6BEG[11] ,
    \Tile_X9Y2_E6BEG[10] ,
    \Tile_X9Y2_E6BEG[9] ,
    \Tile_X9Y2_E6BEG[8] ,
    \Tile_X9Y2_E6BEG[7] ,
    \Tile_X9Y2_E6BEG[6] ,
    \Tile_X9Y2_E6BEG[5] ,
    \Tile_X9Y2_E6BEG[4] ,
    \Tile_X9Y2_E6BEG[3] ,
    \Tile_X9Y2_E6BEG[2] ,
    \Tile_X9Y2_E6BEG[1] ,
    \Tile_X9Y2_E6BEG[0] }),
    .E6END({\Tile_X8Y2_E6BEG[11] ,
    \Tile_X8Y2_E6BEG[10] ,
    \Tile_X8Y2_E6BEG[9] ,
    \Tile_X8Y2_E6BEG[8] ,
    \Tile_X8Y2_E6BEG[7] ,
    \Tile_X8Y2_E6BEG[6] ,
    \Tile_X8Y2_E6BEG[5] ,
    \Tile_X8Y2_E6BEG[4] ,
    \Tile_X8Y2_E6BEG[3] ,
    \Tile_X8Y2_E6BEG[2] ,
    \Tile_X8Y2_E6BEG[1] ,
    \Tile_X8Y2_E6BEG[0] }),
    .EE4BEG({\Tile_X9Y2_EE4BEG[15] ,
    \Tile_X9Y2_EE4BEG[14] ,
    \Tile_X9Y2_EE4BEG[13] ,
    \Tile_X9Y2_EE4BEG[12] ,
    \Tile_X9Y2_EE4BEG[11] ,
    \Tile_X9Y2_EE4BEG[10] ,
    \Tile_X9Y2_EE4BEG[9] ,
    \Tile_X9Y2_EE4BEG[8] ,
    \Tile_X9Y2_EE4BEG[7] ,
    \Tile_X9Y2_EE4BEG[6] ,
    \Tile_X9Y2_EE4BEG[5] ,
    \Tile_X9Y2_EE4BEG[4] ,
    \Tile_X9Y2_EE4BEG[3] ,
    \Tile_X9Y2_EE4BEG[2] ,
    \Tile_X9Y2_EE4BEG[1] ,
    \Tile_X9Y2_EE4BEG[0] }),
    .EE4END({\Tile_X8Y2_EE4BEG[15] ,
    \Tile_X8Y2_EE4BEG[14] ,
    \Tile_X8Y2_EE4BEG[13] ,
    \Tile_X8Y2_EE4BEG[12] ,
    \Tile_X8Y2_EE4BEG[11] ,
    \Tile_X8Y2_EE4BEG[10] ,
    \Tile_X8Y2_EE4BEG[9] ,
    \Tile_X8Y2_EE4BEG[8] ,
    \Tile_X8Y2_EE4BEG[7] ,
    \Tile_X8Y2_EE4BEG[6] ,
    \Tile_X8Y2_EE4BEG[5] ,
    \Tile_X8Y2_EE4BEG[4] ,
    \Tile_X8Y2_EE4BEG[3] ,
    \Tile_X8Y2_EE4BEG[2] ,
    \Tile_X8Y2_EE4BEG[1] ,
    \Tile_X8Y2_EE4BEG[0] }),
    .FrameData({\Tile_X8Y2_FrameData_O[31] ,
    \Tile_X8Y2_FrameData_O[30] ,
    \Tile_X8Y2_FrameData_O[29] ,
    \Tile_X8Y2_FrameData_O[28] ,
    \Tile_X8Y2_FrameData_O[27] ,
    \Tile_X8Y2_FrameData_O[26] ,
    \Tile_X8Y2_FrameData_O[25] ,
    \Tile_X8Y2_FrameData_O[24] ,
    \Tile_X8Y2_FrameData_O[23] ,
    \Tile_X8Y2_FrameData_O[22] ,
    \Tile_X8Y2_FrameData_O[21] ,
    \Tile_X8Y2_FrameData_O[20] ,
    \Tile_X8Y2_FrameData_O[19] ,
    \Tile_X8Y2_FrameData_O[18] ,
    \Tile_X8Y2_FrameData_O[17] ,
    \Tile_X8Y2_FrameData_O[16] ,
    \Tile_X8Y2_FrameData_O[15] ,
    \Tile_X8Y2_FrameData_O[14] ,
    \Tile_X8Y2_FrameData_O[13] ,
    \Tile_X8Y2_FrameData_O[12] ,
    \Tile_X8Y2_FrameData_O[11] ,
    \Tile_X8Y2_FrameData_O[10] ,
    \Tile_X8Y2_FrameData_O[9] ,
    \Tile_X8Y2_FrameData_O[8] ,
    \Tile_X8Y2_FrameData_O[7] ,
    \Tile_X8Y2_FrameData_O[6] ,
    \Tile_X8Y2_FrameData_O[5] ,
    \Tile_X8Y2_FrameData_O[4] ,
    \Tile_X8Y2_FrameData_O[3] ,
    \Tile_X8Y2_FrameData_O[2] ,
    \Tile_X8Y2_FrameData_O[1] ,
    \Tile_X8Y2_FrameData_O[0] }),
    .FrameData_O({\Tile_X9Y2_FrameData_O[31] ,
    \Tile_X9Y2_FrameData_O[30] ,
    \Tile_X9Y2_FrameData_O[29] ,
    \Tile_X9Y2_FrameData_O[28] ,
    \Tile_X9Y2_FrameData_O[27] ,
    \Tile_X9Y2_FrameData_O[26] ,
    \Tile_X9Y2_FrameData_O[25] ,
    \Tile_X9Y2_FrameData_O[24] ,
    \Tile_X9Y2_FrameData_O[23] ,
    \Tile_X9Y2_FrameData_O[22] ,
    \Tile_X9Y2_FrameData_O[21] ,
    \Tile_X9Y2_FrameData_O[20] ,
    \Tile_X9Y2_FrameData_O[19] ,
    \Tile_X9Y2_FrameData_O[18] ,
    \Tile_X9Y2_FrameData_O[17] ,
    \Tile_X9Y2_FrameData_O[16] ,
    \Tile_X9Y2_FrameData_O[15] ,
    \Tile_X9Y2_FrameData_O[14] ,
    \Tile_X9Y2_FrameData_O[13] ,
    \Tile_X9Y2_FrameData_O[12] ,
    \Tile_X9Y2_FrameData_O[11] ,
    \Tile_X9Y2_FrameData_O[10] ,
    \Tile_X9Y2_FrameData_O[9] ,
    \Tile_X9Y2_FrameData_O[8] ,
    \Tile_X9Y2_FrameData_O[7] ,
    \Tile_X9Y2_FrameData_O[6] ,
    \Tile_X9Y2_FrameData_O[5] ,
    \Tile_X9Y2_FrameData_O[4] ,
    \Tile_X9Y2_FrameData_O[3] ,
    \Tile_X9Y2_FrameData_O[2] ,
    \Tile_X9Y2_FrameData_O[1] ,
    \Tile_X9Y2_FrameData_O[0] }),
    .FrameStrobe({\Tile_X9Y3_FrameStrobe_O[19] ,
    \Tile_X9Y3_FrameStrobe_O[18] ,
    \Tile_X9Y3_FrameStrobe_O[17] ,
    \Tile_X9Y3_FrameStrobe_O[16] ,
    \Tile_X9Y3_FrameStrobe_O[15] ,
    \Tile_X9Y3_FrameStrobe_O[14] ,
    \Tile_X9Y3_FrameStrobe_O[13] ,
    \Tile_X9Y3_FrameStrobe_O[12] ,
    \Tile_X9Y3_FrameStrobe_O[11] ,
    \Tile_X9Y3_FrameStrobe_O[10] ,
    \Tile_X9Y3_FrameStrobe_O[9] ,
    \Tile_X9Y3_FrameStrobe_O[8] ,
    \Tile_X9Y3_FrameStrobe_O[7] ,
    \Tile_X9Y3_FrameStrobe_O[6] ,
    \Tile_X9Y3_FrameStrobe_O[5] ,
    \Tile_X9Y3_FrameStrobe_O[4] ,
    \Tile_X9Y3_FrameStrobe_O[3] ,
    \Tile_X9Y3_FrameStrobe_O[2] ,
    \Tile_X9Y3_FrameStrobe_O[1] ,
    \Tile_X9Y3_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X9Y2_FrameStrobe_O[19] ,
    \Tile_X9Y2_FrameStrobe_O[18] ,
    \Tile_X9Y2_FrameStrobe_O[17] ,
    \Tile_X9Y2_FrameStrobe_O[16] ,
    \Tile_X9Y2_FrameStrobe_O[15] ,
    \Tile_X9Y2_FrameStrobe_O[14] ,
    \Tile_X9Y2_FrameStrobe_O[13] ,
    \Tile_X9Y2_FrameStrobe_O[12] ,
    \Tile_X9Y2_FrameStrobe_O[11] ,
    \Tile_X9Y2_FrameStrobe_O[10] ,
    \Tile_X9Y2_FrameStrobe_O[9] ,
    \Tile_X9Y2_FrameStrobe_O[8] ,
    \Tile_X9Y2_FrameStrobe_O[7] ,
    \Tile_X9Y2_FrameStrobe_O[6] ,
    \Tile_X9Y2_FrameStrobe_O[5] ,
    \Tile_X9Y2_FrameStrobe_O[4] ,
    \Tile_X9Y2_FrameStrobe_O[3] ,
    \Tile_X9Y2_FrameStrobe_O[2] ,
    \Tile_X9Y2_FrameStrobe_O[1] ,
    \Tile_X9Y2_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X9Y2_N1BEG[3] ,
    \Tile_X9Y2_N1BEG[2] ,
    \Tile_X9Y2_N1BEG[1] ,
    \Tile_X9Y2_N1BEG[0] }),
    .N1END({\Tile_X9Y3_N1BEG[3] ,
    \Tile_X9Y3_N1BEG[2] ,
    \Tile_X9Y3_N1BEG[1] ,
    \Tile_X9Y3_N1BEG[0] }),
    .N2BEG({\Tile_X9Y2_N2BEG[7] ,
    \Tile_X9Y2_N2BEG[6] ,
    \Tile_X9Y2_N2BEG[5] ,
    \Tile_X9Y2_N2BEG[4] ,
    \Tile_X9Y2_N2BEG[3] ,
    \Tile_X9Y2_N2BEG[2] ,
    \Tile_X9Y2_N2BEG[1] ,
    \Tile_X9Y2_N2BEG[0] }),
    .N2BEGb({\Tile_X9Y2_N2BEGb[7] ,
    \Tile_X9Y2_N2BEGb[6] ,
    \Tile_X9Y2_N2BEGb[5] ,
    \Tile_X9Y2_N2BEGb[4] ,
    \Tile_X9Y2_N2BEGb[3] ,
    \Tile_X9Y2_N2BEGb[2] ,
    \Tile_X9Y2_N2BEGb[1] ,
    \Tile_X9Y2_N2BEGb[0] }),
    .N2END({\Tile_X9Y3_N2BEGb[7] ,
    \Tile_X9Y3_N2BEGb[6] ,
    \Tile_X9Y3_N2BEGb[5] ,
    \Tile_X9Y3_N2BEGb[4] ,
    \Tile_X9Y3_N2BEGb[3] ,
    \Tile_X9Y3_N2BEGb[2] ,
    \Tile_X9Y3_N2BEGb[1] ,
    \Tile_X9Y3_N2BEGb[0] }),
    .N2MID({\Tile_X9Y3_N2BEG[7] ,
    \Tile_X9Y3_N2BEG[6] ,
    \Tile_X9Y3_N2BEG[5] ,
    \Tile_X9Y3_N2BEG[4] ,
    \Tile_X9Y3_N2BEG[3] ,
    \Tile_X9Y3_N2BEG[2] ,
    \Tile_X9Y3_N2BEG[1] ,
    \Tile_X9Y3_N2BEG[0] }),
    .N4BEG({\Tile_X9Y2_N4BEG[15] ,
    \Tile_X9Y2_N4BEG[14] ,
    \Tile_X9Y2_N4BEG[13] ,
    \Tile_X9Y2_N4BEG[12] ,
    \Tile_X9Y2_N4BEG[11] ,
    \Tile_X9Y2_N4BEG[10] ,
    \Tile_X9Y2_N4BEG[9] ,
    \Tile_X9Y2_N4BEG[8] ,
    \Tile_X9Y2_N4BEG[7] ,
    \Tile_X9Y2_N4BEG[6] ,
    \Tile_X9Y2_N4BEG[5] ,
    \Tile_X9Y2_N4BEG[4] ,
    \Tile_X9Y2_N4BEG[3] ,
    \Tile_X9Y2_N4BEG[2] ,
    \Tile_X9Y2_N4BEG[1] ,
    \Tile_X9Y2_N4BEG[0] }),
    .N4END({\Tile_X9Y3_N4BEG[15] ,
    \Tile_X9Y3_N4BEG[14] ,
    \Tile_X9Y3_N4BEG[13] ,
    \Tile_X9Y3_N4BEG[12] ,
    \Tile_X9Y3_N4BEG[11] ,
    \Tile_X9Y3_N4BEG[10] ,
    \Tile_X9Y3_N4BEG[9] ,
    \Tile_X9Y3_N4BEG[8] ,
    \Tile_X9Y3_N4BEG[7] ,
    \Tile_X9Y3_N4BEG[6] ,
    \Tile_X9Y3_N4BEG[5] ,
    \Tile_X9Y3_N4BEG[4] ,
    \Tile_X9Y3_N4BEG[3] ,
    \Tile_X9Y3_N4BEG[2] ,
    \Tile_X9Y3_N4BEG[1] ,
    \Tile_X9Y3_N4BEG[0] }),
    .NN4BEG({\Tile_X9Y2_NN4BEG[15] ,
    \Tile_X9Y2_NN4BEG[14] ,
    \Tile_X9Y2_NN4BEG[13] ,
    \Tile_X9Y2_NN4BEG[12] ,
    \Tile_X9Y2_NN4BEG[11] ,
    \Tile_X9Y2_NN4BEG[10] ,
    \Tile_X9Y2_NN4BEG[9] ,
    \Tile_X9Y2_NN4BEG[8] ,
    \Tile_X9Y2_NN4BEG[7] ,
    \Tile_X9Y2_NN4BEG[6] ,
    \Tile_X9Y2_NN4BEG[5] ,
    \Tile_X9Y2_NN4BEG[4] ,
    \Tile_X9Y2_NN4BEG[3] ,
    \Tile_X9Y2_NN4BEG[2] ,
    \Tile_X9Y2_NN4BEG[1] ,
    \Tile_X9Y2_NN4BEG[0] }),
    .NN4END({\Tile_X9Y3_NN4BEG[15] ,
    \Tile_X9Y3_NN4BEG[14] ,
    \Tile_X9Y3_NN4BEG[13] ,
    \Tile_X9Y3_NN4BEG[12] ,
    \Tile_X9Y3_NN4BEG[11] ,
    \Tile_X9Y3_NN4BEG[10] ,
    \Tile_X9Y3_NN4BEG[9] ,
    \Tile_X9Y3_NN4BEG[8] ,
    \Tile_X9Y3_NN4BEG[7] ,
    \Tile_X9Y3_NN4BEG[6] ,
    \Tile_X9Y3_NN4BEG[5] ,
    \Tile_X9Y3_NN4BEG[4] ,
    \Tile_X9Y3_NN4BEG[3] ,
    \Tile_X9Y3_NN4BEG[2] ,
    \Tile_X9Y3_NN4BEG[1] ,
    \Tile_X9Y3_NN4BEG[0] }),
    .S1BEG({\Tile_X9Y2_S1BEG[3] ,
    \Tile_X9Y2_S1BEG[2] ,
    \Tile_X9Y2_S1BEG[1] ,
    \Tile_X9Y2_S1BEG[0] }),
    .S1END({\Tile_X9Y1_S1BEG[3] ,
    \Tile_X9Y1_S1BEG[2] ,
    \Tile_X9Y1_S1BEG[1] ,
    \Tile_X9Y1_S1BEG[0] }),
    .S2BEG({\Tile_X9Y2_S2BEG[7] ,
    \Tile_X9Y2_S2BEG[6] ,
    \Tile_X9Y2_S2BEG[5] ,
    \Tile_X9Y2_S2BEG[4] ,
    \Tile_X9Y2_S2BEG[3] ,
    \Tile_X9Y2_S2BEG[2] ,
    \Tile_X9Y2_S2BEG[1] ,
    \Tile_X9Y2_S2BEG[0] }),
    .S2BEGb({\Tile_X9Y2_S2BEGb[7] ,
    \Tile_X9Y2_S2BEGb[6] ,
    \Tile_X9Y2_S2BEGb[5] ,
    \Tile_X9Y2_S2BEGb[4] ,
    \Tile_X9Y2_S2BEGb[3] ,
    \Tile_X9Y2_S2BEGb[2] ,
    \Tile_X9Y2_S2BEGb[1] ,
    \Tile_X9Y2_S2BEGb[0] }),
    .S2END({\Tile_X9Y1_S2BEGb[7] ,
    \Tile_X9Y1_S2BEGb[6] ,
    \Tile_X9Y1_S2BEGb[5] ,
    \Tile_X9Y1_S2BEGb[4] ,
    \Tile_X9Y1_S2BEGb[3] ,
    \Tile_X9Y1_S2BEGb[2] ,
    \Tile_X9Y1_S2BEGb[1] ,
    \Tile_X9Y1_S2BEGb[0] }),
    .S2MID({\Tile_X9Y1_S2BEG[7] ,
    \Tile_X9Y1_S2BEG[6] ,
    \Tile_X9Y1_S2BEG[5] ,
    \Tile_X9Y1_S2BEG[4] ,
    \Tile_X9Y1_S2BEG[3] ,
    \Tile_X9Y1_S2BEG[2] ,
    \Tile_X9Y1_S2BEG[1] ,
    \Tile_X9Y1_S2BEG[0] }),
    .S4BEG({\Tile_X9Y2_S4BEG[15] ,
    \Tile_X9Y2_S4BEG[14] ,
    \Tile_X9Y2_S4BEG[13] ,
    \Tile_X9Y2_S4BEG[12] ,
    \Tile_X9Y2_S4BEG[11] ,
    \Tile_X9Y2_S4BEG[10] ,
    \Tile_X9Y2_S4BEG[9] ,
    \Tile_X9Y2_S4BEG[8] ,
    \Tile_X9Y2_S4BEG[7] ,
    \Tile_X9Y2_S4BEG[6] ,
    \Tile_X9Y2_S4BEG[5] ,
    \Tile_X9Y2_S4BEG[4] ,
    \Tile_X9Y2_S4BEG[3] ,
    \Tile_X9Y2_S4BEG[2] ,
    \Tile_X9Y2_S4BEG[1] ,
    \Tile_X9Y2_S4BEG[0] }),
    .S4END({\Tile_X9Y1_S4BEG[15] ,
    \Tile_X9Y1_S4BEG[14] ,
    \Tile_X9Y1_S4BEG[13] ,
    \Tile_X9Y1_S4BEG[12] ,
    \Tile_X9Y1_S4BEG[11] ,
    \Tile_X9Y1_S4BEG[10] ,
    \Tile_X9Y1_S4BEG[9] ,
    \Tile_X9Y1_S4BEG[8] ,
    \Tile_X9Y1_S4BEG[7] ,
    \Tile_X9Y1_S4BEG[6] ,
    \Tile_X9Y1_S4BEG[5] ,
    \Tile_X9Y1_S4BEG[4] ,
    \Tile_X9Y1_S4BEG[3] ,
    \Tile_X9Y1_S4BEG[2] ,
    \Tile_X9Y1_S4BEG[1] ,
    \Tile_X9Y1_S4BEG[0] }),
    .SS4BEG({\Tile_X9Y2_SS4BEG[15] ,
    \Tile_X9Y2_SS4BEG[14] ,
    \Tile_X9Y2_SS4BEG[13] ,
    \Tile_X9Y2_SS4BEG[12] ,
    \Tile_X9Y2_SS4BEG[11] ,
    \Tile_X9Y2_SS4BEG[10] ,
    \Tile_X9Y2_SS4BEG[9] ,
    \Tile_X9Y2_SS4BEG[8] ,
    \Tile_X9Y2_SS4BEG[7] ,
    \Tile_X9Y2_SS4BEG[6] ,
    \Tile_X9Y2_SS4BEG[5] ,
    \Tile_X9Y2_SS4BEG[4] ,
    \Tile_X9Y2_SS4BEG[3] ,
    \Tile_X9Y2_SS4BEG[2] ,
    \Tile_X9Y2_SS4BEG[1] ,
    \Tile_X9Y2_SS4BEG[0] }),
    .SS4END({\Tile_X9Y1_SS4BEG[15] ,
    \Tile_X9Y1_SS4BEG[14] ,
    \Tile_X9Y1_SS4BEG[13] ,
    \Tile_X9Y1_SS4BEG[12] ,
    \Tile_X9Y1_SS4BEG[11] ,
    \Tile_X9Y1_SS4BEG[10] ,
    \Tile_X9Y1_SS4BEG[9] ,
    \Tile_X9Y1_SS4BEG[8] ,
    \Tile_X9Y1_SS4BEG[7] ,
    \Tile_X9Y1_SS4BEG[6] ,
    \Tile_X9Y1_SS4BEG[5] ,
    \Tile_X9Y1_SS4BEG[4] ,
    \Tile_X9Y1_SS4BEG[3] ,
    \Tile_X9Y1_SS4BEG[2] ,
    \Tile_X9Y1_SS4BEG[1] ,
    \Tile_X9Y1_SS4BEG[0] }),
    .W1BEG({\Tile_X9Y2_W1BEG[3] ,
    \Tile_X9Y2_W1BEG[2] ,
    \Tile_X9Y2_W1BEG[1] ,
    \Tile_X9Y2_W1BEG[0] }),
    .W1END({\Tile_X10Y2_W1BEG[3] ,
    \Tile_X10Y2_W1BEG[2] ,
    \Tile_X10Y2_W1BEG[1] ,
    \Tile_X10Y2_W1BEG[0] }),
    .W2BEG({\Tile_X9Y2_W2BEG[7] ,
    \Tile_X9Y2_W2BEG[6] ,
    \Tile_X9Y2_W2BEG[5] ,
    \Tile_X9Y2_W2BEG[4] ,
    \Tile_X9Y2_W2BEG[3] ,
    \Tile_X9Y2_W2BEG[2] ,
    \Tile_X9Y2_W2BEG[1] ,
    \Tile_X9Y2_W2BEG[0] }),
    .W2BEGb({\Tile_X9Y2_W2BEGb[7] ,
    \Tile_X9Y2_W2BEGb[6] ,
    \Tile_X9Y2_W2BEGb[5] ,
    \Tile_X9Y2_W2BEGb[4] ,
    \Tile_X9Y2_W2BEGb[3] ,
    \Tile_X9Y2_W2BEGb[2] ,
    \Tile_X9Y2_W2BEGb[1] ,
    \Tile_X9Y2_W2BEGb[0] }),
    .W2END({\Tile_X10Y2_W2BEGb[7] ,
    \Tile_X10Y2_W2BEGb[6] ,
    \Tile_X10Y2_W2BEGb[5] ,
    \Tile_X10Y2_W2BEGb[4] ,
    \Tile_X10Y2_W2BEGb[3] ,
    \Tile_X10Y2_W2BEGb[2] ,
    \Tile_X10Y2_W2BEGb[1] ,
    \Tile_X10Y2_W2BEGb[0] }),
    .W2MID({\Tile_X10Y2_W2BEG[7] ,
    \Tile_X10Y2_W2BEG[6] ,
    \Tile_X10Y2_W2BEG[5] ,
    \Tile_X10Y2_W2BEG[4] ,
    \Tile_X10Y2_W2BEG[3] ,
    \Tile_X10Y2_W2BEG[2] ,
    \Tile_X10Y2_W2BEG[1] ,
    \Tile_X10Y2_W2BEG[0] }),
    .W6BEG({\Tile_X9Y2_W6BEG[11] ,
    \Tile_X9Y2_W6BEG[10] ,
    \Tile_X9Y2_W6BEG[9] ,
    \Tile_X9Y2_W6BEG[8] ,
    \Tile_X9Y2_W6BEG[7] ,
    \Tile_X9Y2_W6BEG[6] ,
    \Tile_X9Y2_W6BEG[5] ,
    \Tile_X9Y2_W6BEG[4] ,
    \Tile_X9Y2_W6BEG[3] ,
    \Tile_X9Y2_W6BEG[2] ,
    \Tile_X9Y2_W6BEG[1] ,
    \Tile_X9Y2_W6BEG[0] }),
    .W6END({\Tile_X10Y2_W6BEG[11] ,
    \Tile_X10Y2_W6BEG[10] ,
    \Tile_X10Y2_W6BEG[9] ,
    \Tile_X10Y2_W6BEG[8] ,
    \Tile_X10Y2_W6BEG[7] ,
    \Tile_X10Y2_W6BEG[6] ,
    \Tile_X10Y2_W6BEG[5] ,
    \Tile_X10Y2_W6BEG[4] ,
    \Tile_X10Y2_W6BEG[3] ,
    \Tile_X10Y2_W6BEG[2] ,
    \Tile_X10Y2_W6BEG[1] ,
    \Tile_X10Y2_W6BEG[0] }),
    .WW4BEG({\Tile_X9Y2_WW4BEG[15] ,
    \Tile_X9Y2_WW4BEG[14] ,
    \Tile_X9Y2_WW4BEG[13] ,
    \Tile_X9Y2_WW4BEG[12] ,
    \Tile_X9Y2_WW4BEG[11] ,
    \Tile_X9Y2_WW4BEG[10] ,
    \Tile_X9Y2_WW4BEG[9] ,
    \Tile_X9Y2_WW4BEG[8] ,
    \Tile_X9Y2_WW4BEG[7] ,
    \Tile_X9Y2_WW4BEG[6] ,
    \Tile_X9Y2_WW4BEG[5] ,
    \Tile_X9Y2_WW4BEG[4] ,
    \Tile_X9Y2_WW4BEG[3] ,
    \Tile_X9Y2_WW4BEG[2] ,
    \Tile_X9Y2_WW4BEG[1] ,
    \Tile_X9Y2_WW4BEG[0] }),
    .WW4END({\Tile_X10Y2_WW4BEG[15] ,
    \Tile_X10Y2_WW4BEG[14] ,
    \Tile_X10Y2_WW4BEG[13] ,
    \Tile_X10Y2_WW4BEG[12] ,
    \Tile_X10Y2_WW4BEG[11] ,
    \Tile_X10Y2_WW4BEG[10] ,
    \Tile_X10Y2_WW4BEG[9] ,
    \Tile_X10Y2_WW4BEG[8] ,
    \Tile_X10Y2_WW4BEG[7] ,
    \Tile_X10Y2_WW4BEG[6] ,
    \Tile_X10Y2_WW4BEG[5] ,
    \Tile_X10Y2_WW4BEG[4] ,
    \Tile_X10Y2_WW4BEG[3] ,
    \Tile_X10Y2_WW4BEG[2] ,
    \Tile_X10Y2_WW4BEG[1] ,
    \Tile_X10Y2_WW4BEG[0] }));
 LUT4AB Tile_X9Y3_LUT4AB (.Ci(Tile_X9Y4_Co),
    .Co(Tile_X9Y3_Co),
    .UserCLK(Tile_X9Y4_UserCLKo),
    .UserCLKo(Tile_X9Y3_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X9Y3_E1BEG[3] ,
    \Tile_X9Y3_E1BEG[2] ,
    \Tile_X9Y3_E1BEG[1] ,
    \Tile_X9Y3_E1BEG[0] }),
    .E1END({\Tile_X8Y3_E1BEG[3] ,
    \Tile_X8Y3_E1BEG[2] ,
    \Tile_X8Y3_E1BEG[1] ,
    \Tile_X8Y3_E1BEG[0] }),
    .E2BEG({\Tile_X9Y3_E2BEG[7] ,
    \Tile_X9Y3_E2BEG[6] ,
    \Tile_X9Y3_E2BEG[5] ,
    \Tile_X9Y3_E2BEG[4] ,
    \Tile_X9Y3_E2BEG[3] ,
    \Tile_X9Y3_E2BEG[2] ,
    \Tile_X9Y3_E2BEG[1] ,
    \Tile_X9Y3_E2BEG[0] }),
    .E2BEGb({\Tile_X9Y3_E2BEGb[7] ,
    \Tile_X9Y3_E2BEGb[6] ,
    \Tile_X9Y3_E2BEGb[5] ,
    \Tile_X9Y3_E2BEGb[4] ,
    \Tile_X9Y3_E2BEGb[3] ,
    \Tile_X9Y3_E2BEGb[2] ,
    \Tile_X9Y3_E2BEGb[1] ,
    \Tile_X9Y3_E2BEGb[0] }),
    .E2END({\Tile_X8Y3_E2BEGb[7] ,
    \Tile_X8Y3_E2BEGb[6] ,
    \Tile_X8Y3_E2BEGb[5] ,
    \Tile_X8Y3_E2BEGb[4] ,
    \Tile_X8Y3_E2BEGb[3] ,
    \Tile_X8Y3_E2BEGb[2] ,
    \Tile_X8Y3_E2BEGb[1] ,
    \Tile_X8Y3_E2BEGb[0] }),
    .E2MID({\Tile_X8Y3_E2BEG[7] ,
    \Tile_X8Y3_E2BEG[6] ,
    \Tile_X8Y3_E2BEG[5] ,
    \Tile_X8Y3_E2BEG[4] ,
    \Tile_X8Y3_E2BEG[3] ,
    \Tile_X8Y3_E2BEG[2] ,
    \Tile_X8Y3_E2BEG[1] ,
    \Tile_X8Y3_E2BEG[0] }),
    .E6BEG({\Tile_X9Y3_E6BEG[11] ,
    \Tile_X9Y3_E6BEG[10] ,
    \Tile_X9Y3_E6BEG[9] ,
    \Tile_X9Y3_E6BEG[8] ,
    \Tile_X9Y3_E6BEG[7] ,
    \Tile_X9Y3_E6BEG[6] ,
    \Tile_X9Y3_E6BEG[5] ,
    \Tile_X9Y3_E6BEG[4] ,
    \Tile_X9Y3_E6BEG[3] ,
    \Tile_X9Y3_E6BEG[2] ,
    \Tile_X9Y3_E6BEG[1] ,
    \Tile_X9Y3_E6BEG[0] }),
    .E6END({\Tile_X8Y3_E6BEG[11] ,
    \Tile_X8Y3_E6BEG[10] ,
    \Tile_X8Y3_E6BEG[9] ,
    \Tile_X8Y3_E6BEG[8] ,
    \Tile_X8Y3_E6BEG[7] ,
    \Tile_X8Y3_E6BEG[6] ,
    \Tile_X8Y3_E6BEG[5] ,
    \Tile_X8Y3_E6BEG[4] ,
    \Tile_X8Y3_E6BEG[3] ,
    \Tile_X8Y3_E6BEG[2] ,
    \Tile_X8Y3_E6BEG[1] ,
    \Tile_X8Y3_E6BEG[0] }),
    .EE4BEG({\Tile_X9Y3_EE4BEG[15] ,
    \Tile_X9Y3_EE4BEG[14] ,
    \Tile_X9Y3_EE4BEG[13] ,
    \Tile_X9Y3_EE4BEG[12] ,
    \Tile_X9Y3_EE4BEG[11] ,
    \Tile_X9Y3_EE4BEG[10] ,
    \Tile_X9Y3_EE4BEG[9] ,
    \Tile_X9Y3_EE4BEG[8] ,
    \Tile_X9Y3_EE4BEG[7] ,
    \Tile_X9Y3_EE4BEG[6] ,
    \Tile_X9Y3_EE4BEG[5] ,
    \Tile_X9Y3_EE4BEG[4] ,
    \Tile_X9Y3_EE4BEG[3] ,
    \Tile_X9Y3_EE4BEG[2] ,
    \Tile_X9Y3_EE4BEG[1] ,
    \Tile_X9Y3_EE4BEG[0] }),
    .EE4END({\Tile_X8Y3_EE4BEG[15] ,
    \Tile_X8Y3_EE4BEG[14] ,
    \Tile_X8Y3_EE4BEG[13] ,
    \Tile_X8Y3_EE4BEG[12] ,
    \Tile_X8Y3_EE4BEG[11] ,
    \Tile_X8Y3_EE4BEG[10] ,
    \Tile_X8Y3_EE4BEG[9] ,
    \Tile_X8Y3_EE4BEG[8] ,
    \Tile_X8Y3_EE4BEG[7] ,
    \Tile_X8Y3_EE4BEG[6] ,
    \Tile_X8Y3_EE4BEG[5] ,
    \Tile_X8Y3_EE4BEG[4] ,
    \Tile_X8Y3_EE4BEG[3] ,
    \Tile_X8Y3_EE4BEG[2] ,
    \Tile_X8Y3_EE4BEG[1] ,
    \Tile_X8Y3_EE4BEG[0] }),
    .FrameData({\Tile_X8Y3_FrameData_O[31] ,
    \Tile_X8Y3_FrameData_O[30] ,
    \Tile_X8Y3_FrameData_O[29] ,
    \Tile_X8Y3_FrameData_O[28] ,
    \Tile_X8Y3_FrameData_O[27] ,
    \Tile_X8Y3_FrameData_O[26] ,
    \Tile_X8Y3_FrameData_O[25] ,
    \Tile_X8Y3_FrameData_O[24] ,
    \Tile_X8Y3_FrameData_O[23] ,
    \Tile_X8Y3_FrameData_O[22] ,
    \Tile_X8Y3_FrameData_O[21] ,
    \Tile_X8Y3_FrameData_O[20] ,
    \Tile_X8Y3_FrameData_O[19] ,
    \Tile_X8Y3_FrameData_O[18] ,
    \Tile_X8Y3_FrameData_O[17] ,
    \Tile_X8Y3_FrameData_O[16] ,
    \Tile_X8Y3_FrameData_O[15] ,
    \Tile_X8Y3_FrameData_O[14] ,
    \Tile_X8Y3_FrameData_O[13] ,
    \Tile_X8Y3_FrameData_O[12] ,
    \Tile_X8Y3_FrameData_O[11] ,
    \Tile_X8Y3_FrameData_O[10] ,
    \Tile_X8Y3_FrameData_O[9] ,
    \Tile_X8Y3_FrameData_O[8] ,
    \Tile_X8Y3_FrameData_O[7] ,
    \Tile_X8Y3_FrameData_O[6] ,
    \Tile_X8Y3_FrameData_O[5] ,
    \Tile_X8Y3_FrameData_O[4] ,
    \Tile_X8Y3_FrameData_O[3] ,
    \Tile_X8Y3_FrameData_O[2] ,
    \Tile_X8Y3_FrameData_O[1] ,
    \Tile_X8Y3_FrameData_O[0] }),
    .FrameData_O({\Tile_X9Y3_FrameData_O[31] ,
    \Tile_X9Y3_FrameData_O[30] ,
    \Tile_X9Y3_FrameData_O[29] ,
    \Tile_X9Y3_FrameData_O[28] ,
    \Tile_X9Y3_FrameData_O[27] ,
    \Tile_X9Y3_FrameData_O[26] ,
    \Tile_X9Y3_FrameData_O[25] ,
    \Tile_X9Y3_FrameData_O[24] ,
    \Tile_X9Y3_FrameData_O[23] ,
    \Tile_X9Y3_FrameData_O[22] ,
    \Tile_X9Y3_FrameData_O[21] ,
    \Tile_X9Y3_FrameData_O[20] ,
    \Tile_X9Y3_FrameData_O[19] ,
    \Tile_X9Y3_FrameData_O[18] ,
    \Tile_X9Y3_FrameData_O[17] ,
    \Tile_X9Y3_FrameData_O[16] ,
    \Tile_X9Y3_FrameData_O[15] ,
    \Tile_X9Y3_FrameData_O[14] ,
    \Tile_X9Y3_FrameData_O[13] ,
    \Tile_X9Y3_FrameData_O[12] ,
    \Tile_X9Y3_FrameData_O[11] ,
    \Tile_X9Y3_FrameData_O[10] ,
    \Tile_X9Y3_FrameData_O[9] ,
    \Tile_X9Y3_FrameData_O[8] ,
    \Tile_X9Y3_FrameData_O[7] ,
    \Tile_X9Y3_FrameData_O[6] ,
    \Tile_X9Y3_FrameData_O[5] ,
    \Tile_X9Y3_FrameData_O[4] ,
    \Tile_X9Y3_FrameData_O[3] ,
    \Tile_X9Y3_FrameData_O[2] ,
    \Tile_X9Y3_FrameData_O[1] ,
    \Tile_X9Y3_FrameData_O[0] }),
    .FrameStrobe({\Tile_X9Y4_FrameStrobe_O[19] ,
    \Tile_X9Y4_FrameStrobe_O[18] ,
    \Tile_X9Y4_FrameStrobe_O[17] ,
    \Tile_X9Y4_FrameStrobe_O[16] ,
    \Tile_X9Y4_FrameStrobe_O[15] ,
    \Tile_X9Y4_FrameStrobe_O[14] ,
    \Tile_X9Y4_FrameStrobe_O[13] ,
    \Tile_X9Y4_FrameStrobe_O[12] ,
    \Tile_X9Y4_FrameStrobe_O[11] ,
    \Tile_X9Y4_FrameStrobe_O[10] ,
    \Tile_X9Y4_FrameStrobe_O[9] ,
    \Tile_X9Y4_FrameStrobe_O[8] ,
    \Tile_X9Y4_FrameStrobe_O[7] ,
    \Tile_X9Y4_FrameStrobe_O[6] ,
    \Tile_X9Y4_FrameStrobe_O[5] ,
    \Tile_X9Y4_FrameStrobe_O[4] ,
    \Tile_X9Y4_FrameStrobe_O[3] ,
    \Tile_X9Y4_FrameStrobe_O[2] ,
    \Tile_X9Y4_FrameStrobe_O[1] ,
    \Tile_X9Y4_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X9Y3_FrameStrobe_O[19] ,
    \Tile_X9Y3_FrameStrobe_O[18] ,
    \Tile_X9Y3_FrameStrobe_O[17] ,
    \Tile_X9Y3_FrameStrobe_O[16] ,
    \Tile_X9Y3_FrameStrobe_O[15] ,
    \Tile_X9Y3_FrameStrobe_O[14] ,
    \Tile_X9Y3_FrameStrobe_O[13] ,
    \Tile_X9Y3_FrameStrobe_O[12] ,
    \Tile_X9Y3_FrameStrobe_O[11] ,
    \Tile_X9Y3_FrameStrobe_O[10] ,
    \Tile_X9Y3_FrameStrobe_O[9] ,
    \Tile_X9Y3_FrameStrobe_O[8] ,
    \Tile_X9Y3_FrameStrobe_O[7] ,
    \Tile_X9Y3_FrameStrobe_O[6] ,
    \Tile_X9Y3_FrameStrobe_O[5] ,
    \Tile_X9Y3_FrameStrobe_O[4] ,
    \Tile_X9Y3_FrameStrobe_O[3] ,
    \Tile_X9Y3_FrameStrobe_O[2] ,
    \Tile_X9Y3_FrameStrobe_O[1] ,
    \Tile_X9Y3_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X9Y3_N1BEG[3] ,
    \Tile_X9Y3_N1BEG[2] ,
    \Tile_X9Y3_N1BEG[1] ,
    \Tile_X9Y3_N1BEG[0] }),
    .N1END({\Tile_X9Y4_N1BEG[3] ,
    \Tile_X9Y4_N1BEG[2] ,
    \Tile_X9Y4_N1BEG[1] ,
    \Tile_X9Y4_N1BEG[0] }),
    .N2BEG({\Tile_X9Y3_N2BEG[7] ,
    \Tile_X9Y3_N2BEG[6] ,
    \Tile_X9Y3_N2BEG[5] ,
    \Tile_X9Y3_N2BEG[4] ,
    \Tile_X9Y3_N2BEG[3] ,
    \Tile_X9Y3_N2BEG[2] ,
    \Tile_X9Y3_N2BEG[1] ,
    \Tile_X9Y3_N2BEG[0] }),
    .N2BEGb({\Tile_X9Y3_N2BEGb[7] ,
    \Tile_X9Y3_N2BEGb[6] ,
    \Tile_X9Y3_N2BEGb[5] ,
    \Tile_X9Y3_N2BEGb[4] ,
    \Tile_X9Y3_N2BEGb[3] ,
    \Tile_X9Y3_N2BEGb[2] ,
    \Tile_X9Y3_N2BEGb[1] ,
    \Tile_X9Y3_N2BEGb[0] }),
    .N2END({\Tile_X9Y4_N2BEGb[7] ,
    \Tile_X9Y4_N2BEGb[6] ,
    \Tile_X9Y4_N2BEGb[5] ,
    \Tile_X9Y4_N2BEGb[4] ,
    \Tile_X9Y4_N2BEGb[3] ,
    \Tile_X9Y4_N2BEGb[2] ,
    \Tile_X9Y4_N2BEGb[1] ,
    \Tile_X9Y4_N2BEGb[0] }),
    .N2MID({\Tile_X9Y4_N2BEG[7] ,
    \Tile_X9Y4_N2BEG[6] ,
    \Tile_X9Y4_N2BEG[5] ,
    \Tile_X9Y4_N2BEG[4] ,
    \Tile_X9Y4_N2BEG[3] ,
    \Tile_X9Y4_N2BEG[2] ,
    \Tile_X9Y4_N2BEG[1] ,
    \Tile_X9Y4_N2BEG[0] }),
    .N4BEG({\Tile_X9Y3_N4BEG[15] ,
    \Tile_X9Y3_N4BEG[14] ,
    \Tile_X9Y3_N4BEG[13] ,
    \Tile_X9Y3_N4BEG[12] ,
    \Tile_X9Y3_N4BEG[11] ,
    \Tile_X9Y3_N4BEG[10] ,
    \Tile_X9Y3_N4BEG[9] ,
    \Tile_X9Y3_N4BEG[8] ,
    \Tile_X9Y3_N4BEG[7] ,
    \Tile_X9Y3_N4BEG[6] ,
    \Tile_X9Y3_N4BEG[5] ,
    \Tile_X9Y3_N4BEG[4] ,
    \Tile_X9Y3_N4BEG[3] ,
    \Tile_X9Y3_N4BEG[2] ,
    \Tile_X9Y3_N4BEG[1] ,
    \Tile_X9Y3_N4BEG[0] }),
    .N4END({\Tile_X9Y4_N4BEG[15] ,
    \Tile_X9Y4_N4BEG[14] ,
    \Tile_X9Y4_N4BEG[13] ,
    \Tile_X9Y4_N4BEG[12] ,
    \Tile_X9Y4_N4BEG[11] ,
    \Tile_X9Y4_N4BEG[10] ,
    \Tile_X9Y4_N4BEG[9] ,
    \Tile_X9Y4_N4BEG[8] ,
    \Tile_X9Y4_N4BEG[7] ,
    \Tile_X9Y4_N4BEG[6] ,
    \Tile_X9Y4_N4BEG[5] ,
    \Tile_X9Y4_N4BEG[4] ,
    \Tile_X9Y4_N4BEG[3] ,
    \Tile_X9Y4_N4BEG[2] ,
    \Tile_X9Y4_N4BEG[1] ,
    \Tile_X9Y4_N4BEG[0] }),
    .NN4BEG({\Tile_X9Y3_NN4BEG[15] ,
    \Tile_X9Y3_NN4BEG[14] ,
    \Tile_X9Y3_NN4BEG[13] ,
    \Tile_X9Y3_NN4BEG[12] ,
    \Tile_X9Y3_NN4BEG[11] ,
    \Tile_X9Y3_NN4BEG[10] ,
    \Tile_X9Y3_NN4BEG[9] ,
    \Tile_X9Y3_NN4BEG[8] ,
    \Tile_X9Y3_NN4BEG[7] ,
    \Tile_X9Y3_NN4BEG[6] ,
    \Tile_X9Y3_NN4BEG[5] ,
    \Tile_X9Y3_NN4BEG[4] ,
    \Tile_X9Y3_NN4BEG[3] ,
    \Tile_X9Y3_NN4BEG[2] ,
    \Tile_X9Y3_NN4BEG[1] ,
    \Tile_X9Y3_NN4BEG[0] }),
    .NN4END({\Tile_X9Y4_NN4BEG[15] ,
    \Tile_X9Y4_NN4BEG[14] ,
    \Tile_X9Y4_NN4BEG[13] ,
    \Tile_X9Y4_NN4BEG[12] ,
    \Tile_X9Y4_NN4BEG[11] ,
    \Tile_X9Y4_NN4BEG[10] ,
    \Tile_X9Y4_NN4BEG[9] ,
    \Tile_X9Y4_NN4BEG[8] ,
    \Tile_X9Y4_NN4BEG[7] ,
    \Tile_X9Y4_NN4BEG[6] ,
    \Tile_X9Y4_NN4BEG[5] ,
    \Tile_X9Y4_NN4BEG[4] ,
    \Tile_X9Y4_NN4BEG[3] ,
    \Tile_X9Y4_NN4BEG[2] ,
    \Tile_X9Y4_NN4BEG[1] ,
    \Tile_X9Y4_NN4BEG[0] }),
    .S1BEG({\Tile_X9Y3_S1BEG[3] ,
    \Tile_X9Y3_S1BEG[2] ,
    \Tile_X9Y3_S1BEG[1] ,
    \Tile_X9Y3_S1BEG[0] }),
    .S1END({\Tile_X9Y2_S1BEG[3] ,
    \Tile_X9Y2_S1BEG[2] ,
    \Tile_X9Y2_S1BEG[1] ,
    \Tile_X9Y2_S1BEG[0] }),
    .S2BEG({\Tile_X9Y3_S2BEG[7] ,
    \Tile_X9Y3_S2BEG[6] ,
    \Tile_X9Y3_S2BEG[5] ,
    \Tile_X9Y3_S2BEG[4] ,
    \Tile_X9Y3_S2BEG[3] ,
    \Tile_X9Y3_S2BEG[2] ,
    \Tile_X9Y3_S2BEG[1] ,
    \Tile_X9Y3_S2BEG[0] }),
    .S2BEGb({\Tile_X9Y3_S2BEGb[7] ,
    \Tile_X9Y3_S2BEGb[6] ,
    \Tile_X9Y3_S2BEGb[5] ,
    \Tile_X9Y3_S2BEGb[4] ,
    \Tile_X9Y3_S2BEGb[3] ,
    \Tile_X9Y3_S2BEGb[2] ,
    \Tile_X9Y3_S2BEGb[1] ,
    \Tile_X9Y3_S2BEGb[0] }),
    .S2END({\Tile_X9Y2_S2BEGb[7] ,
    \Tile_X9Y2_S2BEGb[6] ,
    \Tile_X9Y2_S2BEGb[5] ,
    \Tile_X9Y2_S2BEGb[4] ,
    \Tile_X9Y2_S2BEGb[3] ,
    \Tile_X9Y2_S2BEGb[2] ,
    \Tile_X9Y2_S2BEGb[1] ,
    \Tile_X9Y2_S2BEGb[0] }),
    .S2MID({\Tile_X9Y2_S2BEG[7] ,
    \Tile_X9Y2_S2BEG[6] ,
    \Tile_X9Y2_S2BEG[5] ,
    \Tile_X9Y2_S2BEG[4] ,
    \Tile_X9Y2_S2BEG[3] ,
    \Tile_X9Y2_S2BEG[2] ,
    \Tile_X9Y2_S2BEG[1] ,
    \Tile_X9Y2_S2BEG[0] }),
    .S4BEG({\Tile_X9Y3_S4BEG[15] ,
    \Tile_X9Y3_S4BEG[14] ,
    \Tile_X9Y3_S4BEG[13] ,
    \Tile_X9Y3_S4BEG[12] ,
    \Tile_X9Y3_S4BEG[11] ,
    \Tile_X9Y3_S4BEG[10] ,
    \Tile_X9Y3_S4BEG[9] ,
    \Tile_X9Y3_S4BEG[8] ,
    \Tile_X9Y3_S4BEG[7] ,
    \Tile_X9Y3_S4BEG[6] ,
    \Tile_X9Y3_S4BEG[5] ,
    \Tile_X9Y3_S4BEG[4] ,
    \Tile_X9Y3_S4BEG[3] ,
    \Tile_X9Y3_S4BEG[2] ,
    \Tile_X9Y3_S4BEG[1] ,
    \Tile_X9Y3_S4BEG[0] }),
    .S4END({\Tile_X9Y2_S4BEG[15] ,
    \Tile_X9Y2_S4BEG[14] ,
    \Tile_X9Y2_S4BEG[13] ,
    \Tile_X9Y2_S4BEG[12] ,
    \Tile_X9Y2_S4BEG[11] ,
    \Tile_X9Y2_S4BEG[10] ,
    \Tile_X9Y2_S4BEG[9] ,
    \Tile_X9Y2_S4BEG[8] ,
    \Tile_X9Y2_S4BEG[7] ,
    \Tile_X9Y2_S4BEG[6] ,
    \Tile_X9Y2_S4BEG[5] ,
    \Tile_X9Y2_S4BEG[4] ,
    \Tile_X9Y2_S4BEG[3] ,
    \Tile_X9Y2_S4BEG[2] ,
    \Tile_X9Y2_S4BEG[1] ,
    \Tile_X9Y2_S4BEG[0] }),
    .SS4BEG({\Tile_X9Y3_SS4BEG[15] ,
    \Tile_X9Y3_SS4BEG[14] ,
    \Tile_X9Y3_SS4BEG[13] ,
    \Tile_X9Y3_SS4BEG[12] ,
    \Tile_X9Y3_SS4BEG[11] ,
    \Tile_X9Y3_SS4BEG[10] ,
    \Tile_X9Y3_SS4BEG[9] ,
    \Tile_X9Y3_SS4BEG[8] ,
    \Tile_X9Y3_SS4BEG[7] ,
    \Tile_X9Y3_SS4BEG[6] ,
    \Tile_X9Y3_SS4BEG[5] ,
    \Tile_X9Y3_SS4BEG[4] ,
    \Tile_X9Y3_SS4BEG[3] ,
    \Tile_X9Y3_SS4BEG[2] ,
    \Tile_X9Y3_SS4BEG[1] ,
    \Tile_X9Y3_SS4BEG[0] }),
    .SS4END({\Tile_X9Y2_SS4BEG[15] ,
    \Tile_X9Y2_SS4BEG[14] ,
    \Tile_X9Y2_SS4BEG[13] ,
    \Tile_X9Y2_SS4BEG[12] ,
    \Tile_X9Y2_SS4BEG[11] ,
    \Tile_X9Y2_SS4BEG[10] ,
    \Tile_X9Y2_SS4BEG[9] ,
    \Tile_X9Y2_SS4BEG[8] ,
    \Tile_X9Y2_SS4BEG[7] ,
    \Tile_X9Y2_SS4BEG[6] ,
    \Tile_X9Y2_SS4BEG[5] ,
    \Tile_X9Y2_SS4BEG[4] ,
    \Tile_X9Y2_SS4BEG[3] ,
    \Tile_X9Y2_SS4BEG[2] ,
    \Tile_X9Y2_SS4BEG[1] ,
    \Tile_X9Y2_SS4BEG[0] }),
    .W1BEG({\Tile_X9Y3_W1BEG[3] ,
    \Tile_X9Y3_W1BEG[2] ,
    \Tile_X9Y3_W1BEG[1] ,
    \Tile_X9Y3_W1BEG[0] }),
    .W1END({\Tile_X10Y3_W1BEG[3] ,
    \Tile_X10Y3_W1BEG[2] ,
    \Tile_X10Y3_W1BEG[1] ,
    \Tile_X10Y3_W1BEG[0] }),
    .W2BEG({\Tile_X9Y3_W2BEG[7] ,
    \Tile_X9Y3_W2BEG[6] ,
    \Tile_X9Y3_W2BEG[5] ,
    \Tile_X9Y3_W2BEG[4] ,
    \Tile_X9Y3_W2BEG[3] ,
    \Tile_X9Y3_W2BEG[2] ,
    \Tile_X9Y3_W2BEG[1] ,
    \Tile_X9Y3_W2BEG[0] }),
    .W2BEGb({\Tile_X9Y3_W2BEGb[7] ,
    \Tile_X9Y3_W2BEGb[6] ,
    \Tile_X9Y3_W2BEGb[5] ,
    \Tile_X9Y3_W2BEGb[4] ,
    \Tile_X9Y3_W2BEGb[3] ,
    \Tile_X9Y3_W2BEGb[2] ,
    \Tile_X9Y3_W2BEGb[1] ,
    \Tile_X9Y3_W2BEGb[0] }),
    .W2END({\Tile_X10Y3_W2BEGb[7] ,
    \Tile_X10Y3_W2BEGb[6] ,
    \Tile_X10Y3_W2BEGb[5] ,
    \Tile_X10Y3_W2BEGb[4] ,
    \Tile_X10Y3_W2BEGb[3] ,
    \Tile_X10Y3_W2BEGb[2] ,
    \Tile_X10Y3_W2BEGb[1] ,
    \Tile_X10Y3_W2BEGb[0] }),
    .W2MID({\Tile_X10Y3_W2BEG[7] ,
    \Tile_X10Y3_W2BEG[6] ,
    \Tile_X10Y3_W2BEG[5] ,
    \Tile_X10Y3_W2BEG[4] ,
    \Tile_X10Y3_W2BEG[3] ,
    \Tile_X10Y3_W2BEG[2] ,
    \Tile_X10Y3_W2BEG[1] ,
    \Tile_X10Y3_W2BEG[0] }),
    .W6BEG({\Tile_X9Y3_W6BEG[11] ,
    \Tile_X9Y3_W6BEG[10] ,
    \Tile_X9Y3_W6BEG[9] ,
    \Tile_X9Y3_W6BEG[8] ,
    \Tile_X9Y3_W6BEG[7] ,
    \Tile_X9Y3_W6BEG[6] ,
    \Tile_X9Y3_W6BEG[5] ,
    \Tile_X9Y3_W6BEG[4] ,
    \Tile_X9Y3_W6BEG[3] ,
    \Tile_X9Y3_W6BEG[2] ,
    \Tile_X9Y3_W6BEG[1] ,
    \Tile_X9Y3_W6BEG[0] }),
    .W6END({\Tile_X10Y3_W6BEG[11] ,
    \Tile_X10Y3_W6BEG[10] ,
    \Tile_X10Y3_W6BEG[9] ,
    \Tile_X10Y3_W6BEG[8] ,
    \Tile_X10Y3_W6BEG[7] ,
    \Tile_X10Y3_W6BEG[6] ,
    \Tile_X10Y3_W6BEG[5] ,
    \Tile_X10Y3_W6BEG[4] ,
    \Tile_X10Y3_W6BEG[3] ,
    \Tile_X10Y3_W6BEG[2] ,
    \Tile_X10Y3_W6BEG[1] ,
    \Tile_X10Y3_W6BEG[0] }),
    .WW4BEG({\Tile_X9Y3_WW4BEG[15] ,
    \Tile_X9Y3_WW4BEG[14] ,
    \Tile_X9Y3_WW4BEG[13] ,
    \Tile_X9Y3_WW4BEG[12] ,
    \Tile_X9Y3_WW4BEG[11] ,
    \Tile_X9Y3_WW4BEG[10] ,
    \Tile_X9Y3_WW4BEG[9] ,
    \Tile_X9Y3_WW4BEG[8] ,
    \Tile_X9Y3_WW4BEG[7] ,
    \Tile_X9Y3_WW4BEG[6] ,
    \Tile_X9Y3_WW4BEG[5] ,
    \Tile_X9Y3_WW4BEG[4] ,
    \Tile_X9Y3_WW4BEG[3] ,
    \Tile_X9Y3_WW4BEG[2] ,
    \Tile_X9Y3_WW4BEG[1] ,
    \Tile_X9Y3_WW4BEG[0] }),
    .WW4END({\Tile_X10Y3_WW4BEG[15] ,
    \Tile_X10Y3_WW4BEG[14] ,
    \Tile_X10Y3_WW4BEG[13] ,
    \Tile_X10Y3_WW4BEG[12] ,
    \Tile_X10Y3_WW4BEG[11] ,
    \Tile_X10Y3_WW4BEG[10] ,
    \Tile_X10Y3_WW4BEG[9] ,
    \Tile_X10Y3_WW4BEG[8] ,
    \Tile_X10Y3_WW4BEG[7] ,
    \Tile_X10Y3_WW4BEG[6] ,
    \Tile_X10Y3_WW4BEG[5] ,
    \Tile_X10Y3_WW4BEG[4] ,
    \Tile_X10Y3_WW4BEG[3] ,
    \Tile_X10Y3_WW4BEG[2] ,
    \Tile_X10Y3_WW4BEG[1] ,
    \Tile_X10Y3_WW4BEG[0] }));
 LUT4AB Tile_X9Y4_LUT4AB (.Ci(Tile_X9Y5_Co),
    .Co(Tile_X9Y4_Co),
    .UserCLK(Tile_X9Y5_UserCLKo),
    .UserCLKo(Tile_X9Y4_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X9Y4_E1BEG[3] ,
    \Tile_X9Y4_E1BEG[2] ,
    \Tile_X9Y4_E1BEG[1] ,
    \Tile_X9Y4_E1BEG[0] }),
    .E1END({\Tile_X8Y4_E1BEG[3] ,
    \Tile_X8Y4_E1BEG[2] ,
    \Tile_X8Y4_E1BEG[1] ,
    \Tile_X8Y4_E1BEG[0] }),
    .E2BEG({\Tile_X9Y4_E2BEG[7] ,
    \Tile_X9Y4_E2BEG[6] ,
    \Tile_X9Y4_E2BEG[5] ,
    \Tile_X9Y4_E2BEG[4] ,
    \Tile_X9Y4_E2BEG[3] ,
    \Tile_X9Y4_E2BEG[2] ,
    \Tile_X9Y4_E2BEG[1] ,
    \Tile_X9Y4_E2BEG[0] }),
    .E2BEGb({\Tile_X9Y4_E2BEGb[7] ,
    \Tile_X9Y4_E2BEGb[6] ,
    \Tile_X9Y4_E2BEGb[5] ,
    \Tile_X9Y4_E2BEGb[4] ,
    \Tile_X9Y4_E2BEGb[3] ,
    \Tile_X9Y4_E2BEGb[2] ,
    \Tile_X9Y4_E2BEGb[1] ,
    \Tile_X9Y4_E2BEGb[0] }),
    .E2END({\Tile_X8Y4_E2BEGb[7] ,
    \Tile_X8Y4_E2BEGb[6] ,
    \Tile_X8Y4_E2BEGb[5] ,
    \Tile_X8Y4_E2BEGb[4] ,
    \Tile_X8Y4_E2BEGb[3] ,
    \Tile_X8Y4_E2BEGb[2] ,
    \Tile_X8Y4_E2BEGb[1] ,
    \Tile_X8Y4_E2BEGb[0] }),
    .E2MID({\Tile_X8Y4_E2BEG[7] ,
    \Tile_X8Y4_E2BEG[6] ,
    \Tile_X8Y4_E2BEG[5] ,
    \Tile_X8Y4_E2BEG[4] ,
    \Tile_X8Y4_E2BEG[3] ,
    \Tile_X8Y4_E2BEG[2] ,
    \Tile_X8Y4_E2BEG[1] ,
    \Tile_X8Y4_E2BEG[0] }),
    .E6BEG({\Tile_X9Y4_E6BEG[11] ,
    \Tile_X9Y4_E6BEG[10] ,
    \Tile_X9Y4_E6BEG[9] ,
    \Tile_X9Y4_E6BEG[8] ,
    \Tile_X9Y4_E6BEG[7] ,
    \Tile_X9Y4_E6BEG[6] ,
    \Tile_X9Y4_E6BEG[5] ,
    \Tile_X9Y4_E6BEG[4] ,
    \Tile_X9Y4_E6BEG[3] ,
    \Tile_X9Y4_E6BEG[2] ,
    \Tile_X9Y4_E6BEG[1] ,
    \Tile_X9Y4_E6BEG[0] }),
    .E6END({\Tile_X8Y4_E6BEG[11] ,
    \Tile_X8Y4_E6BEG[10] ,
    \Tile_X8Y4_E6BEG[9] ,
    \Tile_X8Y4_E6BEG[8] ,
    \Tile_X8Y4_E6BEG[7] ,
    \Tile_X8Y4_E6BEG[6] ,
    \Tile_X8Y4_E6BEG[5] ,
    \Tile_X8Y4_E6BEG[4] ,
    \Tile_X8Y4_E6BEG[3] ,
    \Tile_X8Y4_E6BEG[2] ,
    \Tile_X8Y4_E6BEG[1] ,
    \Tile_X8Y4_E6BEG[0] }),
    .EE4BEG({\Tile_X9Y4_EE4BEG[15] ,
    \Tile_X9Y4_EE4BEG[14] ,
    \Tile_X9Y4_EE4BEG[13] ,
    \Tile_X9Y4_EE4BEG[12] ,
    \Tile_X9Y4_EE4BEG[11] ,
    \Tile_X9Y4_EE4BEG[10] ,
    \Tile_X9Y4_EE4BEG[9] ,
    \Tile_X9Y4_EE4BEG[8] ,
    \Tile_X9Y4_EE4BEG[7] ,
    \Tile_X9Y4_EE4BEG[6] ,
    \Tile_X9Y4_EE4BEG[5] ,
    \Tile_X9Y4_EE4BEG[4] ,
    \Tile_X9Y4_EE4BEG[3] ,
    \Tile_X9Y4_EE4BEG[2] ,
    \Tile_X9Y4_EE4BEG[1] ,
    \Tile_X9Y4_EE4BEG[0] }),
    .EE4END({\Tile_X8Y4_EE4BEG[15] ,
    \Tile_X8Y4_EE4BEG[14] ,
    \Tile_X8Y4_EE4BEG[13] ,
    \Tile_X8Y4_EE4BEG[12] ,
    \Tile_X8Y4_EE4BEG[11] ,
    \Tile_X8Y4_EE4BEG[10] ,
    \Tile_X8Y4_EE4BEG[9] ,
    \Tile_X8Y4_EE4BEG[8] ,
    \Tile_X8Y4_EE4BEG[7] ,
    \Tile_X8Y4_EE4BEG[6] ,
    \Tile_X8Y4_EE4BEG[5] ,
    \Tile_X8Y4_EE4BEG[4] ,
    \Tile_X8Y4_EE4BEG[3] ,
    \Tile_X8Y4_EE4BEG[2] ,
    \Tile_X8Y4_EE4BEG[1] ,
    \Tile_X8Y4_EE4BEG[0] }),
    .FrameData({\Tile_X8Y4_FrameData_O[31] ,
    \Tile_X8Y4_FrameData_O[30] ,
    \Tile_X8Y4_FrameData_O[29] ,
    \Tile_X8Y4_FrameData_O[28] ,
    \Tile_X8Y4_FrameData_O[27] ,
    \Tile_X8Y4_FrameData_O[26] ,
    \Tile_X8Y4_FrameData_O[25] ,
    \Tile_X8Y4_FrameData_O[24] ,
    \Tile_X8Y4_FrameData_O[23] ,
    \Tile_X8Y4_FrameData_O[22] ,
    \Tile_X8Y4_FrameData_O[21] ,
    \Tile_X8Y4_FrameData_O[20] ,
    \Tile_X8Y4_FrameData_O[19] ,
    \Tile_X8Y4_FrameData_O[18] ,
    \Tile_X8Y4_FrameData_O[17] ,
    \Tile_X8Y4_FrameData_O[16] ,
    \Tile_X8Y4_FrameData_O[15] ,
    \Tile_X8Y4_FrameData_O[14] ,
    \Tile_X8Y4_FrameData_O[13] ,
    \Tile_X8Y4_FrameData_O[12] ,
    \Tile_X8Y4_FrameData_O[11] ,
    \Tile_X8Y4_FrameData_O[10] ,
    \Tile_X8Y4_FrameData_O[9] ,
    \Tile_X8Y4_FrameData_O[8] ,
    \Tile_X8Y4_FrameData_O[7] ,
    \Tile_X8Y4_FrameData_O[6] ,
    \Tile_X8Y4_FrameData_O[5] ,
    \Tile_X8Y4_FrameData_O[4] ,
    \Tile_X8Y4_FrameData_O[3] ,
    \Tile_X8Y4_FrameData_O[2] ,
    \Tile_X8Y4_FrameData_O[1] ,
    \Tile_X8Y4_FrameData_O[0] }),
    .FrameData_O({\Tile_X9Y4_FrameData_O[31] ,
    \Tile_X9Y4_FrameData_O[30] ,
    \Tile_X9Y4_FrameData_O[29] ,
    \Tile_X9Y4_FrameData_O[28] ,
    \Tile_X9Y4_FrameData_O[27] ,
    \Tile_X9Y4_FrameData_O[26] ,
    \Tile_X9Y4_FrameData_O[25] ,
    \Tile_X9Y4_FrameData_O[24] ,
    \Tile_X9Y4_FrameData_O[23] ,
    \Tile_X9Y4_FrameData_O[22] ,
    \Tile_X9Y4_FrameData_O[21] ,
    \Tile_X9Y4_FrameData_O[20] ,
    \Tile_X9Y4_FrameData_O[19] ,
    \Tile_X9Y4_FrameData_O[18] ,
    \Tile_X9Y4_FrameData_O[17] ,
    \Tile_X9Y4_FrameData_O[16] ,
    \Tile_X9Y4_FrameData_O[15] ,
    \Tile_X9Y4_FrameData_O[14] ,
    \Tile_X9Y4_FrameData_O[13] ,
    \Tile_X9Y4_FrameData_O[12] ,
    \Tile_X9Y4_FrameData_O[11] ,
    \Tile_X9Y4_FrameData_O[10] ,
    \Tile_X9Y4_FrameData_O[9] ,
    \Tile_X9Y4_FrameData_O[8] ,
    \Tile_X9Y4_FrameData_O[7] ,
    \Tile_X9Y4_FrameData_O[6] ,
    \Tile_X9Y4_FrameData_O[5] ,
    \Tile_X9Y4_FrameData_O[4] ,
    \Tile_X9Y4_FrameData_O[3] ,
    \Tile_X9Y4_FrameData_O[2] ,
    \Tile_X9Y4_FrameData_O[1] ,
    \Tile_X9Y4_FrameData_O[0] }),
    .FrameStrobe({\Tile_X9Y5_FrameStrobe_O[19] ,
    \Tile_X9Y5_FrameStrobe_O[18] ,
    \Tile_X9Y5_FrameStrobe_O[17] ,
    \Tile_X9Y5_FrameStrobe_O[16] ,
    \Tile_X9Y5_FrameStrobe_O[15] ,
    \Tile_X9Y5_FrameStrobe_O[14] ,
    \Tile_X9Y5_FrameStrobe_O[13] ,
    \Tile_X9Y5_FrameStrobe_O[12] ,
    \Tile_X9Y5_FrameStrobe_O[11] ,
    \Tile_X9Y5_FrameStrobe_O[10] ,
    \Tile_X9Y5_FrameStrobe_O[9] ,
    \Tile_X9Y5_FrameStrobe_O[8] ,
    \Tile_X9Y5_FrameStrobe_O[7] ,
    \Tile_X9Y5_FrameStrobe_O[6] ,
    \Tile_X9Y5_FrameStrobe_O[5] ,
    \Tile_X9Y5_FrameStrobe_O[4] ,
    \Tile_X9Y5_FrameStrobe_O[3] ,
    \Tile_X9Y5_FrameStrobe_O[2] ,
    \Tile_X9Y5_FrameStrobe_O[1] ,
    \Tile_X9Y5_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X9Y4_FrameStrobe_O[19] ,
    \Tile_X9Y4_FrameStrobe_O[18] ,
    \Tile_X9Y4_FrameStrobe_O[17] ,
    \Tile_X9Y4_FrameStrobe_O[16] ,
    \Tile_X9Y4_FrameStrobe_O[15] ,
    \Tile_X9Y4_FrameStrobe_O[14] ,
    \Tile_X9Y4_FrameStrobe_O[13] ,
    \Tile_X9Y4_FrameStrobe_O[12] ,
    \Tile_X9Y4_FrameStrobe_O[11] ,
    \Tile_X9Y4_FrameStrobe_O[10] ,
    \Tile_X9Y4_FrameStrobe_O[9] ,
    \Tile_X9Y4_FrameStrobe_O[8] ,
    \Tile_X9Y4_FrameStrobe_O[7] ,
    \Tile_X9Y4_FrameStrobe_O[6] ,
    \Tile_X9Y4_FrameStrobe_O[5] ,
    \Tile_X9Y4_FrameStrobe_O[4] ,
    \Tile_X9Y4_FrameStrobe_O[3] ,
    \Tile_X9Y4_FrameStrobe_O[2] ,
    \Tile_X9Y4_FrameStrobe_O[1] ,
    \Tile_X9Y4_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X9Y4_N1BEG[3] ,
    \Tile_X9Y4_N1BEG[2] ,
    \Tile_X9Y4_N1BEG[1] ,
    \Tile_X9Y4_N1BEG[0] }),
    .N1END({\Tile_X9Y5_N1BEG[3] ,
    \Tile_X9Y5_N1BEG[2] ,
    \Tile_X9Y5_N1BEG[1] ,
    \Tile_X9Y5_N1BEG[0] }),
    .N2BEG({\Tile_X9Y4_N2BEG[7] ,
    \Tile_X9Y4_N2BEG[6] ,
    \Tile_X9Y4_N2BEG[5] ,
    \Tile_X9Y4_N2BEG[4] ,
    \Tile_X9Y4_N2BEG[3] ,
    \Tile_X9Y4_N2BEG[2] ,
    \Tile_X9Y4_N2BEG[1] ,
    \Tile_X9Y4_N2BEG[0] }),
    .N2BEGb({\Tile_X9Y4_N2BEGb[7] ,
    \Tile_X9Y4_N2BEGb[6] ,
    \Tile_X9Y4_N2BEGb[5] ,
    \Tile_X9Y4_N2BEGb[4] ,
    \Tile_X9Y4_N2BEGb[3] ,
    \Tile_X9Y4_N2BEGb[2] ,
    \Tile_X9Y4_N2BEGb[1] ,
    \Tile_X9Y4_N2BEGb[0] }),
    .N2END({\Tile_X9Y5_N2BEGb[7] ,
    \Tile_X9Y5_N2BEGb[6] ,
    \Tile_X9Y5_N2BEGb[5] ,
    \Tile_X9Y5_N2BEGb[4] ,
    \Tile_X9Y5_N2BEGb[3] ,
    \Tile_X9Y5_N2BEGb[2] ,
    \Tile_X9Y5_N2BEGb[1] ,
    \Tile_X9Y5_N2BEGb[0] }),
    .N2MID({\Tile_X9Y5_N2BEG[7] ,
    \Tile_X9Y5_N2BEG[6] ,
    \Tile_X9Y5_N2BEG[5] ,
    \Tile_X9Y5_N2BEG[4] ,
    \Tile_X9Y5_N2BEG[3] ,
    \Tile_X9Y5_N2BEG[2] ,
    \Tile_X9Y5_N2BEG[1] ,
    \Tile_X9Y5_N2BEG[0] }),
    .N4BEG({\Tile_X9Y4_N4BEG[15] ,
    \Tile_X9Y4_N4BEG[14] ,
    \Tile_X9Y4_N4BEG[13] ,
    \Tile_X9Y4_N4BEG[12] ,
    \Tile_X9Y4_N4BEG[11] ,
    \Tile_X9Y4_N4BEG[10] ,
    \Tile_X9Y4_N4BEG[9] ,
    \Tile_X9Y4_N4BEG[8] ,
    \Tile_X9Y4_N4BEG[7] ,
    \Tile_X9Y4_N4BEG[6] ,
    \Tile_X9Y4_N4BEG[5] ,
    \Tile_X9Y4_N4BEG[4] ,
    \Tile_X9Y4_N4BEG[3] ,
    \Tile_X9Y4_N4BEG[2] ,
    \Tile_X9Y4_N4BEG[1] ,
    \Tile_X9Y4_N4BEG[0] }),
    .N4END({\Tile_X9Y5_N4BEG[15] ,
    \Tile_X9Y5_N4BEG[14] ,
    \Tile_X9Y5_N4BEG[13] ,
    \Tile_X9Y5_N4BEG[12] ,
    \Tile_X9Y5_N4BEG[11] ,
    \Tile_X9Y5_N4BEG[10] ,
    \Tile_X9Y5_N4BEG[9] ,
    \Tile_X9Y5_N4BEG[8] ,
    \Tile_X9Y5_N4BEG[7] ,
    \Tile_X9Y5_N4BEG[6] ,
    \Tile_X9Y5_N4BEG[5] ,
    \Tile_X9Y5_N4BEG[4] ,
    \Tile_X9Y5_N4BEG[3] ,
    \Tile_X9Y5_N4BEG[2] ,
    \Tile_X9Y5_N4BEG[1] ,
    \Tile_X9Y5_N4BEG[0] }),
    .NN4BEG({\Tile_X9Y4_NN4BEG[15] ,
    \Tile_X9Y4_NN4BEG[14] ,
    \Tile_X9Y4_NN4BEG[13] ,
    \Tile_X9Y4_NN4BEG[12] ,
    \Tile_X9Y4_NN4BEG[11] ,
    \Tile_X9Y4_NN4BEG[10] ,
    \Tile_X9Y4_NN4BEG[9] ,
    \Tile_X9Y4_NN4BEG[8] ,
    \Tile_X9Y4_NN4BEG[7] ,
    \Tile_X9Y4_NN4BEG[6] ,
    \Tile_X9Y4_NN4BEG[5] ,
    \Tile_X9Y4_NN4BEG[4] ,
    \Tile_X9Y4_NN4BEG[3] ,
    \Tile_X9Y4_NN4BEG[2] ,
    \Tile_X9Y4_NN4BEG[1] ,
    \Tile_X9Y4_NN4BEG[0] }),
    .NN4END({\Tile_X9Y5_NN4BEG[15] ,
    \Tile_X9Y5_NN4BEG[14] ,
    \Tile_X9Y5_NN4BEG[13] ,
    \Tile_X9Y5_NN4BEG[12] ,
    \Tile_X9Y5_NN4BEG[11] ,
    \Tile_X9Y5_NN4BEG[10] ,
    \Tile_X9Y5_NN4BEG[9] ,
    \Tile_X9Y5_NN4BEG[8] ,
    \Tile_X9Y5_NN4BEG[7] ,
    \Tile_X9Y5_NN4BEG[6] ,
    \Tile_X9Y5_NN4BEG[5] ,
    \Tile_X9Y5_NN4BEG[4] ,
    \Tile_X9Y5_NN4BEG[3] ,
    \Tile_X9Y5_NN4BEG[2] ,
    \Tile_X9Y5_NN4BEG[1] ,
    \Tile_X9Y5_NN4BEG[0] }),
    .S1BEG({\Tile_X9Y4_S1BEG[3] ,
    \Tile_X9Y4_S1BEG[2] ,
    \Tile_X9Y4_S1BEG[1] ,
    \Tile_X9Y4_S1BEG[0] }),
    .S1END({\Tile_X9Y3_S1BEG[3] ,
    \Tile_X9Y3_S1BEG[2] ,
    \Tile_X9Y3_S1BEG[1] ,
    \Tile_X9Y3_S1BEG[0] }),
    .S2BEG({\Tile_X9Y4_S2BEG[7] ,
    \Tile_X9Y4_S2BEG[6] ,
    \Tile_X9Y4_S2BEG[5] ,
    \Tile_X9Y4_S2BEG[4] ,
    \Tile_X9Y4_S2BEG[3] ,
    \Tile_X9Y4_S2BEG[2] ,
    \Tile_X9Y4_S2BEG[1] ,
    \Tile_X9Y4_S2BEG[0] }),
    .S2BEGb({\Tile_X9Y4_S2BEGb[7] ,
    \Tile_X9Y4_S2BEGb[6] ,
    \Tile_X9Y4_S2BEGb[5] ,
    \Tile_X9Y4_S2BEGb[4] ,
    \Tile_X9Y4_S2BEGb[3] ,
    \Tile_X9Y4_S2BEGb[2] ,
    \Tile_X9Y4_S2BEGb[1] ,
    \Tile_X9Y4_S2BEGb[0] }),
    .S2END({\Tile_X9Y3_S2BEGb[7] ,
    \Tile_X9Y3_S2BEGb[6] ,
    \Tile_X9Y3_S2BEGb[5] ,
    \Tile_X9Y3_S2BEGb[4] ,
    \Tile_X9Y3_S2BEGb[3] ,
    \Tile_X9Y3_S2BEGb[2] ,
    \Tile_X9Y3_S2BEGb[1] ,
    \Tile_X9Y3_S2BEGb[0] }),
    .S2MID({\Tile_X9Y3_S2BEG[7] ,
    \Tile_X9Y3_S2BEG[6] ,
    \Tile_X9Y3_S2BEG[5] ,
    \Tile_X9Y3_S2BEG[4] ,
    \Tile_X9Y3_S2BEG[3] ,
    \Tile_X9Y3_S2BEG[2] ,
    \Tile_X9Y3_S2BEG[1] ,
    \Tile_X9Y3_S2BEG[0] }),
    .S4BEG({\Tile_X9Y4_S4BEG[15] ,
    \Tile_X9Y4_S4BEG[14] ,
    \Tile_X9Y4_S4BEG[13] ,
    \Tile_X9Y4_S4BEG[12] ,
    \Tile_X9Y4_S4BEG[11] ,
    \Tile_X9Y4_S4BEG[10] ,
    \Tile_X9Y4_S4BEG[9] ,
    \Tile_X9Y4_S4BEG[8] ,
    \Tile_X9Y4_S4BEG[7] ,
    \Tile_X9Y4_S4BEG[6] ,
    \Tile_X9Y4_S4BEG[5] ,
    \Tile_X9Y4_S4BEG[4] ,
    \Tile_X9Y4_S4BEG[3] ,
    \Tile_X9Y4_S4BEG[2] ,
    \Tile_X9Y4_S4BEG[1] ,
    \Tile_X9Y4_S4BEG[0] }),
    .S4END({\Tile_X9Y3_S4BEG[15] ,
    \Tile_X9Y3_S4BEG[14] ,
    \Tile_X9Y3_S4BEG[13] ,
    \Tile_X9Y3_S4BEG[12] ,
    \Tile_X9Y3_S4BEG[11] ,
    \Tile_X9Y3_S4BEG[10] ,
    \Tile_X9Y3_S4BEG[9] ,
    \Tile_X9Y3_S4BEG[8] ,
    \Tile_X9Y3_S4BEG[7] ,
    \Tile_X9Y3_S4BEG[6] ,
    \Tile_X9Y3_S4BEG[5] ,
    \Tile_X9Y3_S4BEG[4] ,
    \Tile_X9Y3_S4BEG[3] ,
    \Tile_X9Y3_S4BEG[2] ,
    \Tile_X9Y3_S4BEG[1] ,
    \Tile_X9Y3_S4BEG[0] }),
    .SS4BEG({\Tile_X9Y4_SS4BEG[15] ,
    \Tile_X9Y4_SS4BEG[14] ,
    \Tile_X9Y4_SS4BEG[13] ,
    \Tile_X9Y4_SS4BEG[12] ,
    \Tile_X9Y4_SS4BEG[11] ,
    \Tile_X9Y4_SS4BEG[10] ,
    \Tile_X9Y4_SS4BEG[9] ,
    \Tile_X9Y4_SS4BEG[8] ,
    \Tile_X9Y4_SS4BEG[7] ,
    \Tile_X9Y4_SS4BEG[6] ,
    \Tile_X9Y4_SS4BEG[5] ,
    \Tile_X9Y4_SS4BEG[4] ,
    \Tile_X9Y4_SS4BEG[3] ,
    \Tile_X9Y4_SS4BEG[2] ,
    \Tile_X9Y4_SS4BEG[1] ,
    \Tile_X9Y4_SS4BEG[0] }),
    .SS4END({\Tile_X9Y3_SS4BEG[15] ,
    \Tile_X9Y3_SS4BEG[14] ,
    \Tile_X9Y3_SS4BEG[13] ,
    \Tile_X9Y3_SS4BEG[12] ,
    \Tile_X9Y3_SS4BEG[11] ,
    \Tile_X9Y3_SS4BEG[10] ,
    \Tile_X9Y3_SS4BEG[9] ,
    \Tile_X9Y3_SS4BEG[8] ,
    \Tile_X9Y3_SS4BEG[7] ,
    \Tile_X9Y3_SS4BEG[6] ,
    \Tile_X9Y3_SS4BEG[5] ,
    \Tile_X9Y3_SS4BEG[4] ,
    \Tile_X9Y3_SS4BEG[3] ,
    \Tile_X9Y3_SS4BEG[2] ,
    \Tile_X9Y3_SS4BEG[1] ,
    \Tile_X9Y3_SS4BEG[0] }),
    .W1BEG({\Tile_X9Y4_W1BEG[3] ,
    \Tile_X9Y4_W1BEG[2] ,
    \Tile_X9Y4_W1BEG[1] ,
    \Tile_X9Y4_W1BEG[0] }),
    .W1END({\Tile_X10Y4_W1BEG[3] ,
    \Tile_X10Y4_W1BEG[2] ,
    \Tile_X10Y4_W1BEG[1] ,
    \Tile_X10Y4_W1BEG[0] }),
    .W2BEG({\Tile_X9Y4_W2BEG[7] ,
    \Tile_X9Y4_W2BEG[6] ,
    \Tile_X9Y4_W2BEG[5] ,
    \Tile_X9Y4_W2BEG[4] ,
    \Tile_X9Y4_W2BEG[3] ,
    \Tile_X9Y4_W2BEG[2] ,
    \Tile_X9Y4_W2BEG[1] ,
    \Tile_X9Y4_W2BEG[0] }),
    .W2BEGb({\Tile_X9Y4_W2BEGb[7] ,
    \Tile_X9Y4_W2BEGb[6] ,
    \Tile_X9Y4_W2BEGb[5] ,
    \Tile_X9Y4_W2BEGb[4] ,
    \Tile_X9Y4_W2BEGb[3] ,
    \Tile_X9Y4_W2BEGb[2] ,
    \Tile_X9Y4_W2BEGb[1] ,
    \Tile_X9Y4_W2BEGb[0] }),
    .W2END({\Tile_X10Y4_W2BEGb[7] ,
    \Tile_X10Y4_W2BEGb[6] ,
    \Tile_X10Y4_W2BEGb[5] ,
    \Tile_X10Y4_W2BEGb[4] ,
    \Tile_X10Y4_W2BEGb[3] ,
    \Tile_X10Y4_W2BEGb[2] ,
    \Tile_X10Y4_W2BEGb[1] ,
    \Tile_X10Y4_W2BEGb[0] }),
    .W2MID({\Tile_X10Y4_W2BEG[7] ,
    \Tile_X10Y4_W2BEG[6] ,
    \Tile_X10Y4_W2BEG[5] ,
    \Tile_X10Y4_W2BEG[4] ,
    \Tile_X10Y4_W2BEG[3] ,
    \Tile_X10Y4_W2BEG[2] ,
    \Tile_X10Y4_W2BEG[1] ,
    \Tile_X10Y4_W2BEG[0] }),
    .W6BEG({\Tile_X9Y4_W6BEG[11] ,
    \Tile_X9Y4_W6BEG[10] ,
    \Tile_X9Y4_W6BEG[9] ,
    \Tile_X9Y4_W6BEG[8] ,
    \Tile_X9Y4_W6BEG[7] ,
    \Tile_X9Y4_W6BEG[6] ,
    \Tile_X9Y4_W6BEG[5] ,
    \Tile_X9Y4_W6BEG[4] ,
    \Tile_X9Y4_W6BEG[3] ,
    \Tile_X9Y4_W6BEG[2] ,
    \Tile_X9Y4_W6BEG[1] ,
    \Tile_X9Y4_W6BEG[0] }),
    .W6END({\Tile_X10Y4_W6BEG[11] ,
    \Tile_X10Y4_W6BEG[10] ,
    \Tile_X10Y4_W6BEG[9] ,
    \Tile_X10Y4_W6BEG[8] ,
    \Tile_X10Y4_W6BEG[7] ,
    \Tile_X10Y4_W6BEG[6] ,
    \Tile_X10Y4_W6BEG[5] ,
    \Tile_X10Y4_W6BEG[4] ,
    \Tile_X10Y4_W6BEG[3] ,
    \Tile_X10Y4_W6BEG[2] ,
    \Tile_X10Y4_W6BEG[1] ,
    \Tile_X10Y4_W6BEG[0] }),
    .WW4BEG({\Tile_X9Y4_WW4BEG[15] ,
    \Tile_X9Y4_WW4BEG[14] ,
    \Tile_X9Y4_WW4BEG[13] ,
    \Tile_X9Y4_WW4BEG[12] ,
    \Tile_X9Y4_WW4BEG[11] ,
    \Tile_X9Y4_WW4BEG[10] ,
    \Tile_X9Y4_WW4BEG[9] ,
    \Tile_X9Y4_WW4BEG[8] ,
    \Tile_X9Y4_WW4BEG[7] ,
    \Tile_X9Y4_WW4BEG[6] ,
    \Tile_X9Y4_WW4BEG[5] ,
    \Tile_X9Y4_WW4BEG[4] ,
    \Tile_X9Y4_WW4BEG[3] ,
    \Tile_X9Y4_WW4BEG[2] ,
    \Tile_X9Y4_WW4BEG[1] ,
    \Tile_X9Y4_WW4BEG[0] }),
    .WW4END({\Tile_X10Y4_WW4BEG[15] ,
    \Tile_X10Y4_WW4BEG[14] ,
    \Tile_X10Y4_WW4BEG[13] ,
    \Tile_X10Y4_WW4BEG[12] ,
    \Tile_X10Y4_WW4BEG[11] ,
    \Tile_X10Y4_WW4BEG[10] ,
    \Tile_X10Y4_WW4BEG[9] ,
    \Tile_X10Y4_WW4BEG[8] ,
    \Tile_X10Y4_WW4BEG[7] ,
    \Tile_X10Y4_WW4BEG[6] ,
    \Tile_X10Y4_WW4BEG[5] ,
    \Tile_X10Y4_WW4BEG[4] ,
    \Tile_X10Y4_WW4BEG[3] ,
    \Tile_X10Y4_WW4BEG[2] ,
    \Tile_X10Y4_WW4BEG[1] ,
    \Tile_X10Y4_WW4BEG[0] }));
 LUT4AB Tile_X9Y5_LUT4AB (.Ci(Tile_X9Y6_Co),
    .Co(Tile_X9Y5_Co),
    .UserCLK(Tile_X9Y6_UserCLKo),
    .UserCLKo(Tile_X9Y5_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X9Y5_E1BEG[3] ,
    \Tile_X9Y5_E1BEG[2] ,
    \Tile_X9Y5_E1BEG[1] ,
    \Tile_X9Y5_E1BEG[0] }),
    .E1END({\Tile_X8Y5_E1BEG[3] ,
    \Tile_X8Y5_E1BEG[2] ,
    \Tile_X8Y5_E1BEG[1] ,
    \Tile_X8Y5_E1BEG[0] }),
    .E2BEG({\Tile_X9Y5_E2BEG[7] ,
    \Tile_X9Y5_E2BEG[6] ,
    \Tile_X9Y5_E2BEG[5] ,
    \Tile_X9Y5_E2BEG[4] ,
    \Tile_X9Y5_E2BEG[3] ,
    \Tile_X9Y5_E2BEG[2] ,
    \Tile_X9Y5_E2BEG[1] ,
    \Tile_X9Y5_E2BEG[0] }),
    .E2BEGb({\Tile_X9Y5_E2BEGb[7] ,
    \Tile_X9Y5_E2BEGb[6] ,
    \Tile_X9Y5_E2BEGb[5] ,
    \Tile_X9Y5_E2BEGb[4] ,
    \Tile_X9Y5_E2BEGb[3] ,
    \Tile_X9Y5_E2BEGb[2] ,
    \Tile_X9Y5_E2BEGb[1] ,
    \Tile_X9Y5_E2BEGb[0] }),
    .E2END({\Tile_X8Y5_E2BEGb[7] ,
    \Tile_X8Y5_E2BEGb[6] ,
    \Tile_X8Y5_E2BEGb[5] ,
    \Tile_X8Y5_E2BEGb[4] ,
    \Tile_X8Y5_E2BEGb[3] ,
    \Tile_X8Y5_E2BEGb[2] ,
    \Tile_X8Y5_E2BEGb[1] ,
    \Tile_X8Y5_E2BEGb[0] }),
    .E2MID({\Tile_X8Y5_E2BEG[7] ,
    \Tile_X8Y5_E2BEG[6] ,
    \Tile_X8Y5_E2BEG[5] ,
    \Tile_X8Y5_E2BEG[4] ,
    \Tile_X8Y5_E2BEG[3] ,
    \Tile_X8Y5_E2BEG[2] ,
    \Tile_X8Y5_E2BEG[1] ,
    \Tile_X8Y5_E2BEG[0] }),
    .E6BEG({\Tile_X9Y5_E6BEG[11] ,
    \Tile_X9Y5_E6BEG[10] ,
    \Tile_X9Y5_E6BEG[9] ,
    \Tile_X9Y5_E6BEG[8] ,
    \Tile_X9Y5_E6BEG[7] ,
    \Tile_X9Y5_E6BEG[6] ,
    \Tile_X9Y5_E6BEG[5] ,
    \Tile_X9Y5_E6BEG[4] ,
    \Tile_X9Y5_E6BEG[3] ,
    \Tile_X9Y5_E6BEG[2] ,
    \Tile_X9Y5_E6BEG[1] ,
    \Tile_X9Y5_E6BEG[0] }),
    .E6END({\Tile_X8Y5_E6BEG[11] ,
    \Tile_X8Y5_E6BEG[10] ,
    \Tile_X8Y5_E6BEG[9] ,
    \Tile_X8Y5_E6BEG[8] ,
    \Tile_X8Y5_E6BEG[7] ,
    \Tile_X8Y5_E6BEG[6] ,
    \Tile_X8Y5_E6BEG[5] ,
    \Tile_X8Y5_E6BEG[4] ,
    \Tile_X8Y5_E6BEG[3] ,
    \Tile_X8Y5_E6BEG[2] ,
    \Tile_X8Y5_E6BEG[1] ,
    \Tile_X8Y5_E6BEG[0] }),
    .EE4BEG({\Tile_X9Y5_EE4BEG[15] ,
    \Tile_X9Y5_EE4BEG[14] ,
    \Tile_X9Y5_EE4BEG[13] ,
    \Tile_X9Y5_EE4BEG[12] ,
    \Tile_X9Y5_EE4BEG[11] ,
    \Tile_X9Y5_EE4BEG[10] ,
    \Tile_X9Y5_EE4BEG[9] ,
    \Tile_X9Y5_EE4BEG[8] ,
    \Tile_X9Y5_EE4BEG[7] ,
    \Tile_X9Y5_EE4BEG[6] ,
    \Tile_X9Y5_EE4BEG[5] ,
    \Tile_X9Y5_EE4BEG[4] ,
    \Tile_X9Y5_EE4BEG[3] ,
    \Tile_X9Y5_EE4BEG[2] ,
    \Tile_X9Y5_EE4BEG[1] ,
    \Tile_X9Y5_EE4BEG[0] }),
    .EE4END({\Tile_X8Y5_EE4BEG[15] ,
    \Tile_X8Y5_EE4BEG[14] ,
    \Tile_X8Y5_EE4BEG[13] ,
    \Tile_X8Y5_EE4BEG[12] ,
    \Tile_X8Y5_EE4BEG[11] ,
    \Tile_X8Y5_EE4BEG[10] ,
    \Tile_X8Y5_EE4BEG[9] ,
    \Tile_X8Y5_EE4BEG[8] ,
    \Tile_X8Y5_EE4BEG[7] ,
    \Tile_X8Y5_EE4BEG[6] ,
    \Tile_X8Y5_EE4BEG[5] ,
    \Tile_X8Y5_EE4BEG[4] ,
    \Tile_X8Y5_EE4BEG[3] ,
    \Tile_X8Y5_EE4BEG[2] ,
    \Tile_X8Y5_EE4BEG[1] ,
    \Tile_X8Y5_EE4BEG[0] }),
    .FrameData({\Tile_X8Y5_FrameData_O[31] ,
    \Tile_X8Y5_FrameData_O[30] ,
    \Tile_X8Y5_FrameData_O[29] ,
    \Tile_X8Y5_FrameData_O[28] ,
    \Tile_X8Y5_FrameData_O[27] ,
    \Tile_X8Y5_FrameData_O[26] ,
    \Tile_X8Y5_FrameData_O[25] ,
    \Tile_X8Y5_FrameData_O[24] ,
    \Tile_X8Y5_FrameData_O[23] ,
    \Tile_X8Y5_FrameData_O[22] ,
    \Tile_X8Y5_FrameData_O[21] ,
    \Tile_X8Y5_FrameData_O[20] ,
    \Tile_X8Y5_FrameData_O[19] ,
    \Tile_X8Y5_FrameData_O[18] ,
    \Tile_X8Y5_FrameData_O[17] ,
    \Tile_X8Y5_FrameData_O[16] ,
    \Tile_X8Y5_FrameData_O[15] ,
    \Tile_X8Y5_FrameData_O[14] ,
    \Tile_X8Y5_FrameData_O[13] ,
    \Tile_X8Y5_FrameData_O[12] ,
    \Tile_X8Y5_FrameData_O[11] ,
    \Tile_X8Y5_FrameData_O[10] ,
    \Tile_X8Y5_FrameData_O[9] ,
    \Tile_X8Y5_FrameData_O[8] ,
    \Tile_X8Y5_FrameData_O[7] ,
    \Tile_X8Y5_FrameData_O[6] ,
    \Tile_X8Y5_FrameData_O[5] ,
    \Tile_X8Y5_FrameData_O[4] ,
    \Tile_X8Y5_FrameData_O[3] ,
    \Tile_X8Y5_FrameData_O[2] ,
    \Tile_X8Y5_FrameData_O[1] ,
    \Tile_X8Y5_FrameData_O[0] }),
    .FrameData_O({\Tile_X9Y5_FrameData_O[31] ,
    \Tile_X9Y5_FrameData_O[30] ,
    \Tile_X9Y5_FrameData_O[29] ,
    \Tile_X9Y5_FrameData_O[28] ,
    \Tile_X9Y5_FrameData_O[27] ,
    \Tile_X9Y5_FrameData_O[26] ,
    \Tile_X9Y5_FrameData_O[25] ,
    \Tile_X9Y5_FrameData_O[24] ,
    \Tile_X9Y5_FrameData_O[23] ,
    \Tile_X9Y5_FrameData_O[22] ,
    \Tile_X9Y5_FrameData_O[21] ,
    \Tile_X9Y5_FrameData_O[20] ,
    \Tile_X9Y5_FrameData_O[19] ,
    \Tile_X9Y5_FrameData_O[18] ,
    \Tile_X9Y5_FrameData_O[17] ,
    \Tile_X9Y5_FrameData_O[16] ,
    \Tile_X9Y5_FrameData_O[15] ,
    \Tile_X9Y5_FrameData_O[14] ,
    \Tile_X9Y5_FrameData_O[13] ,
    \Tile_X9Y5_FrameData_O[12] ,
    \Tile_X9Y5_FrameData_O[11] ,
    \Tile_X9Y5_FrameData_O[10] ,
    \Tile_X9Y5_FrameData_O[9] ,
    \Tile_X9Y5_FrameData_O[8] ,
    \Tile_X9Y5_FrameData_O[7] ,
    \Tile_X9Y5_FrameData_O[6] ,
    \Tile_X9Y5_FrameData_O[5] ,
    \Tile_X9Y5_FrameData_O[4] ,
    \Tile_X9Y5_FrameData_O[3] ,
    \Tile_X9Y5_FrameData_O[2] ,
    \Tile_X9Y5_FrameData_O[1] ,
    \Tile_X9Y5_FrameData_O[0] }),
    .FrameStrobe({\Tile_X9Y6_FrameStrobe_O[19] ,
    \Tile_X9Y6_FrameStrobe_O[18] ,
    \Tile_X9Y6_FrameStrobe_O[17] ,
    \Tile_X9Y6_FrameStrobe_O[16] ,
    \Tile_X9Y6_FrameStrobe_O[15] ,
    \Tile_X9Y6_FrameStrobe_O[14] ,
    \Tile_X9Y6_FrameStrobe_O[13] ,
    \Tile_X9Y6_FrameStrobe_O[12] ,
    \Tile_X9Y6_FrameStrobe_O[11] ,
    \Tile_X9Y6_FrameStrobe_O[10] ,
    \Tile_X9Y6_FrameStrobe_O[9] ,
    \Tile_X9Y6_FrameStrobe_O[8] ,
    \Tile_X9Y6_FrameStrobe_O[7] ,
    \Tile_X9Y6_FrameStrobe_O[6] ,
    \Tile_X9Y6_FrameStrobe_O[5] ,
    \Tile_X9Y6_FrameStrobe_O[4] ,
    \Tile_X9Y6_FrameStrobe_O[3] ,
    \Tile_X9Y6_FrameStrobe_O[2] ,
    \Tile_X9Y6_FrameStrobe_O[1] ,
    \Tile_X9Y6_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X9Y5_FrameStrobe_O[19] ,
    \Tile_X9Y5_FrameStrobe_O[18] ,
    \Tile_X9Y5_FrameStrobe_O[17] ,
    \Tile_X9Y5_FrameStrobe_O[16] ,
    \Tile_X9Y5_FrameStrobe_O[15] ,
    \Tile_X9Y5_FrameStrobe_O[14] ,
    \Tile_X9Y5_FrameStrobe_O[13] ,
    \Tile_X9Y5_FrameStrobe_O[12] ,
    \Tile_X9Y5_FrameStrobe_O[11] ,
    \Tile_X9Y5_FrameStrobe_O[10] ,
    \Tile_X9Y5_FrameStrobe_O[9] ,
    \Tile_X9Y5_FrameStrobe_O[8] ,
    \Tile_X9Y5_FrameStrobe_O[7] ,
    \Tile_X9Y5_FrameStrobe_O[6] ,
    \Tile_X9Y5_FrameStrobe_O[5] ,
    \Tile_X9Y5_FrameStrobe_O[4] ,
    \Tile_X9Y5_FrameStrobe_O[3] ,
    \Tile_X9Y5_FrameStrobe_O[2] ,
    \Tile_X9Y5_FrameStrobe_O[1] ,
    \Tile_X9Y5_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X9Y5_N1BEG[3] ,
    \Tile_X9Y5_N1BEG[2] ,
    \Tile_X9Y5_N1BEG[1] ,
    \Tile_X9Y5_N1BEG[0] }),
    .N1END({\Tile_X9Y6_N1BEG[3] ,
    \Tile_X9Y6_N1BEG[2] ,
    \Tile_X9Y6_N1BEG[1] ,
    \Tile_X9Y6_N1BEG[0] }),
    .N2BEG({\Tile_X9Y5_N2BEG[7] ,
    \Tile_X9Y5_N2BEG[6] ,
    \Tile_X9Y5_N2BEG[5] ,
    \Tile_X9Y5_N2BEG[4] ,
    \Tile_X9Y5_N2BEG[3] ,
    \Tile_X9Y5_N2BEG[2] ,
    \Tile_X9Y5_N2BEG[1] ,
    \Tile_X9Y5_N2BEG[0] }),
    .N2BEGb({\Tile_X9Y5_N2BEGb[7] ,
    \Tile_X9Y5_N2BEGb[6] ,
    \Tile_X9Y5_N2BEGb[5] ,
    \Tile_X9Y5_N2BEGb[4] ,
    \Tile_X9Y5_N2BEGb[3] ,
    \Tile_X9Y5_N2BEGb[2] ,
    \Tile_X9Y5_N2BEGb[1] ,
    \Tile_X9Y5_N2BEGb[0] }),
    .N2END({\Tile_X9Y6_N2BEGb[7] ,
    \Tile_X9Y6_N2BEGb[6] ,
    \Tile_X9Y6_N2BEGb[5] ,
    \Tile_X9Y6_N2BEGb[4] ,
    \Tile_X9Y6_N2BEGb[3] ,
    \Tile_X9Y6_N2BEGb[2] ,
    \Tile_X9Y6_N2BEGb[1] ,
    \Tile_X9Y6_N2BEGb[0] }),
    .N2MID({\Tile_X9Y6_N2BEG[7] ,
    \Tile_X9Y6_N2BEG[6] ,
    \Tile_X9Y6_N2BEG[5] ,
    \Tile_X9Y6_N2BEG[4] ,
    \Tile_X9Y6_N2BEG[3] ,
    \Tile_X9Y6_N2BEG[2] ,
    \Tile_X9Y6_N2BEG[1] ,
    \Tile_X9Y6_N2BEG[0] }),
    .N4BEG({\Tile_X9Y5_N4BEG[15] ,
    \Tile_X9Y5_N4BEG[14] ,
    \Tile_X9Y5_N4BEG[13] ,
    \Tile_X9Y5_N4BEG[12] ,
    \Tile_X9Y5_N4BEG[11] ,
    \Tile_X9Y5_N4BEG[10] ,
    \Tile_X9Y5_N4BEG[9] ,
    \Tile_X9Y5_N4BEG[8] ,
    \Tile_X9Y5_N4BEG[7] ,
    \Tile_X9Y5_N4BEG[6] ,
    \Tile_X9Y5_N4BEG[5] ,
    \Tile_X9Y5_N4BEG[4] ,
    \Tile_X9Y5_N4BEG[3] ,
    \Tile_X9Y5_N4BEG[2] ,
    \Tile_X9Y5_N4BEG[1] ,
    \Tile_X9Y5_N4BEG[0] }),
    .N4END({\Tile_X9Y6_N4BEG[15] ,
    \Tile_X9Y6_N4BEG[14] ,
    \Tile_X9Y6_N4BEG[13] ,
    \Tile_X9Y6_N4BEG[12] ,
    \Tile_X9Y6_N4BEG[11] ,
    \Tile_X9Y6_N4BEG[10] ,
    \Tile_X9Y6_N4BEG[9] ,
    \Tile_X9Y6_N4BEG[8] ,
    \Tile_X9Y6_N4BEG[7] ,
    \Tile_X9Y6_N4BEG[6] ,
    \Tile_X9Y6_N4BEG[5] ,
    \Tile_X9Y6_N4BEG[4] ,
    \Tile_X9Y6_N4BEG[3] ,
    \Tile_X9Y6_N4BEG[2] ,
    \Tile_X9Y6_N4BEG[1] ,
    \Tile_X9Y6_N4BEG[0] }),
    .NN4BEG({\Tile_X9Y5_NN4BEG[15] ,
    \Tile_X9Y5_NN4BEG[14] ,
    \Tile_X9Y5_NN4BEG[13] ,
    \Tile_X9Y5_NN4BEG[12] ,
    \Tile_X9Y5_NN4BEG[11] ,
    \Tile_X9Y5_NN4BEG[10] ,
    \Tile_X9Y5_NN4BEG[9] ,
    \Tile_X9Y5_NN4BEG[8] ,
    \Tile_X9Y5_NN4BEG[7] ,
    \Tile_X9Y5_NN4BEG[6] ,
    \Tile_X9Y5_NN4BEG[5] ,
    \Tile_X9Y5_NN4BEG[4] ,
    \Tile_X9Y5_NN4BEG[3] ,
    \Tile_X9Y5_NN4BEG[2] ,
    \Tile_X9Y5_NN4BEG[1] ,
    \Tile_X9Y5_NN4BEG[0] }),
    .NN4END({\Tile_X9Y6_NN4BEG[15] ,
    \Tile_X9Y6_NN4BEG[14] ,
    \Tile_X9Y6_NN4BEG[13] ,
    \Tile_X9Y6_NN4BEG[12] ,
    \Tile_X9Y6_NN4BEG[11] ,
    \Tile_X9Y6_NN4BEG[10] ,
    \Tile_X9Y6_NN4BEG[9] ,
    \Tile_X9Y6_NN4BEG[8] ,
    \Tile_X9Y6_NN4BEG[7] ,
    \Tile_X9Y6_NN4BEG[6] ,
    \Tile_X9Y6_NN4BEG[5] ,
    \Tile_X9Y6_NN4BEG[4] ,
    \Tile_X9Y6_NN4BEG[3] ,
    \Tile_X9Y6_NN4BEG[2] ,
    \Tile_X9Y6_NN4BEG[1] ,
    \Tile_X9Y6_NN4BEG[0] }),
    .S1BEG({\Tile_X9Y5_S1BEG[3] ,
    \Tile_X9Y5_S1BEG[2] ,
    \Tile_X9Y5_S1BEG[1] ,
    \Tile_X9Y5_S1BEG[0] }),
    .S1END({\Tile_X9Y4_S1BEG[3] ,
    \Tile_X9Y4_S1BEG[2] ,
    \Tile_X9Y4_S1BEG[1] ,
    \Tile_X9Y4_S1BEG[0] }),
    .S2BEG({\Tile_X9Y5_S2BEG[7] ,
    \Tile_X9Y5_S2BEG[6] ,
    \Tile_X9Y5_S2BEG[5] ,
    \Tile_X9Y5_S2BEG[4] ,
    \Tile_X9Y5_S2BEG[3] ,
    \Tile_X9Y5_S2BEG[2] ,
    \Tile_X9Y5_S2BEG[1] ,
    \Tile_X9Y5_S2BEG[0] }),
    .S2BEGb({\Tile_X9Y5_S2BEGb[7] ,
    \Tile_X9Y5_S2BEGb[6] ,
    \Tile_X9Y5_S2BEGb[5] ,
    \Tile_X9Y5_S2BEGb[4] ,
    \Tile_X9Y5_S2BEGb[3] ,
    \Tile_X9Y5_S2BEGb[2] ,
    \Tile_X9Y5_S2BEGb[1] ,
    \Tile_X9Y5_S2BEGb[0] }),
    .S2END({\Tile_X9Y4_S2BEGb[7] ,
    \Tile_X9Y4_S2BEGb[6] ,
    \Tile_X9Y4_S2BEGb[5] ,
    \Tile_X9Y4_S2BEGb[4] ,
    \Tile_X9Y4_S2BEGb[3] ,
    \Tile_X9Y4_S2BEGb[2] ,
    \Tile_X9Y4_S2BEGb[1] ,
    \Tile_X9Y4_S2BEGb[0] }),
    .S2MID({\Tile_X9Y4_S2BEG[7] ,
    \Tile_X9Y4_S2BEG[6] ,
    \Tile_X9Y4_S2BEG[5] ,
    \Tile_X9Y4_S2BEG[4] ,
    \Tile_X9Y4_S2BEG[3] ,
    \Tile_X9Y4_S2BEG[2] ,
    \Tile_X9Y4_S2BEG[1] ,
    \Tile_X9Y4_S2BEG[0] }),
    .S4BEG({\Tile_X9Y5_S4BEG[15] ,
    \Tile_X9Y5_S4BEG[14] ,
    \Tile_X9Y5_S4BEG[13] ,
    \Tile_X9Y5_S4BEG[12] ,
    \Tile_X9Y5_S4BEG[11] ,
    \Tile_X9Y5_S4BEG[10] ,
    \Tile_X9Y5_S4BEG[9] ,
    \Tile_X9Y5_S4BEG[8] ,
    \Tile_X9Y5_S4BEG[7] ,
    \Tile_X9Y5_S4BEG[6] ,
    \Tile_X9Y5_S4BEG[5] ,
    \Tile_X9Y5_S4BEG[4] ,
    \Tile_X9Y5_S4BEG[3] ,
    \Tile_X9Y5_S4BEG[2] ,
    \Tile_X9Y5_S4BEG[1] ,
    \Tile_X9Y5_S4BEG[0] }),
    .S4END({\Tile_X9Y4_S4BEG[15] ,
    \Tile_X9Y4_S4BEG[14] ,
    \Tile_X9Y4_S4BEG[13] ,
    \Tile_X9Y4_S4BEG[12] ,
    \Tile_X9Y4_S4BEG[11] ,
    \Tile_X9Y4_S4BEG[10] ,
    \Tile_X9Y4_S4BEG[9] ,
    \Tile_X9Y4_S4BEG[8] ,
    \Tile_X9Y4_S4BEG[7] ,
    \Tile_X9Y4_S4BEG[6] ,
    \Tile_X9Y4_S4BEG[5] ,
    \Tile_X9Y4_S4BEG[4] ,
    \Tile_X9Y4_S4BEG[3] ,
    \Tile_X9Y4_S4BEG[2] ,
    \Tile_X9Y4_S4BEG[1] ,
    \Tile_X9Y4_S4BEG[0] }),
    .SS4BEG({\Tile_X9Y5_SS4BEG[15] ,
    \Tile_X9Y5_SS4BEG[14] ,
    \Tile_X9Y5_SS4BEG[13] ,
    \Tile_X9Y5_SS4BEG[12] ,
    \Tile_X9Y5_SS4BEG[11] ,
    \Tile_X9Y5_SS4BEG[10] ,
    \Tile_X9Y5_SS4BEG[9] ,
    \Tile_X9Y5_SS4BEG[8] ,
    \Tile_X9Y5_SS4BEG[7] ,
    \Tile_X9Y5_SS4BEG[6] ,
    \Tile_X9Y5_SS4BEG[5] ,
    \Tile_X9Y5_SS4BEG[4] ,
    \Tile_X9Y5_SS4BEG[3] ,
    \Tile_X9Y5_SS4BEG[2] ,
    \Tile_X9Y5_SS4BEG[1] ,
    \Tile_X9Y5_SS4BEG[0] }),
    .SS4END({\Tile_X9Y4_SS4BEG[15] ,
    \Tile_X9Y4_SS4BEG[14] ,
    \Tile_X9Y4_SS4BEG[13] ,
    \Tile_X9Y4_SS4BEG[12] ,
    \Tile_X9Y4_SS4BEG[11] ,
    \Tile_X9Y4_SS4BEG[10] ,
    \Tile_X9Y4_SS4BEG[9] ,
    \Tile_X9Y4_SS4BEG[8] ,
    \Tile_X9Y4_SS4BEG[7] ,
    \Tile_X9Y4_SS4BEG[6] ,
    \Tile_X9Y4_SS4BEG[5] ,
    \Tile_X9Y4_SS4BEG[4] ,
    \Tile_X9Y4_SS4BEG[3] ,
    \Tile_X9Y4_SS4BEG[2] ,
    \Tile_X9Y4_SS4BEG[1] ,
    \Tile_X9Y4_SS4BEG[0] }),
    .W1BEG({\Tile_X9Y5_W1BEG[3] ,
    \Tile_X9Y5_W1BEG[2] ,
    \Tile_X9Y5_W1BEG[1] ,
    \Tile_X9Y5_W1BEG[0] }),
    .W1END({\Tile_X10Y5_W1BEG[3] ,
    \Tile_X10Y5_W1BEG[2] ,
    \Tile_X10Y5_W1BEG[1] ,
    \Tile_X10Y5_W1BEG[0] }),
    .W2BEG({\Tile_X9Y5_W2BEG[7] ,
    \Tile_X9Y5_W2BEG[6] ,
    \Tile_X9Y5_W2BEG[5] ,
    \Tile_X9Y5_W2BEG[4] ,
    \Tile_X9Y5_W2BEG[3] ,
    \Tile_X9Y5_W2BEG[2] ,
    \Tile_X9Y5_W2BEG[1] ,
    \Tile_X9Y5_W2BEG[0] }),
    .W2BEGb({\Tile_X9Y5_W2BEGb[7] ,
    \Tile_X9Y5_W2BEGb[6] ,
    \Tile_X9Y5_W2BEGb[5] ,
    \Tile_X9Y5_W2BEGb[4] ,
    \Tile_X9Y5_W2BEGb[3] ,
    \Tile_X9Y5_W2BEGb[2] ,
    \Tile_X9Y5_W2BEGb[1] ,
    \Tile_X9Y5_W2BEGb[0] }),
    .W2END({\Tile_X10Y5_W2BEGb[7] ,
    \Tile_X10Y5_W2BEGb[6] ,
    \Tile_X10Y5_W2BEGb[5] ,
    \Tile_X10Y5_W2BEGb[4] ,
    \Tile_X10Y5_W2BEGb[3] ,
    \Tile_X10Y5_W2BEGb[2] ,
    \Tile_X10Y5_W2BEGb[1] ,
    \Tile_X10Y5_W2BEGb[0] }),
    .W2MID({\Tile_X10Y5_W2BEG[7] ,
    \Tile_X10Y5_W2BEG[6] ,
    \Tile_X10Y5_W2BEG[5] ,
    \Tile_X10Y5_W2BEG[4] ,
    \Tile_X10Y5_W2BEG[3] ,
    \Tile_X10Y5_W2BEG[2] ,
    \Tile_X10Y5_W2BEG[1] ,
    \Tile_X10Y5_W2BEG[0] }),
    .W6BEG({\Tile_X9Y5_W6BEG[11] ,
    \Tile_X9Y5_W6BEG[10] ,
    \Tile_X9Y5_W6BEG[9] ,
    \Tile_X9Y5_W6BEG[8] ,
    \Tile_X9Y5_W6BEG[7] ,
    \Tile_X9Y5_W6BEG[6] ,
    \Tile_X9Y5_W6BEG[5] ,
    \Tile_X9Y5_W6BEG[4] ,
    \Tile_X9Y5_W6BEG[3] ,
    \Tile_X9Y5_W6BEG[2] ,
    \Tile_X9Y5_W6BEG[1] ,
    \Tile_X9Y5_W6BEG[0] }),
    .W6END({\Tile_X10Y5_W6BEG[11] ,
    \Tile_X10Y5_W6BEG[10] ,
    \Tile_X10Y5_W6BEG[9] ,
    \Tile_X10Y5_W6BEG[8] ,
    \Tile_X10Y5_W6BEG[7] ,
    \Tile_X10Y5_W6BEG[6] ,
    \Tile_X10Y5_W6BEG[5] ,
    \Tile_X10Y5_W6BEG[4] ,
    \Tile_X10Y5_W6BEG[3] ,
    \Tile_X10Y5_W6BEG[2] ,
    \Tile_X10Y5_W6BEG[1] ,
    \Tile_X10Y5_W6BEG[0] }),
    .WW4BEG({\Tile_X9Y5_WW4BEG[15] ,
    \Tile_X9Y5_WW4BEG[14] ,
    \Tile_X9Y5_WW4BEG[13] ,
    \Tile_X9Y5_WW4BEG[12] ,
    \Tile_X9Y5_WW4BEG[11] ,
    \Tile_X9Y5_WW4BEG[10] ,
    \Tile_X9Y5_WW4BEG[9] ,
    \Tile_X9Y5_WW4BEG[8] ,
    \Tile_X9Y5_WW4BEG[7] ,
    \Tile_X9Y5_WW4BEG[6] ,
    \Tile_X9Y5_WW4BEG[5] ,
    \Tile_X9Y5_WW4BEG[4] ,
    \Tile_X9Y5_WW4BEG[3] ,
    \Tile_X9Y5_WW4BEG[2] ,
    \Tile_X9Y5_WW4BEG[1] ,
    \Tile_X9Y5_WW4BEG[0] }),
    .WW4END({\Tile_X10Y5_WW4BEG[15] ,
    \Tile_X10Y5_WW4BEG[14] ,
    \Tile_X10Y5_WW4BEG[13] ,
    \Tile_X10Y5_WW4BEG[12] ,
    \Tile_X10Y5_WW4BEG[11] ,
    \Tile_X10Y5_WW4BEG[10] ,
    \Tile_X10Y5_WW4BEG[9] ,
    \Tile_X10Y5_WW4BEG[8] ,
    \Tile_X10Y5_WW4BEG[7] ,
    \Tile_X10Y5_WW4BEG[6] ,
    \Tile_X10Y5_WW4BEG[5] ,
    \Tile_X10Y5_WW4BEG[4] ,
    \Tile_X10Y5_WW4BEG[3] ,
    \Tile_X10Y5_WW4BEG[2] ,
    \Tile_X10Y5_WW4BEG[1] ,
    \Tile_X10Y5_WW4BEG[0] }));
 LUT4AB Tile_X9Y6_LUT4AB (.Ci(Tile_X9Y7_Co),
    .Co(Tile_X9Y6_Co),
    .UserCLK(Tile_X9Y7_UserCLKo),
    .UserCLKo(Tile_X9Y6_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X9Y6_E1BEG[3] ,
    \Tile_X9Y6_E1BEG[2] ,
    \Tile_X9Y6_E1BEG[1] ,
    \Tile_X9Y6_E1BEG[0] }),
    .E1END({\Tile_X8Y6_E1BEG[3] ,
    \Tile_X8Y6_E1BEG[2] ,
    \Tile_X8Y6_E1BEG[1] ,
    \Tile_X8Y6_E1BEG[0] }),
    .E2BEG({\Tile_X9Y6_E2BEG[7] ,
    \Tile_X9Y6_E2BEG[6] ,
    \Tile_X9Y6_E2BEG[5] ,
    \Tile_X9Y6_E2BEG[4] ,
    \Tile_X9Y6_E2BEG[3] ,
    \Tile_X9Y6_E2BEG[2] ,
    \Tile_X9Y6_E2BEG[1] ,
    \Tile_X9Y6_E2BEG[0] }),
    .E2BEGb({\Tile_X9Y6_E2BEGb[7] ,
    \Tile_X9Y6_E2BEGb[6] ,
    \Tile_X9Y6_E2BEGb[5] ,
    \Tile_X9Y6_E2BEGb[4] ,
    \Tile_X9Y6_E2BEGb[3] ,
    \Tile_X9Y6_E2BEGb[2] ,
    \Tile_X9Y6_E2BEGb[1] ,
    \Tile_X9Y6_E2BEGb[0] }),
    .E2END({\Tile_X8Y6_E2BEGb[7] ,
    \Tile_X8Y6_E2BEGb[6] ,
    \Tile_X8Y6_E2BEGb[5] ,
    \Tile_X8Y6_E2BEGb[4] ,
    \Tile_X8Y6_E2BEGb[3] ,
    \Tile_X8Y6_E2BEGb[2] ,
    \Tile_X8Y6_E2BEGb[1] ,
    \Tile_X8Y6_E2BEGb[0] }),
    .E2MID({\Tile_X8Y6_E2BEG[7] ,
    \Tile_X8Y6_E2BEG[6] ,
    \Tile_X8Y6_E2BEG[5] ,
    \Tile_X8Y6_E2BEG[4] ,
    \Tile_X8Y6_E2BEG[3] ,
    \Tile_X8Y6_E2BEG[2] ,
    \Tile_X8Y6_E2BEG[1] ,
    \Tile_X8Y6_E2BEG[0] }),
    .E6BEG({\Tile_X9Y6_E6BEG[11] ,
    \Tile_X9Y6_E6BEG[10] ,
    \Tile_X9Y6_E6BEG[9] ,
    \Tile_X9Y6_E6BEG[8] ,
    \Tile_X9Y6_E6BEG[7] ,
    \Tile_X9Y6_E6BEG[6] ,
    \Tile_X9Y6_E6BEG[5] ,
    \Tile_X9Y6_E6BEG[4] ,
    \Tile_X9Y6_E6BEG[3] ,
    \Tile_X9Y6_E6BEG[2] ,
    \Tile_X9Y6_E6BEG[1] ,
    \Tile_X9Y6_E6BEG[0] }),
    .E6END({\Tile_X8Y6_E6BEG[11] ,
    \Tile_X8Y6_E6BEG[10] ,
    \Tile_X8Y6_E6BEG[9] ,
    \Tile_X8Y6_E6BEG[8] ,
    \Tile_X8Y6_E6BEG[7] ,
    \Tile_X8Y6_E6BEG[6] ,
    \Tile_X8Y6_E6BEG[5] ,
    \Tile_X8Y6_E6BEG[4] ,
    \Tile_X8Y6_E6BEG[3] ,
    \Tile_X8Y6_E6BEG[2] ,
    \Tile_X8Y6_E6BEG[1] ,
    \Tile_X8Y6_E6BEG[0] }),
    .EE4BEG({\Tile_X9Y6_EE4BEG[15] ,
    \Tile_X9Y6_EE4BEG[14] ,
    \Tile_X9Y6_EE4BEG[13] ,
    \Tile_X9Y6_EE4BEG[12] ,
    \Tile_X9Y6_EE4BEG[11] ,
    \Tile_X9Y6_EE4BEG[10] ,
    \Tile_X9Y6_EE4BEG[9] ,
    \Tile_X9Y6_EE4BEG[8] ,
    \Tile_X9Y6_EE4BEG[7] ,
    \Tile_X9Y6_EE4BEG[6] ,
    \Tile_X9Y6_EE4BEG[5] ,
    \Tile_X9Y6_EE4BEG[4] ,
    \Tile_X9Y6_EE4BEG[3] ,
    \Tile_X9Y6_EE4BEG[2] ,
    \Tile_X9Y6_EE4BEG[1] ,
    \Tile_X9Y6_EE4BEG[0] }),
    .EE4END({\Tile_X8Y6_EE4BEG[15] ,
    \Tile_X8Y6_EE4BEG[14] ,
    \Tile_X8Y6_EE4BEG[13] ,
    \Tile_X8Y6_EE4BEG[12] ,
    \Tile_X8Y6_EE4BEG[11] ,
    \Tile_X8Y6_EE4BEG[10] ,
    \Tile_X8Y6_EE4BEG[9] ,
    \Tile_X8Y6_EE4BEG[8] ,
    \Tile_X8Y6_EE4BEG[7] ,
    \Tile_X8Y6_EE4BEG[6] ,
    \Tile_X8Y6_EE4BEG[5] ,
    \Tile_X8Y6_EE4BEG[4] ,
    \Tile_X8Y6_EE4BEG[3] ,
    \Tile_X8Y6_EE4BEG[2] ,
    \Tile_X8Y6_EE4BEG[1] ,
    \Tile_X8Y6_EE4BEG[0] }),
    .FrameData({\Tile_X8Y6_FrameData_O[31] ,
    \Tile_X8Y6_FrameData_O[30] ,
    \Tile_X8Y6_FrameData_O[29] ,
    \Tile_X8Y6_FrameData_O[28] ,
    \Tile_X8Y6_FrameData_O[27] ,
    \Tile_X8Y6_FrameData_O[26] ,
    \Tile_X8Y6_FrameData_O[25] ,
    \Tile_X8Y6_FrameData_O[24] ,
    \Tile_X8Y6_FrameData_O[23] ,
    \Tile_X8Y6_FrameData_O[22] ,
    \Tile_X8Y6_FrameData_O[21] ,
    \Tile_X8Y6_FrameData_O[20] ,
    \Tile_X8Y6_FrameData_O[19] ,
    \Tile_X8Y6_FrameData_O[18] ,
    \Tile_X8Y6_FrameData_O[17] ,
    \Tile_X8Y6_FrameData_O[16] ,
    \Tile_X8Y6_FrameData_O[15] ,
    \Tile_X8Y6_FrameData_O[14] ,
    \Tile_X8Y6_FrameData_O[13] ,
    \Tile_X8Y6_FrameData_O[12] ,
    \Tile_X8Y6_FrameData_O[11] ,
    \Tile_X8Y6_FrameData_O[10] ,
    \Tile_X8Y6_FrameData_O[9] ,
    \Tile_X8Y6_FrameData_O[8] ,
    \Tile_X8Y6_FrameData_O[7] ,
    \Tile_X8Y6_FrameData_O[6] ,
    \Tile_X8Y6_FrameData_O[5] ,
    \Tile_X8Y6_FrameData_O[4] ,
    \Tile_X8Y6_FrameData_O[3] ,
    \Tile_X8Y6_FrameData_O[2] ,
    \Tile_X8Y6_FrameData_O[1] ,
    \Tile_X8Y6_FrameData_O[0] }),
    .FrameData_O({\Tile_X9Y6_FrameData_O[31] ,
    \Tile_X9Y6_FrameData_O[30] ,
    \Tile_X9Y6_FrameData_O[29] ,
    \Tile_X9Y6_FrameData_O[28] ,
    \Tile_X9Y6_FrameData_O[27] ,
    \Tile_X9Y6_FrameData_O[26] ,
    \Tile_X9Y6_FrameData_O[25] ,
    \Tile_X9Y6_FrameData_O[24] ,
    \Tile_X9Y6_FrameData_O[23] ,
    \Tile_X9Y6_FrameData_O[22] ,
    \Tile_X9Y6_FrameData_O[21] ,
    \Tile_X9Y6_FrameData_O[20] ,
    \Tile_X9Y6_FrameData_O[19] ,
    \Tile_X9Y6_FrameData_O[18] ,
    \Tile_X9Y6_FrameData_O[17] ,
    \Tile_X9Y6_FrameData_O[16] ,
    \Tile_X9Y6_FrameData_O[15] ,
    \Tile_X9Y6_FrameData_O[14] ,
    \Tile_X9Y6_FrameData_O[13] ,
    \Tile_X9Y6_FrameData_O[12] ,
    \Tile_X9Y6_FrameData_O[11] ,
    \Tile_X9Y6_FrameData_O[10] ,
    \Tile_X9Y6_FrameData_O[9] ,
    \Tile_X9Y6_FrameData_O[8] ,
    \Tile_X9Y6_FrameData_O[7] ,
    \Tile_X9Y6_FrameData_O[6] ,
    \Tile_X9Y6_FrameData_O[5] ,
    \Tile_X9Y6_FrameData_O[4] ,
    \Tile_X9Y6_FrameData_O[3] ,
    \Tile_X9Y6_FrameData_O[2] ,
    \Tile_X9Y6_FrameData_O[1] ,
    \Tile_X9Y6_FrameData_O[0] }),
    .FrameStrobe({\Tile_X9Y7_FrameStrobe_O[19] ,
    \Tile_X9Y7_FrameStrobe_O[18] ,
    \Tile_X9Y7_FrameStrobe_O[17] ,
    \Tile_X9Y7_FrameStrobe_O[16] ,
    \Tile_X9Y7_FrameStrobe_O[15] ,
    \Tile_X9Y7_FrameStrobe_O[14] ,
    \Tile_X9Y7_FrameStrobe_O[13] ,
    \Tile_X9Y7_FrameStrobe_O[12] ,
    \Tile_X9Y7_FrameStrobe_O[11] ,
    \Tile_X9Y7_FrameStrobe_O[10] ,
    \Tile_X9Y7_FrameStrobe_O[9] ,
    \Tile_X9Y7_FrameStrobe_O[8] ,
    \Tile_X9Y7_FrameStrobe_O[7] ,
    \Tile_X9Y7_FrameStrobe_O[6] ,
    \Tile_X9Y7_FrameStrobe_O[5] ,
    \Tile_X9Y7_FrameStrobe_O[4] ,
    \Tile_X9Y7_FrameStrobe_O[3] ,
    \Tile_X9Y7_FrameStrobe_O[2] ,
    \Tile_X9Y7_FrameStrobe_O[1] ,
    \Tile_X9Y7_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X9Y6_FrameStrobe_O[19] ,
    \Tile_X9Y6_FrameStrobe_O[18] ,
    \Tile_X9Y6_FrameStrobe_O[17] ,
    \Tile_X9Y6_FrameStrobe_O[16] ,
    \Tile_X9Y6_FrameStrobe_O[15] ,
    \Tile_X9Y6_FrameStrobe_O[14] ,
    \Tile_X9Y6_FrameStrobe_O[13] ,
    \Tile_X9Y6_FrameStrobe_O[12] ,
    \Tile_X9Y6_FrameStrobe_O[11] ,
    \Tile_X9Y6_FrameStrobe_O[10] ,
    \Tile_X9Y6_FrameStrobe_O[9] ,
    \Tile_X9Y6_FrameStrobe_O[8] ,
    \Tile_X9Y6_FrameStrobe_O[7] ,
    \Tile_X9Y6_FrameStrobe_O[6] ,
    \Tile_X9Y6_FrameStrobe_O[5] ,
    \Tile_X9Y6_FrameStrobe_O[4] ,
    \Tile_X9Y6_FrameStrobe_O[3] ,
    \Tile_X9Y6_FrameStrobe_O[2] ,
    \Tile_X9Y6_FrameStrobe_O[1] ,
    \Tile_X9Y6_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X9Y6_N1BEG[3] ,
    \Tile_X9Y6_N1BEG[2] ,
    \Tile_X9Y6_N1BEG[1] ,
    \Tile_X9Y6_N1BEG[0] }),
    .N1END({\Tile_X9Y7_N1BEG[3] ,
    \Tile_X9Y7_N1BEG[2] ,
    \Tile_X9Y7_N1BEG[1] ,
    \Tile_X9Y7_N1BEG[0] }),
    .N2BEG({\Tile_X9Y6_N2BEG[7] ,
    \Tile_X9Y6_N2BEG[6] ,
    \Tile_X9Y6_N2BEG[5] ,
    \Tile_X9Y6_N2BEG[4] ,
    \Tile_X9Y6_N2BEG[3] ,
    \Tile_X9Y6_N2BEG[2] ,
    \Tile_X9Y6_N2BEG[1] ,
    \Tile_X9Y6_N2BEG[0] }),
    .N2BEGb({\Tile_X9Y6_N2BEGb[7] ,
    \Tile_X9Y6_N2BEGb[6] ,
    \Tile_X9Y6_N2BEGb[5] ,
    \Tile_X9Y6_N2BEGb[4] ,
    \Tile_X9Y6_N2BEGb[3] ,
    \Tile_X9Y6_N2BEGb[2] ,
    \Tile_X9Y6_N2BEGb[1] ,
    \Tile_X9Y6_N2BEGb[0] }),
    .N2END({\Tile_X9Y7_N2BEGb[7] ,
    \Tile_X9Y7_N2BEGb[6] ,
    \Tile_X9Y7_N2BEGb[5] ,
    \Tile_X9Y7_N2BEGb[4] ,
    \Tile_X9Y7_N2BEGb[3] ,
    \Tile_X9Y7_N2BEGb[2] ,
    \Tile_X9Y7_N2BEGb[1] ,
    \Tile_X9Y7_N2BEGb[0] }),
    .N2MID({\Tile_X9Y7_N2BEG[7] ,
    \Tile_X9Y7_N2BEG[6] ,
    \Tile_X9Y7_N2BEG[5] ,
    \Tile_X9Y7_N2BEG[4] ,
    \Tile_X9Y7_N2BEG[3] ,
    \Tile_X9Y7_N2BEG[2] ,
    \Tile_X9Y7_N2BEG[1] ,
    \Tile_X9Y7_N2BEG[0] }),
    .N4BEG({\Tile_X9Y6_N4BEG[15] ,
    \Tile_X9Y6_N4BEG[14] ,
    \Tile_X9Y6_N4BEG[13] ,
    \Tile_X9Y6_N4BEG[12] ,
    \Tile_X9Y6_N4BEG[11] ,
    \Tile_X9Y6_N4BEG[10] ,
    \Tile_X9Y6_N4BEG[9] ,
    \Tile_X9Y6_N4BEG[8] ,
    \Tile_X9Y6_N4BEG[7] ,
    \Tile_X9Y6_N4BEG[6] ,
    \Tile_X9Y6_N4BEG[5] ,
    \Tile_X9Y6_N4BEG[4] ,
    \Tile_X9Y6_N4BEG[3] ,
    \Tile_X9Y6_N4BEG[2] ,
    \Tile_X9Y6_N4BEG[1] ,
    \Tile_X9Y6_N4BEG[0] }),
    .N4END({\Tile_X9Y7_N4BEG[15] ,
    \Tile_X9Y7_N4BEG[14] ,
    \Tile_X9Y7_N4BEG[13] ,
    \Tile_X9Y7_N4BEG[12] ,
    \Tile_X9Y7_N4BEG[11] ,
    \Tile_X9Y7_N4BEG[10] ,
    \Tile_X9Y7_N4BEG[9] ,
    \Tile_X9Y7_N4BEG[8] ,
    \Tile_X9Y7_N4BEG[7] ,
    \Tile_X9Y7_N4BEG[6] ,
    \Tile_X9Y7_N4BEG[5] ,
    \Tile_X9Y7_N4BEG[4] ,
    \Tile_X9Y7_N4BEG[3] ,
    \Tile_X9Y7_N4BEG[2] ,
    \Tile_X9Y7_N4BEG[1] ,
    \Tile_X9Y7_N4BEG[0] }),
    .NN4BEG({\Tile_X9Y6_NN4BEG[15] ,
    \Tile_X9Y6_NN4BEG[14] ,
    \Tile_X9Y6_NN4BEG[13] ,
    \Tile_X9Y6_NN4BEG[12] ,
    \Tile_X9Y6_NN4BEG[11] ,
    \Tile_X9Y6_NN4BEG[10] ,
    \Tile_X9Y6_NN4BEG[9] ,
    \Tile_X9Y6_NN4BEG[8] ,
    \Tile_X9Y6_NN4BEG[7] ,
    \Tile_X9Y6_NN4BEG[6] ,
    \Tile_X9Y6_NN4BEG[5] ,
    \Tile_X9Y6_NN4BEG[4] ,
    \Tile_X9Y6_NN4BEG[3] ,
    \Tile_X9Y6_NN4BEG[2] ,
    \Tile_X9Y6_NN4BEG[1] ,
    \Tile_X9Y6_NN4BEG[0] }),
    .NN4END({\Tile_X9Y7_NN4BEG[15] ,
    \Tile_X9Y7_NN4BEG[14] ,
    \Tile_X9Y7_NN4BEG[13] ,
    \Tile_X9Y7_NN4BEG[12] ,
    \Tile_X9Y7_NN4BEG[11] ,
    \Tile_X9Y7_NN4BEG[10] ,
    \Tile_X9Y7_NN4BEG[9] ,
    \Tile_X9Y7_NN4BEG[8] ,
    \Tile_X9Y7_NN4BEG[7] ,
    \Tile_X9Y7_NN4BEG[6] ,
    \Tile_X9Y7_NN4BEG[5] ,
    \Tile_X9Y7_NN4BEG[4] ,
    \Tile_X9Y7_NN4BEG[3] ,
    \Tile_X9Y7_NN4BEG[2] ,
    \Tile_X9Y7_NN4BEG[1] ,
    \Tile_X9Y7_NN4BEG[0] }),
    .S1BEG({\Tile_X9Y6_S1BEG[3] ,
    \Tile_X9Y6_S1BEG[2] ,
    \Tile_X9Y6_S1BEG[1] ,
    \Tile_X9Y6_S1BEG[0] }),
    .S1END({\Tile_X9Y5_S1BEG[3] ,
    \Tile_X9Y5_S1BEG[2] ,
    \Tile_X9Y5_S1BEG[1] ,
    \Tile_X9Y5_S1BEG[0] }),
    .S2BEG({\Tile_X9Y6_S2BEG[7] ,
    \Tile_X9Y6_S2BEG[6] ,
    \Tile_X9Y6_S2BEG[5] ,
    \Tile_X9Y6_S2BEG[4] ,
    \Tile_X9Y6_S2BEG[3] ,
    \Tile_X9Y6_S2BEG[2] ,
    \Tile_X9Y6_S2BEG[1] ,
    \Tile_X9Y6_S2BEG[0] }),
    .S2BEGb({\Tile_X9Y6_S2BEGb[7] ,
    \Tile_X9Y6_S2BEGb[6] ,
    \Tile_X9Y6_S2BEGb[5] ,
    \Tile_X9Y6_S2BEGb[4] ,
    \Tile_X9Y6_S2BEGb[3] ,
    \Tile_X9Y6_S2BEGb[2] ,
    \Tile_X9Y6_S2BEGb[1] ,
    \Tile_X9Y6_S2BEGb[0] }),
    .S2END({\Tile_X9Y5_S2BEGb[7] ,
    \Tile_X9Y5_S2BEGb[6] ,
    \Tile_X9Y5_S2BEGb[5] ,
    \Tile_X9Y5_S2BEGb[4] ,
    \Tile_X9Y5_S2BEGb[3] ,
    \Tile_X9Y5_S2BEGb[2] ,
    \Tile_X9Y5_S2BEGb[1] ,
    \Tile_X9Y5_S2BEGb[0] }),
    .S2MID({\Tile_X9Y5_S2BEG[7] ,
    \Tile_X9Y5_S2BEG[6] ,
    \Tile_X9Y5_S2BEG[5] ,
    \Tile_X9Y5_S2BEG[4] ,
    \Tile_X9Y5_S2BEG[3] ,
    \Tile_X9Y5_S2BEG[2] ,
    \Tile_X9Y5_S2BEG[1] ,
    \Tile_X9Y5_S2BEG[0] }),
    .S4BEG({\Tile_X9Y6_S4BEG[15] ,
    \Tile_X9Y6_S4BEG[14] ,
    \Tile_X9Y6_S4BEG[13] ,
    \Tile_X9Y6_S4BEG[12] ,
    \Tile_X9Y6_S4BEG[11] ,
    \Tile_X9Y6_S4BEG[10] ,
    \Tile_X9Y6_S4BEG[9] ,
    \Tile_X9Y6_S4BEG[8] ,
    \Tile_X9Y6_S4BEG[7] ,
    \Tile_X9Y6_S4BEG[6] ,
    \Tile_X9Y6_S4BEG[5] ,
    \Tile_X9Y6_S4BEG[4] ,
    \Tile_X9Y6_S4BEG[3] ,
    \Tile_X9Y6_S4BEG[2] ,
    \Tile_X9Y6_S4BEG[1] ,
    \Tile_X9Y6_S4BEG[0] }),
    .S4END({\Tile_X9Y5_S4BEG[15] ,
    \Tile_X9Y5_S4BEG[14] ,
    \Tile_X9Y5_S4BEG[13] ,
    \Tile_X9Y5_S4BEG[12] ,
    \Tile_X9Y5_S4BEG[11] ,
    \Tile_X9Y5_S4BEG[10] ,
    \Tile_X9Y5_S4BEG[9] ,
    \Tile_X9Y5_S4BEG[8] ,
    \Tile_X9Y5_S4BEG[7] ,
    \Tile_X9Y5_S4BEG[6] ,
    \Tile_X9Y5_S4BEG[5] ,
    \Tile_X9Y5_S4BEG[4] ,
    \Tile_X9Y5_S4BEG[3] ,
    \Tile_X9Y5_S4BEG[2] ,
    \Tile_X9Y5_S4BEG[1] ,
    \Tile_X9Y5_S4BEG[0] }),
    .SS4BEG({\Tile_X9Y6_SS4BEG[15] ,
    \Tile_X9Y6_SS4BEG[14] ,
    \Tile_X9Y6_SS4BEG[13] ,
    \Tile_X9Y6_SS4BEG[12] ,
    \Tile_X9Y6_SS4BEG[11] ,
    \Tile_X9Y6_SS4BEG[10] ,
    \Tile_X9Y6_SS4BEG[9] ,
    \Tile_X9Y6_SS4BEG[8] ,
    \Tile_X9Y6_SS4BEG[7] ,
    \Tile_X9Y6_SS4BEG[6] ,
    \Tile_X9Y6_SS4BEG[5] ,
    \Tile_X9Y6_SS4BEG[4] ,
    \Tile_X9Y6_SS4BEG[3] ,
    \Tile_X9Y6_SS4BEG[2] ,
    \Tile_X9Y6_SS4BEG[1] ,
    \Tile_X9Y6_SS4BEG[0] }),
    .SS4END({\Tile_X9Y5_SS4BEG[15] ,
    \Tile_X9Y5_SS4BEG[14] ,
    \Tile_X9Y5_SS4BEG[13] ,
    \Tile_X9Y5_SS4BEG[12] ,
    \Tile_X9Y5_SS4BEG[11] ,
    \Tile_X9Y5_SS4BEG[10] ,
    \Tile_X9Y5_SS4BEG[9] ,
    \Tile_X9Y5_SS4BEG[8] ,
    \Tile_X9Y5_SS4BEG[7] ,
    \Tile_X9Y5_SS4BEG[6] ,
    \Tile_X9Y5_SS4BEG[5] ,
    \Tile_X9Y5_SS4BEG[4] ,
    \Tile_X9Y5_SS4BEG[3] ,
    \Tile_X9Y5_SS4BEG[2] ,
    \Tile_X9Y5_SS4BEG[1] ,
    \Tile_X9Y5_SS4BEG[0] }),
    .W1BEG({\Tile_X9Y6_W1BEG[3] ,
    \Tile_X9Y6_W1BEG[2] ,
    \Tile_X9Y6_W1BEG[1] ,
    \Tile_X9Y6_W1BEG[0] }),
    .W1END({\Tile_X10Y6_W1BEG[3] ,
    \Tile_X10Y6_W1BEG[2] ,
    \Tile_X10Y6_W1BEG[1] ,
    \Tile_X10Y6_W1BEG[0] }),
    .W2BEG({\Tile_X9Y6_W2BEG[7] ,
    \Tile_X9Y6_W2BEG[6] ,
    \Tile_X9Y6_W2BEG[5] ,
    \Tile_X9Y6_W2BEG[4] ,
    \Tile_X9Y6_W2BEG[3] ,
    \Tile_X9Y6_W2BEG[2] ,
    \Tile_X9Y6_W2BEG[1] ,
    \Tile_X9Y6_W2BEG[0] }),
    .W2BEGb({\Tile_X9Y6_W2BEGb[7] ,
    \Tile_X9Y6_W2BEGb[6] ,
    \Tile_X9Y6_W2BEGb[5] ,
    \Tile_X9Y6_W2BEGb[4] ,
    \Tile_X9Y6_W2BEGb[3] ,
    \Tile_X9Y6_W2BEGb[2] ,
    \Tile_X9Y6_W2BEGb[1] ,
    \Tile_X9Y6_W2BEGb[0] }),
    .W2END({\Tile_X10Y6_W2BEGb[7] ,
    \Tile_X10Y6_W2BEGb[6] ,
    \Tile_X10Y6_W2BEGb[5] ,
    \Tile_X10Y6_W2BEGb[4] ,
    \Tile_X10Y6_W2BEGb[3] ,
    \Tile_X10Y6_W2BEGb[2] ,
    \Tile_X10Y6_W2BEGb[1] ,
    \Tile_X10Y6_W2BEGb[0] }),
    .W2MID({\Tile_X10Y6_W2BEG[7] ,
    \Tile_X10Y6_W2BEG[6] ,
    \Tile_X10Y6_W2BEG[5] ,
    \Tile_X10Y6_W2BEG[4] ,
    \Tile_X10Y6_W2BEG[3] ,
    \Tile_X10Y6_W2BEG[2] ,
    \Tile_X10Y6_W2BEG[1] ,
    \Tile_X10Y6_W2BEG[0] }),
    .W6BEG({\Tile_X9Y6_W6BEG[11] ,
    \Tile_X9Y6_W6BEG[10] ,
    \Tile_X9Y6_W6BEG[9] ,
    \Tile_X9Y6_W6BEG[8] ,
    \Tile_X9Y6_W6BEG[7] ,
    \Tile_X9Y6_W6BEG[6] ,
    \Tile_X9Y6_W6BEG[5] ,
    \Tile_X9Y6_W6BEG[4] ,
    \Tile_X9Y6_W6BEG[3] ,
    \Tile_X9Y6_W6BEG[2] ,
    \Tile_X9Y6_W6BEG[1] ,
    \Tile_X9Y6_W6BEG[0] }),
    .W6END({\Tile_X10Y6_W6BEG[11] ,
    \Tile_X10Y6_W6BEG[10] ,
    \Tile_X10Y6_W6BEG[9] ,
    \Tile_X10Y6_W6BEG[8] ,
    \Tile_X10Y6_W6BEG[7] ,
    \Tile_X10Y6_W6BEG[6] ,
    \Tile_X10Y6_W6BEG[5] ,
    \Tile_X10Y6_W6BEG[4] ,
    \Tile_X10Y6_W6BEG[3] ,
    \Tile_X10Y6_W6BEG[2] ,
    \Tile_X10Y6_W6BEG[1] ,
    \Tile_X10Y6_W6BEG[0] }),
    .WW4BEG({\Tile_X9Y6_WW4BEG[15] ,
    \Tile_X9Y6_WW4BEG[14] ,
    \Tile_X9Y6_WW4BEG[13] ,
    \Tile_X9Y6_WW4BEG[12] ,
    \Tile_X9Y6_WW4BEG[11] ,
    \Tile_X9Y6_WW4BEG[10] ,
    \Tile_X9Y6_WW4BEG[9] ,
    \Tile_X9Y6_WW4BEG[8] ,
    \Tile_X9Y6_WW4BEG[7] ,
    \Tile_X9Y6_WW4BEG[6] ,
    \Tile_X9Y6_WW4BEG[5] ,
    \Tile_X9Y6_WW4BEG[4] ,
    \Tile_X9Y6_WW4BEG[3] ,
    \Tile_X9Y6_WW4BEG[2] ,
    \Tile_X9Y6_WW4BEG[1] ,
    \Tile_X9Y6_WW4BEG[0] }),
    .WW4END({\Tile_X10Y6_WW4BEG[15] ,
    \Tile_X10Y6_WW4BEG[14] ,
    \Tile_X10Y6_WW4BEG[13] ,
    \Tile_X10Y6_WW4BEG[12] ,
    \Tile_X10Y6_WW4BEG[11] ,
    \Tile_X10Y6_WW4BEG[10] ,
    \Tile_X10Y6_WW4BEG[9] ,
    \Tile_X10Y6_WW4BEG[8] ,
    \Tile_X10Y6_WW4BEG[7] ,
    \Tile_X10Y6_WW4BEG[6] ,
    \Tile_X10Y6_WW4BEG[5] ,
    \Tile_X10Y6_WW4BEG[4] ,
    \Tile_X10Y6_WW4BEG[3] ,
    \Tile_X10Y6_WW4BEG[2] ,
    \Tile_X10Y6_WW4BEG[1] ,
    \Tile_X10Y6_WW4BEG[0] }));
 LUT4AB Tile_X9Y7_LUT4AB (.Ci(Tile_X9Y8_Co),
    .Co(Tile_X9Y7_Co),
    .UserCLK(Tile_X9Y8_UserCLKo),
    .UserCLKo(Tile_X9Y7_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X9Y7_E1BEG[3] ,
    \Tile_X9Y7_E1BEG[2] ,
    \Tile_X9Y7_E1BEG[1] ,
    \Tile_X9Y7_E1BEG[0] }),
    .E1END({\Tile_X8Y7_E1BEG[3] ,
    \Tile_X8Y7_E1BEG[2] ,
    \Tile_X8Y7_E1BEG[1] ,
    \Tile_X8Y7_E1BEG[0] }),
    .E2BEG({\Tile_X9Y7_E2BEG[7] ,
    \Tile_X9Y7_E2BEG[6] ,
    \Tile_X9Y7_E2BEG[5] ,
    \Tile_X9Y7_E2BEG[4] ,
    \Tile_X9Y7_E2BEG[3] ,
    \Tile_X9Y7_E2BEG[2] ,
    \Tile_X9Y7_E2BEG[1] ,
    \Tile_X9Y7_E2BEG[0] }),
    .E2BEGb({\Tile_X9Y7_E2BEGb[7] ,
    \Tile_X9Y7_E2BEGb[6] ,
    \Tile_X9Y7_E2BEGb[5] ,
    \Tile_X9Y7_E2BEGb[4] ,
    \Tile_X9Y7_E2BEGb[3] ,
    \Tile_X9Y7_E2BEGb[2] ,
    \Tile_X9Y7_E2BEGb[1] ,
    \Tile_X9Y7_E2BEGb[0] }),
    .E2END({\Tile_X8Y7_E2BEGb[7] ,
    \Tile_X8Y7_E2BEGb[6] ,
    \Tile_X8Y7_E2BEGb[5] ,
    \Tile_X8Y7_E2BEGb[4] ,
    \Tile_X8Y7_E2BEGb[3] ,
    \Tile_X8Y7_E2BEGb[2] ,
    \Tile_X8Y7_E2BEGb[1] ,
    \Tile_X8Y7_E2BEGb[0] }),
    .E2MID({\Tile_X8Y7_E2BEG[7] ,
    \Tile_X8Y7_E2BEG[6] ,
    \Tile_X8Y7_E2BEG[5] ,
    \Tile_X8Y7_E2BEG[4] ,
    \Tile_X8Y7_E2BEG[3] ,
    \Tile_X8Y7_E2BEG[2] ,
    \Tile_X8Y7_E2BEG[1] ,
    \Tile_X8Y7_E2BEG[0] }),
    .E6BEG({\Tile_X9Y7_E6BEG[11] ,
    \Tile_X9Y7_E6BEG[10] ,
    \Tile_X9Y7_E6BEG[9] ,
    \Tile_X9Y7_E6BEG[8] ,
    \Tile_X9Y7_E6BEG[7] ,
    \Tile_X9Y7_E6BEG[6] ,
    \Tile_X9Y7_E6BEG[5] ,
    \Tile_X9Y7_E6BEG[4] ,
    \Tile_X9Y7_E6BEG[3] ,
    \Tile_X9Y7_E6BEG[2] ,
    \Tile_X9Y7_E6BEG[1] ,
    \Tile_X9Y7_E6BEG[0] }),
    .E6END({\Tile_X8Y7_E6BEG[11] ,
    \Tile_X8Y7_E6BEG[10] ,
    \Tile_X8Y7_E6BEG[9] ,
    \Tile_X8Y7_E6BEG[8] ,
    \Tile_X8Y7_E6BEG[7] ,
    \Tile_X8Y7_E6BEG[6] ,
    \Tile_X8Y7_E6BEG[5] ,
    \Tile_X8Y7_E6BEG[4] ,
    \Tile_X8Y7_E6BEG[3] ,
    \Tile_X8Y7_E6BEG[2] ,
    \Tile_X8Y7_E6BEG[1] ,
    \Tile_X8Y7_E6BEG[0] }),
    .EE4BEG({\Tile_X9Y7_EE4BEG[15] ,
    \Tile_X9Y7_EE4BEG[14] ,
    \Tile_X9Y7_EE4BEG[13] ,
    \Tile_X9Y7_EE4BEG[12] ,
    \Tile_X9Y7_EE4BEG[11] ,
    \Tile_X9Y7_EE4BEG[10] ,
    \Tile_X9Y7_EE4BEG[9] ,
    \Tile_X9Y7_EE4BEG[8] ,
    \Tile_X9Y7_EE4BEG[7] ,
    \Tile_X9Y7_EE4BEG[6] ,
    \Tile_X9Y7_EE4BEG[5] ,
    \Tile_X9Y7_EE4BEG[4] ,
    \Tile_X9Y7_EE4BEG[3] ,
    \Tile_X9Y7_EE4BEG[2] ,
    \Tile_X9Y7_EE4BEG[1] ,
    \Tile_X9Y7_EE4BEG[0] }),
    .EE4END({\Tile_X8Y7_EE4BEG[15] ,
    \Tile_X8Y7_EE4BEG[14] ,
    \Tile_X8Y7_EE4BEG[13] ,
    \Tile_X8Y7_EE4BEG[12] ,
    \Tile_X8Y7_EE4BEG[11] ,
    \Tile_X8Y7_EE4BEG[10] ,
    \Tile_X8Y7_EE4BEG[9] ,
    \Tile_X8Y7_EE4BEG[8] ,
    \Tile_X8Y7_EE4BEG[7] ,
    \Tile_X8Y7_EE4BEG[6] ,
    \Tile_X8Y7_EE4BEG[5] ,
    \Tile_X8Y7_EE4BEG[4] ,
    \Tile_X8Y7_EE4BEG[3] ,
    \Tile_X8Y7_EE4BEG[2] ,
    \Tile_X8Y7_EE4BEG[1] ,
    \Tile_X8Y7_EE4BEG[0] }),
    .FrameData({\Tile_X8Y7_FrameData_O[31] ,
    \Tile_X8Y7_FrameData_O[30] ,
    \Tile_X8Y7_FrameData_O[29] ,
    \Tile_X8Y7_FrameData_O[28] ,
    \Tile_X8Y7_FrameData_O[27] ,
    \Tile_X8Y7_FrameData_O[26] ,
    \Tile_X8Y7_FrameData_O[25] ,
    \Tile_X8Y7_FrameData_O[24] ,
    \Tile_X8Y7_FrameData_O[23] ,
    \Tile_X8Y7_FrameData_O[22] ,
    \Tile_X8Y7_FrameData_O[21] ,
    \Tile_X8Y7_FrameData_O[20] ,
    \Tile_X8Y7_FrameData_O[19] ,
    \Tile_X8Y7_FrameData_O[18] ,
    \Tile_X8Y7_FrameData_O[17] ,
    \Tile_X8Y7_FrameData_O[16] ,
    \Tile_X8Y7_FrameData_O[15] ,
    \Tile_X8Y7_FrameData_O[14] ,
    \Tile_X8Y7_FrameData_O[13] ,
    \Tile_X8Y7_FrameData_O[12] ,
    \Tile_X8Y7_FrameData_O[11] ,
    \Tile_X8Y7_FrameData_O[10] ,
    \Tile_X8Y7_FrameData_O[9] ,
    \Tile_X8Y7_FrameData_O[8] ,
    \Tile_X8Y7_FrameData_O[7] ,
    \Tile_X8Y7_FrameData_O[6] ,
    \Tile_X8Y7_FrameData_O[5] ,
    \Tile_X8Y7_FrameData_O[4] ,
    \Tile_X8Y7_FrameData_O[3] ,
    \Tile_X8Y7_FrameData_O[2] ,
    \Tile_X8Y7_FrameData_O[1] ,
    \Tile_X8Y7_FrameData_O[0] }),
    .FrameData_O({\Tile_X9Y7_FrameData_O[31] ,
    \Tile_X9Y7_FrameData_O[30] ,
    \Tile_X9Y7_FrameData_O[29] ,
    \Tile_X9Y7_FrameData_O[28] ,
    \Tile_X9Y7_FrameData_O[27] ,
    \Tile_X9Y7_FrameData_O[26] ,
    \Tile_X9Y7_FrameData_O[25] ,
    \Tile_X9Y7_FrameData_O[24] ,
    \Tile_X9Y7_FrameData_O[23] ,
    \Tile_X9Y7_FrameData_O[22] ,
    \Tile_X9Y7_FrameData_O[21] ,
    \Tile_X9Y7_FrameData_O[20] ,
    \Tile_X9Y7_FrameData_O[19] ,
    \Tile_X9Y7_FrameData_O[18] ,
    \Tile_X9Y7_FrameData_O[17] ,
    \Tile_X9Y7_FrameData_O[16] ,
    \Tile_X9Y7_FrameData_O[15] ,
    \Tile_X9Y7_FrameData_O[14] ,
    \Tile_X9Y7_FrameData_O[13] ,
    \Tile_X9Y7_FrameData_O[12] ,
    \Tile_X9Y7_FrameData_O[11] ,
    \Tile_X9Y7_FrameData_O[10] ,
    \Tile_X9Y7_FrameData_O[9] ,
    \Tile_X9Y7_FrameData_O[8] ,
    \Tile_X9Y7_FrameData_O[7] ,
    \Tile_X9Y7_FrameData_O[6] ,
    \Tile_X9Y7_FrameData_O[5] ,
    \Tile_X9Y7_FrameData_O[4] ,
    \Tile_X9Y7_FrameData_O[3] ,
    \Tile_X9Y7_FrameData_O[2] ,
    \Tile_X9Y7_FrameData_O[1] ,
    \Tile_X9Y7_FrameData_O[0] }),
    .FrameStrobe({\Tile_X9Y8_FrameStrobe_O[19] ,
    \Tile_X9Y8_FrameStrobe_O[18] ,
    \Tile_X9Y8_FrameStrobe_O[17] ,
    \Tile_X9Y8_FrameStrobe_O[16] ,
    \Tile_X9Y8_FrameStrobe_O[15] ,
    \Tile_X9Y8_FrameStrobe_O[14] ,
    \Tile_X9Y8_FrameStrobe_O[13] ,
    \Tile_X9Y8_FrameStrobe_O[12] ,
    \Tile_X9Y8_FrameStrobe_O[11] ,
    \Tile_X9Y8_FrameStrobe_O[10] ,
    \Tile_X9Y8_FrameStrobe_O[9] ,
    \Tile_X9Y8_FrameStrobe_O[8] ,
    \Tile_X9Y8_FrameStrobe_O[7] ,
    \Tile_X9Y8_FrameStrobe_O[6] ,
    \Tile_X9Y8_FrameStrobe_O[5] ,
    \Tile_X9Y8_FrameStrobe_O[4] ,
    \Tile_X9Y8_FrameStrobe_O[3] ,
    \Tile_X9Y8_FrameStrobe_O[2] ,
    \Tile_X9Y8_FrameStrobe_O[1] ,
    \Tile_X9Y8_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X9Y7_FrameStrobe_O[19] ,
    \Tile_X9Y7_FrameStrobe_O[18] ,
    \Tile_X9Y7_FrameStrobe_O[17] ,
    \Tile_X9Y7_FrameStrobe_O[16] ,
    \Tile_X9Y7_FrameStrobe_O[15] ,
    \Tile_X9Y7_FrameStrobe_O[14] ,
    \Tile_X9Y7_FrameStrobe_O[13] ,
    \Tile_X9Y7_FrameStrobe_O[12] ,
    \Tile_X9Y7_FrameStrobe_O[11] ,
    \Tile_X9Y7_FrameStrobe_O[10] ,
    \Tile_X9Y7_FrameStrobe_O[9] ,
    \Tile_X9Y7_FrameStrobe_O[8] ,
    \Tile_X9Y7_FrameStrobe_O[7] ,
    \Tile_X9Y7_FrameStrobe_O[6] ,
    \Tile_X9Y7_FrameStrobe_O[5] ,
    \Tile_X9Y7_FrameStrobe_O[4] ,
    \Tile_X9Y7_FrameStrobe_O[3] ,
    \Tile_X9Y7_FrameStrobe_O[2] ,
    \Tile_X9Y7_FrameStrobe_O[1] ,
    \Tile_X9Y7_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X9Y7_N1BEG[3] ,
    \Tile_X9Y7_N1BEG[2] ,
    \Tile_X9Y7_N1BEG[1] ,
    \Tile_X9Y7_N1BEG[0] }),
    .N1END({\Tile_X9Y8_N1BEG[3] ,
    \Tile_X9Y8_N1BEG[2] ,
    \Tile_X9Y8_N1BEG[1] ,
    \Tile_X9Y8_N1BEG[0] }),
    .N2BEG({\Tile_X9Y7_N2BEG[7] ,
    \Tile_X9Y7_N2BEG[6] ,
    \Tile_X9Y7_N2BEG[5] ,
    \Tile_X9Y7_N2BEG[4] ,
    \Tile_X9Y7_N2BEG[3] ,
    \Tile_X9Y7_N2BEG[2] ,
    \Tile_X9Y7_N2BEG[1] ,
    \Tile_X9Y7_N2BEG[0] }),
    .N2BEGb({\Tile_X9Y7_N2BEGb[7] ,
    \Tile_X9Y7_N2BEGb[6] ,
    \Tile_X9Y7_N2BEGb[5] ,
    \Tile_X9Y7_N2BEGb[4] ,
    \Tile_X9Y7_N2BEGb[3] ,
    \Tile_X9Y7_N2BEGb[2] ,
    \Tile_X9Y7_N2BEGb[1] ,
    \Tile_X9Y7_N2BEGb[0] }),
    .N2END({\Tile_X9Y8_N2BEGb[7] ,
    \Tile_X9Y8_N2BEGb[6] ,
    \Tile_X9Y8_N2BEGb[5] ,
    \Tile_X9Y8_N2BEGb[4] ,
    \Tile_X9Y8_N2BEGb[3] ,
    \Tile_X9Y8_N2BEGb[2] ,
    \Tile_X9Y8_N2BEGb[1] ,
    \Tile_X9Y8_N2BEGb[0] }),
    .N2MID({\Tile_X9Y8_N2BEG[7] ,
    \Tile_X9Y8_N2BEG[6] ,
    \Tile_X9Y8_N2BEG[5] ,
    \Tile_X9Y8_N2BEG[4] ,
    \Tile_X9Y8_N2BEG[3] ,
    \Tile_X9Y8_N2BEG[2] ,
    \Tile_X9Y8_N2BEG[1] ,
    \Tile_X9Y8_N2BEG[0] }),
    .N4BEG({\Tile_X9Y7_N4BEG[15] ,
    \Tile_X9Y7_N4BEG[14] ,
    \Tile_X9Y7_N4BEG[13] ,
    \Tile_X9Y7_N4BEG[12] ,
    \Tile_X9Y7_N4BEG[11] ,
    \Tile_X9Y7_N4BEG[10] ,
    \Tile_X9Y7_N4BEG[9] ,
    \Tile_X9Y7_N4BEG[8] ,
    \Tile_X9Y7_N4BEG[7] ,
    \Tile_X9Y7_N4BEG[6] ,
    \Tile_X9Y7_N4BEG[5] ,
    \Tile_X9Y7_N4BEG[4] ,
    \Tile_X9Y7_N4BEG[3] ,
    \Tile_X9Y7_N4BEG[2] ,
    \Tile_X9Y7_N4BEG[1] ,
    \Tile_X9Y7_N4BEG[0] }),
    .N4END({\Tile_X9Y8_N4BEG[15] ,
    \Tile_X9Y8_N4BEG[14] ,
    \Tile_X9Y8_N4BEG[13] ,
    \Tile_X9Y8_N4BEG[12] ,
    \Tile_X9Y8_N4BEG[11] ,
    \Tile_X9Y8_N4BEG[10] ,
    \Tile_X9Y8_N4BEG[9] ,
    \Tile_X9Y8_N4BEG[8] ,
    \Tile_X9Y8_N4BEG[7] ,
    \Tile_X9Y8_N4BEG[6] ,
    \Tile_X9Y8_N4BEG[5] ,
    \Tile_X9Y8_N4BEG[4] ,
    \Tile_X9Y8_N4BEG[3] ,
    \Tile_X9Y8_N4BEG[2] ,
    \Tile_X9Y8_N4BEG[1] ,
    \Tile_X9Y8_N4BEG[0] }),
    .NN4BEG({\Tile_X9Y7_NN4BEG[15] ,
    \Tile_X9Y7_NN4BEG[14] ,
    \Tile_X9Y7_NN4BEG[13] ,
    \Tile_X9Y7_NN4BEG[12] ,
    \Tile_X9Y7_NN4BEG[11] ,
    \Tile_X9Y7_NN4BEG[10] ,
    \Tile_X9Y7_NN4BEG[9] ,
    \Tile_X9Y7_NN4BEG[8] ,
    \Tile_X9Y7_NN4BEG[7] ,
    \Tile_X9Y7_NN4BEG[6] ,
    \Tile_X9Y7_NN4BEG[5] ,
    \Tile_X9Y7_NN4BEG[4] ,
    \Tile_X9Y7_NN4BEG[3] ,
    \Tile_X9Y7_NN4BEG[2] ,
    \Tile_X9Y7_NN4BEG[1] ,
    \Tile_X9Y7_NN4BEG[0] }),
    .NN4END({\Tile_X9Y8_NN4BEG[15] ,
    \Tile_X9Y8_NN4BEG[14] ,
    \Tile_X9Y8_NN4BEG[13] ,
    \Tile_X9Y8_NN4BEG[12] ,
    \Tile_X9Y8_NN4BEG[11] ,
    \Tile_X9Y8_NN4BEG[10] ,
    \Tile_X9Y8_NN4BEG[9] ,
    \Tile_X9Y8_NN4BEG[8] ,
    \Tile_X9Y8_NN4BEG[7] ,
    \Tile_X9Y8_NN4BEG[6] ,
    \Tile_X9Y8_NN4BEG[5] ,
    \Tile_X9Y8_NN4BEG[4] ,
    \Tile_X9Y8_NN4BEG[3] ,
    \Tile_X9Y8_NN4BEG[2] ,
    \Tile_X9Y8_NN4BEG[1] ,
    \Tile_X9Y8_NN4BEG[0] }),
    .S1BEG({\Tile_X9Y7_S1BEG[3] ,
    \Tile_X9Y7_S1BEG[2] ,
    \Tile_X9Y7_S1BEG[1] ,
    \Tile_X9Y7_S1BEG[0] }),
    .S1END({\Tile_X9Y6_S1BEG[3] ,
    \Tile_X9Y6_S1BEG[2] ,
    \Tile_X9Y6_S1BEG[1] ,
    \Tile_X9Y6_S1BEG[0] }),
    .S2BEG({\Tile_X9Y7_S2BEG[7] ,
    \Tile_X9Y7_S2BEG[6] ,
    \Tile_X9Y7_S2BEG[5] ,
    \Tile_X9Y7_S2BEG[4] ,
    \Tile_X9Y7_S2BEG[3] ,
    \Tile_X9Y7_S2BEG[2] ,
    \Tile_X9Y7_S2BEG[1] ,
    \Tile_X9Y7_S2BEG[0] }),
    .S2BEGb({\Tile_X9Y7_S2BEGb[7] ,
    \Tile_X9Y7_S2BEGb[6] ,
    \Tile_X9Y7_S2BEGb[5] ,
    \Tile_X9Y7_S2BEGb[4] ,
    \Tile_X9Y7_S2BEGb[3] ,
    \Tile_X9Y7_S2BEGb[2] ,
    \Tile_X9Y7_S2BEGb[1] ,
    \Tile_X9Y7_S2BEGb[0] }),
    .S2END({\Tile_X9Y6_S2BEGb[7] ,
    \Tile_X9Y6_S2BEGb[6] ,
    \Tile_X9Y6_S2BEGb[5] ,
    \Tile_X9Y6_S2BEGb[4] ,
    \Tile_X9Y6_S2BEGb[3] ,
    \Tile_X9Y6_S2BEGb[2] ,
    \Tile_X9Y6_S2BEGb[1] ,
    \Tile_X9Y6_S2BEGb[0] }),
    .S2MID({\Tile_X9Y6_S2BEG[7] ,
    \Tile_X9Y6_S2BEG[6] ,
    \Tile_X9Y6_S2BEG[5] ,
    \Tile_X9Y6_S2BEG[4] ,
    \Tile_X9Y6_S2BEG[3] ,
    \Tile_X9Y6_S2BEG[2] ,
    \Tile_X9Y6_S2BEG[1] ,
    \Tile_X9Y6_S2BEG[0] }),
    .S4BEG({\Tile_X9Y7_S4BEG[15] ,
    \Tile_X9Y7_S4BEG[14] ,
    \Tile_X9Y7_S4BEG[13] ,
    \Tile_X9Y7_S4BEG[12] ,
    \Tile_X9Y7_S4BEG[11] ,
    \Tile_X9Y7_S4BEG[10] ,
    \Tile_X9Y7_S4BEG[9] ,
    \Tile_X9Y7_S4BEG[8] ,
    \Tile_X9Y7_S4BEG[7] ,
    \Tile_X9Y7_S4BEG[6] ,
    \Tile_X9Y7_S4BEG[5] ,
    \Tile_X9Y7_S4BEG[4] ,
    \Tile_X9Y7_S4BEG[3] ,
    \Tile_X9Y7_S4BEG[2] ,
    \Tile_X9Y7_S4BEG[1] ,
    \Tile_X9Y7_S4BEG[0] }),
    .S4END({\Tile_X9Y6_S4BEG[15] ,
    \Tile_X9Y6_S4BEG[14] ,
    \Tile_X9Y6_S4BEG[13] ,
    \Tile_X9Y6_S4BEG[12] ,
    \Tile_X9Y6_S4BEG[11] ,
    \Tile_X9Y6_S4BEG[10] ,
    \Tile_X9Y6_S4BEG[9] ,
    \Tile_X9Y6_S4BEG[8] ,
    \Tile_X9Y6_S4BEG[7] ,
    \Tile_X9Y6_S4BEG[6] ,
    \Tile_X9Y6_S4BEG[5] ,
    \Tile_X9Y6_S4BEG[4] ,
    \Tile_X9Y6_S4BEG[3] ,
    \Tile_X9Y6_S4BEG[2] ,
    \Tile_X9Y6_S4BEG[1] ,
    \Tile_X9Y6_S4BEG[0] }),
    .SS4BEG({\Tile_X9Y7_SS4BEG[15] ,
    \Tile_X9Y7_SS4BEG[14] ,
    \Tile_X9Y7_SS4BEG[13] ,
    \Tile_X9Y7_SS4BEG[12] ,
    \Tile_X9Y7_SS4BEG[11] ,
    \Tile_X9Y7_SS4BEG[10] ,
    \Tile_X9Y7_SS4BEG[9] ,
    \Tile_X9Y7_SS4BEG[8] ,
    \Tile_X9Y7_SS4BEG[7] ,
    \Tile_X9Y7_SS4BEG[6] ,
    \Tile_X9Y7_SS4BEG[5] ,
    \Tile_X9Y7_SS4BEG[4] ,
    \Tile_X9Y7_SS4BEG[3] ,
    \Tile_X9Y7_SS4BEG[2] ,
    \Tile_X9Y7_SS4BEG[1] ,
    \Tile_X9Y7_SS4BEG[0] }),
    .SS4END({\Tile_X9Y6_SS4BEG[15] ,
    \Tile_X9Y6_SS4BEG[14] ,
    \Tile_X9Y6_SS4BEG[13] ,
    \Tile_X9Y6_SS4BEG[12] ,
    \Tile_X9Y6_SS4BEG[11] ,
    \Tile_X9Y6_SS4BEG[10] ,
    \Tile_X9Y6_SS4BEG[9] ,
    \Tile_X9Y6_SS4BEG[8] ,
    \Tile_X9Y6_SS4BEG[7] ,
    \Tile_X9Y6_SS4BEG[6] ,
    \Tile_X9Y6_SS4BEG[5] ,
    \Tile_X9Y6_SS4BEG[4] ,
    \Tile_X9Y6_SS4BEG[3] ,
    \Tile_X9Y6_SS4BEG[2] ,
    \Tile_X9Y6_SS4BEG[1] ,
    \Tile_X9Y6_SS4BEG[0] }),
    .W1BEG({\Tile_X9Y7_W1BEG[3] ,
    \Tile_X9Y7_W1BEG[2] ,
    \Tile_X9Y7_W1BEG[1] ,
    \Tile_X9Y7_W1BEG[0] }),
    .W1END({\Tile_X10Y7_W1BEG[3] ,
    \Tile_X10Y7_W1BEG[2] ,
    \Tile_X10Y7_W1BEG[1] ,
    \Tile_X10Y7_W1BEG[0] }),
    .W2BEG({\Tile_X9Y7_W2BEG[7] ,
    \Tile_X9Y7_W2BEG[6] ,
    \Tile_X9Y7_W2BEG[5] ,
    \Tile_X9Y7_W2BEG[4] ,
    \Tile_X9Y7_W2BEG[3] ,
    \Tile_X9Y7_W2BEG[2] ,
    \Tile_X9Y7_W2BEG[1] ,
    \Tile_X9Y7_W2BEG[0] }),
    .W2BEGb({\Tile_X9Y7_W2BEGb[7] ,
    \Tile_X9Y7_W2BEGb[6] ,
    \Tile_X9Y7_W2BEGb[5] ,
    \Tile_X9Y7_W2BEGb[4] ,
    \Tile_X9Y7_W2BEGb[3] ,
    \Tile_X9Y7_W2BEGb[2] ,
    \Tile_X9Y7_W2BEGb[1] ,
    \Tile_X9Y7_W2BEGb[0] }),
    .W2END({\Tile_X10Y7_W2BEGb[7] ,
    \Tile_X10Y7_W2BEGb[6] ,
    \Tile_X10Y7_W2BEGb[5] ,
    \Tile_X10Y7_W2BEGb[4] ,
    \Tile_X10Y7_W2BEGb[3] ,
    \Tile_X10Y7_W2BEGb[2] ,
    \Tile_X10Y7_W2BEGb[1] ,
    \Tile_X10Y7_W2BEGb[0] }),
    .W2MID({\Tile_X10Y7_W2BEG[7] ,
    \Tile_X10Y7_W2BEG[6] ,
    \Tile_X10Y7_W2BEG[5] ,
    \Tile_X10Y7_W2BEG[4] ,
    \Tile_X10Y7_W2BEG[3] ,
    \Tile_X10Y7_W2BEG[2] ,
    \Tile_X10Y7_W2BEG[1] ,
    \Tile_X10Y7_W2BEG[0] }),
    .W6BEG({\Tile_X9Y7_W6BEG[11] ,
    \Tile_X9Y7_W6BEG[10] ,
    \Tile_X9Y7_W6BEG[9] ,
    \Tile_X9Y7_W6BEG[8] ,
    \Tile_X9Y7_W6BEG[7] ,
    \Tile_X9Y7_W6BEG[6] ,
    \Tile_X9Y7_W6BEG[5] ,
    \Tile_X9Y7_W6BEG[4] ,
    \Tile_X9Y7_W6BEG[3] ,
    \Tile_X9Y7_W6BEG[2] ,
    \Tile_X9Y7_W6BEG[1] ,
    \Tile_X9Y7_W6BEG[0] }),
    .W6END({\Tile_X10Y7_W6BEG[11] ,
    \Tile_X10Y7_W6BEG[10] ,
    \Tile_X10Y7_W6BEG[9] ,
    \Tile_X10Y7_W6BEG[8] ,
    \Tile_X10Y7_W6BEG[7] ,
    \Tile_X10Y7_W6BEG[6] ,
    \Tile_X10Y7_W6BEG[5] ,
    \Tile_X10Y7_W6BEG[4] ,
    \Tile_X10Y7_W6BEG[3] ,
    \Tile_X10Y7_W6BEG[2] ,
    \Tile_X10Y7_W6BEG[1] ,
    \Tile_X10Y7_W6BEG[0] }),
    .WW4BEG({\Tile_X9Y7_WW4BEG[15] ,
    \Tile_X9Y7_WW4BEG[14] ,
    \Tile_X9Y7_WW4BEG[13] ,
    \Tile_X9Y7_WW4BEG[12] ,
    \Tile_X9Y7_WW4BEG[11] ,
    \Tile_X9Y7_WW4BEG[10] ,
    \Tile_X9Y7_WW4BEG[9] ,
    \Tile_X9Y7_WW4BEG[8] ,
    \Tile_X9Y7_WW4BEG[7] ,
    \Tile_X9Y7_WW4BEG[6] ,
    \Tile_X9Y7_WW4BEG[5] ,
    \Tile_X9Y7_WW4BEG[4] ,
    \Tile_X9Y7_WW4BEG[3] ,
    \Tile_X9Y7_WW4BEG[2] ,
    \Tile_X9Y7_WW4BEG[1] ,
    \Tile_X9Y7_WW4BEG[0] }),
    .WW4END({\Tile_X10Y7_WW4BEG[15] ,
    \Tile_X10Y7_WW4BEG[14] ,
    \Tile_X10Y7_WW4BEG[13] ,
    \Tile_X10Y7_WW4BEG[12] ,
    \Tile_X10Y7_WW4BEG[11] ,
    \Tile_X10Y7_WW4BEG[10] ,
    \Tile_X10Y7_WW4BEG[9] ,
    \Tile_X10Y7_WW4BEG[8] ,
    \Tile_X10Y7_WW4BEG[7] ,
    \Tile_X10Y7_WW4BEG[6] ,
    \Tile_X10Y7_WW4BEG[5] ,
    \Tile_X10Y7_WW4BEG[4] ,
    \Tile_X10Y7_WW4BEG[3] ,
    \Tile_X10Y7_WW4BEG[2] ,
    \Tile_X10Y7_WW4BEG[1] ,
    \Tile_X10Y7_WW4BEG[0] }));
 LUT4AB Tile_X9Y8_LUT4AB (.Ci(Tile_X9Y9_Co),
    .Co(Tile_X9Y8_Co),
    .UserCLK(Tile_X9Y9_UserCLKo),
    .UserCLKo(Tile_X9Y8_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X9Y8_E1BEG[3] ,
    \Tile_X9Y8_E1BEG[2] ,
    \Tile_X9Y8_E1BEG[1] ,
    \Tile_X9Y8_E1BEG[0] }),
    .E1END({\Tile_X8Y8_E1BEG[3] ,
    \Tile_X8Y8_E1BEG[2] ,
    \Tile_X8Y8_E1BEG[1] ,
    \Tile_X8Y8_E1BEG[0] }),
    .E2BEG({\Tile_X9Y8_E2BEG[7] ,
    \Tile_X9Y8_E2BEG[6] ,
    \Tile_X9Y8_E2BEG[5] ,
    \Tile_X9Y8_E2BEG[4] ,
    \Tile_X9Y8_E2BEG[3] ,
    \Tile_X9Y8_E2BEG[2] ,
    \Tile_X9Y8_E2BEG[1] ,
    \Tile_X9Y8_E2BEG[0] }),
    .E2BEGb({\Tile_X9Y8_E2BEGb[7] ,
    \Tile_X9Y8_E2BEGb[6] ,
    \Tile_X9Y8_E2BEGb[5] ,
    \Tile_X9Y8_E2BEGb[4] ,
    \Tile_X9Y8_E2BEGb[3] ,
    \Tile_X9Y8_E2BEGb[2] ,
    \Tile_X9Y8_E2BEGb[1] ,
    \Tile_X9Y8_E2BEGb[0] }),
    .E2END({\Tile_X8Y8_E2BEGb[7] ,
    \Tile_X8Y8_E2BEGb[6] ,
    \Tile_X8Y8_E2BEGb[5] ,
    \Tile_X8Y8_E2BEGb[4] ,
    \Tile_X8Y8_E2BEGb[3] ,
    \Tile_X8Y8_E2BEGb[2] ,
    \Tile_X8Y8_E2BEGb[1] ,
    \Tile_X8Y8_E2BEGb[0] }),
    .E2MID({\Tile_X8Y8_E2BEG[7] ,
    \Tile_X8Y8_E2BEG[6] ,
    \Tile_X8Y8_E2BEG[5] ,
    \Tile_X8Y8_E2BEG[4] ,
    \Tile_X8Y8_E2BEG[3] ,
    \Tile_X8Y8_E2BEG[2] ,
    \Tile_X8Y8_E2BEG[1] ,
    \Tile_X8Y8_E2BEG[0] }),
    .E6BEG({\Tile_X9Y8_E6BEG[11] ,
    \Tile_X9Y8_E6BEG[10] ,
    \Tile_X9Y8_E6BEG[9] ,
    \Tile_X9Y8_E6BEG[8] ,
    \Tile_X9Y8_E6BEG[7] ,
    \Tile_X9Y8_E6BEG[6] ,
    \Tile_X9Y8_E6BEG[5] ,
    \Tile_X9Y8_E6BEG[4] ,
    \Tile_X9Y8_E6BEG[3] ,
    \Tile_X9Y8_E6BEG[2] ,
    \Tile_X9Y8_E6BEG[1] ,
    \Tile_X9Y8_E6BEG[0] }),
    .E6END({\Tile_X8Y8_E6BEG[11] ,
    \Tile_X8Y8_E6BEG[10] ,
    \Tile_X8Y8_E6BEG[9] ,
    \Tile_X8Y8_E6BEG[8] ,
    \Tile_X8Y8_E6BEG[7] ,
    \Tile_X8Y8_E6BEG[6] ,
    \Tile_X8Y8_E6BEG[5] ,
    \Tile_X8Y8_E6BEG[4] ,
    \Tile_X8Y8_E6BEG[3] ,
    \Tile_X8Y8_E6BEG[2] ,
    \Tile_X8Y8_E6BEG[1] ,
    \Tile_X8Y8_E6BEG[0] }),
    .EE4BEG({\Tile_X9Y8_EE4BEG[15] ,
    \Tile_X9Y8_EE4BEG[14] ,
    \Tile_X9Y8_EE4BEG[13] ,
    \Tile_X9Y8_EE4BEG[12] ,
    \Tile_X9Y8_EE4BEG[11] ,
    \Tile_X9Y8_EE4BEG[10] ,
    \Tile_X9Y8_EE4BEG[9] ,
    \Tile_X9Y8_EE4BEG[8] ,
    \Tile_X9Y8_EE4BEG[7] ,
    \Tile_X9Y8_EE4BEG[6] ,
    \Tile_X9Y8_EE4BEG[5] ,
    \Tile_X9Y8_EE4BEG[4] ,
    \Tile_X9Y8_EE4BEG[3] ,
    \Tile_X9Y8_EE4BEG[2] ,
    \Tile_X9Y8_EE4BEG[1] ,
    \Tile_X9Y8_EE4BEG[0] }),
    .EE4END({\Tile_X8Y8_EE4BEG[15] ,
    \Tile_X8Y8_EE4BEG[14] ,
    \Tile_X8Y8_EE4BEG[13] ,
    \Tile_X8Y8_EE4BEG[12] ,
    \Tile_X8Y8_EE4BEG[11] ,
    \Tile_X8Y8_EE4BEG[10] ,
    \Tile_X8Y8_EE4BEG[9] ,
    \Tile_X8Y8_EE4BEG[8] ,
    \Tile_X8Y8_EE4BEG[7] ,
    \Tile_X8Y8_EE4BEG[6] ,
    \Tile_X8Y8_EE4BEG[5] ,
    \Tile_X8Y8_EE4BEG[4] ,
    \Tile_X8Y8_EE4BEG[3] ,
    \Tile_X8Y8_EE4BEG[2] ,
    \Tile_X8Y8_EE4BEG[1] ,
    \Tile_X8Y8_EE4BEG[0] }),
    .FrameData({\Tile_X8Y8_FrameData_O[31] ,
    \Tile_X8Y8_FrameData_O[30] ,
    \Tile_X8Y8_FrameData_O[29] ,
    \Tile_X8Y8_FrameData_O[28] ,
    \Tile_X8Y8_FrameData_O[27] ,
    \Tile_X8Y8_FrameData_O[26] ,
    \Tile_X8Y8_FrameData_O[25] ,
    \Tile_X8Y8_FrameData_O[24] ,
    \Tile_X8Y8_FrameData_O[23] ,
    \Tile_X8Y8_FrameData_O[22] ,
    \Tile_X8Y8_FrameData_O[21] ,
    \Tile_X8Y8_FrameData_O[20] ,
    \Tile_X8Y8_FrameData_O[19] ,
    \Tile_X8Y8_FrameData_O[18] ,
    \Tile_X8Y8_FrameData_O[17] ,
    \Tile_X8Y8_FrameData_O[16] ,
    \Tile_X8Y8_FrameData_O[15] ,
    \Tile_X8Y8_FrameData_O[14] ,
    \Tile_X8Y8_FrameData_O[13] ,
    \Tile_X8Y8_FrameData_O[12] ,
    \Tile_X8Y8_FrameData_O[11] ,
    \Tile_X8Y8_FrameData_O[10] ,
    \Tile_X8Y8_FrameData_O[9] ,
    \Tile_X8Y8_FrameData_O[8] ,
    \Tile_X8Y8_FrameData_O[7] ,
    \Tile_X8Y8_FrameData_O[6] ,
    \Tile_X8Y8_FrameData_O[5] ,
    \Tile_X8Y8_FrameData_O[4] ,
    \Tile_X8Y8_FrameData_O[3] ,
    \Tile_X8Y8_FrameData_O[2] ,
    \Tile_X8Y8_FrameData_O[1] ,
    \Tile_X8Y8_FrameData_O[0] }),
    .FrameData_O({\Tile_X9Y8_FrameData_O[31] ,
    \Tile_X9Y8_FrameData_O[30] ,
    \Tile_X9Y8_FrameData_O[29] ,
    \Tile_X9Y8_FrameData_O[28] ,
    \Tile_X9Y8_FrameData_O[27] ,
    \Tile_X9Y8_FrameData_O[26] ,
    \Tile_X9Y8_FrameData_O[25] ,
    \Tile_X9Y8_FrameData_O[24] ,
    \Tile_X9Y8_FrameData_O[23] ,
    \Tile_X9Y8_FrameData_O[22] ,
    \Tile_X9Y8_FrameData_O[21] ,
    \Tile_X9Y8_FrameData_O[20] ,
    \Tile_X9Y8_FrameData_O[19] ,
    \Tile_X9Y8_FrameData_O[18] ,
    \Tile_X9Y8_FrameData_O[17] ,
    \Tile_X9Y8_FrameData_O[16] ,
    \Tile_X9Y8_FrameData_O[15] ,
    \Tile_X9Y8_FrameData_O[14] ,
    \Tile_X9Y8_FrameData_O[13] ,
    \Tile_X9Y8_FrameData_O[12] ,
    \Tile_X9Y8_FrameData_O[11] ,
    \Tile_X9Y8_FrameData_O[10] ,
    \Tile_X9Y8_FrameData_O[9] ,
    \Tile_X9Y8_FrameData_O[8] ,
    \Tile_X9Y8_FrameData_O[7] ,
    \Tile_X9Y8_FrameData_O[6] ,
    \Tile_X9Y8_FrameData_O[5] ,
    \Tile_X9Y8_FrameData_O[4] ,
    \Tile_X9Y8_FrameData_O[3] ,
    \Tile_X9Y8_FrameData_O[2] ,
    \Tile_X9Y8_FrameData_O[1] ,
    \Tile_X9Y8_FrameData_O[0] }),
    .FrameStrobe({\Tile_X9Y9_FrameStrobe_O[19] ,
    \Tile_X9Y9_FrameStrobe_O[18] ,
    \Tile_X9Y9_FrameStrobe_O[17] ,
    \Tile_X9Y9_FrameStrobe_O[16] ,
    \Tile_X9Y9_FrameStrobe_O[15] ,
    \Tile_X9Y9_FrameStrobe_O[14] ,
    \Tile_X9Y9_FrameStrobe_O[13] ,
    \Tile_X9Y9_FrameStrobe_O[12] ,
    \Tile_X9Y9_FrameStrobe_O[11] ,
    \Tile_X9Y9_FrameStrobe_O[10] ,
    \Tile_X9Y9_FrameStrobe_O[9] ,
    \Tile_X9Y9_FrameStrobe_O[8] ,
    \Tile_X9Y9_FrameStrobe_O[7] ,
    \Tile_X9Y9_FrameStrobe_O[6] ,
    \Tile_X9Y9_FrameStrobe_O[5] ,
    \Tile_X9Y9_FrameStrobe_O[4] ,
    \Tile_X9Y9_FrameStrobe_O[3] ,
    \Tile_X9Y9_FrameStrobe_O[2] ,
    \Tile_X9Y9_FrameStrobe_O[1] ,
    \Tile_X9Y9_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X9Y8_FrameStrobe_O[19] ,
    \Tile_X9Y8_FrameStrobe_O[18] ,
    \Tile_X9Y8_FrameStrobe_O[17] ,
    \Tile_X9Y8_FrameStrobe_O[16] ,
    \Tile_X9Y8_FrameStrobe_O[15] ,
    \Tile_X9Y8_FrameStrobe_O[14] ,
    \Tile_X9Y8_FrameStrobe_O[13] ,
    \Tile_X9Y8_FrameStrobe_O[12] ,
    \Tile_X9Y8_FrameStrobe_O[11] ,
    \Tile_X9Y8_FrameStrobe_O[10] ,
    \Tile_X9Y8_FrameStrobe_O[9] ,
    \Tile_X9Y8_FrameStrobe_O[8] ,
    \Tile_X9Y8_FrameStrobe_O[7] ,
    \Tile_X9Y8_FrameStrobe_O[6] ,
    \Tile_X9Y8_FrameStrobe_O[5] ,
    \Tile_X9Y8_FrameStrobe_O[4] ,
    \Tile_X9Y8_FrameStrobe_O[3] ,
    \Tile_X9Y8_FrameStrobe_O[2] ,
    \Tile_X9Y8_FrameStrobe_O[1] ,
    \Tile_X9Y8_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X9Y8_N1BEG[3] ,
    \Tile_X9Y8_N1BEG[2] ,
    \Tile_X9Y8_N1BEG[1] ,
    \Tile_X9Y8_N1BEG[0] }),
    .N1END({\Tile_X9Y9_N1BEG[3] ,
    \Tile_X9Y9_N1BEG[2] ,
    \Tile_X9Y9_N1BEG[1] ,
    \Tile_X9Y9_N1BEG[0] }),
    .N2BEG({\Tile_X9Y8_N2BEG[7] ,
    \Tile_X9Y8_N2BEG[6] ,
    \Tile_X9Y8_N2BEG[5] ,
    \Tile_X9Y8_N2BEG[4] ,
    \Tile_X9Y8_N2BEG[3] ,
    \Tile_X9Y8_N2BEG[2] ,
    \Tile_X9Y8_N2BEG[1] ,
    \Tile_X9Y8_N2BEG[0] }),
    .N2BEGb({\Tile_X9Y8_N2BEGb[7] ,
    \Tile_X9Y8_N2BEGb[6] ,
    \Tile_X9Y8_N2BEGb[5] ,
    \Tile_X9Y8_N2BEGb[4] ,
    \Tile_X9Y8_N2BEGb[3] ,
    \Tile_X9Y8_N2BEGb[2] ,
    \Tile_X9Y8_N2BEGb[1] ,
    \Tile_X9Y8_N2BEGb[0] }),
    .N2END({\Tile_X9Y9_N2BEGb[7] ,
    \Tile_X9Y9_N2BEGb[6] ,
    \Tile_X9Y9_N2BEGb[5] ,
    \Tile_X9Y9_N2BEGb[4] ,
    \Tile_X9Y9_N2BEGb[3] ,
    \Tile_X9Y9_N2BEGb[2] ,
    \Tile_X9Y9_N2BEGb[1] ,
    \Tile_X9Y9_N2BEGb[0] }),
    .N2MID({\Tile_X9Y9_N2BEG[7] ,
    \Tile_X9Y9_N2BEG[6] ,
    \Tile_X9Y9_N2BEG[5] ,
    \Tile_X9Y9_N2BEG[4] ,
    \Tile_X9Y9_N2BEG[3] ,
    \Tile_X9Y9_N2BEG[2] ,
    \Tile_X9Y9_N2BEG[1] ,
    \Tile_X9Y9_N2BEG[0] }),
    .N4BEG({\Tile_X9Y8_N4BEG[15] ,
    \Tile_X9Y8_N4BEG[14] ,
    \Tile_X9Y8_N4BEG[13] ,
    \Tile_X9Y8_N4BEG[12] ,
    \Tile_X9Y8_N4BEG[11] ,
    \Tile_X9Y8_N4BEG[10] ,
    \Tile_X9Y8_N4BEG[9] ,
    \Tile_X9Y8_N4BEG[8] ,
    \Tile_X9Y8_N4BEG[7] ,
    \Tile_X9Y8_N4BEG[6] ,
    \Tile_X9Y8_N4BEG[5] ,
    \Tile_X9Y8_N4BEG[4] ,
    \Tile_X9Y8_N4BEG[3] ,
    \Tile_X9Y8_N4BEG[2] ,
    \Tile_X9Y8_N4BEG[1] ,
    \Tile_X9Y8_N4BEG[0] }),
    .N4END({\Tile_X9Y9_N4BEG[15] ,
    \Tile_X9Y9_N4BEG[14] ,
    \Tile_X9Y9_N4BEG[13] ,
    \Tile_X9Y9_N4BEG[12] ,
    \Tile_X9Y9_N4BEG[11] ,
    \Tile_X9Y9_N4BEG[10] ,
    \Tile_X9Y9_N4BEG[9] ,
    \Tile_X9Y9_N4BEG[8] ,
    \Tile_X9Y9_N4BEG[7] ,
    \Tile_X9Y9_N4BEG[6] ,
    \Tile_X9Y9_N4BEG[5] ,
    \Tile_X9Y9_N4BEG[4] ,
    \Tile_X9Y9_N4BEG[3] ,
    \Tile_X9Y9_N4BEG[2] ,
    \Tile_X9Y9_N4BEG[1] ,
    \Tile_X9Y9_N4BEG[0] }),
    .NN4BEG({\Tile_X9Y8_NN4BEG[15] ,
    \Tile_X9Y8_NN4BEG[14] ,
    \Tile_X9Y8_NN4BEG[13] ,
    \Tile_X9Y8_NN4BEG[12] ,
    \Tile_X9Y8_NN4BEG[11] ,
    \Tile_X9Y8_NN4BEG[10] ,
    \Tile_X9Y8_NN4BEG[9] ,
    \Tile_X9Y8_NN4BEG[8] ,
    \Tile_X9Y8_NN4BEG[7] ,
    \Tile_X9Y8_NN4BEG[6] ,
    \Tile_X9Y8_NN4BEG[5] ,
    \Tile_X9Y8_NN4BEG[4] ,
    \Tile_X9Y8_NN4BEG[3] ,
    \Tile_X9Y8_NN4BEG[2] ,
    \Tile_X9Y8_NN4BEG[1] ,
    \Tile_X9Y8_NN4BEG[0] }),
    .NN4END({\Tile_X9Y9_NN4BEG[15] ,
    \Tile_X9Y9_NN4BEG[14] ,
    \Tile_X9Y9_NN4BEG[13] ,
    \Tile_X9Y9_NN4BEG[12] ,
    \Tile_X9Y9_NN4BEG[11] ,
    \Tile_X9Y9_NN4BEG[10] ,
    \Tile_X9Y9_NN4BEG[9] ,
    \Tile_X9Y9_NN4BEG[8] ,
    \Tile_X9Y9_NN4BEG[7] ,
    \Tile_X9Y9_NN4BEG[6] ,
    \Tile_X9Y9_NN4BEG[5] ,
    \Tile_X9Y9_NN4BEG[4] ,
    \Tile_X9Y9_NN4BEG[3] ,
    \Tile_X9Y9_NN4BEG[2] ,
    \Tile_X9Y9_NN4BEG[1] ,
    \Tile_X9Y9_NN4BEG[0] }),
    .S1BEG({\Tile_X9Y8_S1BEG[3] ,
    \Tile_X9Y8_S1BEG[2] ,
    \Tile_X9Y8_S1BEG[1] ,
    \Tile_X9Y8_S1BEG[0] }),
    .S1END({\Tile_X9Y7_S1BEG[3] ,
    \Tile_X9Y7_S1BEG[2] ,
    \Tile_X9Y7_S1BEG[1] ,
    \Tile_X9Y7_S1BEG[0] }),
    .S2BEG({\Tile_X9Y8_S2BEG[7] ,
    \Tile_X9Y8_S2BEG[6] ,
    \Tile_X9Y8_S2BEG[5] ,
    \Tile_X9Y8_S2BEG[4] ,
    \Tile_X9Y8_S2BEG[3] ,
    \Tile_X9Y8_S2BEG[2] ,
    \Tile_X9Y8_S2BEG[1] ,
    \Tile_X9Y8_S2BEG[0] }),
    .S2BEGb({\Tile_X9Y8_S2BEGb[7] ,
    \Tile_X9Y8_S2BEGb[6] ,
    \Tile_X9Y8_S2BEGb[5] ,
    \Tile_X9Y8_S2BEGb[4] ,
    \Tile_X9Y8_S2BEGb[3] ,
    \Tile_X9Y8_S2BEGb[2] ,
    \Tile_X9Y8_S2BEGb[1] ,
    \Tile_X9Y8_S2BEGb[0] }),
    .S2END({\Tile_X9Y7_S2BEGb[7] ,
    \Tile_X9Y7_S2BEGb[6] ,
    \Tile_X9Y7_S2BEGb[5] ,
    \Tile_X9Y7_S2BEGb[4] ,
    \Tile_X9Y7_S2BEGb[3] ,
    \Tile_X9Y7_S2BEGb[2] ,
    \Tile_X9Y7_S2BEGb[1] ,
    \Tile_X9Y7_S2BEGb[0] }),
    .S2MID({\Tile_X9Y7_S2BEG[7] ,
    \Tile_X9Y7_S2BEG[6] ,
    \Tile_X9Y7_S2BEG[5] ,
    \Tile_X9Y7_S2BEG[4] ,
    \Tile_X9Y7_S2BEG[3] ,
    \Tile_X9Y7_S2BEG[2] ,
    \Tile_X9Y7_S2BEG[1] ,
    \Tile_X9Y7_S2BEG[0] }),
    .S4BEG({\Tile_X9Y8_S4BEG[15] ,
    \Tile_X9Y8_S4BEG[14] ,
    \Tile_X9Y8_S4BEG[13] ,
    \Tile_X9Y8_S4BEG[12] ,
    \Tile_X9Y8_S4BEG[11] ,
    \Tile_X9Y8_S4BEG[10] ,
    \Tile_X9Y8_S4BEG[9] ,
    \Tile_X9Y8_S4BEG[8] ,
    \Tile_X9Y8_S4BEG[7] ,
    \Tile_X9Y8_S4BEG[6] ,
    \Tile_X9Y8_S4BEG[5] ,
    \Tile_X9Y8_S4BEG[4] ,
    \Tile_X9Y8_S4BEG[3] ,
    \Tile_X9Y8_S4BEG[2] ,
    \Tile_X9Y8_S4BEG[1] ,
    \Tile_X9Y8_S4BEG[0] }),
    .S4END({\Tile_X9Y7_S4BEG[15] ,
    \Tile_X9Y7_S4BEG[14] ,
    \Tile_X9Y7_S4BEG[13] ,
    \Tile_X9Y7_S4BEG[12] ,
    \Tile_X9Y7_S4BEG[11] ,
    \Tile_X9Y7_S4BEG[10] ,
    \Tile_X9Y7_S4BEG[9] ,
    \Tile_X9Y7_S4BEG[8] ,
    \Tile_X9Y7_S4BEG[7] ,
    \Tile_X9Y7_S4BEG[6] ,
    \Tile_X9Y7_S4BEG[5] ,
    \Tile_X9Y7_S4BEG[4] ,
    \Tile_X9Y7_S4BEG[3] ,
    \Tile_X9Y7_S4BEG[2] ,
    \Tile_X9Y7_S4BEG[1] ,
    \Tile_X9Y7_S4BEG[0] }),
    .SS4BEG({\Tile_X9Y8_SS4BEG[15] ,
    \Tile_X9Y8_SS4BEG[14] ,
    \Tile_X9Y8_SS4BEG[13] ,
    \Tile_X9Y8_SS4BEG[12] ,
    \Tile_X9Y8_SS4BEG[11] ,
    \Tile_X9Y8_SS4BEG[10] ,
    \Tile_X9Y8_SS4BEG[9] ,
    \Tile_X9Y8_SS4BEG[8] ,
    \Tile_X9Y8_SS4BEG[7] ,
    \Tile_X9Y8_SS4BEG[6] ,
    \Tile_X9Y8_SS4BEG[5] ,
    \Tile_X9Y8_SS4BEG[4] ,
    \Tile_X9Y8_SS4BEG[3] ,
    \Tile_X9Y8_SS4BEG[2] ,
    \Tile_X9Y8_SS4BEG[1] ,
    \Tile_X9Y8_SS4BEG[0] }),
    .SS4END({\Tile_X9Y7_SS4BEG[15] ,
    \Tile_X9Y7_SS4BEG[14] ,
    \Tile_X9Y7_SS4BEG[13] ,
    \Tile_X9Y7_SS4BEG[12] ,
    \Tile_X9Y7_SS4BEG[11] ,
    \Tile_X9Y7_SS4BEG[10] ,
    \Tile_X9Y7_SS4BEG[9] ,
    \Tile_X9Y7_SS4BEG[8] ,
    \Tile_X9Y7_SS4BEG[7] ,
    \Tile_X9Y7_SS4BEG[6] ,
    \Tile_X9Y7_SS4BEG[5] ,
    \Tile_X9Y7_SS4BEG[4] ,
    \Tile_X9Y7_SS4BEG[3] ,
    \Tile_X9Y7_SS4BEG[2] ,
    \Tile_X9Y7_SS4BEG[1] ,
    \Tile_X9Y7_SS4BEG[0] }),
    .W1BEG({\Tile_X9Y8_W1BEG[3] ,
    \Tile_X9Y8_W1BEG[2] ,
    \Tile_X9Y8_W1BEG[1] ,
    \Tile_X9Y8_W1BEG[0] }),
    .W1END({\Tile_X10Y8_W1BEG[3] ,
    \Tile_X10Y8_W1BEG[2] ,
    \Tile_X10Y8_W1BEG[1] ,
    \Tile_X10Y8_W1BEG[0] }),
    .W2BEG({\Tile_X9Y8_W2BEG[7] ,
    \Tile_X9Y8_W2BEG[6] ,
    \Tile_X9Y8_W2BEG[5] ,
    \Tile_X9Y8_W2BEG[4] ,
    \Tile_X9Y8_W2BEG[3] ,
    \Tile_X9Y8_W2BEG[2] ,
    \Tile_X9Y8_W2BEG[1] ,
    \Tile_X9Y8_W2BEG[0] }),
    .W2BEGb({\Tile_X9Y8_W2BEGb[7] ,
    \Tile_X9Y8_W2BEGb[6] ,
    \Tile_X9Y8_W2BEGb[5] ,
    \Tile_X9Y8_W2BEGb[4] ,
    \Tile_X9Y8_W2BEGb[3] ,
    \Tile_X9Y8_W2BEGb[2] ,
    \Tile_X9Y8_W2BEGb[1] ,
    \Tile_X9Y8_W2BEGb[0] }),
    .W2END({\Tile_X10Y8_W2BEGb[7] ,
    \Tile_X10Y8_W2BEGb[6] ,
    \Tile_X10Y8_W2BEGb[5] ,
    \Tile_X10Y8_W2BEGb[4] ,
    \Tile_X10Y8_W2BEGb[3] ,
    \Tile_X10Y8_W2BEGb[2] ,
    \Tile_X10Y8_W2BEGb[1] ,
    \Tile_X10Y8_W2BEGb[0] }),
    .W2MID({\Tile_X10Y8_W2BEG[7] ,
    \Tile_X10Y8_W2BEG[6] ,
    \Tile_X10Y8_W2BEG[5] ,
    \Tile_X10Y8_W2BEG[4] ,
    \Tile_X10Y8_W2BEG[3] ,
    \Tile_X10Y8_W2BEG[2] ,
    \Tile_X10Y8_W2BEG[1] ,
    \Tile_X10Y8_W2BEG[0] }),
    .W6BEG({\Tile_X9Y8_W6BEG[11] ,
    \Tile_X9Y8_W6BEG[10] ,
    \Tile_X9Y8_W6BEG[9] ,
    \Tile_X9Y8_W6BEG[8] ,
    \Tile_X9Y8_W6BEG[7] ,
    \Tile_X9Y8_W6BEG[6] ,
    \Tile_X9Y8_W6BEG[5] ,
    \Tile_X9Y8_W6BEG[4] ,
    \Tile_X9Y8_W6BEG[3] ,
    \Tile_X9Y8_W6BEG[2] ,
    \Tile_X9Y8_W6BEG[1] ,
    \Tile_X9Y8_W6BEG[0] }),
    .W6END({\Tile_X10Y8_W6BEG[11] ,
    \Tile_X10Y8_W6BEG[10] ,
    \Tile_X10Y8_W6BEG[9] ,
    \Tile_X10Y8_W6BEG[8] ,
    \Tile_X10Y8_W6BEG[7] ,
    \Tile_X10Y8_W6BEG[6] ,
    \Tile_X10Y8_W6BEG[5] ,
    \Tile_X10Y8_W6BEG[4] ,
    \Tile_X10Y8_W6BEG[3] ,
    \Tile_X10Y8_W6BEG[2] ,
    \Tile_X10Y8_W6BEG[1] ,
    \Tile_X10Y8_W6BEG[0] }),
    .WW4BEG({\Tile_X9Y8_WW4BEG[15] ,
    \Tile_X9Y8_WW4BEG[14] ,
    \Tile_X9Y8_WW4BEG[13] ,
    \Tile_X9Y8_WW4BEG[12] ,
    \Tile_X9Y8_WW4BEG[11] ,
    \Tile_X9Y8_WW4BEG[10] ,
    \Tile_X9Y8_WW4BEG[9] ,
    \Tile_X9Y8_WW4BEG[8] ,
    \Tile_X9Y8_WW4BEG[7] ,
    \Tile_X9Y8_WW4BEG[6] ,
    \Tile_X9Y8_WW4BEG[5] ,
    \Tile_X9Y8_WW4BEG[4] ,
    \Tile_X9Y8_WW4BEG[3] ,
    \Tile_X9Y8_WW4BEG[2] ,
    \Tile_X9Y8_WW4BEG[1] ,
    \Tile_X9Y8_WW4BEG[0] }),
    .WW4END({\Tile_X10Y8_WW4BEG[15] ,
    \Tile_X10Y8_WW4BEG[14] ,
    \Tile_X10Y8_WW4BEG[13] ,
    \Tile_X10Y8_WW4BEG[12] ,
    \Tile_X10Y8_WW4BEG[11] ,
    \Tile_X10Y8_WW4BEG[10] ,
    \Tile_X10Y8_WW4BEG[9] ,
    \Tile_X10Y8_WW4BEG[8] ,
    \Tile_X10Y8_WW4BEG[7] ,
    \Tile_X10Y8_WW4BEG[6] ,
    \Tile_X10Y8_WW4BEG[5] ,
    \Tile_X10Y8_WW4BEG[4] ,
    \Tile_X10Y8_WW4BEG[3] ,
    \Tile_X10Y8_WW4BEG[2] ,
    \Tile_X10Y8_WW4BEG[1] ,
    \Tile_X10Y8_WW4BEG[0] }));
 LUT4AB Tile_X9Y9_LUT4AB (.Ci(Tile_X9Y10_Co),
    .Co(Tile_X9Y9_Co),
    .UserCLK(Tile_X9Y10_UserCLKo),
    .UserCLKo(Tile_X9Y9_UserCLKo),
    .VGND(VGND),
    .VPWR(VPWR),
    .E1BEG({\Tile_X9Y9_E1BEG[3] ,
    \Tile_X9Y9_E1BEG[2] ,
    \Tile_X9Y9_E1BEG[1] ,
    \Tile_X9Y9_E1BEG[0] }),
    .E1END({\Tile_X8Y9_E1BEG[3] ,
    \Tile_X8Y9_E1BEG[2] ,
    \Tile_X8Y9_E1BEG[1] ,
    \Tile_X8Y9_E1BEG[0] }),
    .E2BEG({\Tile_X9Y9_E2BEG[7] ,
    \Tile_X9Y9_E2BEG[6] ,
    \Tile_X9Y9_E2BEG[5] ,
    \Tile_X9Y9_E2BEG[4] ,
    \Tile_X9Y9_E2BEG[3] ,
    \Tile_X9Y9_E2BEG[2] ,
    \Tile_X9Y9_E2BEG[1] ,
    \Tile_X9Y9_E2BEG[0] }),
    .E2BEGb({\Tile_X9Y9_E2BEGb[7] ,
    \Tile_X9Y9_E2BEGb[6] ,
    \Tile_X9Y9_E2BEGb[5] ,
    \Tile_X9Y9_E2BEGb[4] ,
    \Tile_X9Y9_E2BEGb[3] ,
    \Tile_X9Y9_E2BEGb[2] ,
    \Tile_X9Y9_E2BEGb[1] ,
    \Tile_X9Y9_E2BEGb[0] }),
    .E2END({\Tile_X8Y9_E2BEGb[7] ,
    \Tile_X8Y9_E2BEGb[6] ,
    \Tile_X8Y9_E2BEGb[5] ,
    \Tile_X8Y9_E2BEGb[4] ,
    \Tile_X8Y9_E2BEGb[3] ,
    \Tile_X8Y9_E2BEGb[2] ,
    \Tile_X8Y9_E2BEGb[1] ,
    \Tile_X8Y9_E2BEGb[0] }),
    .E2MID({\Tile_X8Y9_E2BEG[7] ,
    \Tile_X8Y9_E2BEG[6] ,
    \Tile_X8Y9_E2BEG[5] ,
    \Tile_X8Y9_E2BEG[4] ,
    \Tile_X8Y9_E2BEG[3] ,
    \Tile_X8Y9_E2BEG[2] ,
    \Tile_X8Y9_E2BEG[1] ,
    \Tile_X8Y9_E2BEG[0] }),
    .E6BEG({\Tile_X9Y9_E6BEG[11] ,
    \Tile_X9Y9_E6BEG[10] ,
    \Tile_X9Y9_E6BEG[9] ,
    \Tile_X9Y9_E6BEG[8] ,
    \Tile_X9Y9_E6BEG[7] ,
    \Tile_X9Y9_E6BEG[6] ,
    \Tile_X9Y9_E6BEG[5] ,
    \Tile_X9Y9_E6BEG[4] ,
    \Tile_X9Y9_E6BEG[3] ,
    \Tile_X9Y9_E6BEG[2] ,
    \Tile_X9Y9_E6BEG[1] ,
    \Tile_X9Y9_E6BEG[0] }),
    .E6END({\Tile_X8Y9_E6BEG[11] ,
    \Tile_X8Y9_E6BEG[10] ,
    \Tile_X8Y9_E6BEG[9] ,
    \Tile_X8Y9_E6BEG[8] ,
    \Tile_X8Y9_E6BEG[7] ,
    \Tile_X8Y9_E6BEG[6] ,
    \Tile_X8Y9_E6BEG[5] ,
    \Tile_X8Y9_E6BEG[4] ,
    \Tile_X8Y9_E6BEG[3] ,
    \Tile_X8Y9_E6BEG[2] ,
    \Tile_X8Y9_E6BEG[1] ,
    \Tile_X8Y9_E6BEG[0] }),
    .EE4BEG({\Tile_X9Y9_EE4BEG[15] ,
    \Tile_X9Y9_EE4BEG[14] ,
    \Tile_X9Y9_EE4BEG[13] ,
    \Tile_X9Y9_EE4BEG[12] ,
    \Tile_X9Y9_EE4BEG[11] ,
    \Tile_X9Y9_EE4BEG[10] ,
    \Tile_X9Y9_EE4BEG[9] ,
    \Tile_X9Y9_EE4BEG[8] ,
    \Tile_X9Y9_EE4BEG[7] ,
    \Tile_X9Y9_EE4BEG[6] ,
    \Tile_X9Y9_EE4BEG[5] ,
    \Tile_X9Y9_EE4BEG[4] ,
    \Tile_X9Y9_EE4BEG[3] ,
    \Tile_X9Y9_EE4BEG[2] ,
    \Tile_X9Y9_EE4BEG[1] ,
    \Tile_X9Y9_EE4BEG[0] }),
    .EE4END({\Tile_X8Y9_EE4BEG[15] ,
    \Tile_X8Y9_EE4BEG[14] ,
    \Tile_X8Y9_EE4BEG[13] ,
    \Tile_X8Y9_EE4BEG[12] ,
    \Tile_X8Y9_EE4BEG[11] ,
    \Tile_X8Y9_EE4BEG[10] ,
    \Tile_X8Y9_EE4BEG[9] ,
    \Tile_X8Y9_EE4BEG[8] ,
    \Tile_X8Y9_EE4BEG[7] ,
    \Tile_X8Y9_EE4BEG[6] ,
    \Tile_X8Y9_EE4BEG[5] ,
    \Tile_X8Y9_EE4BEG[4] ,
    \Tile_X8Y9_EE4BEG[3] ,
    \Tile_X8Y9_EE4BEG[2] ,
    \Tile_X8Y9_EE4BEG[1] ,
    \Tile_X8Y9_EE4BEG[0] }),
    .FrameData({\Tile_X8Y9_FrameData_O[31] ,
    \Tile_X8Y9_FrameData_O[30] ,
    \Tile_X8Y9_FrameData_O[29] ,
    \Tile_X8Y9_FrameData_O[28] ,
    \Tile_X8Y9_FrameData_O[27] ,
    \Tile_X8Y9_FrameData_O[26] ,
    \Tile_X8Y9_FrameData_O[25] ,
    \Tile_X8Y9_FrameData_O[24] ,
    \Tile_X8Y9_FrameData_O[23] ,
    \Tile_X8Y9_FrameData_O[22] ,
    \Tile_X8Y9_FrameData_O[21] ,
    \Tile_X8Y9_FrameData_O[20] ,
    \Tile_X8Y9_FrameData_O[19] ,
    \Tile_X8Y9_FrameData_O[18] ,
    \Tile_X8Y9_FrameData_O[17] ,
    \Tile_X8Y9_FrameData_O[16] ,
    \Tile_X8Y9_FrameData_O[15] ,
    \Tile_X8Y9_FrameData_O[14] ,
    \Tile_X8Y9_FrameData_O[13] ,
    \Tile_X8Y9_FrameData_O[12] ,
    \Tile_X8Y9_FrameData_O[11] ,
    \Tile_X8Y9_FrameData_O[10] ,
    \Tile_X8Y9_FrameData_O[9] ,
    \Tile_X8Y9_FrameData_O[8] ,
    \Tile_X8Y9_FrameData_O[7] ,
    \Tile_X8Y9_FrameData_O[6] ,
    \Tile_X8Y9_FrameData_O[5] ,
    \Tile_X8Y9_FrameData_O[4] ,
    \Tile_X8Y9_FrameData_O[3] ,
    \Tile_X8Y9_FrameData_O[2] ,
    \Tile_X8Y9_FrameData_O[1] ,
    \Tile_X8Y9_FrameData_O[0] }),
    .FrameData_O({\Tile_X9Y9_FrameData_O[31] ,
    \Tile_X9Y9_FrameData_O[30] ,
    \Tile_X9Y9_FrameData_O[29] ,
    \Tile_X9Y9_FrameData_O[28] ,
    \Tile_X9Y9_FrameData_O[27] ,
    \Tile_X9Y9_FrameData_O[26] ,
    \Tile_X9Y9_FrameData_O[25] ,
    \Tile_X9Y9_FrameData_O[24] ,
    \Tile_X9Y9_FrameData_O[23] ,
    \Tile_X9Y9_FrameData_O[22] ,
    \Tile_X9Y9_FrameData_O[21] ,
    \Tile_X9Y9_FrameData_O[20] ,
    \Tile_X9Y9_FrameData_O[19] ,
    \Tile_X9Y9_FrameData_O[18] ,
    \Tile_X9Y9_FrameData_O[17] ,
    \Tile_X9Y9_FrameData_O[16] ,
    \Tile_X9Y9_FrameData_O[15] ,
    \Tile_X9Y9_FrameData_O[14] ,
    \Tile_X9Y9_FrameData_O[13] ,
    \Tile_X9Y9_FrameData_O[12] ,
    \Tile_X9Y9_FrameData_O[11] ,
    \Tile_X9Y9_FrameData_O[10] ,
    \Tile_X9Y9_FrameData_O[9] ,
    \Tile_X9Y9_FrameData_O[8] ,
    \Tile_X9Y9_FrameData_O[7] ,
    \Tile_X9Y9_FrameData_O[6] ,
    \Tile_X9Y9_FrameData_O[5] ,
    \Tile_X9Y9_FrameData_O[4] ,
    \Tile_X9Y9_FrameData_O[3] ,
    \Tile_X9Y9_FrameData_O[2] ,
    \Tile_X9Y9_FrameData_O[1] ,
    \Tile_X9Y9_FrameData_O[0] }),
    .FrameStrobe({\Tile_X9Y10_FrameStrobe_O[19] ,
    \Tile_X9Y10_FrameStrobe_O[18] ,
    \Tile_X9Y10_FrameStrobe_O[17] ,
    \Tile_X9Y10_FrameStrobe_O[16] ,
    \Tile_X9Y10_FrameStrobe_O[15] ,
    \Tile_X9Y10_FrameStrobe_O[14] ,
    \Tile_X9Y10_FrameStrobe_O[13] ,
    \Tile_X9Y10_FrameStrobe_O[12] ,
    \Tile_X9Y10_FrameStrobe_O[11] ,
    \Tile_X9Y10_FrameStrobe_O[10] ,
    \Tile_X9Y10_FrameStrobe_O[9] ,
    \Tile_X9Y10_FrameStrobe_O[8] ,
    \Tile_X9Y10_FrameStrobe_O[7] ,
    \Tile_X9Y10_FrameStrobe_O[6] ,
    \Tile_X9Y10_FrameStrobe_O[5] ,
    \Tile_X9Y10_FrameStrobe_O[4] ,
    \Tile_X9Y10_FrameStrobe_O[3] ,
    \Tile_X9Y10_FrameStrobe_O[2] ,
    \Tile_X9Y10_FrameStrobe_O[1] ,
    \Tile_X9Y10_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Tile_X9Y9_FrameStrobe_O[19] ,
    \Tile_X9Y9_FrameStrobe_O[18] ,
    \Tile_X9Y9_FrameStrobe_O[17] ,
    \Tile_X9Y9_FrameStrobe_O[16] ,
    \Tile_X9Y9_FrameStrobe_O[15] ,
    \Tile_X9Y9_FrameStrobe_O[14] ,
    \Tile_X9Y9_FrameStrobe_O[13] ,
    \Tile_X9Y9_FrameStrobe_O[12] ,
    \Tile_X9Y9_FrameStrobe_O[11] ,
    \Tile_X9Y9_FrameStrobe_O[10] ,
    \Tile_X9Y9_FrameStrobe_O[9] ,
    \Tile_X9Y9_FrameStrobe_O[8] ,
    \Tile_X9Y9_FrameStrobe_O[7] ,
    \Tile_X9Y9_FrameStrobe_O[6] ,
    \Tile_X9Y9_FrameStrobe_O[5] ,
    \Tile_X9Y9_FrameStrobe_O[4] ,
    \Tile_X9Y9_FrameStrobe_O[3] ,
    \Tile_X9Y9_FrameStrobe_O[2] ,
    \Tile_X9Y9_FrameStrobe_O[1] ,
    \Tile_X9Y9_FrameStrobe_O[0] }),
    .N1BEG({\Tile_X9Y9_N1BEG[3] ,
    \Tile_X9Y9_N1BEG[2] ,
    \Tile_X9Y9_N1BEG[1] ,
    \Tile_X9Y9_N1BEG[0] }),
    .N1END({\Tile_X9Y10_N1BEG[3] ,
    \Tile_X9Y10_N1BEG[2] ,
    \Tile_X9Y10_N1BEG[1] ,
    \Tile_X9Y10_N1BEG[0] }),
    .N2BEG({\Tile_X9Y9_N2BEG[7] ,
    \Tile_X9Y9_N2BEG[6] ,
    \Tile_X9Y9_N2BEG[5] ,
    \Tile_X9Y9_N2BEG[4] ,
    \Tile_X9Y9_N2BEG[3] ,
    \Tile_X9Y9_N2BEG[2] ,
    \Tile_X9Y9_N2BEG[1] ,
    \Tile_X9Y9_N2BEG[0] }),
    .N2BEGb({\Tile_X9Y9_N2BEGb[7] ,
    \Tile_X9Y9_N2BEGb[6] ,
    \Tile_X9Y9_N2BEGb[5] ,
    \Tile_X9Y9_N2BEGb[4] ,
    \Tile_X9Y9_N2BEGb[3] ,
    \Tile_X9Y9_N2BEGb[2] ,
    \Tile_X9Y9_N2BEGb[1] ,
    \Tile_X9Y9_N2BEGb[0] }),
    .N2END({\Tile_X9Y10_N2BEGb[7] ,
    \Tile_X9Y10_N2BEGb[6] ,
    \Tile_X9Y10_N2BEGb[5] ,
    \Tile_X9Y10_N2BEGb[4] ,
    \Tile_X9Y10_N2BEGb[3] ,
    \Tile_X9Y10_N2BEGb[2] ,
    \Tile_X9Y10_N2BEGb[1] ,
    \Tile_X9Y10_N2BEGb[0] }),
    .N2MID({\Tile_X9Y10_N2BEG[7] ,
    \Tile_X9Y10_N2BEG[6] ,
    \Tile_X9Y10_N2BEG[5] ,
    \Tile_X9Y10_N2BEG[4] ,
    \Tile_X9Y10_N2BEG[3] ,
    \Tile_X9Y10_N2BEG[2] ,
    \Tile_X9Y10_N2BEG[1] ,
    \Tile_X9Y10_N2BEG[0] }),
    .N4BEG({\Tile_X9Y9_N4BEG[15] ,
    \Tile_X9Y9_N4BEG[14] ,
    \Tile_X9Y9_N4BEG[13] ,
    \Tile_X9Y9_N4BEG[12] ,
    \Tile_X9Y9_N4BEG[11] ,
    \Tile_X9Y9_N4BEG[10] ,
    \Tile_X9Y9_N4BEG[9] ,
    \Tile_X9Y9_N4BEG[8] ,
    \Tile_X9Y9_N4BEG[7] ,
    \Tile_X9Y9_N4BEG[6] ,
    \Tile_X9Y9_N4BEG[5] ,
    \Tile_X9Y9_N4BEG[4] ,
    \Tile_X9Y9_N4BEG[3] ,
    \Tile_X9Y9_N4BEG[2] ,
    \Tile_X9Y9_N4BEG[1] ,
    \Tile_X9Y9_N4BEG[0] }),
    .N4END({\Tile_X9Y10_N4BEG[15] ,
    \Tile_X9Y10_N4BEG[14] ,
    \Tile_X9Y10_N4BEG[13] ,
    \Tile_X9Y10_N4BEG[12] ,
    \Tile_X9Y10_N4BEG[11] ,
    \Tile_X9Y10_N4BEG[10] ,
    \Tile_X9Y10_N4BEG[9] ,
    \Tile_X9Y10_N4BEG[8] ,
    \Tile_X9Y10_N4BEG[7] ,
    \Tile_X9Y10_N4BEG[6] ,
    \Tile_X9Y10_N4BEG[5] ,
    \Tile_X9Y10_N4BEG[4] ,
    \Tile_X9Y10_N4BEG[3] ,
    \Tile_X9Y10_N4BEG[2] ,
    \Tile_X9Y10_N4BEG[1] ,
    \Tile_X9Y10_N4BEG[0] }),
    .NN4BEG({\Tile_X9Y9_NN4BEG[15] ,
    \Tile_X9Y9_NN4BEG[14] ,
    \Tile_X9Y9_NN4BEG[13] ,
    \Tile_X9Y9_NN4BEG[12] ,
    \Tile_X9Y9_NN4BEG[11] ,
    \Tile_X9Y9_NN4BEG[10] ,
    \Tile_X9Y9_NN4BEG[9] ,
    \Tile_X9Y9_NN4BEG[8] ,
    \Tile_X9Y9_NN4BEG[7] ,
    \Tile_X9Y9_NN4BEG[6] ,
    \Tile_X9Y9_NN4BEG[5] ,
    \Tile_X9Y9_NN4BEG[4] ,
    \Tile_X9Y9_NN4BEG[3] ,
    \Tile_X9Y9_NN4BEG[2] ,
    \Tile_X9Y9_NN4BEG[1] ,
    \Tile_X9Y9_NN4BEG[0] }),
    .NN4END({\Tile_X9Y10_NN4BEG[15] ,
    \Tile_X9Y10_NN4BEG[14] ,
    \Tile_X9Y10_NN4BEG[13] ,
    \Tile_X9Y10_NN4BEG[12] ,
    \Tile_X9Y10_NN4BEG[11] ,
    \Tile_X9Y10_NN4BEG[10] ,
    \Tile_X9Y10_NN4BEG[9] ,
    \Tile_X9Y10_NN4BEG[8] ,
    \Tile_X9Y10_NN4BEG[7] ,
    \Tile_X9Y10_NN4BEG[6] ,
    \Tile_X9Y10_NN4BEG[5] ,
    \Tile_X9Y10_NN4BEG[4] ,
    \Tile_X9Y10_NN4BEG[3] ,
    \Tile_X9Y10_NN4BEG[2] ,
    \Tile_X9Y10_NN4BEG[1] ,
    \Tile_X9Y10_NN4BEG[0] }),
    .S1BEG({\Tile_X9Y9_S1BEG[3] ,
    \Tile_X9Y9_S1BEG[2] ,
    \Tile_X9Y9_S1BEG[1] ,
    \Tile_X9Y9_S1BEG[0] }),
    .S1END({\Tile_X9Y8_S1BEG[3] ,
    \Tile_X9Y8_S1BEG[2] ,
    \Tile_X9Y8_S1BEG[1] ,
    \Tile_X9Y8_S1BEG[0] }),
    .S2BEG({\Tile_X9Y9_S2BEG[7] ,
    \Tile_X9Y9_S2BEG[6] ,
    \Tile_X9Y9_S2BEG[5] ,
    \Tile_X9Y9_S2BEG[4] ,
    \Tile_X9Y9_S2BEG[3] ,
    \Tile_X9Y9_S2BEG[2] ,
    \Tile_X9Y9_S2BEG[1] ,
    \Tile_X9Y9_S2BEG[0] }),
    .S2BEGb({\Tile_X9Y9_S2BEGb[7] ,
    \Tile_X9Y9_S2BEGb[6] ,
    \Tile_X9Y9_S2BEGb[5] ,
    \Tile_X9Y9_S2BEGb[4] ,
    \Tile_X9Y9_S2BEGb[3] ,
    \Tile_X9Y9_S2BEGb[2] ,
    \Tile_X9Y9_S2BEGb[1] ,
    \Tile_X9Y9_S2BEGb[0] }),
    .S2END({\Tile_X9Y8_S2BEGb[7] ,
    \Tile_X9Y8_S2BEGb[6] ,
    \Tile_X9Y8_S2BEGb[5] ,
    \Tile_X9Y8_S2BEGb[4] ,
    \Tile_X9Y8_S2BEGb[3] ,
    \Tile_X9Y8_S2BEGb[2] ,
    \Tile_X9Y8_S2BEGb[1] ,
    \Tile_X9Y8_S2BEGb[0] }),
    .S2MID({\Tile_X9Y8_S2BEG[7] ,
    \Tile_X9Y8_S2BEG[6] ,
    \Tile_X9Y8_S2BEG[5] ,
    \Tile_X9Y8_S2BEG[4] ,
    \Tile_X9Y8_S2BEG[3] ,
    \Tile_X9Y8_S2BEG[2] ,
    \Tile_X9Y8_S2BEG[1] ,
    \Tile_X9Y8_S2BEG[0] }),
    .S4BEG({\Tile_X9Y9_S4BEG[15] ,
    \Tile_X9Y9_S4BEG[14] ,
    \Tile_X9Y9_S4BEG[13] ,
    \Tile_X9Y9_S4BEG[12] ,
    \Tile_X9Y9_S4BEG[11] ,
    \Tile_X9Y9_S4BEG[10] ,
    \Tile_X9Y9_S4BEG[9] ,
    \Tile_X9Y9_S4BEG[8] ,
    \Tile_X9Y9_S4BEG[7] ,
    \Tile_X9Y9_S4BEG[6] ,
    \Tile_X9Y9_S4BEG[5] ,
    \Tile_X9Y9_S4BEG[4] ,
    \Tile_X9Y9_S4BEG[3] ,
    \Tile_X9Y9_S4BEG[2] ,
    \Tile_X9Y9_S4BEG[1] ,
    \Tile_X9Y9_S4BEG[0] }),
    .S4END({\Tile_X9Y8_S4BEG[15] ,
    \Tile_X9Y8_S4BEG[14] ,
    \Tile_X9Y8_S4BEG[13] ,
    \Tile_X9Y8_S4BEG[12] ,
    \Tile_X9Y8_S4BEG[11] ,
    \Tile_X9Y8_S4BEG[10] ,
    \Tile_X9Y8_S4BEG[9] ,
    \Tile_X9Y8_S4BEG[8] ,
    \Tile_X9Y8_S4BEG[7] ,
    \Tile_X9Y8_S4BEG[6] ,
    \Tile_X9Y8_S4BEG[5] ,
    \Tile_X9Y8_S4BEG[4] ,
    \Tile_X9Y8_S4BEG[3] ,
    \Tile_X9Y8_S4BEG[2] ,
    \Tile_X9Y8_S4BEG[1] ,
    \Tile_X9Y8_S4BEG[0] }),
    .SS4BEG({\Tile_X9Y9_SS4BEG[15] ,
    \Tile_X9Y9_SS4BEG[14] ,
    \Tile_X9Y9_SS4BEG[13] ,
    \Tile_X9Y9_SS4BEG[12] ,
    \Tile_X9Y9_SS4BEG[11] ,
    \Tile_X9Y9_SS4BEG[10] ,
    \Tile_X9Y9_SS4BEG[9] ,
    \Tile_X9Y9_SS4BEG[8] ,
    \Tile_X9Y9_SS4BEG[7] ,
    \Tile_X9Y9_SS4BEG[6] ,
    \Tile_X9Y9_SS4BEG[5] ,
    \Tile_X9Y9_SS4BEG[4] ,
    \Tile_X9Y9_SS4BEG[3] ,
    \Tile_X9Y9_SS4BEG[2] ,
    \Tile_X9Y9_SS4BEG[1] ,
    \Tile_X9Y9_SS4BEG[0] }),
    .SS4END({\Tile_X9Y8_SS4BEG[15] ,
    \Tile_X9Y8_SS4BEG[14] ,
    \Tile_X9Y8_SS4BEG[13] ,
    \Tile_X9Y8_SS4BEG[12] ,
    \Tile_X9Y8_SS4BEG[11] ,
    \Tile_X9Y8_SS4BEG[10] ,
    \Tile_X9Y8_SS4BEG[9] ,
    \Tile_X9Y8_SS4BEG[8] ,
    \Tile_X9Y8_SS4BEG[7] ,
    \Tile_X9Y8_SS4BEG[6] ,
    \Tile_X9Y8_SS4BEG[5] ,
    \Tile_X9Y8_SS4BEG[4] ,
    \Tile_X9Y8_SS4BEG[3] ,
    \Tile_X9Y8_SS4BEG[2] ,
    \Tile_X9Y8_SS4BEG[1] ,
    \Tile_X9Y8_SS4BEG[0] }),
    .W1BEG({\Tile_X9Y9_W1BEG[3] ,
    \Tile_X9Y9_W1BEG[2] ,
    \Tile_X9Y9_W1BEG[1] ,
    \Tile_X9Y9_W1BEG[0] }),
    .W1END({\Tile_X10Y9_W1BEG[3] ,
    \Tile_X10Y9_W1BEG[2] ,
    \Tile_X10Y9_W1BEG[1] ,
    \Tile_X10Y9_W1BEG[0] }),
    .W2BEG({\Tile_X9Y9_W2BEG[7] ,
    \Tile_X9Y9_W2BEG[6] ,
    \Tile_X9Y9_W2BEG[5] ,
    \Tile_X9Y9_W2BEG[4] ,
    \Tile_X9Y9_W2BEG[3] ,
    \Tile_X9Y9_W2BEG[2] ,
    \Tile_X9Y9_W2BEG[1] ,
    \Tile_X9Y9_W2BEG[0] }),
    .W2BEGb({\Tile_X9Y9_W2BEGb[7] ,
    \Tile_X9Y9_W2BEGb[6] ,
    \Tile_X9Y9_W2BEGb[5] ,
    \Tile_X9Y9_W2BEGb[4] ,
    \Tile_X9Y9_W2BEGb[3] ,
    \Tile_X9Y9_W2BEGb[2] ,
    \Tile_X9Y9_W2BEGb[1] ,
    \Tile_X9Y9_W2BEGb[0] }),
    .W2END({\Tile_X10Y9_W2BEGb[7] ,
    \Tile_X10Y9_W2BEGb[6] ,
    \Tile_X10Y9_W2BEGb[5] ,
    \Tile_X10Y9_W2BEGb[4] ,
    \Tile_X10Y9_W2BEGb[3] ,
    \Tile_X10Y9_W2BEGb[2] ,
    \Tile_X10Y9_W2BEGb[1] ,
    \Tile_X10Y9_W2BEGb[0] }),
    .W2MID({\Tile_X10Y9_W2BEG[7] ,
    \Tile_X10Y9_W2BEG[6] ,
    \Tile_X10Y9_W2BEG[5] ,
    \Tile_X10Y9_W2BEG[4] ,
    \Tile_X10Y9_W2BEG[3] ,
    \Tile_X10Y9_W2BEG[2] ,
    \Tile_X10Y9_W2BEG[1] ,
    \Tile_X10Y9_W2BEG[0] }),
    .W6BEG({\Tile_X9Y9_W6BEG[11] ,
    \Tile_X9Y9_W6BEG[10] ,
    \Tile_X9Y9_W6BEG[9] ,
    \Tile_X9Y9_W6BEG[8] ,
    \Tile_X9Y9_W6BEG[7] ,
    \Tile_X9Y9_W6BEG[6] ,
    \Tile_X9Y9_W6BEG[5] ,
    \Tile_X9Y9_W6BEG[4] ,
    \Tile_X9Y9_W6BEG[3] ,
    \Tile_X9Y9_W6BEG[2] ,
    \Tile_X9Y9_W6BEG[1] ,
    \Tile_X9Y9_W6BEG[0] }),
    .W6END({\Tile_X10Y9_W6BEG[11] ,
    \Tile_X10Y9_W6BEG[10] ,
    \Tile_X10Y9_W6BEG[9] ,
    \Tile_X10Y9_W6BEG[8] ,
    \Tile_X10Y9_W6BEG[7] ,
    \Tile_X10Y9_W6BEG[6] ,
    \Tile_X10Y9_W6BEG[5] ,
    \Tile_X10Y9_W6BEG[4] ,
    \Tile_X10Y9_W6BEG[3] ,
    \Tile_X10Y9_W6BEG[2] ,
    \Tile_X10Y9_W6BEG[1] ,
    \Tile_X10Y9_W6BEG[0] }),
    .WW4BEG({\Tile_X9Y9_WW4BEG[15] ,
    \Tile_X9Y9_WW4BEG[14] ,
    \Tile_X9Y9_WW4BEG[13] ,
    \Tile_X9Y9_WW4BEG[12] ,
    \Tile_X9Y9_WW4BEG[11] ,
    \Tile_X9Y9_WW4BEG[10] ,
    \Tile_X9Y9_WW4BEG[9] ,
    \Tile_X9Y9_WW4BEG[8] ,
    \Tile_X9Y9_WW4BEG[7] ,
    \Tile_X9Y9_WW4BEG[6] ,
    \Tile_X9Y9_WW4BEG[5] ,
    \Tile_X9Y9_WW4BEG[4] ,
    \Tile_X9Y9_WW4BEG[3] ,
    \Tile_X9Y9_WW4BEG[2] ,
    \Tile_X9Y9_WW4BEG[1] ,
    \Tile_X9Y9_WW4BEG[0] }),
    .WW4END({\Tile_X10Y9_WW4BEG[15] ,
    \Tile_X10Y9_WW4BEG[14] ,
    \Tile_X10Y9_WW4BEG[13] ,
    \Tile_X10Y9_WW4BEG[12] ,
    \Tile_X10Y9_WW4BEG[11] ,
    \Tile_X10Y9_WW4BEG[10] ,
    \Tile_X10Y9_WW4BEG[9] ,
    \Tile_X10Y9_WW4BEG[8] ,
    \Tile_X10Y9_WW4BEG[7] ,
    \Tile_X10Y9_WW4BEG[6] ,
    \Tile_X10Y9_WW4BEG[5] ,
    \Tile_X10Y9_WW4BEG[4] ,
    \Tile_X10Y9_WW4BEG[3] ,
    \Tile_X10Y9_WW4BEG[2] ,
    \Tile_X10Y9_WW4BEG[1] ,
    \Tile_X10Y9_WW4BEG[0] }));
endmodule
