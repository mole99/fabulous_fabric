VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO eFPGA
  CLASS BLOCK ;
  FOREIGN eFPGA ;
  ORIGIN 0.000 0.000 ;
  SIZE 2435.000 BY 3782.500 ;
  PIN FrameData[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 38.730 3778.500 39.010 3782.500 ;
    END
  END FrameData[0]
  PIN FrameData[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3104.240 4.000 3104.840 ;
    END
  END FrameData[100]
  PIN FrameData[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3107.640 4.000 3108.240 ;
    END
  END FrameData[101]
  PIN FrameData[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3114.440 4.000 3115.040 ;
    END
  END FrameData[102]
  PIN FrameData[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3117.840 4.000 3118.440 ;
    END
  END FrameData[103]
  PIN FrameData[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3121.240 4.000 3121.840 ;
    END
  END FrameData[104]
  PIN FrameData[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3124.640 4.000 3125.240 ;
    END
  END FrameData[105]
  PIN FrameData[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3128.040 4.000 3128.640 ;
    END
  END FrameData[106]
  PIN FrameData[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3134.840 4.000 3135.440 ;
    END
  END FrameData[107]
  PIN FrameData[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3138.240 4.000 3138.840 ;
    END
  END FrameData[108]
  PIN FrameData[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3141.640 4.000 3142.240 ;
    END
  END FrameData[109]
  PIN FrameData[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 106.350 3778.500 106.630 3782.500 ;
    END
  END FrameData[10]
  PIN FrameData[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3145.040 4.000 3145.640 ;
    END
  END FrameData[110]
  PIN FrameData[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3148.440 4.000 3149.040 ;
    END
  END FrameData[111]
  PIN FrameData[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3155.240 4.000 3155.840 ;
    END
  END FrameData[112]
  PIN FrameData[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3158.640 4.000 3159.240 ;
    END
  END FrameData[113]
  PIN FrameData[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3162.040 4.000 3162.640 ;
    END
  END FrameData[114]
  PIN FrameData[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3165.440 4.000 3166.040 ;
    END
  END FrameData[115]
  PIN FrameData[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3168.840 4.000 3169.440 ;
    END
  END FrameData[116]
  PIN FrameData[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3175.640 4.000 3176.240 ;
    END
  END FrameData[117]
  PIN FrameData[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3179.040 4.000 3179.640 ;
    END
  END FrameData[118]
  PIN FrameData[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3182.440 4.000 3183.040 ;
    END
  END FrameData[119]
  PIN FrameData[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 77.370 3778.500 77.650 3782.500 ;
    END
  END FrameData[11]
  PIN FrameData[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3185.840 4.000 3186.440 ;
    END
  END FrameData[120]
  PIN FrameData[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3189.240 4.000 3189.840 ;
    END
  END FrameData[121]
  PIN FrameData[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3196.040 4.000 3196.640 ;
    END
  END FrameData[122]
  PIN FrameData[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3199.440 4.000 3200.040 ;
    END
  END FrameData[123]
  PIN FrameData[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3202.840 4.000 3203.440 ;
    END
  END FrameData[124]
  PIN FrameData[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3206.240 4.000 3206.840 ;
    END
  END FrameData[125]
  PIN FrameData[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3209.640 4.000 3210.240 ;
    END
  END FrameData[126]
  PIN FrameData[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3216.440 4.000 3217.040 ;
    END
  END FrameData[127]
  PIN FrameData[128]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2862.840 4.000 2863.440 ;
    END
  END FrameData[128]
  PIN FrameData[129]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2866.240 4.000 2866.840 ;
    END
  END FrameData[129]
  PIN FrameData[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 61.270 3778.500 61.550 3782.500 ;
    END
  END FrameData[12]
  PIN FrameData[130]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2873.040 4.000 2873.640 ;
    END
  END FrameData[130]
  PIN FrameData[131]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2876.440 4.000 2877.040 ;
    END
  END FrameData[131]
  PIN FrameData[132]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2879.840 4.000 2880.440 ;
    END
  END FrameData[132]
  PIN FrameData[133]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2883.240 4.000 2883.840 ;
    END
  END FrameData[133]
  PIN FrameData[134]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2886.640 4.000 2887.240 ;
    END
  END FrameData[134]
  PIN FrameData[135]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2893.440 4.000 2894.040 ;
    END
  END FrameData[135]
  PIN FrameData[136]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2896.840 4.000 2897.440 ;
    END
  END FrameData[136]
  PIN FrameData[137]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2900.240 4.000 2900.840 ;
    END
  END FrameData[137]
  PIN FrameData[138]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2903.640 4.000 2904.240 ;
    END
  END FrameData[138]
  PIN FrameData[139]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2907.040 4.000 2907.640 ;
    END
  END FrameData[139]
  PIN FrameData[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 99.910 3778.500 100.190 3782.500 ;
    END
  END FrameData[13]
  PIN FrameData[140]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2913.840 4.000 2914.440 ;
    END
  END FrameData[140]
  PIN FrameData[141]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2917.240 4.000 2917.840 ;
    END
  END FrameData[141]
  PIN FrameData[142]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2920.640 4.000 2921.240 ;
    END
  END FrameData[142]
  PIN FrameData[143]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2924.040 4.000 2924.640 ;
    END
  END FrameData[143]
  PIN FrameData[144]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2927.440 4.000 2928.040 ;
    END
  END FrameData[144]
  PIN FrameData[145]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2934.240 4.000 2934.840 ;
    END
  END FrameData[145]
  PIN FrameData[146]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2937.640 4.000 2938.240 ;
    END
  END FrameData[146]
  PIN FrameData[147]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2941.040 4.000 2941.640 ;
    END
  END FrameData[147]
  PIN FrameData[148]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2944.440 4.000 2945.040 ;
    END
  END FrameData[148]
  PIN FrameData[149]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2947.840 4.000 2948.440 ;
    END
  END FrameData[149]
  PIN FrameData[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 103.130 3778.500 103.410 3782.500 ;
    END
  END FrameData[14]
  PIN FrameData[150]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2954.640 4.000 2955.240 ;
    END
  END FrameData[150]
  PIN FrameData[151]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2958.040 4.000 2958.640 ;
    END
  END FrameData[151]
  PIN FrameData[152]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2961.440 4.000 2962.040 ;
    END
  END FrameData[152]
  PIN FrameData[153]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2964.840 4.000 2965.440 ;
    END
  END FrameData[153]
  PIN FrameData[154]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2968.240 4.000 2968.840 ;
    END
  END FrameData[154]
  PIN FrameData[155]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2975.040 4.000 2975.640 ;
    END
  END FrameData[155]
  PIN FrameData[156]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2978.440 4.000 2979.040 ;
    END
  END FrameData[156]
  PIN FrameData[157]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2981.840 4.000 2982.440 ;
    END
  END FrameData[157]
  PIN FrameData[158]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2985.240 4.000 2985.840 ;
    END
  END FrameData[158]
  PIN FrameData[159]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2988.640 4.000 2989.240 ;
    END
  END FrameData[159]
  PIN FrameData[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 74.150 3778.500 74.430 3782.500 ;
    END
  END FrameData[15]
  PIN FrameData[160]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2638.440 4.000 2639.040 ;
    END
  END FrameData[160]
  PIN FrameData[161]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2641.840 4.000 2642.440 ;
    END
  END FrameData[161]
  PIN FrameData[162]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2648.640 4.000 2649.240 ;
    END
  END FrameData[162]
  PIN FrameData[163]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2652.040 4.000 2652.640 ;
    END
  END FrameData[163]
  PIN FrameData[164]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2655.440 4.000 2656.040 ;
    END
  END FrameData[164]
  PIN FrameData[165]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2658.840 4.000 2659.440 ;
    END
  END FrameData[165]
  PIN FrameData[166]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2662.240 4.000 2662.840 ;
    END
  END FrameData[166]
  PIN FrameData[167]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2669.040 4.000 2669.640 ;
    END
  END FrameData[167]
  PIN FrameData[168]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2672.440 4.000 2673.040 ;
    END
  END FrameData[168]
  PIN FrameData[169]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2675.840 4.000 2676.440 ;
    END
  END FrameData[169]
  PIN FrameData[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 51.610 3778.500 51.890 3782.500 ;
    END
  END FrameData[16]
  PIN FrameData[170]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2679.240 4.000 2679.840 ;
    END
  END FrameData[170]
  PIN FrameData[171]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2682.640 4.000 2683.240 ;
    END
  END FrameData[171]
  PIN FrameData[172]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2689.440 4.000 2690.040 ;
    END
  END FrameData[172]
  PIN FrameData[173]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2692.840 4.000 2693.440 ;
    END
  END FrameData[173]
  PIN FrameData[174]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2696.240 4.000 2696.840 ;
    END
  END FrameData[174]
  PIN FrameData[175]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2699.640 4.000 2700.240 ;
    END
  END FrameData[175]
  PIN FrameData[176]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2703.040 4.000 2703.640 ;
    END
  END FrameData[176]
  PIN FrameData[177]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2709.840 4.000 2710.440 ;
    END
  END FrameData[177]
  PIN FrameData[178]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2713.240 4.000 2713.840 ;
    END
  END FrameData[178]
  PIN FrameData[179]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2716.640 4.000 2717.240 ;
    END
  END FrameData[179]
  PIN FrameData[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 141.770 3778.500 142.050 3782.500 ;
    END
  END FrameData[17]
  PIN FrameData[180]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2720.040 4.000 2720.640 ;
    END
  END FrameData[180]
  PIN FrameData[181]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2723.440 4.000 2724.040 ;
    END
  END FrameData[181]
  PIN FrameData[182]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2730.240 4.000 2730.840 ;
    END
  END FrameData[182]
  PIN FrameData[183]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2733.640 4.000 2734.240 ;
    END
  END FrameData[183]
  PIN FrameData[184]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2737.040 4.000 2737.640 ;
    END
  END FrameData[184]
  PIN FrameData[185]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2740.440 4.000 2741.040 ;
    END
  END FrameData[185]
  PIN FrameData[186]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2743.840 4.000 2744.440 ;
    END
  END FrameData[186]
  PIN FrameData[187]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2750.640 4.000 2751.240 ;
    END
  END FrameData[187]
  PIN FrameData[188]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2754.040 4.000 2754.640 ;
    END
  END FrameData[188]
  PIN FrameData[189]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2757.440 4.000 2758.040 ;
    END
  END FrameData[189]
  PIN FrameData[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 87.030 3778.500 87.310 3782.500 ;
    END
  END FrameData[18]
  PIN FrameData[190]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2760.840 4.000 2761.440 ;
    END
  END FrameData[190]
  PIN FrameData[191]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2764.240 4.000 2764.840 ;
    END
  END FrameData[191]
  PIN FrameData[192]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2414.040 4.000 2414.640 ;
    END
  END FrameData[192]
  PIN FrameData[193]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2417.440 4.000 2418.040 ;
    END
  END FrameData[193]
  PIN FrameData[194]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2420.840 4.000 2421.440 ;
    END
  END FrameData[194]
  PIN FrameData[195]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2427.640 4.000 2428.240 ;
    END
  END FrameData[195]
  PIN FrameData[196]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2431.040 4.000 2431.640 ;
    END
  END FrameData[196]
  PIN FrameData[197]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2434.440 4.000 2435.040 ;
    END
  END FrameData[197]
  PIN FrameData[198]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2437.840 4.000 2438.440 ;
    END
  END FrameData[198]
  PIN FrameData[199]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2441.240 4.000 2441.840 ;
    END
  END FrameData[199]
  PIN FrameData[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 58.050 3778.500 58.330 3782.500 ;
    END
  END FrameData[19]
  PIN FrameData[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 70.930 3778.500 71.210 3782.500 ;
    END
  END FrameData[1]
  PIN FrameData[200]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2448.040 4.000 2448.640 ;
    END
  END FrameData[200]
  PIN FrameData[201]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2451.440 4.000 2452.040 ;
    END
  END FrameData[201]
  PIN FrameData[202]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2454.840 4.000 2455.440 ;
    END
  END FrameData[202]
  PIN FrameData[203]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2458.240 4.000 2458.840 ;
    END
  END FrameData[203]
  PIN FrameData[204]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2461.640 4.000 2462.240 ;
    END
  END FrameData[204]
  PIN FrameData[205]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2468.440 4.000 2469.040 ;
    END
  END FrameData[205]
  PIN FrameData[206]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2471.840 4.000 2472.440 ;
    END
  END FrameData[206]
  PIN FrameData[207]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2475.240 4.000 2475.840 ;
    END
  END FrameData[207]
  PIN FrameData[208]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2478.640 4.000 2479.240 ;
    END
  END FrameData[208]
  PIN FrameData[209]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2482.040 4.000 2482.640 ;
    END
  END FrameData[209]
  PIN FrameData[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 96.690 3778.500 96.970 3782.500 ;
    END
  END FrameData[20]
  PIN FrameData[210]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2488.840 4.000 2489.440 ;
    END
  END FrameData[210]
  PIN FrameData[211]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2492.240 4.000 2492.840 ;
    END
  END FrameData[211]
  PIN FrameData[212]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2495.640 4.000 2496.240 ;
    END
  END FrameData[212]
  PIN FrameData[213]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2499.040 4.000 2499.640 ;
    END
  END FrameData[213]
  PIN FrameData[214]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2502.440 4.000 2503.040 ;
    END
  END FrameData[214]
  PIN FrameData[215]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2509.240 4.000 2509.840 ;
    END
  END FrameData[215]
  PIN FrameData[216]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2512.640 4.000 2513.240 ;
    END
  END FrameData[216]
  PIN FrameData[217]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2516.040 4.000 2516.640 ;
    END
  END FrameData[217]
  PIN FrameData[218]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2519.440 4.000 2520.040 ;
    END
  END FrameData[218]
  PIN FrameData[219]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2522.840 4.000 2523.440 ;
    END
  END FrameData[219]
  PIN FrameData[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 112.790 3778.500 113.070 3782.500 ;
    END
  END FrameData[21]
  PIN FrameData[220]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2529.640 4.000 2530.240 ;
    END
  END FrameData[220]
  PIN FrameData[221]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2533.040 4.000 2533.640 ;
    END
  END FrameData[221]
  PIN FrameData[222]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2536.440 4.000 2537.040 ;
    END
  END FrameData[222]
  PIN FrameData[223]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2539.840 4.000 2540.440 ;
    END
  END FrameData[223]
  PIN FrameData[224]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2189.640 4.000 2190.240 ;
    END
  END FrameData[224]
  PIN FrameData[225]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2193.040 4.000 2193.640 ;
    END
  END FrameData[225]
  PIN FrameData[226]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2196.440 4.000 2197.040 ;
    END
  END FrameData[226]
  PIN FrameData[227]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2199.840 4.000 2200.440 ;
    END
  END FrameData[227]
  PIN FrameData[228]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2206.640 4.000 2207.240 ;
    END
  END FrameData[228]
  PIN FrameData[229]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2210.040 4.000 2210.640 ;
    END
  END FrameData[229]
  PIN FrameData[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 119.230 3778.500 119.510 3782.500 ;
    END
  END FrameData[22]
  PIN FrameData[230]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2213.440 4.000 2214.040 ;
    END
  END FrameData[230]
  PIN FrameData[231]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2216.840 4.000 2217.440 ;
    END
  END FrameData[231]
  PIN FrameData[232]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2220.240 4.000 2220.840 ;
    END
  END FrameData[232]
  PIN FrameData[233]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2227.040 4.000 2227.640 ;
    END
  END FrameData[233]
  PIN FrameData[234]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2230.440 4.000 2231.040 ;
    END
  END FrameData[234]
  PIN FrameData[235]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2233.840 4.000 2234.440 ;
    END
  END FrameData[235]
  PIN FrameData[236]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2237.240 4.000 2237.840 ;
    END
  END FrameData[236]
  PIN FrameData[237]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2240.640 4.000 2241.240 ;
    END
  END FrameData[237]
  PIN FrameData[238]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2247.440 4.000 2248.040 ;
    END
  END FrameData[238]
  PIN FrameData[239]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2250.840 4.000 2251.440 ;
    END
  END FrameData[239]
  PIN FrameData[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 67.710 3778.500 67.990 3782.500 ;
    END
  END FrameData[23]
  PIN FrameData[240]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2254.240 4.000 2254.840 ;
    END
  END FrameData[240]
  PIN FrameData[241]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2257.640 4.000 2258.240 ;
    END
  END FrameData[241]
  PIN FrameData[242]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2261.040 4.000 2261.640 ;
    END
  END FrameData[242]
  PIN FrameData[243]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2267.840 4.000 2268.440 ;
    END
  END FrameData[243]
  PIN FrameData[244]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2271.240 4.000 2271.840 ;
    END
  END FrameData[244]
  PIN FrameData[245]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2274.640 4.000 2275.240 ;
    END
  END FrameData[245]
  PIN FrameData[246]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2278.040 4.000 2278.640 ;
    END
  END FrameData[246]
  PIN FrameData[247]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2281.440 4.000 2282.040 ;
    END
  END FrameData[247]
  PIN FrameData[248]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2288.240 4.000 2288.840 ;
    END
  END FrameData[248]
  PIN FrameData[249]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2291.640 4.000 2292.240 ;
    END
  END FrameData[249]
  PIN FrameData[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 93.470 3778.500 93.750 3782.500 ;
    END
  END FrameData[24]
  PIN FrameData[250]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2295.040 4.000 2295.640 ;
    END
  END FrameData[250]
  PIN FrameData[251]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2298.440 4.000 2299.040 ;
    END
  END FrameData[251]
  PIN FrameData[252]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2301.840 4.000 2302.440 ;
    END
  END FrameData[252]
  PIN FrameData[253]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2308.640 4.000 2309.240 ;
    END
  END FrameData[253]
  PIN FrameData[254]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2312.040 4.000 2312.640 ;
    END
  END FrameData[254]
  PIN FrameData[255]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2315.440 4.000 2316.040 ;
    END
  END FrameData[255]
  PIN FrameData[256]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1965.240 4.000 1965.840 ;
    END
  END FrameData[256]
  PIN FrameData[257]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1968.640 4.000 1969.240 ;
    END
  END FrameData[257]
  PIN FrameData[258]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1972.040 4.000 1972.640 ;
    END
  END FrameData[258]
  PIN FrameData[259]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1975.440 4.000 1976.040 ;
    END
  END FrameData[259]
  PIN FrameData[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 41.950 3778.500 42.230 3782.500 ;
    END
  END FrameData[25]
  PIN FrameData[260]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1978.840 4.000 1979.440 ;
    END
  END FrameData[260]
  PIN FrameData[261]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1985.640 4.000 1986.240 ;
    END
  END FrameData[261]
  PIN FrameData[262]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1989.040 4.000 1989.640 ;
    END
  END FrameData[262]
  PIN FrameData[263]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1992.440 4.000 1993.040 ;
    END
  END FrameData[263]
  PIN FrameData[264]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1995.840 4.000 1996.440 ;
    END
  END FrameData[264]
  PIN FrameData[265]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1999.240 4.000 1999.840 ;
    END
  END FrameData[265]
  PIN FrameData[266]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2006.040 4.000 2006.640 ;
    END
  END FrameData[266]
  PIN FrameData[267]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2009.440 4.000 2010.040 ;
    END
  END FrameData[267]
  PIN FrameData[268]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2012.840 4.000 2013.440 ;
    END
  END FrameData[268]
  PIN FrameData[269]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2016.240 4.000 2016.840 ;
    END
  END FrameData[269]
  PIN FrameData[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 157.870 3778.500 158.150 3782.500 ;
    END
  END FrameData[26]
  PIN FrameData[270]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2019.640 4.000 2020.240 ;
    END
  END FrameData[270]
  PIN FrameData[271]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2026.440 4.000 2027.040 ;
    END
  END FrameData[271]
  PIN FrameData[272]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2029.840 4.000 2030.440 ;
    END
  END FrameData[272]
  PIN FrameData[273]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2033.240 4.000 2033.840 ;
    END
  END FrameData[273]
  PIN FrameData[274]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2036.640 4.000 2037.240 ;
    END
  END FrameData[274]
  PIN FrameData[275]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2040.040 4.000 2040.640 ;
    END
  END FrameData[275]
  PIN FrameData[276]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2046.840 4.000 2047.440 ;
    END
  END FrameData[276]
  PIN FrameData[277]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2050.240 4.000 2050.840 ;
    END
  END FrameData[277]
  PIN FrameData[278]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2053.640 4.000 2054.240 ;
    END
  END FrameData[278]
  PIN FrameData[279]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2057.040 4.000 2057.640 ;
    END
  END FrameData[279]
  PIN FrameData[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 90.250 3778.500 90.530 3782.500 ;
    END
  END FrameData[27]
  PIN FrameData[280]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2060.440 4.000 2061.040 ;
    END
  END FrameData[280]
  PIN FrameData[281]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2067.240 4.000 2067.840 ;
    END
  END FrameData[281]
  PIN FrameData[282]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2070.640 4.000 2071.240 ;
    END
  END FrameData[282]
  PIN FrameData[283]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2074.040 4.000 2074.640 ;
    END
  END FrameData[283]
  PIN FrameData[284]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2077.440 4.000 2078.040 ;
    END
  END FrameData[284]
  PIN FrameData[285]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2080.840 4.000 2081.440 ;
    END
  END FrameData[285]
  PIN FrameData[286]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2087.640 4.000 2088.240 ;
    END
  END FrameData[286]
  PIN FrameData[287]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2091.040 4.000 2091.640 ;
    END
  END FrameData[287]
  PIN FrameData[288]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1737.440 4.000 1738.040 ;
    END
  END FrameData[288]
  PIN FrameData[289]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1740.840 4.000 1741.440 ;
    END
  END FrameData[289]
  PIN FrameData[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 48.390 3778.500 48.670 3782.500 ;
    END
  END FrameData[28]
  PIN FrameData[290]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1747.640 4.000 1748.240 ;
    END
  END FrameData[290]
  PIN FrameData[291]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1751.040 4.000 1751.640 ;
    END
  END FrameData[291]
  PIN FrameData[292]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1754.440 4.000 1755.040 ;
    END
  END FrameData[292]
  PIN FrameData[293]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1757.840 4.000 1758.440 ;
    END
  END FrameData[293]
  PIN FrameData[294]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1764.640 4.000 1765.240 ;
    END
  END FrameData[294]
  PIN FrameData[295]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1768.040 4.000 1768.640 ;
    END
  END FrameData[295]
  PIN FrameData[296]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1771.440 4.000 1772.040 ;
    END
  END FrameData[296]
  PIN FrameData[297]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1774.840 4.000 1775.440 ;
    END
  END FrameData[297]
  PIN FrameData[298]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1778.240 4.000 1778.840 ;
    END
  END FrameData[298]
  PIN FrameData[299]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1785.040 4.000 1785.640 ;
    END
  END FrameData[299]
  PIN FrameData[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 64.490 3778.500 64.770 3782.500 ;
    END
  END FrameData[29]
  PIN FrameData[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 54.830 3778.500 55.110 3782.500 ;
    END
  END FrameData[2]
  PIN FrameData[300]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1788.440 4.000 1789.040 ;
    END
  END FrameData[300]
  PIN FrameData[301]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1791.840 4.000 1792.440 ;
    END
  END FrameData[301]
  PIN FrameData[302]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1795.240 4.000 1795.840 ;
    END
  END FrameData[302]
  PIN FrameData[303]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1798.640 4.000 1799.240 ;
    END
  END FrameData[303]
  PIN FrameData[304]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1805.440 4.000 1806.040 ;
    END
  END FrameData[304]
  PIN FrameData[305]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1808.840 4.000 1809.440 ;
    END
  END FrameData[305]
  PIN FrameData[306]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1812.240 4.000 1812.840 ;
    END
  END FrameData[306]
  PIN FrameData[307]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1815.640 4.000 1816.240 ;
    END
  END FrameData[307]
  PIN FrameData[308]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1819.040 4.000 1819.640 ;
    END
  END FrameData[308]
  PIN FrameData[309]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1825.840 4.000 1826.440 ;
    END
  END FrameData[309]
  PIN FrameData[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 135.330 3778.500 135.610 3782.500 ;
    END
  END FrameData[30]
  PIN FrameData[310]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1829.240 4.000 1829.840 ;
    END
  END FrameData[310]
  PIN FrameData[311]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1832.640 4.000 1833.240 ;
    END
  END FrameData[311]
  PIN FrameData[312]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1836.040 4.000 1836.640 ;
    END
  END FrameData[312]
  PIN FrameData[313]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1839.440 4.000 1840.040 ;
    END
  END FrameData[313]
  PIN FrameData[314]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1846.240 4.000 1846.840 ;
    END
  END FrameData[314]
  PIN FrameData[315]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1849.640 4.000 1850.240 ;
    END
  END FrameData[315]
  PIN FrameData[316]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1853.040 4.000 1853.640 ;
    END
  END FrameData[316]
  PIN FrameData[317]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1856.440 4.000 1857.040 ;
    END
  END FrameData[317]
  PIN FrameData[318]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1859.840 4.000 1860.440 ;
    END
  END FrameData[318]
  PIN FrameData[319]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1866.640 4.000 1867.240 ;
    END
  END FrameData[319]
  PIN FrameData[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 45.170 3778.500 45.450 3782.500 ;
    END
  END FrameData[31]
  PIN FrameData[320]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1513.040 4.000 1513.640 ;
    END
  END FrameData[320]
  PIN FrameData[321]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1516.440 4.000 1517.040 ;
    END
  END FrameData[321]
  PIN FrameData[322]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1523.240 4.000 1523.840 ;
    END
  END FrameData[322]
  PIN FrameData[323]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1526.640 4.000 1527.240 ;
    END
  END FrameData[323]
  PIN FrameData[324]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1530.040 4.000 1530.640 ;
    END
  END FrameData[324]
  PIN FrameData[325]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1533.440 4.000 1534.040 ;
    END
  END FrameData[325]
  PIN FrameData[326]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1536.840 4.000 1537.440 ;
    END
  END FrameData[326]
  PIN FrameData[327]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1543.640 4.000 1544.240 ;
    END
  END FrameData[327]
  PIN FrameData[328]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1547.040 4.000 1547.640 ;
    END
  END FrameData[328]
  PIN FrameData[329]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1550.440 4.000 1551.040 ;
    END
  END FrameData[329]
  PIN FrameData[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3539.440 4.000 3540.040 ;
    END
  END FrameData[32]
  PIN FrameData[330]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1553.840 4.000 1554.440 ;
    END
  END FrameData[330]
  PIN FrameData[331]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1557.240 4.000 1557.840 ;
    END
  END FrameData[331]
  PIN FrameData[332]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1564.040 4.000 1564.640 ;
    END
  END FrameData[332]
  PIN FrameData[333]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1567.440 4.000 1568.040 ;
    END
  END FrameData[333]
  PIN FrameData[334]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1570.840 4.000 1571.440 ;
    END
  END FrameData[334]
  PIN FrameData[335]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1574.240 4.000 1574.840 ;
    END
  END FrameData[335]
  PIN FrameData[336]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1577.640 4.000 1578.240 ;
    END
  END FrameData[336]
  PIN FrameData[337]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1584.440 4.000 1585.040 ;
    END
  END FrameData[337]
  PIN FrameData[338]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1587.840 4.000 1588.440 ;
    END
  END FrameData[338]
  PIN FrameData[339]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1591.240 4.000 1591.840 ;
    END
  END FrameData[339]
  PIN FrameData[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3542.840 4.000 3543.440 ;
    END
  END FrameData[33]
  PIN FrameData[340]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1594.640 4.000 1595.240 ;
    END
  END FrameData[340]
  PIN FrameData[341]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1598.040 4.000 1598.640 ;
    END
  END FrameData[341]
  PIN FrameData[342]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1604.840 4.000 1605.440 ;
    END
  END FrameData[342]
  PIN FrameData[343]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1608.240 4.000 1608.840 ;
    END
  END FrameData[343]
  PIN FrameData[344]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1611.640 4.000 1612.240 ;
    END
  END FrameData[344]
  PIN FrameData[345]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1615.040 4.000 1615.640 ;
    END
  END FrameData[345]
  PIN FrameData[346]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1618.440 4.000 1619.040 ;
    END
  END FrameData[346]
  PIN FrameData[347]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1625.240 4.000 1625.840 ;
    END
  END FrameData[347]
  PIN FrameData[348]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1628.640 4.000 1629.240 ;
    END
  END FrameData[348]
  PIN FrameData[349]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1632.040 4.000 1632.640 ;
    END
  END FrameData[349]
  PIN FrameData[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3546.240 4.000 3546.840 ;
    END
  END FrameData[34]
  PIN FrameData[350]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1635.440 4.000 1636.040 ;
    END
  END FrameData[350]
  PIN FrameData[351]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1638.840 4.000 1639.440 ;
    END
  END FrameData[351]
  PIN FrameData[352]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1288.640 4.000 1289.240 ;
    END
  END FrameData[352]
  PIN FrameData[353]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1292.040 4.000 1292.640 ;
    END
  END FrameData[353]
  PIN FrameData[354]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1295.440 4.000 1296.040 ;
    END
  END FrameData[354]
  PIN FrameData[355]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1302.240 4.000 1302.840 ;
    END
  END FrameData[355]
  PIN FrameData[356]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1305.640 4.000 1306.240 ;
    END
  END FrameData[356]
  PIN FrameData[357]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1309.040 4.000 1309.640 ;
    END
  END FrameData[357]
  PIN FrameData[358]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1312.440 4.000 1313.040 ;
    END
  END FrameData[358]
  PIN FrameData[359]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1315.840 4.000 1316.440 ;
    END
  END FrameData[359]
  PIN FrameData[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3549.640 4.000 3550.240 ;
    END
  END FrameData[35]
  PIN FrameData[360]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1322.640 4.000 1323.240 ;
    END
  END FrameData[360]
  PIN FrameData[361]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1326.040 4.000 1326.640 ;
    END
  END FrameData[361]
  PIN FrameData[362]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1329.440 4.000 1330.040 ;
    END
  END FrameData[362]
  PIN FrameData[363]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1332.840 4.000 1333.440 ;
    END
  END FrameData[363]
  PIN FrameData[364]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1336.240 4.000 1336.840 ;
    END
  END FrameData[364]
  PIN FrameData[365]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1343.040 4.000 1343.640 ;
    END
  END FrameData[365]
  PIN FrameData[366]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1346.440 4.000 1347.040 ;
    END
  END FrameData[366]
  PIN FrameData[367]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1349.840 4.000 1350.440 ;
    END
  END FrameData[367]
  PIN FrameData[368]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1353.240 4.000 1353.840 ;
    END
  END FrameData[368]
  PIN FrameData[369]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1356.640 4.000 1357.240 ;
    END
  END FrameData[369]
  PIN FrameData[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3556.440 4.000 3557.040 ;
    END
  END FrameData[36]
  PIN FrameData[370]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1363.440 4.000 1364.040 ;
    END
  END FrameData[370]
  PIN FrameData[371]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1366.840 4.000 1367.440 ;
    END
  END FrameData[371]
  PIN FrameData[372]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1370.240 4.000 1370.840 ;
    END
  END FrameData[372]
  PIN FrameData[373]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1373.640 4.000 1374.240 ;
    END
  END FrameData[373]
  PIN FrameData[374]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1377.040 4.000 1377.640 ;
    END
  END FrameData[374]
  PIN FrameData[375]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1383.840 4.000 1384.440 ;
    END
  END FrameData[375]
  PIN FrameData[376]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1387.240 4.000 1387.840 ;
    END
  END FrameData[376]
  PIN FrameData[377]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1390.640 4.000 1391.240 ;
    END
  END FrameData[377]
  PIN FrameData[378]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1394.040 4.000 1394.640 ;
    END
  END FrameData[378]
  PIN FrameData[379]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1397.440 4.000 1398.040 ;
    END
  END FrameData[379]
  PIN FrameData[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3559.840 4.000 3560.440 ;
    END
  END FrameData[37]
  PIN FrameData[380]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1404.240 4.000 1404.840 ;
    END
  END FrameData[380]
  PIN FrameData[381]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1407.640 4.000 1408.240 ;
    END
  END FrameData[381]
  PIN FrameData[382]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1411.040 4.000 1411.640 ;
    END
  END FrameData[382]
  PIN FrameData[383]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1414.440 4.000 1415.040 ;
    END
  END FrameData[383]
  PIN FrameData[384]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1060.840 4.000 1061.440 ;
    END
  END FrameData[384]
  PIN FrameData[385]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1067.640 4.000 1068.240 ;
    END
  END FrameData[385]
  PIN FrameData[386]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1071.040 4.000 1071.640 ;
    END
  END FrameData[386]
  PIN FrameData[387]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1074.440 4.000 1075.040 ;
    END
  END FrameData[387]
  PIN FrameData[388]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1081.240 4.000 1081.840 ;
    END
  END FrameData[388]
  PIN FrameData[389]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1084.640 4.000 1085.240 ;
    END
  END FrameData[389]
  PIN FrameData[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3563.240 4.000 3563.840 ;
    END
  END FrameData[38]
  PIN FrameData[390]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1088.040 4.000 1088.640 ;
    END
  END FrameData[390]
  PIN FrameData[391]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1091.440 4.000 1092.040 ;
    END
  END FrameData[391]
  PIN FrameData[392]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1094.840 4.000 1095.440 ;
    END
  END FrameData[392]
  PIN FrameData[393]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1101.640 4.000 1102.240 ;
    END
  END FrameData[393]
  PIN FrameData[394]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1105.040 4.000 1105.640 ;
    END
  END FrameData[394]
  PIN FrameData[395]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1108.440 4.000 1109.040 ;
    END
  END FrameData[395]
  PIN FrameData[396]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1111.840 4.000 1112.440 ;
    END
  END FrameData[396]
  PIN FrameData[397]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1115.240 4.000 1115.840 ;
    END
  END FrameData[397]
  PIN FrameData[398]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1122.040 4.000 1122.640 ;
    END
  END FrameData[398]
  PIN FrameData[399]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1125.440 4.000 1126.040 ;
    END
  END FrameData[399]
  PIN FrameData[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3566.640 4.000 3567.240 ;
    END
  END FrameData[39]
  PIN FrameData[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 109.570 3778.500 109.850 3782.500 ;
    END
  END FrameData[3]
  PIN FrameData[400]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1128.840 4.000 1129.440 ;
    END
  END FrameData[400]
  PIN FrameData[401]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1132.240 4.000 1132.840 ;
    END
  END FrameData[401]
  PIN FrameData[402]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1135.640 4.000 1136.240 ;
    END
  END FrameData[402]
  PIN FrameData[403]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1142.440 4.000 1143.040 ;
    END
  END FrameData[403]
  PIN FrameData[404]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1145.840 4.000 1146.440 ;
    END
  END FrameData[404]
  PIN FrameData[405]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1149.240 4.000 1149.840 ;
    END
  END FrameData[405]
  PIN FrameData[406]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1152.640 4.000 1153.240 ;
    END
  END FrameData[406]
  PIN FrameData[407]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1156.040 4.000 1156.640 ;
    END
  END FrameData[407]
  PIN FrameData[408]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1162.840 4.000 1163.440 ;
    END
  END FrameData[408]
  PIN FrameData[409]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1166.240 4.000 1166.840 ;
    END
  END FrameData[409]
  PIN FrameData[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3570.040 4.000 3570.640 ;
    END
  END FrameData[40]
  PIN FrameData[410]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1169.640 4.000 1170.240 ;
    END
  END FrameData[410]
  PIN FrameData[411]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1173.040 4.000 1173.640 ;
    END
  END FrameData[411]
  PIN FrameData[412]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1176.440 4.000 1177.040 ;
    END
  END FrameData[412]
  PIN FrameData[413]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1183.240 4.000 1183.840 ;
    END
  END FrameData[413]
  PIN FrameData[414]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1186.640 4.000 1187.240 ;
    END
  END FrameData[414]
  PIN FrameData[415]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1190.040 4.000 1190.640 ;
    END
  END FrameData[415]
  PIN FrameData[416]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 839.840 4.000 840.440 ;
    END
  END FrameData[416]
  PIN FrameData[417]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 843.240 4.000 843.840 ;
    END
  END FrameData[417]
  PIN FrameData[418]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 846.640 4.000 847.240 ;
    END
  END FrameData[418]
  PIN FrameData[419]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 850.040 4.000 850.640 ;
    END
  END FrameData[419]
  PIN FrameData[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3576.840 4.000 3577.440 ;
    END
  END FrameData[41]
  PIN FrameData[420]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 853.440 4.000 854.040 ;
    END
  END FrameData[420]
  PIN FrameData[421]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 860.240 4.000 860.840 ;
    END
  END FrameData[421]
  PIN FrameData[422]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 863.640 4.000 864.240 ;
    END
  END FrameData[422]
  PIN FrameData[423]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 867.040 4.000 867.640 ;
    END
  END FrameData[423]
  PIN FrameData[424]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 870.440 4.000 871.040 ;
    END
  END FrameData[424]
  PIN FrameData[425]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 873.840 4.000 874.440 ;
    END
  END FrameData[425]
  PIN FrameData[426]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 880.640 4.000 881.240 ;
    END
  END FrameData[426]
  PIN FrameData[427]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 884.040 4.000 884.640 ;
    END
  END FrameData[427]
  PIN FrameData[428]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 887.440 4.000 888.040 ;
    END
  END FrameData[428]
  PIN FrameData[429]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 890.840 4.000 891.440 ;
    END
  END FrameData[429]
  PIN FrameData[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3580.240 4.000 3580.840 ;
    END
  END FrameData[42]
  PIN FrameData[430]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 894.240 4.000 894.840 ;
    END
  END FrameData[430]
  PIN FrameData[431]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 901.040 4.000 901.640 ;
    END
  END FrameData[431]
  PIN FrameData[432]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 904.440 4.000 905.040 ;
    END
  END FrameData[432]
  PIN FrameData[433]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 907.840 4.000 908.440 ;
    END
  END FrameData[433]
  PIN FrameData[434]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 911.240 4.000 911.840 ;
    END
  END FrameData[434]
  PIN FrameData[435]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 914.640 4.000 915.240 ;
    END
  END FrameData[435]
  PIN FrameData[436]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 921.440 4.000 922.040 ;
    END
  END FrameData[436]
  PIN FrameData[437]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 924.840 4.000 925.440 ;
    END
  END FrameData[437]
  PIN FrameData[438]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 928.240 4.000 928.840 ;
    END
  END FrameData[438]
  PIN FrameData[439]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 931.640 4.000 932.240 ;
    END
  END FrameData[439]
  PIN FrameData[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3583.640 4.000 3584.240 ;
    END
  END FrameData[43]
  PIN FrameData[440]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 935.040 4.000 935.640 ;
    END
  END FrameData[440]
  PIN FrameData[441]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 941.840 4.000 942.440 ;
    END
  END FrameData[441]
  PIN FrameData[442]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 945.240 4.000 945.840 ;
    END
  END FrameData[442]
  PIN FrameData[443]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 948.640 4.000 949.240 ;
    END
  END FrameData[443]
  PIN FrameData[444]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 952.040 4.000 952.640 ;
    END
  END FrameData[444]
  PIN FrameData[445]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 955.440 4.000 956.040 ;
    END
  END FrameData[445]
  PIN FrameData[446]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 962.240 4.000 962.840 ;
    END
  END FrameData[446]
  PIN FrameData[447]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 965.640 4.000 966.240 ;
    END
  END FrameData[447]
  PIN FrameData[448]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 615.440 4.000 616.040 ;
    END
  END FrameData[448]
  PIN FrameData[449]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 618.840 4.000 619.440 ;
    END
  END FrameData[449]
  PIN FrameData[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3587.040 4.000 3587.640 ;
    END
  END FrameData[44]
  PIN FrameData[450]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 622.240 4.000 622.840 ;
    END
  END FrameData[450]
  PIN FrameData[451]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 625.640 4.000 626.240 ;
    END
  END FrameData[451]
  PIN FrameData[452]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 629.040 4.000 629.640 ;
    END
  END FrameData[452]
  PIN FrameData[453]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 635.840 4.000 636.440 ;
    END
  END FrameData[453]
  PIN FrameData[454]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 639.240 4.000 639.840 ;
    END
  END FrameData[454]
  PIN FrameData[455]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 642.640 4.000 643.240 ;
    END
  END FrameData[455]
  PIN FrameData[456]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 646.040 4.000 646.640 ;
    END
  END FrameData[456]
  PIN FrameData[457]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 649.440 4.000 650.040 ;
    END
  END FrameData[457]
  PIN FrameData[458]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 656.240 4.000 656.840 ;
    END
  END FrameData[458]
  PIN FrameData[459]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 659.640 4.000 660.240 ;
    END
  END FrameData[459]
  PIN FrameData[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3590.440 4.000 3591.040 ;
    END
  END FrameData[45]
  PIN FrameData[460]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 663.040 4.000 663.640 ;
    END
  END FrameData[460]
  PIN FrameData[461]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 666.440 4.000 667.040 ;
    END
  END FrameData[461]
  PIN FrameData[462]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 669.840 4.000 670.440 ;
    END
  END FrameData[462]
  PIN FrameData[463]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 676.640 4.000 677.240 ;
    END
  END FrameData[463]
  PIN FrameData[464]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 680.040 4.000 680.640 ;
    END
  END FrameData[464]
  PIN FrameData[465]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 683.440 4.000 684.040 ;
    END
  END FrameData[465]
  PIN FrameData[466]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 686.840 4.000 687.440 ;
    END
  END FrameData[466]
  PIN FrameData[467]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 690.240 4.000 690.840 ;
    END
  END FrameData[467]
  PIN FrameData[468]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 697.040 4.000 697.640 ;
    END
  END FrameData[468]
  PIN FrameData[469]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 700.440 4.000 701.040 ;
    END
  END FrameData[469]
  PIN FrameData[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3597.240 4.000 3597.840 ;
    END
  END FrameData[46]
  PIN FrameData[470]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 703.840 4.000 704.440 ;
    END
  END FrameData[470]
  PIN FrameData[471]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 707.240 4.000 707.840 ;
    END
  END FrameData[471]
  PIN FrameData[472]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 710.640 4.000 711.240 ;
    END
  END FrameData[472]
  PIN FrameData[473]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 717.440 4.000 718.040 ;
    END
  END FrameData[473]
  PIN FrameData[474]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 720.840 4.000 721.440 ;
    END
  END FrameData[474]
  PIN FrameData[475]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 724.240 4.000 724.840 ;
    END
  END FrameData[475]
  PIN FrameData[476]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 727.640 4.000 728.240 ;
    END
  END FrameData[476]
  PIN FrameData[477]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 731.040 4.000 731.640 ;
    END
  END FrameData[477]
  PIN FrameData[478]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 737.840 4.000 738.440 ;
    END
  END FrameData[478]
  PIN FrameData[479]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 741.240 4.000 741.840 ;
    END
  END FrameData[479]
  PIN FrameData[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3600.640 4.000 3601.240 ;
    END
  END FrameData[47]
  PIN FrameData[480]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 221.040 4.000 221.640 ;
    END
  END FrameData[480]
  PIN FrameData[481]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 302.640 4.000 303.240 ;
    END
  END FrameData[481]
  PIN FrameData[482]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 312.840 4.000 313.440 ;
    END
  END FrameData[482]
  PIN FrameData[483]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 343.440 4.000 344.040 ;
    END
  END FrameData[483]
  PIN FrameData[484]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 370.640 4.000 371.240 ;
    END
  END FrameData[484]
  PIN FrameData[485]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 299.240 4.000 299.840 ;
    END
  END FrameData[485]
  PIN FrameData[486]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 367.240 4.000 367.840 ;
    END
  END FrameData[486]
  PIN FrameData[487]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 295.840 4.000 296.440 ;
    END
  END FrameData[487]
  PIN FrameData[488]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 374.040 4.000 374.640 ;
    END
  END FrameData[488]
  PIN FrameData[489]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 292.440 4.000 293.040 ;
    END
  END FrameData[489]
  PIN FrameData[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3604.040 4.000 3604.640 ;
    END
  END FrameData[48]
  PIN FrameData[490]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 333.240 4.000 333.840 ;
    END
  END FrameData[490]
  PIN FrameData[491]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 363.840 4.000 364.440 ;
    END
  END FrameData[491]
  PIN FrameData[492]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 360.440 4.000 361.040 ;
    END
  END FrameData[492]
  PIN FrameData[493]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 282.240 4.000 282.840 ;
    END
  END FrameData[493]
  PIN FrameData[494]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 377.440 4.000 378.040 ;
    END
  END FrameData[494]
  PIN FrameData[495]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 336.640 4.000 337.240 ;
    END
  END FrameData[495]
  PIN FrameData[496]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 380.840 4.000 381.440 ;
    END
  END FrameData[496]
  PIN FrameData[497]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 459.040 4.000 459.640 ;
    END
  END FrameData[497]
  PIN FrameData[498]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 462.440 4.000 463.040 ;
    END
  END FrameData[498]
  PIN FrameData[499]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 465.840 4.000 466.440 ;
    END
  END FrameData[499]
  PIN FrameData[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3607.440 4.000 3608.040 ;
    END
  END FrameData[49]
  PIN FrameData[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 83.810 3778.500 84.090 3782.500 ;
    END
  END FrameData[4]
  PIN FrameData[500]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 469.240 4.000 469.840 ;
    END
  END FrameData[500]
  PIN FrameData[501]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 476.040 4.000 476.640 ;
    END
  END FrameData[501]
  PIN FrameData[502]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 479.440 4.000 480.040 ;
    END
  END FrameData[502]
  PIN FrameData[503]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 482.840 4.000 483.440 ;
    END
  END FrameData[503]
  PIN FrameData[504]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 486.240 4.000 486.840 ;
    END
  END FrameData[504]
  PIN FrameData[505]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 489.640 4.000 490.240 ;
    END
  END FrameData[505]
  PIN FrameData[506]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 496.440 4.000 497.040 ;
    END
  END FrameData[506]
  PIN FrameData[507]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 499.840 4.000 500.440 ;
    END
  END FrameData[507]
  PIN FrameData[508]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 503.240 4.000 503.840 ;
    END
  END FrameData[508]
  PIN FrameData[509]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 506.640 4.000 507.240 ;
    END
  END FrameData[509]
  PIN FrameData[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3610.840 4.000 3611.440 ;
    END
  END FrameData[50]
  PIN FrameData[510]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 510.040 4.000 510.640 ;
    END
  END FrameData[510]
  PIN FrameData[511]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 516.840 4.000 517.440 ;
    END
  END FrameData[511]
  PIN FrameData[512]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 183.640 4.000 184.240 ;
    END
  END FrameData[512]
  PIN FrameData[513]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 170.040 4.000 170.640 ;
    END
  END FrameData[513]
  PIN FrameData[514]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 173.440 4.000 174.040 ;
    END
  END FrameData[514]
  PIN FrameData[515]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 176.840 4.000 177.440 ;
    END
  END FrameData[515]
  PIN FrameData[516]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 180.240 4.000 180.840 ;
    END
  END FrameData[516]
  PIN FrameData[517]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 187.040 4.000 187.640 ;
    END
  END FrameData[517]
  PIN FrameData[518]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 190.440 4.000 191.040 ;
    END
  END FrameData[518]
  PIN FrameData[519]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 193.840 4.000 194.440 ;
    END
  END FrameData[519]
  PIN FrameData[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3617.640 4.000 3618.240 ;
    END
  END FrameData[51]
  PIN FrameData[520]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 197.240 4.000 197.840 ;
    END
  END FrameData[520]
  PIN FrameData[521]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 200.640 4.000 201.240 ;
    END
  END FrameData[521]
  PIN FrameData[522]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 204.040 4.000 204.640 ;
    END
  END FrameData[522]
  PIN FrameData[523]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 207.440 4.000 208.040 ;
    END
  END FrameData[523]
  PIN FrameData[524]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 210.840 4.000 211.440 ;
    END
  END FrameData[524]
  PIN FrameData[525]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 214.240 4.000 214.840 ;
    END
  END FrameData[525]
  PIN FrameData[526]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 217.640 4.000 218.240 ;
    END
  END FrameData[526]
  PIN FrameData[527]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 224.440 4.000 225.040 ;
    END
  END FrameData[527]
  PIN FrameData[528]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 227.840 4.000 228.440 ;
    END
  END FrameData[528]
  PIN FrameData[529]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 231.240 4.000 231.840 ;
    END
  END FrameData[529]
  PIN FrameData[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3621.040 4.000 3621.640 ;
    END
  END FrameData[52]
  PIN FrameData[530]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 234.640 4.000 235.240 ;
    END
  END FrameData[530]
  PIN FrameData[531]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 238.040 4.000 238.640 ;
    END
  END FrameData[531]
  PIN FrameData[532]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 244.840 4.000 245.440 ;
    END
  END FrameData[532]
  PIN FrameData[533]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 248.240 4.000 248.840 ;
    END
  END FrameData[533]
  PIN FrameData[534]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 251.640 4.000 252.240 ;
    END
  END FrameData[534]
  PIN FrameData[535]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 255.040 4.000 255.640 ;
    END
  END FrameData[535]
  PIN FrameData[536]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 258.440 4.000 259.040 ;
    END
  END FrameData[536]
  PIN FrameData[537]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 265.240 4.000 265.840 ;
    END
  END FrameData[537]
  PIN FrameData[538]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 268.640 4.000 269.240 ;
    END
  END FrameData[538]
  PIN FrameData[539]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 272.040 4.000 272.640 ;
    END
  END FrameData[539]
  PIN FrameData[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3624.440 4.000 3625.040 ;
    END
  END FrameData[53]
  PIN FrameData[540]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 275.440 4.000 276.040 ;
    END
  END FrameData[540]
  PIN FrameData[541]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 278.840 4.000 279.440 ;
    END
  END FrameData[541]
  PIN FrameData[542]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 285.640 4.000 286.240 ;
    END
  END FrameData[542]
  PIN FrameData[543]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 289.040 4.000 289.640 ;
    END
  END FrameData[543]
  PIN FrameData[544]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 112.790 0.000 113.070 4.000 ;
    END
  END FrameData[544]
  PIN FrameData[545]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 106.350 0.000 106.630 4.000 ;
    END
  END FrameData[545]
  PIN FrameData[546]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 103.130 0.000 103.410 4.000 ;
    END
  END FrameData[546]
  PIN FrameData[547]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 109.570 0.000 109.850 4.000 ;
    END
  END FrameData[547]
  PIN FrameData[548]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.840 4.000 24.440 ;
    END
  END FrameData[548]
  PIN FrameData[549]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 37.440 4.000 38.040 ;
    END
  END FrameData[549]
  PIN FrameData[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3627.840 4.000 3628.440 ;
    END
  END FrameData[54]
  PIN FrameData[550]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 0.040 4.000 0.640 ;
    END
  END FrameData[550]
  PIN FrameData[551]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3.440 4.000 4.040 ;
    END
  END FrameData[551]
  PIN FrameData[552]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 4.000 48.240 ;
    END
  END FrameData[552]
  PIN FrameData[553]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.040 4.000 17.640 ;
    END
  END FrameData[553]
  PIN FrameData[554]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 4.000 27.840 ;
    END
  END FrameData[554]
  PIN FrameData[555]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.040 4.000 51.640 ;
    END
  END FrameData[555]
  PIN FrameData[556]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 30.640 4.000 31.240 ;
    END
  END FrameData[556]
  PIN FrameData[557]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 4.000 34.640 ;
    END
  END FrameData[557]
  PIN FrameData[558]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.240 4.000 10.840 ;
    END
  END FrameData[558]
  PIN FrameData[559]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 4.000 55.040 ;
    END
  END FrameData[559]
  PIN FrameData[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3631.240 4.000 3631.840 ;
    END
  END FrameData[55]
  PIN FrameData[560]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 4.000 41.440 ;
    END
  END FrameData[560]
  PIN FrameData[561]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.840 4.000 58.440 ;
    END
  END FrameData[561]
  PIN FrameData[562]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.840 4.000 7.440 ;
    END
  END FrameData[562]
  PIN FrameData[563]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.240 4.000 44.840 ;
    END
  END FrameData[563]
  PIN FrameData[564]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.240 4.000 61.840 ;
    END
  END FrameData[564]
  PIN FrameData[565]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 20.440 4.000 21.040 ;
    END
  END FrameData[565]
  PIN FrameData[566]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 13.640 4.000 14.240 ;
    END
  END FrameData[566]
  PIN FrameData[567]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 64.640 4.000 65.240 ;
    END
  END FrameData[567]
  PIN FrameData[568]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 4.000 68.640 ;
    END
  END FrameData[568]
  PIN FrameData[569]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 71.440 4.000 72.040 ;
    END
  END FrameData[569]
  PIN FrameData[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3638.040 4.000 3638.640 ;
    END
  END FrameData[56]
  PIN FrameData[570]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 166.640 4.000 167.240 ;
    END
  END FrameData[570]
  PIN FrameData[571]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 4.000 75.440 ;
    END
  END FrameData[571]
  PIN FrameData[572]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 163.240 4.000 163.840 ;
    END
  END FrameData[572]
  PIN FrameData[573]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.040 4.000 85.640 ;
    END
  END FrameData[573]
  PIN FrameData[574]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.240 4.000 78.840 ;
    END
  END FrameData[574]
  PIN FrameData[575]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 81.640 4.000 82.240 ;
    END
  END FrameData[575]
  PIN FrameData[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3641.440 4.000 3642.040 ;
    END
  END FrameData[57]
  PIN FrameData[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3644.840 4.000 3645.440 ;
    END
  END FrameData[58]
  PIN FrameData[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3648.240 4.000 3648.840 ;
    END
  END FrameData[59]
  PIN FrameData[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 128.890 3778.500 129.170 3782.500 ;
    END
  END FrameData[5]
  PIN FrameData[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3651.640 4.000 3652.240 ;
    END
  END FrameData[60]
  PIN FrameData[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3658.440 4.000 3659.040 ;
    END
  END FrameData[61]
  PIN FrameData[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3661.840 4.000 3662.440 ;
    END
  END FrameData[62]
  PIN FrameData[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3665.240 4.000 3665.840 ;
    END
  END FrameData[63]
  PIN FrameData[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3315.040 4.000 3315.640 ;
    END
  END FrameData[64]
  PIN FrameData[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3318.440 4.000 3319.040 ;
    END
  END FrameData[65]
  PIN FrameData[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3321.840 4.000 3322.440 ;
    END
  END FrameData[66]
  PIN FrameData[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3325.240 4.000 3325.840 ;
    END
  END FrameData[67]
  PIN FrameData[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3328.640 4.000 3329.240 ;
    END
  END FrameData[68]
  PIN FrameData[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3335.440 4.000 3336.040 ;
    END
  END FrameData[69]
  PIN FrameData[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 173.970 3778.500 174.250 3782.500 ;
    END
  END FrameData[6]
  PIN FrameData[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3338.840 4.000 3339.440 ;
    END
  END FrameData[70]
  PIN FrameData[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3342.240 4.000 3342.840 ;
    END
  END FrameData[71]
  PIN FrameData[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3345.640 4.000 3346.240 ;
    END
  END FrameData[72]
  PIN FrameData[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3349.040 4.000 3349.640 ;
    END
  END FrameData[73]
  PIN FrameData[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3355.840 4.000 3356.440 ;
    END
  END FrameData[74]
  PIN FrameData[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3359.240 4.000 3359.840 ;
    END
  END FrameData[75]
  PIN FrameData[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3362.640 4.000 3363.240 ;
    END
  END FrameData[76]
  PIN FrameData[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3366.040 4.000 3366.640 ;
    END
  END FrameData[77]
  PIN FrameData[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3369.440 4.000 3370.040 ;
    END
  END FrameData[78]
  PIN FrameData[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3376.240 4.000 3376.840 ;
    END
  END FrameData[79]
  PIN FrameData[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 80.590 3778.500 80.870 3782.500 ;
    END
  END FrameData[7]
  PIN FrameData[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3379.640 4.000 3380.240 ;
    END
  END FrameData[80]
  PIN FrameData[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3383.040 4.000 3383.640 ;
    END
  END FrameData[81]
  PIN FrameData[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3386.440 4.000 3387.040 ;
    END
  END FrameData[82]
  PIN FrameData[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3389.840 4.000 3390.440 ;
    END
  END FrameData[83]
  PIN FrameData[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3396.640 4.000 3397.240 ;
    END
  END FrameData[84]
  PIN FrameData[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3400.040 4.000 3400.640 ;
    END
  END FrameData[85]
  PIN FrameData[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3403.440 4.000 3404.040 ;
    END
  END FrameData[86]
  PIN FrameData[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3406.840 4.000 3407.440 ;
    END
  END FrameData[87]
  PIN FrameData[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3410.240 4.000 3410.840 ;
    END
  END FrameData[88]
  PIN FrameData[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3417.040 4.000 3417.640 ;
    END
  END FrameData[89]
  PIN FrameData[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 151.430 3778.500 151.710 3782.500 ;
    END
  END FrameData[8]
  PIN FrameData[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3420.440 4.000 3421.040 ;
    END
  END FrameData[90]
  PIN FrameData[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3423.840 4.000 3424.440 ;
    END
  END FrameData[91]
  PIN FrameData[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3427.240 4.000 3427.840 ;
    END
  END FrameData[92]
  PIN FrameData[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3430.640 4.000 3431.240 ;
    END
  END FrameData[93]
  PIN FrameData[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3437.440 4.000 3438.040 ;
    END
  END FrameData[94]
  PIN FrameData[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3440.840 4.000 3441.440 ;
    END
  END FrameData[95]
  PIN FrameData[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3087.240 4.000 3087.840 ;
    END
  END FrameData[96]
  PIN FrameData[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3094.040 4.000 3094.640 ;
    END
  END FrameData[97]
  PIN FrameData[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3097.440 4.000 3098.040 ;
    END
  END FrameData[98]
  PIN FrameData[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3100.840 4.000 3101.440 ;
    END
  END FrameData[99]
  PIN FrameData[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 167.530 3778.500 167.810 3782.500 ;
    END
  END FrameData[9]
  PIN FrameStrobe[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.409500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 159.840 4.000 160.440 ;
    END
  END FrameStrobe[0]
  PIN FrameStrobe[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 1094.890 0.000 1095.170 4.000 ;
    END
  END FrameStrobe[100]
  PIN FrameStrobe[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 1098.110 0.000 1098.390 4.000 ;
    END
  END FrameStrobe[101]
  PIN FrameStrobe[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 1101.330 0.000 1101.610 4.000 ;
    END
  END FrameStrobe[102]
  PIN FrameStrobe[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1104.550 0.000 1104.830 4.000 ;
    END
  END FrameStrobe[103]
  PIN FrameStrobe[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1107.770 0.000 1108.050 4.000 ;
    END
  END FrameStrobe[104]
  PIN FrameStrobe[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1114.210 0.000 1114.490 4.000 ;
    END
  END FrameStrobe[105]
  PIN FrameStrobe[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1117.430 0.000 1117.710 4.000 ;
    END
  END FrameStrobe[106]
  PIN FrameStrobe[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1120.650 0.000 1120.930 4.000 ;
    END
  END FrameStrobe[107]
  PIN FrameStrobe[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1123.870 0.000 1124.150 4.000 ;
    END
  END FrameStrobe[108]
  PIN FrameStrobe[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1127.090 0.000 1127.370 4.000 ;
    END
  END FrameStrobe[109]
  PIN FrameStrobe[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 125.840 4.000 126.440 ;
    END
  END FrameStrobe[10]
  PIN FrameStrobe[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1130.310 0.000 1130.590 4.000 ;
    END
  END FrameStrobe[110]
  PIN FrameStrobe[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1133.530 0.000 1133.810 4.000 ;
    END
  END FrameStrobe[111]
  PIN FrameStrobe[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1139.970 0.000 1140.250 4.000 ;
    END
  END FrameStrobe[112]
  PIN FrameStrobe[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1143.190 0.000 1143.470 4.000 ;
    END
  END FrameStrobe[113]
  PIN FrameStrobe[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1146.410 0.000 1146.690 4.000 ;
    END
  END FrameStrobe[114]
  PIN FrameStrobe[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1149.630 0.000 1149.910 4.000 ;
    END
  END FrameStrobe[115]
  PIN FrameStrobe[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1152.850 0.000 1153.130 4.000 ;
    END
  END FrameStrobe[116]
  PIN FrameStrobe[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1156.070 0.000 1156.350 4.000 ;
    END
  END FrameStrobe[117]
  PIN FrameStrobe[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1159.290 0.000 1159.570 4.000 ;
    END
  END FrameStrobe[118]
  PIN FrameStrobe[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1165.730 0.000 1166.010 4.000 ;
    END
  END FrameStrobe[119]
  PIN FrameStrobe[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 156.440 4.000 157.040 ;
    END
  END FrameStrobe[11]
  PIN FrameStrobe[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 1297.750 0.000 1298.030 4.000 ;
    END
  END FrameStrobe[120]
  PIN FrameStrobe[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 1304.190 0.000 1304.470 4.000 ;
    END
  END FrameStrobe[121]
  PIN FrameStrobe[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 1307.410 0.000 1307.690 4.000 ;
    END
  END FrameStrobe[122]
  PIN FrameStrobe[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1310.630 0.000 1310.910 4.000 ;
    END
  END FrameStrobe[123]
  PIN FrameStrobe[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1313.850 0.000 1314.130 4.000 ;
    END
  END FrameStrobe[124]
  PIN FrameStrobe[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1317.070 0.000 1317.350 4.000 ;
    END
  END FrameStrobe[125]
  PIN FrameStrobe[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1320.290 0.000 1320.570 4.000 ;
    END
  END FrameStrobe[126]
  PIN FrameStrobe[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1323.510 0.000 1323.790 4.000 ;
    END
  END FrameStrobe[127]
  PIN FrameStrobe[128]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1329.950 0.000 1330.230 4.000 ;
    END
  END FrameStrobe[128]
  PIN FrameStrobe[129]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1333.170 0.000 1333.450 4.000 ;
    END
  END FrameStrobe[129]
  PIN FrameStrobe[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.240 4.000 95.840 ;
    END
  END FrameStrobe[12]
  PIN FrameStrobe[130]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1336.390 0.000 1336.670 4.000 ;
    END
  END FrameStrobe[130]
  PIN FrameStrobe[131]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1339.610 0.000 1339.890 4.000 ;
    END
  END FrameStrobe[131]
  PIN FrameStrobe[132]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1342.830 0.000 1343.110 4.000 ;
    END
  END FrameStrobe[132]
  PIN FrameStrobe[133]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1346.050 0.000 1346.330 4.000 ;
    END
  END FrameStrobe[133]
  PIN FrameStrobe[134]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1349.270 0.000 1349.550 4.000 ;
    END
  END FrameStrobe[134]
  PIN FrameStrobe[135]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1355.710 0.000 1355.990 4.000 ;
    END
  END FrameStrobe[135]
  PIN FrameStrobe[136]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1358.930 0.000 1359.210 4.000 ;
    END
  END FrameStrobe[136]
  PIN FrameStrobe[137]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1362.150 0.000 1362.430 4.000 ;
    END
  END FrameStrobe[137]
  PIN FrameStrobe[138]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1365.370 0.000 1365.650 4.000 ;
    END
  END FrameStrobe[138]
  PIN FrameStrobe[139]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1368.590 0.000 1368.870 4.000 ;
    END
  END FrameStrobe[139]
  PIN FrameStrobe[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 102.040 4.000 102.640 ;
    END
  END FrameStrobe[13]
  PIN FrameStrobe[140]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1394.350 0.000 1394.630 4.000 ;
    END
  END FrameStrobe[140]
  PIN FrameStrobe[141]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1404.010 0.000 1404.290 4.000 ;
    END
  END FrameStrobe[141]
  PIN FrameStrobe[142]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1413.670 0.000 1413.950 4.000 ;
    END
  END FrameStrobe[142]
  PIN FrameStrobe[143]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1426.550 0.000 1426.830 4.000 ;
    END
  END FrameStrobe[143]
  PIN FrameStrobe[144]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1436.210 0.000 1436.490 4.000 ;
    END
  END FrameStrobe[144]
  PIN FrameStrobe[145]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1445.870 0.000 1446.150 4.000 ;
    END
  END FrameStrobe[145]
  PIN FrameStrobe[146]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1455.530 0.000 1455.810 4.000 ;
    END
  END FrameStrobe[146]
  PIN FrameStrobe[147]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1468.410 0.000 1468.690 4.000 ;
    END
  END FrameStrobe[147]
  PIN FrameStrobe[148]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1478.070 0.000 1478.350 4.000 ;
    END
  END FrameStrobe[148]
  PIN FrameStrobe[149]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1487.730 0.000 1488.010 4.000 ;
    END
  END FrameStrobe[149]
  PIN FrameStrobe[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 105.440 4.000 106.040 ;
    END
  END FrameStrobe[14]
  PIN FrameStrobe[150]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1500.610 0.000 1500.890 4.000 ;
    END
  END FrameStrobe[150]
  PIN FrameStrobe[151]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1510.270 0.000 1510.550 4.000 ;
    END
  END FrameStrobe[151]
  PIN FrameStrobe[152]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1519.930 0.000 1520.210 4.000 ;
    END
  END FrameStrobe[152]
  PIN FrameStrobe[153]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1529.590 0.000 1529.870 4.000 ;
    END
  END FrameStrobe[153]
  PIN FrameStrobe[154]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1542.470 0.000 1542.750 4.000 ;
    END
  END FrameStrobe[154]
  PIN FrameStrobe[155]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1552.130 0.000 1552.410 4.000 ;
    END
  END FrameStrobe[155]
  PIN FrameStrobe[156]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1561.790 0.000 1562.070 4.000 ;
    END
  END FrameStrobe[156]
  PIN FrameStrobe[157]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1574.670 0.000 1574.950 4.000 ;
    END
  END FrameStrobe[157]
  PIN FrameStrobe[158]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1584.330 0.000 1584.610 4.000 ;
    END
  END FrameStrobe[158]
  PIN FrameStrobe[159]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1593.990 0.000 1594.270 4.000 ;
    END
  END FrameStrobe[159]
  PIN FrameStrobe[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 132.640 4.000 133.240 ;
    END
  END FrameStrobe[15]
  PIN FrameStrobe[160]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 1729.230 0.000 1729.510 4.000 ;
    END
  END FrameStrobe[160]
  PIN FrameStrobe[161]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 1732.450 0.000 1732.730 4.000 ;
    END
  END FrameStrobe[161]
  PIN FrameStrobe[162]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 1735.670 0.000 1735.950 4.000 ;
    END
  END FrameStrobe[162]
  PIN FrameStrobe[163]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1738.890 0.000 1739.170 4.000 ;
    END
  END FrameStrobe[163]
  PIN FrameStrobe[164]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1745.330 0.000 1745.610 4.000 ;
    END
  END FrameStrobe[164]
  PIN FrameStrobe[165]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1748.550 0.000 1748.830 4.000 ;
    END
  END FrameStrobe[165]
  PIN FrameStrobe[166]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1751.770 0.000 1752.050 4.000 ;
    END
  END FrameStrobe[166]
  PIN FrameStrobe[167]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1754.990 0.000 1755.270 4.000 ;
    END
  END FrameStrobe[167]
  PIN FrameStrobe[168]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1758.210 0.000 1758.490 4.000 ;
    END
  END FrameStrobe[168]
  PIN FrameStrobe[169]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1761.430 0.000 1761.710 4.000 ;
    END
  END FrameStrobe[169]
  PIN FrameStrobe[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.240 4.000 112.840 ;
    END
  END FrameStrobe[16]
  PIN FrameStrobe[170]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1764.650 0.000 1764.930 4.000 ;
    END
  END FrameStrobe[170]
  PIN FrameStrobe[171]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1771.090 0.000 1771.370 4.000 ;
    END
  END FrameStrobe[171]
  PIN FrameStrobe[172]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1774.310 0.000 1774.590 4.000 ;
    END
  END FrameStrobe[172]
  PIN FrameStrobe[173]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1777.530 0.000 1777.810 4.000 ;
    END
  END FrameStrobe[173]
  PIN FrameStrobe[174]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1780.750 0.000 1781.030 4.000 ;
    END
  END FrameStrobe[174]
  PIN FrameStrobe[175]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1783.970 0.000 1784.250 4.000 ;
    END
  END FrameStrobe[175]
  PIN FrameStrobe[176]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1787.190 0.000 1787.470 4.000 ;
    END
  END FrameStrobe[176]
  PIN FrameStrobe[177]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1790.410 0.000 1790.690 4.000 ;
    END
  END FrameStrobe[177]
  PIN FrameStrobe[178]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1796.850 0.000 1797.130 4.000 ;
    END
  END FrameStrobe[178]
  PIN FrameStrobe[179]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1800.070 0.000 1800.350 4.000 ;
    END
  END FrameStrobe[179]
  PIN FrameStrobe[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 139.440 4.000 140.040 ;
    END
  END FrameStrobe[17]
  PIN FrameStrobe[180]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.568500 ;
    PORT
      LAYER met2 ;
        RECT 1970.730 0.000 1971.010 4.000 ;
    END
  END FrameStrobe[180]
  PIN FrameStrobe[181]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1935.310 0.000 1935.590 4.000 ;
    END
  END FrameStrobe[181]
  PIN FrameStrobe[182]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1941.750 0.000 1942.030 4.000 ;
    END
  END FrameStrobe[182]
  PIN FrameStrobe[183]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1964.290 0.000 1964.570 4.000 ;
    END
  END FrameStrobe[183]
  PIN FrameStrobe[184]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1938.530 0.000 1938.810 4.000 ;
    END
  END FrameStrobe[184]
  PIN FrameStrobe[185]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1932.090 0.000 1932.370 4.000 ;
    END
  END FrameStrobe[185]
  PIN FrameStrobe[186]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1954.630 0.000 1954.910 4.000 ;
    END
  END FrameStrobe[186]
  PIN FrameStrobe[187]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1944.970 0.000 1945.250 4.000 ;
    END
  END FrameStrobe[187]
  PIN FrameStrobe[188]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1948.190 0.000 1948.470 4.000 ;
    END
  END FrameStrobe[188]
  PIN FrameStrobe[189]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1951.410 0.000 1951.690 4.000 ;
    END
  END FrameStrobe[189]
  PIN FrameStrobe[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 142.840 4.000 143.440 ;
    END
  END FrameStrobe[18]
  PIN FrameStrobe[190]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1957.850 0.000 1958.130 4.000 ;
    END
  END FrameStrobe[190]
  PIN FrameStrobe[191]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1961.070 0.000 1961.350 4.000 ;
    END
  END FrameStrobe[191]
  PIN FrameStrobe[192]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1967.510 0.000 1967.790 4.000 ;
    END
  END FrameStrobe[192]
  PIN FrameStrobe[193]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1973.950 0.000 1974.230 4.000 ;
    END
  END FrameStrobe[193]
  PIN FrameStrobe[194]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1977.170 0.000 1977.450 4.000 ;
    END
  END FrameStrobe[194]
  PIN FrameStrobe[195]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1983.610 0.000 1983.890 4.000 ;
    END
  END FrameStrobe[195]
  PIN FrameStrobe[196]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1990.050 0.000 1990.330 4.000 ;
    END
  END FrameStrobe[196]
  PIN FrameStrobe[197]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1993.270 0.000 1993.550 4.000 ;
    END
  END FrameStrobe[197]
  PIN FrameStrobe[198]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1999.710 0.000 1999.990 4.000 ;
    END
  END FrameStrobe[198]
  PIN FrameStrobe[199]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 2006.150 0.000 2006.430 4.000 ;
    END
  END FrameStrobe[199]
  PIN FrameStrobe[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 149.640 4.000 150.240 ;
    END
  END FrameStrobe[19]
  PIN FrameStrobe[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 146.240 4.000 146.840 ;
    END
  END FrameStrobe[1]
  PIN FrameStrobe[200]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 2080.210 0.000 2080.490 4.000 ;
    END
  END FrameStrobe[200]
  PIN FrameStrobe[201]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.339000 ;
    PORT
      LAYER met2 ;
        RECT 2086.650 0.000 2086.930 4.000 ;
    END
  END FrameStrobe[201]
  PIN FrameStrobe[202]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 2093.090 0.000 2093.370 4.000 ;
    END
  END FrameStrobe[202]
  PIN FrameStrobe[203]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 2099.530 0.000 2099.810 4.000 ;
    END
  END FrameStrobe[203]
  PIN FrameStrobe[204]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 2105.970 0.000 2106.250 4.000 ;
    END
  END FrameStrobe[204]
  PIN FrameStrobe[205]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 2112.410 0.000 2112.690 4.000 ;
    END
  END FrameStrobe[205]
  PIN FrameStrobe[206]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 2118.850 0.000 2119.130 4.000 ;
    END
  END FrameStrobe[206]
  PIN FrameStrobe[207]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 2128.510 0.000 2128.790 4.000 ;
    END
  END FrameStrobe[207]
  PIN FrameStrobe[208]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 2134.950 0.000 2135.230 4.000 ;
    END
  END FrameStrobe[208]
  PIN FrameStrobe[209]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 2141.390 0.000 2141.670 4.000 ;
    END
  END FrameStrobe[209]
  PIN FrameStrobe[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 154.650 0.000 154.930 4.000 ;
    END
  END FrameStrobe[20]
  PIN FrameStrobe[210]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 2147.830 0.000 2148.110 4.000 ;
    END
  END FrameStrobe[210]
  PIN FrameStrobe[211]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 2154.270 0.000 2154.550 4.000 ;
    END
  END FrameStrobe[211]
  PIN FrameStrobe[212]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 2160.710 0.000 2160.990 4.000 ;
    END
  END FrameStrobe[212]
  PIN FrameStrobe[213]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 2167.150 0.000 2167.430 4.000 ;
    END
  END FrameStrobe[213]
  PIN FrameStrobe[214]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 2176.810 0.000 2177.090 4.000 ;
    END
  END FrameStrobe[214]
  PIN FrameStrobe[215]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 2183.250 0.000 2183.530 4.000 ;
    END
  END FrameStrobe[215]
  PIN FrameStrobe[216]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 2189.690 0.000 2189.970 4.000 ;
    END
  END FrameStrobe[216]
  PIN FrameStrobe[217]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 2196.130 0.000 2196.410 4.000 ;
    END
  END FrameStrobe[217]
  PIN FrameStrobe[218]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 2202.570 0.000 2202.850 4.000 ;
    END
  END FrameStrobe[218]
  PIN FrameStrobe[219]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 2209.010 0.000 2209.290 4.000 ;
    END
  END FrameStrobe[219]
  PIN FrameStrobe[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 161.090 0.000 161.370 4.000 ;
    END
  END FrameStrobe[21]
  PIN FrameStrobe[220]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 2231.550 0.000 2231.830 4.000 ;
    END
  END FrameStrobe[220]
  PIN FrameStrobe[221]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 2237.990 0.000 2238.270 4.000 ;
    END
  END FrameStrobe[221]
  PIN FrameStrobe[222]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 2244.430 0.000 2244.710 4.000 ;
    END
  END FrameStrobe[222]
  PIN FrameStrobe[223]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 2254.090 0.000 2254.370 4.000 ;
    END
  END FrameStrobe[223]
  PIN FrameStrobe[224]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 2260.530 0.000 2260.810 4.000 ;
    END
  END FrameStrobe[224]
  PIN FrameStrobe[225]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 2270.190 0.000 2270.470 4.000 ;
    END
  END FrameStrobe[225]
  PIN FrameStrobe[226]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 2276.630 0.000 2276.910 4.000 ;
    END
  END FrameStrobe[226]
  PIN FrameStrobe[227]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 2286.290 0.000 2286.570 4.000 ;
    END
  END FrameStrobe[227]
  PIN FrameStrobe[228]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 2292.730 0.000 2293.010 4.000 ;
    END
  END FrameStrobe[228]
  PIN FrameStrobe[229]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 2299.170 0.000 2299.450 4.000 ;
    END
  END FrameStrobe[229]
  PIN FrameStrobe[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 170.750 0.000 171.030 4.000 ;
    END
  END FrameStrobe[22]
  PIN FrameStrobe[230]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 2308.830 0.000 2309.110 4.000 ;
    END
  END FrameStrobe[230]
  PIN FrameStrobe[231]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 2315.270 0.000 2315.550 4.000 ;
    END
  END FrameStrobe[231]
  PIN FrameStrobe[232]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 2324.930 0.000 2325.210 4.000 ;
    END
  END FrameStrobe[232]
  PIN FrameStrobe[233]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 2331.370 0.000 2331.650 4.000 ;
    END
  END FrameStrobe[233]
  PIN FrameStrobe[234]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 2341.030 0.000 2341.310 4.000 ;
    END
  END FrameStrobe[234]
  PIN FrameStrobe[235]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 2347.470 0.000 2347.750 4.000 ;
    END
  END FrameStrobe[235]
  PIN FrameStrobe[236]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 2353.910 0.000 2354.190 4.000 ;
    END
  END FrameStrobe[236]
  PIN FrameStrobe[237]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 2363.570 0.000 2363.850 4.000 ;
    END
  END FrameStrobe[237]
  PIN FrameStrobe[238]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 2370.010 0.000 2370.290 4.000 ;
    END
  END FrameStrobe[238]
  PIN FrameStrobe[239]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 2379.670 0.000 2379.950 4.000 ;
    END
  END FrameStrobe[239]
  PIN FrameStrobe[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 177.190 0.000 177.470 4.000 ;
    END
  END FrameStrobe[23]
  PIN FrameStrobe[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 183.630 0.000 183.910 4.000 ;
    END
  END FrameStrobe[24]
  PIN FrameStrobe[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 193.290 0.000 193.570 4.000 ;
    END
  END FrameStrobe[25]
  PIN FrameStrobe[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 199.730 0.000 200.010 4.000 ;
    END
  END FrameStrobe[26]
  PIN FrameStrobe[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 209.390 0.000 209.670 4.000 ;
    END
  END FrameStrobe[27]
  PIN FrameStrobe[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 215.830 0.000 216.110 4.000 ;
    END
  END FrameStrobe[28]
  PIN FrameStrobe[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 225.490 0.000 225.770 4.000 ;
    END
  END FrameStrobe[29]
  PIN FrameStrobe[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 98.640 4.000 99.240 ;
    END
  END FrameStrobe[2]
  PIN FrameStrobe[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 231.930 0.000 232.210 4.000 ;
    END
  END FrameStrobe[30]
  PIN FrameStrobe[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 238.370 0.000 238.650 4.000 ;
    END
  END FrameStrobe[31]
  PIN FrameStrobe[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 248.030 0.000 248.310 4.000 ;
    END
  END FrameStrobe[32]
  PIN FrameStrobe[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 254.470 0.000 254.750 4.000 ;
    END
  END FrameStrobe[33]
  PIN FrameStrobe[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 264.130 0.000 264.410 4.000 ;
    END
  END FrameStrobe[34]
  PIN FrameStrobe[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 270.570 0.000 270.850 4.000 ;
    END
  END FrameStrobe[35]
  PIN FrameStrobe[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 280.230 0.000 280.510 4.000 ;
    END
  END FrameStrobe[36]
  PIN FrameStrobe[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 286.670 0.000 286.950 4.000 ;
    END
  END FrameStrobe[37]
  PIN FrameStrobe[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 293.110 0.000 293.390 4.000 ;
    END
  END FrameStrobe[38]
  PIN FrameStrobe[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 302.770 0.000 303.050 4.000 ;
    END
  END FrameStrobe[39]
  PIN FrameStrobe[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.840 4.000 92.440 ;
    END
  END FrameStrobe[3]
  PIN FrameStrobe[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 370.390 0.000 370.670 4.000 ;
    END
  END FrameStrobe[40]
  PIN FrameStrobe[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 376.830 0.000 377.110 4.000 ;
    END
  END FrameStrobe[41]
  PIN FrameStrobe[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 383.270 0.000 383.550 4.000 ;
    END
  END FrameStrobe[42]
  PIN FrameStrobe[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 392.930 0.000 393.210 4.000 ;
    END
  END FrameStrobe[43]
  PIN FrameStrobe[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 399.370 0.000 399.650 4.000 ;
    END
  END FrameStrobe[44]
  PIN FrameStrobe[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 405.810 0.000 406.090 4.000 ;
    END
  END FrameStrobe[45]
  PIN FrameStrobe[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 412.250 0.000 412.530 4.000 ;
    END
  END FrameStrobe[46]
  PIN FrameStrobe[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 421.910 0.000 422.190 4.000 ;
    END
  END FrameStrobe[47]
  PIN FrameStrobe[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 428.350 0.000 428.630 4.000 ;
    END
  END FrameStrobe[48]
  PIN FrameStrobe[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 434.790 0.000 435.070 4.000 ;
    END
  END FrameStrobe[49]
  PIN FrameStrobe[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.440 4.000 89.040 ;
    END
  END FrameStrobe[4]
  PIN FrameStrobe[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 444.450 0.000 444.730 4.000 ;
    END
  END FrameStrobe[50]
  PIN FrameStrobe[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 450.890 0.000 451.170 4.000 ;
    END
  END FrameStrobe[51]
  PIN FrameStrobe[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 457.330 0.000 457.610 4.000 ;
    END
  END FrameStrobe[52]
  PIN FrameStrobe[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 463.770 0.000 464.050 4.000 ;
    END
  END FrameStrobe[53]
  PIN FrameStrobe[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 473.430 0.000 473.710 4.000 ;
    END
  END FrameStrobe[54]
  PIN FrameStrobe[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 479.870 0.000 480.150 4.000 ;
    END
  END FrameStrobe[55]
  PIN FrameStrobe[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 486.310 0.000 486.590 4.000 ;
    END
  END FrameStrobe[56]
  PIN FrameStrobe[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 495.970 0.000 496.250 4.000 ;
    END
  END FrameStrobe[57]
  PIN FrameStrobe[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 502.410 0.000 502.690 4.000 ;
    END
  END FrameStrobe[58]
  PIN FrameStrobe[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 508.850 0.000 509.130 4.000 ;
    END
  END FrameStrobe[59]
  PIN FrameStrobe[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.240 4.000 129.840 ;
    END
  END FrameStrobe[5]
  PIN FrameStrobe[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 534.610 0.000 534.890 4.000 ;
    END
  END FrameStrobe[60]
  PIN FrameStrobe[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 547.490 0.000 547.770 4.000 ;
    END
  END FrameStrobe[61]
  PIN FrameStrobe[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 557.150 0.000 557.430 4.000 ;
    END
  END FrameStrobe[62]
  PIN FrameStrobe[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 570.030 0.000 570.310 4.000 ;
    END
  END FrameStrobe[63]
  PIN FrameStrobe[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 579.690 0.000 579.970 4.000 ;
    END
  END FrameStrobe[64]
  PIN FrameStrobe[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 592.570 0.000 592.850 4.000 ;
    END
  END FrameStrobe[65]
  PIN FrameStrobe[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 602.230 0.000 602.510 4.000 ;
    END
  END FrameStrobe[66]
  PIN FrameStrobe[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 615.110 0.000 615.390 4.000 ;
    END
  END FrameStrobe[67]
  PIN FrameStrobe[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 627.990 0.000 628.270 4.000 ;
    END
  END FrameStrobe[68]
  PIN FrameStrobe[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 637.650 0.000 637.930 4.000 ;
    END
  END FrameStrobe[69]
  PIN FrameStrobe[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 115.640 4.000 116.240 ;
    END
  END FrameStrobe[6]
  PIN FrameStrobe[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 650.530 0.000 650.810 4.000 ;
    END
  END FrameStrobe[70]
  PIN FrameStrobe[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 660.190 0.000 660.470 4.000 ;
    END
  END FrameStrobe[71]
  PIN FrameStrobe[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 673.070 0.000 673.350 4.000 ;
    END
  END FrameStrobe[72]
  PIN FrameStrobe[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 682.730 0.000 683.010 4.000 ;
    END
  END FrameStrobe[73]
  PIN FrameStrobe[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 695.610 0.000 695.890 4.000 ;
    END
  END FrameStrobe[74]
  PIN FrameStrobe[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 708.490 0.000 708.770 4.000 ;
    END
  END FrameStrobe[75]
  PIN FrameStrobe[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 718.150 0.000 718.430 4.000 ;
    END
  END FrameStrobe[76]
  PIN FrameStrobe[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 731.030 0.000 731.310 4.000 ;
    END
  END FrameStrobe[77]
  PIN FrameStrobe[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 740.690 0.000 740.970 4.000 ;
    END
  END FrameStrobe[78]
  PIN FrameStrobe[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 753.570 0.000 753.850 4.000 ;
    END
  END FrameStrobe[79]
  PIN FrameStrobe[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.065900 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 0.000 153.040 4.000 153.640 ;
    END
  END FrameStrobe[7]
  PIN FrameStrobe[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 888.810 0.000 889.090 4.000 ;
    END
  END FrameStrobe[80]
  PIN FrameStrobe[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 892.030 0.000 892.310 4.000 ;
    END
  END FrameStrobe[81]
  PIN FrameStrobe[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 895.250 0.000 895.530 4.000 ;
    END
  END FrameStrobe[82]
  PIN FrameStrobe[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 901.690 0.000 901.970 4.000 ;
    END
  END FrameStrobe[83]
  PIN FrameStrobe[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 904.910 0.000 905.190 4.000 ;
    END
  END FrameStrobe[84]
  PIN FrameStrobe[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 908.130 0.000 908.410 4.000 ;
    END
  END FrameStrobe[85]
  PIN FrameStrobe[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 911.350 0.000 911.630 4.000 ;
    END
  END FrameStrobe[86]
  PIN FrameStrobe[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 914.570 0.000 914.850 4.000 ;
    END
  END FrameStrobe[87]
  PIN FrameStrobe[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 917.790 0.000 918.070 4.000 ;
    END
  END FrameStrobe[88]
  PIN FrameStrobe[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 921.010 0.000 921.290 4.000 ;
    END
  END FrameStrobe[89]
  PIN FrameStrobe[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 136.040 4.000 136.640 ;
    END
  END FrameStrobe[8]
  PIN FrameStrobe[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 927.450 0.000 927.730 4.000 ;
    END
  END FrameStrobe[90]
  PIN FrameStrobe[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 930.670 0.000 930.950 4.000 ;
    END
  END FrameStrobe[91]
  PIN FrameStrobe[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 933.890 0.000 934.170 4.000 ;
    END
  END FrameStrobe[92]
  PIN FrameStrobe[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 937.110 0.000 937.390 4.000 ;
    END
  END FrameStrobe[93]
  PIN FrameStrobe[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 940.330 0.000 940.610 4.000 ;
    END
  END FrameStrobe[94]
  PIN FrameStrobe[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 943.550 0.000 943.830 4.000 ;
    END
  END FrameStrobe[95]
  PIN FrameStrobe[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 946.770 0.000 947.050 4.000 ;
    END
  END FrameStrobe[96]
  PIN FrameStrobe[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 953.210 0.000 953.490 4.000 ;
    END
  END FrameStrobe[97]
  PIN FrameStrobe[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 956.430 0.000 956.710 4.000 ;
    END
  END FrameStrobe[98]
  PIN FrameStrobe[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 959.650 0.000 959.930 4.000 ;
    END
  END FrameStrobe[99]
  PIN FrameStrobe[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.040 4.000 119.640 ;
    END
  END FrameStrobe[9]
  PIN Tile_X0Y10_A_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1462.040 4.000 1462.640 ;
    END
  END Tile_X0Y10_A_I_top
  PIN Tile_X0Y10_A_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1455.240 4.000 1455.840 ;
    END
  END Tile_X0Y10_A_O_top
  PIN Tile_X0Y10_A_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1465.440 4.000 1466.040 ;
    END
  END Tile_X0Y10_A_T_top
  PIN Tile_X0Y10_A_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1482.440 4.000 1483.040 ;
    END
  END Tile_X0Y10_A_config_C_bit0
  PIN Tile_X0Y10_A_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1485.840 4.000 1486.440 ;
    END
  END Tile_X0Y10_A_config_C_bit1
  PIN Tile_X0Y10_A_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1489.240 4.000 1489.840 ;
    END
  END Tile_X0Y10_A_config_C_bit2
  PIN Tile_X0Y10_A_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1492.640 4.000 1493.240 ;
    END
  END Tile_X0Y10_A_config_C_bit3
  PIN Tile_X0Y10_B_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1472.240 4.000 1472.840 ;
    END
  END Tile_X0Y10_B_I_top
  PIN Tile_X0Y10_B_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1468.840 4.000 1469.440 ;
    END
  END Tile_X0Y10_B_O_top
  PIN Tile_X0Y10_B_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1475.640 4.000 1476.240 ;
    END
  END Tile_X0Y10_B_T_top
  PIN Tile_X0Y10_B_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1496.040 4.000 1496.640 ;
    END
  END Tile_X0Y10_B_config_C_bit0
  PIN Tile_X0Y10_B_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1502.840 4.000 1503.440 ;
    END
  END Tile_X0Y10_B_config_C_bit1
  PIN Tile_X0Y10_B_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1506.240 4.000 1506.840 ;
    END
  END Tile_X0Y10_B_config_C_bit2
  PIN Tile_X0Y10_B_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1509.640 4.000 1510.240 ;
    END
  END Tile_X0Y10_B_config_C_bit3
  PIN Tile_X0Y11_A_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1234.240 4.000 1234.840 ;
    END
  END Tile_X0Y11_A_I_top
  PIN Tile_X0Y11_A_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1230.840 4.000 1231.440 ;
    END
  END Tile_X0Y11_A_O_top
  PIN Tile_X0Y11_A_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1241.040 4.000 1241.640 ;
    END
  END Tile_X0Y11_A_T_top
  PIN Tile_X0Y11_A_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1254.640 4.000 1255.240 ;
    END
  END Tile_X0Y11_A_config_C_bit0
  PIN Tile_X0Y11_A_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1261.440 4.000 1262.040 ;
    END
  END Tile_X0Y11_A_config_C_bit1
  PIN Tile_X0Y11_A_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1264.840 4.000 1265.440 ;
    END
  END Tile_X0Y11_A_config_C_bit2
  PIN Tile_X0Y11_A_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1268.240 4.000 1268.840 ;
    END
  END Tile_X0Y11_A_config_C_bit3
  PIN Tile_X0Y11_B_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1247.840 4.000 1248.440 ;
    END
  END Tile_X0Y11_B_I_top
  PIN Tile_X0Y11_B_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1244.440 4.000 1245.040 ;
    END
  END Tile_X0Y11_B_O_top
  PIN Tile_X0Y11_B_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1251.240 4.000 1251.840 ;
    END
  END Tile_X0Y11_B_T_top
  PIN Tile_X0Y11_B_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1271.640 4.000 1272.240 ;
    END
  END Tile_X0Y11_B_config_C_bit0
  PIN Tile_X0Y11_B_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1275.040 4.000 1275.640 ;
    END
  END Tile_X0Y11_B_config_C_bit1
  PIN Tile_X0Y11_B_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1281.840 4.000 1282.440 ;
    END
  END Tile_X0Y11_B_config_C_bit2
  PIN Tile_X0Y11_B_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1285.240 4.000 1285.840 ;
    END
  END Tile_X0Y11_B_config_C_bit3
  PIN Tile_X0Y12_A_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1009.840 4.000 1010.440 ;
    END
  END Tile_X0Y12_A_I_top
  PIN Tile_X0Y12_A_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1006.440 4.000 1007.040 ;
    END
  END Tile_X0Y12_A_O_top
  PIN Tile_X0Y12_A_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1013.240 4.000 1013.840 ;
    END
  END Tile_X0Y12_A_T_top
  PIN Tile_X0Y12_A_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1030.240 4.000 1030.840 ;
    END
  END Tile_X0Y12_A_config_C_bit0
  PIN Tile_X0Y12_A_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1033.640 4.000 1034.240 ;
    END
  END Tile_X0Y12_A_config_C_bit1
  PIN Tile_X0Y12_A_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1040.440 4.000 1041.040 ;
    END
  END Tile_X0Y12_A_config_C_bit2
  PIN Tile_X0Y12_A_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1043.840 4.000 1044.440 ;
    END
  END Tile_X0Y12_A_config_C_bit3
  PIN Tile_X0Y12_B_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1023.440 4.000 1024.040 ;
    END
  END Tile_X0Y12_B_I_top
  PIN Tile_X0Y12_B_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1020.040 4.000 1020.640 ;
    END
  END Tile_X0Y12_B_O_top
  PIN Tile_X0Y12_B_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1026.840 4.000 1027.440 ;
    END
  END Tile_X0Y12_B_T_top
  PIN Tile_X0Y12_B_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1047.240 4.000 1047.840 ;
    END
  END Tile_X0Y12_B_config_C_bit0
  PIN Tile_X0Y12_B_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1050.640 4.000 1051.240 ;
    END
  END Tile_X0Y12_B_config_C_bit1
  PIN Tile_X0Y12_B_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1054.040 4.000 1054.640 ;
    END
  END Tile_X0Y12_B_config_C_bit2
  PIN Tile_X0Y12_B_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1057.440 4.000 1058.040 ;
    END
  END Tile_X0Y12_B_config_C_bit3
  PIN Tile_X0Y13_A_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 785.440 4.000 786.040 ;
    END
  END Tile_X0Y13_A_I_top
  PIN Tile_X0Y13_A_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 782.040 4.000 782.640 ;
    END
  END Tile_X0Y13_A_O_top
  PIN Tile_X0Y13_A_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 788.840 4.000 789.440 ;
    END
  END Tile_X0Y13_A_T_top
  PIN Tile_X0Y13_A_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 805.840 4.000 806.440 ;
    END
  END Tile_X0Y13_A_config_C_bit0
  PIN Tile_X0Y13_A_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 809.240 4.000 809.840 ;
    END
  END Tile_X0Y13_A_config_C_bit1
  PIN Tile_X0Y13_A_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 812.640 4.000 813.240 ;
    END
  END Tile_X0Y13_A_config_C_bit2
  PIN Tile_X0Y13_A_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 819.440 4.000 820.040 ;
    END
  END Tile_X0Y13_A_config_C_bit3
  PIN Tile_X0Y13_B_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 799.040 4.000 799.640 ;
    END
  END Tile_X0Y13_B_I_top
  PIN Tile_X0Y13_B_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 792.240 4.000 792.840 ;
    END
  END Tile_X0Y13_B_O_top
  PIN Tile_X0Y13_B_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 802.440 4.000 803.040 ;
    END
  END Tile_X0Y13_B_T_top
  PIN Tile_X0Y13_B_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 822.840 4.000 823.440 ;
    END
  END Tile_X0Y13_B_config_C_bit0
  PIN Tile_X0Y13_B_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 826.240 4.000 826.840 ;
    END
  END Tile_X0Y13_B_config_C_bit1
  PIN Tile_X0Y13_B_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 829.640 4.000 830.240 ;
    END
  END Tile_X0Y13_B_config_C_bit2
  PIN Tile_X0Y13_B_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 833.040 4.000 833.640 ;
    END
  END Tile_X0Y13_B_config_C_bit3
  PIN Tile_X0Y14_A_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 561.040 4.000 561.640 ;
    END
  END Tile_X0Y14_A_I_top
  PIN Tile_X0Y14_A_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 557.640 4.000 558.240 ;
    END
  END Tile_X0Y14_A_O_top
  PIN Tile_X0Y14_A_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 564.440 4.000 565.040 ;
    END
  END Tile_X0Y14_A_T_top
  PIN Tile_X0Y14_A_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 581.440 4.000 582.040 ;
    END
  END Tile_X0Y14_A_config_C_bit0
  PIN Tile_X0Y14_A_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 584.840 4.000 585.440 ;
    END
  END Tile_X0Y14_A_config_C_bit1
  PIN Tile_X0Y14_A_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 588.240 4.000 588.840 ;
    END
  END Tile_X0Y14_A_config_C_bit2
  PIN Tile_X0Y14_A_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 595.040 4.000 595.640 ;
    END
  END Tile_X0Y14_A_config_C_bit3
  PIN Tile_X0Y14_B_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 574.640 4.000 575.240 ;
    END
  END Tile_X0Y14_B_I_top
  PIN Tile_X0Y14_B_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 567.840 4.000 568.440 ;
    END
  END Tile_X0Y14_B_O_top
  PIN Tile_X0Y14_B_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 578.040 4.000 578.640 ;
    END
  END Tile_X0Y14_B_T_top
  PIN Tile_X0Y14_B_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 598.440 4.000 599.040 ;
    END
  END Tile_X0Y14_B_config_C_bit0
  PIN Tile_X0Y14_B_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 601.840 4.000 602.440 ;
    END
  END Tile_X0Y14_B_config_C_bit1
  PIN Tile_X0Y14_B_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 605.240 4.000 605.840 ;
    END
  END Tile_X0Y14_B_config_C_bit2
  PIN Tile_X0Y14_B_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 608.640 4.000 609.240 ;
    END
  END Tile_X0Y14_B_config_C_bit3
  PIN Tile_X0Y15_A_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 329.840 4.000 330.440 ;
    END
  END Tile_X0Y15_A_I_top
  PIN Tile_X0Y15_A_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 261.840 4.000 262.440 ;
    END
  END Tile_X0Y15_A_O_top
  PIN Tile_X0Y15_A_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 323.040 4.000 323.640 ;
    END
  END Tile_X0Y15_A_T_top
  PIN Tile_X0Y15_A_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 353.640 4.000 354.240 ;
    END
  END Tile_X0Y15_A_config_C_bit0
  PIN Tile_X0Y15_A_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 319.640 4.000 320.240 ;
    END
  END Tile_X0Y15_A_config_C_bit1
  PIN Tile_X0Y15_A_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 326.440 4.000 327.040 ;
    END
  END Tile_X0Y15_A_config_C_bit2
  PIN Tile_X0Y15_A_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 316.240 4.000 316.840 ;
    END
  END Tile_X0Y15_A_config_C_bit3
  PIN Tile_X0Y15_B_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 346.840 4.000 347.440 ;
    END
  END Tile_X0Y15_B_I_top
  PIN Tile_X0Y15_B_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 241.440 4.000 242.040 ;
    END
  END Tile_X0Y15_B_O_top
  PIN Tile_X0Y15_B_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 350.240 4.000 350.840 ;
    END
  END Tile_X0Y15_B_T_top
  PIN Tile_X0Y15_B_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 309.440 4.000 310.040 ;
    END
  END Tile_X0Y15_B_config_C_bit0
  PIN Tile_X0Y15_B_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 357.040 4.000 357.640 ;
    END
  END Tile_X0Y15_B_config_C_bit1
  PIN Tile_X0Y15_B_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 306.040 4.000 306.640 ;
    END
  END Tile_X0Y15_B_config_C_bit2
  PIN Tile_X0Y15_B_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 340.040 4.000 340.640 ;
    END
  END Tile_X0Y15_B_config_C_bit3
  PIN Tile_X0Y16_A_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 122.440 4.000 123.040 ;
    END
  END Tile_X0Y16_A_I_top
  PIN Tile_X0Y16_A_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.840 4.000 109.440 ;
    END
  END Tile_X0Y16_A_O_top
  PIN Tile_X0Y16_A_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 32.290 0.000 32.570 4.000 ;
    END
  END Tile_X0Y16_A_T_top
  PIN Tile_X0Y16_A_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 51.610 0.000 51.890 4.000 ;
    END
  END Tile_X0Y16_A_config_C_bit0
  PIN Tile_X0Y16_A_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 61.270 0.000 61.550 4.000 ;
    END
  END Tile_X0Y16_A_config_C_bit1
  PIN Tile_X0Y16_A_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 67.710 0.000 67.990 4.000 ;
    END
  END Tile_X0Y16_A_config_C_bit2
  PIN Tile_X0Y16_A_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 54.830 0.000 55.110 4.000 ;
    END
  END Tile_X0Y16_A_config_C_bit3
  PIN Tile_X0Y16_B_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 45.170 0.000 45.450 4.000 ;
    END
  END Tile_X0Y16_B_I_top
  PIN Tile_X0Y16_B_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 38.730 0.000 39.010 4.000 ;
    END
  END Tile_X0Y16_B_O_top
  PIN Tile_X0Y16_B_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 58.050 0.000 58.330 4.000 ;
    END
  END Tile_X0Y16_B_T_top
  PIN Tile_X0Y16_B_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 48.390 0.000 48.670 4.000 ;
    END
  END Tile_X0Y16_B_config_C_bit0
  PIN Tile_X0Y16_B_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 64.490 0.000 64.770 4.000 ;
    END
  END Tile_X0Y16_B_config_C_bit1
  PIN Tile_X0Y16_B_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 35.510 0.000 35.790 4.000 ;
    END
  END Tile_X0Y16_B_config_C_bit2
  PIN Tile_X0Y16_B_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 41.950 0.000 42.230 4.000 ;
    END
  END Tile_X0Y16_B_config_C_bit3
  PIN Tile_X0Y1_A_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3485.040 4.000 3485.640 ;
    END
  END Tile_X0Y1_A_I_top
  PIN Tile_X0Y1_A_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3481.640 4.000 3482.240 ;
    END
  END Tile_X0Y1_A_O_top
  PIN Tile_X0Y1_A_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3488.440 4.000 3489.040 ;
    END
  END Tile_X0Y1_A_T_top
  PIN Tile_X0Y1_A_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3505.440 4.000 3506.040 ;
    END
  END Tile_X0Y1_A_config_C_bit0
  PIN Tile_X0Y1_A_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3508.840 4.000 3509.440 ;
    END
  END Tile_X0Y1_A_config_C_bit1
  PIN Tile_X0Y1_A_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3515.640 4.000 3516.240 ;
    END
  END Tile_X0Y1_A_config_C_bit2
  PIN Tile_X0Y1_A_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3519.040 4.000 3519.640 ;
    END
  END Tile_X0Y1_A_config_C_bit3
  PIN Tile_X0Y1_B_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3498.640 4.000 3499.240 ;
    END
  END Tile_X0Y1_B_I_top
  PIN Tile_X0Y1_B_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3495.240 4.000 3495.840 ;
    END
  END Tile_X0Y1_B_O_top
  PIN Tile_X0Y1_B_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3502.040 4.000 3502.640 ;
    END
  END Tile_X0Y1_B_T_top
  PIN Tile_X0Y1_B_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3522.440 4.000 3523.040 ;
    END
  END Tile_X0Y1_B_config_C_bit0
  PIN Tile_X0Y1_B_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3525.840 4.000 3526.440 ;
    END
  END Tile_X0Y1_B_config_C_bit1
  PIN Tile_X0Y1_B_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3529.240 4.000 3529.840 ;
    END
  END Tile_X0Y1_B_config_C_bit2
  PIN Tile_X0Y1_B_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3536.040 4.000 3536.640 ;
    END
  END Tile_X0Y1_B_config_C_bit3
  PIN Tile_X0Y2_A_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3260.640 4.000 3261.240 ;
    END
  END Tile_X0Y2_A_I_top
  PIN Tile_X0Y2_A_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3257.240 4.000 3257.840 ;
    END
  END Tile_X0Y2_A_O_top
  PIN Tile_X0Y2_A_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3264.040 4.000 3264.640 ;
    END
  END Tile_X0Y2_A_T_top
  PIN Tile_X0Y2_A_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3281.040 4.000 3281.640 ;
    END
  END Tile_X0Y2_A_config_C_bit0
  PIN Tile_X0Y2_A_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3284.440 4.000 3285.040 ;
    END
  END Tile_X0Y2_A_config_C_bit1
  PIN Tile_X0Y2_A_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3287.840 4.000 3288.440 ;
    END
  END Tile_X0Y2_A_config_C_bit2
  PIN Tile_X0Y2_A_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3294.640 4.000 3295.240 ;
    END
  END Tile_X0Y2_A_config_C_bit3
  PIN Tile_X0Y2_B_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3274.240 4.000 3274.840 ;
    END
  END Tile_X0Y2_B_I_top
  PIN Tile_X0Y2_B_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3267.440 4.000 3268.040 ;
    END
  END Tile_X0Y2_B_O_top
  PIN Tile_X0Y2_B_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3277.640 4.000 3278.240 ;
    END
  END Tile_X0Y2_B_T_top
  PIN Tile_X0Y2_B_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3298.040 4.000 3298.640 ;
    END
  END Tile_X0Y2_B_config_C_bit0
  PIN Tile_X0Y2_B_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3301.440 4.000 3302.040 ;
    END
  END Tile_X0Y2_B_config_C_bit1
  PIN Tile_X0Y2_B_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3304.840 4.000 3305.440 ;
    END
  END Tile_X0Y2_B_config_C_bit2
  PIN Tile_X0Y2_B_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3308.240 4.000 3308.840 ;
    END
  END Tile_X0Y2_B_config_C_bit3
  PIN Tile_X0Y3_A_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3036.240 4.000 3036.840 ;
    END
  END Tile_X0Y3_A_I_top
  PIN Tile_X0Y3_A_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3032.840 4.000 3033.440 ;
    END
  END Tile_X0Y3_A_O_top
  PIN Tile_X0Y3_A_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3039.640 4.000 3040.240 ;
    END
  END Tile_X0Y3_A_T_top
  PIN Tile_X0Y3_A_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3056.640 4.000 3057.240 ;
    END
  END Tile_X0Y3_A_config_C_bit0
  PIN Tile_X0Y3_A_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3060.040 4.000 3060.640 ;
    END
  END Tile_X0Y3_A_config_C_bit1
  PIN Tile_X0Y3_A_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3063.440 4.000 3064.040 ;
    END
  END Tile_X0Y3_A_config_C_bit2
  PIN Tile_X0Y3_A_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3066.840 4.000 3067.440 ;
    END
  END Tile_X0Y3_A_config_C_bit3
  PIN Tile_X0Y3_B_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3046.440 4.000 3047.040 ;
    END
  END Tile_X0Y3_B_I_top
  PIN Tile_X0Y3_B_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3043.040 4.000 3043.640 ;
    END
  END Tile_X0Y3_B_O_top
  PIN Tile_X0Y3_B_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3053.240 4.000 3053.840 ;
    END
  END Tile_X0Y3_B_T_top
  PIN Tile_X0Y3_B_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3073.640 4.000 3074.240 ;
    END
  END Tile_X0Y3_B_config_C_bit0
  PIN Tile_X0Y3_B_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3077.040 4.000 3077.640 ;
    END
  END Tile_X0Y3_B_config_C_bit1
  PIN Tile_X0Y3_B_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3080.440 4.000 3081.040 ;
    END
  END Tile_X0Y3_B_config_C_bit2
  PIN Tile_X0Y3_B_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3083.840 4.000 3084.440 ;
    END
  END Tile_X0Y3_B_config_C_bit3
  PIN Tile_X0Y4_A_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2811.840 4.000 2812.440 ;
    END
  END Tile_X0Y4_A_I_top
  PIN Tile_X0Y4_A_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2805.040 4.000 2805.640 ;
    END
  END Tile_X0Y4_A_O_top
  PIN Tile_X0Y4_A_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2815.240 4.000 2815.840 ;
    END
  END Tile_X0Y4_A_T_top
  PIN Tile_X0Y4_A_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2832.240 4.000 2832.840 ;
    END
  END Tile_X0Y4_A_config_C_bit0
  PIN Tile_X0Y4_A_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2835.640 4.000 2836.240 ;
    END
  END Tile_X0Y4_A_config_C_bit1
  PIN Tile_X0Y4_A_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2839.040 4.000 2839.640 ;
    END
  END Tile_X0Y4_A_config_C_bit2
  PIN Tile_X0Y4_A_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2842.440 4.000 2843.040 ;
    END
  END Tile_X0Y4_A_config_C_bit3
  PIN Tile_X0Y4_B_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2822.040 4.000 2822.640 ;
    END
  END Tile_X0Y4_B_I_top
  PIN Tile_X0Y4_B_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2818.640 4.000 2819.240 ;
    END
  END Tile_X0Y4_B_O_top
  PIN Tile_X0Y4_B_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2825.440 4.000 2826.040 ;
    END
  END Tile_X0Y4_B_T_top
  PIN Tile_X0Y4_B_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2845.840 4.000 2846.440 ;
    END
  END Tile_X0Y4_B_config_C_bit0
  PIN Tile_X0Y4_B_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2852.640 4.000 2853.240 ;
    END
  END Tile_X0Y4_B_config_C_bit1
  PIN Tile_X0Y4_B_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2856.040 4.000 2856.640 ;
    END
  END Tile_X0Y4_B_config_C_bit2
  PIN Tile_X0Y4_B_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2859.440 4.000 2860.040 ;
    END
  END Tile_X0Y4_B_config_C_bit3
  PIN Tile_X0Y5_A_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2587.440 4.000 2588.040 ;
    END
  END Tile_X0Y5_A_I_top
  PIN Tile_X0Y5_A_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2580.640 4.000 2581.240 ;
    END
  END Tile_X0Y5_A_O_top
  PIN Tile_X0Y5_A_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2590.840 4.000 2591.440 ;
    END
  END Tile_X0Y5_A_T_top
  PIN Tile_X0Y5_A_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2607.840 4.000 2608.440 ;
    END
  END Tile_X0Y5_A_config_C_bit0
  PIN Tile_X0Y5_A_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2611.240 4.000 2611.840 ;
    END
  END Tile_X0Y5_A_config_C_bit1
  PIN Tile_X0Y5_A_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2614.640 4.000 2615.240 ;
    END
  END Tile_X0Y5_A_config_C_bit2
  PIN Tile_X0Y5_A_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2618.040 4.000 2618.640 ;
    END
  END Tile_X0Y5_A_config_C_bit3
  PIN Tile_X0Y5_B_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2597.640 4.000 2598.240 ;
    END
  END Tile_X0Y5_B_I_top
  PIN Tile_X0Y5_B_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2594.240 4.000 2594.840 ;
    END
  END Tile_X0Y5_B_O_top
  PIN Tile_X0Y5_B_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2601.040 4.000 2601.640 ;
    END
  END Tile_X0Y5_B_T_top
  PIN Tile_X0Y5_B_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2621.440 4.000 2622.040 ;
    END
  END Tile_X0Y5_B_config_C_bit0
  PIN Tile_X0Y5_B_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2628.240 4.000 2628.840 ;
    END
  END Tile_X0Y5_B_config_C_bit1
  PIN Tile_X0Y5_B_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2631.640 4.000 2632.240 ;
    END
  END Tile_X0Y5_B_config_C_bit2
  PIN Tile_X0Y5_B_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2635.040 4.000 2635.640 ;
    END
  END Tile_X0Y5_B_config_C_bit3
  PIN Tile_X0Y6_A_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2359.640 4.000 2360.240 ;
    END
  END Tile_X0Y6_A_I_top
  PIN Tile_X0Y6_A_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2356.240 4.000 2356.840 ;
    END
  END Tile_X0Y6_A_O_top
  PIN Tile_X0Y6_A_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2366.440 4.000 2367.040 ;
    END
  END Tile_X0Y6_A_T_top
  PIN Tile_X0Y6_A_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2380.040 4.000 2380.640 ;
    END
  END Tile_X0Y6_A_config_C_bit0
  PIN Tile_X0Y6_A_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2386.840 4.000 2387.440 ;
    END
  END Tile_X0Y6_A_config_C_bit1
  PIN Tile_X0Y6_A_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2390.240 4.000 2390.840 ;
    END
  END Tile_X0Y6_A_config_C_bit2
  PIN Tile_X0Y6_A_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2393.640 4.000 2394.240 ;
    END
  END Tile_X0Y6_A_config_C_bit3
  PIN Tile_X0Y6_B_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2373.240 4.000 2373.840 ;
    END
  END Tile_X0Y6_B_I_top
  PIN Tile_X0Y6_B_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2369.840 4.000 2370.440 ;
    END
  END Tile_X0Y6_B_O_top
  PIN Tile_X0Y6_B_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2376.640 4.000 2377.240 ;
    END
  END Tile_X0Y6_B_T_top
  PIN Tile_X0Y6_B_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2397.040 4.000 2397.640 ;
    END
  END Tile_X0Y6_B_config_C_bit0
  PIN Tile_X0Y6_B_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2400.440 4.000 2401.040 ;
    END
  END Tile_X0Y6_B_config_C_bit1
  PIN Tile_X0Y6_B_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2407.240 4.000 2407.840 ;
    END
  END Tile_X0Y6_B_config_C_bit2
  PIN Tile_X0Y6_B_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2410.640 4.000 2411.240 ;
    END
  END Tile_X0Y6_B_config_C_bit3
  PIN Tile_X0Y7_A_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2135.240 4.000 2135.840 ;
    END
  END Tile_X0Y7_A_I_top
  PIN Tile_X0Y7_A_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2131.840 4.000 2132.440 ;
    END
  END Tile_X0Y7_A_O_top
  PIN Tile_X0Y7_A_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2138.640 4.000 2139.240 ;
    END
  END Tile_X0Y7_A_T_top
  PIN Tile_X0Y7_A_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2155.640 4.000 2156.240 ;
    END
  END Tile_X0Y7_A_config_C_bit0
  PIN Tile_X0Y7_A_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2159.040 4.000 2159.640 ;
    END
  END Tile_X0Y7_A_config_C_bit1
  PIN Tile_X0Y7_A_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2165.840 4.000 2166.440 ;
    END
  END Tile_X0Y7_A_config_C_bit2
  PIN Tile_X0Y7_A_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2169.240 4.000 2169.840 ;
    END
  END Tile_X0Y7_A_config_C_bit3
  PIN Tile_X0Y7_B_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2148.840 4.000 2149.440 ;
    END
  END Tile_X0Y7_B_I_top
  PIN Tile_X0Y7_B_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2145.440 4.000 2146.040 ;
    END
  END Tile_X0Y7_B_O_top
  PIN Tile_X0Y7_B_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2152.240 4.000 2152.840 ;
    END
  END Tile_X0Y7_B_T_top
  PIN Tile_X0Y7_B_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2172.640 4.000 2173.240 ;
    END
  END Tile_X0Y7_B_config_C_bit0
  PIN Tile_X0Y7_B_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2176.040 4.000 2176.640 ;
    END
  END Tile_X0Y7_B_config_C_bit1
  PIN Tile_X0Y7_B_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2179.440 4.000 2180.040 ;
    END
  END Tile_X0Y7_B_config_C_bit2
  PIN Tile_X0Y7_B_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2186.240 4.000 2186.840 ;
    END
  END Tile_X0Y7_B_config_C_bit3
  PIN Tile_X0Y8_A_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1910.840 4.000 1911.440 ;
    END
  END Tile_X0Y8_A_I_top
  PIN Tile_X0Y8_A_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1907.440 4.000 1908.040 ;
    END
  END Tile_X0Y8_A_O_top
  PIN Tile_X0Y8_A_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1914.240 4.000 1914.840 ;
    END
  END Tile_X0Y8_A_T_top
  PIN Tile_X0Y8_A_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1931.240 4.000 1931.840 ;
    END
  END Tile_X0Y8_A_config_C_bit0
  PIN Tile_X0Y8_A_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1934.640 4.000 1935.240 ;
    END
  END Tile_X0Y8_A_config_C_bit1
  PIN Tile_X0Y8_A_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1938.040 4.000 1938.640 ;
    END
  END Tile_X0Y8_A_config_C_bit2
  PIN Tile_X0Y8_A_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1944.840 4.000 1945.440 ;
    END
  END Tile_X0Y8_A_config_C_bit3
  PIN Tile_X0Y8_B_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1924.440 4.000 1925.040 ;
    END
  END Tile_X0Y8_B_I_top
  PIN Tile_X0Y8_B_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1917.640 4.000 1918.240 ;
    END
  END Tile_X0Y8_B_O_top
  PIN Tile_X0Y8_B_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1927.840 4.000 1928.440 ;
    END
  END Tile_X0Y8_B_T_top
  PIN Tile_X0Y8_B_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1948.240 4.000 1948.840 ;
    END
  END Tile_X0Y8_B_config_C_bit0
  PIN Tile_X0Y8_B_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1951.640 4.000 1952.240 ;
    END
  END Tile_X0Y8_B_config_C_bit1
  PIN Tile_X0Y8_B_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1955.040 4.000 1955.640 ;
    END
  END Tile_X0Y8_B_config_C_bit2
  PIN Tile_X0Y8_B_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1958.440 4.000 1959.040 ;
    END
  END Tile_X0Y8_B_config_C_bit3
  PIN Tile_X0Y9_A_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1686.440 4.000 1687.040 ;
    END
  END Tile_X0Y9_A_I_top
  PIN Tile_X0Y9_A_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1683.040 4.000 1683.640 ;
    END
  END Tile_X0Y9_A_O_top
  PIN Tile_X0Y9_A_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1689.840 4.000 1690.440 ;
    END
  END Tile_X0Y9_A_T_top
  PIN Tile_X0Y9_A_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1706.840 4.000 1707.440 ;
    END
  END Tile_X0Y9_A_config_C_bit0
  PIN Tile_X0Y9_A_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1710.240 4.000 1710.840 ;
    END
  END Tile_X0Y9_A_config_C_bit1
  PIN Tile_X0Y9_A_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1713.640 4.000 1714.240 ;
    END
  END Tile_X0Y9_A_config_C_bit2
  PIN Tile_X0Y9_A_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1717.040 4.000 1717.640 ;
    END
  END Tile_X0Y9_A_config_C_bit3
  PIN Tile_X0Y9_B_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1696.640 4.000 1697.240 ;
    END
  END Tile_X0Y9_B_I_top
  PIN Tile_X0Y9_B_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1693.240 4.000 1693.840 ;
    END
  END Tile_X0Y9_B_O_top
  PIN Tile_X0Y9_B_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1703.440 4.000 1704.040 ;
    END
  END Tile_X0Y9_B_T_top
  PIN Tile_X0Y9_B_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1723.840 4.000 1724.440 ;
    END
  END Tile_X0Y9_B_config_C_bit0
  PIN Tile_X0Y9_B_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1727.240 4.000 1727.840 ;
    END
  END Tile_X0Y9_B_config_C_bit1
  PIN Tile_X0Y9_B_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1730.640 4.000 1731.240 ;
    END
  END Tile_X0Y9_B_config_C_bit2
  PIN Tile_X0Y9_B_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1734.040 4.000 1734.640 ;
    END
  END Tile_X0Y9_B_config_C_bit3
  PIN Tile_X10Y0_A_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 2025.470 3778.500 2025.750 3782.500 ;
    END
  END Tile_X10Y0_A_I_top
  PIN Tile_X10Y0_A_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 2019.030 3778.500 2019.310 3782.500 ;
    END
  END Tile_X10Y0_A_O_top
  PIN Tile_X10Y0_A_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 2031.910 3778.500 2032.190 3782.500 ;
    END
  END Tile_X10Y0_A_T_top
  PIN Tile_X10Y0_A_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 2051.230 3778.500 2051.510 3782.500 ;
    END
  END Tile_X10Y0_A_config_C_bit0
  PIN Tile_X10Y0_A_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 2057.670 3778.500 2057.950 3782.500 ;
    END
  END Tile_X10Y0_A_config_C_bit1
  PIN Tile_X10Y0_A_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 2064.110 3778.500 2064.390 3782.500 ;
    END
  END Tile_X10Y0_A_config_C_bit2
  PIN Tile_X10Y0_A_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 2070.550 3778.500 2070.830 3782.500 ;
    END
  END Tile_X10Y0_A_config_C_bit3
  PIN Tile_X10Y0_B_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 2041.570 3778.500 2041.850 3782.500 ;
    END
  END Tile_X10Y0_B_I_top
  PIN Tile_X10Y0_B_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 2035.130 3778.500 2035.410 3782.500 ;
    END
  END Tile_X10Y0_B_O_top
  PIN Tile_X10Y0_B_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 2048.010 3778.500 2048.290 3782.500 ;
    END
  END Tile_X10Y0_B_T_top
  PIN Tile_X10Y0_B_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 2073.770 3778.500 2074.050 3782.500 ;
    END
  END Tile_X10Y0_B_config_C_bit0
  PIN Tile_X10Y0_B_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 2080.210 3778.500 2080.490 3782.500 ;
    END
  END Tile_X10Y0_B_config_C_bit1
  PIN Tile_X10Y0_B_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 2086.650 3778.500 2086.930 3782.500 ;
    END
  END Tile_X10Y0_B_config_C_bit2
  PIN Tile_X10Y0_B_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 2089.870 3778.500 2090.150 3782.500 ;
    END
  END Tile_X10Y0_B_config_C_bit3
  PIN Tile_X10Y17_VALUE_top0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 2015.810 0.000 2016.090 4.000 ;
    END
  END Tile_X10Y17_VALUE_top0
  PIN Tile_X10Y17_VALUE_top1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 2022.250 0.000 2022.530 4.000 ;
    END
  END Tile_X10Y17_VALUE_top1
  PIN Tile_X10Y17_VALUE_top2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 2031.910 0.000 2032.190 4.000 ;
    END
  END Tile_X10Y17_VALUE_top2
  PIN Tile_X10Y17_VALUE_top3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 2038.350 0.000 2038.630 4.000 ;
    END
  END Tile_X10Y17_VALUE_top3
  PIN Tile_X10Y17_VALUE_top4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 2044.790 0.000 2045.070 4.000 ;
    END
  END Tile_X10Y17_VALUE_top4
  PIN Tile_X10Y17_VALUE_top5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 2051.230 0.000 2051.510 4.000 ;
    END
  END Tile_X10Y17_VALUE_top5
  PIN Tile_X10Y17_VALUE_top6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 2057.670 0.000 2057.950 4.000 ;
    END
  END Tile_X10Y17_VALUE_top6
  PIN Tile_X10Y17_VALUE_top7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 2064.110 0.000 2064.390 4.000 ;
    END
  END Tile_X10Y17_VALUE_top7
  PIN Tile_X11Y10_AD_SRAM0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1434.840 2435.000 1435.440 ;
    END
  END Tile_X11Y10_AD_SRAM0
  PIN Tile_X11Y10_AD_SRAM1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1587.840 2435.000 1588.440 ;
    END
  END Tile_X11Y10_AD_SRAM1
  PIN Tile_X11Y10_AD_SRAM2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1475.640 2435.000 1476.240 ;
    END
  END Tile_X11Y10_AD_SRAM2
  PIN Tile_X11Y10_AD_SRAM3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1591.240 2435.000 1591.840 ;
    END
  END Tile_X11Y10_AD_SRAM3
  PIN Tile_X11Y10_AD_SRAM4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1472.240 2435.000 1472.840 ;
    END
  END Tile_X11Y10_AD_SRAM4
  PIN Tile_X11Y10_AD_SRAM5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1468.840 2435.000 1469.440 ;
    END
  END Tile_X11Y10_AD_SRAM5
  PIN Tile_X11Y10_AD_SRAM6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1594.640 2435.000 1595.240 ;
    END
  END Tile_X11Y10_AD_SRAM6
  PIN Tile_X11Y10_AD_SRAM7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1465.440 2435.000 1466.040 ;
    END
  END Tile_X11Y10_AD_SRAM7
  PIN Tile_X11Y10_AD_SRAM8
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1598.040 2435.000 1598.640 ;
    END
  END Tile_X11Y10_AD_SRAM8
  PIN Tile_X11Y10_AD_SRAM9
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1462.040 2435.000 1462.640 ;
    END
  END Tile_X11Y10_AD_SRAM9
  PIN Tile_X11Y10_BEN_SRAM0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1458.640 2435.000 1459.240 ;
    END
  END Tile_X11Y10_BEN_SRAM0
  PIN Tile_X11Y10_BEN_SRAM1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1601.440 2435.000 1602.040 ;
    END
  END Tile_X11Y10_BEN_SRAM1
  PIN Tile_X11Y10_BEN_SRAM10
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1438.240 2435.000 1438.840 ;
    END
  END Tile_X11Y10_BEN_SRAM10
  PIN Tile_X11Y10_BEN_SRAM11
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1615.040 2435.000 1615.640 ;
    END
  END Tile_X11Y10_BEN_SRAM11
  PIN Tile_X11Y10_BEN_SRAM12
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1618.440 2435.000 1619.040 ;
    END
  END Tile_X11Y10_BEN_SRAM12
  PIN Tile_X11Y10_BEN_SRAM13
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1802.040 2435.000 1802.640 ;
    END
  END Tile_X11Y10_BEN_SRAM13
  PIN Tile_X11Y10_BEN_SRAM14
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1798.640 2435.000 1799.240 ;
    END
  END Tile_X11Y10_BEN_SRAM14
  PIN Tile_X11Y10_BEN_SRAM15
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1621.840 2435.000 1622.440 ;
    END
  END Tile_X11Y10_BEN_SRAM15
  PIN Tile_X11Y10_BEN_SRAM16
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1795.240 2435.000 1795.840 ;
    END
  END Tile_X11Y10_BEN_SRAM16
  PIN Tile_X11Y10_BEN_SRAM17
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1625.240 2435.000 1625.840 ;
    END
  END Tile_X11Y10_BEN_SRAM17
  PIN Tile_X11Y10_BEN_SRAM18
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1791.840 2435.000 1792.440 ;
    END
  END Tile_X11Y10_BEN_SRAM18
  PIN Tile_X11Y10_BEN_SRAM19
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1788.440 2435.000 1789.040 ;
    END
  END Tile_X11Y10_BEN_SRAM19
  PIN Tile_X11Y10_BEN_SRAM2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1455.240 2435.000 1455.840 ;
    END
  END Tile_X11Y10_BEN_SRAM2
  PIN Tile_X11Y10_BEN_SRAM20
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1628.640 2435.000 1629.240 ;
    END
  END Tile_X11Y10_BEN_SRAM20
  PIN Tile_X11Y10_BEN_SRAM21
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1785.040 2435.000 1785.640 ;
    END
  END Tile_X11Y10_BEN_SRAM21
  PIN Tile_X11Y10_BEN_SRAM22
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1632.040 2435.000 1632.640 ;
    END
  END Tile_X11Y10_BEN_SRAM22
  PIN Tile_X11Y10_BEN_SRAM23
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1781.640 2435.000 1782.240 ;
    END
  END Tile_X11Y10_BEN_SRAM23
  PIN Tile_X11Y10_BEN_SRAM24
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1778.240 2435.000 1778.840 ;
    END
  END Tile_X11Y10_BEN_SRAM24
  PIN Tile_X11Y10_BEN_SRAM25
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1635.440 2435.000 1636.040 ;
    END
  END Tile_X11Y10_BEN_SRAM25
  PIN Tile_X11Y10_BEN_SRAM26
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1774.840 2435.000 1775.440 ;
    END
  END Tile_X11Y10_BEN_SRAM26
  PIN Tile_X11Y10_BEN_SRAM27
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1638.840 2435.000 1639.440 ;
    END
  END Tile_X11Y10_BEN_SRAM27
  PIN Tile_X11Y10_BEN_SRAM28
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1771.440 2435.000 1772.040 ;
    END
  END Tile_X11Y10_BEN_SRAM28
  PIN Tile_X11Y10_BEN_SRAM29
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1768.040 2435.000 1768.640 ;
    END
  END Tile_X11Y10_BEN_SRAM29
  PIN Tile_X11Y10_BEN_SRAM3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1604.840 2435.000 1605.440 ;
    END
  END Tile_X11Y10_BEN_SRAM3
  PIN Tile_X11Y10_BEN_SRAM30
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1642.240 2435.000 1642.840 ;
    END
  END Tile_X11Y10_BEN_SRAM30
  PIN Tile_X11Y10_BEN_SRAM31
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1764.640 2435.000 1765.240 ;
    END
  END Tile_X11Y10_BEN_SRAM31
  PIN Tile_X11Y10_BEN_SRAM4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1451.840 2435.000 1452.440 ;
    END
  END Tile_X11Y10_BEN_SRAM4
  PIN Tile_X11Y10_BEN_SRAM5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1448.440 2435.000 1449.040 ;
    END
  END Tile_X11Y10_BEN_SRAM5
  PIN Tile_X11Y10_BEN_SRAM6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1608.240 2435.000 1608.840 ;
    END
  END Tile_X11Y10_BEN_SRAM6
  PIN Tile_X11Y10_BEN_SRAM7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1445.040 2435.000 1445.640 ;
    END
  END Tile_X11Y10_BEN_SRAM7
  PIN Tile_X11Y10_BEN_SRAM8
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1611.640 2435.000 1612.240 ;
    END
  END Tile_X11Y10_BEN_SRAM8
  PIN Tile_X11Y10_BEN_SRAM9
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1441.640 2435.000 1442.240 ;
    END
  END Tile_X11Y10_BEN_SRAM9
  PIN Tile_X11Y10_CLOCK_SRAM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1645.640 2435.000 1646.240 ;
    END
  END Tile_X11Y10_CLOCK_SRAM
  PIN Tile_X11Y10_DI_SRAM0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1761.240 2435.000 1761.840 ;
    END
  END Tile_X11Y10_DI_SRAM0
  PIN Tile_X11Y10_DI_SRAM1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1757.840 2435.000 1758.440 ;
    END
  END Tile_X11Y10_DI_SRAM1
  PIN Tile_X11Y10_DI_SRAM10
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1754.440 2435.000 1755.040 ;
    END
  END Tile_X11Y10_DI_SRAM10
  PIN Tile_X11Y10_DI_SRAM11
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1737.440 2435.000 1738.040 ;
    END
  END Tile_X11Y10_DI_SRAM11
  PIN Tile_X11Y10_DI_SRAM12
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1672.840 2435.000 1673.440 ;
    END
  END Tile_X11Y10_DI_SRAM12
  PIN Tile_X11Y10_DI_SRAM13
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1734.040 2435.000 1734.640 ;
    END
  END Tile_X11Y10_DI_SRAM13
  PIN Tile_X11Y10_DI_SRAM14
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1676.240 2435.000 1676.840 ;
    END
  END Tile_X11Y10_DI_SRAM14
  PIN Tile_X11Y10_DI_SRAM15
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1730.640 2435.000 1731.240 ;
    END
  END Tile_X11Y10_DI_SRAM15
  PIN Tile_X11Y10_DI_SRAM16
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1727.240 2435.000 1727.840 ;
    END
  END Tile_X11Y10_DI_SRAM16
  PIN Tile_X11Y10_DI_SRAM17
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1679.640 2435.000 1680.240 ;
    END
  END Tile_X11Y10_DI_SRAM17
  PIN Tile_X11Y10_DI_SRAM18
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1723.840 2435.000 1724.440 ;
    END
  END Tile_X11Y10_DI_SRAM18
  PIN Tile_X11Y10_DI_SRAM19
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1683.040 2435.000 1683.640 ;
    END
  END Tile_X11Y10_DI_SRAM19
  PIN Tile_X11Y10_DI_SRAM2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1649.040 2435.000 1649.640 ;
    END
  END Tile_X11Y10_DI_SRAM2
  PIN Tile_X11Y10_DI_SRAM20
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1720.440 2435.000 1721.040 ;
    END
  END Tile_X11Y10_DI_SRAM20
  PIN Tile_X11Y10_DI_SRAM21
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1717.040 2435.000 1717.640 ;
    END
  END Tile_X11Y10_DI_SRAM21
  PIN Tile_X11Y10_DI_SRAM22
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1751.040 2435.000 1751.640 ;
    END
  END Tile_X11Y10_DI_SRAM22
  PIN Tile_X11Y10_DI_SRAM23
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1713.640 2435.000 1714.240 ;
    END
  END Tile_X11Y10_DI_SRAM23
  PIN Tile_X11Y10_DI_SRAM24
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1747.640 2435.000 1748.240 ;
    END
  END Tile_X11Y10_DI_SRAM24
  PIN Tile_X11Y10_DI_SRAM25
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1744.240 2435.000 1744.840 ;
    END
  END Tile_X11Y10_DI_SRAM25
  PIN Tile_X11Y10_DI_SRAM26
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1706.840 2435.000 1707.440 ;
    END
  END Tile_X11Y10_DI_SRAM26
  PIN Tile_X11Y10_DI_SRAM27
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1740.840 2435.000 1741.440 ;
    END
  END Tile_X11Y10_DI_SRAM27
  PIN Tile_X11Y10_DI_SRAM28
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1703.440 2435.000 1704.040 ;
    END
  END Tile_X11Y10_DI_SRAM28
  PIN Tile_X11Y10_DI_SRAM29
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1686.440 2435.000 1687.040 ;
    END
  END Tile_X11Y10_DI_SRAM29
  PIN Tile_X11Y10_DI_SRAM3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1652.440 2435.000 1653.040 ;
    END
  END Tile_X11Y10_DI_SRAM3
  PIN Tile_X11Y10_DI_SRAM30
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1700.040 2435.000 1700.640 ;
    END
  END Tile_X11Y10_DI_SRAM30
  PIN Tile_X11Y10_DI_SRAM31
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1696.640 2435.000 1697.240 ;
    END
  END Tile_X11Y10_DI_SRAM31
  PIN Tile_X11Y10_DI_SRAM4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1655.840 2435.000 1656.440 ;
    END
  END Tile_X11Y10_DI_SRAM4
  PIN Tile_X11Y10_DI_SRAM5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1659.240 2435.000 1659.840 ;
    END
  END Tile_X11Y10_DI_SRAM5
  PIN Tile_X11Y10_DI_SRAM6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1693.240 2435.000 1693.840 ;
    END
  END Tile_X11Y10_DI_SRAM6
  PIN Tile_X11Y10_DI_SRAM7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1662.640 2435.000 1663.240 ;
    END
  END Tile_X11Y10_DI_SRAM7
  PIN Tile_X11Y10_DI_SRAM8
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1666.040 2435.000 1666.640 ;
    END
  END Tile_X11Y10_DI_SRAM8
  PIN Tile_X11Y10_DI_SRAM9
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1669.440 2435.000 1670.040 ;
    END
  END Tile_X11Y10_DI_SRAM9
  PIN Tile_X11Y10_DO_SRAM0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1479.040 2435.000 1479.640 ;
    END
  END Tile_X11Y10_DO_SRAM0
  PIN Tile_X11Y10_DO_SRAM1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1543.640 2435.000 1544.240 ;
    END
  END Tile_X11Y10_DO_SRAM1
  PIN Tile_X11Y10_DO_SRAM10
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1557.240 2435.000 1557.840 ;
    END
  END Tile_X11Y10_DO_SRAM10
  PIN Tile_X11Y10_DO_SRAM11
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1523.240 2435.000 1523.840 ;
    END
  END Tile_X11Y10_DO_SRAM11
  PIN Tile_X11Y10_DO_SRAM12
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1519.840 2435.000 1520.440 ;
    END
  END Tile_X11Y10_DO_SRAM12
  PIN Tile_X11Y10_DO_SRAM13
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1560.640 2435.000 1561.240 ;
    END
  END Tile_X11Y10_DO_SRAM13
  PIN Tile_X11Y10_DO_SRAM14
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1516.440 2435.000 1517.040 ;
    END
  END Tile_X11Y10_DO_SRAM14
  PIN Tile_X11Y10_DO_SRAM15
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1564.040 2435.000 1564.640 ;
    END
  END Tile_X11Y10_DO_SRAM15
  PIN Tile_X11Y10_DO_SRAM16
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1513.040 2435.000 1513.640 ;
    END
  END Tile_X11Y10_DO_SRAM16
  PIN Tile_X11Y10_DO_SRAM17
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1509.640 2435.000 1510.240 ;
    END
  END Tile_X11Y10_DO_SRAM17
  PIN Tile_X11Y10_DO_SRAM18
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1567.440 2435.000 1568.040 ;
    END
  END Tile_X11Y10_DO_SRAM18
  PIN Tile_X11Y10_DO_SRAM19
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1506.240 2435.000 1506.840 ;
    END
  END Tile_X11Y10_DO_SRAM19
  PIN Tile_X11Y10_DO_SRAM2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1540.240 2435.000 1540.840 ;
    END
  END Tile_X11Y10_DO_SRAM2
  PIN Tile_X11Y10_DO_SRAM20
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1570.840 2435.000 1571.440 ;
    END
  END Tile_X11Y10_DO_SRAM20
  PIN Tile_X11Y10_DO_SRAM21
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1502.840 2435.000 1503.440 ;
    END
  END Tile_X11Y10_DO_SRAM21
  PIN Tile_X11Y10_DO_SRAM22
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1499.440 2435.000 1500.040 ;
    END
  END Tile_X11Y10_DO_SRAM22
  PIN Tile_X11Y10_DO_SRAM23
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1574.240 2435.000 1574.840 ;
    END
  END Tile_X11Y10_DO_SRAM23
  PIN Tile_X11Y10_DO_SRAM24
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1496.040 2435.000 1496.640 ;
    END
  END Tile_X11Y10_DO_SRAM24
  PIN Tile_X11Y10_DO_SRAM25
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1577.640 2435.000 1578.240 ;
    END
  END Tile_X11Y10_DO_SRAM25
  PIN Tile_X11Y10_DO_SRAM26
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1492.640 2435.000 1493.240 ;
    END
  END Tile_X11Y10_DO_SRAM26
  PIN Tile_X11Y10_DO_SRAM27
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1489.240 2435.000 1489.840 ;
    END
  END Tile_X11Y10_DO_SRAM27
  PIN Tile_X11Y10_DO_SRAM28
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1581.040 2435.000 1581.640 ;
    END
  END Tile_X11Y10_DO_SRAM28
  PIN Tile_X11Y10_DO_SRAM29
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1485.840 2435.000 1486.440 ;
    END
  END Tile_X11Y10_DO_SRAM29
  PIN Tile_X11Y10_DO_SRAM3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1547.040 2435.000 1547.640 ;
    END
  END Tile_X11Y10_DO_SRAM3
  PIN Tile_X11Y10_DO_SRAM30
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1584.440 2435.000 1585.040 ;
    END
  END Tile_X11Y10_DO_SRAM30
  PIN Tile_X11Y10_DO_SRAM31
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1482.440 2435.000 1483.040 ;
    END
  END Tile_X11Y10_DO_SRAM31
  PIN Tile_X11Y10_DO_SRAM4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1536.840 2435.000 1537.440 ;
    END
  END Tile_X11Y10_DO_SRAM4
  PIN Tile_X11Y10_DO_SRAM5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1550.440 2435.000 1551.040 ;
    END
  END Tile_X11Y10_DO_SRAM5
  PIN Tile_X11Y10_DO_SRAM6
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1533.440 2435.000 1534.040 ;
    END
  END Tile_X11Y10_DO_SRAM6
  PIN Tile_X11Y10_DO_SRAM7
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1530.040 2435.000 1530.640 ;
    END
  END Tile_X11Y10_DO_SRAM7
  PIN Tile_X11Y10_DO_SRAM8
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1553.840 2435.000 1554.440 ;
    END
  END Tile_X11Y10_DO_SRAM8
  PIN Tile_X11Y10_DO_SRAM9
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1526.640 2435.000 1527.240 ;
    END
  END Tile_X11Y10_DO_SRAM9
  PIN Tile_X11Y10_EN_SRAM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1689.840 2435.000 1690.440 ;
    END
  END Tile_X11Y10_EN_SRAM
  PIN Tile_X11Y10_R_WB_SRAM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1710.240 2435.000 1710.840 ;
    END
  END Tile_X11Y10_R_WB_SRAM
  PIN Tile_X11Y12_AD_SRAM0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 982.640 2435.000 983.240 ;
    END
  END Tile_X11Y12_AD_SRAM0
  PIN Tile_X11Y12_AD_SRAM1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1026.840 2435.000 1027.440 ;
    END
  END Tile_X11Y12_AD_SRAM1
  PIN Tile_X11Y12_AD_SRAM2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1139.040 2435.000 1139.640 ;
    END
  END Tile_X11Y12_AD_SRAM2
  PIN Tile_X11Y12_AD_SRAM3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1023.440 2435.000 1024.040 ;
    END
  END Tile_X11Y12_AD_SRAM3
  PIN Tile_X11Y12_AD_SRAM4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1142.440 2435.000 1143.040 ;
    END
  END Tile_X11Y12_AD_SRAM4
  PIN Tile_X11Y12_AD_SRAM5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1020.040 2435.000 1020.640 ;
    END
  END Tile_X11Y12_AD_SRAM5
  PIN Tile_X11Y12_AD_SRAM6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1016.640 2435.000 1017.240 ;
    END
  END Tile_X11Y12_AD_SRAM6
  PIN Tile_X11Y12_AD_SRAM7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1145.840 2435.000 1146.440 ;
    END
  END Tile_X11Y12_AD_SRAM7
  PIN Tile_X11Y12_AD_SRAM8
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1013.240 2435.000 1013.840 ;
    END
  END Tile_X11Y12_AD_SRAM8
  PIN Tile_X11Y12_AD_SRAM9
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1149.240 2435.000 1149.840 ;
    END
  END Tile_X11Y12_AD_SRAM9
  PIN Tile_X11Y12_BEN_SRAM0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1009.840 2435.000 1010.440 ;
    END
  END Tile_X11Y12_BEN_SRAM0
  PIN Tile_X11Y12_BEN_SRAM1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1006.440 2435.000 1007.040 ;
    END
  END Tile_X11Y12_BEN_SRAM1
  PIN Tile_X11Y12_BEN_SRAM10
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1162.840 2435.000 1163.440 ;
    END
  END Tile_X11Y12_BEN_SRAM10
  PIN Tile_X11Y12_BEN_SRAM11
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 986.040 2435.000 986.640 ;
    END
  END Tile_X11Y12_BEN_SRAM11
  PIN Tile_X11Y12_BEN_SRAM12
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1166.240 2435.000 1166.840 ;
    END
  END Tile_X11Y12_BEN_SRAM12
  PIN Tile_X11Y12_BEN_SRAM13
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1169.640 2435.000 1170.240 ;
    END
  END Tile_X11Y12_BEN_SRAM13
  PIN Tile_X11Y12_BEN_SRAM14
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1349.840 2435.000 1350.440 ;
    END
  END Tile_X11Y12_BEN_SRAM14
  PIN Tile_X11Y12_BEN_SRAM15
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1346.440 2435.000 1347.040 ;
    END
  END Tile_X11Y12_BEN_SRAM15
  PIN Tile_X11Y12_BEN_SRAM16
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1173.040 2435.000 1173.640 ;
    END
  END Tile_X11Y12_BEN_SRAM16
  PIN Tile_X11Y12_BEN_SRAM17
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1343.040 2435.000 1343.640 ;
    END
  END Tile_X11Y12_BEN_SRAM17
  PIN Tile_X11Y12_BEN_SRAM18
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1176.440 2435.000 1177.040 ;
    END
  END Tile_X11Y12_BEN_SRAM18
  PIN Tile_X11Y12_BEN_SRAM19
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1339.640 2435.000 1340.240 ;
    END
  END Tile_X11Y12_BEN_SRAM19
  PIN Tile_X11Y12_BEN_SRAM2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1152.640 2435.000 1153.240 ;
    END
  END Tile_X11Y12_BEN_SRAM2
  PIN Tile_X11Y12_BEN_SRAM20
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1336.240 2435.000 1336.840 ;
    END
  END Tile_X11Y12_BEN_SRAM20
  PIN Tile_X11Y12_BEN_SRAM21
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1179.840 2435.000 1180.440 ;
    END
  END Tile_X11Y12_BEN_SRAM21
  PIN Tile_X11Y12_BEN_SRAM22
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1332.840 2435.000 1333.440 ;
    END
  END Tile_X11Y12_BEN_SRAM22
  PIN Tile_X11Y12_BEN_SRAM23
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1183.240 2435.000 1183.840 ;
    END
  END Tile_X11Y12_BEN_SRAM23
  PIN Tile_X11Y12_BEN_SRAM24
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1329.440 2435.000 1330.040 ;
    END
  END Tile_X11Y12_BEN_SRAM24
  PIN Tile_X11Y12_BEN_SRAM25
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1326.040 2435.000 1326.640 ;
    END
  END Tile_X11Y12_BEN_SRAM25
  PIN Tile_X11Y12_BEN_SRAM26
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1186.640 2435.000 1187.240 ;
    END
  END Tile_X11Y12_BEN_SRAM26
  PIN Tile_X11Y12_BEN_SRAM27
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1322.640 2435.000 1323.240 ;
    END
  END Tile_X11Y12_BEN_SRAM27
  PIN Tile_X11Y12_BEN_SRAM28
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1190.040 2435.000 1190.640 ;
    END
  END Tile_X11Y12_BEN_SRAM28
  PIN Tile_X11Y12_BEN_SRAM29
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1319.240 2435.000 1319.840 ;
    END
  END Tile_X11Y12_BEN_SRAM29
  PIN Tile_X11Y12_BEN_SRAM3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1003.040 2435.000 1003.640 ;
    END
  END Tile_X11Y12_BEN_SRAM3
  PIN Tile_X11Y12_BEN_SRAM30
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1315.840 2435.000 1316.440 ;
    END
  END Tile_X11Y12_BEN_SRAM30
  PIN Tile_X11Y12_BEN_SRAM31
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1193.440 2435.000 1194.040 ;
    END
  END Tile_X11Y12_BEN_SRAM31
  PIN Tile_X11Y12_BEN_SRAM4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1156.040 2435.000 1156.640 ;
    END
  END Tile_X11Y12_BEN_SRAM4
  PIN Tile_X11Y12_BEN_SRAM5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 999.640 2435.000 1000.240 ;
    END
  END Tile_X11Y12_BEN_SRAM5
  PIN Tile_X11Y12_BEN_SRAM6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 996.240 2435.000 996.840 ;
    END
  END Tile_X11Y12_BEN_SRAM6
  PIN Tile_X11Y12_BEN_SRAM7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1159.440 2435.000 1160.040 ;
    END
  END Tile_X11Y12_BEN_SRAM7
  PIN Tile_X11Y12_BEN_SRAM8
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 992.840 2435.000 993.440 ;
    END
  END Tile_X11Y12_BEN_SRAM8
  PIN Tile_X11Y12_BEN_SRAM9
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 989.440 2435.000 990.040 ;
    END
  END Tile_X11Y12_BEN_SRAM9
  PIN Tile_X11Y12_CLOCK_SRAM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1312.440 2435.000 1313.040 ;
    END
  END Tile_X11Y12_CLOCK_SRAM
  PIN Tile_X11Y12_DI_SRAM0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1196.840 2435.000 1197.440 ;
    END
  END Tile_X11Y12_DI_SRAM0
  PIN Tile_X11Y12_DI_SRAM1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1309.040 2435.000 1309.640 ;
    END
  END Tile_X11Y12_DI_SRAM1
  PIN Tile_X11Y12_DI_SRAM10
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1305.640 2435.000 1306.240 ;
    END
  END Tile_X11Y12_DI_SRAM10
  PIN Tile_X11Y12_DI_SRAM11
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1288.640 2435.000 1289.240 ;
    END
  END Tile_X11Y12_DI_SRAM11
  PIN Tile_X11Y12_DI_SRAM12
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1285.240 2435.000 1285.840 ;
    END
  END Tile_X11Y12_DI_SRAM12
  PIN Tile_X11Y12_DI_SRAM13
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1224.040 2435.000 1224.640 ;
    END
  END Tile_X11Y12_DI_SRAM13
  PIN Tile_X11Y12_DI_SRAM14
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1281.840 2435.000 1282.440 ;
    END
  END Tile_X11Y12_DI_SRAM14
  PIN Tile_X11Y12_DI_SRAM15
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1227.440 2435.000 1228.040 ;
    END
  END Tile_X11Y12_DI_SRAM15
  PIN Tile_X11Y12_DI_SRAM16
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1302.240 2435.000 1302.840 ;
    END
  END Tile_X11Y12_DI_SRAM16
  PIN Tile_X11Y12_DI_SRAM17
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1275.040 2435.000 1275.640 ;
    END
  END Tile_X11Y12_DI_SRAM17
  PIN Tile_X11Y12_DI_SRAM18
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1298.840 2435.000 1299.440 ;
    END
  END Tile_X11Y12_DI_SRAM18
  PIN Tile_X11Y12_DI_SRAM19
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1271.640 2435.000 1272.240 ;
    END
  END Tile_X11Y12_DI_SRAM19
  PIN Tile_X11Y12_DI_SRAM2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1200.240 2435.000 1200.840 ;
    END
  END Tile_X11Y12_DI_SRAM2
  PIN Tile_X11Y12_DI_SRAM20
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1230.840 2435.000 1231.440 ;
    END
  END Tile_X11Y12_DI_SRAM20
  PIN Tile_X11Y12_DI_SRAM21
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1268.240 2435.000 1268.840 ;
    END
  END Tile_X11Y12_DI_SRAM21
  PIN Tile_X11Y12_DI_SRAM22
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1264.840 2435.000 1265.440 ;
    END
  END Tile_X11Y12_DI_SRAM22
  PIN Tile_X11Y12_DI_SRAM23
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1234.240 2435.000 1234.840 ;
    END
  END Tile_X11Y12_DI_SRAM23
  PIN Tile_X11Y12_DI_SRAM24
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1295.440 2435.000 1296.040 ;
    END
  END Tile_X11Y12_DI_SRAM24
  PIN Tile_X11Y12_DI_SRAM25
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1237.640 2435.000 1238.240 ;
    END
  END Tile_X11Y12_DI_SRAM25
  PIN Tile_X11Y12_DI_SRAM26
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1292.040 2435.000 1292.640 ;
    END
  END Tile_X11Y12_DI_SRAM26
  PIN Tile_X11Y12_DI_SRAM27
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1254.640 2435.000 1255.240 ;
    END
  END Tile_X11Y12_DI_SRAM27
  PIN Tile_X11Y12_DI_SRAM28
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1241.040 2435.000 1241.640 ;
    END
  END Tile_X11Y12_DI_SRAM28
  PIN Tile_X11Y12_DI_SRAM29
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1251.240 2435.000 1251.840 ;
    END
  END Tile_X11Y12_DI_SRAM29
  PIN Tile_X11Y12_DI_SRAM3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1203.640 2435.000 1204.240 ;
    END
  END Tile_X11Y12_DI_SRAM3
  PIN Tile_X11Y12_DI_SRAM30
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1244.440 2435.000 1245.040 ;
    END
  END Tile_X11Y12_DI_SRAM30
  PIN Tile_X11Y12_DI_SRAM31
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1247.840 2435.000 1248.440 ;
    END
  END Tile_X11Y12_DI_SRAM31
  PIN Tile_X11Y12_DI_SRAM4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1207.040 2435.000 1207.640 ;
    END
  END Tile_X11Y12_DI_SRAM4
  PIN Tile_X11Y12_DI_SRAM5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1210.440 2435.000 1211.040 ;
    END
  END Tile_X11Y12_DI_SRAM5
  PIN Tile_X11Y12_DI_SRAM6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1213.840 2435.000 1214.440 ;
    END
  END Tile_X11Y12_DI_SRAM6
  PIN Tile_X11Y12_DI_SRAM7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1217.240 2435.000 1217.840 ;
    END
  END Tile_X11Y12_DI_SRAM7
  PIN Tile_X11Y12_DI_SRAM8
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1220.640 2435.000 1221.240 ;
    END
  END Tile_X11Y12_DI_SRAM8
  PIN Tile_X11Y12_DI_SRAM9
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1278.440 2435.000 1279.040 ;
    END
  END Tile_X11Y12_DI_SRAM9
  PIN Tile_X11Y12_DO_SRAM0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1030.240 2435.000 1030.840 ;
    END
  END Tile_X11Y12_DO_SRAM0
  PIN Tile_X11Y12_DO_SRAM1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1094.840 2435.000 1095.440 ;
    END
  END Tile_X11Y12_DO_SRAM1
  PIN Tile_X11Y12_DO_SRAM10
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1074.440 2435.000 1075.040 ;
    END
  END Tile_X11Y12_DO_SRAM10
  PIN Tile_X11Y12_DO_SRAM11
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1108.440 2435.000 1109.040 ;
    END
  END Tile_X11Y12_DO_SRAM11
  PIN Tile_X11Y12_DO_SRAM12
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1071.040 2435.000 1071.640 ;
    END
  END Tile_X11Y12_DO_SRAM12
  PIN Tile_X11Y12_DO_SRAM13
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1067.640 2435.000 1068.240 ;
    END
  END Tile_X11Y12_DO_SRAM13
  PIN Tile_X11Y12_DO_SRAM14
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1111.840 2435.000 1112.440 ;
    END
  END Tile_X11Y12_DO_SRAM14
  PIN Tile_X11Y12_DO_SRAM15
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1064.240 2435.000 1064.840 ;
    END
  END Tile_X11Y12_DO_SRAM15
  PIN Tile_X11Y12_DO_SRAM16
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1115.240 2435.000 1115.840 ;
    END
  END Tile_X11Y12_DO_SRAM16
  PIN Tile_X11Y12_DO_SRAM17
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1060.840 2435.000 1061.440 ;
    END
  END Tile_X11Y12_DO_SRAM17
  PIN Tile_X11Y12_DO_SRAM18
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1057.440 2435.000 1058.040 ;
    END
  END Tile_X11Y12_DO_SRAM18
  PIN Tile_X11Y12_DO_SRAM19
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1118.640 2435.000 1119.240 ;
    END
  END Tile_X11Y12_DO_SRAM19
  PIN Tile_X11Y12_DO_SRAM2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1091.440 2435.000 1092.040 ;
    END
  END Tile_X11Y12_DO_SRAM2
  PIN Tile_X11Y12_DO_SRAM20
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1054.040 2435.000 1054.640 ;
    END
  END Tile_X11Y12_DO_SRAM20
  PIN Tile_X11Y12_DO_SRAM21
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1122.040 2435.000 1122.640 ;
    END
  END Tile_X11Y12_DO_SRAM21
  PIN Tile_X11Y12_DO_SRAM22
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1050.640 2435.000 1051.240 ;
    END
  END Tile_X11Y12_DO_SRAM22
  PIN Tile_X11Y12_DO_SRAM23
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1047.240 2435.000 1047.840 ;
    END
  END Tile_X11Y12_DO_SRAM23
  PIN Tile_X11Y12_DO_SRAM24
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1125.440 2435.000 1126.040 ;
    END
  END Tile_X11Y12_DO_SRAM24
  PIN Tile_X11Y12_DO_SRAM25
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1043.840 2435.000 1044.440 ;
    END
  END Tile_X11Y12_DO_SRAM25
  PIN Tile_X11Y12_DO_SRAM26
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1128.840 2435.000 1129.440 ;
    END
  END Tile_X11Y12_DO_SRAM26
  PIN Tile_X11Y12_DO_SRAM27
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1040.440 2435.000 1041.040 ;
    END
  END Tile_X11Y12_DO_SRAM27
  PIN Tile_X11Y12_DO_SRAM28
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1037.040 2435.000 1037.640 ;
    END
  END Tile_X11Y12_DO_SRAM28
  PIN Tile_X11Y12_DO_SRAM29
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1132.240 2435.000 1132.840 ;
    END
  END Tile_X11Y12_DO_SRAM29
  PIN Tile_X11Y12_DO_SRAM3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1088.040 2435.000 1088.640 ;
    END
  END Tile_X11Y12_DO_SRAM3
  PIN Tile_X11Y12_DO_SRAM30
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1033.640 2435.000 1034.240 ;
    END
  END Tile_X11Y12_DO_SRAM30
  PIN Tile_X11Y12_DO_SRAM31
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1135.640 2435.000 1136.240 ;
    END
  END Tile_X11Y12_DO_SRAM31
  PIN Tile_X11Y12_DO_SRAM4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1098.240 2435.000 1098.840 ;
    END
  END Tile_X11Y12_DO_SRAM4
  PIN Tile_X11Y12_DO_SRAM5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1084.640 2435.000 1085.240 ;
    END
  END Tile_X11Y12_DO_SRAM5
  PIN Tile_X11Y12_DO_SRAM6
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1101.640 2435.000 1102.240 ;
    END
  END Tile_X11Y12_DO_SRAM6
  PIN Tile_X11Y12_DO_SRAM7
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1081.240 2435.000 1081.840 ;
    END
  END Tile_X11Y12_DO_SRAM7
  PIN Tile_X11Y12_DO_SRAM8
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1077.840 2435.000 1078.440 ;
    END
  END Tile_X11Y12_DO_SRAM8
  PIN Tile_X11Y12_DO_SRAM9
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1105.040 2435.000 1105.640 ;
    END
  END Tile_X11Y12_DO_SRAM9
  PIN Tile_X11Y12_EN_SRAM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1261.440 2435.000 1262.040 ;
    END
  END Tile_X11Y12_EN_SRAM
  PIN Tile_X11Y12_R_WB_SRAM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1258.040 2435.000 1258.640 ;
    END
  END Tile_X11Y12_R_WB_SRAM
  PIN Tile_X11Y14_AD_SRAM0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 962.240 2435.000 962.840 ;
    END
  END Tile_X11Y14_AD_SRAM0
  PIN Tile_X11Y14_AD_SRAM1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 945.240 2435.000 945.840 ;
    END
  END Tile_X11Y14_AD_SRAM1
  PIN Tile_X11Y14_AD_SRAM2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 690.240 2435.000 690.840 ;
    END
  END Tile_X11Y14_AD_SRAM2
  PIN Tile_X11Y14_AD_SRAM3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 941.840 2435.000 942.440 ;
    END
  END Tile_X11Y14_AD_SRAM3
  PIN Tile_X11Y14_AD_SRAM4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 744.640 2435.000 745.240 ;
    END
  END Tile_X11Y14_AD_SRAM4
  PIN Tile_X11Y14_AD_SRAM5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 938.440 2435.000 939.040 ;
    END
  END Tile_X11Y14_AD_SRAM5
  PIN Tile_X11Y14_AD_SRAM6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 935.040 2435.000 935.640 ;
    END
  END Tile_X11Y14_AD_SRAM6
  PIN Tile_X11Y14_AD_SRAM7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 697.040 2435.000 697.640 ;
    END
  END Tile_X11Y14_AD_SRAM7
  PIN Tile_X11Y14_AD_SRAM8
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 931.640 2435.000 932.240 ;
    END
  END Tile_X11Y14_AD_SRAM8
  PIN Tile_X11Y14_AD_SRAM9
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 700.440 2435.000 701.040 ;
    END
  END Tile_X11Y14_AD_SRAM9
  PIN Tile_X11Y14_BEN_SRAM0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 928.240 2435.000 928.840 ;
    END
  END Tile_X11Y14_BEN_SRAM0
  PIN Tile_X11Y14_BEN_SRAM1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 924.840 2435.000 925.440 ;
    END
  END Tile_X11Y14_BEN_SRAM1
  PIN Tile_X11Y14_BEN_SRAM10
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 921.440 2435.000 922.040 ;
    END
  END Tile_X11Y14_BEN_SRAM10
  PIN Tile_X11Y14_BEN_SRAM11
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 904.440 2435.000 905.040 ;
    END
  END Tile_X11Y14_BEN_SRAM11
  PIN Tile_X11Y14_BEN_SRAM12
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 727.640 2435.000 728.240 ;
    END
  END Tile_X11Y14_BEN_SRAM12
  PIN Tile_X11Y14_BEN_SRAM13
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 901.040 2435.000 901.640 ;
    END
  END Tile_X11Y14_BEN_SRAM13
  PIN Tile_X11Y14_BEN_SRAM14
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 731.040 2435.000 731.640 ;
    END
  END Tile_X11Y14_BEN_SRAM14
  PIN Tile_X11Y14_BEN_SRAM15
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 897.640 2435.000 898.240 ;
    END
  END Tile_X11Y14_BEN_SRAM15
  PIN Tile_X11Y14_BEN_SRAM16
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 958.840 2435.000 959.440 ;
    END
  END Tile_X11Y14_BEN_SRAM16
  PIN Tile_X11Y14_BEN_SRAM17
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 724.240 2435.000 724.840 ;
    END
  END Tile_X11Y14_BEN_SRAM17
  PIN Tile_X11Y14_BEN_SRAM18
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 890.840 2435.000 891.440 ;
    END
  END Tile_X11Y14_BEN_SRAM18
  PIN Tile_X11Y14_BEN_SRAM19
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 955.440 2435.000 956.040 ;
    END
  END Tile_X11Y14_BEN_SRAM19
  PIN Tile_X11Y14_BEN_SRAM2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 703.840 2435.000 704.440 ;
    END
  END Tile_X11Y14_BEN_SRAM2
  PIN Tile_X11Y14_BEN_SRAM20
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 887.440 2435.000 888.040 ;
    END
  END Tile_X11Y14_BEN_SRAM20
  PIN Tile_X11Y14_BEN_SRAM21
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 884.040 2435.000 884.640 ;
    END
  END Tile_X11Y14_BEN_SRAM21
  PIN Tile_X11Y14_BEN_SRAM22
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 952.040 2435.000 952.640 ;
    END
  END Tile_X11Y14_BEN_SRAM22
  PIN Tile_X11Y14_BEN_SRAM23
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 880.640 2435.000 881.240 ;
    END
  END Tile_X11Y14_BEN_SRAM23
  PIN Tile_X11Y14_BEN_SRAM24
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 741.240 2435.000 741.840 ;
    END
  END Tile_X11Y14_BEN_SRAM24
  PIN Tile_X11Y14_BEN_SRAM25
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 948.640 2435.000 949.240 ;
    END
  END Tile_X11Y14_BEN_SRAM25
  PIN Tile_X11Y14_BEN_SRAM26
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 873.840 2435.000 874.440 ;
    END
  END Tile_X11Y14_BEN_SRAM26
  PIN Tile_X11Y14_BEN_SRAM27
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 737.840 2435.000 738.440 ;
    END
  END Tile_X11Y14_BEN_SRAM27
  PIN Tile_X11Y14_BEN_SRAM28
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 870.440 2435.000 871.040 ;
    END
  END Tile_X11Y14_BEN_SRAM28
  PIN Tile_X11Y14_BEN_SRAM29
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 748.040 2435.000 748.640 ;
    END
  END Tile_X11Y14_BEN_SRAM29
  PIN Tile_X11Y14_BEN_SRAM3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 710.640 2435.000 711.240 ;
    END
  END Tile_X11Y14_BEN_SRAM3
  PIN Tile_X11Y14_BEN_SRAM30
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 867.040 2435.000 867.640 ;
    END
  END Tile_X11Y14_BEN_SRAM30
  PIN Tile_X11Y14_BEN_SRAM31
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 863.640 2435.000 864.240 ;
    END
  END Tile_X11Y14_BEN_SRAM31
  PIN Tile_X11Y14_BEN_SRAM4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 707.240 2435.000 707.840 ;
    END
  END Tile_X11Y14_BEN_SRAM4
  PIN Tile_X11Y14_BEN_SRAM5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 717.440 2435.000 718.040 ;
    END
  END Tile_X11Y14_BEN_SRAM5
  PIN Tile_X11Y14_BEN_SRAM6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 714.040 2435.000 714.640 ;
    END
  END Tile_X11Y14_BEN_SRAM6
  PIN Tile_X11Y14_BEN_SRAM7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 765.040 2435.000 765.640 ;
    END
  END Tile_X11Y14_BEN_SRAM7
  PIN Tile_X11Y14_BEN_SRAM8
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 751.440 2435.000 752.040 ;
    END
  END Tile_X11Y14_BEN_SRAM8
  PIN Tile_X11Y14_BEN_SRAM9
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 720.840 2435.000 721.440 ;
    END
  END Tile_X11Y14_BEN_SRAM9
  PIN Tile_X11Y14_CLOCK_SRAM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 805.840 2435.000 806.440 ;
    END
  END Tile_X11Y14_CLOCK_SRAM
  PIN Tile_X11Y14_DI_SRAM0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 860.240 2435.000 860.840 ;
    END
  END Tile_X11Y14_DI_SRAM0
  PIN Tile_X11Y14_DI_SRAM1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 768.440 2435.000 769.040 ;
    END
  END Tile_X11Y14_DI_SRAM1
  PIN Tile_X11Y14_DI_SRAM10
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 856.840 2435.000 857.440 ;
    END
  END Tile_X11Y14_DI_SRAM10
  PIN Tile_X11Y14_DI_SRAM11
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 771.840 2435.000 772.440 ;
    END
  END Tile_X11Y14_DI_SRAM11
  PIN Tile_X11Y14_DI_SRAM12
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 836.440 2435.000 837.040 ;
    END
  END Tile_X11Y14_DI_SRAM12
  PIN Tile_X11Y14_DI_SRAM13
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 833.040 2435.000 833.640 ;
    END
  END Tile_X11Y14_DI_SRAM13
  PIN Tile_X11Y14_DI_SRAM14
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 795.640 2435.000 796.240 ;
    END
  END Tile_X11Y14_DI_SRAM14
  PIN Tile_X11Y14_DI_SRAM15
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 829.640 2435.000 830.240 ;
    END
  END Tile_X11Y14_DI_SRAM15
  PIN Tile_X11Y14_DI_SRAM16
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 775.240 2435.000 775.840 ;
    END
  END Tile_X11Y14_DI_SRAM16
  PIN Tile_X11Y14_DI_SRAM17
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 826.240 2435.000 826.840 ;
    END
  END Tile_X11Y14_DI_SRAM17
  PIN Tile_X11Y14_DI_SRAM18
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 918.040 2435.000 918.640 ;
    END
  END Tile_X11Y14_DI_SRAM18
  PIN Tile_X11Y14_DI_SRAM19
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 778.640 2435.000 779.240 ;
    END
  END Tile_X11Y14_DI_SRAM19
  PIN Tile_X11Y14_DI_SRAM2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 792.240 2435.000 792.840 ;
    END
  END Tile_X11Y14_DI_SRAM2
  PIN Tile_X11Y14_DI_SRAM20
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 914.640 2435.000 915.240 ;
    END
  END Tile_X11Y14_DI_SRAM20
  PIN Tile_X11Y14_DI_SRAM21
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 839.840 2435.000 840.440 ;
    END
  END Tile_X11Y14_DI_SRAM21
  PIN Tile_X11Y14_DI_SRAM22
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 816.040 2435.000 816.640 ;
    END
  END Tile_X11Y14_DI_SRAM22
  PIN Tile_X11Y14_DI_SRAM23
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 812.640 2435.000 813.240 ;
    END
  END Tile_X11Y14_DI_SRAM23
  PIN Tile_X11Y14_DI_SRAM24
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 850.040 2435.000 850.640 ;
    END
  END Tile_X11Y14_DI_SRAM24
  PIN Tile_X11Y14_DI_SRAM25
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 809.240 2435.000 809.840 ;
    END
  END Tile_X11Y14_DI_SRAM25
  PIN Tile_X11Y14_DI_SRAM26
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 782.040 2435.000 782.640 ;
    END
  END Tile_X11Y14_DI_SRAM26
  PIN Tile_X11Y14_DI_SRAM27
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 843.240 2435.000 843.840 ;
    END
  END Tile_X11Y14_DI_SRAM27
  PIN Tile_X11Y14_DI_SRAM28
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 802.440 2435.000 803.040 ;
    END
  END Tile_X11Y14_DI_SRAM28
  PIN Tile_X11Y14_DI_SRAM29
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 785.440 2435.000 786.040 ;
    END
  END Tile_X11Y14_DI_SRAM29
  PIN Tile_X11Y14_DI_SRAM3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 911.240 2435.000 911.840 ;
    END
  END Tile_X11Y14_DI_SRAM3
  PIN Tile_X11Y14_DI_SRAM30
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 799.040 2435.000 799.640 ;
    END
  END Tile_X11Y14_DI_SRAM30
  PIN Tile_X11Y14_DI_SRAM31
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 788.840 2435.000 789.440 ;
    END
  END Tile_X11Y14_DI_SRAM31
  PIN Tile_X11Y14_DI_SRAM4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 853.440 2435.000 854.040 ;
    END
  END Tile_X11Y14_DI_SRAM4
  PIN Tile_X11Y14_DI_SRAM5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 754.840 2435.000 755.440 ;
    END
  END Tile_X11Y14_DI_SRAM5
  PIN Tile_X11Y14_DI_SRAM6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 758.240 2435.000 758.840 ;
    END
  END Tile_X11Y14_DI_SRAM6
  PIN Tile_X11Y14_DI_SRAM7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 761.640 2435.000 762.240 ;
    END
  END Tile_X11Y14_DI_SRAM7
  PIN Tile_X11Y14_DI_SRAM8
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 907.840 2435.000 908.440 ;
    END
  END Tile_X11Y14_DI_SRAM8
  PIN Tile_X11Y14_DI_SRAM9
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 819.440 2435.000 820.040 ;
    END
  END Tile_X11Y14_DI_SRAM9
  PIN Tile_X11Y14_DO_SRAM0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 595.040 2435.000 595.640 ;
    END
  END Tile_X11Y14_DO_SRAM0
  PIN Tile_X11Y14_DO_SRAM1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 642.640 2435.000 643.240 ;
    END
  END Tile_X11Y14_DO_SRAM1
  PIN Tile_X11Y14_DO_SRAM10
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 656.240 2435.000 656.840 ;
    END
  END Tile_X11Y14_DO_SRAM10
  PIN Tile_X11Y14_DO_SRAM11
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 622.240 2435.000 622.840 ;
    END
  END Tile_X11Y14_DO_SRAM11
  PIN Tile_X11Y14_DO_SRAM12
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 659.640 2435.000 660.240 ;
    END
  END Tile_X11Y14_DO_SRAM12
  PIN Tile_X11Y14_DO_SRAM13
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 618.840 2435.000 619.440 ;
    END
  END Tile_X11Y14_DO_SRAM13
  PIN Tile_X11Y14_DO_SRAM14
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 615.440 2435.000 616.040 ;
    END
  END Tile_X11Y14_DO_SRAM14
  PIN Tile_X11Y14_DO_SRAM15
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 663.040 2435.000 663.640 ;
    END
  END Tile_X11Y14_DO_SRAM15
  PIN Tile_X11Y14_DO_SRAM16
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 612.040 2435.000 612.640 ;
    END
  END Tile_X11Y14_DO_SRAM16
  PIN Tile_X11Y14_DO_SRAM17
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 666.440 2435.000 667.040 ;
    END
  END Tile_X11Y14_DO_SRAM17
  PIN Tile_X11Y14_DO_SRAM18
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 608.640 2435.000 609.240 ;
    END
  END Tile_X11Y14_DO_SRAM18
  PIN Tile_X11Y14_DO_SRAM19
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 605.240 2435.000 605.840 ;
    END
  END Tile_X11Y14_DO_SRAM19
  PIN Tile_X11Y14_DO_SRAM2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 646.040 2435.000 646.640 ;
    END
  END Tile_X11Y14_DO_SRAM2
  PIN Tile_X11Y14_DO_SRAM20
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 669.840 2435.000 670.440 ;
    END
  END Tile_X11Y14_DO_SRAM20
  PIN Tile_X11Y14_DO_SRAM21
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 601.840 2435.000 602.440 ;
    END
  END Tile_X11Y14_DO_SRAM21
  PIN Tile_X11Y14_DO_SRAM22
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 673.240 2435.000 673.840 ;
    END
  END Tile_X11Y14_DO_SRAM22
  PIN Tile_X11Y14_DO_SRAM23
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 598.440 2435.000 599.040 ;
    END
  END Tile_X11Y14_DO_SRAM23
  PIN Tile_X11Y14_DO_SRAM24
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 676.640 2435.000 677.240 ;
    END
  END Tile_X11Y14_DO_SRAM24
  PIN Tile_X11Y14_DO_SRAM25
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 680.040 2435.000 680.640 ;
    END
  END Tile_X11Y14_DO_SRAM25
  PIN Tile_X11Y14_DO_SRAM26
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 734.440 2435.000 735.040 ;
    END
  END Tile_X11Y14_DO_SRAM26
  PIN Tile_X11Y14_DO_SRAM27
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 894.240 2435.000 894.840 ;
    END
  END Tile_X11Y14_DO_SRAM27
  PIN Tile_X11Y14_DO_SRAM28
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 686.840 2435.000 687.440 ;
    END
  END Tile_X11Y14_DO_SRAM28
  PIN Tile_X11Y14_DO_SRAM29
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 683.440 2435.000 684.040 ;
    END
  END Tile_X11Y14_DO_SRAM29
  PIN Tile_X11Y14_DO_SRAM3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 639.240 2435.000 639.840 ;
    END
  END Tile_X11Y14_DO_SRAM3
  PIN Tile_X11Y14_DO_SRAM30
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 693.640 2435.000 694.240 ;
    END
  END Tile_X11Y14_DO_SRAM30
  PIN Tile_X11Y14_DO_SRAM31
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 877.240 2435.000 877.840 ;
    END
  END Tile_X11Y14_DO_SRAM31
  PIN Tile_X11Y14_DO_SRAM4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 635.840 2435.000 636.440 ;
    END
  END Tile_X11Y14_DO_SRAM4
  PIN Tile_X11Y14_DO_SRAM5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 649.440 2435.000 650.040 ;
    END
  END Tile_X11Y14_DO_SRAM5
  PIN Tile_X11Y14_DO_SRAM6
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 632.440 2435.000 633.040 ;
    END
  END Tile_X11Y14_DO_SRAM6
  PIN Tile_X11Y14_DO_SRAM7
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 652.840 2435.000 653.440 ;
    END
  END Tile_X11Y14_DO_SRAM7
  PIN Tile_X11Y14_DO_SRAM8
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 629.040 2435.000 629.640 ;
    END
  END Tile_X11Y14_DO_SRAM8
  PIN Tile_X11Y14_DO_SRAM9
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 625.640 2435.000 626.240 ;
    END
  END Tile_X11Y14_DO_SRAM9
  PIN Tile_X11Y14_EN_SRAM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 846.640 2435.000 847.240 ;
    END
  END Tile_X11Y14_EN_SRAM
  PIN Tile_X11Y14_R_WB_SRAM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 822.840 2435.000 823.440 ;
    END
  END Tile_X11Y14_R_WB_SRAM
  PIN Tile_X11Y16_AD_SRAM0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 85.040 2435.000 85.640 ;
    END
  END Tile_X11Y16_AD_SRAM0
  PIN Tile_X11Y16_AD_SRAM1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 238.040 2435.000 238.640 ;
    END
  END Tile_X11Y16_AD_SRAM1
  PIN Tile_X11Y16_AD_SRAM2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 125.840 2435.000 126.440 ;
    END
  END Tile_X11Y16_AD_SRAM2
  PIN Tile_X11Y16_AD_SRAM3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 122.440 2435.000 123.040 ;
    END
  END Tile_X11Y16_AD_SRAM3
  PIN Tile_X11Y16_AD_SRAM4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 241.440 2435.000 242.040 ;
    END
  END Tile_X11Y16_AD_SRAM4
  PIN Tile_X11Y16_AD_SRAM5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 119.040 2435.000 119.640 ;
    END
  END Tile_X11Y16_AD_SRAM5
  PIN Tile_X11Y16_AD_SRAM6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 244.840 2435.000 245.440 ;
    END
  END Tile_X11Y16_AD_SRAM6
  PIN Tile_X11Y16_AD_SRAM7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 115.640 2435.000 116.240 ;
    END
  END Tile_X11Y16_AD_SRAM7
  PIN Tile_X11Y16_AD_SRAM8
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 112.240 2435.000 112.840 ;
    END
  END Tile_X11Y16_AD_SRAM8
  PIN Tile_X11Y16_AD_SRAM9
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 248.240 2435.000 248.840 ;
    END
  END Tile_X11Y16_AD_SRAM9
  PIN Tile_X11Y16_BEN_SRAM0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 108.840 2435.000 109.440 ;
    END
  END Tile_X11Y16_BEN_SRAM0
  PIN Tile_X11Y16_BEN_SRAM1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 251.640 2435.000 252.240 ;
    END
  END Tile_X11Y16_BEN_SRAM1
  PIN Tile_X11Y16_BEN_SRAM10
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 88.440 2435.000 89.040 ;
    END
  END Tile_X11Y16_BEN_SRAM10
  PIN Tile_X11Y16_BEN_SRAM11
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 265.240 2435.000 265.840 ;
    END
  END Tile_X11Y16_BEN_SRAM11
  PIN Tile_X11Y16_BEN_SRAM12
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 452.240 2435.000 452.840 ;
    END
  END Tile_X11Y16_BEN_SRAM12
  PIN Tile_X11Y16_BEN_SRAM13
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 268.640 2435.000 269.240 ;
    END
  END Tile_X11Y16_BEN_SRAM13
  PIN Tile_X11Y16_BEN_SRAM14
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 448.840 2435.000 449.440 ;
    END
  END Tile_X11Y16_BEN_SRAM14
  PIN Tile_X11Y16_BEN_SRAM15
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 272.040 2435.000 272.640 ;
    END
  END Tile_X11Y16_BEN_SRAM15
  PIN Tile_X11Y16_BEN_SRAM16
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 445.440 2435.000 446.040 ;
    END
  END Tile_X11Y16_BEN_SRAM16
  PIN Tile_X11Y16_BEN_SRAM17
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 442.040 2435.000 442.640 ;
    END
  END Tile_X11Y16_BEN_SRAM17
  PIN Tile_X11Y16_BEN_SRAM18
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 275.440 2435.000 276.040 ;
    END
  END Tile_X11Y16_BEN_SRAM18
  PIN Tile_X11Y16_BEN_SRAM19
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 438.640 2435.000 439.240 ;
    END
  END Tile_X11Y16_BEN_SRAM19
  PIN Tile_X11Y16_BEN_SRAM2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 105.440 2435.000 106.040 ;
    END
  END Tile_X11Y16_BEN_SRAM2
  PIN Tile_X11Y16_BEN_SRAM20
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 278.840 2435.000 279.440 ;
    END
  END Tile_X11Y16_BEN_SRAM20
  PIN Tile_X11Y16_BEN_SRAM21
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 435.240 2435.000 435.840 ;
    END
  END Tile_X11Y16_BEN_SRAM21
  PIN Tile_X11Y16_BEN_SRAM22
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 431.840 2435.000 432.440 ;
    END
  END Tile_X11Y16_BEN_SRAM22
  PIN Tile_X11Y16_BEN_SRAM23
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 282.240 2435.000 282.840 ;
    END
  END Tile_X11Y16_BEN_SRAM23
  PIN Tile_X11Y16_BEN_SRAM24
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 428.440 2435.000 429.040 ;
    END
  END Tile_X11Y16_BEN_SRAM24
  PIN Tile_X11Y16_BEN_SRAM25
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 285.640 2435.000 286.240 ;
    END
  END Tile_X11Y16_BEN_SRAM25
  PIN Tile_X11Y16_BEN_SRAM26
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 425.040 2435.000 425.640 ;
    END
  END Tile_X11Y16_BEN_SRAM26
  PIN Tile_X11Y16_BEN_SRAM27
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 421.640 2435.000 422.240 ;
    END
  END Tile_X11Y16_BEN_SRAM27
  PIN Tile_X11Y16_BEN_SRAM28
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 289.040 2435.000 289.640 ;
    END
  END Tile_X11Y16_BEN_SRAM28
  PIN Tile_X11Y16_BEN_SRAM29
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 418.240 2435.000 418.840 ;
    END
  END Tile_X11Y16_BEN_SRAM29
  PIN Tile_X11Y16_BEN_SRAM3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 102.040 2435.000 102.640 ;
    END
  END Tile_X11Y16_BEN_SRAM3
  PIN Tile_X11Y16_BEN_SRAM30
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 292.440 2435.000 293.040 ;
    END
  END Tile_X11Y16_BEN_SRAM30
  PIN Tile_X11Y16_BEN_SRAM31
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 414.840 2435.000 415.440 ;
    END
  END Tile_X11Y16_BEN_SRAM31
  PIN Tile_X11Y16_BEN_SRAM4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 255.040 2435.000 255.640 ;
    END
  END Tile_X11Y16_BEN_SRAM4
  PIN Tile_X11Y16_BEN_SRAM5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 98.640 2435.000 99.240 ;
    END
  END Tile_X11Y16_BEN_SRAM5
  PIN Tile_X11Y16_BEN_SRAM6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 258.440 2435.000 259.040 ;
    END
  END Tile_X11Y16_BEN_SRAM6
  PIN Tile_X11Y16_BEN_SRAM7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 95.240 2435.000 95.840 ;
    END
  END Tile_X11Y16_BEN_SRAM7
  PIN Tile_X11Y16_BEN_SRAM8
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 91.840 2435.000 92.440 ;
    END
  END Tile_X11Y16_BEN_SRAM8
  PIN Tile_X11Y16_BEN_SRAM9
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 261.840 2435.000 262.440 ;
    END
  END Tile_X11Y16_BEN_SRAM9
  PIN Tile_X11Y16_CLOCK_SRAM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 411.440 2435.000 412.040 ;
    END
  END Tile_X11Y16_CLOCK_SRAM
  PIN Tile_X11Y16_DI_SRAM0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 295.840 2435.000 296.440 ;
    END
  END Tile_X11Y16_DI_SRAM0
  PIN Tile_X11Y16_DI_SRAM1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 408.040 2435.000 408.640 ;
    END
  END Tile_X11Y16_DI_SRAM1
  PIN Tile_X11Y16_DI_SRAM10
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 404.640 2435.000 405.240 ;
    END
  END Tile_X11Y16_DI_SRAM10
  PIN Tile_X11Y16_DI_SRAM11
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 401.240 2435.000 401.840 ;
    END
  END Tile_X11Y16_DI_SRAM11
  PIN Tile_X11Y16_DI_SRAM12
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 326.440 2435.000 327.040 ;
    END
  END Tile_X11Y16_DI_SRAM12
  PIN Tile_X11Y16_DI_SRAM13
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 384.240 2435.000 384.840 ;
    END
  END Tile_X11Y16_DI_SRAM13
  PIN Tile_X11Y16_DI_SRAM14
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 380.840 2435.000 381.440 ;
    END
  END Tile_X11Y16_DI_SRAM14
  PIN Tile_X11Y16_DI_SRAM15
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 319.640 2435.000 320.240 ;
    END
  END Tile_X11Y16_DI_SRAM15
  PIN Tile_X11Y16_DI_SRAM16
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 377.440 2435.000 378.040 ;
    END
  END Tile_X11Y16_DI_SRAM16
  PIN Tile_X11Y16_DI_SRAM17
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 329.840 2435.000 330.440 ;
    END
  END Tile_X11Y16_DI_SRAM17
  PIN Tile_X11Y16_DI_SRAM18
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 397.840 2435.000 398.440 ;
    END
  END Tile_X11Y16_DI_SRAM18
  PIN Tile_X11Y16_DI_SRAM19
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 370.640 2435.000 371.240 ;
    END
  END Tile_X11Y16_DI_SRAM19
  PIN Tile_X11Y16_DI_SRAM2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 299.240 2435.000 299.840 ;
    END
  END Tile_X11Y16_DI_SRAM2
  PIN Tile_X11Y16_DI_SRAM20
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 336.640 2435.000 337.240 ;
    END
  END Tile_X11Y16_DI_SRAM20
  PIN Tile_X11Y16_DI_SRAM21
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 367.240 2435.000 367.840 ;
    END
  END Tile_X11Y16_DI_SRAM21
  PIN Tile_X11Y16_DI_SRAM22
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 340.040 2435.000 340.640 ;
    END
  END Tile_X11Y16_DI_SRAM22
  PIN Tile_X11Y16_DI_SRAM23
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 394.440 2435.000 395.040 ;
    END
  END Tile_X11Y16_DI_SRAM23
  PIN Tile_X11Y16_DI_SRAM24
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 360.440 2435.000 361.040 ;
    END
  END Tile_X11Y16_DI_SRAM24
  PIN Tile_X11Y16_DI_SRAM25
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 333.240 2435.000 333.840 ;
    END
  END Tile_X11Y16_DI_SRAM25
  PIN Tile_X11Y16_DI_SRAM26
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 357.040 2435.000 357.640 ;
    END
  END Tile_X11Y16_DI_SRAM26
  PIN Tile_X11Y16_DI_SRAM27
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 391.040 2435.000 391.640 ;
    END
  END Tile_X11Y16_DI_SRAM27
  PIN Tile_X11Y16_DI_SRAM28
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 353.640 2435.000 354.240 ;
    END
  END Tile_X11Y16_DI_SRAM28
  PIN Tile_X11Y16_DI_SRAM29
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 350.240 2435.000 350.840 ;
    END
  END Tile_X11Y16_DI_SRAM29
  PIN Tile_X11Y16_DI_SRAM3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 302.640 2435.000 303.240 ;
    END
  END Tile_X11Y16_DI_SRAM3
  PIN Tile_X11Y16_DI_SRAM30
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 343.440 2435.000 344.040 ;
    END
  END Tile_X11Y16_DI_SRAM30
  PIN Tile_X11Y16_DI_SRAM31
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 346.840 2435.000 347.440 ;
    END
  END Tile_X11Y16_DI_SRAM31
  PIN Tile_X11Y16_DI_SRAM4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 316.240 2435.000 316.840 ;
    END
  END Tile_X11Y16_DI_SRAM4
  PIN Tile_X11Y16_DI_SRAM5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 309.440 2435.000 310.040 ;
    END
  END Tile_X11Y16_DI_SRAM5
  PIN Tile_X11Y16_DI_SRAM6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 312.840 2435.000 313.440 ;
    END
  END Tile_X11Y16_DI_SRAM6
  PIN Tile_X11Y16_DI_SRAM7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 306.040 2435.000 306.640 ;
    END
  END Tile_X11Y16_DI_SRAM7
  PIN Tile_X11Y16_DI_SRAM8
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 387.640 2435.000 388.240 ;
    END
  END Tile_X11Y16_DI_SRAM8
  PIN Tile_X11Y16_DI_SRAM9
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 323.040 2435.000 323.640 ;
    END
  END Tile_X11Y16_DI_SRAM9
  PIN Tile_X11Y16_DO_SRAM0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 129.240 2435.000 129.840 ;
    END
  END Tile_X11Y16_DO_SRAM0
  PIN Tile_X11Y16_DO_SRAM1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 193.840 2435.000 194.440 ;
    END
  END Tile_X11Y16_DO_SRAM1
  PIN Tile_X11Y16_DO_SRAM10
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 173.440 2435.000 174.040 ;
    END
  END Tile_X11Y16_DO_SRAM10
  PIN Tile_X11Y16_DO_SRAM11
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 207.440 2435.000 208.040 ;
    END
  END Tile_X11Y16_DO_SRAM11
  PIN Tile_X11Y16_DO_SRAM12
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 170.040 2435.000 170.640 ;
    END
  END Tile_X11Y16_DO_SRAM12
  PIN Tile_X11Y16_DO_SRAM13
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 210.840 2435.000 211.440 ;
    END
  END Tile_X11Y16_DO_SRAM13
  PIN Tile_X11Y16_DO_SRAM14
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 166.640 2435.000 167.240 ;
    END
  END Tile_X11Y16_DO_SRAM14
  PIN Tile_X11Y16_DO_SRAM15
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 163.240 2435.000 163.840 ;
    END
  END Tile_X11Y16_DO_SRAM15
  PIN Tile_X11Y16_DO_SRAM16
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 214.240 2435.000 214.840 ;
    END
  END Tile_X11Y16_DO_SRAM16
  PIN Tile_X11Y16_DO_SRAM17
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 159.840 2435.000 160.440 ;
    END
  END Tile_X11Y16_DO_SRAM17
  PIN Tile_X11Y16_DO_SRAM18
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 217.640 2435.000 218.240 ;
    END
  END Tile_X11Y16_DO_SRAM18
  PIN Tile_X11Y16_DO_SRAM19
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 156.440 2435.000 157.040 ;
    END
  END Tile_X11Y16_DO_SRAM19
  PIN Tile_X11Y16_DO_SRAM2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 190.440 2435.000 191.040 ;
    END
  END Tile_X11Y16_DO_SRAM2
  PIN Tile_X11Y16_DO_SRAM20
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 153.040 2435.000 153.640 ;
    END
  END Tile_X11Y16_DO_SRAM20
  PIN Tile_X11Y16_DO_SRAM21
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 221.040 2435.000 221.640 ;
    END
  END Tile_X11Y16_DO_SRAM21
  PIN Tile_X11Y16_DO_SRAM22
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 149.640 2435.000 150.240 ;
    END
  END Tile_X11Y16_DO_SRAM22
  PIN Tile_X11Y16_DO_SRAM23
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 224.440 2435.000 225.040 ;
    END
  END Tile_X11Y16_DO_SRAM23
  PIN Tile_X11Y16_DO_SRAM24
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 146.240 2435.000 146.840 ;
    END
  END Tile_X11Y16_DO_SRAM24
  PIN Tile_X11Y16_DO_SRAM25
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 142.840 2435.000 143.440 ;
    END
  END Tile_X11Y16_DO_SRAM25
  PIN Tile_X11Y16_DO_SRAM26
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 227.840 2435.000 228.440 ;
    END
  END Tile_X11Y16_DO_SRAM26
  PIN Tile_X11Y16_DO_SRAM27
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 139.440 2435.000 140.040 ;
    END
  END Tile_X11Y16_DO_SRAM27
  PIN Tile_X11Y16_DO_SRAM28
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 231.240 2435.000 231.840 ;
    END
  END Tile_X11Y16_DO_SRAM28
  PIN Tile_X11Y16_DO_SRAM29
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 136.040 2435.000 136.640 ;
    END
  END Tile_X11Y16_DO_SRAM29
  PIN Tile_X11Y16_DO_SRAM3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 197.240 2435.000 197.840 ;
    END
  END Tile_X11Y16_DO_SRAM3
  PIN Tile_X11Y16_DO_SRAM30
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 132.640 2435.000 133.240 ;
    END
  END Tile_X11Y16_DO_SRAM30
  PIN Tile_X11Y16_DO_SRAM31
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 234.640 2435.000 235.240 ;
    END
  END Tile_X11Y16_DO_SRAM31
  PIN Tile_X11Y16_DO_SRAM4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 187.040 2435.000 187.640 ;
    END
  END Tile_X11Y16_DO_SRAM4
  PIN Tile_X11Y16_DO_SRAM5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 183.640 2435.000 184.240 ;
    END
  END Tile_X11Y16_DO_SRAM5
  PIN Tile_X11Y16_DO_SRAM6
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 200.640 2435.000 201.240 ;
    END
  END Tile_X11Y16_DO_SRAM6
  PIN Tile_X11Y16_DO_SRAM7
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 180.240 2435.000 180.840 ;
    END
  END Tile_X11Y16_DO_SRAM7
  PIN Tile_X11Y16_DO_SRAM8
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 204.040 2435.000 204.640 ;
    END
  END Tile_X11Y16_DO_SRAM8
  PIN Tile_X11Y16_DO_SRAM9
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 176.840 2435.000 177.440 ;
    END
  END Tile_X11Y16_DO_SRAM9
  PIN Tile_X11Y16_EN_SRAM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 374.040 2435.000 374.640 ;
    END
  END Tile_X11Y16_EN_SRAM
  PIN Tile_X11Y16_R_WB_SRAM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 363.840 2435.000 364.440 ;
    END
  END Tile_X11Y16_R_WB_SRAM
  PIN Tile_X11Y2_AD_SRAM0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3767.240 2435.000 3767.840 ;
    END
  END Tile_X11Y2_AD_SRAM0
  PIN Tile_X11Y2_AD_SRAM1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3403.440 2435.000 3404.040 ;
    END
  END Tile_X11Y2_AD_SRAM1
  PIN Tile_X11Y2_AD_SRAM2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3695.840 2435.000 3696.440 ;
    END
  END Tile_X11Y2_AD_SRAM2
  PIN Tile_X11Y2_AD_SRAM3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3474.840 2435.000 3475.440 ;
    END
  END Tile_X11Y2_AD_SRAM3
  PIN Tile_X11Y2_AD_SRAM4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3743.440 2435.000 3744.040 ;
    END
  END Tile_X11Y2_AD_SRAM4
  PIN Tile_X11Y2_AD_SRAM5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3621.040 2435.000 3621.640 ;
    END
  END Tile_X11Y2_AD_SRAM5
  PIN Tile_X11Y2_AD_SRAM6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3536.040 2435.000 3536.640 ;
    END
  END Tile_X11Y2_AD_SRAM6
  PIN Tile_X11Y2_AD_SRAM7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3457.840 2435.000 3458.440 ;
    END
  END Tile_X11Y2_AD_SRAM7
  PIN Tile_X11Y2_AD_SRAM8
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3699.240 2435.000 3699.840 ;
    END
  END Tile_X11Y2_AD_SRAM8
  PIN Tile_X11Y2_AD_SRAM9
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3634.640 2435.000 3635.240 ;
    END
  END Tile_X11Y2_AD_SRAM9
  PIN Tile_X11Y2_BEN_SRAM0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3757.040 2435.000 3757.640 ;
    END
  END Tile_X11Y2_BEN_SRAM0
  PIN Tile_X11Y2_BEN_SRAM1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3427.240 2435.000 3427.840 ;
    END
  END Tile_X11Y2_BEN_SRAM1
  PIN Tile_X11Y2_BEN_SRAM10
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3624.440 2435.000 3625.040 ;
    END
  END Tile_X11Y2_BEN_SRAM10
  PIN Tile_X11Y2_BEN_SRAM11
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3454.440 2435.000 3455.040 ;
    END
  END Tile_X11Y2_BEN_SRAM11
  PIN Tile_X11Y2_BEN_SRAM12
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3610.840 2435.000 3611.440 ;
    END
  END Tile_X11Y2_BEN_SRAM12
  PIN Tile_X11Y2_BEN_SRAM13
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3702.640 2435.000 3703.240 ;
    END
  END Tile_X11Y2_BEN_SRAM13
  PIN Tile_X11Y2_BEN_SRAM14
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3502.040 2435.000 3502.640 ;
    END
  END Tile_X11Y2_BEN_SRAM14
  PIN Tile_X11Y2_BEN_SRAM15
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3746.840 2435.000 3747.440 ;
    END
  END Tile_X11Y2_BEN_SRAM15
  PIN Tile_X11Y2_BEN_SRAM16
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3430.640 2435.000 3431.240 ;
    END
  END Tile_X11Y2_BEN_SRAM16
  PIN Tile_X11Y2_BEN_SRAM17
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3706.040 2435.000 3706.640 ;
    END
  END Tile_X11Y2_BEN_SRAM17
  PIN Tile_X11Y2_BEN_SRAM18
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3590.440 2435.000 3591.040 ;
    END
  END Tile_X11Y2_BEN_SRAM18
  PIN Tile_X11Y2_BEN_SRAM19
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3512.240 2435.000 3512.840 ;
    END
  END Tile_X11Y2_BEN_SRAM19
  PIN Tile_X11Y2_BEN_SRAM2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3464.640 2435.000 3465.240 ;
    END
  END Tile_X11Y2_BEN_SRAM2
  PIN Tile_X11Y2_BEN_SRAM20
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3587.040 2435.000 3587.640 ;
    END
  END Tile_X11Y2_BEN_SRAM20
  PIN Tile_X11Y2_BEN_SRAM21
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3709.440 2435.000 3710.040 ;
    END
  END Tile_X11Y2_BEN_SRAM21
  PIN Tile_X11Y2_BEN_SRAM22
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3648.240 2435.000 3648.840 ;
    END
  END Tile_X11Y2_BEN_SRAM22
  PIN Tile_X11Y2_BEN_SRAM23
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3580.240 2435.000 3580.840 ;
    END
  END Tile_X11Y2_BEN_SRAM23
  PIN Tile_X11Y2_BEN_SRAM24
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3491.840 2435.000 3492.440 ;
    END
  END Tile_X11Y2_BEN_SRAM24
  PIN Tile_X11Y2_BEN_SRAM25
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3576.840 2435.000 3577.440 ;
    END
  END Tile_X11Y2_BEN_SRAM25
  PIN Tile_X11Y2_BEN_SRAM26
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3437.440 2435.000 3438.040 ;
    END
  END Tile_X11Y2_BEN_SRAM26
  PIN Tile_X11Y2_BEN_SRAM27
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3573.440 2435.000 3574.040 ;
    END
  END Tile_X11Y2_BEN_SRAM27
  PIN Tile_X11Y2_BEN_SRAM28
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3712.840 2435.000 3713.440 ;
    END
  END Tile_X11Y2_BEN_SRAM28
  PIN Tile_X11Y2_BEN_SRAM29
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3478.240 2435.000 3478.840 ;
    END
  END Tile_X11Y2_BEN_SRAM29
  PIN Tile_X11Y2_BEN_SRAM3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3638.040 2435.000 3638.640 ;
    END
  END Tile_X11Y2_BEN_SRAM3
  PIN Tile_X11Y2_BEN_SRAM30
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3760.440 2435.000 3761.040 ;
    END
  END Tile_X11Y2_BEN_SRAM30
  PIN Tile_X11Y2_BEN_SRAM31
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3444.240 2435.000 3444.840 ;
    END
  END Tile_X11Y2_BEN_SRAM31
  PIN Tile_X11Y2_BEN_SRAM4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3410.240 2435.000 3410.840 ;
    END
  END Tile_X11Y2_BEN_SRAM4
  PIN Tile_X11Y2_BEN_SRAM5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3641.440 2435.000 3642.040 ;
    END
  END Tile_X11Y2_BEN_SRAM5
  PIN Tile_X11Y2_BEN_SRAM6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3417.040 2435.000 3417.640 ;
    END
  END Tile_X11Y2_BEN_SRAM6
  PIN Tile_X11Y2_BEN_SRAM7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3716.240 2435.000 3716.840 ;
    END
  END Tile_X11Y2_BEN_SRAM7
  PIN Tile_X11Y2_BEN_SRAM8
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3644.840 2435.000 3645.440 ;
    END
  END Tile_X11Y2_BEN_SRAM8
  PIN Tile_X11Y2_BEN_SRAM9
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3525.840 2435.000 3526.440 ;
    END
  END Tile_X11Y2_BEN_SRAM9
  PIN Tile_X11Y2_CLOCK_SRAM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3661.840 2435.000 3662.440 ;
    END
  END Tile_X11Y2_CLOCK_SRAM
  PIN Tile_X11Y2_DI_SRAM0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3559.840 2435.000 3560.440 ;
    END
  END Tile_X11Y2_DI_SRAM0
  PIN Tile_X11Y2_DI_SRAM1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3447.640 2435.000 3448.240 ;
    END
  END Tile_X11Y2_DI_SRAM1
  PIN Tile_X11Y2_DI_SRAM10
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3556.440 2435.000 3557.040 ;
    END
  END Tile_X11Y2_DI_SRAM10
  PIN Tile_X11Y2_DI_SRAM11
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3505.440 2435.000 3506.040 ;
    END
  END Tile_X11Y2_DI_SRAM11
  PIN Tile_X11Y2_DI_SRAM12
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3750.240 2435.000 3750.840 ;
    END
  END Tile_X11Y2_DI_SRAM12
  PIN Tile_X11Y2_DI_SRAM13
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3719.640 2435.000 3720.240 ;
    END
  END Tile_X11Y2_DI_SRAM13
  PIN Tile_X11Y2_DI_SRAM14
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3631.240 2435.000 3631.840 ;
    END
  END Tile_X11Y2_DI_SRAM14
  PIN Tile_X11Y2_DI_SRAM15
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3549.640 2435.000 3550.240 ;
    END
  END Tile_X11Y2_DI_SRAM15
  PIN Tile_X11Y2_DI_SRAM16
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3468.040 2435.000 3468.640 ;
    END
  END Tile_X11Y2_DI_SRAM16
  PIN Tile_X11Y2_DI_SRAM17
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3542.840 2435.000 3543.440 ;
    END
  END Tile_X11Y2_DI_SRAM17
  PIN Tile_X11Y2_DI_SRAM18
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3723.040 2435.000 3723.640 ;
    END
  END Tile_X11Y2_DI_SRAM18
  PIN Tile_X11Y2_DI_SRAM19
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3522.440 2435.000 3523.040 ;
    END
  END Tile_X11Y2_DI_SRAM19
  PIN Tile_X11Y2_DI_SRAM2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3617.640 2435.000 3618.240 ;
    END
  END Tile_X11Y2_DI_SRAM2
  PIN Tile_X11Y2_DI_SRAM20
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3651.640 2435.000 3652.240 ;
    END
  END Tile_X11Y2_DI_SRAM20
  PIN Tile_X11Y2_DI_SRAM21
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3546.240 2435.000 3546.840 ;
    END
  END Tile_X11Y2_DI_SRAM21
  PIN Tile_X11Y2_DI_SRAM22
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3515.640 2435.000 3516.240 ;
    END
  END Tile_X11Y2_DI_SRAM22
  PIN Tile_X11Y2_DI_SRAM23
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3655.040 2435.000 3655.640 ;
    END
  END Tile_X11Y2_DI_SRAM23
  PIN Tile_X11Y2_DI_SRAM24
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3566.640 2435.000 3567.240 ;
    END
  END Tile_X11Y2_DI_SRAM24
  PIN Tile_X11Y2_DI_SRAM25
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3726.440 2435.000 3727.040 ;
    END
  END Tile_X11Y2_DI_SRAM25
  PIN Tile_X11Y2_DI_SRAM26
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3495.240 2435.000 3495.840 ;
    END
  END Tile_X11Y2_DI_SRAM26
  PIN Tile_X11Y2_DI_SRAM27
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3539.440 2435.000 3540.040 ;
    END
  END Tile_X11Y2_DI_SRAM27
  PIN Tile_X11Y2_DI_SRAM28
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3597.240 2435.000 3597.840 ;
    END
  END Tile_X11Y2_DI_SRAM28
  PIN Tile_X11Y2_DI_SRAM29
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3614.240 2435.000 3614.840 ;
    END
  END Tile_X11Y2_DI_SRAM29
  PIN Tile_X11Y2_DI_SRAM3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3553.040 2435.000 3553.640 ;
    END
  END Tile_X11Y2_DI_SRAM3
  PIN Tile_X11Y2_DI_SRAM30
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3627.840 2435.000 3628.440 ;
    END
  END Tile_X11Y2_DI_SRAM30
  PIN Tile_X11Y2_DI_SRAM31
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3488.440 2435.000 3489.040 ;
    END
  END Tile_X11Y2_DI_SRAM31
  PIN Tile_X11Y2_DI_SRAM4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3729.840 2435.000 3730.440 ;
    END
  END Tile_X11Y2_DI_SRAM4
  PIN Tile_X11Y2_DI_SRAM5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3658.440 2435.000 3659.040 ;
    END
  END Tile_X11Y2_DI_SRAM5
  PIN Tile_X11Y2_DI_SRAM6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3665.240 2435.000 3665.840 ;
    END
  END Tile_X11Y2_DI_SRAM6
  PIN Tile_X11Y2_DI_SRAM7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3461.240 2435.000 3461.840 ;
    END
  END Tile_X11Y2_DI_SRAM7
  PIN Tile_X11Y2_DI_SRAM8
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3753.640 2435.000 3754.240 ;
    END
  END Tile_X11Y2_DI_SRAM8
  PIN Tile_X11Y2_DI_SRAM9
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3481.640 2435.000 3482.240 ;
    END
  END Tile_X11Y2_DI_SRAM9
  PIN Tile_X11Y2_DO_SRAM0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3508.840 2435.000 3509.440 ;
    END
  END Tile_X11Y2_DO_SRAM0
  PIN Tile_X11Y2_DO_SRAM1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3682.240 2435.000 3682.840 ;
    END
  END Tile_X11Y2_DO_SRAM1
  PIN Tile_X11Y2_DO_SRAM10
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3451.040 2435.000 3451.640 ;
    END
  END Tile_X11Y2_DO_SRAM10
  PIN Tile_X11Y2_DO_SRAM11
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3733.240 2435.000 3733.840 ;
    END
  END Tile_X11Y2_DO_SRAM11
  PIN Tile_X11Y2_DO_SRAM12
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3668.640 2435.000 3669.240 ;
    END
  END Tile_X11Y2_DO_SRAM12
  PIN Tile_X11Y2_DO_SRAM13
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3406.840 2435.000 3407.440 ;
    END
  END Tile_X11Y2_DO_SRAM13
  PIN Tile_X11Y2_DO_SRAM14
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3440.840 2435.000 3441.440 ;
    END
  END Tile_X11Y2_DO_SRAM14
  PIN Tile_X11Y2_DO_SRAM15
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3593.840 2435.000 3594.440 ;
    END
  END Tile_X11Y2_DO_SRAM15
  PIN Tile_X11Y2_DO_SRAM16
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3672.040 2435.000 3672.640 ;
    END
  END Tile_X11Y2_DO_SRAM16
  PIN Tile_X11Y2_DO_SRAM17
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3600.640 2435.000 3601.240 ;
    END
  END Tile_X11Y2_DO_SRAM17
  PIN Tile_X11Y2_DO_SRAM18
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3736.640 2435.000 3737.240 ;
    END
  END Tile_X11Y2_DO_SRAM18
  PIN Tile_X11Y2_DO_SRAM19
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3570.040 2435.000 3570.640 ;
    END
  END Tile_X11Y2_DO_SRAM19
  PIN Tile_X11Y2_DO_SRAM2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3675.440 2435.000 3676.040 ;
    END
  END Tile_X11Y2_DO_SRAM2
  PIN Tile_X11Y2_DO_SRAM20
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3400.040 2435.000 3400.640 ;
    END
  END Tile_X11Y2_DO_SRAM20
  PIN Tile_X11Y2_DO_SRAM21
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3413.640 2435.000 3414.240 ;
    END
  END Tile_X11Y2_DO_SRAM21
  PIN Tile_X11Y2_DO_SRAM22
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3420.440 2435.000 3421.040 ;
    END
  END Tile_X11Y2_DO_SRAM22
  PIN Tile_X11Y2_DO_SRAM23
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3678.840 2435.000 3679.440 ;
    END
  END Tile_X11Y2_DO_SRAM23
  PIN Tile_X11Y2_DO_SRAM24
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3498.640 2435.000 3499.240 ;
    END
  END Tile_X11Y2_DO_SRAM24
  PIN Tile_X11Y2_DO_SRAM25
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3519.040 2435.000 3519.640 ;
    END
  END Tile_X11Y2_DO_SRAM25
  PIN Tile_X11Y2_DO_SRAM26
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3423.840 2435.000 3424.440 ;
    END
  END Tile_X11Y2_DO_SRAM26
  PIN Tile_X11Y2_DO_SRAM27
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3740.040 2435.000 3740.640 ;
    END
  END Tile_X11Y2_DO_SRAM27
  PIN Tile_X11Y2_DO_SRAM28
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3485.040 2435.000 3485.640 ;
    END
  END Tile_X11Y2_DO_SRAM28
  PIN Tile_X11Y2_DO_SRAM29
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3434.040 2435.000 3434.640 ;
    END
  END Tile_X11Y2_DO_SRAM29
  PIN Tile_X11Y2_DO_SRAM3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3685.640 2435.000 3686.240 ;
    END
  END Tile_X11Y2_DO_SRAM3
  PIN Tile_X11Y2_DO_SRAM30
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3763.840 2435.000 3764.440 ;
    END
  END Tile_X11Y2_DO_SRAM30
  PIN Tile_X11Y2_DO_SRAM31
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3563.240 2435.000 3563.840 ;
    END
  END Tile_X11Y2_DO_SRAM31
  PIN Tile_X11Y2_DO_SRAM4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3689.040 2435.000 3689.640 ;
    END
  END Tile_X11Y2_DO_SRAM4
  PIN Tile_X11Y2_DO_SRAM5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3471.440 2435.000 3472.040 ;
    END
  END Tile_X11Y2_DO_SRAM5
  PIN Tile_X11Y2_DO_SRAM6
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3583.640 2435.000 3584.240 ;
    END
  END Tile_X11Y2_DO_SRAM6
  PIN Tile_X11Y2_DO_SRAM7
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3607.440 2435.000 3608.040 ;
    END
  END Tile_X11Y2_DO_SRAM7
  PIN Tile_X11Y2_DO_SRAM8
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3532.640 2435.000 3533.240 ;
    END
  END Tile_X11Y2_DO_SRAM8
  PIN Tile_X11Y2_DO_SRAM9
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3692.440 2435.000 3693.040 ;
    END
  END Tile_X11Y2_DO_SRAM9
  PIN Tile_X11Y2_EN_SRAM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3529.240 2435.000 3529.840 ;
    END
  END Tile_X11Y2_EN_SRAM
  PIN Tile_X11Y2_R_WB_SRAM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3604.040 2435.000 3604.640 ;
    END
  END Tile_X11Y2_R_WB_SRAM
  PIN Tile_X11Y4_AD_SRAM0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2784.640 2435.000 2785.240 ;
    END
  END Tile_X11Y4_AD_SRAM0
  PIN Tile_X11Y4_AD_SRAM1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2937.640 2435.000 2938.240 ;
    END
  END Tile_X11Y4_AD_SRAM1
  PIN Tile_X11Y4_AD_SRAM2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2825.440 2435.000 2826.040 ;
    END
  END Tile_X11Y4_AD_SRAM2
  PIN Tile_X11Y4_AD_SRAM3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2941.040 2435.000 2941.640 ;
    END
  END Tile_X11Y4_AD_SRAM3
  PIN Tile_X11Y4_AD_SRAM4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2822.040 2435.000 2822.640 ;
    END
  END Tile_X11Y4_AD_SRAM4
  PIN Tile_X11Y4_AD_SRAM5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2818.640 2435.000 2819.240 ;
    END
  END Tile_X11Y4_AD_SRAM5
  PIN Tile_X11Y4_AD_SRAM6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2944.440 2435.000 2945.040 ;
    END
  END Tile_X11Y4_AD_SRAM6
  PIN Tile_X11Y4_AD_SRAM7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2815.240 2435.000 2815.840 ;
    END
  END Tile_X11Y4_AD_SRAM7
  PIN Tile_X11Y4_AD_SRAM8
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2947.840 2435.000 2948.440 ;
    END
  END Tile_X11Y4_AD_SRAM8
  PIN Tile_X11Y4_AD_SRAM9
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2811.840 2435.000 2812.440 ;
    END
  END Tile_X11Y4_AD_SRAM9
  PIN Tile_X11Y4_BEN_SRAM0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2808.440 2435.000 2809.040 ;
    END
  END Tile_X11Y4_BEN_SRAM0
  PIN Tile_X11Y4_BEN_SRAM1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2951.240 2435.000 2951.840 ;
    END
  END Tile_X11Y4_BEN_SRAM1
  PIN Tile_X11Y4_BEN_SRAM10
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2788.040 2435.000 2788.640 ;
    END
  END Tile_X11Y4_BEN_SRAM10
  PIN Tile_X11Y4_BEN_SRAM11
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2964.840 2435.000 2965.440 ;
    END
  END Tile_X11Y4_BEN_SRAM11
  PIN Tile_X11Y4_BEN_SRAM12
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2968.240 2435.000 2968.840 ;
    END
  END Tile_X11Y4_BEN_SRAM12
  PIN Tile_X11Y4_BEN_SRAM13
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3151.840 2435.000 3152.440 ;
    END
  END Tile_X11Y4_BEN_SRAM13
  PIN Tile_X11Y4_BEN_SRAM14
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3148.440 2435.000 3149.040 ;
    END
  END Tile_X11Y4_BEN_SRAM14
  PIN Tile_X11Y4_BEN_SRAM15
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2971.640 2435.000 2972.240 ;
    END
  END Tile_X11Y4_BEN_SRAM15
  PIN Tile_X11Y4_BEN_SRAM16
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3145.040 2435.000 3145.640 ;
    END
  END Tile_X11Y4_BEN_SRAM16
  PIN Tile_X11Y4_BEN_SRAM17
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2975.040 2435.000 2975.640 ;
    END
  END Tile_X11Y4_BEN_SRAM17
  PIN Tile_X11Y4_BEN_SRAM18
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3141.640 2435.000 3142.240 ;
    END
  END Tile_X11Y4_BEN_SRAM18
  PIN Tile_X11Y4_BEN_SRAM19
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3138.240 2435.000 3138.840 ;
    END
  END Tile_X11Y4_BEN_SRAM19
  PIN Tile_X11Y4_BEN_SRAM2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2805.040 2435.000 2805.640 ;
    END
  END Tile_X11Y4_BEN_SRAM2
  PIN Tile_X11Y4_BEN_SRAM20
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2978.440 2435.000 2979.040 ;
    END
  END Tile_X11Y4_BEN_SRAM20
  PIN Tile_X11Y4_BEN_SRAM21
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3134.840 2435.000 3135.440 ;
    END
  END Tile_X11Y4_BEN_SRAM21
  PIN Tile_X11Y4_BEN_SRAM22
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2981.840 2435.000 2982.440 ;
    END
  END Tile_X11Y4_BEN_SRAM22
  PIN Tile_X11Y4_BEN_SRAM23
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3131.440 2435.000 3132.040 ;
    END
  END Tile_X11Y4_BEN_SRAM23
  PIN Tile_X11Y4_BEN_SRAM24
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3128.040 2435.000 3128.640 ;
    END
  END Tile_X11Y4_BEN_SRAM24
  PIN Tile_X11Y4_BEN_SRAM25
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2985.240 2435.000 2985.840 ;
    END
  END Tile_X11Y4_BEN_SRAM25
  PIN Tile_X11Y4_BEN_SRAM26
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3124.640 2435.000 3125.240 ;
    END
  END Tile_X11Y4_BEN_SRAM26
  PIN Tile_X11Y4_BEN_SRAM27
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2988.640 2435.000 2989.240 ;
    END
  END Tile_X11Y4_BEN_SRAM27
  PIN Tile_X11Y4_BEN_SRAM28
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3121.240 2435.000 3121.840 ;
    END
  END Tile_X11Y4_BEN_SRAM28
  PIN Tile_X11Y4_BEN_SRAM29
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3117.840 2435.000 3118.440 ;
    END
  END Tile_X11Y4_BEN_SRAM29
  PIN Tile_X11Y4_BEN_SRAM3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2954.640 2435.000 2955.240 ;
    END
  END Tile_X11Y4_BEN_SRAM3
  PIN Tile_X11Y4_BEN_SRAM30
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2992.040 2435.000 2992.640 ;
    END
  END Tile_X11Y4_BEN_SRAM30
  PIN Tile_X11Y4_BEN_SRAM31
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3114.440 2435.000 3115.040 ;
    END
  END Tile_X11Y4_BEN_SRAM31
  PIN Tile_X11Y4_BEN_SRAM4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2801.640 2435.000 2802.240 ;
    END
  END Tile_X11Y4_BEN_SRAM4
  PIN Tile_X11Y4_BEN_SRAM5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2798.240 2435.000 2798.840 ;
    END
  END Tile_X11Y4_BEN_SRAM5
  PIN Tile_X11Y4_BEN_SRAM6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2958.040 2435.000 2958.640 ;
    END
  END Tile_X11Y4_BEN_SRAM6
  PIN Tile_X11Y4_BEN_SRAM7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2794.840 2435.000 2795.440 ;
    END
  END Tile_X11Y4_BEN_SRAM7
  PIN Tile_X11Y4_BEN_SRAM8
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2961.440 2435.000 2962.040 ;
    END
  END Tile_X11Y4_BEN_SRAM8
  PIN Tile_X11Y4_BEN_SRAM9
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2791.440 2435.000 2792.040 ;
    END
  END Tile_X11Y4_BEN_SRAM9
  PIN Tile_X11Y4_CLOCK_SRAM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2995.440 2435.000 2996.040 ;
    END
  END Tile_X11Y4_CLOCK_SRAM
  PIN Tile_X11Y4_DI_SRAM0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3111.040 2435.000 3111.640 ;
    END
  END Tile_X11Y4_DI_SRAM0
  PIN Tile_X11Y4_DI_SRAM1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3107.640 2435.000 3108.240 ;
    END
  END Tile_X11Y4_DI_SRAM1
  PIN Tile_X11Y4_DI_SRAM10
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3104.240 2435.000 3104.840 ;
    END
  END Tile_X11Y4_DI_SRAM10
  PIN Tile_X11Y4_DI_SRAM11
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3087.240 2435.000 3087.840 ;
    END
  END Tile_X11Y4_DI_SRAM11
  PIN Tile_X11Y4_DI_SRAM12
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3060.040 2435.000 3060.640 ;
    END
  END Tile_X11Y4_DI_SRAM12
  PIN Tile_X11Y4_DI_SRAM13
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3083.840 2435.000 3084.440 ;
    END
  END Tile_X11Y4_DI_SRAM13
  PIN Tile_X11Y4_DI_SRAM14
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3022.640 2435.000 3023.240 ;
    END
  END Tile_X11Y4_DI_SRAM14
  PIN Tile_X11Y4_DI_SRAM15
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3097.440 2435.000 3098.040 ;
    END
  END Tile_X11Y4_DI_SRAM15
  PIN Tile_X11Y4_DI_SRAM16
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3077.040 2435.000 3077.640 ;
    END
  END Tile_X11Y4_DI_SRAM16
  PIN Tile_X11Y4_DI_SRAM17
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3019.240 2435.000 3019.840 ;
    END
  END Tile_X11Y4_DI_SRAM17
  PIN Tile_X11Y4_DI_SRAM18
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3073.640 2435.000 3074.240 ;
    END
  END Tile_X11Y4_DI_SRAM18
  PIN Tile_X11Y4_DI_SRAM19
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3039.640 2435.000 3040.240 ;
    END
  END Tile_X11Y4_DI_SRAM19
  PIN Tile_X11Y4_DI_SRAM2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2998.840 2435.000 2999.440 ;
    END
  END Tile_X11Y4_DI_SRAM2
  PIN Tile_X11Y4_DI_SRAM20
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3070.240 2435.000 3070.840 ;
    END
  END Tile_X11Y4_DI_SRAM20
  PIN Tile_X11Y4_DI_SRAM21
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3066.840 2435.000 3067.440 ;
    END
  END Tile_X11Y4_DI_SRAM21
  PIN Tile_X11Y4_DI_SRAM22
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3026.040 2435.000 3026.640 ;
    END
  END Tile_X11Y4_DI_SRAM22
  PIN Tile_X11Y4_DI_SRAM23
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3094.040 2435.000 3094.640 ;
    END
  END Tile_X11Y4_DI_SRAM23
  PIN Tile_X11Y4_DI_SRAM24
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3036.240 2435.000 3036.840 ;
    END
  END Tile_X11Y4_DI_SRAM24
  PIN Tile_X11Y4_DI_SRAM25
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3090.640 2435.000 3091.240 ;
    END
  END Tile_X11Y4_DI_SRAM25
  PIN Tile_X11Y4_DI_SRAM26
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3056.640 2435.000 3057.240 ;
    END
  END Tile_X11Y4_DI_SRAM26
  PIN Tile_X11Y4_DI_SRAM27
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3032.840 2435.000 3033.440 ;
    END
  END Tile_X11Y4_DI_SRAM27
  PIN Tile_X11Y4_DI_SRAM28
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3053.240 2435.000 3053.840 ;
    END
  END Tile_X11Y4_DI_SRAM28
  PIN Tile_X11Y4_DI_SRAM29
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3100.840 2435.000 3101.440 ;
    END
  END Tile_X11Y4_DI_SRAM29
  PIN Tile_X11Y4_DI_SRAM3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3002.240 2435.000 3002.840 ;
    END
  END Tile_X11Y4_DI_SRAM3
  PIN Tile_X11Y4_DI_SRAM30
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3049.840 2435.000 3050.440 ;
    END
  END Tile_X11Y4_DI_SRAM30
  PIN Tile_X11Y4_DI_SRAM31
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3046.440 2435.000 3047.040 ;
    END
  END Tile_X11Y4_DI_SRAM31
  PIN Tile_X11Y4_DI_SRAM4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3043.040 2435.000 3043.640 ;
    END
  END Tile_X11Y4_DI_SRAM4
  PIN Tile_X11Y4_DI_SRAM5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3005.640 2435.000 3006.240 ;
    END
  END Tile_X11Y4_DI_SRAM5
  PIN Tile_X11Y4_DI_SRAM6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3009.040 2435.000 3009.640 ;
    END
  END Tile_X11Y4_DI_SRAM6
  PIN Tile_X11Y4_DI_SRAM7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3012.440 2435.000 3013.040 ;
    END
  END Tile_X11Y4_DI_SRAM7
  PIN Tile_X11Y4_DI_SRAM8
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3015.840 2435.000 3016.440 ;
    END
  END Tile_X11Y4_DI_SRAM8
  PIN Tile_X11Y4_DI_SRAM9
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3029.440 2435.000 3030.040 ;
    END
  END Tile_X11Y4_DI_SRAM9
  PIN Tile_X11Y4_DO_SRAM0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2828.840 2435.000 2829.440 ;
    END
  END Tile_X11Y4_DO_SRAM0
  PIN Tile_X11Y4_DO_SRAM1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2893.440 2435.000 2894.040 ;
    END
  END Tile_X11Y4_DO_SRAM1
  PIN Tile_X11Y4_DO_SRAM10
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2907.040 2435.000 2907.640 ;
    END
  END Tile_X11Y4_DO_SRAM10
  PIN Tile_X11Y4_DO_SRAM11
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2873.040 2435.000 2873.640 ;
    END
  END Tile_X11Y4_DO_SRAM11
  PIN Tile_X11Y4_DO_SRAM12
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2869.640 2435.000 2870.240 ;
    END
  END Tile_X11Y4_DO_SRAM12
  PIN Tile_X11Y4_DO_SRAM13
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2910.440 2435.000 2911.040 ;
    END
  END Tile_X11Y4_DO_SRAM13
  PIN Tile_X11Y4_DO_SRAM14
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2866.240 2435.000 2866.840 ;
    END
  END Tile_X11Y4_DO_SRAM14
  PIN Tile_X11Y4_DO_SRAM15
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2913.840 2435.000 2914.440 ;
    END
  END Tile_X11Y4_DO_SRAM15
  PIN Tile_X11Y4_DO_SRAM16
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2862.840 2435.000 2863.440 ;
    END
  END Tile_X11Y4_DO_SRAM16
  PIN Tile_X11Y4_DO_SRAM17
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2859.440 2435.000 2860.040 ;
    END
  END Tile_X11Y4_DO_SRAM17
  PIN Tile_X11Y4_DO_SRAM18
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2917.240 2435.000 2917.840 ;
    END
  END Tile_X11Y4_DO_SRAM18
  PIN Tile_X11Y4_DO_SRAM19
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2856.040 2435.000 2856.640 ;
    END
  END Tile_X11Y4_DO_SRAM19
  PIN Tile_X11Y4_DO_SRAM2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2890.040 2435.000 2890.640 ;
    END
  END Tile_X11Y4_DO_SRAM2
  PIN Tile_X11Y4_DO_SRAM20
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2920.640 2435.000 2921.240 ;
    END
  END Tile_X11Y4_DO_SRAM20
  PIN Tile_X11Y4_DO_SRAM21
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2852.640 2435.000 2853.240 ;
    END
  END Tile_X11Y4_DO_SRAM21
  PIN Tile_X11Y4_DO_SRAM22
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2849.240 2435.000 2849.840 ;
    END
  END Tile_X11Y4_DO_SRAM22
  PIN Tile_X11Y4_DO_SRAM23
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2924.040 2435.000 2924.640 ;
    END
  END Tile_X11Y4_DO_SRAM23
  PIN Tile_X11Y4_DO_SRAM24
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2845.840 2435.000 2846.440 ;
    END
  END Tile_X11Y4_DO_SRAM24
  PIN Tile_X11Y4_DO_SRAM25
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2927.440 2435.000 2928.040 ;
    END
  END Tile_X11Y4_DO_SRAM25
  PIN Tile_X11Y4_DO_SRAM26
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2842.440 2435.000 2843.040 ;
    END
  END Tile_X11Y4_DO_SRAM26
  PIN Tile_X11Y4_DO_SRAM27
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2839.040 2435.000 2839.640 ;
    END
  END Tile_X11Y4_DO_SRAM27
  PIN Tile_X11Y4_DO_SRAM28
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2930.840 2435.000 2931.440 ;
    END
  END Tile_X11Y4_DO_SRAM28
  PIN Tile_X11Y4_DO_SRAM29
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2835.640 2435.000 2836.240 ;
    END
  END Tile_X11Y4_DO_SRAM29
  PIN Tile_X11Y4_DO_SRAM3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2896.840 2435.000 2897.440 ;
    END
  END Tile_X11Y4_DO_SRAM3
  PIN Tile_X11Y4_DO_SRAM30
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2934.240 2435.000 2934.840 ;
    END
  END Tile_X11Y4_DO_SRAM30
  PIN Tile_X11Y4_DO_SRAM31
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2832.240 2435.000 2832.840 ;
    END
  END Tile_X11Y4_DO_SRAM31
  PIN Tile_X11Y4_DO_SRAM4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2886.640 2435.000 2887.240 ;
    END
  END Tile_X11Y4_DO_SRAM4
  PIN Tile_X11Y4_DO_SRAM5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2900.240 2435.000 2900.840 ;
    END
  END Tile_X11Y4_DO_SRAM5
  PIN Tile_X11Y4_DO_SRAM6
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2883.240 2435.000 2883.840 ;
    END
  END Tile_X11Y4_DO_SRAM6
  PIN Tile_X11Y4_DO_SRAM7
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2879.840 2435.000 2880.440 ;
    END
  END Tile_X11Y4_DO_SRAM7
  PIN Tile_X11Y4_DO_SRAM8
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2903.640 2435.000 2904.240 ;
    END
  END Tile_X11Y4_DO_SRAM8
  PIN Tile_X11Y4_DO_SRAM9
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2876.440 2435.000 2877.040 ;
    END
  END Tile_X11Y4_DO_SRAM9
  PIN Tile_X11Y4_EN_SRAM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3080.440 2435.000 3081.040 ;
    END
  END Tile_X11Y4_EN_SRAM
  PIN Tile_X11Y4_R_WB_SRAM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 3063.440 2435.000 3064.040 ;
    END
  END Tile_X11Y4_R_WB_SRAM
  PIN Tile_X11Y6_AD_SRAM0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2332.440 2435.000 2333.040 ;
    END
  END Tile_X11Y6_AD_SRAM0
  PIN Tile_X11Y6_AD_SRAM1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2376.640 2435.000 2377.240 ;
    END
  END Tile_X11Y6_AD_SRAM1
  PIN Tile_X11Y6_AD_SRAM2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2488.840 2435.000 2489.440 ;
    END
  END Tile_X11Y6_AD_SRAM2
  PIN Tile_X11Y6_AD_SRAM3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2373.240 2435.000 2373.840 ;
    END
  END Tile_X11Y6_AD_SRAM3
  PIN Tile_X11Y6_AD_SRAM4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2492.240 2435.000 2492.840 ;
    END
  END Tile_X11Y6_AD_SRAM4
  PIN Tile_X11Y6_AD_SRAM5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2369.840 2435.000 2370.440 ;
    END
  END Tile_X11Y6_AD_SRAM5
  PIN Tile_X11Y6_AD_SRAM6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2366.440 2435.000 2367.040 ;
    END
  END Tile_X11Y6_AD_SRAM6
  PIN Tile_X11Y6_AD_SRAM7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2495.640 2435.000 2496.240 ;
    END
  END Tile_X11Y6_AD_SRAM7
  PIN Tile_X11Y6_AD_SRAM8
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2363.040 2435.000 2363.640 ;
    END
  END Tile_X11Y6_AD_SRAM8
  PIN Tile_X11Y6_AD_SRAM9
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2499.040 2435.000 2499.640 ;
    END
  END Tile_X11Y6_AD_SRAM9
  PIN Tile_X11Y6_BEN_SRAM0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2359.640 2435.000 2360.240 ;
    END
  END Tile_X11Y6_BEN_SRAM0
  PIN Tile_X11Y6_BEN_SRAM1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2356.240 2435.000 2356.840 ;
    END
  END Tile_X11Y6_BEN_SRAM1
  PIN Tile_X11Y6_BEN_SRAM10
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2339.240 2435.000 2339.840 ;
    END
  END Tile_X11Y6_BEN_SRAM10
  PIN Tile_X11Y6_BEN_SRAM11
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2335.840 2435.000 2336.440 ;
    END
  END Tile_X11Y6_BEN_SRAM11
  PIN Tile_X11Y6_BEN_SRAM12
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2516.040 2435.000 2516.640 ;
    END
  END Tile_X11Y6_BEN_SRAM12
  PIN Tile_X11Y6_BEN_SRAM13
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2519.440 2435.000 2520.040 ;
    END
  END Tile_X11Y6_BEN_SRAM13
  PIN Tile_X11Y6_BEN_SRAM14
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2699.640 2435.000 2700.240 ;
    END
  END Tile_X11Y6_BEN_SRAM14
  PIN Tile_X11Y6_BEN_SRAM15
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2696.240 2435.000 2696.840 ;
    END
  END Tile_X11Y6_BEN_SRAM15
  PIN Tile_X11Y6_BEN_SRAM16
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2522.840 2435.000 2523.440 ;
    END
  END Tile_X11Y6_BEN_SRAM16
  PIN Tile_X11Y6_BEN_SRAM17
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2692.840 2435.000 2693.440 ;
    END
  END Tile_X11Y6_BEN_SRAM17
  PIN Tile_X11Y6_BEN_SRAM18
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2526.240 2435.000 2526.840 ;
    END
  END Tile_X11Y6_BEN_SRAM18
  PIN Tile_X11Y6_BEN_SRAM19
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2689.440 2435.000 2690.040 ;
    END
  END Tile_X11Y6_BEN_SRAM19
  PIN Tile_X11Y6_BEN_SRAM2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2502.440 2435.000 2503.040 ;
    END
  END Tile_X11Y6_BEN_SRAM2
  PIN Tile_X11Y6_BEN_SRAM20
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2686.040 2435.000 2686.640 ;
    END
  END Tile_X11Y6_BEN_SRAM20
  PIN Tile_X11Y6_BEN_SRAM21
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2529.640 2435.000 2530.240 ;
    END
  END Tile_X11Y6_BEN_SRAM21
  PIN Tile_X11Y6_BEN_SRAM22
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2682.640 2435.000 2683.240 ;
    END
  END Tile_X11Y6_BEN_SRAM22
  PIN Tile_X11Y6_BEN_SRAM23
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2533.040 2435.000 2533.640 ;
    END
  END Tile_X11Y6_BEN_SRAM23
  PIN Tile_X11Y6_BEN_SRAM24
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2679.240 2435.000 2679.840 ;
    END
  END Tile_X11Y6_BEN_SRAM24
  PIN Tile_X11Y6_BEN_SRAM25
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2675.840 2435.000 2676.440 ;
    END
  END Tile_X11Y6_BEN_SRAM25
  PIN Tile_X11Y6_BEN_SRAM26
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2536.440 2435.000 2537.040 ;
    END
  END Tile_X11Y6_BEN_SRAM26
  PIN Tile_X11Y6_BEN_SRAM27
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2672.440 2435.000 2673.040 ;
    END
  END Tile_X11Y6_BEN_SRAM27
  PIN Tile_X11Y6_BEN_SRAM28
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2539.840 2435.000 2540.440 ;
    END
  END Tile_X11Y6_BEN_SRAM28
  PIN Tile_X11Y6_BEN_SRAM29
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2669.040 2435.000 2669.640 ;
    END
  END Tile_X11Y6_BEN_SRAM29
  PIN Tile_X11Y6_BEN_SRAM3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2352.840 2435.000 2353.440 ;
    END
  END Tile_X11Y6_BEN_SRAM3
  PIN Tile_X11Y6_BEN_SRAM30
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2665.640 2435.000 2666.240 ;
    END
  END Tile_X11Y6_BEN_SRAM30
  PIN Tile_X11Y6_BEN_SRAM31
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2543.240 2435.000 2543.840 ;
    END
  END Tile_X11Y6_BEN_SRAM31
  PIN Tile_X11Y6_BEN_SRAM4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2505.840 2435.000 2506.440 ;
    END
  END Tile_X11Y6_BEN_SRAM4
  PIN Tile_X11Y6_BEN_SRAM5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2349.440 2435.000 2350.040 ;
    END
  END Tile_X11Y6_BEN_SRAM5
  PIN Tile_X11Y6_BEN_SRAM6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2346.040 2435.000 2346.640 ;
    END
  END Tile_X11Y6_BEN_SRAM6
  PIN Tile_X11Y6_BEN_SRAM7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2509.240 2435.000 2509.840 ;
    END
  END Tile_X11Y6_BEN_SRAM7
  PIN Tile_X11Y6_BEN_SRAM8
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2342.640 2435.000 2343.240 ;
    END
  END Tile_X11Y6_BEN_SRAM8
  PIN Tile_X11Y6_BEN_SRAM9
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2512.640 2435.000 2513.240 ;
    END
  END Tile_X11Y6_BEN_SRAM9
  PIN Tile_X11Y6_CLOCK_SRAM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2662.240 2435.000 2662.840 ;
    END
  END Tile_X11Y6_CLOCK_SRAM
  PIN Tile_X11Y6_DI_SRAM0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2546.640 2435.000 2547.240 ;
    END
  END Tile_X11Y6_DI_SRAM0
  PIN Tile_X11Y6_DI_SRAM1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2658.840 2435.000 2659.440 ;
    END
  END Tile_X11Y6_DI_SRAM1
  PIN Tile_X11Y6_DI_SRAM10
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2655.440 2435.000 2656.040 ;
    END
  END Tile_X11Y6_DI_SRAM10
  PIN Tile_X11Y6_DI_SRAM11
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2638.440 2435.000 2639.040 ;
    END
  END Tile_X11Y6_DI_SRAM11
  PIN Tile_X11Y6_DI_SRAM12
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2635.040 2435.000 2635.640 ;
    END
  END Tile_X11Y6_DI_SRAM12
  PIN Tile_X11Y6_DI_SRAM13
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2570.440 2435.000 2571.040 ;
    END
  END Tile_X11Y6_DI_SRAM13
  PIN Tile_X11Y6_DI_SRAM14
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2631.640 2435.000 2632.240 ;
    END
  END Tile_X11Y6_DI_SRAM14
  PIN Tile_X11Y6_DI_SRAM15
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2590.840 2435.000 2591.440 ;
    END
  END Tile_X11Y6_DI_SRAM15
  PIN Tile_X11Y6_DI_SRAM16
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2645.240 2435.000 2645.840 ;
    END
  END Tile_X11Y6_DI_SRAM16
  PIN Tile_X11Y6_DI_SRAM17
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2624.840 2435.000 2625.440 ;
    END
  END Tile_X11Y6_DI_SRAM17
  PIN Tile_X11Y6_DI_SRAM18
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2577.240 2435.000 2577.840 ;
    END
  END Tile_X11Y6_DI_SRAM18
  PIN Tile_X11Y6_DI_SRAM19
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2621.440 2435.000 2622.040 ;
    END
  END Tile_X11Y6_DI_SRAM19
  PIN Tile_X11Y6_DI_SRAM2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2550.040 2435.000 2550.640 ;
    END
  END Tile_X11Y6_DI_SRAM2
  PIN Tile_X11Y6_DI_SRAM20
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2573.840 2435.000 2574.440 ;
    END
  END Tile_X11Y6_DI_SRAM20
  PIN Tile_X11Y6_DI_SRAM21
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2618.040 2435.000 2618.640 ;
    END
  END Tile_X11Y6_DI_SRAM21
  PIN Tile_X11Y6_DI_SRAM22
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2614.640 2435.000 2615.240 ;
    END
  END Tile_X11Y6_DI_SRAM22
  PIN Tile_X11Y6_DI_SRAM23
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2594.240 2435.000 2594.840 ;
    END
  END Tile_X11Y6_DI_SRAM23
  PIN Tile_X11Y6_DI_SRAM24
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2641.840 2435.000 2642.440 ;
    END
  END Tile_X11Y6_DI_SRAM24
  PIN Tile_X11Y6_DI_SRAM25
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2580.640 2435.000 2581.240 ;
    END
  END Tile_X11Y6_DI_SRAM25
  PIN Tile_X11Y6_DI_SRAM26
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2652.040 2435.000 2652.640 ;
    END
  END Tile_X11Y6_DI_SRAM26
  PIN Tile_X11Y6_DI_SRAM27
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2604.440 2435.000 2605.040 ;
    END
  END Tile_X11Y6_DI_SRAM27
  PIN Tile_X11Y6_DI_SRAM28
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2611.240 2435.000 2611.840 ;
    END
  END Tile_X11Y6_DI_SRAM28
  PIN Tile_X11Y6_DI_SRAM29
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2601.040 2435.000 2601.640 ;
    END
  END Tile_X11Y6_DI_SRAM29
  PIN Tile_X11Y6_DI_SRAM3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2556.840 2435.000 2557.440 ;
    END
  END Tile_X11Y6_DI_SRAM3
  PIN Tile_X11Y6_DI_SRAM30
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2587.440 2435.000 2588.040 ;
    END
  END Tile_X11Y6_DI_SRAM30
  PIN Tile_X11Y6_DI_SRAM31
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2597.640 2435.000 2598.240 ;
    END
  END Tile_X11Y6_DI_SRAM31
  PIN Tile_X11Y6_DI_SRAM4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2553.440 2435.000 2554.040 ;
    END
  END Tile_X11Y6_DI_SRAM4
  PIN Tile_X11Y6_DI_SRAM5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2563.640 2435.000 2564.240 ;
    END
  END Tile_X11Y6_DI_SRAM5
  PIN Tile_X11Y6_DI_SRAM6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2567.040 2435.000 2567.640 ;
    END
  END Tile_X11Y6_DI_SRAM6
  PIN Tile_X11Y6_DI_SRAM7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2560.240 2435.000 2560.840 ;
    END
  END Tile_X11Y6_DI_SRAM7
  PIN Tile_X11Y6_DI_SRAM8
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2607.840 2435.000 2608.440 ;
    END
  END Tile_X11Y6_DI_SRAM8
  PIN Tile_X11Y6_DI_SRAM9
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2584.040 2435.000 2584.640 ;
    END
  END Tile_X11Y6_DI_SRAM9
  PIN Tile_X11Y6_DO_SRAM0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2380.040 2435.000 2380.640 ;
    END
  END Tile_X11Y6_DO_SRAM0
  PIN Tile_X11Y6_DO_SRAM1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2444.640 2435.000 2445.240 ;
    END
  END Tile_X11Y6_DO_SRAM1
  PIN Tile_X11Y6_DO_SRAM10
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2424.240 2435.000 2424.840 ;
    END
  END Tile_X11Y6_DO_SRAM10
  PIN Tile_X11Y6_DO_SRAM11
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2458.240 2435.000 2458.840 ;
    END
  END Tile_X11Y6_DO_SRAM11
  PIN Tile_X11Y6_DO_SRAM12
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2420.840 2435.000 2421.440 ;
    END
  END Tile_X11Y6_DO_SRAM12
  PIN Tile_X11Y6_DO_SRAM13
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2417.440 2435.000 2418.040 ;
    END
  END Tile_X11Y6_DO_SRAM13
  PIN Tile_X11Y6_DO_SRAM14
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2461.640 2435.000 2462.240 ;
    END
  END Tile_X11Y6_DO_SRAM14
  PIN Tile_X11Y6_DO_SRAM15
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2414.040 2435.000 2414.640 ;
    END
  END Tile_X11Y6_DO_SRAM15
  PIN Tile_X11Y6_DO_SRAM16
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2465.040 2435.000 2465.640 ;
    END
  END Tile_X11Y6_DO_SRAM16
  PIN Tile_X11Y6_DO_SRAM17
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2410.640 2435.000 2411.240 ;
    END
  END Tile_X11Y6_DO_SRAM17
  PIN Tile_X11Y6_DO_SRAM18
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2407.240 2435.000 2407.840 ;
    END
  END Tile_X11Y6_DO_SRAM18
  PIN Tile_X11Y6_DO_SRAM19
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2468.440 2435.000 2469.040 ;
    END
  END Tile_X11Y6_DO_SRAM19
  PIN Tile_X11Y6_DO_SRAM2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2441.240 2435.000 2441.840 ;
    END
  END Tile_X11Y6_DO_SRAM2
  PIN Tile_X11Y6_DO_SRAM20
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2403.840 2435.000 2404.440 ;
    END
  END Tile_X11Y6_DO_SRAM20
  PIN Tile_X11Y6_DO_SRAM21
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2471.840 2435.000 2472.440 ;
    END
  END Tile_X11Y6_DO_SRAM21
  PIN Tile_X11Y6_DO_SRAM22
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2400.440 2435.000 2401.040 ;
    END
  END Tile_X11Y6_DO_SRAM22
  PIN Tile_X11Y6_DO_SRAM23
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2397.040 2435.000 2397.640 ;
    END
  END Tile_X11Y6_DO_SRAM23
  PIN Tile_X11Y6_DO_SRAM24
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2475.240 2435.000 2475.840 ;
    END
  END Tile_X11Y6_DO_SRAM24
  PIN Tile_X11Y6_DO_SRAM25
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2393.640 2435.000 2394.240 ;
    END
  END Tile_X11Y6_DO_SRAM25
  PIN Tile_X11Y6_DO_SRAM26
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2478.640 2435.000 2479.240 ;
    END
  END Tile_X11Y6_DO_SRAM26
  PIN Tile_X11Y6_DO_SRAM27
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2390.240 2435.000 2390.840 ;
    END
  END Tile_X11Y6_DO_SRAM27
  PIN Tile_X11Y6_DO_SRAM28
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2386.840 2435.000 2387.440 ;
    END
  END Tile_X11Y6_DO_SRAM28
  PIN Tile_X11Y6_DO_SRAM29
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2482.040 2435.000 2482.640 ;
    END
  END Tile_X11Y6_DO_SRAM29
  PIN Tile_X11Y6_DO_SRAM3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2437.840 2435.000 2438.440 ;
    END
  END Tile_X11Y6_DO_SRAM3
  PIN Tile_X11Y6_DO_SRAM30
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2383.440 2435.000 2384.040 ;
    END
  END Tile_X11Y6_DO_SRAM30
  PIN Tile_X11Y6_DO_SRAM31
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2485.440 2435.000 2486.040 ;
    END
  END Tile_X11Y6_DO_SRAM31
  PIN Tile_X11Y6_DO_SRAM4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2448.040 2435.000 2448.640 ;
    END
  END Tile_X11Y6_DO_SRAM4
  PIN Tile_X11Y6_DO_SRAM5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2434.440 2435.000 2435.040 ;
    END
  END Tile_X11Y6_DO_SRAM5
  PIN Tile_X11Y6_DO_SRAM6
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2451.440 2435.000 2452.040 ;
    END
  END Tile_X11Y6_DO_SRAM6
  PIN Tile_X11Y6_DO_SRAM7
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2431.040 2435.000 2431.640 ;
    END
  END Tile_X11Y6_DO_SRAM7
  PIN Tile_X11Y6_DO_SRAM8
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2427.640 2435.000 2428.240 ;
    END
  END Tile_X11Y6_DO_SRAM8
  PIN Tile_X11Y6_DO_SRAM9
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2454.840 2435.000 2455.440 ;
    END
  END Tile_X11Y6_DO_SRAM9
  PIN Tile_X11Y6_EN_SRAM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2628.240 2435.000 2628.840 ;
    END
  END Tile_X11Y6_EN_SRAM
  PIN Tile_X11Y6_R_WB_SRAM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2648.640 2435.000 2649.240 ;
    END
  END Tile_X11Y6_R_WB_SRAM
  PIN Tile_X11Y8_AD_SRAM0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2298.440 2435.000 2299.040 ;
    END
  END Tile_X11Y8_AD_SRAM0
  PIN Tile_X11Y8_AD_SRAM1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2043.440 2435.000 2044.040 ;
    END
  END Tile_X11Y8_AD_SRAM1
  PIN Tile_X11Y8_AD_SRAM2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2040.040 2435.000 2040.640 ;
    END
  END Tile_X11Y8_AD_SRAM2
  PIN Tile_X11Y8_AD_SRAM3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2291.640 2435.000 2292.240 ;
    END
  END Tile_X11Y8_AD_SRAM3
  PIN Tile_X11Y8_AD_SRAM4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2050.240 2435.000 2050.840 ;
    END
  END Tile_X11Y8_AD_SRAM4
  PIN Tile_X11Y8_AD_SRAM5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2288.240 2435.000 2288.840 ;
    END
  END Tile_X11Y8_AD_SRAM5
  PIN Tile_X11Y8_AD_SRAM6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2284.840 2435.000 2285.440 ;
    END
  END Tile_X11Y8_AD_SRAM6
  PIN Tile_X11Y8_AD_SRAM7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2046.840 2435.000 2047.440 ;
    END
  END Tile_X11Y8_AD_SRAM7
  PIN Tile_X11Y8_AD_SRAM8
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2281.440 2435.000 2282.040 ;
    END
  END Tile_X11Y8_AD_SRAM8
  PIN Tile_X11Y8_AD_SRAM9
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2057.040 2435.000 2057.640 ;
    END
  END Tile_X11Y8_AD_SRAM9
  PIN Tile_X11Y8_BEN_SRAM0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2278.040 2435.000 2278.640 ;
    END
  END Tile_X11Y8_BEN_SRAM0
  PIN Tile_X11Y8_BEN_SRAM1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2274.640 2435.000 2275.240 ;
    END
  END Tile_X11Y8_BEN_SRAM1
  PIN Tile_X11Y8_BEN_SRAM10
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2271.240 2435.000 2271.840 ;
    END
  END Tile_X11Y8_BEN_SRAM10
  PIN Tile_X11Y8_BEN_SRAM11
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2254.240 2435.000 2254.840 ;
    END
  END Tile_X11Y8_BEN_SRAM11
  PIN Tile_X11Y8_BEN_SRAM12
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2097.840 2435.000 2098.440 ;
    END
  END Tile_X11Y8_BEN_SRAM12
  PIN Tile_X11Y8_BEN_SRAM13
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2250.840 2435.000 2251.440 ;
    END
  END Tile_X11Y8_BEN_SRAM13
  PIN Tile_X11Y8_BEN_SRAM14
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2080.840 2435.000 2081.440 ;
    END
  END Tile_X11Y8_BEN_SRAM14
  PIN Tile_X11Y8_BEN_SRAM15
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2247.440 2435.000 2248.040 ;
    END
  END Tile_X11Y8_BEN_SRAM15
  PIN Tile_X11Y8_BEN_SRAM16
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2244.040 2435.000 2244.640 ;
    END
  END Tile_X11Y8_BEN_SRAM16
  PIN Tile_X11Y8_BEN_SRAM17
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2074.040 2435.000 2074.640 ;
    END
  END Tile_X11Y8_BEN_SRAM17
  PIN Tile_X11Y8_BEN_SRAM18
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2240.640 2435.000 2241.240 ;
    END
  END Tile_X11Y8_BEN_SRAM18
  PIN Tile_X11Y8_BEN_SRAM19
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2084.240 2435.000 2084.840 ;
    END
  END Tile_X11Y8_BEN_SRAM19
  PIN Tile_X11Y8_BEN_SRAM2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2053.640 2435.000 2054.240 ;
    END
  END Tile_X11Y8_BEN_SRAM2
  PIN Tile_X11Y8_BEN_SRAM20
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2237.240 2435.000 2237.840 ;
    END
  END Tile_X11Y8_BEN_SRAM20
  PIN Tile_X11Y8_BEN_SRAM21
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2233.840 2435.000 2234.440 ;
    END
  END Tile_X11Y8_BEN_SRAM21
  PIN Tile_X11Y8_BEN_SRAM22
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2193.040 2435.000 2193.640 ;
    END
  END Tile_X11Y8_BEN_SRAM22
  PIN Tile_X11Y8_BEN_SRAM23
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2230.440 2435.000 2231.040 ;
    END
  END Tile_X11Y8_BEN_SRAM23
  PIN Tile_X11Y8_BEN_SRAM24
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2091.040 2435.000 2091.640 ;
    END
  END Tile_X11Y8_BEN_SRAM24
  PIN Tile_X11Y8_BEN_SRAM25
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2227.040 2435.000 2227.640 ;
    END
  END Tile_X11Y8_BEN_SRAM25
  PIN Tile_X11Y8_BEN_SRAM26
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2223.640 2435.000 2224.240 ;
    END
  END Tile_X11Y8_BEN_SRAM26
  PIN Tile_X11Y8_BEN_SRAM27
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2087.640 2435.000 2088.240 ;
    END
  END Tile_X11Y8_BEN_SRAM27
  PIN Tile_X11Y8_BEN_SRAM28
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2220.240 2435.000 2220.840 ;
    END
  END Tile_X11Y8_BEN_SRAM28
  PIN Tile_X11Y8_BEN_SRAM29
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2295.040 2435.000 2295.640 ;
    END
  END Tile_X11Y8_BEN_SRAM29
  PIN Tile_X11Y8_BEN_SRAM3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2060.440 2435.000 2061.040 ;
    END
  END Tile_X11Y8_BEN_SRAM3
  PIN Tile_X11Y8_BEN_SRAM30
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2216.840 2435.000 2217.440 ;
    END
  END Tile_X11Y8_BEN_SRAM30
  PIN Tile_X11Y8_BEN_SRAM31
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2213.440 2435.000 2214.040 ;
    END
  END Tile_X11Y8_BEN_SRAM31
  PIN Tile_X11Y8_BEN_SRAM4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2067.240 2435.000 2067.840 ;
    END
  END Tile_X11Y8_BEN_SRAM4
  PIN Tile_X11Y8_BEN_SRAM5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2070.640 2435.000 2071.240 ;
    END
  END Tile_X11Y8_BEN_SRAM5
  PIN Tile_X11Y8_BEN_SRAM6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2063.840 2435.000 2064.440 ;
    END
  END Tile_X11Y8_BEN_SRAM6
  PIN Tile_X11Y8_BEN_SRAM7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2114.840 2435.000 2115.440 ;
    END
  END Tile_X11Y8_BEN_SRAM7
  PIN Tile_X11Y8_BEN_SRAM8
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2101.240 2435.000 2101.840 ;
    END
  END Tile_X11Y8_BEN_SRAM8
  PIN Tile_X11Y8_BEN_SRAM9
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2077.440 2435.000 2078.040 ;
    END
  END Tile_X11Y8_BEN_SRAM9
  PIN Tile_X11Y8_CLOCK_SRAM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2094.440 2435.000 2095.040 ;
    END
  END Tile_X11Y8_CLOCK_SRAM
  PIN Tile_X11Y8_DI_SRAM0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2210.040 2435.000 2210.640 ;
    END
  END Tile_X11Y8_DI_SRAM0
  PIN Tile_X11Y8_DI_SRAM1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2118.240 2435.000 2118.840 ;
    END
  END Tile_X11Y8_DI_SRAM1
  PIN Tile_X11Y8_DI_SRAM10
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2206.640 2435.000 2207.240 ;
    END
  END Tile_X11Y8_DI_SRAM10
  PIN Tile_X11Y8_DI_SRAM11
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2121.640 2435.000 2122.240 ;
    END
  END Tile_X11Y8_DI_SRAM11
  PIN Tile_X11Y8_DI_SRAM12
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2186.240 2435.000 2186.840 ;
    END
  END Tile_X11Y8_DI_SRAM12
  PIN Tile_X11Y8_DI_SRAM13
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2182.840 2435.000 2183.440 ;
    END
  END Tile_X11Y8_DI_SRAM13
  PIN Tile_X11Y8_DI_SRAM14
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2145.440 2435.000 2146.040 ;
    END
  END Tile_X11Y8_DI_SRAM14
  PIN Tile_X11Y8_DI_SRAM15
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2179.440 2435.000 2180.040 ;
    END
  END Tile_X11Y8_DI_SRAM15
  PIN Tile_X11Y8_DI_SRAM16
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2125.040 2435.000 2125.640 ;
    END
  END Tile_X11Y8_DI_SRAM16
  PIN Tile_X11Y8_DI_SRAM17
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2176.040 2435.000 2176.640 ;
    END
  END Tile_X11Y8_DI_SRAM17
  PIN Tile_X11Y8_DI_SRAM18
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2267.840 2435.000 2268.440 ;
    END
  END Tile_X11Y8_DI_SRAM18
  PIN Tile_X11Y8_DI_SRAM19
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2128.440 2435.000 2129.040 ;
    END
  END Tile_X11Y8_DI_SRAM19
  PIN Tile_X11Y8_DI_SRAM2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2142.040 2435.000 2142.640 ;
    END
  END Tile_X11Y8_DI_SRAM2
  PIN Tile_X11Y8_DI_SRAM20
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2264.440 2435.000 2265.040 ;
    END
  END Tile_X11Y8_DI_SRAM20
  PIN Tile_X11Y8_DI_SRAM21
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2189.640 2435.000 2190.240 ;
    END
  END Tile_X11Y8_DI_SRAM21
  PIN Tile_X11Y8_DI_SRAM22
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2165.840 2435.000 2166.440 ;
    END
  END Tile_X11Y8_DI_SRAM22
  PIN Tile_X11Y8_DI_SRAM23
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2162.440 2435.000 2163.040 ;
    END
  END Tile_X11Y8_DI_SRAM23
  PIN Tile_X11Y8_DI_SRAM24
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2199.840 2435.000 2200.440 ;
    END
  END Tile_X11Y8_DI_SRAM24
  PIN Tile_X11Y8_DI_SRAM25
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2159.040 2435.000 2159.640 ;
    END
  END Tile_X11Y8_DI_SRAM25
  PIN Tile_X11Y8_DI_SRAM26
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2131.840 2435.000 2132.440 ;
    END
  END Tile_X11Y8_DI_SRAM26
  PIN Tile_X11Y8_DI_SRAM27
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2155.640 2435.000 2156.240 ;
    END
  END Tile_X11Y8_DI_SRAM27
  PIN Tile_X11Y8_DI_SRAM28
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2152.240 2435.000 2152.840 ;
    END
  END Tile_X11Y8_DI_SRAM28
  PIN Tile_X11Y8_DI_SRAM29
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2135.240 2435.000 2135.840 ;
    END
  END Tile_X11Y8_DI_SRAM29
  PIN Tile_X11Y8_DI_SRAM3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2261.040 2435.000 2261.640 ;
    END
  END Tile_X11Y8_DI_SRAM3
  PIN Tile_X11Y8_DI_SRAM30
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2148.840 2435.000 2149.440 ;
    END
  END Tile_X11Y8_DI_SRAM30
  PIN Tile_X11Y8_DI_SRAM31
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2138.640 2435.000 2139.240 ;
    END
  END Tile_X11Y8_DI_SRAM31
  PIN Tile_X11Y8_DI_SRAM4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2203.240 2435.000 2203.840 ;
    END
  END Tile_X11Y8_DI_SRAM4
  PIN Tile_X11Y8_DI_SRAM5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2104.640 2435.000 2105.240 ;
    END
  END Tile_X11Y8_DI_SRAM5
  PIN Tile_X11Y8_DI_SRAM6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2108.040 2435.000 2108.640 ;
    END
  END Tile_X11Y8_DI_SRAM6
  PIN Tile_X11Y8_DI_SRAM7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2111.440 2435.000 2112.040 ;
    END
  END Tile_X11Y8_DI_SRAM7
  PIN Tile_X11Y8_DI_SRAM8
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2257.640 2435.000 2258.240 ;
    END
  END Tile_X11Y8_DI_SRAM8
  PIN Tile_X11Y8_DI_SRAM9
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2169.240 2435.000 2169.840 ;
    END
  END Tile_X11Y8_DI_SRAM9
  PIN Tile_X11Y8_DO_SRAM0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1931.240 2435.000 1931.840 ;
    END
  END Tile_X11Y8_DO_SRAM0
  PIN Tile_X11Y8_DO_SRAM1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1992.440 2435.000 1993.040 ;
    END
  END Tile_X11Y8_DO_SRAM1
  PIN Tile_X11Y8_DO_SRAM10
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2006.040 2435.000 2006.640 ;
    END
  END Tile_X11Y8_DO_SRAM10
  PIN Tile_X11Y8_DO_SRAM11
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1972.040 2435.000 1972.640 ;
    END
  END Tile_X11Y8_DO_SRAM11
  PIN Tile_X11Y8_DO_SRAM12
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2009.440 2435.000 2010.040 ;
    END
  END Tile_X11Y8_DO_SRAM12
  PIN Tile_X11Y8_DO_SRAM13
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1968.640 2435.000 1969.240 ;
    END
  END Tile_X11Y8_DO_SRAM13
  PIN Tile_X11Y8_DO_SRAM14
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1965.240 2435.000 1965.840 ;
    END
  END Tile_X11Y8_DO_SRAM14
  PIN Tile_X11Y8_DO_SRAM15
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2012.840 2435.000 2013.440 ;
    END
  END Tile_X11Y8_DO_SRAM15
  PIN Tile_X11Y8_DO_SRAM16
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1961.840 2435.000 1962.440 ;
    END
  END Tile_X11Y8_DO_SRAM16
  PIN Tile_X11Y8_DO_SRAM17
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2016.240 2435.000 2016.840 ;
    END
  END Tile_X11Y8_DO_SRAM17
  PIN Tile_X11Y8_DO_SRAM18
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1958.440 2435.000 1959.040 ;
    END
  END Tile_X11Y8_DO_SRAM18
  PIN Tile_X11Y8_DO_SRAM19
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1955.040 2435.000 1955.640 ;
    END
  END Tile_X11Y8_DO_SRAM19
  PIN Tile_X11Y8_DO_SRAM2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1995.840 2435.000 1996.440 ;
    END
  END Tile_X11Y8_DO_SRAM2
  PIN Tile_X11Y8_DO_SRAM20
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2019.640 2435.000 2020.240 ;
    END
  END Tile_X11Y8_DO_SRAM20
  PIN Tile_X11Y8_DO_SRAM21
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1951.640 2435.000 1952.240 ;
    END
  END Tile_X11Y8_DO_SRAM21
  PIN Tile_X11Y8_DO_SRAM22
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2023.040 2435.000 2023.640 ;
    END
  END Tile_X11Y8_DO_SRAM22
  PIN Tile_X11Y8_DO_SRAM23
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1948.240 2435.000 1948.840 ;
    END
  END Tile_X11Y8_DO_SRAM23
  PIN Tile_X11Y8_DO_SRAM24
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1944.840 2435.000 1945.440 ;
    END
  END Tile_X11Y8_DO_SRAM24
  PIN Tile_X11Y8_DO_SRAM25
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2026.440 2435.000 2027.040 ;
    END
  END Tile_X11Y8_DO_SRAM25
  PIN Tile_X11Y8_DO_SRAM26
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1941.440 2435.000 1942.040 ;
    END
  END Tile_X11Y8_DO_SRAM26
  PIN Tile_X11Y8_DO_SRAM27
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2029.840 2435.000 2030.440 ;
    END
  END Tile_X11Y8_DO_SRAM27
  PIN Tile_X11Y8_DO_SRAM28
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1938.040 2435.000 1938.640 ;
    END
  END Tile_X11Y8_DO_SRAM28
  PIN Tile_X11Y8_DO_SRAM29
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1934.640 2435.000 1935.240 ;
    END
  END Tile_X11Y8_DO_SRAM29
  PIN Tile_X11Y8_DO_SRAM3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1989.040 2435.000 1989.640 ;
    END
  END Tile_X11Y8_DO_SRAM3
  PIN Tile_X11Y8_DO_SRAM30
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2033.240 2435.000 2033.840 ;
    END
  END Tile_X11Y8_DO_SRAM30
  PIN Tile_X11Y8_DO_SRAM31
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2036.640 2435.000 2037.240 ;
    END
  END Tile_X11Y8_DO_SRAM31
  PIN Tile_X11Y8_DO_SRAM4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1985.640 2435.000 1986.240 ;
    END
  END Tile_X11Y8_DO_SRAM4
  PIN Tile_X11Y8_DO_SRAM5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1999.240 2435.000 1999.840 ;
    END
  END Tile_X11Y8_DO_SRAM5
  PIN Tile_X11Y8_DO_SRAM6
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1982.240 2435.000 1982.840 ;
    END
  END Tile_X11Y8_DO_SRAM6
  PIN Tile_X11Y8_DO_SRAM7
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2002.640 2435.000 2003.240 ;
    END
  END Tile_X11Y8_DO_SRAM7
  PIN Tile_X11Y8_DO_SRAM8
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1978.840 2435.000 1979.440 ;
    END
  END Tile_X11Y8_DO_SRAM8
  PIN Tile_X11Y8_DO_SRAM9
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 1975.440 2435.000 1976.040 ;
    END
  END Tile_X11Y8_DO_SRAM9
  PIN Tile_X11Y8_EN_SRAM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2196.440 2435.000 2197.040 ;
    END
  END Tile_X11Y8_EN_SRAM
  PIN Tile_X11Y8_R_WB_SRAM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 2431.000 2172.640 2435.000 2173.240 ;
    END
  END Tile_X11Y8_R_WB_SRAM
  PIN Tile_X1Y0_A_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 122.450 3778.500 122.730 3782.500 ;
    END
  END Tile_X1Y0_A_I_top
  PIN Tile_X1Y0_A_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 116.010 3778.500 116.290 3782.500 ;
    END
  END Tile_X1Y0_A_O_top
  PIN Tile_X1Y0_A_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 125.670 3778.500 125.950 3782.500 ;
    END
  END Tile_X1Y0_A_T_top
  PIN Tile_X1Y0_A_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 148.210 3778.500 148.490 3782.500 ;
    END
  END Tile_X1Y0_A_config_C_bit0
  PIN Tile_X1Y0_A_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 154.650 3778.500 154.930 3782.500 ;
    END
  END Tile_X1Y0_A_config_C_bit1
  PIN Tile_X1Y0_A_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 161.090 3778.500 161.370 3782.500 ;
    END
  END Tile_X1Y0_A_config_C_bit2
  PIN Tile_X1Y0_A_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 164.310 3778.500 164.590 3782.500 ;
    END
  END Tile_X1Y0_A_config_C_bit3
  PIN Tile_X1Y0_B_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 138.550 3778.500 138.830 3782.500 ;
    END
  END Tile_X1Y0_B_I_top
  PIN Tile_X1Y0_B_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 132.110 3778.500 132.390 3782.500 ;
    END
  END Tile_X1Y0_B_O_top
  PIN Tile_X1Y0_B_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 144.990 3778.500 145.270 3782.500 ;
    END
  END Tile_X1Y0_B_T_top
  PIN Tile_X1Y0_B_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 170.750 3778.500 171.030 3782.500 ;
    END
  END Tile_X1Y0_B_config_C_bit0
  PIN Tile_X1Y0_B_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 177.190 3778.500 177.470 3782.500 ;
    END
  END Tile_X1Y0_B_config_C_bit1
  PIN Tile_X1Y0_B_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 180.410 3778.500 180.690 3782.500 ;
    END
  END Tile_X1Y0_B_config_C_bit2
  PIN Tile_X1Y0_B_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 186.850 3778.500 187.130 3782.500 ;
    END
  END Tile_X1Y0_B_config_C_bit3
  PIN Tile_X1Y17_IRQ_top0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 116.010 0.000 116.290 4.000 ;
    END
  END Tile_X1Y17_IRQ_top0
  PIN Tile_X1Y17_IRQ_top1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 122.450 0.000 122.730 4.000 ;
    END
  END Tile_X1Y17_IRQ_top1
  PIN Tile_X1Y17_IRQ_top2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 128.890 0.000 129.170 4.000 ;
    END
  END Tile_X1Y17_IRQ_top2
  PIN Tile_X1Y17_IRQ_top3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 138.550 0.000 138.830 4.000 ;
    END
  END Tile_X1Y17_IRQ_top3
  PIN Tile_X2Y0_A_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 325.310 3778.500 325.590 3782.500 ;
    END
  END Tile_X2Y0_A_I_top
  PIN Tile_X2Y0_A_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 318.870 3778.500 319.150 3782.500 ;
    END
  END Tile_X2Y0_A_O_top
  PIN Tile_X2Y0_A_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 331.750 3778.500 332.030 3782.500 ;
    END
  END Tile_X2Y0_A_T_top
  PIN Tile_X2Y0_A_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 354.290 3778.500 354.570 3782.500 ;
    END
  END Tile_X2Y0_A_config_C_bit0
  PIN Tile_X2Y0_A_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 357.510 3778.500 357.790 3782.500 ;
    END
  END Tile_X2Y0_A_config_C_bit1
  PIN Tile_X2Y0_A_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 363.950 3778.500 364.230 3782.500 ;
    END
  END Tile_X2Y0_A_config_C_bit2
  PIN Tile_X2Y0_A_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 370.390 3778.500 370.670 3782.500 ;
    END
  END Tile_X2Y0_A_config_C_bit3
  PIN Tile_X2Y0_B_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 341.410 3778.500 341.690 3782.500 ;
    END
  END Tile_X2Y0_B_I_top
  PIN Tile_X2Y0_B_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 334.970 3778.500 335.250 3782.500 ;
    END
  END Tile_X2Y0_B_O_top
  PIN Tile_X2Y0_B_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 347.850 3778.500 348.130 3782.500 ;
    END
  END Tile_X2Y0_B_T_top
  PIN Tile_X2Y0_B_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 373.610 3778.500 373.890 3782.500 ;
    END
  END Tile_X2Y0_B_config_C_bit0
  PIN Tile_X2Y0_B_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 380.050 3778.500 380.330 3782.500 ;
    END
  END Tile_X2Y0_B_config_C_bit1
  PIN Tile_X2Y0_B_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 386.490 3778.500 386.770 3782.500 ;
    END
  END Tile_X2Y0_B_config_C_bit2
  PIN Tile_X2Y0_B_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 392.930 3778.500 393.210 3782.500 ;
    END
  END Tile_X2Y0_B_config_C_bit3
  PIN Tile_X2Y17_BOOT_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 325.310 0.000 325.590 4.000 ;
    END
  END Tile_X2Y17_BOOT_top
  PIN Tile_X2Y17_RESET_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 318.870 0.000 319.150 4.000 ;
    END
  END Tile_X2Y17_RESET_top
  PIN Tile_X2Y17_SLOT_top0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 331.750 0.000 332.030 4.000 ;
    END
  END Tile_X2Y17_SLOT_top0
  PIN Tile_X2Y17_SLOT_top1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 341.410 0.000 341.690 4.000 ;
    END
  END Tile_X2Y17_SLOT_top1
  PIN Tile_X2Y17_SLOT_top2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 347.850 0.000 348.130 4.000 ;
    END
  END Tile_X2Y17_SLOT_top2
  PIN Tile_X2Y17_SLOT_top3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 354.290 0.000 354.570 4.000 ;
    END
  END Tile_X2Y17_SLOT_top3
  PIN Tile_X4Y0_A_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 776.110 3778.500 776.390 3782.500 ;
    END
  END Tile_X4Y0_A_I_top
  PIN Tile_X4Y0_A_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 769.670 3778.500 769.950 3782.500 ;
    END
  END Tile_X4Y0_A_O_top
  PIN Tile_X4Y0_A_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 779.330 3778.500 779.610 3782.500 ;
    END
  END Tile_X4Y0_A_T_top
  PIN Tile_X4Y0_A_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 801.870 3778.500 802.150 3782.500 ;
    END
  END Tile_X4Y0_A_config_C_bit0
  PIN Tile_X4Y0_A_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 808.310 3778.500 808.590 3782.500 ;
    END
  END Tile_X4Y0_A_config_C_bit1
  PIN Tile_X4Y0_A_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 814.750 3778.500 815.030 3782.500 ;
    END
  END Tile_X4Y0_A_config_C_bit2
  PIN Tile_X4Y0_A_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 817.970 3778.500 818.250 3782.500 ;
    END
  END Tile_X4Y0_A_config_C_bit3
  PIN Tile_X4Y0_B_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 792.210 3778.500 792.490 3782.500 ;
    END
  END Tile_X4Y0_B_I_top
  PIN Tile_X4Y0_B_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 785.770 3778.500 786.050 3782.500 ;
    END
  END Tile_X4Y0_B_O_top
  PIN Tile_X4Y0_B_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 798.650 3778.500 798.930 3782.500 ;
    END
  END Tile_X4Y0_B_T_top
  PIN Tile_X4Y0_B_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 824.410 3778.500 824.690 3782.500 ;
    END
  END Tile_X4Y0_B_config_C_bit0
  PIN Tile_X4Y0_B_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 830.850 3778.500 831.130 3782.500 ;
    END
  END Tile_X4Y0_B_config_C_bit1
  PIN Tile_X4Y0_B_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 837.290 3778.500 837.570 3782.500 ;
    END
  END Tile_X4Y0_B_config_C_bit2
  PIN Tile_X4Y0_B_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 840.510 3778.500 840.790 3782.500 ;
    END
  END Tile_X4Y0_B_config_C_bit3
  PIN Tile_X4Y17_I_top0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 827.630 0.000 827.910 4.000 ;
    END
  END Tile_X4Y17_I_top0
  PIN Tile_X4Y17_I_top1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 830.850 0.000 831.130 4.000 ;
    END
  END Tile_X4Y17_I_top1
  PIN Tile_X4Y17_I_top10
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 863.050 0.000 863.330 4.000 ;
    END
  END Tile_X4Y17_I_top10
  PIN Tile_X4Y17_I_top11
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 866.270 0.000 866.550 4.000 ;
    END
  END Tile_X4Y17_I_top11
  PIN Tile_X4Y17_I_top12
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 869.490 0.000 869.770 4.000 ;
    END
  END Tile_X4Y17_I_top12
  PIN Tile_X4Y17_I_top13
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 875.930 0.000 876.210 4.000 ;
    END
  END Tile_X4Y17_I_top13
  PIN Tile_X4Y17_I_top14
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 879.150 0.000 879.430 4.000 ;
    END
  END Tile_X4Y17_I_top14
  PIN Tile_X4Y17_I_top15
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 882.370 0.000 882.650 4.000 ;
    END
  END Tile_X4Y17_I_top15
  PIN Tile_X4Y17_I_top2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 834.070 0.000 834.350 4.000 ;
    END
  END Tile_X4Y17_I_top2
  PIN Tile_X4Y17_I_top3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 837.290 0.000 837.570 4.000 ;
    END
  END Tile_X4Y17_I_top3
  PIN Tile_X4Y17_I_top4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 840.510 0.000 840.790 4.000 ;
    END
  END Tile_X4Y17_I_top4
  PIN Tile_X4Y17_I_top5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 843.730 0.000 844.010 4.000 ;
    END
  END Tile_X4Y17_I_top5
  PIN Tile_X4Y17_I_top6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 850.170 0.000 850.450 4.000 ;
    END
  END Tile_X4Y17_I_top6
  PIN Tile_X4Y17_I_top7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 853.390 0.000 853.670 4.000 ;
    END
  END Tile_X4Y17_I_top7
  PIN Tile_X4Y17_I_top8
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 856.610 0.000 856.890 4.000 ;
    END
  END Tile_X4Y17_I_top8
  PIN Tile_X4Y17_I_top9
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 859.830 0.000 860.110 4.000 ;
    END
  END Tile_X4Y17_I_top9
  PIN Tile_X4Y17_O_top0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 766.450 0.000 766.730 4.000 ;
    END
  END Tile_X4Y17_O_top0
  PIN Tile_X4Y17_O_top1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 772.890 0.000 773.170 4.000 ;
    END
  END Tile_X4Y17_O_top1
  PIN Tile_X4Y17_O_top10
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 805.090 0.000 805.370 4.000 ;
    END
  END Tile_X4Y17_O_top10
  PIN Tile_X4Y17_O_top11
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 808.310 0.000 808.590 4.000 ;
    END
  END Tile_X4Y17_O_top11
  PIN Tile_X4Y17_O_top12
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 811.530 0.000 811.810 4.000 ;
    END
  END Tile_X4Y17_O_top12
  PIN Tile_X4Y17_O_top13
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 814.750 0.000 815.030 4.000 ;
    END
  END Tile_X4Y17_O_top13
  PIN Tile_X4Y17_O_top14
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 817.970 0.000 818.250 4.000 ;
    END
  END Tile_X4Y17_O_top14
  PIN Tile_X4Y17_O_top15
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 824.410 0.000 824.690 4.000 ;
    END
  END Tile_X4Y17_O_top15
  PIN Tile_X4Y17_O_top2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 776.110 0.000 776.390 4.000 ;
    END
  END Tile_X4Y17_O_top2
  PIN Tile_X4Y17_O_top3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 779.330 0.000 779.610 4.000 ;
    END
  END Tile_X4Y17_O_top3
  PIN Tile_X4Y17_O_top4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 782.550 0.000 782.830 4.000 ;
    END
  END Tile_X4Y17_O_top4
  PIN Tile_X4Y17_O_top5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 785.770 0.000 786.050 4.000 ;
    END
  END Tile_X4Y17_O_top5
  PIN Tile_X4Y17_O_top6
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 788.990 0.000 789.270 4.000 ;
    END
  END Tile_X4Y17_O_top6
  PIN Tile_X4Y17_O_top7
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 792.210 0.000 792.490 4.000 ;
    END
  END Tile_X4Y17_O_top7
  PIN Tile_X4Y17_O_top8
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 798.650 0.000 798.930 4.000 ;
    END
  END Tile_X4Y17_O_top8
  PIN Tile_X4Y17_O_top9
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 801.870 0.000 802.150 4.000 ;
    END
  END Tile_X4Y17_O_top9
  PIN Tile_X5Y0_A_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 978.970 3778.500 979.250 3782.500 ;
    END
  END Tile_X5Y0_A_I_top
  PIN Tile_X5Y0_A_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 975.750 3778.500 976.030 3782.500 ;
    END
  END Tile_X5Y0_A_O_top
  PIN Tile_X5Y0_A_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 985.410 3778.500 985.690 3782.500 ;
    END
  END Tile_X5Y0_A_T_top
  PIN Tile_X5Y0_A_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1007.950 3778.500 1008.230 3782.500 ;
    END
  END Tile_X5Y0_A_config_C_bit0
  PIN Tile_X5Y0_A_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1014.390 3778.500 1014.670 3782.500 ;
    END
  END Tile_X5Y0_A_config_C_bit1
  PIN Tile_X5Y0_A_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1017.610 3778.500 1017.890 3782.500 ;
    END
  END Tile_X5Y0_A_config_C_bit2
  PIN Tile_X5Y0_A_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1024.050 3778.500 1024.330 3782.500 ;
    END
  END Tile_X5Y0_A_config_C_bit3
  PIN Tile_X5Y0_B_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 998.290 3778.500 998.570 3782.500 ;
    END
  END Tile_X5Y0_B_I_top
  PIN Tile_X5Y0_B_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 991.850 3778.500 992.130 3782.500 ;
    END
  END Tile_X5Y0_B_O_top
  PIN Tile_X5Y0_B_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1001.510 3778.500 1001.790 3782.500 ;
    END
  END Tile_X5Y0_B_T_top
  PIN Tile_X5Y0_B_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1030.490 3778.500 1030.770 3782.500 ;
    END
  END Tile_X5Y0_B_config_C_bit0
  PIN Tile_X5Y0_B_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1036.930 3778.500 1037.210 3782.500 ;
    END
  END Tile_X5Y0_B_config_C_bit1
  PIN Tile_X5Y0_B_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1040.150 3778.500 1040.430 3782.500 ;
    END
  END Tile_X5Y0_B_config_C_bit2
  PIN Tile_X5Y0_B_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1046.590 3778.500 1046.870 3782.500 ;
    END
  END Tile_X5Y0_B_config_C_bit3
  PIN Tile_X5Y17_I_top0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1030.490 0.000 1030.770 4.000 ;
    END
  END Tile_X5Y17_I_top0
  PIN Tile_X5Y17_I_top1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1036.930 0.000 1037.210 4.000 ;
    END
  END Tile_X5Y17_I_top1
  PIN Tile_X5Y17_I_top10
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1069.130 0.000 1069.410 4.000 ;
    END
  END Tile_X5Y17_I_top10
  PIN Tile_X5Y17_I_top11
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1072.350 0.000 1072.630 4.000 ;
    END
  END Tile_X5Y17_I_top11
  PIN Tile_X5Y17_I_top12
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1075.570 0.000 1075.850 4.000 ;
    END
  END Tile_X5Y17_I_top12
  PIN Tile_X5Y17_I_top13
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1078.790 0.000 1079.070 4.000 ;
    END
  END Tile_X5Y17_I_top13
  PIN Tile_X5Y17_I_top14
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1082.010 0.000 1082.290 4.000 ;
    END
  END Tile_X5Y17_I_top14
  PIN Tile_X5Y17_I_top15
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1088.450 0.000 1088.730 4.000 ;
    END
  END Tile_X5Y17_I_top15
  PIN Tile_X5Y17_I_top2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1040.150 0.000 1040.430 4.000 ;
    END
  END Tile_X5Y17_I_top2
  PIN Tile_X5Y17_I_top3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1043.370 0.000 1043.650 4.000 ;
    END
  END Tile_X5Y17_I_top3
  PIN Tile_X5Y17_I_top4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1046.590 0.000 1046.870 4.000 ;
    END
  END Tile_X5Y17_I_top4
  PIN Tile_X5Y17_I_top5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1049.810 0.000 1050.090 4.000 ;
    END
  END Tile_X5Y17_I_top5
  PIN Tile_X5Y17_I_top6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1053.030 0.000 1053.310 4.000 ;
    END
  END Tile_X5Y17_I_top6
  PIN Tile_X5Y17_I_top7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1056.250 0.000 1056.530 4.000 ;
    END
  END Tile_X5Y17_I_top7
  PIN Tile_X5Y17_I_top8
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1062.690 0.000 1062.970 4.000 ;
    END
  END Tile_X5Y17_I_top8
  PIN Tile_X5Y17_I_top9
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1065.910 0.000 1066.190 4.000 ;
    END
  END Tile_X5Y17_I_top9
  PIN Tile_X5Y17_O_top0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 972.530 0.000 972.810 4.000 ;
    END
  END Tile_X5Y17_O_top0
  PIN Tile_X5Y17_O_top1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 975.750 0.000 976.030 4.000 ;
    END
  END Tile_X5Y17_O_top1
  PIN Tile_X5Y17_O_top10
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 1011.170 0.000 1011.450 4.000 ;
    END
  END Tile_X5Y17_O_top10
  PIN Tile_X5Y17_O_top11
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1014.390 0.000 1014.670 4.000 ;
    END
  END Tile_X5Y17_O_top11
  PIN Tile_X5Y17_O_top12
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1017.610 0.000 1017.890 4.000 ;
    END
  END Tile_X5Y17_O_top12
  PIN Tile_X5Y17_O_top13
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1020.830 0.000 1021.110 4.000 ;
    END
  END Tile_X5Y17_O_top13
  PIN Tile_X5Y17_O_top14
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 1024.050 0.000 1024.330 4.000 ;
    END
  END Tile_X5Y17_O_top14
  PIN Tile_X5Y17_O_top15
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1027.270 0.000 1027.550 4.000 ;
    END
  END Tile_X5Y17_O_top15
  PIN Tile_X5Y17_O_top2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 978.970 0.000 979.250 4.000 ;
    END
  END Tile_X5Y17_O_top2
  PIN Tile_X5Y17_O_top3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 985.410 0.000 985.690 4.000 ;
    END
  END Tile_X5Y17_O_top3
  PIN Tile_X5Y17_O_top4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 988.630 0.000 988.910 4.000 ;
    END
  END Tile_X5Y17_O_top4
  PIN Tile_X5Y17_O_top5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 991.850 0.000 992.130 4.000 ;
    END
  END Tile_X5Y17_O_top5
  PIN Tile_X5Y17_O_top6
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 995.070 0.000 995.350 4.000 ;
    END
  END Tile_X5Y17_O_top6
  PIN Tile_X5Y17_O_top7
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 998.290 0.000 998.570 4.000 ;
    END
  END Tile_X5Y17_O_top7
  PIN Tile_X5Y17_O_top8
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1001.510 0.000 1001.790 4.000 ;
    END
  END Tile_X5Y17_O_top8
  PIN Tile_X5Y17_O_top9
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1004.730 0.000 1005.010 4.000 ;
    END
  END Tile_X5Y17_O_top9
  PIN Tile_X6Y0_A_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1185.050 3778.500 1185.330 3782.500 ;
    END
  END Tile_X6Y0_A_I_top
  PIN Tile_X6Y0_A_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 1178.610 3778.500 1178.890 3782.500 ;
    END
  END Tile_X6Y0_A_O_top
  PIN Tile_X6Y0_A_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1191.490 3778.500 1191.770 3782.500 ;
    END
  END Tile_X6Y0_A_T_top
  PIN Tile_X6Y0_A_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1214.030 3778.500 1214.310 3782.500 ;
    END
  END Tile_X6Y0_A_config_C_bit0
  PIN Tile_X6Y0_A_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1217.250 3778.500 1217.530 3782.500 ;
    END
  END Tile_X6Y0_A_config_C_bit1
  PIN Tile_X6Y0_A_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1223.690 3778.500 1223.970 3782.500 ;
    END
  END Tile_X6Y0_A_config_C_bit2
  PIN Tile_X6Y0_A_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1230.130 3778.500 1230.410 3782.500 ;
    END
  END Tile_X6Y0_A_config_C_bit3
  PIN Tile_X6Y0_B_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1201.150 3778.500 1201.430 3782.500 ;
    END
  END Tile_X6Y0_B_I_top
  PIN Tile_X6Y0_B_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 1194.710 3778.500 1194.990 3782.500 ;
    END
  END Tile_X6Y0_B_O_top
  PIN Tile_X6Y0_B_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1207.590 3778.500 1207.870 3782.500 ;
    END
  END Tile_X6Y0_B_T_top
  PIN Tile_X6Y0_B_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1233.350 3778.500 1233.630 3782.500 ;
    END
  END Tile_X6Y0_B_config_C_bit0
  PIN Tile_X6Y0_B_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1239.790 3778.500 1240.070 3782.500 ;
    END
  END Tile_X6Y0_B_config_C_bit1
  PIN Tile_X6Y0_B_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1246.230 3778.500 1246.510 3782.500 ;
    END
  END Tile_X6Y0_B_config_C_bit2
  PIN Tile_X6Y0_B_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1252.670 3778.500 1252.950 3782.500 ;
    END
  END Tile_X6Y0_B_config_C_bit3
  PIN Tile_X6Y17_I_top0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1236.570 0.000 1236.850 4.000 ;
    END
  END Tile_X6Y17_I_top0
  PIN Tile_X6Y17_I_top1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1239.790 0.000 1240.070 4.000 ;
    END
  END Tile_X6Y17_I_top1
  PIN Tile_X6Y17_I_top10
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1271.990 0.000 1272.270 4.000 ;
    END
  END Tile_X6Y17_I_top10
  PIN Tile_X6Y17_I_top11
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1278.430 0.000 1278.710 4.000 ;
    END
  END Tile_X6Y17_I_top11
  PIN Tile_X6Y17_I_top12
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1281.650 0.000 1281.930 4.000 ;
    END
  END Tile_X6Y17_I_top12
  PIN Tile_X6Y17_I_top13
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1284.870 0.000 1285.150 4.000 ;
    END
  END Tile_X6Y17_I_top13
  PIN Tile_X6Y17_I_top14
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1288.090 0.000 1288.370 4.000 ;
    END
  END Tile_X6Y17_I_top14
  PIN Tile_X6Y17_I_top15
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1291.310 0.000 1291.590 4.000 ;
    END
  END Tile_X6Y17_I_top15
  PIN Tile_X6Y17_I_top2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1243.010 0.000 1243.290 4.000 ;
    END
  END Tile_X6Y17_I_top2
  PIN Tile_X6Y17_I_top3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1246.230 0.000 1246.510 4.000 ;
    END
  END Tile_X6Y17_I_top3
  PIN Tile_X6Y17_I_top4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1252.670 0.000 1252.950 4.000 ;
    END
  END Tile_X6Y17_I_top4
  PIN Tile_X6Y17_I_top5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1255.890 0.000 1256.170 4.000 ;
    END
  END Tile_X6Y17_I_top5
  PIN Tile_X6Y17_I_top6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1259.110 0.000 1259.390 4.000 ;
    END
  END Tile_X6Y17_I_top6
  PIN Tile_X6Y17_I_top7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1262.330 0.000 1262.610 4.000 ;
    END
  END Tile_X6Y17_I_top7
  PIN Tile_X6Y17_I_top8
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1265.550 0.000 1265.830 4.000 ;
    END
  END Tile_X6Y17_I_top8
  PIN Tile_X6Y17_I_top9
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1268.770 0.000 1269.050 4.000 ;
    END
  END Tile_X6Y17_I_top9
  PIN Tile_X6Y17_O_top0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1178.610 0.000 1178.890 4.000 ;
    END
  END Tile_X6Y17_O_top0
  PIN Tile_X6Y17_O_top1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1181.830 0.000 1182.110 4.000 ;
    END
  END Tile_X6Y17_O_top1
  PIN Tile_X6Y17_O_top10
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 1214.030 0.000 1214.310 4.000 ;
    END
  END Tile_X6Y17_O_top10
  PIN Tile_X6Y17_O_top11
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1217.250 0.000 1217.530 4.000 ;
    END
  END Tile_X6Y17_O_top11
  PIN Tile_X6Y17_O_top12
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1220.470 0.000 1220.750 4.000 ;
    END
  END Tile_X6Y17_O_top12
  PIN Tile_X6Y17_O_top13
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1226.910 0.000 1227.190 4.000 ;
    END
  END Tile_X6Y17_O_top13
  PIN Tile_X6Y17_O_top14
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 1230.130 0.000 1230.410 4.000 ;
    END
  END Tile_X6Y17_O_top14
  PIN Tile_X6Y17_O_top15
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1233.350 0.000 1233.630 4.000 ;
    END
  END Tile_X6Y17_O_top15
  PIN Tile_X6Y17_O_top2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 1185.050 0.000 1185.330 4.000 ;
    END
  END Tile_X6Y17_O_top2
  PIN Tile_X6Y17_O_top3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 1188.270 0.000 1188.550 4.000 ;
    END
  END Tile_X6Y17_O_top3
  PIN Tile_X6Y17_O_top4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1191.490 0.000 1191.770 4.000 ;
    END
  END Tile_X6Y17_O_top4
  PIN Tile_X6Y17_O_top5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1194.710 0.000 1194.990 4.000 ;
    END
  END Tile_X6Y17_O_top5
  PIN Tile_X6Y17_O_top6
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 1201.150 0.000 1201.430 4.000 ;
    END
  END Tile_X6Y17_O_top6
  PIN Tile_X6Y17_O_top7
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1204.370 0.000 1204.650 4.000 ;
    END
  END Tile_X6Y17_O_top7
  PIN Tile_X6Y17_O_top8
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1207.590 0.000 1207.870 4.000 ;
    END
  END Tile_X6Y17_O_top8
  PIN Tile_X6Y17_O_top9
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1210.810 0.000 1211.090 4.000 ;
    END
  END Tile_X6Y17_O_top9
  PIN Tile_X8Y0_A_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1616.530 3778.500 1616.810 3782.500 ;
    END
  END Tile_X8Y0_A_I_top
  PIN Tile_X8Y0_A_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 1610.090 3778.500 1610.370 3782.500 ;
    END
  END Tile_X8Y0_A_O_top
  PIN Tile_X8Y0_A_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1619.750 3778.500 1620.030 3782.500 ;
    END
  END Tile_X8Y0_A_T_top
  PIN Tile_X8Y0_A_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1642.290 3778.500 1642.570 3782.500 ;
    END
  END Tile_X8Y0_A_config_C_bit0
  PIN Tile_X8Y0_A_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1648.730 3778.500 1649.010 3782.500 ;
    END
  END Tile_X8Y0_A_config_C_bit1
  PIN Tile_X8Y0_A_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1655.170 3778.500 1655.450 3782.500 ;
    END
  END Tile_X8Y0_A_config_C_bit2
  PIN Tile_X8Y0_A_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1658.390 3778.500 1658.670 3782.500 ;
    END
  END Tile_X8Y0_A_config_C_bit3
  PIN Tile_X8Y0_B_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1632.630 3778.500 1632.910 3782.500 ;
    END
  END Tile_X8Y0_B_I_top
  PIN Tile_X8Y0_B_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 1626.190 3778.500 1626.470 3782.500 ;
    END
  END Tile_X8Y0_B_O_top
  PIN Tile_X8Y0_B_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1635.850 3778.500 1636.130 3782.500 ;
    END
  END Tile_X8Y0_B_T_top
  PIN Tile_X8Y0_B_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1664.830 3778.500 1665.110 3782.500 ;
    END
  END Tile_X8Y0_B_config_C_bit0
  PIN Tile_X8Y0_B_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1671.270 3778.500 1671.550 3782.500 ;
    END
  END Tile_X8Y0_B_config_C_bit1
  PIN Tile_X8Y0_B_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1674.490 3778.500 1674.770 3782.500 ;
    END
  END Tile_X8Y0_B_config_C_bit2
  PIN Tile_X8Y0_B_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1680.930 3778.500 1681.210 3782.500 ;
    END
  END Tile_X8Y0_B_config_C_bit3
  PIN Tile_X8Y17_I_top0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1668.050 0.000 1668.330 4.000 ;
    END
  END Tile_X8Y17_I_top0
  PIN Tile_X8Y17_I_top1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1671.270 0.000 1671.550 4.000 ;
    END
  END Tile_X8Y17_I_top1
  PIN Tile_X8Y17_I_top10
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1703.470 0.000 1703.750 4.000 ;
    END
  END Tile_X8Y17_I_top10
  PIN Tile_X8Y17_I_top11
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1706.690 0.000 1706.970 4.000 ;
    END
  END Tile_X8Y17_I_top11
  PIN Tile_X8Y17_I_top12
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1709.910 0.000 1710.190 4.000 ;
    END
  END Tile_X8Y17_I_top12
  PIN Tile_X8Y17_I_top13
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1713.130 0.000 1713.410 4.000 ;
    END
  END Tile_X8Y17_I_top13
  PIN Tile_X8Y17_I_top14
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1719.570 0.000 1719.850 4.000 ;
    END
  END Tile_X8Y17_I_top14
  PIN Tile_X8Y17_I_top15
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1722.790 0.000 1723.070 4.000 ;
    END
  END Tile_X8Y17_I_top15
  PIN Tile_X8Y17_I_top2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1674.490 0.000 1674.770 4.000 ;
    END
  END Tile_X8Y17_I_top2
  PIN Tile_X8Y17_I_top3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1677.710 0.000 1677.990 4.000 ;
    END
  END Tile_X8Y17_I_top3
  PIN Tile_X8Y17_I_top4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1680.930 0.000 1681.210 4.000 ;
    END
  END Tile_X8Y17_I_top4
  PIN Tile_X8Y17_I_top5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1684.150 0.000 1684.430 4.000 ;
    END
  END Tile_X8Y17_I_top5
  PIN Tile_X8Y17_I_top6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1687.370 0.000 1687.650 4.000 ;
    END
  END Tile_X8Y17_I_top6
  PIN Tile_X8Y17_I_top7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1693.810 0.000 1694.090 4.000 ;
    END
  END Tile_X8Y17_I_top7
  PIN Tile_X8Y17_I_top8
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1697.030 0.000 1697.310 4.000 ;
    END
  END Tile_X8Y17_I_top8
  PIN Tile_X8Y17_I_top9
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1700.250 0.000 1700.530 4.000 ;
    END
  END Tile_X8Y17_I_top9
  PIN Tile_X8Y17_O_top0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1606.870 0.000 1607.150 4.000 ;
    END
  END Tile_X8Y17_O_top0
  PIN Tile_X8Y17_O_top1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1610.090 0.000 1610.370 4.000 ;
    END
  END Tile_X8Y17_O_top1
  PIN Tile_X8Y17_O_top10
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 1645.510 0.000 1645.790 4.000 ;
    END
  END Tile_X8Y17_O_top10
  PIN Tile_X8Y17_O_top11
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1648.730 0.000 1649.010 4.000 ;
    END
  END Tile_X8Y17_O_top11
  PIN Tile_X8Y17_O_top12
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1651.950 0.000 1652.230 4.000 ;
    END
  END Tile_X8Y17_O_top12
  PIN Tile_X8Y17_O_top13
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1655.170 0.000 1655.450 4.000 ;
    END
  END Tile_X8Y17_O_top13
  PIN Tile_X8Y17_O_top14
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 1658.390 0.000 1658.670 4.000 ;
    END
  END Tile_X8Y17_O_top14
  PIN Tile_X8Y17_O_top15
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1661.610 0.000 1661.890 4.000 ;
    END
  END Tile_X8Y17_O_top15
  PIN Tile_X8Y17_O_top2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 1616.530 0.000 1616.810 4.000 ;
    END
  END Tile_X8Y17_O_top2
  PIN Tile_X8Y17_O_top3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 1619.750 0.000 1620.030 4.000 ;
    END
  END Tile_X8Y17_O_top3
  PIN Tile_X8Y17_O_top4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1622.970 0.000 1623.250 4.000 ;
    END
  END Tile_X8Y17_O_top4
  PIN Tile_X8Y17_O_top5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1626.190 0.000 1626.470 4.000 ;
    END
  END Tile_X8Y17_O_top5
  PIN Tile_X8Y17_O_top6
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 1629.410 0.000 1629.690 4.000 ;
    END
  END Tile_X8Y17_O_top6
  PIN Tile_X8Y17_O_top7
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1632.630 0.000 1632.910 4.000 ;
    END
  END Tile_X8Y17_O_top7
  PIN Tile_X8Y17_O_top8
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1635.850 0.000 1636.130 4.000 ;
    END
  END Tile_X8Y17_O_top8
  PIN Tile_X8Y17_O_top9
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1642.290 0.000 1642.570 4.000 ;
    END
  END Tile_X8Y17_O_top9
  PIN Tile_X9Y0_A_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1819.390 3778.500 1819.670 3782.500 ;
    END
  END Tile_X9Y0_A_I_top
  PIN Tile_X9Y0_A_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 1816.170 3778.500 1816.450 3782.500 ;
    END
  END Tile_X9Y0_A_O_top
  PIN Tile_X9Y0_A_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1825.830 3778.500 1826.110 3782.500 ;
    END
  END Tile_X9Y0_A_T_top
  PIN Tile_X9Y0_A_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1848.370 3778.500 1848.650 3782.500 ;
    END
  END Tile_X9Y0_A_config_C_bit0
  PIN Tile_X9Y0_A_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1854.810 3778.500 1855.090 3782.500 ;
    END
  END Tile_X9Y0_A_config_C_bit1
  PIN Tile_X9Y0_A_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1858.030 3778.500 1858.310 3782.500 ;
    END
  END Tile_X9Y0_A_config_C_bit2
  PIN Tile_X9Y0_A_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1864.470 3778.500 1864.750 3782.500 ;
    END
  END Tile_X9Y0_A_config_C_bit3
  PIN Tile_X9Y0_B_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1835.490 3778.500 1835.770 3782.500 ;
    END
  END Tile_X9Y0_B_I_top
  PIN Tile_X9Y0_B_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 1832.270 3778.500 1832.550 3782.500 ;
    END
  END Tile_X9Y0_B_O_top
  PIN Tile_X9Y0_B_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1841.930 3778.500 1842.210 3782.500 ;
    END
  END Tile_X9Y0_B_T_top
  PIN Tile_X9Y0_B_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1870.910 3778.500 1871.190 3782.500 ;
    END
  END Tile_X9Y0_B_config_C_bit0
  PIN Tile_X9Y0_B_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1874.130 3778.500 1874.410 3782.500 ;
    END
  END Tile_X9Y0_B_config_C_bit1
  PIN Tile_X9Y0_B_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1880.570 3778.500 1880.850 3782.500 ;
    END
  END Tile_X9Y0_B_config_C_bit2
  PIN Tile_X9Y0_B_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1887.010 3778.500 1887.290 3782.500 ;
    END
  END Tile_X9Y0_B_config_C_bit3
  PIN Tile_X9Y17_CMP_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1812.950 0.000 1813.230 4.000 ;
    END
  END Tile_X9Y17_CMP_top
  PIN Tile_X9Y17_HOLD_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1816.170 0.000 1816.450 4.000 ;
    END
  END Tile_X9Y17_HOLD_top
  PIN Tile_X9Y17_RESET_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1822.610 0.000 1822.890 4.000 ;
    END
  END Tile_X9Y17_RESET_top
  PIN Tile_X9Y17_VALUE_top0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1829.050 0.000 1829.330 4.000 ;
    END
  END Tile_X9Y17_VALUE_top0
  PIN Tile_X9Y17_VALUE_top1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1835.490 0.000 1835.770 4.000 ;
    END
  END Tile_X9Y17_VALUE_top1
  PIN Tile_X9Y17_VALUE_top10
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1883.790 0.000 1884.070 4.000 ;
    END
  END Tile_X9Y17_VALUE_top10
  PIN Tile_X9Y17_VALUE_top11
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1890.230 0.000 1890.510 4.000 ;
    END
  END Tile_X9Y17_VALUE_top11
  PIN Tile_X9Y17_VALUE_top2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1838.710 0.000 1838.990 4.000 ;
    END
  END Tile_X9Y17_VALUE_top2
  PIN Tile_X9Y17_VALUE_top3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1845.150 0.000 1845.430 4.000 ;
    END
  END Tile_X9Y17_VALUE_top3
  PIN Tile_X9Y17_VALUE_top4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1851.590 0.000 1851.870 4.000 ;
    END
  END Tile_X9Y17_VALUE_top4
  PIN Tile_X9Y17_VALUE_top5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1854.810 0.000 1855.090 4.000 ;
    END
  END Tile_X9Y17_VALUE_top5
  PIN Tile_X9Y17_VALUE_top6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1861.250 0.000 1861.530 4.000 ;
    END
  END Tile_X9Y17_VALUE_top6
  PIN Tile_X9Y17_VALUE_top7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1867.690 0.000 1867.970 4.000 ;
    END
  END Tile_X9Y17_VALUE_top7
  PIN Tile_X9Y17_VALUE_top8
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1874.130 0.000 1874.410 4.000 ;
    END
  END Tile_X9Y17_VALUE_top8
  PIN Tile_X9Y17_VALUE_top9
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1877.350 0.000 1877.630 4.000 ;
    END
  END Tile_X9Y17_VALUE_top9
  PIN UserCLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.998000 ;
    PORT
      LAYER met2 ;
        RECT 70.930 0.000 71.210 4.000 ;
    END
  END UserCLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 65.020 30.000 66.620 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 95.020 30.000 96.620 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 121.270 30.000 122.870 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 151.270 30.000 152.870 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 181.270 30.000 182.870 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 211.270 30.000 212.870 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 241.270 30.000 242.870 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 271.270 30.000 272.870 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 301.270 30.000 302.870 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 326.270 30.000 327.870 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 356.270 30.000 357.870 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 386.270 30.000 387.870 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 416.270 30.000 417.870 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 446.270 30.000 447.870 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 476.270 30.000 477.870 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 506.270 30.000 507.870 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 531.270 30.000 532.870 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 561.270 30.000 562.870 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 591.270 30.000 592.870 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 621.270 30.000 622.870 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 651.270 30.000 652.870 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 681.270 30.000 682.870 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 711.270 30.000 712.870 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 741.270 30.000 742.870 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 776.270 30.000 777.870 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 806.270 30.000 807.870 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 836.270 30.000 837.870 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 866.270 30.000 867.870 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 896.270 30.000 897.870 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 926.270 30.000 927.870 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 956.270 30.000 957.870 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 981.270 30.000 982.870 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1011.270 30.000 1012.870 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1041.270 30.000 1042.870 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1071.270 30.000 1072.870 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1101.270 30.000 1102.870 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1131.270 30.000 1132.870 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1161.270 30.000 1162.870 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1186.270 30.000 1187.870 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1216.270 30.000 1217.870 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1246.270 30.000 1247.870 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1276.270 30.000 1277.870 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1306.270 30.000 1307.870 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1336.270 30.000 1337.870 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1366.270 30.000 1367.870 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1391.270 30.000 1392.870 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1421.270 30.000 1422.870 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1451.270 30.000 1452.870 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1481.270 30.000 1482.870 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1511.270 30.000 1512.870 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1541.270 30.000 1542.870 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1571.270 30.000 1572.870 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1616.270 30.000 1617.870 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1646.270 30.000 1647.870 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1676.270 30.000 1677.870 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1706.270 30.000 1707.870 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1736.270 30.000 1737.870 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1766.270 30.000 1767.870 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1796.270 30.000 1797.870 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1821.270 30.000 1822.870 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1851.270 30.000 1852.870 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1881.270 30.000 1882.870 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1911.270 30.000 1912.870 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1941.270 30.000 1942.870 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1971.270 30.000 1972.870 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 2001.270 30.000 2002.870 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 2026.270 30.000 2027.870 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 2056.270 30.000 2057.870 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 2086.270 30.000 2087.870 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 2116.270 30.000 2117.870 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 2146.270 30.000 2147.870 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 2176.270 30.000 2177.870 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 2206.270 30.000 2207.870 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 2231.270 30.000 2232.870 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 2261.270 30.000 2262.870 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 2291.270 30.000 2292.870 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 2321.270 30.000 2322.870 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 2351.270 30.000 2352.870 3742.500 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 59.720 30.000 61.320 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 89.720 30.000 91.320 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 115.970 30.000 117.570 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 145.970 30.000 147.570 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 175.970 30.000 177.570 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 205.970 30.000 207.570 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 235.970 30.000 237.570 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 265.970 30.000 267.570 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 295.970 30.000 297.570 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 320.970 30.000 322.570 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 350.970 30.000 352.570 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 380.970 30.000 382.570 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 410.970 30.000 412.570 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 440.970 30.000 442.570 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 470.970 30.000 472.570 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 500.970 30.000 502.570 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 525.970 30.000 527.570 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 555.970 30.000 557.570 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 585.970 30.000 587.570 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 615.970 30.000 617.570 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 645.970 30.000 647.570 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 675.970 30.000 677.570 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 705.970 30.000 707.570 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 735.970 30.000 737.570 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 770.970 30.000 772.570 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 800.970 30.000 802.570 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 830.970 30.000 832.570 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 860.970 30.000 862.570 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 890.970 30.000 892.570 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 920.970 30.000 922.570 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 950.970 30.000 952.570 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 975.970 30.000 977.570 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1005.970 30.000 1007.570 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1035.970 30.000 1037.570 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1065.970 30.000 1067.570 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1095.970 30.000 1097.570 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1125.970 30.000 1127.570 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1155.970 30.000 1157.570 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1180.970 30.000 1182.570 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1210.970 30.000 1212.570 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1240.970 30.000 1242.570 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1270.970 30.000 1272.570 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1300.970 30.000 1302.570 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1330.970 30.000 1332.570 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1360.970 30.000 1362.570 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1385.970 30.000 1387.570 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1415.970 30.000 1417.570 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1445.970 30.000 1447.570 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1475.970 30.000 1477.570 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1505.970 30.000 1507.570 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1535.970 30.000 1537.570 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1565.970 30.000 1567.570 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1610.970 30.000 1612.570 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1640.970 30.000 1642.570 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1670.970 30.000 1672.570 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1700.970 30.000 1702.570 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1730.970 30.000 1732.570 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1760.970 30.000 1762.570 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1790.970 30.000 1792.570 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1815.970 30.000 1817.570 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1845.970 30.000 1847.570 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1875.970 30.000 1877.570 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1905.970 30.000 1907.570 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1935.970 30.000 1937.570 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1965.970 30.000 1967.570 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1995.970 30.000 1997.570 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 2020.970 30.000 2022.570 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 2050.970 30.000 2052.570 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 2080.970 30.000 2082.570 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 2110.970 30.000 2112.570 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 2140.970 30.000 2142.570 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 2170.970 30.000 2172.570 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 2200.970 30.000 2202.570 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 2225.970 30.000 2227.570 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 2255.970 30.000 2257.570 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 2285.970 30.000 2287.570 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 2315.970 30.000 2317.570 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 2345.970 30.000 2347.570 3742.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 2375.970 30.000 2377.570 3742.500 ;
    END
  END VPWR
  OBS
      LAYER nwell ;
        RECT 55.330 40.795 2379.280 3729.855 ;
      LAYER li1 ;
        RECT 55.520 40.795 2379.090 3729.855 ;
      LAYER met1 ;
        RECT 30.890 30.040 2414.930 3740.610 ;
      LAYER met2 ;
        RECT 1.010 3778.220 38.450 3779.285 ;
        RECT 39.290 3778.220 41.670 3779.285 ;
        RECT 42.510 3778.220 44.890 3779.285 ;
        RECT 45.730 3778.220 48.110 3779.285 ;
        RECT 48.950 3778.220 51.330 3779.285 ;
        RECT 52.170 3778.220 54.550 3779.285 ;
        RECT 55.390 3778.220 57.770 3779.285 ;
        RECT 58.610 3778.220 60.990 3779.285 ;
        RECT 61.830 3778.220 64.210 3779.285 ;
        RECT 65.050 3778.220 67.430 3779.285 ;
        RECT 68.270 3778.220 70.650 3779.285 ;
        RECT 71.490 3778.220 73.870 3779.285 ;
        RECT 74.710 3778.220 77.090 3779.285 ;
        RECT 77.930 3778.220 80.310 3779.285 ;
        RECT 81.150 3778.220 83.530 3779.285 ;
        RECT 84.370 3778.220 86.750 3779.285 ;
        RECT 87.590 3778.220 89.970 3779.285 ;
        RECT 90.810 3778.220 93.190 3779.285 ;
        RECT 94.030 3778.220 96.410 3779.285 ;
        RECT 97.250 3778.220 99.630 3779.285 ;
        RECT 100.470 3778.220 102.850 3779.285 ;
        RECT 103.690 3778.220 106.070 3779.285 ;
        RECT 106.910 3778.220 109.290 3779.285 ;
        RECT 110.130 3778.220 112.510 3779.285 ;
        RECT 113.350 3778.220 115.730 3779.285 ;
        RECT 116.570 3778.220 118.950 3779.285 ;
        RECT 119.790 3778.220 122.170 3779.285 ;
        RECT 123.010 3778.220 125.390 3779.285 ;
        RECT 126.230 3778.220 128.610 3779.285 ;
        RECT 129.450 3778.220 131.830 3779.285 ;
        RECT 132.670 3778.220 135.050 3779.285 ;
        RECT 135.890 3778.220 138.270 3779.285 ;
        RECT 139.110 3778.220 141.490 3779.285 ;
        RECT 142.330 3778.220 144.710 3779.285 ;
        RECT 145.550 3778.220 147.930 3779.285 ;
        RECT 148.770 3778.220 151.150 3779.285 ;
        RECT 151.990 3778.220 154.370 3779.285 ;
        RECT 155.210 3778.220 157.590 3779.285 ;
        RECT 158.430 3778.220 160.810 3779.285 ;
        RECT 161.650 3778.220 164.030 3779.285 ;
        RECT 164.870 3778.220 167.250 3779.285 ;
        RECT 168.090 3778.220 170.470 3779.285 ;
        RECT 171.310 3778.220 173.690 3779.285 ;
        RECT 174.530 3778.220 176.910 3779.285 ;
        RECT 177.750 3778.220 180.130 3779.285 ;
        RECT 180.970 3778.220 186.570 3779.285 ;
        RECT 187.410 3778.220 318.590 3779.285 ;
        RECT 319.430 3778.220 325.030 3779.285 ;
        RECT 325.870 3778.220 331.470 3779.285 ;
        RECT 332.310 3778.220 334.690 3779.285 ;
        RECT 335.530 3778.220 341.130 3779.285 ;
        RECT 341.970 3778.220 347.570 3779.285 ;
        RECT 348.410 3778.220 354.010 3779.285 ;
        RECT 354.850 3778.220 357.230 3779.285 ;
        RECT 358.070 3778.220 363.670 3779.285 ;
        RECT 364.510 3778.220 370.110 3779.285 ;
        RECT 370.950 3778.220 373.330 3779.285 ;
        RECT 374.170 3778.220 379.770 3779.285 ;
        RECT 380.610 3778.220 386.210 3779.285 ;
        RECT 387.050 3778.220 392.650 3779.285 ;
        RECT 393.490 3778.220 769.390 3779.285 ;
        RECT 770.230 3778.220 775.830 3779.285 ;
        RECT 776.670 3778.220 779.050 3779.285 ;
        RECT 779.890 3778.220 785.490 3779.285 ;
        RECT 786.330 3778.220 791.930 3779.285 ;
        RECT 792.770 3778.220 798.370 3779.285 ;
        RECT 799.210 3778.220 801.590 3779.285 ;
        RECT 802.430 3778.220 808.030 3779.285 ;
        RECT 808.870 3778.220 814.470 3779.285 ;
        RECT 815.310 3778.220 817.690 3779.285 ;
        RECT 818.530 3778.220 824.130 3779.285 ;
        RECT 824.970 3778.220 830.570 3779.285 ;
        RECT 831.410 3778.220 837.010 3779.285 ;
        RECT 837.850 3778.220 840.230 3779.285 ;
        RECT 841.070 3778.220 975.470 3779.285 ;
        RECT 976.310 3778.220 978.690 3779.285 ;
        RECT 979.530 3778.220 985.130 3779.285 ;
        RECT 985.970 3778.220 991.570 3779.285 ;
        RECT 992.410 3778.220 998.010 3779.285 ;
        RECT 998.850 3778.220 1001.230 3779.285 ;
        RECT 1002.070 3778.220 1007.670 3779.285 ;
        RECT 1008.510 3778.220 1014.110 3779.285 ;
        RECT 1014.950 3778.220 1017.330 3779.285 ;
        RECT 1018.170 3778.220 1023.770 3779.285 ;
        RECT 1024.610 3778.220 1030.210 3779.285 ;
        RECT 1031.050 3778.220 1036.650 3779.285 ;
        RECT 1037.490 3778.220 1039.870 3779.285 ;
        RECT 1040.710 3778.220 1046.310 3779.285 ;
        RECT 1047.150 3778.220 1178.330 3779.285 ;
        RECT 1179.170 3778.220 1184.770 3779.285 ;
        RECT 1185.610 3778.220 1191.210 3779.285 ;
        RECT 1192.050 3778.220 1194.430 3779.285 ;
        RECT 1195.270 3778.220 1200.870 3779.285 ;
        RECT 1201.710 3778.220 1207.310 3779.285 ;
        RECT 1208.150 3778.220 1213.750 3779.285 ;
        RECT 1214.590 3778.220 1216.970 3779.285 ;
        RECT 1217.810 3778.220 1223.410 3779.285 ;
        RECT 1224.250 3778.220 1229.850 3779.285 ;
        RECT 1230.690 3778.220 1233.070 3779.285 ;
        RECT 1233.910 3778.220 1239.510 3779.285 ;
        RECT 1240.350 3778.220 1245.950 3779.285 ;
        RECT 1246.790 3778.220 1252.390 3779.285 ;
        RECT 1253.230 3778.220 1609.810 3779.285 ;
        RECT 1610.650 3778.220 1616.250 3779.285 ;
        RECT 1617.090 3778.220 1619.470 3779.285 ;
        RECT 1620.310 3778.220 1625.910 3779.285 ;
        RECT 1626.750 3778.220 1632.350 3779.285 ;
        RECT 1633.190 3778.220 1635.570 3779.285 ;
        RECT 1636.410 3778.220 1642.010 3779.285 ;
        RECT 1642.850 3778.220 1648.450 3779.285 ;
        RECT 1649.290 3778.220 1654.890 3779.285 ;
        RECT 1655.730 3778.220 1658.110 3779.285 ;
        RECT 1658.950 3778.220 1664.550 3779.285 ;
        RECT 1665.390 3778.220 1670.990 3779.285 ;
        RECT 1671.830 3778.220 1674.210 3779.285 ;
        RECT 1675.050 3778.220 1680.650 3779.285 ;
        RECT 1681.490 3778.220 1815.890 3779.285 ;
        RECT 1816.730 3778.220 1819.110 3779.285 ;
        RECT 1819.950 3778.220 1825.550 3779.285 ;
        RECT 1826.390 3778.220 1831.990 3779.285 ;
        RECT 1832.830 3778.220 1835.210 3779.285 ;
        RECT 1836.050 3778.220 1841.650 3779.285 ;
        RECT 1842.490 3778.220 1848.090 3779.285 ;
        RECT 1848.930 3778.220 1854.530 3779.285 ;
        RECT 1855.370 3778.220 1857.750 3779.285 ;
        RECT 1858.590 3778.220 1864.190 3779.285 ;
        RECT 1865.030 3778.220 1870.630 3779.285 ;
        RECT 1871.470 3778.220 1873.850 3779.285 ;
        RECT 1874.690 3778.220 1880.290 3779.285 ;
        RECT 1881.130 3778.220 1886.730 3779.285 ;
        RECT 1887.570 3778.220 2018.750 3779.285 ;
        RECT 2019.590 3778.220 2025.190 3779.285 ;
        RECT 2026.030 3778.220 2031.630 3779.285 ;
        RECT 2032.470 3778.220 2034.850 3779.285 ;
        RECT 2035.690 3778.220 2041.290 3779.285 ;
        RECT 2042.130 3778.220 2047.730 3779.285 ;
        RECT 2048.570 3778.220 2050.950 3779.285 ;
        RECT 2051.790 3778.220 2057.390 3779.285 ;
        RECT 2058.230 3778.220 2063.830 3779.285 ;
        RECT 2064.670 3778.220 2070.270 3779.285 ;
        RECT 2071.110 3778.220 2073.490 3779.285 ;
        RECT 2074.330 3778.220 2079.930 3779.285 ;
        RECT 2080.770 3778.220 2086.370 3779.285 ;
        RECT 2087.210 3778.220 2089.590 3779.285 ;
        RECT 2090.430 3778.220 2432.390 3779.285 ;
        RECT 1.010 4.280 2432.390 3778.220 ;
        RECT 1.010 0.835 32.010 4.280 ;
        RECT 32.850 0.835 35.230 4.280 ;
        RECT 36.070 0.835 38.450 4.280 ;
        RECT 39.290 0.835 41.670 4.280 ;
        RECT 42.510 0.835 44.890 4.280 ;
        RECT 45.730 0.835 48.110 4.280 ;
        RECT 48.950 0.835 51.330 4.280 ;
        RECT 52.170 0.835 54.550 4.280 ;
        RECT 55.390 0.835 57.770 4.280 ;
        RECT 58.610 0.835 60.990 4.280 ;
        RECT 61.830 0.835 64.210 4.280 ;
        RECT 65.050 0.835 67.430 4.280 ;
        RECT 68.270 0.835 70.650 4.280 ;
        RECT 71.490 0.835 102.850 4.280 ;
        RECT 103.690 0.835 106.070 4.280 ;
        RECT 106.910 0.835 109.290 4.280 ;
        RECT 110.130 0.835 112.510 4.280 ;
        RECT 113.350 0.835 115.730 4.280 ;
        RECT 116.570 0.835 122.170 4.280 ;
        RECT 123.010 0.835 128.610 4.280 ;
        RECT 129.450 0.835 138.270 4.280 ;
        RECT 139.110 0.835 154.370 4.280 ;
        RECT 155.210 0.835 160.810 4.280 ;
        RECT 161.650 0.835 170.470 4.280 ;
        RECT 171.310 0.835 176.910 4.280 ;
        RECT 177.750 0.835 183.350 4.280 ;
        RECT 184.190 0.835 193.010 4.280 ;
        RECT 193.850 0.835 199.450 4.280 ;
        RECT 200.290 0.835 209.110 4.280 ;
        RECT 209.950 0.835 215.550 4.280 ;
        RECT 216.390 0.835 225.210 4.280 ;
        RECT 226.050 0.835 231.650 4.280 ;
        RECT 232.490 0.835 238.090 4.280 ;
        RECT 238.930 0.835 247.750 4.280 ;
        RECT 248.590 0.835 254.190 4.280 ;
        RECT 255.030 0.835 263.850 4.280 ;
        RECT 264.690 0.835 270.290 4.280 ;
        RECT 271.130 0.835 279.950 4.280 ;
        RECT 280.790 0.835 286.390 4.280 ;
        RECT 287.230 0.835 292.830 4.280 ;
        RECT 293.670 0.835 302.490 4.280 ;
        RECT 303.330 0.835 318.590 4.280 ;
        RECT 319.430 0.835 325.030 4.280 ;
        RECT 325.870 0.835 331.470 4.280 ;
        RECT 332.310 0.835 341.130 4.280 ;
        RECT 341.970 0.835 347.570 4.280 ;
        RECT 348.410 0.835 354.010 4.280 ;
        RECT 354.850 0.835 370.110 4.280 ;
        RECT 370.950 0.835 376.550 4.280 ;
        RECT 377.390 0.835 382.990 4.280 ;
        RECT 383.830 0.835 392.650 4.280 ;
        RECT 393.490 0.835 399.090 4.280 ;
        RECT 399.930 0.835 405.530 4.280 ;
        RECT 406.370 0.835 411.970 4.280 ;
        RECT 412.810 0.835 421.630 4.280 ;
        RECT 422.470 0.835 428.070 4.280 ;
        RECT 428.910 0.835 434.510 4.280 ;
        RECT 435.350 0.835 444.170 4.280 ;
        RECT 445.010 0.835 450.610 4.280 ;
        RECT 451.450 0.835 457.050 4.280 ;
        RECT 457.890 0.835 463.490 4.280 ;
        RECT 464.330 0.835 473.150 4.280 ;
        RECT 473.990 0.835 479.590 4.280 ;
        RECT 480.430 0.835 486.030 4.280 ;
        RECT 486.870 0.835 495.690 4.280 ;
        RECT 496.530 0.835 502.130 4.280 ;
        RECT 502.970 0.835 508.570 4.280 ;
        RECT 509.410 0.835 534.330 4.280 ;
        RECT 535.170 0.835 547.210 4.280 ;
        RECT 548.050 0.835 556.870 4.280 ;
        RECT 557.710 0.835 569.750 4.280 ;
        RECT 570.590 0.835 579.410 4.280 ;
        RECT 580.250 0.835 592.290 4.280 ;
        RECT 593.130 0.835 601.950 4.280 ;
        RECT 602.790 0.835 614.830 4.280 ;
        RECT 615.670 0.835 627.710 4.280 ;
        RECT 628.550 0.835 637.370 4.280 ;
        RECT 638.210 0.835 650.250 4.280 ;
        RECT 651.090 0.835 659.910 4.280 ;
        RECT 660.750 0.835 672.790 4.280 ;
        RECT 673.630 0.835 682.450 4.280 ;
        RECT 683.290 0.835 695.330 4.280 ;
        RECT 696.170 0.835 708.210 4.280 ;
        RECT 709.050 0.835 717.870 4.280 ;
        RECT 718.710 0.835 730.750 4.280 ;
        RECT 731.590 0.835 740.410 4.280 ;
        RECT 741.250 0.835 753.290 4.280 ;
        RECT 754.130 0.835 766.170 4.280 ;
        RECT 767.010 0.835 772.610 4.280 ;
        RECT 773.450 0.835 775.830 4.280 ;
        RECT 776.670 0.835 779.050 4.280 ;
        RECT 779.890 0.835 782.270 4.280 ;
        RECT 783.110 0.835 785.490 4.280 ;
        RECT 786.330 0.835 788.710 4.280 ;
        RECT 789.550 0.835 791.930 4.280 ;
        RECT 792.770 0.835 798.370 4.280 ;
        RECT 799.210 0.835 801.590 4.280 ;
        RECT 802.430 0.835 804.810 4.280 ;
        RECT 805.650 0.835 808.030 4.280 ;
        RECT 808.870 0.835 811.250 4.280 ;
        RECT 812.090 0.835 814.470 4.280 ;
        RECT 815.310 0.835 817.690 4.280 ;
        RECT 818.530 0.835 824.130 4.280 ;
        RECT 824.970 0.835 827.350 4.280 ;
        RECT 828.190 0.835 830.570 4.280 ;
        RECT 831.410 0.835 833.790 4.280 ;
        RECT 834.630 0.835 837.010 4.280 ;
        RECT 837.850 0.835 840.230 4.280 ;
        RECT 841.070 0.835 843.450 4.280 ;
        RECT 844.290 0.835 849.890 4.280 ;
        RECT 850.730 0.835 853.110 4.280 ;
        RECT 853.950 0.835 856.330 4.280 ;
        RECT 857.170 0.835 859.550 4.280 ;
        RECT 860.390 0.835 862.770 4.280 ;
        RECT 863.610 0.835 865.990 4.280 ;
        RECT 866.830 0.835 869.210 4.280 ;
        RECT 870.050 0.835 875.650 4.280 ;
        RECT 876.490 0.835 878.870 4.280 ;
        RECT 879.710 0.835 882.090 4.280 ;
        RECT 882.930 0.835 888.530 4.280 ;
        RECT 889.370 0.835 891.750 4.280 ;
        RECT 892.590 0.835 894.970 4.280 ;
        RECT 895.810 0.835 901.410 4.280 ;
        RECT 902.250 0.835 904.630 4.280 ;
        RECT 905.470 0.835 907.850 4.280 ;
        RECT 908.690 0.835 911.070 4.280 ;
        RECT 911.910 0.835 914.290 4.280 ;
        RECT 915.130 0.835 917.510 4.280 ;
        RECT 918.350 0.835 920.730 4.280 ;
        RECT 921.570 0.835 927.170 4.280 ;
        RECT 928.010 0.835 930.390 4.280 ;
        RECT 931.230 0.835 933.610 4.280 ;
        RECT 934.450 0.835 936.830 4.280 ;
        RECT 937.670 0.835 940.050 4.280 ;
        RECT 940.890 0.835 943.270 4.280 ;
        RECT 944.110 0.835 946.490 4.280 ;
        RECT 947.330 0.835 952.930 4.280 ;
        RECT 953.770 0.835 956.150 4.280 ;
        RECT 956.990 0.835 959.370 4.280 ;
        RECT 960.210 0.835 972.250 4.280 ;
        RECT 973.090 0.835 975.470 4.280 ;
        RECT 976.310 0.835 978.690 4.280 ;
        RECT 979.530 0.835 985.130 4.280 ;
        RECT 985.970 0.835 988.350 4.280 ;
        RECT 989.190 0.835 991.570 4.280 ;
        RECT 992.410 0.835 994.790 4.280 ;
        RECT 995.630 0.835 998.010 4.280 ;
        RECT 998.850 0.835 1001.230 4.280 ;
        RECT 1002.070 0.835 1004.450 4.280 ;
        RECT 1005.290 0.835 1010.890 4.280 ;
        RECT 1011.730 0.835 1014.110 4.280 ;
        RECT 1014.950 0.835 1017.330 4.280 ;
        RECT 1018.170 0.835 1020.550 4.280 ;
        RECT 1021.390 0.835 1023.770 4.280 ;
        RECT 1024.610 0.835 1026.990 4.280 ;
        RECT 1027.830 0.835 1030.210 4.280 ;
        RECT 1031.050 0.835 1036.650 4.280 ;
        RECT 1037.490 0.835 1039.870 4.280 ;
        RECT 1040.710 0.835 1043.090 4.280 ;
        RECT 1043.930 0.835 1046.310 4.280 ;
        RECT 1047.150 0.835 1049.530 4.280 ;
        RECT 1050.370 0.835 1052.750 4.280 ;
        RECT 1053.590 0.835 1055.970 4.280 ;
        RECT 1056.810 0.835 1062.410 4.280 ;
        RECT 1063.250 0.835 1065.630 4.280 ;
        RECT 1066.470 0.835 1068.850 4.280 ;
        RECT 1069.690 0.835 1072.070 4.280 ;
        RECT 1072.910 0.835 1075.290 4.280 ;
        RECT 1076.130 0.835 1078.510 4.280 ;
        RECT 1079.350 0.835 1081.730 4.280 ;
        RECT 1082.570 0.835 1088.170 4.280 ;
        RECT 1089.010 0.835 1094.610 4.280 ;
        RECT 1095.450 0.835 1097.830 4.280 ;
        RECT 1098.670 0.835 1101.050 4.280 ;
        RECT 1101.890 0.835 1104.270 4.280 ;
        RECT 1105.110 0.835 1107.490 4.280 ;
        RECT 1108.330 0.835 1113.930 4.280 ;
        RECT 1114.770 0.835 1117.150 4.280 ;
        RECT 1117.990 0.835 1120.370 4.280 ;
        RECT 1121.210 0.835 1123.590 4.280 ;
        RECT 1124.430 0.835 1126.810 4.280 ;
        RECT 1127.650 0.835 1130.030 4.280 ;
        RECT 1130.870 0.835 1133.250 4.280 ;
        RECT 1134.090 0.835 1139.690 4.280 ;
        RECT 1140.530 0.835 1142.910 4.280 ;
        RECT 1143.750 0.835 1146.130 4.280 ;
        RECT 1146.970 0.835 1149.350 4.280 ;
        RECT 1150.190 0.835 1152.570 4.280 ;
        RECT 1153.410 0.835 1155.790 4.280 ;
        RECT 1156.630 0.835 1159.010 4.280 ;
        RECT 1159.850 0.835 1165.450 4.280 ;
        RECT 1166.290 0.835 1178.330 4.280 ;
        RECT 1179.170 0.835 1181.550 4.280 ;
        RECT 1182.390 0.835 1184.770 4.280 ;
        RECT 1185.610 0.835 1187.990 4.280 ;
        RECT 1188.830 0.835 1191.210 4.280 ;
        RECT 1192.050 0.835 1194.430 4.280 ;
        RECT 1195.270 0.835 1200.870 4.280 ;
        RECT 1201.710 0.835 1204.090 4.280 ;
        RECT 1204.930 0.835 1207.310 4.280 ;
        RECT 1208.150 0.835 1210.530 4.280 ;
        RECT 1211.370 0.835 1213.750 4.280 ;
        RECT 1214.590 0.835 1216.970 4.280 ;
        RECT 1217.810 0.835 1220.190 4.280 ;
        RECT 1221.030 0.835 1226.630 4.280 ;
        RECT 1227.470 0.835 1229.850 4.280 ;
        RECT 1230.690 0.835 1233.070 4.280 ;
        RECT 1233.910 0.835 1236.290 4.280 ;
        RECT 1237.130 0.835 1239.510 4.280 ;
        RECT 1240.350 0.835 1242.730 4.280 ;
        RECT 1243.570 0.835 1245.950 4.280 ;
        RECT 1246.790 0.835 1252.390 4.280 ;
        RECT 1253.230 0.835 1255.610 4.280 ;
        RECT 1256.450 0.835 1258.830 4.280 ;
        RECT 1259.670 0.835 1262.050 4.280 ;
        RECT 1262.890 0.835 1265.270 4.280 ;
        RECT 1266.110 0.835 1268.490 4.280 ;
        RECT 1269.330 0.835 1271.710 4.280 ;
        RECT 1272.550 0.835 1278.150 4.280 ;
        RECT 1278.990 0.835 1281.370 4.280 ;
        RECT 1282.210 0.835 1284.590 4.280 ;
        RECT 1285.430 0.835 1287.810 4.280 ;
        RECT 1288.650 0.835 1291.030 4.280 ;
        RECT 1291.870 0.835 1297.470 4.280 ;
        RECT 1298.310 0.835 1303.910 4.280 ;
        RECT 1304.750 0.835 1307.130 4.280 ;
        RECT 1307.970 0.835 1310.350 4.280 ;
        RECT 1311.190 0.835 1313.570 4.280 ;
        RECT 1314.410 0.835 1316.790 4.280 ;
        RECT 1317.630 0.835 1320.010 4.280 ;
        RECT 1320.850 0.835 1323.230 4.280 ;
        RECT 1324.070 0.835 1329.670 4.280 ;
        RECT 1330.510 0.835 1332.890 4.280 ;
        RECT 1333.730 0.835 1336.110 4.280 ;
        RECT 1336.950 0.835 1339.330 4.280 ;
        RECT 1340.170 0.835 1342.550 4.280 ;
        RECT 1343.390 0.835 1345.770 4.280 ;
        RECT 1346.610 0.835 1348.990 4.280 ;
        RECT 1349.830 0.835 1355.430 4.280 ;
        RECT 1356.270 0.835 1358.650 4.280 ;
        RECT 1359.490 0.835 1361.870 4.280 ;
        RECT 1362.710 0.835 1365.090 4.280 ;
        RECT 1365.930 0.835 1368.310 4.280 ;
        RECT 1369.150 0.835 1394.070 4.280 ;
        RECT 1394.910 0.835 1403.730 4.280 ;
        RECT 1404.570 0.835 1413.390 4.280 ;
        RECT 1414.230 0.835 1426.270 4.280 ;
        RECT 1427.110 0.835 1435.930 4.280 ;
        RECT 1436.770 0.835 1445.590 4.280 ;
        RECT 1446.430 0.835 1455.250 4.280 ;
        RECT 1456.090 0.835 1468.130 4.280 ;
        RECT 1468.970 0.835 1477.790 4.280 ;
        RECT 1478.630 0.835 1487.450 4.280 ;
        RECT 1488.290 0.835 1500.330 4.280 ;
        RECT 1501.170 0.835 1509.990 4.280 ;
        RECT 1510.830 0.835 1519.650 4.280 ;
        RECT 1520.490 0.835 1529.310 4.280 ;
        RECT 1530.150 0.835 1542.190 4.280 ;
        RECT 1543.030 0.835 1551.850 4.280 ;
        RECT 1552.690 0.835 1561.510 4.280 ;
        RECT 1562.350 0.835 1574.390 4.280 ;
        RECT 1575.230 0.835 1584.050 4.280 ;
        RECT 1584.890 0.835 1593.710 4.280 ;
        RECT 1594.550 0.835 1606.590 4.280 ;
        RECT 1607.430 0.835 1609.810 4.280 ;
        RECT 1610.650 0.835 1616.250 4.280 ;
        RECT 1617.090 0.835 1619.470 4.280 ;
        RECT 1620.310 0.835 1622.690 4.280 ;
        RECT 1623.530 0.835 1625.910 4.280 ;
        RECT 1626.750 0.835 1629.130 4.280 ;
        RECT 1629.970 0.835 1632.350 4.280 ;
        RECT 1633.190 0.835 1635.570 4.280 ;
        RECT 1636.410 0.835 1642.010 4.280 ;
        RECT 1642.850 0.835 1645.230 4.280 ;
        RECT 1646.070 0.835 1648.450 4.280 ;
        RECT 1649.290 0.835 1651.670 4.280 ;
        RECT 1652.510 0.835 1654.890 4.280 ;
        RECT 1655.730 0.835 1658.110 4.280 ;
        RECT 1658.950 0.835 1661.330 4.280 ;
        RECT 1662.170 0.835 1667.770 4.280 ;
        RECT 1668.610 0.835 1670.990 4.280 ;
        RECT 1671.830 0.835 1674.210 4.280 ;
        RECT 1675.050 0.835 1677.430 4.280 ;
        RECT 1678.270 0.835 1680.650 4.280 ;
        RECT 1681.490 0.835 1683.870 4.280 ;
        RECT 1684.710 0.835 1687.090 4.280 ;
        RECT 1687.930 0.835 1693.530 4.280 ;
        RECT 1694.370 0.835 1696.750 4.280 ;
        RECT 1697.590 0.835 1699.970 4.280 ;
        RECT 1700.810 0.835 1703.190 4.280 ;
        RECT 1704.030 0.835 1706.410 4.280 ;
        RECT 1707.250 0.835 1709.630 4.280 ;
        RECT 1710.470 0.835 1712.850 4.280 ;
        RECT 1713.690 0.835 1719.290 4.280 ;
        RECT 1720.130 0.835 1722.510 4.280 ;
        RECT 1723.350 0.835 1728.950 4.280 ;
        RECT 1729.790 0.835 1732.170 4.280 ;
        RECT 1733.010 0.835 1735.390 4.280 ;
        RECT 1736.230 0.835 1738.610 4.280 ;
        RECT 1739.450 0.835 1745.050 4.280 ;
        RECT 1745.890 0.835 1748.270 4.280 ;
        RECT 1749.110 0.835 1751.490 4.280 ;
        RECT 1752.330 0.835 1754.710 4.280 ;
        RECT 1755.550 0.835 1757.930 4.280 ;
        RECT 1758.770 0.835 1761.150 4.280 ;
        RECT 1761.990 0.835 1764.370 4.280 ;
        RECT 1765.210 0.835 1770.810 4.280 ;
        RECT 1771.650 0.835 1774.030 4.280 ;
        RECT 1774.870 0.835 1777.250 4.280 ;
        RECT 1778.090 0.835 1780.470 4.280 ;
        RECT 1781.310 0.835 1783.690 4.280 ;
        RECT 1784.530 0.835 1786.910 4.280 ;
        RECT 1787.750 0.835 1790.130 4.280 ;
        RECT 1790.970 0.835 1796.570 4.280 ;
        RECT 1797.410 0.835 1799.790 4.280 ;
        RECT 1800.630 0.835 1812.670 4.280 ;
        RECT 1813.510 0.835 1815.890 4.280 ;
        RECT 1816.730 0.835 1822.330 4.280 ;
        RECT 1823.170 0.835 1828.770 4.280 ;
        RECT 1829.610 0.835 1835.210 4.280 ;
        RECT 1836.050 0.835 1838.430 4.280 ;
        RECT 1839.270 0.835 1844.870 4.280 ;
        RECT 1845.710 0.835 1851.310 4.280 ;
        RECT 1852.150 0.835 1854.530 4.280 ;
        RECT 1855.370 0.835 1860.970 4.280 ;
        RECT 1861.810 0.835 1867.410 4.280 ;
        RECT 1868.250 0.835 1873.850 4.280 ;
        RECT 1874.690 0.835 1877.070 4.280 ;
        RECT 1877.910 0.835 1883.510 4.280 ;
        RECT 1884.350 0.835 1889.950 4.280 ;
        RECT 1890.790 0.835 1931.810 4.280 ;
        RECT 1932.650 0.835 1935.030 4.280 ;
        RECT 1935.870 0.835 1938.250 4.280 ;
        RECT 1939.090 0.835 1941.470 4.280 ;
        RECT 1942.310 0.835 1944.690 4.280 ;
        RECT 1945.530 0.835 1947.910 4.280 ;
        RECT 1948.750 0.835 1951.130 4.280 ;
        RECT 1951.970 0.835 1954.350 4.280 ;
        RECT 1955.190 0.835 1957.570 4.280 ;
        RECT 1958.410 0.835 1960.790 4.280 ;
        RECT 1961.630 0.835 1964.010 4.280 ;
        RECT 1964.850 0.835 1967.230 4.280 ;
        RECT 1968.070 0.835 1970.450 4.280 ;
        RECT 1971.290 0.835 1973.670 4.280 ;
        RECT 1974.510 0.835 1976.890 4.280 ;
        RECT 1977.730 0.835 1983.330 4.280 ;
        RECT 1984.170 0.835 1989.770 4.280 ;
        RECT 1990.610 0.835 1992.990 4.280 ;
        RECT 1993.830 0.835 1999.430 4.280 ;
        RECT 2000.270 0.835 2005.870 4.280 ;
        RECT 2006.710 0.835 2015.530 4.280 ;
        RECT 2016.370 0.835 2021.970 4.280 ;
        RECT 2022.810 0.835 2031.630 4.280 ;
        RECT 2032.470 0.835 2038.070 4.280 ;
        RECT 2038.910 0.835 2044.510 4.280 ;
        RECT 2045.350 0.835 2050.950 4.280 ;
        RECT 2051.790 0.835 2057.390 4.280 ;
        RECT 2058.230 0.835 2063.830 4.280 ;
        RECT 2064.670 0.835 2079.930 4.280 ;
        RECT 2080.770 0.835 2086.370 4.280 ;
        RECT 2087.210 0.835 2092.810 4.280 ;
        RECT 2093.650 0.835 2099.250 4.280 ;
        RECT 2100.090 0.835 2105.690 4.280 ;
        RECT 2106.530 0.835 2112.130 4.280 ;
        RECT 2112.970 0.835 2118.570 4.280 ;
        RECT 2119.410 0.835 2128.230 4.280 ;
        RECT 2129.070 0.835 2134.670 4.280 ;
        RECT 2135.510 0.835 2141.110 4.280 ;
        RECT 2141.950 0.835 2147.550 4.280 ;
        RECT 2148.390 0.835 2153.990 4.280 ;
        RECT 2154.830 0.835 2160.430 4.280 ;
        RECT 2161.270 0.835 2166.870 4.280 ;
        RECT 2167.710 0.835 2176.530 4.280 ;
        RECT 2177.370 0.835 2182.970 4.280 ;
        RECT 2183.810 0.835 2189.410 4.280 ;
        RECT 2190.250 0.835 2195.850 4.280 ;
        RECT 2196.690 0.835 2202.290 4.280 ;
        RECT 2203.130 0.835 2208.730 4.280 ;
        RECT 2209.570 0.835 2231.270 4.280 ;
        RECT 2232.110 0.835 2237.710 4.280 ;
        RECT 2238.550 0.835 2244.150 4.280 ;
        RECT 2244.990 0.835 2253.810 4.280 ;
        RECT 2254.650 0.835 2260.250 4.280 ;
        RECT 2261.090 0.835 2269.910 4.280 ;
        RECT 2270.750 0.835 2276.350 4.280 ;
        RECT 2277.190 0.835 2286.010 4.280 ;
        RECT 2286.850 0.835 2292.450 4.280 ;
        RECT 2293.290 0.835 2298.890 4.280 ;
        RECT 2299.730 0.835 2308.550 4.280 ;
        RECT 2309.390 0.835 2314.990 4.280 ;
        RECT 2315.830 0.835 2324.650 4.280 ;
        RECT 2325.490 0.835 2331.090 4.280 ;
        RECT 2331.930 0.835 2340.750 4.280 ;
        RECT 2341.590 0.835 2347.190 4.280 ;
        RECT 2348.030 0.835 2353.630 4.280 ;
        RECT 2354.470 0.835 2363.290 4.280 ;
        RECT 2364.130 0.835 2369.730 4.280 ;
        RECT 2370.570 0.835 2379.390 4.280 ;
        RECT 2380.230 0.835 2432.390 4.280 ;
      LAYER met3 ;
        RECT 0.270 3768.240 2432.415 3779.265 ;
        RECT 0.270 3766.840 2430.600 3768.240 ;
        RECT 0.270 3764.840 2432.415 3766.840 ;
        RECT 0.270 3763.440 2430.600 3764.840 ;
        RECT 0.270 3761.440 2432.415 3763.440 ;
        RECT 0.270 3760.040 2430.600 3761.440 ;
        RECT 0.270 3758.040 2432.415 3760.040 ;
        RECT 0.270 3756.640 2430.600 3758.040 ;
        RECT 0.270 3754.640 2432.415 3756.640 ;
        RECT 0.270 3753.240 2430.600 3754.640 ;
        RECT 0.270 3751.240 2432.415 3753.240 ;
        RECT 0.270 3749.840 2430.600 3751.240 ;
        RECT 0.270 3747.840 2432.415 3749.840 ;
        RECT 0.270 3746.440 2430.600 3747.840 ;
        RECT 0.270 3744.440 2432.415 3746.440 ;
        RECT 0.270 3743.040 2430.600 3744.440 ;
        RECT 0.270 3741.040 2432.415 3743.040 ;
        RECT 0.270 3739.640 2430.600 3741.040 ;
        RECT 0.270 3737.640 2432.415 3739.640 ;
        RECT 0.270 3736.240 2430.600 3737.640 ;
        RECT 0.270 3734.240 2432.415 3736.240 ;
        RECT 0.270 3732.840 2430.600 3734.240 ;
        RECT 0.270 3730.840 2432.415 3732.840 ;
        RECT 0.270 3729.440 2430.600 3730.840 ;
        RECT 0.270 3727.440 2432.415 3729.440 ;
        RECT 0.270 3726.040 2430.600 3727.440 ;
        RECT 0.270 3724.040 2432.415 3726.040 ;
        RECT 0.270 3722.640 2430.600 3724.040 ;
        RECT 0.270 3720.640 2432.415 3722.640 ;
        RECT 0.270 3719.240 2430.600 3720.640 ;
        RECT 0.270 3717.240 2432.415 3719.240 ;
        RECT 0.270 3715.840 2430.600 3717.240 ;
        RECT 0.270 3713.840 2432.415 3715.840 ;
        RECT 0.270 3712.440 2430.600 3713.840 ;
        RECT 0.270 3710.440 2432.415 3712.440 ;
        RECT 0.270 3709.040 2430.600 3710.440 ;
        RECT 0.270 3707.040 2432.415 3709.040 ;
        RECT 0.270 3705.640 2430.600 3707.040 ;
        RECT 0.270 3703.640 2432.415 3705.640 ;
        RECT 0.270 3702.240 2430.600 3703.640 ;
        RECT 0.270 3700.240 2432.415 3702.240 ;
        RECT 0.270 3698.840 2430.600 3700.240 ;
        RECT 0.270 3696.840 2432.415 3698.840 ;
        RECT 0.270 3695.440 2430.600 3696.840 ;
        RECT 0.270 3693.440 2432.415 3695.440 ;
        RECT 0.270 3692.040 2430.600 3693.440 ;
        RECT 0.270 3690.040 2432.415 3692.040 ;
        RECT 0.270 3688.640 2430.600 3690.040 ;
        RECT 0.270 3686.640 2432.415 3688.640 ;
        RECT 0.270 3685.240 2430.600 3686.640 ;
        RECT 0.270 3683.240 2432.415 3685.240 ;
        RECT 0.270 3681.840 2430.600 3683.240 ;
        RECT 0.270 3679.840 2432.415 3681.840 ;
        RECT 0.270 3678.440 2430.600 3679.840 ;
        RECT 0.270 3676.440 2432.415 3678.440 ;
        RECT 0.270 3675.040 2430.600 3676.440 ;
        RECT 0.270 3673.040 2432.415 3675.040 ;
        RECT 0.270 3671.640 2430.600 3673.040 ;
        RECT 0.270 3669.640 2432.415 3671.640 ;
        RECT 0.270 3668.240 2430.600 3669.640 ;
        RECT 0.270 3666.240 2432.415 3668.240 ;
        RECT 4.400 3664.840 2430.600 3666.240 ;
        RECT 0.270 3662.840 2432.415 3664.840 ;
        RECT 4.400 3661.440 2430.600 3662.840 ;
        RECT 0.270 3659.440 2432.415 3661.440 ;
        RECT 4.400 3658.040 2430.600 3659.440 ;
        RECT 0.270 3656.040 2432.415 3658.040 ;
        RECT 0.270 3654.640 2430.600 3656.040 ;
        RECT 0.270 3652.640 2432.415 3654.640 ;
        RECT 4.400 3651.240 2430.600 3652.640 ;
        RECT 0.270 3649.240 2432.415 3651.240 ;
        RECT 4.400 3647.840 2430.600 3649.240 ;
        RECT 0.270 3645.840 2432.415 3647.840 ;
        RECT 4.400 3644.440 2430.600 3645.840 ;
        RECT 0.270 3642.440 2432.415 3644.440 ;
        RECT 4.400 3641.040 2430.600 3642.440 ;
        RECT 0.270 3639.040 2432.415 3641.040 ;
        RECT 4.400 3637.640 2430.600 3639.040 ;
        RECT 0.270 3635.640 2432.415 3637.640 ;
        RECT 0.270 3634.240 2430.600 3635.640 ;
        RECT 0.270 3632.240 2432.415 3634.240 ;
        RECT 4.400 3630.840 2430.600 3632.240 ;
        RECT 0.270 3628.840 2432.415 3630.840 ;
        RECT 4.400 3627.440 2430.600 3628.840 ;
        RECT 0.270 3625.440 2432.415 3627.440 ;
        RECT 4.400 3624.040 2430.600 3625.440 ;
        RECT 0.270 3622.040 2432.415 3624.040 ;
        RECT 4.400 3620.640 2430.600 3622.040 ;
        RECT 0.270 3618.640 2432.415 3620.640 ;
        RECT 4.400 3617.240 2430.600 3618.640 ;
        RECT 0.270 3615.240 2432.415 3617.240 ;
        RECT 0.270 3613.840 2430.600 3615.240 ;
        RECT 0.270 3611.840 2432.415 3613.840 ;
        RECT 4.400 3610.440 2430.600 3611.840 ;
        RECT 0.270 3608.440 2432.415 3610.440 ;
        RECT 4.400 3607.040 2430.600 3608.440 ;
        RECT 0.270 3605.040 2432.415 3607.040 ;
        RECT 4.400 3603.640 2430.600 3605.040 ;
        RECT 0.270 3601.640 2432.415 3603.640 ;
        RECT 4.400 3600.240 2430.600 3601.640 ;
        RECT 0.270 3598.240 2432.415 3600.240 ;
        RECT 4.400 3596.840 2430.600 3598.240 ;
        RECT 0.270 3594.840 2432.415 3596.840 ;
        RECT 0.270 3593.440 2430.600 3594.840 ;
        RECT 0.270 3591.440 2432.415 3593.440 ;
        RECT 4.400 3590.040 2430.600 3591.440 ;
        RECT 0.270 3588.040 2432.415 3590.040 ;
        RECT 4.400 3586.640 2430.600 3588.040 ;
        RECT 0.270 3584.640 2432.415 3586.640 ;
        RECT 4.400 3583.240 2430.600 3584.640 ;
        RECT 0.270 3581.240 2432.415 3583.240 ;
        RECT 4.400 3579.840 2430.600 3581.240 ;
        RECT 0.270 3577.840 2432.415 3579.840 ;
        RECT 4.400 3576.440 2430.600 3577.840 ;
        RECT 0.270 3574.440 2432.415 3576.440 ;
        RECT 0.270 3573.040 2430.600 3574.440 ;
        RECT 0.270 3571.040 2432.415 3573.040 ;
        RECT 4.400 3569.640 2430.600 3571.040 ;
        RECT 0.270 3567.640 2432.415 3569.640 ;
        RECT 4.400 3566.240 2430.600 3567.640 ;
        RECT 0.270 3564.240 2432.415 3566.240 ;
        RECT 4.400 3562.840 2430.600 3564.240 ;
        RECT 0.270 3560.840 2432.415 3562.840 ;
        RECT 4.400 3559.440 2430.600 3560.840 ;
        RECT 0.270 3557.440 2432.415 3559.440 ;
        RECT 4.400 3556.040 2430.600 3557.440 ;
        RECT 0.270 3554.040 2432.415 3556.040 ;
        RECT 0.270 3552.640 2430.600 3554.040 ;
        RECT 0.270 3550.640 2432.415 3552.640 ;
        RECT 4.400 3549.240 2430.600 3550.640 ;
        RECT 0.270 3547.240 2432.415 3549.240 ;
        RECT 4.400 3545.840 2430.600 3547.240 ;
        RECT 0.270 3543.840 2432.415 3545.840 ;
        RECT 4.400 3542.440 2430.600 3543.840 ;
        RECT 0.270 3540.440 2432.415 3542.440 ;
        RECT 4.400 3539.040 2430.600 3540.440 ;
        RECT 0.270 3537.040 2432.415 3539.040 ;
        RECT 4.400 3535.640 2430.600 3537.040 ;
        RECT 0.270 3533.640 2432.415 3535.640 ;
        RECT 0.270 3532.240 2430.600 3533.640 ;
        RECT 0.270 3530.240 2432.415 3532.240 ;
        RECT 4.400 3528.840 2430.600 3530.240 ;
        RECT 0.270 3526.840 2432.415 3528.840 ;
        RECT 4.400 3525.440 2430.600 3526.840 ;
        RECT 0.270 3523.440 2432.415 3525.440 ;
        RECT 4.400 3522.040 2430.600 3523.440 ;
        RECT 0.270 3520.040 2432.415 3522.040 ;
        RECT 4.400 3518.640 2430.600 3520.040 ;
        RECT 0.270 3516.640 2432.415 3518.640 ;
        RECT 4.400 3515.240 2430.600 3516.640 ;
        RECT 0.270 3513.240 2432.415 3515.240 ;
        RECT 0.270 3511.840 2430.600 3513.240 ;
        RECT 0.270 3509.840 2432.415 3511.840 ;
        RECT 4.400 3508.440 2430.600 3509.840 ;
        RECT 0.270 3506.440 2432.415 3508.440 ;
        RECT 4.400 3505.040 2430.600 3506.440 ;
        RECT 0.270 3503.040 2432.415 3505.040 ;
        RECT 4.400 3501.640 2430.600 3503.040 ;
        RECT 0.270 3499.640 2432.415 3501.640 ;
        RECT 4.400 3498.240 2430.600 3499.640 ;
        RECT 0.270 3496.240 2432.415 3498.240 ;
        RECT 4.400 3494.840 2430.600 3496.240 ;
        RECT 0.270 3492.840 2432.415 3494.840 ;
        RECT 0.270 3491.440 2430.600 3492.840 ;
        RECT 0.270 3489.440 2432.415 3491.440 ;
        RECT 4.400 3488.040 2430.600 3489.440 ;
        RECT 0.270 3486.040 2432.415 3488.040 ;
        RECT 4.400 3484.640 2430.600 3486.040 ;
        RECT 0.270 3482.640 2432.415 3484.640 ;
        RECT 4.400 3481.240 2430.600 3482.640 ;
        RECT 0.270 3479.240 2432.415 3481.240 ;
        RECT 0.270 3477.840 2430.600 3479.240 ;
        RECT 0.270 3475.840 2432.415 3477.840 ;
        RECT 0.270 3474.440 2430.600 3475.840 ;
        RECT 0.270 3472.440 2432.415 3474.440 ;
        RECT 0.270 3471.040 2430.600 3472.440 ;
        RECT 0.270 3469.040 2432.415 3471.040 ;
        RECT 0.270 3467.640 2430.600 3469.040 ;
        RECT 0.270 3465.640 2432.415 3467.640 ;
        RECT 0.270 3464.240 2430.600 3465.640 ;
        RECT 0.270 3462.240 2432.415 3464.240 ;
        RECT 0.270 3460.840 2430.600 3462.240 ;
        RECT 0.270 3458.840 2432.415 3460.840 ;
        RECT 0.270 3457.440 2430.600 3458.840 ;
        RECT 0.270 3455.440 2432.415 3457.440 ;
        RECT 0.270 3454.040 2430.600 3455.440 ;
        RECT 0.270 3452.040 2432.415 3454.040 ;
        RECT 0.270 3450.640 2430.600 3452.040 ;
        RECT 0.270 3448.640 2432.415 3450.640 ;
        RECT 0.270 3447.240 2430.600 3448.640 ;
        RECT 0.270 3445.240 2432.415 3447.240 ;
        RECT 0.270 3443.840 2430.600 3445.240 ;
        RECT 0.270 3441.840 2432.415 3443.840 ;
        RECT 4.400 3440.440 2430.600 3441.840 ;
        RECT 0.270 3438.440 2432.415 3440.440 ;
        RECT 4.400 3437.040 2430.600 3438.440 ;
        RECT 0.270 3435.040 2432.415 3437.040 ;
        RECT 0.270 3433.640 2430.600 3435.040 ;
        RECT 0.270 3431.640 2432.415 3433.640 ;
        RECT 4.400 3430.240 2430.600 3431.640 ;
        RECT 0.270 3428.240 2432.415 3430.240 ;
        RECT 4.400 3426.840 2430.600 3428.240 ;
        RECT 0.270 3424.840 2432.415 3426.840 ;
        RECT 4.400 3423.440 2430.600 3424.840 ;
        RECT 0.270 3421.440 2432.415 3423.440 ;
        RECT 4.400 3420.040 2430.600 3421.440 ;
        RECT 0.270 3418.040 2432.415 3420.040 ;
        RECT 4.400 3416.640 2430.600 3418.040 ;
        RECT 0.270 3414.640 2432.415 3416.640 ;
        RECT 0.270 3413.240 2430.600 3414.640 ;
        RECT 0.270 3411.240 2432.415 3413.240 ;
        RECT 4.400 3409.840 2430.600 3411.240 ;
        RECT 0.270 3407.840 2432.415 3409.840 ;
        RECT 4.400 3406.440 2430.600 3407.840 ;
        RECT 0.270 3404.440 2432.415 3406.440 ;
        RECT 4.400 3403.040 2430.600 3404.440 ;
        RECT 0.270 3401.040 2432.415 3403.040 ;
        RECT 4.400 3399.640 2430.600 3401.040 ;
        RECT 0.270 3397.640 2432.415 3399.640 ;
        RECT 4.400 3396.240 2432.415 3397.640 ;
        RECT 0.270 3390.840 2432.415 3396.240 ;
        RECT 4.400 3389.440 2432.415 3390.840 ;
        RECT 0.270 3387.440 2432.415 3389.440 ;
        RECT 4.400 3386.040 2432.415 3387.440 ;
        RECT 0.270 3384.040 2432.415 3386.040 ;
        RECT 4.400 3382.640 2432.415 3384.040 ;
        RECT 0.270 3380.640 2432.415 3382.640 ;
        RECT 4.400 3379.240 2432.415 3380.640 ;
        RECT 0.270 3377.240 2432.415 3379.240 ;
        RECT 4.400 3375.840 2432.415 3377.240 ;
        RECT 0.270 3370.440 2432.415 3375.840 ;
        RECT 4.400 3369.040 2432.415 3370.440 ;
        RECT 0.270 3367.040 2432.415 3369.040 ;
        RECT 4.400 3365.640 2432.415 3367.040 ;
        RECT 0.270 3363.640 2432.415 3365.640 ;
        RECT 4.400 3362.240 2432.415 3363.640 ;
        RECT 0.270 3360.240 2432.415 3362.240 ;
        RECT 4.400 3358.840 2432.415 3360.240 ;
        RECT 0.270 3356.840 2432.415 3358.840 ;
        RECT 4.400 3355.440 2432.415 3356.840 ;
        RECT 0.270 3350.040 2432.415 3355.440 ;
        RECT 4.400 3348.640 2432.415 3350.040 ;
        RECT 0.270 3346.640 2432.415 3348.640 ;
        RECT 4.400 3345.240 2432.415 3346.640 ;
        RECT 0.270 3343.240 2432.415 3345.240 ;
        RECT 4.400 3341.840 2432.415 3343.240 ;
        RECT 0.270 3339.840 2432.415 3341.840 ;
        RECT 4.400 3338.440 2432.415 3339.840 ;
        RECT 0.270 3336.440 2432.415 3338.440 ;
        RECT 4.400 3335.040 2432.415 3336.440 ;
        RECT 0.270 3329.640 2432.415 3335.040 ;
        RECT 4.400 3328.240 2432.415 3329.640 ;
        RECT 0.270 3326.240 2432.415 3328.240 ;
        RECT 4.400 3324.840 2432.415 3326.240 ;
        RECT 0.270 3322.840 2432.415 3324.840 ;
        RECT 4.400 3321.440 2432.415 3322.840 ;
        RECT 0.270 3319.440 2432.415 3321.440 ;
        RECT 4.400 3318.040 2432.415 3319.440 ;
        RECT 0.270 3316.040 2432.415 3318.040 ;
        RECT 4.400 3314.640 2432.415 3316.040 ;
        RECT 0.270 3309.240 2432.415 3314.640 ;
        RECT 4.400 3307.840 2432.415 3309.240 ;
        RECT 0.270 3305.840 2432.415 3307.840 ;
        RECT 4.400 3304.440 2432.415 3305.840 ;
        RECT 0.270 3302.440 2432.415 3304.440 ;
        RECT 4.400 3301.040 2432.415 3302.440 ;
        RECT 0.270 3299.040 2432.415 3301.040 ;
        RECT 4.400 3297.640 2432.415 3299.040 ;
        RECT 0.270 3295.640 2432.415 3297.640 ;
        RECT 4.400 3294.240 2432.415 3295.640 ;
        RECT 0.270 3288.840 2432.415 3294.240 ;
        RECT 4.400 3287.440 2432.415 3288.840 ;
        RECT 0.270 3285.440 2432.415 3287.440 ;
        RECT 4.400 3284.040 2432.415 3285.440 ;
        RECT 0.270 3282.040 2432.415 3284.040 ;
        RECT 4.400 3280.640 2432.415 3282.040 ;
        RECT 0.270 3278.640 2432.415 3280.640 ;
        RECT 4.400 3277.240 2432.415 3278.640 ;
        RECT 0.270 3275.240 2432.415 3277.240 ;
        RECT 4.400 3273.840 2432.415 3275.240 ;
        RECT 0.270 3268.440 2432.415 3273.840 ;
        RECT 4.400 3267.040 2432.415 3268.440 ;
        RECT 0.270 3265.040 2432.415 3267.040 ;
        RECT 4.400 3263.640 2432.415 3265.040 ;
        RECT 0.270 3261.640 2432.415 3263.640 ;
        RECT 4.400 3260.240 2432.415 3261.640 ;
        RECT 0.270 3258.240 2432.415 3260.240 ;
        RECT 4.400 3256.840 2432.415 3258.240 ;
        RECT 0.270 3217.440 2432.415 3256.840 ;
        RECT 4.400 3216.040 2432.415 3217.440 ;
        RECT 0.270 3210.640 2432.415 3216.040 ;
        RECT 4.400 3209.240 2432.415 3210.640 ;
        RECT 0.270 3207.240 2432.415 3209.240 ;
        RECT 4.400 3205.840 2432.415 3207.240 ;
        RECT 0.270 3203.840 2432.415 3205.840 ;
        RECT 4.400 3202.440 2432.415 3203.840 ;
        RECT 0.270 3200.440 2432.415 3202.440 ;
        RECT 4.400 3199.040 2432.415 3200.440 ;
        RECT 0.270 3197.040 2432.415 3199.040 ;
        RECT 4.400 3195.640 2432.415 3197.040 ;
        RECT 0.270 3190.240 2432.415 3195.640 ;
        RECT 4.400 3188.840 2432.415 3190.240 ;
        RECT 0.270 3186.840 2432.415 3188.840 ;
        RECT 4.400 3185.440 2432.415 3186.840 ;
        RECT 0.270 3183.440 2432.415 3185.440 ;
        RECT 4.400 3182.040 2432.415 3183.440 ;
        RECT 0.270 3180.040 2432.415 3182.040 ;
        RECT 4.400 3178.640 2432.415 3180.040 ;
        RECT 0.270 3176.640 2432.415 3178.640 ;
        RECT 4.400 3175.240 2432.415 3176.640 ;
        RECT 0.270 3169.840 2432.415 3175.240 ;
        RECT 4.400 3168.440 2432.415 3169.840 ;
        RECT 0.270 3166.440 2432.415 3168.440 ;
        RECT 4.400 3165.040 2432.415 3166.440 ;
        RECT 0.270 3163.040 2432.415 3165.040 ;
        RECT 4.400 3161.640 2432.415 3163.040 ;
        RECT 0.270 3159.640 2432.415 3161.640 ;
        RECT 4.400 3158.240 2432.415 3159.640 ;
        RECT 0.270 3156.240 2432.415 3158.240 ;
        RECT 4.400 3154.840 2432.415 3156.240 ;
        RECT 0.270 3152.840 2432.415 3154.840 ;
        RECT 0.270 3151.440 2430.600 3152.840 ;
        RECT 0.270 3149.440 2432.415 3151.440 ;
        RECT 4.400 3148.040 2430.600 3149.440 ;
        RECT 0.270 3146.040 2432.415 3148.040 ;
        RECT 4.400 3144.640 2430.600 3146.040 ;
        RECT 0.270 3142.640 2432.415 3144.640 ;
        RECT 4.400 3141.240 2430.600 3142.640 ;
        RECT 0.270 3139.240 2432.415 3141.240 ;
        RECT 4.400 3137.840 2430.600 3139.240 ;
        RECT 0.270 3135.840 2432.415 3137.840 ;
        RECT 4.400 3134.440 2430.600 3135.840 ;
        RECT 0.270 3132.440 2432.415 3134.440 ;
        RECT 0.270 3131.040 2430.600 3132.440 ;
        RECT 0.270 3129.040 2432.415 3131.040 ;
        RECT 4.400 3127.640 2430.600 3129.040 ;
        RECT 0.270 3125.640 2432.415 3127.640 ;
        RECT 4.400 3124.240 2430.600 3125.640 ;
        RECT 0.270 3122.240 2432.415 3124.240 ;
        RECT 4.400 3120.840 2430.600 3122.240 ;
        RECT 0.270 3118.840 2432.415 3120.840 ;
        RECT 4.400 3117.440 2430.600 3118.840 ;
        RECT 0.270 3115.440 2432.415 3117.440 ;
        RECT 4.400 3114.040 2430.600 3115.440 ;
        RECT 0.270 3112.040 2432.415 3114.040 ;
        RECT 0.270 3110.640 2430.600 3112.040 ;
        RECT 0.270 3108.640 2432.415 3110.640 ;
        RECT 4.400 3107.240 2430.600 3108.640 ;
        RECT 0.270 3105.240 2432.415 3107.240 ;
        RECT 4.400 3103.840 2430.600 3105.240 ;
        RECT 0.270 3101.840 2432.415 3103.840 ;
        RECT 4.400 3100.440 2430.600 3101.840 ;
        RECT 0.270 3098.440 2432.415 3100.440 ;
        RECT 4.400 3097.040 2430.600 3098.440 ;
        RECT 0.270 3095.040 2432.415 3097.040 ;
        RECT 4.400 3093.640 2430.600 3095.040 ;
        RECT 0.270 3091.640 2432.415 3093.640 ;
        RECT 0.270 3090.240 2430.600 3091.640 ;
        RECT 0.270 3088.240 2432.415 3090.240 ;
        RECT 4.400 3086.840 2430.600 3088.240 ;
        RECT 0.270 3084.840 2432.415 3086.840 ;
        RECT 4.400 3083.440 2430.600 3084.840 ;
        RECT 0.270 3081.440 2432.415 3083.440 ;
        RECT 4.400 3080.040 2430.600 3081.440 ;
        RECT 0.270 3078.040 2432.415 3080.040 ;
        RECT 4.400 3076.640 2430.600 3078.040 ;
        RECT 0.270 3074.640 2432.415 3076.640 ;
        RECT 4.400 3073.240 2430.600 3074.640 ;
        RECT 0.270 3071.240 2432.415 3073.240 ;
        RECT 0.270 3069.840 2430.600 3071.240 ;
        RECT 0.270 3067.840 2432.415 3069.840 ;
        RECT 4.400 3066.440 2430.600 3067.840 ;
        RECT 0.270 3064.440 2432.415 3066.440 ;
        RECT 4.400 3063.040 2430.600 3064.440 ;
        RECT 0.270 3061.040 2432.415 3063.040 ;
        RECT 4.400 3059.640 2430.600 3061.040 ;
        RECT 0.270 3057.640 2432.415 3059.640 ;
        RECT 4.400 3056.240 2430.600 3057.640 ;
        RECT 0.270 3054.240 2432.415 3056.240 ;
        RECT 4.400 3052.840 2430.600 3054.240 ;
        RECT 0.270 3050.840 2432.415 3052.840 ;
        RECT 0.270 3049.440 2430.600 3050.840 ;
        RECT 0.270 3047.440 2432.415 3049.440 ;
        RECT 4.400 3046.040 2430.600 3047.440 ;
        RECT 0.270 3044.040 2432.415 3046.040 ;
        RECT 4.400 3042.640 2430.600 3044.040 ;
        RECT 0.270 3040.640 2432.415 3042.640 ;
        RECT 4.400 3039.240 2430.600 3040.640 ;
        RECT 0.270 3037.240 2432.415 3039.240 ;
        RECT 4.400 3035.840 2430.600 3037.240 ;
        RECT 0.270 3033.840 2432.415 3035.840 ;
        RECT 4.400 3032.440 2430.600 3033.840 ;
        RECT 0.270 3030.440 2432.415 3032.440 ;
        RECT 0.270 3029.040 2430.600 3030.440 ;
        RECT 0.270 3027.040 2432.415 3029.040 ;
        RECT 0.270 3025.640 2430.600 3027.040 ;
        RECT 0.270 3023.640 2432.415 3025.640 ;
        RECT 0.270 3022.240 2430.600 3023.640 ;
        RECT 0.270 3020.240 2432.415 3022.240 ;
        RECT 0.270 3018.840 2430.600 3020.240 ;
        RECT 0.270 3016.840 2432.415 3018.840 ;
        RECT 0.270 3015.440 2430.600 3016.840 ;
        RECT 0.270 3013.440 2432.415 3015.440 ;
        RECT 0.270 3012.040 2430.600 3013.440 ;
        RECT 0.270 3010.040 2432.415 3012.040 ;
        RECT 0.270 3008.640 2430.600 3010.040 ;
        RECT 0.270 3006.640 2432.415 3008.640 ;
        RECT 0.270 3005.240 2430.600 3006.640 ;
        RECT 0.270 3003.240 2432.415 3005.240 ;
        RECT 0.270 3001.840 2430.600 3003.240 ;
        RECT 0.270 2999.840 2432.415 3001.840 ;
        RECT 0.270 2998.440 2430.600 2999.840 ;
        RECT 0.270 2996.440 2432.415 2998.440 ;
        RECT 0.270 2995.040 2430.600 2996.440 ;
        RECT 0.270 2993.040 2432.415 2995.040 ;
        RECT 0.270 2991.640 2430.600 2993.040 ;
        RECT 0.270 2989.640 2432.415 2991.640 ;
        RECT 4.400 2988.240 2430.600 2989.640 ;
        RECT 0.270 2986.240 2432.415 2988.240 ;
        RECT 4.400 2984.840 2430.600 2986.240 ;
        RECT 0.270 2982.840 2432.415 2984.840 ;
        RECT 4.400 2981.440 2430.600 2982.840 ;
        RECT 0.270 2979.440 2432.415 2981.440 ;
        RECT 4.400 2978.040 2430.600 2979.440 ;
        RECT 0.270 2976.040 2432.415 2978.040 ;
        RECT 4.400 2974.640 2430.600 2976.040 ;
        RECT 0.270 2972.640 2432.415 2974.640 ;
        RECT 0.270 2971.240 2430.600 2972.640 ;
        RECT 0.270 2969.240 2432.415 2971.240 ;
        RECT 4.400 2967.840 2430.600 2969.240 ;
        RECT 0.270 2965.840 2432.415 2967.840 ;
        RECT 4.400 2964.440 2430.600 2965.840 ;
        RECT 0.270 2962.440 2432.415 2964.440 ;
        RECT 4.400 2961.040 2430.600 2962.440 ;
        RECT 0.270 2959.040 2432.415 2961.040 ;
        RECT 4.400 2957.640 2430.600 2959.040 ;
        RECT 0.270 2955.640 2432.415 2957.640 ;
        RECT 4.400 2954.240 2430.600 2955.640 ;
        RECT 0.270 2952.240 2432.415 2954.240 ;
        RECT 0.270 2950.840 2430.600 2952.240 ;
        RECT 0.270 2948.840 2432.415 2950.840 ;
        RECT 4.400 2947.440 2430.600 2948.840 ;
        RECT 0.270 2945.440 2432.415 2947.440 ;
        RECT 4.400 2944.040 2430.600 2945.440 ;
        RECT 0.270 2942.040 2432.415 2944.040 ;
        RECT 4.400 2940.640 2430.600 2942.040 ;
        RECT 0.270 2938.640 2432.415 2940.640 ;
        RECT 4.400 2937.240 2430.600 2938.640 ;
        RECT 0.270 2935.240 2432.415 2937.240 ;
        RECT 4.400 2933.840 2430.600 2935.240 ;
        RECT 0.270 2931.840 2432.415 2933.840 ;
        RECT 0.270 2930.440 2430.600 2931.840 ;
        RECT 0.270 2928.440 2432.415 2930.440 ;
        RECT 4.400 2927.040 2430.600 2928.440 ;
        RECT 0.270 2925.040 2432.415 2927.040 ;
        RECT 4.400 2923.640 2430.600 2925.040 ;
        RECT 0.270 2921.640 2432.415 2923.640 ;
        RECT 4.400 2920.240 2430.600 2921.640 ;
        RECT 0.270 2918.240 2432.415 2920.240 ;
        RECT 4.400 2916.840 2430.600 2918.240 ;
        RECT 0.270 2914.840 2432.415 2916.840 ;
        RECT 4.400 2913.440 2430.600 2914.840 ;
        RECT 0.270 2911.440 2432.415 2913.440 ;
        RECT 0.270 2910.040 2430.600 2911.440 ;
        RECT 0.270 2908.040 2432.415 2910.040 ;
        RECT 4.400 2906.640 2430.600 2908.040 ;
        RECT 0.270 2904.640 2432.415 2906.640 ;
        RECT 4.400 2903.240 2430.600 2904.640 ;
        RECT 0.270 2901.240 2432.415 2903.240 ;
        RECT 4.400 2899.840 2430.600 2901.240 ;
        RECT 0.270 2897.840 2432.415 2899.840 ;
        RECT 4.400 2896.440 2430.600 2897.840 ;
        RECT 0.270 2894.440 2432.415 2896.440 ;
        RECT 4.400 2893.040 2430.600 2894.440 ;
        RECT 0.270 2891.040 2432.415 2893.040 ;
        RECT 0.270 2889.640 2430.600 2891.040 ;
        RECT 0.270 2887.640 2432.415 2889.640 ;
        RECT 4.400 2886.240 2430.600 2887.640 ;
        RECT 0.270 2884.240 2432.415 2886.240 ;
        RECT 4.400 2882.840 2430.600 2884.240 ;
        RECT 0.270 2880.840 2432.415 2882.840 ;
        RECT 4.400 2879.440 2430.600 2880.840 ;
        RECT 0.270 2877.440 2432.415 2879.440 ;
        RECT 4.400 2876.040 2430.600 2877.440 ;
        RECT 0.270 2874.040 2432.415 2876.040 ;
        RECT 4.400 2872.640 2430.600 2874.040 ;
        RECT 0.270 2870.640 2432.415 2872.640 ;
        RECT 0.270 2869.240 2430.600 2870.640 ;
        RECT 0.270 2867.240 2432.415 2869.240 ;
        RECT 4.400 2865.840 2430.600 2867.240 ;
        RECT 0.270 2863.840 2432.415 2865.840 ;
        RECT 4.400 2862.440 2430.600 2863.840 ;
        RECT 0.270 2860.440 2432.415 2862.440 ;
        RECT 4.400 2859.040 2430.600 2860.440 ;
        RECT 0.270 2857.040 2432.415 2859.040 ;
        RECT 4.400 2855.640 2430.600 2857.040 ;
        RECT 0.270 2853.640 2432.415 2855.640 ;
        RECT 4.400 2852.240 2430.600 2853.640 ;
        RECT 0.270 2850.240 2432.415 2852.240 ;
        RECT 0.270 2848.840 2430.600 2850.240 ;
        RECT 0.270 2846.840 2432.415 2848.840 ;
        RECT 4.400 2845.440 2430.600 2846.840 ;
        RECT 0.270 2843.440 2432.415 2845.440 ;
        RECT 4.400 2842.040 2430.600 2843.440 ;
        RECT 0.270 2840.040 2432.415 2842.040 ;
        RECT 4.400 2838.640 2430.600 2840.040 ;
        RECT 0.270 2836.640 2432.415 2838.640 ;
        RECT 4.400 2835.240 2430.600 2836.640 ;
        RECT 0.270 2833.240 2432.415 2835.240 ;
        RECT 4.400 2831.840 2430.600 2833.240 ;
        RECT 0.270 2829.840 2432.415 2831.840 ;
        RECT 0.270 2828.440 2430.600 2829.840 ;
        RECT 0.270 2826.440 2432.415 2828.440 ;
        RECT 4.400 2825.040 2430.600 2826.440 ;
        RECT 0.270 2823.040 2432.415 2825.040 ;
        RECT 4.400 2821.640 2430.600 2823.040 ;
        RECT 0.270 2819.640 2432.415 2821.640 ;
        RECT 4.400 2818.240 2430.600 2819.640 ;
        RECT 0.270 2816.240 2432.415 2818.240 ;
        RECT 4.400 2814.840 2430.600 2816.240 ;
        RECT 0.270 2812.840 2432.415 2814.840 ;
        RECT 4.400 2811.440 2430.600 2812.840 ;
        RECT 0.270 2809.440 2432.415 2811.440 ;
        RECT 0.270 2808.040 2430.600 2809.440 ;
        RECT 0.270 2806.040 2432.415 2808.040 ;
        RECT 4.400 2804.640 2430.600 2806.040 ;
        RECT 0.270 2802.640 2432.415 2804.640 ;
        RECT 0.270 2801.240 2430.600 2802.640 ;
        RECT 0.270 2799.240 2432.415 2801.240 ;
        RECT 0.270 2797.840 2430.600 2799.240 ;
        RECT 0.270 2795.840 2432.415 2797.840 ;
        RECT 0.270 2794.440 2430.600 2795.840 ;
        RECT 0.270 2792.440 2432.415 2794.440 ;
        RECT 0.270 2791.040 2430.600 2792.440 ;
        RECT 0.270 2789.040 2432.415 2791.040 ;
        RECT 0.270 2787.640 2430.600 2789.040 ;
        RECT 0.270 2785.640 2432.415 2787.640 ;
        RECT 0.270 2784.240 2430.600 2785.640 ;
        RECT 0.270 2765.240 2432.415 2784.240 ;
        RECT 4.400 2763.840 2432.415 2765.240 ;
        RECT 0.270 2761.840 2432.415 2763.840 ;
        RECT 4.400 2760.440 2432.415 2761.840 ;
        RECT 0.270 2758.440 2432.415 2760.440 ;
        RECT 4.400 2757.040 2432.415 2758.440 ;
        RECT 0.270 2755.040 2432.415 2757.040 ;
        RECT 4.400 2753.640 2432.415 2755.040 ;
        RECT 0.270 2751.640 2432.415 2753.640 ;
        RECT 4.400 2750.240 2432.415 2751.640 ;
        RECT 0.270 2744.840 2432.415 2750.240 ;
        RECT 4.400 2743.440 2432.415 2744.840 ;
        RECT 0.270 2741.440 2432.415 2743.440 ;
        RECT 4.400 2740.040 2432.415 2741.440 ;
        RECT 0.270 2738.040 2432.415 2740.040 ;
        RECT 4.400 2736.640 2432.415 2738.040 ;
        RECT 0.270 2734.640 2432.415 2736.640 ;
        RECT 4.400 2733.240 2432.415 2734.640 ;
        RECT 0.270 2731.240 2432.415 2733.240 ;
        RECT 4.400 2729.840 2432.415 2731.240 ;
        RECT 0.270 2724.440 2432.415 2729.840 ;
        RECT 4.400 2723.040 2432.415 2724.440 ;
        RECT 0.270 2721.040 2432.415 2723.040 ;
        RECT 4.400 2719.640 2432.415 2721.040 ;
        RECT 0.270 2717.640 2432.415 2719.640 ;
        RECT 4.400 2716.240 2432.415 2717.640 ;
        RECT 0.270 2714.240 2432.415 2716.240 ;
        RECT 4.400 2712.840 2432.415 2714.240 ;
        RECT 0.270 2710.840 2432.415 2712.840 ;
        RECT 4.400 2709.440 2432.415 2710.840 ;
        RECT 0.270 2704.040 2432.415 2709.440 ;
        RECT 4.400 2702.640 2432.415 2704.040 ;
        RECT 0.270 2700.640 2432.415 2702.640 ;
        RECT 4.400 2699.240 2430.600 2700.640 ;
        RECT 0.270 2697.240 2432.415 2699.240 ;
        RECT 4.400 2695.840 2430.600 2697.240 ;
        RECT 0.270 2693.840 2432.415 2695.840 ;
        RECT 4.400 2692.440 2430.600 2693.840 ;
        RECT 0.270 2690.440 2432.415 2692.440 ;
        RECT 4.400 2689.040 2430.600 2690.440 ;
        RECT 0.270 2687.040 2432.415 2689.040 ;
        RECT 0.270 2685.640 2430.600 2687.040 ;
        RECT 0.270 2683.640 2432.415 2685.640 ;
        RECT 4.400 2682.240 2430.600 2683.640 ;
        RECT 0.270 2680.240 2432.415 2682.240 ;
        RECT 4.400 2678.840 2430.600 2680.240 ;
        RECT 0.270 2676.840 2432.415 2678.840 ;
        RECT 4.400 2675.440 2430.600 2676.840 ;
        RECT 0.270 2673.440 2432.415 2675.440 ;
        RECT 4.400 2672.040 2430.600 2673.440 ;
        RECT 0.270 2670.040 2432.415 2672.040 ;
        RECT 4.400 2668.640 2430.600 2670.040 ;
        RECT 0.270 2666.640 2432.415 2668.640 ;
        RECT 0.270 2665.240 2430.600 2666.640 ;
        RECT 0.270 2663.240 2432.415 2665.240 ;
        RECT 4.400 2661.840 2430.600 2663.240 ;
        RECT 0.270 2659.840 2432.415 2661.840 ;
        RECT 4.400 2658.440 2430.600 2659.840 ;
        RECT 0.270 2656.440 2432.415 2658.440 ;
        RECT 4.400 2655.040 2430.600 2656.440 ;
        RECT 0.270 2653.040 2432.415 2655.040 ;
        RECT 4.400 2651.640 2430.600 2653.040 ;
        RECT 0.270 2649.640 2432.415 2651.640 ;
        RECT 4.400 2648.240 2430.600 2649.640 ;
        RECT 0.270 2646.240 2432.415 2648.240 ;
        RECT 0.270 2644.840 2430.600 2646.240 ;
        RECT 0.270 2642.840 2432.415 2644.840 ;
        RECT 4.400 2641.440 2430.600 2642.840 ;
        RECT 0.270 2639.440 2432.415 2641.440 ;
        RECT 4.400 2638.040 2430.600 2639.440 ;
        RECT 0.270 2636.040 2432.415 2638.040 ;
        RECT 4.400 2634.640 2430.600 2636.040 ;
        RECT 0.270 2632.640 2432.415 2634.640 ;
        RECT 4.400 2631.240 2430.600 2632.640 ;
        RECT 0.270 2629.240 2432.415 2631.240 ;
        RECT 4.400 2627.840 2430.600 2629.240 ;
        RECT 0.270 2625.840 2432.415 2627.840 ;
        RECT 0.270 2624.440 2430.600 2625.840 ;
        RECT 0.270 2622.440 2432.415 2624.440 ;
        RECT 4.400 2621.040 2430.600 2622.440 ;
        RECT 0.270 2619.040 2432.415 2621.040 ;
        RECT 4.400 2617.640 2430.600 2619.040 ;
        RECT 0.270 2615.640 2432.415 2617.640 ;
        RECT 4.400 2614.240 2430.600 2615.640 ;
        RECT 0.270 2612.240 2432.415 2614.240 ;
        RECT 4.400 2610.840 2430.600 2612.240 ;
        RECT 0.270 2608.840 2432.415 2610.840 ;
        RECT 4.400 2607.440 2430.600 2608.840 ;
        RECT 0.270 2605.440 2432.415 2607.440 ;
        RECT 0.270 2604.040 2430.600 2605.440 ;
        RECT 0.270 2602.040 2432.415 2604.040 ;
        RECT 4.400 2600.640 2430.600 2602.040 ;
        RECT 0.270 2598.640 2432.415 2600.640 ;
        RECT 4.400 2597.240 2430.600 2598.640 ;
        RECT 0.270 2595.240 2432.415 2597.240 ;
        RECT 4.400 2593.840 2430.600 2595.240 ;
        RECT 0.270 2591.840 2432.415 2593.840 ;
        RECT 4.400 2590.440 2430.600 2591.840 ;
        RECT 0.270 2588.440 2432.415 2590.440 ;
        RECT 4.400 2587.040 2430.600 2588.440 ;
        RECT 0.270 2585.040 2432.415 2587.040 ;
        RECT 0.270 2583.640 2430.600 2585.040 ;
        RECT 0.270 2581.640 2432.415 2583.640 ;
        RECT 4.400 2580.240 2430.600 2581.640 ;
        RECT 0.270 2578.240 2432.415 2580.240 ;
        RECT 0.270 2576.840 2430.600 2578.240 ;
        RECT 0.270 2574.840 2432.415 2576.840 ;
        RECT 0.270 2573.440 2430.600 2574.840 ;
        RECT 0.270 2571.440 2432.415 2573.440 ;
        RECT 0.270 2570.040 2430.600 2571.440 ;
        RECT 0.270 2568.040 2432.415 2570.040 ;
        RECT 0.270 2566.640 2430.600 2568.040 ;
        RECT 0.270 2564.640 2432.415 2566.640 ;
        RECT 0.270 2563.240 2430.600 2564.640 ;
        RECT 0.270 2561.240 2432.415 2563.240 ;
        RECT 0.270 2559.840 2430.600 2561.240 ;
        RECT 0.270 2557.840 2432.415 2559.840 ;
        RECT 0.270 2556.440 2430.600 2557.840 ;
        RECT 0.270 2554.440 2432.415 2556.440 ;
        RECT 0.270 2553.040 2430.600 2554.440 ;
        RECT 0.270 2551.040 2432.415 2553.040 ;
        RECT 0.270 2549.640 2430.600 2551.040 ;
        RECT 0.270 2547.640 2432.415 2549.640 ;
        RECT 0.270 2546.240 2430.600 2547.640 ;
        RECT 0.270 2544.240 2432.415 2546.240 ;
        RECT 0.270 2542.840 2430.600 2544.240 ;
        RECT 0.270 2540.840 2432.415 2542.840 ;
        RECT 4.400 2539.440 2430.600 2540.840 ;
        RECT 0.270 2537.440 2432.415 2539.440 ;
        RECT 4.400 2536.040 2430.600 2537.440 ;
        RECT 0.270 2534.040 2432.415 2536.040 ;
        RECT 4.400 2532.640 2430.600 2534.040 ;
        RECT 0.270 2530.640 2432.415 2532.640 ;
        RECT 4.400 2529.240 2430.600 2530.640 ;
        RECT 0.270 2527.240 2432.415 2529.240 ;
        RECT 0.270 2525.840 2430.600 2527.240 ;
        RECT 0.270 2523.840 2432.415 2525.840 ;
        RECT 4.400 2522.440 2430.600 2523.840 ;
        RECT 0.270 2520.440 2432.415 2522.440 ;
        RECT 4.400 2519.040 2430.600 2520.440 ;
        RECT 0.270 2517.040 2432.415 2519.040 ;
        RECT 4.400 2515.640 2430.600 2517.040 ;
        RECT 0.270 2513.640 2432.415 2515.640 ;
        RECT 4.400 2512.240 2430.600 2513.640 ;
        RECT 0.270 2510.240 2432.415 2512.240 ;
        RECT 4.400 2508.840 2430.600 2510.240 ;
        RECT 0.270 2506.840 2432.415 2508.840 ;
        RECT 0.270 2505.440 2430.600 2506.840 ;
        RECT 0.270 2503.440 2432.415 2505.440 ;
        RECT 4.400 2502.040 2430.600 2503.440 ;
        RECT 0.270 2500.040 2432.415 2502.040 ;
        RECT 4.400 2498.640 2430.600 2500.040 ;
        RECT 0.270 2496.640 2432.415 2498.640 ;
        RECT 4.400 2495.240 2430.600 2496.640 ;
        RECT 0.270 2493.240 2432.415 2495.240 ;
        RECT 4.400 2491.840 2430.600 2493.240 ;
        RECT 0.270 2489.840 2432.415 2491.840 ;
        RECT 4.400 2488.440 2430.600 2489.840 ;
        RECT 0.270 2486.440 2432.415 2488.440 ;
        RECT 0.270 2485.040 2430.600 2486.440 ;
        RECT 0.270 2483.040 2432.415 2485.040 ;
        RECT 4.400 2481.640 2430.600 2483.040 ;
        RECT 0.270 2479.640 2432.415 2481.640 ;
        RECT 4.400 2478.240 2430.600 2479.640 ;
        RECT 0.270 2476.240 2432.415 2478.240 ;
        RECT 4.400 2474.840 2430.600 2476.240 ;
        RECT 0.270 2472.840 2432.415 2474.840 ;
        RECT 4.400 2471.440 2430.600 2472.840 ;
        RECT 0.270 2469.440 2432.415 2471.440 ;
        RECT 4.400 2468.040 2430.600 2469.440 ;
        RECT 0.270 2466.040 2432.415 2468.040 ;
        RECT 0.270 2464.640 2430.600 2466.040 ;
        RECT 0.270 2462.640 2432.415 2464.640 ;
        RECT 4.400 2461.240 2430.600 2462.640 ;
        RECT 0.270 2459.240 2432.415 2461.240 ;
        RECT 4.400 2457.840 2430.600 2459.240 ;
        RECT 0.270 2455.840 2432.415 2457.840 ;
        RECT 4.400 2454.440 2430.600 2455.840 ;
        RECT 0.270 2452.440 2432.415 2454.440 ;
        RECT 4.400 2451.040 2430.600 2452.440 ;
        RECT 0.270 2449.040 2432.415 2451.040 ;
        RECT 4.400 2447.640 2430.600 2449.040 ;
        RECT 0.270 2445.640 2432.415 2447.640 ;
        RECT 0.270 2444.240 2430.600 2445.640 ;
        RECT 0.270 2442.240 2432.415 2444.240 ;
        RECT 4.400 2440.840 2430.600 2442.240 ;
        RECT 0.270 2438.840 2432.415 2440.840 ;
        RECT 4.400 2437.440 2430.600 2438.840 ;
        RECT 0.270 2435.440 2432.415 2437.440 ;
        RECT 4.400 2434.040 2430.600 2435.440 ;
        RECT 0.270 2432.040 2432.415 2434.040 ;
        RECT 4.400 2430.640 2430.600 2432.040 ;
        RECT 0.270 2428.640 2432.415 2430.640 ;
        RECT 4.400 2427.240 2430.600 2428.640 ;
        RECT 0.270 2425.240 2432.415 2427.240 ;
        RECT 0.270 2423.840 2430.600 2425.240 ;
        RECT 0.270 2421.840 2432.415 2423.840 ;
        RECT 4.400 2420.440 2430.600 2421.840 ;
        RECT 0.270 2418.440 2432.415 2420.440 ;
        RECT 4.400 2417.040 2430.600 2418.440 ;
        RECT 0.270 2415.040 2432.415 2417.040 ;
        RECT 4.400 2413.640 2430.600 2415.040 ;
        RECT 0.270 2411.640 2432.415 2413.640 ;
        RECT 4.400 2410.240 2430.600 2411.640 ;
        RECT 0.270 2408.240 2432.415 2410.240 ;
        RECT 4.400 2406.840 2430.600 2408.240 ;
        RECT 0.270 2404.840 2432.415 2406.840 ;
        RECT 0.270 2403.440 2430.600 2404.840 ;
        RECT 0.270 2401.440 2432.415 2403.440 ;
        RECT 4.400 2400.040 2430.600 2401.440 ;
        RECT 0.270 2398.040 2432.415 2400.040 ;
        RECT 4.400 2396.640 2430.600 2398.040 ;
        RECT 0.270 2394.640 2432.415 2396.640 ;
        RECT 4.400 2393.240 2430.600 2394.640 ;
        RECT 0.270 2391.240 2432.415 2393.240 ;
        RECT 4.400 2389.840 2430.600 2391.240 ;
        RECT 0.270 2387.840 2432.415 2389.840 ;
        RECT 4.400 2386.440 2430.600 2387.840 ;
        RECT 0.270 2384.440 2432.415 2386.440 ;
        RECT 0.270 2383.040 2430.600 2384.440 ;
        RECT 0.270 2381.040 2432.415 2383.040 ;
        RECT 4.400 2379.640 2430.600 2381.040 ;
        RECT 0.270 2377.640 2432.415 2379.640 ;
        RECT 4.400 2376.240 2430.600 2377.640 ;
        RECT 0.270 2374.240 2432.415 2376.240 ;
        RECT 4.400 2372.840 2430.600 2374.240 ;
        RECT 0.270 2370.840 2432.415 2372.840 ;
        RECT 4.400 2369.440 2430.600 2370.840 ;
        RECT 0.270 2367.440 2432.415 2369.440 ;
        RECT 4.400 2366.040 2430.600 2367.440 ;
        RECT 0.270 2364.040 2432.415 2366.040 ;
        RECT 0.270 2362.640 2430.600 2364.040 ;
        RECT 0.270 2360.640 2432.415 2362.640 ;
        RECT 4.400 2359.240 2430.600 2360.640 ;
        RECT 0.270 2357.240 2432.415 2359.240 ;
        RECT 4.400 2355.840 2430.600 2357.240 ;
        RECT 0.270 2353.840 2432.415 2355.840 ;
        RECT 0.270 2352.440 2430.600 2353.840 ;
        RECT 0.270 2350.440 2432.415 2352.440 ;
        RECT 0.270 2349.040 2430.600 2350.440 ;
        RECT 0.270 2347.040 2432.415 2349.040 ;
        RECT 0.270 2345.640 2430.600 2347.040 ;
        RECT 0.270 2343.640 2432.415 2345.640 ;
        RECT 0.270 2342.240 2430.600 2343.640 ;
        RECT 0.270 2340.240 2432.415 2342.240 ;
        RECT 0.270 2338.840 2430.600 2340.240 ;
        RECT 0.270 2336.840 2432.415 2338.840 ;
        RECT 0.270 2335.440 2430.600 2336.840 ;
        RECT 0.270 2333.440 2432.415 2335.440 ;
        RECT 0.270 2332.040 2430.600 2333.440 ;
        RECT 0.270 2316.440 2432.415 2332.040 ;
        RECT 4.400 2315.040 2432.415 2316.440 ;
        RECT 0.270 2313.040 2432.415 2315.040 ;
        RECT 4.400 2311.640 2432.415 2313.040 ;
        RECT 0.270 2309.640 2432.415 2311.640 ;
        RECT 4.400 2308.240 2432.415 2309.640 ;
        RECT 0.270 2302.840 2432.415 2308.240 ;
        RECT 4.400 2301.440 2432.415 2302.840 ;
        RECT 0.270 2299.440 2432.415 2301.440 ;
        RECT 4.400 2298.040 2430.600 2299.440 ;
        RECT 0.270 2296.040 2432.415 2298.040 ;
        RECT 4.400 2294.640 2430.600 2296.040 ;
        RECT 0.270 2292.640 2432.415 2294.640 ;
        RECT 4.400 2291.240 2430.600 2292.640 ;
        RECT 0.270 2289.240 2432.415 2291.240 ;
        RECT 4.400 2287.840 2430.600 2289.240 ;
        RECT 0.270 2285.840 2432.415 2287.840 ;
        RECT 0.270 2284.440 2430.600 2285.840 ;
        RECT 0.270 2282.440 2432.415 2284.440 ;
        RECT 4.400 2281.040 2430.600 2282.440 ;
        RECT 0.270 2279.040 2432.415 2281.040 ;
        RECT 4.400 2277.640 2430.600 2279.040 ;
        RECT 0.270 2275.640 2432.415 2277.640 ;
        RECT 4.400 2274.240 2430.600 2275.640 ;
        RECT 0.270 2272.240 2432.415 2274.240 ;
        RECT 4.400 2270.840 2430.600 2272.240 ;
        RECT 0.270 2268.840 2432.415 2270.840 ;
        RECT 4.400 2267.440 2430.600 2268.840 ;
        RECT 0.270 2265.440 2432.415 2267.440 ;
        RECT 0.270 2264.040 2430.600 2265.440 ;
        RECT 0.270 2262.040 2432.415 2264.040 ;
        RECT 4.400 2260.640 2430.600 2262.040 ;
        RECT 0.270 2258.640 2432.415 2260.640 ;
        RECT 4.400 2257.240 2430.600 2258.640 ;
        RECT 0.270 2255.240 2432.415 2257.240 ;
        RECT 4.400 2253.840 2430.600 2255.240 ;
        RECT 0.270 2251.840 2432.415 2253.840 ;
        RECT 4.400 2250.440 2430.600 2251.840 ;
        RECT 0.270 2248.440 2432.415 2250.440 ;
        RECT 4.400 2247.040 2430.600 2248.440 ;
        RECT 0.270 2245.040 2432.415 2247.040 ;
        RECT 0.270 2243.640 2430.600 2245.040 ;
        RECT 0.270 2241.640 2432.415 2243.640 ;
        RECT 4.400 2240.240 2430.600 2241.640 ;
        RECT 0.270 2238.240 2432.415 2240.240 ;
        RECT 4.400 2236.840 2430.600 2238.240 ;
        RECT 0.270 2234.840 2432.415 2236.840 ;
        RECT 4.400 2233.440 2430.600 2234.840 ;
        RECT 0.270 2231.440 2432.415 2233.440 ;
        RECT 4.400 2230.040 2430.600 2231.440 ;
        RECT 0.270 2228.040 2432.415 2230.040 ;
        RECT 4.400 2226.640 2430.600 2228.040 ;
        RECT 0.270 2224.640 2432.415 2226.640 ;
        RECT 0.270 2223.240 2430.600 2224.640 ;
        RECT 0.270 2221.240 2432.415 2223.240 ;
        RECT 4.400 2219.840 2430.600 2221.240 ;
        RECT 0.270 2217.840 2432.415 2219.840 ;
        RECT 4.400 2216.440 2430.600 2217.840 ;
        RECT 0.270 2214.440 2432.415 2216.440 ;
        RECT 4.400 2213.040 2430.600 2214.440 ;
        RECT 0.270 2211.040 2432.415 2213.040 ;
        RECT 4.400 2209.640 2430.600 2211.040 ;
        RECT 0.270 2207.640 2432.415 2209.640 ;
        RECT 4.400 2206.240 2430.600 2207.640 ;
        RECT 0.270 2204.240 2432.415 2206.240 ;
        RECT 0.270 2202.840 2430.600 2204.240 ;
        RECT 0.270 2200.840 2432.415 2202.840 ;
        RECT 4.400 2199.440 2430.600 2200.840 ;
        RECT 0.270 2197.440 2432.415 2199.440 ;
        RECT 4.400 2196.040 2430.600 2197.440 ;
        RECT 0.270 2194.040 2432.415 2196.040 ;
        RECT 4.400 2192.640 2430.600 2194.040 ;
        RECT 0.270 2190.640 2432.415 2192.640 ;
        RECT 4.400 2189.240 2430.600 2190.640 ;
        RECT 0.270 2187.240 2432.415 2189.240 ;
        RECT 4.400 2185.840 2430.600 2187.240 ;
        RECT 0.270 2183.840 2432.415 2185.840 ;
        RECT 0.270 2182.440 2430.600 2183.840 ;
        RECT 0.270 2180.440 2432.415 2182.440 ;
        RECT 4.400 2179.040 2430.600 2180.440 ;
        RECT 0.270 2177.040 2432.415 2179.040 ;
        RECT 4.400 2175.640 2430.600 2177.040 ;
        RECT 0.270 2173.640 2432.415 2175.640 ;
        RECT 4.400 2172.240 2430.600 2173.640 ;
        RECT 0.270 2170.240 2432.415 2172.240 ;
        RECT 4.400 2168.840 2430.600 2170.240 ;
        RECT 0.270 2166.840 2432.415 2168.840 ;
        RECT 4.400 2165.440 2430.600 2166.840 ;
        RECT 0.270 2163.440 2432.415 2165.440 ;
        RECT 0.270 2162.040 2430.600 2163.440 ;
        RECT 0.270 2160.040 2432.415 2162.040 ;
        RECT 4.400 2158.640 2430.600 2160.040 ;
        RECT 0.270 2156.640 2432.415 2158.640 ;
        RECT 4.400 2155.240 2430.600 2156.640 ;
        RECT 0.270 2153.240 2432.415 2155.240 ;
        RECT 4.400 2151.840 2430.600 2153.240 ;
        RECT 0.270 2149.840 2432.415 2151.840 ;
        RECT 4.400 2148.440 2430.600 2149.840 ;
        RECT 0.270 2146.440 2432.415 2148.440 ;
        RECT 4.400 2145.040 2430.600 2146.440 ;
        RECT 0.270 2143.040 2432.415 2145.040 ;
        RECT 0.270 2141.640 2430.600 2143.040 ;
        RECT 0.270 2139.640 2432.415 2141.640 ;
        RECT 4.400 2138.240 2430.600 2139.640 ;
        RECT 0.270 2136.240 2432.415 2138.240 ;
        RECT 4.400 2134.840 2430.600 2136.240 ;
        RECT 0.270 2132.840 2432.415 2134.840 ;
        RECT 4.400 2131.440 2430.600 2132.840 ;
        RECT 0.270 2129.440 2432.415 2131.440 ;
        RECT 0.270 2128.040 2430.600 2129.440 ;
        RECT 0.270 2126.040 2432.415 2128.040 ;
        RECT 0.270 2124.640 2430.600 2126.040 ;
        RECT 0.270 2122.640 2432.415 2124.640 ;
        RECT 0.270 2121.240 2430.600 2122.640 ;
        RECT 0.270 2119.240 2432.415 2121.240 ;
        RECT 0.270 2117.840 2430.600 2119.240 ;
        RECT 0.270 2115.840 2432.415 2117.840 ;
        RECT 0.270 2114.440 2430.600 2115.840 ;
        RECT 0.270 2112.440 2432.415 2114.440 ;
        RECT 0.270 2111.040 2430.600 2112.440 ;
        RECT 0.270 2109.040 2432.415 2111.040 ;
        RECT 0.270 2107.640 2430.600 2109.040 ;
        RECT 0.270 2105.640 2432.415 2107.640 ;
        RECT 0.270 2104.240 2430.600 2105.640 ;
        RECT 0.270 2102.240 2432.415 2104.240 ;
        RECT 0.270 2100.840 2430.600 2102.240 ;
        RECT 0.270 2098.840 2432.415 2100.840 ;
        RECT 0.270 2097.440 2430.600 2098.840 ;
        RECT 0.270 2095.440 2432.415 2097.440 ;
        RECT 0.270 2094.040 2430.600 2095.440 ;
        RECT 0.270 2092.040 2432.415 2094.040 ;
        RECT 4.400 2090.640 2430.600 2092.040 ;
        RECT 0.270 2088.640 2432.415 2090.640 ;
        RECT 4.400 2087.240 2430.600 2088.640 ;
        RECT 0.270 2085.240 2432.415 2087.240 ;
        RECT 0.270 2083.840 2430.600 2085.240 ;
        RECT 0.270 2081.840 2432.415 2083.840 ;
        RECT 4.400 2080.440 2430.600 2081.840 ;
        RECT 0.270 2078.440 2432.415 2080.440 ;
        RECT 4.400 2077.040 2430.600 2078.440 ;
        RECT 0.270 2075.040 2432.415 2077.040 ;
        RECT 4.400 2073.640 2430.600 2075.040 ;
        RECT 0.270 2071.640 2432.415 2073.640 ;
        RECT 4.400 2070.240 2430.600 2071.640 ;
        RECT 0.270 2068.240 2432.415 2070.240 ;
        RECT 4.400 2066.840 2430.600 2068.240 ;
        RECT 0.270 2064.840 2432.415 2066.840 ;
        RECT 0.270 2063.440 2430.600 2064.840 ;
        RECT 0.270 2061.440 2432.415 2063.440 ;
        RECT 4.400 2060.040 2430.600 2061.440 ;
        RECT 0.270 2058.040 2432.415 2060.040 ;
        RECT 4.400 2056.640 2430.600 2058.040 ;
        RECT 0.270 2054.640 2432.415 2056.640 ;
        RECT 4.400 2053.240 2430.600 2054.640 ;
        RECT 0.270 2051.240 2432.415 2053.240 ;
        RECT 4.400 2049.840 2430.600 2051.240 ;
        RECT 0.270 2047.840 2432.415 2049.840 ;
        RECT 4.400 2046.440 2430.600 2047.840 ;
        RECT 0.270 2044.440 2432.415 2046.440 ;
        RECT 0.270 2043.040 2430.600 2044.440 ;
        RECT 0.270 2041.040 2432.415 2043.040 ;
        RECT 4.400 2039.640 2430.600 2041.040 ;
        RECT 0.270 2037.640 2432.415 2039.640 ;
        RECT 4.400 2036.240 2430.600 2037.640 ;
        RECT 0.270 2034.240 2432.415 2036.240 ;
        RECT 4.400 2032.840 2430.600 2034.240 ;
        RECT 0.270 2030.840 2432.415 2032.840 ;
        RECT 4.400 2029.440 2430.600 2030.840 ;
        RECT 0.270 2027.440 2432.415 2029.440 ;
        RECT 4.400 2026.040 2430.600 2027.440 ;
        RECT 0.270 2024.040 2432.415 2026.040 ;
        RECT 0.270 2022.640 2430.600 2024.040 ;
        RECT 0.270 2020.640 2432.415 2022.640 ;
        RECT 4.400 2019.240 2430.600 2020.640 ;
        RECT 0.270 2017.240 2432.415 2019.240 ;
        RECT 4.400 2015.840 2430.600 2017.240 ;
        RECT 0.270 2013.840 2432.415 2015.840 ;
        RECT 4.400 2012.440 2430.600 2013.840 ;
        RECT 0.270 2010.440 2432.415 2012.440 ;
        RECT 4.400 2009.040 2430.600 2010.440 ;
        RECT 0.270 2007.040 2432.415 2009.040 ;
        RECT 4.400 2005.640 2430.600 2007.040 ;
        RECT 0.270 2003.640 2432.415 2005.640 ;
        RECT 0.270 2002.240 2430.600 2003.640 ;
        RECT 0.270 2000.240 2432.415 2002.240 ;
        RECT 4.400 1998.840 2430.600 2000.240 ;
        RECT 0.270 1996.840 2432.415 1998.840 ;
        RECT 4.400 1995.440 2430.600 1996.840 ;
        RECT 0.270 1993.440 2432.415 1995.440 ;
        RECT 4.400 1992.040 2430.600 1993.440 ;
        RECT 0.270 1990.040 2432.415 1992.040 ;
        RECT 4.400 1988.640 2430.600 1990.040 ;
        RECT 0.270 1986.640 2432.415 1988.640 ;
        RECT 4.400 1985.240 2430.600 1986.640 ;
        RECT 0.270 1983.240 2432.415 1985.240 ;
        RECT 0.270 1981.840 2430.600 1983.240 ;
        RECT 0.270 1979.840 2432.415 1981.840 ;
        RECT 4.400 1978.440 2430.600 1979.840 ;
        RECT 0.270 1976.440 2432.415 1978.440 ;
        RECT 4.400 1975.040 2430.600 1976.440 ;
        RECT 0.270 1973.040 2432.415 1975.040 ;
        RECT 4.400 1971.640 2430.600 1973.040 ;
        RECT 0.270 1969.640 2432.415 1971.640 ;
        RECT 4.400 1968.240 2430.600 1969.640 ;
        RECT 0.270 1966.240 2432.415 1968.240 ;
        RECT 4.400 1964.840 2430.600 1966.240 ;
        RECT 0.270 1962.840 2432.415 1964.840 ;
        RECT 0.270 1961.440 2430.600 1962.840 ;
        RECT 0.270 1959.440 2432.415 1961.440 ;
        RECT 4.400 1958.040 2430.600 1959.440 ;
        RECT 0.270 1956.040 2432.415 1958.040 ;
        RECT 4.400 1954.640 2430.600 1956.040 ;
        RECT 0.270 1952.640 2432.415 1954.640 ;
        RECT 4.400 1951.240 2430.600 1952.640 ;
        RECT 0.270 1949.240 2432.415 1951.240 ;
        RECT 4.400 1947.840 2430.600 1949.240 ;
        RECT 0.270 1945.840 2432.415 1947.840 ;
        RECT 4.400 1944.440 2430.600 1945.840 ;
        RECT 0.270 1942.440 2432.415 1944.440 ;
        RECT 0.270 1941.040 2430.600 1942.440 ;
        RECT 0.270 1939.040 2432.415 1941.040 ;
        RECT 4.400 1937.640 2430.600 1939.040 ;
        RECT 0.270 1935.640 2432.415 1937.640 ;
        RECT 4.400 1934.240 2430.600 1935.640 ;
        RECT 0.270 1932.240 2432.415 1934.240 ;
        RECT 4.400 1930.840 2430.600 1932.240 ;
        RECT 0.270 1928.840 2432.415 1930.840 ;
        RECT 4.400 1927.440 2432.415 1928.840 ;
        RECT 0.270 1925.440 2432.415 1927.440 ;
        RECT 4.400 1924.040 2432.415 1925.440 ;
        RECT 0.270 1918.640 2432.415 1924.040 ;
        RECT 4.400 1917.240 2432.415 1918.640 ;
        RECT 0.270 1915.240 2432.415 1917.240 ;
        RECT 4.400 1913.840 2432.415 1915.240 ;
        RECT 0.270 1911.840 2432.415 1913.840 ;
        RECT 4.400 1910.440 2432.415 1911.840 ;
        RECT 0.270 1908.440 2432.415 1910.440 ;
        RECT 4.400 1907.040 2432.415 1908.440 ;
        RECT 0.270 1867.640 2432.415 1907.040 ;
        RECT 4.400 1866.240 2432.415 1867.640 ;
        RECT 0.270 1860.840 2432.415 1866.240 ;
        RECT 4.400 1859.440 2432.415 1860.840 ;
        RECT 0.270 1857.440 2432.415 1859.440 ;
        RECT 4.400 1856.040 2432.415 1857.440 ;
        RECT 0.270 1854.040 2432.415 1856.040 ;
        RECT 4.400 1852.640 2432.415 1854.040 ;
        RECT 0.270 1850.640 2432.415 1852.640 ;
        RECT 4.400 1849.240 2432.415 1850.640 ;
        RECT 0.270 1847.240 2432.415 1849.240 ;
        RECT 4.400 1845.840 2432.415 1847.240 ;
        RECT 0.270 1840.440 2432.415 1845.840 ;
        RECT 4.400 1839.040 2432.415 1840.440 ;
        RECT 0.270 1837.040 2432.415 1839.040 ;
        RECT 4.400 1835.640 2432.415 1837.040 ;
        RECT 0.270 1833.640 2432.415 1835.640 ;
        RECT 4.400 1832.240 2432.415 1833.640 ;
        RECT 0.270 1830.240 2432.415 1832.240 ;
        RECT 4.400 1828.840 2432.415 1830.240 ;
        RECT 0.270 1826.840 2432.415 1828.840 ;
        RECT 4.400 1825.440 2432.415 1826.840 ;
        RECT 0.270 1820.040 2432.415 1825.440 ;
        RECT 4.400 1818.640 2432.415 1820.040 ;
        RECT 0.270 1816.640 2432.415 1818.640 ;
        RECT 4.400 1815.240 2432.415 1816.640 ;
        RECT 0.270 1813.240 2432.415 1815.240 ;
        RECT 4.400 1811.840 2432.415 1813.240 ;
        RECT 0.270 1809.840 2432.415 1811.840 ;
        RECT 4.400 1808.440 2432.415 1809.840 ;
        RECT 0.270 1806.440 2432.415 1808.440 ;
        RECT 4.400 1805.040 2432.415 1806.440 ;
        RECT 0.270 1803.040 2432.415 1805.040 ;
        RECT 0.270 1801.640 2430.600 1803.040 ;
        RECT 0.270 1799.640 2432.415 1801.640 ;
        RECT 4.400 1798.240 2430.600 1799.640 ;
        RECT 0.270 1796.240 2432.415 1798.240 ;
        RECT 4.400 1794.840 2430.600 1796.240 ;
        RECT 0.270 1792.840 2432.415 1794.840 ;
        RECT 4.400 1791.440 2430.600 1792.840 ;
        RECT 0.270 1789.440 2432.415 1791.440 ;
        RECT 4.400 1788.040 2430.600 1789.440 ;
        RECT 0.270 1786.040 2432.415 1788.040 ;
        RECT 4.400 1784.640 2430.600 1786.040 ;
        RECT 0.270 1782.640 2432.415 1784.640 ;
        RECT 0.270 1781.240 2430.600 1782.640 ;
        RECT 0.270 1779.240 2432.415 1781.240 ;
        RECT 4.400 1777.840 2430.600 1779.240 ;
        RECT 0.270 1775.840 2432.415 1777.840 ;
        RECT 4.400 1774.440 2430.600 1775.840 ;
        RECT 0.270 1772.440 2432.415 1774.440 ;
        RECT 4.400 1771.040 2430.600 1772.440 ;
        RECT 0.270 1769.040 2432.415 1771.040 ;
        RECT 4.400 1767.640 2430.600 1769.040 ;
        RECT 0.270 1765.640 2432.415 1767.640 ;
        RECT 4.400 1764.240 2430.600 1765.640 ;
        RECT 0.270 1762.240 2432.415 1764.240 ;
        RECT 0.270 1760.840 2430.600 1762.240 ;
        RECT 0.270 1758.840 2432.415 1760.840 ;
        RECT 4.400 1757.440 2430.600 1758.840 ;
        RECT 0.270 1755.440 2432.415 1757.440 ;
        RECT 4.400 1754.040 2430.600 1755.440 ;
        RECT 0.270 1752.040 2432.415 1754.040 ;
        RECT 4.400 1750.640 2430.600 1752.040 ;
        RECT 0.270 1748.640 2432.415 1750.640 ;
        RECT 4.400 1747.240 2430.600 1748.640 ;
        RECT 0.270 1745.240 2432.415 1747.240 ;
        RECT 0.270 1743.840 2430.600 1745.240 ;
        RECT 0.270 1741.840 2432.415 1743.840 ;
        RECT 4.400 1740.440 2430.600 1741.840 ;
        RECT 0.270 1738.440 2432.415 1740.440 ;
        RECT 4.400 1737.040 2430.600 1738.440 ;
        RECT 0.270 1735.040 2432.415 1737.040 ;
        RECT 4.400 1733.640 2430.600 1735.040 ;
        RECT 0.270 1731.640 2432.415 1733.640 ;
        RECT 4.400 1730.240 2430.600 1731.640 ;
        RECT 0.270 1728.240 2432.415 1730.240 ;
        RECT 4.400 1726.840 2430.600 1728.240 ;
        RECT 0.270 1724.840 2432.415 1726.840 ;
        RECT 4.400 1723.440 2430.600 1724.840 ;
        RECT 0.270 1721.440 2432.415 1723.440 ;
        RECT 0.270 1720.040 2430.600 1721.440 ;
        RECT 0.270 1718.040 2432.415 1720.040 ;
        RECT 4.400 1716.640 2430.600 1718.040 ;
        RECT 0.270 1714.640 2432.415 1716.640 ;
        RECT 4.400 1713.240 2430.600 1714.640 ;
        RECT 0.270 1711.240 2432.415 1713.240 ;
        RECT 4.400 1709.840 2430.600 1711.240 ;
        RECT 0.270 1707.840 2432.415 1709.840 ;
        RECT 4.400 1706.440 2430.600 1707.840 ;
        RECT 0.270 1704.440 2432.415 1706.440 ;
        RECT 4.400 1703.040 2430.600 1704.440 ;
        RECT 0.270 1701.040 2432.415 1703.040 ;
        RECT 0.270 1699.640 2430.600 1701.040 ;
        RECT 0.270 1697.640 2432.415 1699.640 ;
        RECT 4.400 1696.240 2430.600 1697.640 ;
        RECT 0.270 1694.240 2432.415 1696.240 ;
        RECT 4.400 1692.840 2430.600 1694.240 ;
        RECT 0.270 1690.840 2432.415 1692.840 ;
        RECT 4.400 1689.440 2430.600 1690.840 ;
        RECT 0.270 1687.440 2432.415 1689.440 ;
        RECT 4.400 1686.040 2430.600 1687.440 ;
        RECT 0.270 1684.040 2432.415 1686.040 ;
        RECT 4.400 1682.640 2430.600 1684.040 ;
        RECT 0.270 1680.640 2432.415 1682.640 ;
        RECT 0.270 1679.240 2430.600 1680.640 ;
        RECT 0.270 1677.240 2432.415 1679.240 ;
        RECT 0.270 1675.840 2430.600 1677.240 ;
        RECT 0.270 1673.840 2432.415 1675.840 ;
        RECT 0.270 1672.440 2430.600 1673.840 ;
        RECT 0.270 1670.440 2432.415 1672.440 ;
        RECT 0.270 1669.040 2430.600 1670.440 ;
        RECT 0.270 1667.040 2432.415 1669.040 ;
        RECT 0.270 1665.640 2430.600 1667.040 ;
        RECT 0.270 1663.640 2432.415 1665.640 ;
        RECT 0.270 1662.240 2430.600 1663.640 ;
        RECT 0.270 1660.240 2432.415 1662.240 ;
        RECT 0.270 1658.840 2430.600 1660.240 ;
        RECT 0.270 1656.840 2432.415 1658.840 ;
        RECT 0.270 1655.440 2430.600 1656.840 ;
        RECT 0.270 1653.440 2432.415 1655.440 ;
        RECT 0.270 1652.040 2430.600 1653.440 ;
        RECT 0.270 1650.040 2432.415 1652.040 ;
        RECT 0.270 1648.640 2430.600 1650.040 ;
        RECT 0.270 1646.640 2432.415 1648.640 ;
        RECT 0.270 1645.240 2430.600 1646.640 ;
        RECT 0.270 1643.240 2432.415 1645.240 ;
        RECT 0.270 1641.840 2430.600 1643.240 ;
        RECT 0.270 1639.840 2432.415 1641.840 ;
        RECT 4.400 1638.440 2430.600 1639.840 ;
        RECT 0.270 1636.440 2432.415 1638.440 ;
        RECT 4.400 1635.040 2430.600 1636.440 ;
        RECT 0.270 1633.040 2432.415 1635.040 ;
        RECT 4.400 1631.640 2430.600 1633.040 ;
        RECT 0.270 1629.640 2432.415 1631.640 ;
        RECT 4.400 1628.240 2430.600 1629.640 ;
        RECT 0.270 1626.240 2432.415 1628.240 ;
        RECT 4.400 1624.840 2430.600 1626.240 ;
        RECT 0.270 1622.840 2432.415 1624.840 ;
        RECT 0.270 1621.440 2430.600 1622.840 ;
        RECT 0.270 1619.440 2432.415 1621.440 ;
        RECT 4.400 1618.040 2430.600 1619.440 ;
        RECT 0.270 1616.040 2432.415 1618.040 ;
        RECT 4.400 1614.640 2430.600 1616.040 ;
        RECT 0.270 1612.640 2432.415 1614.640 ;
        RECT 4.400 1611.240 2430.600 1612.640 ;
        RECT 0.270 1609.240 2432.415 1611.240 ;
        RECT 4.400 1607.840 2430.600 1609.240 ;
        RECT 0.270 1605.840 2432.415 1607.840 ;
        RECT 4.400 1604.440 2430.600 1605.840 ;
        RECT 0.270 1602.440 2432.415 1604.440 ;
        RECT 0.270 1601.040 2430.600 1602.440 ;
        RECT 0.270 1599.040 2432.415 1601.040 ;
        RECT 4.400 1597.640 2430.600 1599.040 ;
        RECT 0.270 1595.640 2432.415 1597.640 ;
        RECT 4.400 1594.240 2430.600 1595.640 ;
        RECT 0.270 1592.240 2432.415 1594.240 ;
        RECT 4.400 1590.840 2430.600 1592.240 ;
        RECT 0.270 1588.840 2432.415 1590.840 ;
        RECT 4.400 1587.440 2430.600 1588.840 ;
        RECT 0.270 1585.440 2432.415 1587.440 ;
        RECT 4.400 1584.040 2430.600 1585.440 ;
        RECT 0.270 1582.040 2432.415 1584.040 ;
        RECT 0.270 1580.640 2430.600 1582.040 ;
        RECT 0.270 1578.640 2432.415 1580.640 ;
        RECT 4.400 1577.240 2430.600 1578.640 ;
        RECT 0.270 1575.240 2432.415 1577.240 ;
        RECT 4.400 1573.840 2430.600 1575.240 ;
        RECT 0.270 1571.840 2432.415 1573.840 ;
        RECT 4.400 1570.440 2430.600 1571.840 ;
        RECT 0.270 1568.440 2432.415 1570.440 ;
        RECT 4.400 1567.040 2430.600 1568.440 ;
        RECT 0.270 1565.040 2432.415 1567.040 ;
        RECT 4.400 1563.640 2430.600 1565.040 ;
        RECT 0.270 1561.640 2432.415 1563.640 ;
        RECT 0.270 1560.240 2430.600 1561.640 ;
        RECT 0.270 1558.240 2432.415 1560.240 ;
        RECT 4.400 1556.840 2430.600 1558.240 ;
        RECT 0.270 1554.840 2432.415 1556.840 ;
        RECT 4.400 1553.440 2430.600 1554.840 ;
        RECT 0.270 1551.440 2432.415 1553.440 ;
        RECT 4.400 1550.040 2430.600 1551.440 ;
        RECT 0.270 1548.040 2432.415 1550.040 ;
        RECT 4.400 1546.640 2430.600 1548.040 ;
        RECT 0.270 1544.640 2432.415 1546.640 ;
        RECT 4.400 1543.240 2430.600 1544.640 ;
        RECT 0.270 1541.240 2432.415 1543.240 ;
        RECT 0.270 1539.840 2430.600 1541.240 ;
        RECT 0.270 1537.840 2432.415 1539.840 ;
        RECT 4.400 1536.440 2430.600 1537.840 ;
        RECT 0.270 1534.440 2432.415 1536.440 ;
        RECT 4.400 1533.040 2430.600 1534.440 ;
        RECT 0.270 1531.040 2432.415 1533.040 ;
        RECT 4.400 1529.640 2430.600 1531.040 ;
        RECT 0.270 1527.640 2432.415 1529.640 ;
        RECT 4.400 1526.240 2430.600 1527.640 ;
        RECT 0.270 1524.240 2432.415 1526.240 ;
        RECT 4.400 1522.840 2430.600 1524.240 ;
        RECT 0.270 1520.840 2432.415 1522.840 ;
        RECT 0.270 1519.440 2430.600 1520.840 ;
        RECT 0.270 1517.440 2432.415 1519.440 ;
        RECT 4.400 1516.040 2430.600 1517.440 ;
        RECT 0.270 1514.040 2432.415 1516.040 ;
        RECT 4.400 1512.640 2430.600 1514.040 ;
        RECT 0.270 1510.640 2432.415 1512.640 ;
        RECT 4.400 1509.240 2430.600 1510.640 ;
        RECT 0.270 1507.240 2432.415 1509.240 ;
        RECT 4.400 1505.840 2430.600 1507.240 ;
        RECT 0.270 1503.840 2432.415 1505.840 ;
        RECT 4.400 1502.440 2430.600 1503.840 ;
        RECT 0.270 1500.440 2432.415 1502.440 ;
        RECT 0.270 1499.040 2430.600 1500.440 ;
        RECT 0.270 1497.040 2432.415 1499.040 ;
        RECT 4.400 1495.640 2430.600 1497.040 ;
        RECT 0.270 1493.640 2432.415 1495.640 ;
        RECT 4.400 1492.240 2430.600 1493.640 ;
        RECT 0.270 1490.240 2432.415 1492.240 ;
        RECT 4.400 1488.840 2430.600 1490.240 ;
        RECT 0.270 1486.840 2432.415 1488.840 ;
        RECT 4.400 1485.440 2430.600 1486.840 ;
        RECT 0.270 1483.440 2432.415 1485.440 ;
        RECT 4.400 1482.040 2430.600 1483.440 ;
        RECT 0.270 1480.040 2432.415 1482.040 ;
        RECT 0.270 1478.640 2430.600 1480.040 ;
        RECT 0.270 1476.640 2432.415 1478.640 ;
        RECT 4.400 1475.240 2430.600 1476.640 ;
        RECT 0.270 1473.240 2432.415 1475.240 ;
        RECT 4.400 1471.840 2430.600 1473.240 ;
        RECT 0.270 1469.840 2432.415 1471.840 ;
        RECT 4.400 1468.440 2430.600 1469.840 ;
        RECT 0.270 1466.440 2432.415 1468.440 ;
        RECT 4.400 1465.040 2430.600 1466.440 ;
        RECT 0.270 1463.040 2432.415 1465.040 ;
        RECT 4.400 1461.640 2430.600 1463.040 ;
        RECT 0.270 1459.640 2432.415 1461.640 ;
        RECT 0.270 1458.240 2430.600 1459.640 ;
        RECT 0.270 1456.240 2432.415 1458.240 ;
        RECT 4.400 1454.840 2430.600 1456.240 ;
        RECT 0.270 1452.840 2432.415 1454.840 ;
        RECT 0.270 1451.440 2430.600 1452.840 ;
        RECT 0.270 1449.440 2432.415 1451.440 ;
        RECT 0.270 1448.040 2430.600 1449.440 ;
        RECT 0.270 1446.040 2432.415 1448.040 ;
        RECT 0.270 1444.640 2430.600 1446.040 ;
        RECT 0.270 1442.640 2432.415 1444.640 ;
        RECT 0.270 1441.240 2430.600 1442.640 ;
        RECT 0.270 1439.240 2432.415 1441.240 ;
        RECT 0.270 1437.840 2430.600 1439.240 ;
        RECT 0.270 1435.840 2432.415 1437.840 ;
        RECT 0.270 1434.440 2430.600 1435.840 ;
        RECT 0.270 1415.440 2432.415 1434.440 ;
        RECT 4.400 1414.040 2432.415 1415.440 ;
        RECT 0.270 1412.040 2432.415 1414.040 ;
        RECT 4.400 1410.640 2432.415 1412.040 ;
        RECT 0.270 1408.640 2432.415 1410.640 ;
        RECT 4.400 1407.240 2432.415 1408.640 ;
        RECT 0.270 1405.240 2432.415 1407.240 ;
        RECT 4.400 1403.840 2432.415 1405.240 ;
        RECT 0.270 1398.440 2432.415 1403.840 ;
        RECT 4.400 1397.040 2432.415 1398.440 ;
        RECT 0.270 1395.040 2432.415 1397.040 ;
        RECT 4.400 1393.640 2432.415 1395.040 ;
        RECT 0.270 1391.640 2432.415 1393.640 ;
        RECT 4.400 1390.240 2432.415 1391.640 ;
        RECT 0.270 1388.240 2432.415 1390.240 ;
        RECT 4.400 1386.840 2432.415 1388.240 ;
        RECT 0.270 1384.840 2432.415 1386.840 ;
        RECT 4.400 1383.440 2432.415 1384.840 ;
        RECT 0.270 1378.040 2432.415 1383.440 ;
        RECT 4.400 1376.640 2432.415 1378.040 ;
        RECT 0.270 1374.640 2432.415 1376.640 ;
        RECT 4.400 1373.240 2432.415 1374.640 ;
        RECT 0.270 1371.240 2432.415 1373.240 ;
        RECT 4.400 1369.840 2432.415 1371.240 ;
        RECT 0.270 1367.840 2432.415 1369.840 ;
        RECT 4.400 1366.440 2432.415 1367.840 ;
        RECT 0.270 1364.440 2432.415 1366.440 ;
        RECT 4.400 1363.040 2432.415 1364.440 ;
        RECT 0.270 1357.640 2432.415 1363.040 ;
        RECT 4.400 1356.240 2432.415 1357.640 ;
        RECT 0.270 1354.240 2432.415 1356.240 ;
        RECT 4.400 1352.840 2432.415 1354.240 ;
        RECT 0.270 1350.840 2432.415 1352.840 ;
        RECT 4.400 1349.440 2430.600 1350.840 ;
        RECT 0.270 1347.440 2432.415 1349.440 ;
        RECT 4.400 1346.040 2430.600 1347.440 ;
        RECT 0.270 1344.040 2432.415 1346.040 ;
        RECT 4.400 1342.640 2430.600 1344.040 ;
        RECT 0.270 1340.640 2432.415 1342.640 ;
        RECT 0.270 1339.240 2430.600 1340.640 ;
        RECT 0.270 1337.240 2432.415 1339.240 ;
        RECT 4.400 1335.840 2430.600 1337.240 ;
        RECT 0.270 1333.840 2432.415 1335.840 ;
        RECT 4.400 1332.440 2430.600 1333.840 ;
        RECT 0.270 1330.440 2432.415 1332.440 ;
        RECT 4.400 1329.040 2430.600 1330.440 ;
        RECT 0.270 1327.040 2432.415 1329.040 ;
        RECT 4.400 1325.640 2430.600 1327.040 ;
        RECT 0.270 1323.640 2432.415 1325.640 ;
        RECT 4.400 1322.240 2430.600 1323.640 ;
        RECT 0.270 1320.240 2432.415 1322.240 ;
        RECT 0.270 1318.840 2430.600 1320.240 ;
        RECT 0.270 1316.840 2432.415 1318.840 ;
        RECT 4.400 1315.440 2430.600 1316.840 ;
        RECT 0.270 1313.440 2432.415 1315.440 ;
        RECT 4.400 1312.040 2430.600 1313.440 ;
        RECT 0.270 1310.040 2432.415 1312.040 ;
        RECT 4.400 1308.640 2430.600 1310.040 ;
        RECT 0.270 1306.640 2432.415 1308.640 ;
        RECT 4.400 1305.240 2430.600 1306.640 ;
        RECT 0.270 1303.240 2432.415 1305.240 ;
        RECT 4.400 1301.840 2430.600 1303.240 ;
        RECT 0.270 1299.840 2432.415 1301.840 ;
        RECT 0.270 1298.440 2430.600 1299.840 ;
        RECT 0.270 1296.440 2432.415 1298.440 ;
        RECT 4.400 1295.040 2430.600 1296.440 ;
        RECT 0.270 1293.040 2432.415 1295.040 ;
        RECT 4.400 1291.640 2430.600 1293.040 ;
        RECT 0.270 1289.640 2432.415 1291.640 ;
        RECT 4.400 1288.240 2430.600 1289.640 ;
        RECT 0.270 1286.240 2432.415 1288.240 ;
        RECT 4.400 1284.840 2430.600 1286.240 ;
        RECT 0.270 1282.840 2432.415 1284.840 ;
        RECT 4.400 1281.440 2430.600 1282.840 ;
        RECT 0.270 1279.440 2432.415 1281.440 ;
        RECT 0.270 1278.040 2430.600 1279.440 ;
        RECT 0.270 1276.040 2432.415 1278.040 ;
        RECT 4.400 1274.640 2430.600 1276.040 ;
        RECT 0.270 1272.640 2432.415 1274.640 ;
        RECT 4.400 1271.240 2430.600 1272.640 ;
        RECT 0.270 1269.240 2432.415 1271.240 ;
        RECT 4.400 1267.840 2430.600 1269.240 ;
        RECT 0.270 1265.840 2432.415 1267.840 ;
        RECT 4.400 1264.440 2430.600 1265.840 ;
        RECT 0.270 1262.440 2432.415 1264.440 ;
        RECT 4.400 1261.040 2430.600 1262.440 ;
        RECT 0.270 1259.040 2432.415 1261.040 ;
        RECT 0.270 1257.640 2430.600 1259.040 ;
        RECT 0.270 1255.640 2432.415 1257.640 ;
        RECT 4.400 1254.240 2430.600 1255.640 ;
        RECT 0.270 1252.240 2432.415 1254.240 ;
        RECT 4.400 1250.840 2430.600 1252.240 ;
        RECT 0.270 1248.840 2432.415 1250.840 ;
        RECT 4.400 1247.440 2430.600 1248.840 ;
        RECT 0.270 1245.440 2432.415 1247.440 ;
        RECT 4.400 1244.040 2430.600 1245.440 ;
        RECT 0.270 1242.040 2432.415 1244.040 ;
        RECT 4.400 1240.640 2430.600 1242.040 ;
        RECT 0.270 1238.640 2432.415 1240.640 ;
        RECT 0.270 1237.240 2430.600 1238.640 ;
        RECT 0.270 1235.240 2432.415 1237.240 ;
        RECT 4.400 1233.840 2430.600 1235.240 ;
        RECT 0.270 1231.840 2432.415 1233.840 ;
        RECT 4.400 1230.440 2430.600 1231.840 ;
        RECT 0.270 1228.440 2432.415 1230.440 ;
        RECT 0.270 1227.040 2430.600 1228.440 ;
        RECT 0.270 1225.040 2432.415 1227.040 ;
        RECT 0.270 1223.640 2430.600 1225.040 ;
        RECT 0.270 1221.640 2432.415 1223.640 ;
        RECT 0.270 1220.240 2430.600 1221.640 ;
        RECT 0.270 1218.240 2432.415 1220.240 ;
        RECT 0.270 1216.840 2430.600 1218.240 ;
        RECT 0.270 1214.840 2432.415 1216.840 ;
        RECT 0.270 1213.440 2430.600 1214.840 ;
        RECT 0.270 1211.440 2432.415 1213.440 ;
        RECT 0.270 1210.040 2430.600 1211.440 ;
        RECT 0.270 1208.040 2432.415 1210.040 ;
        RECT 0.270 1206.640 2430.600 1208.040 ;
        RECT 0.270 1204.640 2432.415 1206.640 ;
        RECT 0.270 1203.240 2430.600 1204.640 ;
        RECT 0.270 1201.240 2432.415 1203.240 ;
        RECT 0.270 1199.840 2430.600 1201.240 ;
        RECT 0.270 1197.840 2432.415 1199.840 ;
        RECT 0.270 1196.440 2430.600 1197.840 ;
        RECT 0.270 1194.440 2432.415 1196.440 ;
        RECT 0.270 1193.040 2430.600 1194.440 ;
        RECT 0.270 1191.040 2432.415 1193.040 ;
        RECT 4.400 1189.640 2430.600 1191.040 ;
        RECT 0.270 1187.640 2432.415 1189.640 ;
        RECT 4.400 1186.240 2430.600 1187.640 ;
        RECT 0.270 1184.240 2432.415 1186.240 ;
        RECT 4.400 1182.840 2430.600 1184.240 ;
        RECT 0.270 1180.840 2432.415 1182.840 ;
        RECT 0.270 1179.440 2430.600 1180.840 ;
        RECT 0.270 1177.440 2432.415 1179.440 ;
        RECT 4.400 1176.040 2430.600 1177.440 ;
        RECT 0.270 1174.040 2432.415 1176.040 ;
        RECT 4.400 1172.640 2430.600 1174.040 ;
        RECT 0.270 1170.640 2432.415 1172.640 ;
        RECT 4.400 1169.240 2430.600 1170.640 ;
        RECT 0.270 1167.240 2432.415 1169.240 ;
        RECT 4.400 1165.840 2430.600 1167.240 ;
        RECT 0.270 1163.840 2432.415 1165.840 ;
        RECT 4.400 1162.440 2430.600 1163.840 ;
        RECT 0.270 1160.440 2432.415 1162.440 ;
        RECT 0.270 1159.040 2430.600 1160.440 ;
        RECT 0.270 1157.040 2432.415 1159.040 ;
        RECT 4.400 1155.640 2430.600 1157.040 ;
        RECT 0.270 1153.640 2432.415 1155.640 ;
        RECT 4.400 1152.240 2430.600 1153.640 ;
        RECT 0.270 1150.240 2432.415 1152.240 ;
        RECT 4.400 1148.840 2430.600 1150.240 ;
        RECT 0.270 1146.840 2432.415 1148.840 ;
        RECT 4.400 1145.440 2430.600 1146.840 ;
        RECT 0.270 1143.440 2432.415 1145.440 ;
        RECT 4.400 1142.040 2430.600 1143.440 ;
        RECT 0.270 1140.040 2432.415 1142.040 ;
        RECT 0.270 1138.640 2430.600 1140.040 ;
        RECT 0.270 1136.640 2432.415 1138.640 ;
        RECT 4.400 1135.240 2430.600 1136.640 ;
        RECT 0.270 1133.240 2432.415 1135.240 ;
        RECT 4.400 1131.840 2430.600 1133.240 ;
        RECT 0.270 1129.840 2432.415 1131.840 ;
        RECT 4.400 1128.440 2430.600 1129.840 ;
        RECT 0.270 1126.440 2432.415 1128.440 ;
        RECT 4.400 1125.040 2430.600 1126.440 ;
        RECT 0.270 1123.040 2432.415 1125.040 ;
        RECT 4.400 1121.640 2430.600 1123.040 ;
        RECT 0.270 1119.640 2432.415 1121.640 ;
        RECT 0.270 1118.240 2430.600 1119.640 ;
        RECT 0.270 1116.240 2432.415 1118.240 ;
        RECT 4.400 1114.840 2430.600 1116.240 ;
        RECT 0.270 1112.840 2432.415 1114.840 ;
        RECT 4.400 1111.440 2430.600 1112.840 ;
        RECT 0.270 1109.440 2432.415 1111.440 ;
        RECT 4.400 1108.040 2430.600 1109.440 ;
        RECT 0.270 1106.040 2432.415 1108.040 ;
        RECT 4.400 1104.640 2430.600 1106.040 ;
        RECT 0.270 1102.640 2432.415 1104.640 ;
        RECT 4.400 1101.240 2430.600 1102.640 ;
        RECT 0.270 1099.240 2432.415 1101.240 ;
        RECT 0.270 1097.840 2430.600 1099.240 ;
        RECT 0.270 1095.840 2432.415 1097.840 ;
        RECT 4.400 1094.440 2430.600 1095.840 ;
        RECT 0.270 1092.440 2432.415 1094.440 ;
        RECT 4.400 1091.040 2430.600 1092.440 ;
        RECT 0.270 1089.040 2432.415 1091.040 ;
        RECT 4.400 1087.640 2430.600 1089.040 ;
        RECT 0.270 1085.640 2432.415 1087.640 ;
        RECT 4.400 1084.240 2430.600 1085.640 ;
        RECT 0.270 1082.240 2432.415 1084.240 ;
        RECT 4.400 1080.840 2430.600 1082.240 ;
        RECT 0.270 1078.840 2432.415 1080.840 ;
        RECT 0.270 1077.440 2430.600 1078.840 ;
        RECT 0.270 1075.440 2432.415 1077.440 ;
        RECT 4.400 1074.040 2430.600 1075.440 ;
        RECT 0.270 1072.040 2432.415 1074.040 ;
        RECT 4.400 1070.640 2430.600 1072.040 ;
        RECT 0.270 1068.640 2432.415 1070.640 ;
        RECT 4.400 1067.240 2430.600 1068.640 ;
        RECT 0.270 1065.240 2432.415 1067.240 ;
        RECT 0.270 1063.840 2430.600 1065.240 ;
        RECT 0.270 1061.840 2432.415 1063.840 ;
        RECT 4.400 1060.440 2430.600 1061.840 ;
        RECT 0.270 1058.440 2432.415 1060.440 ;
        RECT 4.400 1057.040 2430.600 1058.440 ;
        RECT 0.270 1055.040 2432.415 1057.040 ;
        RECT 4.400 1053.640 2430.600 1055.040 ;
        RECT 0.270 1051.640 2432.415 1053.640 ;
        RECT 4.400 1050.240 2430.600 1051.640 ;
        RECT 0.270 1048.240 2432.415 1050.240 ;
        RECT 4.400 1046.840 2430.600 1048.240 ;
        RECT 0.270 1044.840 2432.415 1046.840 ;
        RECT 4.400 1043.440 2430.600 1044.840 ;
        RECT 0.270 1041.440 2432.415 1043.440 ;
        RECT 4.400 1040.040 2430.600 1041.440 ;
        RECT 0.270 1038.040 2432.415 1040.040 ;
        RECT 0.270 1036.640 2430.600 1038.040 ;
        RECT 0.270 1034.640 2432.415 1036.640 ;
        RECT 4.400 1033.240 2430.600 1034.640 ;
        RECT 0.270 1031.240 2432.415 1033.240 ;
        RECT 4.400 1029.840 2430.600 1031.240 ;
        RECT 0.270 1027.840 2432.415 1029.840 ;
        RECT 4.400 1026.440 2430.600 1027.840 ;
        RECT 0.270 1024.440 2432.415 1026.440 ;
        RECT 4.400 1023.040 2430.600 1024.440 ;
        RECT 0.270 1021.040 2432.415 1023.040 ;
        RECT 4.400 1019.640 2430.600 1021.040 ;
        RECT 0.270 1017.640 2432.415 1019.640 ;
        RECT 0.270 1016.240 2430.600 1017.640 ;
        RECT 0.270 1014.240 2432.415 1016.240 ;
        RECT 4.400 1012.840 2430.600 1014.240 ;
        RECT 0.270 1010.840 2432.415 1012.840 ;
        RECT 4.400 1009.440 2430.600 1010.840 ;
        RECT 0.270 1007.440 2432.415 1009.440 ;
        RECT 4.400 1006.040 2430.600 1007.440 ;
        RECT 0.270 1004.040 2432.415 1006.040 ;
        RECT 0.270 1002.640 2430.600 1004.040 ;
        RECT 0.270 1000.640 2432.415 1002.640 ;
        RECT 0.270 999.240 2430.600 1000.640 ;
        RECT 0.270 997.240 2432.415 999.240 ;
        RECT 0.270 995.840 2430.600 997.240 ;
        RECT 0.270 993.840 2432.415 995.840 ;
        RECT 0.270 992.440 2430.600 993.840 ;
        RECT 0.270 990.440 2432.415 992.440 ;
        RECT 0.270 989.040 2430.600 990.440 ;
        RECT 0.270 987.040 2432.415 989.040 ;
        RECT 0.270 985.640 2430.600 987.040 ;
        RECT 0.270 983.640 2432.415 985.640 ;
        RECT 0.270 982.240 2430.600 983.640 ;
        RECT 0.270 966.640 2432.415 982.240 ;
        RECT 4.400 965.240 2432.415 966.640 ;
        RECT 0.270 963.240 2432.415 965.240 ;
        RECT 4.400 961.840 2430.600 963.240 ;
        RECT 0.270 959.840 2432.415 961.840 ;
        RECT 0.270 958.440 2430.600 959.840 ;
        RECT 0.270 956.440 2432.415 958.440 ;
        RECT 4.400 955.040 2430.600 956.440 ;
        RECT 0.270 953.040 2432.415 955.040 ;
        RECT 4.400 951.640 2430.600 953.040 ;
        RECT 0.270 949.640 2432.415 951.640 ;
        RECT 4.400 948.240 2430.600 949.640 ;
        RECT 0.270 946.240 2432.415 948.240 ;
        RECT 4.400 944.840 2430.600 946.240 ;
        RECT 0.270 942.840 2432.415 944.840 ;
        RECT 4.400 941.440 2430.600 942.840 ;
        RECT 0.270 939.440 2432.415 941.440 ;
        RECT 0.270 938.040 2430.600 939.440 ;
        RECT 0.270 936.040 2432.415 938.040 ;
        RECT 4.400 934.640 2430.600 936.040 ;
        RECT 0.270 932.640 2432.415 934.640 ;
        RECT 4.400 931.240 2430.600 932.640 ;
        RECT 0.270 929.240 2432.415 931.240 ;
        RECT 4.400 927.840 2430.600 929.240 ;
        RECT 0.270 925.840 2432.415 927.840 ;
        RECT 4.400 924.440 2430.600 925.840 ;
        RECT 0.270 922.440 2432.415 924.440 ;
        RECT 4.400 921.040 2430.600 922.440 ;
        RECT 0.270 919.040 2432.415 921.040 ;
        RECT 0.270 917.640 2430.600 919.040 ;
        RECT 0.270 915.640 2432.415 917.640 ;
        RECT 4.400 914.240 2430.600 915.640 ;
        RECT 0.270 912.240 2432.415 914.240 ;
        RECT 4.400 910.840 2430.600 912.240 ;
        RECT 0.270 908.840 2432.415 910.840 ;
        RECT 4.400 907.440 2430.600 908.840 ;
        RECT 0.270 905.440 2432.415 907.440 ;
        RECT 4.400 904.040 2430.600 905.440 ;
        RECT 0.270 902.040 2432.415 904.040 ;
        RECT 4.400 900.640 2430.600 902.040 ;
        RECT 0.270 898.640 2432.415 900.640 ;
        RECT 0.270 897.240 2430.600 898.640 ;
        RECT 0.270 895.240 2432.415 897.240 ;
        RECT 4.400 893.840 2430.600 895.240 ;
        RECT 0.270 891.840 2432.415 893.840 ;
        RECT 4.400 890.440 2430.600 891.840 ;
        RECT 0.270 888.440 2432.415 890.440 ;
        RECT 4.400 887.040 2430.600 888.440 ;
        RECT 0.270 885.040 2432.415 887.040 ;
        RECT 4.400 883.640 2430.600 885.040 ;
        RECT 0.270 881.640 2432.415 883.640 ;
        RECT 4.400 880.240 2430.600 881.640 ;
        RECT 0.270 878.240 2432.415 880.240 ;
        RECT 0.270 876.840 2430.600 878.240 ;
        RECT 0.270 874.840 2432.415 876.840 ;
        RECT 4.400 873.440 2430.600 874.840 ;
        RECT 0.270 871.440 2432.415 873.440 ;
        RECT 4.400 870.040 2430.600 871.440 ;
        RECT 0.270 868.040 2432.415 870.040 ;
        RECT 4.400 866.640 2430.600 868.040 ;
        RECT 0.270 864.640 2432.415 866.640 ;
        RECT 4.400 863.240 2430.600 864.640 ;
        RECT 0.270 861.240 2432.415 863.240 ;
        RECT 4.400 859.840 2430.600 861.240 ;
        RECT 0.270 857.840 2432.415 859.840 ;
        RECT 0.270 856.440 2430.600 857.840 ;
        RECT 0.270 854.440 2432.415 856.440 ;
        RECT 4.400 853.040 2430.600 854.440 ;
        RECT 0.270 851.040 2432.415 853.040 ;
        RECT 4.400 849.640 2430.600 851.040 ;
        RECT 0.270 847.640 2432.415 849.640 ;
        RECT 4.400 846.240 2430.600 847.640 ;
        RECT 0.270 844.240 2432.415 846.240 ;
        RECT 4.400 842.840 2430.600 844.240 ;
        RECT 0.270 840.840 2432.415 842.840 ;
        RECT 4.400 839.440 2430.600 840.840 ;
        RECT 0.270 837.440 2432.415 839.440 ;
        RECT 0.270 836.040 2430.600 837.440 ;
        RECT 0.270 834.040 2432.415 836.040 ;
        RECT 4.400 832.640 2430.600 834.040 ;
        RECT 0.270 830.640 2432.415 832.640 ;
        RECT 4.400 829.240 2430.600 830.640 ;
        RECT 0.270 827.240 2432.415 829.240 ;
        RECT 4.400 825.840 2430.600 827.240 ;
        RECT 0.270 823.840 2432.415 825.840 ;
        RECT 4.400 822.440 2430.600 823.840 ;
        RECT 0.270 820.440 2432.415 822.440 ;
        RECT 4.400 819.040 2430.600 820.440 ;
        RECT 0.270 817.040 2432.415 819.040 ;
        RECT 0.270 815.640 2430.600 817.040 ;
        RECT 0.270 813.640 2432.415 815.640 ;
        RECT 4.400 812.240 2430.600 813.640 ;
        RECT 0.270 810.240 2432.415 812.240 ;
        RECT 4.400 808.840 2430.600 810.240 ;
        RECT 0.270 806.840 2432.415 808.840 ;
        RECT 4.400 805.440 2430.600 806.840 ;
        RECT 0.270 803.440 2432.415 805.440 ;
        RECT 4.400 802.040 2430.600 803.440 ;
        RECT 0.270 800.040 2432.415 802.040 ;
        RECT 4.400 798.640 2430.600 800.040 ;
        RECT 0.270 796.640 2432.415 798.640 ;
        RECT 0.270 795.240 2430.600 796.640 ;
        RECT 0.270 793.240 2432.415 795.240 ;
        RECT 4.400 791.840 2430.600 793.240 ;
        RECT 0.270 789.840 2432.415 791.840 ;
        RECT 4.400 788.440 2430.600 789.840 ;
        RECT 0.270 786.440 2432.415 788.440 ;
        RECT 4.400 785.040 2430.600 786.440 ;
        RECT 0.270 783.040 2432.415 785.040 ;
        RECT 4.400 781.640 2430.600 783.040 ;
        RECT 0.270 779.640 2432.415 781.640 ;
        RECT 0.270 778.240 2430.600 779.640 ;
        RECT 0.270 776.240 2432.415 778.240 ;
        RECT 0.270 774.840 2430.600 776.240 ;
        RECT 0.270 772.840 2432.415 774.840 ;
        RECT 0.270 771.440 2430.600 772.840 ;
        RECT 0.270 769.440 2432.415 771.440 ;
        RECT 0.270 768.040 2430.600 769.440 ;
        RECT 0.270 766.040 2432.415 768.040 ;
        RECT 0.270 764.640 2430.600 766.040 ;
        RECT 0.270 762.640 2432.415 764.640 ;
        RECT 0.270 761.240 2430.600 762.640 ;
        RECT 0.270 759.240 2432.415 761.240 ;
        RECT 0.270 757.840 2430.600 759.240 ;
        RECT 0.270 755.840 2432.415 757.840 ;
        RECT 0.270 754.440 2430.600 755.840 ;
        RECT 0.270 752.440 2432.415 754.440 ;
        RECT 0.270 751.040 2430.600 752.440 ;
        RECT 0.270 749.040 2432.415 751.040 ;
        RECT 0.270 747.640 2430.600 749.040 ;
        RECT 0.270 745.640 2432.415 747.640 ;
        RECT 0.270 744.240 2430.600 745.640 ;
        RECT 0.270 742.240 2432.415 744.240 ;
        RECT 4.400 740.840 2430.600 742.240 ;
        RECT 0.270 738.840 2432.415 740.840 ;
        RECT 4.400 737.440 2430.600 738.840 ;
        RECT 0.270 735.440 2432.415 737.440 ;
        RECT 0.270 734.040 2430.600 735.440 ;
        RECT 0.270 732.040 2432.415 734.040 ;
        RECT 4.400 730.640 2430.600 732.040 ;
        RECT 0.270 728.640 2432.415 730.640 ;
        RECT 4.400 727.240 2430.600 728.640 ;
        RECT 0.270 725.240 2432.415 727.240 ;
        RECT 4.400 723.840 2430.600 725.240 ;
        RECT 0.270 721.840 2432.415 723.840 ;
        RECT 4.400 720.440 2430.600 721.840 ;
        RECT 0.270 718.440 2432.415 720.440 ;
        RECT 4.400 717.040 2430.600 718.440 ;
        RECT 0.270 715.040 2432.415 717.040 ;
        RECT 0.270 713.640 2430.600 715.040 ;
        RECT 0.270 711.640 2432.415 713.640 ;
        RECT 4.400 710.240 2430.600 711.640 ;
        RECT 0.270 708.240 2432.415 710.240 ;
        RECT 4.400 706.840 2430.600 708.240 ;
        RECT 0.270 704.840 2432.415 706.840 ;
        RECT 4.400 703.440 2430.600 704.840 ;
        RECT 0.270 701.440 2432.415 703.440 ;
        RECT 4.400 700.040 2430.600 701.440 ;
        RECT 0.270 698.040 2432.415 700.040 ;
        RECT 4.400 696.640 2430.600 698.040 ;
        RECT 0.270 694.640 2432.415 696.640 ;
        RECT 0.270 693.240 2430.600 694.640 ;
        RECT 0.270 691.240 2432.415 693.240 ;
        RECT 4.400 689.840 2430.600 691.240 ;
        RECT 0.270 687.840 2432.415 689.840 ;
        RECT 4.400 686.440 2430.600 687.840 ;
        RECT 0.270 684.440 2432.415 686.440 ;
        RECT 4.400 683.040 2430.600 684.440 ;
        RECT 0.270 681.040 2432.415 683.040 ;
        RECT 4.400 679.640 2430.600 681.040 ;
        RECT 0.270 677.640 2432.415 679.640 ;
        RECT 4.400 676.240 2430.600 677.640 ;
        RECT 0.270 674.240 2432.415 676.240 ;
        RECT 0.270 672.840 2430.600 674.240 ;
        RECT 0.270 670.840 2432.415 672.840 ;
        RECT 4.400 669.440 2430.600 670.840 ;
        RECT 0.270 667.440 2432.415 669.440 ;
        RECT 4.400 666.040 2430.600 667.440 ;
        RECT 0.270 664.040 2432.415 666.040 ;
        RECT 4.400 662.640 2430.600 664.040 ;
        RECT 0.270 660.640 2432.415 662.640 ;
        RECT 4.400 659.240 2430.600 660.640 ;
        RECT 0.270 657.240 2432.415 659.240 ;
        RECT 4.400 655.840 2430.600 657.240 ;
        RECT 0.270 653.840 2432.415 655.840 ;
        RECT 0.270 652.440 2430.600 653.840 ;
        RECT 0.270 650.440 2432.415 652.440 ;
        RECT 4.400 649.040 2430.600 650.440 ;
        RECT 0.270 647.040 2432.415 649.040 ;
        RECT 4.400 645.640 2430.600 647.040 ;
        RECT 0.270 643.640 2432.415 645.640 ;
        RECT 4.400 642.240 2430.600 643.640 ;
        RECT 0.270 640.240 2432.415 642.240 ;
        RECT 4.400 638.840 2430.600 640.240 ;
        RECT 0.270 636.840 2432.415 638.840 ;
        RECT 4.400 635.440 2430.600 636.840 ;
        RECT 0.270 633.440 2432.415 635.440 ;
        RECT 0.270 632.040 2430.600 633.440 ;
        RECT 0.270 630.040 2432.415 632.040 ;
        RECT 4.400 628.640 2430.600 630.040 ;
        RECT 0.270 626.640 2432.415 628.640 ;
        RECT 4.400 625.240 2430.600 626.640 ;
        RECT 0.270 623.240 2432.415 625.240 ;
        RECT 4.400 621.840 2430.600 623.240 ;
        RECT 0.270 619.840 2432.415 621.840 ;
        RECT 4.400 618.440 2430.600 619.840 ;
        RECT 0.270 616.440 2432.415 618.440 ;
        RECT 4.400 615.040 2430.600 616.440 ;
        RECT 0.270 613.040 2432.415 615.040 ;
        RECT 0.270 611.640 2430.600 613.040 ;
        RECT 0.270 609.640 2432.415 611.640 ;
        RECT 4.400 608.240 2430.600 609.640 ;
        RECT 0.270 606.240 2432.415 608.240 ;
        RECT 4.400 604.840 2430.600 606.240 ;
        RECT 0.270 602.840 2432.415 604.840 ;
        RECT 4.400 601.440 2430.600 602.840 ;
        RECT 0.270 599.440 2432.415 601.440 ;
        RECT 4.400 598.040 2430.600 599.440 ;
        RECT 0.270 596.040 2432.415 598.040 ;
        RECT 4.400 594.640 2430.600 596.040 ;
        RECT 0.270 589.240 2432.415 594.640 ;
        RECT 4.400 587.840 2432.415 589.240 ;
        RECT 0.270 585.840 2432.415 587.840 ;
        RECT 4.400 584.440 2432.415 585.840 ;
        RECT 0.270 582.440 2432.415 584.440 ;
        RECT 4.400 581.040 2432.415 582.440 ;
        RECT 0.270 579.040 2432.415 581.040 ;
        RECT 4.400 577.640 2432.415 579.040 ;
        RECT 0.270 575.640 2432.415 577.640 ;
        RECT 4.400 574.240 2432.415 575.640 ;
        RECT 0.270 568.840 2432.415 574.240 ;
        RECT 4.400 567.440 2432.415 568.840 ;
        RECT 0.270 565.440 2432.415 567.440 ;
        RECT 4.400 564.040 2432.415 565.440 ;
        RECT 0.270 562.040 2432.415 564.040 ;
        RECT 4.400 560.640 2432.415 562.040 ;
        RECT 0.270 558.640 2432.415 560.640 ;
        RECT 4.400 557.240 2432.415 558.640 ;
        RECT 0.270 517.840 2432.415 557.240 ;
        RECT 4.400 516.440 2432.415 517.840 ;
        RECT 0.270 511.040 2432.415 516.440 ;
        RECT 4.400 509.640 2432.415 511.040 ;
        RECT 0.270 507.640 2432.415 509.640 ;
        RECT 4.400 506.240 2432.415 507.640 ;
        RECT 0.270 504.240 2432.415 506.240 ;
        RECT 4.400 502.840 2432.415 504.240 ;
        RECT 0.270 500.840 2432.415 502.840 ;
        RECT 4.400 499.440 2432.415 500.840 ;
        RECT 0.270 497.440 2432.415 499.440 ;
        RECT 4.400 496.040 2432.415 497.440 ;
        RECT 0.270 490.640 2432.415 496.040 ;
        RECT 4.400 489.240 2432.415 490.640 ;
        RECT 0.270 487.240 2432.415 489.240 ;
        RECT 4.400 485.840 2432.415 487.240 ;
        RECT 0.270 483.840 2432.415 485.840 ;
        RECT 4.400 482.440 2432.415 483.840 ;
        RECT 0.270 480.440 2432.415 482.440 ;
        RECT 4.400 479.040 2432.415 480.440 ;
        RECT 0.270 477.040 2432.415 479.040 ;
        RECT 4.400 475.640 2432.415 477.040 ;
        RECT 0.270 470.240 2432.415 475.640 ;
        RECT 4.400 468.840 2432.415 470.240 ;
        RECT 0.270 466.840 2432.415 468.840 ;
        RECT 4.400 465.440 2432.415 466.840 ;
        RECT 0.270 463.440 2432.415 465.440 ;
        RECT 4.400 462.040 2432.415 463.440 ;
        RECT 0.270 460.040 2432.415 462.040 ;
        RECT 4.400 458.640 2432.415 460.040 ;
        RECT 0.270 453.240 2432.415 458.640 ;
        RECT 0.270 451.840 2430.600 453.240 ;
        RECT 0.270 449.840 2432.415 451.840 ;
        RECT 0.270 448.440 2430.600 449.840 ;
        RECT 0.270 446.440 2432.415 448.440 ;
        RECT 0.270 445.040 2430.600 446.440 ;
        RECT 0.270 443.040 2432.415 445.040 ;
        RECT 0.270 441.640 2430.600 443.040 ;
        RECT 0.270 439.640 2432.415 441.640 ;
        RECT 0.270 438.240 2430.600 439.640 ;
        RECT 0.270 436.240 2432.415 438.240 ;
        RECT 0.270 434.840 2430.600 436.240 ;
        RECT 0.270 432.840 2432.415 434.840 ;
        RECT 0.270 431.440 2430.600 432.840 ;
        RECT 0.270 429.440 2432.415 431.440 ;
        RECT 0.270 428.040 2430.600 429.440 ;
        RECT 0.270 426.040 2432.415 428.040 ;
        RECT 0.270 424.640 2430.600 426.040 ;
        RECT 0.270 422.640 2432.415 424.640 ;
        RECT 0.270 421.240 2430.600 422.640 ;
        RECT 0.270 419.240 2432.415 421.240 ;
        RECT 0.270 417.840 2430.600 419.240 ;
        RECT 0.270 415.840 2432.415 417.840 ;
        RECT 0.270 414.440 2430.600 415.840 ;
        RECT 0.270 412.440 2432.415 414.440 ;
        RECT 0.270 411.040 2430.600 412.440 ;
        RECT 0.270 409.040 2432.415 411.040 ;
        RECT 0.270 407.640 2430.600 409.040 ;
        RECT 0.270 405.640 2432.415 407.640 ;
        RECT 0.270 404.240 2430.600 405.640 ;
        RECT 0.270 402.240 2432.415 404.240 ;
        RECT 0.270 400.840 2430.600 402.240 ;
        RECT 0.270 398.840 2432.415 400.840 ;
        RECT 0.270 397.440 2430.600 398.840 ;
        RECT 0.270 395.440 2432.415 397.440 ;
        RECT 0.270 394.040 2430.600 395.440 ;
        RECT 0.270 392.040 2432.415 394.040 ;
        RECT 0.270 390.640 2430.600 392.040 ;
        RECT 0.270 388.640 2432.415 390.640 ;
        RECT 0.270 387.240 2430.600 388.640 ;
        RECT 0.270 385.240 2432.415 387.240 ;
        RECT 0.270 383.840 2430.600 385.240 ;
        RECT 0.270 381.840 2432.415 383.840 ;
        RECT 4.400 380.440 2430.600 381.840 ;
        RECT 0.270 378.440 2432.415 380.440 ;
        RECT 4.400 377.040 2430.600 378.440 ;
        RECT 0.270 375.040 2432.415 377.040 ;
        RECT 4.400 373.640 2430.600 375.040 ;
        RECT 0.270 371.640 2432.415 373.640 ;
        RECT 4.400 370.240 2430.600 371.640 ;
        RECT 0.270 368.240 2432.415 370.240 ;
        RECT 4.400 366.840 2430.600 368.240 ;
        RECT 0.270 364.840 2432.415 366.840 ;
        RECT 4.400 363.440 2430.600 364.840 ;
        RECT 0.270 361.440 2432.415 363.440 ;
        RECT 4.400 360.040 2430.600 361.440 ;
        RECT 0.270 358.040 2432.415 360.040 ;
        RECT 4.400 356.640 2430.600 358.040 ;
        RECT 0.270 354.640 2432.415 356.640 ;
        RECT 4.400 353.240 2430.600 354.640 ;
        RECT 0.270 351.240 2432.415 353.240 ;
        RECT 4.400 349.840 2430.600 351.240 ;
        RECT 0.270 347.840 2432.415 349.840 ;
        RECT 4.400 346.440 2430.600 347.840 ;
        RECT 0.270 344.440 2432.415 346.440 ;
        RECT 4.400 343.040 2430.600 344.440 ;
        RECT 0.270 341.040 2432.415 343.040 ;
        RECT 4.400 339.640 2430.600 341.040 ;
        RECT 0.270 337.640 2432.415 339.640 ;
        RECT 4.400 336.240 2430.600 337.640 ;
        RECT 0.270 334.240 2432.415 336.240 ;
        RECT 4.400 332.840 2430.600 334.240 ;
        RECT 0.270 330.840 2432.415 332.840 ;
        RECT 4.400 329.440 2430.600 330.840 ;
        RECT 0.270 327.440 2432.415 329.440 ;
        RECT 4.400 326.040 2430.600 327.440 ;
        RECT 0.270 324.040 2432.415 326.040 ;
        RECT 4.400 322.640 2430.600 324.040 ;
        RECT 0.270 320.640 2432.415 322.640 ;
        RECT 4.400 319.240 2430.600 320.640 ;
        RECT 0.270 317.240 2432.415 319.240 ;
        RECT 4.400 315.840 2430.600 317.240 ;
        RECT 0.270 313.840 2432.415 315.840 ;
        RECT 4.400 312.440 2430.600 313.840 ;
        RECT 0.270 310.440 2432.415 312.440 ;
        RECT 4.400 309.040 2430.600 310.440 ;
        RECT 0.270 307.040 2432.415 309.040 ;
        RECT 4.400 305.640 2430.600 307.040 ;
        RECT 0.270 303.640 2432.415 305.640 ;
        RECT 4.400 302.240 2430.600 303.640 ;
        RECT 0.270 300.240 2432.415 302.240 ;
        RECT 4.400 298.840 2430.600 300.240 ;
        RECT 0.270 296.840 2432.415 298.840 ;
        RECT 4.400 295.440 2430.600 296.840 ;
        RECT 0.270 293.440 2432.415 295.440 ;
        RECT 4.400 292.040 2430.600 293.440 ;
        RECT 0.270 290.040 2432.415 292.040 ;
        RECT 4.400 288.640 2430.600 290.040 ;
        RECT 0.270 286.640 2432.415 288.640 ;
        RECT 4.400 285.240 2430.600 286.640 ;
        RECT 0.270 283.240 2432.415 285.240 ;
        RECT 4.400 281.840 2430.600 283.240 ;
        RECT 0.270 279.840 2432.415 281.840 ;
        RECT 4.400 278.440 2430.600 279.840 ;
        RECT 0.270 276.440 2432.415 278.440 ;
        RECT 4.400 275.040 2430.600 276.440 ;
        RECT 0.270 273.040 2432.415 275.040 ;
        RECT 4.400 271.640 2430.600 273.040 ;
        RECT 0.270 269.640 2432.415 271.640 ;
        RECT 4.400 268.240 2430.600 269.640 ;
        RECT 0.270 266.240 2432.415 268.240 ;
        RECT 4.400 264.840 2430.600 266.240 ;
        RECT 0.270 262.840 2432.415 264.840 ;
        RECT 4.400 261.440 2430.600 262.840 ;
        RECT 0.270 259.440 2432.415 261.440 ;
        RECT 4.400 258.040 2430.600 259.440 ;
        RECT 0.270 256.040 2432.415 258.040 ;
        RECT 4.400 254.640 2430.600 256.040 ;
        RECT 0.270 252.640 2432.415 254.640 ;
        RECT 4.400 251.240 2430.600 252.640 ;
        RECT 0.270 249.240 2432.415 251.240 ;
        RECT 4.400 247.840 2430.600 249.240 ;
        RECT 0.270 245.840 2432.415 247.840 ;
        RECT 4.400 244.440 2430.600 245.840 ;
        RECT 0.270 242.440 2432.415 244.440 ;
        RECT 4.400 241.040 2430.600 242.440 ;
        RECT 0.270 239.040 2432.415 241.040 ;
        RECT 4.400 237.640 2430.600 239.040 ;
        RECT 0.270 235.640 2432.415 237.640 ;
        RECT 4.400 234.240 2430.600 235.640 ;
        RECT 0.270 232.240 2432.415 234.240 ;
        RECT 4.400 230.840 2430.600 232.240 ;
        RECT 0.270 228.840 2432.415 230.840 ;
        RECT 4.400 227.440 2430.600 228.840 ;
        RECT 0.270 225.440 2432.415 227.440 ;
        RECT 4.400 224.040 2430.600 225.440 ;
        RECT 0.270 222.040 2432.415 224.040 ;
        RECT 4.400 220.640 2430.600 222.040 ;
        RECT 0.270 218.640 2432.415 220.640 ;
        RECT 4.400 217.240 2430.600 218.640 ;
        RECT 0.270 215.240 2432.415 217.240 ;
        RECT 4.400 213.840 2430.600 215.240 ;
        RECT 0.270 211.840 2432.415 213.840 ;
        RECT 4.400 210.440 2430.600 211.840 ;
        RECT 0.270 208.440 2432.415 210.440 ;
        RECT 4.400 207.040 2430.600 208.440 ;
        RECT 0.270 205.040 2432.415 207.040 ;
        RECT 4.400 203.640 2430.600 205.040 ;
        RECT 0.270 201.640 2432.415 203.640 ;
        RECT 4.400 200.240 2430.600 201.640 ;
        RECT 0.270 198.240 2432.415 200.240 ;
        RECT 4.400 196.840 2430.600 198.240 ;
        RECT 0.270 194.840 2432.415 196.840 ;
        RECT 4.400 193.440 2430.600 194.840 ;
        RECT 0.270 191.440 2432.415 193.440 ;
        RECT 4.400 190.040 2430.600 191.440 ;
        RECT 0.270 188.040 2432.415 190.040 ;
        RECT 4.400 186.640 2430.600 188.040 ;
        RECT 0.270 184.640 2432.415 186.640 ;
        RECT 4.400 183.240 2430.600 184.640 ;
        RECT 0.270 181.240 2432.415 183.240 ;
        RECT 4.400 179.840 2430.600 181.240 ;
        RECT 0.270 177.840 2432.415 179.840 ;
        RECT 4.400 176.440 2430.600 177.840 ;
        RECT 0.270 174.440 2432.415 176.440 ;
        RECT 4.400 173.040 2430.600 174.440 ;
        RECT 0.270 171.040 2432.415 173.040 ;
        RECT 4.400 169.640 2430.600 171.040 ;
        RECT 0.270 167.640 2432.415 169.640 ;
        RECT 4.400 166.240 2430.600 167.640 ;
        RECT 0.270 164.240 2432.415 166.240 ;
        RECT 4.400 162.840 2430.600 164.240 ;
        RECT 0.270 160.840 2432.415 162.840 ;
        RECT 4.400 159.440 2430.600 160.840 ;
        RECT 0.270 157.440 2432.415 159.440 ;
        RECT 4.400 156.040 2430.600 157.440 ;
        RECT 0.270 154.040 2432.415 156.040 ;
        RECT 4.400 152.640 2430.600 154.040 ;
        RECT 0.270 150.640 2432.415 152.640 ;
        RECT 4.400 149.240 2430.600 150.640 ;
        RECT 0.270 147.240 2432.415 149.240 ;
        RECT 4.400 145.840 2430.600 147.240 ;
        RECT 0.270 143.840 2432.415 145.840 ;
        RECT 4.400 142.440 2430.600 143.840 ;
        RECT 0.270 140.440 2432.415 142.440 ;
        RECT 4.400 139.040 2430.600 140.440 ;
        RECT 0.270 137.040 2432.415 139.040 ;
        RECT 4.400 135.640 2430.600 137.040 ;
        RECT 0.270 133.640 2432.415 135.640 ;
        RECT 4.400 132.240 2430.600 133.640 ;
        RECT 0.270 130.240 2432.415 132.240 ;
        RECT 4.400 128.840 2430.600 130.240 ;
        RECT 0.270 126.840 2432.415 128.840 ;
        RECT 4.400 125.440 2430.600 126.840 ;
        RECT 0.270 123.440 2432.415 125.440 ;
        RECT 4.400 122.040 2430.600 123.440 ;
        RECT 0.270 120.040 2432.415 122.040 ;
        RECT 4.400 118.640 2430.600 120.040 ;
        RECT 0.270 116.640 2432.415 118.640 ;
        RECT 4.400 115.240 2430.600 116.640 ;
        RECT 0.270 113.240 2432.415 115.240 ;
        RECT 4.400 111.840 2430.600 113.240 ;
        RECT 0.270 109.840 2432.415 111.840 ;
        RECT 4.400 108.440 2430.600 109.840 ;
        RECT 0.270 106.440 2432.415 108.440 ;
        RECT 4.400 105.040 2430.600 106.440 ;
        RECT 0.270 103.040 2432.415 105.040 ;
        RECT 4.400 101.640 2430.600 103.040 ;
        RECT 0.270 99.640 2432.415 101.640 ;
        RECT 4.400 98.240 2430.600 99.640 ;
        RECT 0.270 96.240 2432.415 98.240 ;
        RECT 4.400 94.840 2430.600 96.240 ;
        RECT 0.270 92.840 2432.415 94.840 ;
        RECT 4.400 91.440 2430.600 92.840 ;
        RECT 0.270 89.440 2432.415 91.440 ;
        RECT 4.400 88.040 2430.600 89.440 ;
        RECT 0.270 86.040 2432.415 88.040 ;
        RECT 4.400 84.640 2430.600 86.040 ;
        RECT 0.270 82.640 2432.415 84.640 ;
        RECT 4.400 81.240 2432.415 82.640 ;
        RECT 0.270 79.240 2432.415 81.240 ;
        RECT 4.400 77.840 2432.415 79.240 ;
        RECT 0.270 75.840 2432.415 77.840 ;
        RECT 4.400 74.440 2432.415 75.840 ;
        RECT 0.270 72.440 2432.415 74.440 ;
        RECT 4.400 71.040 2432.415 72.440 ;
        RECT 0.270 69.040 2432.415 71.040 ;
        RECT 4.400 67.640 2432.415 69.040 ;
        RECT 0.270 65.640 2432.415 67.640 ;
        RECT 4.400 64.240 2432.415 65.640 ;
        RECT 0.270 62.240 2432.415 64.240 ;
        RECT 4.400 60.840 2432.415 62.240 ;
        RECT 0.270 58.840 2432.415 60.840 ;
        RECT 4.400 57.440 2432.415 58.840 ;
        RECT 0.270 55.440 2432.415 57.440 ;
        RECT 4.400 54.040 2432.415 55.440 ;
        RECT 0.270 52.040 2432.415 54.040 ;
        RECT 4.400 50.640 2432.415 52.040 ;
        RECT 0.270 48.640 2432.415 50.640 ;
        RECT 4.400 47.240 2432.415 48.640 ;
        RECT 0.270 45.240 2432.415 47.240 ;
        RECT 4.400 43.840 2432.415 45.240 ;
        RECT 0.270 41.840 2432.415 43.840 ;
        RECT 4.400 40.440 2432.415 41.840 ;
        RECT 0.270 38.440 2432.415 40.440 ;
        RECT 4.400 37.040 2432.415 38.440 ;
        RECT 0.270 35.040 2432.415 37.040 ;
        RECT 4.400 33.640 2432.415 35.040 ;
        RECT 0.270 31.640 2432.415 33.640 ;
        RECT 4.400 30.240 2432.415 31.640 ;
        RECT 0.270 28.240 2432.415 30.240 ;
        RECT 4.400 26.840 2432.415 28.240 ;
        RECT 0.270 24.840 2432.415 26.840 ;
        RECT 4.400 23.440 2432.415 24.840 ;
        RECT 0.270 21.440 2432.415 23.440 ;
        RECT 4.400 20.040 2432.415 21.440 ;
        RECT 0.270 18.040 2432.415 20.040 ;
        RECT 4.400 16.640 2432.415 18.040 ;
        RECT 0.270 14.640 2432.415 16.640 ;
        RECT 4.400 13.240 2432.415 14.640 ;
        RECT 0.270 11.240 2432.415 13.240 ;
        RECT 4.400 9.840 2432.415 11.240 ;
        RECT 0.270 7.840 2432.415 9.840 ;
        RECT 4.400 6.440 2432.415 7.840 ;
        RECT 0.270 4.440 2432.415 6.440 ;
        RECT 4.400 3.040 2432.415 4.440 ;
        RECT 0.270 1.040 2432.415 3.040 ;
        RECT 4.400 0.190 2432.415 1.040 ;
      LAYER met4 ;
        RECT 0.295 3742.900 2433.105 3779.265 ;
        RECT 0.295 29.600 59.320 3742.900 ;
        RECT 61.720 29.600 64.620 3742.900 ;
        RECT 67.020 29.600 89.320 3742.900 ;
        RECT 91.720 29.600 94.620 3742.900 ;
        RECT 97.020 29.600 115.570 3742.900 ;
        RECT 117.970 29.600 120.870 3742.900 ;
        RECT 123.270 29.600 145.570 3742.900 ;
        RECT 147.970 29.600 150.870 3742.900 ;
        RECT 153.270 29.600 175.570 3742.900 ;
        RECT 177.970 29.600 180.870 3742.900 ;
        RECT 183.270 29.600 205.570 3742.900 ;
        RECT 207.970 29.600 210.870 3742.900 ;
        RECT 213.270 29.600 235.570 3742.900 ;
        RECT 237.970 29.600 240.870 3742.900 ;
        RECT 243.270 29.600 265.570 3742.900 ;
        RECT 267.970 29.600 270.870 3742.900 ;
        RECT 273.270 29.600 295.570 3742.900 ;
        RECT 297.970 29.600 300.870 3742.900 ;
        RECT 303.270 29.600 320.570 3742.900 ;
        RECT 322.970 29.600 325.870 3742.900 ;
        RECT 328.270 29.600 350.570 3742.900 ;
        RECT 352.970 29.600 355.870 3742.900 ;
        RECT 358.270 29.600 380.570 3742.900 ;
        RECT 382.970 29.600 385.870 3742.900 ;
        RECT 388.270 29.600 410.570 3742.900 ;
        RECT 412.970 29.600 415.870 3742.900 ;
        RECT 418.270 29.600 440.570 3742.900 ;
        RECT 442.970 29.600 445.870 3742.900 ;
        RECT 448.270 29.600 470.570 3742.900 ;
        RECT 472.970 29.600 475.870 3742.900 ;
        RECT 478.270 29.600 500.570 3742.900 ;
        RECT 502.970 29.600 505.870 3742.900 ;
        RECT 508.270 29.600 525.570 3742.900 ;
        RECT 527.970 29.600 530.870 3742.900 ;
        RECT 533.270 29.600 555.570 3742.900 ;
        RECT 557.970 29.600 560.870 3742.900 ;
        RECT 563.270 29.600 585.570 3742.900 ;
        RECT 587.970 29.600 590.870 3742.900 ;
        RECT 593.270 29.600 615.570 3742.900 ;
        RECT 617.970 29.600 620.870 3742.900 ;
        RECT 623.270 29.600 645.570 3742.900 ;
        RECT 647.970 29.600 650.870 3742.900 ;
        RECT 653.270 29.600 675.570 3742.900 ;
        RECT 677.970 29.600 680.870 3742.900 ;
        RECT 683.270 29.600 705.570 3742.900 ;
        RECT 707.970 29.600 710.870 3742.900 ;
        RECT 713.270 29.600 735.570 3742.900 ;
        RECT 737.970 29.600 740.870 3742.900 ;
        RECT 743.270 29.600 770.570 3742.900 ;
        RECT 772.970 29.600 775.870 3742.900 ;
        RECT 778.270 29.600 800.570 3742.900 ;
        RECT 802.970 29.600 805.870 3742.900 ;
        RECT 808.270 29.600 830.570 3742.900 ;
        RECT 832.970 29.600 835.870 3742.900 ;
        RECT 838.270 29.600 860.570 3742.900 ;
        RECT 862.970 29.600 865.870 3742.900 ;
        RECT 868.270 29.600 890.570 3742.900 ;
        RECT 892.970 29.600 895.870 3742.900 ;
        RECT 898.270 29.600 920.570 3742.900 ;
        RECT 922.970 29.600 925.870 3742.900 ;
        RECT 928.270 29.600 950.570 3742.900 ;
        RECT 952.970 29.600 955.870 3742.900 ;
        RECT 958.270 29.600 975.570 3742.900 ;
        RECT 977.970 29.600 980.870 3742.900 ;
        RECT 983.270 29.600 1005.570 3742.900 ;
        RECT 1007.970 29.600 1010.870 3742.900 ;
        RECT 1013.270 29.600 1035.570 3742.900 ;
        RECT 1037.970 29.600 1040.870 3742.900 ;
        RECT 1043.270 29.600 1065.570 3742.900 ;
        RECT 1067.970 29.600 1070.870 3742.900 ;
        RECT 1073.270 29.600 1095.570 3742.900 ;
        RECT 1097.970 29.600 1100.870 3742.900 ;
        RECT 1103.270 29.600 1125.570 3742.900 ;
        RECT 1127.970 29.600 1130.870 3742.900 ;
        RECT 1133.270 29.600 1155.570 3742.900 ;
        RECT 1157.970 29.600 1160.870 3742.900 ;
        RECT 1163.270 29.600 1180.570 3742.900 ;
        RECT 1182.970 29.600 1185.870 3742.900 ;
        RECT 1188.270 29.600 1210.570 3742.900 ;
        RECT 1212.970 29.600 1215.870 3742.900 ;
        RECT 1218.270 29.600 1240.570 3742.900 ;
        RECT 1242.970 29.600 1245.870 3742.900 ;
        RECT 1248.270 29.600 1270.570 3742.900 ;
        RECT 1272.970 29.600 1275.870 3742.900 ;
        RECT 1278.270 29.600 1300.570 3742.900 ;
        RECT 1302.970 29.600 1305.870 3742.900 ;
        RECT 1308.270 29.600 1330.570 3742.900 ;
        RECT 1332.970 29.600 1335.870 3742.900 ;
        RECT 1338.270 29.600 1360.570 3742.900 ;
        RECT 1362.970 29.600 1365.870 3742.900 ;
        RECT 1368.270 29.600 1385.570 3742.900 ;
        RECT 1387.970 29.600 1390.870 3742.900 ;
        RECT 1393.270 29.600 1415.570 3742.900 ;
        RECT 1417.970 29.600 1420.870 3742.900 ;
        RECT 1423.270 29.600 1445.570 3742.900 ;
        RECT 1447.970 29.600 1450.870 3742.900 ;
        RECT 1453.270 29.600 1475.570 3742.900 ;
        RECT 1477.970 29.600 1480.870 3742.900 ;
        RECT 1483.270 29.600 1505.570 3742.900 ;
        RECT 1507.970 29.600 1510.870 3742.900 ;
        RECT 1513.270 29.600 1535.570 3742.900 ;
        RECT 1537.970 29.600 1540.870 3742.900 ;
        RECT 1543.270 29.600 1565.570 3742.900 ;
        RECT 1567.970 29.600 1570.870 3742.900 ;
        RECT 1573.270 29.600 1610.570 3742.900 ;
        RECT 1612.970 29.600 1615.870 3742.900 ;
        RECT 1618.270 29.600 1640.570 3742.900 ;
        RECT 1642.970 29.600 1645.870 3742.900 ;
        RECT 1648.270 29.600 1670.570 3742.900 ;
        RECT 1672.970 29.600 1675.870 3742.900 ;
        RECT 1678.270 29.600 1700.570 3742.900 ;
        RECT 1702.970 29.600 1705.870 3742.900 ;
        RECT 1708.270 29.600 1730.570 3742.900 ;
        RECT 1732.970 29.600 1735.870 3742.900 ;
        RECT 1738.270 29.600 1760.570 3742.900 ;
        RECT 1762.970 29.600 1765.870 3742.900 ;
        RECT 1768.270 29.600 1790.570 3742.900 ;
        RECT 1792.970 29.600 1795.870 3742.900 ;
        RECT 1798.270 29.600 1815.570 3742.900 ;
        RECT 1817.970 29.600 1820.870 3742.900 ;
        RECT 1823.270 29.600 1845.570 3742.900 ;
        RECT 1847.970 29.600 1850.870 3742.900 ;
        RECT 1853.270 29.600 1875.570 3742.900 ;
        RECT 1877.970 29.600 1880.870 3742.900 ;
        RECT 1883.270 29.600 1905.570 3742.900 ;
        RECT 1907.970 29.600 1910.870 3742.900 ;
        RECT 1913.270 29.600 1935.570 3742.900 ;
        RECT 1937.970 29.600 1940.870 3742.900 ;
        RECT 1943.270 29.600 1965.570 3742.900 ;
        RECT 1967.970 29.600 1970.870 3742.900 ;
        RECT 1973.270 29.600 1995.570 3742.900 ;
        RECT 1997.970 29.600 2000.870 3742.900 ;
        RECT 2003.270 29.600 2020.570 3742.900 ;
        RECT 2022.970 29.600 2025.870 3742.900 ;
        RECT 2028.270 29.600 2050.570 3742.900 ;
        RECT 2052.970 29.600 2055.870 3742.900 ;
        RECT 2058.270 29.600 2080.570 3742.900 ;
        RECT 2082.970 29.600 2085.870 3742.900 ;
        RECT 2088.270 29.600 2110.570 3742.900 ;
        RECT 2112.970 29.600 2115.870 3742.900 ;
        RECT 2118.270 29.600 2140.570 3742.900 ;
        RECT 2142.970 29.600 2145.870 3742.900 ;
        RECT 2148.270 29.600 2170.570 3742.900 ;
        RECT 2172.970 29.600 2175.870 3742.900 ;
        RECT 2178.270 29.600 2200.570 3742.900 ;
        RECT 2202.970 29.600 2205.870 3742.900 ;
        RECT 2208.270 29.600 2225.570 3742.900 ;
        RECT 2227.970 29.600 2230.870 3742.900 ;
        RECT 2233.270 29.600 2255.570 3742.900 ;
        RECT 2257.970 29.600 2260.870 3742.900 ;
        RECT 2263.270 29.600 2285.570 3742.900 ;
        RECT 2287.970 29.600 2290.870 3742.900 ;
        RECT 2293.270 29.600 2315.570 3742.900 ;
        RECT 2317.970 29.600 2320.870 3742.900 ;
        RECT 2323.270 29.600 2345.570 3742.900 ;
        RECT 2347.970 29.600 2350.870 3742.900 ;
        RECT 2353.270 29.600 2375.570 3742.900 ;
        RECT 2377.970 29.600 2433.105 3742.900 ;
        RECT 0.295 0.855 2433.105 29.600 ;
  END
END eFPGA
END LIBRARY

